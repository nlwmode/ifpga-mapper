module top( \G0_pad  , \G10_pad  , \G11_pad  , \G12_pad  , \G13_pad  , \G1_pad  , \G29_reg/NET0131  , \G2_pad  , \G30_reg/NET0131  , \G31_reg/NET0131  , \G32_reg/NET0131  , \G33_reg/NET0131  , \G34_reg/NET0131  , \G35_reg/NET0131  , \G36_reg/NET0131  , \G37_reg/NET0131  , \G38_reg/NET0131  , \G39_reg/NET0131  , \G3_pad  , \G40_reg/NET0131  , \G41_reg/NET0131  , \G42_reg/NET0131  , \G43_reg/NET0131  , \G44_reg/NET0131  , \G46_reg/NET0131  , \G4_pad  , \G5_pad  , \G6_pad  , \G7_pad  , \G8_pad  , \G9_pad  , \G532_pad  , \G537_pad  , \G539_pad  , \G542_pad  , \G546_pad  , \G547_pad  , \G548_pad  , \G549_pad  , \G550_pad  , \G551_pad  , \G552_pad  , \_al_n0  , \_al_n1  , \g1667/_3_  , \g1737/_0_  , \g1744/_0_  , \g1787/_0_  , \g1811/_0_  , \g1830/_0_  , \g1831/_0_  , \g1846/_0_  , \g1852/_0_  , \g1866/_0_  , \g19/_2_  , \g1931/_0_  , \g1945/_0_  , \g2014/_0_  , \g2015/_0_  , \g2643/_0_  , \g2859/_1_  , \g3397/_2_  , \g3546/_0_  , \g3606/_3_  );
  input \G0_pad  ;
  input \G10_pad  ;
  input \G11_pad  ;
  input \G12_pad  ;
  input \G13_pad  ;
  input \G1_pad  ;
  input \G29_reg/NET0131  ;
  input \G2_pad  ;
  input \G30_reg/NET0131  ;
  input \G31_reg/NET0131  ;
  input \G32_reg/NET0131  ;
  input \G33_reg/NET0131  ;
  input \G34_reg/NET0131  ;
  input \G35_reg/NET0131  ;
  input \G36_reg/NET0131  ;
  input \G37_reg/NET0131  ;
  input \G38_reg/NET0131  ;
  input \G39_reg/NET0131  ;
  input \G3_pad  ;
  input \G40_reg/NET0131  ;
  input \G41_reg/NET0131  ;
  input \G42_reg/NET0131  ;
  input \G43_reg/NET0131  ;
  input \G44_reg/NET0131  ;
  input \G46_reg/NET0131  ;
  input \G4_pad  ;
  input \G5_pad  ;
  input \G6_pad  ;
  input \G7_pad  ;
  input \G8_pad  ;
  input \G9_pad  ;
  output \G532_pad  ;
  output \G537_pad  ;
  output \G539_pad  ;
  output \G542_pad  ;
  output \G546_pad  ;
  output \G547_pad  ;
  output \G548_pad  ;
  output \G549_pad  ;
  output \G550_pad  ;
  output \G551_pad  ;
  output \G552_pad  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1667/_3_  ;
  output \g1737/_0_  ;
  output \g1744/_0_  ;
  output \g1787/_0_  ;
  output \g1811/_0_  ;
  output \g1830/_0_  ;
  output \g1831/_0_  ;
  output \g1846/_0_  ;
  output \g1852/_0_  ;
  output \g1866/_0_  ;
  output \g19/_2_  ;
  output \g1931/_0_  ;
  output \g1945/_0_  ;
  output \g2014/_0_  ;
  output \g2015/_0_  ;
  output \g2643/_0_  ;
  output \g2859/_1_  ;
  output \g3397/_2_  ;
  output \g3546/_0_  ;
  output \g3606/_3_  ;
  wire n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 ;
  assign n34 = \G11_pad  & \G9_pad  ;
  assign n35 = \G8_pad  & n34 ;
  assign n36 = \G10_pad  & \G7_pad  ;
  assign n37 = ~n35 & n36 ;
  assign n32 = ~\G7_pad  & \G8_pad  ;
  assign n33 = \G30_reg/NET0131  & n32 ;
  assign n38 = ~\G10_pad  & \G9_pad  ;
  assign n39 = \G7_pad  & n38 ;
  assign n40 = ~n33 & ~n39 ;
  assign n41 = ~n37 & n40 ;
  assign n42 = \G32_reg/NET0131  & ~n41 ;
  assign n43 = ~\G13_pad  & ~n42 ;
  assign n44 = ~\G5_pad  & \G6_pad  ;
  assign n45 = \G3_pad  & \G4_pad  ;
  assign n46 = n44 & n45 ;
  assign n47 = \G11_pad  & n46 ;
  assign n48 = \G7_pad  & ~\G8_pad  ;
  assign n49 = \G8_pad  & \G9_pad  ;
  assign n52 = ~n48 & ~n49 ;
  assign n50 = \G10_pad  & ~\G9_pad  ;
  assign n51 = ~\G10_pad  & ~\G7_pad  ;
  assign n53 = ~n50 & ~n51 ;
  assign n54 = n52 & n53 ;
  assign n55 = ~\G7_pad  & n38 ;
  assign n56 = \G8_pad  & n55 ;
  assign n57 = ~n54 & ~n56 ;
  assign n58 = n47 & ~n57 ;
  assign n59 = \G36_reg/NET0131  & ~\G6_pad  ;
  assign n60 = \G4_pad  & \G6_pad  ;
  assign n61 = \G5_pad  & n60 ;
  assign n62 = \G11_pad  & n61 ;
  assign n63 = n54 & n62 ;
  assign n64 = ~n59 & ~n63 ;
  assign n65 = ~\G3_pad  & ~n64 ;
  assign n66 = ~n58 & ~n65 ;
  assign n67 = ~\G2_pad  & ~n66 ;
  assign n68 = n43 & n67 ;
  assign n69 = \G3_pad  & n68 ;
  assign n70 = ~\G1_pad  & \G2_pad  ;
  assign n71 = \G3_pad  & \G5_pad  ;
  assign n72 = \G4_pad  & ~n71 ;
  assign n73 = \G2_pad  & ~\G3_pad  ;
  assign n74 = ~\G2_pad  & \G3_pad  ;
  assign n75 = ~n73 & ~n74 ;
  assign n76 = ~n72 & n75 ;
  assign n77 = \G6_pad  & ~n76 ;
  assign n78 = \G4_pad  & ~\G5_pad  ;
  assign n79 = ~\G3_pad  & n78 ;
  assign n80 = ~n77 & ~n79 ;
  assign n81 = \G1_pad  & ~n80 ;
  assign n90 = \G1_pad  & ~\G4_pad  ;
  assign n91 = ~\G2_pad  & ~n90 ;
  assign n88 = \G1_pad  & \G4_pad  ;
  assign n89 = ~\G5_pad  & ~n88 ;
  assign n92 = ~\G6_pad  & ~n89 ;
  assign n93 = ~n91 & n92 ;
  assign n82 = ~\G4_pad  & \G6_pad  ;
  assign n83 = ~\G5_pad  & ~n82 ;
  assign n84 = n70 & ~n83 ;
  assign n85 = \G1_pad  & \G3_pad  ;
  assign n86 = \G5_pad  & ~n60 ;
  assign n87 = n85 & n86 ;
  assign n94 = ~n84 & ~n87 ;
  assign n95 = ~n93 & n94 ;
  assign n96 = ~n81 & n95 ;
  assign n97 = ~n41 & ~n96 ;
  assign n98 = \G11_pad  & ~\G9_pad  ;
  assign n99 = ~\G10_pad  & \G7_pad  ;
  assign n100 = \G8_pad  & n99 ;
  assign n101 = n98 & n100 ;
  assign n102 = ~\G7_pad  & ~\G8_pad  ;
  assign n103 = \G10_pad  & n34 ;
  assign n104 = n102 & n103 ;
  assign n105 = ~n101 & ~n104 ;
  assign n106 = \G3_pad  & \G6_pad  ;
  assign n107 = ~\G1_pad  & \G4_pad  ;
  assign n108 = ~n90 & ~n107 ;
  assign n109 = n106 & ~n108 ;
  assign n110 = ~n105 & n109 ;
  assign n111 = ~\G1_pad  & \G3_pad  ;
  assign n112 = n51 & n60 ;
  assign n113 = n35 & n112 ;
  assign n114 = ~\G8_pad  & n99 ;
  assign n115 = ~\G4_pad  & ~\G6_pad  ;
  assign n116 = n98 & n115 ;
  assign n117 = n114 & n116 ;
  assign n118 = ~n113 & ~n117 ;
  assign n119 = n111 & ~n118 ;
  assign n120 = ~n110 & ~n119 ;
  assign n121 = \G2_pad  & ~\G5_pad  ;
  assign n122 = ~n120 & n121 ;
  assign n123 = ~\G10_pad  & ~\G11_pad  ;
  assign n124 = n102 & n123 ;
  assign n125 = \G9_pad  & n124 ;
  assign n126 = n35 & n36 ;
  assign n127 = ~n125 & ~n126 ;
  assign n128 = n60 & n71 ;
  assign n129 = ~n127 & n128 ;
  assign n130 = \G1_pad  & \G2_pad  ;
  assign n131 = n129 & n130 ;
  assign n132 = ~n122 & ~n131 ;
  assign n133 = ~n97 & ~n132 ;
  assign n134 = \G13_pad  & n133 ;
  assign n135 = n70 & n134 ;
  assign n136 = ~n69 & ~n135 ;
  assign n137 = \G6_pad  & n78 ;
  assign n138 = n104 & n137 ;
  assign n139 = ~n136 & n138 ;
  assign n147 = ~\G4_pad  & ~\G5_pad  ;
  assign n148 = \G11_pad  & n147 ;
  assign n149 = \G35_reg/NET0131  & \G3_pad  ;
  assign n150 = n148 & n149 ;
  assign n151 = ~n129 & ~n150 ;
  assign n152 = \G2_pad  & ~n151 ;
  assign n153 = ~n67 & ~n152 ;
  assign n154 = n43 & ~n153 ;
  assign n155 = \G13_pad  & \G1_pad  ;
  assign n156 = n133 & n155 ;
  assign n157 = ~n154 & ~n156 ;
  assign n158 = \G4_pad  & \G5_pad  ;
  assign n159 = n125 & n158 ;
  assign n160 = n54 & n148 ;
  assign n161 = ~n159 & ~n160 ;
  assign n162 = \G2_pad  & n106 ;
  assign n163 = ~n161 & n162 ;
  assign n164 = ~n157 & n163 ;
  assign n140 = \G13_pad  & ~\G43_reg/NET0131  ;
  assign n141 = n97 & n140 ;
  assign n142 = n61 & n101 ;
  assign n143 = \G36_reg/NET0131  & n115 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = ~\G3_pad  & ~n144 ;
  assign n146 = n68 & n145 ;
  assign n165 = ~n141 & ~n146 ;
  assign n166 = ~n164 & n165 ;
  assign n167 = ~n139 & n166 ;
  assign n168 = ~\G12_pad  & ~n167 ;
  assign n169 = \G12_pad  & ~\G13_pad  ;
  assign n178 = ~\G6_pad  & \G7_pad  ;
  assign n179 = \G30_reg/NET0131  & n178 ;
  assign n180 = ~\G10_pad  & ~n179 ;
  assign n181 = ~\G9_pad  & ~n180 ;
  assign n174 = \G31_reg/NET0131  & \G8_pad  ;
  assign n175 = ~\G10_pad  & ~\G8_pad  ;
  assign n176 = ~\G7_pad  & ~n175 ;
  assign n177 = \G9_pad  & ~n176 ;
  assign n182 = ~n174 & ~n177 ;
  assign n183 = ~n181 & n182 ;
  assign n184 = ~\G11_pad  & ~n183 ;
  assign n186 = ~\G31_reg/NET0131  & ~n179 ;
  assign n187 = \G8_pad  & ~n186 ;
  assign n188 = \G10_pad  & \G8_pad  ;
  assign n189 = \G9_pad  & ~n188 ;
  assign n190 = ~n48 & ~n189 ;
  assign n191 = ~n187 & n190 ;
  assign n185 = ~\G30_reg/NET0131  & ~\G6_pad  ;
  assign n192 = \G11_pad  & ~n185 ;
  assign n193 = ~n191 & n192 ;
  assign n194 = ~n184 & ~n193 ;
  assign n170 = \G0_pad  & \G3_pad  ;
  assign n171 = ~\G3_pad  & \G5_pad  ;
  assign n172 = ~\G4_pad  & ~n171 ;
  assign n173 = ~n170 & n172 ;
  assign n195 = \G46_reg/NET0131  & ~n173 ;
  assign n196 = ~n194 & n195 ;
  assign n197 = n169 & n196 ;
  assign n198 = \G3_pad  & ~\G4_pad  ;
  assign n199 = ~\G2_pad  & \G5_pad  ;
  assign n200 = ~n198 & ~n199 ;
  assign n201 = \G1_pad  & ~n200 ;
  assign n204 = ~\G2_pad  & n71 ;
  assign n202 = ~\G3_pad  & ~\G5_pad  ;
  assign n203 = \G2_pad  & ~n85 ;
  assign n205 = ~n202 & ~n203 ;
  assign n206 = ~n204 & n205 ;
  assign n207 = \G4_pad  & ~n206 ;
  assign n208 = ~n201 & ~n207 ;
  assign n209 = \G0_pad  & ~n208 ;
  assign n210 = n197 & n209 ;
  assign n211 = ~n168 & ~n210 ;
  assign n212 = ~\G5_pad  & n115 ;
  assign n213 = n123 & n212 ;
  assign n214 = n61 & n103 ;
  assign n215 = ~n213 & ~n214 ;
  assign n216 = n102 & ~n215 ;
  assign n217 = ~\G6_pad  & n36 ;
  assign n218 = n35 & n78 ;
  assign n219 = n217 & n218 ;
  assign n220 = ~n216 & ~n219 ;
  assign n221 = ~\G3_pad  & ~n220 ;
  assign n222 = n46 & n54 ;
  assign n223 = \G11_pad  & n222 ;
  assign n224 = ~n221 & ~n223 ;
  assign n225 = ~\G12_pad  & n68 ;
  assign n226 = ~n224 & n225 ;
  assign n227 = \G11_pad  & \G2_pad  ;
  assign n228 = \G6_pad  & \G9_pad  ;
  assign n229 = \G4_pad  & n36 ;
  assign n230 = n228 & n229 ;
  assign n231 = n71 & n230 ;
  assign n232 = ~\G9_pad  & n99 ;
  assign n233 = n106 & n147 ;
  assign n234 = n232 & n233 ;
  assign n235 = ~n231 & ~n234 ;
  assign n236 = \G8_pad  & ~n235 ;
  assign n237 = ~n157 & n236 ;
  assign n238 = ~\G1_pad  & n134 ;
  assign n239 = n222 & n238 ;
  assign n240 = ~n237 & ~n239 ;
  assign n241 = ~\G12_pad  & ~n240 ;
  assign n242 = n169 & ~n196 ;
  assign n243 = ~\G0_pad  & ~\G4_pad  ;
  assign n246 = \G10_pad  & ~\G8_pad  ;
  assign n247 = n202 & n246 ;
  assign n244 = \G6_pad  & ~\G9_pad  ;
  assign n245 = \G11_pad  & ~\G7_pad  ;
  assign n248 = n244 & n245 ;
  assign n249 = n247 & n248 ;
  assign n250 = \G11_pad  & \G37_reg/NET0131  ;
  assign n251 = n71 & n250 ;
  assign n252 = n100 & n251 ;
  assign n253 = ~n249 & ~n252 ;
  assign n254 = n243 & ~n253 ;
  assign n255 = n61 & n170 ;
  assign n256 = n126 & n255 ;
  assign n257 = ~n254 & ~n256 ;
  assign n258 = n130 & ~n257 ;
  assign n259 = n242 & n258 ;
  assign n260 = \G0_pad  & n230 ;
  assign n261 = \G38_reg/NET0131  & n244 ;
  assign n262 = ~n260 & ~n261 ;
  assign n263 = \G1_pad  & \G8_pad  ;
  assign n264 = n71 & n263 ;
  assign n265 = ~n262 & n264 ;
  assign n266 = n259 & n265 ;
  assign n267 = ~n241 & ~n266 ;
  assign n268 = n227 & ~n267 ;
  assign n269 = ~n226 & ~n268 ;
  assign n274 = ~\G12_pad  & n43 ;
  assign n275 = n153 & n274 ;
  assign n270 = n242 & ~n258 ;
  assign n271 = ~\G12_pad  & \G13_pad  ;
  assign n272 = ~n97 & n271 ;
  assign n273 = n132 & n272 ;
  assign n276 = ~n270 & ~n273 ;
  assign n277 = ~n275 & n276 ;
  assign n280 = \G34_reg/NET0131  & \G8_pad  ;
  assign n281 = \G6_pad  & n197 ;
  assign n282 = ~n280 & ~n281 ;
  assign n283 = n39 & ~n282 ;
  assign n278 = \G34_reg/NET0131  & n36 ;
  assign n279 = ~n49 & n278 ;
  assign n289 = ~\G8_pad  & n103 ;
  assign n284 = \G11_pad  & ~n48 ;
  assign n285 = ~\G9_pad  & ~n123 ;
  assign n286 = ~n284 & n285 ;
  assign n287 = \G7_pad  & \G9_pad  ;
  assign n288 = n188 & ~n287 ;
  assign n290 = ~n286 & ~n288 ;
  assign n291 = ~n289 & n290 ;
  assign n292 = n281 & ~n291 ;
  assign n293 = ~n279 & ~n292 ;
  assign n294 = ~n283 & n293 ;
  assign n295 = n197 & n217 ;
  assign n297 = ~\G7_pad  & ~n188 ;
  assign n296 = \G8_pad  & n36 ;
  assign n298 = \G34_reg/NET0131  & ~n296 ;
  assign n299 = ~n297 & n298 ;
  assign n300 = ~n295 & ~n299 ;
  assign n301 = \G9_pad  & ~n300 ;
  assign n304 = n32 & ~n50 ;
  assign n305 = ~n123 & n304 ;
  assign n302 = ~n34 & ~n38 ;
  assign n303 = ~\G8_pad  & ~n302 ;
  assign n306 = ~n39 & ~n303 ;
  assign n307 = ~n305 & n306 ;
  assign n308 = n281 & ~n307 ;
  assign n309 = ~n301 & ~n308 ;
  assign n310 = ~\G42_reg/NET0131  & n197 ;
  assign n311 = \G7_pad  & ~n50 ;
  assign n312 = ~n189 & n311 ;
  assign n313 = \G11_pad  & \G34_reg/NET0131  ;
  assign n314 = ~n102 & n313 ;
  assign n315 = ~n55 & n314 ;
  assign n316 = ~n312 & n315 ;
  assign n317 = ~n310 & ~n316 ;
  assign n318 = n97 & n271 ;
  assign n319 = \G1_pad  & n318 ;
  assign n326 = ~\G5_pad  & ~\G6_pad  ;
  assign n325 = ~\G2_pad  & \G6_pad  ;
  assign n327 = ~n106 & ~n325 ;
  assign n328 = ~n326 & n327 ;
  assign n329 = ~n71 & ~n328 ;
  assign n330 = ~\G4_pad  & ~n329 ;
  assign n320 = ~\G3_pad  & n60 ;
  assign n321 = ~n74 & ~n320 ;
  assign n322 = \G5_pad  & ~n321 ;
  assign n323 = \G2_pad  & \G4_pad  ;
  assign n324 = ~\G5_pad  & n323 ;
  assign n331 = ~n322 & ~n324 ;
  assign n332 = ~n330 & n331 ;
  assign n333 = n319 & ~n332 ;
  assign n334 = n88 & ~n170 ;
  assign n335 = n197 & n334 ;
  assign n336 = ~\G13_pad  & ~\G33_reg/NET0131  ;
  assign n337 = \G3_pad  & n336 ;
  assign n339 = ~\G12_pad  & n42 ;
  assign n340 = ~\G13_pad  & n339 ;
  assign n338 = \G2_pad  & \G5_pad  ;
  assign n341 = ~n45 & n338 ;
  assign n342 = n340 & n341 ;
  assign n343 = ~n337 & ~n342 ;
  assign n344 = ~n335 & n343 ;
  assign n345 = ~n333 & n344 ;
  assign n353 = \G5_pad  & n88 ;
  assign n354 = \G2_pad  & ~n89 ;
  assign n355 = ~n353 & n354 ;
  assign n356 = n318 & n355 ;
  assign n346 = \G0_pad  & ~\G29_reg/NET0131  ;
  assign n347 = ~\G0_pad  & n88 ;
  assign n348 = \G3_pad  & n347 ;
  assign n349 = ~n346 & ~n348 ;
  assign n350 = n197 & ~n349 ;
  assign n351 = n71 & ~n323 ;
  assign n352 = n340 & n351 ;
  assign n357 = ~n337 & ~n352 ;
  assign n358 = ~n350 & n357 ;
  assign n359 = ~n356 & n358 ;
  assign n361 = \G0_pad  & \G2_pad  ;
  assign n363 = ~\G4_pad  & n361 ;
  assign n362 = ~\G1_pad  & ~n361 ;
  assign n364 = ~\G3_pad  & ~n362 ;
  assign n365 = ~n363 & n364 ;
  assign n360 = ~n88 & n170 ;
  assign n366 = ~n347 & ~n360 ;
  assign n367 = ~n365 & n366 ;
  assign n368 = n197 & ~n367 ;
  assign n369 = ~\G2_pad  & ~n85 ;
  assign n370 = \G4_pad  & ~n130 ;
  assign n371 = ~n369 & n370 ;
  assign n372 = n318 & n371 ;
  assign n373 = ~n368 & ~n372 ;
  assign n374 = \G5_pad  & ~n373 ;
  assign n376 = n44 & n74 ;
  assign n375 = ~n74 & n78 ;
  assign n377 = ~n320 & ~n375 ;
  assign n378 = ~n376 & n377 ;
  assign n379 = n319 & ~n378 ;
  assign n380 = \G39_reg/NET0131  & \G4_pad  ;
  assign n381 = n340 & n380 ;
  assign n382 = ~n379 & ~n381 ;
  assign n383 = ~n374 & n382 ;
  assign n384 = ~\G1_pad  & \G5_pad  ;
  assign n385 = \G4_pad  & ~n384 ;
  assign n386 = n203 & ~n385 ;
  assign n387 = ~\G4_pad  & \G5_pad  ;
  assign n388 = n85 & n387 ;
  assign n389 = ~n386 & ~n388 ;
  assign n390 = n318 & ~n389 ;
  assign n391 = n74 & ~n78 ;
  assign n392 = \G2_pad  & ~n147 ;
  assign n393 = \G5_pad  & n45 ;
  assign n394 = n392 & ~n393 ;
  assign n395 = ~n391 & ~n394 ;
  assign n396 = n340 & ~n395 ;
  assign n397 = ~n390 & ~n396 ;
  assign n398 = \G6_pad  & ~n397 ;
  assign n399 = ~\G40_reg/NET0131  & n197 ;
  assign n400 = n60 & ~n338 ;
  assign n401 = n319 & n400 ;
  assign n402 = ~n399 & ~n401 ;
  assign n403 = ~n398 & n402 ;
  assign n404 = n65 & n225 ;
  assign n406 = ~\G0_pad  & n172 ;
  assign n405 = \G0_pad  & ~n198 ;
  assign n407 = \G1_pad  & ~n405 ;
  assign n408 = ~n406 & n407 ;
  assign n409 = ~n72 & ~n384 ;
  assign n410 = \G0_pad  & ~n409 ;
  assign n411 = ~n408 & ~n410 ;
  assign n412 = \G2_pad  & ~n411 ;
  assign n413 = n197 & n412 ;
  assign n414 = ~n404 & ~n413 ;
  assign n415 = \G3_pad  & ~n78 ;
  assign n416 = ~n338 & ~n375 ;
  assign n417 = ~n415 & n416 ;
  assign n418 = \G0_pad  & ~n417 ;
  assign n419 = ~\G1_pad  & ~n418 ;
  assign n420 = ~\G10_pad  & ~\G30_reg/NET0131  ;
  assign n421 = \G7_pad  & ~n420 ;
  assign n422 = ~\G6_pad  & ~n421 ;
  assign n423 = n111 & ~n387 ;
  assign n424 = ~n78 & n405 ;
  assign n425 = ~n423 & ~n424 ;
  assign n426 = \G2_pad  & n409 ;
  assign n427 = ~n425 & n426 ;
  assign n428 = ~n422 & ~n427 ;
  assign n429 = ~n419 & n428 ;
  assign n430 = ~n318 & ~n340 ;
  assign n432 = \G10_pad  & \G11_pad  ;
  assign n431 = ~\G11_pad  & ~\G7_pad  ;
  assign n433 = \G9_pad  & ~n431 ;
  assign n434 = ~n432 & n433 ;
  assign n435 = ~\G31_reg/NET0131  & ~n434 ;
  assign n436 = \G6_pad  & ~n435 ;
  assign n437 = ~n179 & ~n436 ;
  assign n438 = \G8_pad  & ~n437 ;
  assign n440 = \G6_pad  & n188 ;
  assign n441 = ~n48 & ~n440 ;
  assign n442 = ~\G9_pad  & ~n441 ;
  assign n439 = ~n36 & n228 ;
  assign n443 = ~n38 & n178 ;
  assign n444 = ~n439 & ~n443 ;
  assign n445 = ~n442 & n444 ;
  assign n446 = \G11_pad  & ~n445 ;
  assign n447 = ~n86 & ~n325 ;
  assign n448 = ~n324 & n447 ;
  assign n449 = \G1_pad  & ~n448 ;
  assign n450 = ~n84 & ~n449 ;
  assign n451 = \G3_pad  & ~n450 ;
  assign n453 = n61 & n104 ;
  assign n452 = n126 & n212 ;
  assign n454 = ~\G9_pad  & n326 ;
  assign n455 = n124 & n454 ;
  assign n456 = ~n452 & ~n455 ;
  assign n457 = ~n453 & n456 ;
  assign n458 = ~n124 & ~n126 ;
  assign n459 = ~\G5_pad  & ~n458 ;
  assign n460 = n74 & ~n83 ;
  assign n461 = ~n128 & n392 ;
  assign n462 = ~n460 & ~n461 ;
  assign n463 = ~n45 & ~n387 ;
  assign n464 = n70 & ~n463 ;
  assign n465 = ~n391 & ~n464 ;
  assign n466 = n99 & n243 ;
  assign n467 = \G2_pad  & ~n71 ;
  assign n468 = ~n204 & ~n467 ;
  assign n469 = \G10_pad  & ~n34 ;
  assign n470 = ~n245 & ~n469 ;
  assign n471 = ~\G10_pad  & ~n98 ;
  assign n472 = ~\G6_pad  & ~\G9_pad  ;
  assign n473 = ~n228 & ~n472 ;
  assign n474 = ~n134 & ~n154 ;
  assign n475 = ~\G12_pad  & ~n474 ;
  assign n476 = ~n259 & ~n475 ;
  assign n477 = ~n55 & ~n232 ;
  assign n478 = \G8_pad  & ~n477 ;
  assign n479 = n47 & n478 ;
  assign n480 = ~\G3_pad  & ~\G44_reg/NET0131  ;
  assign n481 = ~n479 & ~n480 ;
  assign n482 = n225 & ~n481 ;
  assign n483 = n54 & n147 ;
  assign n484 = ~n157 & n483 ;
  assign n485 = n238 & n478 ;
  assign n486 = ~n484 & ~n485 ;
  assign n487 = ~\G12_pad  & n106 ;
  assign n488 = ~n486 & n487 ;
  assign n489 = \G37_reg/NET0131  & \G38_reg/NET0131  ;
  assign n490 = n264 & n489 ;
  assign n491 = n259 & n490 ;
  assign n492 = ~n488 & ~n491 ;
  assign n493 = n227 & ~n492 ;
  assign n494 = ~n482 & ~n493 ;
  assign n495 = n36 & ~n228 ;
  assign n496 = n197 & n495 ;
  assign n497 = \G34_reg/NET0131  & n288 ;
  assign n498 = ~n496 & ~n497 ;
  assign n499 = ~n283 & n498 ;
  assign n500 = n324 & n339 ;
  assign n501 = \G0_pad  & \G12_pad  ;
  assign n502 = n90 & n501 ;
  assign n503 = n196 & n502 ;
  assign n504 = ~n500 & ~n503 ;
  assign n505 = \G6_pad  & n54 ;
  assign n506 = n114 & n472 ;
  assign n507 = ~n505 & ~n506 ;
  assign \G532_pad  = ~n211 ;
  assign \G537_pad  = ~n269 ;
  assign \G539_pad  = ~n277 ;
  assign \G542_pad  = ~n294 ;
  assign \G546_pad  = ~\G41_reg/NET0131  ;
  assign \G547_pad  = ~n309 ;
  assign \G548_pad  = ~n317 ;
  assign \G549_pad  = ~n345 ;
  assign \G550_pad  = ~n359 ;
  assign \G551_pad  = ~n383 ;
  assign \G552_pad  = ~n403 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1667/_3_  = ~n414 ;
  assign \g1737/_0_  = n429 ;
  assign \g1744/_0_  = ~n430 ;
  assign \g1787/_0_  = ~n438 ;
  assign \g1811/_0_  = ~n446 ;
  assign \g1830/_0_  = ~n451 ;
  assign \g1831/_0_  = n457 ;
  assign \g1846/_0_  = n459 ;
  assign \g1852/_0_  = ~n462 ;
  assign \g1866/_0_  = n465 ;
  assign \g19/_2_  = n466 ;
  assign \g1931/_0_  = ~n468 ;
  assign \g1945/_0_  = ~n470 ;
  assign \g2014/_0_  = ~n471 ;
  assign \g2015/_0_  = n473 ;
  assign \g2643/_0_  = ~n476 ;
  assign \g2859/_1_  = ~n494 ;
  assign \g3397/_2_  = n499 ;
  assign \g3546/_0_  = n504 ;
  assign \g3606/_3_  = ~n507 ;
endmodule
