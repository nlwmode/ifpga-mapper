module top( \g1002_reg/NET0131  , \g1008_reg/NET0131  , \g10122_pad  , \g1018_reg/NET0131  , \g1024_reg/NET0131  , \g10306_pad  , \g1030_reg/NET0131  , \g1036_reg/NET0131  , \g1041_reg/NET0131  , \g1046_reg/NET0131  , \g10500_pad  , \g10527_pad  , \g1052_reg/NET0131  , \g1061_reg/NET0131  , \g1070_reg/NET0131  , \g1087_reg/NET0131  , \g1094_reg/NET0131  , \g1099_reg/NET0131  , \g1105_reg/NET0131  , \g1111_reg/NET0131  , \g1124_reg/NET0131  , \g1129_reg/NET0131  , \g1135_reg/NET0131  , \g1141_reg/NET0131  , \g11447_pad  , \g1146_reg/NET0131  , \g1152_reg/NET0131  , \g1171_reg/NET0131  , \g11770_pad  , \g1178_reg/NET0131  , \g1183_reg/NET0131  , \g1189_reg/NET0131  , \g1193_reg/NET0131  , \g1199_reg/NET0131  , \g1205_reg/NET0131  , \g1211_reg/NET0131  , \g1216_reg/NET0131  , \g12184_pad  , \g1221_reg/NET0131  , \g1236_reg/NET0131  , \g1242_reg/NET0131  , \g1246_reg/NET0131  , \g12919_pad  , \g12923_pad  , \g1300_reg/NET0131  , \g13039_pad  , \g1306_reg/NET0131  , \g1312_reg/NET0131  , \g1319_reg/NET0131  , \g1322_reg/NET0131  , \g13259_pad  , \g13272_pad  , \g1333_reg/NET0131  , \g1339_reg/NET0131  , \g1345_reg/NET0131  , \g1351_reg/NET0131  , \g1361_reg/NET0131  , \g1367_reg/NET0131  , \g1373_reg/NET0131  , \g1379_reg/NET0131  , \g1384_reg/NET0131  , \g13865_pad  , \g13895_pad  , \g1389_reg/NET0131  , \g1395_reg/NET0131  , \g1404_reg/NET0131  , \g14096_pad  , \g14125_pad  , \g1413_reg/NET0131  , \g14147_pad  , \g14167_pad  , \g14189_pad  , \g14201_pad  , \g14217_pad  , \g142_reg/NET0131  , \g1430_reg/NET0131  , \g1437_reg/NET0131  , \g1442_reg/NET0131  , \g1448_reg/NET0131  , \g1454_reg/NET0131  , \g1467_reg/NET0131  , \g146_reg/NET0131  , \g1472_reg/NET0131  , \g1478_reg/NET0131  , \g1484_reg/NET0131  , \g1489_reg/NET0131  , \g1495_reg/NET0131  , \g150_reg/NET0131  , \g1514_reg/NET0131  , \g1521_reg/NET0131  , \g1526_reg/NET0131  , \g1532_reg/NET0131  , \g1536_reg/NET0131  , \g153_reg/NET0131  , \g1542_reg/NET0131  , \g1548_reg/NET0131  , \g1554_reg/NET0131  , \g1559_reg/NET0131  , \g1564_reg/NET0131  , \g1579_reg/NET0131  , \g157_reg/NET0131  , \g1585_reg/NET0131  , \g1589_reg/NET0131  , \g1592_reg/NET0131  , \g1600_reg/NET0131  , \g1604_reg/NET0131  , \g1608_reg/NET0131  , \g160_reg/NET0131  , \g1612_reg/NET0131  , \g1616_reg/NET0131  , \g1620_reg/NET0131  , \g1624_reg/NET0131  , \g1632_reg/NET0131  , \g1636_reg/NET0131  , \g1644_reg/NET0131  , \g1648_reg/NET0131  , \g164_reg/NET0131  , \g1657_reg/NET0131  , \g16603_pad  , \g16624_pad  , \g1664_reg/NET0131  , \g16686_pad  , \g1668_reg/NET0131  , \g16718_pad  , \g1677_reg/NET0131  , \g1682_reg/NET0131  , \g16874_pad  , \g1687_reg/NET0131  , \g168_reg/NET0131  , \g1691_reg/NET0131  , \g1696_reg/NET0131  , \g1700_reg/NET0131  , \g1706_reg/NET0131  , \g1710_reg/NET0131  , \g1714_reg/NET0131  , \g1720_reg/NET0131  , \g1724_reg/NET0131  , \g1728_reg/NET0131  , \g17291_pad  , \g17316_pad  , \g17320_pad  , \g1736_reg/NET0131  , \g17400_pad  , \g17404_pad  , \g1740_reg/NET0131  , \g17423_pad  , \g1744_reg/NET0131  , \g1748_reg/NET0131  , \g174_reg/NET0131  , \g1752_reg/NET0131  , \g1756_reg/NET0131  , \g1760_reg/NET0131  , \g1768_reg/NET0131  , \g1772_reg/NET0131  , \g1779_reg/NET0131  , \g1783_reg/NET0131  , \g1792_reg/NET0131  , \g1798_reg/NET0131  , \g1802_reg/NET0131  , \g18094_pad  , \g18095_pad  , \g18096_pad  , \g18098_pad  , \g18099_pad  , \g1811_reg/NET0131  , \g1816_reg/NET0131  , \g1821_reg/NET0131  , \g1825_reg/NET0131  , \g182_reg/NET0131  , \g1830_reg/NET0131  , \g1834_reg/NET0131  , \g1840_reg/NET0131  , \g1844_reg/NET0131  , \g1848_reg/NET0131  , \g1854_reg/NET0131  , \g1858_reg/NET0131  , \g1862_reg/NET0131  , \g1870_reg/NET0131  , \g1874_reg/NET0131  , \g1878_reg/NET0131  , \g1882_reg/NET0131  , \g1886_reg/NET0131  , \g1890_reg/NET0131  , \g1894_reg/NET0131  , \g1902_reg/NET0131  , \g1906_reg/NET0131  , \g1913_reg/NET0131  , \g1917_reg/NET0131  , \g191_reg/NET0131  , \g1926_reg/NET0131  , \g1932_reg/NET0131  , \g19334_pad  , \g19357_pad  , \g1936_reg/NET0131  , \g1945_reg/NET0131  , \g1950_reg/NET0131  , \g1955_reg/NET0131  , \g1959_reg/NET0131  , \g1964_reg/NET0131  , \g1968_reg/NET0131  , \g1974_reg/NET0131  , \g1978_reg/NET0131  , \g1982_reg/NET0131  , \g1988_reg/NET0131  , \g1992_reg/NET0131  , \g1996_reg/NET0131  , \g2004_reg/NET0131  , \g2008_reg/NET0131  , \g2012_reg/NET0131  , \g2016_reg/NET0131  , \g2020_reg/NET0131  , \g2024_reg/NET0131  , \g2028_reg/NET0131  , \g2036_reg/NET0131  , \g203_reg/NET0131  , \g2040_reg/NET0131  , \g2047_reg/NET0131  , \g2051_reg/NET0131  , \g2060_reg/NET0131  , \g2066_reg/NET0131  , \g2070_reg/NET0131  , \g2079_reg/NET0131  , \g2084_reg/NET0131  , \g2089_reg/NET0131  , \g2093_reg/NET0131  , \g2098_reg/NET0131  , \g209_reg/NET0131  , \g2102_reg/NET0131  , \g2108_reg/NET0131  , \g2112_reg/NET0131  , \g2116_reg/NET0131  , \g2122_reg/NET0131  , \g2126_reg/NET0131  , \g2153_reg/NET0131  , \g2161_reg/NET0131  , \g2165_reg/NET0131  , \g2169_reg/NET0131  , \g2173_reg/NET0131  , \g2177_reg/NET0131  , \g2181_reg/NET0131  , \g2185_reg/NET0131  , \g218_reg/NET0131  , \g2193_reg/NET0131  , \g2197_reg/NET0131  , \g2204_reg/NET0131  , \g2208_reg/NET0131  , \g2217_reg/NET0131  , \g2223_reg/NET0131  , \g2227_reg/NET0131  , \g222_reg/NET0131  , \g2236_reg/NET0131  , \g2241_reg/NET0131  , \g2246_reg/NET0131  , \g2250_reg/NET0131  , \g2255_reg/NET0131  , \g2259_reg/NET0131  , \g225_reg/NET0131  , \g2265_reg/NET0131  , \g2269_reg/NET0131  , \g2273_reg/NET0131  , \g2279_reg/NET0131  , \g2283_reg/NET0131  , \g2287_reg/NET0131  , \g2295_reg/NET0131  , \g2299_reg/NET0131  , \g2303_reg/NET0131  , \g2307_reg/NET0131  , \g2311_reg/NET0131  , \g2315_reg/NET0131  , \g2319_reg/NET0131  , \g2327_reg/NET0131  , \g232_reg/NET0131  , \g2331_reg/NET0131  , \g2338_reg/NET0131  , \g2342_reg/NET0131  , \g2351_reg/NET0131  , \g2357_reg/NET0131  , \g2361_reg/NET0131  , \g2370_reg/NET0131  , \g2375_reg/NET0131  , \g2380_reg/NET0131  , \g2384_reg/NET0131  , \g2389_reg/NET0131  , \g2393_reg/NET0131  , \g2399_reg/NET0131  , \g239_reg/NET0131  , \g2403_reg/NET0131  , \g2407_reg/NET0131  , \g2413_reg/NET0131  , \g2417_reg/NET0131  , \g2421_reg/NET0131  , \g2429_reg/NET0131  , \g2433_reg/NET0131  , \g2437_reg/NET0131  , \g2441_reg/NET0131  , \g2445_reg/NET0131  , \g2449_reg/NET0131  , \g2453_reg/NET0131  , \g2461_reg/NET0131  , \g2465_reg/NET0131  , \g246_reg/NET0131  , \g2472_reg/NET0131  , \g2476_reg/NET0131  , \g2485_reg/NET0131  , \g2491_reg/NET0131  , \g2495_reg/NET0131  , \g2504_reg/NET0131  , \g2509_reg/NET0131  , \g2514_reg/NET0131  , \g2518_reg/NET0131  , \g2523_reg/NET0131  , \g2527_reg/NET0131  , \g2533_reg/NET0131  , \g2537_reg/NET0131  , \g2541_reg/NET0131  , \g2547_reg/NET0131  , \g2551_reg/NET0131  , \g2555_reg/NET0131  , \g255_reg/NET0131  , \g2563_reg/NET0131  , \g2567_reg/NET0131  , \g2571_reg/NET0131  , \g2575_reg/NET0131  , \g2579_reg/NET0131  , \g2583_reg/NET0131  , \g2587_reg/NET0131  , \g2595_reg/NET0131  , \g2599_reg/NET0131  , \g2606_reg/NET0131  , \g2610_reg/NET0131  , \g2619_reg/NET0131  , \g2625_reg/NET0131  , \g2629_reg/NET0131  , \g262_reg/NET0131  , \g2638_reg/NET0131  , \g2643_reg/NET0131  , \g2648_reg/NET0131  , \g2652_reg/NET0131  , \g2657_reg/NET0131  , \g2661_reg/NET0131  , \g2667_reg/NET0131  , \g2671_reg/NET0131  , \g2675_reg/NET0131  , \g2681_reg/NET0131  , \g2685_reg/NET0131  , \g269_reg/NET0131  , \g2715_reg/NET0131  , \g2719_reg/NET0131  , \g2724_reg/NET0131  , \g2729_reg/NET0131  , \g2735_reg/NET0131  , \g2741_reg/NET0131  , \g2748_reg/NET0131  , \g2756_reg/NET0131  , \g2759_reg/NET0131  , \g2763_reg/NET0131  , \g2767_reg/NET0131  , \g2771_reg/NET0131  , \g2775_reg/NET0131  , \g2779_reg/NET0131  , \g2783_reg/NET0131  , \g2787_reg/NET0131  , \g278_reg/NET0131  , \g2791_reg/NET0131  , \g2795_reg/NET0131  , \g2799_reg/NET0131  , \g2803_reg/NET0131  , \g2807_reg/NET0131  , \g2811_reg/NET0131  , \g2815_reg/NET0131  , \g2819_reg/NET0131  , \g2823_reg/NET0131  , \g2827_reg/NET0131  , \g2831_reg/NET0131  , \g2834_reg/NET0131  , \g283_reg/NET0131  , \g2848_reg/NET0131  , \g2856_reg/NET0131  , \g2864_reg/NET0131  , \g2873_reg/NET0131  , \g2878_reg/NET0131  , \g287_reg/NET0131  , \g2882_reg/NET0131  , \g2886_reg/NET0131  , \g2898_reg/NET0131  , \g2902_reg/NET0131  , \g2907_reg/NET0131  , \g2912_reg/NET0131  , \g2917_reg/NET0131  , \g291_reg/NET0131  , \g29211_pad  , \g29212_pad  , \g29213_pad  , \g29214_pad  , \g29215_pad  , \g29216_pad  , \g29218_pad  , \g29219_pad  , \g29220_pad  , \g29221_pad  , \g2922_reg/NET0131  , \g2927_reg/NET0131  , \g2932_reg/NET0131  , \g2936_reg/NET0131  , \g2941_reg/NET0131  , \g2946_reg/NET0131  , \g294_reg/NET0131  , \g2950_reg/NET0131  , \g2955_reg/NET0131  , \g2960_reg/NET0131  , \g2965_reg/NET0131  , \g2970_reg/NET0131  , \g2975_reg/NET0131  , \g2980_reg/NET0131  , \g2984_reg/NET0131  , \g2988_reg/NET0131  , \g298_reg/NET0131  , \g2999_reg/NET0131  , \g3003_reg/NET0131  , \g301_reg/NET0131  , \g3050_reg/NET0131  , \g305_reg/NET0131  , \g3096_reg/NET0131  , \g3100_reg/NET0131  , \g3106_reg/NET0131  , \g3111_reg/NET0131  , \g3115_reg/NET0131  , \g3119_reg/NET0131  , \g311_reg/NET0131  , \g3125_reg/NET0131  , \g3129_reg/NET0131  , \g3133_reg/NET0131  , \g3139_reg/NET0131  , \g3143_reg/NET0131  , \g3147_reg/NET0131  , \g3155_reg/NET0131  , \g3161_reg/NET0131  , \g3167_reg/NET0131  , \g316_reg/NET0131  , \g3171_reg/NET0131  , \g3179_reg/NET0131  , \g3187_reg/NET0131  , \g3191_reg/NET0131  , \g3195_reg/NET0131  , \g3199_reg/NET0131  , \g319_reg/NET0131  , \g3203_reg/NET0131  , \g3207_reg/NET0131  , \g3211_reg/NET0131  , \g3215_reg/NET0131  , \g3219_reg/NET0131  , \g3223_reg/NET0131  , \g3227_reg/NET0131  , \g3231_reg/NET0131  , \g3235_reg/NET0131  , \g3239_reg/NET0131  , \g3243_reg/NET0131  , \g3247_reg/NET0131  , \g324_reg/NET0131  , \g3251_reg/NET0131  , \g3255_reg/NET0131  , \g3259_reg/NET0131  , \g3263_reg/NET0131  , \g3288_reg/NET0131  , \g329_reg/NET0131  , \g3303_reg/NET0131  , \g3329_reg/NET0131  , \g3333_reg/NET0131  , \g3338_reg/NET0131  , \g333_reg/NET0131  , \g3343_reg/NET0131  , \g3347_reg/NET0131  , \g3352_reg/NET0131  , \g336_reg/NET0131  , \g341_reg/NET0131  , \g3457_reg/NET0131  , \g3466_reg/NET0131  , \g3470_reg/NET0131  , \g3476_reg/NET0131  , \g347_reg/NET0131  , \g3480_reg/NET0131  , \g3484_reg/NET0131  , \g3490_reg/NET0131  , \g3494_reg/NET0131  , \g34_reg/NET0131  , \g351_reg/NET0131  , \g355_reg/NET0131  , \g358_reg/NET0131  , \g35_pad  , \g3639_reg/NET0131  , \g3684_reg/NET0131  , \g3703_reg/NET0131  , \g370_reg/NET0131  , \g376_reg/NET0131  , \g37_reg/NET0131  , \g3808_reg/NET0131  , \g3817_reg/NET0131  , \g3821_reg/NET0131  , \g3827_reg/NET0131  , \g3831_reg/NET0131  , \g3835_reg/NET0131  , \g3841_reg/NET0131  , \g3845_reg/NET0131  , \g385_reg/NET0131  , \g392_reg/NET0131  , \g3990_reg/NET0131  , \g401_reg/NET0131  , \g4035_reg/NET0131  , \g4054_reg/NET0131  , \g4057_reg/NET0131  , \g405_reg/NET0131  , \g4064_reg/NET0131  , \g4072_reg/NET0131  , \g4076_reg/NET0131  , \g4082_reg/NET0131  , \g4087_reg/NET0131  , \g4093_reg/NET0131  , \g4098_reg/NET0131  , \g4104_reg/NET0131  , \g4108_reg/NET0131  , \g4112_reg/NET0131  , \g4116_reg/NET0131  , \g4119_reg/NET0131  , \g411_reg/NET0131  , \g4122_reg/NET0131  , \g4141_reg/NET0131  , \g4145_reg/NET0131  , \g4146_reg/NET0131  , \g4153_reg/NET0131  , \g4157_reg/NET0131  , \g4164_reg/NET0131  , \g4172_reg/NET0131  , \g4176_reg/NET0131  , \g417_reg/NET0131  , \g4180_reg/NET0131  , \g4235_reg/NET0131  , \g4239_reg/NET0131  , \g4242_reg/NET0131  , \g4245_reg/NET0131  , \g424_reg/NET0131  , \g4253_reg/NET0131  , \g4258_reg/NET0131  , \g4264_reg/NET0131  , \g4269_reg/NET0131  , \g4273_reg/NET0131  , \g4281_reg/NET0131  , \g4284_reg/NET0131  , \g4291_reg/NET0131  , \g4297_reg/NET0131  , \g4300_reg/NET0131  , \g4308_reg/NET0131  , \g4311_reg/NET0131  , \g4322_reg/NET0131  , \g4332_reg/NET0131  , \g433_reg/NET0131  , \g4340_reg/NET0131  , \g4349_reg/NET0131  , \g4358_reg/NET0131  , \g4366_reg/NET0131  , \g4369_reg/NET0131  , \g4372_reg/NET0131  , \g4375_reg/NET0131  , \g437_reg/NET0131  , \g4382_reg/NET0131  , \g4388_reg/NET0131  , \g4392_reg/NET0131  , \g4401_reg/NET0131  , \g4405_reg/NET0131  , \g4411_reg/NET0131  , \g4417_reg/NET0131  , \g441_reg/NET0131  , \g4420_reg/NET0131  , \g4423_reg/NET0131  , \g4427_reg/NET0131  , \g4430_reg/NET0131  , \g4434_reg/NET0131  , \g4438_reg/NET0131  , \g4443_reg/NET0131  , \g4452_reg/NET0131  , \g4455_reg/NET0131  , \g4459_reg/NET0131  , \g4462_reg/NET0131  , \g4467_reg/NET0131  , \g446_reg/NET0131  , \g4473_reg/NET0131  , \g4477_reg/NET0131  , \g4480_reg/NET0131  , \g4483_reg/NET0131  , \g4486_reg/NET0131  , \g4489_reg/NET0131  , \g4492_reg/NET0131  , \g4495_reg/NET0131  , \g4498_reg/NET0131  , \g4501_reg/NET0131  , \g4504_reg/NET0131  , \g4512_reg/NET0131  , \g4515_reg/NET0131  , \g4521_reg/NET0131  , \g4527_reg/NET0131  , \g452_reg/NET0131  , \g4531_reg/NET0131  , \g4534_reg/NET0131  , \g4540_reg/NET0131  , \g4543_reg/NET0131  , \g4546_reg/NET0131  , \g4549_reg/NET0131  , \g4552_reg/NET0131  , \g4555_reg/NET0131  , \g4558_reg/NET0131  , \g4561_reg/NET0131  , \g4564_reg/NET0131  , \g4567_reg/NET0131  , \g4572_reg/NET0131  , \g4575_reg/NET0131  , \g4581_reg/NET0131  , \g4584_reg/NET0131  , \g4593_reg/NET0131  , \g4601_reg/NET0131  , \g4608_reg/NET0131  , \g460_reg/NET0131  , \g4616_reg/NET0131  , \g4621_reg/NET0131  , \g4628_reg/NET0131  , \g4633_reg/NET0131  , \g4639_reg/NET0131  , \g4643_reg/NET0131  , \g4646_reg/NET0131  , \g4653_reg/NET0131  , \g4659_reg/NET0131  , \g4664_reg/NET0131  , \g4669_reg/NET0131  , \g4674_reg/NET0131  , \g4681_reg/NET0131  , \g4688_reg/NET0131  , \g4698_reg/NET0131  , \g4704_reg/NET0131  , \g4709_reg/NET0131  , \g4743_reg/NET0131  , \g4749_reg/NET0131  , \g4754_reg/NET0131  , \g475_reg/NET0131  , \g4760_reg/NET0131  , \g4765_reg/NET0131  , \g4771_reg/NET0131  , \g4776_reg/NET0131  , \g4785_reg/NET0131  , \g4793_reg/NET0131  , \g479_reg/NET0131  , \g4801_reg/NET0131  , \g482_reg/NET0131  , \g490_reg/NET0131  , \g496_reg/NET0131  , \g499_reg/NET0131  , \g5016_reg/NET0131  , \g5022_reg/NET0131  , \g5029_reg/NET0131  , \g5033_reg/NET0131  , \g5037_reg/NET0131  , \g5041_reg/NET0131  , \g5046_reg/NET0131  , \g504_reg/NET0131  , \g5052_reg/NET0131  , \g5057_reg/NET0131  , \g5069_reg/NET0131  , \g5073_reg/NET0131  , \g5077_reg/NET0131  , \g5080_reg/NET0131  , \g5084_reg/NET0131  , \g5092_reg/NET0131  , \g5097_reg/NET0131  , \g5101_reg/NET0131  , \g5112_reg/NET0131  , \g5115_reg/NET0131  , \g5124_reg/NET0131  , \g5128_reg/NET0131  , \g5134_reg/NET0131  , \g5138_reg/NET0131  , \g513_reg/NET0131  , \g5142_reg/NET0131  , \g5148_reg/NET0131  , \g5152_reg/NET0131  , \g518_reg/NET0131  , \g528_reg/NET0131  , \g5297_reg/NET0131  , \g534_reg/NET0131  , \g5357_reg/NET0131  , \g538_reg/NET0131  , \g542_reg/NET0131  , \g546_reg/NET0131  , \g550_reg/NET0131  , \g554_reg/NET0131  , \g645_reg/NET0131  , \g650_reg/NET0131  , \g655_reg/NET0131  , \g661_reg/NET0131  , \g667_reg/NET0131  , \g671_reg/NET0131  , \g676_reg/NET0131  , \g681_reg/NET0131  , \g686_reg/NET0131  , \g691_reg/NET0131  , \g699_reg/NET0131  , \g703_reg/NET0131  , \g714_reg/NET0131  , \g718_reg/NET0131  , \g723_reg/NET0131  , \g7243_pad  , \g7245_pad  , \g7257_pad  , \g7260_pad  , \g728_reg/NET0131  , \g732_reg/NET0131  , \g736_reg/NET0131  , \g739_reg/NET0131  , \g744_reg/NET0131  , \g749_reg/NET0131  , \g753_reg/NET0131  , \g7540_pad  , \g758_reg/NET0131  , \g763_reg/NET0131  , \g767_reg/NET0131  , \g772_reg/NET0131  , \g776_reg/NET0131  , \g781_reg/NET0131  , \g785_reg/NET0131  , \g790_reg/NET0131  , \g7916_pad  , \g7946_pad  , \g794_reg/NET0131  , \g802_reg/NET0131  , \g807_reg/NET0131  , \g812_reg/NET0131  , \g817_reg/NET0131  , \g822_reg/NET0131  , \g827_reg/NET0131  , \g8291_pad  , \g832_reg/NET0131  , \g8358_pad  , \g837_reg/NET0131  , \g8416_pad  , \g843_reg/NET0131  , \g8475_pad  , \g847_reg/NET0131  , \g854_reg/NET0131  , \g862_reg/NET0131  , \g8719_pad  , \g872_reg/NET0131  , \g8783_pad  , \g8784_pad  , \g8785_pad  , \g8786_pad  , \g8787_pad  , \g8788_pad  , \g8789_pad  , \g8839_pad  , \g8870_pad  , \g890_reg/NET0131  , \g8915_pad  , \g8916_pad  , \g8917_pad  , \g8918_pad  , \g8919_pad  , \g8920_pad  , \g896_reg/NET0131  , \g9019_pad  , \g9251_pad  , \g956_reg/NET0131  , \g962_reg/NET0131  , \g969_reg/NET0131  , \g976_reg/NET0131  , \g979_reg/NET0131  , \g990_reg/NET0131  , \g996_reg/NET0131  , \g136_reg/P0001  , \g21727_pad  , \g23190_pad  , \g26875_pad  , \g26876_pad  , \g26877_pad  , \g28041_pad  , \g28042_pad  , \g30327_pad  , \g30330_pad  , \g30331_pad  , \g31793_pad  , \g31860_pad  , \g31862_pad  , \g31863_pad  , \g32185_pad  , \g33079_pad  , \g33435_pad  , \g33959_pad  , \g34435_pad  , \g34788_pad  , \g34956_pad  , \g34_reg/P0001  , \g35_syn_2  , \g37/_0_  , \g41/_0_  , \g60853/_3_  , \g60856/_3_  , \g60879/_3_  , \g60882/_0_  , \g60888/_0_  , \g60891/_0_  , \g60896/_0_  , \g60899/_0_  , \g60900/_3_  , \g60909/_3_  , \g60911/_0_  , \g60915/_0_  , \g60918/_0_  , \g60919/_0_  , \g60928/_0_  , \g60929/_0_  , \g60936/_0_  , \g60937/_0_  , \g60939/_0_  , \g60940/_0_  , \g60941/_0_  , \g60942/_0_  , \g60943/_0_  , \g60944/_0_  , \g60952/_0_  , \g60954/_0_  , \g60958/_0_  , \g60962/_3_  , \g60972/_0_  , \g60980/_0_  , \g60984/_0_  , \g60986/_0_  , \g60989/_0_  , \g60991/_3_  , \g61006/_0_  , \g61008/_0_  , \g61013/_0_  , \g61014/_0_  , \g61015/_0_  , \g61016/_0_  , \g61017/_0_  , \g61026/_3_  , \g61027/_3_  , \g61030/_0_  , \g61031/_0_  , \g61037/_0_  , \g61038/_0_  , \g61042/_0_  , \g61044/_0_  , \g61045/_0_  , \g61046/_0_  , \g61050/_0_  , \g61051/_0_  , \g61052/_0_  , \g61078/_0_  , \g61131/_0_  , \g61137/_3_  , \g61142/_3_  , \g61143/_3_  , \g61151/_0_  , \g61152/_0_  , \g61161/_0_  , \g61168/_3_  , \g61169/_3_  , \g61170/_0_  , \g61171/_3_  , \g61172/_0_  , \g61173/_0_  , \g61174/_0_  , \g61175/_0_  , \g61176/_0_  , \g61177/_3_  , \g61178/_0_  , \g61179/_0_  , \g61180/_0_  , \g61181/_0_  , \g61182/_3_  , \g61183/_0_  , \g61184/_3_  , \g61185/_0_  , \g61186/_0_  , \g61187/_0_  , \g61188/_0_  , \g61189/_0_  , \g61190/_3_  , \g61191/_0_  , \g61192/_0_  , \g61193/_0_  , \g61194/_0_  , \g61221/_0_  , \g61222/_0_  , \g61223/_3_  , \g61224/_3_  , \g61261/_0_  , \g61295/_3_  , \g61308/_0_  , \g61316/_0_  , \g61327/_0_  , \g61329/_0_  , \g61330/_0_  , \g61331/_0_  , \g61332/_3_  , \g61333/_0_  , \g61334/_0_  , \g61335/_0_  , \g61336/_0_  , \g61337/_0_  , \g61338/_3_  , \g61339/_0_  , \g61340/_0_  , \g61341/_0_  , \g61342/_0_  , \g61343/_0_  , \g61344/_3_  , \g61345/_0_  , \g61346/_0_  , \g61347/_0_  , \g61348/_0_  , \g61349/_0_  , \g61350/_3_  , \g61351/_0_  , \g61352/_0_  , \g61353/_0_  , \g61354/_0_  , \g61367/_0_  , \g61372/_0_  , \g61373/_0_  , \g61375/_0_  , \g61382/_0_  , \g61385/_3_  , \g61386/_0_  , \g61399/_0_  , \g61400/_0_  , \g61402/_0_  , \g61405/_0_  , \g61435/_3_  , \g61449/_0_  , \g61468/_0_  , \g61475/_0_  , \g61480/_0_  , \g61482/_0_  , \g61483/_0_  , \g61484/_0_  , \g61486/_3_  , \g61494/_0_  , \g61496/_0_  , \g61497/_0_  , \g61514/_0_  , \g61517/_0_  , \g61519/_3_  , \g61520/_3_  , \g61527/_0_  , \g61541/_0_  , \g61544/_0_  , \g61550/_0_  , \g61551/_0_  , \g61554/_0_  , \g61556/_3_  , \g61567/_0_  , \g61571/_0_  , \g61574/_0_  , \g61587/_0_  , \g61592/_0_  , \g61632/_0_  , \g61634/_0_  , \g61635/_0_  , \g61639/_0_  , \g61644/_0_  , \g61652/_3_  , \g61709/_0_  , \g61714/_0_  , \g61720/_0_  , \g61721/_0_  , \g61723/_0_  , \g61725/_0_  , \g61726/_0_  , \g61734/_0_  , \g61739/_0_  , \g61744/_0_  , \g61746/_3_  , \g61747/_3_  , \g61748/_3_  , \g61750/u3_syn_7  , \g61802/_0_  , \g61804/_0_  , \g61808/_0_  , \g61811/_0_  , \g61816/_0_  , \g61818/_0_  , \g61820/_0_  , \g61823/_0_  , \g61824/_0_  , \g61841/_0_  , \g61842/_3_  , \g61844/_3_  , \g61845/_3_  , \g61846/_3_  , \g61847/u3_syn_7  , \g61848/_0_  , \g61849/_3_  , \g61850/_0_  , \g61851/u3_syn_7  , \g61852/_0_  , \g61853/_3_  , \g61854/_3_  , \g61855/_0_  , \g61856/u3_syn_7  , \g61857/_0_  , \g61858/_3_  , \g61859/_3_  , \g61860/u3_syn_7  , \g61861/_0_  , \g61862/_3_  , \g61863/_3_  , \g61864/u3_syn_7  , \g61865/_0_  , \g61866/_3_  , \g61867/_3_  , \g61868/u3_syn_7  , \g61869/_0_  , \g61870/_0_  , \g61871/_3_  , \g61872/_3_  , \g61873/u3_syn_7  , \g61874/_0_  , \g61875/_0_  , \g61877/_3_  , \g61878/_3_  , \g61879/u3_syn_7  , \g61880/_0_  , \g61881/_0_  , \g61882/_0_  , \g61883/_0_  , \g61884/_0_  , \g61914/_0_  , \g61915/_0_  , \g61917/_0_  , \g61918/_0_  , \g61922/_0_  , \g61923/_0_  , \g61924/_0_  , \g61932/_0_  , \g61936/_0_  , \g61945/_0_  , \g61947/_0_  , \g61959/_0_  , \g61960/_0_  , \g61962/_0_  , \g61973/_3_  , \g61974/u3_syn_7  , \g61975/_3_  , \g61976/u3_syn_7  , \g61977/_3_  , \g61978/_3_  , \g61979/u3_syn_7  , \g61980/_3_  , \g61981/_3_  , \g61982/_3_  , \g61983/u3_syn_7  , \g61984/_3_  , \g61985/_3_  , \g61986/u3_syn_7  , \g61987/_3_  , \g61988/_3_  , \g61989/u3_syn_7  , \g61990/_3_  , \g61991/_3_  , \g61992/u3_syn_7  , \g61993/_3_  , \g61994/u3_syn_7  , \g61995/_3_  , \g61996/_3_  , \g61997/_3_  , \g62022/_0_  , \g62028/_0_  , \g62029/_0_  , \g62031/_0_  , \g62033/_0_  , \g62038/_0_  , \g62042/_0_  , \g62046/_0_  , \g62048/_0_  , \g62049/_0_  , \g62051/_0_  , \g62053/_0_  , \g62085/_0_  , \g62101/_0_  , \g62102/_0_  , \g62103/_0_  , \g62105/_0_  , \g62108/_3_  , \g62112/_0_  , \g62137/_3_  , \g62207/_0_  , \g62239/_0_  , \g62240/_0_  , \g62267/_0_  , \g62273/_0_  , \g62284/_0_  , \g62291/_0_  , \g62293/_0_  , \g62298/_0_  , \g62303/_3_  , \g62322/_3_  , \g62323/_3_  , \g62324/_3_  , \g62325/_3_  , \g62583/_0_  , \g62598/_0_  , \g62609/_0_  , \g62636/_0_  , \g62646/_0_  , \g62649/_0_  , \g62658/_0_  , \g62663/_0_  , \g62664/_0_  , \g62667/_0_  , \g62676/_0_  , \g62677/_0_  , \g62678/_3_  , \g62679/_0_  , \g62687/u3_syn_7  , \g62688/u3_syn_7  , \g62689/_0_  , \g62690/_3_  , \g62691/_3_  , \g62693/_0_  , \g62694/_3_  , \g62695/_3_  , \g62696/_3_  , \g62697/_3_  , \g62698/_3_  , \g62699/_3_  , \g62700/_3_  , \g62701/_3_  , \g62702/_3_  , \g62703/_3_  , \g62704/u3_syn_7  , \g62705/_0_  , \g62706/_3_  , \g62707/_3_  , \g62708/u3_syn_7  , \g62709/_0_  , \g62710/_3_  , \g62711/_3_  , \g62712/u3_syn_7  , \g62713/_0_  , \g62714/_3_  , \g62715/_0_  , \g62716/u3_syn_7  , \g62717/_0_  , \g62718/_3_  , \g62719/_0_  , \g62720/u3_syn_7  , \g62721/_0_  , \g62722/_3_  , \g62723/_0_  , \g62724/u3_syn_7  , \g62725/_0_  , \g62726/_3_  , \g62728/_0_  , \g62790/_0_  , \g62791/_0_  , \g62793/_0_  , \g62794/_0_  , \g62795/_0_  , \g62796/_0_  , \g62797/_0_  , \g62807/_0_  , \g62823/_0_  , \g62824/_0_  , \g62833/_0_  , \g62846/_0_  , \g62859/_0_  , \g62860/_0_  , \g62897/_0_  , \g62898/_0_  , \g62922/_3_  , \g62923/_0_  , \g62927/_0_  , \g62938/_3_  , \g62939/_3_  , \g62940/_3_  , \g62941/u3_syn_7  , \g62942/_0_  , \g62943/_3_  , \g62987/_3_  , \g62991/_3_  , \g63015/u3_syn_7  , \g63016/_0_  , \g63017/_3_  , \g63018/_3_  , \g63019/_3_  , \g63020/_3_  , \g63021/_3_  , \g63022/_3_  , \g63025/_3_  , \g63026/_3_  , \g63027/_3_  , \g63029/_3_  , \g63030/_3_  , \g63031/_3_  , \g63033/_3_  , \g63034/_3_  , \g63043/_3_  , \g63044/_3_  , \g63051/_3_  , \g63057/_3_  , \g63068/_3_  , \g63070/_3_  , \g63073/_3_  , \g63081/_3_  , \g63082/_3_  , \g63083/u3_syn_7  , \g63084/_3_  , \g63085/_0_  , \g63086/_3_  , \g63107/_3_  , \g63108/u3_syn_7  , \g63109/u3_syn_7  , \g63110/_0_  , \g63111/_3_  , \g63132/_3_  , \g63133/_3_  , \g63134/_3_  , \g63135/_3_  , \g63136/_3_  , \g63137/_3_  , \g63138/_3_  , \g63139/u3_syn_7  , \g63140/_3_  , \g63141/_3_  , \g63142/_3_  , \g63143/_3_  , \g63144/_3_  , \g63145/_3_  , \g63146/u3_syn_7  , \g63198/_0_  , \g63205/_0_  , \g63208/_0_  , \g63212/_0_  , \g63215/_0_  , \g63219/_0_  , \g63244/_0_  , \g63246/_0_  , \g63254/_0_  , \g63255/_0_  , \g63272/_0_  , \g63276/_0_  , \g63278/_0_  , \g63279/_0_  , \g63280/_0_  , \g63327/_0_  , \g63345/_0_  , \g63346/_3_  , \g63347/_3_  , \g63354/_3_  , \g63358/_3_  , \g63359/u3_syn_7  , \g63361/_3_  , \g63365/_3_  , \g63366/_3_  , \g63367/_3_  , \g63368/_3_  , \g63370/_3_  , \g63479/_0_  , \g63484/_0_  , \g63499/_1_  , \g63520/_0_  , \g63523/_0_  , \g63526/_0_  , \g63538/_0_  , \g63539/_0_  , \g63541/_0_  , \g63555/_0_  , \g63642/_0_  , \g63645/_0_  , \g63648/_3_  , \g63777/_3_  , \g63778/_3_  , \g63781/_0_  , \g63786/u3_syn_7  , \g63787/_3_  , \g63788/_3_  , \g63790/_3_  , \g63791/_3_  , \g63792/u3_syn_7  , \g63794/_0_  , \g63795/_0_  , \g63796/_0_  , \g63798/_3_  , \g63800/_3_  , \g63804/_3_  , \g63805/_3_  , \g63806/_3_  , \g63807/_3_  , \g63808/_3_  , \g63809/_3_  , \g63870/_0_  , \g63883/_0_  , \g63934/_0_  , \g63936/_0_  , \g63938/_0_  , \g63939/_0_  , \g63966/_0_  , \g63970/_0_  , \g63999/_0_  , \g64039/_0_  , \g64040/_0_  , \g64043/_0_  , \g64062/_3_  , \g64078/_0_  , \g64091/_0_  , \g64095/_3_  , \g64096/_3_  , \g64097/u3_syn_7  , \g64098/u3_syn_7  , \g64099/u3_syn_7  , \g64100/u3_syn_7  , \g64134/_0_  , \g64135/_0_  , \g64153/_0_  , \g64155/_0_  , \g64179/_0_  , \g64229/_0_  , \g64235/_0_  , \g64236/_0_  , \g64280/_0_  , \g64315/_0_  , \g64365/_0_  , \g64426/_3_  , \g64438/_3_  , \g64442/u3_syn_7  , \g64445/_3_  , \g64447/_3_  , \g64449/_3_  , \g64451/_3_  , \g64453/_3_  , \g64454/_3_  , \g64460/_3_  , \g64461/_3_  , \g64510/_0_  , \g64527/_0_  , \g64528/_0_  , \g64544/_0_  , \g64549/_0_  , \g64566/_0_  , \g64576/_0_  , \g64602/_0_  , \g64691/_0_  , \g64697/_0_  , \g64707/_3_  , \g64778/_3_  , \g64790/_3_  , \g64791/_3_  , \g64792/_3_  , \g64793/_3_  , \g64794/_3_  , \g64795/_3_  , \g64796/_3_  , \g64797/_3_  , \g64877/_0_  , \g64912/_0_  , \g64973/_0_  , \g65047/_3_  , \g65081/_3_  , \g65088/_3_  , \g65097/_3_  , \g65100/_3_  , \g65101/_3_  , \g65104/_3_  , \g65105/_3_  , \g65107/_3_  , \g65110/_3_  , \g65111/_3_  , \g65113/_3_  , \g65114/_3_  , \g65266/_0_  , \g65267/_0_  , \g65294/_1_  , \g65328/_1_  , \g65495/_0_  , \g65499/_0_  , \g65503/_0_  , \g65529/_0_  , \g65530/_3_  , \g65531/_3_  , \g65532/_3_  , \g65533/_3_  , \g65624/_0_  , \g65625/_1_  , \g65641/_0_  , \g65701/_0_  , \g65704/_0_  , \g65853/_0_  , \g65891/_0_  , \g65901/_0_  , \g65986/_0_  , \g66029/_0_  , \g66066/_0_  , \g66067/_0_  , \g66068/_0_  , \g66154/_3_  , \g66362/_0_  , \g66369/_0_  , \g66398/_0_  , \g66409/_0_  , \g66419/_0_  , \g66439/_0_  , \g66443/_0_  , \g66464/_0_  , \g66471/_0_  , \g66512/_0_  , \g66528/_0_  , \g66541/_0_  , \g66558/_0_  , \g66644/_0_  , \g66684/_0_  , \g66697/_0_  , \g66698/_0_  , \g66701/_0_  , \g66714/_0_  , \g66715/_0_  , \g66745/_0_  , \g66750/_0_  , \g66751/_0_  , \g66810/_0_  , \g66844/_0_  , \g66853/_0_  , \g66897/_0_  , \g66905/_0_  , \g69743/_0_  , \g69750/_0_  , \g69773/_1_  , \g69792/_1_  , \g69858/_0_  , \g69938/_0_  , \g69949/_0_  , \g70167/_0_  , \g71190/_0_  , \g71198/_0_  , \g71284/_0_  , \g72369/_1_  , \g72467/_0_  , \g72476/_0_  , \g72477/_1_  , \g72648/_0_  , \g72741/_0_  , \g72772/_0_  , \g8132_pad  );
  input \g1002_reg/NET0131  ;
  input \g1008_reg/NET0131  ;
  input \g10122_pad  ;
  input \g1018_reg/NET0131  ;
  input \g1024_reg/NET0131  ;
  input \g10306_pad  ;
  input \g1030_reg/NET0131  ;
  input \g1036_reg/NET0131  ;
  input \g1041_reg/NET0131  ;
  input \g1046_reg/NET0131  ;
  input \g10500_pad  ;
  input \g10527_pad  ;
  input \g1052_reg/NET0131  ;
  input \g1061_reg/NET0131  ;
  input \g1070_reg/NET0131  ;
  input \g1087_reg/NET0131  ;
  input \g1094_reg/NET0131  ;
  input \g1099_reg/NET0131  ;
  input \g1105_reg/NET0131  ;
  input \g1111_reg/NET0131  ;
  input \g1124_reg/NET0131  ;
  input \g1129_reg/NET0131  ;
  input \g1135_reg/NET0131  ;
  input \g1141_reg/NET0131  ;
  input \g11447_pad  ;
  input \g1146_reg/NET0131  ;
  input \g1152_reg/NET0131  ;
  input \g1171_reg/NET0131  ;
  input \g11770_pad  ;
  input \g1178_reg/NET0131  ;
  input \g1183_reg/NET0131  ;
  input \g1189_reg/NET0131  ;
  input \g1193_reg/NET0131  ;
  input \g1199_reg/NET0131  ;
  input \g1205_reg/NET0131  ;
  input \g1211_reg/NET0131  ;
  input \g1216_reg/NET0131  ;
  input \g12184_pad  ;
  input \g1221_reg/NET0131  ;
  input \g1236_reg/NET0131  ;
  input \g1242_reg/NET0131  ;
  input \g1246_reg/NET0131  ;
  input \g12919_pad  ;
  input \g12923_pad  ;
  input \g1300_reg/NET0131  ;
  input \g13039_pad  ;
  input \g1306_reg/NET0131  ;
  input \g1312_reg/NET0131  ;
  input \g1319_reg/NET0131  ;
  input \g1322_reg/NET0131  ;
  input \g13259_pad  ;
  input \g13272_pad  ;
  input \g1333_reg/NET0131  ;
  input \g1339_reg/NET0131  ;
  input \g1345_reg/NET0131  ;
  input \g1351_reg/NET0131  ;
  input \g1361_reg/NET0131  ;
  input \g1367_reg/NET0131  ;
  input \g1373_reg/NET0131  ;
  input \g1379_reg/NET0131  ;
  input \g1384_reg/NET0131  ;
  input \g13865_pad  ;
  input \g13895_pad  ;
  input \g1389_reg/NET0131  ;
  input \g1395_reg/NET0131  ;
  input \g1404_reg/NET0131  ;
  input \g14096_pad  ;
  input \g14125_pad  ;
  input \g1413_reg/NET0131  ;
  input \g14147_pad  ;
  input \g14167_pad  ;
  input \g14189_pad  ;
  input \g14201_pad  ;
  input \g14217_pad  ;
  input \g142_reg/NET0131  ;
  input \g1430_reg/NET0131  ;
  input \g1437_reg/NET0131  ;
  input \g1442_reg/NET0131  ;
  input \g1448_reg/NET0131  ;
  input \g1454_reg/NET0131  ;
  input \g1467_reg/NET0131  ;
  input \g146_reg/NET0131  ;
  input \g1472_reg/NET0131  ;
  input \g1478_reg/NET0131  ;
  input \g1484_reg/NET0131  ;
  input \g1489_reg/NET0131  ;
  input \g1495_reg/NET0131  ;
  input \g150_reg/NET0131  ;
  input \g1514_reg/NET0131  ;
  input \g1521_reg/NET0131  ;
  input \g1526_reg/NET0131  ;
  input \g1532_reg/NET0131  ;
  input \g1536_reg/NET0131  ;
  input \g153_reg/NET0131  ;
  input \g1542_reg/NET0131  ;
  input \g1548_reg/NET0131  ;
  input \g1554_reg/NET0131  ;
  input \g1559_reg/NET0131  ;
  input \g1564_reg/NET0131  ;
  input \g1579_reg/NET0131  ;
  input \g157_reg/NET0131  ;
  input \g1585_reg/NET0131  ;
  input \g1589_reg/NET0131  ;
  input \g1592_reg/NET0131  ;
  input \g1600_reg/NET0131  ;
  input \g1604_reg/NET0131  ;
  input \g1608_reg/NET0131  ;
  input \g160_reg/NET0131  ;
  input \g1612_reg/NET0131  ;
  input \g1616_reg/NET0131  ;
  input \g1620_reg/NET0131  ;
  input \g1624_reg/NET0131  ;
  input \g1632_reg/NET0131  ;
  input \g1636_reg/NET0131  ;
  input \g1644_reg/NET0131  ;
  input \g1648_reg/NET0131  ;
  input \g164_reg/NET0131  ;
  input \g1657_reg/NET0131  ;
  input \g16603_pad  ;
  input \g16624_pad  ;
  input \g1664_reg/NET0131  ;
  input \g16686_pad  ;
  input \g1668_reg/NET0131  ;
  input \g16718_pad  ;
  input \g1677_reg/NET0131  ;
  input \g1682_reg/NET0131  ;
  input \g16874_pad  ;
  input \g1687_reg/NET0131  ;
  input \g168_reg/NET0131  ;
  input \g1691_reg/NET0131  ;
  input \g1696_reg/NET0131  ;
  input \g1700_reg/NET0131  ;
  input \g1706_reg/NET0131  ;
  input \g1710_reg/NET0131  ;
  input \g1714_reg/NET0131  ;
  input \g1720_reg/NET0131  ;
  input \g1724_reg/NET0131  ;
  input \g1728_reg/NET0131  ;
  input \g17291_pad  ;
  input \g17316_pad  ;
  input \g17320_pad  ;
  input \g1736_reg/NET0131  ;
  input \g17400_pad  ;
  input \g17404_pad  ;
  input \g1740_reg/NET0131  ;
  input \g17423_pad  ;
  input \g1744_reg/NET0131  ;
  input \g1748_reg/NET0131  ;
  input \g174_reg/NET0131  ;
  input \g1752_reg/NET0131  ;
  input \g1756_reg/NET0131  ;
  input \g1760_reg/NET0131  ;
  input \g1768_reg/NET0131  ;
  input \g1772_reg/NET0131  ;
  input \g1779_reg/NET0131  ;
  input \g1783_reg/NET0131  ;
  input \g1792_reg/NET0131  ;
  input \g1798_reg/NET0131  ;
  input \g1802_reg/NET0131  ;
  input \g18094_pad  ;
  input \g18095_pad  ;
  input \g18096_pad  ;
  input \g18098_pad  ;
  input \g18099_pad  ;
  input \g1811_reg/NET0131  ;
  input \g1816_reg/NET0131  ;
  input \g1821_reg/NET0131  ;
  input \g1825_reg/NET0131  ;
  input \g182_reg/NET0131  ;
  input \g1830_reg/NET0131  ;
  input \g1834_reg/NET0131  ;
  input \g1840_reg/NET0131  ;
  input \g1844_reg/NET0131  ;
  input \g1848_reg/NET0131  ;
  input \g1854_reg/NET0131  ;
  input \g1858_reg/NET0131  ;
  input \g1862_reg/NET0131  ;
  input \g1870_reg/NET0131  ;
  input \g1874_reg/NET0131  ;
  input \g1878_reg/NET0131  ;
  input \g1882_reg/NET0131  ;
  input \g1886_reg/NET0131  ;
  input \g1890_reg/NET0131  ;
  input \g1894_reg/NET0131  ;
  input \g1902_reg/NET0131  ;
  input \g1906_reg/NET0131  ;
  input \g1913_reg/NET0131  ;
  input \g1917_reg/NET0131  ;
  input \g191_reg/NET0131  ;
  input \g1926_reg/NET0131  ;
  input \g1932_reg/NET0131  ;
  input \g19334_pad  ;
  input \g19357_pad  ;
  input \g1936_reg/NET0131  ;
  input \g1945_reg/NET0131  ;
  input \g1950_reg/NET0131  ;
  input \g1955_reg/NET0131  ;
  input \g1959_reg/NET0131  ;
  input \g1964_reg/NET0131  ;
  input \g1968_reg/NET0131  ;
  input \g1974_reg/NET0131  ;
  input \g1978_reg/NET0131  ;
  input \g1982_reg/NET0131  ;
  input \g1988_reg/NET0131  ;
  input \g1992_reg/NET0131  ;
  input \g1996_reg/NET0131  ;
  input \g2004_reg/NET0131  ;
  input \g2008_reg/NET0131  ;
  input \g2012_reg/NET0131  ;
  input \g2016_reg/NET0131  ;
  input \g2020_reg/NET0131  ;
  input \g2024_reg/NET0131  ;
  input \g2028_reg/NET0131  ;
  input \g2036_reg/NET0131  ;
  input \g203_reg/NET0131  ;
  input \g2040_reg/NET0131  ;
  input \g2047_reg/NET0131  ;
  input \g2051_reg/NET0131  ;
  input \g2060_reg/NET0131  ;
  input \g2066_reg/NET0131  ;
  input \g2070_reg/NET0131  ;
  input \g2079_reg/NET0131  ;
  input \g2084_reg/NET0131  ;
  input \g2089_reg/NET0131  ;
  input \g2093_reg/NET0131  ;
  input \g2098_reg/NET0131  ;
  input \g209_reg/NET0131  ;
  input \g2102_reg/NET0131  ;
  input \g2108_reg/NET0131  ;
  input \g2112_reg/NET0131  ;
  input \g2116_reg/NET0131  ;
  input \g2122_reg/NET0131  ;
  input \g2126_reg/NET0131  ;
  input \g2153_reg/NET0131  ;
  input \g2161_reg/NET0131  ;
  input \g2165_reg/NET0131  ;
  input \g2169_reg/NET0131  ;
  input \g2173_reg/NET0131  ;
  input \g2177_reg/NET0131  ;
  input \g2181_reg/NET0131  ;
  input \g2185_reg/NET0131  ;
  input \g218_reg/NET0131  ;
  input \g2193_reg/NET0131  ;
  input \g2197_reg/NET0131  ;
  input \g2204_reg/NET0131  ;
  input \g2208_reg/NET0131  ;
  input \g2217_reg/NET0131  ;
  input \g2223_reg/NET0131  ;
  input \g2227_reg/NET0131  ;
  input \g222_reg/NET0131  ;
  input \g2236_reg/NET0131  ;
  input \g2241_reg/NET0131  ;
  input \g2246_reg/NET0131  ;
  input \g2250_reg/NET0131  ;
  input \g2255_reg/NET0131  ;
  input \g2259_reg/NET0131  ;
  input \g225_reg/NET0131  ;
  input \g2265_reg/NET0131  ;
  input \g2269_reg/NET0131  ;
  input \g2273_reg/NET0131  ;
  input \g2279_reg/NET0131  ;
  input \g2283_reg/NET0131  ;
  input \g2287_reg/NET0131  ;
  input \g2295_reg/NET0131  ;
  input \g2299_reg/NET0131  ;
  input \g2303_reg/NET0131  ;
  input \g2307_reg/NET0131  ;
  input \g2311_reg/NET0131  ;
  input \g2315_reg/NET0131  ;
  input \g2319_reg/NET0131  ;
  input \g2327_reg/NET0131  ;
  input \g232_reg/NET0131  ;
  input \g2331_reg/NET0131  ;
  input \g2338_reg/NET0131  ;
  input \g2342_reg/NET0131  ;
  input \g2351_reg/NET0131  ;
  input \g2357_reg/NET0131  ;
  input \g2361_reg/NET0131  ;
  input \g2370_reg/NET0131  ;
  input \g2375_reg/NET0131  ;
  input \g2380_reg/NET0131  ;
  input \g2384_reg/NET0131  ;
  input \g2389_reg/NET0131  ;
  input \g2393_reg/NET0131  ;
  input \g2399_reg/NET0131  ;
  input \g239_reg/NET0131  ;
  input \g2403_reg/NET0131  ;
  input \g2407_reg/NET0131  ;
  input \g2413_reg/NET0131  ;
  input \g2417_reg/NET0131  ;
  input \g2421_reg/NET0131  ;
  input \g2429_reg/NET0131  ;
  input \g2433_reg/NET0131  ;
  input \g2437_reg/NET0131  ;
  input \g2441_reg/NET0131  ;
  input \g2445_reg/NET0131  ;
  input \g2449_reg/NET0131  ;
  input \g2453_reg/NET0131  ;
  input \g2461_reg/NET0131  ;
  input \g2465_reg/NET0131  ;
  input \g246_reg/NET0131  ;
  input \g2472_reg/NET0131  ;
  input \g2476_reg/NET0131  ;
  input \g2485_reg/NET0131  ;
  input \g2491_reg/NET0131  ;
  input \g2495_reg/NET0131  ;
  input \g2504_reg/NET0131  ;
  input \g2509_reg/NET0131  ;
  input \g2514_reg/NET0131  ;
  input \g2518_reg/NET0131  ;
  input \g2523_reg/NET0131  ;
  input \g2527_reg/NET0131  ;
  input \g2533_reg/NET0131  ;
  input \g2537_reg/NET0131  ;
  input \g2541_reg/NET0131  ;
  input \g2547_reg/NET0131  ;
  input \g2551_reg/NET0131  ;
  input \g2555_reg/NET0131  ;
  input \g255_reg/NET0131  ;
  input \g2563_reg/NET0131  ;
  input \g2567_reg/NET0131  ;
  input \g2571_reg/NET0131  ;
  input \g2575_reg/NET0131  ;
  input \g2579_reg/NET0131  ;
  input \g2583_reg/NET0131  ;
  input \g2587_reg/NET0131  ;
  input \g2595_reg/NET0131  ;
  input \g2599_reg/NET0131  ;
  input \g2606_reg/NET0131  ;
  input \g2610_reg/NET0131  ;
  input \g2619_reg/NET0131  ;
  input \g2625_reg/NET0131  ;
  input \g2629_reg/NET0131  ;
  input \g262_reg/NET0131  ;
  input \g2638_reg/NET0131  ;
  input \g2643_reg/NET0131  ;
  input \g2648_reg/NET0131  ;
  input \g2652_reg/NET0131  ;
  input \g2657_reg/NET0131  ;
  input \g2661_reg/NET0131  ;
  input \g2667_reg/NET0131  ;
  input \g2671_reg/NET0131  ;
  input \g2675_reg/NET0131  ;
  input \g2681_reg/NET0131  ;
  input \g2685_reg/NET0131  ;
  input \g269_reg/NET0131  ;
  input \g2715_reg/NET0131  ;
  input \g2719_reg/NET0131  ;
  input \g2724_reg/NET0131  ;
  input \g2729_reg/NET0131  ;
  input \g2735_reg/NET0131  ;
  input \g2741_reg/NET0131  ;
  input \g2748_reg/NET0131  ;
  input \g2756_reg/NET0131  ;
  input \g2759_reg/NET0131  ;
  input \g2763_reg/NET0131  ;
  input \g2767_reg/NET0131  ;
  input \g2771_reg/NET0131  ;
  input \g2775_reg/NET0131  ;
  input \g2779_reg/NET0131  ;
  input \g2783_reg/NET0131  ;
  input \g2787_reg/NET0131  ;
  input \g278_reg/NET0131  ;
  input \g2791_reg/NET0131  ;
  input \g2795_reg/NET0131  ;
  input \g2799_reg/NET0131  ;
  input \g2803_reg/NET0131  ;
  input \g2807_reg/NET0131  ;
  input \g2811_reg/NET0131  ;
  input \g2815_reg/NET0131  ;
  input \g2819_reg/NET0131  ;
  input \g2823_reg/NET0131  ;
  input \g2827_reg/NET0131  ;
  input \g2831_reg/NET0131  ;
  input \g2834_reg/NET0131  ;
  input \g283_reg/NET0131  ;
  input \g2848_reg/NET0131  ;
  input \g2856_reg/NET0131  ;
  input \g2864_reg/NET0131  ;
  input \g2873_reg/NET0131  ;
  input \g2878_reg/NET0131  ;
  input \g287_reg/NET0131  ;
  input \g2882_reg/NET0131  ;
  input \g2886_reg/NET0131  ;
  input \g2898_reg/NET0131  ;
  input \g2902_reg/NET0131  ;
  input \g2907_reg/NET0131  ;
  input \g2912_reg/NET0131  ;
  input \g2917_reg/NET0131  ;
  input \g291_reg/NET0131  ;
  input \g29211_pad  ;
  input \g29212_pad  ;
  input \g29213_pad  ;
  input \g29214_pad  ;
  input \g29215_pad  ;
  input \g29216_pad  ;
  input \g29218_pad  ;
  input \g29219_pad  ;
  input \g29220_pad  ;
  input \g29221_pad  ;
  input \g2922_reg/NET0131  ;
  input \g2927_reg/NET0131  ;
  input \g2932_reg/NET0131  ;
  input \g2936_reg/NET0131  ;
  input \g2941_reg/NET0131  ;
  input \g2946_reg/NET0131  ;
  input \g294_reg/NET0131  ;
  input \g2950_reg/NET0131  ;
  input \g2955_reg/NET0131  ;
  input \g2960_reg/NET0131  ;
  input \g2965_reg/NET0131  ;
  input \g2970_reg/NET0131  ;
  input \g2975_reg/NET0131  ;
  input \g2980_reg/NET0131  ;
  input \g2984_reg/NET0131  ;
  input \g2988_reg/NET0131  ;
  input \g298_reg/NET0131  ;
  input \g2999_reg/NET0131  ;
  input \g3003_reg/NET0131  ;
  input \g301_reg/NET0131  ;
  input \g3050_reg/NET0131  ;
  input \g305_reg/NET0131  ;
  input \g3096_reg/NET0131  ;
  input \g3100_reg/NET0131  ;
  input \g3106_reg/NET0131  ;
  input \g3111_reg/NET0131  ;
  input \g3115_reg/NET0131  ;
  input \g3119_reg/NET0131  ;
  input \g311_reg/NET0131  ;
  input \g3125_reg/NET0131  ;
  input \g3129_reg/NET0131  ;
  input \g3133_reg/NET0131  ;
  input \g3139_reg/NET0131  ;
  input \g3143_reg/NET0131  ;
  input \g3147_reg/NET0131  ;
  input \g3155_reg/NET0131  ;
  input \g3161_reg/NET0131  ;
  input \g3167_reg/NET0131  ;
  input \g316_reg/NET0131  ;
  input \g3171_reg/NET0131  ;
  input \g3179_reg/NET0131  ;
  input \g3187_reg/NET0131  ;
  input \g3191_reg/NET0131  ;
  input \g3195_reg/NET0131  ;
  input \g3199_reg/NET0131  ;
  input \g319_reg/NET0131  ;
  input \g3203_reg/NET0131  ;
  input \g3207_reg/NET0131  ;
  input \g3211_reg/NET0131  ;
  input \g3215_reg/NET0131  ;
  input \g3219_reg/NET0131  ;
  input \g3223_reg/NET0131  ;
  input \g3227_reg/NET0131  ;
  input \g3231_reg/NET0131  ;
  input \g3235_reg/NET0131  ;
  input \g3239_reg/NET0131  ;
  input \g3243_reg/NET0131  ;
  input \g3247_reg/NET0131  ;
  input \g324_reg/NET0131  ;
  input \g3251_reg/NET0131  ;
  input \g3255_reg/NET0131  ;
  input \g3259_reg/NET0131  ;
  input \g3263_reg/NET0131  ;
  input \g3288_reg/NET0131  ;
  input \g329_reg/NET0131  ;
  input \g3303_reg/NET0131  ;
  input \g3329_reg/NET0131  ;
  input \g3333_reg/NET0131  ;
  input \g3338_reg/NET0131  ;
  input \g333_reg/NET0131  ;
  input \g3343_reg/NET0131  ;
  input \g3347_reg/NET0131  ;
  input \g3352_reg/NET0131  ;
  input \g336_reg/NET0131  ;
  input \g341_reg/NET0131  ;
  input \g3457_reg/NET0131  ;
  input \g3466_reg/NET0131  ;
  input \g3470_reg/NET0131  ;
  input \g3476_reg/NET0131  ;
  input \g347_reg/NET0131  ;
  input \g3480_reg/NET0131  ;
  input \g3484_reg/NET0131  ;
  input \g3490_reg/NET0131  ;
  input \g3494_reg/NET0131  ;
  input \g34_reg/NET0131  ;
  input \g351_reg/NET0131  ;
  input \g355_reg/NET0131  ;
  input \g358_reg/NET0131  ;
  input \g35_pad  ;
  input \g3639_reg/NET0131  ;
  input \g3684_reg/NET0131  ;
  input \g3703_reg/NET0131  ;
  input \g370_reg/NET0131  ;
  input \g376_reg/NET0131  ;
  input \g37_reg/NET0131  ;
  input \g3808_reg/NET0131  ;
  input \g3817_reg/NET0131  ;
  input \g3821_reg/NET0131  ;
  input \g3827_reg/NET0131  ;
  input \g3831_reg/NET0131  ;
  input \g3835_reg/NET0131  ;
  input \g3841_reg/NET0131  ;
  input \g3845_reg/NET0131  ;
  input \g385_reg/NET0131  ;
  input \g392_reg/NET0131  ;
  input \g3990_reg/NET0131  ;
  input \g401_reg/NET0131  ;
  input \g4035_reg/NET0131  ;
  input \g4054_reg/NET0131  ;
  input \g4057_reg/NET0131  ;
  input \g405_reg/NET0131  ;
  input \g4064_reg/NET0131  ;
  input \g4072_reg/NET0131  ;
  input \g4076_reg/NET0131  ;
  input \g4082_reg/NET0131  ;
  input \g4087_reg/NET0131  ;
  input \g4093_reg/NET0131  ;
  input \g4098_reg/NET0131  ;
  input \g4104_reg/NET0131  ;
  input \g4108_reg/NET0131  ;
  input \g4112_reg/NET0131  ;
  input \g4116_reg/NET0131  ;
  input \g4119_reg/NET0131  ;
  input \g411_reg/NET0131  ;
  input \g4122_reg/NET0131  ;
  input \g4141_reg/NET0131  ;
  input \g4145_reg/NET0131  ;
  input \g4146_reg/NET0131  ;
  input \g4153_reg/NET0131  ;
  input \g4157_reg/NET0131  ;
  input \g4164_reg/NET0131  ;
  input \g4172_reg/NET0131  ;
  input \g4176_reg/NET0131  ;
  input \g417_reg/NET0131  ;
  input \g4180_reg/NET0131  ;
  input \g4235_reg/NET0131  ;
  input \g4239_reg/NET0131  ;
  input \g4242_reg/NET0131  ;
  input \g4245_reg/NET0131  ;
  input \g424_reg/NET0131  ;
  input \g4253_reg/NET0131  ;
  input \g4258_reg/NET0131  ;
  input \g4264_reg/NET0131  ;
  input \g4269_reg/NET0131  ;
  input \g4273_reg/NET0131  ;
  input \g4281_reg/NET0131  ;
  input \g4284_reg/NET0131  ;
  input \g4291_reg/NET0131  ;
  input \g4297_reg/NET0131  ;
  input \g4300_reg/NET0131  ;
  input \g4308_reg/NET0131  ;
  input \g4311_reg/NET0131  ;
  input \g4322_reg/NET0131  ;
  input \g4332_reg/NET0131  ;
  input \g433_reg/NET0131  ;
  input \g4340_reg/NET0131  ;
  input \g4349_reg/NET0131  ;
  input \g4358_reg/NET0131  ;
  input \g4366_reg/NET0131  ;
  input \g4369_reg/NET0131  ;
  input \g4372_reg/NET0131  ;
  input \g4375_reg/NET0131  ;
  input \g437_reg/NET0131  ;
  input \g4382_reg/NET0131  ;
  input \g4388_reg/NET0131  ;
  input \g4392_reg/NET0131  ;
  input \g4401_reg/NET0131  ;
  input \g4405_reg/NET0131  ;
  input \g4411_reg/NET0131  ;
  input \g4417_reg/NET0131  ;
  input \g441_reg/NET0131  ;
  input \g4420_reg/NET0131  ;
  input \g4423_reg/NET0131  ;
  input \g4427_reg/NET0131  ;
  input \g4430_reg/NET0131  ;
  input \g4434_reg/NET0131  ;
  input \g4438_reg/NET0131  ;
  input \g4443_reg/NET0131  ;
  input \g4452_reg/NET0131  ;
  input \g4455_reg/NET0131  ;
  input \g4459_reg/NET0131  ;
  input \g4462_reg/NET0131  ;
  input \g4467_reg/NET0131  ;
  input \g446_reg/NET0131  ;
  input \g4473_reg/NET0131  ;
  input \g4477_reg/NET0131  ;
  input \g4480_reg/NET0131  ;
  input \g4483_reg/NET0131  ;
  input \g4486_reg/NET0131  ;
  input \g4489_reg/NET0131  ;
  input \g4492_reg/NET0131  ;
  input \g4495_reg/NET0131  ;
  input \g4498_reg/NET0131  ;
  input \g4501_reg/NET0131  ;
  input \g4504_reg/NET0131  ;
  input \g4512_reg/NET0131  ;
  input \g4515_reg/NET0131  ;
  input \g4521_reg/NET0131  ;
  input \g4527_reg/NET0131  ;
  input \g452_reg/NET0131  ;
  input \g4531_reg/NET0131  ;
  input \g4534_reg/NET0131  ;
  input \g4540_reg/NET0131  ;
  input \g4543_reg/NET0131  ;
  input \g4546_reg/NET0131  ;
  input \g4549_reg/NET0131  ;
  input \g4552_reg/NET0131  ;
  input \g4555_reg/NET0131  ;
  input \g4558_reg/NET0131  ;
  input \g4561_reg/NET0131  ;
  input \g4564_reg/NET0131  ;
  input \g4567_reg/NET0131  ;
  input \g4572_reg/NET0131  ;
  input \g4575_reg/NET0131  ;
  input \g4581_reg/NET0131  ;
  input \g4584_reg/NET0131  ;
  input \g4593_reg/NET0131  ;
  input \g4601_reg/NET0131  ;
  input \g4608_reg/NET0131  ;
  input \g460_reg/NET0131  ;
  input \g4616_reg/NET0131  ;
  input \g4621_reg/NET0131  ;
  input \g4628_reg/NET0131  ;
  input \g4633_reg/NET0131  ;
  input \g4639_reg/NET0131  ;
  input \g4643_reg/NET0131  ;
  input \g4646_reg/NET0131  ;
  input \g4653_reg/NET0131  ;
  input \g4659_reg/NET0131  ;
  input \g4664_reg/NET0131  ;
  input \g4669_reg/NET0131  ;
  input \g4674_reg/NET0131  ;
  input \g4681_reg/NET0131  ;
  input \g4688_reg/NET0131  ;
  input \g4698_reg/NET0131  ;
  input \g4704_reg/NET0131  ;
  input \g4709_reg/NET0131  ;
  input \g4743_reg/NET0131  ;
  input \g4749_reg/NET0131  ;
  input \g4754_reg/NET0131  ;
  input \g475_reg/NET0131  ;
  input \g4760_reg/NET0131  ;
  input \g4765_reg/NET0131  ;
  input \g4771_reg/NET0131  ;
  input \g4776_reg/NET0131  ;
  input \g4785_reg/NET0131  ;
  input \g4793_reg/NET0131  ;
  input \g479_reg/NET0131  ;
  input \g4801_reg/NET0131  ;
  input \g482_reg/NET0131  ;
  input \g490_reg/NET0131  ;
  input \g496_reg/NET0131  ;
  input \g499_reg/NET0131  ;
  input \g5016_reg/NET0131  ;
  input \g5022_reg/NET0131  ;
  input \g5029_reg/NET0131  ;
  input \g5033_reg/NET0131  ;
  input \g5037_reg/NET0131  ;
  input \g5041_reg/NET0131  ;
  input \g5046_reg/NET0131  ;
  input \g504_reg/NET0131  ;
  input \g5052_reg/NET0131  ;
  input \g5057_reg/NET0131  ;
  input \g5069_reg/NET0131  ;
  input \g5073_reg/NET0131  ;
  input \g5077_reg/NET0131  ;
  input \g5080_reg/NET0131  ;
  input \g5084_reg/NET0131  ;
  input \g5092_reg/NET0131  ;
  input \g5097_reg/NET0131  ;
  input \g5101_reg/NET0131  ;
  input \g5112_reg/NET0131  ;
  input \g5115_reg/NET0131  ;
  input \g5124_reg/NET0131  ;
  input \g5128_reg/NET0131  ;
  input \g5134_reg/NET0131  ;
  input \g5138_reg/NET0131  ;
  input \g513_reg/NET0131  ;
  input \g5142_reg/NET0131  ;
  input \g5148_reg/NET0131  ;
  input \g5152_reg/NET0131  ;
  input \g518_reg/NET0131  ;
  input \g528_reg/NET0131  ;
  input \g5297_reg/NET0131  ;
  input \g534_reg/NET0131  ;
  input \g5357_reg/NET0131  ;
  input \g538_reg/NET0131  ;
  input \g542_reg/NET0131  ;
  input \g546_reg/NET0131  ;
  input \g550_reg/NET0131  ;
  input \g554_reg/NET0131  ;
  input \g645_reg/NET0131  ;
  input \g650_reg/NET0131  ;
  input \g655_reg/NET0131  ;
  input \g661_reg/NET0131  ;
  input \g667_reg/NET0131  ;
  input \g671_reg/NET0131  ;
  input \g676_reg/NET0131  ;
  input \g681_reg/NET0131  ;
  input \g686_reg/NET0131  ;
  input \g691_reg/NET0131  ;
  input \g699_reg/NET0131  ;
  input \g703_reg/NET0131  ;
  input \g714_reg/NET0131  ;
  input \g718_reg/NET0131  ;
  input \g723_reg/NET0131  ;
  input \g7243_pad  ;
  input \g7245_pad  ;
  input \g7257_pad  ;
  input \g7260_pad  ;
  input \g728_reg/NET0131  ;
  input \g732_reg/NET0131  ;
  input \g736_reg/NET0131  ;
  input \g739_reg/NET0131  ;
  input \g744_reg/NET0131  ;
  input \g749_reg/NET0131  ;
  input \g753_reg/NET0131  ;
  input \g7540_pad  ;
  input \g758_reg/NET0131  ;
  input \g763_reg/NET0131  ;
  input \g767_reg/NET0131  ;
  input \g772_reg/NET0131  ;
  input \g776_reg/NET0131  ;
  input \g781_reg/NET0131  ;
  input \g785_reg/NET0131  ;
  input \g790_reg/NET0131  ;
  input \g7916_pad  ;
  input \g7946_pad  ;
  input \g794_reg/NET0131  ;
  input \g802_reg/NET0131  ;
  input \g807_reg/NET0131  ;
  input \g812_reg/NET0131  ;
  input \g817_reg/NET0131  ;
  input \g822_reg/NET0131  ;
  input \g827_reg/NET0131  ;
  input \g8291_pad  ;
  input \g832_reg/NET0131  ;
  input \g8358_pad  ;
  input \g837_reg/NET0131  ;
  input \g8416_pad  ;
  input \g843_reg/NET0131  ;
  input \g8475_pad  ;
  input \g847_reg/NET0131  ;
  input \g854_reg/NET0131  ;
  input \g862_reg/NET0131  ;
  input \g8719_pad  ;
  input \g872_reg/NET0131  ;
  input \g8783_pad  ;
  input \g8784_pad  ;
  input \g8785_pad  ;
  input \g8786_pad  ;
  input \g8787_pad  ;
  input \g8788_pad  ;
  input \g8789_pad  ;
  input \g8839_pad  ;
  input \g8870_pad  ;
  input \g890_reg/NET0131  ;
  input \g8915_pad  ;
  input \g8916_pad  ;
  input \g8917_pad  ;
  input \g8918_pad  ;
  input \g8919_pad  ;
  input \g8920_pad  ;
  input \g896_reg/NET0131  ;
  input \g9019_pad  ;
  input \g9251_pad  ;
  input \g956_reg/NET0131  ;
  input \g962_reg/NET0131  ;
  input \g969_reg/NET0131  ;
  input \g976_reg/NET0131  ;
  input \g979_reg/NET0131  ;
  input \g990_reg/NET0131  ;
  input \g996_reg/NET0131  ;
  output \g136_reg/P0001  ;
  output \g21727_pad  ;
  output \g23190_pad  ;
  output \g26875_pad  ;
  output \g26876_pad  ;
  output \g26877_pad  ;
  output \g28041_pad  ;
  output \g28042_pad  ;
  output \g30327_pad  ;
  output \g30330_pad  ;
  output \g30331_pad  ;
  output \g31793_pad  ;
  output \g31860_pad  ;
  output \g31862_pad  ;
  output \g31863_pad  ;
  output \g32185_pad  ;
  output \g33079_pad  ;
  output \g33435_pad  ;
  output \g33959_pad  ;
  output \g34435_pad  ;
  output \g34788_pad  ;
  output \g34956_pad  ;
  output \g34_reg/P0001  ;
  output \g35_syn_2  ;
  output \g37/_0_  ;
  output \g41/_0_  ;
  output \g60853/_3_  ;
  output \g60856/_3_  ;
  output \g60879/_3_  ;
  output \g60882/_0_  ;
  output \g60888/_0_  ;
  output \g60891/_0_  ;
  output \g60896/_0_  ;
  output \g60899/_0_  ;
  output \g60900/_3_  ;
  output \g60909/_3_  ;
  output \g60911/_0_  ;
  output \g60915/_0_  ;
  output \g60918/_0_  ;
  output \g60919/_0_  ;
  output \g60928/_0_  ;
  output \g60929/_0_  ;
  output \g60936/_0_  ;
  output \g60937/_0_  ;
  output \g60939/_0_  ;
  output \g60940/_0_  ;
  output \g60941/_0_  ;
  output \g60942/_0_  ;
  output \g60943/_0_  ;
  output \g60944/_0_  ;
  output \g60952/_0_  ;
  output \g60954/_0_  ;
  output \g60958/_0_  ;
  output \g60962/_3_  ;
  output \g60972/_0_  ;
  output \g60980/_0_  ;
  output \g60984/_0_  ;
  output \g60986/_0_  ;
  output \g60989/_0_  ;
  output \g60991/_3_  ;
  output \g61006/_0_  ;
  output \g61008/_0_  ;
  output \g61013/_0_  ;
  output \g61014/_0_  ;
  output \g61015/_0_  ;
  output \g61016/_0_  ;
  output \g61017/_0_  ;
  output \g61026/_3_  ;
  output \g61027/_3_  ;
  output \g61030/_0_  ;
  output \g61031/_0_  ;
  output \g61037/_0_  ;
  output \g61038/_0_  ;
  output \g61042/_0_  ;
  output \g61044/_0_  ;
  output \g61045/_0_  ;
  output \g61046/_0_  ;
  output \g61050/_0_  ;
  output \g61051/_0_  ;
  output \g61052/_0_  ;
  output \g61078/_0_  ;
  output \g61131/_0_  ;
  output \g61137/_3_  ;
  output \g61142/_3_  ;
  output \g61143/_3_  ;
  output \g61151/_0_  ;
  output \g61152/_0_  ;
  output \g61161/_0_  ;
  output \g61168/_3_  ;
  output \g61169/_3_  ;
  output \g61170/_0_  ;
  output \g61171/_3_  ;
  output \g61172/_0_  ;
  output \g61173/_0_  ;
  output \g61174/_0_  ;
  output \g61175/_0_  ;
  output \g61176/_0_  ;
  output \g61177/_3_  ;
  output \g61178/_0_  ;
  output \g61179/_0_  ;
  output \g61180/_0_  ;
  output \g61181/_0_  ;
  output \g61182/_3_  ;
  output \g61183/_0_  ;
  output \g61184/_3_  ;
  output \g61185/_0_  ;
  output \g61186/_0_  ;
  output \g61187/_0_  ;
  output \g61188/_0_  ;
  output \g61189/_0_  ;
  output \g61190/_3_  ;
  output \g61191/_0_  ;
  output \g61192/_0_  ;
  output \g61193/_0_  ;
  output \g61194/_0_  ;
  output \g61221/_0_  ;
  output \g61222/_0_  ;
  output \g61223/_3_  ;
  output \g61224/_3_  ;
  output \g61261/_0_  ;
  output \g61295/_3_  ;
  output \g61308/_0_  ;
  output \g61316/_0_  ;
  output \g61327/_0_  ;
  output \g61329/_0_  ;
  output \g61330/_0_  ;
  output \g61331/_0_  ;
  output \g61332/_3_  ;
  output \g61333/_0_  ;
  output \g61334/_0_  ;
  output \g61335/_0_  ;
  output \g61336/_0_  ;
  output \g61337/_0_  ;
  output \g61338/_3_  ;
  output \g61339/_0_  ;
  output \g61340/_0_  ;
  output \g61341/_0_  ;
  output \g61342/_0_  ;
  output \g61343/_0_  ;
  output \g61344/_3_  ;
  output \g61345/_0_  ;
  output \g61346/_0_  ;
  output \g61347/_0_  ;
  output \g61348/_0_  ;
  output \g61349/_0_  ;
  output \g61350/_3_  ;
  output \g61351/_0_  ;
  output \g61352/_0_  ;
  output \g61353/_0_  ;
  output \g61354/_0_  ;
  output \g61367/_0_  ;
  output \g61372/_0_  ;
  output \g61373/_0_  ;
  output \g61375/_0_  ;
  output \g61382/_0_  ;
  output \g61385/_3_  ;
  output \g61386/_0_  ;
  output \g61399/_0_  ;
  output \g61400/_0_  ;
  output \g61402/_0_  ;
  output \g61405/_0_  ;
  output \g61435/_3_  ;
  output \g61449/_0_  ;
  output \g61468/_0_  ;
  output \g61475/_0_  ;
  output \g61480/_0_  ;
  output \g61482/_0_  ;
  output \g61483/_0_  ;
  output \g61484/_0_  ;
  output \g61486/_3_  ;
  output \g61494/_0_  ;
  output \g61496/_0_  ;
  output \g61497/_0_  ;
  output \g61514/_0_  ;
  output \g61517/_0_  ;
  output \g61519/_3_  ;
  output \g61520/_3_  ;
  output \g61527/_0_  ;
  output \g61541/_0_  ;
  output \g61544/_0_  ;
  output \g61550/_0_  ;
  output \g61551/_0_  ;
  output \g61554/_0_  ;
  output \g61556/_3_  ;
  output \g61567/_0_  ;
  output \g61571/_0_  ;
  output \g61574/_0_  ;
  output \g61587/_0_  ;
  output \g61592/_0_  ;
  output \g61632/_0_  ;
  output \g61634/_0_  ;
  output \g61635/_0_  ;
  output \g61639/_0_  ;
  output \g61644/_0_  ;
  output \g61652/_3_  ;
  output \g61709/_0_  ;
  output \g61714/_0_  ;
  output \g61720/_0_  ;
  output \g61721/_0_  ;
  output \g61723/_0_  ;
  output \g61725/_0_  ;
  output \g61726/_0_  ;
  output \g61734/_0_  ;
  output \g61739/_0_  ;
  output \g61744/_0_  ;
  output \g61746/_3_  ;
  output \g61747/_3_  ;
  output \g61748/_3_  ;
  output \g61750/u3_syn_7  ;
  output \g61802/_0_  ;
  output \g61804/_0_  ;
  output \g61808/_0_  ;
  output \g61811/_0_  ;
  output \g61816/_0_  ;
  output \g61818/_0_  ;
  output \g61820/_0_  ;
  output \g61823/_0_  ;
  output \g61824/_0_  ;
  output \g61841/_0_  ;
  output \g61842/_3_  ;
  output \g61844/_3_  ;
  output \g61845/_3_  ;
  output \g61846/_3_  ;
  output \g61847/u3_syn_7  ;
  output \g61848/_0_  ;
  output \g61849/_3_  ;
  output \g61850/_0_  ;
  output \g61851/u3_syn_7  ;
  output \g61852/_0_  ;
  output \g61853/_3_  ;
  output \g61854/_3_  ;
  output \g61855/_0_  ;
  output \g61856/u3_syn_7  ;
  output \g61857/_0_  ;
  output \g61858/_3_  ;
  output \g61859/_3_  ;
  output \g61860/u3_syn_7  ;
  output \g61861/_0_  ;
  output \g61862/_3_  ;
  output \g61863/_3_  ;
  output \g61864/u3_syn_7  ;
  output \g61865/_0_  ;
  output \g61866/_3_  ;
  output \g61867/_3_  ;
  output \g61868/u3_syn_7  ;
  output \g61869/_0_  ;
  output \g61870/_0_  ;
  output \g61871/_3_  ;
  output \g61872/_3_  ;
  output \g61873/u3_syn_7  ;
  output \g61874/_0_  ;
  output \g61875/_0_  ;
  output \g61877/_3_  ;
  output \g61878/_3_  ;
  output \g61879/u3_syn_7  ;
  output \g61880/_0_  ;
  output \g61881/_0_  ;
  output \g61882/_0_  ;
  output \g61883/_0_  ;
  output \g61884/_0_  ;
  output \g61914/_0_  ;
  output \g61915/_0_  ;
  output \g61917/_0_  ;
  output \g61918/_0_  ;
  output \g61922/_0_  ;
  output \g61923/_0_  ;
  output \g61924/_0_  ;
  output \g61932/_0_  ;
  output \g61936/_0_  ;
  output \g61945/_0_  ;
  output \g61947/_0_  ;
  output \g61959/_0_  ;
  output \g61960/_0_  ;
  output \g61962/_0_  ;
  output \g61973/_3_  ;
  output \g61974/u3_syn_7  ;
  output \g61975/_3_  ;
  output \g61976/u3_syn_7  ;
  output \g61977/_3_  ;
  output \g61978/_3_  ;
  output \g61979/u3_syn_7  ;
  output \g61980/_3_  ;
  output \g61981/_3_  ;
  output \g61982/_3_  ;
  output \g61983/u3_syn_7  ;
  output \g61984/_3_  ;
  output \g61985/_3_  ;
  output \g61986/u3_syn_7  ;
  output \g61987/_3_  ;
  output \g61988/_3_  ;
  output \g61989/u3_syn_7  ;
  output \g61990/_3_  ;
  output \g61991/_3_  ;
  output \g61992/u3_syn_7  ;
  output \g61993/_3_  ;
  output \g61994/u3_syn_7  ;
  output \g61995/_3_  ;
  output \g61996/_3_  ;
  output \g61997/_3_  ;
  output \g62022/_0_  ;
  output \g62028/_0_  ;
  output \g62029/_0_  ;
  output \g62031/_0_  ;
  output \g62033/_0_  ;
  output \g62038/_0_  ;
  output \g62042/_0_  ;
  output \g62046/_0_  ;
  output \g62048/_0_  ;
  output \g62049/_0_  ;
  output \g62051/_0_  ;
  output \g62053/_0_  ;
  output \g62085/_0_  ;
  output \g62101/_0_  ;
  output \g62102/_0_  ;
  output \g62103/_0_  ;
  output \g62105/_0_  ;
  output \g62108/_3_  ;
  output \g62112/_0_  ;
  output \g62137/_3_  ;
  output \g62207/_0_  ;
  output \g62239/_0_  ;
  output \g62240/_0_  ;
  output \g62267/_0_  ;
  output \g62273/_0_  ;
  output \g62284/_0_  ;
  output \g62291/_0_  ;
  output \g62293/_0_  ;
  output \g62298/_0_  ;
  output \g62303/_3_  ;
  output \g62322/_3_  ;
  output \g62323/_3_  ;
  output \g62324/_3_  ;
  output \g62325/_3_  ;
  output \g62583/_0_  ;
  output \g62598/_0_  ;
  output \g62609/_0_  ;
  output \g62636/_0_  ;
  output \g62646/_0_  ;
  output \g62649/_0_  ;
  output \g62658/_0_  ;
  output \g62663/_0_  ;
  output \g62664/_0_  ;
  output \g62667/_0_  ;
  output \g62676/_0_  ;
  output \g62677/_0_  ;
  output \g62678/_3_  ;
  output \g62679/_0_  ;
  output \g62687/u3_syn_7  ;
  output \g62688/u3_syn_7  ;
  output \g62689/_0_  ;
  output \g62690/_3_  ;
  output \g62691/_3_  ;
  output \g62693/_0_  ;
  output \g62694/_3_  ;
  output \g62695/_3_  ;
  output \g62696/_3_  ;
  output \g62697/_3_  ;
  output \g62698/_3_  ;
  output \g62699/_3_  ;
  output \g62700/_3_  ;
  output \g62701/_3_  ;
  output \g62702/_3_  ;
  output \g62703/_3_  ;
  output \g62704/u3_syn_7  ;
  output \g62705/_0_  ;
  output \g62706/_3_  ;
  output \g62707/_3_  ;
  output \g62708/u3_syn_7  ;
  output \g62709/_0_  ;
  output \g62710/_3_  ;
  output \g62711/_3_  ;
  output \g62712/u3_syn_7  ;
  output \g62713/_0_  ;
  output \g62714/_3_  ;
  output \g62715/_0_  ;
  output \g62716/u3_syn_7  ;
  output \g62717/_0_  ;
  output \g62718/_3_  ;
  output \g62719/_0_  ;
  output \g62720/u3_syn_7  ;
  output \g62721/_0_  ;
  output \g62722/_3_  ;
  output \g62723/_0_  ;
  output \g62724/u3_syn_7  ;
  output \g62725/_0_  ;
  output \g62726/_3_  ;
  output \g62728/_0_  ;
  output \g62790/_0_  ;
  output \g62791/_0_  ;
  output \g62793/_0_  ;
  output \g62794/_0_  ;
  output \g62795/_0_  ;
  output \g62796/_0_  ;
  output \g62797/_0_  ;
  output \g62807/_0_  ;
  output \g62823/_0_  ;
  output \g62824/_0_  ;
  output \g62833/_0_  ;
  output \g62846/_0_  ;
  output \g62859/_0_  ;
  output \g62860/_0_  ;
  output \g62897/_0_  ;
  output \g62898/_0_  ;
  output \g62922/_3_  ;
  output \g62923/_0_  ;
  output \g62927/_0_  ;
  output \g62938/_3_  ;
  output \g62939/_3_  ;
  output \g62940/_3_  ;
  output \g62941/u3_syn_7  ;
  output \g62942/_0_  ;
  output \g62943/_3_  ;
  output \g62987/_3_  ;
  output \g62991/_3_  ;
  output \g63015/u3_syn_7  ;
  output \g63016/_0_  ;
  output \g63017/_3_  ;
  output \g63018/_3_  ;
  output \g63019/_3_  ;
  output \g63020/_3_  ;
  output \g63021/_3_  ;
  output \g63022/_3_  ;
  output \g63025/_3_  ;
  output \g63026/_3_  ;
  output \g63027/_3_  ;
  output \g63029/_3_  ;
  output \g63030/_3_  ;
  output \g63031/_3_  ;
  output \g63033/_3_  ;
  output \g63034/_3_  ;
  output \g63043/_3_  ;
  output \g63044/_3_  ;
  output \g63051/_3_  ;
  output \g63057/_3_  ;
  output \g63068/_3_  ;
  output \g63070/_3_  ;
  output \g63073/_3_  ;
  output \g63081/_3_  ;
  output \g63082/_3_  ;
  output \g63083/u3_syn_7  ;
  output \g63084/_3_  ;
  output \g63085/_0_  ;
  output \g63086/_3_  ;
  output \g63107/_3_  ;
  output \g63108/u3_syn_7  ;
  output \g63109/u3_syn_7  ;
  output \g63110/_0_  ;
  output \g63111/_3_  ;
  output \g63132/_3_  ;
  output \g63133/_3_  ;
  output \g63134/_3_  ;
  output \g63135/_3_  ;
  output \g63136/_3_  ;
  output \g63137/_3_  ;
  output \g63138/_3_  ;
  output \g63139/u3_syn_7  ;
  output \g63140/_3_  ;
  output \g63141/_3_  ;
  output \g63142/_3_  ;
  output \g63143/_3_  ;
  output \g63144/_3_  ;
  output \g63145/_3_  ;
  output \g63146/u3_syn_7  ;
  output \g63198/_0_  ;
  output \g63205/_0_  ;
  output \g63208/_0_  ;
  output \g63212/_0_  ;
  output \g63215/_0_  ;
  output \g63219/_0_  ;
  output \g63244/_0_  ;
  output \g63246/_0_  ;
  output \g63254/_0_  ;
  output \g63255/_0_  ;
  output \g63272/_0_  ;
  output \g63276/_0_  ;
  output \g63278/_0_  ;
  output \g63279/_0_  ;
  output \g63280/_0_  ;
  output \g63327/_0_  ;
  output \g63345/_0_  ;
  output \g63346/_3_  ;
  output \g63347/_3_  ;
  output \g63354/_3_  ;
  output \g63358/_3_  ;
  output \g63359/u3_syn_7  ;
  output \g63361/_3_  ;
  output \g63365/_3_  ;
  output \g63366/_3_  ;
  output \g63367/_3_  ;
  output \g63368/_3_  ;
  output \g63370/_3_  ;
  output \g63479/_0_  ;
  output \g63484/_0_  ;
  output \g63499/_1_  ;
  output \g63520/_0_  ;
  output \g63523/_0_  ;
  output \g63526/_0_  ;
  output \g63538/_0_  ;
  output \g63539/_0_  ;
  output \g63541/_0_  ;
  output \g63555/_0_  ;
  output \g63642/_0_  ;
  output \g63645/_0_  ;
  output \g63648/_3_  ;
  output \g63777/_3_  ;
  output \g63778/_3_  ;
  output \g63781/_0_  ;
  output \g63786/u3_syn_7  ;
  output \g63787/_3_  ;
  output \g63788/_3_  ;
  output \g63790/_3_  ;
  output \g63791/_3_  ;
  output \g63792/u3_syn_7  ;
  output \g63794/_0_  ;
  output \g63795/_0_  ;
  output \g63796/_0_  ;
  output \g63798/_3_  ;
  output \g63800/_3_  ;
  output \g63804/_3_  ;
  output \g63805/_3_  ;
  output \g63806/_3_  ;
  output \g63807/_3_  ;
  output \g63808/_3_  ;
  output \g63809/_3_  ;
  output \g63870/_0_  ;
  output \g63883/_0_  ;
  output \g63934/_0_  ;
  output \g63936/_0_  ;
  output \g63938/_0_  ;
  output \g63939/_0_  ;
  output \g63966/_0_  ;
  output \g63970/_0_  ;
  output \g63999/_0_  ;
  output \g64039/_0_  ;
  output \g64040/_0_  ;
  output \g64043/_0_  ;
  output \g64062/_3_  ;
  output \g64078/_0_  ;
  output \g64091/_0_  ;
  output \g64095/_3_  ;
  output \g64096/_3_  ;
  output \g64097/u3_syn_7  ;
  output \g64098/u3_syn_7  ;
  output \g64099/u3_syn_7  ;
  output \g64100/u3_syn_7  ;
  output \g64134/_0_  ;
  output \g64135/_0_  ;
  output \g64153/_0_  ;
  output \g64155/_0_  ;
  output \g64179/_0_  ;
  output \g64229/_0_  ;
  output \g64235/_0_  ;
  output \g64236/_0_  ;
  output \g64280/_0_  ;
  output \g64315/_0_  ;
  output \g64365/_0_  ;
  output \g64426/_3_  ;
  output \g64438/_3_  ;
  output \g64442/u3_syn_7  ;
  output \g64445/_3_  ;
  output \g64447/_3_  ;
  output \g64449/_3_  ;
  output \g64451/_3_  ;
  output \g64453/_3_  ;
  output \g64454/_3_  ;
  output \g64460/_3_  ;
  output \g64461/_3_  ;
  output \g64510/_0_  ;
  output \g64527/_0_  ;
  output \g64528/_0_  ;
  output \g64544/_0_  ;
  output \g64549/_0_  ;
  output \g64566/_0_  ;
  output \g64576/_0_  ;
  output \g64602/_0_  ;
  output \g64691/_0_  ;
  output \g64697/_0_  ;
  output \g64707/_3_  ;
  output \g64778/_3_  ;
  output \g64790/_3_  ;
  output \g64791/_3_  ;
  output \g64792/_3_  ;
  output \g64793/_3_  ;
  output \g64794/_3_  ;
  output \g64795/_3_  ;
  output \g64796/_3_  ;
  output \g64797/_3_  ;
  output \g64877/_0_  ;
  output \g64912/_0_  ;
  output \g64973/_0_  ;
  output \g65047/_3_  ;
  output \g65081/_3_  ;
  output \g65088/_3_  ;
  output \g65097/_3_  ;
  output \g65100/_3_  ;
  output \g65101/_3_  ;
  output \g65104/_3_  ;
  output \g65105/_3_  ;
  output \g65107/_3_  ;
  output \g65110/_3_  ;
  output \g65111/_3_  ;
  output \g65113/_3_  ;
  output \g65114/_3_  ;
  output \g65266/_0_  ;
  output \g65267/_0_  ;
  output \g65294/_1_  ;
  output \g65328/_1_  ;
  output \g65495/_0_  ;
  output \g65499/_0_  ;
  output \g65503/_0_  ;
  output \g65529/_0_  ;
  output \g65530/_3_  ;
  output \g65531/_3_  ;
  output \g65532/_3_  ;
  output \g65533/_3_  ;
  output \g65624/_0_  ;
  output \g65625/_1_  ;
  output \g65641/_0_  ;
  output \g65701/_0_  ;
  output \g65704/_0_  ;
  output \g65853/_0_  ;
  output \g65891/_0_  ;
  output \g65901/_0_  ;
  output \g65986/_0_  ;
  output \g66029/_0_  ;
  output \g66066/_0_  ;
  output \g66067/_0_  ;
  output \g66068/_0_  ;
  output \g66154/_3_  ;
  output \g66362/_0_  ;
  output \g66369/_0_  ;
  output \g66398/_0_  ;
  output \g66409/_0_  ;
  output \g66419/_0_  ;
  output \g66439/_0_  ;
  output \g66443/_0_  ;
  output \g66464/_0_  ;
  output \g66471/_0_  ;
  output \g66512/_0_  ;
  output \g66528/_0_  ;
  output \g66541/_0_  ;
  output \g66558/_0_  ;
  output \g66644/_0_  ;
  output \g66684/_0_  ;
  output \g66697/_0_  ;
  output \g66698/_0_  ;
  output \g66701/_0_  ;
  output \g66714/_0_  ;
  output \g66715/_0_  ;
  output \g66745/_0_  ;
  output \g66750/_0_  ;
  output \g66751/_0_  ;
  output \g66810/_0_  ;
  output \g66844/_0_  ;
  output \g66853/_0_  ;
  output \g66897/_0_  ;
  output \g66905/_0_  ;
  output \g69743/_0_  ;
  output \g69750/_0_  ;
  output \g69773/_1_  ;
  output \g69792/_1_  ;
  output \g69858/_0_  ;
  output \g69938/_0_  ;
  output \g69949/_0_  ;
  output \g70167/_0_  ;
  output \g71190/_0_  ;
  output \g71198/_0_  ;
  output \g71284/_0_  ;
  output \g72369/_1_  ;
  output \g72467/_0_  ;
  output \g72476/_0_  ;
  output \g72477/_1_  ;
  output \g72648/_0_  ;
  output \g72741/_0_  ;
  output \g72772/_0_  ;
  output \g8132_pad  ;
  wire n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 ;
  assign n774 = \g3003_reg/NET0131  & ~\g35_pad  ;
  assign n775 = ~\g2255_reg/NET0131  & ~\g2389_reg/NET0131  ;
  assign n776 = ~\g2523_reg/NET0131  & ~\g2657_reg/NET0131  ;
  assign n777 = n775 & n776 ;
  assign n778 = ~\g1696_reg/NET0131  & ~\g1830_reg/NET0131  ;
  assign n779 = ~\g1964_reg/NET0131  & ~\g2098_reg/NET0131  ;
  assign n780 = n778 & n779 ;
  assign n781 = \g35_pad  & ~n780 ;
  assign n782 = ~n777 & n781 ;
  assign n783 = ~\g1978_reg/NET0131  & ~\g1992_reg/NET0131  ;
  assign n784 = ~\g2112_reg/NET0131  & ~\g2126_reg/NET0131  ;
  assign n785 = n783 & n784 ;
  assign n786 = ~\g1710_reg/NET0131  & ~\g1724_reg/NET0131  ;
  assign n787 = ~\g1844_reg/NET0131  & ~\g1858_reg/NET0131  ;
  assign n788 = n786 & n787 ;
  assign n789 = n785 & n788 ;
  assign n790 = \g35_pad  & ~n789 ;
  assign n791 = ~\g2537_reg/NET0131  & ~\g2551_reg/NET0131  ;
  assign n792 = ~\g2671_reg/NET0131  & ~\g2685_reg/NET0131  ;
  assign n793 = n791 & n792 ;
  assign n794 = ~\g2269_reg/NET0131  & ~\g2283_reg/NET0131  ;
  assign n795 = ~\g2403_reg/NET0131  & ~\g2417_reg/NET0131  ;
  assign n796 = n794 & n795 ;
  assign n797 = n793 & n796 ;
  assign n798 = n790 & ~n797 ;
  assign n799 = ~\g2472_reg/NET0131  & ~\g2491_reg/NET0131  ;
  assign n800 = ~\g2606_reg/NET0131  & ~\g2625_reg/NET0131  ;
  assign n801 = n799 & n800 ;
  assign n802 = ~\g2204_reg/NET0131  & ~\g2223_reg/NET0131  ;
  assign n803 = ~\g2338_reg/NET0131  & ~\g2357_reg/NET0131  ;
  assign n804 = n802 & n803 ;
  assign n805 = n801 & n804 ;
  assign n806 = \g35_pad  & ~n805 ;
  assign n807 = ~\g1913_reg/NET0131  & ~\g1932_reg/NET0131  ;
  assign n808 = ~\g2047_reg/NET0131  & ~\g2066_reg/NET0131  ;
  assign n809 = n807 & n808 ;
  assign n810 = ~\g1644_reg/NET0131  & ~\g1664_reg/NET0131  ;
  assign n811 = ~\g1779_reg/NET0131  & ~\g1798_reg/NET0131  ;
  assign n812 = n810 & n811 ;
  assign n813 = n809 & n812 ;
  assign n814 = n806 & ~n813 ;
  assign n815 = ~\g1312_reg/NET0131  & ~\g1351_reg/NET0131  ;
  assign n816 = \g1536_reg/NET0131  & ~n815 ;
  assign n817 = ~\g1008_reg/NET0131  & ~\g969_reg/NET0131  ;
  assign n818 = \g1193_reg/NET0131  & ~n817 ;
  assign n819 = \g35_pad  & ~n818 ;
  assign n820 = ~n816 & n819 ;
  assign n821 = ~\g1306_reg/NET0131  & \g35_pad  ;
  assign n822 = ~\g962_reg/NET0131  & n821 ;
  assign n823 = ~\g3115_reg/NET0131  & ~\g3466_reg/NET0131  ;
  assign n824 = ~\g3817_reg/NET0131  & ~\g5124_reg/NET0131  ;
  assign n825 = n823 & n824 ;
  assign n826 = \g35_pad  & ~n825 ;
  assign n827 = \g5297_reg/NET0131  & \g5357_reg/NET0131  ;
  assign n828 = ~\g1636_reg/NET0131  & \g1668_reg/NET0131  ;
  assign n829 = \g1648_reg/NET0131  & ~\g1657_reg/NET0131  ;
  assign n830 = \g2902_reg/NET0131  & \g2907_reg/NET0131  ;
  assign n831 = \g2912_reg/NET0131  & \g2917_reg/NET0131  ;
  assign n832 = \g2936_reg/NET0131  & \g2941_reg/NET0131  ;
  assign n833 = ~n831 & ~n832 ;
  assign n834 = ~n830 & n833 ;
  assign n835 = \g2970_reg/NET0131  & \g2975_reg/NET0131  ;
  assign n836 = \g2960_reg/NET0131  & \g2965_reg/NET0131  ;
  assign n837 = ~n835 & ~n836 ;
  assign n838 = \g2922_reg/NET0131  & \g2927_reg/NET0131  ;
  assign n839 = \g2950_reg/NET0131  & \g2955_reg/NET0131  ;
  assign n840 = ~n838 & ~n839 ;
  assign n841 = n837 & n840 ;
  assign n842 = n834 & n841 ;
  assign n843 = \g2724_reg/NET0131  & \g2819_reg/NET0131  ;
  assign n844 = ~\g2724_reg/NET0131  & \g2815_reg/NET0131  ;
  assign n845 = \g2729_reg/NET0131  & ~n844 ;
  assign n846 = ~n843 & n845 ;
  assign n847 = \g2724_reg/NET0131  & \g2807_reg/NET0131  ;
  assign n848 = ~\g2724_reg/NET0131  & \g2803_reg/NET0131  ;
  assign n849 = ~\g2729_reg/NET0131  & ~n848 ;
  assign n850 = ~n847 & n849 ;
  assign n851 = ~n846 & ~n850 ;
  assign n852 = \g2724_reg/NET0131  & \g2787_reg/NET0131  ;
  assign n853 = ~\g2724_reg/NET0131  & \g2783_reg/NET0131  ;
  assign n854 = \g2729_reg/NET0131  & ~n853 ;
  assign n855 = ~n852 & n854 ;
  assign n856 = \g2724_reg/NET0131  & \g2775_reg/NET0131  ;
  assign n857 = ~\g2724_reg/NET0131  & \g2771_reg/NET0131  ;
  assign n858 = ~\g2729_reg/NET0131  & ~n857 ;
  assign n859 = ~n856 & n858 ;
  assign n860 = ~n855 & ~n859 ;
  assign n861 = ~\g4709_reg/NET0131  & ~\g4785_reg/NET0131  ;
  assign n862 = \g4698_reg/NET0131  & n861 ;
  assign n863 = \g4776_reg/NET0131  & ~\g4801_reg/NET0131  ;
  assign n864 = ~\g4793_reg/NET0131  & n863 ;
  assign n865 = \g4659_reg/NET0131  & \g4669_reg/NET0131  ;
  assign n866 = \g4653_reg/NET0131  & n865 ;
  assign n867 = n864 & n866 ;
  assign n868 = n862 & n867 ;
  assign n869 = \g4646_reg/NET0131  & ~n868 ;
  assign n870 = ~\g4057_reg/NET0131  & ~\g4064_reg/NET0131  ;
  assign n871 = ~\g4082_reg/NET0131  & ~\g4141_reg/NET0131  ;
  assign n872 = n870 & ~n871 ;
  assign n873 = ~\g4087_reg/NET0131  & ~\g4093_reg/NET0131  ;
  assign n874 = ~\g4098_reg/NET0131  & n873 ;
  assign n875 = \g4076_reg/NET0131  & \g4112_reg/NET0131  ;
  assign n876 = n870 & n875 ;
  assign n877 = n874 & n876 ;
  assign n878 = ~n872 & ~n877 ;
  assign n879 = ~\g482_reg/NET0131  & ~\g490_reg/NET0131  ;
  assign n880 = \g479_reg/NET0131  & ~\g528_reg/NET0131  ;
  assign n881 = n879 & n880 ;
  assign n882 = \g890_reg/NET0131  & ~n881 ;
  assign n883 = ~\g4311_reg/NET0131  & ~\g4322_reg/NET0131  ;
  assign n884 = ~\g4332_reg/NET0131  & ~\g4366_reg/NET0131  ;
  assign n885 = n883 & n884 ;
  assign n886 = \g4369_reg/NET0131  & ~n885 ;
  assign n887 = \g16686_pad  & \g3247_reg/NET0131  ;
  assign n888 = \g16624_pad  & \g3263_reg/NET0131  ;
  assign n889 = ~n887 & ~n888 ;
  assign n890 = \g3338_reg/NET0131  & ~n889 ;
  assign n891 = \g16874_pad  & \g3223_reg/NET0131  ;
  assign n892 = \g3207_reg/NET0131  & \g3303_reg/NET0131  ;
  assign n893 = ~n891 & ~n892 ;
  assign n894 = ~\g3338_reg/NET0131  & ~n893 ;
  assign n895 = ~n890 & ~n894 ;
  assign n896 = ~\g3303_reg/NET0131  & ~\g3338_reg/NET0131  ;
  assign n897 = \g3303_reg/NET0131  & \g3338_reg/NET0131  ;
  assign n898 = ~n896 & ~n897 ;
  assign n899 = \g16718_pad  & \g3235_reg/NET0131  ;
  assign n900 = ~n898 & n899 ;
  assign n901 = \g3990_reg/NET0131  & ~n900 ;
  assign n902 = n895 & n901 ;
  assign n903 = \g3191_reg/NET0131  & \g3303_reg/NET0131  ;
  assign n904 = \g16874_pad  & \g3215_reg/NET0131  ;
  assign n905 = ~n903 & ~n904 ;
  assign n906 = \g3338_reg/NET0131  & ~n905 ;
  assign n907 = \g16686_pad  & \g3255_reg/NET0131  ;
  assign n908 = \g16624_pad  & \g3203_reg/NET0131  ;
  assign n909 = ~n907 & ~n908 ;
  assign n910 = ~\g3338_reg/NET0131  & ~n909 ;
  assign n911 = ~n906 & ~n910 ;
  assign n912 = \g16718_pad  & \g3243_reg/NET0131  ;
  assign n913 = n898 & n912 ;
  assign n914 = ~\g3990_reg/NET0131  & ~n913 ;
  assign n915 = n911 & n914 ;
  assign n916 = \g4054_reg/NET0131  & ~n915 ;
  assign n917 = ~n902 & n916 ;
  assign n918 = \g16603_pad  & \g3259_reg/NET0131  ;
  assign n919 = n898 & ~n918 ;
  assign n920 = \g13895_pad  & \g3219_reg/NET0131  ;
  assign n921 = ~n898 & ~n920 ;
  assign n922 = ~n919 & ~n921 ;
  assign n923 = \g13039_pad  & \g3199_reg/NET0131  ;
  assign n924 = \g3211_reg/NET0131  & \g3329_reg/NET0131  ;
  assign n925 = ~n923 & ~n924 ;
  assign n926 = ~\g3338_reg/NET0131  & ~n925 ;
  assign n927 = \g13865_pad  & \g3231_reg/NET0131  ;
  assign n928 = \g3338_reg/NET0131  & n927 ;
  assign n929 = \g3990_reg/NET0131  & ~n928 ;
  assign n930 = ~n926 & n929 ;
  assign n931 = ~n922 & n930 ;
  assign n932 = \g13895_pad  & \g3227_reg/NET0131  ;
  assign n933 = n898 & ~n932 ;
  assign n934 = \g16603_pad  & \g3251_reg/NET0131  ;
  assign n935 = ~n898 & ~n934 ;
  assign n936 = ~n933 & ~n935 ;
  assign n937 = \g13039_pad  & \g3187_reg/NET0131  ;
  assign n938 = \g3195_reg/NET0131  & \g3329_reg/NET0131  ;
  assign n939 = ~n937 & ~n938 ;
  assign n940 = \g3338_reg/NET0131  & ~n939 ;
  assign n941 = \g13865_pad  & \g3239_reg/NET0131  ;
  assign n942 = ~\g3338_reg/NET0131  & n941 ;
  assign n943 = ~\g3990_reg/NET0131  & ~n942 ;
  assign n944 = ~n940 & n943 ;
  assign n945 = ~n936 & n944 ;
  assign n946 = ~\g4054_reg/NET0131  & ~n945 ;
  assign n947 = ~n931 & n946 ;
  assign n948 = ~n917 & ~n947 ;
  assign n949 = \g4709_reg/NET0131  & \g4785_reg/NET0131  ;
  assign n950 = \g4765_reg/NET0131  & n949 ;
  assign n951 = n867 & n950 ;
  assign n952 = \g35_pad  & \g4688_reg/NET0131  ;
  assign n953 = ~n951 & n952 ;
  assign n954 = \g16624_pad  & \g3338_reg/NET0131  ;
  assign n955 = \g3990_reg/NET0131  & \g4054_reg/NET0131  ;
  assign n956 = n954 & n955 ;
  assign n957 = \g3808_reg/NET0131  & ~n956 ;
  assign n958 = n953 & ~n957 ;
  assign n959 = ~n948 & n958 ;
  assign n960 = n953 & n957 ;
  assign n961 = n948 & n960 ;
  assign n962 = ~n959 & ~n961 ;
  assign n963 = \g3111_reg/NET0131  & ~\g35_pad  ;
  assign n964 = \g35_pad  & ~\g4688_reg/NET0131  ;
  assign n965 = \g35_pad  & n950 ;
  assign n966 = n867 & n965 ;
  assign n967 = ~n964 & ~n966 ;
  assign n968 = \g3808_reg/NET0131  & ~n967 ;
  assign n969 = ~n963 & ~n968 ;
  assign n970 = n962 & n969 ;
  assign n971 = ~\g528_reg/NET0131  & n879 ;
  assign n972 = \g554_reg/NET0131  & \g807_reg/NET0131  ;
  assign n973 = ~\g499_reg/NET0131  & ~\g518_reg/NET0131  ;
  assign n974 = ~n972 & n973 ;
  assign n975 = n971 & n974 ;
  assign n976 = ~\g736_reg/NET0131  & \g802_reg/NET0131  ;
  assign n977 = \g749_reg/NET0131  & \g758_reg/NET0131  ;
  assign n978 = ~n976 & n977 ;
  assign n979 = \g739_reg/NET0131  & \g744_reg/NET0131  ;
  assign n980 = \g763_reg/NET0131  & \g767_reg/NET0131  ;
  assign n981 = n979 & n980 ;
  assign n982 = \g358_reg/NET0131  & \g376_reg/NET0131  ;
  assign n983 = ~n976 & n982 ;
  assign n984 = n981 & n983 ;
  assign n985 = n978 & n984 ;
  assign n986 = n975 & n985 ;
  assign n987 = \g655_reg/NET0131  & \g718_reg/NET0131  ;
  assign n988 = \g753_reg/NET0131  & n987 ;
  assign n989 = ~\g370_reg/NET0131  & \g385_reg/NET0131  ;
  assign n990 = ~n988 & n989 ;
  assign n991 = \g12184_pad  & ~\g802_reg/NET0131  ;
  assign n992 = ~\g655_reg/NET0131  & ~\g718_reg/NET0131  ;
  assign n993 = ~\g753_reg/NET0131  & n992 ;
  assign n994 = ~n991 & ~n993 ;
  assign n995 = n990 & n994 ;
  assign n996 = \g772_reg/NET0131  & ~n976 ;
  assign n997 = \g776_reg/NET0131  & n996 ;
  assign n998 = n995 & n997 ;
  assign n999 = n986 & n998 ;
  assign n1000 = \g785_reg/NET0131  & ~n976 ;
  assign n1001 = \g781_reg/NET0131  & \g790_reg/NET0131  ;
  assign n1002 = n1000 & n1001 ;
  assign n1003 = \g794_reg/NET0131  & n1002 ;
  assign n1004 = \g35_pad  & \g807_reg/NET0131  ;
  assign n1005 = ~n976 & n1004 ;
  assign n1006 = ~\g554_reg/NET0131  & n1005 ;
  assign n1007 = n1003 & n1006 ;
  assign n1008 = n999 & n1007 ;
  assign n1009 = \g35_pad  & \g554_reg/NET0131  ;
  assign n1010 = ~n976 & n1009 ;
  assign n1011 = ~\g35_pad  & \g807_reg/NET0131  ;
  assign n1012 = ~n1010 & ~n1011 ;
  assign n1013 = ~n1008 & n1012 ;
  assign n1014 = ~\g2941_reg/NET0131  & ~\g35_pad  ;
  assign n1015 = \g35_pad  & n780 ;
  assign n1016 = n777 & n1015 ;
  assign n1017 = ~\g4420_reg/NET0131  & ~\g4427_reg/NET0131  ;
  assign n1018 = ~\g2946_reg/NET0131  & ~\g2955_reg/NET0131  ;
  assign n1019 = n1017 & n1018 ;
  assign n1020 = n825 & n1019 ;
  assign n1021 = n789 & n1020 ;
  assign n1022 = ~\g3831_reg/NET0131  & ~\g3845_reg/NET0131  ;
  assign n1023 = ~\g5138_reg/NET0131  & ~\g5152_reg/NET0131  ;
  assign n1024 = n1022 & n1023 ;
  assign n1025 = ~\g3129_reg/NET0131  & ~\g3143_reg/NET0131  ;
  assign n1026 = ~\g3480_reg/NET0131  & ~\g3494_reg/NET0131  ;
  assign n1027 = n1025 & n1026 ;
  assign n1028 = n1024 & n1027 ;
  assign n1029 = n797 & n1028 ;
  assign n1030 = n1021 & n1029 ;
  assign n1031 = n1016 & n1030 ;
  assign n1032 = ~n1014 & ~n1031 ;
  assign n1033 = ~\g2856_reg/NET0131  & ~\g35_pad  ;
  assign n1034 = ~\g2864_reg/NET0131  & \g35_pad  ;
  assign n1035 = n1017 & n1034 ;
  assign n1036 = n825 & n1035 ;
  assign n1037 = ~n1033 & ~n1036 ;
  assign n1038 = \g10306_pad  & \g35_pad  ;
  assign n1039 = ~\g4534_reg/NET0131  & ~n1038 ;
  assign n1040 = \g4534_reg/NET0131  & n1038 ;
  assign n1041 = ~n1039 & ~n1040 ;
  assign n1042 = ~\g35_pad  & \g4564_reg/NET0131  ;
  assign n1043 = \g4555_reg/NET0131  & \g4558_reg/NET0131  ;
  assign n1044 = \g4561_reg/NET0131  & \g4564_reg/NET0131  ;
  assign n1045 = n1043 & n1044 ;
  assign n1046 = ~n1042 & ~n1045 ;
  assign n1047 = \g2988_reg/NET0131  & \g35_pad  ;
  assign n1048 = n1046 & ~n1047 ;
  assign n1049 = ~\g35_pad  & \g4561_reg/NET0131  ;
  assign n1050 = \g18096_pad  & \g35_pad  ;
  assign n1051 = ~n1049 & ~n1050 ;
  assign n1052 = ~\g35_pad  & \g4558_reg/NET0131  ;
  assign n1053 = \g18095_pad  & \g35_pad  ;
  assign n1054 = ~n1052 & ~n1053 ;
  assign n1055 = ~\g35_pad  & \g4555_reg/NET0131  ;
  assign n1056 = \g18094_pad  & \g35_pad  ;
  assign n1057 = ~n1055 & ~n1056 ;
  assign n1058 = \g4483_reg/NET0131  & \g4486_reg/NET0131  ;
  assign n1059 = \g4489_reg/NET0131  & \g4492_reg/NET0131  ;
  assign n1060 = n1058 & n1059 ;
  assign n1061 = \g35_pad  & ~\g4527_reg/NET0131  ;
  assign n1062 = ~n1060 & n1061 ;
  assign n1063 = \g35_pad  & \g4527_reg/NET0131  ;
  assign n1064 = n1060 & n1063 ;
  assign n1065 = ~n1062 & ~n1064 ;
  assign n1066 = \g4521_reg/NET0131  & n1065 ;
  assign n1067 = ~\g4584_reg/NET0131  & \g4608_reg/NET0131  ;
  assign n1068 = \g4593_reg/NET0131  & ~\g4601_reg/NET0131  ;
  assign n1069 = ~n1067 & ~n1068 ;
  assign n1070 = \g4584_reg/NET0131  & ~\g4608_reg/NET0131  ;
  assign n1071 = \g4593_reg/NET0131  & ~n1070 ;
  assign n1072 = ~n1069 & ~n1071 ;
  assign n1073 = \g35_pad  & ~\g4521_reg/NET0131  ;
  assign n1074 = n1072 & n1073 ;
  assign n1075 = ~\g4593_reg/NET0131  & \g4601_reg/NET0131  ;
  assign n1076 = ~\g4616_reg/NET0131  & ~n1070 ;
  assign n1077 = ~n1075 & n1076 ;
  assign n1078 = n1069 & n1073 ;
  assign n1079 = n1077 & n1078 ;
  assign n1080 = ~n1074 & ~n1079 ;
  assign n1081 = ~n1066 & n1080 ;
  assign n1082 = ~\g35_pad  & \g4527_reg/NET0131  ;
  assign n1083 = ~\g35_pad  & ~n1082 ;
  assign n1084 = ~\g4521_reg/NET0131  & \g4527_reg/NET0131  ;
  assign n1085 = ~n1060 & n1084 ;
  assign n1086 = ~\g4521_reg/NET0131  & ~\g4527_reg/NET0131  ;
  assign n1087 = n1060 & n1086 ;
  assign n1088 = ~n1085 & ~n1087 ;
  assign n1089 = \g4515_reg/NET0131  & \g4521_reg/NET0131  ;
  assign n1090 = ~n1082 & ~n1089 ;
  assign n1091 = n1088 & n1090 ;
  assign n1092 = ~n1083 & ~n1091 ;
  assign n1093 = \g35_pad  & \g4572_reg/NET0131  ;
  assign n1094 = \g4581_reg/NET0131  & n1093 ;
  assign n1095 = \g35_pad  & \g4512_reg/NET0131  ;
  assign n1096 = ~\g4581_reg/NET0131  & n1095 ;
  assign n1097 = ~\g35_pad  & \g4515_reg/NET0131  ;
  assign n1098 = ~n1096 & ~n1097 ;
  assign n1099 = ~n1094 & n1098 ;
  assign n1100 = \g35_pad  & \g4581_reg/NET0131  ;
  assign n1101 = \g4552_reg/NET0131  & ~n1100 ;
  assign n1102 = \g4575_reg/NET0131  & n1100 ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = ~\g35_pad  & ~\g4512_reg/NET0131  ;
  assign n1105 = \g4531_reg/NET0131  & n1100 ;
  assign n1106 = ~n1104 & ~n1105 ;
  assign n1107 = ~\g1322_reg/NET0131  & ~\g1339_reg/NET0131  ;
  assign n1108 = \g1322_reg/NET0131  & \g1339_reg/NET0131  ;
  assign n1109 = ~n1107 & ~n1108 ;
  assign n1110 = \g1351_reg/NET0131  & ~\g1389_reg/NET0131  ;
  assign n1111 = n1109 & ~n1110 ;
  assign n1112 = ~\g1312_reg/NET0131  & ~n1111 ;
  assign n1113 = \g1361_reg/NET0131  & \g1373_reg/NET0131  ;
  assign n1114 = \g1351_reg/NET0131  & n1113 ;
  assign n1115 = ~n1109 & n1114 ;
  assign n1116 = \g1345_reg/NET0131  & \g1361_reg/NET0131  ;
  assign n1117 = \g1367_reg/NET0131  & n1116 ;
  assign n1118 = ~n1115 & ~n1117 ;
  assign n1119 = n1112 & n1118 ;
  assign n1120 = ~\g1322_reg/NET0131  & ~\g1333_reg/NET0131  ;
  assign n1121 = ~\g1312_reg/NET0131  & ~\g1373_reg/NET0131  ;
  assign n1122 = ~n1111 & n1121 ;
  assign n1123 = ~n1120 & ~n1122 ;
  assign n1124 = ~n1119 & n1123 ;
  assign n1125 = ~\g1379_reg/NET0131  & ~n1115 ;
  assign n1126 = n1112 & n1125 ;
  assign n1127 = \g35_pad  & ~n1126 ;
  assign n1128 = n1124 & n1127 ;
  assign n1129 = ~\g1379_reg/NET0131  & \g35_pad  ;
  assign n1130 = ~n1124 & n1129 ;
  assign n1131 = ~n1128 & ~n1130 ;
  assign n1132 = ~\g1373_reg/NET0131  & ~\g35_pad  ;
  assign n1133 = n1131 & ~n1132 ;
  assign n1134 = ~\g1514_reg/NET0131  & ~\g1526_reg/NET0131  ;
  assign n1135 = ~\g1526_reg/NET0131  & ~\g7946_pad  ;
  assign n1136 = \g35_pad  & n1135 ;
  assign n1137 = \g1514_reg/NET0131  & \g7946_pad  ;
  assign n1138 = \g1526_reg/NET0131  & \g35_pad  ;
  assign n1139 = n1137 & n1138 ;
  assign n1140 = ~n1136 & ~n1139 ;
  assign n1141 = ~n1134 & n1140 ;
  assign n1142 = ~\g1514_reg/NET0131  & ~\g35_pad  ;
  assign n1143 = n1141 & ~n1142 ;
  assign n1144 = \g1339_reg/NET0131  & \g1521_reg/NET0131  ;
  assign n1145 = ~\g1532_reg/NET0131  & \g7946_pad  ;
  assign n1146 = n1144 & n1145 ;
  assign n1147 = ~n815 & n1146 ;
  assign n1148 = ~n1109 & ~n1120 ;
  assign n1149 = \g1345_reg/NET0131  & \g1367_reg/NET0131  ;
  assign n1150 = \g1379_reg/NET0131  & n1149 ;
  assign n1151 = n1146 & n1150 ;
  assign n1152 = n1148 & n1151 ;
  assign n1153 = ~n1147 & ~n1152 ;
  assign n1154 = ~\g1514_reg/NET0131  & \g1526_reg/NET0131  ;
  assign n1155 = \g1536_reg/NET0131  & ~n1154 ;
  assign n1156 = ~n1142 & ~n1155 ;
  assign n1157 = ~n1153 & n1156 ;
  assign n1158 = ~n1143 & ~n1157 ;
  assign n1159 = \g1367_reg/NET0131  & ~\g35_pad  ;
  assign n1160 = ~n1119 & ~n1120 ;
  assign n1161 = ~\g1373_reg/NET0131  & ~n1160 ;
  assign n1162 = \g35_pad  & ~n1124 ;
  assign n1163 = ~n1161 & n1162 ;
  assign n1164 = ~n1159 & ~n1163 ;
  assign n1165 = \g4549_reg/NET0131  & ~n1100 ;
  assign n1166 = ~n1102 & ~n1165 ;
  assign n1167 = ~\g1514_reg/NET0131  & ~\g7946_pad  ;
  assign n1168 = ~n1137 & ~n1167 ;
  assign n1169 = \g35_pad  & n1168 ;
  assign n1170 = \g35_pad  & ~n1155 ;
  assign n1171 = ~n1153 & n1170 ;
  assign n1172 = ~n1169 & ~n1171 ;
  assign n1173 = \g1345_reg/NET0131  & ~\g1367_reg/NET0131  ;
  assign n1174 = ~n1120 & n1173 ;
  assign n1175 = ~n1115 & n1174 ;
  assign n1176 = n1112 & n1175 ;
  assign n1177 = \g35_pad  & ~n1176 ;
  assign n1178 = \g1361_reg/NET0131  & ~n1177 ;
  assign n1179 = ~n1115 & ~n1116 ;
  assign n1180 = n1112 & n1179 ;
  assign n1181 = ~n1120 & ~n1180 ;
  assign n1182 = \g1367_reg/NET0131  & \g35_pad  ;
  assign n1183 = ~n1181 & n1182 ;
  assign n1184 = ~n1178 & ~n1183 ;
  assign n1185 = ~n1153 & ~n1155 ;
  assign n1186 = ~\g1532_reg/NET0131  & n1144 ;
  assign n1187 = \g1542_reg/NET0131  & \g7946_pad  ;
  assign n1188 = n1154 & n1187 ;
  assign n1189 = ~n1186 & n1188 ;
  assign n1190 = \g35_pad  & ~n1189 ;
  assign n1191 = \g1413_reg/NET0131  & n1190 ;
  assign n1192 = ~n1185 & n1191 ;
  assign n1193 = ~\g1413_reg/NET0131  & \g7946_pad  ;
  assign n1194 = n1154 & n1193 ;
  assign n1195 = ~n1186 & n1194 ;
  assign n1196 = \g35_pad  & ~n1195 ;
  assign n1197 = \g1542_reg/NET0131  & ~n1196 ;
  assign n1198 = ~n1192 & ~n1197 ;
  assign n1199 = \g1514_reg/NET0131  & ~\g1526_reg/NET0131  ;
  assign n1200 = \g13272_pad  & n1199 ;
  assign n1201 = ~\g1442_reg/NET0131  & ~\g1489_reg/NET0131  ;
  assign n1202 = n1200 & n1201 ;
  assign n1203 = ~\g1437_reg/NET0131  & ~n1202 ;
  assign n1204 = ~\g1319_reg/NET0131  & \g1536_reg/NET0131  ;
  assign n1205 = ~n815 & n1204 ;
  assign n1206 = \g13272_pad  & ~\g1478_reg/NET0131  ;
  assign n1207 = n1199 & n1206 ;
  assign n1208 = ~n1205 & n1207 ;
  assign n1209 = \g13272_pad  & \g1478_reg/NET0131  ;
  assign n1210 = n1199 & n1209 ;
  assign n1211 = n1205 & n1210 ;
  assign n1212 = ~n1208 & ~n1211 ;
  assign n1213 = ~n1203 & n1212 ;
  assign n1214 = \g35_pad  & ~n1213 ;
  assign n1215 = ~\g1442_reg/NET0131  & ~\g35_pad  ;
  assign n1216 = ~n1214 & ~n1215 ;
  assign n1217 = \g13272_pad  & n1154 ;
  assign n1218 = n1201 & n1217 ;
  assign n1219 = ~\g1454_reg/NET0131  & ~n1218 ;
  assign n1220 = \g13272_pad  & ~\g1448_reg/NET0131  ;
  assign n1221 = n1154 & n1220 ;
  assign n1222 = ~n1205 & n1221 ;
  assign n1223 = \g13272_pad  & \g1448_reg/NET0131  ;
  assign n1224 = n1154 & n1223 ;
  assign n1225 = n1205 & n1224 ;
  assign n1226 = ~n1222 & ~n1225 ;
  assign n1227 = ~n1219 & n1226 ;
  assign n1228 = \g35_pad  & ~n1227 ;
  assign n1229 = ~\g1478_reg/NET0131  & ~\g35_pad  ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = \g1514_reg/NET0131  & \g1526_reg/NET0131  ;
  assign n1232 = \g13272_pad  & n1231 ;
  assign n1233 = n1201 & n1232 ;
  assign n1234 = ~\g1467_reg/NET0131  & ~n1233 ;
  assign n1235 = \g13272_pad  & ~\g1472_reg/NET0131  ;
  assign n1236 = n1231 & n1235 ;
  assign n1237 = ~n1205 & n1236 ;
  assign n1238 = \g13272_pad  & \g1472_reg/NET0131  ;
  assign n1239 = n1231 & n1238 ;
  assign n1240 = n1205 & n1239 ;
  assign n1241 = ~n1237 & ~n1240 ;
  assign n1242 = ~n1234 & n1241 ;
  assign n1243 = \g35_pad  & ~n1242 ;
  assign n1244 = ~\g1448_reg/NET0131  & ~\g35_pad  ;
  assign n1245 = ~n1243 & ~n1244 ;
  assign n1246 = \g13272_pad  & n1134 ;
  assign n1247 = n1201 & n1246 ;
  assign n1248 = ~\g1484_reg/NET0131  & ~n1247 ;
  assign n1249 = ~\g1300_reg/NET0131  & \g13272_pad  ;
  assign n1250 = n1134 & n1249 ;
  assign n1251 = ~n1205 & n1250 ;
  assign n1252 = \g1300_reg/NET0131  & \g13272_pad  ;
  assign n1253 = n1134 & n1252 ;
  assign n1254 = n1205 & n1253 ;
  assign n1255 = ~n1251 & ~n1254 ;
  assign n1256 = ~n1248 & n1255 ;
  assign n1257 = \g35_pad  & ~n1256 ;
  assign n1258 = ~\g1472_reg/NET0131  & ~\g35_pad  ;
  assign n1259 = ~n1257 & ~n1258 ;
  assign n1260 = \g4504_reg/NET0131  & ~n1100 ;
  assign n1261 = ~n1094 & ~n1260 ;
  assign n1262 = ~\g1345_reg/NET0131  & ~n1115 ;
  assign n1263 = n1112 & n1262 ;
  assign n1264 = ~n1120 & ~n1263 ;
  assign n1265 = \g1361_reg/NET0131  & \g35_pad  ;
  assign n1266 = ~n1264 & n1265 ;
  assign n1267 = ~\g1361_reg/NET0131  & ~n1120 ;
  assign n1268 = ~n1115 & n1267 ;
  assign n1269 = n1112 & n1268 ;
  assign n1270 = \g35_pad  & ~n1269 ;
  assign n1271 = \g1345_reg/NET0131  & ~n1270 ;
  assign n1272 = ~n1266 & ~n1271 ;
  assign n1273 = ~\g1532_reg/NET0131  & ~\g35_pad  ;
  assign n1274 = \g1413_reg/NET0131  & \g1536_reg/NET0131  ;
  assign n1275 = n1189 & n1274 ;
  assign n1276 = \g35_pad  & n1275 ;
  assign n1277 = ~\g1536_reg/NET0131  & \g35_pad  ;
  assign n1278 = n1153 & n1277 ;
  assign n1279 = ~n1276 & ~n1278 ;
  assign n1280 = ~n1273 & n1279 ;
  assign n1281 = \g1536_reg/NET0131  & ~\g35_pad  ;
  assign n1282 = \g7946_pad  & n1154 ;
  assign n1283 = ~n1186 & n1282 ;
  assign n1284 = ~\g1542_reg/NET0131  & ~n1283 ;
  assign n1285 = n1190 & ~n1284 ;
  assign n1286 = ~n1185 & n1285 ;
  assign n1287 = ~n1281 & ~n1286 ;
  assign n1288 = ~\g333_reg/NET0131  & \g351_reg/NET0131  ;
  assign n1289 = \g35_pad  & ~n1288 ;
  assign n1290 = ~\g355_reg/NET0131  & ~n1289 ;
  assign n1291 = ~\g29211_pad  & ~\g351_reg/NET0131  ;
  assign n1292 = \g35_pad  & n1291 ;
  assign n1293 = ~n1290 & ~n1292 ;
  assign n1294 = ~\g1351_reg/NET0131  & \g1379_reg/NET0131  ;
  assign n1295 = n1149 & n1294 ;
  assign n1296 = ~n1109 & n1295 ;
  assign n1297 = ~n1120 & n1296 ;
  assign n1298 = \g1389_reg/NET0131  & n1109 ;
  assign n1299 = n1114 & ~n1120 ;
  assign n1300 = ~n1298 & n1299 ;
  assign n1301 = ~n1297 & ~n1300 ;
  assign n1302 = n1109 & ~n1120 ;
  assign n1303 = \g1312_reg/NET0131  & ~n1302 ;
  assign n1304 = n1301 & ~n1303 ;
  assign n1305 = \g35_pad  & ~n1304 ;
  assign n1306 = \g1312_reg/NET0131  & ~\g35_pad  ;
  assign n1307 = \g1312_reg/NET0131  & ~n1120 ;
  assign n1308 = n1109 & n1307 ;
  assign n1309 = ~n1306 & ~n1308 ;
  assign n1310 = n1113 & ~n1120 ;
  assign n1311 = \g1389_reg/NET0131  & ~n1120 ;
  assign n1312 = n1109 & n1311 ;
  assign n1313 = ~n1310 & ~n1312 ;
  assign n1314 = \g1351_reg/NET0131  & \g35_pad  ;
  assign n1315 = n1313 & n1314 ;
  assign n1316 = n1309 & ~n1315 ;
  assign n1317 = ~\g333_reg/NET0131  & ~\g355_reg/NET0131  ;
  assign n1318 = ~\g351_reg/NET0131  & \g35_pad  ;
  assign n1319 = ~n1317 & n1318 ;
  assign n1320 = \g351_reg/NET0131  & ~\g35_pad  ;
  assign n1321 = ~n1319 & ~n1320 ;
  assign n1322 = ~\g4546_reg/NET0131  & ~n1100 ;
  assign n1323 = n815 & ~n1120 ;
  assign n1324 = n1109 & n1323 ;
  assign n1325 = \g1322_reg/NET0131  & ~\g1579_reg/NET0131  ;
  assign n1326 = ~\g1322_reg/NET0131  & \g1579_reg/NET0131  ;
  assign n1327 = ~n1325 & ~n1326 ;
  assign n1328 = n1324 & ~n1327 ;
  assign n1329 = ~\g1333_reg/NET0131  & ~\g19357_pad  ;
  assign n1330 = ~\g7946_pad  & n1329 ;
  assign n1331 = ~\g13272_pad  & ~\g8475_pad  ;
  assign n1332 = n1330 & n1331 ;
  assign n1333 = \g35_pad  & ~n1332 ;
  assign n1334 = n1328 & n1333 ;
  assign n1335 = \g35_pad  & n1332 ;
  assign n1336 = ~n1328 & n1335 ;
  assign n1337 = ~n1334 & ~n1336 ;
  assign n1338 = \g1339_reg/NET0131  & ~\g35_pad  ;
  assign n1339 = n1337 & ~n1338 ;
  assign n1340 = \g35_pad  & ~n1327 ;
  assign n1341 = n1324 & n1340 ;
  assign n1342 = ~\g1333_reg/NET0131  & ~n1341 ;
  assign n1343 = \g1333_reg/NET0131  & \g35_pad  ;
  assign n1344 = ~n1327 & n1343 ;
  assign n1345 = n1324 & n1344 ;
  assign n1346 = ~n1342 & ~n1345 ;
  assign n1347 = \g1351_reg/NET0131  & ~\g35_pad  ;
  assign n1348 = ~\g1345_reg/NET0131  & n1120 ;
  assign n1349 = \g35_pad  & ~n1348 ;
  assign n1350 = ~n1264 & n1349 ;
  assign n1351 = ~n1347 & ~n1350 ;
  assign n1352 = ~\g4411_reg/NET0131  & ~\g7243_pad  ;
  assign n1353 = ~\g7257_pad  & n1352 ;
  assign n1354 = ~\g4375_reg/NET0131  & ~\g4405_reg/NET0131  ;
  assign n1355 = \g35_pad  & ~\g4392_reg/NET0131  ;
  assign n1356 = n1354 & n1355 ;
  assign n1357 = n1353 & n1356 ;
  assign n1358 = ~\g4417_reg/NET0131  & n1357 ;
  assign n1359 = n1353 & n1354 ;
  assign n1360 = \g4375_reg/NET0131  & ~\g4382_reg/NET0131  ;
  assign n1361 = ~\g4375_reg/NET0131  & \g4382_reg/NET0131  ;
  assign n1362 = ~n1360 & ~n1361 ;
  assign n1363 = \g35_pad  & ~n1362 ;
  assign n1364 = ~n1359 & n1363 ;
  assign n1365 = ~\g35_pad  & \g4388_reg/NET0131  ;
  assign n1366 = ~n1364 & ~n1365 ;
  assign n1367 = ~n1358 & n1366 ;
  assign n1368 = \g1171_reg/NET0131  & ~\g1183_reg/NET0131  ;
  assign n1369 = \g13259_pad  & n1368 ;
  assign n1370 = ~\g1099_reg/NET0131  & ~\g1146_reg/NET0131  ;
  assign n1371 = n1369 & n1370 ;
  assign n1372 = ~\g1094_reg/NET0131  & ~n1371 ;
  assign n1373 = \g1193_reg/NET0131  & ~\g976_reg/NET0131  ;
  assign n1374 = ~n817 & n1373 ;
  assign n1375 = ~\g1135_reg/NET0131  & \g13259_pad  ;
  assign n1376 = n1368 & n1375 ;
  assign n1377 = ~n1374 & n1376 ;
  assign n1378 = \g1135_reg/NET0131  & \g13259_pad  ;
  assign n1379 = n1368 & n1378 ;
  assign n1380 = n1374 & n1379 ;
  assign n1381 = ~n1377 & ~n1380 ;
  assign n1382 = ~n1372 & n1381 ;
  assign n1383 = \g35_pad  & ~n1382 ;
  assign n1384 = ~\g1099_reg/NET0131  & ~\g35_pad  ;
  assign n1385 = ~n1383 & ~n1384 ;
  assign n1386 = ~\g1171_reg/NET0131  & \g1183_reg/NET0131  ;
  assign n1387 = \g13259_pad  & n1386 ;
  assign n1388 = n1370 & n1387 ;
  assign n1389 = ~\g1111_reg/NET0131  & ~n1388 ;
  assign n1390 = ~\g1105_reg/NET0131  & \g13259_pad  ;
  assign n1391 = n1386 & n1390 ;
  assign n1392 = ~n1374 & n1391 ;
  assign n1393 = \g1105_reg/NET0131  & \g13259_pad  ;
  assign n1394 = n1386 & n1393 ;
  assign n1395 = n1374 & n1394 ;
  assign n1396 = ~n1392 & ~n1395 ;
  assign n1397 = ~n1389 & n1396 ;
  assign n1398 = \g35_pad  & ~n1397 ;
  assign n1399 = ~\g1135_reg/NET0131  & ~\g35_pad  ;
  assign n1400 = ~n1398 & ~n1399 ;
  assign n1401 = \g1171_reg/NET0131  & \g1183_reg/NET0131  ;
  assign n1402 = \g13259_pad  & n1401 ;
  assign n1403 = n1370 & n1402 ;
  assign n1404 = ~\g1124_reg/NET0131  & ~n1403 ;
  assign n1405 = ~\g1129_reg/NET0131  & \g13259_pad  ;
  assign n1406 = n1401 & n1405 ;
  assign n1407 = ~n1374 & n1406 ;
  assign n1408 = \g1129_reg/NET0131  & \g13259_pad  ;
  assign n1409 = n1401 & n1408 ;
  assign n1410 = n1374 & n1409 ;
  assign n1411 = ~n1407 & ~n1410 ;
  assign n1412 = ~n1404 & n1411 ;
  assign n1413 = \g35_pad  & ~n1412 ;
  assign n1414 = ~\g1105_reg/NET0131  & ~\g35_pad  ;
  assign n1415 = ~n1413 & ~n1414 ;
  assign n1416 = ~\g1171_reg/NET0131  & ~\g1183_reg/NET0131  ;
  assign n1417 = \g13259_pad  & n1416 ;
  assign n1418 = n1370 & n1417 ;
  assign n1419 = ~\g1141_reg/NET0131  & ~n1418 ;
  assign n1420 = \g13259_pad  & ~\g956_reg/NET0131  ;
  assign n1421 = n1416 & n1420 ;
  assign n1422 = ~n1374 & n1421 ;
  assign n1423 = \g13259_pad  & \g956_reg/NET0131  ;
  assign n1424 = n1416 & n1423 ;
  assign n1425 = n1374 & n1424 ;
  assign n1426 = ~n1422 & ~n1425 ;
  assign n1427 = ~n1419 & n1426 ;
  assign n1428 = \g35_pad  & ~n1427 ;
  assign n1429 = ~\g1129_reg/NET0131  & ~\g35_pad  ;
  assign n1430 = ~n1428 & ~n1429 ;
  assign n1431 = ~\g4501_reg/NET0131  & ~n1100 ;
  assign n1432 = \g35_pad  & \g4411_reg/NET0131  ;
  assign n1433 = ~\g4401_reg/NET0131  & ~n1432 ;
  assign n1434 = \g4392_reg/NET0131  & n1354 ;
  assign n1435 = n1353 & n1434 ;
  assign n1436 = \g35_pad  & ~n1432 ;
  assign n1437 = ~n1435 & n1436 ;
  assign n1438 = ~n1433 & ~n1437 ;
  assign n1439 = \g4388_reg/NET0131  & n1357 ;
  assign n1440 = ~\g4405_reg/NET0131  & ~n1439 ;
  assign n1441 = \g35_pad  & ~\g4382_reg/NET0131  ;
  assign n1442 = \g4375_reg/NET0131  & ~n1441 ;
  assign n1443 = \g35_pad  & \g4392_reg/NET0131  ;
  assign n1444 = n1354 & n1443 ;
  assign n1445 = n1353 & n1444 ;
  assign n1446 = ~n1442 & ~n1445 ;
  assign n1447 = ~\g35_pad  & \g4455_reg/NET0131  ;
  assign n1448 = ~n1359 & n1443 ;
  assign n1449 = ~n1358 & ~n1448 ;
  assign n1450 = ~n1447 & n1449 ;
  assign n1451 = n1110 & ~n1120 ;
  assign n1452 = n1109 & n1451 ;
  assign n1453 = \g35_pad  & ~n1452 ;
  assign n1454 = \g1384_reg/NET0131  & ~n1453 ;
  assign n1455 = \g1351_reg/NET0131  & ~\g1384_reg/NET0131  ;
  assign n1456 = ~n1120 & ~n1455 ;
  assign n1457 = n1109 & n1456 ;
  assign n1458 = \g1389_reg/NET0131  & \g35_pad  ;
  assign n1459 = ~n1457 & n1458 ;
  assign n1460 = ~n1454 & ~n1459 ;
  assign n1461 = \g1430_reg/NET0131  & \g1548_reg/NET0131  ;
  assign n1462 = \g1554_reg/NET0131  & \g1564_reg/NET0131  ;
  assign n1463 = n1461 & n1462 ;
  assign n1464 = ~n1324 & n1463 ;
  assign n1465 = ~\g17320_pad  & ~\g17404_pad  ;
  assign n1466 = ~\g17423_pad  & \g35_pad  ;
  assign n1467 = n1465 & n1466 ;
  assign n1468 = ~n1464 & n1467 ;
  assign n1469 = ~\g209_reg/NET0131  & \g691_reg/NET0131  ;
  assign n1470 = ~\g1478_reg/NET0131  & n1469 ;
  assign n1471 = n816 & n1470 ;
  assign n1472 = \g35_pad  & ~n1471 ;
  assign n1473 = ~\g1548_reg/NET0131  & ~\g1554_reg/NET0131  ;
  assign n1474 = ~\g1559_reg/NET0131  & ~\g1564_reg/NET0131  ;
  assign n1475 = n1473 & n1474 ;
  assign n1476 = \g1322_reg/NET0131  & \g1404_reg/NET0131  ;
  assign n1477 = n1199 & n1476 ;
  assign n1478 = n1475 & n1477 ;
  assign n1479 = \g17320_pad  & \g35_pad  ;
  assign n1480 = ~n1478 & n1479 ;
  assign n1481 = ~n1472 & ~n1480 ;
  assign n1482 = ~\g2153_reg/NET0131  & ~\g2227_reg/NET0131  ;
  assign n1483 = \g2241_reg/NET0131  & ~n1482 ;
  assign n1484 = ~\g1478_reg/NET0131  & ~\g1589_reg/NET0131  ;
  assign n1485 = n1469 & n1484 ;
  assign n1486 = n816 & n1485 ;
  assign n1487 = ~n1483 & n1486 ;
  assign n1488 = n1483 & ~n1486 ;
  assign n1489 = ~n1487 & ~n1488 ;
  assign n1490 = ~n1481 & n1489 ;
  assign n1491 = \g17320_pad  & ~n1478 ;
  assign n1492 = \g2241_reg/NET0131  & \g35_pad  ;
  assign n1493 = n1471 & n1492 ;
  assign n1494 = ~n1491 & n1493 ;
  assign n1495 = \g2227_reg/NET0131  & ~\g35_pad  ;
  assign n1496 = ~n1494 & ~n1495 ;
  assign n1497 = ~n1490 & n1496 ;
  assign n1498 = ~\g1448_reg/NET0131  & n1469 ;
  assign n1499 = n816 & n1498 ;
  assign n1500 = \g35_pad  & ~n1499 ;
  assign n1501 = n1154 & n1476 ;
  assign n1502 = n1475 & n1501 ;
  assign n1503 = \g17404_pad  & \g35_pad  ;
  assign n1504 = ~n1502 & n1503 ;
  assign n1505 = ~n1500 & ~n1504 ;
  assign n1506 = ~\g2287_reg/NET0131  & ~\g2361_reg/NET0131  ;
  assign n1507 = \g2375_reg/NET0131  & ~n1506 ;
  assign n1508 = ~\g1448_reg/NET0131  & \g1589_reg/NET0131  ;
  assign n1509 = n1469 & n1508 ;
  assign n1510 = n816 & n1509 ;
  assign n1511 = ~n1507 & n1510 ;
  assign n1512 = n1507 & ~n1510 ;
  assign n1513 = ~n1511 & ~n1512 ;
  assign n1514 = ~n1505 & n1513 ;
  assign n1515 = \g17404_pad  & ~n1502 ;
  assign n1516 = \g2375_reg/NET0131  & \g35_pad  ;
  assign n1517 = n1499 & n1516 ;
  assign n1518 = ~n1515 & n1517 ;
  assign n1519 = \g2361_reg/NET0131  & ~\g35_pad  ;
  assign n1520 = ~n1518 & ~n1519 ;
  assign n1521 = ~n1514 & n1520 ;
  assign n1522 = ~\g1472_reg/NET0131  & n1469 ;
  assign n1523 = n816 & n1522 ;
  assign n1524 = \g35_pad  & ~n1523 ;
  assign n1525 = n1231 & n1476 ;
  assign n1526 = n1475 & n1525 ;
  assign n1527 = \g17423_pad  & \g35_pad  ;
  assign n1528 = ~n1526 & n1527 ;
  assign n1529 = ~n1524 & ~n1528 ;
  assign n1530 = ~\g2421_reg/NET0131  & ~\g2495_reg/NET0131  ;
  assign n1531 = \g2509_reg/NET0131  & ~n1530 ;
  assign n1532 = ~\g1472_reg/NET0131  & ~\g1589_reg/NET0131  ;
  assign n1533 = n1469 & n1532 ;
  assign n1534 = n816 & n1533 ;
  assign n1535 = ~n1531 & n1534 ;
  assign n1536 = n1531 & ~n1534 ;
  assign n1537 = ~n1535 & ~n1536 ;
  assign n1538 = ~n1529 & n1537 ;
  assign n1539 = \g17423_pad  & ~n1526 ;
  assign n1540 = \g2509_reg/NET0131  & \g35_pad  ;
  assign n1541 = n1523 & n1540 ;
  assign n1542 = ~n1539 & n1541 ;
  assign n1543 = \g2495_reg/NET0131  & ~\g35_pad  ;
  assign n1544 = ~n1542 & ~n1543 ;
  assign n1545 = ~n1538 & n1544 ;
  assign n1546 = ~\g1300_reg/NET0131  & n1469 ;
  assign n1547 = n816 & n1546 ;
  assign n1548 = \g35_pad  & ~n1547 ;
  assign n1549 = n1134 & n1476 ;
  assign n1550 = n1475 & n1549 ;
  assign n1551 = \g1430_reg/NET0131  & \g35_pad  ;
  assign n1552 = ~n1550 & n1551 ;
  assign n1553 = ~n1548 & ~n1552 ;
  assign n1554 = ~\g2555_reg/NET0131  & ~\g2629_reg/NET0131  ;
  assign n1555 = \g2643_reg/NET0131  & ~n1554 ;
  assign n1556 = ~\g1300_reg/NET0131  & \g1589_reg/NET0131  ;
  assign n1557 = n1469 & n1556 ;
  assign n1558 = n816 & n1557 ;
  assign n1559 = ~n1555 & n1558 ;
  assign n1560 = n1555 & ~n1558 ;
  assign n1561 = ~n1559 & ~n1560 ;
  assign n1562 = ~n1553 & n1561 ;
  assign n1563 = \g1430_reg/NET0131  & ~n1550 ;
  assign n1564 = \g2643_reg/NET0131  & \g35_pad  ;
  assign n1565 = n1547 & n1564 ;
  assign n1566 = ~n1563 & n1565 ;
  assign n1567 = \g2629_reg/NET0131  & ~\g35_pad  ;
  assign n1568 = ~n1566 & ~n1567 ;
  assign n1569 = ~n1562 & n1568 ;
  assign n1570 = ~\g35_pad  & \g4417_reg/NET0131  ;
  assign n1571 = n1449 & ~n1570 ;
  assign n1572 = ~\g35_pad  & \g4411_reg/NET0131  ;
  assign n1573 = \g35_pad  & n1360 ;
  assign n1574 = ~n1572 & ~n1573 ;
  assign n1575 = ~n1357 & n1574 ;
  assign n1576 = \g1379_reg/NET0131  & ~\g35_pad  ;
  assign n1577 = \g35_pad  & ~n1457 ;
  assign n1578 = ~\g1384_reg/NET0131  & ~n1302 ;
  assign n1579 = n1577 & ~n1578 ;
  assign n1580 = ~n1576 & ~n1579 ;
  assign n1581 = ~\g4567_reg/NET0131  & ~n1100 ;
  assign n1582 = ~\g4498_reg/NET0131  & ~n1100 ;
  assign n1583 = \g218_reg/NET0131  & \g8291_pad  ;
  assign n1584 = \g35_pad  & \g8358_pad  ;
  assign n1585 = ~n1583 & n1584 ;
  assign n1586 = ~\g191_reg/NET0131  & \g35_pad  ;
  assign n1587 = n1583 & n1586 ;
  assign n1588 = ~n1585 & ~n1587 ;
  assign n1589 = \g222_reg/NET0131  & ~\g35_pad  ;
  assign n1590 = n1588 & ~n1589 ;
  assign n1591 = \g347_reg/NET0131  & ~\g35_pad  ;
  assign n1592 = ~\g347_reg/NET0131  & \g35_pad  ;
  assign n1593 = \g7540_pad  & n1592 ;
  assign n1594 = ~n1591 & ~n1593 ;
  assign n1595 = ~\g4242_reg/NET0131  & ~\g4300_reg/NET0131  ;
  assign n1596 = \g35_pad  & ~n1595 ;
  assign n1597 = ~\g35_pad  & \g4297_reg/NET0131  ;
  assign n1598 = ~n1596 & ~n1597 ;
  assign n1599 = ~\g1105_reg/NET0131  & n1469 ;
  assign n1600 = n818 & n1599 ;
  assign n1601 = \g35_pad  & ~n1600 ;
  assign n1602 = \g1061_reg/NET0131  & ~\g1205_reg/NET0131  ;
  assign n1603 = ~\g1221_reg/NET0131  & \g979_reg/NET0131  ;
  assign n1604 = n1602 & n1603 ;
  assign n1605 = ~\g1211_reg/NET0131  & ~\g1216_reg/NET0131  ;
  assign n1606 = n1386 & n1605 ;
  assign n1607 = n1604 & n1606 ;
  assign n1608 = \g17316_pad  & \g35_pad  ;
  assign n1609 = ~n1607 & n1608 ;
  assign n1610 = ~n1601 & ~n1609 ;
  assign n1611 = ~\g1728_reg/NET0131  & ~\g1802_reg/NET0131  ;
  assign n1612 = \g1816_reg/NET0131  & ~n1611 ;
  assign n1613 = ~\g1105_reg/NET0131  & \g1246_reg/NET0131  ;
  assign n1614 = n1469 & n1613 ;
  assign n1615 = n818 & n1614 ;
  assign n1616 = ~n1612 & n1615 ;
  assign n1617 = n1612 & ~n1615 ;
  assign n1618 = ~n1616 & ~n1617 ;
  assign n1619 = ~n1610 & n1618 ;
  assign n1620 = \g17316_pad  & ~n1607 ;
  assign n1621 = \g1816_reg/NET0131  & \g35_pad  ;
  assign n1622 = n1600 & n1621 ;
  assign n1623 = ~n1620 & n1622 ;
  assign n1624 = \g1802_reg/NET0131  & ~\g35_pad  ;
  assign n1625 = ~n1623 & ~n1624 ;
  assign n1626 = ~n1619 & n1625 ;
  assign n1627 = ~\g1129_reg/NET0131  & n1469 ;
  assign n1628 = n818 & n1627 ;
  assign n1629 = \g35_pad  & ~n1628 ;
  assign n1630 = n1401 & n1605 ;
  assign n1631 = n1604 & n1630 ;
  assign n1632 = \g17400_pad  & \g35_pad  ;
  assign n1633 = ~n1631 & n1632 ;
  assign n1634 = ~n1629 & ~n1633 ;
  assign n1635 = ~\g1862_reg/NET0131  & ~\g1936_reg/NET0131  ;
  assign n1636 = \g1950_reg/NET0131  & ~n1635 ;
  assign n1637 = ~\g1129_reg/NET0131  & ~\g1246_reg/NET0131  ;
  assign n1638 = n1469 & n1637 ;
  assign n1639 = n818 & n1638 ;
  assign n1640 = ~n1636 & n1639 ;
  assign n1641 = n1636 & ~n1639 ;
  assign n1642 = ~n1640 & ~n1641 ;
  assign n1643 = ~n1634 & n1642 ;
  assign n1644 = \g17400_pad  & ~n1631 ;
  assign n1645 = \g1950_reg/NET0131  & \g35_pad  ;
  assign n1646 = n1628 & n1645 ;
  assign n1647 = ~n1644 & n1646 ;
  assign n1648 = \g1936_reg/NET0131  & ~\g35_pad  ;
  assign n1649 = ~n1647 & ~n1648 ;
  assign n1650 = ~n1643 & n1649 ;
  assign n1651 = ~\g956_reg/NET0131  & n1469 ;
  assign n1652 = n818 & n1651 ;
  assign n1653 = \g35_pad  & ~n1652 ;
  assign n1654 = n1416 & n1605 ;
  assign n1655 = n1604 & n1654 ;
  assign n1656 = \g1087_reg/NET0131  & \g35_pad  ;
  assign n1657 = ~n1655 & n1656 ;
  assign n1658 = ~n1653 & ~n1657 ;
  assign n1659 = ~\g1996_reg/NET0131  & ~\g2070_reg/NET0131  ;
  assign n1660 = \g2084_reg/NET0131  & ~n1659 ;
  assign n1661 = \g1246_reg/NET0131  & ~\g956_reg/NET0131  ;
  assign n1662 = n1469 & n1661 ;
  assign n1663 = n818 & n1662 ;
  assign n1664 = ~n1660 & n1663 ;
  assign n1665 = n1660 & ~n1663 ;
  assign n1666 = ~n1664 & ~n1665 ;
  assign n1667 = ~n1658 & n1666 ;
  assign n1668 = \g1087_reg/NET0131  & ~n1655 ;
  assign n1669 = \g2084_reg/NET0131  & \g35_pad  ;
  assign n1670 = n1652 & n1669 ;
  assign n1671 = ~n1668 & n1670 ;
  assign n1672 = \g2070_reg/NET0131  & ~\g35_pad  ;
  assign n1673 = ~n1671 & ~n1672 ;
  assign n1674 = ~n1667 & n1673 ;
  assign n1675 = ~\g2970_reg/NET0131  & ~\g35_pad  ;
  assign n1676 = ~\g301_reg/NET0131  & \g35_pad  ;
  assign n1677 = ~\g2902_reg/NET0131  & n1469 ;
  assign n1678 = n1676 & n1677 ;
  assign n1679 = ~n1675 & ~n1678 ;
  assign n1680 = \g1339_reg/NET0131  & \g7946_pad  ;
  assign n1681 = n1231 & n1680 ;
  assign n1682 = \g35_pad  & n1681 ;
  assign n1683 = \g1526_reg/NET0131  & n1137 ;
  assign n1684 = \g1306_reg/NET0131  & \g35_pad  ;
  assign n1685 = ~n1683 & n1684 ;
  assign n1686 = ~n1682 & ~n1685 ;
  assign n1687 = \g1521_reg/NET0131  & ~\g35_pad  ;
  assign n1688 = n1686 & ~n1687 ;
  assign n1689 = ~\g2197_reg/NET0131  & ~n1471 ;
  assign n1690 = \g17320_pad  & ~\g2197_reg/NET0131  ;
  assign n1691 = ~n1478 & n1690 ;
  assign n1692 = ~n1689 & ~n1691 ;
  assign n1693 = ~\g1478_reg/NET0131  & ~\g1585_reg/NET0131  ;
  assign n1694 = n1469 & n1693 ;
  assign n1695 = n816 & n1694 ;
  assign n1696 = \g2153_reg/NET0131  & ~n1695 ;
  assign n1697 = ~n1692 & n1696 ;
  assign n1698 = \g35_pad  & n1697 ;
  assign n1699 = \g2153_reg/NET0131  & ~n1692 ;
  assign n1700 = \g2161_reg/NET0131  & \g35_pad  ;
  assign n1701 = ~n1699 & n1700 ;
  assign n1702 = ~n1698 & ~n1701 ;
  assign n1703 = \g2165_reg/NET0131  & ~\g35_pad  ;
  assign n1704 = n1702 & ~n1703 ;
  assign n1705 = ~n1471 & n1482 ;
  assign n1706 = \g17320_pad  & n1482 ;
  assign n1707 = ~n1478 & n1706 ;
  assign n1708 = ~n1705 & ~n1707 ;
  assign n1709 = \g2165_reg/NET0131  & \g35_pad  ;
  assign n1710 = n1708 & n1709 ;
  assign n1711 = \g35_pad  & ~n1695 ;
  assign n1712 = ~n1708 & n1711 ;
  assign n1713 = ~n1710 & ~n1712 ;
  assign n1714 = \g2246_reg/NET0131  & ~\g35_pad  ;
  assign n1715 = n1713 & ~n1714 ;
  assign n1716 = \g2197_reg/NET0131  & ~n1471 ;
  assign n1717 = \g17320_pad  & \g2197_reg/NET0131  ;
  assign n1718 = ~n1478 & n1717 ;
  assign n1719 = ~n1716 & ~n1718 ;
  assign n1720 = ~\g2227_reg/NET0131  & ~n1695 ;
  assign n1721 = ~n1719 & n1720 ;
  assign n1722 = \g35_pad  & n1721 ;
  assign n1723 = ~\g2227_reg/NET0131  & ~n1719 ;
  assign n1724 = \g2169_reg/NET0131  & \g35_pad  ;
  assign n1725 = ~n1723 & n1724 ;
  assign n1726 = ~n1722 & ~n1725 ;
  assign n1727 = \g2161_reg/NET0131  & ~\g35_pad  ;
  assign n1728 = n1726 & ~n1727 ;
  assign n1729 = \g2153_reg/NET0131  & ~n1471 ;
  assign n1730 = \g17320_pad  & \g2153_reg/NET0131  ;
  assign n1731 = ~n1478 & n1730 ;
  assign n1732 = ~n1729 & ~n1731 ;
  assign n1733 = \g2227_reg/NET0131  & ~n1695 ;
  assign n1734 = ~n1732 & n1733 ;
  assign n1735 = \g35_pad  & n1734 ;
  assign n1736 = \g2227_reg/NET0131  & ~n1732 ;
  assign n1737 = \g2173_reg/NET0131  & \g35_pad  ;
  assign n1738 = ~n1736 & n1737 ;
  assign n1739 = ~n1735 & ~n1738 ;
  assign n1740 = \g2177_reg/NET0131  & ~\g35_pad  ;
  assign n1741 = n1739 & ~n1740 ;
  assign n1742 = ~\g2153_reg/NET0131  & ~n1695 ;
  assign n1743 = ~n1719 & n1742 ;
  assign n1744 = \g35_pad  & n1743 ;
  assign n1745 = ~\g2153_reg/NET0131  & ~n1719 ;
  assign n1746 = \g2177_reg/NET0131  & \g35_pad  ;
  assign n1747 = ~n1745 & n1746 ;
  assign n1748 = ~n1744 & ~n1747 ;
  assign n1749 = \g2181_reg/NET0131  & ~\g35_pad  ;
  assign n1750 = n1748 & ~n1749 ;
  assign n1751 = ~n1692 & n1733 ;
  assign n1752 = \g35_pad  & n1751 ;
  assign n1753 = \g2227_reg/NET0131  & ~n1692 ;
  assign n1754 = \g2181_reg/NET0131  & \g35_pad  ;
  assign n1755 = ~n1753 & n1754 ;
  assign n1756 = ~n1752 & ~n1755 ;
  assign n1757 = \g2169_reg/NET0131  & ~\g35_pad  ;
  assign n1758 = n1756 & ~n1757 ;
  assign n1759 = ~\g2331_reg/NET0131  & ~n1499 ;
  assign n1760 = \g17404_pad  & ~\g2331_reg/NET0131  ;
  assign n1761 = ~n1502 & n1760 ;
  assign n1762 = ~n1759 & ~n1761 ;
  assign n1763 = ~\g1448_reg/NET0131  & \g1585_reg/NET0131  ;
  assign n1764 = n1469 & n1763 ;
  assign n1765 = n816 & n1764 ;
  assign n1766 = \g2287_reg/NET0131  & ~n1765 ;
  assign n1767 = ~n1762 & n1766 ;
  assign n1768 = \g35_pad  & n1767 ;
  assign n1769 = \g2287_reg/NET0131  & ~n1762 ;
  assign n1770 = \g2295_reg/NET0131  & \g35_pad  ;
  assign n1771 = ~n1769 & n1770 ;
  assign n1772 = ~n1768 & ~n1771 ;
  assign n1773 = \g2299_reg/NET0131  & ~\g35_pad  ;
  assign n1774 = n1772 & ~n1773 ;
  assign n1775 = ~n1499 & n1506 ;
  assign n1776 = \g17404_pad  & n1506 ;
  assign n1777 = ~n1502 & n1776 ;
  assign n1778 = ~n1775 & ~n1777 ;
  assign n1779 = \g2299_reg/NET0131  & \g35_pad  ;
  assign n1780 = n1778 & n1779 ;
  assign n1781 = \g35_pad  & ~n1765 ;
  assign n1782 = ~n1778 & n1781 ;
  assign n1783 = ~n1780 & ~n1782 ;
  assign n1784 = \g2380_reg/NET0131  & ~\g35_pad  ;
  assign n1785 = n1783 & ~n1784 ;
  assign n1786 = \g2331_reg/NET0131  & ~n1499 ;
  assign n1787 = \g17404_pad  & \g2331_reg/NET0131  ;
  assign n1788 = ~n1502 & n1787 ;
  assign n1789 = ~n1786 & ~n1788 ;
  assign n1790 = ~\g2361_reg/NET0131  & ~n1765 ;
  assign n1791 = ~n1789 & n1790 ;
  assign n1792 = \g35_pad  & n1791 ;
  assign n1793 = ~\g2361_reg/NET0131  & ~n1789 ;
  assign n1794 = \g2303_reg/NET0131  & \g35_pad  ;
  assign n1795 = ~n1793 & n1794 ;
  assign n1796 = ~n1792 & ~n1795 ;
  assign n1797 = \g2295_reg/NET0131  & ~\g35_pad  ;
  assign n1798 = n1796 & ~n1797 ;
  assign n1799 = \g2287_reg/NET0131  & ~n1499 ;
  assign n1800 = \g17404_pad  & \g2287_reg/NET0131  ;
  assign n1801 = ~n1502 & n1800 ;
  assign n1802 = ~n1799 & ~n1801 ;
  assign n1803 = \g2361_reg/NET0131  & ~n1765 ;
  assign n1804 = ~n1802 & n1803 ;
  assign n1805 = \g35_pad  & n1804 ;
  assign n1806 = \g2361_reg/NET0131  & ~n1802 ;
  assign n1807 = \g2307_reg/NET0131  & \g35_pad  ;
  assign n1808 = ~n1806 & n1807 ;
  assign n1809 = ~n1805 & ~n1808 ;
  assign n1810 = \g2311_reg/NET0131  & ~\g35_pad  ;
  assign n1811 = n1809 & ~n1810 ;
  assign n1812 = ~\g2287_reg/NET0131  & ~n1765 ;
  assign n1813 = ~n1789 & n1812 ;
  assign n1814 = \g35_pad  & n1813 ;
  assign n1815 = ~\g2287_reg/NET0131  & ~n1789 ;
  assign n1816 = \g2311_reg/NET0131  & \g35_pad  ;
  assign n1817 = ~n1815 & n1816 ;
  assign n1818 = ~n1814 & ~n1817 ;
  assign n1819 = \g2315_reg/NET0131  & ~\g35_pad  ;
  assign n1820 = n1818 & ~n1819 ;
  assign n1821 = ~n1762 & n1803 ;
  assign n1822 = \g35_pad  & n1821 ;
  assign n1823 = \g2361_reg/NET0131  & ~n1762 ;
  assign n1824 = \g2315_reg/NET0131  & \g35_pad  ;
  assign n1825 = ~n1823 & n1824 ;
  assign n1826 = ~n1822 & ~n1825 ;
  assign n1827 = \g2303_reg/NET0131  & ~\g35_pad  ;
  assign n1828 = n1826 & ~n1827 ;
  assign n1829 = \g1521_reg/NET0131  & ~\g7946_pad  ;
  assign n1830 = ~n1680 & ~n1829 ;
  assign n1831 = \g35_pad  & ~n1830 ;
  assign n1832 = \g1526_reg/NET0131  & ~\g35_pad  ;
  assign n1833 = ~n1831 & ~n1832 ;
  assign n1834 = ~\g2465_reg/NET0131  & ~n1523 ;
  assign n1835 = \g17423_pad  & ~\g2465_reg/NET0131  ;
  assign n1836 = ~n1526 & n1835 ;
  assign n1837 = ~n1834 & ~n1836 ;
  assign n1838 = ~\g1472_reg/NET0131  & ~\g1585_reg/NET0131  ;
  assign n1839 = n1469 & n1838 ;
  assign n1840 = n816 & n1839 ;
  assign n1841 = \g2421_reg/NET0131  & ~n1840 ;
  assign n1842 = ~n1837 & n1841 ;
  assign n1843 = \g35_pad  & n1842 ;
  assign n1844 = \g2421_reg/NET0131  & ~n1837 ;
  assign n1845 = \g2429_reg/NET0131  & \g35_pad  ;
  assign n1846 = ~n1844 & n1845 ;
  assign n1847 = ~n1843 & ~n1846 ;
  assign n1848 = \g2433_reg/NET0131  & ~\g35_pad  ;
  assign n1849 = n1847 & ~n1848 ;
  assign n1850 = ~n1523 & n1530 ;
  assign n1851 = \g17423_pad  & n1530 ;
  assign n1852 = ~n1526 & n1851 ;
  assign n1853 = ~n1850 & ~n1852 ;
  assign n1854 = \g2433_reg/NET0131  & \g35_pad  ;
  assign n1855 = n1853 & n1854 ;
  assign n1856 = \g35_pad  & ~n1840 ;
  assign n1857 = ~n1853 & n1856 ;
  assign n1858 = ~n1855 & ~n1857 ;
  assign n1859 = \g2514_reg/NET0131  & ~\g35_pad  ;
  assign n1860 = n1858 & ~n1859 ;
  assign n1861 = \g2465_reg/NET0131  & ~n1523 ;
  assign n1862 = \g17423_pad  & \g2465_reg/NET0131  ;
  assign n1863 = ~n1526 & n1862 ;
  assign n1864 = ~n1861 & ~n1863 ;
  assign n1865 = ~\g2495_reg/NET0131  & ~n1840 ;
  assign n1866 = ~n1864 & n1865 ;
  assign n1867 = \g35_pad  & n1866 ;
  assign n1868 = ~\g2495_reg/NET0131  & ~n1864 ;
  assign n1869 = \g2437_reg/NET0131  & \g35_pad  ;
  assign n1870 = ~n1868 & n1869 ;
  assign n1871 = ~n1867 & ~n1870 ;
  assign n1872 = \g2429_reg/NET0131  & ~\g35_pad  ;
  assign n1873 = n1871 & ~n1872 ;
  assign n1874 = \g2421_reg/NET0131  & ~n1523 ;
  assign n1875 = \g17423_pad  & \g2421_reg/NET0131  ;
  assign n1876 = ~n1526 & n1875 ;
  assign n1877 = ~n1874 & ~n1876 ;
  assign n1878 = \g2495_reg/NET0131  & ~n1840 ;
  assign n1879 = ~n1877 & n1878 ;
  assign n1880 = \g35_pad  & n1879 ;
  assign n1881 = \g2495_reg/NET0131  & ~n1877 ;
  assign n1882 = \g2441_reg/NET0131  & \g35_pad  ;
  assign n1883 = ~n1881 & n1882 ;
  assign n1884 = ~n1880 & ~n1883 ;
  assign n1885 = \g2445_reg/NET0131  & ~\g35_pad  ;
  assign n1886 = n1884 & ~n1885 ;
  assign n1887 = ~\g2421_reg/NET0131  & ~n1840 ;
  assign n1888 = ~n1864 & n1887 ;
  assign n1889 = \g35_pad  & n1888 ;
  assign n1890 = ~\g2421_reg/NET0131  & ~n1864 ;
  assign n1891 = \g2445_reg/NET0131  & \g35_pad  ;
  assign n1892 = ~n1890 & n1891 ;
  assign n1893 = ~n1889 & ~n1892 ;
  assign n1894 = \g2449_reg/NET0131  & ~\g35_pad  ;
  assign n1895 = n1893 & ~n1894 ;
  assign n1896 = ~n1837 & n1878 ;
  assign n1897 = \g35_pad  & n1896 ;
  assign n1898 = \g2495_reg/NET0131  & ~n1837 ;
  assign n1899 = \g2449_reg/NET0131  & \g35_pad  ;
  assign n1900 = ~n1898 & n1899 ;
  assign n1901 = ~n1897 & ~n1900 ;
  assign n1902 = \g2437_reg/NET0131  & ~\g35_pad  ;
  assign n1903 = n1901 & ~n1902 ;
  assign n1904 = ~\g2599_reg/NET0131  & ~n1547 ;
  assign n1905 = \g1430_reg/NET0131  & ~\g2599_reg/NET0131  ;
  assign n1906 = ~n1550 & n1905 ;
  assign n1907 = ~n1904 & ~n1906 ;
  assign n1908 = ~\g1300_reg/NET0131  & \g1585_reg/NET0131  ;
  assign n1909 = n1469 & n1908 ;
  assign n1910 = n816 & n1909 ;
  assign n1911 = \g2555_reg/NET0131  & ~n1910 ;
  assign n1912 = ~n1907 & n1911 ;
  assign n1913 = \g35_pad  & n1912 ;
  assign n1914 = \g2555_reg/NET0131  & ~n1907 ;
  assign n1915 = \g2563_reg/NET0131  & \g35_pad  ;
  assign n1916 = ~n1914 & n1915 ;
  assign n1917 = ~n1913 & ~n1916 ;
  assign n1918 = \g2567_reg/NET0131  & ~\g35_pad  ;
  assign n1919 = n1917 & ~n1918 ;
  assign n1920 = ~n1547 & n1554 ;
  assign n1921 = \g1430_reg/NET0131  & n1554 ;
  assign n1922 = ~n1550 & n1921 ;
  assign n1923 = ~n1920 & ~n1922 ;
  assign n1924 = \g2567_reg/NET0131  & \g35_pad  ;
  assign n1925 = n1923 & n1924 ;
  assign n1926 = \g35_pad  & ~n1910 ;
  assign n1927 = ~n1923 & n1926 ;
  assign n1928 = ~n1925 & ~n1927 ;
  assign n1929 = \g2648_reg/NET0131  & ~\g35_pad  ;
  assign n1930 = n1928 & ~n1929 ;
  assign n1931 = \g2599_reg/NET0131  & ~n1547 ;
  assign n1932 = \g1430_reg/NET0131  & \g2599_reg/NET0131  ;
  assign n1933 = ~n1550 & n1932 ;
  assign n1934 = ~n1931 & ~n1933 ;
  assign n1935 = ~\g2629_reg/NET0131  & ~n1910 ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1937 = \g35_pad  & n1936 ;
  assign n1938 = ~\g2629_reg/NET0131  & ~n1934 ;
  assign n1939 = \g2571_reg/NET0131  & \g35_pad  ;
  assign n1940 = ~n1938 & n1939 ;
  assign n1941 = ~n1937 & ~n1940 ;
  assign n1942 = \g2563_reg/NET0131  & ~\g35_pad  ;
  assign n1943 = n1941 & ~n1942 ;
  assign n1944 = \g2629_reg/NET0131  & ~n1547 ;
  assign n1945 = \g1430_reg/NET0131  & \g2629_reg/NET0131  ;
  assign n1946 = ~n1550 & n1945 ;
  assign n1947 = ~n1944 & ~n1946 ;
  assign n1948 = n1911 & ~n1947 ;
  assign n1949 = \g35_pad  & n1948 ;
  assign n1950 = \g2555_reg/NET0131  & ~n1947 ;
  assign n1951 = \g2575_reg/NET0131  & \g35_pad  ;
  assign n1952 = ~n1950 & n1951 ;
  assign n1953 = ~n1949 & ~n1952 ;
  assign n1954 = \g2579_reg/NET0131  & ~\g35_pad  ;
  assign n1955 = n1953 & ~n1954 ;
  assign n1956 = ~\g2555_reg/NET0131  & ~n1910 ;
  assign n1957 = ~n1934 & n1956 ;
  assign n1958 = \g35_pad  & n1957 ;
  assign n1959 = ~\g2555_reg/NET0131  & ~n1934 ;
  assign n1960 = \g2579_reg/NET0131  & \g35_pad  ;
  assign n1961 = ~n1959 & n1960 ;
  assign n1962 = ~n1958 & ~n1961 ;
  assign n1963 = \g2583_reg/NET0131  & ~\g35_pad  ;
  assign n1964 = n1962 & ~n1963 ;
  assign n1965 = \g2629_reg/NET0131  & ~n1910 ;
  assign n1966 = ~n1907 & n1965 ;
  assign n1967 = \g35_pad  & n1966 ;
  assign n1968 = \g2629_reg/NET0131  & ~n1907 ;
  assign n1969 = \g2583_reg/NET0131  & \g35_pad  ;
  assign n1970 = ~n1968 & n1969 ;
  assign n1971 = ~n1967 & ~n1970 ;
  assign n1972 = \g2571_reg/NET0131  & ~\g35_pad  ;
  assign n1973 = n1971 & ~n1972 ;
  assign n1974 = ~\g4543_reg/NET0131  & ~n1100 ;
  assign n1975 = \g1395_reg/NET0131  & ~\g35_pad  ;
  assign n1976 = \g12923_pad  & \g1395_reg/NET0131  ;
  assign n1977 = ~n1330 & n1976 ;
  assign n1978 = ~\g1404_reg/NET0131  & ~n1977 ;
  assign n1979 = ~\g1322_reg/NET0131  & \g35_pad  ;
  assign n1980 = \g12923_pad  & \g1404_reg/NET0131  ;
  assign n1981 = \g1395_reg/NET0131  & n1980 ;
  assign n1982 = ~n1330 & n1981 ;
  assign n1983 = n1979 & ~n1982 ;
  assign n1984 = ~n1978 & n1983 ;
  assign n1985 = ~n1975 & ~n1984 ;
  assign n1986 = \g10527_pad  & ~\g17423_pad  ;
  assign n1987 = \g12923_pad  & \g17423_pad  ;
  assign n1988 = ~n1986 & ~n1987 ;
  assign n1989 = \g35_pad  & ~n1988 ;
  assign n1990 = \g1589_reg/NET0131  & ~\g35_pad  ;
  assign n1991 = ~n1989 & ~n1990 ;
  assign n1992 = ~\g35_pad  & ~\g542_reg/NET0131  ;
  assign n1993 = ~\g534_reg/NET0131  & n1676 ;
  assign n1994 = ~n1992 & ~n1993 ;
  assign n1995 = ~\g4495_reg/NET0131  & ~n1100 ;
  assign n1996 = ~\g1404_reg/NET0131  & ~\g35_pad  ;
  assign n1997 = \g12923_pad  & ~\g1395_reg/NET0131  ;
  assign n1998 = ~\g1404_reg/NET0131  & \g19357_pad  ;
  assign n1999 = n1997 & n1998 ;
  assign n2000 = ~n1996 & ~n1999 ;
  assign n2001 = ~\g12923_pad  & \g1404_reg/NET0131  ;
  assign n2002 = \g19357_pad  & \g35_pad  ;
  assign n2003 = n2001 & n2002 ;
  assign n2004 = n2000 & ~n2003 ;
  assign n2005 = n999 & n1003 ;
  assign n2006 = n1005 & ~n2005 ;
  assign n2007 = ~\g807_reg/NET0131  & n1002 ;
  assign n2008 = n999 & n2007 ;
  assign n2009 = \g35_pad  & ~n2008 ;
  assign n2010 = \g794_reg/NET0131  & ~n2009 ;
  assign n2011 = ~n2006 & ~n2010 ;
  assign n2012 = ~\g35_pad  & \g4427_reg/NET0131  ;
  assign n2013 = \g35_pad  & \g4423_reg/NET0131  ;
  assign n2014 = ~n2012 & ~n2013 ;
  assign n2015 = ~\g12923_pad  & ~\g1395_reg/NET0131  ;
  assign n2016 = ~\g1395_reg/NET0131  & ~\g7946_pad  ;
  assign n2017 = n1329 & n2016 ;
  assign n2018 = ~n2015 & ~n2017 ;
  assign n2019 = ~n1977 & n1979 ;
  assign n2020 = n2018 & n2019 ;
  assign n2021 = ~\g8918_pad  & ~\g8919_pad  ;
  assign n2022 = ~\g8920_pad  & n2021 ;
  assign n2023 = ~\g11770_pad  & ~\g8915_pad  ;
  assign n2024 = ~\g8916_pad  & ~\g8917_pad  ;
  assign n2025 = n2023 & n2024 ;
  assign n2026 = n2022 & n2025 ;
  assign n2027 = ~\g4164_reg/NET0131  & \g4253_reg/NET0131  ;
  assign n2028 = ~\g4145_reg/NET0131  & ~\g4253_reg/NET0131  ;
  assign n2029 = ~n2027 & ~n2028 ;
  assign n2030 = ~\g4235_reg/NET0131  & n2029 ;
  assign n2031 = n2026 & n2030 ;
  assign n2032 = \g4235_reg/NET0131  & ~\g8870_pad  ;
  assign n2033 = n2029 & n2032 ;
  assign n2034 = ~\g4235_reg/NET0131  & \g8870_pad  ;
  assign n2035 = n2029 & n2034 ;
  assign n2036 = ~n2033 & ~n2035 ;
  assign n2037 = ~n2031 & n2036 ;
  assign n2038 = \g4235_reg/NET0131  & \g8870_pad  ;
  assign n2039 = ~n2029 & n2038 ;
  assign n2040 = ~\g4235_reg/NET0131  & ~\g8870_pad  ;
  assign n2041 = ~n2029 & n2040 ;
  assign n2042 = ~n2026 & n2041 ;
  assign n2043 = ~n2039 & ~n2042 ;
  assign n2044 = n2037 & n2043 ;
  assign n2045 = \g35_pad  & ~n2044 ;
  assign n2046 = ~\g35_pad  & \g4235_reg/NET0131  ;
  assign n2047 = ~n2045 & ~n2046 ;
  assign n2048 = \g333_reg/NET0131  & ~\g35_pad  ;
  assign n2049 = ~n1592 & ~n2048 ;
  assign n2050 = ~\g1772_reg/NET0131  & ~n1600 ;
  assign n2051 = \g17316_pad  & ~\g1772_reg/NET0131  ;
  assign n2052 = ~n1607 & n2051 ;
  assign n2053 = ~n2050 & ~n2052 ;
  assign n2054 = ~\g1105_reg/NET0131  & \g1242_reg/NET0131  ;
  assign n2055 = n1469 & n2054 ;
  assign n2056 = n818 & n2055 ;
  assign n2057 = \g1728_reg/NET0131  & ~n2056 ;
  assign n2058 = ~n2053 & n2057 ;
  assign n2059 = \g35_pad  & n2058 ;
  assign n2060 = \g1728_reg/NET0131  & ~n2053 ;
  assign n2061 = \g1736_reg/NET0131  & \g35_pad  ;
  assign n2062 = ~n2060 & n2061 ;
  assign n2063 = ~n2059 & ~n2062 ;
  assign n2064 = \g1740_reg/NET0131  & ~\g35_pad  ;
  assign n2065 = n2063 & ~n2064 ;
  assign n2066 = ~n1600 & n1611 ;
  assign n2067 = \g17316_pad  & n1611 ;
  assign n2068 = ~n1607 & n2067 ;
  assign n2069 = ~n2066 & ~n2068 ;
  assign n2070 = \g1740_reg/NET0131  & \g35_pad  ;
  assign n2071 = n2069 & n2070 ;
  assign n2072 = \g35_pad  & ~n2056 ;
  assign n2073 = ~n2069 & n2072 ;
  assign n2074 = ~n2071 & ~n2073 ;
  assign n2075 = \g1821_reg/NET0131  & ~\g35_pad  ;
  assign n2076 = n2074 & ~n2075 ;
  assign n2077 = \g1728_reg/NET0131  & ~n1600 ;
  assign n2078 = \g1728_reg/NET0131  & \g17316_pad  ;
  assign n2079 = ~n1607 & n2078 ;
  assign n2080 = ~n2077 & ~n2079 ;
  assign n2081 = \g1802_reg/NET0131  & ~n2056 ;
  assign n2082 = ~n2080 & n2081 ;
  assign n2083 = \g35_pad  & n2082 ;
  assign n2084 = \g1802_reg/NET0131  & ~n2080 ;
  assign n2085 = \g1748_reg/NET0131  & \g35_pad  ;
  assign n2086 = ~n2084 & n2085 ;
  assign n2087 = ~n2083 & ~n2086 ;
  assign n2088 = \g1752_reg/NET0131  & ~\g35_pad  ;
  assign n2089 = n2087 & ~n2088 ;
  assign n2090 = \g1772_reg/NET0131  & ~n1600 ;
  assign n2091 = \g17316_pad  & \g1772_reg/NET0131  ;
  assign n2092 = ~n1607 & n2091 ;
  assign n2093 = ~n2090 & ~n2092 ;
  assign n2094 = ~\g1802_reg/NET0131  & ~n2056 ;
  assign n2095 = ~n2093 & n2094 ;
  assign n2096 = \g35_pad  & n2095 ;
  assign n2097 = ~\g1802_reg/NET0131  & ~n2093 ;
  assign n2098 = \g1744_reg/NET0131  & \g35_pad  ;
  assign n2099 = ~n2097 & n2098 ;
  assign n2100 = ~n2096 & ~n2099 ;
  assign n2101 = \g1736_reg/NET0131  & ~\g35_pad  ;
  assign n2102 = n2100 & ~n2101 ;
  assign n2103 = ~\g1728_reg/NET0131  & ~n2056 ;
  assign n2104 = ~n2093 & n2103 ;
  assign n2105 = \g35_pad  & n2104 ;
  assign n2106 = ~\g1728_reg/NET0131  & ~n2093 ;
  assign n2107 = \g1752_reg/NET0131  & \g35_pad  ;
  assign n2108 = ~n2106 & n2107 ;
  assign n2109 = ~n2105 & ~n2108 ;
  assign n2110 = \g1756_reg/NET0131  & ~\g35_pad  ;
  assign n2111 = n2109 & ~n2110 ;
  assign n2112 = ~n2053 & n2081 ;
  assign n2113 = \g35_pad  & n2112 ;
  assign n2114 = \g1802_reg/NET0131  & ~n2053 ;
  assign n2115 = \g1756_reg/NET0131  & \g35_pad  ;
  assign n2116 = ~n2114 & n2115 ;
  assign n2117 = ~n2113 & ~n2116 ;
  assign n2118 = \g1744_reg/NET0131  & ~\g35_pad  ;
  assign n2119 = n2117 & ~n2118 ;
  assign n2120 = ~\g1906_reg/NET0131  & ~n1628 ;
  assign n2121 = \g17400_pad  & ~\g1906_reg/NET0131  ;
  assign n2122 = ~n1631 & n2121 ;
  assign n2123 = ~n2120 & ~n2122 ;
  assign n2124 = ~\g1129_reg/NET0131  & ~\g1242_reg/NET0131  ;
  assign n2125 = n1469 & n2124 ;
  assign n2126 = n818 & n2125 ;
  assign n2127 = \g1862_reg/NET0131  & ~n2126 ;
  assign n2128 = ~n2123 & n2127 ;
  assign n2129 = \g35_pad  & n2128 ;
  assign n2130 = \g1862_reg/NET0131  & ~n2123 ;
  assign n2131 = \g1870_reg/NET0131  & \g35_pad  ;
  assign n2132 = ~n2130 & n2131 ;
  assign n2133 = ~n2129 & ~n2132 ;
  assign n2134 = \g1874_reg/NET0131  & ~\g35_pad  ;
  assign n2135 = n2133 & ~n2134 ;
  assign n2136 = ~n1628 & n1635 ;
  assign n2137 = \g17400_pad  & n1635 ;
  assign n2138 = ~n1631 & n2137 ;
  assign n2139 = ~n2136 & ~n2138 ;
  assign n2140 = \g1874_reg/NET0131  & \g35_pad  ;
  assign n2141 = n2139 & n2140 ;
  assign n2142 = \g35_pad  & ~n2126 ;
  assign n2143 = ~n2139 & n2142 ;
  assign n2144 = ~n2141 & ~n2143 ;
  assign n2145 = \g1955_reg/NET0131  & ~\g35_pad  ;
  assign n2146 = n2144 & ~n2145 ;
  assign n2147 = \g1906_reg/NET0131  & ~n1628 ;
  assign n2148 = \g17400_pad  & \g1906_reg/NET0131  ;
  assign n2149 = ~n1631 & n2148 ;
  assign n2150 = ~n2147 & ~n2149 ;
  assign n2151 = ~\g1936_reg/NET0131  & ~n2126 ;
  assign n2152 = ~n2150 & n2151 ;
  assign n2153 = \g35_pad  & n2152 ;
  assign n2154 = ~\g1936_reg/NET0131  & ~n2150 ;
  assign n2155 = \g1878_reg/NET0131  & \g35_pad  ;
  assign n2156 = ~n2154 & n2155 ;
  assign n2157 = ~n2153 & ~n2156 ;
  assign n2158 = \g1870_reg/NET0131  & ~\g35_pad  ;
  assign n2159 = n2157 & ~n2158 ;
  assign n2160 = \g1862_reg/NET0131  & ~n1628 ;
  assign n2161 = \g17400_pad  & \g1862_reg/NET0131  ;
  assign n2162 = ~n1631 & n2161 ;
  assign n2163 = ~n2160 & ~n2162 ;
  assign n2164 = \g1936_reg/NET0131  & ~n2126 ;
  assign n2165 = ~n2163 & n2164 ;
  assign n2166 = \g35_pad  & n2165 ;
  assign n2167 = \g1936_reg/NET0131  & ~n2163 ;
  assign n2168 = \g1882_reg/NET0131  & \g35_pad  ;
  assign n2169 = ~n2167 & n2168 ;
  assign n2170 = ~n2166 & ~n2169 ;
  assign n2171 = \g1886_reg/NET0131  & ~\g35_pad  ;
  assign n2172 = n2170 & ~n2171 ;
  assign n2173 = ~\g1862_reg/NET0131  & ~n2126 ;
  assign n2174 = ~n2150 & n2173 ;
  assign n2175 = \g35_pad  & n2174 ;
  assign n2176 = ~\g1862_reg/NET0131  & ~n2150 ;
  assign n2177 = \g1886_reg/NET0131  & \g35_pad  ;
  assign n2178 = ~n2176 & n2177 ;
  assign n2179 = ~n2175 & ~n2178 ;
  assign n2180 = \g1890_reg/NET0131  & ~\g35_pad  ;
  assign n2181 = n2179 & ~n2180 ;
  assign n2182 = ~n2123 & n2164 ;
  assign n2183 = \g35_pad  & n2182 ;
  assign n2184 = \g1936_reg/NET0131  & ~n2123 ;
  assign n2185 = \g1890_reg/NET0131  & \g35_pad  ;
  assign n2186 = ~n2184 & n2185 ;
  assign n2187 = ~n2183 & ~n2186 ;
  assign n2188 = \g1878_reg/NET0131  & ~\g35_pad  ;
  assign n2189 = n2187 & ~n2188 ;
  assign n2190 = \g1996_reg/NET0131  & ~n1652 ;
  assign n2191 = \g1087_reg/NET0131  & \g1996_reg/NET0131  ;
  assign n2192 = ~n1655 & n2191 ;
  assign n2193 = ~n2190 & ~n2192 ;
  assign n2194 = \g1242_reg/NET0131  & ~\g956_reg/NET0131  ;
  assign n2195 = n1469 & n2194 ;
  assign n2196 = n818 & n2195 ;
  assign n2197 = ~\g2040_reg/NET0131  & ~n2196 ;
  assign n2198 = ~n2193 & n2197 ;
  assign n2199 = \g35_pad  & n2198 ;
  assign n2200 = ~\g2040_reg/NET0131  & ~n2193 ;
  assign n2201 = \g2004_reg/NET0131  & \g35_pad  ;
  assign n2202 = ~n2200 & n2201 ;
  assign n2203 = ~n2199 & ~n2202 ;
  assign n2204 = \g2008_reg/NET0131  & ~\g35_pad  ;
  assign n2205 = n2203 & ~n2204 ;
  assign n2206 = ~n1652 & n1659 ;
  assign n2207 = \g1087_reg/NET0131  & n1659 ;
  assign n2208 = ~n1655 & n2207 ;
  assign n2209 = ~n2206 & ~n2208 ;
  assign n2210 = \g2008_reg/NET0131  & \g35_pad  ;
  assign n2211 = n2209 & n2210 ;
  assign n2212 = \g35_pad  & ~n2196 ;
  assign n2213 = ~n2209 & n2212 ;
  assign n2214 = ~n2211 & ~n2213 ;
  assign n2215 = \g2089_reg/NET0131  & ~\g35_pad  ;
  assign n2216 = n2214 & ~n2215 ;
  assign n2217 = \g2040_reg/NET0131  & ~n1652 ;
  assign n2218 = \g1087_reg/NET0131  & \g2040_reg/NET0131  ;
  assign n2219 = ~n1655 & n2218 ;
  assign n2220 = ~n2217 & ~n2219 ;
  assign n2221 = ~\g2070_reg/NET0131  & ~n2196 ;
  assign n2222 = ~n2220 & n2221 ;
  assign n2223 = \g35_pad  & n2222 ;
  assign n2224 = ~\g2070_reg/NET0131  & ~n2220 ;
  assign n2225 = \g2012_reg/NET0131  & \g35_pad  ;
  assign n2226 = ~n2224 & n2225 ;
  assign n2227 = ~n2223 & ~n2226 ;
  assign n2228 = \g2004_reg/NET0131  & ~\g35_pad  ;
  assign n2229 = n2227 & ~n2228 ;
  assign n2230 = \g2070_reg/NET0131  & ~n2196 ;
  assign n2231 = ~n2193 & n2230 ;
  assign n2232 = \g35_pad  & n2231 ;
  assign n2233 = \g2070_reg/NET0131  & ~n2193 ;
  assign n2234 = \g2016_reg/NET0131  & \g35_pad  ;
  assign n2235 = ~n2233 & n2234 ;
  assign n2236 = ~n2232 & ~n2235 ;
  assign n2237 = \g2020_reg/NET0131  & ~\g35_pad  ;
  assign n2238 = n2236 & ~n2237 ;
  assign n2239 = ~\g1996_reg/NET0131  & ~n2196 ;
  assign n2240 = ~n2220 & n2239 ;
  assign n2241 = \g35_pad  & n2240 ;
  assign n2242 = ~\g1996_reg/NET0131  & ~n2220 ;
  assign n2243 = \g2020_reg/NET0131  & \g35_pad  ;
  assign n2244 = ~n2242 & n2243 ;
  assign n2245 = ~n2241 & ~n2244 ;
  assign n2246 = \g2024_reg/NET0131  & ~\g35_pad  ;
  assign n2247 = n2245 & ~n2246 ;
  assign n2248 = ~\g2040_reg/NET0131  & ~n1652 ;
  assign n2249 = \g1087_reg/NET0131  & ~\g2040_reg/NET0131  ;
  assign n2250 = ~n1655 & n2249 ;
  assign n2251 = ~n2248 & ~n2250 ;
  assign n2252 = n2230 & ~n2251 ;
  assign n2253 = \g35_pad  & n2252 ;
  assign n2254 = \g2070_reg/NET0131  & ~n2251 ;
  assign n2255 = \g2024_reg/NET0131  & \g35_pad  ;
  assign n2256 = ~n2254 & n2255 ;
  assign n2257 = ~n2253 & ~n2256 ;
  assign n2258 = \g2012_reg/NET0131  & ~\g35_pad  ;
  assign n2259 = n2257 & ~n2258 ;
  assign n2260 = ~\g1135_reg/NET0131  & n1469 ;
  assign n2261 = n818 & n2260 ;
  assign n2262 = \g1592_reg/NET0131  & ~n2261 ;
  assign n2263 = n1368 & n1605 ;
  assign n2264 = n1604 & n2263 ;
  assign n2265 = \g1592_reg/NET0131  & \g17291_pad  ;
  assign n2266 = ~n2264 & n2265 ;
  assign n2267 = ~n2262 & ~n2266 ;
  assign n2268 = ~\g1135_reg/NET0131  & ~\g1242_reg/NET0131  ;
  assign n2269 = n1469 & n2268 ;
  assign n2270 = n818 & n2269 ;
  assign n2271 = ~\g1636_reg/NET0131  & ~n2270 ;
  assign n2272 = ~n2267 & n2271 ;
  assign n2273 = \g35_pad  & n2272 ;
  assign n2274 = ~\g1636_reg/NET0131  & ~n2267 ;
  assign n2275 = \g1600_reg/NET0131  & \g35_pad  ;
  assign n2276 = ~n2274 & n2275 ;
  assign n2277 = ~n2273 & ~n2276 ;
  assign n2278 = \g1604_reg/NET0131  & ~\g35_pad  ;
  assign n2279 = n2277 & ~n2278 ;
  assign n2280 = ~\g1592_reg/NET0131  & ~\g1668_reg/NET0131  ;
  assign n2281 = ~n2261 & n2280 ;
  assign n2282 = \g17291_pad  & n2280 ;
  assign n2283 = ~n2264 & n2282 ;
  assign n2284 = ~n2281 & ~n2283 ;
  assign n2285 = \g1604_reg/NET0131  & \g35_pad  ;
  assign n2286 = n2284 & n2285 ;
  assign n2287 = \g35_pad  & ~n2270 ;
  assign n2288 = ~n2284 & n2287 ;
  assign n2289 = ~n2286 & ~n2288 ;
  assign n2290 = \g1687_reg/NET0131  & ~\g35_pad  ;
  assign n2291 = n2289 & ~n2290 ;
  assign n2292 = \g1636_reg/NET0131  & ~n2261 ;
  assign n2293 = \g1636_reg/NET0131  & \g17291_pad  ;
  assign n2294 = ~n2264 & n2293 ;
  assign n2295 = ~n2292 & ~n2294 ;
  assign n2296 = ~\g1668_reg/NET0131  & ~n2270 ;
  assign n2297 = ~n2295 & n2296 ;
  assign n2298 = \g35_pad  & n2297 ;
  assign n2299 = ~\g1668_reg/NET0131  & ~n2295 ;
  assign n2300 = \g1608_reg/NET0131  & \g35_pad  ;
  assign n2301 = ~n2299 & n2300 ;
  assign n2302 = ~n2298 & ~n2301 ;
  assign n2303 = \g1600_reg/NET0131  & ~\g35_pad  ;
  assign n2304 = n2302 & ~n2303 ;
  assign n2305 = \g1668_reg/NET0131  & ~n2270 ;
  assign n2306 = ~n2267 & n2305 ;
  assign n2307 = \g35_pad  & n2306 ;
  assign n2308 = \g1668_reg/NET0131  & ~n2267 ;
  assign n2309 = \g1612_reg/NET0131  & \g35_pad  ;
  assign n2310 = ~n2308 & n2309 ;
  assign n2311 = ~n2307 & ~n2310 ;
  assign n2312 = \g1616_reg/NET0131  & ~\g35_pad  ;
  assign n2313 = n2311 & ~n2312 ;
  assign n2314 = ~\g1592_reg/NET0131  & ~n2270 ;
  assign n2315 = ~n2295 & n2314 ;
  assign n2316 = \g35_pad  & n2315 ;
  assign n2317 = ~\g1592_reg/NET0131  & ~n2295 ;
  assign n2318 = \g1616_reg/NET0131  & \g35_pad  ;
  assign n2319 = ~n2317 & n2318 ;
  assign n2320 = ~n2316 & ~n2319 ;
  assign n2321 = \g1620_reg/NET0131  & ~\g35_pad  ;
  assign n2322 = n2320 & ~n2321 ;
  assign n2323 = n828 & ~n2261 ;
  assign n2324 = \g17291_pad  & n828 ;
  assign n2325 = ~n2264 & n2324 ;
  assign n2326 = ~n2323 & ~n2325 ;
  assign n2327 = \g1620_reg/NET0131  & \g35_pad  ;
  assign n2328 = n2326 & n2327 ;
  assign n2329 = n2287 & ~n2326 ;
  assign n2330 = ~n2328 & ~n2329 ;
  assign n2331 = \g1608_reg/NET0131  & ~\g35_pad  ;
  assign n2332 = n2330 & ~n2331 ;
  assign n2333 = ~\g35_pad  & \g790_reg/NET0131  ;
  assign n2334 = n999 & n1002 ;
  assign n2335 = \g794_reg/NET0131  & ~n976 ;
  assign n2336 = ~n2334 & ~n2335 ;
  assign n2337 = \g35_pad  & ~n2005 ;
  assign n2338 = ~n2336 & n2337 ;
  assign n2339 = ~n2333 & ~n2338 ;
  assign n2340 = \g1585_reg/NET0131  & ~\g35_pad  ;
  assign n2341 = \g12923_pad  & \g35_pad  ;
  assign n2342 = ~n2340 & ~n2341 ;
  assign n2343 = ~\g513_reg/NET0131  & \g518_reg/NET0131  ;
  assign n2344 = \g203_reg/NET0131  & n2343 ;
  assign n2345 = ~\g174_reg/NET0131  & ~\g182_reg/NET0131  ;
  assign n2346 = ~\g168_reg/NET0131  & n2345 ;
  assign n2347 = n2344 & ~n2346 ;
  assign n2348 = \g691_reg/NET0131  & ~n2347 ;
  assign n2349 = n990 & ~n993 ;
  assign n2350 = n975 & n982 ;
  assign n2351 = n2349 & n2350 ;
  assign n2352 = n2348 & ~n2351 ;
  assign n2353 = \g146_reg/NET0131  & \g203_reg/NET0131  ;
  assign n2354 = n2343 & n2353 ;
  assign n2355 = \g164_reg/NET0131  & \g691_reg/NET0131  ;
  assign n2356 = n2354 & n2355 ;
  assign n2357 = ~n2347 & n2356 ;
  assign n2358 = \g150_reg/NET0131  & \g153_reg/NET0131  ;
  assign n2359 = n2357 & n2358 ;
  assign n2360 = ~\g160_reg/NET0131  & n2359 ;
  assign n2361 = n2352 & n2360 ;
  assign n2362 = \g35_pad  & ~n2361 ;
  assign n2363 = \g157_reg/NET0131  & ~n2362 ;
  assign n2364 = \g157_reg/NET0131  & n2359 ;
  assign n2365 = n2352 & n2364 ;
  assign n2366 = \g160_reg/NET0131  & \g35_pad  ;
  assign n2367 = n2348 & n2366 ;
  assign n2368 = ~n2351 & n2367 ;
  assign n2369 = ~n2365 & n2368 ;
  assign n2370 = ~n2363 & ~n2369 ;
  assign n2371 = ~\g232_reg/NET0131  & \g255_reg/NET0131  ;
  assign n2372 = ~\g225_reg/NET0131  & n2371 ;
  assign n2373 = ~\g239_reg/NET0131  & \g262_reg/NET0131  ;
  assign n2374 = ~\g246_reg/NET0131  & \g269_reg/NET0131  ;
  assign n2375 = n2373 & n2374 ;
  assign n2376 = n2372 & n2375 ;
  assign n2377 = ~\g278_reg/NET0131  & \g691_reg/NET0131  ;
  assign n2378 = n2376 & n2377 ;
  assign n2379 = \g246_reg/NET0131  & ~\g269_reg/NET0131  ;
  assign n2380 = \g225_reg/NET0131  & n2379 ;
  assign n2381 = \g239_reg/NET0131  & ~\g262_reg/NET0131  ;
  assign n2382 = \g232_reg/NET0131  & ~\g255_reg/NET0131  ;
  assign n2383 = n2381 & n2382 ;
  assign n2384 = n2380 & n2383 ;
  assign n2385 = \g278_reg/NET0131  & \g691_reg/NET0131  ;
  assign n2386 = n2384 & n2385 ;
  assign n2387 = ~n2378 & ~n2386 ;
  assign n2388 = ~n2351 & ~n2387 ;
  assign n2389 = \g283_reg/NET0131  & \g287_reg/NET0131  ;
  assign n2390 = \g291_reg/NET0131  & n2389 ;
  assign n2391 = \g294_reg/NET0131  & \g298_reg/NET0131  ;
  assign n2392 = n2390 & n2391 ;
  assign n2393 = n2388 & n2392 ;
  assign n2394 = \g142_reg/NET0131  & \g35_pad  ;
  assign n2395 = n2388 & n2394 ;
  assign n2396 = ~n2393 & n2395 ;
  assign n2397 = ~\g142_reg/NET0131  & \g35_pad  ;
  assign n2398 = n2393 & n2397 ;
  assign n2399 = \g298_reg/NET0131  & ~\g35_pad  ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = ~n2396 & n2400 ;
  assign n2402 = ~\g4540_reg/NET0131  & ~n1100 ;
  assign n2403 = \g10500_pad  & ~\g17400_pad  ;
  assign n2404 = \g12919_pad  & \g17400_pad  ;
  assign n2405 = ~n2403 & ~n2404 ;
  assign n2406 = \g35_pad  & ~n2405 ;
  assign n2407 = \g1246_reg/NET0131  & ~\g35_pad  ;
  assign n2408 = ~n2406 & ~n2407 ;
  assign n2409 = \g1052_reg/NET0131  & ~\g35_pad  ;
  assign n2410 = ~\g19334_pad  & ~\g7916_pad  ;
  assign n2411 = ~\g990_reg/NET0131  & n2410 ;
  assign n2412 = \g1052_reg/NET0131  & \g12919_pad  ;
  assign n2413 = ~n2411 & n2412 ;
  assign n2414 = ~\g1061_reg/NET0131  & ~n2413 ;
  assign n2415 = \g35_pad  & ~\g979_reg/NET0131  ;
  assign n2416 = \g1061_reg/NET0131  & n2412 ;
  assign n2417 = ~n2411 & n2416 ;
  assign n2418 = n2415 & ~n2417 ;
  assign n2419 = ~n2414 & n2418 ;
  assign n2420 = ~n2409 & ~n2419 ;
  assign n2421 = \g1579_reg/NET0131  & ~\g35_pad  ;
  assign n2422 = ~n2341 & ~n2421 ;
  assign n2423 = \g781_reg/NET0131  & ~n976 ;
  assign n2424 = ~\g790_reg/NET0131  & n2423 ;
  assign n2425 = n999 & n2424 ;
  assign n2426 = \g35_pad  & ~n2425 ;
  assign n2427 = \g785_reg/NET0131  & ~n2426 ;
  assign n2428 = \g785_reg/NET0131  & n2423 ;
  assign n2429 = n999 & n2428 ;
  assign n2430 = \g35_pad  & \g790_reg/NET0131  ;
  assign n2431 = ~n976 & n2430 ;
  assign n2432 = ~n2429 & n2431 ;
  assign n2433 = ~n2427 & ~n2432 ;
  assign n2434 = \g35_pad  & ~n2365 ;
  assign n2435 = \g160_reg/NET0131  & ~n2434 ;
  assign n2436 = ~\g4480_reg/NET0131  & ~n1100 ;
  assign n2437 = ~\g1061_reg/NET0131  & ~\g35_pad  ;
  assign n2438 = ~\g1052_reg/NET0131  & \g12919_pad  ;
  assign n2439 = ~\g1061_reg/NET0131  & \g19334_pad  ;
  assign n2440 = n2438 & n2439 ;
  assign n2441 = ~n2437 & ~n2440 ;
  assign n2442 = \g1061_reg/NET0131  & ~\g12919_pad  ;
  assign n2443 = \g19334_pad  & \g35_pad  ;
  assign n2444 = n2442 & n2443 ;
  assign n2445 = n2441 & ~n2444 ;
  assign n2446 = ~n2371 & ~n2382 ;
  assign n2447 = \g225_reg/NET0131  & n2446 ;
  assign n2448 = ~\g225_reg/NET0131  & ~n2446 ;
  assign n2449 = ~n2447 & ~n2448 ;
  assign n2450 = ~n2374 & ~n2379 ;
  assign n2451 = n2449 & n2450 ;
  assign n2452 = ~n2449 & ~n2450 ;
  assign n2453 = ~n2451 & ~n2452 ;
  assign n2454 = n971 & n973 ;
  assign n2455 = n982 & n989 ;
  assign n2456 = n2454 & n2455 ;
  assign n2457 = ~n2373 & ~n2381 ;
  assign n2458 = \g732_reg/NET0131  & n2457 ;
  assign n2459 = ~n2456 & n2458 ;
  assign n2460 = ~\g732_reg/NET0131  & ~n2457 ;
  assign n2461 = n2455 & ~n2457 ;
  assign n2462 = n2454 & n2461 ;
  assign n2463 = ~n2460 & ~n2462 ;
  assign n2464 = ~n2459 & n2463 ;
  assign n2465 = n2453 & ~n2464 ;
  assign n2466 = ~n2453 & n2464 ;
  assign n2467 = \g35_pad  & ~n2466 ;
  assign n2468 = ~n2465 & n2467 ;
  assign n2469 = \g153_reg/NET0131  & ~\g35_pad  ;
  assign n2470 = \g150_reg/NET0131  & n2357 ;
  assign n2471 = ~n2351 & n2470 ;
  assign n2472 = ~\g157_reg/NET0131  & \g691_reg/NET0131  ;
  assign n2473 = ~n2347 & n2472 ;
  assign n2474 = \g153_reg/NET0131  & n2473 ;
  assign n2475 = n2471 & n2474 ;
  assign n2476 = ~n2469 & ~n2475 ;
  assign n2477 = \g157_reg/NET0131  & \g35_pad  ;
  assign n2478 = ~n2359 & n2477 ;
  assign n2479 = n2352 & n2478 ;
  assign n2480 = n2476 & ~n2479 ;
  assign n2481 = \g35_pad  & n2429 ;
  assign n2482 = n999 & n2423 ;
  assign n2483 = \g35_pad  & ~n1000 ;
  assign n2484 = ~n2482 & n2483 ;
  assign n2485 = ~n2481 & ~n2484 ;
  assign n2486 = ~\g35_pad  & ~\g781_reg/NET0131  ;
  assign n2487 = n2485 & ~n2486 ;
  assign n2488 = ~\g1052_reg/NET0131  & ~\g12919_pad  ;
  assign n2489 = ~\g1052_reg/NET0131  & ~\g990_reg/NET0131  ;
  assign n2490 = n2410 & n2489 ;
  assign n2491 = ~n2488 & ~n2490 ;
  assign n2492 = ~n2413 & n2415 ;
  assign n2493 = n2491 & n2492 ;
  assign n2494 = \g35_pad  & \g4443_reg/NET0131  ;
  assign n2495 = ~\g4434_reg/NET0131  & ~n2494 ;
  assign n2496 = ~\g4452_reg/NET0131  & ~\g7245_pad  ;
  assign n2497 = ~\g7260_pad  & n2496 ;
  assign n2498 = ~\g4438_reg/NET0131  & ~\g4443_reg/NET0131  ;
  assign n2499 = \g4392_reg/NET0131  & n2498 ;
  assign n2500 = n2497 & n2499 ;
  assign n2501 = \g35_pad  & ~n2494 ;
  assign n2502 = ~n2500 & n2501 ;
  assign n2503 = ~n2495 & ~n2502 ;
  assign n2504 = \g329_reg/NET0131  & ~\g35_pad  ;
  assign n2505 = ~\g305_reg/NET0131  & ~\g311_reg/NET0131  ;
  assign n2506 = ~\g319_reg/NET0131  & ~\g329_reg/NET0131  ;
  assign n2507 = n2505 & n2506 ;
  assign n2508 = \g35_pad  & n2507 ;
  assign n2509 = \g305_reg/NET0131  & \g336_reg/NET0131  ;
  assign n2510 = \g311_reg/NET0131  & ~\g336_reg/NET0131  ;
  assign n2511 = ~\g319_reg/NET0131  & ~n2510 ;
  assign n2512 = ~n2509 & n2511 ;
  assign n2513 = ~\g305_reg/NET0131  & \g324_reg/NET0131  ;
  assign n2514 = ~\g311_reg/NET0131  & ~\g324_reg/NET0131  ;
  assign n2515 = ~n2513 & ~n2514 ;
  assign n2516 = \g35_pad  & n2515 ;
  assign n2517 = ~n2512 & n2516 ;
  assign n2518 = ~n2508 & ~n2517 ;
  assign n2519 = ~n2504 & n2518 ;
  assign n2520 = \g4621_reg/NET0131  & ~\g4639_reg/NET0131  ;
  assign n2521 = \g4628_reg/NET0131  & n2520 ;
  assign n2522 = \g4340_reg/NET0131  & \g4349_reg/NET0131  ;
  assign n2523 = \g4358_reg/NET0131  & n2522 ;
  assign n2524 = n2521 & n2523 ;
  assign n2525 = \g4322_reg/NET0131  & \g4332_reg/NET0131  ;
  assign n2526 = \g4584_reg/NET0131  & \g4593_reg/NET0131  ;
  assign n2527 = n2525 & n2526 ;
  assign n2528 = n2524 & n2527 ;
  assign n2529 = \g4601_reg/NET0131  & \g4608_reg/NET0131  ;
  assign n2530 = n2528 & n2529 ;
  assign n2531 = \g4584_reg/NET0131  & n2525 ;
  assign n2532 = n2524 & n2531 ;
  assign n2533 = \g35_pad  & \g4616_reg/NET0131  ;
  assign n2534 = ~n2532 & n2533 ;
  assign n2535 = ~n2530 & n2534 ;
  assign n2536 = \g4601_reg/NET0131  & ~\g4616_reg/NET0131  ;
  assign n2537 = n2528 & n2536 ;
  assign n2538 = \g35_pad  & ~n2537 ;
  assign n2539 = \g4608_reg/NET0131  & ~n2538 ;
  assign n2540 = ~n2535 & ~n2539 ;
  assign n2541 = \g4401_reg/NET0131  & ~\g4434_reg/NET0131  ;
  assign n2542 = ~\g4401_reg/NET0131  & \g4434_reg/NET0131  ;
  assign n2543 = ~n2541 & ~n2542 ;
  assign n2544 = \g35_pad  & ~n2543 ;
  assign n2545 = \g35_pad  & \g4388_reg/NET0131  ;
  assign n2546 = \g4430_reg/NET0131  & ~n2545 ;
  assign n2547 = ~\g4430_reg/NET0131  & n2545 ;
  assign n2548 = ~n2546 & ~n2547 ;
  assign n2549 = ~n2544 & n2548 ;
  assign n2550 = \g1242_reg/NET0131  & ~\g35_pad  ;
  assign n2551 = \g12919_pad  & \g35_pad  ;
  assign n2552 = ~n2550 & ~n2551 ;
  assign n2553 = \g291_reg/NET0131  & ~\g298_reg/NET0131  ;
  assign n2554 = n2389 & n2553 ;
  assign n2555 = n2388 & n2554 ;
  assign n2556 = \g35_pad  & ~n2555 ;
  assign n2557 = \g294_reg/NET0131  & ~n2556 ;
  assign n2558 = \g291_reg/NET0131  & \g294_reg/NET0131  ;
  assign n2559 = n2389 & n2558 ;
  assign n2560 = n2388 & n2559 ;
  assign n2561 = \g298_reg/NET0131  & \g35_pad  ;
  assign n2562 = n2388 & n2561 ;
  assign n2563 = ~n2560 & n2562 ;
  assign n2564 = ~n2557 & ~n2563 ;
  assign n2565 = ~\g781_reg/NET0131  & n996 ;
  assign n2566 = n995 & n2565 ;
  assign n2567 = n986 & n2566 ;
  assign n2568 = \g35_pad  & ~n2567 ;
  assign n2569 = \g776_reg/NET0131  & ~n2568 ;
  assign n2570 = \g35_pad  & \g781_reg/NET0131  ;
  assign n2571 = ~n976 & n2570 ;
  assign n2572 = ~n999 & n2571 ;
  assign n2573 = ~n2569 & ~n2572 ;
  assign n2574 = ~\g35_pad  & \g4423_reg/NET0131  ;
  assign n2575 = ~\g4372_reg/NET0131  & ~\g4581_reg/NET0131  ;
  assign n2576 = \g35_pad  & ~n2575 ;
  assign n2577 = ~n2574 & ~n2576 ;
  assign n2578 = \g370_reg/NET0131  & \g385_reg/NET0131  ;
  assign n2579 = n982 & n2578 ;
  assign n2580 = \g817_reg/NET0131  & \g832_reg/NET0131  ;
  assign n2581 = \g822_reg/NET0131  & n2580 ;
  assign n2582 = n2579 & n2581 ;
  assign n2583 = \g827_reg/NET0131  & n2582 ;
  assign n2584 = ~\g812_reg/NET0131  & \g837_reg/NET0131  ;
  assign n2585 = \g847_reg/NET0131  & ~n2584 ;
  assign n2586 = \g35_pad  & ~n2585 ;
  assign n2587 = \g723_reg/NET0131  & n2586 ;
  assign n2588 = ~n2583 & n2587 ;
  assign n2589 = ~\g723_reg/NET0131  & ~n2585 ;
  assign n2590 = n2582 & n2589 ;
  assign n2591 = \g35_pad  & ~n2590 ;
  assign n2592 = \g827_reg/NET0131  & ~n2591 ;
  assign n2593 = ~n2588 & ~n2592 ;
  assign n2594 = \g3263_reg/NET0131  & ~\g35_pad  ;
  assign n2595 = ~\g3333_reg/NET0131  & ~\g4674_reg/NET0131  ;
  assign n2596 = ~\g4709_reg/NET0131  & \g4785_reg/NET0131  ;
  assign n2597 = \g4743_reg/NET0131  & n2596 ;
  assign n2598 = ~\g3333_reg/NET0131  & n2597 ;
  assign n2599 = n867 & n2598 ;
  assign n2600 = ~n2595 & ~n2599 ;
  assign n2601 = \g35_pad  & n2600 ;
  assign n2602 = ~n2594 & ~n2601 ;
  assign n2603 = \g3288_reg/NET0131  & ~n900 ;
  assign n2604 = n895 & n2603 ;
  assign n2605 = ~\g3288_reg/NET0131  & ~n913 ;
  assign n2606 = n911 & n2605 ;
  assign n2607 = \g3352_reg/NET0131  & ~n2606 ;
  assign n2608 = ~n2604 & n2607 ;
  assign n2609 = \g3288_reg/NET0131  & ~n928 ;
  assign n2610 = ~n926 & n2609 ;
  assign n2611 = ~n922 & n2610 ;
  assign n2612 = ~\g3288_reg/NET0131  & ~n942 ;
  assign n2613 = ~n940 & n2612 ;
  assign n2614 = ~n936 & n2613 ;
  assign n2615 = ~\g3352_reg/NET0131  & ~n2614 ;
  assign n2616 = ~n2611 & n2615 ;
  assign n2617 = ~n2608 & ~n2616 ;
  assign n2618 = n867 & n2597 ;
  assign n2619 = \g4674_reg/NET0131  & ~n2618 ;
  assign n2620 = ~n2594 & n2619 ;
  assign n2621 = n2617 & n2620 ;
  assign n2622 = ~n2602 & ~n2621 ;
  assign n2623 = ~\g3684_reg/NET0131  & ~\g4681_reg/NET0131  ;
  assign n2624 = \g4709_reg/NET0131  & ~\g4785_reg/NET0131  ;
  assign n2625 = \g4754_reg/NET0131  & n2624 ;
  assign n2626 = ~\g3684_reg/NET0131  & n2625 ;
  assign n2627 = n867 & n2626 ;
  assign n2628 = ~n2623 & ~n2627 ;
  assign n2629 = \g35_pad  & n2628 ;
  assign n2630 = ~n2594 & ~n2629 ;
  assign n2631 = \g3703_reg/NET0131  & ~n900 ;
  assign n2632 = n895 & n2631 ;
  assign n2633 = ~\g3703_reg/NET0131  & ~n928 ;
  assign n2634 = ~n926 & n2633 ;
  assign n2635 = ~n922 & n2634 ;
  assign n2636 = \g3639_reg/NET0131  & ~n2635 ;
  assign n2637 = ~n2632 & n2636 ;
  assign n2638 = \g3703_reg/NET0131  & ~n913 ;
  assign n2639 = n911 & n2638 ;
  assign n2640 = ~\g3703_reg/NET0131  & ~n942 ;
  assign n2641 = ~n940 & n2640 ;
  assign n2642 = ~n936 & n2641 ;
  assign n2643 = ~\g3639_reg/NET0131  & ~n2642 ;
  assign n2644 = ~n2639 & n2643 ;
  assign n2645 = ~n2637 & ~n2644 ;
  assign n2646 = n867 & n2625 ;
  assign n2647 = \g4681_reg/NET0131  & ~n2646 ;
  assign n2648 = ~n2594 & n2647 ;
  assign n2649 = n2645 & n2648 ;
  assign n2650 = ~n2630 & ~n2649 ;
  assign n2651 = ~\g35_pad  & \g4477_reg/NET0131  ;
  assign n2652 = ~n2576 & ~n2651 ;
  assign n2653 = ~\g153_reg/NET0131  & \g164_reg/NET0131  ;
  assign n2654 = n2354 & n2653 ;
  assign n2655 = n2348 & n2654 ;
  assign n2656 = ~n2351 & n2655 ;
  assign n2657 = \g35_pad  & ~n2656 ;
  assign n2658 = \g150_reg/NET0131  & ~n2657 ;
  assign n2659 = \g35_pad  & n2348 ;
  assign n2660 = ~n2351 & n2659 ;
  assign n2661 = \g153_reg/NET0131  & ~n2471 ;
  assign n2662 = n2660 & n2661 ;
  assign n2663 = ~n2658 & ~n2662 ;
  assign n2664 = ~\g776_reg/NET0131  & ~n976 ;
  assign n2665 = n995 & n2664 ;
  assign n2666 = n986 & n2665 ;
  assign n2667 = \g35_pad  & ~n2666 ;
  assign n2668 = \g772_reg/NET0131  & ~n2667 ;
  assign n2669 = n995 & n996 ;
  assign n2670 = n986 & n2669 ;
  assign n2671 = \g35_pad  & \g776_reg/NET0131  ;
  assign n2672 = ~n976 & n2671 ;
  assign n2673 = ~n2670 & n2672 ;
  assign n2674 = ~n2668 & ~n2673 ;
  assign n2675 = \g1236_reg/NET0131  & ~\g35_pad  ;
  assign n2676 = ~n2551 & ~n2675 ;
  assign n2677 = \g1554_reg/NET0131  & ~\g35_pad  ;
  assign n2678 = \g35_pad  & \g496_reg/NET0131  ;
  assign n2679 = ~n2677 & ~n2678 ;
  assign n2680 = ~\g35_pad  & \g4601_reg/NET0131  ;
  assign n2681 = \g4584_reg/NET0131  & \g4616_reg/NET0131  ;
  assign n2682 = n2525 & n2681 ;
  assign n2683 = n2524 & n2682 ;
  assign n2684 = \g35_pad  & ~n2683 ;
  assign n2685 = ~n2530 & n2684 ;
  assign n2686 = \g4601_reg/NET0131  & n2528 ;
  assign n2687 = ~\g4608_reg/NET0131  & ~n2686 ;
  assign n2688 = n2685 & ~n2687 ;
  assign n2689 = ~n2680 & ~n2688 ;
  assign n2690 = ~\g4035_reg/NET0131  & ~\g4688_reg/NET0131  ;
  assign n2691 = ~\g4035_reg/NET0131  & n950 ;
  assign n2692 = n867 & n2691 ;
  assign n2693 = ~n2690 & ~n2692 ;
  assign n2694 = \g35_pad  & n2693 ;
  assign n2695 = ~n2594 & ~n2694 ;
  assign n2696 = \g4688_reg/NET0131  & ~n951 ;
  assign n2697 = ~n2594 & n2696 ;
  assign n2698 = n948 & n2697 ;
  assign n2699 = ~n2695 & ~n2698 ;
  assign n2700 = \g29219_pad  & ~\g35_pad  ;
  assign n2701 = ~\g2748_reg/NET0131  & ~\g2756_reg/NET0131  ;
  assign n2702 = \g2741_reg/NET0131  & n2701 ;
  assign n2703 = \g35_pad  & ~n2702 ;
  assign n2704 = ~n2700 & ~n2703 ;
  assign n2705 = \g2735_reg/NET0131  & \g2741_reg/NET0131  ;
  assign n2706 = \g2748_reg/NET0131  & \g2756_reg/NET0131  ;
  assign n2707 = n2705 & n2706 ;
  assign n2708 = ~\g2193_reg/NET0131  & ~n2701 ;
  assign n2709 = ~n2707 & n2708 ;
  assign n2710 = ~\g2799_reg/NET0131  & ~n2700 ;
  assign n2711 = ~n2709 & n2710 ;
  assign n2712 = ~n2704 & ~n2711 ;
  assign n2713 = ~\g294_reg/NET0131  & n2389 ;
  assign n2714 = n2388 & n2713 ;
  assign n2715 = \g35_pad  & ~n2714 ;
  assign n2716 = \g291_reg/NET0131  & ~n2715 ;
  assign n2717 = n2388 & n2390 ;
  assign n2718 = \g294_reg/NET0131  & \g35_pad  ;
  assign n2719 = n2388 & n2718 ;
  assign n2720 = ~n2717 & n2719 ;
  assign n2721 = ~n2716 & ~n2720 ;
  assign n2722 = \g772_reg/NET0131  & n995 ;
  assign n2723 = n986 & n2722 ;
  assign n2724 = \g35_pad  & n2723 ;
  assign n2725 = n986 & n995 ;
  assign n2726 = \g35_pad  & ~n996 ;
  assign n2727 = ~n2725 & n2726 ;
  assign n2728 = ~n2724 & ~n2727 ;
  assign n2729 = ~\g35_pad  & ~\g767_reg/NET0131  ;
  assign n2730 = n2728 & ~n2729 ;
  assign n2731 = \g29211_pad  & ~\g35_pad  ;
  assign n2732 = \g329_reg/NET0131  & ~\g341_reg/NET0131  ;
  assign n2733 = \g35_pad  & n2732 ;
  assign n2734 = ~n2515 & n2733 ;
  assign n2735 = ~n2731 & ~n2734 ;
  assign n2736 = ~\g35_pad  & \g822_reg/NET0131  ;
  assign n2737 = \g35_pad  & \g827_reg/NET0131  ;
  assign n2738 = ~n2585 & n2737 ;
  assign n2739 = ~n2582 & n2738 ;
  assign n2740 = \g35_pad  & ~\g827_reg/NET0131  ;
  assign n2741 = ~n2585 & n2740 ;
  assign n2742 = n2582 & n2741 ;
  assign n2743 = ~n2739 & ~n2742 ;
  assign n2744 = ~n2736 & n2743 ;
  assign n2745 = \g164_reg/NET0131  & ~\g35_pad  ;
  assign n2746 = ~\g35_pad  & ~n2745 ;
  assign n2747 = \g164_reg/NET0131  & n2354 ;
  assign n2748 = \g150_reg/NET0131  & ~n2747 ;
  assign n2749 = n2348 & n2748 ;
  assign n2750 = ~n2351 & n2749 ;
  assign n2751 = ~\g150_reg/NET0131  & n2357 ;
  assign n2752 = ~n2745 & ~n2751 ;
  assign n2753 = ~n2750 & n2752 ;
  assign n2754 = ~n2746 & ~n2753 ;
  assign n2755 = \g35_pad  & ~\g4674_reg/NET0131  ;
  assign n2756 = \g35_pad  & n2597 ;
  assign n2757 = n867 & n2756 ;
  assign n2758 = ~n2755 & ~n2757 ;
  assign n2759 = \g4749_reg/NET0131  & ~n2758 ;
  assign n2760 = \g35_pad  & \g4674_reg/NET0131  ;
  assign n2761 = ~n2618 & n2760 ;
  assign n2762 = \g4793_reg/NET0131  & n863 ;
  assign n2763 = n861 & n2762 ;
  assign n2764 = \g3343_reg/NET0131  & ~\g3352_reg/NET0131  ;
  assign n2765 = \g3347_reg/NET0131  & \g3352_reg/NET0131  ;
  assign n2766 = ~n2764 & ~n2765 ;
  assign n2767 = ~\g3288_reg/NET0131  & ~\g4749_reg/NET0131  ;
  assign n2768 = ~n2766 & n2767 ;
  assign n2769 = \g3288_reg/NET0131  & ~\g4749_reg/NET0131  ;
  assign n2770 = n2766 & n2769 ;
  assign n2771 = ~n2768 & ~n2770 ;
  assign n2772 = n2763 & n2771 ;
  assign n2773 = n2761 & n2772 ;
  assign n2774 = ~n2759 & ~n2773 ;
  assign n2775 = \g4771_reg/NET0131  & ~n967 ;
  assign n2776 = n2624 & n2762 ;
  assign n2777 = \g3343_reg/NET0131  & ~\g4054_reg/NET0131  ;
  assign n2778 = \g3347_reg/NET0131  & \g4054_reg/NET0131  ;
  assign n2779 = ~n2777 & ~n2778 ;
  assign n2780 = ~\g3990_reg/NET0131  & ~\g4771_reg/NET0131  ;
  assign n2781 = ~n2779 & n2780 ;
  assign n2782 = \g3990_reg/NET0131  & ~\g4771_reg/NET0131  ;
  assign n2783 = n2779 & n2782 ;
  assign n2784 = ~n2781 & ~n2783 ;
  assign n2785 = n2776 & n2784 ;
  assign n2786 = n953 & n2785 ;
  assign n2787 = ~n2775 & ~n2786 ;
  assign n2788 = \g739_reg/NET0131  & ~n976 ;
  assign n2789 = n982 & n2788 ;
  assign n2790 = n975 & n2789 ;
  assign n2791 = n995 & n2790 ;
  assign n2792 = \g744_reg/NET0131  & n978 ;
  assign n2793 = ~\g767_reg/NET0131  & ~n976 ;
  assign n2794 = n2792 & n2793 ;
  assign n2795 = n2791 & n2794 ;
  assign n2796 = \g35_pad  & ~n2795 ;
  assign n2797 = \g763_reg/NET0131  & ~n2796 ;
  assign n2798 = \g744_reg/NET0131  & \g763_reg/NET0131  ;
  assign n2799 = n978 & n2798 ;
  assign n2800 = n2791 & n2799 ;
  assign n2801 = \g35_pad  & \g767_reg/NET0131  ;
  assign n2802 = ~n976 & n2801 ;
  assign n2803 = ~n2800 & n2802 ;
  assign n2804 = ~n2797 & ~n2803 ;
  assign n2805 = ~\g1099_reg/NET0131  & \g13259_pad  ;
  assign n2806 = n1416 & n2805 ;
  assign n2807 = \g35_pad  & n2806 ;
  assign n2808 = \g1152_reg/NET0131  & \g13259_pad  ;
  assign n2809 = n1416 & n2808 ;
  assign n2810 = \g1146_reg/NET0131  & \g35_pad  ;
  assign n2811 = ~n2809 & n2810 ;
  assign n2812 = ~n2807 & ~n2811 ;
  assign n2813 = \g979_reg/NET0131  & ~\g996_reg/NET0131  ;
  assign n2814 = ~\g979_reg/NET0131  & \g996_reg/NET0131  ;
  assign n2815 = ~n2813 & ~n2814 ;
  assign n2816 = ~\g979_reg/NET0131  & ~\g990_reg/NET0131  ;
  assign n2817 = n817 & ~n2816 ;
  assign n2818 = ~n2815 & n2817 ;
  assign n2819 = \g1236_reg/NET0131  & ~\g979_reg/NET0131  ;
  assign n2820 = ~\g1236_reg/NET0131  & \g979_reg/NET0131  ;
  assign n2821 = ~n2819 & ~n2820 ;
  assign n2822 = n2818 & ~n2821 ;
  assign n2823 = \g35_pad  & \g990_reg/NET0131  ;
  assign n2824 = n2822 & n2823 ;
  assign n2825 = ~\g13259_pad  & ~\g8416_pad  ;
  assign n2826 = n2410 & n2825 ;
  assign n2827 = \g35_pad  & ~n2826 ;
  assign n2828 = n2822 & n2827 ;
  assign n2829 = \g35_pad  & ~\g990_reg/NET0131  ;
  assign n2830 = n2826 & n2829 ;
  assign n2831 = ~n2822 & n2830 ;
  assign n2832 = ~n2828 & ~n2831 ;
  assign n2833 = ~n2824 & n2832 ;
  assign n2834 = ~\g35_pad  & \g996_reg/NET0131  ;
  assign n2835 = n2833 & ~n2834 ;
  assign n2836 = ~\g35_pad  & \g4664_reg/NET0131  ;
  assign n2837 = \g4653_reg/NET0131  & \g4688_reg/NET0131  ;
  assign n2838 = n865 & n2837 ;
  assign n2839 = \g35_pad  & ~n2838 ;
  assign n2840 = \g4659_reg/NET0131  & \g4664_reg/NET0131  ;
  assign n2841 = n2837 & n2840 ;
  assign n2842 = ~\g4669_reg/NET0131  & ~n2841 ;
  assign n2843 = n2839 & ~n2842 ;
  assign n2844 = ~n2836 & ~n2843 ;
  assign n2845 = \g287_reg/NET0131  & ~\g35_pad  ;
  assign n2846 = \g283_reg/NET0131  & ~\g291_reg/NET0131  ;
  assign n2847 = \g287_reg/NET0131  & n2846 ;
  assign n2848 = n2388 & n2847 ;
  assign n2849 = ~n2845 & ~n2848 ;
  assign n2850 = \g291_reg/NET0131  & \g35_pad  ;
  assign n2851 = ~n2389 & n2850 ;
  assign n2852 = n2388 & n2851 ;
  assign n2853 = n2849 & ~n2852 ;
  assign n2854 = \g35_pad  & n2800 ;
  assign n2855 = n2791 & n2792 ;
  assign n2856 = \g763_reg/NET0131  & ~n976 ;
  assign n2857 = \g35_pad  & ~n2856 ;
  assign n2858 = ~n2855 & n2857 ;
  assign n2859 = ~n2854 & ~n2858 ;
  assign n2860 = ~\g35_pad  & ~\g758_reg/NET0131  ;
  assign n2861 = n2859 & ~n2860 ;
  assign n2862 = \g35_pad  & \g956_reg/NET0131  ;
  assign n2863 = \g1141_reg/NET0131  & ~\g35_pad  ;
  assign n2864 = \g1099_reg/NET0131  & ~\g1152_reg/NET0131  ;
  assign n2865 = \g1141_reg/NET0131  & n2864 ;
  assign n2866 = n1417 & n2865 ;
  assign n2867 = ~n2863 & ~n2866 ;
  assign n2868 = n2862 & n2867 ;
  assign n2869 = ~n2862 & ~n2867 ;
  assign n2870 = ~n2868 & ~n2869 ;
  assign n2871 = \g1105_reg/NET0131  & \g35_pad  ;
  assign n2872 = \g1111_reg/NET0131  & ~\g35_pad  ;
  assign n2873 = \g1111_reg/NET0131  & n2864 ;
  assign n2874 = n1387 & n2873 ;
  assign n2875 = ~n2872 & ~n2874 ;
  assign n2876 = n2871 & n2875 ;
  assign n2877 = ~n2871 & ~n2875 ;
  assign n2878 = ~n2876 & ~n2877 ;
  assign n2879 = \g1129_reg/NET0131  & \g35_pad  ;
  assign n2880 = \g1124_reg/NET0131  & ~\g35_pad  ;
  assign n2881 = \g1124_reg/NET0131  & n2864 ;
  assign n2882 = n1402 & n2881 ;
  assign n2883 = ~n2880 & ~n2882 ;
  assign n2884 = n2879 & n2883 ;
  assign n2885 = ~n2879 & ~n2883 ;
  assign n2886 = ~n2884 & ~n2885 ;
  assign n2887 = \g1135_reg/NET0131  & \g35_pad  ;
  assign n2888 = \g1094_reg/NET0131  & ~\g35_pad  ;
  assign n2889 = \g1094_reg/NET0131  & n2864 ;
  assign n2890 = n1369 & n2889 ;
  assign n2891 = ~n2888 & ~n2890 ;
  assign n2892 = n2887 & n2891 ;
  assign n2893 = ~n2887 & ~n2891 ;
  assign n2894 = ~n2892 & ~n2893 ;
  assign n2895 = \g35_pad  & ~\g4681_reg/NET0131  ;
  assign n2896 = \g35_pad  & n2625 ;
  assign n2897 = n867 & n2896 ;
  assign n2898 = ~n2895 & ~n2897 ;
  assign n2899 = \g4760_reg/NET0131  & ~n2898 ;
  assign n2900 = \g35_pad  & \g4681_reg/NET0131  ;
  assign n2901 = ~n2646 & n2900 ;
  assign n2902 = n2596 & n2762 ;
  assign n2903 = \g3343_reg/NET0131  & ~\g3703_reg/NET0131  ;
  assign n2904 = \g3347_reg/NET0131  & \g3703_reg/NET0131  ;
  assign n2905 = ~n2903 & ~n2904 ;
  assign n2906 = ~\g3639_reg/NET0131  & ~\g4760_reg/NET0131  ;
  assign n2907 = ~n2905 & n2906 ;
  assign n2908 = \g3639_reg/NET0131  & ~\g4760_reg/NET0131  ;
  assign n2909 = n2905 & n2908 ;
  assign n2910 = ~n2907 & ~n2909 ;
  assign n2911 = n2902 & n2910 ;
  assign n2912 = n2901 & n2911 ;
  assign n2913 = ~n2899 & ~n2912 ;
  assign n2914 = ~\g35_pad  & \g676_reg/NET0131  ;
  assign n2915 = \g482_reg/NET0131  & \g490_reg/NET0131  ;
  assign n2916 = \g499_reg/NET0131  & ~\g504_reg/NET0131  ;
  assign n2917 = ~\g528_reg/NET0131  & n2916 ;
  assign n2918 = n2915 & n2917 ;
  assign n2919 = n2579 & n2918 ;
  assign n2920 = ~n987 & ~n992 ;
  assign n2921 = ~\g661_reg/NET0131  & ~\g728_reg/NET0131  ;
  assign n2922 = \g661_reg/NET0131  & \g728_reg/NET0131  ;
  assign n2923 = ~n2921 & ~n2922 ;
  assign n2924 = ~\g645_reg/NET0131  & ~\g650_reg/NET0131  ;
  assign n2925 = \g681_reg/NET0131  & \g699_reg/NET0131  ;
  assign n2926 = n2924 & n2925 ;
  assign n2927 = ~n2923 & n2926 ;
  assign n2928 = ~n2920 & n2927 ;
  assign n2929 = n2919 & n2928 ;
  assign n2930 = \g35_pad  & \g703_reg/NET0131  ;
  assign n2931 = ~n2929 & n2930 ;
  assign n2932 = \g671_reg/NET0131  & \g676_reg/NET0131  ;
  assign n2933 = n2579 & n2932 ;
  assign n2934 = n2918 & n2933 ;
  assign n2935 = ~\g714_reg/NET0131  & ~n2934 ;
  assign n2936 = \g714_reg/NET0131  & n2934 ;
  assign n2937 = ~n2935 & ~n2936 ;
  assign n2938 = n2931 & n2937 ;
  assign n2939 = ~n2914 & ~n2938 ;
  assign n2940 = ~\g35_pad  & \g4593_reg/NET0131  ;
  assign n2941 = ~n2684 & ~n2940 ;
  assign n2942 = ~\g4601_reg/NET0131  & ~n2940 ;
  assign n2943 = ~n2528 & n2942 ;
  assign n2944 = \g4601_reg/NET0131  & ~n2940 ;
  assign n2945 = n2528 & n2944 ;
  assign n2946 = ~n2943 & ~n2945 ;
  assign n2947 = ~n2941 & n2946 ;
  assign n2948 = \g269_reg/NET0131  & \g35_pad  ;
  assign n2949 = \g29215_pad  & ~\g35_pad  ;
  assign n2950 = ~n2948 & ~n2949 ;
  assign n2951 = \g1146_reg/NET0131  & ~\g35_pad  ;
  assign n2952 = \g1146_reg/NET0131  & \g13259_pad  ;
  assign n2953 = n1416 & n2952 ;
  assign n2954 = ~n2951 & ~n2953 ;
  assign n2955 = \g1152_reg/NET0131  & \g35_pad  ;
  assign n2956 = ~n1417 & n2955 ;
  assign n2957 = n2954 & ~n2956 ;
  assign n2958 = \g29215_pad  & \g35_pad  ;
  assign n2959 = \g1211_reg/NET0131  & ~\g35_pad  ;
  assign n2960 = ~n2958 & ~n2959 ;
  assign n2961 = \g35_pad  & ~n1417 ;
  assign n2962 = ~\g2715_reg/NET0131  & \g2719_reg/NET0131  ;
  assign n2963 = ~\g2724_reg/NET0131  & ~\g2729_reg/NET0131  ;
  assign n2964 = n2962 & ~n2963 ;
  assign n2965 = ~\g2741_reg/NET0131  & ~\g2748_reg/NET0131  ;
  assign n2966 = \g2735_reg/NET0131  & ~\g2756_reg/NET0131  ;
  assign n2967 = n2965 & n2966 ;
  assign n2968 = ~\g2783_reg/NET0131  & n2962 ;
  assign n2969 = n2967 & n2968 ;
  assign n2970 = ~n2964 & ~n2969 ;
  assign n2971 = ~\g1862_reg/NET0131  & \g1906_reg/NET0131  ;
  assign n2972 = \g1917_reg/NET0131  & ~\g1926_reg/NET0131  ;
  assign n2973 = \g35_pad  & n2972 ;
  assign n2974 = ~n2971 & n2973 ;
  assign n2975 = ~n2970 & n2974 ;
  assign n2976 = ~n2970 & n2973 ;
  assign n2977 = ~\g1882_reg/NET0131  & ~\g35_pad  ;
  assign n2978 = ~\g1902_reg/NET0131  & \g35_pad  ;
  assign n2979 = ~n2977 & ~n2978 ;
  assign n2980 = ~n2976 & n2979 ;
  assign n2981 = ~n2975 & ~n2980 ;
  assign n2982 = \g376_reg/NET0131  & \g8719_pad  ;
  assign n2983 = \g385_reg/NET0131  & n2982 ;
  assign n2984 = \g896_reg/NET0131  & n2983 ;
  assign n2985 = \g370_reg/NET0131  & ~\g385_reg/NET0131  ;
  assign n2986 = n2982 & n2985 ;
  assign n2987 = \g392_reg/NET0131  & \g452_reg/NET0131  ;
  assign n2988 = \g174_reg/NET0131  & ~\g392_reg/NET0131  ;
  assign n2989 = ~n2987 & ~n2988 ;
  assign n2990 = ~\g182_reg/NET0131  & n2989 ;
  assign n2991 = \g182_reg/NET0131  & ~n2989 ;
  assign n2992 = ~\g392_reg/NET0131  & \g411_reg/NET0131  ;
  assign n2993 = \g392_reg/NET0131  & \g441_reg/NET0131  ;
  assign n2994 = ~\g417_reg/NET0131  & ~\g691_reg/NET0131  ;
  assign n2995 = ~n2993 & n2994 ;
  assign n2996 = ~n2992 & n2995 ;
  assign n2997 = ~n2991 & n2996 ;
  assign n2998 = ~n2990 & n2997 ;
  assign n2999 = n2986 & n2998 ;
  assign n3000 = ~\g392_reg/NET0131  & ~\g405_reg/NET0131  ;
  assign n3001 = \g392_reg/NET0131  & \g405_reg/NET0131  ;
  assign n3002 = ~n3000 & ~n3001 ;
  assign n3003 = ~\g437_reg/NET0131  & n3002 ;
  assign n3004 = \g392_reg/NET0131  & ~\g401_reg/NET0131  ;
  assign n3005 = ~\g392_reg/NET0131  & ~\g424_reg/NET0131  ;
  assign n3006 = ~n3004 & ~n3005 ;
  assign n3007 = ~n3002 & ~n3006 ;
  assign n3008 = ~n3003 & ~n3007 ;
  assign n3009 = ~\g417_reg/NET0131  & n2986 ;
  assign n3010 = ~n3008 & n3009 ;
  assign n3011 = \g417_reg/NET0131  & n2986 ;
  assign n3012 = n3008 & n3011 ;
  assign n3013 = ~n3010 & ~n3012 ;
  assign n3014 = ~n2999 & n3013 ;
  assign n3015 = ~\g703_reg/NET0131  & \g896_reg/NET0131  ;
  assign n3016 = ~n3014 & n3015 ;
  assign n3017 = ~n2984 & ~n3016 ;
  assign n3018 = \g35_pad  & \g862_reg/NET0131  ;
  assign n3019 = n3017 & n3018 ;
  assign n3020 = ~\g35_pad  & \g446_reg/NET0131  ;
  assign n3021 = \g35_pad  & \g890_reg/NET0131  ;
  assign n3022 = \g896_reg/NET0131  & n3021 ;
  assign n3023 = ~n3020 & ~n3022 ;
  assign n3024 = ~n3019 & n3023 ;
  assign n3025 = ~\g2715_reg/NET0131  & ~\g2719_reg/NET0131  ;
  assign n3026 = ~n2963 & n3025 ;
  assign n3027 = ~\g2803_reg/NET0131  & n3025 ;
  assign n3028 = n2967 & n3027 ;
  assign n3029 = ~n3026 & ~n3028 ;
  assign n3030 = ~\g2153_reg/NET0131  & \g2197_reg/NET0131  ;
  assign n3031 = \g2208_reg/NET0131  & ~\g2217_reg/NET0131  ;
  assign n3032 = \g35_pad  & n3031 ;
  assign n3033 = ~n3030 & n3032 ;
  assign n3034 = ~n3029 & n3033 ;
  assign n3035 = ~n3029 & n3032 ;
  assign n3036 = ~\g2173_reg/NET0131  & ~\g35_pad  ;
  assign n3037 = ~\g2193_reg/NET0131  & \g35_pad  ;
  assign n3038 = ~n3036 & ~n3037 ;
  assign n3039 = ~n3035 & n3038 ;
  assign n3040 = ~n3034 & ~n3039 ;
  assign n3041 = \g2715_reg/NET0131  & ~\g2807_reg/NET0131  ;
  assign n3042 = ~\g2719_reg/NET0131  & n3041 ;
  assign n3043 = n2967 & n3042 ;
  assign n3044 = \g2715_reg/NET0131  & ~\g2719_reg/NET0131  ;
  assign n3045 = ~n2963 & n3044 ;
  assign n3046 = ~n3043 & ~n3045 ;
  assign n3047 = ~\g2287_reg/NET0131  & \g2331_reg/NET0131  ;
  assign n3048 = \g2342_reg/NET0131  & ~\g2351_reg/NET0131  ;
  assign n3049 = \g35_pad  & n3048 ;
  assign n3050 = ~n3047 & n3049 ;
  assign n3051 = ~n3046 & n3050 ;
  assign n3052 = ~\g2307_reg/NET0131  & ~\g35_pad  ;
  assign n3053 = ~\g2327_reg/NET0131  & \g35_pad  ;
  assign n3054 = ~n3052 & ~n3053 ;
  assign n3055 = ~n3049 & n3054 ;
  assign n3056 = ~n3045 & n3054 ;
  assign n3057 = ~n3043 & n3056 ;
  assign n3058 = ~n3055 & ~n3057 ;
  assign n3059 = ~n3051 & n3058 ;
  assign n3060 = \g35_pad  & ~\g4646_reg/NET0131  ;
  assign n3061 = \g35_pad  & n862 ;
  assign n3062 = n867 & n3061 ;
  assign n3063 = ~n3060 & ~n3062 ;
  assign n3064 = \g4704_reg/NET0131  & ~n3063 ;
  assign n3065 = \g35_pad  & \g4646_reg/NET0131  ;
  assign n3066 = ~n868 & n3065 ;
  assign n3067 = n949 & n2762 ;
  assign n3068 = \g3343_reg/NET0131  & ~\g5357_reg/NET0131  ;
  assign n3069 = \g3347_reg/NET0131  & \g5357_reg/NET0131  ;
  assign n3070 = ~n3068 & ~n3069 ;
  assign n3071 = ~\g4704_reg/NET0131  & ~\g5297_reg/NET0131  ;
  assign n3072 = ~n3070 & n3071 ;
  assign n3073 = ~\g4704_reg/NET0131  & \g5297_reg/NET0131  ;
  assign n3074 = n3070 & n3073 ;
  assign n3075 = ~n3072 & ~n3074 ;
  assign n3076 = n3067 & n3075 ;
  assign n3077 = n3066 & n3076 ;
  assign n3078 = ~n3064 & ~n3077 ;
  assign n3079 = ~\g2815_reg/NET0131  & n2962 ;
  assign n3080 = n2967 & n3079 ;
  assign n3081 = ~n2964 & ~n3080 ;
  assign n3082 = ~\g2421_reg/NET0131  & \g2465_reg/NET0131  ;
  assign n3083 = \g2476_reg/NET0131  & ~\g2485_reg/NET0131  ;
  assign n3084 = \g35_pad  & n3083 ;
  assign n3085 = ~n3082 & n3084 ;
  assign n3086 = ~n3081 & n3085 ;
  assign n3087 = ~n3081 & n3084 ;
  assign n3088 = ~\g2441_reg/NET0131  & ~\g35_pad  ;
  assign n3089 = ~\g2461_reg/NET0131  & \g35_pad  ;
  assign n3090 = ~n3088 & ~n3089 ;
  assign n3091 = ~n3087 & n3090 ;
  assign n3092 = ~n3086 & ~n3091 ;
  assign n3093 = ~\g2771_reg/NET0131  & n3025 ;
  assign n3094 = n2967 & n3093 ;
  assign n3095 = ~n3026 & ~n3094 ;
  assign n3096 = ~\g1592_reg/NET0131  & \g1636_reg/NET0131  ;
  assign n3097 = n829 & ~n3096 ;
  assign n3098 = ~n3095 & n3097 ;
  assign n3099 = \g35_pad  & n3098 ;
  assign n3100 = n829 & ~n3095 ;
  assign n3101 = \g1632_reg/NET0131  & \g35_pad  ;
  assign n3102 = ~n3100 & n3101 ;
  assign n3103 = ~n3099 & ~n3102 ;
  assign n3104 = \g1612_reg/NET0131  & ~\g35_pad  ;
  assign n3105 = n3103 & ~n3104 ;
  assign n3106 = \g146_reg/NET0131  & ~\g35_pad  ;
  assign n3107 = ~\g164_reg/NET0131  & ~n2354 ;
  assign n3108 = ~n2747 & ~n3107 ;
  assign n3109 = n2660 & n3108 ;
  assign n3110 = ~n3106 & ~n3109 ;
  assign n3111 = \g744_reg/NET0131  & ~\g758_reg/NET0131  ;
  assign n3112 = n2791 & n3111 ;
  assign n3113 = \g35_pad  & ~n3112 ;
  assign n3114 = \g749_reg/NET0131  & ~n3113 ;
  assign n3115 = \g744_reg/NET0131  & \g749_reg/NET0131  ;
  assign n3116 = n2791 & n3115 ;
  assign n3117 = \g35_pad  & \g758_reg/NET0131  ;
  assign n3118 = ~n976 & n3117 ;
  assign n3119 = ~n3116 & n3118 ;
  assign n3120 = ~n3114 & ~n3119 ;
  assign n3121 = ~\g35_pad  & \g832_reg/NET0131  ;
  assign n3122 = n2579 & n2580 ;
  assign n3123 = ~\g822_reg/NET0131  & ~n3122 ;
  assign n3124 = ~n2582 & n2586 ;
  assign n3125 = ~n3123 & n3124 ;
  assign n3126 = ~n3121 & ~n3125 ;
  assign n3127 = n1355 & n2498 ;
  assign n3128 = n2497 & n3127 ;
  assign n3129 = \g4430_reg/NET0131  & n3128 ;
  assign n3130 = ~\g4452_reg/NET0131  & ~n3129 ;
  assign n3131 = \g2715_reg/NET0131  & \g2719_reg/NET0131  ;
  assign n3132 = ~n2963 & n3131 ;
  assign n3133 = ~\g2819_reg/NET0131  & n3131 ;
  assign n3134 = n2967 & n3133 ;
  assign n3135 = ~n3132 & ~n3134 ;
  assign n3136 = ~\g2587_reg/NET0131  & \g2610_reg/NET0131  ;
  assign n3137 = \g2648_reg/NET0131  & ~\g2652_reg/NET0131  ;
  assign n3138 = ~\g2648_reg/NET0131  & \g2652_reg/NET0131  ;
  assign n3139 = ~n3137 & ~n3138 ;
  assign n3140 = n3136 & ~n3139 ;
  assign n3141 = ~n3135 & n3140 ;
  assign n3142 = \g35_pad  & n3141 ;
  assign n3143 = ~n3135 & n3136 ;
  assign n3144 = \g2657_reg/NET0131  & \g35_pad  ;
  assign n3145 = ~n3143 & n3144 ;
  assign n3146 = ~n3142 & ~n3145 ;
  assign n3147 = \g2652_reg/NET0131  & ~\g35_pad  ;
  assign n3148 = n3146 & ~n3147 ;
  assign n3149 = \g2587_reg/NET0131  & \g2619_reg/NET0131  ;
  assign n3150 = ~n3135 & n3149 ;
  assign n3151 = \g2661_reg/NET0131  & \g35_pad  ;
  assign n3152 = ~n3150 & n3151 ;
  assign n3153 = ~\g2661_reg/NET0131  & \g35_pad  ;
  assign n3154 = n3150 & n3153 ;
  assign n3155 = ~n3152 & ~n3154 ;
  assign n3156 = \g2657_reg/NET0131  & ~\g35_pad  ;
  assign n3157 = n3155 & ~n3156 ;
  assign n3158 = ~\g1624_reg/NET0131  & \g1648_reg/NET0131  ;
  assign n3159 = \g1687_reg/NET0131  & ~\g1691_reg/NET0131  ;
  assign n3160 = ~\g1687_reg/NET0131  & \g1691_reg/NET0131  ;
  assign n3161 = ~n3159 & ~n3160 ;
  assign n3162 = n3158 & ~n3161 ;
  assign n3163 = ~n3095 & n3162 ;
  assign n3164 = \g35_pad  & n3163 ;
  assign n3165 = ~n3095 & n3158 ;
  assign n3166 = \g1696_reg/NET0131  & \g35_pad  ;
  assign n3167 = ~n3165 & n3166 ;
  assign n3168 = ~n3164 & ~n3167 ;
  assign n3169 = \g1691_reg/NET0131  & ~\g35_pad  ;
  assign n3170 = n3168 & ~n3169 ;
  assign n3171 = \g35_pad  & ~n3150 ;
  assign n3172 = \g2587_reg/NET0131  & \g2675_reg/NET0131  ;
  assign n3173 = \g2619_reg/NET0131  & n3172 ;
  assign n3174 = ~n3135 & n3173 ;
  assign n3175 = \g35_pad  & ~n3174 ;
  assign n3176 = ~\g2681_reg/NET0131  & ~n3175 ;
  assign n3177 = ~\g2675_reg/NET0131  & \g2681_reg/NET0131  ;
  assign n3178 = n3149 & n3177 ;
  assign n3179 = ~n3135 & n3178 ;
  assign n3180 = \g35_pad  & n3179 ;
  assign n3181 = ~\g2685_reg/NET0131  & \g35_pad  ;
  assign n3182 = ~n3150 & n3181 ;
  assign n3183 = ~n3180 & ~n3182 ;
  assign n3184 = ~n3176 & n3183 ;
  assign n3185 = \g1624_reg/NET0131  & \g1657_reg/NET0131  ;
  assign n3186 = ~n3095 & n3185 ;
  assign n3187 = \g1700_reg/NET0131  & \g35_pad  ;
  assign n3188 = ~n3186 & n3187 ;
  assign n3189 = ~\g1700_reg/NET0131  & \g35_pad  ;
  assign n3190 = n3186 & n3189 ;
  assign n3191 = ~n3188 & ~n3190 ;
  assign n3192 = \g1696_reg/NET0131  & ~\g35_pad  ;
  assign n3193 = n3191 & ~n3192 ;
  assign n3194 = \g1624_reg/NET0131  & \g1714_reg/NET0131  ;
  assign n3195 = \g1657_reg/NET0131  & n3194 ;
  assign n3196 = ~n3095 & n3195 ;
  assign n3197 = \g35_pad  & ~n3196 ;
  assign n3198 = ~\g1720_reg/NET0131  & ~n3197 ;
  assign n3199 = ~\g1714_reg/NET0131  & \g1720_reg/NET0131  ;
  assign n3200 = n3185 & n3199 ;
  assign n3201 = ~n3095 & n3200 ;
  assign n3202 = \g35_pad  & n3201 ;
  assign n3203 = ~\g1724_reg/NET0131  & \g35_pad  ;
  assign n3204 = ~n3186 & n3203 ;
  assign n3205 = ~n3202 & ~n3204 ;
  assign n3206 = ~n3198 & n3205 ;
  assign n3207 = \g35_pad  & ~n3186 ;
  assign n3208 = \g2715_reg/NET0131  & ~\g2775_reg/NET0131  ;
  assign n3209 = ~\g2719_reg/NET0131  & n3208 ;
  assign n3210 = n2967 & n3209 ;
  assign n3211 = ~n3045 & ~n3210 ;
  assign n3212 = \g1792_reg/NET0131  & ~n3211 ;
  assign n3213 = ~\g1760_reg/NET0131  & \g1783_reg/NET0131  ;
  assign n3214 = ~\g1760_reg/NET0131  & ~n3045 ;
  assign n3215 = ~n3210 & n3214 ;
  assign n3216 = ~n3213 & ~n3215 ;
  assign n3217 = ~n3212 & n3216 ;
  assign n3218 = \g35_pad  & ~n3217 ;
  assign n3219 = ~\g1768_reg/NET0131  & ~\g35_pad  ;
  assign n3220 = ~n3218 & ~n3219 ;
  assign n3221 = \g1821_reg/NET0131  & ~\g1825_reg/NET0131  ;
  assign n3222 = ~\g1821_reg/NET0131  & \g1825_reg/NET0131  ;
  assign n3223 = ~n3221 & ~n3222 ;
  assign n3224 = n3213 & ~n3223 ;
  assign n3225 = ~n3211 & n3224 ;
  assign n3226 = \g35_pad  & n3225 ;
  assign n3227 = ~n3211 & n3213 ;
  assign n3228 = \g1830_reg/NET0131  & \g35_pad  ;
  assign n3229 = ~n3227 & n3228 ;
  assign n3230 = ~n3226 & ~n3229 ;
  assign n3231 = \g1825_reg/NET0131  & ~\g35_pad  ;
  assign n3232 = n3230 & ~n3231 ;
  assign n3233 = \g1760_reg/NET0131  & \g1792_reg/NET0131  ;
  assign n3234 = ~n3211 & n3233 ;
  assign n3235 = \g1834_reg/NET0131  & \g35_pad  ;
  assign n3236 = ~n3234 & n3235 ;
  assign n3237 = ~\g1834_reg/NET0131  & \g35_pad  ;
  assign n3238 = n3234 & n3237 ;
  assign n3239 = ~n3236 & ~n3238 ;
  assign n3240 = \g1830_reg/NET0131  & ~\g35_pad  ;
  assign n3241 = n3239 & ~n3240 ;
  assign n3242 = \g1760_reg/NET0131  & \g1848_reg/NET0131  ;
  assign n3243 = \g1792_reg/NET0131  & n3242 ;
  assign n3244 = ~n3211 & n3243 ;
  assign n3245 = \g35_pad  & ~n3244 ;
  assign n3246 = ~\g1854_reg/NET0131  & ~n3245 ;
  assign n3247 = ~\g1848_reg/NET0131  & \g1854_reg/NET0131  ;
  assign n3248 = n3233 & n3247 ;
  assign n3249 = ~n3211 & n3248 ;
  assign n3250 = \g35_pad  & n3249 ;
  assign n3251 = ~\g1858_reg/NET0131  & \g35_pad  ;
  assign n3252 = ~n3234 & n3251 ;
  assign n3253 = ~n3250 & ~n3252 ;
  assign n3254 = ~n3246 & n3253 ;
  assign n3255 = \g35_pad  & ~n3234 ;
  assign n3256 = \g1926_reg/NET0131  & ~n2970 ;
  assign n3257 = \g35_pad  & n3256 ;
  assign n3258 = ~\g1917_reg/NET0131  & ~n2970 ;
  assign n3259 = ~\g1894_reg/NET0131  & \g35_pad  ;
  assign n3260 = ~n3258 & n3259 ;
  assign n3261 = ~n3257 & ~n3260 ;
  assign n3262 = ~\g1902_reg/NET0131  & ~\g35_pad  ;
  assign n3263 = n3261 & ~n3262 ;
  assign n3264 = ~\g1894_reg/NET0131  & \g1917_reg/NET0131  ;
  assign n3265 = \g1955_reg/NET0131  & ~\g1959_reg/NET0131  ;
  assign n3266 = ~\g1955_reg/NET0131  & \g1959_reg/NET0131  ;
  assign n3267 = ~n3265 & ~n3266 ;
  assign n3268 = n3264 & ~n3267 ;
  assign n3269 = ~n2970 & n3268 ;
  assign n3270 = \g35_pad  & n3269 ;
  assign n3271 = ~n2970 & n3264 ;
  assign n3272 = \g1964_reg/NET0131  & \g35_pad  ;
  assign n3273 = ~n3271 & n3272 ;
  assign n3274 = ~n3270 & ~n3273 ;
  assign n3275 = \g1959_reg/NET0131  & ~\g35_pad  ;
  assign n3276 = n3274 & ~n3275 ;
  assign n3277 = \g1894_reg/NET0131  & \g1926_reg/NET0131  ;
  assign n3278 = ~n2970 & n3277 ;
  assign n3279 = \g1968_reg/NET0131  & \g35_pad  ;
  assign n3280 = ~n3278 & n3279 ;
  assign n3281 = ~\g1968_reg/NET0131  & \g35_pad  ;
  assign n3282 = n3278 & n3281 ;
  assign n3283 = ~n3280 & ~n3282 ;
  assign n3284 = \g1964_reg/NET0131  & ~\g35_pad  ;
  assign n3285 = n3283 & ~n3284 ;
  assign n3286 = \g35_pad  & ~n3278 ;
  assign n3287 = \g1894_reg/NET0131  & \g1982_reg/NET0131  ;
  assign n3288 = \g1926_reg/NET0131  & n3287 ;
  assign n3289 = ~n2970 & n3288 ;
  assign n3290 = \g35_pad  & ~n3289 ;
  assign n3291 = ~\g1988_reg/NET0131  & ~n3290 ;
  assign n3292 = ~\g1982_reg/NET0131  & \g1988_reg/NET0131  ;
  assign n3293 = n3277 & n3292 ;
  assign n3294 = ~n2970 & n3293 ;
  assign n3295 = \g35_pad  & n3294 ;
  assign n3296 = ~\g1992_reg/NET0131  & \g35_pad  ;
  assign n3297 = ~n3278 & n3296 ;
  assign n3298 = ~n3295 & ~n3297 ;
  assign n3299 = ~n3291 & n3298 ;
  assign n3300 = ~\g2787_reg/NET0131  & n3131 ;
  assign n3301 = n2967 & n3300 ;
  assign n3302 = ~n3132 & ~n3301 ;
  assign n3303 = ~\g2028_reg/NET0131  & \g2051_reg/NET0131  ;
  assign n3304 = \g2089_reg/NET0131  & ~\g2093_reg/NET0131  ;
  assign n3305 = ~\g2089_reg/NET0131  & \g2093_reg/NET0131  ;
  assign n3306 = ~n3304 & ~n3305 ;
  assign n3307 = n3303 & ~n3306 ;
  assign n3308 = ~n3302 & n3307 ;
  assign n3309 = \g35_pad  & n3308 ;
  assign n3310 = ~n3302 & n3303 ;
  assign n3311 = \g2098_reg/NET0131  & \g35_pad  ;
  assign n3312 = ~n3310 & n3311 ;
  assign n3313 = ~n3309 & ~n3312 ;
  assign n3314 = \g2093_reg/NET0131  & ~\g35_pad  ;
  assign n3315 = n3313 & ~n3314 ;
  assign n3316 = \g2028_reg/NET0131  & \g2060_reg/NET0131  ;
  assign n3317 = ~n3302 & n3316 ;
  assign n3318 = \g2102_reg/NET0131  & \g35_pad  ;
  assign n3319 = ~n3317 & n3318 ;
  assign n3320 = ~\g2102_reg/NET0131  & \g35_pad  ;
  assign n3321 = n3317 & n3320 ;
  assign n3322 = ~n3319 & ~n3321 ;
  assign n3323 = \g2098_reg/NET0131  & ~\g35_pad  ;
  assign n3324 = n3322 & ~n3323 ;
  assign n3325 = \g35_pad  & ~n3317 ;
  assign n3326 = \g2028_reg/NET0131  & \g2116_reg/NET0131  ;
  assign n3327 = \g2060_reg/NET0131  & n3326 ;
  assign n3328 = ~n3302 & n3327 ;
  assign n3329 = \g35_pad  & ~n3328 ;
  assign n3330 = ~\g2122_reg/NET0131  & ~n3329 ;
  assign n3331 = ~\g2116_reg/NET0131  & \g2122_reg/NET0131  ;
  assign n3332 = n3316 & n3331 ;
  assign n3333 = ~n3302 & n3332 ;
  assign n3334 = \g35_pad  & n3333 ;
  assign n3335 = ~\g2126_reg/NET0131  & \g35_pad  ;
  assign n3336 = ~n3317 & n3335 ;
  assign n3337 = ~n3334 & ~n3336 ;
  assign n3338 = ~n3330 & n3337 ;
  assign n3339 = ~\g2185_reg/NET0131  & \g2208_reg/NET0131  ;
  assign n3340 = \g2246_reg/NET0131  & ~\g2250_reg/NET0131  ;
  assign n3341 = ~\g2246_reg/NET0131  & \g2250_reg/NET0131  ;
  assign n3342 = ~n3340 & ~n3341 ;
  assign n3343 = n3339 & ~n3342 ;
  assign n3344 = ~n3029 & n3343 ;
  assign n3345 = \g35_pad  & n3344 ;
  assign n3346 = ~n3029 & n3339 ;
  assign n3347 = \g2255_reg/NET0131  & \g35_pad  ;
  assign n3348 = ~n3346 & n3347 ;
  assign n3349 = ~n3345 & ~n3348 ;
  assign n3350 = \g2250_reg/NET0131  & ~\g35_pad  ;
  assign n3351 = n3349 & ~n3350 ;
  assign n3352 = \g2185_reg/NET0131  & \g2217_reg/NET0131  ;
  assign n3353 = ~n3029 & n3352 ;
  assign n3354 = \g2259_reg/NET0131  & \g35_pad  ;
  assign n3355 = ~n3353 & n3354 ;
  assign n3356 = ~\g2259_reg/NET0131  & \g35_pad  ;
  assign n3357 = n3353 & n3356 ;
  assign n3358 = ~n3355 & ~n3357 ;
  assign n3359 = \g2255_reg/NET0131  & ~\g35_pad  ;
  assign n3360 = n3358 & ~n3359 ;
  assign n3361 = \g35_pad  & ~n3353 ;
  assign n3362 = \g2185_reg/NET0131  & \g2273_reg/NET0131  ;
  assign n3363 = \g2217_reg/NET0131  & n3362 ;
  assign n3364 = ~n3029 & n3363 ;
  assign n3365 = \g35_pad  & ~n3364 ;
  assign n3366 = ~\g2279_reg/NET0131  & ~n3365 ;
  assign n3367 = ~\g2273_reg/NET0131  & \g2279_reg/NET0131  ;
  assign n3368 = n3352 & n3367 ;
  assign n3369 = ~n3029 & n3368 ;
  assign n3370 = \g35_pad  & n3369 ;
  assign n3371 = ~\g2283_reg/NET0131  & \g35_pad  ;
  assign n3372 = ~n3353 & n3371 ;
  assign n3373 = ~n3370 & ~n3372 ;
  assign n3374 = ~n3366 & n3373 ;
  assign n3375 = \g2351_reg/NET0131  & ~n3046 ;
  assign n3376 = ~\g2319_reg/NET0131  & \g2342_reg/NET0131  ;
  assign n3377 = ~\g2319_reg/NET0131  & ~n3045 ;
  assign n3378 = ~n3043 & n3377 ;
  assign n3379 = ~n3376 & ~n3378 ;
  assign n3380 = ~n3375 & n3379 ;
  assign n3381 = \g35_pad  & ~n3380 ;
  assign n3382 = ~\g2327_reg/NET0131  & ~\g35_pad  ;
  assign n3383 = ~n3381 & ~n3382 ;
  assign n3384 = \g2380_reg/NET0131  & ~\g2384_reg/NET0131  ;
  assign n3385 = ~\g2380_reg/NET0131  & \g2384_reg/NET0131  ;
  assign n3386 = ~n3384 & ~n3385 ;
  assign n3387 = n3376 & ~n3386 ;
  assign n3388 = ~n3046 & n3387 ;
  assign n3389 = \g2389_reg/NET0131  & ~n3376 ;
  assign n3390 = \g2389_reg/NET0131  & ~n3045 ;
  assign n3391 = ~n3043 & n3390 ;
  assign n3392 = ~n3389 & ~n3391 ;
  assign n3393 = ~n3388 & n3392 ;
  assign n3394 = \g35_pad  & ~n3393 ;
  assign n3395 = \g2384_reg/NET0131  & ~\g35_pad  ;
  assign n3396 = ~n3394 & ~n3395 ;
  assign n3397 = \g2319_reg/NET0131  & \g2351_reg/NET0131  ;
  assign n3398 = ~n3046 & n3397 ;
  assign n3399 = \g2393_reg/NET0131  & \g35_pad  ;
  assign n3400 = ~n3398 & n3399 ;
  assign n3401 = ~\g2393_reg/NET0131  & \g35_pad  ;
  assign n3402 = n3398 & n3401 ;
  assign n3403 = ~n3400 & ~n3402 ;
  assign n3404 = \g2389_reg/NET0131  & ~\g35_pad  ;
  assign n3405 = n3403 & ~n3404 ;
  assign n3406 = \g35_pad  & ~n3398 ;
  assign n3407 = \g2319_reg/NET0131  & \g2407_reg/NET0131  ;
  assign n3408 = \g2351_reg/NET0131  & n3407 ;
  assign n3409 = ~n3046 & n3408 ;
  assign n3410 = \g35_pad  & ~n3409 ;
  assign n3411 = ~\g2413_reg/NET0131  & ~n3410 ;
  assign n3412 = ~\g2407_reg/NET0131  & \g2413_reg/NET0131  ;
  assign n3413 = n3397 & n3412 ;
  assign n3414 = ~n3046 & n3413 ;
  assign n3415 = \g35_pad  & n3414 ;
  assign n3416 = ~\g2417_reg/NET0131  & \g35_pad  ;
  assign n3417 = ~n3398 & n3416 ;
  assign n3418 = ~n3415 & ~n3417 ;
  assign n3419 = ~n3411 & n3418 ;
  assign n3420 = \g2485_reg/NET0131  & ~n3081 ;
  assign n3421 = \g35_pad  & n3420 ;
  assign n3422 = ~\g2476_reg/NET0131  & ~n3081 ;
  assign n3423 = ~\g2453_reg/NET0131  & \g35_pad  ;
  assign n3424 = ~n3422 & n3423 ;
  assign n3425 = ~n3421 & ~n3424 ;
  assign n3426 = ~\g2461_reg/NET0131  & ~\g35_pad  ;
  assign n3427 = n3425 & ~n3426 ;
  assign n3428 = ~\g2453_reg/NET0131  & \g2476_reg/NET0131  ;
  assign n3429 = \g2514_reg/NET0131  & ~\g2518_reg/NET0131  ;
  assign n3430 = ~\g2514_reg/NET0131  & \g2518_reg/NET0131  ;
  assign n3431 = ~n3429 & ~n3430 ;
  assign n3432 = n3428 & ~n3431 ;
  assign n3433 = ~n3081 & n3432 ;
  assign n3434 = \g35_pad  & n3433 ;
  assign n3435 = ~n3081 & n3428 ;
  assign n3436 = \g2523_reg/NET0131  & \g35_pad  ;
  assign n3437 = ~n3435 & n3436 ;
  assign n3438 = ~n3434 & ~n3437 ;
  assign n3439 = \g2518_reg/NET0131  & ~\g35_pad  ;
  assign n3440 = n3438 & ~n3439 ;
  assign n3441 = \g2453_reg/NET0131  & \g2485_reg/NET0131  ;
  assign n3442 = ~n3081 & n3441 ;
  assign n3443 = \g2527_reg/NET0131  & \g35_pad  ;
  assign n3444 = ~n3442 & n3443 ;
  assign n3445 = ~\g2527_reg/NET0131  & \g35_pad  ;
  assign n3446 = n3442 & n3445 ;
  assign n3447 = ~n3444 & ~n3446 ;
  assign n3448 = \g2523_reg/NET0131  & ~\g35_pad  ;
  assign n3449 = n3447 & ~n3448 ;
  assign n3450 = \g35_pad  & ~n3442 ;
  assign n3451 = \g2453_reg/NET0131  & \g2541_reg/NET0131  ;
  assign n3452 = \g2485_reg/NET0131  & n3451 ;
  assign n3453 = ~n3081 & n3452 ;
  assign n3454 = \g35_pad  & ~n3453 ;
  assign n3455 = ~\g2547_reg/NET0131  & ~n3454 ;
  assign n3456 = ~\g2541_reg/NET0131  & \g2547_reg/NET0131  ;
  assign n3457 = n3441 & n3456 ;
  assign n3458 = ~n3081 & n3457 ;
  assign n3459 = \g35_pad  & n3458 ;
  assign n3460 = ~\g2551_reg/NET0131  & \g35_pad  ;
  assign n3461 = ~n3442 & n3460 ;
  assign n3462 = ~n3459 & ~n3461 ;
  assign n3463 = ~n3455 & n3462 ;
  assign n3464 = \g2060_reg/NET0131  & ~n3302 ;
  assign n3465 = \g35_pad  & n3464 ;
  assign n3466 = ~\g2051_reg/NET0131  & ~n3302 ;
  assign n3467 = ~\g2028_reg/NET0131  & \g35_pad  ;
  assign n3468 = ~n3466 & n3467 ;
  assign n3469 = ~n3465 & ~n3468 ;
  assign n3470 = ~\g2036_reg/NET0131  & ~\g35_pad  ;
  assign n3471 = n3469 & ~n3470 ;
  assign n3472 = \g2217_reg/NET0131  & ~n3029 ;
  assign n3473 = \g35_pad  & n3472 ;
  assign n3474 = ~\g2208_reg/NET0131  & ~n3029 ;
  assign n3475 = ~\g2185_reg/NET0131  & \g35_pad  ;
  assign n3476 = ~n3474 & n3475 ;
  assign n3477 = ~n3473 & ~n3476 ;
  assign n3478 = ~\g2193_reg/NET0131  & ~\g35_pad  ;
  assign n3479 = n3477 & ~n3478 ;
  assign n3480 = \g1657_reg/NET0131  & ~n3095 ;
  assign n3481 = \g35_pad  & n3480 ;
  assign n3482 = ~\g1648_reg/NET0131  & ~n3095 ;
  assign n3483 = ~\g1624_reg/NET0131  & \g35_pad  ;
  assign n3484 = ~n3482 & n3483 ;
  assign n3485 = ~n3481 & ~n3484 ;
  assign n3486 = ~\g1632_reg/NET0131  & ~\g35_pad  ;
  assign n3487 = n3485 & ~n3486 ;
  assign n3488 = \g2619_reg/NET0131  & ~n3135 ;
  assign n3489 = \g35_pad  & n3488 ;
  assign n3490 = ~\g2610_reg/NET0131  & ~n3135 ;
  assign n3491 = ~\g2587_reg/NET0131  & \g35_pad  ;
  assign n3492 = ~n3490 & n3491 ;
  assign n3493 = ~n3489 & ~n3492 ;
  assign n3494 = ~\g2595_reg/NET0131  & ~\g35_pad  ;
  assign n3495 = n3493 & ~n3494 ;
  assign n3496 = \g4438_reg/NET0131  & ~n1441 ;
  assign n3497 = n1443 & n2498 ;
  assign n3498 = n2497 & n3497 ;
  assign n3499 = ~n3496 & ~n3498 ;
  assign n3500 = \g35_pad  & ~\g5084_reg/NET0131  ;
  assign n3501 = \g5080_reg/NET0131  & ~n3500 ;
  assign n3502 = ~\g5073_reg/NET0131  & \g5077_reg/NET0131  ;
  assign n3503 = ~\g5069_reg/NET0131  & \g5077_reg/NET0131  ;
  assign n3504 = ~\g5080_reg/NET0131  & ~\g5084_reg/NET0131  ;
  assign n3505 = ~n3503 & n3504 ;
  assign n3506 = ~n3502 & ~n3505 ;
  assign n3507 = \g35_pad  & ~n3506 ;
  assign n3508 = ~n3501 & ~n3507 ;
  assign n3509 = \g2831_reg/NET0131  & ~\g35_pad  ;
  assign n3510 = ~\g2715_reg/NET0131  & ~\g2783_reg/NET0131  ;
  assign n3511 = \g2715_reg/NET0131  & ~\g2787_reg/NET0131  ;
  assign n3512 = \g2719_reg/NET0131  & ~n3511 ;
  assign n3513 = ~n3510 & n3512 ;
  assign n3514 = ~\g2715_reg/NET0131  & ~\g2771_reg/NET0131  ;
  assign n3515 = ~\g2719_reg/NET0131  & ~n3208 ;
  assign n3516 = ~n3514 & n3515 ;
  assign n3517 = ~n3513 & ~n3516 ;
  assign n3518 = ~\g2756_reg/NET0131  & n2965 ;
  assign n3519 = ~\g2735_reg/NET0131  & n2963 ;
  assign n3520 = n3518 & n3519 ;
  assign n3521 = \g35_pad  & n3520 ;
  assign n3522 = n3517 & n3521 ;
  assign n3523 = \g2079_reg/NET0131  & \g2715_reg/NET0131  ;
  assign n3524 = \g1945_reg/NET0131  & ~\g2715_reg/NET0131  ;
  assign n3525 = \g2719_reg/NET0131  & ~n3524 ;
  assign n3526 = ~n3523 & n3525 ;
  assign n3527 = \g1811_reg/NET0131  & \g2715_reg/NET0131  ;
  assign n3528 = \g1677_reg/NET0131  & ~\g2715_reg/NET0131  ;
  assign n3529 = ~\g2719_reg/NET0131  & ~n3528 ;
  assign n3530 = ~n3527 & n3529 ;
  assign n3531 = ~n3526 & ~n3530 ;
  assign n3532 = \g35_pad  & ~n3520 ;
  assign n3533 = n3531 & n3532 ;
  assign n3534 = ~n3522 & ~n3533 ;
  assign n3535 = ~n3509 & n3534 ;
  assign n3536 = \g35_pad  & ~n2388 ;
  assign n3537 = \g35_pad  & n2389 ;
  assign n3538 = ~\g283_reg/NET0131  & ~\g35_pad  ;
  assign n3539 = ~\g283_reg/NET0131  & ~\g287_reg/NET0131  ;
  assign n3540 = ~n3538 & ~n3539 ;
  assign n3541 = ~n3537 & n3540 ;
  assign n3542 = ~n3536 & n3541 ;
  assign n3543 = ~\g1792_reg/NET0131  & \g35_pad  ;
  assign n3544 = ~\g1728_reg/NET0131  & \g1772_reg/NET0131  ;
  assign n3545 = \g1783_reg/NET0131  & ~n3544 ;
  assign n3546 = n3543 & n3545 ;
  assign n3547 = ~n3211 & n3546 ;
  assign n3548 = \g1783_reg/NET0131  & n3543 ;
  assign n3549 = ~n3211 & n3548 ;
  assign n3550 = ~\g1748_reg/NET0131  & ~\g35_pad  ;
  assign n3551 = ~\g1768_reg/NET0131  & \g35_pad  ;
  assign n3552 = ~n3550 & ~n3551 ;
  assign n3553 = ~n3549 & n3552 ;
  assign n3554 = ~n3547 & ~n3553 ;
  assign n3555 = ~\g35_pad  & \g744_reg/NET0131  ;
  assign n3556 = \g744_reg/NET0131  & ~\g749_reg/NET0131  ;
  assign n3557 = n2791 & n3556 ;
  assign n3558 = ~n3555 & ~n3557 ;
  assign n3559 = \g744_reg/NET0131  & n2791 ;
  assign n3560 = \g749_reg/NET0131  & ~n976 ;
  assign n3561 = \g35_pad  & n3560 ;
  assign n3562 = ~n3559 & n3561 ;
  assign n3563 = n3558 & ~n3562 ;
  assign n3564 = \g2051_reg/NET0131  & ~\g2060_reg/NET0131  ;
  assign n3565 = ~\g1996_reg/NET0131  & \g2040_reg/NET0131  ;
  assign n3566 = n3564 & n3565 ;
  assign n3567 = ~n3302 & n3566 ;
  assign n3568 = \g35_pad  & n3567 ;
  assign n3569 = ~n3302 & n3564 ;
  assign n3570 = ~\g2036_reg/NET0131  & \g35_pad  ;
  assign n3571 = ~n3569 & n3570 ;
  assign n3572 = ~n3568 & ~n3571 ;
  assign n3573 = ~\g2016_reg/NET0131  & ~\g35_pad  ;
  assign n3574 = n3572 & ~n3573 ;
  assign n3575 = \g2834_reg/NET0131  & ~\g35_pad  ;
  assign n3576 = ~\g2715_reg/NET0131  & ~\g2815_reg/NET0131  ;
  assign n3577 = \g2715_reg/NET0131  & ~\g2819_reg/NET0131  ;
  assign n3578 = \g2719_reg/NET0131  & ~n3577 ;
  assign n3579 = ~n3576 & n3578 ;
  assign n3580 = ~\g2715_reg/NET0131  & ~\g2803_reg/NET0131  ;
  assign n3581 = ~\g2719_reg/NET0131  & ~n3041 ;
  assign n3582 = ~n3580 & n3581 ;
  assign n3583 = ~n3579 & ~n3582 ;
  assign n3584 = n3521 & n3583 ;
  assign n3585 = \g2638_reg/NET0131  & \g2715_reg/NET0131  ;
  assign n3586 = \g2504_reg/NET0131  & ~\g2715_reg/NET0131  ;
  assign n3587 = \g2719_reg/NET0131  & ~n3586 ;
  assign n3588 = ~n3585 & n3587 ;
  assign n3589 = \g2370_reg/NET0131  & \g2715_reg/NET0131  ;
  assign n3590 = \g2236_reg/NET0131  & ~\g2715_reg/NET0131  ;
  assign n3591 = ~\g2719_reg/NET0131  & ~n3590 ;
  assign n3592 = ~n3589 & n3591 ;
  assign n3593 = ~n3588 & ~n3592 ;
  assign n3594 = n3532 & n3593 ;
  assign n3595 = ~n3584 & ~n3594 ;
  assign n3596 = ~n3575 & n3595 ;
  assign n3597 = \g2610_reg/NET0131  & ~\g2619_reg/NET0131  ;
  assign n3598 = ~\g2555_reg/NET0131  & \g2599_reg/NET0131  ;
  assign n3599 = n3597 & n3598 ;
  assign n3600 = ~n3135 & n3599 ;
  assign n3601 = \g35_pad  & n3600 ;
  assign n3602 = ~n3135 & n3597 ;
  assign n3603 = ~\g2595_reg/NET0131  & \g35_pad  ;
  assign n3604 = ~n3602 & n3603 ;
  assign n3605 = ~n3601 & ~n3604 ;
  assign n3606 = ~\g2575_reg/NET0131  & ~\g35_pad  ;
  assign n3607 = n3605 & ~n3606 ;
  assign n3608 = \g142_reg/NET0131  & ~\g35_pad  ;
  assign n3609 = ~\g146_reg/NET0131  & ~n2344 ;
  assign n3610 = ~n2354 & ~n3609 ;
  assign n3611 = n2660 & n3610 ;
  assign n3612 = ~n3608 & ~n3611 ;
  assign n3613 = ~\g35_pad  & \g4443_reg/NET0131  ;
  assign n3614 = \g4438_reg/NET0131  & n1441 ;
  assign n3615 = ~n3613 & ~n3614 ;
  assign n3616 = ~n3128 & n3615 ;
  assign n3617 = ~\g35_pad  & \g4801_reg/NET0131  ;
  assign n3618 = \g4776_reg/NET0131  & \g4793_reg/NET0131  ;
  assign n3619 = n2838 & n3618 ;
  assign n3620 = \g35_pad  & ~n3619 ;
  assign n3621 = \g4793_reg/NET0131  & \g4801_reg/NET0131  ;
  assign n3622 = n2838 & n3621 ;
  assign n3623 = ~\g4776_reg/NET0131  & ~n3622 ;
  assign n3624 = n3620 & ~n3623 ;
  assign n3625 = ~n3617 & ~n3624 ;
  assign n3626 = ~\g35_pad  & \g671_reg/NET0131  ;
  assign n3627 = \g671_reg/NET0131  & n2579 ;
  assign n3628 = n2918 & n3627 ;
  assign n3629 = ~\g676_reg/NET0131  & ~n3628 ;
  assign n3630 = n2930 & ~n2934 ;
  assign n3631 = ~n2929 & n3630 ;
  assign n3632 = ~n3629 & n3631 ;
  assign n3633 = ~n3626 & ~n3632 ;
  assign n3634 = ~\g35_pad  & \g4659_reg/NET0131  ;
  assign n3635 = ~n2839 & ~n3634 ;
  assign n3636 = \g4659_reg/NET0131  & n2837 ;
  assign n3637 = ~\g4664_reg/NET0131  & ~n3634 ;
  assign n3638 = ~n3636 & n3637 ;
  assign n3639 = \g4664_reg/NET0131  & ~n3634 ;
  assign n3640 = n3636 & n3639 ;
  assign n3641 = ~n3638 & ~n3640 ;
  assign n3642 = ~n3635 & n3641 ;
  assign n3643 = \g1798_reg/NET0131  & ~\g35_pad  ;
  assign n3644 = ~\g1792_reg/NET0131  & ~n3045 ;
  assign n3645 = ~n3210 & n3644 ;
  assign n3646 = \g1783_reg/NET0131  & \g35_pad  ;
  assign n3647 = \g35_pad  & ~n3045 ;
  assign n3648 = ~n3210 & n3647 ;
  assign n3649 = ~n3646 & ~n3648 ;
  assign n3650 = ~n3645 & ~n3649 ;
  assign n3651 = ~n3643 & ~n3650 ;
  assign n3652 = \g1811_reg/NET0131  & ~n3045 ;
  assign n3653 = ~n3210 & n3652 ;
  assign n3654 = \g35_pad  & n3653 ;
  assign n3655 = \g1740_reg/NET0131  & \g1792_reg/NET0131  ;
  assign n3656 = \g1752_reg/NET0131  & ~\g1783_reg/NET0131  ;
  assign n3657 = ~n3655 & ~n3656 ;
  assign n3658 = \g1760_reg/NET0131  & ~n3657 ;
  assign n3659 = \g1748_reg/NET0131  & ~\g1760_reg/NET0131  ;
  assign n3660 = \g1756_reg/NET0131  & \g1783_reg/NET0131  ;
  assign n3661 = ~n3659 & ~n3660 ;
  assign n3662 = ~\g1792_reg/NET0131  & ~n3661 ;
  assign n3663 = \g1736_reg/NET0131  & n3213 ;
  assign n3664 = \g1744_reg/NET0131  & ~\g1783_reg/NET0131  ;
  assign n3665 = \g1792_reg/NET0131  & n3664 ;
  assign n3666 = ~n3663 & ~n3665 ;
  assign n3667 = ~n3662 & n3666 ;
  assign n3668 = ~n3658 & n3667 ;
  assign n3669 = \g35_pad  & ~n3211 ;
  assign n3670 = ~n3668 & n3669 ;
  assign n3671 = ~n3654 & ~n3670 ;
  assign n3672 = \g1792_reg/NET0131  & ~\g35_pad  ;
  assign n3673 = n3671 & ~n3672 ;
  assign n3674 = \g35_pad  & n2970 ;
  assign n3675 = ~\g1926_reg/NET0131  & \g35_pad  ;
  assign n3676 = n2970 & n3675 ;
  assign n3677 = ~\g1917_reg/NET0131  & \g35_pad  ;
  assign n3678 = ~n2970 & n3677 ;
  assign n3679 = ~n3676 & ~n3678 ;
  assign n3680 = ~\g1932_reg/NET0131  & ~\g35_pad  ;
  assign n3681 = n3679 & ~n3680 ;
  assign n3682 = \g1945_reg/NET0131  & n2970 ;
  assign n3683 = \g35_pad  & n3682 ;
  assign n3684 = \g1874_reg/NET0131  & \g1926_reg/NET0131  ;
  assign n3685 = \g1886_reg/NET0131  & ~\g1917_reg/NET0131  ;
  assign n3686 = ~n3684 & ~n3685 ;
  assign n3687 = \g1894_reg/NET0131  & ~n3686 ;
  assign n3688 = \g1882_reg/NET0131  & ~\g1894_reg/NET0131  ;
  assign n3689 = \g1890_reg/NET0131  & \g1917_reg/NET0131  ;
  assign n3690 = ~n3688 & ~n3689 ;
  assign n3691 = ~\g1926_reg/NET0131  & ~n3690 ;
  assign n3692 = \g1870_reg/NET0131  & n3264 ;
  assign n3693 = \g1878_reg/NET0131  & ~\g1917_reg/NET0131  ;
  assign n3694 = \g1926_reg/NET0131  & n3693 ;
  assign n3695 = ~n3692 & ~n3694 ;
  assign n3696 = ~n3691 & n3695 ;
  assign n3697 = ~n3687 & n3696 ;
  assign n3698 = \g35_pad  & ~n2970 ;
  assign n3699 = ~n3697 & n3698 ;
  assign n3700 = ~n3683 & ~n3699 ;
  assign n3701 = \g1926_reg/NET0131  & ~\g35_pad  ;
  assign n3702 = n3700 & ~n3701 ;
  assign n3703 = \g35_pad  & n3302 ;
  assign n3704 = \g2066_reg/NET0131  & ~\g35_pad  ;
  assign n3705 = \g2060_reg/NET0131  & \g35_pad  ;
  assign n3706 = n3302 & n3705 ;
  assign n3707 = \g2051_reg/NET0131  & \g35_pad  ;
  assign n3708 = ~n3302 & n3707 ;
  assign n3709 = ~n3706 & ~n3708 ;
  assign n3710 = ~n3704 & n3709 ;
  assign n3711 = \g2079_reg/NET0131  & n3302 ;
  assign n3712 = \g35_pad  & n3711 ;
  assign n3713 = \g2008_reg/NET0131  & \g2060_reg/NET0131  ;
  assign n3714 = \g2020_reg/NET0131  & ~\g2051_reg/NET0131  ;
  assign n3715 = ~n3713 & ~n3714 ;
  assign n3716 = \g2028_reg/NET0131  & ~n3715 ;
  assign n3717 = \g2016_reg/NET0131  & ~\g2028_reg/NET0131  ;
  assign n3718 = \g2024_reg/NET0131  & \g2051_reg/NET0131  ;
  assign n3719 = ~n3717 & ~n3718 ;
  assign n3720 = ~\g2060_reg/NET0131  & ~n3719 ;
  assign n3721 = \g2004_reg/NET0131  & n3303 ;
  assign n3722 = \g2012_reg/NET0131  & ~\g2051_reg/NET0131  ;
  assign n3723 = \g2060_reg/NET0131  & n3722 ;
  assign n3724 = ~n3721 & ~n3723 ;
  assign n3725 = ~n3720 & n3724 ;
  assign n3726 = ~n3716 & n3725 ;
  assign n3727 = \g35_pad  & ~n3302 ;
  assign n3728 = ~n3726 & n3727 ;
  assign n3729 = ~n3712 & ~n3728 ;
  assign n3730 = \g2060_reg/NET0131  & ~\g35_pad  ;
  assign n3731 = n3729 & ~n3730 ;
  assign n3732 = \g411_reg/NET0131  & ~n2579 ;
  assign n3733 = \g35_pad  & n3732 ;
  assign n3734 = \g35_pad  & n2579 ;
  assign n3735 = ~n3008 & n3734 ;
  assign n3736 = ~n3733 & ~n3735 ;
  assign n3737 = ~\g35_pad  & \g417_reg/NET0131  ;
  assign n3738 = n3736 & ~n3737 ;
  assign n3739 = \g35_pad  & n3029 ;
  assign n3740 = ~\g2217_reg/NET0131  & \g35_pad  ;
  assign n3741 = n3029 & n3740 ;
  assign n3742 = ~\g2208_reg/NET0131  & \g35_pad  ;
  assign n3743 = ~n3029 & n3742 ;
  assign n3744 = ~n3741 & ~n3743 ;
  assign n3745 = ~\g2223_reg/NET0131  & ~\g35_pad  ;
  assign n3746 = n3744 & ~n3745 ;
  assign n3747 = \g2236_reg/NET0131  & n3029 ;
  assign n3748 = \g35_pad  & n3747 ;
  assign n3749 = \g2169_reg/NET0131  & ~\g2208_reg/NET0131  ;
  assign n3750 = \g2165_reg/NET0131  & \g2185_reg/NET0131  ;
  assign n3751 = ~n3749 & ~n3750 ;
  assign n3752 = \g2217_reg/NET0131  & ~n3751 ;
  assign n3753 = \g2173_reg/NET0131  & ~\g2217_reg/NET0131  ;
  assign n3754 = \g2161_reg/NET0131  & \g2208_reg/NET0131  ;
  assign n3755 = ~n3753 & ~n3754 ;
  assign n3756 = ~\g2185_reg/NET0131  & ~n3755 ;
  assign n3757 = \g2181_reg/NET0131  & n3031 ;
  assign n3758 = \g2177_reg/NET0131  & \g2185_reg/NET0131  ;
  assign n3759 = ~\g2208_reg/NET0131  & n3758 ;
  assign n3760 = ~n3757 & ~n3759 ;
  assign n3761 = ~n3756 & n3760 ;
  assign n3762 = ~n3752 & n3761 ;
  assign n3763 = \g35_pad  & ~n3029 ;
  assign n3764 = ~n3762 & n3763 ;
  assign n3765 = ~n3748 & ~n3764 ;
  assign n3766 = \g2217_reg/NET0131  & ~\g35_pad  ;
  assign n3767 = n3765 & ~n3766 ;
  assign n3768 = ~n3043 & n3647 ;
  assign n3769 = ~\g2351_reg/NET0131  & ~n3045 ;
  assign n3770 = ~n3043 & n3769 ;
  assign n3771 = \g35_pad  & n3770 ;
  assign n3772 = ~\g2342_reg/NET0131  & \g35_pad  ;
  assign n3773 = ~n3046 & n3772 ;
  assign n3774 = ~n3771 & ~n3773 ;
  assign n3775 = ~\g2357_reg/NET0131  & ~\g35_pad  ;
  assign n3776 = n3774 & ~n3775 ;
  assign n3777 = \g2370_reg/NET0131  & ~n3045 ;
  assign n3778 = ~n3043 & n3777 ;
  assign n3779 = \g35_pad  & n3778 ;
  assign n3780 = \g2303_reg/NET0131  & ~\g2342_reg/NET0131  ;
  assign n3781 = \g2299_reg/NET0131  & \g2319_reg/NET0131  ;
  assign n3782 = ~n3780 & ~n3781 ;
  assign n3783 = \g2351_reg/NET0131  & ~n3782 ;
  assign n3784 = \g2307_reg/NET0131  & ~\g2351_reg/NET0131  ;
  assign n3785 = \g2295_reg/NET0131  & \g2342_reg/NET0131  ;
  assign n3786 = ~n3784 & ~n3785 ;
  assign n3787 = ~\g2319_reg/NET0131  & ~n3786 ;
  assign n3788 = \g2315_reg/NET0131  & n3048 ;
  assign n3789 = \g2311_reg/NET0131  & \g2319_reg/NET0131  ;
  assign n3790 = ~\g2342_reg/NET0131  & n3789 ;
  assign n3791 = ~n3788 & ~n3790 ;
  assign n3792 = ~n3787 & n3791 ;
  assign n3793 = ~n3783 & n3792 ;
  assign n3794 = \g35_pad  & ~n3046 ;
  assign n3795 = ~n3793 & n3794 ;
  assign n3796 = ~n3779 & ~n3795 ;
  assign n3797 = \g2351_reg/NET0131  & ~\g35_pad  ;
  assign n3798 = n3796 & ~n3797 ;
  assign n3799 = \g35_pad  & n3081 ;
  assign n3800 = ~\g2485_reg/NET0131  & \g35_pad  ;
  assign n3801 = n3081 & n3800 ;
  assign n3802 = ~\g2476_reg/NET0131  & \g35_pad  ;
  assign n3803 = ~n3081 & n3802 ;
  assign n3804 = ~n3801 & ~n3803 ;
  assign n3805 = ~\g2491_reg/NET0131  & ~\g35_pad  ;
  assign n3806 = n3804 & ~n3805 ;
  assign n3807 = \g2504_reg/NET0131  & n3081 ;
  assign n3808 = \g35_pad  & n3807 ;
  assign n3809 = \g2437_reg/NET0131  & ~\g2476_reg/NET0131  ;
  assign n3810 = \g2433_reg/NET0131  & \g2453_reg/NET0131  ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3812 = \g2485_reg/NET0131  & ~n3811 ;
  assign n3813 = \g2441_reg/NET0131  & ~\g2485_reg/NET0131  ;
  assign n3814 = \g2429_reg/NET0131  & \g2476_reg/NET0131  ;
  assign n3815 = ~n3813 & ~n3814 ;
  assign n3816 = ~\g2453_reg/NET0131  & ~n3815 ;
  assign n3817 = \g2449_reg/NET0131  & n3083 ;
  assign n3818 = \g2445_reg/NET0131  & \g2453_reg/NET0131  ;
  assign n3819 = ~\g2476_reg/NET0131  & n3818 ;
  assign n3820 = ~n3817 & ~n3819 ;
  assign n3821 = ~n3816 & n3820 ;
  assign n3822 = ~n3812 & n3821 ;
  assign n3823 = \g35_pad  & ~n3081 ;
  assign n3824 = ~n3822 & n3823 ;
  assign n3825 = ~n3808 & ~n3824 ;
  assign n3826 = \g2485_reg/NET0131  & ~\g35_pad  ;
  assign n3827 = n3825 & ~n3826 ;
  assign n3828 = \g35_pad  & n3095 ;
  assign n3829 = ~\g1657_reg/NET0131  & \g35_pad  ;
  assign n3830 = n3095 & n3829 ;
  assign n3831 = ~\g1648_reg/NET0131  & \g35_pad  ;
  assign n3832 = ~n3095 & n3831 ;
  assign n3833 = ~n3830 & ~n3832 ;
  assign n3834 = ~\g1664_reg/NET0131  & ~\g35_pad  ;
  assign n3835 = n3833 & ~n3834 ;
  assign n3836 = \g35_pad  & n3135 ;
  assign n3837 = \g1677_reg/NET0131  & n3095 ;
  assign n3838 = \g35_pad  & n3837 ;
  assign n3839 = \g1604_reg/NET0131  & \g1657_reg/NET0131  ;
  assign n3840 = \g1616_reg/NET0131  & ~\g1648_reg/NET0131  ;
  assign n3841 = ~n3839 & ~n3840 ;
  assign n3842 = \g1624_reg/NET0131  & ~n3841 ;
  assign n3843 = \g1612_reg/NET0131  & ~\g1624_reg/NET0131  ;
  assign n3844 = \g1620_reg/NET0131  & \g1648_reg/NET0131  ;
  assign n3845 = ~n3843 & ~n3844 ;
  assign n3846 = ~\g1657_reg/NET0131  & ~n3845 ;
  assign n3847 = \g1600_reg/NET0131  & n3158 ;
  assign n3848 = \g1608_reg/NET0131  & ~\g1648_reg/NET0131  ;
  assign n3849 = \g1657_reg/NET0131  & n3848 ;
  assign n3850 = ~n3847 & ~n3849 ;
  assign n3851 = ~n3846 & n3850 ;
  assign n3852 = ~n3842 & n3851 ;
  assign n3853 = \g35_pad  & ~n3095 ;
  assign n3854 = ~n3852 & n3853 ;
  assign n3855 = ~n3838 & ~n3854 ;
  assign n3856 = \g1657_reg/NET0131  & ~\g35_pad  ;
  assign n3857 = n3855 & ~n3856 ;
  assign n3858 = \g2625_reg/NET0131  & ~\g35_pad  ;
  assign n3859 = \g2619_reg/NET0131  & \g35_pad  ;
  assign n3860 = n3135 & n3859 ;
  assign n3861 = \g2610_reg/NET0131  & \g35_pad  ;
  assign n3862 = ~n3135 & n3861 ;
  assign n3863 = ~n3860 & ~n3862 ;
  assign n3864 = ~n3858 & n3863 ;
  assign n3865 = \g2638_reg/NET0131  & n3135 ;
  assign n3866 = \g35_pad  & n3865 ;
  assign n3867 = \g2579_reg/NET0131  & \g2587_reg/NET0131  ;
  assign n3868 = \g2571_reg/NET0131  & \g2619_reg/NET0131  ;
  assign n3869 = ~n3867 & ~n3868 ;
  assign n3870 = ~\g2610_reg/NET0131  & ~n3869 ;
  assign n3871 = \g2575_reg/NET0131  & ~\g2587_reg/NET0131  ;
  assign n3872 = \g2583_reg/NET0131  & \g2610_reg/NET0131  ;
  assign n3873 = ~n3871 & ~n3872 ;
  assign n3874 = ~\g2619_reg/NET0131  & ~n3873 ;
  assign n3875 = \g2563_reg/NET0131  & n3136 ;
  assign n3876 = \g2567_reg/NET0131  & \g2587_reg/NET0131  ;
  assign n3877 = \g2619_reg/NET0131  & n3876 ;
  assign n3878 = ~n3875 & ~n3877 ;
  assign n3879 = ~n3874 & n3878 ;
  assign n3880 = ~n3870 & n3879 ;
  assign n3881 = \g35_pad  & ~n3135 ;
  assign n3882 = ~n3880 & n3881 ;
  assign n3883 = ~n3866 & ~n3882 ;
  assign n3884 = \g2619_reg/NET0131  & ~\g35_pad  ;
  assign n3885 = n3883 & ~n3884 ;
  assign n3886 = \g1691_reg/NET0131  & \g35_pad  ;
  assign n3887 = n3095 & n3886 ;
  assign n3888 = ~n3158 & n3886 ;
  assign n3889 = ~\g1677_reg/NET0131  & ~n3888 ;
  assign n3890 = \g1677_reg/NET0131  & n3888 ;
  assign n3891 = ~n3889 & ~n3890 ;
  assign n3892 = ~n3828 & n3891 ;
  assign n3893 = ~n3887 & ~n3892 ;
  assign n3894 = \g1825_reg/NET0131  & \g35_pad  ;
  assign n3895 = ~n3045 & n3894 ;
  assign n3896 = ~n3210 & n3895 ;
  assign n3897 = ~n3213 & n3894 ;
  assign n3898 = ~\g1811_reg/NET0131  & ~n3897 ;
  assign n3899 = \g1811_reg/NET0131  & n3897 ;
  assign n3900 = ~n3898 & ~n3899 ;
  assign n3901 = ~n3648 & n3900 ;
  assign n3902 = ~n3896 & ~n3901 ;
  assign n3903 = \g35_pad  & ~n2505 ;
  assign n3904 = \g316_reg/NET0131  & ~\g35_pad  ;
  assign n3905 = ~n3903 & ~n3904 ;
  assign n3906 = \g1008_reg/NET0131  & ~\g1046_reg/NET0131  ;
  assign n3907 = ~n2815 & ~n3906 ;
  assign n3908 = ~\g969_reg/NET0131  & ~n3907 ;
  assign n3909 = \g1018_reg/NET0131  & \g1030_reg/NET0131  ;
  assign n3910 = \g1008_reg/NET0131  & n3909 ;
  assign n3911 = n2815 & n3910 ;
  assign n3912 = \g1002_reg/NET0131  & \g1018_reg/NET0131  ;
  assign n3913 = ~n3911 & ~n3912 ;
  assign n3914 = n3908 & n3913 ;
  assign n3915 = ~n2816 & ~n3914 ;
  assign n3916 = ~\g1024_reg/NET0131  & ~n3911 ;
  assign n3917 = n3908 & n3916 ;
  assign n3918 = ~\g1030_reg/NET0131  & ~\g969_reg/NET0131  ;
  assign n3919 = ~n3907 & n3918 ;
  assign n3920 = ~n3917 & ~n3919 ;
  assign n3921 = n3915 & n3920 ;
  assign n3922 = ~\g1036_reg/NET0131  & ~n3911 ;
  assign n3923 = n3908 & n3922 ;
  assign n3924 = \g35_pad  & ~n3923 ;
  assign n3925 = n3921 & n3924 ;
  assign n3926 = ~\g1036_reg/NET0131  & \g35_pad  ;
  assign n3927 = ~n3921 & n3926 ;
  assign n3928 = ~n3925 & ~n3927 ;
  assign n3929 = ~\g1030_reg/NET0131  & ~\g35_pad  ;
  assign n3930 = n3928 & ~n3929 ;
  assign n3931 = \g1959_reg/NET0131  & \g35_pad  ;
  assign n3932 = n2970 & n3931 ;
  assign n3933 = ~n3264 & n3931 ;
  assign n3934 = ~\g1945_reg/NET0131  & ~n3933 ;
  assign n3935 = \g1945_reg/NET0131  & n3933 ;
  assign n3936 = ~n3934 & ~n3935 ;
  assign n3937 = ~n3674 & n3936 ;
  assign n3938 = ~n3932 & ~n3937 ;
  assign n3939 = \g2250_reg/NET0131  & \g35_pad  ;
  assign n3940 = n3029 & n3939 ;
  assign n3941 = ~n3339 & n3939 ;
  assign n3942 = ~\g2236_reg/NET0131  & ~n3941 ;
  assign n3943 = \g2236_reg/NET0131  & n3941 ;
  assign n3944 = ~n3942 & ~n3943 ;
  assign n3945 = ~n3739 & n3944 ;
  assign n3946 = ~n3940 & ~n3945 ;
  assign n3947 = \g2384_reg/NET0131  & \g35_pad  ;
  assign n3948 = ~n3045 & n3947 ;
  assign n3949 = ~n3043 & n3948 ;
  assign n3950 = ~n3376 & n3947 ;
  assign n3951 = ~\g2370_reg/NET0131  & ~n3950 ;
  assign n3952 = \g2370_reg/NET0131  & n3950 ;
  assign n3953 = ~n3951 & ~n3952 ;
  assign n3954 = ~n3768 & n3953 ;
  assign n3955 = ~n3949 & ~n3954 ;
  assign n3956 = \g2518_reg/NET0131  & \g35_pad  ;
  assign n3957 = n3081 & n3956 ;
  assign n3958 = ~n3428 & n3956 ;
  assign n3959 = ~\g2504_reg/NET0131  & ~n3958 ;
  assign n3960 = \g2504_reg/NET0131  & n3958 ;
  assign n3961 = ~n3959 & ~n3960 ;
  assign n3962 = ~n3799 & n3961 ;
  assign n3963 = ~n3957 & ~n3962 ;
  assign n3964 = ~\g35_pad  & \g739_reg/NET0131  ;
  assign n3965 = \g35_pad  & ~n3559 ;
  assign n3966 = \g739_reg/NET0131  & n982 ;
  assign n3967 = n975 & n3966 ;
  assign n3968 = n995 & n3967 ;
  assign n3969 = ~\g744_reg/NET0131  & ~n3968 ;
  assign n3970 = ~n976 & ~n3969 ;
  assign n3971 = n3965 & n3970 ;
  assign n3972 = ~n3964 & ~n3971 ;
  assign n3973 = \g2093_reg/NET0131  & \g35_pad  ;
  assign n3974 = n3302 & n3973 ;
  assign n3975 = ~n3303 & n3973 ;
  assign n3976 = ~\g2079_reg/NET0131  & ~n3975 ;
  assign n3977 = \g2079_reg/NET0131  & n3975 ;
  assign n3978 = ~n3976 & ~n3977 ;
  assign n3979 = ~n3703 & n3978 ;
  assign n3980 = ~n3974 & ~n3979 ;
  assign n3981 = \g2652_reg/NET0131  & \g35_pad  ;
  assign n3982 = n3135 & n3981 ;
  assign n3983 = ~n3136 & n3981 ;
  assign n3984 = ~\g2638_reg/NET0131  & ~n3983 ;
  assign n3985 = \g2638_reg/NET0131  & n3983 ;
  assign n3986 = ~n3984 & ~n3985 ;
  assign n3987 = ~n3836 & n3986 ;
  assign n3988 = ~n3982 & ~n3987 ;
  assign n3989 = \g358_reg/NET0131  & ~\g376_reg/NET0131  ;
  assign n3990 = \g385_reg/NET0131  & n3989 ;
  assign n3991 = n2343 & n3990 ;
  assign n3992 = ~\g528_reg/NET0131  & ~n2915 ;
  assign n3993 = \g667_reg/NET0131  & ~\g686_reg/NET0131  ;
  assign n3994 = \g490_reg/NET0131  & ~n3993 ;
  assign n3995 = ~n3992 & ~n3994 ;
  assign n3996 = n3991 & n3995 ;
  assign n3997 = \g35_pad  & ~n3996 ;
  assign n3998 = \g482_reg/NET0131  & ~n3997 ;
  assign n3999 = \g482_reg/NET0131  & ~n3992 ;
  assign n4000 = n3991 & n3999 ;
  assign n4001 = ~\g490_reg/NET0131  & ~n3993 ;
  assign n4002 = \g35_pad  & ~n4001 ;
  assign n4003 = ~n4000 & n4002 ;
  assign n4004 = ~n3998 & ~n4003 ;
  assign n4005 = ~\g35_pad  & \g736_reg/NET0131  ;
  assign n4006 = n995 & n2350 ;
  assign n4007 = ~\g739_reg/NET0131  & ~n4006 ;
  assign n4008 = \g35_pad  & ~n976 ;
  assign n4009 = ~n3968 & n4008 ;
  assign n4010 = ~n4007 & n4009 ;
  assign n4011 = ~n4005 & ~n4010 ;
  assign n4012 = \g1087_reg/NET0131  & \g1205_reg/NET0131  ;
  assign n4013 = \g1221_reg/NET0131  & n4012 ;
  assign n4014 = \g1211_reg/NET0131  & \g35_pad  ;
  assign n4015 = ~n4013 & n4014 ;
  assign n4016 = ~\g1211_reg/NET0131  & \g1221_reg/NET0131  ;
  assign n4017 = n4012 & n4016 ;
  assign n4018 = \g35_pad  & ~n4017 ;
  assign n4019 = \g1216_reg/NET0131  & ~n4018 ;
  assign n4020 = ~n4015 & ~n4019 ;
  assign n4021 = n2524 & n2525 ;
  assign n4022 = \g35_pad  & ~n4021 ;
  assign n4023 = \g4311_reg/NET0131  & \g4628_reg/NET0131  ;
  assign n4024 = n2520 & n4023 ;
  assign n4025 = n2523 & n4024 ;
  assign n4026 = \g4322_reg/NET0131  & n4025 ;
  assign n4027 = \g4332_reg/NET0131  & ~n4026 ;
  assign n4028 = n4022 & n4027 ;
  assign n4029 = ~\g35_pad  & \g4322_reg/NET0131  ;
  assign n4030 = \g4322_reg/NET0131  & ~\g4332_reg/NET0131  ;
  assign n4031 = n4025 & n4030 ;
  assign n4032 = ~n4029 & ~n4031 ;
  assign n4033 = ~n4028 & n4032 ;
  assign n4034 = \g1559_reg/NET0131  & ~\g35_pad  ;
  assign n4035 = \g35_pad  & ~n1463 ;
  assign n4036 = \g1559_reg/NET0131  & \g1564_reg/NET0131  ;
  assign n4037 = n1461 & n4036 ;
  assign n4038 = ~\g1554_reg/NET0131  & ~n4037 ;
  assign n4039 = n4035 & ~n4038 ;
  assign n4040 = ~n4034 & ~n4039 ;
  assign n4041 = ~\g5069_reg/NET0131  & \g5084_reg/NET0131  ;
  assign n4042 = ~\g5073_reg/NET0131  & ~\g5084_reg/NET0131  ;
  assign n4043 = \g35_pad  & ~n4042 ;
  assign n4044 = ~n4041 & n4043 ;
  assign n4045 = \g5077_reg/NET0131  & ~n4044 ;
  assign n4046 = \g246_reg/NET0131  & \g35_pad  ;
  assign n4047 = ~\g35_pad  & \g479_reg/NET0131  ;
  assign n4048 = ~n4046 & ~n4047 ;
  assign n4049 = ~\g35_pad  & \g4584_reg/NET0131  ;
  assign n4050 = \g35_pad  & \g4593_reg/NET0131  ;
  assign n4051 = ~n2532 & n4050 ;
  assign n4052 = \g35_pad  & ~\g4616_reg/NET0131  ;
  assign n4053 = ~\g4593_reg/NET0131  & n4052 ;
  assign n4054 = n2532 & n4053 ;
  assign n4055 = ~n4051 & ~n4054 ;
  assign n4056 = ~n4049 & n4055 ;
  assign n4057 = ~\g862_reg/NET0131  & \g890_reg/NET0131  ;
  assign n4058 = \g872_reg/NET0131  & ~\g896_reg/NET0131  ;
  assign n4059 = n4057 & n4058 ;
  assign n4060 = \g35_pad  & n4059 ;
  assign n4061 = ~\g896_reg/NET0131  & n4057 ;
  assign n4062 = \g35_pad  & \g446_reg/NET0131  ;
  assign n4063 = ~n4061 & n4062 ;
  assign n4064 = ~n4060 & ~n4063 ;
  assign n4065 = \g246_reg/NET0131  & ~\g35_pad  ;
  assign n4066 = n4064 & ~n4065 ;
  assign n4067 = \g854_reg/NET0131  & ~n2986 ;
  assign n4068 = n3014 & ~n4067 ;
  assign n4069 = \g35_pad  & ~n4068 ;
  assign n4070 = ~\g4340_reg/NET0131  & n1072 ;
  assign n4071 = ~\g4340_reg/NET0131  & n1069 ;
  assign n4072 = n1077 & n4071 ;
  assign n4073 = ~n4070 & ~n4072 ;
  assign n4074 = \g4349_reg/NET0131  & n4073 ;
  assign n4075 = \g4311_reg/NET0131  & ~\g4322_reg/NET0131  ;
  assign n4076 = \g4332_reg/NET0131  & n4075 ;
  assign n4077 = ~\g4515_reg/NET0131  & n4030 ;
  assign n4078 = ~\g4340_reg/NET0131  & ~\g4349_reg/NET0131  ;
  assign n4079 = ~n4077 & n4078 ;
  assign n4080 = ~n4076 & n4079 ;
  assign n4081 = \g35_pad  & ~\g4358_reg/NET0131  ;
  assign n4082 = ~n4080 & n4081 ;
  assign n4083 = ~n4074 & n4082 ;
  assign n4084 = ~\g35_pad  & \g4366_reg/NET0131  ;
  assign n4085 = \g35_pad  & \g4358_reg/NET0131  ;
  assign n4086 = ~n4084 & ~n4085 ;
  assign n4087 = ~n2522 & ~n4084 ;
  assign n4088 = n4073 & n4087 ;
  assign n4089 = ~n4086 & ~n4088 ;
  assign n4090 = ~n4083 & ~n4089 ;
  assign n4091 = \g1024_reg/NET0131  & ~\g35_pad  ;
  assign n4092 = n3915 & ~n3917 ;
  assign n4093 = ~\g1030_reg/NET0131  & ~n4092 ;
  assign n4094 = \g35_pad  & ~n3921 ;
  assign n4095 = ~n4093 & n4094 ;
  assign n4096 = ~n4091 & ~n4095 ;
  assign n4097 = \g4785_reg/NET0131  & n3618 ;
  assign n4098 = n2838 & n4097 ;
  assign n4099 = \g35_pad  & \g4709_reg/NET0131  ;
  assign n4100 = ~n4098 & n4099 ;
  assign n4101 = \g4785_reg/NET0131  & ~n4099 ;
  assign n4102 = ~n3620 & n4101 ;
  assign n4103 = ~n4100 & ~n4102 ;
  assign n4104 = ~\g35_pad  & ~\g843_reg/NET0131  ;
  assign n4105 = \g843_reg/NET0131  & \g847_reg/NET0131  ;
  assign n4106 = n2579 & n4105 ;
  assign n4107 = ~\g812_reg/NET0131  & ~n4106 ;
  assign n4108 = \g812_reg/NET0131  & \g847_reg/NET0131  ;
  assign n4109 = \g843_reg/NET0131  & n4108 ;
  assign n4110 = n2579 & n4109 ;
  assign n4111 = \g837_reg/NET0131  & ~n4110 ;
  assign n4112 = ~n4107 & n4111 ;
  assign n4113 = \g35_pad  & ~n4112 ;
  assign n4114 = ~n4104 & ~n4113 ;
  assign n4115 = ~\g35_pad  & \g667_reg/NET0131  ;
  assign n4116 = ~\g671_reg/NET0131  & ~n2919 ;
  assign n4117 = ~n3628 & ~n4116 ;
  assign n4118 = n2931 & n4117 ;
  assign n4119 = ~n4115 & ~n4118 ;
  assign n4120 = ~\g283_reg/NET0131  & \g35_pad  ;
  assign n4121 = n2388 & n4120 ;
  assign n4122 = \g278_reg/NET0131  & ~\g35_pad  ;
  assign n4123 = ~n4121 & ~n4122 ;
  assign n4124 = ~\g35_pad  & \g817_reg/NET0131  ;
  assign n4125 = \g817_reg/NET0131  & n2579 ;
  assign n4126 = ~\g832_reg/NET0131  & ~n4125 ;
  assign n4127 = n2586 & ~n3122 ;
  assign n4128 = ~n4126 & n4127 ;
  assign n4129 = ~n4124 & ~n4128 ;
  assign n4130 = ~\g35_pad  & \g4793_reg/NET0131  ;
  assign n4131 = \g4793_reg/NET0131  & n2838 ;
  assign n4132 = \g35_pad  & \g4801_reg/NET0131  ;
  assign n4133 = ~n4131 & n4132 ;
  assign n4134 = \g35_pad  & ~\g4801_reg/NET0131  ;
  assign n4135 = ~\g4776_reg/NET0131  & n4134 ;
  assign n4136 = n4131 & n4135 ;
  assign n4137 = ~n4133 & ~n4136 ;
  assign n4138 = ~n4130 & n4137 ;
  assign n4139 = ~\g5016_reg/NET0131  & \g5022_reg/NET0131  ;
  assign n4140 = ~\g5029_reg/NET0131  & ~\g5033_reg/NET0131  ;
  assign n4141 = n4139 & n4140 ;
  assign n4142 = ~\g5037_reg/NET0131  & ~\g5046_reg/NET0131  ;
  assign n4143 = ~\g5041_reg/NET0131  & n4142 ;
  assign n4144 = n4141 & n4143 ;
  assign n4145 = \g3050_reg/NET0131  & \g5016_reg/NET0131  ;
  assign n4146 = \g5029_reg/NET0131  & \g5033_reg/NET0131  ;
  assign n4147 = n4145 & n4146 ;
  assign n4148 = \g5037_reg/NET0131  & \g5046_reg/NET0131  ;
  assign n4149 = \g5041_reg/NET0131  & n4148 ;
  assign n4150 = n4147 & n4149 ;
  assign n4151 = ~n4144 & ~n4150 ;
  assign n4152 = \g3050_reg/NET0131  & \g5046_reg/NET0131  ;
  assign n4153 = \g5052_reg/NET0131  & ~\g5057_reg/NET0131  ;
  assign n4154 = n4152 & n4153 ;
  assign n4155 = \g5052_reg/NET0131  & ~n4154 ;
  assign n4156 = \g35_pad  & n4155 ;
  assign n4157 = n4151 & n4156 ;
  assign n4158 = \g35_pad  & ~\g5052_reg/NET0131  ;
  assign n4159 = ~n4151 & n4158 ;
  assign n4160 = ~n4157 & ~n4159 ;
  assign n4161 = ~\g35_pad  & \g5046_reg/NET0131  ;
  assign n4162 = n4160 & ~n4161 ;
  assign n4163 = \g686_reg/NET0131  & ~n3990 ;
  assign n4164 = \g35_pad  & n4163 ;
  assign n4165 = ~\g691_reg/NET0131  & \g703_reg/NET0131  ;
  assign n4166 = ~n2920 & n4165 ;
  assign n4167 = n2927 & n4166 ;
  assign n4168 = \g35_pad  & n3990 ;
  assign n4169 = ~n4167 & n4168 ;
  assign n4170 = ~n4164 & ~n4169 ;
  assign n4171 = ~\g35_pad  & \g691_reg/NET0131  ;
  assign n4172 = n4170 & ~n4171 ;
  assign n4173 = \g316_reg/NET0131  & \g35_pad  ;
  assign n4174 = \g29216_pad  & ~\g35_pad  ;
  assign n4175 = ~n4173 & ~n4174 ;
  assign n4176 = ~\g35_pad  & \g4776_reg/NET0131  ;
  assign n4177 = \g35_pad  & ~n4098 ;
  assign n4178 = ~\g4785_reg/NET0131  & ~n3619 ;
  assign n4179 = n4177 & ~n4178 ;
  assign n4180 = ~n4176 & ~n4179 ;
  assign n4181 = \g14167_pad  & ~\g896_reg/NET0131  ;
  assign n4182 = n4057 & n4181 ;
  assign n4183 = \g35_pad  & n4182 ;
  assign n4184 = n4046 & ~n4061 ;
  assign n4185 = ~n4183 & ~n4184 ;
  assign n4186 = \g269_reg/NET0131  & ~\g35_pad  ;
  assign n4187 = n4185 & ~n4186 ;
  assign n4188 = ~\g1171_reg/NET0131  & ~\g7916_pad  ;
  assign n4189 = \g1171_reg/NET0131  & \g7916_pad  ;
  assign n4190 = ~n4188 & ~n4189 ;
  assign n4191 = \g35_pad  & n4190 ;
  assign n4192 = \g1178_reg/NET0131  & ~\g1189_reg/NET0131  ;
  assign n4193 = \g7916_pad  & \g996_reg/NET0131  ;
  assign n4194 = n4192 & n4193 ;
  assign n4195 = ~n817 & n4194 ;
  assign n4196 = n2815 & ~n2816 ;
  assign n4197 = \g1002_reg/NET0131  & \g1024_reg/NET0131  ;
  assign n4198 = \g1036_reg/NET0131  & n4197 ;
  assign n4199 = n4194 & n4198 ;
  assign n4200 = n4196 & n4199 ;
  assign n4201 = ~n4195 & ~n4200 ;
  assign n4202 = \g1193_reg/NET0131  & ~n1386 ;
  assign n4203 = \g35_pad  & ~n4202 ;
  assign n4204 = ~n4201 & n4203 ;
  assign n4205 = ~n4191 & ~n4204 ;
  assign n4206 = \g1018_reg/NET0131  & ~\g35_pad  ;
  assign n4207 = \g1024_reg/NET0131  & \g35_pad  ;
  assign n4208 = ~n3915 & n4207 ;
  assign n4209 = \g35_pad  & n3917 ;
  assign n4210 = n3915 & n4209 ;
  assign n4211 = ~n4208 & ~n4210 ;
  assign n4212 = ~n4206 & n4211 ;
  assign n4213 = ~n4201 & ~n4202 ;
  assign n4214 = \g996_reg/NET0131  & n4192 ;
  assign n4215 = \g1199_reg/NET0131  & \g7916_pad  ;
  assign n4216 = n1386 & n4215 ;
  assign n4217 = ~n4214 & n4216 ;
  assign n4218 = \g35_pad  & ~n4217 ;
  assign n4219 = \g1070_reg/NET0131  & n4218 ;
  assign n4220 = ~n4213 & n4219 ;
  assign n4221 = ~\g1070_reg/NET0131  & \g7916_pad  ;
  assign n4222 = n1386 & n4221 ;
  assign n4223 = ~n4214 & n4222 ;
  assign n4224 = \g35_pad  & ~n4223 ;
  assign n4225 = \g1199_reg/NET0131  & ~n4224 ;
  assign n4226 = ~n4220 & ~n4225 ;
  assign n4227 = ~\g5052_reg/NET0131  & n4144 ;
  assign n4228 = \g5052_reg/NET0131  & n4150 ;
  assign n4229 = ~n4227 & ~n4228 ;
  assign n4230 = \g35_pad  & ~n4154 ;
  assign n4231 = \g5022_reg/NET0131  & ~\g5046_reg/NET0131  ;
  assign n4232 = ~\g5052_reg/NET0131  & \g5057_reg/NET0131  ;
  assign n4233 = n4231 & n4232 ;
  assign n4234 = \g5057_reg/NET0131  & ~n4233 ;
  assign n4235 = n4230 & n4234 ;
  assign n4236 = n4229 & n4235 ;
  assign n4237 = ~\g35_pad  & \g5052_reg/NET0131  ;
  assign n4238 = \g35_pad  & ~\g5057_reg/NET0131  ;
  assign n4239 = \g5052_reg/NET0131  & n4238 ;
  assign n4240 = n4150 & n4239 ;
  assign n4241 = ~\g5052_reg/NET0131  & n4238 ;
  assign n4242 = n4144 & n4241 ;
  assign n4243 = ~n4240 & ~n4242 ;
  assign n4244 = ~n4237 & n4243 ;
  assign n4245 = ~n4236 & n4244 ;
  assign n4246 = ~\g1216_reg/NET0131  & \g35_pad  ;
  assign n4247 = ~n4013 & n4246 ;
  assign n4248 = \g35_pad  & ~n1605 ;
  assign n4249 = n4013 & n4248 ;
  assign n4250 = ~n4247 & ~n4249 ;
  assign n4251 = ~\g1221_reg/NET0131  & ~\g35_pad  ;
  assign n4252 = n4250 & ~n4251 ;
  assign n4253 = \g3338_reg/NET0131  & \g35_pad  ;
  assign n4254 = \g13895_pad  & \g3303_reg/NET0131  ;
  assign n4255 = \g16603_pad  & \g16718_pad  ;
  assign n4256 = n4254 & n4255 ;
  assign n4257 = n4253 & n4256 ;
  assign n4258 = \g3343_reg/NET0131  & ~n4257 ;
  assign n4259 = \g1564_reg/NET0131  & ~\g35_pad  ;
  assign n4260 = \g1564_reg/NET0131  & n1461 ;
  assign n4261 = \g1559_reg/NET0131  & \g35_pad  ;
  assign n4262 = ~n4260 & n4261 ;
  assign n4263 = ~\g1554_reg/NET0131  & \g35_pad  ;
  assign n4264 = ~\g1559_reg/NET0131  & n4263 ;
  assign n4265 = n4260 & n4264 ;
  assign n4266 = ~n4262 & ~n4265 ;
  assign n4267 = ~n4259 & n4266 ;
  assign n4268 = \g2771_reg/NET0131  & ~\g35_pad  ;
  assign n4269 = n3534 & ~n4268 ;
  assign n4270 = \g2803_reg/NET0131  & ~\g35_pad  ;
  assign n4271 = n3595 & ~n4270 ;
  assign n4272 = n2521 & n2522 ;
  assign n4273 = n4085 & ~n4272 ;
  assign n4274 = \g4340_reg/NET0131  & \g4628_reg/NET0131  ;
  assign n4275 = n2520 & n4274 ;
  assign n4276 = \g35_pad  & ~n4275 ;
  assign n4277 = \g4349_reg/NET0131  & ~n4085 ;
  assign n4278 = ~n4276 & n4277 ;
  assign n4279 = ~n4273 & ~n4278 ;
  assign n4280 = \g305_reg/NET0131  & ~n2514 ;
  assign n4281 = \g35_pad  & n4280 ;
  assign n4282 = \g336_reg/NET0131  & \g35_pad  ;
  assign n4283 = ~n2515 & n4282 ;
  assign n4284 = ~n4281 & ~n4283 ;
  assign n4285 = \g311_reg/NET0131  & ~\g35_pad  ;
  assign n4286 = n4284 & ~n4285 ;
  assign n4287 = ~\g35_pad  & \g4311_reg/NET0131  ;
  assign n4288 = ~\g4322_reg/NET0131  & ~n4025 ;
  assign n4289 = ~n4026 & ~n4288 ;
  assign n4290 = n4022 & n4289 ;
  assign n4291 = ~n4287 & ~n4290 ;
  assign n4292 = \g14189_pad  & ~\g896_reg/NET0131  ;
  assign n4293 = n4057 & n4292 ;
  assign n4294 = \g35_pad  & n4293 ;
  assign n4295 = \g225_reg/NET0131  & \g35_pad  ;
  assign n4296 = ~n4061 & n4295 ;
  assign n4297 = ~n4294 & ~n4296 ;
  assign n4298 = ~\g35_pad  & \g872_reg/NET0131  ;
  assign n4299 = n4297 & ~n4298 ;
  assign n4300 = ~\g35_pad  & \g4653_reg/NET0131  ;
  assign n4301 = \g35_pad  & \g4659_reg/NET0131  ;
  assign n4302 = ~n2837 & n4301 ;
  assign n4303 = \g35_pad  & ~\g4659_reg/NET0131  ;
  assign n4304 = n2837 & n4303 ;
  assign n4305 = ~n4302 & ~n4304 ;
  assign n4306 = ~n4300 & n4305 ;
  assign n4307 = \g35_pad  & n2284 ;
  assign n4308 = \g35_pad  & n1923 ;
  assign n4309 = ~\g2667_reg/NET0131  & ~\g35_pad  ;
  assign n4310 = \g2661_reg/NET0131  & ~\g2667_reg/NET0131  ;
  assign n4311 = ~n1923 & n4310 ;
  assign n4312 = ~n4309 & ~n4311 ;
  assign n4313 = ~\g2661_reg/NET0131  & \g2667_reg/NET0131  ;
  assign n4314 = \g35_pad  & n4313 ;
  assign n4315 = ~n1923 & n4314 ;
  assign n4316 = ~\g2671_reg/NET0131  & \g35_pad  ;
  assign n4317 = n1923 & n4316 ;
  assign n4318 = ~n4315 & ~n4317 ;
  assign n4319 = n4312 & n4318 ;
  assign n4320 = \g2675_reg/NET0131  & \g35_pad  ;
  assign n4321 = n1923 & n4320 ;
  assign n4322 = ~\g2675_reg/NET0131  & \g35_pad  ;
  assign n4323 = ~n1923 & n4322 ;
  assign n4324 = ~n4321 & ~n4323 ;
  assign n4325 = \g2671_reg/NET0131  & ~\g35_pad  ;
  assign n4326 = n4324 & ~n4325 ;
  assign n4327 = \g14147_pad  & ~\g896_reg/NET0131  ;
  assign n4328 = n4057 & n4327 ;
  assign n4329 = \g35_pad  & n4328 ;
  assign n4330 = \g269_reg/NET0131  & \g35_pad  ;
  assign n4331 = ~n4061 & n4330 ;
  assign n4332 = ~n4329 & ~n4331 ;
  assign n4333 = \g239_reg/NET0131  & ~\g35_pad  ;
  assign n4334 = n4332 & ~n4333 ;
  assign n4335 = ~\g1706_reg/NET0131  & ~\g35_pad  ;
  assign n4336 = \g1700_reg/NET0131  & ~\g1706_reg/NET0131  ;
  assign n4337 = ~n2284 & n4336 ;
  assign n4338 = ~n4335 & ~n4337 ;
  assign n4339 = ~\g1700_reg/NET0131  & \g1706_reg/NET0131  ;
  assign n4340 = \g35_pad  & n4339 ;
  assign n4341 = ~n2284 & n4340 ;
  assign n4342 = ~\g1710_reg/NET0131  & \g35_pad  ;
  assign n4343 = n2284 & n4342 ;
  assign n4344 = ~n4341 & ~n4343 ;
  assign n4345 = n4338 & n4344 ;
  assign n4346 = ~\g2767_reg/NET0131  & n2963 ;
  assign n4347 = n2707 & n4346 ;
  assign n4348 = \g35_pad  & n4347 ;
  assign n4349 = n2707 & n2963 ;
  assign n4350 = \g2771_reg/NET0131  & \g35_pad  ;
  assign n4351 = ~n4349 & n4350 ;
  assign n4352 = ~n4348 & ~n4351 ;
  assign n4353 = \g2775_reg/NET0131  & ~\g35_pad  ;
  assign n4354 = n4352 & ~n4353 ;
  assign n4355 = \g2724_reg/NET0131  & ~\g2729_reg/NET0131  ;
  assign n4356 = ~\g2779_reg/NET0131  & n4355 ;
  assign n4357 = n2707 & n4356 ;
  assign n4358 = \g35_pad  & n4357 ;
  assign n4359 = n2707 & n4355 ;
  assign n4360 = \g2775_reg/NET0131  & \g35_pad  ;
  assign n4361 = ~n4359 & n4360 ;
  assign n4362 = ~n4358 & ~n4361 ;
  assign n4363 = \g2783_reg/NET0131  & ~\g35_pad  ;
  assign n4364 = n4362 & ~n4363 ;
  assign n4365 = ~\g2724_reg/NET0131  & ~\g2791_reg/NET0131  ;
  assign n4366 = \g2729_reg/NET0131  & n4365 ;
  assign n4367 = n2707 & n4366 ;
  assign n4368 = \g35_pad  & n4367 ;
  assign n4369 = ~\g2724_reg/NET0131  & \g2729_reg/NET0131  ;
  assign n4370 = n2707 & n4369 ;
  assign n4371 = \g2783_reg/NET0131  & \g35_pad  ;
  assign n4372 = ~n4370 & n4371 ;
  assign n4373 = ~n4368 & ~n4372 ;
  assign n4374 = \g2787_reg/NET0131  & ~\g35_pad  ;
  assign n4375 = n4373 & ~n4374 ;
  assign n4376 = \g2724_reg/NET0131  & ~\g2795_reg/NET0131  ;
  assign n4377 = \g2729_reg/NET0131  & n4376 ;
  assign n4378 = n2707 & n4377 ;
  assign n4379 = \g35_pad  & n4378 ;
  assign n4380 = \g2724_reg/NET0131  & \g2729_reg/NET0131  ;
  assign n4381 = n2707 & n4380 ;
  assign n4382 = \g2787_reg/NET0131  & \g35_pad  ;
  assign n4383 = ~n4381 & n4382 ;
  assign n4384 = ~n4379 & ~n4383 ;
  assign n4385 = \g2795_reg/NET0131  & ~\g35_pad  ;
  assign n4386 = n4384 & ~n4385 ;
  assign n4387 = \g1714_reg/NET0131  & \g35_pad  ;
  assign n4388 = n2284 & n4387 ;
  assign n4389 = ~\g1714_reg/NET0131  & \g35_pad  ;
  assign n4390 = ~n2284 & n4389 ;
  assign n4391 = ~n4388 & ~n4390 ;
  assign n4392 = \g1710_reg/NET0131  & ~\g35_pad  ;
  assign n4393 = n4391 & ~n4392 ;
  assign n4394 = ~\g2799_reg/NET0131  & n2963 ;
  assign n4395 = n2707 & n4394 ;
  assign n4396 = \g35_pad  & n4395 ;
  assign n4397 = \g2803_reg/NET0131  & \g35_pad  ;
  assign n4398 = ~n4349 & n4397 ;
  assign n4399 = ~n4396 & ~n4398 ;
  assign n4400 = \g2807_reg/NET0131  & ~\g35_pad  ;
  assign n4401 = n4399 & ~n4400 ;
  assign n4402 = ~\g2811_reg/NET0131  & n4355 ;
  assign n4403 = n2707 & n4402 ;
  assign n4404 = \g35_pad  & n4403 ;
  assign n4405 = \g2807_reg/NET0131  & \g35_pad  ;
  assign n4406 = ~n4359 & n4405 ;
  assign n4407 = ~n4404 & ~n4406 ;
  assign n4408 = \g2815_reg/NET0131  & ~\g35_pad  ;
  assign n4409 = n4407 & ~n4408 ;
  assign n4410 = ~\g2724_reg/NET0131  & ~\g2823_reg/NET0131  ;
  assign n4411 = \g2729_reg/NET0131  & n4410 ;
  assign n4412 = n2707 & n4411 ;
  assign n4413 = \g35_pad  & n4412 ;
  assign n4414 = \g2815_reg/NET0131  & \g35_pad  ;
  assign n4415 = ~n4370 & n4414 ;
  assign n4416 = ~n4413 & ~n4415 ;
  assign n4417 = \g2819_reg/NET0131  & ~\g35_pad  ;
  assign n4418 = n4416 & ~n4417 ;
  assign n4419 = \g2724_reg/NET0131  & ~\g2827_reg/NET0131  ;
  assign n4420 = \g2729_reg/NET0131  & n4419 ;
  assign n4421 = n2707 & n4420 ;
  assign n4422 = \g35_pad  & n4421 ;
  assign n4423 = \g2819_reg/NET0131  & \g35_pad  ;
  assign n4424 = ~n4381 & n4423 ;
  assign n4425 = ~n4422 & ~n4424 ;
  assign n4426 = \g2827_reg/NET0131  & ~\g35_pad  ;
  assign n4427 = n4425 & ~n4426 ;
  assign n4428 = \g35_pad  & n2069 ;
  assign n4429 = \g1816_reg/NET0131  & ~n4428 ;
  assign n4430 = \g1821_reg/NET0131  & \g35_pad  ;
  assign n4431 = n2069 & n4430 ;
  assign n4432 = ~n4429 & ~n4431 ;
  assign n4433 = ~\g1840_reg/NET0131  & ~\g35_pad  ;
  assign n4434 = \g1834_reg/NET0131  & ~\g1840_reg/NET0131  ;
  assign n4435 = ~n2069 & n4434 ;
  assign n4436 = ~n4433 & ~n4435 ;
  assign n4437 = ~\g1834_reg/NET0131  & \g1840_reg/NET0131  ;
  assign n4438 = \g35_pad  & n4437 ;
  assign n4439 = ~n2069 & n4438 ;
  assign n4440 = ~\g1844_reg/NET0131  & \g35_pad  ;
  assign n4441 = n2069 & n4440 ;
  assign n4442 = ~n4439 & ~n4441 ;
  assign n4443 = n4436 & n4442 ;
  assign n4444 = \g1848_reg/NET0131  & \g35_pad  ;
  assign n4445 = n2069 & n4444 ;
  assign n4446 = ~\g1848_reg/NET0131  & \g35_pad  ;
  assign n4447 = ~n2069 & n4446 ;
  assign n4448 = ~n4445 & ~n4447 ;
  assign n4449 = \g1844_reg/NET0131  & ~\g35_pad  ;
  assign n4450 = n4448 & ~n4449 ;
  assign n4451 = \g35_pad  & n2139 ;
  assign n4452 = \g1950_reg/NET0131  & ~n4451 ;
  assign n4453 = \g1955_reg/NET0131  & \g35_pad  ;
  assign n4454 = n2139 & n4453 ;
  assign n4455 = ~n4452 & ~n4454 ;
  assign n4456 = ~\g1974_reg/NET0131  & ~\g35_pad  ;
  assign n4457 = \g1968_reg/NET0131  & ~\g1974_reg/NET0131  ;
  assign n4458 = ~n2139 & n4457 ;
  assign n4459 = ~n4456 & ~n4458 ;
  assign n4460 = ~\g1968_reg/NET0131  & \g1974_reg/NET0131  ;
  assign n4461 = \g35_pad  & n4460 ;
  assign n4462 = ~n2139 & n4461 ;
  assign n4463 = ~\g1978_reg/NET0131  & \g35_pad  ;
  assign n4464 = n2139 & n4463 ;
  assign n4465 = ~n4462 & ~n4464 ;
  assign n4466 = n4459 & n4465 ;
  assign n4467 = \g1982_reg/NET0131  & \g35_pad  ;
  assign n4468 = n2139 & n4467 ;
  assign n4469 = ~\g1982_reg/NET0131  & \g35_pad  ;
  assign n4470 = ~n2139 & n4469 ;
  assign n4471 = ~n4468 & ~n4470 ;
  assign n4472 = \g1978_reg/NET0131  & ~\g35_pad  ;
  assign n4473 = n4471 & ~n4472 ;
  assign n4474 = \g35_pad  & n2209 ;
  assign n4475 = \g2084_reg/NET0131  & ~n4474 ;
  assign n4476 = \g2089_reg/NET0131  & \g35_pad  ;
  assign n4477 = n2209 & n4476 ;
  assign n4478 = ~n4475 & ~n4477 ;
  assign n4479 = ~\g2108_reg/NET0131  & ~\g35_pad  ;
  assign n4480 = \g2102_reg/NET0131  & ~\g2108_reg/NET0131  ;
  assign n4481 = ~n2209 & n4480 ;
  assign n4482 = ~n4479 & ~n4481 ;
  assign n4483 = ~\g2102_reg/NET0131  & \g2108_reg/NET0131  ;
  assign n4484 = \g35_pad  & n4483 ;
  assign n4485 = ~n2209 & n4484 ;
  assign n4486 = ~\g2112_reg/NET0131  & \g35_pad  ;
  assign n4487 = n2209 & n4486 ;
  assign n4488 = ~n4485 & ~n4487 ;
  assign n4489 = n4482 & n4488 ;
  assign n4490 = \g2116_reg/NET0131  & \g35_pad  ;
  assign n4491 = n2209 & n4490 ;
  assign n4492 = ~\g2116_reg/NET0131  & \g35_pad  ;
  assign n4493 = ~n2209 & n4492 ;
  assign n4494 = ~n4491 & ~n4493 ;
  assign n4495 = \g2112_reg/NET0131  & ~\g35_pad  ;
  assign n4496 = n4494 & ~n4495 ;
  assign n4497 = \g35_pad  & n1708 ;
  assign n4498 = \g2241_reg/NET0131  & ~n4497 ;
  assign n4499 = \g2246_reg/NET0131  & \g35_pad  ;
  assign n4500 = n1708 & n4499 ;
  assign n4501 = ~n4498 & ~n4500 ;
  assign n4502 = ~\g2265_reg/NET0131  & ~\g35_pad  ;
  assign n4503 = \g2259_reg/NET0131  & ~\g2265_reg/NET0131  ;
  assign n4504 = ~n1708 & n4503 ;
  assign n4505 = ~n4502 & ~n4504 ;
  assign n4506 = ~\g2259_reg/NET0131  & \g2265_reg/NET0131  ;
  assign n4507 = \g35_pad  & n4506 ;
  assign n4508 = ~n1708 & n4507 ;
  assign n4509 = ~\g2269_reg/NET0131  & \g35_pad  ;
  assign n4510 = n1708 & n4509 ;
  assign n4511 = ~n4508 & ~n4510 ;
  assign n4512 = n4505 & n4511 ;
  assign n4513 = \g2273_reg/NET0131  & \g35_pad  ;
  assign n4514 = n1708 & n4513 ;
  assign n4515 = ~\g2273_reg/NET0131  & \g35_pad  ;
  assign n4516 = ~n1708 & n4515 ;
  assign n4517 = ~n4514 & ~n4516 ;
  assign n4518 = \g2269_reg/NET0131  & ~\g35_pad  ;
  assign n4519 = n4517 & ~n4518 ;
  assign n4520 = \g35_pad  & n1778 ;
  assign n4521 = \g2375_reg/NET0131  & ~n4520 ;
  assign n4522 = \g2380_reg/NET0131  & \g35_pad  ;
  assign n4523 = n1778 & n4522 ;
  assign n4524 = ~n4521 & ~n4523 ;
  assign n4525 = ~\g2399_reg/NET0131  & ~\g35_pad  ;
  assign n4526 = \g2393_reg/NET0131  & ~\g2399_reg/NET0131  ;
  assign n4527 = ~n1778 & n4526 ;
  assign n4528 = ~n4525 & ~n4527 ;
  assign n4529 = ~\g2393_reg/NET0131  & \g2399_reg/NET0131  ;
  assign n4530 = \g35_pad  & n4529 ;
  assign n4531 = ~n1778 & n4530 ;
  assign n4532 = ~\g2403_reg/NET0131  & \g35_pad  ;
  assign n4533 = n1778 & n4532 ;
  assign n4534 = ~n4531 & ~n4533 ;
  assign n4535 = n4528 & n4534 ;
  assign n4536 = \g2407_reg/NET0131  & \g35_pad  ;
  assign n4537 = n1778 & n4536 ;
  assign n4538 = ~\g2407_reg/NET0131  & \g35_pad  ;
  assign n4539 = ~n1778 & n4538 ;
  assign n4540 = ~n4537 & ~n4539 ;
  assign n4541 = \g2403_reg/NET0131  & ~\g35_pad  ;
  assign n4542 = n4540 & ~n4541 ;
  assign n4543 = \g35_pad  & n1853 ;
  assign n4544 = \g2509_reg/NET0131  & ~n4543 ;
  assign n4545 = \g2514_reg/NET0131  & \g35_pad  ;
  assign n4546 = n1853 & n4545 ;
  assign n4547 = ~n4544 & ~n4546 ;
  assign n4548 = ~\g2533_reg/NET0131  & ~\g35_pad  ;
  assign n4549 = \g2527_reg/NET0131  & ~\g2533_reg/NET0131  ;
  assign n4550 = ~n1853 & n4549 ;
  assign n4551 = ~n4548 & ~n4550 ;
  assign n4552 = ~\g2527_reg/NET0131  & \g2533_reg/NET0131  ;
  assign n4553 = \g35_pad  & n4552 ;
  assign n4554 = ~n1853 & n4553 ;
  assign n4555 = ~\g2537_reg/NET0131  & \g35_pad  ;
  assign n4556 = n1853 & n4555 ;
  assign n4557 = ~n4554 & ~n4556 ;
  assign n4558 = n4551 & n4557 ;
  assign n4559 = \g2541_reg/NET0131  & \g35_pad  ;
  assign n4560 = n1853 & n4559 ;
  assign n4561 = ~\g2541_reg/NET0131  & \g35_pad  ;
  assign n4562 = ~n1853 & n4561 ;
  assign n4563 = ~n4560 & ~n4562 ;
  assign n4564 = \g2537_reg/NET0131  & ~\g35_pad  ;
  assign n4565 = n4563 & ~n4564 ;
  assign n4566 = \g2643_reg/NET0131  & ~n4308 ;
  assign n4567 = \g2648_reg/NET0131  & \g35_pad  ;
  assign n4568 = n1923 & n4567 ;
  assign n4569 = ~n4566 & ~n4568 ;
  assign n4570 = ~\g1636_reg/NET0131  & ~n2261 ;
  assign n4571 = ~\g1636_reg/NET0131  & \g17291_pad  ;
  assign n4572 = ~n2264 & n4571 ;
  assign n4573 = ~n4570 & ~n4572 ;
  assign n4574 = ~\g1592_reg/NET0131  & n4573 ;
  assign n4575 = \g1668_reg/NET0131  & ~n2261 ;
  assign n4576 = \g1668_reg/NET0131  & \g17291_pad  ;
  assign n4577 = ~n2264 & n4576 ;
  assign n4578 = ~n4575 & ~n4577 ;
  assign n4579 = \g35_pad  & n4578 ;
  assign n4580 = ~n4574 & n4579 ;
  assign n4581 = ~\g1008_reg/NET0131  & \g1036_reg/NET0131  ;
  assign n4582 = n4197 & n4581 ;
  assign n4583 = n2815 & n4582 ;
  assign n4584 = ~n2816 & n4583 ;
  assign n4585 = \g1046_reg/NET0131  & ~n2815 ;
  assign n4586 = ~n2816 & n3910 ;
  assign n4587 = ~n4585 & n4586 ;
  assign n4588 = ~n4584 & ~n4587 ;
  assign n4589 = ~n2815 & ~n2816 ;
  assign n4590 = \g969_reg/NET0131  & ~n4589 ;
  assign n4591 = n4588 & ~n4590 ;
  assign n4592 = \g35_pad  & ~n4591 ;
  assign n4593 = \g2763_reg/NET0131  & ~\g35_pad  ;
  assign n4594 = ~n2703 & ~n4593 ;
  assign n4595 = ~\g1632_reg/NET0131  & ~n2701 ;
  assign n4596 = ~n2707 & n4595 ;
  assign n4597 = ~\g2767_reg/NET0131  & ~n4593 ;
  assign n4598 = ~n4596 & n4597 ;
  assign n4599 = ~n4594 & ~n4598 ;
  assign n4600 = \g2767_reg/NET0131  & ~\g35_pad  ;
  assign n4601 = ~n2703 & ~n4600 ;
  assign n4602 = ~\g1768_reg/NET0131  & ~n2701 ;
  assign n4603 = ~n2707 & n4602 ;
  assign n4604 = ~\g2779_reg/NET0131  & ~n4600 ;
  assign n4605 = ~n4603 & n4604 ;
  assign n4606 = ~n4601 & ~n4605 ;
  assign n4607 = \g2779_reg/NET0131  & ~\g35_pad  ;
  assign n4608 = ~n2703 & ~n4607 ;
  assign n4609 = ~\g1902_reg/NET0131  & ~n2701 ;
  assign n4610 = ~n2707 & n4609 ;
  assign n4611 = ~\g2791_reg/NET0131  & ~n4607 ;
  assign n4612 = ~n4610 & n4611 ;
  assign n4613 = ~n4608 & ~n4612 ;
  assign n4614 = \g2791_reg/NET0131  & ~\g35_pad  ;
  assign n4615 = ~n2703 & ~n4614 ;
  assign n4616 = ~\g2036_reg/NET0131  & ~n2701 ;
  assign n4617 = ~n2707 & n4616 ;
  assign n4618 = ~\g2795_reg/NET0131  & ~n4614 ;
  assign n4619 = ~n4617 & n4618 ;
  assign n4620 = ~n4615 & ~n4619 ;
  assign n4621 = \g2799_reg/NET0131  & ~\g35_pad  ;
  assign n4622 = ~n2703 & ~n4621 ;
  assign n4623 = ~\g2327_reg/NET0131  & ~n2701 ;
  assign n4624 = ~n2707 & n4623 ;
  assign n4625 = ~\g2811_reg/NET0131  & ~n4621 ;
  assign n4626 = ~n4624 & n4625 ;
  assign n4627 = ~n4622 & ~n4626 ;
  assign n4628 = ~\g1002_reg/NET0131  & ~n3911 ;
  assign n4629 = n3908 & n4628 ;
  assign n4630 = ~n2816 & ~n4629 ;
  assign n4631 = \g1018_reg/NET0131  & \g35_pad  ;
  assign n4632 = ~n4630 & n4631 ;
  assign n4633 = ~\g1018_reg/NET0131  & ~n2816 ;
  assign n4634 = ~n3911 & n4633 ;
  assign n4635 = n3908 & n4634 ;
  assign n4636 = \g35_pad  & ~n4635 ;
  assign n4637 = \g1002_reg/NET0131  & ~n4636 ;
  assign n4638 = ~n4632 & ~n4637 ;
  assign n4639 = \g35_pad  & \g4793_reg/NET0131  ;
  assign n4640 = ~n2838 & n4639 ;
  assign n4641 = \g35_pad  & ~\g4793_reg/NET0131  ;
  assign n4642 = n2838 & n4641 ;
  assign n4643 = ~n4640 & ~n4642 ;
  assign n4644 = \g174_reg/NET0131  & \g182_reg/NET0131  ;
  assign n4645 = ~\g168_reg/NET0131  & ~n4644 ;
  assign n4646 = \g35_pad  & ~n2345 ;
  assign n4647 = n2344 & n4646 ;
  assign n4648 = ~n4645 & n4647 ;
  assign n4649 = \g1189_reg/NET0131  & ~\g35_pad  ;
  assign n4650 = \g1070_reg/NET0131  & n4217 ;
  assign n4651 = \g1193_reg/NET0131  & ~n4650 ;
  assign n4652 = \g35_pad  & n4651 ;
  assign n4653 = ~\g1193_reg/NET0131  & \g35_pad  ;
  assign n4654 = ~n4201 & n4653 ;
  assign n4655 = ~n4652 & ~n4654 ;
  assign n4656 = ~n4649 & n4655 ;
  assign n4657 = \g29218_pad  & ~\g35_pad  ;
  assign n4658 = ~\g4349_reg/NET0131  & ~\g4358_reg/NET0131  ;
  assign n4659 = n883 & n4658 ;
  assign n4660 = \g35_pad  & ~\g4332_reg/NET0131  ;
  assign n4661 = ~\g4340_reg/NET0131  & \g4643_reg/NET0131  ;
  assign n4662 = n4660 & n4661 ;
  assign n4663 = n4659 & n4662 ;
  assign n4664 = ~n4657 & ~n4663 ;
  assign n4665 = \g2811_reg/NET0131  & ~\g35_pad  ;
  assign n4666 = ~n2703 & ~n4665 ;
  assign n4667 = ~\g2461_reg/NET0131  & ~n2701 ;
  assign n4668 = ~n2707 & n4667 ;
  assign n4669 = ~\g2823_reg/NET0131  & ~n4665 ;
  assign n4670 = ~n4668 & n4669 ;
  assign n4671 = ~n4666 & ~n4670 ;
  assign n4672 = \g2823_reg/NET0131  & ~\g35_pad  ;
  assign n4673 = ~n2703 & ~n4672 ;
  assign n4674 = ~\g2595_reg/NET0131  & ~n2701 ;
  assign n4675 = ~n2707 & n4674 ;
  assign n4676 = ~\g2827_reg/NET0131  & ~n4672 ;
  assign n4677 = ~n4675 & n4676 ;
  assign n4678 = ~n4673 & ~n4677 ;
  assign n4679 = ~\g2927_reg/NET0131  & ~\g35_pad  ;
  assign n4680 = \g35_pad  & ~\g4072_reg/NET0131  ;
  assign n4681 = ~\g2941_reg/NET0131  & ~\g4153_reg/NET0131  ;
  assign n4682 = n4680 & n4681 ;
  assign n4683 = ~n4679 & ~n4682 ;
  assign n4684 = \g1193_reg/NET0131  & ~\g35_pad  ;
  assign n4685 = \g7916_pad  & n1386 ;
  assign n4686 = ~n4214 & n4685 ;
  assign n4687 = ~\g1199_reg/NET0131  & ~n4686 ;
  assign n4688 = n4218 & ~n4687 ;
  assign n4689 = ~n4213 & n4688 ;
  assign n4690 = ~n4684 & ~n4689 ;
  assign n4691 = \g3329_reg/NET0131  & ~\g35_pad  ;
  assign n4692 = n4253 & ~n4256 ;
  assign n4693 = ~\g3338_reg/NET0131  & \g35_pad  ;
  assign n4694 = n4256 & n4693 ;
  assign n4695 = ~n4692 & ~n4694 ;
  assign n4696 = ~n4691 & n4695 ;
  assign n4697 = \g847_reg/NET0131  & n2579 ;
  assign n4698 = \g35_pad  & ~\g843_reg/NET0131  ;
  assign n4699 = ~n4697 & n4698 ;
  assign n4700 = \g35_pad  & \g843_reg/NET0131  ;
  assign n4701 = n4697 & n4700 ;
  assign n4702 = ~n4699 & ~n4701 ;
  assign n4703 = \g837_reg/NET0131  & n4702 ;
  assign n4704 = ~\g4584_reg/NET0131  & ~n4021 ;
  assign n4705 = \g35_pad  & ~n2532 ;
  assign n4706 = ~n4704 & n4705 ;
  assign n4707 = ~\g35_pad  & \g4332_reg/NET0131  ;
  assign n4708 = ~n4706 & ~n4707 ;
  assign n4709 = ~\g2856_reg/NET0131  & n797 ;
  assign n4710 = \g35_pad  & ~n4709 ;
  assign n4711 = \g2848_reg/NET0131  & ~\g35_pad  ;
  assign n4712 = ~n790 & ~n4711 ;
  assign n4713 = ~n4710 & n4712 ;
  assign n4714 = ~\g5037_reg/NET0131  & n4141 ;
  assign n4715 = \g5037_reg/NET0131  & n4147 ;
  assign n4716 = ~n4714 & ~n4715 ;
  assign n4717 = \g35_pad  & ~\g5041_reg/NET0131  ;
  assign n4718 = ~n4716 & n4717 ;
  assign n4719 = ~n4154 & ~n4233 ;
  assign n4720 = \g35_pad  & \g5041_reg/NET0131  ;
  assign n4721 = n4719 & n4720 ;
  assign n4722 = n4716 & n4721 ;
  assign n4723 = ~n4718 & ~n4722 ;
  assign n4724 = ~\g35_pad  & \g5037_reg/NET0131  ;
  assign n4725 = n4723 & ~n4724 ;
  assign n4726 = ~\g2882_reg/NET0131  & n813 ;
  assign n4727 = \g35_pad  & ~n4726 ;
  assign n4728 = \g2898_reg/NET0131  & ~\g35_pad  ;
  assign n4729 = ~n806 & ~n4728 ;
  assign n4730 = ~n4727 & n4729 ;
  assign n4731 = n827 & n954 ;
  assign n4732 = \g4646_reg/NET0131  & n4731 ;
  assign n4733 = ~n868 & n4732 ;
  assign n4734 = \g35_pad  & ~n4733 ;
  assign n4735 = \g4646_reg/NET0131  & \g5128_reg/NET0131  ;
  assign n4736 = n4731 & n4735 ;
  assign n4737 = ~n868 & n4736 ;
  assign n4738 = \g35_pad  & ~n4737 ;
  assign n4739 = ~\g5134_reg/NET0131  & ~n4738 ;
  assign n4740 = ~\g5128_reg/NET0131  & \g5134_reg/NET0131  ;
  assign n4741 = \g4646_reg/NET0131  & n4740 ;
  assign n4742 = n4731 & n4741 ;
  assign n4743 = ~n868 & n4742 ;
  assign n4744 = \g35_pad  & n4743 ;
  assign n4745 = \g35_pad  & ~\g5138_reg/NET0131  ;
  assign n4746 = ~n4733 & n4745 ;
  assign n4747 = ~n4744 & ~n4746 ;
  assign n4748 = ~n4739 & n4747 ;
  assign n4749 = \g35_pad  & \g5142_reg/NET0131  ;
  assign n4750 = ~n4733 & n4749 ;
  assign n4751 = \g35_pad  & ~\g5142_reg/NET0131  ;
  assign n4752 = n4733 & n4751 ;
  assign n4753 = ~n4750 & ~n4752 ;
  assign n4754 = ~\g35_pad  & \g5138_reg/NET0131  ;
  assign n4755 = n4753 & ~n4754 ;
  assign n4756 = \g1772_reg/NET0131  & n1600 ;
  assign n4757 = ~n1620 & n4756 ;
  assign n4758 = n2080 & ~n4757 ;
  assign n4759 = \g35_pad  & ~n4758 ;
  assign n4760 = \g1779_reg/NET0131  & ~\g35_pad  ;
  assign n4761 = ~n4759 & ~n4760 ;
  assign n4762 = \g35_pad  & n1600 ;
  assign n4763 = ~n1620 & n4762 ;
  assign n4764 = \g1772_reg/NET0131  & ~n4763 ;
  assign n4765 = \g1802_reg/NET0131  & \g35_pad  ;
  assign n4766 = n1600 & n4765 ;
  assign n4767 = ~n1620 & n4766 ;
  assign n4768 = ~n4764 & ~n4767 ;
  assign n4769 = \g3352_reg/NET0131  & \g4674_reg/NET0131  ;
  assign n4770 = \g3288_reg/NET0131  & n954 ;
  assign n4771 = n4769 & n4770 ;
  assign n4772 = ~n2618 & n4771 ;
  assign n4773 = \g35_pad  & ~n4772 ;
  assign n4774 = ~\g3125_reg/NET0131  & ~\g35_pad  ;
  assign n4775 = \g3119_reg/NET0131  & ~\g3125_reg/NET0131  ;
  assign n4776 = n4772 & n4775 ;
  assign n4777 = ~n4774 & ~n4776 ;
  assign n4778 = ~\g3119_reg/NET0131  & \g3125_reg/NET0131  ;
  assign n4779 = \g35_pad  & n4778 ;
  assign n4780 = n4772 & n4779 ;
  assign n4781 = ~\g3129_reg/NET0131  & \g35_pad  ;
  assign n4782 = ~n4772 & n4781 ;
  assign n4783 = ~n4780 & ~n4782 ;
  assign n4784 = n4777 & n4783 ;
  assign n4785 = ~\g3155_reg/NET0131  & ~\g3161_reg/NET0131  ;
  assign n4786 = ~\g3167_reg/NET0131  & n4785 ;
  assign n4787 = ~\g3171_reg/NET0131  & ~\g3179_reg/NET0131  ;
  assign n4788 = \g4180_reg/NET0131  & ~\g4284_reg/NET0131  ;
  assign n4789 = n4787 & ~n4788 ;
  assign n4790 = n4786 & n4789 ;
  assign n4791 = \g35_pad  & n4790 ;
  assign n4792 = n4786 & n4787 ;
  assign n4793 = \g3187_reg/NET0131  & \g35_pad  ;
  assign n4794 = ~n4792 & n4793 ;
  assign n4795 = ~n4791 & ~n4794 ;
  assign n4796 = \g3179_reg/NET0131  & ~\g35_pad  ;
  assign n4797 = n4795 & ~n4796 ;
  assign n4798 = \g3171_reg/NET0131  & ~\g3179_reg/NET0131  ;
  assign n4799 = ~n4788 & n4798 ;
  assign n4800 = n4786 & n4799 ;
  assign n4801 = \g35_pad  & n4800 ;
  assign n4802 = n4786 & n4798 ;
  assign n4803 = \g3191_reg/NET0131  & \g35_pad  ;
  assign n4804 = ~n4802 & n4803 ;
  assign n4805 = ~n4801 & ~n4804 ;
  assign n4806 = \g3195_reg/NET0131  & ~\g35_pad  ;
  assign n4807 = n4805 & ~n4806 ;
  assign n4808 = \g3133_reg/NET0131  & \g35_pad  ;
  assign n4809 = ~n4772 & n4808 ;
  assign n4810 = ~\g3133_reg/NET0131  & \g35_pad  ;
  assign n4811 = n4772 & n4810 ;
  assign n4812 = ~n4809 & ~n4811 ;
  assign n4813 = \g3129_reg/NET0131  & ~\g35_pad  ;
  assign n4814 = n4812 & ~n4813 ;
  assign n4815 = \g3167_reg/NET0131  & n4787 ;
  assign n4816 = \g3195_reg/NET0131  & \g35_pad  ;
  assign n4817 = ~n4815 & n4816 ;
  assign n4818 = \g35_pad  & ~n4788 ;
  assign n4819 = n4815 & n4818 ;
  assign n4820 = ~n4817 & ~n4819 ;
  assign n4821 = \g3247_reg/NET0131  & ~\g35_pad  ;
  assign n4822 = n4820 & ~n4821 ;
  assign n4823 = ~\g3171_reg/NET0131  & \g3179_reg/NET0131  ;
  assign n4824 = ~n4788 & n4823 ;
  assign n4825 = n4786 & n4824 ;
  assign n4826 = \g35_pad  & n4825 ;
  assign n4827 = n4786 & n4823 ;
  assign n4828 = \g3199_reg/NET0131  & \g35_pad  ;
  assign n4829 = ~n4827 & n4828 ;
  assign n4830 = ~n4826 & ~n4829 ;
  assign n4831 = \g3203_reg/NET0131  & ~\g35_pad  ;
  assign n4832 = n4830 & ~n4831 ;
  assign n4833 = \g3167_reg/NET0131  & n4798 ;
  assign n4834 = \g3203_reg/NET0131  & \g35_pad  ;
  assign n4835 = ~n4833 & n4834 ;
  assign n4836 = n4818 & n4833 ;
  assign n4837 = ~n4835 & ~n4836 ;
  assign n4838 = \g3251_reg/NET0131  & ~\g35_pad  ;
  assign n4839 = n4837 & ~n4838 ;
  assign n4840 = \g3155_reg/NET0131  & ~\g3161_reg/NET0131  ;
  assign n4841 = n4787 & n4840 ;
  assign n4842 = \g3215_reg/NET0131  & \g35_pad  ;
  assign n4843 = ~n4841 & n4842 ;
  assign n4844 = n4818 & n4841 ;
  assign n4845 = ~n4843 & ~n4844 ;
  assign n4846 = \g3187_reg/NET0131  & ~\g35_pad  ;
  assign n4847 = n4845 & ~n4846 ;
  assign n4848 = n4798 & n4840 ;
  assign n4849 = \g3219_reg/NET0131  & \g35_pad  ;
  assign n4850 = ~n4848 & n4849 ;
  assign n4851 = n4818 & n4848 ;
  assign n4852 = ~n4850 & ~n4851 ;
  assign n4853 = \g3191_reg/NET0131  & ~\g35_pad  ;
  assign n4854 = n4852 & ~n4853 ;
  assign n4855 = n4823 & n4840 ;
  assign n4856 = \g3223_reg/NET0131  & \g35_pad  ;
  assign n4857 = ~n4855 & n4856 ;
  assign n4858 = n4818 & n4855 ;
  assign n4859 = ~n4857 & ~n4858 ;
  assign n4860 = \g3199_reg/NET0131  & ~\g35_pad  ;
  assign n4861 = n4859 & ~n4860 ;
  assign n4862 = ~\g3155_reg/NET0131  & \g3161_reg/NET0131  ;
  assign n4863 = n4787 & n4862 ;
  assign n4864 = \g3231_reg/NET0131  & \g35_pad  ;
  assign n4865 = ~n4863 & n4864 ;
  assign n4866 = n4818 & n4863 ;
  assign n4867 = ~n4865 & ~n4866 ;
  assign n4868 = \g3215_reg/NET0131  & ~\g35_pad  ;
  assign n4869 = n4867 & ~n4868 ;
  assign n4870 = n4798 & n4862 ;
  assign n4871 = \g3235_reg/NET0131  & \g35_pad  ;
  assign n4872 = ~n4870 & n4871 ;
  assign n4873 = n4818 & n4870 ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4875 = \g3219_reg/NET0131  & ~\g35_pad  ;
  assign n4876 = n4874 & ~n4875 ;
  assign n4877 = n4823 & n4862 ;
  assign n4878 = \g3239_reg/NET0131  & \g35_pad  ;
  assign n4879 = ~n4877 & n4878 ;
  assign n4880 = n4818 & n4877 ;
  assign n4881 = ~n4879 & ~n4880 ;
  assign n4882 = \g3223_reg/NET0131  & ~\g35_pad  ;
  assign n4883 = n4881 & ~n4882 ;
  assign n4884 = \g3155_reg/NET0131  & \g3161_reg/NET0131  ;
  assign n4885 = n4787 & n4884 ;
  assign n4886 = \g3247_reg/NET0131  & \g35_pad  ;
  assign n4887 = ~n4885 & n4886 ;
  assign n4888 = n4818 & n4885 ;
  assign n4889 = ~n4887 & ~n4888 ;
  assign n4890 = \g3231_reg/NET0131  & ~\g35_pad  ;
  assign n4891 = n4889 & ~n4890 ;
  assign n4892 = n4798 & n4884 ;
  assign n4893 = \g3251_reg/NET0131  & \g35_pad  ;
  assign n4894 = ~n4892 & n4893 ;
  assign n4895 = n4818 & n4892 ;
  assign n4896 = ~n4894 & ~n4895 ;
  assign n4897 = \g3235_reg/NET0131  & ~\g35_pad  ;
  assign n4898 = n4896 & ~n4897 ;
  assign n4899 = \g3171_reg/NET0131  & \g3179_reg/NET0131  ;
  assign n4900 = ~n4788 & n4899 ;
  assign n4901 = n4786 & n4900 ;
  assign n4902 = \g35_pad  & n4901 ;
  assign n4903 = n4786 & n4899 ;
  assign n4904 = \g3207_reg/NET0131  & \g35_pad  ;
  assign n4905 = ~n4903 & n4904 ;
  assign n4906 = ~n4902 & ~n4905 ;
  assign n4907 = \g3211_reg/NET0131  & ~\g35_pad  ;
  assign n4908 = n4906 & ~n4907 ;
  assign n4909 = \g3167_reg/NET0131  & n4823 ;
  assign n4910 = \g3211_reg/NET0131  & \g35_pad  ;
  assign n4911 = ~n4909 & n4910 ;
  assign n4912 = n4818 & n4909 ;
  assign n4913 = ~n4911 & ~n4912 ;
  assign n4914 = \g3255_reg/NET0131  & ~\g35_pad  ;
  assign n4915 = n4913 & ~n4914 ;
  assign n4916 = n4840 & n4899 ;
  assign n4917 = \g3227_reg/NET0131  & \g35_pad  ;
  assign n4918 = ~n4916 & n4917 ;
  assign n4919 = n4818 & n4916 ;
  assign n4920 = ~n4918 & ~n4919 ;
  assign n4921 = \g3207_reg/NET0131  & ~\g35_pad  ;
  assign n4922 = n4920 & ~n4921 ;
  assign n4923 = n4862 & n4899 ;
  assign n4924 = \g3243_reg/NET0131  & \g35_pad  ;
  assign n4925 = ~n4923 & n4924 ;
  assign n4926 = n4818 & n4923 ;
  assign n4927 = ~n4925 & ~n4926 ;
  assign n4928 = \g3227_reg/NET0131  & ~\g35_pad  ;
  assign n4929 = n4927 & ~n4928 ;
  assign n4930 = n4823 & n4884 ;
  assign n4931 = \g3255_reg/NET0131  & \g35_pad  ;
  assign n4932 = ~n4930 & n4931 ;
  assign n4933 = n4818 & n4930 ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = \g3239_reg/NET0131  & ~\g35_pad  ;
  assign n4936 = n4934 & ~n4935 ;
  assign n4937 = n4884 & n4899 ;
  assign n4938 = \g3259_reg/NET0131  & \g35_pad  ;
  assign n4939 = ~n4937 & n4938 ;
  assign n4940 = n4818 & n4937 ;
  assign n4941 = ~n4939 & ~n4940 ;
  assign n4942 = \g3243_reg/NET0131  & ~\g35_pad  ;
  assign n4943 = n4941 & ~n4942 ;
  assign n4944 = \g3167_reg/NET0131  & n4899 ;
  assign n4945 = \g3263_reg/NET0131  & \g35_pad  ;
  assign n4946 = ~n4944 & n4945 ;
  assign n4947 = n4818 & n4944 ;
  assign n4948 = ~n4946 & ~n4947 ;
  assign n4949 = \g3259_reg/NET0131  & ~\g35_pad  ;
  assign n4950 = n4948 & ~n4949 ;
  assign n4951 = \g1906_reg/NET0131  & n1628 ;
  assign n4952 = ~n1644 & n4951 ;
  assign n4953 = n2163 & ~n4952 ;
  assign n4954 = \g35_pad  & ~n4953 ;
  assign n4955 = \g1913_reg/NET0131  & ~\g35_pad  ;
  assign n4956 = ~n4954 & ~n4955 ;
  assign n4957 = \g35_pad  & n1628 ;
  assign n4958 = ~n1644 & n4957 ;
  assign n4959 = \g1906_reg/NET0131  & ~n4958 ;
  assign n4960 = \g1936_reg/NET0131  & \g35_pad  ;
  assign n4961 = n1628 & n4960 ;
  assign n4962 = ~n1644 & n4961 ;
  assign n4963 = ~n4959 & ~n4962 ;
  assign n4964 = \g35_pad  & ~n2456 ;
  assign n4965 = \g29213_pad  & \g35_pad  ;
  assign n4966 = ~\g5097_reg/NET0131  & n4965 ;
  assign n4967 = \g5084_reg/NET0131  & \g5092_reg/NET0131  ;
  assign n4968 = n4965 & ~n4967 ;
  assign n4969 = ~n4966 & ~n4968 ;
  assign n4970 = \g35_pad  & ~n4967 ;
  assign n4971 = \g5097_reg/NET0131  & ~n4965 ;
  assign n4972 = ~n4970 & n4971 ;
  assign n4973 = n4969 & ~n4972 ;
  assign n4974 = \g3639_reg/NET0131  & \g3703_reg/NET0131  ;
  assign n4975 = n954 & n4974 ;
  assign n4976 = \g3470_reg/NET0131  & \g4681_reg/NET0131  ;
  assign n4977 = n4975 & n4976 ;
  assign n4978 = ~n2646 & n4977 ;
  assign n4979 = \g35_pad  & ~n4978 ;
  assign n4980 = ~\g3476_reg/NET0131  & ~n4979 ;
  assign n4981 = ~\g3470_reg/NET0131  & \g3476_reg/NET0131  ;
  assign n4982 = \g4681_reg/NET0131  & n4981 ;
  assign n4983 = n4975 & n4982 ;
  assign n4984 = ~n2646 & n4983 ;
  assign n4985 = \g35_pad  & n4984 ;
  assign n4986 = \g4681_reg/NET0131  & n4975 ;
  assign n4987 = ~n2646 & n4986 ;
  assign n4988 = ~\g3480_reg/NET0131  & \g35_pad  ;
  assign n4989 = ~n4987 & n4988 ;
  assign n4990 = ~n4985 & ~n4989 ;
  assign n4991 = ~n4980 & n4990 ;
  assign n4992 = \g3484_reg/NET0131  & \g35_pad  ;
  assign n4993 = ~n4987 & n4992 ;
  assign n4994 = ~\g3484_reg/NET0131  & \g35_pad  ;
  assign n4995 = n4987 & n4994 ;
  assign n4996 = ~n4993 & ~n4995 ;
  assign n4997 = \g3480_reg/NET0131  & ~\g35_pad  ;
  assign n4998 = n4996 & ~n4997 ;
  assign n4999 = \g2040_reg/NET0131  & n1652 ;
  assign n5000 = ~n1668 & n4999 ;
  assign n5001 = n2193 & ~n5000 ;
  assign n5002 = \g35_pad  & ~n5001 ;
  assign n5003 = \g2047_reg/NET0131  & ~\g35_pad  ;
  assign n5004 = ~n5002 & ~n5003 ;
  assign n5005 = \g35_pad  & n1652 ;
  assign n5006 = ~n1668 & n5005 ;
  assign n5007 = \g3990_reg/NET0131  & n954 ;
  assign n5008 = \g4054_reg/NET0131  & \g4688_reg/NET0131  ;
  assign n5009 = n5007 & n5008 ;
  assign n5010 = ~n951 & n5009 ;
  assign n5011 = \g35_pad  & ~n5010 ;
  assign n5012 = ~\g35_pad  & ~\g3827_reg/NET0131  ;
  assign n5013 = \g3821_reg/NET0131  & ~\g3827_reg/NET0131  ;
  assign n5014 = n5010 & n5013 ;
  assign n5015 = ~n5012 & ~n5014 ;
  assign n5016 = ~\g3821_reg/NET0131  & \g3827_reg/NET0131  ;
  assign n5017 = \g35_pad  & n5016 ;
  assign n5018 = n5010 & n5017 ;
  assign n5019 = \g35_pad  & ~\g3831_reg/NET0131  ;
  assign n5020 = ~n5010 & n5019 ;
  assign n5021 = ~n5018 & ~n5020 ;
  assign n5022 = n5015 & n5021 ;
  assign n5023 = \g35_pad  & \g3835_reg/NET0131  ;
  assign n5024 = ~n5010 & n5023 ;
  assign n5025 = \g35_pad  & ~\g3835_reg/NET0131  ;
  assign n5026 = n5010 & n5025 ;
  assign n5027 = ~n5024 & ~n5026 ;
  assign n5028 = ~\g35_pad  & \g3831_reg/NET0131  ;
  assign n5029 = n5027 & ~n5028 ;
  assign n5030 = \g2197_reg/NET0131  & n1471 ;
  assign n5031 = ~n1491 & n5030 ;
  assign n5032 = n1732 & ~n5031 ;
  assign n5033 = \g35_pad  & ~n5032 ;
  assign n5034 = \g2204_reg/NET0131  & ~\g35_pad  ;
  assign n5035 = ~n5033 & ~n5034 ;
  assign n5036 = \g35_pad  & n1471 ;
  assign n5037 = ~n1491 & n5036 ;
  assign n5038 = \g2197_reg/NET0131  & ~n5037 ;
  assign n5039 = \g2227_reg/NET0131  & \g35_pad  ;
  assign n5040 = n1471 & n5039 ;
  assign n5041 = ~n1491 & n5040 ;
  assign n5042 = ~n5038 & ~n5041 ;
  assign n5043 = \g4258_reg/NET0131  & \g4264_reg/NET0131  ;
  assign n5044 = \g35_pad  & \g4273_reg/NET0131  ;
  assign n5045 = ~n5043 & n5044 ;
  assign n5046 = \g35_pad  & ~\g4269_reg/NET0131  ;
  assign n5047 = \g4273_reg/NET0131  & n5046 ;
  assign n5048 = ~n5045 & ~n5047 ;
  assign n5049 = \g35_pad  & ~n5043 ;
  assign n5050 = \g4269_reg/NET0131  & ~n5044 ;
  assign n5051 = ~n5049 & n5050 ;
  assign n5052 = n5048 & ~n5051 ;
  assign n5053 = \g35_pad  & \g4349_reg/NET0131  ;
  assign n5054 = \g4340_reg/NET0131  & n5053 ;
  assign n5055 = n2521 & n5054 ;
  assign n5056 = \g35_pad  & ~\g4349_reg/NET0131  ;
  assign n5057 = ~n2521 & n5056 ;
  assign n5058 = ~\g35_pad  & ~\g4340_reg/NET0131  ;
  assign n5059 = ~n4078 & ~n5058 ;
  assign n5060 = ~n5057 & n5059 ;
  assign n5061 = ~n5055 & n5060 ;
  assign n5062 = \g2331_reg/NET0131  & n1499 ;
  assign n5063 = ~n1515 & n5062 ;
  assign n5064 = n1802 & ~n5063 ;
  assign n5065 = \g35_pad  & ~n5064 ;
  assign n5066 = \g2338_reg/NET0131  & ~\g35_pad  ;
  assign n5067 = ~n5065 & ~n5066 ;
  assign n5068 = \g35_pad  & n1499 ;
  assign n5069 = ~n1515 & n5068 ;
  assign n5070 = \g2331_reg/NET0131  & ~n5069 ;
  assign n5071 = \g2361_reg/NET0131  & \g35_pad  ;
  assign n5072 = n1499 & n5071 ;
  assign n5073 = ~n1515 & n5072 ;
  assign n5074 = ~n5070 & ~n5073 ;
  assign n5075 = \g14125_pad  & ~\g896_reg/NET0131  ;
  assign n5076 = n4057 & n5075 ;
  assign n5077 = \g35_pad  & n5076 ;
  assign n5078 = \g239_reg/NET0131  & \g35_pad  ;
  assign n5079 = ~n4061 & n5078 ;
  assign n5080 = ~n5077 & ~n5079 ;
  assign n5081 = \g262_reg/NET0131  & ~\g35_pad  ;
  assign n5082 = n5080 & ~n5081 ;
  assign n5083 = \g35_pad  & ~n4987 ;
  assign n5084 = \g2465_reg/NET0131  & n1523 ;
  assign n5085 = ~n1539 & n5084 ;
  assign n5086 = n1877 & ~n5085 ;
  assign n5087 = \g35_pad  & ~n5086 ;
  assign n5088 = \g2472_reg/NET0131  & ~\g35_pad  ;
  assign n5089 = ~n5087 & ~n5088 ;
  assign n5090 = \g35_pad  & n1523 ;
  assign n5091 = ~n1539 & n5090 ;
  assign n5092 = \g2465_reg/NET0131  & ~n5091 ;
  assign n5093 = \g2495_reg/NET0131  & \g35_pad  ;
  assign n5094 = n1523 & n5093 ;
  assign n5095 = ~n1539 & n5094 ;
  assign n5096 = ~n5092 & ~n5095 ;
  assign n5097 = ~\g35_pad  & ~\g528_reg/NET0131  ;
  assign n5098 = n3991 & ~n3992 ;
  assign n5099 = \g35_pad  & ~n3993 ;
  assign n5100 = ~\g482_reg/NET0131  & n5099 ;
  assign n5101 = ~n5098 & n5100 ;
  assign n5102 = \g482_reg/NET0131  & n5099 ;
  assign n5103 = n5098 & n5102 ;
  assign n5104 = ~n5101 & ~n5103 ;
  assign n5105 = ~n5097 & n5104 ;
  assign n5106 = \g17291_pad  & ~n2264 ;
  assign n5107 = \g1636_reg/NET0131  & n2261 ;
  assign n5108 = ~n5106 & n5107 ;
  assign n5109 = n2267 & ~n5108 ;
  assign n5110 = \g35_pad  & ~n5109 ;
  assign n5111 = \g1644_reg/NET0131  & ~\g35_pad  ;
  assign n5112 = ~n5110 & ~n5111 ;
  assign n5113 = ~\g2555_reg/NET0131  & ~n1547 ;
  assign n5114 = \g1430_reg/NET0131  & ~\g2555_reg/NET0131  ;
  assign n5115 = ~n1550 & n5114 ;
  assign n5116 = ~n5113 & ~n5115 ;
  assign n5117 = ~\g2599_reg/NET0131  & n1547 ;
  assign n5118 = ~n1563 & n5117 ;
  assign n5119 = n5116 & ~n5118 ;
  assign n5120 = \g35_pad  & ~n5119 ;
  assign n5121 = ~\g2606_reg/NET0131  & ~\g35_pad  ;
  assign n5122 = ~n5120 & ~n5121 ;
  assign n5123 = \g35_pad  & n2261 ;
  assign n5124 = ~n5106 & n5123 ;
  assign n5125 = \g1636_reg/NET0131  & ~n5124 ;
  assign n5126 = \g1668_reg/NET0131  & \g35_pad  ;
  assign n5127 = n2261 & n5126 ;
  assign n5128 = ~n5106 & n5127 ;
  assign n5129 = ~n5125 & ~n5128 ;
  assign n5130 = \g35_pad  & n1547 ;
  assign n5131 = ~n1563 & n5130 ;
  assign n5132 = \g3111_reg/NET0131  & \g35_pad  ;
  assign n5133 = ~\g5115_reg/NET0131  & ~n5132 ;
  assign n5134 = \g5115_reg/NET0131  & n5132 ;
  assign n5135 = ~n5133 & ~n5134 ;
  assign n5136 = ~n4734 & ~n5135 ;
  assign n5137 = \g35_pad  & ~\g5124_reg/NET0131  ;
  assign n5138 = ~n4733 & n5137 ;
  assign n5139 = ~n5136 & ~n5138 ;
  assign n5140 = ~\g3106_reg/NET0131  & ~n5132 ;
  assign n5141 = \g3106_reg/NET0131  & n5132 ;
  assign n5142 = ~n5140 & ~n5141 ;
  assign n5143 = ~n4773 & ~n5142 ;
  assign n5144 = ~\g3115_reg/NET0131  & \g35_pad  ;
  assign n5145 = ~n4772 & n5144 ;
  assign n5146 = ~n5143 & ~n5145 ;
  assign n5147 = ~\g336_reg/NET0131  & ~\g35_pad  ;
  assign n5148 = ~\g311_reg/NET0131  & \g324_reg/NET0131  ;
  assign n5149 = ~\g305_reg/NET0131  & \g35_pad  ;
  assign n5150 = ~n5148 & n5149 ;
  assign n5151 = ~n5147 & ~n5150 ;
  assign n5152 = ~\g661_reg/NET0131  & n2579 ;
  assign n5153 = n2918 & n5152 ;
  assign n5154 = \g35_pad  & ~n5153 ;
  assign n5155 = ~\g728_reg/NET0131  & ~n5154 ;
  assign n5156 = ~\g29212_pad  & \g35_pad  ;
  assign n5157 = ~n2919 & n5156 ;
  assign n5158 = ~n5155 & ~n5157 ;
  assign n5159 = ~\g3457_reg/NET0131  & ~n5132 ;
  assign n5160 = \g3457_reg/NET0131  & n5132 ;
  assign n5161 = ~n5159 & ~n5160 ;
  assign n5162 = ~n5083 & ~n5161 ;
  assign n5163 = ~\g3466_reg/NET0131  & \g35_pad  ;
  assign n5164 = ~n4987 & n5163 ;
  assign n5165 = ~n5162 & ~n5164 ;
  assign n5166 = ~\g3808_reg/NET0131  & ~n5132 ;
  assign n5167 = \g3808_reg/NET0131  & n5132 ;
  assign n5168 = ~n5166 & ~n5167 ;
  assign n5169 = ~n5011 & ~n5168 ;
  assign n5170 = \g35_pad  & ~\g3817_reg/NET0131  ;
  assign n5171 = ~n5010 & n5170 ;
  assign n5172 = ~n5169 & ~n5171 ;
  assign n5173 = ~\g5037_reg/NET0131  & ~\g5041_reg/NET0131  ;
  assign n5174 = n4141 & n5173 ;
  assign n5175 = \g5037_reg/NET0131  & \g5041_reg/NET0131  ;
  assign n5176 = n4147 & n5175 ;
  assign n5177 = ~n5174 & ~n5176 ;
  assign n5178 = ~\g35_pad  & \g5041_reg/NET0131  ;
  assign n5179 = \g35_pad  & ~\g5046_reg/NET0131  ;
  assign n5180 = ~n5178 & ~n5179 ;
  assign n5181 = ~n5177 & n5180 ;
  assign n5182 = \g35_pad  & \g5046_reg/NET0131  ;
  assign n5183 = ~n4154 & n5182 ;
  assign n5184 = ~n5178 & ~n5183 ;
  assign n5185 = n5177 & n5184 ;
  assign n5186 = ~n5181 & ~n5185 ;
  assign n5187 = \g35_pad  & ~\g5069_reg/NET0131  ;
  assign n5188 = \g5073_reg/NET0131  & ~n5187 ;
  assign n5189 = \g3147_reg/NET0131  & ~n4788 ;
  assign n5190 = ~n4944 & n5189 ;
  assign n5191 = \g3147_reg/NET0131  & \g35_pad  ;
  assign n5192 = ~n4944 & n5191 ;
  assign n5193 = ~n4818 & ~n5192 ;
  assign n5194 = ~n5190 & ~n5193 ;
  assign n5195 = ~\g35_pad  & \g969_reg/NET0131  ;
  assign n5196 = \g969_reg/NET0131  & ~n2816 ;
  assign n5197 = ~n2815 & n5196 ;
  assign n5198 = ~n5195 & ~n5197 ;
  assign n5199 = ~n2816 & n3909 ;
  assign n5200 = \g1046_reg/NET0131  & ~n2816 ;
  assign n5201 = ~n2815 & n5200 ;
  assign n5202 = ~n5199 & ~n5201 ;
  assign n5203 = \g1008_reg/NET0131  & \g35_pad  ;
  assign n5204 = n5202 & n5203 ;
  assign n5205 = n5198 & ~n5204 ;
  assign n5206 = \g4646_reg/NET0131  & \g5357_reg/NET0131  ;
  assign n5207 = ~n868 & n5206 ;
  assign n5208 = \g35_pad  & \g5297_reg/NET0131  ;
  assign n5209 = ~n5207 & n5208 ;
  assign n5210 = \g5357_reg/NET0131  & ~n5208 ;
  assign n5211 = n3063 & n5210 ;
  assign n5212 = ~n5209 & ~n5211 ;
  assign n5213 = \g3352_reg/NET0131  & n2758 ;
  assign n5214 = \g3288_reg/NET0131  & \g35_pad  ;
  assign n5215 = ~n5213 & n5214 ;
  assign n5216 = \g3352_reg/NET0131  & ~n5214 ;
  assign n5217 = n2758 & n5216 ;
  assign n5218 = ~n5215 & ~n5217 ;
  assign n5219 = \g3703_reg/NET0131  & \g4681_reg/NET0131  ;
  assign n5220 = ~n2646 & n5219 ;
  assign n5221 = \g35_pad  & \g3639_reg/NET0131  ;
  assign n5222 = ~n5220 & n5221 ;
  assign n5223 = \g3703_reg/NET0131  & ~n5221 ;
  assign n5224 = n2898 & n5223 ;
  assign n5225 = ~n5222 & ~n5224 ;
  assign n5226 = ~n951 & n5008 ;
  assign n5227 = \g35_pad  & \g3990_reg/NET0131  ;
  assign n5228 = ~n5226 & n5227 ;
  assign n5229 = \g4054_reg/NET0131  & ~n5227 ;
  assign n5230 = n967 & n5229 ;
  assign n5231 = ~n5228 & ~n5230 ;
  assign n5232 = ~\g3338_reg/NET0131  & ~\g35_pad  ;
  assign n5233 = \g3347_reg/NET0131  & \g35_pad  ;
  assign n5234 = ~n5232 & ~n5233 ;
  assign n5235 = ~n4257 & n5234 ;
  assign n5236 = ~\g35_pad  & \g812_reg/NET0131  ;
  assign n5237 = ~n2586 & ~n5236 ;
  assign n5238 = ~\g817_reg/NET0131  & ~n5236 ;
  assign n5239 = ~n2579 & n5238 ;
  assign n5240 = \g817_reg/NET0131  & ~n5236 ;
  assign n5241 = n2579 & n5240 ;
  assign n5242 = ~n5239 & ~n5241 ;
  assign n5243 = ~n5237 & n5242 ;
  assign n5244 = ~\g2864_reg/NET0131  & ~\g35_pad  ;
  assign n5245 = ~\g2898_reg/NET0131  & \g35_pad  ;
  assign n5246 = n1028 & n5245 ;
  assign n5247 = ~n5244 & ~n5246 ;
  assign n5248 = ~\g35_pad  & ~\g4172_reg/NET0131  ;
  assign n5249 = ~\g4176_reg/NET0131  & n4680 ;
  assign n5250 = ~n5248 & ~n5249 ;
  assign n5251 = \g5029_reg/NET0131  & ~\g5033_reg/NET0131  ;
  assign n5252 = n4145 & n5251 ;
  assign n5253 = ~\g5029_reg/NET0131  & ~\g5033_reg/NET0131  ;
  assign n5254 = n4139 & n5253 ;
  assign n5255 = ~n5252 & ~n5254 ;
  assign n5256 = \g35_pad  & ~n5255 ;
  assign n5257 = \g5033_reg/NET0131  & n4719 ;
  assign n5258 = ~\g5029_reg/NET0131  & n4139 ;
  assign n5259 = \g5029_reg/NET0131  & n4145 ;
  assign n5260 = ~n5258 & ~n5259 ;
  assign n5261 = \g35_pad  & n5260 ;
  assign n5262 = n5257 & n5261 ;
  assign n5263 = ~n5256 & ~n5262 ;
  assign n5264 = ~\g35_pad  & \g5029_reg/NET0131  ;
  assign n5265 = n5263 & ~n5264 ;
  assign n5266 = \g3347_reg/NET0131  & ~\g35_pad  ;
  assign n5267 = \g35_pad  & ~n5207 ;
  assign n5268 = ~\g4646_reg/NET0131  & ~\g5357_reg/NET0131  ;
  assign n5269 = ~\g5357_reg/NET0131  & n862 ;
  assign n5270 = n867 & n5269 ;
  assign n5271 = ~n5268 & ~n5270 ;
  assign n5272 = n5267 & n5271 ;
  assign n5273 = ~n5266 & ~n5272 ;
  assign n5274 = \g691_reg/NET0131  & n973 ;
  assign n5275 = ~\g411_reg/NET0131  & \g417_reg/NET0131  ;
  assign n5276 = ~\g424_reg/NET0131  & ~\g691_reg/NET0131  ;
  assign n5277 = n5275 & n5276 ;
  assign n5278 = ~n5274 & ~n5277 ;
  assign n5279 = \g681_reg/NET0131  & n2455 ;
  assign n5280 = ~n5278 & n5279 ;
  assign n5281 = \g35_pad  & n5280 ;
  assign n5282 = n2455 & ~n5278 ;
  assign n5283 = \g35_pad  & \g650_reg/NET0131  ;
  assign n5284 = ~n5282 & n5283 ;
  assign n5285 = ~n5281 & ~n5284 ;
  assign n5286 = ~\g35_pad  & \g699_reg/NET0131  ;
  assign n5287 = n5285 & ~n5286 ;
  assign n5288 = \g35_pad  & ~n5282 ;
  assign n5289 = ~\g3352_reg/NET0131  & ~\g4674_reg/NET0131  ;
  assign n5290 = ~\g3352_reg/NET0131  & n2597 ;
  assign n5291 = n867 & n5290 ;
  assign n5292 = ~n5289 & ~n5291 ;
  assign n5293 = ~n2618 & n4769 ;
  assign n5294 = \g35_pad  & ~n5293 ;
  assign n5295 = n5292 & n5294 ;
  assign n5296 = ~n5266 & ~n5295 ;
  assign n5297 = ~\g35_pad  & ~\g990_reg/NET0131  ;
  assign n5298 = ~\g990_reg/NET0131  & n2821 ;
  assign n5299 = ~n5297 & ~n5298 ;
  assign n5300 = ~n2821 & n2823 ;
  assign n5301 = n2818 & n5300 ;
  assign n5302 = ~\g990_reg/NET0131  & ~n2818 ;
  assign n5303 = ~n5301 & ~n5302 ;
  assign n5304 = n5299 & n5303 ;
  assign n5305 = \g35_pad  & ~n5220 ;
  assign n5306 = ~\g3703_reg/NET0131  & ~\g4681_reg/NET0131  ;
  assign n5307 = ~\g3703_reg/NET0131  & n2625 ;
  assign n5308 = n867 & n5307 ;
  assign n5309 = ~n5306 & ~n5308 ;
  assign n5310 = n5305 & n5309 ;
  assign n5311 = ~n5266 & ~n5310 ;
  assign n5312 = \g35_pad  & ~n5226 ;
  assign n5313 = ~\g4054_reg/NET0131  & ~\g4688_reg/NET0131  ;
  assign n5314 = ~\g4054_reg/NET0131  & n950 ;
  assign n5315 = n867 & n5314 ;
  assign n5316 = ~n5313 & ~n5315 ;
  assign n5317 = n5312 & n5316 ;
  assign n5318 = ~n5266 & ~n5317 ;
  assign n5319 = \g311_reg/NET0131  & ~\g324_reg/NET0131  ;
  assign n5320 = \g35_pad  & n5319 ;
  assign n5321 = \g324_reg/NET0131  & ~\g35_pad  ;
  assign n5322 = \g305_reg/NET0131  & \g324_reg/NET0131  ;
  assign n5323 = ~n5321 & ~n5322 ;
  assign n5324 = ~n5320 & n5323 ;
  assign n5325 = \g14096_pad  & ~\g896_reg/NET0131  ;
  assign n5326 = n4057 & n5325 ;
  assign n5327 = \g35_pad  & n5326 ;
  assign n5328 = \g262_reg/NET0131  & \g35_pad  ;
  assign n5329 = ~n4061 & n5328 ;
  assign n5330 = ~n5327 & ~n5329 ;
  assign n5331 = \g232_reg/NET0131  & ~\g35_pad  ;
  assign n5332 = n5330 & ~n5331 ;
  assign n5333 = \g1008_reg/NET0131  & ~\g35_pad  ;
  assign n5334 = ~\g1002_reg/NET0131  & n2816 ;
  assign n5335 = \g35_pad  & ~n5334 ;
  assign n5336 = ~n4630 & n5335 ;
  assign n5337 = ~n5333 & ~n5336 ;
  assign n5338 = ~\g446_reg/NET0131  & n2455 ;
  assign n5339 = ~n5278 & n5338 ;
  assign n5340 = \g35_pad  & \g645_reg/NET0131  ;
  assign n5341 = \g35_pad  & n2455 ;
  assign n5342 = ~n5278 & n5341 ;
  assign n5343 = ~n5340 & ~n5342 ;
  assign n5344 = ~n5339 & ~n5343 ;
  assign n5345 = ~\g35_pad  & \g546_reg/NET0131  ;
  assign n5346 = ~\g542_reg/NET0131  & \g691_reg/NET0131  ;
  assign n5347 = n4008 & ~n5346 ;
  assign n5348 = ~n5345 & ~n5347 ;
  assign n5349 = ~\g13895_pad  & ~\g16718_pad  ;
  assign n5350 = ~n4254 & ~n5349 ;
  assign n5351 = ~\g13039_pad  & ~\g16603_pad  ;
  assign n5352 = ~\g16624_pad  & \g35_pad  ;
  assign n5353 = n5351 & n5352 ;
  assign n5354 = ~n5350 & n5353 ;
  assign n5355 = \g4633_reg/NET0131  & n2520 ;
  assign n5356 = n2523 & n5355 ;
  assign n5357 = \g35_pad  & ~n5356 ;
  assign n5358 = n1069 & n1077 ;
  assign n5359 = \g35_pad  & ~n1072 ;
  assign n5360 = ~n5358 & n5359 ;
  assign n5361 = ~n5357 & ~n5360 ;
  assign n5362 = \g35_pad  & \g4653_reg/NET0131  ;
  assign n5363 = ~\g4688_reg/NET0131  & n5362 ;
  assign n5364 = \g4688_reg/NET0131  & ~n5362 ;
  assign n5365 = ~n5363 & ~n5364 ;
  assign n5366 = \g4621_reg/NET0131  & \g4639_reg/NET0131  ;
  assign n5367 = \g4628_reg/NET0131  & n5366 ;
  assign n5368 = \g35_pad  & ~\g4643_reg/NET0131  ;
  assign n5369 = \g4633_reg/NET0131  & n5368 ;
  assign n5370 = ~n5367 & n5369 ;
  assign n5371 = ~\g4633_reg/NET0131  & ~\g4643_reg/NET0131  ;
  assign n5372 = n5366 & n5371 ;
  assign n5373 = \g35_pad  & ~n5372 ;
  assign n5374 = \g4628_reg/NET0131  & ~n5373 ;
  assign n5375 = ~n5370 & ~n5374 ;
  assign n5376 = ~\g2878_reg/NET0131  & ~\g35_pad  ;
  assign n5377 = ~\g2886_reg/NET0131  & ~\g2946_reg/NET0131  ;
  assign n5378 = \g35_pad  & n5377 ;
  assign n5379 = ~n5376 & ~n5378 ;
  assign n5380 = \g4180_reg/NET0131  & \g8786_pad  ;
  assign n5381 = \g35_pad  & n5380 ;
  assign n5382 = ~\g8787_pad  & ~\g8788_pad  ;
  assign n5383 = ~\g8789_pad  & n5382 ;
  assign n5384 = ~\g11447_pad  & ~\g8783_pad  ;
  assign n5385 = ~\g8784_pad  & ~\g8785_pad  ;
  assign n5386 = n5384 & n5385 ;
  assign n5387 = n5383 & n5386 ;
  assign n5388 = ~\g4180_reg/NET0131  & ~\g8786_pad  ;
  assign n5389 = \g35_pad  & n5388 ;
  assign n5390 = ~n5387 & n5389 ;
  assign n5391 = ~n5381 & ~n5390 ;
  assign n5392 = ~\g2946_reg/NET0131  & ~\g35_pad  ;
  assign n5393 = n5391 & ~n5392 ;
  assign n5394 = ~\g35_pad  & \g4145_reg/NET0131  ;
  assign n5395 = ~\g4076_reg/NET0131  & n871 ;
  assign n5396 = n874 & n5395 ;
  assign n5397 = \g4145_reg/NET0131  & n870 ;
  assign n5398 = n5396 & n5397 ;
  assign n5399 = ~n5394 & ~n5398 ;
  assign n5400 = n870 & n5396 ;
  assign n5401 = \g35_pad  & \g4112_reg/NET0131  ;
  assign n5402 = ~n5400 & n5401 ;
  assign n5403 = n5399 & ~n5402 ;
  assign n5404 = ~\g35_pad  & ~\g4369_reg/NET0131  ;
  assign n5405 = ~\g4462_reg/NET0131  & \g4473_reg/NET0131  ;
  assign n5406 = \g35_pad  & ~\g4459_reg/NET0131  ;
  assign n5407 = ~n5405 & n5406 ;
  assign n5408 = ~n5404 & ~n5407 ;
  assign n5409 = ~\g35_pad  & \g518_reg/NET0131  ;
  assign n5410 = \g528_reg/NET0131  & n5099 ;
  assign n5411 = ~n3991 & n5410 ;
  assign n5412 = n3992 & n5099 ;
  assign n5413 = n3991 & n5412 ;
  assign n5414 = ~n5411 & ~n5413 ;
  assign n5415 = ~n5409 & n5414 ;
  assign n5416 = \g699_reg/NET0131  & ~n2579 ;
  assign n5417 = \g35_pad  & n5416 ;
  assign n5418 = ~n5342 & ~n5417 ;
  assign n5419 = ~\g35_pad  & \g681_reg/NET0131  ;
  assign n5420 = n5418 & ~n5419 ;
  assign n5421 = \g723_reg/NET0131  & \g822_reg/NET0131  ;
  assign n5422 = \g817_reg/NET0131  & ~\g847_reg/NET0131  ;
  assign n5423 = n5421 & n5422 ;
  assign n5424 = n2579 & n5423 ;
  assign n5425 = \g35_pad  & n5424 ;
  assign n5426 = \g837_reg/NET0131  & n4108 ;
  assign n5427 = n2579 & n5426 ;
  assign n5428 = n2930 & ~n5427 ;
  assign n5429 = ~n5425 & ~n5428 ;
  assign n5430 = ~\g35_pad  & \g847_reg/NET0131  ;
  assign n5431 = n5429 & ~n5430 ;
  assign n5432 = \g35_pad  & ~n2579 ;
  assign n5433 = \g854_reg/NET0131  & ~n5432 ;
  assign n5434 = \g35_pad  & \g847_reg/NET0131  ;
  assign n5435 = ~n2579 & n5434 ;
  assign n5436 = ~n5433 & ~n5435 ;
  assign n5437 = \g35_pad  & ~n2455 ;
  assign n5438 = \g35_pad  & \g5097_reg/NET0131  ;
  assign n5439 = ~n4967 & n5438 ;
  assign n5440 = \g5092_reg/NET0131  & ~n3500 ;
  assign n5441 = ~n5438 & n5440 ;
  assign n5442 = ~n5439 & ~n5441 ;
  assign n5443 = \g1205_reg/NET0131  & ~\g35_pad  ;
  assign n5444 = \g1221_reg/NET0131  & \g35_pad  ;
  assign n5445 = ~n4012 & n5444 ;
  assign n5446 = ~\g1221_reg/NET0131  & \g35_pad  ;
  assign n5447 = n4012 & n5446 ;
  assign n5448 = ~n5445 & ~n5447 ;
  assign n5449 = ~n5443 & n5448 ;
  assign n5450 = \g182_reg/NET0131  & \g35_pad  ;
  assign n5451 = ~n2455 & n5450 ;
  assign n5452 = n2455 & n4062 ;
  assign n5453 = ~n5451 & ~n5452 ;
  assign n5454 = ~\g35_pad  & \g405_reg/NET0131  ;
  assign n5455 = n5453 & ~n5454 ;
  assign n5456 = ~\g837_reg/NET0131  & \g847_reg/NET0131  ;
  assign n5457 = n2579 & n5456 ;
  assign n5458 = \g35_pad  & ~n5457 ;
  assign n5459 = \g703_reg/NET0131  & ~n5458 ;
  assign n5460 = \g827_reg/NET0131  & \g832_reg/NET0131  ;
  assign n5461 = ~n4108 & ~n5460 ;
  assign n5462 = n2579 & ~n5461 ;
  assign n5463 = \g35_pad  & \g837_reg/NET0131  ;
  assign n5464 = ~n5462 & n5463 ;
  assign n5465 = ~n5459 & ~n5464 ;
  assign n5466 = \g4064_reg/NET0131  & ~\g4098_reg/NET0131  ;
  assign n5467 = n873 & n5466 ;
  assign n5468 = n5395 & n5467 ;
  assign n5469 = ~\g4057_reg/NET0131  & \g4145_reg/NET0131  ;
  assign n5470 = n5468 & n5469 ;
  assign n5471 = \g35_pad  & n5470 ;
  assign n5472 = ~\g4057_reg/NET0131  & n5468 ;
  assign n5473 = \g35_pad  & \g4116_reg/NET0131  ;
  assign n5474 = ~n5472 & n5473 ;
  assign n5475 = ~n5471 & ~n5474 ;
  assign n5476 = ~\g35_pad  & \g4112_reg/NET0131  ;
  assign n5477 = n5475 & ~n5476 ;
  assign n5478 = \g4057_reg/NET0131  & ~\g4064_reg/NET0131  ;
  assign n5479 = \g4145_reg/NET0131  & n5478 ;
  assign n5480 = n5396 & n5479 ;
  assign n5481 = \g35_pad  & n5480 ;
  assign n5482 = n5396 & n5478 ;
  assign n5483 = \g35_pad  & \g4119_reg/NET0131  ;
  assign n5484 = ~n5482 & n5483 ;
  assign n5485 = ~n5481 & ~n5484 ;
  assign n5486 = ~\g35_pad  & \g4116_reg/NET0131  ;
  assign n5487 = n5485 & ~n5486 ;
  assign n5488 = \g4057_reg/NET0131  & \g4145_reg/NET0131  ;
  assign n5489 = n5468 & n5488 ;
  assign n5490 = \g35_pad  & n5489 ;
  assign n5491 = \g4057_reg/NET0131  & n5468 ;
  assign n5492 = \g35_pad  & \g4122_reg/NET0131  ;
  assign n5493 = ~n5491 & n5492 ;
  assign n5494 = ~n5490 & ~n5493 ;
  assign n5495 = ~\g35_pad  & \g4119_reg/NET0131  ;
  assign n5496 = n5494 & ~n5495 ;
  assign n5497 = \g35_pad  & \g4269_reg/NET0131  ;
  assign n5498 = ~n5043 & n5497 ;
  assign n5499 = \g35_pad  & ~\g4258_reg/NET0131  ;
  assign n5500 = \g4264_reg/NET0131  & ~n5497 ;
  assign n5501 = ~n5499 & n5500 ;
  assign n5502 = ~n5498 & ~n5501 ;
  assign n5503 = \g35_pad  & \g433_reg/NET0131  ;
  assign n5504 = ~n2579 & n5503 ;
  assign n5505 = n2579 & n4330 ;
  assign n5506 = ~n5504 & ~n5505 ;
  assign n5507 = ~\g35_pad  & \g437_reg/NET0131  ;
  assign n5508 = n5506 & ~n5507 ;
  assign n5509 = \g14217_pad  & ~\g896_reg/NET0131  ;
  assign n5510 = n4057 & n5509 ;
  assign n5511 = \g35_pad  & n5510 ;
  assign n5512 = \g232_reg/NET0131  & \g35_pad  ;
  assign n5513 = ~n4061 & n5512 ;
  assign n5514 = ~n5511 & ~n5513 ;
  assign n5515 = \g255_reg/NET0131  & ~\g35_pad  ;
  assign n5516 = n5514 & ~n5515 ;
  assign n5517 = \g35_pad  & \g460_reg/NET0131  ;
  assign n5518 = ~n2455 & n5517 ;
  assign n5519 = n2455 & n4046 ;
  assign n5520 = ~n5518 & ~n5519 ;
  assign n5521 = \g168_reg/NET0131  & ~\g35_pad  ;
  assign n5522 = n5520 & ~n5521 ;
  assign n5523 = \g1548_reg/NET0131  & ~\g35_pad  ;
  assign n5524 = \g1564_reg/NET0131  & \g35_pad  ;
  assign n5525 = ~n1461 & n5524 ;
  assign n5526 = ~\g1564_reg/NET0131  & \g35_pad  ;
  assign n5527 = n1461 & n5526 ;
  assign n5528 = ~n5525 & ~n5527 ;
  assign n5529 = ~n5523 & n5528 ;
  assign n5530 = \g35_pad  & \g475_reg/NET0131  ;
  assign n5531 = ~n2579 & n5530 ;
  assign n5532 = n2579 & n4046 ;
  assign n5533 = ~n5531 & ~n5532 ;
  assign n5534 = ~\g35_pad  & \g424_reg/NET0131  ;
  assign n5535 = n5533 & ~n5534 ;
  assign n5536 = \g14201_pad  & ~\g896_reg/NET0131  ;
  assign n5537 = n4057 & n5536 ;
  assign n5538 = \g35_pad  & n5537 ;
  assign n5539 = \g255_reg/NET0131  & \g35_pad  ;
  assign n5540 = ~n4061 & n5539 ;
  assign n5541 = ~n5538 & ~n5540 ;
  assign n5542 = \g225_reg/NET0131  & ~\g35_pad  ;
  assign n5543 = n5541 & ~n5542 ;
  assign n5544 = ~\g3050_reg/NET0131  & ~\g5022_reg/NET0131  ;
  assign n5545 = \g5016_reg/NET0131  & n5544 ;
  assign n5546 = \g35_pad  & n5545 ;
  assign n5547 = ~\g5016_reg/NET0131  & ~n5544 ;
  assign n5548 = \g35_pad  & n5547 ;
  assign n5549 = n4719 & n5548 ;
  assign n5550 = ~n5546 & ~n5549 ;
  assign n5551 = ~\g35_pad  & \g5022_reg/NET0131  ;
  assign n5552 = n5550 & ~n5551 ;
  assign n5553 = \g3100_reg/NET0131  & ~\g35_pad  ;
  assign n5554 = ~\g3100_reg/NET0131  & \g5101_reg/NET0131  ;
  assign n5555 = ~\g3050_reg/NET0131  & ~n5554 ;
  assign n5556 = ~\g3096_reg/NET0131  & \g35_pad  ;
  assign n5557 = ~n5555 & n5556 ;
  assign n5558 = ~n5553 & ~n5557 ;
  assign n5559 = ~\g2932_reg/NET0131  & ~\g2999_reg/NET0131  ;
  assign n5560 = \g35_pad  & ~n5559 ;
  assign n5561 = \g1211_reg/NET0131  & \g1221_reg/NET0131  ;
  assign n5562 = n4012 & n5561 ;
  assign n5563 = ~n2818 & n5562 ;
  assign n5564 = ~\g17291_pad  & ~\g17316_pad  ;
  assign n5565 = ~\g17400_pad  & \g35_pad  ;
  assign n5566 = n5564 & n5565 ;
  assign n5567 = ~n5563 & n5566 ;
  assign n5568 = ~\g35_pad  & ~\g4072_reg/NET0131  ;
  assign n5569 = \g35_pad  & \g417_reg/NET0131  ;
  assign n5570 = ~n2579 & n5569 ;
  assign n5571 = n2579 & n4062 ;
  assign n5572 = ~n5570 & ~n5571 ;
  assign n5573 = \g35_pad  & ~\g4311_reg/NET0131  ;
  assign n5574 = ~n2525 & n5573 ;
  assign n5575 = n2524 & n5574 ;
  assign n5576 = \g35_pad  & \g4311_reg/NET0131  ;
  assign n5577 = ~n2524 & n5576 ;
  assign n5578 = ~n5575 & ~n5577 ;
  assign n5579 = ~n4141 & ~n4147 ;
  assign n5580 = \g5037_reg/NET0131  & ~n4233 ;
  assign n5581 = n4230 & n5580 ;
  assign n5582 = n5579 & n5581 ;
  assign n5583 = ~\g35_pad  & \g5033_reg/NET0131  ;
  assign n5584 = \g35_pad  & ~\g5037_reg/NET0131  ;
  assign n5585 = ~n5579 & n5584 ;
  assign n5586 = ~n5583 & ~n5585 ;
  assign n5587 = ~n5582 & n5586 ;
  assign n5588 = ~n2816 & n3906 ;
  assign n5589 = ~n2815 & n5588 ;
  assign n5590 = \g35_pad  & ~n5589 ;
  assign n5591 = \g1041_reg/NET0131  & ~n5590 ;
  assign n5592 = \g1008_reg/NET0131  & ~\g1041_reg/NET0131  ;
  assign n5593 = ~n2816 & ~n5592 ;
  assign n5594 = ~n2815 & n5593 ;
  assign n5595 = \g1046_reg/NET0131  & \g35_pad  ;
  assign n5596 = ~n5594 & n5595 ;
  assign n5597 = ~n5591 & ~n5596 ;
  assign n5598 = ~\g703_reg/NET0131  & \g854_reg/NET0131  ;
  assign n5599 = \g35_pad  & ~n5598 ;
  assign n5600 = n2579 & n5599 ;
  assign n5601 = \g35_pad  & ~\g392_reg/NET0131  ;
  assign n5602 = ~n2579 & n5601 ;
  assign n5603 = ~n5600 & ~n5602 ;
  assign n5604 = ~\g35_pad  & ~\g401_reg/NET0131  ;
  assign n5605 = n5603 & ~n5604 ;
  assign n5606 = \g1036_reg/NET0131  & ~\g35_pad  ;
  assign n5607 = \g35_pad  & ~n5594 ;
  assign n5608 = ~\g1041_reg/NET0131  & ~n4589 ;
  assign n5609 = n5607 & ~n5608 ;
  assign n5610 = ~n5606 & ~n5609 ;
  assign n5611 = ~\g35_pad  & \g4358_reg/NET0131  ;
  assign n5612 = ~\g4593_reg/NET0131  & ~\g4601_reg/NET0131  ;
  assign n5613 = ~\g4608_reg/NET0131  & ~\g4616_reg/NET0131  ;
  assign n5614 = n5612 & n5613 ;
  assign n5615 = \g4340_reg/NET0131  & ~\g4584_reg/NET0131  ;
  assign n5616 = n4660 & n5615 ;
  assign n5617 = n5614 & n5616 ;
  assign n5618 = n4659 & n5355 ;
  assign n5619 = n5617 & n5618 ;
  assign n5620 = ~n5611 & ~n5619 ;
  assign n5621 = ~\g35_pad  & \g376_reg/NET0131  ;
  assign n5622 = \g35_pad  & \g385_reg/NET0131  ;
  assign n5623 = ~n982 & n5622 ;
  assign n5624 = \g35_pad  & ~\g385_reg/NET0131  ;
  assign n5625 = n982 & n5624 ;
  assign n5626 = ~n5623 & ~n5625 ;
  assign n5627 = ~n5621 & n5626 ;
  assign n5628 = ~\g35_pad  & \g5069_reg/NET0131  ;
  assign n5629 = ~n4230 & ~n5628 ;
  assign n5630 = ~\g35_pad  & \g4284_reg/NET0131  ;
  assign n5631 = \g35_pad  & ~\g4291_reg/NET0131  ;
  assign n5632 = ~n5630 & ~n5631 ;
  assign n5633 = ~\g2902_reg/NET0131  & ~\g35_pad  ;
  assign n5634 = ~\g2917_reg/NET0131  & \g35_pad  ;
  assign n5635 = n818 & n5634 ;
  assign n5636 = n816 & n5635 ;
  assign n5637 = ~n5633 & ~n5636 ;
  assign n5638 = ~\g29214_pad  & ~\g35_pad  ;
  assign n5639 = ~\g2848_reg/NET0131  & n777 ;
  assign n5640 = n1015 & n5639 ;
  assign n5641 = ~n5638 & ~n5640 ;
  assign n5642 = ~\g35_pad  & \g4643_reg/NET0131  ;
  assign n5643 = ~\g4340_reg/NET0131  & ~n2521 ;
  assign n5644 = n4276 & ~n5643 ;
  assign n5645 = ~n5642 & ~n5644 ;
  assign n5646 = \g35_pad  & ~n3067 ;
  assign n5647 = \g35_pad  & ~n2763 ;
  assign n5648 = \g35_pad  & ~n2902 ;
  assign n5649 = \g35_pad  & ~n2776 ;
  assign n5650 = \g385_reg/NET0131  & \g513_reg/NET0131  ;
  assign n5651 = n3989 & n5650 ;
  assign n5652 = \g499_reg/NET0131  & ~n5651 ;
  assign n5653 = \g518_reg/NET0131  & ~n3993 ;
  assign n5654 = n3990 & ~n5653 ;
  assign n5655 = ~n5652 & ~n5654 ;
  assign n5656 = \g35_pad  & ~n5655 ;
  assign n5657 = ~\g35_pad  & \g5112_reg/NET0131  ;
  assign n5658 = \g3096_reg/NET0131  & ~\g5112_reg/NET0131  ;
  assign n5659 = ~\g5022_reg/NET0131  & ~n5658 ;
  assign n5660 = \g35_pad  & ~\g5101_reg/NET0131  ;
  assign n5661 = ~n5659 & n5660 ;
  assign n5662 = ~n5657 & ~n5661 ;
  assign n5663 = \g35_pad  & \g5152_reg/NET0131  ;
  assign n5664 = ~n4944 & n5663 ;
  assign n5665 = \g35_pad  & ~n4944 ;
  assign n5666 = ~\g5148_reg/NET0131  & ~n4751 ;
  assign n5667 = \g5148_reg/NET0131  & n4751 ;
  assign n5668 = ~n5666 & ~n5667 ;
  assign n5669 = ~n5665 & n5668 ;
  assign n5670 = ~n5664 & ~n5669 ;
  assign n5671 = ~\g278_reg/NET0131  & ~n2376 ;
  assign n5672 = \g35_pad  & ~n2384 ;
  assign n5673 = ~n5671 & n5672 ;
  assign n5674 = \g1300_reg/NET0131  & \g35_pad  ;
  assign n5675 = \g1484_reg/NET0131  & ~\g35_pad  ;
  assign n5676 = \g1442_reg/NET0131  & ~\g1495_reg/NET0131  ;
  assign n5677 = \g1484_reg/NET0131  & n5676 ;
  assign n5678 = n1246 & n5677 ;
  assign n5679 = ~n5675 & ~n5678 ;
  assign n5680 = n5674 & n5679 ;
  assign n5681 = ~n5674 & ~n5679 ;
  assign n5682 = ~n5680 & ~n5681 ;
  assign n5683 = \g1448_reg/NET0131  & \g35_pad  ;
  assign n5684 = \g1454_reg/NET0131  & ~\g35_pad  ;
  assign n5685 = \g1454_reg/NET0131  & n5676 ;
  assign n5686 = n1217 & n5685 ;
  assign n5687 = ~n5684 & ~n5686 ;
  assign n5688 = n5683 & n5687 ;
  assign n5689 = ~n5683 & ~n5687 ;
  assign n5690 = ~n5688 & ~n5689 ;
  assign n5691 = \g1472_reg/NET0131  & \g35_pad  ;
  assign n5692 = \g1467_reg/NET0131  & ~\g35_pad  ;
  assign n5693 = \g1467_reg/NET0131  & n5676 ;
  assign n5694 = n1232 & n5693 ;
  assign n5695 = ~n5692 & ~n5694 ;
  assign n5696 = n5691 & n5695 ;
  assign n5697 = ~n5691 & ~n5695 ;
  assign n5698 = ~n5696 & ~n5697 ;
  assign n5699 = \g1478_reg/NET0131  & \g35_pad  ;
  assign n5700 = \g1437_reg/NET0131  & ~\g35_pad  ;
  assign n5701 = \g1437_reg/NET0131  & n5676 ;
  assign n5702 = n1200 & n5701 ;
  assign n5703 = ~n5700 & ~n5702 ;
  assign n5704 = n5699 & n5703 ;
  assign n5705 = ~n5699 & ~n5703 ;
  assign n5706 = ~n5704 & ~n5705 ;
  assign n5707 = ~n4139 & ~n4145 ;
  assign n5708 = \g35_pad  & \g5029_reg/NET0131  ;
  assign n5709 = n5707 & n5708 ;
  assign n5710 = n4719 & n5709 ;
  assign n5711 = ~\g35_pad  & \g5016_reg/NET0131  ;
  assign n5712 = \g35_pad  & ~\g5029_reg/NET0131  ;
  assign n5713 = ~n5707 & n5712 ;
  assign n5714 = ~n5711 & ~n5713 ;
  assign n5715 = ~n5710 & n5714 ;
  assign n5716 = ~\g4646_reg/NET0131  & ~\g4674_reg/NET0131  ;
  assign n5717 = \g35_pad  & ~\g4681_reg/NET0131  ;
  assign n5718 = n5716 & n5717 ;
  assign n5719 = ~n2838 & n5718 ;
  assign n5720 = ~\g35_pad  & \g4621_reg/NET0131  ;
  assign n5721 = ~n5367 & n5368 ;
  assign n5722 = ~\g4628_reg/NET0131  & ~n5366 ;
  assign n5723 = n5721 & ~n5722 ;
  assign n5724 = ~n5720 & ~n5723 ;
  assign n5725 = \g35_pad  & \g5128_reg/NET0131  ;
  assign n5726 = ~n4944 & n5725 ;
  assign n5727 = \g35_pad  & ~\g5128_reg/NET0131  ;
  assign n5728 = n4944 & n5727 ;
  assign n5729 = ~n5726 & ~n5728 ;
  assign n5730 = ~\g35_pad  & \g5124_reg/NET0131  ;
  assign n5731 = n5729 & ~n5730 ;
  assign n5732 = \g3119_reg/NET0131  & \g35_pad  ;
  assign n5733 = ~n4944 & n5732 ;
  assign n5734 = ~\g3119_reg/NET0131  & \g35_pad  ;
  assign n5735 = n4944 & n5734 ;
  assign n5736 = ~n5733 & ~n5735 ;
  assign n5737 = \g3115_reg/NET0131  & ~\g35_pad  ;
  assign n5738 = n5736 & ~n5737 ;
  assign n5739 = \g35_pad  & ~n3990 ;
  assign n5740 = \g3470_reg/NET0131  & \g35_pad  ;
  assign n5741 = ~n4944 & n5740 ;
  assign n5742 = ~\g3470_reg/NET0131  & \g35_pad  ;
  assign n5743 = n4944 & n5742 ;
  assign n5744 = ~n5741 & ~n5743 ;
  assign n5745 = \g3466_reg/NET0131  & ~\g35_pad  ;
  assign n5746 = n5744 & ~n5745 ;
  assign n5747 = n989 & n2982 ;
  assign n5748 = \g35_pad  & n5747 ;
  assign n5749 = \g35_pad  & \g370_reg/NET0131  ;
  assign n5750 = ~n2983 & n5749 ;
  assign n5751 = ~n5748 & ~n5750 ;
  assign n5752 = \g358_reg/NET0131  & ~\g35_pad  ;
  assign n5753 = n5751 & ~n5752 ;
  assign n5754 = \g35_pad  & \g3821_reg/NET0131  ;
  assign n5755 = ~n4944 & n5754 ;
  assign n5756 = \g35_pad  & ~\g3821_reg/NET0131  ;
  assign n5757 = n4944 & n5756 ;
  assign n5758 = ~n5755 & ~n5757 ;
  assign n5759 = ~\g35_pad  & \g3817_reg/NET0131  ;
  assign n5760 = n5758 & ~n5759 ;
  assign n5761 = \g209_reg/NET0131  & ~n1583 ;
  assign n5762 = ~\g191_reg/NET0131  & \g8358_pad  ;
  assign n5763 = n1583 & n5762 ;
  assign n5764 = ~n5761 & ~n5763 ;
  assign n5765 = \g35_pad  & ~n5764 ;
  assign n5766 = \g191_reg/NET0131  & ~\g35_pad  ;
  assign n5767 = \g191_reg/NET0131  & ~\g8358_pad  ;
  assign n5768 = n1583 & n5767 ;
  assign n5769 = ~n5766 & ~n5768 ;
  assign n5770 = ~n5765 & n5769 ;
  assign n5771 = ~\g35_pad  & \g4180_reg/NET0131  ;
  assign n5772 = \g35_pad  & ~n2029 ;
  assign n5773 = ~n5771 & ~n5772 ;
  assign n5774 = \g35_pad  & ~\g4281_reg/NET0131  ;
  assign n5775 = ~\g35_pad  & \g4245_reg/NET0131  ;
  assign n5776 = ~n5774 & ~n5775 ;
  assign n5777 = \g1183_reg/NET0131  & \g996_reg/NET0131  ;
  assign n5778 = n4189 & n5777 ;
  assign n5779 = \g35_pad  & n5778 ;
  assign n5780 = \g1183_reg/NET0131  & n4189 ;
  assign n5781 = \g35_pad  & \g962_reg/NET0131  ;
  assign n5782 = ~n5780 & n5781 ;
  assign n5783 = ~n5779 & ~n5782 ;
  assign n5784 = \g1178_reg/NET0131  & ~\g35_pad  ;
  assign n5785 = n5783 & ~n5784 ;
  assign n5786 = ~\g35_pad  & ~\g499_reg/NET0131  ;
  assign n5787 = ~\g499_reg/NET0131  & ~n3993 ;
  assign n5788 = n3990 & n5787 ;
  assign n5789 = ~n5786 & ~n5788 ;
  assign n5790 = \g35_pad  & ~\g504_reg/NET0131  ;
  assign n5791 = ~n3990 & n5790 ;
  assign n5792 = n5789 & ~n5791 ;
  assign n5793 = \g35_pad  & ~\g4308_reg/NET0131  ;
  assign n5794 = ~\g35_pad  & \g504_reg/NET0131  ;
  assign n5795 = \g504_reg/NET0131  & ~n3993 ;
  assign n5796 = n3990 & n5795 ;
  assign n5797 = ~n5794 & ~n5796 ;
  assign n5798 = \g35_pad  & \g513_reg/NET0131  ;
  assign n5799 = ~n3990 & n5798 ;
  assign n5800 = n5797 & ~n5799 ;
  assign n5801 = ~\g2748_reg/NET0131  & ~\g35_pad  ;
  assign n5802 = \g3143_reg/NET0131  & \g35_pad  ;
  assign n5803 = ~n4944 & n5802 ;
  assign n5804 = ~\g3139_reg/NET0131  & ~n4810 ;
  assign n5805 = \g3139_reg/NET0131  & n4810 ;
  assign n5806 = ~n5804 & ~n5805 ;
  assign n5807 = ~n5665 & n5806 ;
  assign n5808 = ~n5803 & ~n5807 ;
  assign n5809 = \g3494_reg/NET0131  & \g35_pad  ;
  assign n5810 = ~n4944 & n5809 ;
  assign n5811 = ~\g3490_reg/NET0131  & ~n4994 ;
  assign n5812 = \g3490_reg/NET0131  & n4994 ;
  assign n5813 = ~n5811 & ~n5812 ;
  assign n5814 = ~n5665 & n5813 ;
  assign n5815 = ~n5810 & ~n5814 ;
  assign n5816 = \g35_pad  & \g3845_reg/NET0131  ;
  assign n5817 = ~n4944 & n5816 ;
  assign n5818 = ~\g3841_reg/NET0131  & ~n5025 ;
  assign n5819 = \g3841_reg/NET0131  & n5025 ;
  assign n5820 = ~n5818 & ~n5819 ;
  assign n5821 = ~n5665 & n5820 ;
  assign n5822 = ~n5817 & ~n5821 ;
  assign n5823 = \g4076_reg/NET0131  & \g4087_reg/NET0131  ;
  assign n5824 = ~\g4093_reg/NET0131  & \g4098_reg/NET0131  ;
  assign n5825 = n5823 & n5824 ;
  assign n5826 = n870 & n871 ;
  assign n5827 = n5825 & n5826 ;
  assign n5828 = \g35_pad  & ~n5827 ;
  assign n5829 = ~\g35_pad  & \g4639_reg/NET0131  ;
  assign n5830 = n2520 & n5368 ;
  assign n5831 = ~n5829 & ~n5830 ;
  assign n5832 = ~\g4621_reg/NET0131  & \g4639_reg/NET0131  ;
  assign n5833 = n5368 & n5832 ;
  assign n5834 = n5831 & ~n5833 ;
  assign n5835 = ~\g2965_reg/NET0131  & ~\g35_pad  ;
  assign n5836 = \g1306_reg/NET0131  & ~\g2975_reg/NET0131  ;
  assign n5837 = n5781 & n5836 ;
  assign n5838 = ~n5835 & ~n5837 ;
  assign n5839 = \g35_pad  & \g518_reg/NET0131  ;
  assign n5840 = ~n3990 & n5839 ;
  assign n5841 = ~\g35_pad  & \g513_reg/NET0131  ;
  assign n5842 = \g513_reg/NET0131  & ~n3993 ;
  assign n5843 = n3990 & n5842 ;
  assign n5844 = ~n5841 & ~n5843 ;
  assign n5845 = ~n5840 & n5844 ;
  assign n5846 = \g13272_pad  & ~\g1442_reg/NET0131  ;
  assign n5847 = n1134 & n5846 ;
  assign n5848 = \g35_pad  & n5847 ;
  assign n5849 = \g13272_pad  & \g1495_reg/NET0131  ;
  assign n5850 = n1134 & n5849 ;
  assign n5851 = \g1489_reg/NET0131  & \g35_pad  ;
  assign n5852 = ~n5850 & n5851 ;
  assign n5853 = ~n5848 & ~n5852 ;
  assign n5854 = \g35_pad  & \g4473_reg/NET0131  ;
  assign n5855 = ~\g35_pad  & \g4459_reg/NET0131  ;
  assign n5856 = ~n5854 & ~n5855 ;
  assign n5857 = ~\g35_pad  & ~\g4492_reg/NET0131  ;
  assign n5858 = ~\g2988_reg/NET0131  & \g35_pad  ;
  assign n5859 = ~n1060 & n5858 ;
  assign n5860 = ~n5857 & ~n5859 ;
  assign n5861 = \g35_pad  & ~\g4467_reg/NET0131  ;
  assign n5862 = \g4462_reg/NET0131  & \g4643_reg/NET0131  ;
  assign n5863 = n5861 & n5862 ;
  assign n5864 = \g4473_reg/NET0131  & ~n5863 ;
  assign n5865 = \g35_pad  & \g5092_reg/NET0131  ;
  assign n5866 = ~\g5084_reg/NET0131  & ~n5865 ;
  assign n5867 = \g35_pad  & n4967 ;
  assign n5868 = ~n5866 & ~n5867 ;
  assign n5869 = \g1205_reg/NET0131  & \g35_pad  ;
  assign n5870 = ~\g1087_reg/NET0131  & ~n5869 ;
  assign n5871 = \g35_pad  & n4012 ;
  assign n5872 = ~n5870 & ~n5871 ;
  assign n5873 = ~\g35_pad  & \g370_reg/NET0131  ;
  assign n5874 = ~\g358_reg/NET0131  & ~\g376_reg/NET0131  ;
  assign n5875 = \g35_pad  & ~n982 ;
  assign n5876 = ~n5874 & n5875 ;
  assign n5877 = ~n5873 & ~n5876 ;
  assign n5878 = \g35_pad  & \g4264_reg/NET0131  ;
  assign n5879 = ~\g4258_reg/NET0131  & ~n5878 ;
  assign n5880 = \g35_pad  & n5043 ;
  assign n5881 = ~n5879 & ~n5880 ;
  assign n5882 = \g35_pad  & ~\g890_reg/NET0131  ;
  assign n5883 = ~\g862_reg/NET0131  & ~n5882 ;
  assign n5884 = ~\g890_reg/NET0131  & n3018 ;
  assign n5885 = ~n5883 & ~n5884 ;
  assign n5886 = \g1548_reg/NET0131  & \g35_pad  ;
  assign n5887 = ~\g1430_reg/NET0131  & ~n5886 ;
  assign n5888 = \g35_pad  & n1461 ;
  assign n5889 = ~n5887 & ~n5888 ;
  assign n5890 = \g35_pad  & ~n1028 ;
  assign n5891 = ~\g35_pad  & \g4633_reg/NET0131  ;
  assign n5892 = \g4633_reg/NET0131  & ~\g4643_reg/NET0131  ;
  assign n5893 = n2520 & n5892 ;
  assign n5894 = ~n5891 & ~n5893 ;
  assign n5895 = \g3179_reg/NET0131  & \g35_pad  ;
  assign n5896 = \g3167_reg/NET0131  & \g3171_reg/NET0131  ;
  assign n5897 = n5895 & ~n5896 ;
  assign n5898 = ~\g3167_reg/NET0131  & \g35_pad  ;
  assign n5899 = \g3171_reg/NET0131  & ~n5895 ;
  assign n5900 = ~n5898 & n5899 ;
  assign n5901 = ~n5897 & ~n5900 ;
  assign n5902 = \g18098_pad  & \g35_pad  ;
  assign n5903 = \g305_reg/NET0131  & ~\g35_pad  ;
  assign n5904 = ~n5902 & ~n5903 ;
  assign n5905 = ~\g2886_reg/NET0131  & ~\g35_pad  ;
  assign n5906 = ~\g2980_reg/NET0131  & ~\g34_reg/NET0131  ;
  assign n5907 = \g35_pad  & n5906 ;
  assign n5908 = ~n5905 & ~n5907 ;
  assign n5909 = \g3161_reg/NET0131  & \g35_pad  ;
  assign n5910 = ~\g3155_reg/NET0131  & ~n5909 ;
  assign n5911 = \g35_pad  & n4884 ;
  assign n5912 = ~n5910 & ~n5911 ;
  assign n5913 = \g35_pad  & ~n4233 ;
  assign n5914 = ~\g35_pad  & \g5057_reg/NET0131  ;
  assign n5915 = ~n5913 & ~n5914 ;
  assign n5916 = \g35_pad  & \g9251_pad  ;
  assign n5917 = ~\g4308_reg/NET0131  & ~n5916 ;
  assign n5918 = \g4308_reg/NET0131  & n5916 ;
  assign n5919 = ~n5917 & ~n5918 ;
  assign n5920 = \g3171_reg/NET0131  & \g35_pad  ;
  assign n5921 = ~\g3167_reg/NET0131  & ~n5920 ;
  assign n5922 = \g35_pad  & n5896 ;
  assign n5923 = ~n5921 & ~n5922 ;
  assign n5924 = \g35_pad  & ~\g862_reg/NET0131  ;
  assign n5925 = ~\g896_reg/NET0131  & n5924 ;
  assign n5926 = ~\g35_pad  & ~\g890_reg/NET0131  ;
  assign n5927 = ~n3022 & ~n5926 ;
  assign n5928 = ~n5925 & n5927 ;
  assign n5929 = \g35_pad  & \g9019_pad  ;
  assign n5930 = ~\g4291_reg/NET0131  & ~n5929 ;
  assign n5931 = \g4291_reg/NET0131  & n5929 ;
  assign n5932 = ~n5930 & ~n5931 ;
  assign n5933 = \g35_pad  & ~n2982 ;
  assign n5934 = \g385_reg/NET0131  & ~n5933 ;
  assign n5935 = \g35_pad  & \g8839_pad  ;
  assign n5936 = ~\g4281_reg/NET0131  & ~n5935 ;
  assign n5937 = \g4281_reg/NET0131  & n5935 ;
  assign n5938 = ~n5936 & ~n5937 ;
  assign n5939 = \g1532_reg/NET0131  & ~\g7946_pad  ;
  assign n5940 = \g1521_reg/NET0131  & \g7946_pad  ;
  assign n5941 = ~n5939 & ~n5940 ;
  assign n5942 = \g35_pad  & ~n5941 ;
  assign n5943 = \g1306_reg/NET0131  & ~\g35_pad  ;
  assign n5944 = ~n5942 & ~n5943 ;
  assign n5945 = \g1178_reg/NET0131  & ~\g7916_pad  ;
  assign n5946 = \g7916_pad  & \g996_reg/NET0131  ;
  assign n5947 = ~n5945 & ~n5946 ;
  assign n5948 = \g35_pad  & ~n5947 ;
  assign n5949 = \g1183_reg/NET0131  & ~\g35_pad  ;
  assign n5950 = ~n5948 & ~n5949 ;
  assign n5951 = \g1189_reg/NET0131  & ~\g7916_pad  ;
  assign n5952 = \g1178_reg/NET0131  & \g7916_pad  ;
  assign n5953 = ~n5951 & ~n5952 ;
  assign n5954 = \g35_pad  & ~n5953 ;
  assign n5955 = ~\g35_pad  & \g962_reg/NET0131  ;
  assign n5956 = ~n5954 & ~n5955 ;
  assign n5957 = ~\g2724_reg/NET0131  & ~\g35_pad  ;
  assign n5958 = \g2741_reg/NET0131  & ~\g35_pad  ;
  assign n5959 = \g35_pad  & ~n1246 ;
  assign n5960 = \g3155_reg/NET0131  & ~\g3167_reg/NET0131  ;
  assign n5961 = \g35_pad  & ~n5960 ;
  assign n5962 = \g3161_reg/NET0131  & ~n5961 ;
  assign n5963 = ~\g35_pad  & \g4239_reg/NET0131  ;
  assign n5964 = ~\g10122_pad  & \g35_pad  ;
  assign n5965 = ~\g4297_reg/NET0131  & n5964 ;
  assign n5966 = ~n5963 & ~n5965 ;
  assign n5967 = ~\g35_pad  & \g4462_reg/NET0131  ;
  assign n5968 = ~\g4473_reg/NET0131  & n5861 ;
  assign n5969 = ~n5967 & ~n5968 ;
  assign n5970 = ~\g35_pad  & ~\g534_reg/NET0131  ;
  assign n5971 = \g29212_pad  & \g35_pad  ;
  assign n5972 = ~\g550_reg/NET0131  & n5971 ;
  assign n5973 = ~n5970 & ~n5972 ;
  assign n5974 = ~\g2980_reg/NET0131  & ~\g35_pad  ;
  assign n5975 = ~\g2984_reg/NET0131  & \g34_reg/NET0131  ;
  assign n5976 = \g35_pad  & n5975 ;
  assign n5977 = ~n5974 & ~n5976 ;
  assign n5978 = ~\g35_pad  & ~\g538_reg/NET0131  ;
  assign n5979 = \g35_pad  & ~\g546_reg/NET0131  ;
  assign n5980 = \g691_reg/NET0131  & n5979 ;
  assign n5981 = ~n5978 & ~n5980 ;
  assign n5982 = ~\g218_reg/NET0131  & \g35_pad  ;
  assign n5983 = \g209_reg/NET0131  & ~\g35_pad  ;
  assign n5984 = ~n5982 & ~n5983 ;
  assign n5985 = \g4146_reg/NET0131  & \g4157_reg/NET0131  ;
  assign n5986 = \g35_pad  & ~n5985 ;
  assign n5987 = ~\g35_pad  & \g4122_reg/NET0131  ;
  assign n5988 = ~n5986 & ~n5987 ;
  assign n5989 = ~\g209_reg/NET0131  & ~\g538_reg/NET0131  ;
  assign n5990 = \g35_pad  & ~n5989 ;
  assign n5991 = ~\g4153_reg/NET0131  & ~\g4172_reg/NET0131  ;
  assign n5992 = \g35_pad  & ~n5991 ;
  assign n5993 = \g4467_reg/NET0131  & \g4473_reg/NET0131  ;
  assign n5994 = \g35_pad  & ~\g4462_reg/NET0131  ;
  assign n5995 = ~n5993 & n5994 ;
  assign n5996 = ~\g3155_reg/NET0131  & n5898 ;
  assign n5997 = ~\g2715_reg/NET0131  & ~\g35_pad  ;
  assign n5998 = ~\g4639_reg/NET0131  & n5368 ;
  assign n5999 = ~\g358_reg/NET0131  & \g35_pad  ;
  assign n6000 = ~\g8719_pad  & n5999 ;
  assign n6001 = ~n5861 & ~n5994 ;
  assign n6002 = \g3050_reg/NET0131  & ~\g35_pad  ;
  assign n6003 = ~n4253 & ~n6002 ;
  assign n6004 = ~\g35_pad  & \g4483_reg/NET0131  ;
  assign n6005 = ~n1056 & ~n6004 ;
  assign n6006 = ~\g35_pad  & \g4486_reg/NET0131  ;
  assign n6007 = ~n1053 & ~n6006 ;
  assign n6008 = ~\g35_pad  & \g4489_reg/NET0131  ;
  assign n6009 = ~n1050 & ~n6008 ;
  assign n6010 = \g35_pad  & ~\g4239_reg/NET0131  ;
  assign n6011 = ~\g35_pad  & \g4273_reg/NET0131  ;
  assign n6012 = ~n6010 & ~n6011 ;
  assign n6013 = \g2735_reg/NET0131  & ~\g35_pad  ;
  assign n6014 = ~\g35_pad  & \g4382_reg/NET0131  ;
  assign n6015 = \g2719_reg/NET0131  & ~\g35_pad  ;
  assign n6016 = ~\g35_pad  & \g4392_reg/NET0131  ;
  assign n6017 = ~\g35_pad  & \g4153_reg/NET0131  ;
  assign n6018 = \g2975_reg/NET0131  & ~\g35_pad  ;
  assign n6019 = ~\g35_pad  & \g4104_reg/NET0131  ;
  assign n6020 = ~\g35_pad  & \g4087_reg/NET0131  ;
  assign n6021 = ~\g35_pad  & \g4057_reg/NET0131  ;
  assign n6022 = ~\g35_pad  & \g4076_reg/NET0131  ;
  assign n6023 = ~\g35_pad  & \g4064_reg/NET0131  ;
  assign n6024 = ~\g35_pad  & \g753_reg/NET0131  ;
  assign n6025 = ~\g2759_reg/NET0131  & ~\g35_pad  ;
  assign n6026 = ~\g35_pad  & ~\g4108_reg/NET0131  ;
  assign n6027 = ~\g2756_reg/NET0131  & ~\g35_pad  ;
  assign n6028 = ~\g2917_reg/NET0131  & ~\g35_pad  ;
  assign n6029 = \g18099_pad  & \g35_pad  ;
  assign n6030 = ~\g2882_reg/NET0131  & ~\g35_pad  ;
  assign n6031 = ~\g35_pad  & ~\g4141_reg/NET0131  ;
  assign n6032 = ~\g35_pad  & ~\g4082_reg/NET0131  ;
  assign n6033 = \g29216_pad  & \g35_pad  ;
  assign n6034 = ~\g2955_reg/NET0131  & ~\g35_pad  ;
  assign n6035 = ~\g35_pad  & ~\g4098_reg/NET0131  ;
  assign n6036 = ~\g35_pad  & ~\g4093_reg/NET0131  ;
  assign n6037 = ~\g2873_reg/NET0131  & ~\g35_pad  ;
  assign n6038 = ~\g2729_reg/NET0131  & ~\g35_pad  ;
  assign n6039 = ~\g2421_reg/NET0131  & n1837 ;
  assign n6040 = \g2495_reg/NET0131  & ~n1523 ;
  assign n6041 = \g17423_pad  & \g2495_reg/NET0131  ;
  assign n6042 = ~n1526 & n6041 ;
  assign n6043 = ~n6040 & ~n6042 ;
  assign n6044 = \g35_pad  & n6043 ;
  assign n6045 = ~n6039 & n6044 ;
  assign n6046 = ~\g2287_reg/NET0131  & n1762 ;
  assign n6047 = \g2361_reg/NET0131  & ~n1499 ;
  assign n6048 = \g17404_pad  & \g2361_reg/NET0131  ;
  assign n6049 = ~n1502 & n6048 ;
  assign n6050 = ~n6047 & ~n6049 ;
  assign n6051 = \g35_pad  & n6050 ;
  assign n6052 = ~n6046 & n6051 ;
  assign n6053 = ~\g2555_reg/NET0131  & n1907 ;
  assign n6054 = \g35_pad  & n1947 ;
  assign n6055 = ~n6053 & n6054 ;
  assign n6056 = ~\g1862_reg/NET0131  & n2123 ;
  assign n6057 = \g1936_reg/NET0131  & ~n1628 ;
  assign n6058 = \g17400_pad  & \g1936_reg/NET0131  ;
  assign n6059 = ~n1631 & n6058 ;
  assign n6060 = ~n6057 & ~n6059 ;
  assign n6061 = \g35_pad  & n6060 ;
  assign n6062 = ~n6056 & n6061 ;
  assign n6063 = ~\g1996_reg/NET0131  & n2251 ;
  assign n6064 = \g2070_reg/NET0131  & ~n1652 ;
  assign n6065 = \g1087_reg/NET0131  & \g2070_reg/NET0131  ;
  assign n6066 = ~n1655 & n6065 ;
  assign n6067 = ~n6064 & ~n6066 ;
  assign n6068 = \g35_pad  & n6067 ;
  assign n6069 = ~n6063 & n6068 ;
  assign n6070 = \g35_pad  & ~n2261 ;
  assign n6071 = \g17291_pad  & \g35_pad  ;
  assign n6072 = ~n2264 & n6071 ;
  assign n6073 = ~n6070 & ~n6072 ;
  assign n6074 = \g1682_reg/NET0131  & ~n2280 ;
  assign n6075 = ~\g1135_reg/NET0131  & ~\g1246_reg/NET0131  ;
  assign n6076 = n1469 & n6075 ;
  assign n6077 = n818 & n6076 ;
  assign n6078 = ~n6074 & n6077 ;
  assign n6079 = n6074 & ~n6077 ;
  assign n6080 = ~n6078 & ~n6079 ;
  assign n6081 = ~n6073 & n6080 ;
  assign n6082 = \g1682_reg/NET0131  & \g35_pad  ;
  assign n6083 = n2261 & n6082 ;
  assign n6084 = ~n5106 & n6083 ;
  assign n6085 = \g1668_reg/NET0131  & ~\g35_pad  ;
  assign n6086 = ~n6084 & ~n6085 ;
  assign n6087 = ~n6081 & n6086 ;
  assign n6088 = ~\g1728_reg/NET0131  & n2053 ;
  assign n6089 = \g1802_reg/NET0131  & ~n1600 ;
  assign n6090 = \g17316_pad  & \g1802_reg/NET0131  ;
  assign n6091 = ~n1607 & n6090 ;
  assign n6092 = ~n6089 & ~n6091 ;
  assign n6093 = \g35_pad  & n6092 ;
  assign n6094 = ~n6088 & n6093 ;
  assign n6095 = \g3457_reg/NET0131  & ~n4975 ;
  assign n6096 = n2901 & ~n6095 ;
  assign n6097 = ~n2645 & n6096 ;
  assign n6098 = n2901 & n6095 ;
  assign n6099 = n2645 & n6098 ;
  assign n6100 = ~n6097 & ~n6099 ;
  assign n6101 = \g3457_reg/NET0131  & ~n2898 ;
  assign n6102 = ~n963 & ~n6101 ;
  assign n6103 = n6100 & n6102 ;
  assign n6104 = \g3288_reg/NET0131  & \g3352_reg/NET0131  ;
  assign n6105 = n954 & n6104 ;
  assign n6106 = \g3106_reg/NET0131  & ~n6105 ;
  assign n6107 = n2761 & ~n6106 ;
  assign n6108 = ~n2617 & n6107 ;
  assign n6109 = n2761 & n6106 ;
  assign n6110 = n2617 & n6109 ;
  assign n6111 = ~n6108 & ~n6110 ;
  assign n6112 = \g3106_reg/NET0131  & ~n2758 ;
  assign n6113 = ~n963 & ~n6112 ;
  assign n6114 = n6111 & n6113 ;
  assign n6115 = \g1171_reg/NET0131  & ~\g35_pad  ;
  assign n6116 = \g1171_reg/NET0131  & ~\g1193_reg/NET0131  ;
  assign n6117 = ~n4201 & n6116 ;
  assign n6118 = ~n6115 & ~n6117 ;
  assign n6119 = ~\g1171_reg/NET0131  & ~n4202 ;
  assign n6120 = ~n4201 & n6119 ;
  assign n6121 = ~\g1183_reg/NET0131  & ~n4189 ;
  assign n6122 = ~n5780 & ~n6121 ;
  assign n6123 = ~n6120 & ~n6122 ;
  assign n6124 = \g35_pad  & ~n6123 ;
  assign n6125 = n6118 & ~n6124 ;
  assign n6126 = \g5297_reg/NET0131  & ~n900 ;
  assign n6127 = n895 & n6126 ;
  assign n6128 = ~\g5297_reg/NET0131  & ~n913 ;
  assign n6129 = n911 & n6128 ;
  assign n6130 = \g5357_reg/NET0131  & ~n6129 ;
  assign n6131 = ~n6127 & n6130 ;
  assign n6132 = \g5297_reg/NET0131  & ~n928 ;
  assign n6133 = ~n926 & n6132 ;
  assign n6134 = ~n922 & n6133 ;
  assign n6135 = ~\g5297_reg/NET0131  & ~n942 ;
  assign n6136 = ~n940 & n6135 ;
  assign n6137 = ~n936 & n6136 ;
  assign n6138 = ~\g5357_reg/NET0131  & ~n6137 ;
  assign n6139 = ~n6134 & n6138 ;
  assign n6140 = ~n6131 & ~n6139 ;
  assign n6141 = \g5115_reg/NET0131  & ~n4731 ;
  assign n6142 = n3066 & ~n6141 ;
  assign n6143 = ~n6140 & n6142 ;
  assign n6144 = n3066 & n6141 ;
  assign n6145 = n6140 & n6144 ;
  assign n6146 = ~n6143 & ~n6145 ;
  assign n6147 = \g5115_reg/NET0131  & ~n3063 ;
  assign n6148 = ~n963 & ~n6147 ;
  assign n6149 = n6146 & n6148 ;
  assign n6150 = ~\g2153_reg/NET0131  & n1692 ;
  assign n6151 = \g2227_reg/NET0131  & ~n1471 ;
  assign n6152 = \g17320_pad  & \g2227_reg/NET0131  ;
  assign n6153 = ~n1478 & n6152 ;
  assign n6154 = ~n6151 & ~n6153 ;
  assign n6155 = \g35_pad  & n6154 ;
  assign n6156 = ~n6150 & n6155 ;
  assign n6157 = ~\g35_pad  & \g4572_reg/NET0131  ;
  assign n6158 = ~\g35_pad  & ~n6157 ;
  assign n6159 = ~\g4776_reg/NET0131  & ~\g4793_reg/NET0131  ;
  assign n6160 = ~\g4801_reg/NET0131  & n6159 ;
  assign n6161 = ~n861 & n6160 ;
  assign n6162 = ~n2762 & ~n6161 ;
  assign n6163 = ~\g4681_reg/NET0131  & ~\g4688_reg/NET0131  ;
  assign n6164 = n5716 & n6163 ;
  assign n6165 = ~n6162 & n6164 ;
  assign n6166 = ~n862 & ~n950 ;
  assign n6167 = ~n2597 & ~n2625 ;
  assign n6168 = n6166 & n6167 ;
  assign n6169 = ~\g4776_reg/NET0131  & \g4793_reg/NET0131  ;
  assign n6170 = ~n864 & ~n6169 ;
  assign n6171 = n6164 & ~n6170 ;
  assign n6172 = ~n6168 & n6171 ;
  assign n6173 = ~n6165 & ~n6172 ;
  assign n6174 = \g3684_reg/NET0131  & \g4681_reg/NET0131  ;
  assign n6175 = ~\g4035_reg/NET0131  & \g4688_reg/NET0131  ;
  assign n6176 = ~n6174 & ~n6175 ;
  assign n6177 = \g29220_pad  & \g4646_reg/NET0131  ;
  assign n6178 = ~\g3333_reg/NET0131  & \g4674_reg/NET0131  ;
  assign n6179 = ~n6177 & ~n6178 ;
  assign n6180 = n6176 & n6179 ;
  assign n6181 = ~n6157 & n6180 ;
  assign n6182 = n6173 & n6181 ;
  assign n6183 = ~n6158 & ~n6182 ;
  assign n6184 = n6173 & n6180 ;
  assign n6185 = \g35_pad  & ~n6184 ;
  assign n6186 = \g691_reg/NET0131  & \g703_reg/NET0131  ;
  assign n6187 = ~\g714_reg/NET0131  & n6186 ;
  assign n6188 = ~n4167 & ~n6187 ;
  assign n6189 = n3989 & n5622 ;
  assign n6190 = ~n6188 & n6189 ;
  assign n6191 = \g35_pad  & \g691_reg/NET0131  ;
  assign n6192 = ~n3990 & n6191 ;
  assign n6193 = \g29212_pad  & ~\g35_pad  ;
  assign n6194 = ~n6192 & ~n6193 ;
  assign n6195 = ~n6190 & n6194 ;
  assign n6196 = ~\g29220_pad  & ~\g4646_reg/NET0131  ;
  assign n6197 = ~\g29220_pad  & n862 ;
  assign n6198 = n867 & n6197 ;
  assign n6199 = ~n6196 & ~n6198 ;
  assign n6200 = \g35_pad  & n6199 ;
  assign n6201 = ~n2594 & ~n6200 ;
  assign n6202 = n869 & ~n2594 ;
  assign n6203 = n6140 & n6202 ;
  assign n6204 = ~n6201 & ~n6203 ;
  assign n6205 = \g301_reg/NET0131  & ~\g35_pad  ;
  assign n6206 = n2393 & n2394 ;
  assign n6207 = ~n6205 & ~n6206 ;
  assign \g136_reg/P0001  = ~\g29221_pad  ;
  assign \g21727_pad  = n774 ;
  assign \g23190_pad  = ~1'b0 ;
  assign \g26875_pad  = ~n782 ;
  assign \g26876_pad  = ~n798 ;
  assign \g26877_pad  = ~n814 ;
  assign \g28041_pad  = ~n820 ;
  assign \g28042_pad  = ~n822 ;
  assign \g30327_pad  = ~\g37_reg/NET0131  ;
  assign \g30330_pad  = ~\g2834_reg/NET0131  ;
  assign \g30331_pad  = ~\g2831_reg/NET0131  ;
  assign \g31793_pad  = ~n826 ;
  assign \g31860_pad  = n827 ;
  assign \g31862_pad  = n828 ;
  assign \g31863_pad  = n829 ;
  assign \g32185_pad  = n842 ;
  assign \g33079_pad  = ~n851 ;
  assign \g33435_pad  = ~n860 ;
  assign \g33959_pad  = n869 ;
  assign \g34435_pad  = ~n878 ;
  assign \g34788_pad  = n882 ;
  assign \g34956_pad  = n886 ;
  assign \g34_reg/P0001  = ~\g34_reg/NET0131  ;
  assign \g35_syn_2  = ~\g35_pad  ;
  assign \g37/_0_  = ~n970 ;
  assign \g41/_0_  = ~n1013 ;
  assign \g60853/_3_  = n1032 ;
  assign \g60856/_3_  = n1037 ;
  assign \g60879/_3_  = n1041 ;
  assign \g60882/_0_  = ~n1048 ;
  assign \g60888/_0_  = ~n1051 ;
  assign \g60891/_0_  = ~n1054 ;
  assign \g60896/_0_  = ~n1057 ;
  assign \g60899/_0_  = ~n1081 ;
  assign \g60900/_3_  = n1092 ;
  assign \g60909/_3_  = ~n1099 ;
  assign \g60911/_0_  = ~n1103 ;
  assign \g60915/_0_  = n1106 ;
  assign \g60918/_0_  = n1133 ;
  assign \g60919/_0_  = ~n1158 ;
  assign \g60928/_0_  = ~n1164 ;
  assign \g60929/_0_  = ~n1166 ;
  assign \g60936/_0_  = ~n1172 ;
  assign \g60937/_0_  = ~n1184 ;
  assign \g60939/_0_  = ~n1198 ;
  assign \g60940/_0_  = n1216 ;
  assign \g60941/_0_  = n1230 ;
  assign \g60942/_0_  = n1245 ;
  assign \g60943/_0_  = n1259 ;
  assign \g60944/_0_  = ~n1261 ;
  assign \g60952/_0_  = ~n1272 ;
  assign \g60954/_0_  = n1280 ;
  assign \g60958/_0_  = ~n1287 ;
  assign \g60962/_3_  = n1293 ;
  assign \g60972/_0_  = n1305 ;
  assign \g60980/_0_  = ~n1316 ;
  assign \g60984/_0_  = ~n1321 ;
  assign \g60986/_0_  = ~n1322 ;
  assign \g60989/_0_  = ~n1339 ;
  assign \g60991/_3_  = n1346 ;
  assign \g61006/_0_  = ~n1351 ;
  assign \g61008/_0_  = ~n1367 ;
  assign \g61013/_0_  = n1385 ;
  assign \g61014/_0_  = n1400 ;
  assign \g61015/_0_  = n1415 ;
  assign \g61016/_0_  = n1430 ;
  assign \g61017/_0_  = ~n1431 ;
  assign \g61026/_3_  = n1438 ;
  assign \g61027/_3_  = ~n1440 ;
  assign \g61030/_0_  = ~n1446 ;
  assign \g61031/_0_  = ~n1450 ;
  assign \g61037/_0_  = ~n1460 ;
  assign \g61038/_0_  = n1468 ;
  assign \g61042/_0_  = ~n1497 ;
  assign \g61044/_0_  = ~n1521 ;
  assign \g61045/_0_  = ~n1545 ;
  assign \g61046/_0_  = ~n1569 ;
  assign \g61050/_0_  = ~n1571 ;
  assign \g61051/_0_  = ~n1575 ;
  assign \g61052/_0_  = ~n1580 ;
  assign \g61078/_0_  = ~n1581 ;
  assign \g61131/_0_  = ~n1582 ;
  assign \g61137/_3_  = ~n1590 ;
  assign \g61142/_3_  = ~n1594 ;
  assign \g61143/_3_  = ~n1598 ;
  assign \g61151/_0_  = ~n1626 ;
  assign \g61152/_0_  = ~n1650 ;
  assign \g61161/_0_  = ~n1674 ;
  assign \g61168/_3_  = n1679 ;
  assign \g61169/_3_  = ~n1688 ;
  assign \g61170/_0_  = ~n1704 ;
  assign \g61171/_3_  = ~n1715 ;
  assign \g61172/_0_  = ~n1728 ;
  assign \g61173/_0_  = ~n1741 ;
  assign \g61174/_0_  = ~n1750 ;
  assign \g61175/_0_  = ~n1758 ;
  assign \g61176/_0_  = ~n1774 ;
  assign \g61177/_3_  = ~n1785 ;
  assign \g61178/_0_  = ~n1798 ;
  assign \g61179/_0_  = ~n1811 ;
  assign \g61180/_0_  = ~n1820 ;
  assign \g61181/_0_  = ~n1828 ;
  assign \g61182/_3_  = ~n1833 ;
  assign \g61183/_0_  = ~n1849 ;
  assign \g61184/_3_  = ~n1860 ;
  assign \g61185/_0_  = ~n1873 ;
  assign \g61186/_0_  = ~n1886 ;
  assign \g61187/_0_  = ~n1895 ;
  assign \g61188/_0_  = ~n1903 ;
  assign \g61189/_0_  = ~n1919 ;
  assign \g61190/_3_  = ~n1930 ;
  assign \g61191/_0_  = ~n1943 ;
  assign \g61192/_0_  = ~n1955 ;
  assign \g61193/_0_  = ~n1964 ;
  assign \g61194/_0_  = ~n1973 ;
  assign \g61221/_0_  = ~n1974 ;
  assign \g61222/_0_  = ~n1985 ;
  assign \g61223/_3_  = ~n1991 ;
  assign \g61224/_3_  = n1994 ;
  assign \g61261/_0_  = ~n1995 ;
  assign \g61295/_3_  = n2004 ;
  assign \g61308/_0_  = ~n2011 ;
  assign \g61316/_0_  = ~n2014 ;
  assign \g61327/_0_  = n2020 ;
  assign \g61329/_0_  = ~n2047 ;
  assign \g61330/_0_  = ~n2049 ;
  assign \g61331/_0_  = ~n2065 ;
  assign \g61332/_3_  = ~n2076 ;
  assign \g61333/_0_  = ~n2089 ;
  assign \g61334/_0_  = ~n2102 ;
  assign \g61335/_0_  = ~n2111 ;
  assign \g61336/_0_  = ~n2119 ;
  assign \g61337/_0_  = ~n2135 ;
  assign \g61338/_3_  = ~n2146 ;
  assign \g61339/_0_  = ~n2159 ;
  assign \g61340/_0_  = ~n2172 ;
  assign \g61341/_0_  = ~n2181 ;
  assign \g61342/_0_  = ~n2189 ;
  assign \g61343/_0_  = ~n2205 ;
  assign \g61344/_3_  = ~n2216 ;
  assign \g61345/_0_  = ~n2229 ;
  assign \g61346/_0_  = ~n2238 ;
  assign \g61347/_0_  = ~n2247 ;
  assign \g61348/_0_  = ~n2259 ;
  assign \g61349/_0_  = ~n2279 ;
  assign \g61350/_3_  = ~n2291 ;
  assign \g61351/_0_  = ~n2304 ;
  assign \g61352/_0_  = ~n2313 ;
  assign \g61353/_0_  = ~n2322 ;
  assign \g61354/_0_  = ~n2332 ;
  assign \g61367/_0_  = ~n2339 ;
  assign \g61372/_0_  = ~n2342 ;
  assign \g61373/_0_  = ~n2370 ;
  assign \g61375/_0_  = ~n2401 ;
  assign \g61382/_0_  = ~n2402 ;
  assign \g61385/_3_  = ~n2408 ;
  assign \g61386/_0_  = ~n2420 ;
  assign \g61399/_0_  = ~n2422 ;
  assign \g61400/_0_  = ~n2433 ;
  assign \g61402/_0_  = n2435 ;
  assign \g61405/_0_  = ~n2436 ;
  assign \g61435/_3_  = n2445 ;
  assign \g61449/_0_  = n2468 ;
  assign \g61468/_0_  = ~n2480 ;
  assign \g61475/_0_  = n2487 ;
  assign \g61480/_0_  = n2493 ;
  assign \g61482/_0_  = n2503 ;
  assign \g61483/_0_  = ~n2519 ;
  assign \g61484/_0_  = ~n2540 ;
  assign \g61486/_3_  = ~n2549 ;
  assign \g61494/_0_  = ~n2552 ;
  assign \g61496/_0_  = ~n2564 ;
  assign \g61497/_0_  = ~n2573 ;
  assign \g61514/_0_  = ~n2577 ;
  assign \g61517/_0_  = ~n2593 ;
  assign \g61519/_3_  = n2622 ;
  assign \g61520/_3_  = n2650 ;
  assign \g61527/_0_  = ~n2652 ;
  assign \g61541/_0_  = ~n2663 ;
  assign \g61544/_0_  = ~n2674 ;
  assign \g61550/_0_  = ~n2676 ;
  assign \g61551/_0_  = ~n2679 ;
  assign \g61554/_0_  = ~n2689 ;
  assign \g61556/_3_  = n2699 ;
  assign \g61567/_0_  = n2712 ;
  assign \g61571/_0_  = ~n2721 ;
  assign \g61574/_0_  = n2730 ;
  assign \g61587/_0_  = ~n2735 ;
  assign \g61592/_0_  = ~n2744 ;
  assign \g61632/_0_  = n2754 ;
  assign \g61634/_0_  = ~n2774 ;
  assign \g61635/_0_  = ~n2787 ;
  assign \g61639/_0_  = ~n2804 ;
  assign \g61644/_0_  = ~n2812 ;
  assign \g61652/_3_  = ~n2835 ;
  assign \g61709/_0_  = ~n2844 ;
  assign \g61714/_0_  = ~n2853 ;
  assign \g61720/_0_  = n2861 ;
  assign \g61721/_0_  = ~n2870 ;
  assign \g61723/_0_  = ~n2878 ;
  assign \g61725/_0_  = ~n2886 ;
  assign \g61726/_0_  = ~n2894 ;
  assign \g61734/_0_  = ~n2913 ;
  assign \g61739/_0_  = ~n2939 ;
  assign \g61744/_0_  = n2947 ;
  assign \g61746/_3_  = ~n2950 ;
  assign \g61747/_3_  = ~n2957 ;
  assign \g61748/_3_  = ~n2960 ;
  assign \g61750/u3_syn_7  = ~n2961 ;
  assign \g61802/_0_  = ~n2981 ;
  assign \g61804/_0_  = ~n3024 ;
  assign \g61808/_0_  = ~n3040 ;
  assign \g61811/_0_  = ~n3059 ;
  assign \g61816/_0_  = ~n3078 ;
  assign \g61818/_0_  = ~n3092 ;
  assign \g61820/_0_  = ~n3105 ;
  assign \g61823/_0_  = ~n3110 ;
  assign \g61824/_0_  = ~n3120 ;
  assign \g61841/_0_  = ~n3126 ;
  assign \g61842/_3_  = ~n3130 ;
  assign \g61844/_3_  = ~n3148 ;
  assign \g61845/_3_  = ~n3157 ;
  assign \g61846/_3_  = ~n3170 ;
  assign \g61847/u3_syn_7  = ~n3171 ;
  assign \g61848/_0_  = n3184 ;
  assign \g61849/_3_  = ~n3193 ;
  assign \g61850/_0_  = n3206 ;
  assign \g61851/u3_syn_7  = ~n3207 ;
  assign \g61852/_0_  = n3220 ;
  assign \g61853/_3_  = ~n3232 ;
  assign \g61854/_3_  = ~n3241 ;
  assign \g61855/_0_  = n3254 ;
  assign \g61856/u3_syn_7  = ~n3255 ;
  assign \g61857/_0_  = n3263 ;
  assign \g61858/_3_  = ~n3276 ;
  assign \g61859/_3_  = ~n3285 ;
  assign \g61860/u3_syn_7  = ~n3286 ;
  assign \g61861/_0_  = n3299 ;
  assign \g61862/_3_  = ~n3315 ;
  assign \g61863/_3_  = ~n3324 ;
  assign \g61864/u3_syn_7  = ~n3325 ;
  assign \g61865/_0_  = n3338 ;
  assign \g61866/_3_  = ~n3351 ;
  assign \g61867/_3_  = ~n3360 ;
  assign \g61868/u3_syn_7  = ~n3361 ;
  assign \g61869/_0_  = n3374 ;
  assign \g61870/_0_  = n3383 ;
  assign \g61871/_3_  = ~n3396 ;
  assign \g61872/_3_  = ~n3405 ;
  assign \g61873/u3_syn_7  = ~n3406 ;
  assign \g61874/_0_  = n3419 ;
  assign \g61875/_0_  = n3427 ;
  assign \g61877/_3_  = ~n3440 ;
  assign \g61878/_3_  = ~n3449 ;
  assign \g61879/u3_syn_7  = ~n3450 ;
  assign \g61880/_0_  = n3463 ;
  assign \g61881/_0_  = n3471 ;
  assign \g61882/_0_  = n3479 ;
  assign \g61883/_0_  = n3487 ;
  assign \g61884/_0_  = n3495 ;
  assign \g61914/_0_  = ~n3499 ;
  assign \g61915/_0_  = ~n3508 ;
  assign \g61917/_0_  = ~n3535 ;
  assign \g61918/_0_  = n3542 ;
  assign \g61922/_0_  = ~n3554 ;
  assign \g61923/_0_  = ~n3563 ;
  assign \g61924/_0_  = n3574 ;
  assign \g61932/_0_  = ~n3596 ;
  assign \g61936/_0_  = n3607 ;
  assign \g61945/_0_  = ~n3612 ;
  assign \g61947/_0_  = ~n3616 ;
  assign \g61959/_0_  = ~n3625 ;
  assign \g61960/_0_  = ~n3633 ;
  assign \g61962/_0_  = n3642 ;
  assign \g61973/_3_  = ~n3651 ;
  assign \g61974/u3_syn_7  = ~n3648 ;
  assign \g61975/_3_  = ~n3673 ;
  assign \g61976/u3_syn_7  = ~n3674 ;
  assign \g61977/_3_  = n3681 ;
  assign \g61978/_3_  = ~n3702 ;
  assign \g61979/u3_syn_7  = ~n3703 ;
  assign \g61980/_3_  = ~n3710 ;
  assign \g61981/_3_  = ~n3731 ;
  assign \g61982/_3_  = ~n3738 ;
  assign \g61983/u3_syn_7  = ~n3739 ;
  assign \g61984/_3_  = n3746 ;
  assign \g61985/_3_  = ~n3767 ;
  assign \g61986/u3_syn_7  = ~n3768 ;
  assign \g61987/_3_  = n3776 ;
  assign \g61988/_3_  = ~n3798 ;
  assign \g61989/u3_syn_7  = ~n3799 ;
  assign \g61990/_3_  = n3806 ;
  assign \g61991/_3_  = ~n3827 ;
  assign \g61992/u3_syn_7  = ~n3828 ;
  assign \g61993/_3_  = n3835 ;
  assign \g61994/u3_syn_7  = ~n3836 ;
  assign \g61995/_3_  = ~n3857 ;
  assign \g61996/_3_  = ~n3864 ;
  assign \g61997/_3_  = ~n3885 ;
  assign \g62022/_0_  = ~n3893 ;
  assign \g62028/_0_  = ~n3902 ;
  assign \g62029/_0_  = ~n3905 ;
  assign \g62031/_0_  = n3930 ;
  assign \g62033/_0_  = ~n3938 ;
  assign \g62038/_0_  = ~n3946 ;
  assign \g62042/_0_  = ~n3955 ;
  assign \g62046/_0_  = ~n3963 ;
  assign \g62048/_0_  = ~n3972 ;
  assign \g62049/_0_  = ~n3980 ;
  assign \g62051/_0_  = ~n3988 ;
  assign \g62053/_0_  = ~n4004 ;
  assign \g62085/_0_  = ~n4011 ;
  assign \g62101/_0_  = ~n4020 ;
  assign \g62102/_0_  = ~n4033 ;
  assign \g62103/_0_  = ~n4040 ;
  assign \g62105/_0_  = n4045 ;
  assign \g62108/_3_  = ~n4048 ;
  assign \g62112/_0_  = ~n4056 ;
  assign \g62137/_3_  = ~n4066 ;
  assign \g62207/_0_  = n4069 ;
  assign \g62239/_0_  = ~n4090 ;
  assign \g62240/_0_  = ~n4096 ;
  assign \g62267/_0_  = ~n4103 ;
  assign \g62273/_0_  = n4114 ;
  assign \g62284/_0_  = ~n4119 ;
  assign \g62291/_0_  = ~n4123 ;
  assign \g62293/_0_  = ~n4129 ;
  assign \g62298/_0_  = ~n4138 ;
  assign \g62303/_3_  = ~n4162 ;
  assign \g62322/_3_  = ~n4172 ;
  assign \g62323/_3_  = ~n4175 ;
  assign \g62324/_3_  = ~n4180 ;
  assign \g62325/_3_  = ~n4187 ;
  assign \g62583/_0_  = ~n4205 ;
  assign \g62598/_0_  = ~n4212 ;
  assign \g62609/_0_  = ~n4226 ;
  assign \g62636/_0_  = ~n4245 ;
  assign \g62646/_0_  = n4252 ;
  assign \g62649/_0_  = n4258 ;
  assign \g62658/_0_  = ~n4267 ;
  assign \g62663/_0_  = ~n4269 ;
  assign \g62664/_0_  = ~n4271 ;
  assign \g62667/_0_  = ~n4279 ;
  assign \g62676/_0_  = ~n4286 ;
  assign \g62677/_0_  = ~n4291 ;
  assign \g62678/_3_  = ~n4299 ;
  assign \g62679/_0_  = ~n4306 ;
  assign \g62687/u3_syn_7  = ~n4307 ;
  assign \g62688/u3_syn_7  = ~n4308 ;
  assign \g62689/_0_  = n4319 ;
  assign \g62690/_3_  = ~n4326 ;
  assign \g62691/_3_  = ~n4334 ;
  assign \g62693/_0_  = n4345 ;
  assign \g62694/_3_  = ~n4354 ;
  assign \g62695/_3_  = ~n4364 ;
  assign \g62696/_3_  = ~n4375 ;
  assign \g62697/_3_  = ~n4386 ;
  assign \g62698/_3_  = ~n4393 ;
  assign \g62699/_3_  = ~n4401 ;
  assign \g62700/_3_  = ~n4409 ;
  assign \g62701/_3_  = ~n4418 ;
  assign \g62702/_3_  = ~n4427 ;
  assign \g62703/_3_  = ~n4432 ;
  assign \g62704/u3_syn_7  = ~n4428 ;
  assign \g62705/_0_  = n4443 ;
  assign \g62706/_3_  = ~n4450 ;
  assign \g62707/_3_  = ~n4455 ;
  assign \g62708/u3_syn_7  = ~n4451 ;
  assign \g62709/_0_  = n4466 ;
  assign \g62710/_3_  = ~n4473 ;
  assign \g62711/_3_  = ~n4478 ;
  assign \g62712/u3_syn_7  = ~n4474 ;
  assign \g62713/_0_  = n4489 ;
  assign \g62714/_3_  = ~n4496 ;
  assign \g62715/_0_  = ~n4501 ;
  assign \g62716/u3_syn_7  = ~n4497 ;
  assign \g62717/_0_  = n4512 ;
  assign \g62718/_3_  = ~n4519 ;
  assign \g62719/_0_  = ~n4524 ;
  assign \g62720/u3_syn_7  = ~n4520 ;
  assign \g62721/_0_  = n4535 ;
  assign \g62722/_3_  = ~n4542 ;
  assign \g62723/_0_  = ~n4547 ;
  assign \g62724/u3_syn_7  = ~n4543 ;
  assign \g62725/_0_  = n4558 ;
  assign \g62726/_3_  = ~n4565 ;
  assign \g62728/_0_  = ~n4569 ;
  assign \g62790/_0_  = n4580 ;
  assign \g62791/_0_  = n4592 ;
  assign \g62793/_0_  = n4599 ;
  assign \g62794/_0_  = n4606 ;
  assign \g62795/_0_  = n4613 ;
  assign \g62796/_0_  = n4620 ;
  assign \g62797/_0_  = n4627 ;
  assign \g62807/_0_  = ~n4638 ;
  assign \g62823/_0_  = ~n4643 ;
  assign \g62824/_0_  = n4648 ;
  assign \g62833/_0_  = ~n4656 ;
  assign \g62846/_0_  = ~n4664 ;
  assign \g62859/_0_  = n4671 ;
  assign \g62860/_0_  = n4678 ;
  assign \g62897/_0_  = n4683 ;
  assign \g62898/_0_  = ~n4690 ;
  assign \g62922/_3_  = ~n4696 ;
  assign \g62923/_0_  = n4703 ;
  assign \g62927/_0_  = ~n4708 ;
  assign \g62938/_3_  = ~n4713 ;
  assign \g62939/_3_  = ~n4725 ;
  assign \g62940/_3_  = ~n4730 ;
  assign \g62941/u3_syn_7  = ~n4734 ;
  assign \g62942/_0_  = n4748 ;
  assign \g62943/_3_  = ~n4755 ;
  assign \g62987/_3_  = ~n4761 ;
  assign \g62991/_3_  = ~n4768 ;
  assign \g63015/u3_syn_7  = ~n4773 ;
  assign \g63016/_0_  = n4784 ;
  assign \g63017/_3_  = ~n4797 ;
  assign \g63018/_3_  = ~n4807 ;
  assign \g63019/_3_  = ~n4814 ;
  assign \g63020/_3_  = ~n4822 ;
  assign \g63021/_3_  = ~n4832 ;
  assign \g63022/_3_  = ~n4839 ;
  assign \g63025/_3_  = ~n4847 ;
  assign \g63026/_3_  = ~n4854 ;
  assign \g63027/_3_  = ~n4861 ;
  assign \g63029/_3_  = ~n4869 ;
  assign \g63030/_3_  = ~n4876 ;
  assign \g63031/_3_  = ~n4883 ;
  assign \g63033/_3_  = ~n4891 ;
  assign \g63034/_3_  = ~n4898 ;
  assign \g63043/_3_  = ~n4908 ;
  assign \g63044/_3_  = ~n4915 ;
  assign \g63051/_3_  = ~n4922 ;
  assign \g63057/_3_  = ~n4929 ;
  assign \g63068/_3_  = ~n4936 ;
  assign \g63070/_3_  = ~n4943 ;
  assign \g63073/_3_  = ~n4950 ;
  assign \g63081/_3_  = ~n4956 ;
  assign \g63082/_3_  = ~n4963 ;
  assign \g63083/u3_syn_7  = ~n4964 ;
  assign \g63084/_3_  = ~n4973 ;
  assign \g63085/_0_  = n4991 ;
  assign \g63086/_3_  = ~n4998 ;
  assign \g63107/_3_  = ~n5004 ;
  assign \g63108/u3_syn_7  = ~n5006 ;
  assign \g63109/u3_syn_7  = ~n5011 ;
  assign \g63110/_0_  = n5022 ;
  assign \g63111/_3_  = ~n5029 ;
  assign \g63132/_3_  = ~n5035 ;
  assign \g63133/_3_  = ~n5042 ;
  assign \g63134/_3_  = ~n5052 ;
  assign \g63135/_3_  = n5061 ;
  assign \g63136/_3_  = ~n5067 ;
  assign \g63137/_3_  = ~n5074 ;
  assign \g63138/_3_  = ~n5082 ;
  assign \g63139/u3_syn_7  = ~n5083 ;
  assign \g63140/_3_  = ~n5089 ;
  assign \g63141/_3_  = ~n5096 ;
  assign \g63142/_3_  = n5105 ;
  assign \g63143/_3_  = ~n5112 ;
  assign \g63144/_3_  = n5122 ;
  assign \g63145/_3_  = ~n5129 ;
  assign \g63146/u3_syn_7  = ~n5131 ;
  assign \g63198/_0_  = n5139 ;
  assign \g63205/_0_  = n5146 ;
  assign \g63208/_0_  = n5151 ;
  assign \g63212/_0_  = n5158 ;
  assign \g63215/_0_  = n5165 ;
  assign \g63219/_0_  = n5172 ;
  assign \g63244/_0_  = n5186 ;
  assign \g63246/_0_  = n5188 ;
  assign \g63254/_0_  = n5194 ;
  assign \g63255/_0_  = ~n5205 ;
  assign \g63272/_0_  = ~n5212 ;
  assign \g63276/_0_  = ~n5218 ;
  assign \g63278/_0_  = ~n5225 ;
  assign \g63279/_0_  = ~n5231 ;
  assign \g63280/_0_  = n5235 ;
  assign \g63327/_0_  = n5243 ;
  assign \g63345/_0_  = n5247 ;
  assign \g63346/_3_  = n5250 ;
  assign \g63347/_3_  = ~n5265 ;
  assign \g63354/_3_  = ~n5273 ;
  assign \g63358/_3_  = ~n5287 ;
  assign \g63359/u3_syn_7  = ~n5288 ;
  assign \g63361/_3_  = ~n5296 ;
  assign \g63365/_3_  = n5304 ;
  assign \g63366/_3_  = ~n5311 ;
  assign \g63367/_3_  = ~n5318 ;
  assign \g63368/_3_  = ~n5324 ;
  assign \g63370/_3_  = ~n5332 ;
  assign \g63479/_0_  = ~n5337 ;
  assign \g63484/_0_  = n5344 ;
  assign \g63499/_1_  = n2013 ;
  assign \g63520/_0_  = ~n5348 ;
  assign \g63523/_0_  = n5354 ;
  assign \g63526/_0_  = ~n5361 ;
  assign \g63538/_0_  = ~n5365 ;
  assign \g63539/_0_  = ~n5375 ;
  assign \g63541/_0_  = n5379 ;
  assign \g63555/_0_  = n5393 ;
  assign \g63642/_0_  = ~n5403 ;
  assign \g63645/_0_  = n5408 ;
  assign \g63648/_3_  = ~n5415 ;
  assign \g63777/_3_  = ~n5420 ;
  assign \g63778/_3_  = ~n5431 ;
  assign \g63781/_0_  = ~n5436 ;
  assign \g63786/u3_syn_7  = ~n5437 ;
  assign \g63787/_3_  = ~n5442 ;
  assign \g63788/_3_  = ~n5449 ;
  assign \g63790/_3_  = ~n5455 ;
  assign \g63791/_3_  = ~n5465 ;
  assign \g63792/u3_syn_7  = ~n5432 ;
  assign \g63794/_0_  = ~n5477 ;
  assign \g63795/_0_  = ~n5487 ;
  assign \g63796/_0_  = ~n5496 ;
  assign \g63798/_3_  = ~n5502 ;
  assign \g63800/_3_  = ~n5508 ;
  assign \g63804/_3_  = ~n5516 ;
  assign \g63805/_3_  = ~n5522 ;
  assign \g63806/_3_  = ~n5529 ;
  assign \g63807/_3_  = ~n5535 ;
  assign \g63808/_3_  = ~n5543 ;
  assign \g63809/_3_  = ~n5552 ;
  assign \g63870/_0_  = ~n5558 ;
  assign \g63883/_0_  = n5560 ;
  assign \g63934/_0_  = n5567 ;
  assign \g63936/_0_  = ~n5568 ;
  assign \g63938/_0_  = ~n5572 ;
  assign \g63939/_0_  = ~n5578 ;
  assign \g63966/_0_  = ~n5587 ;
  assign \g63970/_0_  = ~n5597 ;
  assign \g63999/_0_  = n5605 ;
  assign \g64039/_0_  = ~n5610 ;
  assign \g64040/_0_  = ~n5620 ;
  assign \g64043/_0_  = ~n5627 ;
  assign \g64062/_3_  = ~n5629 ;
  assign \g64078/_0_  = ~n5632 ;
  assign \g64091/_0_  = n5637 ;
  assign \g64095/_3_  = n5641 ;
  assign \g64096/_3_  = ~n5645 ;
  assign \g64097/u3_syn_7  = ~n5646 ;
  assign \g64098/u3_syn_7  = ~n5647 ;
  assign \g64099/u3_syn_7  = ~n5648 ;
  assign \g64100/u3_syn_7  = ~n5649 ;
  assign \g64134/_0_  = n5656 ;
  assign \g64135/_0_  = ~n5662 ;
  assign \g64153/_0_  = ~n5670 ;
  assign \g64155/_0_  = n5673 ;
  assign \g64179/_0_  = ~n5682 ;
  assign \g64229/_0_  = ~n5690 ;
  assign \g64235/_0_  = ~n5698 ;
  assign \g64236/_0_  = ~n5706 ;
  assign \g64280/_0_  = ~n5715 ;
  assign \g64315/_0_  = n5719 ;
  assign \g64365/_0_  = ~n5724 ;
  assign \g64426/_3_  = ~n5731 ;
  assign \g64438/_3_  = ~n5738 ;
  assign \g64442/u3_syn_7  = ~n5739 ;
  assign \g64445/_3_  = ~n5746 ;
  assign \g64447/_3_  = ~n5753 ;
  assign \g64449/_3_  = ~n5760 ;
  assign \g64451/_3_  = ~n5770 ;
  assign \g64453/_3_  = ~n5773 ;
  assign \g64454/_3_  = ~n5776 ;
  assign \g64460/_3_  = ~n5785 ;
  assign \g64461/_3_  = n5792 ;
  assign \g64510/_0_  = n5793 ;
  assign \g64527/_0_  = ~n5800 ;
  assign \g64528/_0_  = ~n5801 ;
  assign \g64544/_0_  = ~n5808 ;
  assign \g64549/_0_  = ~n5815 ;
  assign \g64566/_0_  = ~n5822 ;
  assign \g64576/_0_  = n5828 ;
  assign \g64602/_0_  = ~n5834 ;
  assign \g64691/_0_  = n5838 ;
  assign \g64697/_0_  = ~n5845 ;
  assign \g64707/_3_  = ~n5853 ;
  assign \g64778/_3_  = ~n5856 ;
  assign \g64790/_3_  = n5860 ;
  assign \g64791/_3_  = n5864 ;
  assign \g64792/_3_  = n5868 ;
  assign \g64793/_3_  = n5872 ;
  assign \g64794/_3_  = ~n5877 ;
  assign \g64795/_3_  = n5881 ;
  assign \g64796/_3_  = n5885 ;
  assign \g64797/_3_  = n5889 ;
  assign \g64877/_0_  = ~n5890 ;
  assign \g64912/_0_  = ~n5894 ;
  assign \g64973/_0_  = ~n5901 ;
  assign \g65047/_3_  = ~n5904 ;
  assign \g65081/_3_  = n5908 ;
  assign \g65088/_3_  = n5912 ;
  assign \g65097/_3_  = ~n5915 ;
  assign \g65100/_3_  = n5919 ;
  assign \g65101/_3_  = n5923 ;
  assign \g65104/_3_  = n5928 ;
  assign \g65105/_3_  = n5932 ;
  assign \g65107/_3_  = n5934 ;
  assign \g65110/_3_  = n5938 ;
  assign \g65111/_3_  = ~n5944 ;
  assign \g65113/_3_  = ~n5950 ;
  assign \g65114/_3_  = ~n5956 ;
  assign \g65266/_0_  = ~n5957 ;
  assign \g65267/_0_  = n5958 ;
  assign \g65294/_1_  = ~n5665 ;
  assign \g65328/_1_  = ~n5959 ;
  assign \g65495/_0_  = n5962 ;
  assign \g65499/_0_  = ~n5966 ;
  assign \g65503/_0_  = ~n5969 ;
  assign \g65529/_0_  = n5973 ;
  assign \g65530/_3_  = n5977 ;
  assign \g65531/_3_  = n5981 ;
  assign \g65532/_3_  = ~n5984 ;
  assign \g65533/_3_  = ~n5988 ;
  assign \g65624/_0_  = n5990 ;
  assign \g65625/_1_  = n4944 ;
  assign \g65641/_0_  = n5992 ;
  assign \g65701/_0_  = ~n5995 ;
  assign \g65704/_0_  = n5996 ;
  assign \g65853/_0_  = ~n5997 ;
  assign \g65891/_0_  = n5998 ;
  assign \g65901/_0_  = n6000 ;
  assign \g65986/_0_  = ~n6001 ;
  assign \g66029/_0_  = ~n6003 ;
  assign \g66066/_0_  = ~n6005 ;
  assign \g66067/_0_  = ~n6007 ;
  assign \g66068/_0_  = ~n6009 ;
  assign \g66154/_3_  = ~n6012 ;
  assign \g66362/_0_  = n6013 ;
  assign \g66369/_0_  = n6014 ;
  assign \g66398/_0_  = n6015 ;
  assign \g66409/_0_  = n6016 ;
  assign \g66419/_0_  = n6017 ;
  assign \g66439/_0_  = n6018 ;
  assign \g66443/_0_  = n6019 ;
  assign \g66464/_0_  = n6020 ;
  assign \g66471/_0_  = n6021 ;
  assign \g66512/_0_  = n6022 ;
  assign \g66528/_0_  = n6023 ;
  assign \g66541/_0_  = n5499 ;
  assign \g66558/_0_  = n6024 ;
  assign \g66644/_0_  = ~n6025 ;
  assign \g66684/_0_  = ~n6026 ;
  assign \g66697/_0_  = ~n6027 ;
  assign \g66698/_0_  = n5895 ;
  assign \g66701/_0_  = ~n6028 ;
  assign \g66714/_0_  = n6029 ;
  assign \g66715/_0_  = ~n6030 ;
  assign \g66745/_0_  = ~n6031 ;
  assign \g66750/_0_  = ~n6032 ;
  assign \g66751/_0_  = n6033 ;
  assign \g66810/_0_  = ~n6034 ;
  assign \g66844/_0_  = ~n6035 ;
  assign \g66853/_0_  = ~n6036 ;
  assign \g66897/_0_  = ~n6037 ;
  assign \g66905/_0_  = ~n6038 ;
  assign \g69743/_0_  = n6045 ;
  assign \g69750/_0_  = n6052 ;
  assign \g69773/_1_  = n6055 ;
  assign \g69792/_1_  = n6062 ;
  assign \g69858/_0_  = n6069 ;
  assign \g69938/_0_  = ~n6087 ;
  assign \g69949/_0_  = n6094 ;
  assign \g70167/_0_  = ~n6103 ;
  assign \g71190/_0_  = ~n6114 ;
  assign \g71198/_0_  = ~n6125 ;
  assign \g71284/_0_  = ~n6149 ;
  assign \g72369/_1_  = n5106 ;
  assign \g72467/_0_  = n6156 ;
  assign \g72476/_0_  = n6183 ;
  assign \g72477/_1_  = n6185 ;
  assign \g72648/_0_  = ~n6195 ;
  assign \g72741/_0_  = n6204 ;
  assign \g72772/_0_  = ~n6207 ;
  assign \g8132_pad  = 1'b0 ;
endmodule
