module top (\A[0] , \A[1] , \A[2] , \A[3] , \A[4] , \A[5] , \A[6] , \A[7] , \A[8] , \A[9] , \A[10] , \A[11] , \A[12] , \A[13] , \A[14] , \A[15] , \A[16] , \A[17] , \A[18] , \A[19] , \A[20] , \A[21] , \A[22] , \A[23] , \A[24] , \A[25] , \A[26] , \A[27] , \A[28] , \A[29] , \A[30] , \A[31] , \A[32] , \A[33] , \A[34] , \A[35] , \A[36] , \A[37] , \A[38] , \A[39] , \A[40] , \A[41] , \A[42] , \A[43] , \A[44] , \A[45] , \A[46] , \A[47] , \A[48] , \A[49] , \A[50] , \A[51] , \A[52] , \A[53] , \A[54] , \A[55] , \A[56] , \A[57] , \A[58] , \A[59] , \A[60] , \A[61] , \A[62] , \A[63] , \A[64] , \A[65] , \A[66] , \A[67] , \A[68] , \A[69] , \A[70] , \A[71] , \A[72] , \A[73] , \A[74] , \A[75] , \A[76] , \A[77] , \A[78] , \A[79] , \A[80] , \A[81] , \A[82] , \A[83] , \A[84] , \A[85] , \A[86] , \A[87] , \A[88] , \A[89] , \A[90] , \A[91] , \A[92] , \A[93] , \A[94] , \A[95] , \A[96] , \A[97] , \A[98] , \A[99] , \A[100] , \A[101] , \A[102] , \A[103] , \A[104] , \A[105] , \A[106] , \A[107] , \A[108] , \A[109] , \A[110] , \A[111] , \A[112] , \A[113] , \A[114] , \A[115] , \A[116] , \A[117] , \A[118] , \A[119] , \A[120] , \A[121] , \A[122] , \A[123] , \A[124] , \A[125] , \A[126] , \A[127] , \A[128] , \A[129] , \A[130] , \A[131] , \A[132] , \A[133] , \A[134] , \A[135] , \A[136] , \A[137] , \A[138] , \A[139] , \A[140] , \A[141] , \A[142] , \A[143] , \A[144] , \A[145] , \A[146] , \A[147] , \A[148] , \A[149] , \A[150] , \A[151] , \A[152] , \A[153] , \A[154] , \A[155] , \A[156] , \A[157] , \A[158] , \A[159] , \A[160] , \A[161] , \A[162] , \A[163] , \A[164] , \A[165] , \A[166] , \A[167] , \A[168] , \A[169] , \A[170] , \A[171] , \A[172] , \A[173] , \A[174] , \A[175] , \A[176] , \A[177] , \A[178] , \A[179] , \A[180] , \A[181] , \A[182] , \A[183] , \A[184] , \A[185] , \A[186] , \A[187] , \A[188] , \A[189] , \A[190] , \A[191] , \A[192] , \A[193] , \A[194] , \A[195] , \A[196] , \A[197] , \A[198] , \A[199] , \A[200] , \A[201] , \A[202] , \A[203] , \A[204] , \A[205] , \A[206] , \A[207] , \A[208] , \A[209] , \A[210] , \A[211] , \A[212] , \A[213] , \A[214] , \A[215] , \A[216] , \A[217] , \A[218] , \A[219] , \A[220] , \A[221] , \A[222] , \A[223] , \A[224] , \A[225] , \A[226] , \A[227] , \A[228] , \A[229] , \A[230] , \A[231] , \A[232] , \A[233] , \A[234] , \A[235] , \A[236] , \A[237] , \A[238] , \A[239] , \A[240] , \A[241] , \A[242] , \A[243] , \A[244] , \A[245] , \A[246] , \A[247] , \A[248] , \A[249] , \A[250] , \A[251] , \A[252] , \A[253] , \A[254] , \A[255] , \A[256] , \A[257] , \A[258] , \A[259] , \A[260] , \A[261] , \A[262] , \A[263] , \A[264] , \A[265] , \A[266] , \A[267] , \A[268] , \A[269] , \A[270] , \A[271] , \A[272] , \A[273] , \A[274] , \A[275] , \A[276] , \A[277] , \A[278] , \A[279] , \A[280] , \A[281] , \A[282] , \A[283] , \A[284] , \A[285] , \A[286] , \A[287] , \A[288] , \A[289] , \A[290] , \A[291] , \A[292] , \A[293] , \A[294] , \A[295] , \A[296] , \A[297] , \A[298] , \A[299] , \A[300] , \A[301] , \A[302] , \A[303] , \A[304] , \A[305] , \A[306] , \A[307] , \A[308] , \A[309] , \A[310] , \A[311] , \A[312] , \A[313] , \A[314] , \A[315] , \A[316] , \A[317] , \A[318] , \A[319] , \A[320] , \A[321] , \A[322] , \A[323] , \A[324] , \A[325] , \A[326] , \A[327] , \A[328] , \A[329] , \A[330] , \A[331] , \A[332] , \A[333] , \A[334] , \A[335] , \A[336] , \A[337] , \A[338] , \A[339] , \A[340] , \A[341] , \A[342] , \A[343] , \A[344] , \A[345] , \A[346] , \A[347] , \A[348] , \A[349] , \A[350] , \A[351] , \A[352] , \A[353] , \A[354] , \A[355] , \A[356] , \A[357] , \A[358] , \A[359] , \A[360] , \A[361] , \A[362] , \A[363] , \A[364] , \A[365] , \A[366] , \A[367] , \A[368] , \A[369] , \A[370] , \A[371] , \A[372] , \A[373] , \A[374] , \A[375] , \A[376] , \A[377] , \A[378] , \A[379] , \A[380] , \A[381] , \A[382] , \A[383] , \A[384] , \A[385] , \A[386] , \A[387] , \A[388] , \A[389] , \A[390] , \A[391] , \A[392] , \A[393] , \A[394] , \A[395] , \A[396] , \A[397] , \A[398] , \A[399] , \A[400] , \A[401] , \A[402] , \A[403] , \A[404] , \A[405] , \A[406] , \A[407] , \A[408] , \A[409] , \A[410] , \A[411] , \A[412] , \A[413] , \A[414] , \A[415] , \A[416] , \A[417] , \A[418] , \A[419] , \A[420] , \A[421] , \A[422] , \A[423] , \A[424] , \A[425] , \A[426] , \A[427] , \A[428] , \A[429] , \A[430] , \A[431] , \A[432] , \A[433] , \A[434] , \A[435] , \A[436] , \A[437] , \A[438] , \A[439] , \A[440] , \A[441] , \A[442] , \A[443] , \A[444] , \A[445] , \A[446] , \A[447] , \A[448] , \A[449] , \A[450] , \A[451] , \A[452] , \A[453] , \A[454] , \A[455] , \A[456] , \A[457] , \A[458] , \A[459] , \A[460] , \A[461] , \A[462] , \A[463] , \A[464] , \A[465] , \A[466] , \A[467] , \A[468] , \A[469] , \A[470] , \A[471] , \A[472] , \A[473] , \A[474] , \A[475] , \A[476] , \A[477] , \A[478] , \A[479] , \A[480] , \A[481] , \A[482] , \A[483] , \A[484] , \A[485] , \A[486] , \A[487] , \A[488] , \A[489] , \A[490] , \A[491] , \A[492] , \A[493] , \A[494] , \A[495] , \A[496] , \A[497] , \A[498] , \A[499] , \A[500] , \A[501] , \A[502] , \A[503] , \A[504] , \A[505] , \A[506] , \A[507] , \A[508] , \A[509] , \A[510] , \A[511] , \A[512] , \A[513] , \A[514] , \A[515] , \A[516] , \A[517] , \A[518] , \A[519] , \A[520] , \A[521] , \A[522] , \A[523] , \A[524] , \A[525] , \A[526] , \A[527] , \A[528] , \A[529] , \A[530] , \A[531] , \A[532] , \A[533] , \A[534] , \A[535] , \A[536] , \A[537] , \A[538] , \A[539] , \A[540] , \A[541] , \A[542] , \A[543] , \A[544] , \A[545] , \A[546] , \A[547] , \A[548] , \A[549] , \A[550] , \A[551] , \A[552] , \A[553] , \A[554] , \A[555] , \A[556] , \A[557] , \A[558] , \A[559] , \A[560] , \A[561] , \A[562] , \A[563] , \A[564] , \A[565] , \A[566] , \A[567] , \A[568] , \A[569] , \A[570] , \A[571] , \A[572] , \A[573] , \A[574] , \A[575] , \A[576] , \A[577] , \A[578] , \A[579] , \A[580] , \A[581] , \A[582] , \A[583] , \A[584] , \A[585] , \A[586] , \A[587] , \A[588] , \A[589] , \A[590] , \A[591] , \A[592] , \A[593] , \A[594] , \A[595] , \A[596] , \A[597] , \A[598] , \A[599] , \A[600] , \A[601] , \A[602] , \A[603] , \A[604] , \A[605] , \A[606] , \A[607] , \A[608] , \A[609] , \A[610] , \A[611] , \A[612] , \A[613] , \A[614] , \A[615] , \A[616] , \A[617] , \A[618] , \A[619] , \A[620] , \A[621] , \A[622] , \A[623] , \A[624] , \A[625] , \A[626] , \A[627] , \A[628] , \A[629] , \A[630] , \A[631] , \A[632] , \A[633] , \A[634] , \A[635] , \A[636] , \A[637] , \A[638] , \A[639] , \A[640] , \A[641] , \A[642] , \A[643] , \A[644] , \A[645] , \A[646] , \A[647] , \A[648] , \A[649] , \A[650] , \A[651] , \A[652] , \A[653] , \A[654] , \A[655] , \A[656] , \A[657] , \A[658] , \A[659] , \A[660] , \A[661] , \A[662] , \A[663] , \A[664] , \A[665] , \A[666] , \A[667] , \A[668] , \A[669] , \A[670] , \A[671] , \A[672] , \A[673] , \A[674] , \A[675] , \A[676] , \A[677] , \A[678] , \A[679] , \A[680] , \A[681] , \A[682] , \A[683] , \A[684] , \A[685] , \A[686] , \A[687] , \A[688] , \A[689] , \A[690] , \A[691] , \A[692] , \A[693] , \A[694] , \A[695] , \A[696] , \A[697] , \A[698] , \A[699] , \A[700] , \A[701] , \A[702] , \A[703] , \A[704] , \A[705] , \A[706] , \A[707] , \A[708] , \A[709] , \A[710] , \A[711] , \A[712] , \A[713] , \A[714] , \A[715] , \A[716] , \A[717] , \A[718] , \A[719] , \A[720] , \A[721] , \A[722] , \A[723] , \A[724] , \A[725] , \A[726] , \A[727] , \A[728] , \A[729] , \A[730] , \A[731] , \A[732] , \A[733] , \A[734] , \A[735] , \A[736] , \A[737] , \A[738] , \A[739] , \A[740] , \A[741] , \A[742] , \A[743] , \A[744] , \A[745] , \A[746] , \A[747] , \A[748] , \A[749] , \A[750] , \A[751] , \A[752] , \A[753] , \A[754] , \A[755] , \A[756] , \A[757] , \A[758] , \A[759] , \A[760] , \A[761] , \A[762] , \A[763] , \A[764] , \A[765] , \A[766] , \A[767] , \A[768] , \A[769] , \A[770] , \A[771] , \A[772] , \A[773] , \A[774] , \A[775] , \A[776] , \A[777] , \A[778] , \A[779] , \A[780] , \A[781] , \A[782] , \A[783] , \A[784] , \A[785] , \A[786] , \A[787] , \A[788] , \A[789] , \A[790] , \A[791] , \A[792] , \A[793] , \A[794] , \A[795] , \A[796] , \A[797] , \A[798] , \A[799] , \A[800] , \A[801] , \A[802] , \A[803] , \A[804] , \A[805] , \A[806] , \A[807] , \A[808] , \A[809] , \A[810] , \A[811] , \A[812] , \A[813] , \A[814] , \A[815] , \A[816] , \A[817] , \A[818] , \A[819] , \A[820] , \A[821] , \A[822] , \A[823] , \A[824] , \A[825] , \A[826] , \A[827] , \A[828] , \A[829] , \A[830] , \A[831] , \A[832] , \A[833] , \A[834] , \A[835] , \A[836] , \A[837] , \A[838] , \A[839] , \A[840] , \A[841] , \A[842] , \A[843] , \A[844] , \A[845] , \A[846] , \A[847] , \A[848] , \A[849] , \A[850] , \A[851] , \A[852] , \A[853] , \A[854] , \A[855] , \A[856] , \A[857] , \A[858] , \A[859] , \A[860] , \A[861] , \A[862] , \A[863] , \A[864] , \A[865] , \A[866] , \A[867] , \A[868] , \A[869] , \A[870] , \A[871] , \A[872] , \A[873] , \A[874] , \A[875] , \A[876] , \A[877] , \A[878] , \A[879] , \A[880] , \A[881] , \A[882] , \A[883] , \A[884] , \A[885] , \A[886] , \A[887] , \A[888] , \A[889] , \A[890] , \A[891] , \A[892] , \A[893] , \A[894] , \A[895] , \A[896] , \A[897] , \A[898] , \A[899] , \A[900] , \A[901] , \A[902] , \A[903] , \A[904] , \A[905] , \A[906] , \A[907] , \A[908] , \A[909] , \A[910] , \A[911] , \A[912] , \A[913] , \A[914] , \A[915] , \A[916] , \A[917] , \A[918] , \A[919] , \A[920] , \A[921] , \A[922] , \A[923] , \A[924] , \A[925] , \A[926] , \A[927] , \A[928] , \A[929] , \A[930] , \A[931] , \A[932] , \A[933] , \A[934] , \A[935] , \A[936] , \A[937] , \A[938] , \A[939] , \A[940] , \A[941] , \A[942] , \A[943] , \A[944] , \A[945] , \A[946] , \A[947] , \A[948] , \A[949] , \A[950] , \A[951] , \A[952] , \A[953] , \A[954] , \A[955] , \A[956] , \A[957] , \A[958] , \A[959] , \A[960] , \A[961] , \A[962] , \A[963] , \A[964] , \A[965] , \A[966] , \A[967] , \A[968] , \A[969] , \A[970] , \A[971] , \A[972] , \A[973] , \A[974] , \A[975] , \A[976] , \A[977] , \A[978] , \A[979] , \A[980] , \A[981] , \A[982] , \A[983] , \A[984] , \A[985] , \A[986] , \A[987] , \A[988] , \A[989] , \A[990] , \A[991] , \A[992] , \A[993] , \A[994] , \A[995] , \A[996] , \A[997] , \A[998] , \A[999] , \A[1000] , maj);
	input \A[0]  ;
	input \A[1]  ;
	input \A[2]  ;
	input \A[3]  ;
	input \A[4]  ;
	input \A[5]  ;
	input \A[6]  ;
	input \A[7]  ;
	input \A[8]  ;
	input \A[9]  ;
	input \A[10]  ;
	input \A[11]  ;
	input \A[12]  ;
	input \A[13]  ;
	input \A[14]  ;
	input \A[15]  ;
	input \A[16]  ;
	input \A[17]  ;
	input \A[18]  ;
	input \A[19]  ;
	input \A[20]  ;
	input \A[21]  ;
	input \A[22]  ;
	input \A[23]  ;
	input \A[24]  ;
	input \A[25]  ;
	input \A[26]  ;
	input \A[27]  ;
	input \A[28]  ;
	input \A[29]  ;
	input \A[30]  ;
	input \A[31]  ;
	input \A[32]  ;
	input \A[33]  ;
	input \A[34]  ;
	input \A[35]  ;
	input \A[36]  ;
	input \A[37]  ;
	input \A[38]  ;
	input \A[39]  ;
	input \A[40]  ;
	input \A[41]  ;
	input \A[42]  ;
	input \A[43]  ;
	input \A[44]  ;
	input \A[45]  ;
	input \A[46]  ;
	input \A[47]  ;
	input \A[48]  ;
	input \A[49]  ;
	input \A[50]  ;
	input \A[51]  ;
	input \A[52]  ;
	input \A[53]  ;
	input \A[54]  ;
	input \A[55]  ;
	input \A[56]  ;
	input \A[57]  ;
	input \A[58]  ;
	input \A[59]  ;
	input \A[60]  ;
	input \A[61]  ;
	input \A[62]  ;
	input \A[63]  ;
	input \A[64]  ;
	input \A[65]  ;
	input \A[66]  ;
	input \A[67]  ;
	input \A[68]  ;
	input \A[69]  ;
	input \A[70]  ;
	input \A[71]  ;
	input \A[72]  ;
	input \A[73]  ;
	input \A[74]  ;
	input \A[75]  ;
	input \A[76]  ;
	input \A[77]  ;
	input \A[78]  ;
	input \A[79]  ;
	input \A[80]  ;
	input \A[81]  ;
	input \A[82]  ;
	input \A[83]  ;
	input \A[84]  ;
	input \A[85]  ;
	input \A[86]  ;
	input \A[87]  ;
	input \A[88]  ;
	input \A[89]  ;
	input \A[90]  ;
	input \A[91]  ;
	input \A[92]  ;
	input \A[93]  ;
	input \A[94]  ;
	input \A[95]  ;
	input \A[96]  ;
	input \A[97]  ;
	input \A[98]  ;
	input \A[99]  ;
	input \A[100]  ;
	input \A[101]  ;
	input \A[102]  ;
	input \A[103]  ;
	input \A[104]  ;
	input \A[105]  ;
	input \A[106]  ;
	input \A[107]  ;
	input \A[108]  ;
	input \A[109]  ;
	input \A[110]  ;
	input \A[111]  ;
	input \A[112]  ;
	input \A[113]  ;
	input \A[114]  ;
	input \A[115]  ;
	input \A[116]  ;
	input \A[117]  ;
	input \A[118]  ;
	input \A[119]  ;
	input \A[120]  ;
	input \A[121]  ;
	input \A[122]  ;
	input \A[123]  ;
	input \A[124]  ;
	input \A[125]  ;
	input \A[126]  ;
	input \A[127]  ;
	input \A[128]  ;
	input \A[129]  ;
	input \A[130]  ;
	input \A[131]  ;
	input \A[132]  ;
	input \A[133]  ;
	input \A[134]  ;
	input \A[135]  ;
	input \A[136]  ;
	input \A[137]  ;
	input \A[138]  ;
	input \A[139]  ;
	input \A[140]  ;
	input \A[141]  ;
	input \A[142]  ;
	input \A[143]  ;
	input \A[144]  ;
	input \A[145]  ;
	input \A[146]  ;
	input \A[147]  ;
	input \A[148]  ;
	input \A[149]  ;
	input \A[150]  ;
	input \A[151]  ;
	input \A[152]  ;
	input \A[153]  ;
	input \A[154]  ;
	input \A[155]  ;
	input \A[156]  ;
	input \A[157]  ;
	input \A[158]  ;
	input \A[159]  ;
	input \A[160]  ;
	input \A[161]  ;
	input \A[162]  ;
	input \A[163]  ;
	input \A[164]  ;
	input \A[165]  ;
	input \A[166]  ;
	input \A[167]  ;
	input \A[168]  ;
	input \A[169]  ;
	input \A[170]  ;
	input \A[171]  ;
	input \A[172]  ;
	input \A[173]  ;
	input \A[174]  ;
	input \A[175]  ;
	input \A[176]  ;
	input \A[177]  ;
	input \A[178]  ;
	input \A[179]  ;
	input \A[180]  ;
	input \A[181]  ;
	input \A[182]  ;
	input \A[183]  ;
	input \A[184]  ;
	input \A[185]  ;
	input \A[186]  ;
	input \A[187]  ;
	input \A[188]  ;
	input \A[189]  ;
	input \A[190]  ;
	input \A[191]  ;
	input \A[192]  ;
	input \A[193]  ;
	input \A[194]  ;
	input \A[195]  ;
	input \A[196]  ;
	input \A[197]  ;
	input \A[198]  ;
	input \A[199]  ;
	input \A[200]  ;
	input \A[201]  ;
	input \A[202]  ;
	input \A[203]  ;
	input \A[204]  ;
	input \A[205]  ;
	input \A[206]  ;
	input \A[207]  ;
	input \A[208]  ;
	input \A[209]  ;
	input \A[210]  ;
	input \A[211]  ;
	input \A[212]  ;
	input \A[213]  ;
	input \A[214]  ;
	input \A[215]  ;
	input \A[216]  ;
	input \A[217]  ;
	input \A[218]  ;
	input \A[219]  ;
	input \A[220]  ;
	input \A[221]  ;
	input \A[222]  ;
	input \A[223]  ;
	input \A[224]  ;
	input \A[225]  ;
	input \A[226]  ;
	input \A[227]  ;
	input \A[228]  ;
	input \A[229]  ;
	input \A[230]  ;
	input \A[231]  ;
	input \A[232]  ;
	input \A[233]  ;
	input \A[234]  ;
	input \A[235]  ;
	input \A[236]  ;
	input \A[237]  ;
	input \A[238]  ;
	input \A[239]  ;
	input \A[240]  ;
	input \A[241]  ;
	input \A[242]  ;
	input \A[243]  ;
	input \A[244]  ;
	input \A[245]  ;
	input \A[246]  ;
	input \A[247]  ;
	input \A[248]  ;
	input \A[249]  ;
	input \A[250]  ;
	input \A[251]  ;
	input \A[252]  ;
	input \A[253]  ;
	input \A[254]  ;
	input \A[255]  ;
	input \A[256]  ;
	input \A[257]  ;
	input \A[258]  ;
	input \A[259]  ;
	input \A[260]  ;
	input \A[261]  ;
	input \A[262]  ;
	input \A[263]  ;
	input \A[264]  ;
	input \A[265]  ;
	input \A[266]  ;
	input \A[267]  ;
	input \A[268]  ;
	input \A[269]  ;
	input \A[270]  ;
	input \A[271]  ;
	input \A[272]  ;
	input \A[273]  ;
	input \A[274]  ;
	input \A[275]  ;
	input \A[276]  ;
	input \A[277]  ;
	input \A[278]  ;
	input \A[279]  ;
	input \A[280]  ;
	input \A[281]  ;
	input \A[282]  ;
	input \A[283]  ;
	input \A[284]  ;
	input \A[285]  ;
	input \A[286]  ;
	input \A[287]  ;
	input \A[288]  ;
	input \A[289]  ;
	input \A[290]  ;
	input \A[291]  ;
	input \A[292]  ;
	input \A[293]  ;
	input \A[294]  ;
	input \A[295]  ;
	input \A[296]  ;
	input \A[297]  ;
	input \A[298]  ;
	input \A[299]  ;
	input \A[300]  ;
	input \A[301]  ;
	input \A[302]  ;
	input \A[303]  ;
	input \A[304]  ;
	input \A[305]  ;
	input \A[306]  ;
	input \A[307]  ;
	input \A[308]  ;
	input \A[309]  ;
	input \A[310]  ;
	input \A[311]  ;
	input \A[312]  ;
	input \A[313]  ;
	input \A[314]  ;
	input \A[315]  ;
	input \A[316]  ;
	input \A[317]  ;
	input \A[318]  ;
	input \A[319]  ;
	input \A[320]  ;
	input \A[321]  ;
	input \A[322]  ;
	input \A[323]  ;
	input \A[324]  ;
	input \A[325]  ;
	input \A[326]  ;
	input \A[327]  ;
	input \A[328]  ;
	input \A[329]  ;
	input \A[330]  ;
	input \A[331]  ;
	input \A[332]  ;
	input \A[333]  ;
	input \A[334]  ;
	input \A[335]  ;
	input \A[336]  ;
	input \A[337]  ;
	input \A[338]  ;
	input \A[339]  ;
	input \A[340]  ;
	input \A[341]  ;
	input \A[342]  ;
	input \A[343]  ;
	input \A[344]  ;
	input \A[345]  ;
	input \A[346]  ;
	input \A[347]  ;
	input \A[348]  ;
	input \A[349]  ;
	input \A[350]  ;
	input \A[351]  ;
	input \A[352]  ;
	input \A[353]  ;
	input \A[354]  ;
	input \A[355]  ;
	input \A[356]  ;
	input \A[357]  ;
	input \A[358]  ;
	input \A[359]  ;
	input \A[360]  ;
	input \A[361]  ;
	input \A[362]  ;
	input \A[363]  ;
	input \A[364]  ;
	input \A[365]  ;
	input \A[366]  ;
	input \A[367]  ;
	input \A[368]  ;
	input \A[369]  ;
	input \A[370]  ;
	input \A[371]  ;
	input \A[372]  ;
	input \A[373]  ;
	input \A[374]  ;
	input \A[375]  ;
	input \A[376]  ;
	input \A[377]  ;
	input \A[378]  ;
	input \A[379]  ;
	input \A[380]  ;
	input \A[381]  ;
	input \A[382]  ;
	input \A[383]  ;
	input \A[384]  ;
	input \A[385]  ;
	input \A[386]  ;
	input \A[387]  ;
	input \A[388]  ;
	input \A[389]  ;
	input \A[390]  ;
	input \A[391]  ;
	input \A[392]  ;
	input \A[393]  ;
	input \A[394]  ;
	input \A[395]  ;
	input \A[396]  ;
	input \A[397]  ;
	input \A[398]  ;
	input \A[399]  ;
	input \A[400]  ;
	input \A[401]  ;
	input \A[402]  ;
	input \A[403]  ;
	input \A[404]  ;
	input \A[405]  ;
	input \A[406]  ;
	input \A[407]  ;
	input \A[408]  ;
	input \A[409]  ;
	input \A[410]  ;
	input \A[411]  ;
	input \A[412]  ;
	input \A[413]  ;
	input \A[414]  ;
	input \A[415]  ;
	input \A[416]  ;
	input \A[417]  ;
	input \A[418]  ;
	input \A[419]  ;
	input \A[420]  ;
	input \A[421]  ;
	input \A[422]  ;
	input \A[423]  ;
	input \A[424]  ;
	input \A[425]  ;
	input \A[426]  ;
	input \A[427]  ;
	input \A[428]  ;
	input \A[429]  ;
	input \A[430]  ;
	input \A[431]  ;
	input \A[432]  ;
	input \A[433]  ;
	input \A[434]  ;
	input \A[435]  ;
	input \A[436]  ;
	input \A[437]  ;
	input \A[438]  ;
	input \A[439]  ;
	input \A[440]  ;
	input \A[441]  ;
	input \A[442]  ;
	input \A[443]  ;
	input \A[444]  ;
	input \A[445]  ;
	input \A[446]  ;
	input \A[447]  ;
	input \A[448]  ;
	input \A[449]  ;
	input \A[450]  ;
	input \A[451]  ;
	input \A[452]  ;
	input \A[453]  ;
	input \A[454]  ;
	input \A[455]  ;
	input \A[456]  ;
	input \A[457]  ;
	input \A[458]  ;
	input \A[459]  ;
	input \A[460]  ;
	input \A[461]  ;
	input \A[462]  ;
	input \A[463]  ;
	input \A[464]  ;
	input \A[465]  ;
	input \A[466]  ;
	input \A[467]  ;
	input \A[468]  ;
	input \A[469]  ;
	input \A[470]  ;
	input \A[471]  ;
	input \A[472]  ;
	input \A[473]  ;
	input \A[474]  ;
	input \A[475]  ;
	input \A[476]  ;
	input \A[477]  ;
	input \A[478]  ;
	input \A[479]  ;
	input \A[480]  ;
	input \A[481]  ;
	input \A[482]  ;
	input \A[483]  ;
	input \A[484]  ;
	input \A[485]  ;
	input \A[486]  ;
	input \A[487]  ;
	input \A[488]  ;
	input \A[489]  ;
	input \A[490]  ;
	input \A[491]  ;
	input \A[492]  ;
	input \A[493]  ;
	input \A[494]  ;
	input \A[495]  ;
	input \A[496]  ;
	input \A[497]  ;
	input \A[498]  ;
	input \A[499]  ;
	input \A[500]  ;
	input \A[501]  ;
	input \A[502]  ;
	input \A[503]  ;
	input \A[504]  ;
	input \A[505]  ;
	input \A[506]  ;
	input \A[507]  ;
	input \A[508]  ;
	input \A[509]  ;
	input \A[510]  ;
	input \A[511]  ;
	input \A[512]  ;
	input \A[513]  ;
	input \A[514]  ;
	input \A[515]  ;
	input \A[516]  ;
	input \A[517]  ;
	input \A[518]  ;
	input \A[519]  ;
	input \A[520]  ;
	input \A[521]  ;
	input \A[522]  ;
	input \A[523]  ;
	input \A[524]  ;
	input \A[525]  ;
	input \A[526]  ;
	input \A[527]  ;
	input \A[528]  ;
	input \A[529]  ;
	input \A[530]  ;
	input \A[531]  ;
	input \A[532]  ;
	input \A[533]  ;
	input \A[534]  ;
	input \A[535]  ;
	input \A[536]  ;
	input \A[537]  ;
	input \A[538]  ;
	input \A[539]  ;
	input \A[540]  ;
	input \A[541]  ;
	input \A[542]  ;
	input \A[543]  ;
	input \A[544]  ;
	input \A[545]  ;
	input \A[546]  ;
	input \A[547]  ;
	input \A[548]  ;
	input \A[549]  ;
	input \A[550]  ;
	input \A[551]  ;
	input \A[552]  ;
	input \A[553]  ;
	input \A[554]  ;
	input \A[555]  ;
	input \A[556]  ;
	input \A[557]  ;
	input \A[558]  ;
	input \A[559]  ;
	input \A[560]  ;
	input \A[561]  ;
	input \A[562]  ;
	input \A[563]  ;
	input \A[564]  ;
	input \A[565]  ;
	input \A[566]  ;
	input \A[567]  ;
	input \A[568]  ;
	input \A[569]  ;
	input \A[570]  ;
	input \A[571]  ;
	input \A[572]  ;
	input \A[573]  ;
	input \A[574]  ;
	input \A[575]  ;
	input \A[576]  ;
	input \A[577]  ;
	input \A[578]  ;
	input \A[579]  ;
	input \A[580]  ;
	input \A[581]  ;
	input \A[582]  ;
	input \A[583]  ;
	input \A[584]  ;
	input \A[585]  ;
	input \A[586]  ;
	input \A[587]  ;
	input \A[588]  ;
	input \A[589]  ;
	input \A[590]  ;
	input \A[591]  ;
	input \A[592]  ;
	input \A[593]  ;
	input \A[594]  ;
	input \A[595]  ;
	input \A[596]  ;
	input \A[597]  ;
	input \A[598]  ;
	input \A[599]  ;
	input \A[600]  ;
	input \A[601]  ;
	input \A[602]  ;
	input \A[603]  ;
	input \A[604]  ;
	input \A[605]  ;
	input \A[606]  ;
	input \A[607]  ;
	input \A[608]  ;
	input \A[609]  ;
	input \A[610]  ;
	input \A[611]  ;
	input \A[612]  ;
	input \A[613]  ;
	input \A[614]  ;
	input \A[615]  ;
	input \A[616]  ;
	input \A[617]  ;
	input \A[618]  ;
	input \A[619]  ;
	input \A[620]  ;
	input \A[621]  ;
	input \A[622]  ;
	input \A[623]  ;
	input \A[624]  ;
	input \A[625]  ;
	input \A[626]  ;
	input \A[627]  ;
	input \A[628]  ;
	input \A[629]  ;
	input \A[630]  ;
	input \A[631]  ;
	input \A[632]  ;
	input \A[633]  ;
	input \A[634]  ;
	input \A[635]  ;
	input \A[636]  ;
	input \A[637]  ;
	input \A[638]  ;
	input \A[639]  ;
	input \A[640]  ;
	input \A[641]  ;
	input \A[642]  ;
	input \A[643]  ;
	input \A[644]  ;
	input \A[645]  ;
	input \A[646]  ;
	input \A[647]  ;
	input \A[648]  ;
	input \A[649]  ;
	input \A[650]  ;
	input \A[651]  ;
	input \A[652]  ;
	input \A[653]  ;
	input \A[654]  ;
	input \A[655]  ;
	input \A[656]  ;
	input \A[657]  ;
	input \A[658]  ;
	input \A[659]  ;
	input \A[660]  ;
	input \A[661]  ;
	input \A[662]  ;
	input \A[663]  ;
	input \A[664]  ;
	input \A[665]  ;
	input \A[666]  ;
	input \A[667]  ;
	input \A[668]  ;
	input \A[669]  ;
	input \A[670]  ;
	input \A[671]  ;
	input \A[672]  ;
	input \A[673]  ;
	input \A[674]  ;
	input \A[675]  ;
	input \A[676]  ;
	input \A[677]  ;
	input \A[678]  ;
	input \A[679]  ;
	input \A[680]  ;
	input \A[681]  ;
	input \A[682]  ;
	input \A[683]  ;
	input \A[684]  ;
	input \A[685]  ;
	input \A[686]  ;
	input \A[687]  ;
	input \A[688]  ;
	input \A[689]  ;
	input \A[690]  ;
	input \A[691]  ;
	input \A[692]  ;
	input \A[693]  ;
	input \A[694]  ;
	input \A[695]  ;
	input \A[696]  ;
	input \A[697]  ;
	input \A[698]  ;
	input \A[699]  ;
	input \A[700]  ;
	input \A[701]  ;
	input \A[702]  ;
	input \A[703]  ;
	input \A[704]  ;
	input \A[705]  ;
	input \A[706]  ;
	input \A[707]  ;
	input \A[708]  ;
	input \A[709]  ;
	input \A[710]  ;
	input \A[711]  ;
	input \A[712]  ;
	input \A[713]  ;
	input \A[714]  ;
	input \A[715]  ;
	input \A[716]  ;
	input \A[717]  ;
	input \A[718]  ;
	input \A[719]  ;
	input \A[720]  ;
	input \A[721]  ;
	input \A[722]  ;
	input \A[723]  ;
	input \A[724]  ;
	input \A[725]  ;
	input \A[726]  ;
	input \A[727]  ;
	input \A[728]  ;
	input \A[729]  ;
	input \A[730]  ;
	input \A[731]  ;
	input \A[732]  ;
	input \A[733]  ;
	input \A[734]  ;
	input \A[735]  ;
	input \A[736]  ;
	input \A[737]  ;
	input \A[738]  ;
	input \A[739]  ;
	input \A[740]  ;
	input \A[741]  ;
	input \A[742]  ;
	input \A[743]  ;
	input \A[744]  ;
	input \A[745]  ;
	input \A[746]  ;
	input \A[747]  ;
	input \A[748]  ;
	input \A[749]  ;
	input \A[750]  ;
	input \A[751]  ;
	input \A[752]  ;
	input \A[753]  ;
	input \A[754]  ;
	input \A[755]  ;
	input \A[756]  ;
	input \A[757]  ;
	input \A[758]  ;
	input \A[759]  ;
	input \A[760]  ;
	input \A[761]  ;
	input \A[762]  ;
	input \A[763]  ;
	input \A[764]  ;
	input \A[765]  ;
	input \A[766]  ;
	input \A[767]  ;
	input \A[768]  ;
	input \A[769]  ;
	input \A[770]  ;
	input \A[771]  ;
	input \A[772]  ;
	input \A[773]  ;
	input \A[774]  ;
	input \A[775]  ;
	input \A[776]  ;
	input \A[777]  ;
	input \A[778]  ;
	input \A[779]  ;
	input \A[780]  ;
	input \A[781]  ;
	input \A[782]  ;
	input \A[783]  ;
	input \A[784]  ;
	input \A[785]  ;
	input \A[786]  ;
	input \A[787]  ;
	input \A[788]  ;
	input \A[789]  ;
	input \A[790]  ;
	input \A[791]  ;
	input \A[792]  ;
	input \A[793]  ;
	input \A[794]  ;
	input \A[795]  ;
	input \A[796]  ;
	input \A[797]  ;
	input \A[798]  ;
	input \A[799]  ;
	input \A[800]  ;
	input \A[801]  ;
	input \A[802]  ;
	input \A[803]  ;
	input \A[804]  ;
	input \A[805]  ;
	input \A[806]  ;
	input \A[807]  ;
	input \A[808]  ;
	input \A[809]  ;
	input \A[810]  ;
	input \A[811]  ;
	input \A[812]  ;
	input \A[813]  ;
	input \A[814]  ;
	input \A[815]  ;
	input \A[816]  ;
	input \A[817]  ;
	input \A[818]  ;
	input \A[819]  ;
	input \A[820]  ;
	input \A[821]  ;
	input \A[822]  ;
	input \A[823]  ;
	input \A[824]  ;
	input \A[825]  ;
	input \A[826]  ;
	input \A[827]  ;
	input \A[828]  ;
	input \A[829]  ;
	input \A[830]  ;
	input \A[831]  ;
	input \A[832]  ;
	input \A[833]  ;
	input \A[834]  ;
	input \A[835]  ;
	input \A[836]  ;
	input \A[837]  ;
	input \A[838]  ;
	input \A[839]  ;
	input \A[840]  ;
	input \A[841]  ;
	input \A[842]  ;
	input \A[843]  ;
	input \A[844]  ;
	input \A[845]  ;
	input \A[846]  ;
	input \A[847]  ;
	input \A[848]  ;
	input \A[849]  ;
	input \A[850]  ;
	input \A[851]  ;
	input \A[852]  ;
	input \A[853]  ;
	input \A[854]  ;
	input \A[855]  ;
	input \A[856]  ;
	input \A[857]  ;
	input \A[858]  ;
	input \A[859]  ;
	input \A[860]  ;
	input \A[861]  ;
	input \A[862]  ;
	input \A[863]  ;
	input \A[864]  ;
	input \A[865]  ;
	input \A[866]  ;
	input \A[867]  ;
	input \A[868]  ;
	input \A[869]  ;
	input \A[870]  ;
	input \A[871]  ;
	input \A[872]  ;
	input \A[873]  ;
	input \A[874]  ;
	input \A[875]  ;
	input \A[876]  ;
	input \A[877]  ;
	input \A[878]  ;
	input \A[879]  ;
	input \A[880]  ;
	input \A[881]  ;
	input \A[882]  ;
	input \A[883]  ;
	input \A[884]  ;
	input \A[885]  ;
	input \A[886]  ;
	input \A[887]  ;
	input \A[888]  ;
	input \A[889]  ;
	input \A[890]  ;
	input \A[891]  ;
	input \A[892]  ;
	input \A[893]  ;
	input \A[894]  ;
	input \A[895]  ;
	input \A[896]  ;
	input \A[897]  ;
	input \A[898]  ;
	input \A[899]  ;
	input \A[900]  ;
	input \A[901]  ;
	input \A[902]  ;
	input \A[903]  ;
	input \A[904]  ;
	input \A[905]  ;
	input \A[906]  ;
	input \A[907]  ;
	input \A[908]  ;
	input \A[909]  ;
	input \A[910]  ;
	input \A[911]  ;
	input \A[912]  ;
	input \A[913]  ;
	input \A[914]  ;
	input \A[915]  ;
	input \A[916]  ;
	input \A[917]  ;
	input \A[918]  ;
	input \A[919]  ;
	input \A[920]  ;
	input \A[921]  ;
	input \A[922]  ;
	input \A[923]  ;
	input \A[924]  ;
	input \A[925]  ;
	input \A[926]  ;
	input \A[927]  ;
	input \A[928]  ;
	input \A[929]  ;
	input \A[930]  ;
	input \A[931]  ;
	input \A[932]  ;
	input \A[933]  ;
	input \A[934]  ;
	input \A[935]  ;
	input \A[936]  ;
	input \A[937]  ;
	input \A[938]  ;
	input \A[939]  ;
	input \A[940]  ;
	input \A[941]  ;
	input \A[942]  ;
	input \A[943]  ;
	input \A[944]  ;
	input \A[945]  ;
	input \A[946]  ;
	input \A[947]  ;
	input \A[948]  ;
	input \A[949]  ;
	input \A[950]  ;
	input \A[951]  ;
	input \A[952]  ;
	input \A[953]  ;
	input \A[954]  ;
	input \A[955]  ;
	input \A[956]  ;
	input \A[957]  ;
	input \A[958]  ;
	input \A[959]  ;
	input \A[960]  ;
	input \A[961]  ;
	input \A[962]  ;
	input \A[963]  ;
	input \A[964]  ;
	input \A[965]  ;
	input \A[966]  ;
	input \A[967]  ;
	input \A[968]  ;
	input \A[969]  ;
	input \A[970]  ;
	input \A[971]  ;
	input \A[972]  ;
	input \A[973]  ;
	input \A[974]  ;
	input \A[975]  ;
	input \A[976]  ;
	input \A[977]  ;
	input \A[978]  ;
	input \A[979]  ;
	input \A[980]  ;
	input \A[981]  ;
	input \A[982]  ;
	input \A[983]  ;
	input \A[984]  ;
	input \A[985]  ;
	input \A[986]  ;
	input \A[987]  ;
	input \A[988]  ;
	input \A[989]  ;
	input \A[990]  ;
	input \A[991]  ;
	input \A[992]  ;
	input \A[993]  ;
	input \A[994]  ;
	input \A[995]  ;
	input \A[996]  ;
	input \A[997]  ;
	input \A[998]  ;
	input \A[999]  ;
	input \A[1000]  ;
	output maj ;
	wire _w9709_ ;
	wire _w9708_ ;
	wire _w9707_ ;
	wire _w9706_ ;
	wire _w9705_ ;
	wire _w9704_ ;
	wire _w9703_ ;
	wire _w9702_ ;
	wire _w9701_ ;
	wire _w9700_ ;
	wire _w9699_ ;
	wire _w9698_ ;
	wire _w9697_ ;
	wire _w9696_ ;
	wire _w9695_ ;
	wire _w9694_ ;
	wire _w9693_ ;
	wire _w9692_ ;
	wire _w9691_ ;
	wire _w9690_ ;
	wire _w9689_ ;
	wire _w9688_ ;
	wire _w9687_ ;
	wire _w9686_ ;
	wire _w9685_ ;
	wire _w9684_ ;
	wire _w9683_ ;
	wire _w9682_ ;
	wire _w9681_ ;
	wire _w9680_ ;
	wire _w9679_ ;
	wire _w9678_ ;
	wire _w9677_ ;
	wire _w9676_ ;
	wire _w9675_ ;
	wire _w9674_ ;
	wire _w9673_ ;
	wire _w9672_ ;
	wire _w9671_ ;
	wire _w9670_ ;
	wire _w9669_ ;
	wire _w9668_ ;
	wire _w9667_ ;
	wire _w9666_ ;
	wire _w9665_ ;
	wire _w9664_ ;
	wire _w9663_ ;
	wire _w9662_ ;
	wire _w9661_ ;
	wire _w9660_ ;
	wire _w9659_ ;
	wire _w9658_ ;
	wire _w9657_ ;
	wire _w9656_ ;
	wire _w9655_ ;
	wire _w9654_ ;
	wire _w9653_ ;
	wire _w9652_ ;
	wire _w9651_ ;
	wire _w9650_ ;
	wire _w9649_ ;
	wire _w9648_ ;
	wire _w9647_ ;
	wire _w9646_ ;
	wire _w9645_ ;
	wire _w9644_ ;
	wire _w9643_ ;
	wire _w9642_ ;
	wire _w9641_ ;
	wire _w9640_ ;
	wire _w9639_ ;
	wire _w9638_ ;
	wire _w9637_ ;
	wire _w9636_ ;
	wire _w9635_ ;
	wire _w9634_ ;
	wire _w9633_ ;
	wire _w9632_ ;
	wire _w9631_ ;
	wire _w9630_ ;
	wire _w9629_ ;
	wire _w9628_ ;
	wire _w9627_ ;
	wire _w9626_ ;
	wire _w9625_ ;
	wire _w9624_ ;
	wire _w9623_ ;
	wire _w9622_ ;
	wire _w9621_ ;
	wire _w9620_ ;
	wire _w9619_ ;
	wire _w9618_ ;
	wire _w9617_ ;
	wire _w9616_ ;
	wire _w9615_ ;
	wire _w9614_ ;
	wire _w9613_ ;
	wire _w9612_ ;
	wire _w9611_ ;
	wire _w9610_ ;
	wire _w9609_ ;
	wire _w9608_ ;
	wire _w9607_ ;
	wire _w9606_ ;
	wire _w9605_ ;
	wire _w9604_ ;
	wire _w9603_ ;
	wire _w9602_ ;
	wire _w9601_ ;
	wire _w9600_ ;
	wire _w9599_ ;
	wire _w9598_ ;
	wire _w9597_ ;
	wire _w9596_ ;
	wire _w9595_ ;
	wire _w9594_ ;
	wire _w9593_ ;
	wire _w9592_ ;
	wire _w9591_ ;
	wire _w9590_ ;
	wire _w9589_ ;
	wire _w9588_ ;
	wire _w9587_ ;
	wire _w9586_ ;
	wire _w9585_ ;
	wire _w9584_ ;
	wire _w9583_ ;
	wire _w9582_ ;
	wire _w9581_ ;
	wire _w9580_ ;
	wire _w9579_ ;
	wire _w9578_ ;
	wire _w9577_ ;
	wire _w9576_ ;
	wire _w9575_ ;
	wire _w9574_ ;
	wire _w9573_ ;
	wire _w9572_ ;
	wire _w9571_ ;
	wire _w9570_ ;
	wire _w9569_ ;
	wire _w9568_ ;
	wire _w9567_ ;
	wire _w9566_ ;
	wire _w9565_ ;
	wire _w9564_ ;
	wire _w9563_ ;
	wire _w9562_ ;
	wire _w9561_ ;
	wire _w9560_ ;
	wire _w9559_ ;
	wire _w9558_ ;
	wire _w9557_ ;
	wire _w9556_ ;
	wire _w9555_ ;
	wire _w9554_ ;
	wire _w9553_ ;
	wire _w9552_ ;
	wire _w9551_ ;
	wire _w9550_ ;
	wire _w9549_ ;
	wire _w9548_ ;
	wire _w9547_ ;
	wire _w9546_ ;
	wire _w9545_ ;
	wire _w9544_ ;
	wire _w9543_ ;
	wire _w9542_ ;
	wire _w9541_ ;
	wire _w9540_ ;
	wire _w9539_ ;
	wire _w9538_ ;
	wire _w9537_ ;
	wire _w9536_ ;
	wire _w9535_ ;
	wire _w9534_ ;
	wire _w9533_ ;
	wire _w9532_ ;
	wire _w9531_ ;
	wire _w9530_ ;
	wire _w9529_ ;
	wire _w9528_ ;
	wire _w9527_ ;
	wire _w9526_ ;
	wire _w9525_ ;
	wire _w9524_ ;
	wire _w9523_ ;
	wire _w9522_ ;
	wire _w9521_ ;
	wire _w9520_ ;
	wire _w9519_ ;
	wire _w9518_ ;
	wire _w9517_ ;
	wire _w9516_ ;
	wire _w9515_ ;
	wire _w9514_ ;
	wire _w9513_ ;
	wire _w9512_ ;
	wire _w9511_ ;
	wire _w9510_ ;
	wire _w9509_ ;
	wire _w9508_ ;
	wire _w9507_ ;
	wire _w9506_ ;
	wire _w9505_ ;
	wire _w9504_ ;
	wire _w9503_ ;
	wire _w9502_ ;
	wire _w9501_ ;
	wire _w9500_ ;
	wire _w9499_ ;
	wire _w9498_ ;
	wire _w9497_ ;
	wire _w9496_ ;
	wire _w9495_ ;
	wire _w9494_ ;
	wire _w9493_ ;
	wire _w9492_ ;
	wire _w9491_ ;
	wire _w9490_ ;
	wire _w9489_ ;
	wire _w9488_ ;
	wire _w9487_ ;
	wire _w9486_ ;
	wire _w9485_ ;
	wire _w9484_ ;
	wire _w9483_ ;
	wire _w9482_ ;
	wire _w9481_ ;
	wire _w9480_ ;
	wire _w9479_ ;
	wire _w9478_ ;
	wire _w9477_ ;
	wire _w9476_ ;
	wire _w9475_ ;
	wire _w9474_ ;
	wire _w9473_ ;
	wire _w9472_ ;
	wire _w9471_ ;
	wire _w9470_ ;
	wire _w9469_ ;
	wire _w9468_ ;
	wire _w9467_ ;
	wire _w9466_ ;
	wire _w9465_ ;
	wire _w9464_ ;
	wire _w9463_ ;
	wire _w9462_ ;
	wire _w9461_ ;
	wire _w9460_ ;
	wire _w9459_ ;
	wire _w9458_ ;
	wire _w9457_ ;
	wire _w9456_ ;
	wire _w9455_ ;
	wire _w9454_ ;
	wire _w9453_ ;
	wire _w9452_ ;
	wire _w9451_ ;
	wire _w9450_ ;
	wire _w9449_ ;
	wire _w9448_ ;
	wire _w9447_ ;
	wire _w9446_ ;
	wire _w9445_ ;
	wire _w9444_ ;
	wire _w9443_ ;
	wire _w9442_ ;
	wire _w9441_ ;
	wire _w9440_ ;
	wire _w9439_ ;
	wire _w9438_ ;
	wire _w9437_ ;
	wire _w9436_ ;
	wire _w9435_ ;
	wire _w9434_ ;
	wire _w9433_ ;
	wire _w9432_ ;
	wire _w9431_ ;
	wire _w9430_ ;
	wire _w9429_ ;
	wire _w9428_ ;
	wire _w9427_ ;
	wire _w9426_ ;
	wire _w9425_ ;
	wire _w9424_ ;
	wire _w9423_ ;
	wire _w9422_ ;
	wire _w9421_ ;
	wire _w9420_ ;
	wire _w9419_ ;
	wire _w9418_ ;
	wire _w9417_ ;
	wire _w9416_ ;
	wire _w9415_ ;
	wire _w9414_ ;
	wire _w9413_ ;
	wire _w9412_ ;
	wire _w9411_ ;
	wire _w9410_ ;
	wire _w9409_ ;
	wire _w9408_ ;
	wire _w9407_ ;
	wire _w9406_ ;
	wire _w9405_ ;
	wire _w9404_ ;
	wire _w9403_ ;
	wire _w9402_ ;
	wire _w9401_ ;
	wire _w9400_ ;
	wire _w9399_ ;
	wire _w9398_ ;
	wire _w9397_ ;
	wire _w9396_ ;
	wire _w9395_ ;
	wire _w9394_ ;
	wire _w9393_ ;
	wire _w9392_ ;
	wire _w9391_ ;
	wire _w9390_ ;
	wire _w9389_ ;
	wire _w9388_ ;
	wire _w9387_ ;
	wire _w9386_ ;
	wire _w9385_ ;
	wire _w9384_ ;
	wire _w9383_ ;
	wire _w9382_ ;
	wire _w9381_ ;
	wire _w9380_ ;
	wire _w9379_ ;
	wire _w9378_ ;
	wire _w9377_ ;
	wire _w9376_ ;
	wire _w9375_ ;
	wire _w9374_ ;
	wire _w9373_ ;
	wire _w9372_ ;
	wire _w9371_ ;
	wire _w9370_ ;
	wire _w9369_ ;
	wire _w9368_ ;
	wire _w9367_ ;
	wire _w9366_ ;
	wire _w9365_ ;
	wire _w9364_ ;
	wire _w9363_ ;
	wire _w9362_ ;
	wire _w9361_ ;
	wire _w9360_ ;
	wire _w9359_ ;
	wire _w9358_ ;
	wire _w9357_ ;
	wire _w9356_ ;
	wire _w9355_ ;
	wire _w9354_ ;
	wire _w9353_ ;
	wire _w9352_ ;
	wire _w9351_ ;
	wire _w9350_ ;
	wire _w9349_ ;
	wire _w9348_ ;
	wire _w9347_ ;
	wire _w9346_ ;
	wire _w9345_ ;
	wire _w9344_ ;
	wire _w9343_ ;
	wire _w9342_ ;
	wire _w9341_ ;
	wire _w9340_ ;
	wire _w9339_ ;
	wire _w9338_ ;
	wire _w9337_ ;
	wire _w9336_ ;
	wire _w9335_ ;
	wire _w9334_ ;
	wire _w9333_ ;
	wire _w9332_ ;
	wire _w9331_ ;
	wire _w9330_ ;
	wire _w9329_ ;
	wire _w9328_ ;
	wire _w9327_ ;
	wire _w9326_ ;
	wire _w9325_ ;
	wire _w9324_ ;
	wire _w9323_ ;
	wire _w9322_ ;
	wire _w9321_ ;
	wire _w9320_ ;
	wire _w9319_ ;
	wire _w9318_ ;
	wire _w9317_ ;
	wire _w9316_ ;
	wire _w9315_ ;
	wire _w9314_ ;
	wire _w9313_ ;
	wire _w9312_ ;
	wire _w9311_ ;
	wire _w9310_ ;
	wire _w9309_ ;
	wire _w9308_ ;
	wire _w9307_ ;
	wire _w9306_ ;
	wire _w9305_ ;
	wire _w9304_ ;
	wire _w9303_ ;
	wire _w9302_ ;
	wire _w9301_ ;
	wire _w9300_ ;
	wire _w9299_ ;
	wire _w9298_ ;
	wire _w9297_ ;
	wire _w9296_ ;
	wire _w9295_ ;
	wire _w9294_ ;
	wire _w9293_ ;
	wire _w9292_ ;
	wire _w9291_ ;
	wire _w9290_ ;
	wire _w9289_ ;
	wire _w9288_ ;
	wire _w9287_ ;
	wire _w9286_ ;
	wire _w9285_ ;
	wire _w9284_ ;
	wire _w9283_ ;
	wire _w9282_ ;
	wire _w9281_ ;
	wire _w9280_ ;
	wire _w9279_ ;
	wire _w9278_ ;
	wire _w9277_ ;
	wire _w9276_ ;
	wire _w9275_ ;
	wire _w9274_ ;
	wire _w9273_ ;
	wire _w9272_ ;
	wire _w9271_ ;
	wire _w9270_ ;
	wire _w9269_ ;
	wire _w9268_ ;
	wire _w9267_ ;
	wire _w9266_ ;
	wire _w9265_ ;
	wire _w9264_ ;
	wire _w9263_ ;
	wire _w9262_ ;
	wire _w9261_ ;
	wire _w9260_ ;
	wire _w9259_ ;
	wire _w9258_ ;
	wire _w9257_ ;
	wire _w9256_ ;
	wire _w9255_ ;
	wire _w9254_ ;
	wire _w9253_ ;
	wire _w9252_ ;
	wire _w9251_ ;
	wire _w9250_ ;
	wire _w9249_ ;
	wire _w9248_ ;
	wire _w9247_ ;
	wire _w9246_ ;
	wire _w9245_ ;
	wire _w9244_ ;
	wire _w9243_ ;
	wire _w9242_ ;
	wire _w9241_ ;
	wire _w9240_ ;
	wire _w9239_ ;
	wire _w9238_ ;
	wire _w9237_ ;
	wire _w9236_ ;
	wire _w9235_ ;
	wire _w9234_ ;
	wire _w9233_ ;
	wire _w9232_ ;
	wire _w9231_ ;
	wire _w9230_ ;
	wire _w9229_ ;
	wire _w9228_ ;
	wire _w9227_ ;
	wire _w9226_ ;
	wire _w9225_ ;
	wire _w9224_ ;
	wire _w9223_ ;
	wire _w9222_ ;
	wire _w9221_ ;
	wire _w9220_ ;
	wire _w9219_ ;
	wire _w9218_ ;
	wire _w9217_ ;
	wire _w9216_ ;
	wire _w9215_ ;
	wire _w9214_ ;
	wire _w9213_ ;
	wire _w9212_ ;
	wire _w9211_ ;
	wire _w9210_ ;
	wire _w9209_ ;
	wire _w9208_ ;
	wire _w9207_ ;
	wire _w9206_ ;
	wire _w9205_ ;
	wire _w9204_ ;
	wire _w9203_ ;
	wire _w9202_ ;
	wire _w9201_ ;
	wire _w9200_ ;
	wire _w9199_ ;
	wire _w9198_ ;
	wire _w9197_ ;
	wire _w9196_ ;
	wire _w9195_ ;
	wire _w9194_ ;
	wire _w9193_ ;
	wire _w9192_ ;
	wire _w9191_ ;
	wire _w9190_ ;
	wire _w9189_ ;
	wire _w9188_ ;
	wire _w9187_ ;
	wire _w9186_ ;
	wire _w9185_ ;
	wire _w9184_ ;
	wire _w9183_ ;
	wire _w9182_ ;
	wire _w9181_ ;
	wire _w9180_ ;
	wire _w9179_ ;
	wire _w9178_ ;
	wire _w9177_ ;
	wire _w9176_ ;
	wire _w9175_ ;
	wire _w9174_ ;
	wire _w9173_ ;
	wire _w9172_ ;
	wire _w9171_ ;
	wire _w9170_ ;
	wire _w9169_ ;
	wire _w9168_ ;
	wire _w9167_ ;
	wire _w9166_ ;
	wire _w9165_ ;
	wire _w9164_ ;
	wire _w9163_ ;
	wire _w9162_ ;
	wire _w9161_ ;
	wire _w9160_ ;
	wire _w9159_ ;
	wire _w9158_ ;
	wire _w9157_ ;
	wire _w9156_ ;
	wire _w9155_ ;
	wire _w9154_ ;
	wire _w9153_ ;
	wire _w9152_ ;
	wire _w9151_ ;
	wire _w9150_ ;
	wire _w9149_ ;
	wire _w9148_ ;
	wire _w9147_ ;
	wire _w9146_ ;
	wire _w9145_ ;
	wire _w9144_ ;
	wire _w9143_ ;
	wire _w9142_ ;
	wire _w9141_ ;
	wire _w9140_ ;
	wire _w9139_ ;
	wire _w9138_ ;
	wire _w9137_ ;
	wire _w9136_ ;
	wire _w9135_ ;
	wire _w9134_ ;
	wire _w9133_ ;
	wire _w9132_ ;
	wire _w9131_ ;
	wire _w9130_ ;
	wire _w9129_ ;
	wire _w9128_ ;
	wire _w9127_ ;
	wire _w9126_ ;
	wire _w9125_ ;
	wire _w9124_ ;
	wire _w9123_ ;
	wire _w9122_ ;
	wire _w9121_ ;
	wire _w9120_ ;
	wire _w9119_ ;
	wire _w9118_ ;
	wire _w9117_ ;
	wire _w9116_ ;
	wire _w9115_ ;
	wire _w9114_ ;
	wire _w9113_ ;
	wire _w9112_ ;
	wire _w9111_ ;
	wire _w9110_ ;
	wire _w9109_ ;
	wire _w9108_ ;
	wire _w9107_ ;
	wire _w9106_ ;
	wire _w9105_ ;
	wire _w9104_ ;
	wire _w9103_ ;
	wire _w9102_ ;
	wire _w9101_ ;
	wire _w9100_ ;
	wire _w9099_ ;
	wire _w9098_ ;
	wire _w9097_ ;
	wire _w9096_ ;
	wire _w9095_ ;
	wire _w9094_ ;
	wire _w9093_ ;
	wire _w9092_ ;
	wire _w9091_ ;
	wire _w9090_ ;
	wire _w9089_ ;
	wire _w9088_ ;
	wire _w9087_ ;
	wire _w9086_ ;
	wire _w9085_ ;
	wire _w9084_ ;
	wire _w9083_ ;
	wire _w9082_ ;
	wire _w9081_ ;
	wire _w9080_ ;
	wire _w9079_ ;
	wire _w9078_ ;
	wire _w9077_ ;
	wire _w9076_ ;
	wire _w9075_ ;
	wire _w9074_ ;
	wire _w9073_ ;
	wire _w9072_ ;
	wire _w9071_ ;
	wire _w9070_ ;
	wire _w9069_ ;
	wire _w9068_ ;
	wire _w9067_ ;
	wire _w9066_ ;
	wire _w9065_ ;
	wire _w9064_ ;
	wire _w9063_ ;
	wire _w9062_ ;
	wire _w9061_ ;
	wire _w9060_ ;
	wire _w9059_ ;
	wire _w9058_ ;
	wire _w9057_ ;
	wire _w9056_ ;
	wire _w9055_ ;
	wire _w9054_ ;
	wire _w9053_ ;
	wire _w9052_ ;
	wire _w9051_ ;
	wire _w9050_ ;
	wire _w9049_ ;
	wire _w9048_ ;
	wire _w9047_ ;
	wire _w9046_ ;
	wire _w9045_ ;
	wire _w9044_ ;
	wire _w9043_ ;
	wire _w9042_ ;
	wire _w9041_ ;
	wire _w9040_ ;
	wire _w9039_ ;
	wire _w9038_ ;
	wire _w9037_ ;
	wire _w9036_ ;
	wire _w9035_ ;
	wire _w9034_ ;
	wire _w9033_ ;
	wire _w9032_ ;
	wire _w9031_ ;
	wire _w9030_ ;
	wire _w9029_ ;
	wire _w9028_ ;
	wire _w9027_ ;
	wire _w9026_ ;
	wire _w9025_ ;
	wire _w9024_ ;
	wire _w9023_ ;
	wire _w9022_ ;
	wire _w9021_ ;
	wire _w9020_ ;
	wire _w9019_ ;
	wire _w9018_ ;
	wire _w9017_ ;
	wire _w9016_ ;
	wire _w9015_ ;
	wire _w9014_ ;
	wire _w9013_ ;
	wire _w9012_ ;
	wire _w9011_ ;
	wire _w9010_ ;
	wire _w9009_ ;
	wire _w9008_ ;
	wire _w9007_ ;
	wire _w9006_ ;
	wire _w9005_ ;
	wire _w9004_ ;
	wire _w9003_ ;
	wire _w9002_ ;
	wire _w9001_ ;
	wire _w9000_ ;
	wire _w8999_ ;
	wire _w8998_ ;
	wire _w8997_ ;
	wire _w8996_ ;
	wire _w8995_ ;
	wire _w8994_ ;
	wire _w8993_ ;
	wire _w8992_ ;
	wire _w8991_ ;
	wire _w8990_ ;
	wire _w8989_ ;
	wire _w8988_ ;
	wire _w8987_ ;
	wire _w8986_ ;
	wire _w8985_ ;
	wire _w8984_ ;
	wire _w8983_ ;
	wire _w8982_ ;
	wire _w8981_ ;
	wire _w8980_ ;
	wire _w8979_ ;
	wire _w8978_ ;
	wire _w8977_ ;
	wire _w8976_ ;
	wire _w8975_ ;
	wire _w8974_ ;
	wire _w8973_ ;
	wire _w8972_ ;
	wire _w8971_ ;
	wire _w8970_ ;
	wire _w8969_ ;
	wire _w8968_ ;
	wire _w8967_ ;
	wire _w8966_ ;
	wire _w8965_ ;
	wire _w8964_ ;
	wire _w8963_ ;
	wire _w8962_ ;
	wire _w8961_ ;
	wire _w8960_ ;
	wire _w8959_ ;
	wire _w8958_ ;
	wire _w8957_ ;
	wire _w8956_ ;
	wire _w8955_ ;
	wire _w8954_ ;
	wire _w8953_ ;
	wire _w8952_ ;
	wire _w8951_ ;
	wire _w8950_ ;
	wire _w8949_ ;
	wire _w8948_ ;
	wire _w8947_ ;
	wire _w8946_ ;
	wire _w8945_ ;
	wire _w8944_ ;
	wire _w8943_ ;
	wire _w8942_ ;
	wire _w8941_ ;
	wire _w8940_ ;
	wire _w8939_ ;
	wire _w8938_ ;
	wire _w8937_ ;
	wire _w8936_ ;
	wire _w8935_ ;
	wire _w8934_ ;
	wire _w8933_ ;
	wire _w8932_ ;
	wire _w8931_ ;
	wire _w8930_ ;
	wire _w8929_ ;
	wire _w8928_ ;
	wire _w8927_ ;
	wire _w8926_ ;
	wire _w8925_ ;
	wire _w8924_ ;
	wire _w8923_ ;
	wire _w8922_ ;
	wire _w8921_ ;
	wire _w8920_ ;
	wire _w8919_ ;
	wire _w8918_ ;
	wire _w8917_ ;
	wire _w8916_ ;
	wire _w8915_ ;
	wire _w8914_ ;
	wire _w8913_ ;
	wire _w8912_ ;
	wire _w8911_ ;
	wire _w8910_ ;
	wire _w8909_ ;
	wire _w8908_ ;
	wire _w8907_ ;
	wire _w8906_ ;
	wire _w8905_ ;
	wire _w8904_ ;
	wire _w8903_ ;
	wire _w8902_ ;
	wire _w8901_ ;
	wire _w8900_ ;
	wire _w8899_ ;
	wire _w8898_ ;
	wire _w8897_ ;
	wire _w8896_ ;
	wire _w8895_ ;
	wire _w8894_ ;
	wire _w8893_ ;
	wire _w8892_ ;
	wire _w8891_ ;
	wire _w8890_ ;
	wire _w8889_ ;
	wire _w8888_ ;
	wire _w8887_ ;
	wire _w8886_ ;
	wire _w8885_ ;
	wire _w8884_ ;
	wire _w8883_ ;
	wire _w8882_ ;
	wire _w8881_ ;
	wire _w8880_ ;
	wire _w8879_ ;
	wire _w8878_ ;
	wire _w8877_ ;
	wire _w8876_ ;
	wire _w8875_ ;
	wire _w8874_ ;
	wire _w8873_ ;
	wire _w8872_ ;
	wire _w8871_ ;
	wire _w8870_ ;
	wire _w8869_ ;
	wire _w8868_ ;
	wire _w8867_ ;
	wire _w8866_ ;
	wire _w8865_ ;
	wire _w8864_ ;
	wire _w8863_ ;
	wire _w8862_ ;
	wire _w8861_ ;
	wire _w8860_ ;
	wire _w8859_ ;
	wire _w8858_ ;
	wire _w8857_ ;
	wire _w8856_ ;
	wire _w8855_ ;
	wire _w8854_ ;
	wire _w8853_ ;
	wire _w8852_ ;
	wire _w8851_ ;
	wire _w8850_ ;
	wire _w8849_ ;
	wire _w8848_ ;
	wire _w8847_ ;
	wire _w8846_ ;
	wire _w8845_ ;
	wire _w8844_ ;
	wire _w8843_ ;
	wire _w8842_ ;
	wire _w8841_ ;
	wire _w8840_ ;
	wire _w8839_ ;
	wire _w8838_ ;
	wire _w8837_ ;
	wire _w8836_ ;
	wire _w8835_ ;
	wire _w8834_ ;
	wire _w8833_ ;
	wire _w8832_ ;
	wire _w8831_ ;
	wire _w8830_ ;
	wire _w8829_ ;
	wire _w8828_ ;
	wire _w8827_ ;
	wire _w8826_ ;
	wire _w8825_ ;
	wire _w8824_ ;
	wire _w8823_ ;
	wire _w8822_ ;
	wire _w8821_ ;
	wire _w8820_ ;
	wire _w8819_ ;
	wire _w8818_ ;
	wire _w8817_ ;
	wire _w8816_ ;
	wire _w8815_ ;
	wire _w8814_ ;
	wire _w8813_ ;
	wire _w8812_ ;
	wire _w8811_ ;
	wire _w8810_ ;
	wire _w8809_ ;
	wire _w8808_ ;
	wire _w8807_ ;
	wire _w8806_ ;
	wire _w8805_ ;
	wire _w8804_ ;
	wire _w8803_ ;
	wire _w8802_ ;
	wire _w8801_ ;
	wire _w8800_ ;
	wire _w8799_ ;
	wire _w8798_ ;
	wire _w8797_ ;
	wire _w8796_ ;
	wire _w8795_ ;
	wire _w8794_ ;
	wire _w8793_ ;
	wire _w8792_ ;
	wire _w8791_ ;
	wire _w8790_ ;
	wire _w8789_ ;
	wire _w8788_ ;
	wire _w8787_ ;
	wire _w8786_ ;
	wire _w8785_ ;
	wire _w8784_ ;
	wire _w8783_ ;
	wire _w8782_ ;
	wire _w8781_ ;
	wire _w8780_ ;
	wire _w8779_ ;
	wire _w8778_ ;
	wire _w8777_ ;
	wire _w8776_ ;
	wire _w8775_ ;
	wire _w8774_ ;
	wire _w8773_ ;
	wire _w8772_ ;
	wire _w8771_ ;
	wire _w8770_ ;
	wire _w8769_ ;
	wire _w8768_ ;
	wire _w8767_ ;
	wire _w8766_ ;
	wire _w8765_ ;
	wire _w8764_ ;
	wire _w8763_ ;
	wire _w8762_ ;
	wire _w8761_ ;
	wire _w8760_ ;
	wire _w8759_ ;
	wire _w8758_ ;
	wire _w8757_ ;
	wire _w8756_ ;
	wire _w8755_ ;
	wire _w8754_ ;
	wire _w8753_ ;
	wire _w8752_ ;
	wire _w8751_ ;
	wire _w8750_ ;
	wire _w8749_ ;
	wire _w8748_ ;
	wire _w8747_ ;
	wire _w8746_ ;
	wire _w8745_ ;
	wire _w8744_ ;
	wire _w8743_ ;
	wire _w8742_ ;
	wire _w8741_ ;
	wire _w8740_ ;
	wire _w8739_ ;
	wire _w8738_ ;
	wire _w8737_ ;
	wire _w8736_ ;
	wire _w8735_ ;
	wire _w8734_ ;
	wire _w8733_ ;
	wire _w8732_ ;
	wire _w8731_ ;
	wire _w8730_ ;
	wire _w8729_ ;
	wire _w8728_ ;
	wire _w8727_ ;
	wire _w8726_ ;
	wire _w8725_ ;
	wire _w8724_ ;
	wire _w8723_ ;
	wire _w8722_ ;
	wire _w8721_ ;
	wire _w8720_ ;
	wire _w8719_ ;
	wire _w8718_ ;
	wire _w8717_ ;
	wire _w8716_ ;
	wire _w8715_ ;
	wire _w8714_ ;
	wire _w8713_ ;
	wire _w8712_ ;
	wire _w8711_ ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w6594_ ;
	wire _w6593_ ;
	wire _w6592_ ;
	wire _w6591_ ;
	wire _w6590_ ;
	wire _w6589_ ;
	wire _w6588_ ;
	wire _w6587_ ;
	wire _w6586_ ;
	wire _w6585_ ;
	wire _w6584_ ;
	wire _w6583_ ;
	wire _w6582_ ;
	wire _w6581_ ;
	wire _w6580_ ;
	wire _w6579_ ;
	wire _w6578_ ;
	wire _w6577_ ;
	wire _w6576_ ;
	wire _w6575_ ;
	wire _w6574_ ;
	wire _w6573_ ;
	wire _w6572_ ;
	wire _w6571_ ;
	wire _w6570_ ;
	wire _w6569_ ;
	wire _w6568_ ;
	wire _w6567_ ;
	wire _w6566_ ;
	wire _w6565_ ;
	wire _w6564_ ;
	wire _w6563_ ;
	wire _w6562_ ;
	wire _w6561_ ;
	wire _w6560_ ;
	wire _w6559_ ;
	wire _w6558_ ;
	wire _w6557_ ;
	wire _w6556_ ;
	wire _w6555_ ;
	wire _w6554_ ;
	wire _w6553_ ;
	wire _w6552_ ;
	wire _w6551_ ;
	wire _w6550_ ;
	wire _w6549_ ;
	wire _w6548_ ;
	wire _w6547_ ;
	wire _w6546_ ;
	wire _w6545_ ;
	wire _w6544_ ;
	wire _w6543_ ;
	wire _w6542_ ;
	wire _w6541_ ;
	wire _w6540_ ;
	wire _w6539_ ;
	wire _w6538_ ;
	wire _w6537_ ;
	wire _w6536_ ;
	wire _w6535_ ;
	wire _w6534_ ;
	wire _w6533_ ;
	wire _w6532_ ;
	wire _w6531_ ;
	wire _w6530_ ;
	wire _w6529_ ;
	wire _w6528_ ;
	wire _w6527_ ;
	wire _w6526_ ;
	wire _w6525_ ;
	wire _w6524_ ;
	wire _w6523_ ;
	wire _w6522_ ;
	wire _w6521_ ;
	wire _w6520_ ;
	wire _w6519_ ;
	wire _w6518_ ;
	wire _w6517_ ;
	wire _w6516_ ;
	wire _w6515_ ;
	wire _w6514_ ;
	wire _w6513_ ;
	wire _w6512_ ;
	wire _w6511_ ;
	wire _w6510_ ;
	wire _w6509_ ;
	wire _w6508_ ;
	wire _w6507_ ;
	wire _w6506_ ;
	wire _w6505_ ;
	wire _w6504_ ;
	wire _w6503_ ;
	wire _w6502_ ;
	wire _w6501_ ;
	wire _w6500_ ;
	wire _w6499_ ;
	wire _w6498_ ;
	wire _w6497_ ;
	wire _w6496_ ;
	wire _w6495_ ;
	wire _w6494_ ;
	wire _w6493_ ;
	wire _w6492_ ;
	wire _w6491_ ;
	wire _w6490_ ;
	wire _w6489_ ;
	wire _w6488_ ;
	wire _w6487_ ;
	wire _w6486_ ;
	wire _w6485_ ;
	wire _w6484_ ;
	wire _w6483_ ;
	wire _w6482_ ;
	wire _w6481_ ;
	wire _w6480_ ;
	wire _w6479_ ;
	wire _w6478_ ;
	wire _w6477_ ;
	wire _w6476_ ;
	wire _w6475_ ;
	wire _w6474_ ;
	wire _w6473_ ;
	wire _w6472_ ;
	wire _w6471_ ;
	wire _w6470_ ;
	wire _w6469_ ;
	wire _w6468_ ;
	wire _w6467_ ;
	wire _w6466_ ;
	wire _w6465_ ;
	wire _w6464_ ;
	wire _w6463_ ;
	wire _w6462_ ;
	wire _w6461_ ;
	wire _w6460_ ;
	wire _w6459_ ;
	wire _w6458_ ;
	wire _w6457_ ;
	wire _w6456_ ;
	wire _w6455_ ;
	wire _w6454_ ;
	wire _w6453_ ;
	wire _w6452_ ;
	wire _w6451_ ;
	wire _w6450_ ;
	wire _w6449_ ;
	wire _w6448_ ;
	wire _w6447_ ;
	wire _w6446_ ;
	wire _w6445_ ;
	wire _w6444_ ;
	wire _w6443_ ;
	wire _w6442_ ;
	wire _w6441_ ;
	wire _w6440_ ;
	wire _w6439_ ;
	wire _w6438_ ;
	wire _w6437_ ;
	wire _w6436_ ;
	wire _w6435_ ;
	wire _w6434_ ;
	wire _w6433_ ;
	wire _w6432_ ;
	wire _w6431_ ;
	wire _w6430_ ;
	wire _w6429_ ;
	wire _w6428_ ;
	wire _w6427_ ;
	wire _w6426_ ;
	wire _w6425_ ;
	wire _w6424_ ;
	wire _w6423_ ;
	wire _w6422_ ;
	wire _w6421_ ;
	wire _w6420_ ;
	wire _w6419_ ;
	wire _w6418_ ;
	wire _w6417_ ;
	wire _w6416_ ;
	wire _w6415_ ;
	wire _w6414_ ;
	wire _w6413_ ;
	wire _w6412_ ;
	wire _w6411_ ;
	wire _w6410_ ;
	wire _w6409_ ;
	wire _w6408_ ;
	wire _w6407_ ;
	wire _w6406_ ;
	wire _w6405_ ;
	wire _w6404_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w1542_ ;
	wire _w1541_ ;
	wire _w1540_ ;
	wire _w1539_ ;
	wire _w1538_ ;
	wire _w1537_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1520_ ;
	wire _w1519_ ;
	wire _w1518_ ;
	wire _w1517_ ;
	wire _w1516_ ;
	wire _w1515_ ;
	wire _w1514_ ;
	wire _w1513_ ;
	wire _w1512_ ;
	wire _w1511_ ;
	wire _w1510_ ;
	wire _w1509_ ;
	wire _w1508_ ;
	wire _w1507_ ;
	wire _w1506_ ;
	wire _w1505_ ;
	wire _w1504_ ;
	wire _w1503_ ;
	wire _w1502_ ;
	wire _w1501_ ;
	wire _w1500_ ;
	wire _w1499_ ;
	wire _w1498_ ;
	wire _w1497_ ;
	wire _w1496_ ;
	wire _w1495_ ;
	wire _w1494_ ;
	wire _w1493_ ;
	wire _w1492_ ;
	wire _w1491_ ;
	wire _w1490_ ;
	wire _w1489_ ;
	wire _w1488_ ;
	wire _w1487_ ;
	wire _w1486_ ;
	wire _w1485_ ;
	wire _w1484_ ;
	wire _w1483_ ;
	wire _w1482_ ;
	wire _w1481_ ;
	wire _w1480_ ;
	wire _w1479_ ;
	wire _w1478_ ;
	wire _w1477_ ;
	wire _w1476_ ;
	wire _w1475_ ;
	wire _w1474_ ;
	wire _w1473_ ;
	wire _w1472_ ;
	wire _w1471_ ;
	wire _w1470_ ;
	wire _w1469_ ;
	wire _w1468_ ;
	wire _w1467_ ;
	wire _w1466_ ;
	wire _w1465_ ;
	wire _w1464_ ;
	wire _w1463_ ;
	wire _w1462_ ;
	wire _w1461_ ;
	wire _w1460_ ;
	wire _w1459_ ;
	wire _w1458_ ;
	wire _w1457_ ;
	wire _w1456_ ;
	wire _w1455_ ;
	wire _w1454_ ;
	wire _w1453_ ;
	wire _w1452_ ;
	wire _w1451_ ;
	wire _w1450_ ;
	wire _w1449_ ;
	wire _w1448_ ;
	wire _w1447_ ;
	wire _w1446_ ;
	wire _w1445_ ;
	wire _w1444_ ;
	wire _w1443_ ;
	wire _w1442_ ;
	wire _w1441_ ;
	wire _w1440_ ;
	wire _w1439_ ;
	wire _w1438_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1419_ ;
	wire _w1418_ ;
	wire _w1417_ ;
	wire _w1416_ ;
	wire _w1415_ ;
	wire _w1414_ ;
	wire _w1413_ ;
	wire _w1412_ ;
	wire _w1411_ ;
	wire _w1410_ ;
	wire _w1409_ ;
	wire _w1408_ ;
	wire _w1407_ ;
	wire _w1406_ ;
	wire _w1405_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1398_ ;
	wire _w1397_ ;
	wire _w1396_ ;
	wire _w1395_ ;
	wire _w1394_ ;
	wire _w1393_ ;
	wire _w1392_ ;
	wire _w1391_ ;
	wire _w1390_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1387_ ;
	wire _w1386_ ;
	wire _w1385_ ;
	wire _w1384_ ;
	wire _w1383_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1374_ ;
	wire _w1373_ ;
	wire _w1372_ ;
	wire _w1371_ ;
	wire _w1370_ ;
	wire _w1369_ ;
	wire _w1368_ ;
	wire _w1367_ ;
	wire _w1366_ ;
	wire _w1365_ ;
	wire _w1364_ ;
	wire _w1363_ ;
	wire _w1362_ ;
	wire _w1361_ ;
	wire _w1360_ ;
	wire _w1359_ ;
	wire _w1358_ ;
	wire _w1357_ ;
	wire _w1356_ ;
	wire _w1355_ ;
	wire _w1354_ ;
	wire _w1353_ ;
	wire _w1352_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1348_ ;
	wire _w1347_ ;
	wire _w1346_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1343_ ;
	wire _w1342_ ;
	wire _w1341_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1338_ ;
	wire _w1337_ ;
	wire _w1336_ ;
	wire _w1335_ ;
	wire _w1334_ ;
	wire _w1333_ ;
	wire _w1332_ ;
	wire _w1331_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1328_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1325_ ;
	wire _w1324_ ;
	wire _w1323_ ;
	wire _w1322_ ;
	wire _w1321_ ;
	wire _w1320_ ;
	wire _w1319_ ;
	wire _w1318_ ;
	wire _w1317_ ;
	wire _w1316_ ;
	wire _w1315_ ;
	wire _w1314_ ;
	wire _w1313_ ;
	wire _w1312_ ;
	wire _w1311_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1307_ ;
	wire _w1306_ ;
	wire _w1305_ ;
	wire _w1304_ ;
	wire _w1303_ ;
	wire _w1302_ ;
	wire _w1301_ ;
	wire _w1300_ ;
	wire _w1299_ ;
	wire _w1298_ ;
	wire _w1297_ ;
	wire _w1296_ ;
	wire _w1295_ ;
	wire _w1294_ ;
	wire _w1293_ ;
	wire _w1292_ ;
	wire _w1291_ ;
	wire _w1290_ ;
	wire _w1289_ ;
	wire _w1288_ ;
	wire _w1287_ ;
	wire _w1286_ ;
	wire _w1285_ ;
	wire _w1284_ ;
	wire _w1283_ ;
	wire _w1282_ ;
	wire _w1281_ ;
	wire _w1280_ ;
	wire _w1279_ ;
	wire _w1278_ ;
	wire _w1277_ ;
	wire _w1276_ ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1002_ ;
	wire _w1003_ ;
	wire _w1004_ ;
	wire _w1005_ ;
	wire _w1006_ ;
	wire _w1007_ ;
	wire _w1008_ ;
	wire _w1009_ ;
	wire _w1010_ ;
	wire _w1011_ ;
	wire _w1012_ ;
	wire _w1013_ ;
	wire _w1014_ ;
	wire _w1031_ ;
	wire _w1032_ ;
	wire _w1033_ ;
	wire _w1034_ ;
	wire _w1035_ ;
	wire _w1036_ ;
	wire _w1037_ ;
	wire _w1038_ ;
	wire _w1039_ ;
	wire _w1040_ ;
	wire _w1041_ ;
	wire _w1042_ ;
	wire _w1043_ ;
	wire _w1044_ ;
	wire _w1045_ ;
	wire _w1046_ ;
	wire _w1047_ ;
	wire _w1048_ ;
	wire _w1049_ ;
	wire _w1050_ ;
	wire _w1051_ ;
	wire _w1052_ ;
	wire _w1053_ ;
	wire _w1054_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1623_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1626_ ;
	wire _w1627_ ;
	wire _w1628_ ;
	wire _w1629_ ;
	wire _w1630_ ;
	wire _w1631_ ;
	wire _w1632_ ;
	wire _w1633_ ;
	wire _w1634_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w1765_ ;
	wire _w1766_ ;
	wire _w1767_ ;
	wire _w1768_ ;
	wire _w1769_ ;
	wire _w1770_ ;
	wire _w1771_ ;
	wire _w1772_ ;
	wire _w1773_ ;
	wire _w1774_ ;
	wire _w1775_ ;
	wire _w1776_ ;
	wire _w1777_ ;
	wire _w1778_ ;
	wire _w1779_ ;
	wire _w1780_ ;
	wire _w1781_ ;
	wire _w1782_ ;
	wire _w1783_ ;
	wire _w1784_ ;
	wire _w1785_ ;
	wire _w1786_ ;
	wire _w1787_ ;
	wire _w1788_ ;
	wire _w1789_ ;
	wire _w1790_ ;
	wire _w1791_ ;
	wire _w1792_ ;
	wire _w1793_ ;
	wire _w1794_ ;
	wire _w1795_ ;
	wire _w1796_ ;
	wire _w1797_ ;
	wire _w1798_ ;
	wire _w1799_ ;
	wire _w1800_ ;
	wire _w1801_ ;
	wire _w1802_ ;
	wire _w1803_ ;
	wire _w1804_ ;
	wire _w1805_ ;
	wire _w1806_ ;
	wire _w1807_ ;
	wire _w1808_ ;
	wire _w1809_ ;
	wire _w1810_ ;
	wire _w1811_ ;
	wire _w1812_ ;
	wire _w1813_ ;
	wire _w1814_ ;
	wire _w1815_ ;
	wire _w1816_ ;
	wire _w1817_ ;
	wire _w1818_ ;
	wire _w1819_ ;
	wire _w1820_ ;
	wire _w1821_ ;
	wire _w1822_ ;
	wire _w1823_ ;
	wire _w1824_ ;
	wire _w1825_ ;
	wire _w1826_ ;
	wire _w1827_ ;
	wire _w1828_ ;
	wire _w1829_ ;
	wire _w1830_ ;
	wire _w1831_ ;
	wire _w1832_ ;
	wire _w1833_ ;
	wire _w1834_ ;
	wire _w1835_ ;
	wire _w1836_ ;
	wire _w1837_ ;
	wire _w1838_ ;
	wire _w1839_ ;
	wire _w1840_ ;
	wire _w1841_ ;
	wire _w1842_ ;
	wire _w1843_ ;
	wire _w1844_ ;
	wire _w1845_ ;
	wire _w1846_ ;
	wire _w1847_ ;
	wire _w1848_ ;
	wire _w1849_ ;
	wire _w1850_ ;
	wire _w1851_ ;
	wire _w1852_ ;
	wire _w1853_ ;
	wire _w1854_ ;
	wire _w1855_ ;
	wire _w1856_ ;
	wire _w1857_ ;
	wire _w1858_ ;
	wire _w1859_ ;
	wire _w1860_ ;
	wire _w1861_ ;
	wire _w1862_ ;
	wire _w1863_ ;
	wire _w1864_ ;
	wire _w1865_ ;
	wire _w1866_ ;
	wire _w1867_ ;
	wire _w1868_ ;
	wire _w1869_ ;
	wire _w1870_ ;
	wire _w1871_ ;
	wire _w1872_ ;
	wire _w1873_ ;
	wire _w1874_ ;
	wire _w1875_ ;
	wire _w1876_ ;
	wire _w1877_ ;
	wire _w1878_ ;
	wire _w1879_ ;
	wire _w1880_ ;
	wire _w1881_ ;
	wire _w1882_ ;
	wire _w1883_ ;
	wire _w1884_ ;
	wire _w1885_ ;
	wire _w1886_ ;
	wire _w1887_ ;
	wire _w1888_ ;
	wire _w1889_ ;
	wire _w1890_ ;
	wire _w1891_ ;
	wire _w1892_ ;
	wire _w1893_ ;
	wire _w1894_ ;
	wire _w1895_ ;
	wire _w1896_ ;
	wire _w1897_ ;
	wire _w1898_ ;
	wire _w1899_ ;
	wire _w1900_ ;
	wire _w1901_ ;
	wire _w1902_ ;
	wire _w1903_ ;
	wire _w1904_ ;
	wire _w1905_ ;
	wire _w1906_ ;
	wire _w1907_ ;
	wire _w1908_ ;
	wire _w1909_ ;
	wire _w1910_ ;
	wire _w1911_ ;
	wire _w1912_ ;
	wire _w1913_ ;
	wire _w1914_ ;
	wire _w1915_ ;
	wire _w1916_ ;
	wire _w1917_ ;
	wire _w1918_ ;
	wire _w1919_ ;
	wire _w1920_ ;
	wire _w1921_ ;
	wire _w1922_ ;
	wire _w1923_ ;
	wire _w1924_ ;
	wire _w1925_ ;
	wire _w1926_ ;
	wire _w1927_ ;
	wire _w1928_ ;
	wire _w1929_ ;
	wire _w1930_ ;
	wire _w1931_ ;
	wire _w1932_ ;
	wire _w1933_ ;
	wire _w1934_ ;
	wire _w1935_ ;
	wire _w1936_ ;
	wire _w1937_ ;
	wire _w1938_ ;
	wire _w1939_ ;
	wire _w1940_ ;
	wire _w1941_ ;
	wire _w1942_ ;
	wire _w1943_ ;
	wire _w1944_ ;
	wire _w1945_ ;
	wire _w1946_ ;
	wire _w1947_ ;
	wire _w1948_ ;
	wire _w1949_ ;
	wire _w1950_ ;
	wire _w1951_ ;
	wire _w1952_ ;
	wire _w1953_ ;
	wire _w1954_ ;
	wire _w1955_ ;
	wire _w1956_ ;
	wire _w1957_ ;
	wire _w1958_ ;
	wire _w1959_ ;
	wire _w1960_ ;
	wire _w1961_ ;
	wire _w1962_ ;
	wire _w1963_ ;
	wire _w1964_ ;
	wire _w1965_ ;
	wire _w1966_ ;
	wire _w1967_ ;
	wire _w1968_ ;
	wire _w1969_ ;
	wire _w1970_ ;
	wire _w1971_ ;
	wire _w1972_ ;
	wire _w1973_ ;
	wire _w1974_ ;
	wire _w1975_ ;
	wire _w1976_ ;
	wire _w1977_ ;
	wire _w1978_ ;
	wire _w1979_ ;
	wire _w1980_ ;
	wire _w1981_ ;
	wire _w1982_ ;
	wire _w1983_ ;
	wire _w1984_ ;
	wire _w1985_ ;
	wire _w1986_ ;
	wire _w1987_ ;
	wire _w1988_ ;
	wire _w1989_ ;
	wire _w1990_ ;
	wire _w1991_ ;
	wire _w1992_ ;
	wire _w1993_ ;
	wire _w1994_ ;
	wire _w1995_ ;
	wire _w1996_ ;
	wire _w1997_ ;
	wire _w1998_ ;
	wire _w1999_ ;
	wire _w2000_ ;
	wire _w2001_ ;
	wire _w2002_ ;
	wire _w2003_ ;
	wire _w2004_ ;
	wire _w2005_ ;
	wire _w2006_ ;
	wire _w2007_ ;
	wire _w2008_ ;
	wire _w2009_ ;
	wire _w2010_ ;
	wire _w2011_ ;
	wire _w2012_ ;
	wire _w2013_ ;
	wire _w2014_ ;
	wire _w2015_ ;
	wire _w2016_ ;
	wire _w2017_ ;
	wire _w2018_ ;
	wire _w2019_ ;
	wire _w2020_ ;
	wire _w2021_ ;
	wire _w2022_ ;
	wire _w2023_ ;
	wire _w2024_ ;
	wire _w2025_ ;
	wire _w2026_ ;
	wire _w2027_ ;
	wire _w2028_ ;
	wire _w2029_ ;
	wire _w2030_ ;
	wire _w2031_ ;
	wire _w2032_ ;
	wire _w2033_ ;
	wire _w2034_ ;
	wire _w2035_ ;
	wire _w2036_ ;
	wire _w2037_ ;
	wire _w2038_ ;
	wire _w2039_ ;
	wire _w2040_ ;
	wire _w2041_ ;
	wire _w2042_ ;
	wire _w2043_ ;
	wire _w2044_ ;
	wire _w2045_ ;
	wire _w2046_ ;
	wire _w2047_ ;
	wire _w2048_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3369_ ;
	wire _w3370_ ;
	wire _w3371_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3483_ ;
	wire _w3484_ ;
	wire _w3485_ ;
	wire _w3486_ ;
	wire _w3487_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3490_ ;
	wire _w3491_ ;
	wire _w3492_ ;
	wire _w3493_ ;
	wire _w3494_ ;
	wire _w3495_ ;
	wire _w3496_ ;
	wire _w3497_ ;
	wire _w3498_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	wire _w3538_ ;
	wire _w3539_ ;
	wire _w3540_ ;
	wire _w3541_ ;
	wire _w3542_ ;
	wire _w3543_ ;
	wire _w3544_ ;
	wire _w3545_ ;
	wire _w3546_ ;
	wire _w3547_ ;
	wire _w3548_ ;
	wire _w3549_ ;
	wire _w3550_ ;
	wire _w3551_ ;
	wire _w3552_ ;
	wire _w3553_ ;
	wire _w3554_ ;
	wire _w3555_ ;
	wire _w3556_ ;
	wire _w3557_ ;
	wire _w3558_ ;
	wire _w3559_ ;
	wire _w3560_ ;
	wire _w3561_ ;
	wire _w3562_ ;
	wire _w3563_ ;
	wire _w3564_ ;
	wire _w3565_ ;
	wire _w3566_ ;
	wire _w3567_ ;
	wire _w3568_ ;
	wire _w3569_ ;
	wire _w3570_ ;
	wire _w3571_ ;
	wire _w3572_ ;
	wire _w3573_ ;
	wire _w3574_ ;
	wire _w3575_ ;
	wire _w3576_ ;
	wire _w3577_ ;
	wire _w3578_ ;
	wire _w3579_ ;
	wire _w3580_ ;
	wire _w3581_ ;
	wire _w3582_ ;
	wire _w3583_ ;
	wire _w3584_ ;
	wire _w3585_ ;
	wire _w3586_ ;
	wire _w3587_ ;
	wire _w3588_ ;
	wire _w3589_ ;
	wire _w3590_ ;
	wire _w3591_ ;
	wire _w3592_ ;
	wire _w3593_ ;
	wire _w3594_ ;
	wire _w3595_ ;
	wire _w3596_ ;
	wire _w3597_ ;
	wire _w3598_ ;
	wire _w3599_ ;
	wire _w3600_ ;
	wire _w3601_ ;
	wire _w3602_ ;
	wire _w3603_ ;
	wire _w3604_ ;
	wire _w3605_ ;
	wire _w3606_ ;
	wire _w3607_ ;
	wire _w3608_ ;
	wire _w3609_ ;
	wire _w3610_ ;
	wire _w3611_ ;
	wire _w3612_ ;
	wire _w3613_ ;
	wire _w3614_ ;
	wire _w3615_ ;
	wire _w3616_ ;
	wire _w3617_ ;
	wire _w3618_ ;
	wire _w3619_ ;
	wire _w3620_ ;
	wire _w3621_ ;
	wire _w3622_ ;
	wire _w3623_ ;
	wire _w3624_ ;
	wire _w3625_ ;
	wire _w3626_ ;
	wire _w3627_ ;
	wire _w3628_ ;
	wire _w3629_ ;
	wire _w3630_ ;
	wire _w3631_ ;
	wire _w3632_ ;
	wire _w3633_ ;
	wire _w3634_ ;
	wire _w3635_ ;
	wire _w3636_ ;
	wire _w3637_ ;
	wire _w3638_ ;
	wire _w3639_ ;
	wire _w3640_ ;
	wire _w3641_ ;
	wire _w3642_ ;
	wire _w3643_ ;
	wire _w3644_ ;
	wire _w3645_ ;
	wire _w3646_ ;
	wire _w3647_ ;
	wire _w3648_ ;
	wire _w3649_ ;
	wire _w3650_ ;
	wire _w3651_ ;
	wire _w3652_ ;
	wire _w3653_ ;
	wire _w3654_ ;
	wire _w3655_ ;
	wire _w3656_ ;
	wire _w3657_ ;
	wire _w3658_ ;
	wire _w3659_ ;
	wire _w3660_ ;
	wire _w3661_ ;
	wire _w3662_ ;
	wire _w3663_ ;
	wire _w3664_ ;
	wire _w3665_ ;
	wire _w3666_ ;
	wire _w3667_ ;
	wire _w3668_ ;
	wire _w3669_ ;
	wire _w3670_ ;
	wire _w3671_ ;
	wire _w3672_ ;
	wire _w3673_ ;
	wire _w3674_ ;
	wire _w3675_ ;
	wire _w3676_ ;
	wire _w3677_ ;
	wire _w3678_ ;
	wire _w3679_ ;
	wire _w3680_ ;
	wire _w3681_ ;
	wire _w3682_ ;
	wire _w3683_ ;
	wire _w3684_ ;
	wire _w3685_ ;
	wire _w3686_ ;
	wire _w3687_ ;
	wire _w3688_ ;
	wire _w3689_ ;
	wire _w3690_ ;
	wire _w3691_ ;
	wire _w3692_ ;
	wire _w3693_ ;
	wire _w3694_ ;
	wire _w3695_ ;
	wire _w3696_ ;
	wire _w3697_ ;
	wire _w3698_ ;
	wire _w3699_ ;
	wire _w3700_ ;
	wire _w3701_ ;
	wire _w3702_ ;
	wire _w3703_ ;
	wire _w3704_ ;
	wire _w3705_ ;
	wire _w3706_ ;
	wire _w3707_ ;
	wire _w3708_ ;
	wire _w3709_ ;
	wire _w3710_ ;
	wire _w3711_ ;
	wire _w3712_ ;
	wire _w3713_ ;
	wire _w3714_ ;
	wire _w3715_ ;
	wire _w3716_ ;
	wire _w3717_ ;
	wire _w3718_ ;
	wire _w3719_ ;
	wire _w3720_ ;
	wire _w3721_ ;
	wire _w3722_ ;
	wire _w3723_ ;
	wire _w3724_ ;
	wire _w3725_ ;
	wire _w3726_ ;
	wire _w3727_ ;
	wire _w3728_ ;
	wire _w3729_ ;
	wire _w3730_ ;
	wire _w3731_ ;
	wire _w3732_ ;
	wire _w3733_ ;
	wire _w3734_ ;
	wire _w3735_ ;
	wire _w3736_ ;
	wire _w3737_ ;
	wire _w3738_ ;
	wire _w3739_ ;
	wire _w3740_ ;
	wire _w3741_ ;
	wire _w3742_ ;
	wire _w3743_ ;
	wire _w3744_ ;
	wire _w3745_ ;
	wire _w3746_ ;
	wire _w3747_ ;
	wire _w3748_ ;
	wire _w3749_ ;
	wire _w3750_ ;
	wire _w3751_ ;
	wire _w3752_ ;
	wire _w3753_ ;
	wire _w3754_ ;
	wire _w3755_ ;
	wire _w3756_ ;
	wire _w3757_ ;
	wire _w3758_ ;
	wire _w3759_ ;
	wire _w3760_ ;
	wire _w3761_ ;
	wire _w3762_ ;
	wire _w3763_ ;
	wire _w3764_ ;
	wire _w3765_ ;
	wire _w3766_ ;
	wire _w3767_ ;
	wire _w3768_ ;
	wire _w3769_ ;
	wire _w3770_ ;
	wire _w3771_ ;
	wire _w3772_ ;
	wire _w3773_ ;
	wire _w3774_ ;
	wire _w3775_ ;
	wire _w3776_ ;
	wire _w3777_ ;
	wire _w3778_ ;
	wire _w3779_ ;
	wire _w3780_ ;
	wire _w3781_ ;
	wire _w3782_ ;
	wire _w3783_ ;
	wire _w3784_ ;
	wire _w3785_ ;
	wire _w3786_ ;
	wire _w3787_ ;
	wire _w3788_ ;
	wire _w3789_ ;
	wire _w3790_ ;
	wire _w3791_ ;
	wire _w3792_ ;
	wire _w3793_ ;
	wire _w3794_ ;
	wire _w3795_ ;
	wire _w3796_ ;
	wire _w3797_ ;
	wire _w3798_ ;
	wire _w3799_ ;
	wire _w3800_ ;
	wire _w3801_ ;
	wire _w3802_ ;
	wire _w3803_ ;
	wire _w3804_ ;
	wire _w3805_ ;
	wire _w3806_ ;
	wire _w3807_ ;
	wire _w3808_ ;
	wire _w3809_ ;
	wire _w3810_ ;
	wire _w3811_ ;
	wire _w3812_ ;
	wire _w3813_ ;
	wire _w3814_ ;
	wire _w3815_ ;
	wire _w3816_ ;
	wire _w3817_ ;
	wire _w3818_ ;
	wire _w3819_ ;
	wire _w3820_ ;
	wire _w3821_ ;
	wire _w3822_ ;
	wire _w3823_ ;
	wire _w3824_ ;
	wire _w3825_ ;
	wire _w3826_ ;
	wire _w3827_ ;
	wire _w3828_ ;
	wire _w3829_ ;
	wire _w3830_ ;
	wire _w3831_ ;
	wire _w3832_ ;
	wire _w3833_ ;
	wire _w3834_ ;
	wire _w3835_ ;
	wire _w3836_ ;
	wire _w3837_ ;
	wire _w3838_ ;
	wire _w3839_ ;
	wire _w3840_ ;
	wire _w3841_ ;
	wire _w3842_ ;
	wire _w3843_ ;
	wire _w3844_ ;
	wire _w3845_ ;
	wire _w3846_ ;
	wire _w3847_ ;
	wire _w3848_ ;
	wire _w3849_ ;
	wire _w3850_ ;
	wire _w3851_ ;
	wire _w3852_ ;
	wire _w3853_ ;
	wire _w3854_ ;
	wire _w3855_ ;
	wire _w3856_ ;
	wire _w3857_ ;
	wire _w3858_ ;
	wire _w3859_ ;
	wire _w3860_ ;
	wire _w3861_ ;
	wire _w3862_ ;
	wire _w3863_ ;
	wire _w3864_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\A[67] ,
		\A[68] ,
		_w1002_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\A[67] ,
		\A[68] ,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		\A[69] ,
		_w1004_,
		_w1005_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		_w1002_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\A[70] ,
		\A[71] ,
		_w1007_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		\A[69] ,
		_w1004_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name7 (
		_w1005_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		\A[70] ,
		\A[71] ,
		_w1010_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w1007_,
		_w1010_,
		_w1011_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\A[72] ,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		\A[72] ,
		_w1011_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w1012_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w1009_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		_w1007_,
		_w1015_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name15 (
		_w1007_,
		_w1012_,
		_w1017_
	);
	LUT2 #(
		.INIT('h4)
	) name16 (
		_w1015_,
		_w1017_,
		_w1018_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		_w1016_,
		_w1018_,
		_w1019_
	);
	LUT2 #(
		.INIT('h2)
	) name18 (
		_w1006_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w1006_,
		_w1019_,
		_w1021_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w1020_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\A[73] ,
		\A[74] ,
		_w1023_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		\A[73] ,
		\A[74] ,
		_w1024_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		_w1023_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		\A[75] ,
		_w1025_,
		_w1026_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\A[75] ,
		_w1025_,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w1026_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\A[76] ,
		\A[77] ,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		\A[76] ,
		\A[77] ,
		_w1030_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w1029_,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\A[78] ,
		_w1031_,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\A[78] ,
		_w1031_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w1032_,
		_w1033_,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w1028_,
		_w1034_,
		_w1035_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w1029_,
		_w1032_,
		_w1036_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w1023_,
		_w1026_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w1036_,
		_w1037_,
		_w1039_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w1038_,
		_w1039_,
		_w1040_
	);
	LUT2 #(
		.INIT('h4)
	) name39 (
		_w1035_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w1009_,
		_w1014_,
		_w1042_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		_w1015_,
		_w1042_,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w1028_,
		_w1034_,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w1035_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		_w1043_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h2)
	) name45 (
		_w1035_,
		_w1040_,
		_w1047_
	);
	LUT2 #(
		.INIT('h1)
	) name46 (
		_w1041_,
		_w1046_,
		_w1048_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('h2)
	) name48 (
		_w1022_,
		_w1049_,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w1040_,
		_w1046_,
		_w1051_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w1006_,
		_w1016_,
		_w1052_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		_w1051_,
		_w1052_,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w1050_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h4)
	) name53 (
		_w1029_,
		_w1037_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		_w1035_,
		_w1055_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w1038_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w1054_,
		_w1057_,
		_w1058_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		_w1006_,
		_w1018_,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w1016_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w1054_,
		_w1057_,
		_w1061_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w1060_,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w1058_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		\A[61] ,
		\A[62] ,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		\A[61] ,
		\A[62] ,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w1064_,
		_w1065_,
		_w1066_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		\A[63] ,
		_w1066_,
		_w1067_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\A[63] ,
		_w1066_,
		_w1068_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w1067_,
		_w1068_,
		_w1069_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\A[64] ,
		\A[65] ,
		_w1070_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		\A[64] ,
		\A[65] ,
		_w1071_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w1070_,
		_w1071_,
		_w1072_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		\A[66] ,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		\A[66] ,
		_w1072_,
		_w1074_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w1073_,
		_w1074_,
		_w1075_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		_w1069_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w1069_,
		_w1075_,
		_w1077_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w1076_,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\A[55] ,
		\A[56] ,
		_w1079_
	);
	LUT2 #(
		.INIT('h1)
	) name78 (
		\A[55] ,
		\A[56] ,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w1079_,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		\A[57] ,
		_w1081_,
		_w1082_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\A[57] ,
		_w1081_,
		_w1083_
	);
	LUT2 #(
		.INIT('h1)
	) name82 (
		_w1082_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\A[58] ,
		\A[59] ,
		_w1085_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		\A[58] ,
		\A[59] ,
		_w1086_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w1085_,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		\A[60] ,
		_w1087_,
		_w1088_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\A[60] ,
		_w1087_,
		_w1089_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w1088_,
		_w1089_,
		_w1090_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		_w1084_,
		_w1090_,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w1084_,
		_w1090_,
		_w1092_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w1091_,
		_w1092_,
		_w1093_
	);
	LUT2 #(
		.INIT('h8)
	) name92 (
		_w1078_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w1064_,
		_w1067_,
		_w1095_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w1070_,
		_w1073_,
		_w1096_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w1076_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h8)
	) name96 (
		_w1070_,
		_w1076_,
		_w1098_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		_w1097_,
		_w1098_,
		_w1099_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		_w1095_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w1095_,
		_w1099_,
		_w1101_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w1100_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w1094_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		_w1079_,
		_w1082_,
		_w1104_
	);
	LUT2 #(
		.INIT('h8)
	) name103 (
		_w1085_,
		_w1091_,
		_w1105_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w1085_,
		_w1088_,
		_w1106_
	);
	LUT2 #(
		.INIT('h4)
	) name105 (
		_w1091_,
		_w1106_,
		_w1107_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w1105_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		_w1104_,
		_w1108_,
		_w1109_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		_w1104_,
		_w1108_,
		_w1110_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w1109_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w1103_,
		_w1111_,
		_w1112_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w1094_,
		_w1102_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w1095_,
		_w1096_,
		_w1114_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w1104_,
		_w1105_,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		_w1114_,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		_w1113_,
		_w1116_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w1112_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w1095_,
		_w1097_,
		_w1119_
	);
	LUT2 #(
		.INIT('h1)
	) name118 (
		_w1098_,
		_w1119_,
		_w1120_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w1118_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w1104_,
		_w1107_,
		_w1122_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w1105_,
		_w1122_,
		_w1123_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		_w1118_,
		_w1120_,
		_w1124_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w1123_,
		_w1124_,
		_w1125_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w1121_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h8)
	) name125 (
		_w1063_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h1)
	) name126 (
		_w1063_,
		_w1126_,
		_w1128_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w1121_,
		_w1124_,
		_w1129_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		_w1123_,
		_w1129_,
		_w1130_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w1123_,
		_w1129_,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		_w1130_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w1058_,
		_w1061_,
		_w1133_
	);
	LUT2 #(
		.INIT('h2)
	) name132 (
		_w1060_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		_w1060_,
		_w1133_,
		_w1135_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w1134_,
		_w1135_,
		_w1136_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w1132_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w1043_,
		_w1045_,
		_w1138_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w1046_,
		_w1138_,
		_w1139_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w1078_,
		_w1093_,
		_w1140_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w1094_,
		_w1140_,
		_w1141_
	);
	LUT2 #(
		.INIT('h8)
	) name140 (
		_w1139_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		_w1050_,
		_w1053_,
		_w1143_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		_w1049_,
		_w1051_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w1022_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w1143_,
		_w1145_,
		_w1146_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		_w1142_,
		_w1146_,
		_w1147_
	);
	LUT2 #(
		.INIT('h2)
	) name146 (
		_w1112_,
		_w1117_,
		_w1148_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w1103_,
		_w1113_,
		_w1149_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w1111_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w1148_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w1142_,
		_w1146_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w1151_,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w1147_,
		_w1153_,
		_w1154_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w1132_,
		_w1136_,
		_w1155_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w1154_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w1137_,
		_w1156_,
		_w1157_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w1128_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w1127_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		\A[43] ,
		\A[44] ,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		\A[43] ,
		\A[44] ,
		_w1161_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w1160_,
		_w1161_,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\A[45] ,
		_w1162_,
		_w1163_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w1160_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\A[46] ,
		\A[47] ,
		_w1165_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		\A[45] ,
		_w1162_,
		_w1166_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w1163_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		\A[46] ,
		\A[47] ,
		_w1168_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		_w1165_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\A[48] ,
		_w1169_,
		_w1170_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		\A[48] ,
		_w1169_,
		_w1171_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w1170_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w1167_,
		_w1172_,
		_w1173_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		_w1165_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w1165_,
		_w1170_,
		_w1175_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		_w1173_,
		_w1175_,
		_w1176_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		_w1174_,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		_w1164_,
		_w1177_,
		_w1178_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		_w1164_,
		_w1177_,
		_w1179_
	);
	LUT2 #(
		.INIT('h1)
	) name178 (
		_w1178_,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		\A[49] ,
		\A[50] ,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		\A[49] ,
		\A[50] ,
		_w1182_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w1181_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\A[51] ,
		_w1183_,
		_w1184_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		\A[51] ,
		_w1183_,
		_w1185_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w1184_,
		_w1185_,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name185 (
		\A[52] ,
		\A[53] ,
		_w1187_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		\A[52] ,
		\A[53] ,
		_w1188_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w1187_,
		_w1188_,
		_w1189_
	);
	LUT2 #(
		.INIT('h8)
	) name188 (
		\A[54] ,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		\A[54] ,
		_w1189_,
		_w1191_
	);
	LUT2 #(
		.INIT('h1)
	) name190 (
		_w1190_,
		_w1191_,
		_w1192_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w1186_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w1187_,
		_w1190_,
		_w1194_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w1181_,
		_w1184_,
		_w1195_
	);
	LUT2 #(
		.INIT('h1)
	) name194 (
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w1194_,
		_w1195_,
		_w1197_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w1196_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		_w1193_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w1167_,
		_w1172_,
		_w1200_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w1173_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w1186_,
		_w1192_,
		_w1202_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w1193_,
		_w1202_,
		_w1203_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		_w1201_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		_w1193_,
		_w1198_,
		_w1205_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w1199_,
		_w1204_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w1205_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		_w1180_,
		_w1207_,
		_w1208_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		_w1198_,
		_w1204_,
		_w1209_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w1164_,
		_w1174_,
		_w1210_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		_w1209_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w1208_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		_w1187_,
		_w1195_,
		_w1213_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		_w1193_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w1196_,
		_w1214_,
		_w1215_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w1212_,
		_w1215_,
		_w1216_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w1164_,
		_w1176_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w1174_,
		_w1217_,
		_w1218_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		_w1212_,
		_w1215_,
		_w1219_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w1218_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w1216_,
		_w1220_,
		_w1221_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\A[37] ,
		\A[38] ,
		_w1222_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		\A[37] ,
		\A[38] ,
		_w1223_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w1222_,
		_w1223_,
		_w1224_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\A[39] ,
		_w1224_,
		_w1225_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		\A[39] ,
		_w1224_,
		_w1226_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w1225_,
		_w1226_,
		_w1227_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\A[40] ,
		\A[41] ,
		_w1228_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		\A[40] ,
		\A[41] ,
		_w1229_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w1228_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		\A[42] ,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		\A[42] ,
		_w1230_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		_w1227_,
		_w1233_,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		_w1227_,
		_w1233_,
		_w1235_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w1234_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\A[31] ,
		\A[32] ,
		_w1237_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		\A[31] ,
		\A[32] ,
		_w1238_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w1237_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\A[33] ,
		_w1239_,
		_w1240_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		\A[33] ,
		_w1239_,
		_w1241_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w1240_,
		_w1241_,
		_w1242_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		\A[34] ,
		\A[35] ,
		_w1243_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		\A[34] ,
		\A[35] ,
		_w1244_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w1243_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		\A[36] ,
		_w1245_,
		_w1246_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\A[36] ,
		_w1245_,
		_w1247_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w1246_,
		_w1247_,
		_w1248_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w1242_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w1242_,
		_w1248_,
		_w1250_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		_w1249_,
		_w1250_,
		_w1251_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		_w1236_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w1228_,
		_w1231_,
		_w1253_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w1222_,
		_w1225_,
		_w1254_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w1253_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		_w1253_,
		_w1254_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w1255_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		_w1252_,
		_w1257_,
		_w1258_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w1243_,
		_w1246_,
		_w1259_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w1237_,
		_w1240_,
		_w1260_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w1259_,
		_w1260_,
		_w1261_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		_w1259_,
		_w1260_,
		_w1262_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w1261_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name262 (
		_w1249_,
		_w1263_,
		_w1264_
	);
	LUT2 #(
		.INIT('h4)
	) name263 (
		_w1249_,
		_w1263_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w1264_,
		_w1265_,
		_w1266_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		_w1258_,
		_w1266_,
		_w1267_
	);
	LUT2 #(
		.INIT('h4)
	) name266 (
		_w1234_,
		_w1257_,
		_w1268_
	);
	LUT2 #(
		.INIT('h2)
	) name267 (
		_w1234_,
		_w1257_,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w1252_,
		_w1268_,
		_w1270_
	);
	LUT2 #(
		.INIT('h4)
	) name269 (
		_w1269_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w1267_,
		_w1271_,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w1234_,
		_w1255_,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w1256_,
		_w1273_,
		_w1274_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w1272_,
		_w1274_,
		_w1275_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w1272_,
		_w1274_,
		_w1276_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w1249_,
		_w1261_,
		_w1277_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w1262_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w1276_,
		_w1278_,
		_w1279_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w1275_,
		_w1279_,
		_w1280_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		_w1221_,
		_w1280_,
		_w1281_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		_w1221_,
		_w1280_,
		_w1282_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		_w1216_,
		_w1219_,
		_w1283_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		_w1218_,
		_w1283_,
		_w1284_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w1218_,
		_w1283_,
		_w1285_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w1284_,
		_w1285_,
		_w1286_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w1275_,
		_w1276_,
		_w1287_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w1278_,
		_w1287_,
		_w1288_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		_w1278_,
		_w1287_,
		_w1289_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w1288_,
		_w1289_,
		_w1290_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		_w1286_,
		_w1290_,
		_w1291_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		_w1286_,
		_w1290_,
		_w1292_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w1201_,
		_w1203_,
		_w1293_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w1204_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w1236_,
		_w1251_,
		_w1295_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w1252_,
		_w1295_,
		_w1296_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		_w1294_,
		_w1296_,
		_w1297_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		_w1208_,
		_w1211_,
		_w1298_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		_w1207_,
		_w1209_,
		_w1299_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w1180_,
		_w1299_,
		_w1300_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w1298_,
		_w1300_,
		_w1301_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		_w1297_,
		_w1301_,
		_w1302_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w1297_,
		_w1301_,
		_w1303_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w1258_,
		_w1271_,
		_w1304_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		_w1266_,
		_w1304_,
		_w1305_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w1266_,
		_w1304_,
		_w1306_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT2 #(
		.INIT('h1)
	) name306 (
		_w1303_,
		_w1307_,
		_w1308_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w1302_,
		_w1308_,
		_w1309_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w1292_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w1291_,
		_w1310_,
		_w1311_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w1282_,
		_w1311_,
		_w1312_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w1281_,
		_w1312_,
		_w1313_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		_w1159_,
		_w1313_,
		_w1314_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		_w1159_,
		_w1313_,
		_w1315_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w1127_,
		_w1128_,
		_w1316_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		_w1157_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		_w1157_,
		_w1316_,
		_w1318_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w1317_,
		_w1318_,
		_w1319_
	);
	LUT2 #(
		.INIT('h1)
	) name318 (
		_w1281_,
		_w1282_,
		_w1320_
	);
	LUT2 #(
		.INIT('h4)
	) name319 (
		_w1311_,
		_w1320_,
		_w1321_
	);
	LUT2 #(
		.INIT('h2)
	) name320 (
		_w1311_,
		_w1320_,
		_w1322_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w1321_,
		_w1322_,
		_w1323_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		_w1319_,
		_w1323_,
		_w1324_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		_w1319_,
		_w1323_,
		_w1325_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w1137_,
		_w1155_,
		_w1326_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w1154_,
		_w1326_,
		_w1327_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w1154_,
		_w1326_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w1327_,
		_w1328_,
		_w1329_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		_w1291_,
		_w1292_,
		_w1330_
	);
	LUT2 #(
		.INIT('h4)
	) name329 (
		_w1309_,
		_w1330_,
		_w1331_
	);
	LUT2 #(
		.INIT('h2)
	) name330 (
		_w1309_,
		_w1330_,
		_w1332_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w1331_,
		_w1332_,
		_w1333_
	);
	LUT2 #(
		.INIT('h8)
	) name332 (
		_w1329_,
		_w1333_,
		_w1334_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w1329_,
		_w1333_,
		_w1335_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w1139_,
		_w1141_,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w1142_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w1294_,
		_w1296_,
		_w1338_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w1297_,
		_w1338_,
		_w1339_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w1337_,
		_w1339_,
		_w1340_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w1147_,
		_w1152_,
		_w1341_
	);
	LUT2 #(
		.INIT('h2)
	) name340 (
		_w1151_,
		_w1341_,
		_w1342_
	);
	LUT2 #(
		.INIT('h4)
	) name341 (
		_w1151_,
		_w1341_,
		_w1343_
	);
	LUT2 #(
		.INIT('h1)
	) name342 (
		_w1342_,
		_w1343_,
		_w1344_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		_w1340_,
		_w1344_,
		_w1345_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		_w1340_,
		_w1344_,
		_w1346_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		_w1302_,
		_w1303_,
		_w1347_
	);
	LUT2 #(
		.INIT('h4)
	) name346 (
		_w1307_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h2)
	) name347 (
		_w1307_,
		_w1347_,
		_w1349_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w1348_,
		_w1349_,
		_w1350_
	);
	LUT2 #(
		.INIT('h4)
	) name349 (
		_w1346_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w1345_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h1)
	) name351 (
		_w1335_,
		_w1352_,
		_w1353_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		_w1334_,
		_w1353_,
		_w1354_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		_w1325_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h1)
	) name354 (
		_w1324_,
		_w1355_,
		_w1356_
	);
	LUT2 #(
		.INIT('h4)
	) name355 (
		_w1315_,
		_w1356_,
		_w1357_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w1314_,
		_w1357_,
		_w1358_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		\A[3] ,
		\A[4] ,
		_w1359_
	);
	LUT2 #(
		.INIT('h1)
	) name358 (
		\A[3] ,
		\A[4] ,
		_w1360_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w1359_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		\A[5] ,
		_w1361_,
		_w1362_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		_w1359_,
		_w1362_,
		_w1363_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		\A[0] ,
		\A[1] ,
		_w1364_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		\A[0] ,
		\A[1] ,
		_w1365_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w1364_,
		_w1365_,
		_w1366_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		\A[2] ,
		_w1366_,
		_w1367_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w1364_,
		_w1367_,
		_w1368_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w1363_,
		_w1368_,
		_w1369_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		\A[2] ,
		_w1366_,
		_w1370_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w1367_,
		_w1370_,
		_w1371_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		\A[6] ,
		_w1371_,
		_w1372_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		\A[6] ,
		_w1371_,
		_w1373_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w1372_,
		_w1373_,
		_w1374_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		\A[5] ,
		_w1361_,
		_w1375_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w1362_,
		_w1375_,
		_w1376_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w1374_,
		_w1376_,
		_w1377_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w1372_,
		_w1377_,
		_w1378_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		_w1363_,
		_w1368_,
		_w1379_
	);
	LUT2 #(
		.INIT('h1)
	) name378 (
		_w1369_,
		_w1379_,
		_w1380_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		_w1378_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w1369_,
		_w1381_,
		_w1382_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w1374_,
		_w1376_,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w1377_,
		_w1383_,
		_w1384_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		\A[997] ,
		\A[998] ,
		_w1385_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		\A[997] ,
		\A[998] ,
		_w1386_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w1385_,
		_w1386_,
		_w1387_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		\A[999] ,
		_w1387_,
		_w1388_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		\A[999] ,
		_w1387_,
		_w1389_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w1388_,
		_w1389_,
		_w1390_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		_w1384_,
		_w1390_,
		_w1391_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		_w1378_,
		_w1380_,
		_w1392_
	);
	LUT2 #(
		.INIT('h1)
	) name391 (
		_w1381_,
		_w1392_,
		_w1393_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w1391_,
		_w1393_,
		_w1394_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		_w1385_,
		_w1388_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		_w1391_,
		_w1393_,
		_w1396_
	);
	LUT2 #(
		.INIT('h2)
	) name395 (
		_w1395_,
		_w1396_,
		_w1397_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w1394_,
		_w1397_,
		_w1398_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w1382_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w1384_,
		_w1390_,
		_w1400_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w1391_,
		_w1400_,
		_w1401_
	);
	LUT2 #(
		.INIT('h8)
	) name400 (
		\A[991] ,
		\A[992] ,
		_w1402_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		\A[991] ,
		\A[992] ,
		_w1403_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w1402_,
		_w1403_,
		_w1404_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		\A[993] ,
		_w1404_,
		_w1405_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		\A[993] ,
		_w1404_,
		_w1406_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w1405_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		\A[994] ,
		\A[995] ,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		\A[994] ,
		\A[995] ,
		_w1409_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w1408_,
		_w1409_,
		_w1410_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		\A[996] ,
		_w1410_,
		_w1411_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		\A[996] ,
		_w1410_,
		_w1412_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w1411_,
		_w1412_,
		_w1413_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		_w1407_,
		_w1413_,
		_w1414_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w1407_,
		_w1413_,
		_w1415_
	);
	LUT2 #(
		.INIT('h1)
	) name414 (
		_w1414_,
		_w1415_,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		_w1401_,
		_w1416_,
		_w1417_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w1394_,
		_w1396_,
		_w1418_
	);
	LUT2 #(
		.INIT('h2)
	) name417 (
		_w1395_,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h4)
	) name418 (
		_w1395_,
		_w1418_,
		_w1420_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w1419_,
		_w1420_,
		_w1421_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w1417_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		_w1417_,
		_w1421_,
		_w1423_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w1408_,
		_w1411_,
		_w1424_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w1402_,
		_w1405_,
		_w1425_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w1424_,
		_w1425_,
		_w1426_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		_w1424_,
		_w1425_,
		_w1427_
	);
	LUT2 #(
		.INIT('h1)
	) name426 (
		_w1426_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h2)
	) name427 (
		_w1414_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h4)
	) name428 (
		_w1414_,
		_w1428_,
		_w1430_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w1429_,
		_w1430_,
		_w1431_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		_w1423_,
		_w1431_,
		_w1432_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w1422_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w1414_,
		_w1426_,
		_w1434_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w1427_,
		_w1434_,
		_w1435_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w1433_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		_w1399_,
		_w1436_,
		_w1437_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		\A[19] ,
		\A[20] ,
		_w1438_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		\A[19] ,
		\A[20] ,
		_w1439_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w1438_,
		_w1439_,
		_w1440_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		\A[21] ,
		_w1440_,
		_w1441_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		\A[21] ,
		_w1440_,
		_w1442_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w1441_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		\A[22] ,
		\A[23] ,
		_w1444_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		\A[22] ,
		\A[23] ,
		_w1445_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w1444_,
		_w1445_,
		_w1446_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		\A[24] ,
		_w1446_,
		_w1447_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		\A[24] ,
		_w1446_,
		_w1448_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w1447_,
		_w1448_,
		_w1449_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w1443_,
		_w1449_,
		_w1450_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w1443_,
		_w1449_,
		_w1451_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w1450_,
		_w1451_,
		_w1452_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		\A[25] ,
		\A[26] ,
		_w1453_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		\A[25] ,
		\A[26] ,
		_w1454_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		_w1453_,
		_w1454_,
		_w1455_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\A[27] ,
		_w1455_,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		\A[27] ,
		_w1455_,
		_w1457_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		_w1456_,
		_w1457_,
		_w1458_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		\A[28] ,
		\A[29] ,
		_w1459_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		\A[28] ,
		\A[29] ,
		_w1460_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w1459_,
		_w1460_,
		_w1461_
	);
	LUT2 #(
		.INIT('h8)
	) name460 (
		\A[30] ,
		_w1461_,
		_w1462_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		\A[30] ,
		_w1461_,
		_w1463_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w1462_,
		_w1463_,
		_w1464_
	);
	LUT2 #(
		.INIT('h8)
	) name463 (
		_w1458_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w1458_,
		_w1464_,
		_w1466_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w1465_,
		_w1466_,
		_w1467_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		_w1452_,
		_w1467_,
		_w1468_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w1459_,
		_w1462_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w1453_,
		_w1456_,
		_w1470_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		_w1469_,
		_w1470_,
		_w1471_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w1469_,
		_w1470_,
		_w1472_
	);
	LUT2 #(
		.INIT('h1)
	) name471 (
		_w1471_,
		_w1472_,
		_w1473_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		_w1468_,
		_w1473_,
		_w1474_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		_w1444_,
		_w1447_,
		_w1475_
	);
	LUT2 #(
		.INIT('h1)
	) name474 (
		_w1438_,
		_w1441_,
		_w1476_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w1475_,
		_w1476_,
		_w1477_
	);
	LUT2 #(
		.INIT('h8)
	) name476 (
		_w1475_,
		_w1476_,
		_w1478_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w1477_,
		_w1478_,
		_w1479_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		_w1450_,
		_w1479_,
		_w1480_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		_w1450_,
		_w1479_,
		_w1481_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		_w1480_,
		_w1481_,
		_w1482_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		_w1474_,
		_w1482_,
		_w1483_
	);
	LUT2 #(
		.INIT('h4)
	) name482 (
		_w1465_,
		_w1473_,
		_w1484_
	);
	LUT2 #(
		.INIT('h2)
	) name483 (
		_w1465_,
		_w1473_,
		_w1485_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w1468_,
		_w1484_,
		_w1486_
	);
	LUT2 #(
		.INIT('h4)
	) name485 (
		_w1485_,
		_w1486_,
		_w1487_
	);
	LUT2 #(
		.INIT('h1)
	) name486 (
		_w1483_,
		_w1487_,
		_w1488_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		_w1465_,
		_w1471_,
		_w1489_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w1472_,
		_w1489_,
		_w1490_
	);
	LUT2 #(
		.INIT('h4)
	) name489 (
		_w1488_,
		_w1490_,
		_w1491_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		_w1488_,
		_w1490_,
		_w1492_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w1450_,
		_w1477_,
		_w1493_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w1478_,
		_w1493_,
		_w1494_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w1492_,
		_w1494_,
		_w1495_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w1491_,
		_w1495_,
		_w1496_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		\A[7] ,
		\A[8] ,
		_w1497_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		\A[7] ,
		\A[8] ,
		_w1498_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w1497_,
		_w1498_,
		_w1499_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\A[9] ,
		_w1499_,
		_w1500_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		\A[9] ,
		_w1499_,
		_w1501_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		\A[10] ,
		\A[11] ,
		_w1503_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		\A[10] ,
		\A[11] ,
		_w1504_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w1503_,
		_w1504_,
		_w1505_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		\A[12] ,
		_w1505_,
		_w1506_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		\A[12] ,
		_w1505_,
		_w1507_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w1506_,
		_w1507_,
		_w1508_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		_w1502_,
		_w1508_,
		_w1509_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w1502_,
		_w1508_,
		_w1510_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\A[13] ,
		\A[14] ,
		_w1512_
	);
	LUT2 #(
		.INIT('h1)
	) name511 (
		\A[13] ,
		\A[14] ,
		_w1513_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w1512_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		\A[15] ,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		\A[15] ,
		_w1514_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w1515_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		\A[16] ,
		\A[17] ,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		\A[16] ,
		\A[17] ,
		_w1519_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		\A[18] ,
		_w1520_,
		_w1521_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		\A[18] ,
		_w1520_,
		_w1522_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w1517_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w1517_,
		_w1523_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w1524_,
		_w1525_,
		_w1526_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		_w1511_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		_w1518_,
		_w1521_,
		_w1528_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		_w1512_,
		_w1515_,
		_w1529_
	);
	LUT2 #(
		.INIT('h8)
	) name528 (
		_w1528_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w1528_,
		_w1529_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		_w1530_,
		_w1531_,
		_w1532_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		_w1527_,
		_w1532_,
		_w1533_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w1503_,
		_w1506_,
		_w1534_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w1497_,
		_w1500_,
		_w1535_
	);
	LUT2 #(
		.INIT('h1)
	) name534 (
		_w1534_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		_w1534_,
		_w1535_,
		_w1537_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w1536_,
		_w1537_,
		_w1538_
	);
	LUT2 #(
		.INIT('h2)
	) name537 (
		_w1509_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		_w1509_,
		_w1538_,
		_w1540_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h4)
	) name540 (
		_w1533_,
		_w1541_,
		_w1542_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w1524_,
		_w1532_,
		_w1543_
	);
	LUT2 #(
		.INIT('h2)
	) name542 (
		_w1524_,
		_w1532_,
		_w1544_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		_w1527_,
		_w1543_,
		_w1545_
	);
	LUT2 #(
		.INIT('h4)
	) name544 (
		_w1544_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		_w1542_,
		_w1546_,
		_w1547_
	);
	LUT2 #(
		.INIT('h2)
	) name546 (
		_w1524_,
		_w1530_,
		_w1548_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w1531_,
		_w1548_,
		_w1549_
	);
	LUT2 #(
		.INIT('h4)
	) name548 (
		_w1547_,
		_w1549_,
		_w1550_
	);
	LUT2 #(
		.INIT('h2)
	) name549 (
		_w1547_,
		_w1549_,
		_w1551_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w1509_,
		_w1536_,
		_w1552_
	);
	LUT2 #(
		.INIT('h1)
	) name551 (
		_w1537_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w1551_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		_w1550_,
		_w1554_,
		_w1555_
	);
	LUT2 #(
		.INIT('h8)
	) name554 (
		_w1496_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w1496_,
		_w1555_,
		_w1557_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w1550_,
		_w1551_,
		_w1558_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		_w1553_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h2)
	) name558 (
		_w1553_,
		_w1558_,
		_w1560_
	);
	LUT2 #(
		.INIT('h1)
	) name559 (
		_w1559_,
		_w1560_,
		_w1561_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w1491_,
		_w1492_,
		_w1562_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		_w1494_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h2)
	) name562 (
		_w1494_,
		_w1562_,
		_w1564_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		_w1563_,
		_w1564_,
		_w1565_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w1561_,
		_w1565_,
		_w1566_
	);
	LUT2 #(
		.INIT('h8)
	) name565 (
		_w1561_,
		_w1565_,
		_w1567_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		_w1452_,
		_w1467_,
		_w1568_
	);
	LUT2 #(
		.INIT('h1)
	) name567 (
		_w1468_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w1511_,
		_w1526_,
		_w1570_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		_w1527_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		_w1569_,
		_w1571_,
		_w1572_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w1474_,
		_w1487_,
		_w1573_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		_w1482_,
		_w1573_,
		_w1574_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w1482_,
		_w1573_,
		_w1575_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		_w1574_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		_w1572_,
		_w1576_,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name576 (
		_w1572_,
		_w1576_,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name577 (
		_w1533_,
		_w1546_,
		_w1579_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		_w1541_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w1541_,
		_w1579_,
		_w1581_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w1580_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w1578_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h1)
	) name582 (
		_w1577_,
		_w1583_,
		_w1584_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w1567_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w1566_,
		_w1585_,
		_w1586_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		_w1557_,
		_w1586_,
		_w1587_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w1556_,
		_w1587_,
		_w1588_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		_w1437_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h4)
	) name588 (
		_w1437_,
		_w1588_,
		_w1590_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w1399_,
		_w1436_,
		_w1591_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w1437_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h2)
	) name591 (
		_w1382_,
		_w1398_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w1399_,
		_w1593_,
		_w1594_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		_w1433_,
		_w1435_,
		_w1595_
	);
	LUT2 #(
		.INIT('h2)
	) name594 (
		_w1594_,
		_w1595_,
		_w1596_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		_w1592_,
		_w1596_,
		_w1597_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w1556_,
		_w1557_,
		_w1598_
	);
	LUT2 #(
		.INIT('h4)
	) name597 (
		_w1586_,
		_w1598_,
		_w1599_
	);
	LUT2 #(
		.INIT('h2)
	) name598 (
		_w1586_,
		_w1598_,
		_w1600_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		_w1597_,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h4)
	) name601 (
		_w1597_,
		_w1601_,
		_w1603_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		_w1435_,
		_w1594_,
		_w1604_
	);
	LUT2 #(
		.INIT('h2)
	) name603 (
		_w1435_,
		_w1594_,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w1604_,
		_w1605_,
		_w1606_
	);
	LUT2 #(
		.INIT('h8)
	) name605 (
		_w1433_,
		_w1606_,
		_w1607_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		_w1433_,
		_w1606_,
		_w1608_
	);
	LUT2 #(
		.INIT('h1)
	) name607 (
		_w1607_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w1566_,
		_w1567_,
		_w1610_
	);
	LUT2 #(
		.INIT('h4)
	) name609 (
		_w1584_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		_w1584_,
		_w1610_,
		_w1612_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w1611_,
		_w1612_,
		_w1613_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		_w1609_,
		_w1613_,
		_w1614_
	);
	LUT2 #(
		.INIT('h2)
	) name613 (
		_w1609_,
		_w1613_,
		_w1615_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		_w1569_,
		_w1571_,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name615 (
		_w1572_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		_w1401_,
		_w1416_,
		_w1618_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		_w1417_,
		_w1618_,
		_w1619_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		_w1617_,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w1577_,
		_w1578_,
		_w1621_
	);
	LUT2 #(
		.INIT('h4)
	) name620 (
		_w1582_,
		_w1621_,
		_w1622_
	);
	LUT2 #(
		.INIT('h2)
	) name621 (
		_w1582_,
		_w1621_,
		_w1623_
	);
	LUT2 #(
		.INIT('h1)
	) name622 (
		_w1622_,
		_w1623_,
		_w1624_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		_w1620_,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w1620_,
		_w1624_,
		_w1626_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		_w1422_,
		_w1423_,
		_w1627_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		_w1431_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		_w1431_,
		_w1627_,
		_w1629_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		_w1628_,
		_w1629_,
		_w1630_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w1626_,
		_w1630_,
		_w1631_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w1625_,
		_w1631_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w1615_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w1614_,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h4)
	) name633 (
		_w1603_,
		_w1634_,
		_w1635_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w1602_,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('h4)
	) name635 (
		_w1590_,
		_w1636_,
		_w1637_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w1589_,
		_w1637_,
		_w1638_
	);
	LUT2 #(
		.INIT('h8)
	) name637 (
		_w1358_,
		_w1638_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		_w1358_,
		_w1638_,
		_w1640_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w1639_,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		_w1314_,
		_w1315_,
		_w1642_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		_w1356_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h2)
	) name642 (
		_w1356_,
		_w1642_,
		_w1644_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w1643_,
		_w1644_,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w1589_,
		_w1590_,
		_w1646_
	);
	LUT2 #(
		.INIT('h4)
	) name645 (
		_w1636_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		_w1636_,
		_w1646_,
		_w1648_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w1647_,
		_w1648_,
		_w1649_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		_w1645_,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		_w1645_,
		_w1649_,
		_w1651_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w1324_,
		_w1325_,
		_w1652_
	);
	LUT2 #(
		.INIT('h4)
	) name651 (
		_w1354_,
		_w1652_,
		_w1653_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		_w1354_,
		_w1652_,
		_w1654_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w1653_,
		_w1654_,
		_w1655_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w1602_,
		_w1603_,
		_w1656_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		_w1634_,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w1634_,
		_w1656_,
		_w1658_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w1657_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h2)
	) name658 (
		_w1655_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h4)
	) name659 (
		_w1655_,
		_w1659_,
		_w1661_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		_w1614_,
		_w1615_,
		_w1662_
	);
	LUT2 #(
		.INIT('h4)
	) name661 (
		_w1632_,
		_w1662_,
		_w1663_
	);
	LUT2 #(
		.INIT('h2)
	) name662 (
		_w1632_,
		_w1662_,
		_w1664_
	);
	LUT2 #(
		.INIT('h1)
	) name663 (
		_w1663_,
		_w1664_,
		_w1665_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w1334_,
		_w1335_,
		_w1666_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		_w1352_,
		_w1666_,
		_w1667_
	);
	LUT2 #(
		.INIT('h2)
	) name666 (
		_w1352_,
		_w1666_,
		_w1668_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w1667_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w1665_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h8)
	) name669 (
		_w1665_,
		_w1669_,
		_w1671_
	);
	LUT2 #(
		.INIT('h1)
	) name670 (
		_w1617_,
		_w1619_,
		_w1672_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w1620_,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w1337_,
		_w1339_,
		_w1674_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		_w1340_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		_w1673_,
		_w1675_,
		_w1676_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w1345_,
		_w1346_,
		_w1677_
	);
	LUT2 #(
		.INIT('h4)
	) name676 (
		_w1350_,
		_w1677_,
		_w1678_
	);
	LUT2 #(
		.INIT('h2)
	) name677 (
		_w1350_,
		_w1677_,
		_w1679_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w1678_,
		_w1679_,
		_w1680_
	);
	LUT2 #(
		.INIT('h2)
	) name679 (
		_w1676_,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h4)
	) name680 (
		_w1676_,
		_w1680_,
		_w1682_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w1625_,
		_w1626_,
		_w1683_
	);
	LUT2 #(
		.INIT('h4)
	) name682 (
		_w1630_,
		_w1683_,
		_w1684_
	);
	LUT2 #(
		.INIT('h2)
	) name683 (
		_w1630_,
		_w1683_,
		_w1685_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w1684_,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h4)
	) name685 (
		_w1682_,
		_w1686_,
		_w1687_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		_w1681_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h4)
	) name687 (
		_w1671_,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		_w1670_,
		_w1689_,
		_w1690_
	);
	LUT2 #(
		.INIT('h4)
	) name689 (
		_w1661_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h1)
	) name690 (
		_w1660_,
		_w1691_,
		_w1692_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		_w1651_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h1)
	) name692 (
		_w1650_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h2)
	) name693 (
		_w1641_,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		_w1641_,
		_w1694_,
		_w1696_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h8)
	) name696 (
		\A[946] ,
		\A[947] ,
		_w1698_
	);
	LUT2 #(
		.INIT('h8)
	) name697 (
		\A[943] ,
		\A[944] ,
		_w1699_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		\A[943] ,
		\A[944] ,
		_w1700_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w1699_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h8)
	) name700 (
		\A[945] ,
		_w1701_,
		_w1702_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		\A[945] ,
		_w1701_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name702 (
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		\A[946] ,
		\A[947] ,
		_w1705_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w1698_,
		_w1705_,
		_w1706_
	);
	LUT2 #(
		.INIT('h8)
	) name705 (
		\A[948] ,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		\A[948] ,
		_w1706_,
		_w1708_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w1707_,
		_w1708_,
		_w1709_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		_w1704_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h8)
	) name709 (
		_w1698_,
		_w1710_,
		_w1711_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w1699_,
		_w1702_,
		_w1712_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w1698_,
		_w1707_,
		_w1713_
	);
	LUT2 #(
		.INIT('h4)
	) name712 (
		_w1710_,
		_w1713_,
		_w1714_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		_w1712_,
		_w1714_,
		_w1715_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w1711_,
		_w1715_,
		_w1716_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		\A[952] ,
		\A[953] ,
		_w1717_
	);
	LUT2 #(
		.INIT('h1)
	) name716 (
		\A[952] ,
		\A[953] ,
		_w1718_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w1717_,
		_w1718_,
		_w1719_
	);
	LUT2 #(
		.INIT('h8)
	) name718 (
		\A[954] ,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w1717_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('h8)
	) name720 (
		\A[949] ,
		\A[950] ,
		_w1722_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		\A[949] ,
		\A[950] ,
		_w1723_
	);
	LUT2 #(
		.INIT('h1)
	) name722 (
		_w1722_,
		_w1723_,
		_w1724_
	);
	LUT2 #(
		.INIT('h8)
	) name723 (
		\A[951] ,
		_w1724_,
		_w1725_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		_w1722_,
		_w1725_,
		_w1726_
	);
	LUT2 #(
		.INIT('h8)
	) name725 (
		_w1721_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		_w1721_,
		_w1726_,
		_w1728_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		\A[951] ,
		_w1724_,
		_w1729_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		_w1725_,
		_w1729_,
		_w1730_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		\A[954] ,
		_w1719_,
		_w1731_
	);
	LUT2 #(
		.INIT('h1)
	) name730 (
		_w1720_,
		_w1731_,
		_w1732_
	);
	LUT2 #(
		.INIT('h8)
	) name731 (
		_w1730_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w1728_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('h1)
	) name733 (
		_w1727_,
		_w1734_,
		_w1735_
	);
	LUT2 #(
		.INIT('h1)
	) name734 (
		_w1730_,
		_w1732_,
		_w1736_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w1733_,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w1704_,
		_w1709_,
		_w1738_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w1710_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h8)
	) name738 (
		_w1737_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h2)
	) name739 (
		_w1711_,
		_w1712_,
		_w1741_
	);
	LUT2 #(
		.INIT('h2)
	) name740 (
		_w1740_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w1727_,
		_w1728_,
		_w1743_
	);
	LUT2 #(
		.INIT('h2)
	) name742 (
		_w1733_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h4)
	) name743 (
		_w1733_,
		_w1743_,
		_w1745_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w1744_,
		_w1745_,
		_w1746_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		_w1742_,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w1742_,
		_w1746_,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w1711_,
		_w1714_,
		_w1749_
	);
	LUT2 #(
		.INIT('h2)
	) name748 (
		_w1712_,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		_w1712_,
		_w1749_,
		_w1751_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		_w1750_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		_w1748_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w1747_,
		_w1753_,
		_w1754_
	);
	LUT2 #(
		.INIT('h2)
	) name753 (
		_w1735_,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h4)
	) name754 (
		_w1735_,
		_w1754_,
		_w1756_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w1755_,
		_w1756_,
		_w1757_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		_w1716_,
		_w1757_,
		_w1758_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w1716_,
		_w1757_,
		_w1759_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		_w1758_,
		_w1759_,
		_w1760_
	);
	LUT2 #(
		.INIT('h8)
	) name759 (
		\A[958] ,
		\A[959] ,
		_w1761_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		\A[955] ,
		\A[956] ,
		_w1762_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		\A[955] ,
		\A[956] ,
		_w1763_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		_w1762_,
		_w1763_,
		_w1764_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		\A[957] ,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		\A[957] ,
		_w1764_,
		_w1766_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT2 #(
		.INIT('h1)
	) name766 (
		\A[958] ,
		\A[959] ,
		_w1768_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w1761_,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h8)
	) name768 (
		\A[960] ,
		_w1769_,
		_w1770_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		\A[960] ,
		_w1769_,
		_w1771_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w1770_,
		_w1771_,
		_w1772_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		_w1767_,
		_w1772_,
		_w1773_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		_w1761_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w1762_,
		_w1765_,
		_w1775_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w1761_,
		_w1770_,
		_w1776_
	);
	LUT2 #(
		.INIT('h4)
	) name775 (
		_w1773_,
		_w1776_,
		_w1777_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w1775_,
		_w1777_,
		_w1778_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		_w1774_,
		_w1778_,
		_w1779_
	);
	LUT2 #(
		.INIT('h8)
	) name778 (
		\A[964] ,
		\A[965] ,
		_w1780_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		\A[964] ,
		\A[965] ,
		_w1781_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w1780_,
		_w1781_,
		_w1782_
	);
	LUT2 #(
		.INIT('h8)
	) name781 (
		\A[966] ,
		_w1782_,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w1780_,
		_w1783_,
		_w1784_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		\A[961] ,
		\A[962] ,
		_w1785_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		\A[961] ,
		\A[962] ,
		_w1786_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w1785_,
		_w1786_,
		_w1787_
	);
	LUT2 #(
		.INIT('h8)
	) name786 (
		\A[963] ,
		_w1787_,
		_w1788_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		_w1785_,
		_w1788_,
		_w1789_
	);
	LUT2 #(
		.INIT('h8)
	) name788 (
		_w1784_,
		_w1789_,
		_w1790_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		_w1784_,
		_w1789_,
		_w1791_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		\A[963] ,
		_w1787_,
		_w1792_
	);
	LUT2 #(
		.INIT('h1)
	) name791 (
		_w1788_,
		_w1792_,
		_w1793_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		\A[966] ,
		_w1782_,
		_w1794_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w1783_,
		_w1794_,
		_w1795_
	);
	LUT2 #(
		.INIT('h8)
	) name794 (
		_w1793_,
		_w1795_,
		_w1796_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w1791_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h1)
	) name796 (
		_w1790_,
		_w1797_,
		_w1798_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w1793_,
		_w1795_,
		_w1799_
	);
	LUT2 #(
		.INIT('h1)
	) name798 (
		_w1796_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h1)
	) name799 (
		_w1767_,
		_w1772_,
		_w1801_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w1773_,
		_w1801_,
		_w1802_
	);
	LUT2 #(
		.INIT('h8)
	) name801 (
		_w1800_,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h2)
	) name802 (
		_w1774_,
		_w1775_,
		_w1804_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		_w1803_,
		_w1804_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w1790_,
		_w1791_,
		_w1806_
	);
	LUT2 #(
		.INIT('h2)
	) name805 (
		_w1796_,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		_w1796_,
		_w1806_,
		_w1808_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w1807_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h2)
	) name808 (
		_w1805_,
		_w1809_,
		_w1810_
	);
	LUT2 #(
		.INIT('h4)
	) name809 (
		_w1805_,
		_w1809_,
		_w1811_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w1774_,
		_w1777_,
		_w1812_
	);
	LUT2 #(
		.INIT('h2)
	) name811 (
		_w1775_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h4)
	) name812 (
		_w1775_,
		_w1812_,
		_w1814_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		_w1813_,
		_w1814_,
		_w1815_
	);
	LUT2 #(
		.INIT('h4)
	) name814 (
		_w1811_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w1810_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h2)
	) name816 (
		_w1798_,
		_w1817_,
		_w1818_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		_w1798_,
		_w1817_,
		_w1819_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w1818_,
		_w1819_,
		_w1820_
	);
	LUT2 #(
		.INIT('h8)
	) name819 (
		_w1779_,
		_w1820_,
		_w1821_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w1779_,
		_w1820_,
		_w1822_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w1821_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w1760_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h8)
	) name823 (
		_w1760_,
		_w1823_,
		_w1825_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w1800_,
		_w1802_,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		_w1803_,
		_w1826_,
		_w1827_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w1737_,
		_w1739_,
		_w1828_
	);
	LUT2 #(
		.INIT('h1)
	) name827 (
		_w1740_,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h8)
	) name828 (
		_w1827_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w1810_,
		_w1811_,
		_w1831_
	);
	LUT2 #(
		.INIT('h8)
	) name830 (
		_w1815_,
		_w1831_,
		_w1832_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		_w1815_,
		_w1831_,
		_w1833_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		_w1832_,
		_w1833_,
		_w1834_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		_w1830_,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h1)
	) name834 (
		_w1830_,
		_w1834_,
		_w1836_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w1747_,
		_w1748_,
		_w1837_
	);
	LUT2 #(
		.INIT('h8)
	) name836 (
		_w1752_,
		_w1837_,
		_w1838_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w1752_,
		_w1837_,
		_w1839_
	);
	LUT2 #(
		.INIT('h1)
	) name838 (
		_w1838_,
		_w1839_,
		_w1840_
	);
	LUT2 #(
		.INIT('h4)
	) name839 (
		_w1836_,
		_w1840_,
		_w1841_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		_w1835_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w1825_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		_w1824_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w1779_,
		_w1819_,
		_w1845_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		_w1818_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w1844_,
		_w1846_,
		_w1847_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		_w1844_,
		_w1846_,
		_w1848_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w1716_,
		_w1756_,
		_w1849_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w1755_,
		_w1849_,
		_w1850_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		_w1848_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w1847_,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h8)
	) name851 (
		\A[979] ,
		\A[980] ,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		\A[979] ,
		\A[980] ,
		_w1854_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w1853_,
		_w1854_,
		_w1855_
	);
	LUT2 #(
		.INIT('h8)
	) name854 (
		\A[981] ,
		_w1855_,
		_w1856_
	);
	LUT2 #(
		.INIT('h1)
	) name855 (
		\A[981] ,
		_w1855_,
		_w1857_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w1856_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h8)
	) name857 (
		\A[982] ,
		\A[983] ,
		_w1859_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		\A[982] ,
		\A[983] ,
		_w1860_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w1859_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h8)
	) name860 (
		\A[984] ,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		\A[984] ,
		_w1861_,
		_w1863_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w1862_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		_w1858_,
		_w1864_,
		_w1865_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w1858_,
		_w1864_,
		_w1866_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		_w1865_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\A[985] ,
		\A[986] ,
		_w1868_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		\A[985] ,
		\A[986] ,
		_w1869_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h8)
	) name869 (
		\A[987] ,
		_w1870_,
		_w1871_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		\A[987] ,
		_w1870_,
		_w1872_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w1871_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h8)
	) name872 (
		\A[988] ,
		\A[989] ,
		_w1874_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		\A[988] ,
		\A[989] ,
		_w1875_
	);
	LUT2 #(
		.INIT('h1)
	) name874 (
		_w1874_,
		_w1875_,
		_w1876_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		\A[990] ,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		\A[990] ,
		_w1876_,
		_w1878_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w1877_,
		_w1878_,
		_w1879_
	);
	LUT2 #(
		.INIT('h8)
	) name878 (
		_w1873_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h1)
	) name879 (
		_w1873_,
		_w1879_,
		_w1881_
	);
	LUT2 #(
		.INIT('h1)
	) name880 (
		_w1880_,
		_w1881_,
		_w1882_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		_w1867_,
		_w1882_,
		_w1883_
	);
	LUT2 #(
		.INIT('h1)
	) name882 (
		_w1874_,
		_w1877_,
		_w1884_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		_w1868_,
		_w1871_,
		_w1885_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		_w1884_,
		_w1885_,
		_w1887_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		_w1886_,
		_w1887_,
		_w1888_
	);
	LUT2 #(
		.INIT('h8)
	) name887 (
		_w1883_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h1)
	) name888 (
		_w1859_,
		_w1862_,
		_w1890_
	);
	LUT2 #(
		.INIT('h1)
	) name889 (
		_w1853_,
		_w1856_,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		_w1890_,
		_w1891_,
		_w1892_
	);
	LUT2 #(
		.INIT('h8)
	) name891 (
		_w1890_,
		_w1891_,
		_w1893_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1892_,
		_w1893_,
		_w1894_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		_w1865_,
		_w1894_,
		_w1895_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		_w1865_,
		_w1894_,
		_w1896_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w1895_,
		_w1896_,
		_w1897_
	);
	LUT2 #(
		.INIT('h4)
	) name896 (
		_w1889_,
		_w1897_,
		_w1898_
	);
	LUT2 #(
		.INIT('h4)
	) name897 (
		_w1880_,
		_w1888_,
		_w1899_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		_w1880_,
		_w1888_,
		_w1900_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w1883_,
		_w1899_,
		_w1901_
	);
	LUT2 #(
		.INIT('h4)
	) name900 (
		_w1900_,
		_w1901_,
		_w1902_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w1898_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h2)
	) name902 (
		_w1880_,
		_w1886_,
		_w1904_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w1887_,
		_w1904_,
		_w1905_
	);
	LUT2 #(
		.INIT('h4)
	) name904 (
		_w1903_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h2)
	) name905 (
		_w1903_,
		_w1905_,
		_w1907_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w1865_,
		_w1892_,
		_w1908_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w1893_,
		_w1908_,
		_w1909_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		_w1907_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		_w1906_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		\A[967] ,
		\A[968] ,
		_w1912_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		\A[967] ,
		\A[968] ,
		_w1913_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1912_,
		_w1913_,
		_w1914_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		\A[969] ,
		_w1914_,
		_w1915_
	);
	LUT2 #(
		.INIT('h1)
	) name914 (
		\A[969] ,
		_w1914_,
		_w1916_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w1915_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h8)
	) name916 (
		\A[970] ,
		\A[971] ,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		\A[970] ,
		\A[971] ,
		_w1919_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		_w1918_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h8)
	) name919 (
		\A[972] ,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		\A[972] ,
		_w1920_,
		_w1922_
	);
	LUT2 #(
		.INIT('h1)
	) name921 (
		_w1921_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		_w1917_,
		_w1923_,
		_w1924_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		_w1917_,
		_w1923_,
		_w1925_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w1924_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h8)
	) name925 (
		\A[973] ,
		\A[974] ,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		\A[973] ,
		\A[974] ,
		_w1928_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1927_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		\A[975] ,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h1)
	) name929 (
		\A[975] ,
		_w1929_,
		_w1931_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w1930_,
		_w1931_,
		_w1932_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		\A[976] ,
		\A[977] ,
		_w1933_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		\A[976] ,
		\A[977] ,
		_w1934_
	);
	LUT2 #(
		.INIT('h1)
	) name933 (
		_w1933_,
		_w1934_,
		_w1935_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		\A[978] ,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h1)
	) name935 (
		\A[978] ,
		_w1935_,
		_w1937_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1936_,
		_w1937_,
		_w1938_
	);
	LUT2 #(
		.INIT('h8)
	) name937 (
		_w1932_,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h1)
	) name938 (
		_w1932_,
		_w1938_,
		_w1940_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w1939_,
		_w1940_,
		_w1941_
	);
	LUT2 #(
		.INIT('h8)
	) name940 (
		_w1926_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h1)
	) name941 (
		_w1933_,
		_w1936_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name942 (
		_w1927_,
		_w1930_,
		_w1944_
	);
	LUT2 #(
		.INIT('h8)
	) name943 (
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w1943_,
		_w1944_,
		_w1946_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		_w1945_,
		_w1946_,
		_w1947_
	);
	LUT2 #(
		.INIT('h8)
	) name946 (
		_w1942_,
		_w1947_,
		_w1948_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w1918_,
		_w1921_,
		_w1949_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w1912_,
		_w1915_,
		_w1950_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w1949_,
		_w1950_,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		_w1949_,
		_w1950_,
		_w1952_
	);
	LUT2 #(
		.INIT('h1)
	) name951 (
		_w1951_,
		_w1952_,
		_w1953_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		_w1924_,
		_w1953_,
		_w1954_
	);
	LUT2 #(
		.INIT('h4)
	) name953 (
		_w1924_,
		_w1953_,
		_w1955_
	);
	LUT2 #(
		.INIT('h1)
	) name954 (
		_w1954_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		_w1948_,
		_w1956_,
		_w1957_
	);
	LUT2 #(
		.INIT('h4)
	) name956 (
		_w1939_,
		_w1947_,
		_w1958_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		_w1939_,
		_w1947_,
		_w1959_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w1942_,
		_w1958_,
		_w1960_
	);
	LUT2 #(
		.INIT('h4)
	) name959 (
		_w1959_,
		_w1960_,
		_w1961_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w1957_,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h2)
	) name961 (
		_w1939_,
		_w1945_,
		_w1963_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		_w1946_,
		_w1963_,
		_w1964_
	);
	LUT2 #(
		.INIT('h4)
	) name963 (
		_w1962_,
		_w1964_,
		_w1965_
	);
	LUT2 #(
		.INIT('h2)
	) name964 (
		_w1962_,
		_w1964_,
		_w1966_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w1924_,
		_w1951_,
		_w1967_
	);
	LUT2 #(
		.INIT('h1)
	) name966 (
		_w1952_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w1966_,
		_w1968_,
		_w1969_
	);
	LUT2 #(
		.INIT('h1)
	) name968 (
		_w1965_,
		_w1969_,
		_w1970_
	);
	LUT2 #(
		.INIT('h8)
	) name969 (
		_w1911_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1911_,
		_w1970_,
		_w1972_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		_w1965_,
		_w1966_,
		_w1973_
	);
	LUT2 #(
		.INIT('h4)
	) name972 (
		_w1968_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h2)
	) name973 (
		_w1968_,
		_w1973_,
		_w1975_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		_w1974_,
		_w1975_,
		_w1976_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		_w1906_,
		_w1907_,
		_w1977_
	);
	LUT2 #(
		.INIT('h4)
	) name976 (
		_w1909_,
		_w1977_,
		_w1978_
	);
	LUT2 #(
		.INIT('h2)
	) name977 (
		_w1909_,
		_w1977_,
		_w1979_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		_w1978_,
		_w1979_,
		_w1980_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1976_,
		_w1980_,
		_w1981_
	);
	LUT2 #(
		.INIT('h8)
	) name980 (
		_w1976_,
		_w1980_,
		_w1982_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w1867_,
		_w1882_,
		_w1983_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		_w1883_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		_w1926_,
		_w1941_,
		_w1985_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w1942_,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('h8)
	) name985 (
		_w1984_,
		_w1986_,
		_w1987_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		_w1889_,
		_w1902_,
		_w1988_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		_w1897_,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w1897_,
		_w1988_,
		_w1990_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w1989_,
		_w1990_,
		_w1991_
	);
	LUT2 #(
		.INIT('h2)
	) name990 (
		_w1987_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		_w1987_,
		_w1991_,
		_w1993_
	);
	LUT2 #(
		.INIT('h1)
	) name992 (
		_w1948_,
		_w1961_,
		_w1994_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		_w1956_,
		_w1994_,
		_w1995_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w1956_,
		_w1994_,
		_w1996_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w1995_,
		_w1996_,
		_w1997_
	);
	LUT2 #(
		.INIT('h1)
	) name996 (
		_w1993_,
		_w1997_,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w1992_,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		_w1982_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		_w1981_,
		_w2000_,
		_w2001_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w1972_,
		_w2001_,
		_w2002_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		_w1971_,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1852_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h8)
	) name1003 (
		_w1852_,
		_w2003_,
		_w2005_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w1847_,
		_w1848_,
		_w2006_
	);
	LUT2 #(
		.INIT('h4)
	) name1005 (
		_w1850_,
		_w2006_,
		_w2007_
	);
	LUT2 #(
		.INIT('h2)
	) name1006 (
		_w1850_,
		_w2006_,
		_w2008_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		_w2007_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h1)
	) name1008 (
		_w1971_,
		_w1972_,
		_w2010_
	);
	LUT2 #(
		.INIT('h4)
	) name1009 (
		_w2001_,
		_w2010_,
		_w2011_
	);
	LUT2 #(
		.INIT('h2)
	) name1010 (
		_w2001_,
		_w2010_,
		_w2012_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w2011_,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name1012 (
		_w2009_,
		_w2013_,
		_w2014_
	);
	LUT2 #(
		.INIT('h1)
	) name1013 (
		_w2009_,
		_w2013_,
		_w2015_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		_w1824_,
		_w1825_,
		_w2016_
	);
	LUT2 #(
		.INIT('h4)
	) name1015 (
		_w1842_,
		_w2016_,
		_w2017_
	);
	LUT2 #(
		.INIT('h2)
	) name1016 (
		_w1842_,
		_w2016_,
		_w2018_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w1981_,
		_w1982_,
		_w2020_
	);
	LUT2 #(
		.INIT('h4)
	) name1019 (
		_w1999_,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('h2)
	) name1020 (
		_w1999_,
		_w2020_,
		_w2022_
	);
	LUT2 #(
		.INIT('h1)
	) name1021 (
		_w2021_,
		_w2022_,
		_w2023_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		_w2019_,
		_w2023_,
		_w2024_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		_w2019_,
		_w2023_,
		_w2025_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w1984_,
		_w1986_,
		_w2026_
	);
	LUT2 #(
		.INIT('h1)
	) name1025 (
		_w1987_,
		_w2026_,
		_w2027_
	);
	LUT2 #(
		.INIT('h1)
	) name1026 (
		_w1827_,
		_w1829_,
		_w2028_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		_w1830_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h8)
	) name1028 (
		_w2027_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h1)
	) name1029 (
		_w1992_,
		_w1993_,
		_w2031_
	);
	LUT2 #(
		.INIT('h4)
	) name1030 (
		_w1997_,
		_w2031_,
		_w2032_
	);
	LUT2 #(
		.INIT('h2)
	) name1031 (
		_w1997_,
		_w2031_,
		_w2033_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		_w2032_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		_w2030_,
		_w2034_,
		_w2035_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w2030_,
		_w2034_,
		_w2036_
	);
	LUT2 #(
		.INIT('h1)
	) name1035 (
		_w1835_,
		_w1836_,
		_w2037_
	);
	LUT2 #(
		.INIT('h4)
	) name1036 (
		_w1840_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('h2)
	) name1037 (
		_w1840_,
		_w2037_,
		_w2039_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w2038_,
		_w2039_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name1039 (
		_w2036_,
		_w2040_,
		_w2041_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w2035_,
		_w2041_,
		_w2042_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w2025_,
		_w2042_,
		_w2043_
	);
	LUT2 #(
		.INIT('h1)
	) name1042 (
		_w2024_,
		_w2043_,
		_w2044_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		_w2015_,
		_w2044_,
		_w2045_
	);
	LUT2 #(
		.INIT('h1)
	) name1044 (
		_w2014_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h1)
	) name1045 (
		_w2005_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h1)
	) name1046 (
		_w2004_,
		_w2047_,
		_w2048_
	);
	LUT2 #(
		.INIT('h2)
	) name1047 (
		_w1697_,
		_w2048_,
		_w2049_
	);
	LUT2 #(
		.INIT('h4)
	) name1048 (
		_w1697_,
		_w2048_,
		_w2050_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		_w2004_,
		_w2005_,
		_w2051_
	);
	LUT2 #(
		.INIT('h4)
	) name1050 (
		_w2046_,
		_w2051_,
		_w2052_
	);
	LUT2 #(
		.INIT('h2)
	) name1051 (
		_w2046_,
		_w2051_,
		_w2053_
	);
	LUT2 #(
		.INIT('h1)
	) name1052 (
		_w2052_,
		_w2053_,
		_w2054_
	);
	LUT2 #(
		.INIT('h1)
	) name1053 (
		_w1650_,
		_w1651_,
		_w2055_
	);
	LUT2 #(
		.INIT('h4)
	) name1054 (
		_w1692_,
		_w2055_,
		_w2056_
	);
	LUT2 #(
		.INIT('h2)
	) name1055 (
		_w1692_,
		_w2055_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name1056 (
		_w2056_,
		_w2057_,
		_w2058_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		_w2054_,
		_w2058_,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name1058 (
		_w2054_,
		_w2058_,
		_w2060_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		_w1660_,
		_w1661_,
		_w2061_
	);
	LUT2 #(
		.INIT('h8)
	) name1060 (
		_w1690_,
		_w2061_,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name1061 (
		_w1690_,
		_w2061_,
		_w2063_
	);
	LUT2 #(
		.INIT('h1)
	) name1062 (
		_w2062_,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h1)
	) name1063 (
		_w2014_,
		_w2015_,
		_w2065_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w2044_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h2)
	) name1065 (
		_w2044_,
		_w2065_,
		_w2067_
	);
	LUT2 #(
		.INIT('h1)
	) name1066 (
		_w2066_,
		_w2067_,
		_w2068_
	);
	LUT2 #(
		.INIT('h1)
	) name1067 (
		_w2064_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		_w2064_,
		_w2068_,
		_w2070_
	);
	LUT2 #(
		.INIT('h1)
	) name1069 (
		_w2024_,
		_w2025_,
		_w2071_
	);
	LUT2 #(
		.INIT('h4)
	) name1070 (
		_w2042_,
		_w2071_,
		_w2072_
	);
	LUT2 #(
		.INIT('h2)
	) name1071 (
		_w2042_,
		_w2071_,
		_w2073_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w2072_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h1)
	) name1073 (
		_w1670_,
		_w1671_,
		_w2075_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		_w1688_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h2)
	) name1075 (
		_w1688_,
		_w2075_,
		_w2077_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w2076_,
		_w2077_,
		_w2078_
	);
	LUT2 #(
		.INIT('h1)
	) name1077 (
		_w2074_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h8)
	) name1078 (
		_w2074_,
		_w2078_,
		_w2080_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w1673_,
		_w1675_,
		_w2081_
	);
	LUT2 #(
		.INIT('h1)
	) name1080 (
		_w1676_,
		_w2081_,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w2027_,
		_w2029_,
		_w2083_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		_w2030_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		_w2082_,
		_w2084_,
		_w2085_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w1681_,
		_w1682_,
		_w2086_
	);
	LUT2 #(
		.INIT('h4)
	) name1085 (
		_w1686_,
		_w2086_,
		_w2087_
	);
	LUT2 #(
		.INIT('h2)
	) name1086 (
		_w1686_,
		_w2086_,
		_w2088_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		_w2087_,
		_w2088_,
		_w2089_
	);
	LUT2 #(
		.INIT('h2)
	) name1088 (
		_w2085_,
		_w2089_,
		_w2090_
	);
	LUT2 #(
		.INIT('h4)
	) name1089 (
		_w2085_,
		_w2089_,
		_w2091_
	);
	LUT2 #(
		.INIT('h1)
	) name1090 (
		_w2035_,
		_w2036_,
		_w2092_
	);
	LUT2 #(
		.INIT('h4)
	) name1091 (
		_w2040_,
		_w2092_,
		_w2093_
	);
	LUT2 #(
		.INIT('h2)
	) name1092 (
		_w2040_,
		_w2092_,
		_w2094_
	);
	LUT2 #(
		.INIT('h1)
	) name1093 (
		_w2093_,
		_w2094_,
		_w2095_
	);
	LUT2 #(
		.INIT('h4)
	) name1094 (
		_w2091_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h1)
	) name1095 (
		_w2090_,
		_w2096_,
		_w2097_
	);
	LUT2 #(
		.INIT('h4)
	) name1096 (
		_w2080_,
		_w2097_,
		_w2098_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w2079_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h1)
	) name1098 (
		_w2070_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		_w2069_,
		_w2100_,
		_w2101_
	);
	LUT2 #(
		.INIT('h1)
	) name1100 (
		_w2060_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h1)
	) name1101 (
		_w2059_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h4)
	) name1102 (
		_w2050_,
		_w2103_,
		_w2104_
	);
	LUT2 #(
		.INIT('h1)
	) name1103 (
		_w2049_,
		_w2104_,
		_w2105_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		_w1639_,
		_w1694_,
		_w2106_
	);
	LUT2 #(
		.INIT('h1)
	) name1105 (
		_w1640_,
		_w2106_,
		_w2107_
	);
	LUT2 #(
		.INIT('h1)
	) name1106 (
		_w2105_,
		_w2107_,
		_w2108_
	);
	LUT2 #(
		.INIT('h8)
	) name1107 (
		_w2105_,
		_w2107_,
		_w2109_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w2108_,
		_w2109_,
		_w2110_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		\A[874] ,
		\A[875] ,
		_w2111_
	);
	LUT2 #(
		.INIT('h8)
	) name1110 (
		\A[871] ,
		\A[872] ,
		_w2112_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		\A[871] ,
		\A[872] ,
		_w2113_
	);
	LUT2 #(
		.INIT('h1)
	) name1112 (
		_w2112_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h8)
	) name1113 (
		\A[873] ,
		_w2114_,
		_w2115_
	);
	LUT2 #(
		.INIT('h1)
	) name1114 (
		\A[873] ,
		_w2114_,
		_w2116_
	);
	LUT2 #(
		.INIT('h1)
	) name1115 (
		_w2115_,
		_w2116_,
		_w2117_
	);
	LUT2 #(
		.INIT('h1)
	) name1116 (
		\A[874] ,
		\A[875] ,
		_w2118_
	);
	LUT2 #(
		.INIT('h1)
	) name1117 (
		_w2111_,
		_w2118_,
		_w2119_
	);
	LUT2 #(
		.INIT('h8)
	) name1118 (
		\A[876] ,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		\A[876] ,
		_w2119_,
		_w2121_
	);
	LUT2 #(
		.INIT('h1)
	) name1120 (
		_w2120_,
		_w2121_,
		_w2122_
	);
	LUT2 #(
		.INIT('h8)
	) name1121 (
		_w2117_,
		_w2122_,
		_w2123_
	);
	LUT2 #(
		.INIT('h8)
	) name1122 (
		_w2111_,
		_w2123_,
		_w2124_
	);
	LUT2 #(
		.INIT('h1)
	) name1123 (
		_w2112_,
		_w2115_,
		_w2125_
	);
	LUT2 #(
		.INIT('h1)
	) name1124 (
		_w2111_,
		_w2120_,
		_w2126_
	);
	LUT2 #(
		.INIT('h4)
	) name1125 (
		_w2123_,
		_w2126_,
		_w2127_
	);
	LUT2 #(
		.INIT('h1)
	) name1126 (
		_w2125_,
		_w2127_,
		_w2128_
	);
	LUT2 #(
		.INIT('h1)
	) name1127 (
		_w2124_,
		_w2128_,
		_w2129_
	);
	LUT2 #(
		.INIT('h8)
	) name1128 (
		\A[880] ,
		\A[881] ,
		_w2130_
	);
	LUT2 #(
		.INIT('h1)
	) name1129 (
		\A[880] ,
		\A[881] ,
		_w2131_
	);
	LUT2 #(
		.INIT('h1)
	) name1130 (
		_w2130_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h8)
	) name1131 (
		\A[882] ,
		_w2132_,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name1132 (
		_w2130_,
		_w2133_,
		_w2134_
	);
	LUT2 #(
		.INIT('h8)
	) name1133 (
		\A[877] ,
		\A[878] ,
		_w2135_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		\A[877] ,
		\A[878] ,
		_w2136_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		_w2135_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h8)
	) name1136 (
		\A[879] ,
		_w2137_,
		_w2138_
	);
	LUT2 #(
		.INIT('h1)
	) name1137 (
		_w2135_,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h8)
	) name1138 (
		_w2134_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		_w2134_,
		_w2139_,
		_w2141_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		\A[879] ,
		_w2137_,
		_w2142_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w2138_,
		_w2142_,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name1142 (
		\A[882] ,
		_w2132_,
		_w2144_
	);
	LUT2 #(
		.INIT('h1)
	) name1143 (
		_w2133_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h8)
	) name1144 (
		_w2143_,
		_w2145_,
		_w2146_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		_w2141_,
		_w2146_,
		_w2147_
	);
	LUT2 #(
		.INIT('h1)
	) name1146 (
		_w2140_,
		_w2147_,
		_w2148_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		_w2143_,
		_w2145_,
		_w2149_
	);
	LUT2 #(
		.INIT('h1)
	) name1148 (
		_w2146_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w2117_,
		_w2122_,
		_w2151_
	);
	LUT2 #(
		.INIT('h1)
	) name1150 (
		_w2123_,
		_w2151_,
		_w2152_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		_w2150_,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h2)
	) name1152 (
		_w2124_,
		_w2125_,
		_w2154_
	);
	LUT2 #(
		.INIT('h2)
	) name1153 (
		_w2153_,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h1)
	) name1154 (
		_w2140_,
		_w2141_,
		_w2156_
	);
	LUT2 #(
		.INIT('h2)
	) name1155 (
		_w2146_,
		_w2156_,
		_w2157_
	);
	LUT2 #(
		.INIT('h4)
	) name1156 (
		_w2146_,
		_w2156_,
		_w2158_
	);
	LUT2 #(
		.INIT('h1)
	) name1157 (
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h2)
	) name1158 (
		_w2155_,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h4)
	) name1159 (
		_w2155_,
		_w2159_,
		_w2161_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		_w2124_,
		_w2127_,
		_w2162_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		_w2125_,
		_w2162_,
		_w2163_
	);
	LUT2 #(
		.INIT('h4)
	) name1162 (
		_w2125_,
		_w2162_,
		_w2164_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w2163_,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h4)
	) name1164 (
		_w2161_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		_w2160_,
		_w2166_,
		_w2167_
	);
	LUT2 #(
		.INIT('h2)
	) name1166 (
		_w2148_,
		_w2167_,
		_w2168_
	);
	LUT2 #(
		.INIT('h4)
	) name1167 (
		_w2148_,
		_w2167_,
		_w2169_
	);
	LUT2 #(
		.INIT('h1)
	) name1168 (
		_w2168_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h8)
	) name1169 (
		_w2129_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		_w2129_,
		_w2170_,
		_w2172_
	);
	LUT2 #(
		.INIT('h1)
	) name1171 (
		_w2171_,
		_w2172_,
		_w2173_
	);
	LUT2 #(
		.INIT('h8)
	) name1172 (
		\A[886] ,
		\A[887] ,
		_w2174_
	);
	LUT2 #(
		.INIT('h8)
	) name1173 (
		\A[883] ,
		\A[884] ,
		_w2175_
	);
	LUT2 #(
		.INIT('h1)
	) name1174 (
		\A[883] ,
		\A[884] ,
		_w2176_
	);
	LUT2 #(
		.INIT('h1)
	) name1175 (
		_w2175_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		\A[885] ,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h1)
	) name1177 (
		\A[885] ,
		_w2177_,
		_w2179_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		_w2178_,
		_w2179_,
		_w2180_
	);
	LUT2 #(
		.INIT('h1)
	) name1179 (
		\A[886] ,
		\A[887] ,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		_w2174_,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h8)
	) name1181 (
		\A[888] ,
		_w2182_,
		_w2183_
	);
	LUT2 #(
		.INIT('h1)
	) name1182 (
		\A[888] ,
		_w2182_,
		_w2184_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w2183_,
		_w2184_,
		_w2185_
	);
	LUT2 #(
		.INIT('h8)
	) name1184 (
		_w2180_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h8)
	) name1185 (
		_w2174_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h1)
	) name1186 (
		_w2175_,
		_w2178_,
		_w2188_
	);
	LUT2 #(
		.INIT('h1)
	) name1187 (
		_w2174_,
		_w2183_,
		_w2189_
	);
	LUT2 #(
		.INIT('h4)
	) name1188 (
		_w2186_,
		_w2189_,
		_w2190_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		_w2188_,
		_w2190_,
		_w2191_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		_w2187_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name1191 (
		\A[892] ,
		\A[893] ,
		_w2193_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		\A[892] ,
		\A[893] ,
		_w2194_
	);
	LUT2 #(
		.INIT('h1)
	) name1193 (
		_w2193_,
		_w2194_,
		_w2195_
	);
	LUT2 #(
		.INIT('h8)
	) name1194 (
		\A[894] ,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h1)
	) name1195 (
		_w2193_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h8)
	) name1196 (
		\A[889] ,
		\A[890] ,
		_w2198_
	);
	LUT2 #(
		.INIT('h1)
	) name1197 (
		\A[889] ,
		\A[890] ,
		_w2199_
	);
	LUT2 #(
		.INIT('h1)
	) name1198 (
		_w2198_,
		_w2199_,
		_w2200_
	);
	LUT2 #(
		.INIT('h8)
	) name1199 (
		\A[891] ,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h1)
	) name1200 (
		_w2198_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h8)
	) name1201 (
		_w2197_,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		_w2197_,
		_w2202_,
		_w2204_
	);
	LUT2 #(
		.INIT('h1)
	) name1203 (
		\A[891] ,
		_w2200_,
		_w2205_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		_w2201_,
		_w2205_,
		_w2206_
	);
	LUT2 #(
		.INIT('h1)
	) name1205 (
		\A[894] ,
		_w2195_,
		_w2207_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w2196_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h8)
	) name1207 (
		_w2206_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h1)
	) name1208 (
		_w2204_,
		_w2209_,
		_w2210_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w2203_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h1)
	) name1210 (
		_w2206_,
		_w2208_,
		_w2212_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w2209_,
		_w2212_,
		_w2213_
	);
	LUT2 #(
		.INIT('h1)
	) name1212 (
		_w2180_,
		_w2185_,
		_w2214_
	);
	LUT2 #(
		.INIT('h1)
	) name1213 (
		_w2186_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		_w2213_,
		_w2215_,
		_w2216_
	);
	LUT2 #(
		.INIT('h2)
	) name1215 (
		_w2187_,
		_w2188_,
		_w2217_
	);
	LUT2 #(
		.INIT('h2)
	) name1216 (
		_w2216_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h1)
	) name1217 (
		_w2203_,
		_w2204_,
		_w2219_
	);
	LUT2 #(
		.INIT('h2)
	) name1218 (
		_w2209_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h4)
	) name1219 (
		_w2209_,
		_w2219_,
		_w2221_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w2220_,
		_w2221_,
		_w2222_
	);
	LUT2 #(
		.INIT('h2)
	) name1221 (
		_w2218_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h4)
	) name1222 (
		_w2218_,
		_w2222_,
		_w2224_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w2187_,
		_w2190_,
		_w2225_
	);
	LUT2 #(
		.INIT('h2)
	) name1224 (
		_w2188_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h4)
	) name1225 (
		_w2188_,
		_w2225_,
		_w2227_
	);
	LUT2 #(
		.INIT('h1)
	) name1226 (
		_w2226_,
		_w2227_,
		_w2228_
	);
	LUT2 #(
		.INIT('h4)
	) name1227 (
		_w2224_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w2223_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('h2)
	) name1229 (
		_w2211_,
		_w2230_,
		_w2231_
	);
	LUT2 #(
		.INIT('h4)
	) name1230 (
		_w2211_,
		_w2230_,
		_w2232_
	);
	LUT2 #(
		.INIT('h1)
	) name1231 (
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h8)
	) name1232 (
		_w2192_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h1)
	) name1233 (
		_w2192_,
		_w2233_,
		_w2235_
	);
	LUT2 #(
		.INIT('h1)
	) name1234 (
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h1)
	) name1235 (
		_w2173_,
		_w2236_,
		_w2237_
	);
	LUT2 #(
		.INIT('h8)
	) name1236 (
		_w2173_,
		_w2236_,
		_w2238_
	);
	LUT2 #(
		.INIT('h1)
	) name1237 (
		_w2213_,
		_w2215_,
		_w2239_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		_w2216_,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		_w2150_,
		_w2152_,
		_w2241_
	);
	LUT2 #(
		.INIT('h1)
	) name1240 (
		_w2153_,
		_w2241_,
		_w2242_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		_w2240_,
		_w2242_,
		_w2243_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w2223_,
		_w2224_,
		_w2244_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		_w2228_,
		_w2244_,
		_w2245_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w2228_,
		_w2244_,
		_w2246_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h8)
	) name1246 (
		_w2243_,
		_w2247_,
		_w2248_
	);
	LUT2 #(
		.INIT('h1)
	) name1247 (
		_w2243_,
		_w2247_,
		_w2249_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w2160_,
		_w2161_,
		_w2250_
	);
	LUT2 #(
		.INIT('h8)
	) name1249 (
		_w2165_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h1)
	) name1250 (
		_w2165_,
		_w2250_,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name1251 (
		_w2251_,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h4)
	) name1252 (
		_w2249_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		_w2248_,
		_w2254_,
		_w2255_
	);
	LUT2 #(
		.INIT('h1)
	) name1254 (
		_w2238_,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h1)
	) name1255 (
		_w2237_,
		_w2256_,
		_w2257_
	);
	LUT2 #(
		.INIT('h1)
	) name1256 (
		_w2192_,
		_w2232_,
		_w2258_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w2231_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h1)
	) name1258 (
		_w2257_,
		_w2259_,
		_w2260_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		_w2257_,
		_w2259_,
		_w2261_
	);
	LUT2 #(
		.INIT('h1)
	) name1260 (
		_w2129_,
		_w2169_,
		_w2262_
	);
	LUT2 #(
		.INIT('h1)
	) name1261 (
		_w2168_,
		_w2262_,
		_w2263_
	);
	LUT2 #(
		.INIT('h1)
	) name1262 (
		_w2261_,
		_w2263_,
		_w2264_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w2260_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h1)
	) name1264 (
		_w2260_,
		_w2261_,
		_w2266_
	);
	LUT2 #(
		.INIT('h4)
	) name1265 (
		_w2263_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h2)
	) name1266 (
		_w2263_,
		_w2266_,
		_w2268_
	);
	LUT2 #(
		.INIT('h1)
	) name1267 (
		_w2267_,
		_w2268_,
		_w2269_
	);
	LUT2 #(
		.INIT('h8)
	) name1268 (
		\A[850] ,
		\A[851] ,
		_w2270_
	);
	LUT2 #(
		.INIT('h8)
	) name1269 (
		\A[847] ,
		\A[848] ,
		_w2271_
	);
	LUT2 #(
		.INIT('h1)
	) name1270 (
		\A[847] ,
		\A[848] ,
		_w2272_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		_w2271_,
		_w2272_,
		_w2273_
	);
	LUT2 #(
		.INIT('h8)
	) name1272 (
		\A[849] ,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h1)
	) name1273 (
		\A[849] ,
		_w2273_,
		_w2275_
	);
	LUT2 #(
		.INIT('h1)
	) name1274 (
		_w2274_,
		_w2275_,
		_w2276_
	);
	LUT2 #(
		.INIT('h1)
	) name1275 (
		\A[850] ,
		\A[851] ,
		_w2277_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w2270_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		\A[852] ,
		_w2278_,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name1278 (
		\A[852] ,
		_w2278_,
		_w2280_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w2279_,
		_w2280_,
		_w2281_
	);
	LUT2 #(
		.INIT('h8)
	) name1280 (
		_w2276_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h8)
	) name1281 (
		_w2270_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h1)
	) name1282 (
		_w2271_,
		_w2274_,
		_w2284_
	);
	LUT2 #(
		.INIT('h1)
	) name1283 (
		_w2270_,
		_w2279_,
		_w2285_
	);
	LUT2 #(
		.INIT('h4)
	) name1284 (
		_w2282_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h1)
	) name1285 (
		_w2284_,
		_w2286_,
		_w2287_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w2283_,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('h8)
	) name1287 (
		\A[856] ,
		\A[857] ,
		_w2289_
	);
	LUT2 #(
		.INIT('h1)
	) name1288 (
		\A[856] ,
		\A[857] ,
		_w2290_
	);
	LUT2 #(
		.INIT('h1)
	) name1289 (
		_w2289_,
		_w2290_,
		_w2291_
	);
	LUT2 #(
		.INIT('h8)
	) name1290 (
		\A[858] ,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h1)
	) name1291 (
		_w2289_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h8)
	) name1292 (
		\A[853] ,
		\A[854] ,
		_w2294_
	);
	LUT2 #(
		.INIT('h1)
	) name1293 (
		\A[853] ,
		\A[854] ,
		_w2295_
	);
	LUT2 #(
		.INIT('h1)
	) name1294 (
		_w2294_,
		_w2295_,
		_w2296_
	);
	LUT2 #(
		.INIT('h8)
	) name1295 (
		\A[855] ,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		_w2294_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h8)
	) name1297 (
		_w2293_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h1)
	) name1298 (
		_w2293_,
		_w2298_,
		_w2300_
	);
	LUT2 #(
		.INIT('h1)
	) name1299 (
		\A[855] ,
		_w2296_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name1300 (
		_w2297_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h1)
	) name1301 (
		\A[858] ,
		_w2291_,
		_w2303_
	);
	LUT2 #(
		.INIT('h1)
	) name1302 (
		_w2292_,
		_w2303_,
		_w2304_
	);
	LUT2 #(
		.INIT('h8)
	) name1303 (
		_w2302_,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h1)
	) name1304 (
		_w2300_,
		_w2305_,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name1305 (
		_w2299_,
		_w2306_,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		_w2302_,
		_w2304_,
		_w2308_
	);
	LUT2 #(
		.INIT('h1)
	) name1307 (
		_w2305_,
		_w2308_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name1308 (
		_w2276_,
		_w2281_,
		_w2310_
	);
	LUT2 #(
		.INIT('h1)
	) name1309 (
		_w2282_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name1310 (
		_w2309_,
		_w2311_,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name1311 (
		_w2283_,
		_w2284_,
		_w2313_
	);
	LUT2 #(
		.INIT('h2)
	) name1312 (
		_w2312_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h1)
	) name1313 (
		_w2299_,
		_w2300_,
		_w2315_
	);
	LUT2 #(
		.INIT('h2)
	) name1314 (
		_w2305_,
		_w2315_,
		_w2316_
	);
	LUT2 #(
		.INIT('h4)
	) name1315 (
		_w2305_,
		_w2315_,
		_w2317_
	);
	LUT2 #(
		.INIT('h1)
	) name1316 (
		_w2316_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('h2)
	) name1317 (
		_w2314_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h4)
	) name1318 (
		_w2314_,
		_w2318_,
		_w2320_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		_w2283_,
		_w2286_,
		_w2321_
	);
	LUT2 #(
		.INIT('h2)
	) name1320 (
		_w2284_,
		_w2321_,
		_w2322_
	);
	LUT2 #(
		.INIT('h4)
	) name1321 (
		_w2284_,
		_w2321_,
		_w2323_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w2322_,
		_w2323_,
		_w2324_
	);
	LUT2 #(
		.INIT('h4)
	) name1323 (
		_w2320_,
		_w2324_,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name1324 (
		_w2319_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		_w2307_,
		_w2326_,
		_w2327_
	);
	LUT2 #(
		.INIT('h4)
	) name1326 (
		_w2307_,
		_w2326_,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		_w2327_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h8)
	) name1328 (
		_w2288_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		_w2288_,
		_w2329_,
		_w2331_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w2330_,
		_w2331_,
		_w2332_
	);
	LUT2 #(
		.INIT('h8)
	) name1331 (
		\A[862] ,
		\A[863] ,
		_w2333_
	);
	LUT2 #(
		.INIT('h8)
	) name1332 (
		\A[859] ,
		\A[860] ,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name1333 (
		\A[859] ,
		\A[860] ,
		_w2335_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		_w2334_,
		_w2335_,
		_w2336_
	);
	LUT2 #(
		.INIT('h8)
	) name1335 (
		\A[861] ,
		_w2336_,
		_w2337_
	);
	LUT2 #(
		.INIT('h1)
	) name1336 (
		\A[861] ,
		_w2336_,
		_w2338_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT2 #(
		.INIT('h1)
	) name1338 (
		\A[862] ,
		\A[863] ,
		_w2340_
	);
	LUT2 #(
		.INIT('h1)
	) name1339 (
		_w2333_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		\A[864] ,
		_w2341_,
		_w2342_
	);
	LUT2 #(
		.INIT('h1)
	) name1341 (
		\A[864] ,
		_w2341_,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w2342_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h8)
	) name1343 (
		_w2339_,
		_w2344_,
		_w2345_
	);
	LUT2 #(
		.INIT('h8)
	) name1344 (
		_w2333_,
		_w2345_,
		_w2346_
	);
	LUT2 #(
		.INIT('h1)
	) name1345 (
		_w2334_,
		_w2337_,
		_w2347_
	);
	LUT2 #(
		.INIT('h1)
	) name1346 (
		_w2333_,
		_w2342_,
		_w2348_
	);
	LUT2 #(
		.INIT('h4)
	) name1347 (
		_w2345_,
		_w2348_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name1348 (
		_w2347_,
		_w2349_,
		_w2350_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		_w2346_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h8)
	) name1350 (
		\A[868] ,
		\A[869] ,
		_w2352_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		\A[868] ,
		\A[869] ,
		_w2353_
	);
	LUT2 #(
		.INIT('h1)
	) name1352 (
		_w2352_,
		_w2353_,
		_w2354_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		\A[870] ,
		_w2354_,
		_w2355_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		_w2352_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h8)
	) name1355 (
		\A[865] ,
		\A[866] ,
		_w2357_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		\A[865] ,
		\A[866] ,
		_w2358_
	);
	LUT2 #(
		.INIT('h1)
	) name1357 (
		_w2357_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h8)
	) name1358 (
		\A[867] ,
		_w2359_,
		_w2360_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		_w2357_,
		_w2360_,
		_w2361_
	);
	LUT2 #(
		.INIT('h8)
	) name1360 (
		_w2356_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h1)
	) name1361 (
		_w2356_,
		_w2361_,
		_w2363_
	);
	LUT2 #(
		.INIT('h1)
	) name1362 (
		\A[867] ,
		_w2359_,
		_w2364_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		_w2360_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h1)
	) name1364 (
		\A[870] ,
		_w2354_,
		_w2366_
	);
	LUT2 #(
		.INIT('h1)
	) name1365 (
		_w2355_,
		_w2366_,
		_w2367_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		_w2365_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h1)
	) name1367 (
		_w2363_,
		_w2368_,
		_w2369_
	);
	LUT2 #(
		.INIT('h1)
	) name1368 (
		_w2362_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		_w2365_,
		_w2367_,
		_w2371_
	);
	LUT2 #(
		.INIT('h1)
	) name1370 (
		_w2368_,
		_w2371_,
		_w2372_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		_w2339_,
		_w2344_,
		_w2373_
	);
	LUT2 #(
		.INIT('h1)
	) name1372 (
		_w2345_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h8)
	) name1373 (
		_w2372_,
		_w2374_,
		_w2375_
	);
	LUT2 #(
		.INIT('h2)
	) name1374 (
		_w2346_,
		_w2347_,
		_w2376_
	);
	LUT2 #(
		.INIT('h2)
	) name1375 (
		_w2375_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		_w2362_,
		_w2363_,
		_w2378_
	);
	LUT2 #(
		.INIT('h2)
	) name1377 (
		_w2368_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h4)
	) name1378 (
		_w2368_,
		_w2378_,
		_w2380_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		_w2379_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h2)
	) name1380 (
		_w2377_,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h4)
	) name1381 (
		_w2377_,
		_w2381_,
		_w2383_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w2346_,
		_w2349_,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name1383 (
		_w2347_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h4)
	) name1384 (
		_w2347_,
		_w2384_,
		_w2386_
	);
	LUT2 #(
		.INIT('h1)
	) name1385 (
		_w2385_,
		_w2386_,
		_w2387_
	);
	LUT2 #(
		.INIT('h4)
	) name1386 (
		_w2383_,
		_w2387_,
		_w2388_
	);
	LUT2 #(
		.INIT('h1)
	) name1387 (
		_w2382_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name1388 (
		_w2370_,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h4)
	) name1389 (
		_w2370_,
		_w2389_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name1390 (
		_w2390_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h8)
	) name1391 (
		_w2351_,
		_w2392_,
		_w2393_
	);
	LUT2 #(
		.INIT('h1)
	) name1392 (
		_w2351_,
		_w2392_,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		_w2393_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h1)
	) name1394 (
		_w2332_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h8)
	) name1395 (
		_w2332_,
		_w2395_,
		_w2397_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		_w2372_,
		_w2374_,
		_w2398_
	);
	LUT2 #(
		.INIT('h1)
	) name1397 (
		_w2375_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w2309_,
		_w2311_,
		_w2400_
	);
	LUT2 #(
		.INIT('h1)
	) name1399 (
		_w2312_,
		_w2400_,
		_w2401_
	);
	LUT2 #(
		.INIT('h8)
	) name1400 (
		_w2399_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		_w2382_,
		_w2383_,
		_w2403_
	);
	LUT2 #(
		.INIT('h8)
	) name1402 (
		_w2387_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h1)
	) name1403 (
		_w2387_,
		_w2403_,
		_w2405_
	);
	LUT2 #(
		.INIT('h1)
	) name1404 (
		_w2404_,
		_w2405_,
		_w2406_
	);
	LUT2 #(
		.INIT('h8)
	) name1405 (
		_w2402_,
		_w2406_,
		_w2407_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		_w2402_,
		_w2406_,
		_w2408_
	);
	LUT2 #(
		.INIT('h1)
	) name1407 (
		_w2319_,
		_w2320_,
		_w2409_
	);
	LUT2 #(
		.INIT('h8)
	) name1408 (
		_w2324_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h1)
	) name1409 (
		_w2324_,
		_w2409_,
		_w2411_
	);
	LUT2 #(
		.INIT('h1)
	) name1410 (
		_w2410_,
		_w2411_,
		_w2412_
	);
	LUT2 #(
		.INIT('h4)
	) name1411 (
		_w2408_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		_w2407_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		_w2397_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		_w2396_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		_w2351_,
		_w2391_,
		_w2417_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		_w2390_,
		_w2417_,
		_w2418_
	);
	LUT2 #(
		.INIT('h1)
	) name1417 (
		_w2416_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h8)
	) name1418 (
		_w2416_,
		_w2418_,
		_w2420_
	);
	LUT2 #(
		.INIT('h1)
	) name1419 (
		_w2419_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h1)
	) name1420 (
		_w2288_,
		_w2328_,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name1421 (
		_w2327_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		_w2421_,
		_w2423_,
		_w2424_
	);
	LUT2 #(
		.INIT('h4)
	) name1423 (
		_w2421_,
		_w2423_,
		_w2425_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w2424_,
		_w2425_,
		_w2426_
	);
	LUT2 #(
		.INIT('h1)
	) name1425 (
		_w2269_,
		_w2426_,
		_w2427_
	);
	LUT2 #(
		.INIT('h8)
	) name1426 (
		_w2269_,
		_w2426_,
		_w2428_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w2396_,
		_w2397_,
		_w2429_
	);
	LUT2 #(
		.INIT('h4)
	) name1428 (
		_w2414_,
		_w2429_,
		_w2430_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		_w2414_,
		_w2429_,
		_w2431_
	);
	LUT2 #(
		.INIT('h1)
	) name1430 (
		_w2430_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h1)
	) name1431 (
		_w2237_,
		_w2238_,
		_w2433_
	);
	LUT2 #(
		.INIT('h4)
	) name1432 (
		_w2255_,
		_w2433_,
		_w2434_
	);
	LUT2 #(
		.INIT('h2)
	) name1433 (
		_w2255_,
		_w2433_,
		_w2435_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		_w2434_,
		_w2435_,
		_w2436_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w2432_,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h8)
	) name1436 (
		_w2432_,
		_w2436_,
		_w2438_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w2240_,
		_w2242_,
		_w2439_
	);
	LUT2 #(
		.INIT('h1)
	) name1438 (
		_w2243_,
		_w2439_,
		_w2440_
	);
	LUT2 #(
		.INIT('h1)
	) name1439 (
		_w2399_,
		_w2401_,
		_w2441_
	);
	LUT2 #(
		.INIT('h1)
	) name1440 (
		_w2402_,
		_w2441_,
		_w2442_
	);
	LUT2 #(
		.INIT('h8)
	) name1441 (
		_w2440_,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		_w2248_,
		_w2249_,
		_w2444_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		_w2253_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h2)
	) name1444 (
		_w2253_,
		_w2444_,
		_w2446_
	);
	LUT2 #(
		.INIT('h1)
	) name1445 (
		_w2445_,
		_w2446_,
		_w2447_
	);
	LUT2 #(
		.INIT('h2)
	) name1446 (
		_w2443_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('h4)
	) name1447 (
		_w2443_,
		_w2447_,
		_w2449_
	);
	LUT2 #(
		.INIT('h1)
	) name1448 (
		_w2407_,
		_w2408_,
		_w2450_
	);
	LUT2 #(
		.INIT('h4)
	) name1449 (
		_w2412_,
		_w2450_,
		_w2451_
	);
	LUT2 #(
		.INIT('h2)
	) name1450 (
		_w2412_,
		_w2450_,
		_w2452_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w2451_,
		_w2452_,
		_w2453_
	);
	LUT2 #(
		.INIT('h1)
	) name1452 (
		_w2449_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('h1)
	) name1453 (
		_w2448_,
		_w2454_,
		_w2455_
	);
	LUT2 #(
		.INIT('h4)
	) name1454 (
		_w2438_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h1)
	) name1455 (
		_w2437_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h1)
	) name1456 (
		_w2428_,
		_w2457_,
		_w2458_
	);
	LUT2 #(
		.INIT('h1)
	) name1457 (
		_w2427_,
		_w2458_,
		_w2459_
	);
	LUT2 #(
		.INIT('h2)
	) name1458 (
		_w2265_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h4)
	) name1459 (
		_w2265_,
		_w2459_,
		_w2461_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w2460_,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w2420_,
		_w2423_,
		_w2463_
	);
	LUT2 #(
		.INIT('h1)
	) name1462 (
		_w2419_,
		_w2463_,
		_w2464_
	);
	LUT2 #(
		.INIT('h8)
	) name1463 (
		_w2462_,
		_w2464_,
		_w2465_
	);
	LUT2 #(
		.INIT('h1)
	) name1464 (
		_w2462_,
		_w2464_,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name1465 (
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h8)
	) name1466 (
		\A[922] ,
		\A[923] ,
		_w2468_
	);
	LUT2 #(
		.INIT('h8)
	) name1467 (
		\A[919] ,
		\A[920] ,
		_w2469_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		\A[919] ,
		\A[920] ,
		_w2470_
	);
	LUT2 #(
		.INIT('h1)
	) name1469 (
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h8)
	) name1470 (
		\A[921] ,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h1)
	) name1471 (
		\A[921] ,
		_w2471_,
		_w2473_
	);
	LUT2 #(
		.INIT('h1)
	) name1472 (
		_w2472_,
		_w2473_,
		_w2474_
	);
	LUT2 #(
		.INIT('h1)
	) name1473 (
		\A[922] ,
		\A[923] ,
		_w2475_
	);
	LUT2 #(
		.INIT('h1)
	) name1474 (
		_w2468_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h8)
	) name1475 (
		\A[924] ,
		_w2476_,
		_w2477_
	);
	LUT2 #(
		.INIT('h1)
	) name1476 (
		\A[924] ,
		_w2476_,
		_w2478_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		_w2477_,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('h8)
	) name1478 (
		_w2474_,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h8)
	) name1479 (
		_w2468_,
		_w2480_,
		_w2481_
	);
	LUT2 #(
		.INIT('h1)
	) name1480 (
		_w2469_,
		_w2472_,
		_w2482_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		_w2468_,
		_w2477_,
		_w2483_
	);
	LUT2 #(
		.INIT('h4)
	) name1482 (
		_w2480_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h1)
	) name1483 (
		_w2482_,
		_w2484_,
		_w2485_
	);
	LUT2 #(
		.INIT('h1)
	) name1484 (
		_w2481_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h8)
	) name1485 (
		\A[928] ,
		\A[929] ,
		_w2487_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		\A[928] ,
		\A[929] ,
		_w2488_
	);
	LUT2 #(
		.INIT('h1)
	) name1487 (
		_w2487_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h8)
	) name1488 (
		\A[930] ,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		_w2487_,
		_w2490_,
		_w2491_
	);
	LUT2 #(
		.INIT('h8)
	) name1490 (
		\A[925] ,
		\A[926] ,
		_w2492_
	);
	LUT2 #(
		.INIT('h1)
	) name1491 (
		\A[925] ,
		\A[926] ,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name1492 (
		_w2492_,
		_w2493_,
		_w2494_
	);
	LUT2 #(
		.INIT('h8)
	) name1493 (
		\A[927] ,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h1)
	) name1494 (
		_w2492_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h8)
	) name1495 (
		_w2491_,
		_w2496_,
		_w2497_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		_w2491_,
		_w2496_,
		_w2498_
	);
	LUT2 #(
		.INIT('h1)
	) name1497 (
		\A[927] ,
		_w2494_,
		_w2499_
	);
	LUT2 #(
		.INIT('h1)
	) name1498 (
		_w2495_,
		_w2499_,
		_w2500_
	);
	LUT2 #(
		.INIT('h1)
	) name1499 (
		\A[930] ,
		_w2489_,
		_w2501_
	);
	LUT2 #(
		.INIT('h1)
	) name1500 (
		_w2490_,
		_w2501_,
		_w2502_
	);
	LUT2 #(
		.INIT('h8)
	) name1501 (
		_w2500_,
		_w2502_,
		_w2503_
	);
	LUT2 #(
		.INIT('h1)
	) name1502 (
		_w2498_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w2497_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h1)
	) name1504 (
		_w2500_,
		_w2502_,
		_w2506_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		_w2503_,
		_w2506_,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name1506 (
		_w2474_,
		_w2479_,
		_w2508_
	);
	LUT2 #(
		.INIT('h1)
	) name1507 (
		_w2480_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h8)
	) name1508 (
		_w2507_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name1509 (
		_w2481_,
		_w2482_,
		_w2511_
	);
	LUT2 #(
		.INIT('h2)
	) name1510 (
		_w2510_,
		_w2511_,
		_w2512_
	);
	LUT2 #(
		.INIT('h1)
	) name1511 (
		_w2497_,
		_w2498_,
		_w2513_
	);
	LUT2 #(
		.INIT('h2)
	) name1512 (
		_w2503_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h4)
	) name1513 (
		_w2503_,
		_w2513_,
		_w2515_
	);
	LUT2 #(
		.INIT('h1)
	) name1514 (
		_w2514_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h2)
	) name1515 (
		_w2512_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h4)
	) name1516 (
		_w2512_,
		_w2516_,
		_w2518_
	);
	LUT2 #(
		.INIT('h1)
	) name1517 (
		_w2481_,
		_w2484_,
		_w2519_
	);
	LUT2 #(
		.INIT('h2)
	) name1518 (
		_w2482_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h4)
	) name1519 (
		_w2482_,
		_w2519_,
		_w2521_
	);
	LUT2 #(
		.INIT('h1)
	) name1520 (
		_w2520_,
		_w2521_,
		_w2522_
	);
	LUT2 #(
		.INIT('h4)
	) name1521 (
		_w2518_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h1)
	) name1522 (
		_w2517_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h2)
	) name1523 (
		_w2505_,
		_w2524_,
		_w2525_
	);
	LUT2 #(
		.INIT('h4)
	) name1524 (
		_w2505_,
		_w2524_,
		_w2526_
	);
	LUT2 #(
		.INIT('h1)
	) name1525 (
		_w2525_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h8)
	) name1526 (
		_w2486_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h1)
	) name1527 (
		_w2486_,
		_w2527_,
		_w2529_
	);
	LUT2 #(
		.INIT('h1)
	) name1528 (
		_w2528_,
		_w2529_,
		_w2530_
	);
	LUT2 #(
		.INIT('h8)
	) name1529 (
		\A[934] ,
		\A[935] ,
		_w2531_
	);
	LUT2 #(
		.INIT('h8)
	) name1530 (
		\A[931] ,
		\A[932] ,
		_w2532_
	);
	LUT2 #(
		.INIT('h1)
	) name1531 (
		\A[931] ,
		\A[932] ,
		_w2533_
	);
	LUT2 #(
		.INIT('h1)
	) name1532 (
		_w2532_,
		_w2533_,
		_w2534_
	);
	LUT2 #(
		.INIT('h8)
	) name1533 (
		\A[933] ,
		_w2534_,
		_w2535_
	);
	LUT2 #(
		.INIT('h1)
	) name1534 (
		\A[933] ,
		_w2534_,
		_w2536_
	);
	LUT2 #(
		.INIT('h1)
	) name1535 (
		_w2535_,
		_w2536_,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name1536 (
		\A[934] ,
		\A[935] ,
		_w2538_
	);
	LUT2 #(
		.INIT('h1)
	) name1537 (
		_w2531_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h8)
	) name1538 (
		\A[936] ,
		_w2539_,
		_w2540_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		\A[936] ,
		_w2539_,
		_w2541_
	);
	LUT2 #(
		.INIT('h1)
	) name1540 (
		_w2540_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h8)
	) name1541 (
		_w2537_,
		_w2542_,
		_w2543_
	);
	LUT2 #(
		.INIT('h8)
	) name1542 (
		_w2531_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h1)
	) name1543 (
		_w2532_,
		_w2535_,
		_w2545_
	);
	LUT2 #(
		.INIT('h1)
	) name1544 (
		_w2531_,
		_w2540_,
		_w2546_
	);
	LUT2 #(
		.INIT('h4)
	) name1545 (
		_w2543_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h1)
	) name1546 (
		_w2545_,
		_w2547_,
		_w2548_
	);
	LUT2 #(
		.INIT('h1)
	) name1547 (
		_w2544_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h8)
	) name1548 (
		\A[940] ,
		\A[941] ,
		_w2550_
	);
	LUT2 #(
		.INIT('h1)
	) name1549 (
		\A[940] ,
		\A[941] ,
		_w2551_
	);
	LUT2 #(
		.INIT('h1)
	) name1550 (
		_w2550_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h8)
	) name1551 (
		\A[942] ,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h1)
	) name1552 (
		_w2550_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h8)
	) name1553 (
		\A[937] ,
		\A[938] ,
		_w2555_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		\A[937] ,
		\A[938] ,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name1555 (
		_w2555_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h8)
	) name1556 (
		\A[939] ,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('h1)
	) name1557 (
		_w2555_,
		_w2558_,
		_w2559_
	);
	LUT2 #(
		.INIT('h8)
	) name1558 (
		_w2554_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h1)
	) name1559 (
		_w2554_,
		_w2559_,
		_w2561_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		\A[939] ,
		_w2557_,
		_w2562_
	);
	LUT2 #(
		.INIT('h1)
	) name1561 (
		_w2558_,
		_w2562_,
		_w2563_
	);
	LUT2 #(
		.INIT('h1)
	) name1562 (
		\A[942] ,
		_w2552_,
		_w2564_
	);
	LUT2 #(
		.INIT('h1)
	) name1563 (
		_w2553_,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('h8)
	) name1564 (
		_w2563_,
		_w2565_,
		_w2566_
	);
	LUT2 #(
		.INIT('h1)
	) name1565 (
		_w2561_,
		_w2566_,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name1566 (
		_w2560_,
		_w2567_,
		_w2568_
	);
	LUT2 #(
		.INIT('h1)
	) name1567 (
		_w2563_,
		_w2565_,
		_w2569_
	);
	LUT2 #(
		.INIT('h1)
	) name1568 (
		_w2566_,
		_w2569_,
		_w2570_
	);
	LUT2 #(
		.INIT('h1)
	) name1569 (
		_w2537_,
		_w2542_,
		_w2571_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		_w2543_,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('h8)
	) name1571 (
		_w2570_,
		_w2572_,
		_w2573_
	);
	LUT2 #(
		.INIT('h2)
	) name1572 (
		_w2544_,
		_w2545_,
		_w2574_
	);
	LUT2 #(
		.INIT('h2)
	) name1573 (
		_w2573_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		_w2560_,
		_w2561_,
		_w2576_
	);
	LUT2 #(
		.INIT('h2)
	) name1575 (
		_w2566_,
		_w2576_,
		_w2577_
	);
	LUT2 #(
		.INIT('h4)
	) name1576 (
		_w2566_,
		_w2576_,
		_w2578_
	);
	LUT2 #(
		.INIT('h1)
	) name1577 (
		_w2577_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h2)
	) name1578 (
		_w2575_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h4)
	) name1579 (
		_w2575_,
		_w2579_,
		_w2581_
	);
	LUT2 #(
		.INIT('h1)
	) name1580 (
		_w2544_,
		_w2547_,
		_w2582_
	);
	LUT2 #(
		.INIT('h2)
	) name1581 (
		_w2545_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h4)
	) name1582 (
		_w2545_,
		_w2582_,
		_w2584_
	);
	LUT2 #(
		.INIT('h1)
	) name1583 (
		_w2583_,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h4)
	) name1584 (
		_w2581_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		_w2580_,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h2)
	) name1586 (
		_w2568_,
		_w2587_,
		_w2588_
	);
	LUT2 #(
		.INIT('h4)
	) name1587 (
		_w2568_,
		_w2587_,
		_w2589_
	);
	LUT2 #(
		.INIT('h1)
	) name1588 (
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h8)
	) name1589 (
		_w2549_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w2549_,
		_w2590_,
		_w2592_
	);
	LUT2 #(
		.INIT('h1)
	) name1591 (
		_w2591_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h1)
	) name1592 (
		_w2530_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h8)
	) name1593 (
		_w2530_,
		_w2593_,
		_w2595_
	);
	LUT2 #(
		.INIT('h1)
	) name1594 (
		_w2570_,
		_w2572_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name1595 (
		_w2573_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h1)
	) name1596 (
		_w2507_,
		_w2509_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name1597 (
		_w2510_,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h8)
	) name1598 (
		_w2597_,
		_w2599_,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name1599 (
		_w2580_,
		_w2581_,
		_w2601_
	);
	LUT2 #(
		.INIT('h8)
	) name1600 (
		_w2585_,
		_w2601_,
		_w2602_
	);
	LUT2 #(
		.INIT('h1)
	) name1601 (
		_w2585_,
		_w2601_,
		_w2603_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w2602_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h8)
	) name1603 (
		_w2600_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h1)
	) name1604 (
		_w2600_,
		_w2604_,
		_w2606_
	);
	LUT2 #(
		.INIT('h1)
	) name1605 (
		_w2517_,
		_w2518_,
		_w2607_
	);
	LUT2 #(
		.INIT('h8)
	) name1606 (
		_w2522_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w2522_,
		_w2607_,
		_w2609_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w2608_,
		_w2609_,
		_w2610_
	);
	LUT2 #(
		.INIT('h4)
	) name1609 (
		_w2606_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w2605_,
		_w2611_,
		_w2612_
	);
	LUT2 #(
		.INIT('h1)
	) name1611 (
		_w2595_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h1)
	) name1612 (
		_w2594_,
		_w2613_,
		_w2614_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w2549_,
		_w2589_,
		_w2615_
	);
	LUT2 #(
		.INIT('h1)
	) name1614 (
		_w2588_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h1)
	) name1615 (
		_w2614_,
		_w2616_,
		_w2617_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		_w2614_,
		_w2616_,
		_w2618_
	);
	LUT2 #(
		.INIT('h1)
	) name1617 (
		_w2486_,
		_w2526_,
		_w2619_
	);
	LUT2 #(
		.INIT('h1)
	) name1618 (
		_w2525_,
		_w2619_,
		_w2620_
	);
	LUT2 #(
		.INIT('h1)
	) name1619 (
		_w2618_,
		_w2620_,
		_w2621_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w2617_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h1)
	) name1621 (
		_w2617_,
		_w2618_,
		_w2623_
	);
	LUT2 #(
		.INIT('h4)
	) name1622 (
		_w2620_,
		_w2623_,
		_w2624_
	);
	LUT2 #(
		.INIT('h2)
	) name1623 (
		_w2620_,
		_w2623_,
		_w2625_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w2624_,
		_w2625_,
		_w2626_
	);
	LUT2 #(
		.INIT('h8)
	) name1625 (
		\A[898] ,
		\A[899] ,
		_w2627_
	);
	LUT2 #(
		.INIT('h8)
	) name1626 (
		\A[895] ,
		\A[896] ,
		_w2628_
	);
	LUT2 #(
		.INIT('h1)
	) name1627 (
		\A[895] ,
		\A[896] ,
		_w2629_
	);
	LUT2 #(
		.INIT('h1)
	) name1628 (
		_w2628_,
		_w2629_,
		_w2630_
	);
	LUT2 #(
		.INIT('h8)
	) name1629 (
		\A[897] ,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h1)
	) name1630 (
		\A[897] ,
		_w2630_,
		_w2632_
	);
	LUT2 #(
		.INIT('h1)
	) name1631 (
		_w2631_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		\A[898] ,
		\A[899] ,
		_w2634_
	);
	LUT2 #(
		.INIT('h1)
	) name1633 (
		_w2627_,
		_w2634_,
		_w2635_
	);
	LUT2 #(
		.INIT('h8)
	) name1634 (
		\A[900] ,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h1)
	) name1635 (
		\A[900] ,
		_w2635_,
		_w2637_
	);
	LUT2 #(
		.INIT('h1)
	) name1636 (
		_w2636_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h8)
	) name1637 (
		_w2633_,
		_w2638_,
		_w2639_
	);
	LUT2 #(
		.INIT('h8)
	) name1638 (
		_w2627_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		_w2628_,
		_w2631_,
		_w2641_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		_w2627_,
		_w2636_,
		_w2642_
	);
	LUT2 #(
		.INIT('h4)
	) name1641 (
		_w2639_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		_w2641_,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h1)
	) name1643 (
		_w2640_,
		_w2644_,
		_w2645_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		\A[904] ,
		\A[905] ,
		_w2646_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		\A[904] ,
		\A[905] ,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name1646 (
		_w2646_,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h8)
	) name1647 (
		\A[906] ,
		_w2648_,
		_w2649_
	);
	LUT2 #(
		.INIT('h1)
	) name1648 (
		_w2646_,
		_w2649_,
		_w2650_
	);
	LUT2 #(
		.INIT('h8)
	) name1649 (
		\A[901] ,
		\A[902] ,
		_w2651_
	);
	LUT2 #(
		.INIT('h1)
	) name1650 (
		\A[901] ,
		\A[902] ,
		_w2652_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		\A[903] ,
		_w2653_,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name1653 (
		_w2651_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h8)
	) name1654 (
		_w2650_,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h1)
	) name1655 (
		_w2650_,
		_w2655_,
		_w2657_
	);
	LUT2 #(
		.INIT('h1)
	) name1656 (
		\A[903] ,
		_w2653_,
		_w2658_
	);
	LUT2 #(
		.INIT('h1)
	) name1657 (
		_w2654_,
		_w2658_,
		_w2659_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		\A[906] ,
		_w2648_,
		_w2660_
	);
	LUT2 #(
		.INIT('h1)
	) name1659 (
		_w2649_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		_w2659_,
		_w2661_,
		_w2662_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		_w2657_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		_w2656_,
		_w2663_,
		_w2664_
	);
	LUT2 #(
		.INIT('h1)
	) name1663 (
		_w2659_,
		_w2661_,
		_w2665_
	);
	LUT2 #(
		.INIT('h1)
	) name1664 (
		_w2662_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		_w2633_,
		_w2638_,
		_w2667_
	);
	LUT2 #(
		.INIT('h1)
	) name1666 (
		_w2639_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h8)
	) name1667 (
		_w2666_,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('h2)
	) name1668 (
		_w2640_,
		_w2641_,
		_w2670_
	);
	LUT2 #(
		.INIT('h2)
	) name1669 (
		_w2669_,
		_w2670_,
		_w2671_
	);
	LUT2 #(
		.INIT('h1)
	) name1670 (
		_w2656_,
		_w2657_,
		_w2672_
	);
	LUT2 #(
		.INIT('h2)
	) name1671 (
		_w2662_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h4)
	) name1672 (
		_w2662_,
		_w2672_,
		_w2674_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		_w2673_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h2)
	) name1674 (
		_w2671_,
		_w2675_,
		_w2676_
	);
	LUT2 #(
		.INIT('h4)
	) name1675 (
		_w2671_,
		_w2675_,
		_w2677_
	);
	LUT2 #(
		.INIT('h1)
	) name1676 (
		_w2640_,
		_w2643_,
		_w2678_
	);
	LUT2 #(
		.INIT('h2)
	) name1677 (
		_w2641_,
		_w2678_,
		_w2679_
	);
	LUT2 #(
		.INIT('h4)
	) name1678 (
		_w2641_,
		_w2678_,
		_w2680_
	);
	LUT2 #(
		.INIT('h1)
	) name1679 (
		_w2679_,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('h4)
	) name1680 (
		_w2677_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h1)
	) name1681 (
		_w2676_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h2)
	) name1682 (
		_w2664_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h4)
	) name1683 (
		_w2664_,
		_w2683_,
		_w2685_
	);
	LUT2 #(
		.INIT('h1)
	) name1684 (
		_w2684_,
		_w2685_,
		_w2686_
	);
	LUT2 #(
		.INIT('h8)
	) name1685 (
		_w2645_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h1)
	) name1686 (
		_w2645_,
		_w2686_,
		_w2688_
	);
	LUT2 #(
		.INIT('h1)
	) name1687 (
		_w2687_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		\A[910] ,
		\A[911] ,
		_w2690_
	);
	LUT2 #(
		.INIT('h8)
	) name1689 (
		\A[907] ,
		\A[908] ,
		_w2691_
	);
	LUT2 #(
		.INIT('h1)
	) name1690 (
		\A[907] ,
		\A[908] ,
		_w2692_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w2691_,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h8)
	) name1692 (
		\A[909] ,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('h1)
	) name1693 (
		\A[909] ,
		_w2693_,
		_w2695_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w2694_,
		_w2695_,
		_w2696_
	);
	LUT2 #(
		.INIT('h1)
	) name1695 (
		\A[910] ,
		\A[911] ,
		_w2697_
	);
	LUT2 #(
		.INIT('h1)
	) name1696 (
		_w2690_,
		_w2697_,
		_w2698_
	);
	LUT2 #(
		.INIT('h8)
	) name1697 (
		\A[912] ,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h1)
	) name1698 (
		\A[912] ,
		_w2698_,
		_w2700_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name1700 (
		_w2696_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		_w2690_,
		_w2702_,
		_w2703_
	);
	LUT2 #(
		.INIT('h1)
	) name1702 (
		_w2691_,
		_w2694_,
		_w2704_
	);
	LUT2 #(
		.INIT('h1)
	) name1703 (
		_w2690_,
		_w2699_,
		_w2705_
	);
	LUT2 #(
		.INIT('h4)
	) name1704 (
		_w2702_,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('h1)
	) name1705 (
		_w2704_,
		_w2706_,
		_w2707_
	);
	LUT2 #(
		.INIT('h1)
	) name1706 (
		_w2703_,
		_w2707_,
		_w2708_
	);
	LUT2 #(
		.INIT('h8)
	) name1707 (
		\A[916] ,
		\A[917] ,
		_w2709_
	);
	LUT2 #(
		.INIT('h1)
	) name1708 (
		\A[916] ,
		\A[917] ,
		_w2710_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w2709_,
		_w2710_,
		_w2711_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		\A[918] ,
		_w2711_,
		_w2712_
	);
	LUT2 #(
		.INIT('h1)
	) name1711 (
		_w2709_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h8)
	) name1712 (
		\A[913] ,
		\A[914] ,
		_w2714_
	);
	LUT2 #(
		.INIT('h1)
	) name1713 (
		\A[913] ,
		\A[914] ,
		_w2715_
	);
	LUT2 #(
		.INIT('h1)
	) name1714 (
		_w2714_,
		_w2715_,
		_w2716_
	);
	LUT2 #(
		.INIT('h8)
	) name1715 (
		\A[915] ,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h1)
	) name1716 (
		_w2714_,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h8)
	) name1717 (
		_w2713_,
		_w2718_,
		_w2719_
	);
	LUT2 #(
		.INIT('h1)
	) name1718 (
		_w2713_,
		_w2718_,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name1719 (
		\A[915] ,
		_w2716_,
		_w2721_
	);
	LUT2 #(
		.INIT('h1)
	) name1720 (
		_w2717_,
		_w2721_,
		_w2722_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		\A[918] ,
		_w2711_,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w2712_,
		_w2723_,
		_w2724_
	);
	LUT2 #(
		.INIT('h8)
	) name1723 (
		_w2722_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h1)
	) name1724 (
		_w2720_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h1)
	) name1725 (
		_w2719_,
		_w2726_,
		_w2727_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		_w2722_,
		_w2724_,
		_w2728_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w2725_,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h1)
	) name1728 (
		_w2696_,
		_w2701_,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name1729 (
		_w2702_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h8)
	) name1730 (
		_w2729_,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h2)
	) name1731 (
		_w2703_,
		_w2704_,
		_w2733_
	);
	LUT2 #(
		.INIT('h2)
	) name1732 (
		_w2732_,
		_w2733_,
		_w2734_
	);
	LUT2 #(
		.INIT('h1)
	) name1733 (
		_w2719_,
		_w2720_,
		_w2735_
	);
	LUT2 #(
		.INIT('h2)
	) name1734 (
		_w2725_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h4)
	) name1735 (
		_w2725_,
		_w2735_,
		_w2737_
	);
	LUT2 #(
		.INIT('h1)
	) name1736 (
		_w2736_,
		_w2737_,
		_w2738_
	);
	LUT2 #(
		.INIT('h2)
	) name1737 (
		_w2734_,
		_w2738_,
		_w2739_
	);
	LUT2 #(
		.INIT('h4)
	) name1738 (
		_w2734_,
		_w2738_,
		_w2740_
	);
	LUT2 #(
		.INIT('h1)
	) name1739 (
		_w2703_,
		_w2706_,
		_w2741_
	);
	LUT2 #(
		.INIT('h2)
	) name1740 (
		_w2704_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h4)
	) name1741 (
		_w2704_,
		_w2741_,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name1742 (
		_w2742_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h4)
	) name1743 (
		_w2740_,
		_w2744_,
		_w2745_
	);
	LUT2 #(
		.INIT('h1)
	) name1744 (
		_w2739_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h2)
	) name1745 (
		_w2727_,
		_w2746_,
		_w2747_
	);
	LUT2 #(
		.INIT('h4)
	) name1746 (
		_w2727_,
		_w2746_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name1747 (
		_w2747_,
		_w2748_,
		_w2749_
	);
	LUT2 #(
		.INIT('h8)
	) name1748 (
		_w2708_,
		_w2749_,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		_w2708_,
		_w2749_,
		_w2751_
	);
	LUT2 #(
		.INIT('h1)
	) name1750 (
		_w2750_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h1)
	) name1751 (
		_w2689_,
		_w2752_,
		_w2753_
	);
	LUT2 #(
		.INIT('h8)
	) name1752 (
		_w2689_,
		_w2752_,
		_w2754_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		_w2729_,
		_w2731_,
		_w2755_
	);
	LUT2 #(
		.INIT('h1)
	) name1754 (
		_w2732_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h1)
	) name1755 (
		_w2666_,
		_w2668_,
		_w2757_
	);
	LUT2 #(
		.INIT('h1)
	) name1756 (
		_w2669_,
		_w2757_,
		_w2758_
	);
	LUT2 #(
		.INIT('h8)
	) name1757 (
		_w2756_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h1)
	) name1758 (
		_w2739_,
		_w2740_,
		_w2760_
	);
	LUT2 #(
		.INIT('h8)
	) name1759 (
		_w2744_,
		_w2760_,
		_w2761_
	);
	LUT2 #(
		.INIT('h1)
	) name1760 (
		_w2744_,
		_w2760_,
		_w2762_
	);
	LUT2 #(
		.INIT('h1)
	) name1761 (
		_w2761_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		_w2759_,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		_w2759_,
		_w2763_,
		_w2765_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		_w2676_,
		_w2677_,
		_w2766_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		_w2681_,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h1)
	) name1766 (
		_w2681_,
		_w2766_,
		_w2768_
	);
	LUT2 #(
		.INIT('h1)
	) name1767 (
		_w2767_,
		_w2768_,
		_w2769_
	);
	LUT2 #(
		.INIT('h4)
	) name1768 (
		_w2765_,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		_w2764_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		_w2754_,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h1)
	) name1771 (
		_w2753_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name1772 (
		_w2708_,
		_w2748_,
		_w2774_
	);
	LUT2 #(
		.INIT('h1)
	) name1773 (
		_w2747_,
		_w2774_,
		_w2775_
	);
	LUT2 #(
		.INIT('h1)
	) name1774 (
		_w2773_,
		_w2775_,
		_w2776_
	);
	LUT2 #(
		.INIT('h8)
	) name1775 (
		_w2773_,
		_w2775_,
		_w2777_
	);
	LUT2 #(
		.INIT('h1)
	) name1776 (
		_w2776_,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h1)
	) name1777 (
		_w2645_,
		_w2685_,
		_w2779_
	);
	LUT2 #(
		.INIT('h1)
	) name1778 (
		_w2684_,
		_w2779_,
		_w2780_
	);
	LUT2 #(
		.INIT('h2)
	) name1779 (
		_w2778_,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h4)
	) name1780 (
		_w2778_,
		_w2780_,
		_w2782_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w2781_,
		_w2782_,
		_w2783_
	);
	LUT2 #(
		.INIT('h1)
	) name1782 (
		_w2626_,
		_w2783_,
		_w2784_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		_w2626_,
		_w2783_,
		_w2785_
	);
	LUT2 #(
		.INIT('h1)
	) name1784 (
		_w2753_,
		_w2754_,
		_w2786_
	);
	LUT2 #(
		.INIT('h4)
	) name1785 (
		_w2771_,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h2)
	) name1786 (
		_w2771_,
		_w2786_,
		_w2788_
	);
	LUT2 #(
		.INIT('h1)
	) name1787 (
		_w2787_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w2594_,
		_w2595_,
		_w2790_
	);
	LUT2 #(
		.INIT('h4)
	) name1789 (
		_w2612_,
		_w2790_,
		_w2791_
	);
	LUT2 #(
		.INIT('h2)
	) name1790 (
		_w2612_,
		_w2790_,
		_w2792_
	);
	LUT2 #(
		.INIT('h1)
	) name1791 (
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name1792 (
		_w2789_,
		_w2793_,
		_w2794_
	);
	LUT2 #(
		.INIT('h8)
	) name1793 (
		_w2789_,
		_w2793_,
		_w2795_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		_w2597_,
		_w2599_,
		_w2796_
	);
	LUT2 #(
		.INIT('h1)
	) name1795 (
		_w2600_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w2756_,
		_w2758_,
		_w2798_
	);
	LUT2 #(
		.INIT('h1)
	) name1797 (
		_w2759_,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h8)
	) name1798 (
		_w2797_,
		_w2799_,
		_w2800_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		_w2605_,
		_w2606_,
		_w2801_
	);
	LUT2 #(
		.INIT('h4)
	) name1800 (
		_w2610_,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h2)
	) name1801 (
		_w2610_,
		_w2801_,
		_w2803_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		_w2802_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		_w2800_,
		_w2804_,
		_w2805_
	);
	LUT2 #(
		.INIT('h4)
	) name1804 (
		_w2800_,
		_w2804_,
		_w2806_
	);
	LUT2 #(
		.INIT('h1)
	) name1805 (
		_w2764_,
		_w2765_,
		_w2807_
	);
	LUT2 #(
		.INIT('h4)
	) name1806 (
		_w2769_,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		_w2769_,
		_w2807_,
		_w2809_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w2808_,
		_w2809_,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name1809 (
		_w2806_,
		_w2810_,
		_w2811_
	);
	LUT2 #(
		.INIT('h1)
	) name1810 (
		_w2805_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		_w2795_,
		_w2812_,
		_w2813_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w2794_,
		_w2813_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name1813 (
		_w2785_,
		_w2814_,
		_w2815_
	);
	LUT2 #(
		.INIT('h1)
	) name1814 (
		_w2784_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		_w2622_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h4)
	) name1816 (
		_w2622_,
		_w2816_,
		_w2818_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w2817_,
		_w2818_,
		_w2819_
	);
	LUT2 #(
		.INIT('h1)
	) name1818 (
		_w2777_,
		_w2780_,
		_w2820_
	);
	LUT2 #(
		.INIT('h1)
	) name1819 (
		_w2776_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('h8)
	) name1820 (
		_w2819_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h1)
	) name1821 (
		_w2819_,
		_w2821_,
		_w2823_
	);
	LUT2 #(
		.INIT('h1)
	) name1822 (
		_w2822_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h1)
	) name1823 (
		_w2467_,
		_w2824_,
		_w2825_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		_w2467_,
		_w2824_,
		_w2826_
	);
	LUT2 #(
		.INIT('h1)
	) name1825 (
		_w2784_,
		_w2785_,
		_w2827_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		_w2814_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h2)
	) name1827 (
		_w2814_,
		_w2827_,
		_w2829_
	);
	LUT2 #(
		.INIT('h1)
	) name1828 (
		_w2828_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h1)
	) name1829 (
		_w2427_,
		_w2428_,
		_w2831_
	);
	LUT2 #(
		.INIT('h4)
	) name1830 (
		_w2457_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h2)
	) name1831 (
		_w2457_,
		_w2831_,
		_w2833_
	);
	LUT2 #(
		.INIT('h1)
	) name1832 (
		_w2832_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h1)
	) name1833 (
		_w2830_,
		_w2834_,
		_w2835_
	);
	LUT2 #(
		.INIT('h8)
	) name1834 (
		_w2830_,
		_w2834_,
		_w2836_
	);
	LUT2 #(
		.INIT('h1)
	) name1835 (
		_w2437_,
		_w2438_,
		_w2837_
	);
	LUT2 #(
		.INIT('h4)
	) name1836 (
		_w2455_,
		_w2837_,
		_w2838_
	);
	LUT2 #(
		.INIT('h2)
	) name1837 (
		_w2455_,
		_w2837_,
		_w2839_
	);
	LUT2 #(
		.INIT('h1)
	) name1838 (
		_w2838_,
		_w2839_,
		_w2840_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w2794_,
		_w2795_,
		_w2841_
	);
	LUT2 #(
		.INIT('h4)
	) name1840 (
		_w2812_,
		_w2841_,
		_w2842_
	);
	LUT2 #(
		.INIT('h2)
	) name1841 (
		_w2812_,
		_w2841_,
		_w2843_
	);
	LUT2 #(
		.INIT('h1)
	) name1842 (
		_w2842_,
		_w2843_,
		_w2844_
	);
	LUT2 #(
		.INIT('h1)
	) name1843 (
		_w2840_,
		_w2844_,
		_w2845_
	);
	LUT2 #(
		.INIT('h8)
	) name1844 (
		_w2840_,
		_w2844_,
		_w2846_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		_w2797_,
		_w2799_,
		_w2847_
	);
	LUT2 #(
		.INIT('h1)
	) name1846 (
		_w2800_,
		_w2847_,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		_w2440_,
		_w2442_,
		_w2849_
	);
	LUT2 #(
		.INIT('h1)
	) name1848 (
		_w2443_,
		_w2849_,
		_w2850_
	);
	LUT2 #(
		.INIT('h8)
	) name1849 (
		_w2848_,
		_w2850_,
		_w2851_
	);
	LUT2 #(
		.INIT('h1)
	) name1850 (
		_w2805_,
		_w2806_,
		_w2852_
	);
	LUT2 #(
		.INIT('h4)
	) name1851 (
		_w2810_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name1852 (
		_w2810_,
		_w2852_,
		_w2854_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w2853_,
		_w2854_,
		_w2855_
	);
	LUT2 #(
		.INIT('h8)
	) name1854 (
		_w2851_,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('h1)
	) name1855 (
		_w2851_,
		_w2855_,
		_w2857_
	);
	LUT2 #(
		.INIT('h1)
	) name1856 (
		_w2448_,
		_w2449_,
		_w2858_
	);
	LUT2 #(
		.INIT('h4)
	) name1857 (
		_w2453_,
		_w2858_,
		_w2859_
	);
	LUT2 #(
		.INIT('h2)
	) name1858 (
		_w2453_,
		_w2858_,
		_w2860_
	);
	LUT2 #(
		.INIT('h1)
	) name1859 (
		_w2859_,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h4)
	) name1860 (
		_w2857_,
		_w2861_,
		_w2862_
	);
	LUT2 #(
		.INIT('h1)
	) name1861 (
		_w2856_,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('h4)
	) name1862 (
		_w2846_,
		_w2863_,
		_w2864_
	);
	LUT2 #(
		.INIT('h1)
	) name1863 (
		_w2845_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h4)
	) name1864 (
		_w2836_,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h1)
	) name1865 (
		_w2835_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h1)
	) name1866 (
		_w2826_,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h1)
	) name1867 (
		_w2825_,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h4)
	) name1868 (
		_w2818_,
		_w2821_,
		_w2870_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w2817_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h2)
	) name1870 (
		_w2869_,
		_w2871_,
		_w2872_
	);
	LUT2 #(
		.INIT('h4)
	) name1871 (
		_w2869_,
		_w2871_,
		_w2873_
	);
	LUT2 #(
		.INIT('h4)
	) name1872 (
		_w2461_,
		_w2464_,
		_w2874_
	);
	LUT2 #(
		.INIT('h1)
	) name1873 (
		_w2460_,
		_w2874_,
		_w2875_
	);
	LUT2 #(
		.INIT('h1)
	) name1874 (
		_w2873_,
		_w2875_,
		_w2876_
	);
	LUT2 #(
		.INIT('h1)
	) name1875 (
		_w2872_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		_w2110_,
		_w2877_,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w2049_,
		_w2050_,
		_w2879_
	);
	LUT2 #(
		.INIT('h8)
	) name1878 (
		_w2103_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h1)
	) name1879 (
		_w2103_,
		_w2879_,
		_w2881_
	);
	LUT2 #(
		.INIT('h1)
	) name1880 (
		_w2880_,
		_w2881_,
		_w2882_
	);
	LUT2 #(
		.INIT('h1)
	) name1881 (
		_w2872_,
		_w2873_,
		_w2883_
	);
	LUT2 #(
		.INIT('h8)
	) name1882 (
		_w2875_,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h1)
	) name1883 (
		_w2875_,
		_w2883_,
		_w2885_
	);
	LUT2 #(
		.INIT('h1)
	) name1884 (
		_w2884_,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h1)
	) name1885 (
		_w2882_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h8)
	) name1886 (
		_w2882_,
		_w2886_,
		_w2888_
	);
	LUT2 #(
		.INIT('h1)
	) name1887 (
		_w2825_,
		_w2826_,
		_w2889_
	);
	LUT2 #(
		.INIT('h4)
	) name1888 (
		_w2867_,
		_w2889_,
		_w2890_
	);
	LUT2 #(
		.INIT('h2)
	) name1889 (
		_w2867_,
		_w2889_,
		_w2891_
	);
	LUT2 #(
		.INIT('h1)
	) name1890 (
		_w2890_,
		_w2891_,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name1891 (
		_w2059_,
		_w2060_,
		_w2893_
	);
	LUT2 #(
		.INIT('h4)
	) name1892 (
		_w2101_,
		_w2893_,
		_w2894_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		_w2101_,
		_w2893_,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name1894 (
		_w2894_,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h4)
	) name1895 (
		_w2892_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h2)
	) name1896 (
		_w2892_,
		_w2896_,
		_w2898_
	);
	LUT2 #(
		.INIT('h1)
	) name1897 (
		_w2069_,
		_w2070_,
		_w2899_
	);
	LUT2 #(
		.INIT('h4)
	) name1898 (
		_w2099_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('h2)
	) name1899 (
		_w2099_,
		_w2899_,
		_w2901_
	);
	LUT2 #(
		.INIT('h1)
	) name1900 (
		_w2900_,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w2835_,
		_w2836_,
		_w2903_
	);
	LUT2 #(
		.INIT('h8)
	) name1902 (
		_w2865_,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		_w2865_,
		_w2903_,
		_w2905_
	);
	LUT2 #(
		.INIT('h1)
	) name1904 (
		_w2904_,
		_w2905_,
		_w2906_
	);
	LUT2 #(
		.INIT('h2)
	) name1905 (
		_w2902_,
		_w2906_,
		_w2907_
	);
	LUT2 #(
		.INIT('h4)
	) name1906 (
		_w2902_,
		_w2906_,
		_w2908_
	);
	LUT2 #(
		.INIT('h1)
	) name1907 (
		_w2845_,
		_w2846_,
		_w2909_
	);
	LUT2 #(
		.INIT('h4)
	) name1908 (
		_w2863_,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h2)
	) name1909 (
		_w2863_,
		_w2909_,
		_w2911_
	);
	LUT2 #(
		.INIT('h1)
	) name1910 (
		_w2910_,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h1)
	) name1911 (
		_w2079_,
		_w2080_,
		_w2913_
	);
	LUT2 #(
		.INIT('h4)
	) name1912 (
		_w2097_,
		_w2913_,
		_w2914_
	);
	LUT2 #(
		.INIT('h2)
	) name1913 (
		_w2097_,
		_w2913_,
		_w2915_
	);
	LUT2 #(
		.INIT('h1)
	) name1914 (
		_w2914_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h1)
	) name1915 (
		_w2912_,
		_w2916_,
		_w2917_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		_w2912_,
		_w2916_,
		_w2918_
	);
	LUT2 #(
		.INIT('h1)
	) name1917 (
		_w2848_,
		_w2850_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name1918 (
		_w2851_,
		_w2919_,
		_w2920_
	);
	LUT2 #(
		.INIT('h1)
	) name1919 (
		_w2082_,
		_w2084_,
		_w2921_
	);
	LUT2 #(
		.INIT('h1)
	) name1920 (
		_w2085_,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h8)
	) name1921 (
		_w2920_,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name1922 (
		_w2090_,
		_w2091_,
		_w2924_
	);
	LUT2 #(
		.INIT('h4)
	) name1923 (
		_w2095_,
		_w2924_,
		_w2925_
	);
	LUT2 #(
		.INIT('h2)
	) name1924 (
		_w2095_,
		_w2924_,
		_w2926_
	);
	LUT2 #(
		.INIT('h1)
	) name1925 (
		_w2925_,
		_w2926_,
		_w2927_
	);
	LUT2 #(
		.INIT('h2)
	) name1926 (
		_w2923_,
		_w2927_,
		_w2928_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		_w2923_,
		_w2927_,
		_w2929_
	);
	LUT2 #(
		.INIT('h1)
	) name1928 (
		_w2856_,
		_w2857_,
		_w2930_
	);
	LUT2 #(
		.INIT('h4)
	) name1929 (
		_w2861_,
		_w2930_,
		_w2931_
	);
	LUT2 #(
		.INIT('h2)
	) name1930 (
		_w2861_,
		_w2930_,
		_w2932_
	);
	LUT2 #(
		.INIT('h1)
	) name1931 (
		_w2931_,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h1)
	) name1932 (
		_w2929_,
		_w2933_,
		_w2934_
	);
	LUT2 #(
		.INIT('h1)
	) name1933 (
		_w2928_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h4)
	) name1934 (
		_w2918_,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w2917_,
		_w2936_,
		_w2937_
	);
	LUT2 #(
		.INIT('h1)
	) name1936 (
		_w2908_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h1)
	) name1937 (
		_w2907_,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h1)
	) name1938 (
		_w2898_,
		_w2939_,
		_w2940_
	);
	LUT2 #(
		.INIT('h1)
	) name1939 (
		_w2897_,
		_w2940_,
		_w2941_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w2888_,
		_w2941_,
		_w2942_
	);
	LUT2 #(
		.INIT('h1)
	) name1941 (
		_w2887_,
		_w2942_,
		_w2943_
	);
	LUT2 #(
		.INIT('h4)
	) name1942 (
		_w2878_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h8)
	) name1943 (
		_w2108_,
		_w2944_,
		_w2945_
	);
	LUT2 #(
		.INIT('h8)
	) name1944 (
		\A[403] ,
		\A[404] ,
		_w2946_
	);
	LUT2 #(
		.INIT('h1)
	) name1945 (
		\A[403] ,
		\A[404] ,
		_w2947_
	);
	LUT2 #(
		.INIT('h1)
	) name1946 (
		_w2946_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h8)
	) name1947 (
		\A[405] ,
		_w2948_,
		_w2949_
	);
	LUT2 #(
		.INIT('h1)
	) name1948 (
		_w2946_,
		_w2949_,
		_w2950_
	);
	LUT2 #(
		.INIT('h8)
	) name1949 (
		\A[406] ,
		\A[407] ,
		_w2951_
	);
	LUT2 #(
		.INIT('h1)
	) name1950 (
		\A[405] ,
		_w2948_,
		_w2952_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		_w2949_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h1)
	) name1952 (
		\A[406] ,
		\A[407] ,
		_w2954_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		_w2951_,
		_w2954_,
		_w2955_
	);
	LUT2 #(
		.INIT('h8)
	) name1954 (
		\A[408] ,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h1)
	) name1955 (
		\A[408] ,
		_w2955_,
		_w2957_
	);
	LUT2 #(
		.INIT('h1)
	) name1956 (
		_w2956_,
		_w2957_,
		_w2958_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		_w2953_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h8)
	) name1958 (
		_w2951_,
		_w2959_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name1959 (
		_w2951_,
		_w2956_,
		_w2961_
	);
	LUT2 #(
		.INIT('h4)
	) name1960 (
		_w2959_,
		_w2961_,
		_w2962_
	);
	LUT2 #(
		.INIT('h1)
	) name1961 (
		_w2960_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h2)
	) name1962 (
		_w2950_,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h4)
	) name1963 (
		_w2950_,
		_w2963_,
		_w2965_
	);
	LUT2 #(
		.INIT('h1)
	) name1964 (
		_w2964_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h8)
	) name1965 (
		\A[409] ,
		\A[410] ,
		_w2967_
	);
	LUT2 #(
		.INIT('h1)
	) name1966 (
		\A[409] ,
		\A[410] ,
		_w2968_
	);
	LUT2 #(
		.INIT('h1)
	) name1967 (
		_w2967_,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h8)
	) name1968 (
		\A[411] ,
		_w2969_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name1969 (
		\A[411] ,
		_w2969_,
		_w2971_
	);
	LUT2 #(
		.INIT('h1)
	) name1970 (
		_w2970_,
		_w2971_,
		_w2972_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		\A[412] ,
		\A[413] ,
		_w2973_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		\A[412] ,
		\A[413] ,
		_w2974_
	);
	LUT2 #(
		.INIT('h1)
	) name1973 (
		_w2973_,
		_w2974_,
		_w2975_
	);
	LUT2 #(
		.INIT('h8)
	) name1974 (
		\A[414] ,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('h1)
	) name1975 (
		\A[414] ,
		_w2975_,
		_w2977_
	);
	LUT2 #(
		.INIT('h1)
	) name1976 (
		_w2976_,
		_w2977_,
		_w2978_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		_w2972_,
		_w2978_,
		_w2979_
	);
	LUT2 #(
		.INIT('h1)
	) name1978 (
		_w2973_,
		_w2976_,
		_w2980_
	);
	LUT2 #(
		.INIT('h1)
	) name1979 (
		_w2967_,
		_w2970_,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name1980 (
		_w2980_,
		_w2981_,
		_w2982_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		_w2980_,
		_w2981_,
		_w2983_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		_w2982_,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h4)
	) name1983 (
		_w2979_,
		_w2984_,
		_w2985_
	);
	LUT2 #(
		.INIT('h1)
	) name1984 (
		_w2953_,
		_w2958_,
		_w2986_
	);
	LUT2 #(
		.INIT('h1)
	) name1985 (
		_w2959_,
		_w2986_,
		_w2987_
	);
	LUT2 #(
		.INIT('h1)
	) name1986 (
		_w2972_,
		_w2978_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name1987 (
		_w2979_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		_w2987_,
		_w2989_,
		_w2990_
	);
	LUT2 #(
		.INIT('h2)
	) name1989 (
		_w2979_,
		_w2984_,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		_w2985_,
		_w2990_,
		_w2992_
	);
	LUT2 #(
		.INIT('h4)
	) name1991 (
		_w2991_,
		_w2992_,
		_w2993_
	);
	LUT2 #(
		.INIT('h2)
	) name1992 (
		_w2966_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		_w2984_,
		_w2990_,
		_w2995_
	);
	LUT2 #(
		.INIT('h4)
	) name1994 (
		_w2950_,
		_w2960_,
		_w2996_
	);
	LUT2 #(
		.INIT('h2)
	) name1995 (
		_w2995_,
		_w2996_,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name1996 (
		_w2994_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h4)
	) name1997 (
		_w2973_,
		_w2981_,
		_w2999_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		_w2979_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		_w2982_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('h1)
	) name2000 (
		_w2998_,
		_w3001_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name2001 (
		_w2950_,
		_w2962_,
		_w3003_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		_w2960_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h8)
	) name2003 (
		_w2998_,
		_w3001_,
		_w3005_
	);
	LUT2 #(
		.INIT('h1)
	) name2004 (
		_w3004_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('h1)
	) name2005 (
		_w3002_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		\A[397] ,
		\A[398] ,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name2007 (
		\A[397] ,
		\A[398] ,
		_w3009_
	);
	LUT2 #(
		.INIT('h1)
	) name2008 (
		_w3008_,
		_w3009_,
		_w3010_
	);
	LUT2 #(
		.INIT('h8)
	) name2009 (
		\A[399] ,
		_w3010_,
		_w3011_
	);
	LUT2 #(
		.INIT('h1)
	) name2010 (
		\A[399] ,
		_w3010_,
		_w3012_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		_w3011_,
		_w3012_,
		_w3013_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		\A[400] ,
		\A[401] ,
		_w3014_
	);
	LUT2 #(
		.INIT('h1)
	) name2013 (
		\A[400] ,
		\A[401] ,
		_w3015_
	);
	LUT2 #(
		.INIT('h1)
	) name2014 (
		_w3014_,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h8)
	) name2015 (
		\A[402] ,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('h1)
	) name2016 (
		\A[402] ,
		_w3016_,
		_w3018_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h8)
	) name2018 (
		_w3013_,
		_w3019_,
		_w3020_
	);
	LUT2 #(
		.INIT('h1)
	) name2019 (
		_w3013_,
		_w3019_,
		_w3021_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w3020_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		\A[391] ,
		\A[392] ,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name2022 (
		\A[391] ,
		\A[392] ,
		_w3024_
	);
	LUT2 #(
		.INIT('h1)
	) name2023 (
		_w3023_,
		_w3024_,
		_w3025_
	);
	LUT2 #(
		.INIT('h8)
	) name2024 (
		\A[393] ,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h1)
	) name2025 (
		\A[393] ,
		_w3025_,
		_w3027_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		_w3026_,
		_w3027_,
		_w3028_
	);
	LUT2 #(
		.INIT('h8)
	) name2027 (
		\A[394] ,
		\A[395] ,
		_w3029_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		\A[394] ,
		\A[395] ,
		_w3030_
	);
	LUT2 #(
		.INIT('h1)
	) name2029 (
		_w3029_,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h8)
	) name2030 (
		\A[396] ,
		_w3031_,
		_w3032_
	);
	LUT2 #(
		.INIT('h1)
	) name2031 (
		\A[396] ,
		_w3031_,
		_w3033_
	);
	LUT2 #(
		.INIT('h1)
	) name2032 (
		_w3032_,
		_w3033_,
		_w3034_
	);
	LUT2 #(
		.INIT('h8)
	) name2033 (
		_w3028_,
		_w3034_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name2034 (
		_w3028_,
		_w3034_,
		_w3036_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		_w3035_,
		_w3036_,
		_w3037_
	);
	LUT2 #(
		.INIT('h8)
	) name2036 (
		_w3022_,
		_w3037_,
		_w3038_
	);
	LUT2 #(
		.INIT('h1)
	) name2037 (
		_w3008_,
		_w3011_,
		_w3039_
	);
	LUT2 #(
		.INIT('h1)
	) name2038 (
		_w3014_,
		_w3017_,
		_w3040_
	);
	LUT2 #(
		.INIT('h4)
	) name2039 (
		_w3020_,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h8)
	) name2040 (
		_w3014_,
		_w3020_,
		_w3042_
	);
	LUT2 #(
		.INIT('h1)
	) name2041 (
		_w3041_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h2)
	) name2042 (
		_w3039_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h4)
	) name2043 (
		_w3039_,
		_w3043_,
		_w3045_
	);
	LUT2 #(
		.INIT('h1)
	) name2044 (
		_w3044_,
		_w3045_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name2045 (
		_w3038_,
		_w3046_,
		_w3047_
	);
	LUT2 #(
		.INIT('h1)
	) name2046 (
		_w3023_,
		_w3026_,
		_w3048_
	);
	LUT2 #(
		.INIT('h8)
	) name2047 (
		_w3029_,
		_w3035_,
		_w3049_
	);
	LUT2 #(
		.INIT('h1)
	) name2048 (
		_w3029_,
		_w3032_,
		_w3050_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		_w3035_,
		_w3050_,
		_w3051_
	);
	LUT2 #(
		.INIT('h1)
	) name2050 (
		_w3049_,
		_w3051_,
		_w3052_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		_w3048_,
		_w3052_,
		_w3053_
	);
	LUT2 #(
		.INIT('h4)
	) name2052 (
		_w3048_,
		_w3052_,
		_w3054_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w3053_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h4)
	) name2054 (
		_w3047_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h8)
	) name2055 (
		_w3038_,
		_w3046_,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name2056 (
		_w3039_,
		_w3040_,
		_w3058_
	);
	LUT2 #(
		.INIT('h4)
	) name2057 (
		_w3048_,
		_w3049_,
		_w3059_
	);
	LUT2 #(
		.INIT('h1)
	) name2058 (
		_w3058_,
		_w3059_,
		_w3060_
	);
	LUT2 #(
		.INIT('h8)
	) name2059 (
		_w3057_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		_w3056_,
		_w3061_,
		_w3062_
	);
	LUT2 #(
		.INIT('h1)
	) name2061 (
		_w3039_,
		_w3041_,
		_w3063_
	);
	LUT2 #(
		.INIT('h1)
	) name2062 (
		_w3042_,
		_w3063_,
		_w3064_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		_w3062_,
		_w3064_,
		_w3065_
	);
	LUT2 #(
		.INIT('h1)
	) name2064 (
		_w3048_,
		_w3051_,
		_w3066_
	);
	LUT2 #(
		.INIT('h1)
	) name2065 (
		_w3049_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		_w3062_,
		_w3064_,
		_w3068_
	);
	LUT2 #(
		.INIT('h1)
	) name2067 (
		_w3067_,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('h1)
	) name2068 (
		_w3065_,
		_w3069_,
		_w3070_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		_w3007_,
		_w3070_,
		_w3071_
	);
	LUT2 #(
		.INIT('h8)
	) name2070 (
		_w3007_,
		_w3070_,
		_w3072_
	);
	LUT2 #(
		.INIT('h1)
	) name2071 (
		_w3065_,
		_w3068_,
		_w3073_
	);
	LUT2 #(
		.INIT('h2)
	) name2072 (
		_w3067_,
		_w3073_,
		_w3074_
	);
	LUT2 #(
		.INIT('h4)
	) name2073 (
		_w3067_,
		_w3073_,
		_w3075_
	);
	LUT2 #(
		.INIT('h1)
	) name2074 (
		_w3074_,
		_w3075_,
		_w3076_
	);
	LUT2 #(
		.INIT('h1)
	) name2075 (
		_w3002_,
		_w3005_,
		_w3077_
	);
	LUT2 #(
		.INIT('h2)
	) name2076 (
		_w3004_,
		_w3077_,
		_w3078_
	);
	LUT2 #(
		.INIT('h4)
	) name2077 (
		_w3004_,
		_w3077_,
		_w3079_
	);
	LUT2 #(
		.INIT('h1)
	) name2078 (
		_w3078_,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h1)
	) name2079 (
		_w3076_,
		_w3080_,
		_w3081_
	);
	LUT2 #(
		.INIT('h1)
	) name2080 (
		_w2987_,
		_w2989_,
		_w3082_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w2990_,
		_w3082_,
		_w3083_
	);
	LUT2 #(
		.INIT('h1)
	) name2082 (
		_w3022_,
		_w3037_,
		_w3084_
	);
	LUT2 #(
		.INIT('h1)
	) name2083 (
		_w3038_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		_w3083_,
		_w3085_,
		_w3086_
	);
	LUT2 #(
		.INIT('h2)
	) name2085 (
		_w2994_,
		_w2997_,
		_w3087_
	);
	LUT2 #(
		.INIT('h1)
	) name2086 (
		_w2993_,
		_w2995_,
		_w3088_
	);
	LUT2 #(
		.INIT('h1)
	) name2087 (
		_w2966_,
		_w3088_,
		_w3089_
	);
	LUT2 #(
		.INIT('h1)
	) name2088 (
		_w3087_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h1)
	) name2089 (
		_w3086_,
		_w3090_,
		_w3091_
	);
	LUT2 #(
		.INIT('h2)
	) name2090 (
		_w3056_,
		_w3061_,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name2091 (
		_w3047_,
		_w3057_,
		_w3093_
	);
	LUT2 #(
		.INIT('h1)
	) name2092 (
		_w3055_,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h1)
	) name2093 (
		_w3092_,
		_w3094_,
		_w3095_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		_w3086_,
		_w3090_,
		_w3096_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h1)
	) name2096 (
		_w3091_,
		_w3097_,
		_w3098_
	);
	LUT2 #(
		.INIT('h8)
	) name2097 (
		_w3076_,
		_w3080_,
		_w3099_
	);
	LUT2 #(
		.INIT('h1)
	) name2098 (
		_w3098_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h1)
	) name2099 (
		_w3081_,
		_w3100_,
		_w3101_
	);
	LUT2 #(
		.INIT('h4)
	) name2100 (
		_w3072_,
		_w3101_,
		_w3102_
	);
	LUT2 #(
		.INIT('h1)
	) name2101 (
		_w3071_,
		_w3102_,
		_w3103_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		\A[385] ,
		\A[386] ,
		_w3104_
	);
	LUT2 #(
		.INIT('h1)
	) name2103 (
		\A[385] ,
		\A[386] ,
		_w3105_
	);
	LUT2 #(
		.INIT('h1)
	) name2104 (
		_w3104_,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('h8)
	) name2105 (
		\A[387] ,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h1)
	) name2106 (
		\A[387] ,
		_w3106_,
		_w3108_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		_w3107_,
		_w3108_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		\A[388] ,
		\A[389] ,
		_w3110_
	);
	LUT2 #(
		.INIT('h1)
	) name2109 (
		\A[388] ,
		\A[389] ,
		_w3111_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		_w3110_,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h8)
	) name2111 (
		\A[390] ,
		_w3112_,
		_w3113_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		\A[390] ,
		_w3112_,
		_w3114_
	);
	LUT2 #(
		.INIT('h1)
	) name2113 (
		_w3113_,
		_w3114_,
		_w3115_
	);
	LUT2 #(
		.INIT('h8)
	) name2114 (
		_w3109_,
		_w3115_,
		_w3116_
	);
	LUT2 #(
		.INIT('h1)
	) name2115 (
		_w3109_,
		_w3115_,
		_w3117_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		_w3116_,
		_w3117_,
		_w3118_
	);
	LUT2 #(
		.INIT('h8)
	) name2117 (
		\A[379] ,
		\A[380] ,
		_w3119_
	);
	LUT2 #(
		.INIT('h1)
	) name2118 (
		\A[379] ,
		\A[380] ,
		_w3120_
	);
	LUT2 #(
		.INIT('h1)
	) name2119 (
		_w3119_,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h8)
	) name2120 (
		\A[381] ,
		_w3121_,
		_w3122_
	);
	LUT2 #(
		.INIT('h1)
	) name2121 (
		\A[381] ,
		_w3121_,
		_w3123_
	);
	LUT2 #(
		.INIT('h1)
	) name2122 (
		_w3122_,
		_w3123_,
		_w3124_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		\A[382] ,
		\A[383] ,
		_w3125_
	);
	LUT2 #(
		.INIT('h1)
	) name2124 (
		\A[382] ,
		\A[383] ,
		_w3126_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w3125_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		\A[384] ,
		_w3127_,
		_w3128_
	);
	LUT2 #(
		.INIT('h1)
	) name2127 (
		\A[384] ,
		_w3127_,
		_w3129_
	);
	LUT2 #(
		.INIT('h1)
	) name2128 (
		_w3128_,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h8)
	) name2129 (
		_w3124_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h1)
	) name2130 (
		_w3124_,
		_w3130_,
		_w3132_
	);
	LUT2 #(
		.INIT('h1)
	) name2131 (
		_w3131_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name2132 (
		_w3118_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h1)
	) name2133 (
		_w3110_,
		_w3113_,
		_w3135_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w3104_,
		_w3107_,
		_w3136_
	);
	LUT2 #(
		.INIT('h1)
	) name2135 (
		_w3135_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h8)
	) name2136 (
		_w3135_,
		_w3136_,
		_w3138_
	);
	LUT2 #(
		.INIT('h1)
	) name2137 (
		_w3137_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h8)
	) name2138 (
		_w3134_,
		_w3139_,
		_w3140_
	);
	LUT2 #(
		.INIT('h1)
	) name2139 (
		_w3119_,
		_w3122_,
		_w3141_
	);
	LUT2 #(
		.INIT('h1)
	) name2140 (
		_w3125_,
		_w3128_,
		_w3142_
	);
	LUT2 #(
		.INIT('h4)
	) name2141 (
		_w3131_,
		_w3142_,
		_w3143_
	);
	LUT2 #(
		.INIT('h8)
	) name2142 (
		_w3125_,
		_w3131_,
		_w3144_
	);
	LUT2 #(
		.INIT('h1)
	) name2143 (
		_w3143_,
		_w3144_,
		_w3145_
	);
	LUT2 #(
		.INIT('h2)
	) name2144 (
		_w3141_,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('h4)
	) name2145 (
		_w3141_,
		_w3145_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name2146 (
		_w3146_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h1)
	) name2147 (
		_w3140_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h4)
	) name2148 (
		_w3116_,
		_w3139_,
		_w3150_
	);
	LUT2 #(
		.INIT('h2)
	) name2149 (
		_w3116_,
		_w3139_,
		_w3151_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		_w3134_,
		_w3150_,
		_w3152_
	);
	LUT2 #(
		.INIT('h4)
	) name2151 (
		_w3151_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h1)
	) name2152 (
		_w3149_,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h1)
	) name2153 (
		_w3116_,
		_w3137_,
		_w3155_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w3138_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h1)
	) name2155 (
		_w3154_,
		_w3156_,
		_w3157_
	);
	LUT2 #(
		.INIT('h8)
	) name2156 (
		_w3154_,
		_w3156_,
		_w3158_
	);
	LUT2 #(
		.INIT('h1)
	) name2157 (
		_w3141_,
		_w3143_,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name2158 (
		_w3144_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h4)
	) name2159 (
		_w3158_,
		_w3160_,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name2160 (
		_w3157_,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h1)
	) name2161 (
		_w3157_,
		_w3158_,
		_w3163_
	);
	LUT2 #(
		.INIT('h4)
	) name2162 (
		_w3160_,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h2)
	) name2163 (
		_w3160_,
		_w3163_,
		_w3165_
	);
	LUT2 #(
		.INIT('h1)
	) name2164 (
		_w3164_,
		_w3165_,
		_w3166_
	);
	LUT2 #(
		.INIT('h8)
	) name2165 (
		\A[370] ,
		\A[371] ,
		_w3167_
	);
	LUT2 #(
		.INIT('h8)
	) name2166 (
		\A[367] ,
		\A[368] ,
		_w3168_
	);
	LUT2 #(
		.INIT('h1)
	) name2167 (
		\A[367] ,
		\A[368] ,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name2168 (
		_w3168_,
		_w3169_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name2169 (
		\A[369] ,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		\A[369] ,
		_w3170_,
		_w3172_
	);
	LUT2 #(
		.INIT('h1)
	) name2171 (
		_w3171_,
		_w3172_,
		_w3173_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		\A[370] ,
		\A[371] ,
		_w3174_
	);
	LUT2 #(
		.INIT('h1)
	) name2173 (
		_w3167_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h8)
	) name2174 (
		\A[372] ,
		_w3175_,
		_w3176_
	);
	LUT2 #(
		.INIT('h1)
	) name2175 (
		\A[372] ,
		_w3175_,
		_w3177_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w3176_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h8)
	) name2177 (
		_w3173_,
		_w3178_,
		_w3179_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		_w3167_,
		_w3179_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name2179 (
		_w3168_,
		_w3171_,
		_w3181_
	);
	LUT2 #(
		.INIT('h1)
	) name2180 (
		_w3167_,
		_w3176_,
		_w3182_
	);
	LUT2 #(
		.INIT('h4)
	) name2181 (
		_w3179_,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		_w3181_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h1)
	) name2183 (
		_w3180_,
		_w3184_,
		_w3185_
	);
	LUT2 #(
		.INIT('h8)
	) name2184 (
		\A[373] ,
		\A[374] ,
		_w3186_
	);
	LUT2 #(
		.INIT('h1)
	) name2185 (
		\A[373] ,
		\A[374] ,
		_w3187_
	);
	LUT2 #(
		.INIT('h1)
	) name2186 (
		_w3186_,
		_w3187_,
		_w3188_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		\A[375] ,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h1)
	) name2188 (
		\A[375] ,
		_w3188_,
		_w3190_
	);
	LUT2 #(
		.INIT('h1)
	) name2189 (
		_w3189_,
		_w3190_,
		_w3191_
	);
	LUT2 #(
		.INIT('h8)
	) name2190 (
		\A[376] ,
		\A[377] ,
		_w3192_
	);
	LUT2 #(
		.INIT('h1)
	) name2191 (
		\A[376] ,
		\A[377] ,
		_w3193_
	);
	LUT2 #(
		.INIT('h1)
	) name2192 (
		_w3192_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h8)
	) name2193 (
		\A[378] ,
		_w3194_,
		_w3195_
	);
	LUT2 #(
		.INIT('h1)
	) name2194 (
		\A[378] ,
		_w3194_,
		_w3196_
	);
	LUT2 #(
		.INIT('h1)
	) name2195 (
		_w3195_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h8)
	) name2196 (
		_w3191_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('h1)
	) name2197 (
		_w3191_,
		_w3197_,
		_w3199_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		_w3198_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h1)
	) name2199 (
		_w3173_,
		_w3178_,
		_w3201_
	);
	LUT2 #(
		.INIT('h1)
	) name2200 (
		_w3179_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h8)
	) name2201 (
		_w3200_,
		_w3202_,
		_w3203_
	);
	LUT2 #(
		.INIT('h1)
	) name2202 (
		_w3192_,
		_w3195_,
		_w3204_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w3186_,
		_w3189_,
		_w3205_
	);
	LUT2 #(
		.INIT('h1)
	) name2204 (
		_w3204_,
		_w3205_,
		_w3206_
	);
	LUT2 #(
		.INIT('h8)
	) name2205 (
		_w3204_,
		_w3205_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w3206_,
		_w3207_,
		_w3208_
	);
	LUT2 #(
		.INIT('h8)
	) name2207 (
		_w3203_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		_w3180_,
		_w3183_,
		_w3210_
	);
	LUT2 #(
		.INIT('h2)
	) name2209 (
		_w3181_,
		_w3210_,
		_w3211_
	);
	LUT2 #(
		.INIT('h4)
	) name2210 (
		_w3181_,
		_w3210_,
		_w3212_
	);
	LUT2 #(
		.INIT('h1)
	) name2211 (
		_w3211_,
		_w3212_,
		_w3213_
	);
	LUT2 #(
		.INIT('h1)
	) name2212 (
		_w3209_,
		_w3213_,
		_w3214_
	);
	LUT2 #(
		.INIT('h4)
	) name2213 (
		_w3198_,
		_w3208_,
		_w3215_
	);
	LUT2 #(
		.INIT('h2)
	) name2214 (
		_w3198_,
		_w3208_,
		_w3216_
	);
	LUT2 #(
		.INIT('h1)
	) name2215 (
		_w3203_,
		_w3215_,
		_w3217_
	);
	LUT2 #(
		.INIT('h4)
	) name2216 (
		_w3216_,
		_w3217_,
		_w3218_
	);
	LUT2 #(
		.INIT('h1)
	) name2217 (
		_w3214_,
		_w3218_,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w3198_,
		_w3206_,
		_w3220_
	);
	LUT2 #(
		.INIT('h1)
	) name2219 (
		_w3207_,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h8)
	) name2220 (
		_w3219_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h1)
	) name2221 (
		_w3219_,
		_w3221_,
		_w3223_
	);
	LUT2 #(
		.INIT('h1)
	) name2222 (
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		_w3185_,
		_w3224_,
		_w3225_
	);
	LUT2 #(
		.INIT('h4)
	) name2224 (
		_w3185_,
		_w3224_,
		_w3226_
	);
	LUT2 #(
		.INIT('h1)
	) name2225 (
		_w3225_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h8)
	) name2226 (
		_w3166_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		_w3166_,
		_w3227_,
		_w3229_
	);
	LUT2 #(
		.INIT('h1)
	) name2228 (
		_w3118_,
		_w3133_,
		_w3230_
	);
	LUT2 #(
		.INIT('h1)
	) name2229 (
		_w3134_,
		_w3230_,
		_w3231_
	);
	LUT2 #(
		.INIT('h1)
	) name2230 (
		_w3200_,
		_w3202_,
		_w3232_
	);
	LUT2 #(
		.INIT('h1)
	) name2231 (
		_w3203_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h8)
	) name2232 (
		_w3231_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w3140_,
		_w3153_,
		_w3235_
	);
	LUT2 #(
		.INIT('h4)
	) name2234 (
		_w3148_,
		_w3235_,
		_w3236_
	);
	LUT2 #(
		.INIT('h2)
	) name2235 (
		_w3148_,
		_w3235_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name2236 (
		_w3236_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h2)
	) name2237 (
		_w3234_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h4)
	) name2238 (
		_w3234_,
		_w3238_,
		_w3240_
	);
	LUT2 #(
		.INIT('h1)
	) name2239 (
		_w3209_,
		_w3218_,
		_w3241_
	);
	LUT2 #(
		.INIT('h4)
	) name2240 (
		_w3213_,
		_w3241_,
		_w3242_
	);
	LUT2 #(
		.INIT('h2)
	) name2241 (
		_w3213_,
		_w3241_,
		_w3243_
	);
	LUT2 #(
		.INIT('h1)
	) name2242 (
		_w3242_,
		_w3243_,
		_w3244_
	);
	LUT2 #(
		.INIT('h1)
	) name2243 (
		_w3240_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('h1)
	) name2244 (
		_w3239_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name2245 (
		_w3229_,
		_w3246_,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name2246 (
		_w3228_,
		_w3247_,
		_w3248_
	);
	LUT2 #(
		.INIT('h2)
	) name2247 (
		_w3162_,
		_w3248_,
		_w3249_
	);
	LUT2 #(
		.INIT('h4)
	) name2248 (
		_w3162_,
		_w3248_,
		_w3250_
	);
	LUT2 #(
		.INIT('h2)
	) name2249 (
		_w3185_,
		_w3222_,
		_w3251_
	);
	LUT2 #(
		.INIT('h1)
	) name2250 (
		_w3223_,
		_w3251_,
		_w3252_
	);
	LUT2 #(
		.INIT('h4)
	) name2251 (
		_w3250_,
		_w3252_,
		_w3253_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		_w3249_,
		_w3253_,
		_w3254_
	);
	LUT2 #(
		.INIT('h1)
	) name2253 (
		_w3103_,
		_w3254_,
		_w3255_
	);
	LUT2 #(
		.INIT('h8)
	) name2254 (
		_w3103_,
		_w3254_,
		_w3256_
	);
	LUT2 #(
		.INIT('h1)
	) name2255 (
		_w3071_,
		_w3072_,
		_w3257_
	);
	LUT2 #(
		.INIT('h2)
	) name2256 (
		_w3101_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h4)
	) name2257 (
		_w3101_,
		_w3257_,
		_w3259_
	);
	LUT2 #(
		.INIT('h1)
	) name2258 (
		_w3258_,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h1)
	) name2259 (
		_w3249_,
		_w3250_,
		_w3261_
	);
	LUT2 #(
		.INIT('h8)
	) name2260 (
		_w3252_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('h1)
	) name2261 (
		_w3252_,
		_w3261_,
		_w3263_
	);
	LUT2 #(
		.INIT('h1)
	) name2262 (
		_w3262_,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h4)
	) name2263 (
		_w3260_,
		_w3264_,
		_w3265_
	);
	LUT2 #(
		.INIT('h2)
	) name2264 (
		_w3260_,
		_w3264_,
		_w3266_
	);
	LUT2 #(
		.INIT('h1)
	) name2265 (
		_w3081_,
		_w3099_,
		_w3267_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		_w3098_,
		_w3267_,
		_w3268_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		_w3098_,
		_w3267_,
		_w3269_
	);
	LUT2 #(
		.INIT('h1)
	) name2268 (
		_w3268_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h1)
	) name2269 (
		_w3228_,
		_w3229_,
		_w3271_
	);
	LUT2 #(
		.INIT('h4)
	) name2270 (
		_w3246_,
		_w3271_,
		_w3272_
	);
	LUT2 #(
		.INIT('h2)
	) name2271 (
		_w3246_,
		_w3271_,
		_w3273_
	);
	LUT2 #(
		.INIT('h1)
	) name2272 (
		_w3272_,
		_w3273_,
		_w3274_
	);
	LUT2 #(
		.INIT('h8)
	) name2273 (
		_w3270_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h1)
	) name2274 (
		_w3270_,
		_w3274_,
		_w3276_
	);
	LUT2 #(
		.INIT('h1)
	) name2275 (
		_w3083_,
		_w3085_,
		_w3277_
	);
	LUT2 #(
		.INIT('h1)
	) name2276 (
		_w3086_,
		_w3277_,
		_w3278_
	);
	LUT2 #(
		.INIT('h1)
	) name2277 (
		_w3231_,
		_w3233_,
		_w3279_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		_w3234_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h8)
	) name2279 (
		_w3278_,
		_w3280_,
		_w3281_
	);
	LUT2 #(
		.INIT('h1)
	) name2280 (
		_w3091_,
		_w3096_,
		_w3282_
	);
	LUT2 #(
		.INIT('h2)
	) name2281 (
		_w3095_,
		_w3282_,
		_w3283_
	);
	LUT2 #(
		.INIT('h4)
	) name2282 (
		_w3095_,
		_w3282_,
		_w3284_
	);
	LUT2 #(
		.INIT('h1)
	) name2283 (
		_w3283_,
		_w3284_,
		_w3285_
	);
	LUT2 #(
		.INIT('h2)
	) name2284 (
		_w3281_,
		_w3285_,
		_w3286_
	);
	LUT2 #(
		.INIT('h4)
	) name2285 (
		_w3281_,
		_w3285_,
		_w3287_
	);
	LUT2 #(
		.INIT('h1)
	) name2286 (
		_w3239_,
		_w3240_,
		_w3288_
	);
	LUT2 #(
		.INIT('h4)
	) name2287 (
		_w3244_,
		_w3288_,
		_w3289_
	);
	LUT2 #(
		.INIT('h2)
	) name2288 (
		_w3244_,
		_w3288_,
		_w3290_
	);
	LUT2 #(
		.INIT('h1)
	) name2289 (
		_w3289_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('h4)
	) name2290 (
		_w3287_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w3286_,
		_w3292_,
		_w3293_
	);
	LUT2 #(
		.INIT('h1)
	) name2292 (
		_w3276_,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('h1)
	) name2293 (
		_w3275_,
		_w3294_,
		_w3295_
	);
	LUT2 #(
		.INIT('h1)
	) name2294 (
		_w3266_,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w3265_,
		_w3296_,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name2296 (
		_w3256_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h1)
	) name2297 (
		_w3255_,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('h8)
	) name2298 (
		\A[445] ,
		\A[446] ,
		_w3300_
	);
	LUT2 #(
		.INIT('h1)
	) name2299 (
		\A[445] ,
		\A[446] ,
		_w3301_
	);
	LUT2 #(
		.INIT('h1)
	) name2300 (
		_w3300_,
		_w3301_,
		_w3302_
	);
	LUT2 #(
		.INIT('h8)
	) name2301 (
		\A[447] ,
		_w3302_,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		\A[447] ,
		_w3302_,
		_w3304_
	);
	LUT2 #(
		.INIT('h1)
	) name2303 (
		_w3303_,
		_w3304_,
		_w3305_
	);
	LUT2 #(
		.INIT('h8)
	) name2304 (
		\A[448] ,
		\A[449] ,
		_w3306_
	);
	LUT2 #(
		.INIT('h1)
	) name2305 (
		\A[448] ,
		\A[449] ,
		_w3307_
	);
	LUT2 #(
		.INIT('h1)
	) name2306 (
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h8)
	) name2307 (
		\A[450] ,
		_w3308_,
		_w3309_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		\A[450] ,
		_w3308_,
		_w3310_
	);
	LUT2 #(
		.INIT('h1)
	) name2309 (
		_w3309_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h8)
	) name2310 (
		_w3305_,
		_w3311_,
		_w3312_
	);
	LUT2 #(
		.INIT('h1)
	) name2311 (
		_w3305_,
		_w3311_,
		_w3313_
	);
	LUT2 #(
		.INIT('h1)
	) name2312 (
		_w3312_,
		_w3313_,
		_w3314_
	);
	LUT2 #(
		.INIT('h8)
	) name2313 (
		\A[439] ,
		\A[440] ,
		_w3315_
	);
	LUT2 #(
		.INIT('h1)
	) name2314 (
		\A[439] ,
		\A[440] ,
		_w3316_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w3315_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('h8)
	) name2316 (
		\A[441] ,
		_w3317_,
		_w3318_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		\A[441] ,
		_w3317_,
		_w3319_
	);
	LUT2 #(
		.INIT('h1)
	) name2318 (
		_w3318_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h8)
	) name2319 (
		\A[442] ,
		\A[443] ,
		_w3321_
	);
	LUT2 #(
		.INIT('h1)
	) name2320 (
		\A[442] ,
		\A[443] ,
		_w3322_
	);
	LUT2 #(
		.INIT('h1)
	) name2321 (
		_w3321_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h8)
	) name2322 (
		\A[444] ,
		_w3323_,
		_w3324_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		\A[444] ,
		_w3323_,
		_w3325_
	);
	LUT2 #(
		.INIT('h1)
	) name2324 (
		_w3324_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		_w3320_,
		_w3326_,
		_w3327_
	);
	LUT2 #(
		.INIT('h1)
	) name2326 (
		_w3320_,
		_w3326_,
		_w3328_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w3327_,
		_w3328_,
		_w3329_
	);
	LUT2 #(
		.INIT('h8)
	) name2328 (
		_w3314_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h1)
	) name2329 (
		_w3300_,
		_w3303_,
		_w3331_
	);
	LUT2 #(
		.INIT('h1)
	) name2330 (
		_w3306_,
		_w3309_,
		_w3332_
	);
	LUT2 #(
		.INIT('h4)
	) name2331 (
		_w3312_,
		_w3332_,
		_w3333_
	);
	LUT2 #(
		.INIT('h8)
	) name2332 (
		_w3306_,
		_w3312_,
		_w3334_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w3333_,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h2)
	) name2334 (
		_w3331_,
		_w3335_,
		_w3336_
	);
	LUT2 #(
		.INIT('h4)
	) name2335 (
		_w3331_,
		_w3335_,
		_w3337_
	);
	LUT2 #(
		.INIT('h1)
	) name2336 (
		_w3336_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h1)
	) name2337 (
		_w3330_,
		_w3338_,
		_w3339_
	);
	LUT2 #(
		.INIT('h1)
	) name2338 (
		_w3315_,
		_w3318_,
		_w3340_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		_w3321_,
		_w3327_,
		_w3341_
	);
	LUT2 #(
		.INIT('h1)
	) name2340 (
		_w3321_,
		_w3324_,
		_w3342_
	);
	LUT2 #(
		.INIT('h4)
	) name2341 (
		_w3327_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h1)
	) name2342 (
		_w3341_,
		_w3343_,
		_w3344_
	);
	LUT2 #(
		.INIT('h2)
	) name2343 (
		_w3340_,
		_w3344_,
		_w3345_
	);
	LUT2 #(
		.INIT('h4)
	) name2344 (
		_w3340_,
		_w3344_,
		_w3346_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h4)
	) name2346 (
		_w3339_,
		_w3347_,
		_w3348_
	);
	LUT2 #(
		.INIT('h8)
	) name2347 (
		_w3330_,
		_w3338_,
		_w3349_
	);
	LUT2 #(
		.INIT('h1)
	) name2348 (
		_w3331_,
		_w3332_,
		_w3350_
	);
	LUT2 #(
		.INIT('h4)
	) name2349 (
		_w3340_,
		_w3341_,
		_w3351_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		_w3350_,
		_w3351_,
		_w3352_
	);
	LUT2 #(
		.INIT('h8)
	) name2351 (
		_w3349_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h1)
	) name2352 (
		_w3348_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h1)
	) name2353 (
		_w3331_,
		_w3333_,
		_w3355_
	);
	LUT2 #(
		.INIT('h1)
	) name2354 (
		_w3334_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h1)
	) name2355 (
		_w3354_,
		_w3356_,
		_w3357_
	);
	LUT2 #(
		.INIT('h1)
	) name2356 (
		_w3340_,
		_w3343_,
		_w3358_
	);
	LUT2 #(
		.INIT('h1)
	) name2357 (
		_w3341_,
		_w3358_,
		_w3359_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		_w3354_,
		_w3356_,
		_w3360_
	);
	LUT2 #(
		.INIT('h1)
	) name2359 (
		_w3359_,
		_w3360_,
		_w3361_
	);
	LUT2 #(
		.INIT('h1)
	) name2360 (
		_w3357_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h8)
	) name2361 (
		\A[451] ,
		\A[452] ,
		_w3363_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		\A[451] ,
		\A[452] ,
		_w3364_
	);
	LUT2 #(
		.INIT('h1)
	) name2363 (
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h8)
	) name2364 (
		\A[453] ,
		_w3365_,
		_w3366_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		\A[453] ,
		_w3365_,
		_w3367_
	);
	LUT2 #(
		.INIT('h1)
	) name2366 (
		_w3366_,
		_w3367_,
		_w3368_
	);
	LUT2 #(
		.INIT('h8)
	) name2367 (
		\A[454] ,
		\A[455] ,
		_w3369_
	);
	LUT2 #(
		.INIT('h1)
	) name2368 (
		\A[454] ,
		\A[455] ,
		_w3370_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		_w3369_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name2370 (
		\A[456] ,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		\A[456] ,
		_w3371_,
		_w3373_
	);
	LUT2 #(
		.INIT('h1)
	) name2372 (
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		_w3368_,
		_w3374_,
		_w3375_
	);
	LUT2 #(
		.INIT('h1)
	) name2374 (
		_w3369_,
		_w3372_,
		_w3376_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w3363_,
		_w3366_,
		_w3377_
	);
	LUT2 #(
		.INIT('h8)
	) name2376 (
		_w3376_,
		_w3377_,
		_w3378_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		_w3376_,
		_w3377_,
		_w3379_
	);
	LUT2 #(
		.INIT('h1)
	) name2378 (
		_w3378_,
		_w3379_,
		_w3380_
	);
	LUT2 #(
		.INIT('h2)
	) name2379 (
		_w3375_,
		_w3380_,
		_w3381_
	);
	LUT2 #(
		.INIT('h4)
	) name2380 (
		_w3375_,
		_w3380_,
		_w3382_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		_w3381_,
		_w3382_,
		_w3383_
	);
	LUT2 #(
		.INIT('h8)
	) name2382 (
		\A[457] ,
		\A[458] ,
		_w3384_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		\A[457] ,
		\A[458] ,
		_w3385_
	);
	LUT2 #(
		.INIT('h1)
	) name2384 (
		_w3384_,
		_w3385_,
		_w3386_
	);
	LUT2 #(
		.INIT('h8)
	) name2385 (
		\A[459] ,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		\A[459] ,
		_w3386_,
		_w3388_
	);
	LUT2 #(
		.INIT('h1)
	) name2387 (
		_w3387_,
		_w3388_,
		_w3389_
	);
	LUT2 #(
		.INIT('h8)
	) name2388 (
		\A[460] ,
		\A[461] ,
		_w3390_
	);
	LUT2 #(
		.INIT('h1)
	) name2389 (
		\A[460] ,
		\A[461] ,
		_w3391_
	);
	LUT2 #(
		.INIT('h1)
	) name2390 (
		_w3390_,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		\A[462] ,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h1)
	) name2392 (
		\A[462] ,
		_w3392_,
		_w3394_
	);
	LUT2 #(
		.INIT('h1)
	) name2393 (
		_w3393_,
		_w3394_,
		_w3395_
	);
	LUT2 #(
		.INIT('h8)
	) name2394 (
		_w3389_,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h1)
	) name2395 (
		_w3390_,
		_w3393_,
		_w3397_
	);
	LUT2 #(
		.INIT('h1)
	) name2396 (
		_w3384_,
		_w3387_,
		_w3398_
	);
	LUT2 #(
		.INIT('h1)
	) name2397 (
		_w3397_,
		_w3398_,
		_w3399_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		_w3397_,
		_w3398_,
		_w3400_
	);
	LUT2 #(
		.INIT('h1)
	) name2399 (
		_w3399_,
		_w3400_,
		_w3401_
	);
	LUT2 #(
		.INIT('h4)
	) name2400 (
		_w3396_,
		_w3401_,
		_w3402_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		_w3389_,
		_w3395_,
		_w3403_
	);
	LUT2 #(
		.INIT('h1)
	) name2402 (
		_w3396_,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('h1)
	) name2403 (
		_w3368_,
		_w3374_,
		_w3405_
	);
	LUT2 #(
		.INIT('h1)
	) name2404 (
		_w3375_,
		_w3405_,
		_w3406_
	);
	LUT2 #(
		.INIT('h8)
	) name2405 (
		_w3404_,
		_w3406_,
		_w3407_
	);
	LUT2 #(
		.INIT('h2)
	) name2406 (
		_w3396_,
		_w3401_,
		_w3408_
	);
	LUT2 #(
		.INIT('h1)
	) name2407 (
		_w3402_,
		_w3407_,
		_w3409_
	);
	LUT2 #(
		.INIT('h4)
	) name2408 (
		_w3408_,
		_w3409_,
		_w3410_
	);
	LUT2 #(
		.INIT('h1)
	) name2409 (
		_w3383_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h8)
	) name2410 (
		_w3375_,
		_w3379_,
		_w3412_
	);
	LUT2 #(
		.INIT('h8)
	) name2411 (
		_w3401_,
		_w3407_,
		_w3413_
	);
	LUT2 #(
		.INIT('h4)
	) name2412 (
		_w3412_,
		_w3413_,
		_w3414_
	);
	LUT2 #(
		.INIT('h1)
	) name2413 (
		_w3411_,
		_w3414_,
		_w3415_
	);
	LUT2 #(
		.INIT('h4)
	) name2414 (
		_w3390_,
		_w3398_,
		_w3416_
	);
	LUT2 #(
		.INIT('h2)
	) name2415 (
		_w3396_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('h1)
	) name2416 (
		_w3399_,
		_w3417_,
		_w3418_
	);
	LUT2 #(
		.INIT('h8)
	) name2417 (
		_w3415_,
		_w3418_,
		_w3419_
	);
	LUT2 #(
		.INIT('h1)
	) name2418 (
		_w3415_,
		_w3418_,
		_w3420_
	);
	LUT2 #(
		.INIT('h1)
	) name2419 (
		_w3375_,
		_w3379_,
		_w3421_
	);
	LUT2 #(
		.INIT('h1)
	) name2420 (
		_w3378_,
		_w3421_,
		_w3422_
	);
	LUT2 #(
		.INIT('h1)
	) name2421 (
		_w3420_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h1)
	) name2422 (
		_w3419_,
		_w3423_,
		_w3424_
	);
	LUT2 #(
		.INIT('h4)
	) name2423 (
		_w3362_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h2)
	) name2424 (
		_w3362_,
		_w3424_,
		_w3426_
	);
	LUT2 #(
		.INIT('h1)
	) name2425 (
		_w3357_,
		_w3360_,
		_w3427_
	);
	LUT2 #(
		.INIT('h2)
	) name2426 (
		_w3359_,
		_w3427_,
		_w3428_
	);
	LUT2 #(
		.INIT('h4)
	) name2427 (
		_w3359_,
		_w3427_,
		_w3429_
	);
	LUT2 #(
		.INIT('h1)
	) name2428 (
		_w3428_,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w3419_,
		_w3420_,
		_w3431_
	);
	LUT2 #(
		.INIT('h4)
	) name2430 (
		_w3422_,
		_w3431_,
		_w3432_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		_w3422_,
		_w3431_,
		_w3433_
	);
	LUT2 #(
		.INIT('h1)
	) name2432 (
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h2)
	) name2433 (
		_w3430_,
		_w3434_,
		_w3435_
	);
	LUT2 #(
		.INIT('h4)
	) name2434 (
		_w3430_,
		_w3434_,
		_w3436_
	);
	LUT2 #(
		.INIT('h1)
	) name2435 (
		_w3404_,
		_w3406_,
		_w3437_
	);
	LUT2 #(
		.INIT('h1)
	) name2436 (
		_w3407_,
		_w3437_,
		_w3438_
	);
	LUT2 #(
		.INIT('h1)
	) name2437 (
		_w3314_,
		_w3329_,
		_w3439_
	);
	LUT2 #(
		.INIT('h1)
	) name2438 (
		_w3330_,
		_w3439_,
		_w3440_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		_w3438_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h2)
	) name2440 (
		_w3411_,
		_w3414_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name2441 (
		_w3410_,
		_w3413_,
		_w3443_
	);
	LUT2 #(
		.INIT('h2)
	) name2442 (
		_w3383_,
		_w3443_,
		_w3444_
	);
	LUT2 #(
		.INIT('h1)
	) name2443 (
		_w3442_,
		_w3444_,
		_w3445_
	);
	LUT2 #(
		.INIT('h1)
	) name2444 (
		_w3441_,
		_w3445_,
		_w3446_
	);
	LUT2 #(
		.INIT('h2)
	) name2445 (
		_w3348_,
		_w3353_,
		_w3447_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		_w3339_,
		_w3349_,
		_w3448_
	);
	LUT2 #(
		.INIT('h1)
	) name2447 (
		_w3347_,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h1)
	) name2448 (
		_w3447_,
		_w3449_,
		_w3450_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		_w3441_,
		_w3445_,
		_w3451_
	);
	LUT2 #(
		.INIT('h1)
	) name2450 (
		_w3450_,
		_w3451_,
		_w3452_
	);
	LUT2 #(
		.INIT('h1)
	) name2451 (
		_w3446_,
		_w3452_,
		_w3453_
	);
	LUT2 #(
		.INIT('h4)
	) name2452 (
		_w3436_,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('h1)
	) name2453 (
		_w3435_,
		_w3454_,
		_w3455_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		_w3426_,
		_w3455_,
		_w3456_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w3425_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h8)
	) name2456 (
		\A[427] ,
		\A[428] ,
		_w3458_
	);
	LUT2 #(
		.INIT('h1)
	) name2457 (
		\A[427] ,
		\A[428] ,
		_w3459_
	);
	LUT2 #(
		.INIT('h1)
	) name2458 (
		_w3458_,
		_w3459_,
		_w3460_
	);
	LUT2 #(
		.INIT('h8)
	) name2459 (
		\A[429] ,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h1)
	) name2460 (
		_w3458_,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		\A[430] ,
		\A[431] ,
		_w3463_
	);
	LUT2 #(
		.INIT('h1)
	) name2462 (
		\A[429] ,
		_w3460_,
		_w3464_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		_w3461_,
		_w3464_,
		_w3465_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		\A[430] ,
		\A[431] ,
		_w3466_
	);
	LUT2 #(
		.INIT('h1)
	) name2465 (
		_w3463_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h8)
	) name2466 (
		\A[432] ,
		_w3467_,
		_w3468_
	);
	LUT2 #(
		.INIT('h1)
	) name2467 (
		\A[432] ,
		_w3467_,
		_w3469_
	);
	LUT2 #(
		.INIT('h1)
	) name2468 (
		_w3468_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		_w3465_,
		_w3470_,
		_w3471_
	);
	LUT2 #(
		.INIT('h8)
	) name2470 (
		_w3463_,
		_w3471_,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name2471 (
		_w3463_,
		_w3468_,
		_w3473_
	);
	LUT2 #(
		.INIT('h4)
	) name2472 (
		_w3471_,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		_w3472_,
		_w3474_,
		_w3475_
	);
	LUT2 #(
		.INIT('h2)
	) name2474 (
		_w3462_,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h4)
	) name2475 (
		_w3462_,
		_w3475_,
		_w3477_
	);
	LUT2 #(
		.INIT('h1)
	) name2476 (
		_w3476_,
		_w3477_,
		_w3478_
	);
	LUT2 #(
		.INIT('h8)
	) name2477 (
		\A[433] ,
		\A[434] ,
		_w3479_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		\A[433] ,
		\A[434] ,
		_w3480_
	);
	LUT2 #(
		.INIT('h1)
	) name2479 (
		_w3479_,
		_w3480_,
		_w3481_
	);
	LUT2 #(
		.INIT('h8)
	) name2480 (
		\A[435] ,
		_w3481_,
		_w3482_
	);
	LUT2 #(
		.INIT('h1)
	) name2481 (
		\A[435] ,
		_w3481_,
		_w3483_
	);
	LUT2 #(
		.INIT('h1)
	) name2482 (
		_w3482_,
		_w3483_,
		_w3484_
	);
	LUT2 #(
		.INIT('h8)
	) name2483 (
		\A[436] ,
		\A[437] ,
		_w3485_
	);
	LUT2 #(
		.INIT('h1)
	) name2484 (
		\A[436] ,
		\A[437] ,
		_w3486_
	);
	LUT2 #(
		.INIT('h1)
	) name2485 (
		_w3485_,
		_w3486_,
		_w3487_
	);
	LUT2 #(
		.INIT('h8)
	) name2486 (
		\A[438] ,
		_w3487_,
		_w3488_
	);
	LUT2 #(
		.INIT('h1)
	) name2487 (
		\A[438] ,
		_w3487_,
		_w3489_
	);
	LUT2 #(
		.INIT('h1)
	) name2488 (
		_w3488_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('h8)
	) name2489 (
		_w3484_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h1)
	) name2490 (
		_w3485_,
		_w3488_,
		_w3492_
	);
	LUT2 #(
		.INIT('h1)
	) name2491 (
		_w3479_,
		_w3482_,
		_w3493_
	);
	LUT2 #(
		.INIT('h1)
	) name2492 (
		_w3492_,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h8)
	) name2493 (
		_w3492_,
		_w3493_,
		_w3495_
	);
	LUT2 #(
		.INIT('h1)
	) name2494 (
		_w3494_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h4)
	) name2495 (
		_w3491_,
		_w3496_,
		_w3497_
	);
	LUT2 #(
		.INIT('h1)
	) name2496 (
		_w3465_,
		_w3470_,
		_w3498_
	);
	LUT2 #(
		.INIT('h1)
	) name2497 (
		_w3471_,
		_w3498_,
		_w3499_
	);
	LUT2 #(
		.INIT('h1)
	) name2498 (
		_w3484_,
		_w3490_,
		_w3500_
	);
	LUT2 #(
		.INIT('h1)
	) name2499 (
		_w3491_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h8)
	) name2500 (
		_w3499_,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h2)
	) name2501 (
		_w3491_,
		_w3496_,
		_w3503_
	);
	LUT2 #(
		.INIT('h1)
	) name2502 (
		_w3497_,
		_w3502_,
		_w3504_
	);
	LUT2 #(
		.INIT('h4)
	) name2503 (
		_w3503_,
		_w3504_,
		_w3505_
	);
	LUT2 #(
		.INIT('h2)
	) name2504 (
		_w3478_,
		_w3505_,
		_w3506_
	);
	LUT2 #(
		.INIT('h8)
	) name2505 (
		_w3496_,
		_w3502_,
		_w3507_
	);
	LUT2 #(
		.INIT('h4)
	) name2506 (
		_w3462_,
		_w3472_,
		_w3508_
	);
	LUT2 #(
		.INIT('h2)
	) name2507 (
		_w3507_,
		_w3508_,
		_w3509_
	);
	LUT2 #(
		.INIT('h1)
	) name2508 (
		_w3506_,
		_w3509_,
		_w3510_
	);
	LUT2 #(
		.INIT('h4)
	) name2509 (
		_w3485_,
		_w3493_,
		_w3511_
	);
	LUT2 #(
		.INIT('h2)
	) name2510 (
		_w3491_,
		_w3511_,
		_w3512_
	);
	LUT2 #(
		.INIT('h1)
	) name2511 (
		_w3494_,
		_w3512_,
		_w3513_
	);
	LUT2 #(
		.INIT('h1)
	) name2512 (
		_w3510_,
		_w3513_,
		_w3514_
	);
	LUT2 #(
		.INIT('h1)
	) name2513 (
		_w3462_,
		_w3474_,
		_w3515_
	);
	LUT2 #(
		.INIT('h1)
	) name2514 (
		_w3472_,
		_w3515_,
		_w3516_
	);
	LUT2 #(
		.INIT('h8)
	) name2515 (
		_w3510_,
		_w3513_,
		_w3517_
	);
	LUT2 #(
		.INIT('h1)
	) name2516 (
		_w3516_,
		_w3517_,
		_w3518_
	);
	LUT2 #(
		.INIT('h1)
	) name2517 (
		_w3514_,
		_w3518_,
		_w3519_
	);
	LUT2 #(
		.INIT('h8)
	) name2518 (
		\A[421] ,
		\A[422] ,
		_w3520_
	);
	LUT2 #(
		.INIT('h1)
	) name2519 (
		\A[421] ,
		\A[422] ,
		_w3521_
	);
	LUT2 #(
		.INIT('h1)
	) name2520 (
		_w3520_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h8)
	) name2521 (
		\A[423] ,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h1)
	) name2522 (
		\A[423] ,
		_w3522_,
		_w3524_
	);
	LUT2 #(
		.INIT('h1)
	) name2523 (
		_w3523_,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h8)
	) name2524 (
		\A[424] ,
		\A[425] ,
		_w3526_
	);
	LUT2 #(
		.INIT('h1)
	) name2525 (
		\A[424] ,
		\A[425] ,
		_w3527_
	);
	LUT2 #(
		.INIT('h1)
	) name2526 (
		_w3526_,
		_w3527_,
		_w3528_
	);
	LUT2 #(
		.INIT('h8)
	) name2527 (
		\A[426] ,
		_w3528_,
		_w3529_
	);
	LUT2 #(
		.INIT('h1)
	) name2528 (
		\A[426] ,
		_w3528_,
		_w3530_
	);
	LUT2 #(
		.INIT('h1)
	) name2529 (
		_w3529_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h8)
	) name2530 (
		_w3525_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name2531 (
		_w3525_,
		_w3531_,
		_w3533_
	);
	LUT2 #(
		.INIT('h1)
	) name2532 (
		_w3532_,
		_w3533_,
		_w3534_
	);
	LUT2 #(
		.INIT('h8)
	) name2533 (
		\A[415] ,
		\A[416] ,
		_w3535_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		\A[415] ,
		\A[416] ,
		_w3536_
	);
	LUT2 #(
		.INIT('h1)
	) name2535 (
		_w3535_,
		_w3536_,
		_w3537_
	);
	LUT2 #(
		.INIT('h8)
	) name2536 (
		\A[417] ,
		_w3537_,
		_w3538_
	);
	LUT2 #(
		.INIT('h1)
	) name2537 (
		\A[417] ,
		_w3537_,
		_w3539_
	);
	LUT2 #(
		.INIT('h1)
	) name2538 (
		_w3538_,
		_w3539_,
		_w3540_
	);
	LUT2 #(
		.INIT('h8)
	) name2539 (
		\A[418] ,
		\A[419] ,
		_w3541_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		\A[418] ,
		\A[419] ,
		_w3542_
	);
	LUT2 #(
		.INIT('h1)
	) name2541 (
		_w3541_,
		_w3542_,
		_w3543_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		\A[420] ,
		_w3543_,
		_w3544_
	);
	LUT2 #(
		.INIT('h1)
	) name2543 (
		\A[420] ,
		_w3543_,
		_w3545_
	);
	LUT2 #(
		.INIT('h1)
	) name2544 (
		_w3544_,
		_w3545_,
		_w3546_
	);
	LUT2 #(
		.INIT('h8)
	) name2545 (
		_w3540_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h1)
	) name2546 (
		_w3540_,
		_w3546_,
		_w3548_
	);
	LUT2 #(
		.INIT('h1)
	) name2547 (
		_w3547_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h8)
	) name2548 (
		_w3534_,
		_w3549_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name2549 (
		_w3526_,
		_w3529_,
		_w3551_
	);
	LUT2 #(
		.INIT('h1)
	) name2550 (
		_w3520_,
		_w3523_,
		_w3552_
	);
	LUT2 #(
		.INIT('h1)
	) name2551 (
		_w3551_,
		_w3552_,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name2552 (
		_w3551_,
		_w3552_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name2553 (
		_w3553_,
		_w3554_,
		_w3555_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		_w3550_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name2555 (
		_w3541_,
		_w3544_,
		_w3557_
	);
	LUT2 #(
		.INIT('h1)
	) name2556 (
		_w3535_,
		_w3538_,
		_w3558_
	);
	LUT2 #(
		.INIT('h8)
	) name2557 (
		_w3557_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h1)
	) name2558 (
		_w3557_,
		_w3558_,
		_w3560_
	);
	LUT2 #(
		.INIT('h1)
	) name2559 (
		_w3559_,
		_w3560_,
		_w3561_
	);
	LUT2 #(
		.INIT('h2)
	) name2560 (
		_w3547_,
		_w3561_,
		_w3562_
	);
	LUT2 #(
		.INIT('h4)
	) name2561 (
		_w3547_,
		_w3561_,
		_w3563_
	);
	LUT2 #(
		.INIT('h1)
	) name2562 (
		_w3562_,
		_w3563_,
		_w3564_
	);
	LUT2 #(
		.INIT('h4)
	) name2563 (
		_w3556_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h4)
	) name2564 (
		_w3532_,
		_w3555_,
		_w3566_
	);
	LUT2 #(
		.INIT('h2)
	) name2565 (
		_w3532_,
		_w3555_,
		_w3567_
	);
	LUT2 #(
		.INIT('h1)
	) name2566 (
		_w3550_,
		_w3566_,
		_w3568_
	);
	LUT2 #(
		.INIT('h4)
	) name2567 (
		_w3567_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h1)
	) name2568 (
		_w3565_,
		_w3569_,
		_w3570_
	);
	LUT2 #(
		.INIT('h1)
	) name2569 (
		_w3532_,
		_w3553_,
		_w3571_
	);
	LUT2 #(
		.INIT('h1)
	) name2570 (
		_w3554_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h1)
	) name2571 (
		_w3570_,
		_w3572_,
		_w3573_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		_w3570_,
		_w3572_,
		_w3574_
	);
	LUT2 #(
		.INIT('h1)
	) name2573 (
		_w3547_,
		_w3560_,
		_w3575_
	);
	LUT2 #(
		.INIT('h1)
	) name2574 (
		_w3559_,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h1)
	) name2575 (
		_w3574_,
		_w3576_,
		_w3577_
	);
	LUT2 #(
		.INIT('h1)
	) name2576 (
		_w3573_,
		_w3577_,
		_w3578_
	);
	LUT2 #(
		.INIT('h4)
	) name2577 (
		_w3519_,
		_w3578_,
		_w3579_
	);
	LUT2 #(
		.INIT('h2)
	) name2578 (
		_w3519_,
		_w3578_,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w3514_,
		_w3517_,
		_w3581_
	);
	LUT2 #(
		.INIT('h2)
	) name2580 (
		_w3516_,
		_w3581_,
		_w3582_
	);
	LUT2 #(
		.INIT('h4)
	) name2581 (
		_w3516_,
		_w3581_,
		_w3583_
	);
	LUT2 #(
		.INIT('h1)
	) name2582 (
		_w3582_,
		_w3583_,
		_w3584_
	);
	LUT2 #(
		.INIT('h1)
	) name2583 (
		_w3573_,
		_w3574_,
		_w3585_
	);
	LUT2 #(
		.INIT('h4)
	) name2584 (
		_w3576_,
		_w3585_,
		_w3586_
	);
	LUT2 #(
		.INIT('h2)
	) name2585 (
		_w3576_,
		_w3585_,
		_w3587_
	);
	LUT2 #(
		.INIT('h1)
	) name2586 (
		_w3586_,
		_w3587_,
		_w3588_
	);
	LUT2 #(
		.INIT('h2)
	) name2587 (
		_w3584_,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h4)
	) name2588 (
		_w3584_,
		_w3588_,
		_w3590_
	);
	LUT2 #(
		.INIT('h1)
	) name2589 (
		_w3499_,
		_w3501_,
		_w3591_
	);
	LUT2 #(
		.INIT('h1)
	) name2590 (
		_w3502_,
		_w3591_,
		_w3592_
	);
	LUT2 #(
		.INIT('h1)
	) name2591 (
		_w3534_,
		_w3549_,
		_w3593_
	);
	LUT2 #(
		.INIT('h1)
	) name2592 (
		_w3550_,
		_w3593_,
		_w3594_
	);
	LUT2 #(
		.INIT('h8)
	) name2593 (
		_w3592_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h2)
	) name2594 (
		_w3506_,
		_w3509_,
		_w3596_
	);
	LUT2 #(
		.INIT('h1)
	) name2595 (
		_w3505_,
		_w3507_,
		_w3597_
	);
	LUT2 #(
		.INIT('h1)
	) name2596 (
		_w3478_,
		_w3597_,
		_w3598_
	);
	LUT2 #(
		.INIT('h1)
	) name2597 (
		_w3596_,
		_w3598_,
		_w3599_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		_w3595_,
		_w3599_,
		_w3600_
	);
	LUT2 #(
		.INIT('h1)
	) name2599 (
		_w3595_,
		_w3599_,
		_w3601_
	);
	LUT2 #(
		.INIT('h1)
	) name2600 (
		_w3556_,
		_w3569_,
		_w3602_
	);
	LUT2 #(
		.INIT('h8)
	) name2601 (
		_w3564_,
		_w3602_,
		_w3603_
	);
	LUT2 #(
		.INIT('h1)
	) name2602 (
		_w3564_,
		_w3602_,
		_w3604_
	);
	LUT2 #(
		.INIT('h1)
	) name2603 (
		_w3603_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h1)
	) name2604 (
		_w3601_,
		_w3605_,
		_w3606_
	);
	LUT2 #(
		.INIT('h1)
	) name2605 (
		_w3600_,
		_w3606_,
		_w3607_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w3590_,
		_w3607_,
		_w3608_
	);
	LUT2 #(
		.INIT('h1)
	) name2607 (
		_w3589_,
		_w3608_,
		_w3609_
	);
	LUT2 #(
		.INIT('h1)
	) name2608 (
		_w3580_,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h1)
	) name2609 (
		_w3579_,
		_w3610_,
		_w3611_
	);
	LUT2 #(
		.INIT('h1)
	) name2610 (
		_w3457_,
		_w3611_,
		_w3612_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		_w3457_,
		_w3611_,
		_w3613_
	);
	LUT2 #(
		.INIT('h1)
	) name2612 (
		_w3425_,
		_w3426_,
		_w3614_
	);
	LUT2 #(
		.INIT('h4)
	) name2613 (
		_w3455_,
		_w3614_,
		_w3615_
	);
	LUT2 #(
		.INIT('h2)
	) name2614 (
		_w3455_,
		_w3614_,
		_w3616_
	);
	LUT2 #(
		.INIT('h1)
	) name2615 (
		_w3615_,
		_w3616_,
		_w3617_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		_w3579_,
		_w3580_,
		_w3618_
	);
	LUT2 #(
		.INIT('h4)
	) name2617 (
		_w3609_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h2)
	) name2618 (
		_w3609_,
		_w3618_,
		_w3620_
	);
	LUT2 #(
		.INIT('h1)
	) name2619 (
		_w3619_,
		_w3620_,
		_w3621_
	);
	LUT2 #(
		.INIT('h1)
	) name2620 (
		_w3617_,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h8)
	) name2621 (
		_w3617_,
		_w3621_,
		_w3623_
	);
	LUT2 #(
		.INIT('h1)
	) name2622 (
		_w3589_,
		_w3590_,
		_w3624_
	);
	LUT2 #(
		.INIT('h4)
	) name2623 (
		_w3607_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('h2)
	) name2624 (
		_w3607_,
		_w3624_,
		_w3626_
	);
	LUT2 #(
		.INIT('h1)
	) name2625 (
		_w3625_,
		_w3626_,
		_w3627_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		_w3435_,
		_w3436_,
		_w3628_
	);
	LUT2 #(
		.INIT('h8)
	) name2627 (
		_w3453_,
		_w3628_,
		_w3629_
	);
	LUT2 #(
		.INIT('h1)
	) name2628 (
		_w3453_,
		_w3628_,
		_w3630_
	);
	LUT2 #(
		.INIT('h1)
	) name2629 (
		_w3629_,
		_w3630_,
		_w3631_
	);
	LUT2 #(
		.INIT('h8)
	) name2630 (
		_w3627_,
		_w3631_,
		_w3632_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w3627_,
		_w3631_,
		_w3633_
	);
	LUT2 #(
		.INIT('h1)
	) name2632 (
		_w3438_,
		_w3440_,
		_w3634_
	);
	LUT2 #(
		.INIT('h1)
	) name2633 (
		_w3441_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name2634 (
		_w3592_,
		_w3594_,
		_w3636_
	);
	LUT2 #(
		.INIT('h1)
	) name2635 (
		_w3595_,
		_w3636_,
		_w3637_
	);
	LUT2 #(
		.INIT('h8)
	) name2636 (
		_w3635_,
		_w3637_,
		_w3638_
	);
	LUT2 #(
		.INIT('h1)
	) name2637 (
		_w3446_,
		_w3451_,
		_w3639_
	);
	LUT2 #(
		.INIT('h2)
	) name2638 (
		_w3450_,
		_w3639_,
		_w3640_
	);
	LUT2 #(
		.INIT('h4)
	) name2639 (
		_w3450_,
		_w3639_,
		_w3641_
	);
	LUT2 #(
		.INIT('h1)
	) name2640 (
		_w3640_,
		_w3641_,
		_w3642_
	);
	LUT2 #(
		.INIT('h2)
	) name2641 (
		_w3638_,
		_w3642_,
		_w3643_
	);
	LUT2 #(
		.INIT('h4)
	) name2642 (
		_w3638_,
		_w3642_,
		_w3644_
	);
	LUT2 #(
		.INIT('h1)
	) name2643 (
		_w3600_,
		_w3601_,
		_w3645_
	);
	LUT2 #(
		.INIT('h4)
	) name2644 (
		_w3605_,
		_w3645_,
		_w3646_
	);
	LUT2 #(
		.INIT('h2)
	) name2645 (
		_w3605_,
		_w3645_,
		_w3647_
	);
	LUT2 #(
		.INIT('h1)
	) name2646 (
		_w3646_,
		_w3647_,
		_w3648_
	);
	LUT2 #(
		.INIT('h4)
	) name2647 (
		_w3644_,
		_w3648_,
		_w3649_
	);
	LUT2 #(
		.INIT('h1)
	) name2648 (
		_w3643_,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h1)
	) name2649 (
		_w3633_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h1)
	) name2650 (
		_w3632_,
		_w3651_,
		_w3652_
	);
	LUT2 #(
		.INIT('h4)
	) name2651 (
		_w3623_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h1)
	) name2652 (
		_w3622_,
		_w3653_,
		_w3654_
	);
	LUT2 #(
		.INIT('h4)
	) name2653 (
		_w3613_,
		_w3654_,
		_w3655_
	);
	LUT2 #(
		.INIT('h1)
	) name2654 (
		_w3612_,
		_w3655_,
		_w3656_
	);
	LUT2 #(
		.INIT('h1)
	) name2655 (
		_w3299_,
		_w3656_,
		_w3657_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		_w3299_,
		_w3656_,
		_w3658_
	);
	LUT2 #(
		.INIT('h1)
	) name2657 (
		_w3612_,
		_w3613_,
		_w3659_
	);
	LUT2 #(
		.INIT('h4)
	) name2658 (
		_w3654_,
		_w3659_,
		_w3660_
	);
	LUT2 #(
		.INIT('h2)
	) name2659 (
		_w3654_,
		_w3659_,
		_w3661_
	);
	LUT2 #(
		.INIT('h1)
	) name2660 (
		_w3660_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h1)
	) name2661 (
		_w3255_,
		_w3256_,
		_w3663_
	);
	LUT2 #(
		.INIT('h4)
	) name2662 (
		_w3297_,
		_w3663_,
		_w3664_
	);
	LUT2 #(
		.INIT('h2)
	) name2663 (
		_w3297_,
		_w3663_,
		_w3665_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		_w3664_,
		_w3665_,
		_w3666_
	);
	LUT2 #(
		.INIT('h2)
	) name2665 (
		_w3662_,
		_w3666_,
		_w3667_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		_w3662_,
		_w3666_,
		_w3668_
	);
	LUT2 #(
		.INIT('h1)
	) name2667 (
		_w3265_,
		_w3266_,
		_w3669_
	);
	LUT2 #(
		.INIT('h4)
	) name2668 (
		_w3295_,
		_w3669_,
		_w3670_
	);
	LUT2 #(
		.INIT('h2)
	) name2669 (
		_w3295_,
		_w3669_,
		_w3671_
	);
	LUT2 #(
		.INIT('h1)
	) name2670 (
		_w3670_,
		_w3671_,
		_w3672_
	);
	LUT2 #(
		.INIT('h1)
	) name2671 (
		_w3622_,
		_w3623_,
		_w3673_
	);
	LUT2 #(
		.INIT('h4)
	) name2672 (
		_w3652_,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h2)
	) name2673 (
		_w3652_,
		_w3673_,
		_w3675_
	);
	LUT2 #(
		.INIT('h1)
	) name2674 (
		_w3674_,
		_w3675_,
		_w3676_
	);
	LUT2 #(
		.INIT('h1)
	) name2675 (
		_w3672_,
		_w3676_,
		_w3677_
	);
	LUT2 #(
		.INIT('h8)
	) name2676 (
		_w3672_,
		_w3676_,
		_w3678_
	);
	LUT2 #(
		.INIT('h1)
	) name2677 (
		_w3275_,
		_w3276_,
		_w3679_
	);
	LUT2 #(
		.INIT('h4)
	) name2678 (
		_w3293_,
		_w3679_,
		_w3680_
	);
	LUT2 #(
		.INIT('h2)
	) name2679 (
		_w3293_,
		_w3679_,
		_w3681_
	);
	LUT2 #(
		.INIT('h1)
	) name2680 (
		_w3680_,
		_w3681_,
		_w3682_
	);
	LUT2 #(
		.INIT('h1)
	) name2681 (
		_w3632_,
		_w3633_,
		_w3683_
	);
	LUT2 #(
		.INIT('h4)
	) name2682 (
		_w3650_,
		_w3683_,
		_w3684_
	);
	LUT2 #(
		.INIT('h2)
	) name2683 (
		_w3650_,
		_w3683_,
		_w3685_
	);
	LUT2 #(
		.INIT('h1)
	) name2684 (
		_w3684_,
		_w3685_,
		_w3686_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		_w3682_,
		_w3686_,
		_w3687_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		_w3682_,
		_w3686_,
		_w3688_
	);
	LUT2 #(
		.INIT('h1)
	) name2687 (
		_w3635_,
		_w3637_,
		_w3689_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		_w3638_,
		_w3689_,
		_w3690_
	);
	LUT2 #(
		.INIT('h1)
	) name2689 (
		_w3278_,
		_w3280_,
		_w3691_
	);
	LUT2 #(
		.INIT('h1)
	) name2690 (
		_w3281_,
		_w3691_,
		_w3692_
	);
	LUT2 #(
		.INIT('h8)
	) name2691 (
		_w3690_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h1)
	) name2692 (
		_w3643_,
		_w3644_,
		_w3694_
	);
	LUT2 #(
		.INIT('h4)
	) name2693 (
		_w3648_,
		_w3694_,
		_w3695_
	);
	LUT2 #(
		.INIT('h2)
	) name2694 (
		_w3648_,
		_w3694_,
		_w3696_
	);
	LUT2 #(
		.INIT('h1)
	) name2695 (
		_w3695_,
		_w3696_,
		_w3697_
	);
	LUT2 #(
		.INIT('h2)
	) name2696 (
		_w3693_,
		_w3697_,
		_w3698_
	);
	LUT2 #(
		.INIT('h4)
	) name2697 (
		_w3693_,
		_w3697_,
		_w3699_
	);
	LUT2 #(
		.INIT('h1)
	) name2698 (
		_w3286_,
		_w3287_,
		_w3700_
	);
	LUT2 #(
		.INIT('h4)
	) name2699 (
		_w3291_,
		_w3700_,
		_w3701_
	);
	LUT2 #(
		.INIT('h2)
	) name2700 (
		_w3291_,
		_w3700_,
		_w3702_
	);
	LUT2 #(
		.INIT('h1)
	) name2701 (
		_w3701_,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h1)
	) name2702 (
		_w3699_,
		_w3703_,
		_w3704_
	);
	LUT2 #(
		.INIT('h1)
	) name2703 (
		_w3698_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h4)
	) name2704 (
		_w3688_,
		_w3705_,
		_w3706_
	);
	LUT2 #(
		.INIT('h1)
	) name2705 (
		_w3687_,
		_w3706_,
		_w3707_
	);
	LUT2 #(
		.INIT('h1)
	) name2706 (
		_w3678_,
		_w3707_,
		_w3708_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		_w3677_,
		_w3708_,
		_w3709_
	);
	LUT2 #(
		.INIT('h1)
	) name2708 (
		_w3668_,
		_w3709_,
		_w3710_
	);
	LUT2 #(
		.INIT('h1)
	) name2709 (
		_w3667_,
		_w3710_,
		_w3711_
	);
	LUT2 #(
		.INIT('h4)
	) name2710 (
		_w3658_,
		_w3711_,
		_w3712_
	);
	LUT2 #(
		.INIT('h1)
	) name2711 (
		_w3657_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h8)
	) name2712 (
		\A[355] ,
		\A[356] ,
		_w3714_
	);
	LUT2 #(
		.INIT('h1)
	) name2713 (
		\A[355] ,
		\A[356] ,
		_w3715_
	);
	LUT2 #(
		.INIT('h1)
	) name2714 (
		_w3714_,
		_w3715_,
		_w3716_
	);
	LUT2 #(
		.INIT('h8)
	) name2715 (
		\A[357] ,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h1)
	) name2716 (
		_w3714_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h8)
	) name2717 (
		\A[358] ,
		\A[359] ,
		_w3719_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		\A[357] ,
		_w3716_,
		_w3720_
	);
	LUT2 #(
		.INIT('h1)
	) name2719 (
		_w3717_,
		_w3720_,
		_w3721_
	);
	LUT2 #(
		.INIT('h1)
	) name2720 (
		\A[358] ,
		\A[359] ,
		_w3722_
	);
	LUT2 #(
		.INIT('h1)
	) name2721 (
		_w3719_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h8)
	) name2722 (
		\A[360] ,
		_w3723_,
		_w3724_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		\A[360] ,
		_w3723_,
		_w3725_
	);
	LUT2 #(
		.INIT('h1)
	) name2724 (
		_w3724_,
		_w3725_,
		_w3726_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		_w3721_,
		_w3726_,
		_w3727_
	);
	LUT2 #(
		.INIT('h8)
	) name2726 (
		_w3719_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h1)
	) name2727 (
		_w3719_,
		_w3724_,
		_w3729_
	);
	LUT2 #(
		.INIT('h4)
	) name2728 (
		_w3727_,
		_w3729_,
		_w3730_
	);
	LUT2 #(
		.INIT('h1)
	) name2729 (
		_w3728_,
		_w3730_,
		_w3731_
	);
	LUT2 #(
		.INIT('h2)
	) name2730 (
		_w3718_,
		_w3731_,
		_w3732_
	);
	LUT2 #(
		.INIT('h4)
	) name2731 (
		_w3718_,
		_w3731_,
		_w3733_
	);
	LUT2 #(
		.INIT('h1)
	) name2732 (
		_w3732_,
		_w3733_,
		_w3734_
	);
	LUT2 #(
		.INIT('h8)
	) name2733 (
		\A[361] ,
		\A[362] ,
		_w3735_
	);
	LUT2 #(
		.INIT('h1)
	) name2734 (
		\A[361] ,
		\A[362] ,
		_w3736_
	);
	LUT2 #(
		.INIT('h1)
	) name2735 (
		_w3735_,
		_w3736_,
		_w3737_
	);
	LUT2 #(
		.INIT('h8)
	) name2736 (
		\A[363] ,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h1)
	) name2737 (
		\A[363] ,
		_w3737_,
		_w3739_
	);
	LUT2 #(
		.INIT('h1)
	) name2738 (
		_w3738_,
		_w3739_,
		_w3740_
	);
	LUT2 #(
		.INIT('h8)
	) name2739 (
		\A[364] ,
		\A[365] ,
		_w3741_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		\A[364] ,
		\A[365] ,
		_w3742_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		_w3741_,
		_w3742_,
		_w3743_
	);
	LUT2 #(
		.INIT('h8)
	) name2742 (
		\A[366] ,
		_w3743_,
		_w3744_
	);
	LUT2 #(
		.INIT('h1)
	) name2743 (
		\A[366] ,
		_w3743_,
		_w3745_
	);
	LUT2 #(
		.INIT('h1)
	) name2744 (
		_w3744_,
		_w3745_,
		_w3746_
	);
	LUT2 #(
		.INIT('h8)
	) name2745 (
		_w3740_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h1)
	) name2746 (
		_w3741_,
		_w3744_,
		_w3748_
	);
	LUT2 #(
		.INIT('h1)
	) name2747 (
		_w3735_,
		_w3738_,
		_w3749_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w3748_,
		_w3749_,
		_w3750_
	);
	LUT2 #(
		.INIT('h8)
	) name2749 (
		_w3748_,
		_w3749_,
		_w3751_
	);
	LUT2 #(
		.INIT('h1)
	) name2750 (
		_w3750_,
		_w3751_,
		_w3752_
	);
	LUT2 #(
		.INIT('h4)
	) name2751 (
		_w3747_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		_w3721_,
		_w3726_,
		_w3754_
	);
	LUT2 #(
		.INIT('h1)
	) name2753 (
		_w3727_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('h1)
	) name2754 (
		_w3740_,
		_w3746_,
		_w3756_
	);
	LUT2 #(
		.INIT('h1)
	) name2755 (
		_w3747_,
		_w3756_,
		_w3757_
	);
	LUT2 #(
		.INIT('h8)
	) name2756 (
		_w3755_,
		_w3757_,
		_w3758_
	);
	LUT2 #(
		.INIT('h2)
	) name2757 (
		_w3747_,
		_w3752_,
		_w3759_
	);
	LUT2 #(
		.INIT('h1)
	) name2758 (
		_w3753_,
		_w3758_,
		_w3760_
	);
	LUT2 #(
		.INIT('h4)
	) name2759 (
		_w3759_,
		_w3760_,
		_w3761_
	);
	LUT2 #(
		.INIT('h2)
	) name2760 (
		_w3734_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h8)
	) name2761 (
		_w3752_,
		_w3758_,
		_w3763_
	);
	LUT2 #(
		.INIT('h4)
	) name2762 (
		_w3718_,
		_w3728_,
		_w3764_
	);
	LUT2 #(
		.INIT('h2)
	) name2763 (
		_w3763_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h1)
	) name2764 (
		_w3762_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('h4)
	) name2765 (
		_w3741_,
		_w3749_,
		_w3767_
	);
	LUT2 #(
		.INIT('h2)
	) name2766 (
		_w3747_,
		_w3767_,
		_w3768_
	);
	LUT2 #(
		.INIT('h1)
	) name2767 (
		_w3750_,
		_w3768_,
		_w3769_
	);
	LUT2 #(
		.INIT('h1)
	) name2768 (
		_w3766_,
		_w3769_,
		_w3770_
	);
	LUT2 #(
		.INIT('h1)
	) name2769 (
		_w3718_,
		_w3730_,
		_w3771_
	);
	LUT2 #(
		.INIT('h1)
	) name2770 (
		_w3728_,
		_w3771_,
		_w3772_
	);
	LUT2 #(
		.INIT('h8)
	) name2771 (
		_w3766_,
		_w3769_,
		_w3773_
	);
	LUT2 #(
		.INIT('h1)
	) name2772 (
		_w3772_,
		_w3773_,
		_w3774_
	);
	LUT2 #(
		.INIT('h1)
	) name2773 (
		_w3770_,
		_w3774_,
		_w3775_
	);
	LUT2 #(
		.INIT('h8)
	) name2774 (
		\A[349] ,
		\A[350] ,
		_w3776_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		\A[349] ,
		\A[350] ,
		_w3777_
	);
	LUT2 #(
		.INIT('h1)
	) name2776 (
		_w3776_,
		_w3777_,
		_w3778_
	);
	LUT2 #(
		.INIT('h8)
	) name2777 (
		\A[351] ,
		_w3778_,
		_w3779_
	);
	LUT2 #(
		.INIT('h1)
	) name2778 (
		\A[351] ,
		_w3778_,
		_w3780_
	);
	LUT2 #(
		.INIT('h1)
	) name2779 (
		_w3779_,
		_w3780_,
		_w3781_
	);
	LUT2 #(
		.INIT('h8)
	) name2780 (
		\A[352] ,
		\A[353] ,
		_w3782_
	);
	LUT2 #(
		.INIT('h1)
	) name2781 (
		\A[352] ,
		\A[353] ,
		_w3783_
	);
	LUT2 #(
		.INIT('h1)
	) name2782 (
		_w3782_,
		_w3783_,
		_w3784_
	);
	LUT2 #(
		.INIT('h8)
	) name2783 (
		\A[354] ,
		_w3784_,
		_w3785_
	);
	LUT2 #(
		.INIT('h1)
	) name2784 (
		\A[354] ,
		_w3784_,
		_w3786_
	);
	LUT2 #(
		.INIT('h1)
	) name2785 (
		_w3785_,
		_w3786_,
		_w3787_
	);
	LUT2 #(
		.INIT('h8)
	) name2786 (
		_w3781_,
		_w3787_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name2787 (
		_w3781_,
		_w3787_,
		_w3789_
	);
	LUT2 #(
		.INIT('h1)
	) name2788 (
		_w3788_,
		_w3789_,
		_w3790_
	);
	LUT2 #(
		.INIT('h8)
	) name2789 (
		\A[343] ,
		\A[344] ,
		_w3791_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		\A[343] ,
		\A[344] ,
		_w3792_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		_w3791_,
		_w3792_,
		_w3793_
	);
	LUT2 #(
		.INIT('h8)
	) name2792 (
		\A[345] ,
		_w3793_,
		_w3794_
	);
	LUT2 #(
		.INIT('h1)
	) name2793 (
		\A[345] ,
		_w3793_,
		_w3795_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		_w3794_,
		_w3795_,
		_w3796_
	);
	LUT2 #(
		.INIT('h8)
	) name2795 (
		\A[346] ,
		\A[347] ,
		_w3797_
	);
	LUT2 #(
		.INIT('h1)
	) name2796 (
		\A[346] ,
		\A[347] ,
		_w3798_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		_w3797_,
		_w3798_,
		_w3799_
	);
	LUT2 #(
		.INIT('h8)
	) name2798 (
		\A[348] ,
		_w3799_,
		_w3800_
	);
	LUT2 #(
		.INIT('h1)
	) name2799 (
		\A[348] ,
		_w3799_,
		_w3801_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w3800_,
		_w3801_,
		_w3802_
	);
	LUT2 #(
		.INIT('h8)
	) name2801 (
		_w3796_,
		_w3802_,
		_w3803_
	);
	LUT2 #(
		.INIT('h1)
	) name2802 (
		_w3796_,
		_w3802_,
		_w3804_
	);
	LUT2 #(
		.INIT('h1)
	) name2803 (
		_w3803_,
		_w3804_,
		_w3805_
	);
	LUT2 #(
		.INIT('h8)
	) name2804 (
		_w3790_,
		_w3805_,
		_w3806_
	);
	LUT2 #(
		.INIT('h1)
	) name2805 (
		_w3776_,
		_w3779_,
		_w3807_
	);
	LUT2 #(
		.INIT('h1)
	) name2806 (
		_w3782_,
		_w3785_,
		_w3808_
	);
	LUT2 #(
		.INIT('h4)
	) name2807 (
		_w3788_,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h8)
	) name2808 (
		_w3782_,
		_w3788_,
		_w3810_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		_w3809_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h2)
	) name2810 (
		_w3807_,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h4)
	) name2811 (
		_w3807_,
		_w3811_,
		_w3813_
	);
	LUT2 #(
		.INIT('h1)
	) name2812 (
		_w3812_,
		_w3813_,
		_w3814_
	);
	LUT2 #(
		.INIT('h1)
	) name2813 (
		_w3806_,
		_w3814_,
		_w3815_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		_w3791_,
		_w3794_,
		_w3816_
	);
	LUT2 #(
		.INIT('h8)
	) name2815 (
		_w3797_,
		_w3803_,
		_w3817_
	);
	LUT2 #(
		.INIT('h1)
	) name2816 (
		_w3797_,
		_w3800_,
		_w3818_
	);
	LUT2 #(
		.INIT('h4)
	) name2817 (
		_w3803_,
		_w3818_,
		_w3819_
	);
	LUT2 #(
		.INIT('h1)
	) name2818 (
		_w3817_,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h2)
	) name2819 (
		_w3816_,
		_w3820_,
		_w3821_
	);
	LUT2 #(
		.INIT('h4)
	) name2820 (
		_w3816_,
		_w3820_,
		_w3822_
	);
	LUT2 #(
		.INIT('h1)
	) name2821 (
		_w3821_,
		_w3822_,
		_w3823_
	);
	LUT2 #(
		.INIT('h4)
	) name2822 (
		_w3815_,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h8)
	) name2823 (
		_w3806_,
		_w3814_,
		_w3825_
	);
	LUT2 #(
		.INIT('h1)
	) name2824 (
		_w3807_,
		_w3808_,
		_w3826_
	);
	LUT2 #(
		.INIT('h4)
	) name2825 (
		_w3816_,
		_w3817_,
		_w3827_
	);
	LUT2 #(
		.INIT('h1)
	) name2826 (
		_w3826_,
		_w3827_,
		_w3828_
	);
	LUT2 #(
		.INIT('h8)
	) name2827 (
		_w3825_,
		_w3828_,
		_w3829_
	);
	LUT2 #(
		.INIT('h1)
	) name2828 (
		_w3824_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h1)
	) name2829 (
		_w3807_,
		_w3809_,
		_w3831_
	);
	LUT2 #(
		.INIT('h1)
	) name2830 (
		_w3810_,
		_w3831_,
		_w3832_
	);
	LUT2 #(
		.INIT('h1)
	) name2831 (
		_w3830_,
		_w3832_,
		_w3833_
	);
	LUT2 #(
		.INIT('h1)
	) name2832 (
		_w3816_,
		_w3819_,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name2833 (
		_w3817_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h8)
	) name2834 (
		_w3830_,
		_w3832_,
		_w3836_
	);
	LUT2 #(
		.INIT('h1)
	) name2835 (
		_w3835_,
		_w3836_,
		_w3837_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		_w3833_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h1)
	) name2837 (
		_w3775_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h8)
	) name2838 (
		_w3775_,
		_w3838_,
		_w3840_
	);
	LUT2 #(
		.INIT('h1)
	) name2839 (
		_w3833_,
		_w3836_,
		_w3841_
	);
	LUT2 #(
		.INIT('h2)
	) name2840 (
		_w3835_,
		_w3841_,
		_w3842_
	);
	LUT2 #(
		.INIT('h4)
	) name2841 (
		_w3835_,
		_w3841_,
		_w3843_
	);
	LUT2 #(
		.INIT('h1)
	) name2842 (
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h1)
	) name2843 (
		_w3770_,
		_w3773_,
		_w3845_
	);
	LUT2 #(
		.INIT('h2)
	) name2844 (
		_w3772_,
		_w3845_,
		_w3846_
	);
	LUT2 #(
		.INIT('h4)
	) name2845 (
		_w3772_,
		_w3845_,
		_w3847_
	);
	LUT2 #(
		.INIT('h1)
	) name2846 (
		_w3846_,
		_w3847_,
		_w3848_
	);
	LUT2 #(
		.INIT('h1)
	) name2847 (
		_w3844_,
		_w3848_,
		_w3849_
	);
	LUT2 #(
		.INIT('h1)
	) name2848 (
		_w3755_,
		_w3757_,
		_w3850_
	);
	LUT2 #(
		.INIT('h1)
	) name2849 (
		_w3758_,
		_w3850_,
		_w3851_
	);
	LUT2 #(
		.INIT('h1)
	) name2850 (
		_w3790_,
		_w3805_,
		_w3852_
	);
	LUT2 #(
		.INIT('h1)
	) name2851 (
		_w3806_,
		_w3852_,
		_w3853_
	);
	LUT2 #(
		.INIT('h8)
	) name2852 (
		_w3851_,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h2)
	) name2853 (
		_w3762_,
		_w3765_,
		_w3855_
	);
	LUT2 #(
		.INIT('h1)
	) name2854 (
		_w3761_,
		_w3763_,
		_w3856_
	);
	LUT2 #(
		.INIT('h1)
	) name2855 (
		_w3734_,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('h1)
	) name2856 (
		_w3855_,
		_w3857_,
		_w3858_
	);
	LUT2 #(
		.INIT('h1)
	) name2857 (
		_w3854_,
		_w3858_,
		_w3859_
	);
	LUT2 #(
		.INIT('h2)
	) name2858 (
		_w3824_,
		_w3829_,
		_w3860_
	);
	LUT2 #(
		.INIT('h1)
	) name2859 (
		_w3815_,
		_w3825_,
		_w3861_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w3823_,
		_w3861_,
		_w3862_
	);
	LUT2 #(
		.INIT('h1)
	) name2861 (
		_w3860_,
		_w3862_,
		_w3863_
	);
	LUT2 #(
		.INIT('h8)
	) name2862 (
		_w3854_,
		_w3858_,
		_w3864_
	);
	LUT2 #(
		.INIT('h1)
	) name2863 (
		_w3863_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h1)
	) name2864 (
		_w3859_,
		_w3865_,
		_w3866_
	);
	LUT2 #(
		.INIT('h8)
	) name2865 (
		_w3844_,
		_w3848_,
		_w3867_
	);
	LUT2 #(
		.INIT('h1)
	) name2866 (
		_w3866_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h1)
	) name2867 (
		_w3849_,
		_w3868_,
		_w3869_
	);
	LUT2 #(
		.INIT('h4)
	) name2868 (
		_w3840_,
		_w3869_,
		_w3870_
	);
	LUT2 #(
		.INIT('h1)
	) name2869 (
		_w3839_,
		_w3870_,
		_w3871_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		\A[331] ,
		\A[332] ,
		_w3872_
	);
	LUT2 #(
		.INIT('h1)
	) name2871 (
		\A[331] ,
		\A[332] ,
		_w3873_
	);
	LUT2 #(
		.INIT('h1)
	) name2872 (
		_w3872_,
		_w3873_,
		_w3874_
	);
	LUT2 #(
		.INIT('h8)
	) name2873 (
		\A[333] ,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h1)
	) name2874 (
		_w3872_,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h8)
	) name2875 (
		\A[334] ,
		\A[335] ,
		_w3877_
	);
	LUT2 #(
		.INIT('h1)
	) name2876 (
		\A[333] ,
		_w3874_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		_w3875_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h1)
	) name2878 (
		\A[334] ,
		\A[335] ,
		_w3880_
	);
	LUT2 #(
		.INIT('h1)
	) name2879 (
		_w3877_,
		_w3880_,
		_w3881_
	);
	LUT2 #(
		.INIT('h8)
	) name2880 (
		\A[336] ,
		_w3881_,
		_w3882_
	);
	LUT2 #(
		.INIT('h1)
	) name2881 (
		\A[336] ,
		_w3881_,
		_w3883_
	);
	LUT2 #(
		.INIT('h1)
	) name2882 (
		_w3882_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('h8)
	) name2883 (
		_w3879_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h8)
	) name2884 (
		_w3877_,
		_w3885_,
		_w3886_
	);
	LUT2 #(
		.INIT('h1)
	) name2885 (
		_w3877_,
		_w3882_,
		_w3887_
	);
	LUT2 #(
		.INIT('h4)
	) name2886 (
		_w3885_,
		_w3887_,
		_w3888_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		_w3886_,
		_w3888_,
		_w3889_
	);
	LUT2 #(
		.INIT('h2)
	) name2888 (
		_w3876_,
		_w3889_,
		_w3890_
	);
	LUT2 #(
		.INIT('h4)
	) name2889 (
		_w3876_,
		_w3889_,
		_w3891_
	);
	LUT2 #(
		.INIT('h1)
	) name2890 (
		_w3890_,
		_w3891_,
		_w3892_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		\A[337] ,
		\A[338] ,
		_w3893_
	);
	LUT2 #(
		.INIT('h1)
	) name2892 (
		\A[337] ,
		\A[338] ,
		_w3894_
	);
	LUT2 #(
		.INIT('h1)
	) name2893 (
		_w3893_,
		_w3894_,
		_w3895_
	);
	LUT2 #(
		.INIT('h8)
	) name2894 (
		\A[339] ,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h1)
	) name2895 (
		\A[339] ,
		_w3895_,
		_w3897_
	);
	LUT2 #(
		.INIT('h1)
	) name2896 (
		_w3896_,
		_w3897_,
		_w3898_
	);
	LUT2 #(
		.INIT('h8)
	) name2897 (
		\A[340] ,
		\A[341] ,
		_w3899_
	);
	LUT2 #(
		.INIT('h1)
	) name2898 (
		\A[340] ,
		\A[341] ,
		_w3900_
	);
	LUT2 #(
		.INIT('h1)
	) name2899 (
		_w3899_,
		_w3900_,
		_w3901_
	);
	LUT2 #(
		.INIT('h8)
	) name2900 (
		\A[342] ,
		_w3901_,
		_w3902_
	);
	LUT2 #(
		.INIT('h1)
	) name2901 (
		\A[342] ,
		_w3901_,
		_w3903_
	);
	LUT2 #(
		.INIT('h1)
	) name2902 (
		_w3902_,
		_w3903_,
		_w3904_
	);
	LUT2 #(
		.INIT('h8)
	) name2903 (
		_w3898_,
		_w3904_,
		_w3905_
	);
	LUT2 #(
		.INIT('h1)
	) name2904 (
		_w3899_,
		_w3902_,
		_w3906_
	);
	LUT2 #(
		.INIT('h1)
	) name2905 (
		_w3893_,
		_w3896_,
		_w3907_
	);
	LUT2 #(
		.INIT('h1)
	) name2906 (
		_w3906_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h8)
	) name2907 (
		_w3906_,
		_w3907_,
		_w3909_
	);
	LUT2 #(
		.INIT('h1)
	) name2908 (
		_w3908_,
		_w3909_,
		_w3910_
	);
	LUT2 #(
		.INIT('h4)
	) name2909 (
		_w3905_,
		_w3910_,
		_w3911_
	);
	LUT2 #(
		.INIT('h1)
	) name2910 (
		_w3879_,
		_w3884_,
		_w3912_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		_w3885_,
		_w3912_,
		_w3913_
	);
	LUT2 #(
		.INIT('h1)
	) name2912 (
		_w3898_,
		_w3904_,
		_w3914_
	);
	LUT2 #(
		.INIT('h1)
	) name2913 (
		_w3905_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('h8)
	) name2914 (
		_w3913_,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('h2)
	) name2915 (
		_w3905_,
		_w3910_,
		_w3917_
	);
	LUT2 #(
		.INIT('h1)
	) name2916 (
		_w3911_,
		_w3916_,
		_w3918_
	);
	LUT2 #(
		.INIT('h4)
	) name2917 (
		_w3917_,
		_w3918_,
		_w3919_
	);
	LUT2 #(
		.INIT('h2)
	) name2918 (
		_w3892_,
		_w3919_,
		_w3920_
	);
	LUT2 #(
		.INIT('h8)
	) name2919 (
		_w3910_,
		_w3916_,
		_w3921_
	);
	LUT2 #(
		.INIT('h4)
	) name2920 (
		_w3876_,
		_w3886_,
		_w3922_
	);
	LUT2 #(
		.INIT('h2)
	) name2921 (
		_w3921_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h1)
	) name2922 (
		_w3920_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('h4)
	) name2923 (
		_w3899_,
		_w3907_,
		_w3925_
	);
	LUT2 #(
		.INIT('h2)
	) name2924 (
		_w3905_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('h1)
	) name2925 (
		_w3908_,
		_w3926_,
		_w3927_
	);
	LUT2 #(
		.INIT('h1)
	) name2926 (
		_w3924_,
		_w3927_,
		_w3928_
	);
	LUT2 #(
		.INIT('h1)
	) name2927 (
		_w3876_,
		_w3888_,
		_w3929_
	);
	LUT2 #(
		.INIT('h1)
	) name2928 (
		_w3886_,
		_w3929_,
		_w3930_
	);
	LUT2 #(
		.INIT('h8)
	) name2929 (
		_w3924_,
		_w3927_,
		_w3931_
	);
	LUT2 #(
		.INIT('h1)
	) name2930 (
		_w3930_,
		_w3931_,
		_w3932_
	);
	LUT2 #(
		.INIT('h1)
	) name2931 (
		_w3928_,
		_w3932_,
		_w3933_
	);
	LUT2 #(
		.INIT('h8)
	) name2932 (
		\A[325] ,
		\A[326] ,
		_w3934_
	);
	LUT2 #(
		.INIT('h1)
	) name2933 (
		\A[325] ,
		\A[326] ,
		_w3935_
	);
	LUT2 #(
		.INIT('h1)
	) name2934 (
		_w3934_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h8)
	) name2935 (
		\A[327] ,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h1)
	) name2936 (
		\A[327] ,
		_w3936_,
		_w3938_
	);
	LUT2 #(
		.INIT('h1)
	) name2937 (
		_w3937_,
		_w3938_,
		_w3939_
	);
	LUT2 #(
		.INIT('h8)
	) name2938 (
		\A[328] ,
		\A[329] ,
		_w3940_
	);
	LUT2 #(
		.INIT('h1)
	) name2939 (
		\A[328] ,
		\A[329] ,
		_w3941_
	);
	LUT2 #(
		.INIT('h1)
	) name2940 (
		_w3940_,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h8)
	) name2941 (
		\A[330] ,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('h1)
	) name2942 (
		\A[330] ,
		_w3942_,
		_w3944_
	);
	LUT2 #(
		.INIT('h1)
	) name2943 (
		_w3943_,
		_w3944_,
		_w3945_
	);
	LUT2 #(
		.INIT('h8)
	) name2944 (
		_w3939_,
		_w3945_,
		_w3946_
	);
	LUT2 #(
		.INIT('h1)
	) name2945 (
		_w3939_,
		_w3945_,
		_w3947_
	);
	LUT2 #(
		.INIT('h1)
	) name2946 (
		_w3946_,
		_w3947_,
		_w3948_
	);
	LUT2 #(
		.INIT('h8)
	) name2947 (
		\A[319] ,
		\A[320] ,
		_w3949_
	);
	LUT2 #(
		.INIT('h1)
	) name2948 (
		\A[319] ,
		\A[320] ,
		_w3950_
	);
	LUT2 #(
		.INIT('h1)
	) name2949 (
		_w3949_,
		_w3950_,
		_w3951_
	);
	LUT2 #(
		.INIT('h8)
	) name2950 (
		\A[321] ,
		_w3951_,
		_w3952_
	);
	LUT2 #(
		.INIT('h1)
	) name2951 (
		\A[321] ,
		_w3951_,
		_w3953_
	);
	LUT2 #(
		.INIT('h1)
	) name2952 (
		_w3952_,
		_w3953_,
		_w3954_
	);
	LUT2 #(
		.INIT('h8)
	) name2953 (
		\A[322] ,
		\A[323] ,
		_w3955_
	);
	LUT2 #(
		.INIT('h1)
	) name2954 (
		\A[322] ,
		\A[323] ,
		_w3956_
	);
	LUT2 #(
		.INIT('h1)
	) name2955 (
		_w3955_,
		_w3956_,
		_w3957_
	);
	LUT2 #(
		.INIT('h8)
	) name2956 (
		\A[324] ,
		_w3957_,
		_w3958_
	);
	LUT2 #(
		.INIT('h1)
	) name2957 (
		\A[324] ,
		_w3957_,
		_w3959_
	);
	LUT2 #(
		.INIT('h1)
	) name2958 (
		_w3958_,
		_w3959_,
		_w3960_
	);
	LUT2 #(
		.INIT('h8)
	) name2959 (
		_w3954_,
		_w3960_,
		_w3961_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w3954_,
		_w3960_,
		_w3962_
	);
	LUT2 #(
		.INIT('h1)
	) name2961 (
		_w3961_,
		_w3962_,
		_w3963_
	);
	LUT2 #(
		.INIT('h8)
	) name2962 (
		_w3948_,
		_w3963_,
		_w3964_
	);
	LUT2 #(
		.INIT('h1)
	) name2963 (
		_w3940_,
		_w3943_,
		_w3965_
	);
	LUT2 #(
		.INIT('h1)
	) name2964 (
		_w3934_,
		_w3937_,
		_w3966_
	);
	LUT2 #(
		.INIT('h1)
	) name2965 (
		_w3965_,
		_w3966_,
		_w3967_
	);
	LUT2 #(
		.INIT('h8)
	) name2966 (
		_w3965_,
		_w3966_,
		_w3968_
	);
	LUT2 #(
		.INIT('h1)
	) name2967 (
		_w3967_,
		_w3968_,
		_w3969_
	);
	LUT2 #(
		.INIT('h8)
	) name2968 (
		_w3964_,
		_w3969_,
		_w3970_
	);
	LUT2 #(
		.INIT('h1)
	) name2969 (
		_w3955_,
		_w3958_,
		_w3971_
	);
	LUT2 #(
		.INIT('h1)
	) name2970 (
		_w3949_,
		_w3952_,
		_w3972_
	);
	LUT2 #(
		.INIT('h8)
	) name2971 (
		_w3971_,
		_w3972_,
		_w3973_
	);
	LUT2 #(
		.INIT('h1)
	) name2972 (
		_w3971_,
		_w3972_,
		_w3974_
	);
	LUT2 #(
		.INIT('h1)
	) name2973 (
		_w3973_,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('h2)
	) name2974 (
		_w3961_,
		_w3975_,
		_w3976_
	);
	LUT2 #(
		.INIT('h4)
	) name2975 (
		_w3961_,
		_w3975_,
		_w3977_
	);
	LUT2 #(
		.INIT('h1)
	) name2976 (
		_w3976_,
		_w3977_,
		_w3978_
	);
	LUT2 #(
		.INIT('h4)
	) name2977 (
		_w3970_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('h4)
	) name2978 (
		_w3946_,
		_w3969_,
		_w3980_
	);
	LUT2 #(
		.INIT('h2)
	) name2979 (
		_w3946_,
		_w3969_,
		_w3981_
	);
	LUT2 #(
		.INIT('h1)
	) name2980 (
		_w3964_,
		_w3980_,
		_w3982_
	);
	LUT2 #(
		.INIT('h4)
	) name2981 (
		_w3981_,
		_w3982_,
		_w3983_
	);
	LUT2 #(
		.INIT('h1)
	) name2982 (
		_w3979_,
		_w3983_,
		_w3984_
	);
	LUT2 #(
		.INIT('h1)
	) name2983 (
		_w3946_,
		_w3967_,
		_w3985_
	);
	LUT2 #(
		.INIT('h1)
	) name2984 (
		_w3968_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h1)
	) name2985 (
		_w3984_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h8)
	) name2986 (
		_w3984_,
		_w3986_,
		_w3988_
	);
	LUT2 #(
		.INIT('h1)
	) name2987 (
		_w3961_,
		_w3974_,
		_w3989_
	);
	LUT2 #(
		.INIT('h1)
	) name2988 (
		_w3973_,
		_w3989_,
		_w3990_
	);
	LUT2 #(
		.INIT('h1)
	) name2989 (
		_w3988_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('h1)
	) name2990 (
		_w3987_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h4)
	) name2991 (
		_w3933_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h2)
	) name2992 (
		_w3933_,
		_w3992_,
		_w3994_
	);
	LUT2 #(
		.INIT('h1)
	) name2993 (
		_w3928_,
		_w3931_,
		_w3995_
	);
	LUT2 #(
		.INIT('h2)
	) name2994 (
		_w3930_,
		_w3995_,
		_w3996_
	);
	LUT2 #(
		.INIT('h4)
	) name2995 (
		_w3930_,
		_w3995_,
		_w3997_
	);
	LUT2 #(
		.INIT('h1)
	) name2996 (
		_w3996_,
		_w3997_,
		_w3998_
	);
	LUT2 #(
		.INIT('h1)
	) name2997 (
		_w3987_,
		_w3988_,
		_w3999_
	);
	LUT2 #(
		.INIT('h4)
	) name2998 (
		_w3990_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h2)
	) name2999 (
		_w3990_,
		_w3999_,
		_w4001_
	);
	LUT2 #(
		.INIT('h1)
	) name3000 (
		_w4000_,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h2)
	) name3001 (
		_w3998_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h4)
	) name3002 (
		_w3998_,
		_w4002_,
		_w4004_
	);
	LUT2 #(
		.INIT('h1)
	) name3003 (
		_w3913_,
		_w3915_,
		_w4005_
	);
	LUT2 #(
		.INIT('h1)
	) name3004 (
		_w3916_,
		_w4005_,
		_w4006_
	);
	LUT2 #(
		.INIT('h1)
	) name3005 (
		_w3948_,
		_w3963_,
		_w4007_
	);
	LUT2 #(
		.INIT('h1)
	) name3006 (
		_w3964_,
		_w4007_,
		_w4008_
	);
	LUT2 #(
		.INIT('h8)
	) name3007 (
		_w4006_,
		_w4008_,
		_w4009_
	);
	LUT2 #(
		.INIT('h2)
	) name3008 (
		_w3920_,
		_w3923_,
		_w4010_
	);
	LUT2 #(
		.INIT('h1)
	) name3009 (
		_w3919_,
		_w3921_,
		_w4011_
	);
	LUT2 #(
		.INIT('h1)
	) name3010 (
		_w3892_,
		_w4011_,
		_w4012_
	);
	LUT2 #(
		.INIT('h1)
	) name3011 (
		_w4010_,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h8)
	) name3012 (
		_w4009_,
		_w4013_,
		_w4014_
	);
	LUT2 #(
		.INIT('h1)
	) name3013 (
		_w4009_,
		_w4013_,
		_w4015_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		_w3970_,
		_w3983_,
		_w4016_
	);
	LUT2 #(
		.INIT('h8)
	) name3015 (
		_w3978_,
		_w4016_,
		_w4017_
	);
	LUT2 #(
		.INIT('h1)
	) name3016 (
		_w3978_,
		_w4016_,
		_w4018_
	);
	LUT2 #(
		.INIT('h1)
	) name3017 (
		_w4017_,
		_w4018_,
		_w4019_
	);
	LUT2 #(
		.INIT('h1)
	) name3018 (
		_w4015_,
		_w4019_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name3019 (
		_w4014_,
		_w4020_,
		_w4021_
	);
	LUT2 #(
		.INIT('h1)
	) name3020 (
		_w4004_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h1)
	) name3021 (
		_w4003_,
		_w4022_,
		_w4023_
	);
	LUT2 #(
		.INIT('h1)
	) name3022 (
		_w3994_,
		_w4023_,
		_w4024_
	);
	LUT2 #(
		.INIT('h1)
	) name3023 (
		_w3993_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h1)
	) name3024 (
		_w3871_,
		_w4025_,
		_w4026_
	);
	LUT2 #(
		.INIT('h8)
	) name3025 (
		_w3871_,
		_w4025_,
		_w4027_
	);
	LUT2 #(
		.INIT('h1)
	) name3026 (
		_w3839_,
		_w3840_,
		_w4028_
	);
	LUT2 #(
		.INIT('h2)
	) name3027 (
		_w3869_,
		_w4028_,
		_w4029_
	);
	LUT2 #(
		.INIT('h4)
	) name3028 (
		_w3869_,
		_w4028_,
		_w4030_
	);
	LUT2 #(
		.INIT('h1)
	) name3029 (
		_w4029_,
		_w4030_,
		_w4031_
	);
	LUT2 #(
		.INIT('h1)
	) name3030 (
		_w3993_,
		_w3994_,
		_w4032_
	);
	LUT2 #(
		.INIT('h4)
	) name3031 (
		_w4023_,
		_w4032_,
		_w4033_
	);
	LUT2 #(
		.INIT('h2)
	) name3032 (
		_w4023_,
		_w4032_,
		_w4034_
	);
	LUT2 #(
		.INIT('h1)
	) name3033 (
		_w4033_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h2)
	) name3034 (
		_w4031_,
		_w4035_,
		_w4036_
	);
	LUT2 #(
		.INIT('h4)
	) name3035 (
		_w4031_,
		_w4035_,
		_w4037_
	);
	LUT2 #(
		.INIT('h1)
	) name3036 (
		_w3849_,
		_w3867_,
		_w4038_
	);
	LUT2 #(
		.INIT('h8)
	) name3037 (
		_w3866_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h1)
	) name3038 (
		_w3866_,
		_w4038_,
		_w4040_
	);
	LUT2 #(
		.INIT('h1)
	) name3039 (
		_w4039_,
		_w4040_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name3040 (
		_w4003_,
		_w4004_,
		_w4042_
	);
	LUT2 #(
		.INIT('h4)
	) name3041 (
		_w4021_,
		_w4042_,
		_w4043_
	);
	LUT2 #(
		.INIT('h2)
	) name3042 (
		_w4021_,
		_w4042_,
		_w4044_
	);
	LUT2 #(
		.INIT('h1)
	) name3043 (
		_w4043_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('h8)
	) name3044 (
		_w4041_,
		_w4045_,
		_w4046_
	);
	LUT2 #(
		.INIT('h1)
	) name3045 (
		_w4041_,
		_w4045_,
		_w4047_
	);
	LUT2 #(
		.INIT('h1)
	) name3046 (
		_w3851_,
		_w3853_,
		_w4048_
	);
	LUT2 #(
		.INIT('h1)
	) name3047 (
		_w3854_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('h1)
	) name3048 (
		_w4006_,
		_w4008_,
		_w4050_
	);
	LUT2 #(
		.INIT('h1)
	) name3049 (
		_w4009_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h8)
	) name3050 (
		_w4049_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h1)
	) name3051 (
		_w3859_,
		_w3864_,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name3052 (
		_w3863_,
		_w4053_,
		_w4054_
	);
	LUT2 #(
		.INIT('h4)
	) name3053 (
		_w3863_,
		_w4053_,
		_w4055_
	);
	LUT2 #(
		.INIT('h1)
	) name3054 (
		_w4054_,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h2)
	) name3055 (
		_w4052_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h4)
	) name3056 (
		_w4052_,
		_w4056_,
		_w4058_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w4014_,
		_w4015_,
		_w4059_
	);
	LUT2 #(
		.INIT('h4)
	) name3058 (
		_w4019_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h2)
	) name3059 (
		_w4019_,
		_w4059_,
		_w4061_
	);
	LUT2 #(
		.INIT('h1)
	) name3060 (
		_w4060_,
		_w4061_,
		_w4062_
	);
	LUT2 #(
		.INIT('h4)
	) name3061 (
		_w4058_,
		_w4062_,
		_w4063_
	);
	LUT2 #(
		.INIT('h1)
	) name3062 (
		_w4057_,
		_w4063_,
		_w4064_
	);
	LUT2 #(
		.INIT('h1)
	) name3063 (
		_w4047_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h1)
	) name3064 (
		_w4046_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('h4)
	) name3065 (
		_w4037_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h1)
	) name3066 (
		_w4036_,
		_w4067_,
		_w4068_
	);
	LUT2 #(
		.INIT('h4)
	) name3067 (
		_w4027_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		_w4026_,
		_w4069_,
		_w4070_
	);
	LUT2 #(
		.INIT('h8)
	) name3069 (
		\A[301] ,
		\A[302] ,
		_w4071_
	);
	LUT2 #(
		.INIT('h1)
	) name3070 (
		\A[301] ,
		\A[302] ,
		_w4072_
	);
	LUT2 #(
		.INIT('h1)
	) name3071 (
		_w4071_,
		_w4072_,
		_w4073_
	);
	LUT2 #(
		.INIT('h8)
	) name3072 (
		\A[303] ,
		_w4073_,
		_w4074_
	);
	LUT2 #(
		.INIT('h1)
	) name3073 (
		\A[303] ,
		_w4073_,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name3074 (
		_w4074_,
		_w4075_,
		_w4076_
	);
	LUT2 #(
		.INIT('h8)
	) name3075 (
		\A[304] ,
		\A[305] ,
		_w4077_
	);
	LUT2 #(
		.INIT('h1)
	) name3076 (
		\A[304] ,
		\A[305] ,
		_w4078_
	);
	LUT2 #(
		.INIT('h1)
	) name3077 (
		_w4077_,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('h8)
	) name3078 (
		\A[306] ,
		_w4079_,
		_w4080_
	);
	LUT2 #(
		.INIT('h1)
	) name3079 (
		\A[306] ,
		_w4079_,
		_w4081_
	);
	LUT2 #(
		.INIT('h1)
	) name3080 (
		_w4080_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h8)
	) name3081 (
		_w4076_,
		_w4082_,
		_w4083_
	);
	LUT2 #(
		.INIT('h1)
	) name3082 (
		_w4076_,
		_w4082_,
		_w4084_
	);
	LUT2 #(
		.INIT('h1)
	) name3083 (
		_w4083_,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h8)
	) name3084 (
		\A[295] ,
		\A[296] ,
		_w4086_
	);
	LUT2 #(
		.INIT('h1)
	) name3085 (
		\A[295] ,
		\A[296] ,
		_w4087_
	);
	LUT2 #(
		.INIT('h1)
	) name3086 (
		_w4086_,
		_w4087_,
		_w4088_
	);
	LUT2 #(
		.INIT('h8)
	) name3087 (
		\A[297] ,
		_w4088_,
		_w4089_
	);
	LUT2 #(
		.INIT('h1)
	) name3088 (
		\A[297] ,
		_w4088_,
		_w4090_
	);
	LUT2 #(
		.INIT('h1)
	) name3089 (
		_w4089_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h8)
	) name3090 (
		\A[298] ,
		\A[299] ,
		_w4092_
	);
	LUT2 #(
		.INIT('h1)
	) name3091 (
		\A[298] ,
		\A[299] ,
		_w4093_
	);
	LUT2 #(
		.INIT('h1)
	) name3092 (
		_w4092_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h8)
	) name3093 (
		\A[300] ,
		_w4094_,
		_w4095_
	);
	LUT2 #(
		.INIT('h1)
	) name3094 (
		\A[300] ,
		_w4094_,
		_w4096_
	);
	LUT2 #(
		.INIT('h1)
	) name3095 (
		_w4095_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h8)
	) name3096 (
		_w4091_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h1)
	) name3097 (
		_w4091_,
		_w4097_,
		_w4099_
	);
	LUT2 #(
		.INIT('h1)
	) name3098 (
		_w4098_,
		_w4099_,
		_w4100_
	);
	LUT2 #(
		.INIT('h8)
	) name3099 (
		_w4085_,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h1)
	) name3100 (
		_w4077_,
		_w4080_,
		_w4102_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		_w4071_,
		_w4074_,
		_w4103_
	);
	LUT2 #(
		.INIT('h1)
	) name3102 (
		_w4102_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h8)
	) name3103 (
		_w4102_,
		_w4103_,
		_w4105_
	);
	LUT2 #(
		.INIT('h1)
	) name3104 (
		_w4104_,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h8)
	) name3105 (
		_w4101_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h1)
	) name3106 (
		_w4092_,
		_w4095_,
		_w4108_
	);
	LUT2 #(
		.INIT('h1)
	) name3107 (
		_w4086_,
		_w4089_,
		_w4109_
	);
	LUT2 #(
		.INIT('h1)
	) name3108 (
		_w4108_,
		_w4109_,
		_w4110_
	);
	LUT2 #(
		.INIT('h8)
	) name3109 (
		_w4108_,
		_w4109_,
		_w4111_
	);
	LUT2 #(
		.INIT('h1)
	) name3110 (
		_w4110_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h2)
	) name3111 (
		_w4098_,
		_w4112_,
		_w4113_
	);
	LUT2 #(
		.INIT('h4)
	) name3112 (
		_w4098_,
		_w4112_,
		_w4114_
	);
	LUT2 #(
		.INIT('h1)
	) name3113 (
		_w4113_,
		_w4114_,
		_w4115_
	);
	LUT2 #(
		.INIT('h4)
	) name3114 (
		_w4107_,
		_w4115_,
		_w4116_
	);
	LUT2 #(
		.INIT('h4)
	) name3115 (
		_w4083_,
		_w4106_,
		_w4117_
	);
	LUT2 #(
		.INIT('h2)
	) name3116 (
		_w4083_,
		_w4106_,
		_w4118_
	);
	LUT2 #(
		.INIT('h1)
	) name3117 (
		_w4101_,
		_w4117_,
		_w4119_
	);
	LUT2 #(
		.INIT('h4)
	) name3118 (
		_w4118_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h1)
	) name3119 (
		_w4116_,
		_w4120_,
		_w4121_
	);
	LUT2 #(
		.INIT('h1)
	) name3120 (
		_w4083_,
		_w4104_,
		_w4122_
	);
	LUT2 #(
		.INIT('h1)
	) name3121 (
		_w4105_,
		_w4122_,
		_w4123_
	);
	LUT2 #(
		.INIT('h1)
	) name3122 (
		_w4121_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h8)
	) name3123 (
		_w4121_,
		_w4123_,
		_w4125_
	);
	LUT2 #(
		.INIT('h1)
	) name3124 (
		_w4098_,
		_w4110_,
		_w4126_
	);
	LUT2 #(
		.INIT('h1)
	) name3125 (
		_w4111_,
		_w4126_,
		_w4127_
	);
	LUT2 #(
		.INIT('h1)
	) name3126 (
		_w4125_,
		_w4127_,
		_w4128_
	);
	LUT2 #(
		.INIT('h1)
	) name3127 (
		_w4124_,
		_w4128_,
		_w4129_
	);
	LUT2 #(
		.INIT('h1)
	) name3128 (
		_w4124_,
		_w4125_,
		_w4130_
	);
	LUT2 #(
		.INIT('h4)
	) name3129 (
		_w4127_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h2)
	) name3130 (
		_w4127_,
		_w4130_,
		_w4132_
	);
	LUT2 #(
		.INIT('h1)
	) name3131 (
		_w4131_,
		_w4132_,
		_w4133_
	);
	LUT2 #(
		.INIT('h8)
	) name3132 (
		\A[313] ,
		\A[314] ,
		_w4134_
	);
	LUT2 #(
		.INIT('h1)
	) name3133 (
		\A[313] ,
		\A[314] ,
		_w4135_
	);
	LUT2 #(
		.INIT('h1)
	) name3134 (
		_w4134_,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h8)
	) name3135 (
		\A[315] ,
		_w4136_,
		_w4137_
	);
	LUT2 #(
		.INIT('h1)
	) name3136 (
		\A[315] ,
		_w4136_,
		_w4138_
	);
	LUT2 #(
		.INIT('h1)
	) name3137 (
		_w4137_,
		_w4138_,
		_w4139_
	);
	LUT2 #(
		.INIT('h8)
	) name3138 (
		\A[316] ,
		\A[317] ,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name3139 (
		\A[316] ,
		\A[317] ,
		_w4141_
	);
	LUT2 #(
		.INIT('h1)
	) name3140 (
		_w4140_,
		_w4141_,
		_w4142_
	);
	LUT2 #(
		.INIT('h8)
	) name3141 (
		\A[318] ,
		_w4142_,
		_w4143_
	);
	LUT2 #(
		.INIT('h1)
	) name3142 (
		\A[318] ,
		_w4142_,
		_w4144_
	);
	LUT2 #(
		.INIT('h1)
	) name3143 (
		_w4143_,
		_w4144_,
		_w4145_
	);
	LUT2 #(
		.INIT('h8)
	) name3144 (
		_w4139_,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h1)
	) name3145 (
		_w4139_,
		_w4145_,
		_w4147_
	);
	LUT2 #(
		.INIT('h1)
	) name3146 (
		_w4146_,
		_w4147_,
		_w4148_
	);
	LUT2 #(
		.INIT('h8)
	) name3147 (
		\A[307] ,
		\A[308] ,
		_w4149_
	);
	LUT2 #(
		.INIT('h1)
	) name3148 (
		\A[307] ,
		\A[308] ,
		_w4150_
	);
	LUT2 #(
		.INIT('h1)
	) name3149 (
		_w4149_,
		_w4150_,
		_w4151_
	);
	LUT2 #(
		.INIT('h8)
	) name3150 (
		\A[309] ,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h1)
	) name3151 (
		\A[309] ,
		_w4151_,
		_w4153_
	);
	LUT2 #(
		.INIT('h1)
	) name3152 (
		_w4152_,
		_w4153_,
		_w4154_
	);
	LUT2 #(
		.INIT('h8)
	) name3153 (
		\A[310] ,
		\A[311] ,
		_w4155_
	);
	LUT2 #(
		.INIT('h1)
	) name3154 (
		\A[310] ,
		\A[311] ,
		_w4156_
	);
	LUT2 #(
		.INIT('h1)
	) name3155 (
		_w4155_,
		_w4156_,
		_w4157_
	);
	LUT2 #(
		.INIT('h8)
	) name3156 (
		\A[312] ,
		_w4157_,
		_w4158_
	);
	LUT2 #(
		.INIT('h1)
	) name3157 (
		\A[312] ,
		_w4157_,
		_w4159_
	);
	LUT2 #(
		.INIT('h1)
	) name3158 (
		_w4158_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h8)
	) name3159 (
		_w4154_,
		_w4160_,
		_w4161_
	);
	LUT2 #(
		.INIT('h1)
	) name3160 (
		_w4154_,
		_w4160_,
		_w4162_
	);
	LUT2 #(
		.INIT('h1)
	) name3161 (
		_w4161_,
		_w4162_,
		_w4163_
	);
	LUT2 #(
		.INIT('h8)
	) name3162 (
		_w4148_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h1)
	) name3163 (
		_w4140_,
		_w4143_,
		_w4165_
	);
	LUT2 #(
		.INIT('h1)
	) name3164 (
		_w4134_,
		_w4137_,
		_w4166_
	);
	LUT2 #(
		.INIT('h1)
	) name3165 (
		_w4165_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name3166 (
		_w4165_,
		_w4166_,
		_w4168_
	);
	LUT2 #(
		.INIT('h1)
	) name3167 (
		_w4167_,
		_w4168_,
		_w4169_
	);
	LUT2 #(
		.INIT('h8)
	) name3168 (
		_w4164_,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h1)
	) name3169 (
		_w4155_,
		_w4158_,
		_w4171_
	);
	LUT2 #(
		.INIT('h1)
	) name3170 (
		_w4149_,
		_w4152_,
		_w4172_
	);
	LUT2 #(
		.INIT('h1)
	) name3171 (
		_w4171_,
		_w4172_,
		_w4173_
	);
	LUT2 #(
		.INIT('h8)
	) name3172 (
		_w4171_,
		_w4172_,
		_w4174_
	);
	LUT2 #(
		.INIT('h1)
	) name3173 (
		_w4173_,
		_w4174_,
		_w4175_
	);
	LUT2 #(
		.INIT('h2)
	) name3174 (
		_w4161_,
		_w4175_,
		_w4176_
	);
	LUT2 #(
		.INIT('h4)
	) name3175 (
		_w4161_,
		_w4175_,
		_w4177_
	);
	LUT2 #(
		.INIT('h1)
	) name3176 (
		_w4176_,
		_w4177_,
		_w4178_
	);
	LUT2 #(
		.INIT('h4)
	) name3177 (
		_w4170_,
		_w4178_,
		_w4179_
	);
	LUT2 #(
		.INIT('h4)
	) name3178 (
		_w4146_,
		_w4169_,
		_w4180_
	);
	LUT2 #(
		.INIT('h2)
	) name3179 (
		_w4146_,
		_w4169_,
		_w4181_
	);
	LUT2 #(
		.INIT('h1)
	) name3180 (
		_w4164_,
		_w4180_,
		_w4182_
	);
	LUT2 #(
		.INIT('h4)
	) name3181 (
		_w4181_,
		_w4182_,
		_w4183_
	);
	LUT2 #(
		.INIT('h1)
	) name3182 (
		_w4179_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h1)
	) name3183 (
		_w4146_,
		_w4167_,
		_w4185_
	);
	LUT2 #(
		.INIT('h1)
	) name3184 (
		_w4168_,
		_w4185_,
		_w4186_
	);
	LUT2 #(
		.INIT('h1)
	) name3185 (
		_w4184_,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h8)
	) name3186 (
		_w4184_,
		_w4186_,
		_w4188_
	);
	LUT2 #(
		.INIT('h1)
	) name3187 (
		_w4187_,
		_w4188_,
		_w4189_
	);
	LUT2 #(
		.INIT('h1)
	) name3188 (
		_w4161_,
		_w4173_,
		_w4190_
	);
	LUT2 #(
		.INIT('h1)
	) name3189 (
		_w4174_,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h2)
	) name3190 (
		_w4189_,
		_w4191_,
		_w4192_
	);
	LUT2 #(
		.INIT('h4)
	) name3191 (
		_w4189_,
		_w4191_,
		_w4193_
	);
	LUT2 #(
		.INIT('h1)
	) name3192 (
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h1)
	) name3193 (
		_w4133_,
		_w4194_,
		_w4195_
	);
	LUT2 #(
		.INIT('h8)
	) name3194 (
		_w4133_,
		_w4194_,
		_w4196_
	);
	LUT2 #(
		.INIT('h1)
	) name3195 (
		_w4148_,
		_w4163_,
		_w4197_
	);
	LUT2 #(
		.INIT('h1)
	) name3196 (
		_w4164_,
		_w4197_,
		_w4198_
	);
	LUT2 #(
		.INIT('h1)
	) name3197 (
		_w4085_,
		_w4100_,
		_w4199_
	);
	LUT2 #(
		.INIT('h1)
	) name3198 (
		_w4101_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h8)
	) name3199 (
		_w4198_,
		_w4200_,
		_w4201_
	);
	LUT2 #(
		.INIT('h1)
	) name3200 (
		_w4170_,
		_w4183_,
		_w4202_
	);
	LUT2 #(
		.INIT('h8)
	) name3201 (
		_w4178_,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h1)
	) name3202 (
		_w4178_,
		_w4202_,
		_w4204_
	);
	LUT2 #(
		.INIT('h1)
	) name3203 (
		_w4203_,
		_w4204_,
		_w4205_
	);
	LUT2 #(
		.INIT('h2)
	) name3204 (
		_w4201_,
		_w4205_,
		_w4206_
	);
	LUT2 #(
		.INIT('h4)
	) name3205 (
		_w4201_,
		_w4205_,
		_w4207_
	);
	LUT2 #(
		.INIT('h1)
	) name3206 (
		_w4107_,
		_w4120_,
		_w4208_
	);
	LUT2 #(
		.INIT('h8)
	) name3207 (
		_w4115_,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name3208 (
		_w4115_,
		_w4208_,
		_w4210_
	);
	LUT2 #(
		.INIT('h1)
	) name3209 (
		_w4209_,
		_w4210_,
		_w4211_
	);
	LUT2 #(
		.INIT('h1)
	) name3210 (
		_w4207_,
		_w4211_,
		_w4212_
	);
	LUT2 #(
		.INIT('h1)
	) name3211 (
		_w4206_,
		_w4212_,
		_w4213_
	);
	LUT2 #(
		.INIT('h1)
	) name3212 (
		_w4196_,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h1)
	) name3213 (
		_w4195_,
		_w4214_,
		_w4215_
	);
	LUT2 #(
		.INIT('h2)
	) name3214 (
		_w4129_,
		_w4215_,
		_w4216_
	);
	LUT2 #(
		.INIT('h4)
	) name3215 (
		_w4129_,
		_w4215_,
		_w4217_
	);
	LUT2 #(
		.INIT('h1)
	) name3216 (
		_w4188_,
		_w4191_,
		_w4218_
	);
	LUT2 #(
		.INIT('h1)
	) name3217 (
		_w4187_,
		_w4218_,
		_w4219_
	);
	LUT2 #(
		.INIT('h4)
	) name3218 (
		_w4217_,
		_w4219_,
		_w4220_
	);
	LUT2 #(
		.INIT('h1)
	) name3219 (
		_w4216_,
		_w4220_,
		_w4221_
	);
	LUT2 #(
		.INIT('h8)
	) name3220 (
		\A[277] ,
		\A[278] ,
		_w4222_
	);
	LUT2 #(
		.INIT('h1)
	) name3221 (
		\A[277] ,
		\A[278] ,
		_w4223_
	);
	LUT2 #(
		.INIT('h1)
	) name3222 (
		_w4222_,
		_w4223_,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name3223 (
		\A[279] ,
		_w4224_,
		_w4225_
	);
	LUT2 #(
		.INIT('h1)
	) name3224 (
		\A[279] ,
		_w4224_,
		_w4226_
	);
	LUT2 #(
		.INIT('h1)
	) name3225 (
		_w4225_,
		_w4226_,
		_w4227_
	);
	LUT2 #(
		.INIT('h8)
	) name3226 (
		\A[280] ,
		\A[281] ,
		_w4228_
	);
	LUT2 #(
		.INIT('h1)
	) name3227 (
		\A[280] ,
		\A[281] ,
		_w4229_
	);
	LUT2 #(
		.INIT('h1)
	) name3228 (
		_w4228_,
		_w4229_,
		_w4230_
	);
	LUT2 #(
		.INIT('h8)
	) name3229 (
		\A[282] ,
		_w4230_,
		_w4231_
	);
	LUT2 #(
		.INIT('h1)
	) name3230 (
		\A[282] ,
		_w4230_,
		_w4232_
	);
	LUT2 #(
		.INIT('h1)
	) name3231 (
		_w4231_,
		_w4232_,
		_w4233_
	);
	LUT2 #(
		.INIT('h8)
	) name3232 (
		_w4227_,
		_w4233_,
		_w4234_
	);
	LUT2 #(
		.INIT('h1)
	) name3233 (
		_w4227_,
		_w4233_,
		_w4235_
	);
	LUT2 #(
		.INIT('h1)
	) name3234 (
		_w4234_,
		_w4235_,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name3235 (
		\A[271] ,
		\A[272] ,
		_w4237_
	);
	LUT2 #(
		.INIT('h1)
	) name3236 (
		\A[271] ,
		\A[272] ,
		_w4238_
	);
	LUT2 #(
		.INIT('h1)
	) name3237 (
		_w4237_,
		_w4238_,
		_w4239_
	);
	LUT2 #(
		.INIT('h8)
	) name3238 (
		\A[273] ,
		_w4239_,
		_w4240_
	);
	LUT2 #(
		.INIT('h1)
	) name3239 (
		\A[273] ,
		_w4239_,
		_w4241_
	);
	LUT2 #(
		.INIT('h1)
	) name3240 (
		_w4240_,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h8)
	) name3241 (
		\A[274] ,
		\A[275] ,
		_w4243_
	);
	LUT2 #(
		.INIT('h1)
	) name3242 (
		\A[274] ,
		\A[275] ,
		_w4244_
	);
	LUT2 #(
		.INIT('h1)
	) name3243 (
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT2 #(
		.INIT('h8)
	) name3244 (
		\A[276] ,
		_w4245_,
		_w4246_
	);
	LUT2 #(
		.INIT('h1)
	) name3245 (
		\A[276] ,
		_w4245_,
		_w4247_
	);
	LUT2 #(
		.INIT('h1)
	) name3246 (
		_w4246_,
		_w4247_,
		_w4248_
	);
	LUT2 #(
		.INIT('h8)
	) name3247 (
		_w4242_,
		_w4248_,
		_w4249_
	);
	LUT2 #(
		.INIT('h1)
	) name3248 (
		_w4242_,
		_w4248_,
		_w4250_
	);
	LUT2 #(
		.INIT('h1)
	) name3249 (
		_w4249_,
		_w4250_,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name3250 (
		_w4236_,
		_w4251_,
		_w4252_
	);
	LUT2 #(
		.INIT('h1)
	) name3251 (
		_w4228_,
		_w4231_,
		_w4253_
	);
	LUT2 #(
		.INIT('h1)
	) name3252 (
		_w4222_,
		_w4225_,
		_w4254_
	);
	LUT2 #(
		.INIT('h1)
	) name3253 (
		_w4253_,
		_w4254_,
		_w4255_
	);
	LUT2 #(
		.INIT('h8)
	) name3254 (
		_w4253_,
		_w4254_,
		_w4256_
	);
	LUT2 #(
		.INIT('h1)
	) name3255 (
		_w4255_,
		_w4256_,
		_w4257_
	);
	LUT2 #(
		.INIT('h8)
	) name3256 (
		_w4252_,
		_w4257_,
		_w4258_
	);
	LUT2 #(
		.INIT('h1)
	) name3257 (
		_w4243_,
		_w4246_,
		_w4259_
	);
	LUT2 #(
		.INIT('h1)
	) name3258 (
		_w4237_,
		_w4240_,
		_w4260_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w4259_,
		_w4260_,
		_w4261_
	);
	LUT2 #(
		.INIT('h8)
	) name3260 (
		_w4259_,
		_w4260_,
		_w4262_
	);
	LUT2 #(
		.INIT('h1)
	) name3261 (
		_w4261_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('h2)
	) name3262 (
		_w4249_,
		_w4263_,
		_w4264_
	);
	LUT2 #(
		.INIT('h4)
	) name3263 (
		_w4249_,
		_w4263_,
		_w4265_
	);
	LUT2 #(
		.INIT('h1)
	) name3264 (
		_w4264_,
		_w4265_,
		_w4266_
	);
	LUT2 #(
		.INIT('h4)
	) name3265 (
		_w4258_,
		_w4266_,
		_w4267_
	);
	LUT2 #(
		.INIT('h4)
	) name3266 (
		_w4234_,
		_w4257_,
		_w4268_
	);
	LUT2 #(
		.INIT('h2)
	) name3267 (
		_w4234_,
		_w4257_,
		_w4269_
	);
	LUT2 #(
		.INIT('h1)
	) name3268 (
		_w4252_,
		_w4268_,
		_w4270_
	);
	LUT2 #(
		.INIT('h4)
	) name3269 (
		_w4269_,
		_w4270_,
		_w4271_
	);
	LUT2 #(
		.INIT('h1)
	) name3270 (
		_w4267_,
		_w4271_,
		_w4272_
	);
	LUT2 #(
		.INIT('h1)
	) name3271 (
		_w4234_,
		_w4255_,
		_w4273_
	);
	LUT2 #(
		.INIT('h1)
	) name3272 (
		_w4256_,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('h1)
	) name3273 (
		_w4272_,
		_w4274_,
		_w4275_
	);
	LUT2 #(
		.INIT('h8)
	) name3274 (
		_w4272_,
		_w4274_,
		_w4276_
	);
	LUT2 #(
		.INIT('h1)
	) name3275 (
		_w4249_,
		_w4261_,
		_w4277_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		_w4262_,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h1)
	) name3277 (
		_w4276_,
		_w4278_,
		_w4279_
	);
	LUT2 #(
		.INIT('h1)
	) name3278 (
		_w4275_,
		_w4279_,
		_w4280_
	);
	LUT2 #(
		.INIT('h1)
	) name3279 (
		_w4275_,
		_w4276_,
		_w4281_
	);
	LUT2 #(
		.INIT('h4)
	) name3280 (
		_w4278_,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h2)
	) name3281 (
		_w4278_,
		_w4281_,
		_w4283_
	);
	LUT2 #(
		.INIT('h1)
	) name3282 (
		_w4282_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('h8)
	) name3283 (
		\A[289] ,
		\A[290] ,
		_w4285_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		\A[289] ,
		\A[290] ,
		_w4286_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		_w4285_,
		_w4286_,
		_w4287_
	);
	LUT2 #(
		.INIT('h8)
	) name3286 (
		\A[291] ,
		_w4287_,
		_w4288_
	);
	LUT2 #(
		.INIT('h1)
	) name3287 (
		\A[291] ,
		_w4287_,
		_w4289_
	);
	LUT2 #(
		.INIT('h1)
	) name3288 (
		_w4288_,
		_w4289_,
		_w4290_
	);
	LUT2 #(
		.INIT('h8)
	) name3289 (
		\A[292] ,
		\A[293] ,
		_w4291_
	);
	LUT2 #(
		.INIT('h1)
	) name3290 (
		\A[292] ,
		\A[293] ,
		_w4292_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		_w4291_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h8)
	) name3292 (
		\A[294] ,
		_w4293_,
		_w4294_
	);
	LUT2 #(
		.INIT('h1)
	) name3293 (
		\A[294] ,
		_w4293_,
		_w4295_
	);
	LUT2 #(
		.INIT('h1)
	) name3294 (
		_w4294_,
		_w4295_,
		_w4296_
	);
	LUT2 #(
		.INIT('h8)
	) name3295 (
		_w4290_,
		_w4296_,
		_w4297_
	);
	LUT2 #(
		.INIT('h1)
	) name3296 (
		_w4290_,
		_w4296_,
		_w4298_
	);
	LUT2 #(
		.INIT('h1)
	) name3297 (
		_w4297_,
		_w4298_,
		_w4299_
	);
	LUT2 #(
		.INIT('h8)
	) name3298 (
		\A[283] ,
		\A[284] ,
		_w4300_
	);
	LUT2 #(
		.INIT('h1)
	) name3299 (
		\A[283] ,
		\A[284] ,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name3300 (
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('h8)
	) name3301 (
		\A[285] ,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h1)
	) name3302 (
		\A[285] ,
		_w4302_,
		_w4304_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		_w4303_,
		_w4304_,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name3304 (
		\A[286] ,
		\A[287] ,
		_w4306_
	);
	LUT2 #(
		.INIT('h1)
	) name3305 (
		\A[286] ,
		\A[287] ,
		_w4307_
	);
	LUT2 #(
		.INIT('h1)
	) name3306 (
		_w4306_,
		_w4307_,
		_w4308_
	);
	LUT2 #(
		.INIT('h8)
	) name3307 (
		\A[288] ,
		_w4308_,
		_w4309_
	);
	LUT2 #(
		.INIT('h1)
	) name3308 (
		\A[288] ,
		_w4308_,
		_w4310_
	);
	LUT2 #(
		.INIT('h1)
	) name3309 (
		_w4309_,
		_w4310_,
		_w4311_
	);
	LUT2 #(
		.INIT('h8)
	) name3310 (
		_w4305_,
		_w4311_,
		_w4312_
	);
	LUT2 #(
		.INIT('h1)
	) name3311 (
		_w4305_,
		_w4311_,
		_w4313_
	);
	LUT2 #(
		.INIT('h1)
	) name3312 (
		_w4312_,
		_w4313_,
		_w4314_
	);
	LUT2 #(
		.INIT('h8)
	) name3313 (
		_w4299_,
		_w4314_,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name3314 (
		_w4291_,
		_w4294_,
		_w4316_
	);
	LUT2 #(
		.INIT('h1)
	) name3315 (
		_w4285_,
		_w4288_,
		_w4317_
	);
	LUT2 #(
		.INIT('h1)
	) name3316 (
		_w4316_,
		_w4317_,
		_w4318_
	);
	LUT2 #(
		.INIT('h8)
	) name3317 (
		_w4316_,
		_w4317_,
		_w4319_
	);
	LUT2 #(
		.INIT('h1)
	) name3318 (
		_w4318_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name3319 (
		_w4315_,
		_w4320_,
		_w4321_
	);
	LUT2 #(
		.INIT('h1)
	) name3320 (
		_w4306_,
		_w4309_,
		_w4322_
	);
	LUT2 #(
		.INIT('h1)
	) name3321 (
		_w4300_,
		_w4303_,
		_w4323_
	);
	LUT2 #(
		.INIT('h1)
	) name3322 (
		_w4322_,
		_w4323_,
		_w4324_
	);
	LUT2 #(
		.INIT('h8)
	) name3323 (
		_w4322_,
		_w4323_,
		_w4325_
	);
	LUT2 #(
		.INIT('h1)
	) name3324 (
		_w4324_,
		_w4325_,
		_w4326_
	);
	LUT2 #(
		.INIT('h2)
	) name3325 (
		_w4312_,
		_w4326_,
		_w4327_
	);
	LUT2 #(
		.INIT('h4)
	) name3326 (
		_w4312_,
		_w4326_,
		_w4328_
	);
	LUT2 #(
		.INIT('h1)
	) name3327 (
		_w4327_,
		_w4328_,
		_w4329_
	);
	LUT2 #(
		.INIT('h4)
	) name3328 (
		_w4321_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('h4)
	) name3329 (
		_w4297_,
		_w4320_,
		_w4331_
	);
	LUT2 #(
		.INIT('h2)
	) name3330 (
		_w4297_,
		_w4320_,
		_w4332_
	);
	LUT2 #(
		.INIT('h1)
	) name3331 (
		_w4315_,
		_w4331_,
		_w4333_
	);
	LUT2 #(
		.INIT('h4)
	) name3332 (
		_w4332_,
		_w4333_,
		_w4334_
	);
	LUT2 #(
		.INIT('h1)
	) name3333 (
		_w4330_,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h1)
	) name3334 (
		_w4297_,
		_w4318_,
		_w4336_
	);
	LUT2 #(
		.INIT('h1)
	) name3335 (
		_w4319_,
		_w4336_,
		_w4337_
	);
	LUT2 #(
		.INIT('h1)
	) name3336 (
		_w4335_,
		_w4337_,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name3337 (
		_w4335_,
		_w4337_,
		_w4339_
	);
	LUT2 #(
		.INIT('h1)
	) name3338 (
		_w4338_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h1)
	) name3339 (
		_w4312_,
		_w4324_,
		_w4341_
	);
	LUT2 #(
		.INIT('h1)
	) name3340 (
		_w4325_,
		_w4341_,
		_w4342_
	);
	LUT2 #(
		.INIT('h2)
	) name3341 (
		_w4340_,
		_w4342_,
		_w4343_
	);
	LUT2 #(
		.INIT('h4)
	) name3342 (
		_w4340_,
		_w4342_,
		_w4344_
	);
	LUT2 #(
		.INIT('h1)
	) name3343 (
		_w4343_,
		_w4344_,
		_w4345_
	);
	LUT2 #(
		.INIT('h1)
	) name3344 (
		_w4284_,
		_w4345_,
		_w4346_
	);
	LUT2 #(
		.INIT('h8)
	) name3345 (
		_w4284_,
		_w4345_,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name3346 (
		_w4299_,
		_w4314_,
		_w4348_
	);
	LUT2 #(
		.INIT('h1)
	) name3347 (
		_w4315_,
		_w4348_,
		_w4349_
	);
	LUT2 #(
		.INIT('h1)
	) name3348 (
		_w4236_,
		_w4251_,
		_w4350_
	);
	LUT2 #(
		.INIT('h1)
	) name3349 (
		_w4252_,
		_w4350_,
		_w4351_
	);
	LUT2 #(
		.INIT('h8)
	) name3350 (
		_w4349_,
		_w4351_,
		_w4352_
	);
	LUT2 #(
		.INIT('h1)
	) name3351 (
		_w4321_,
		_w4334_,
		_w4353_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		_w4329_,
		_w4353_,
		_w4354_
	);
	LUT2 #(
		.INIT('h1)
	) name3353 (
		_w4329_,
		_w4353_,
		_w4355_
	);
	LUT2 #(
		.INIT('h1)
	) name3354 (
		_w4354_,
		_w4355_,
		_w4356_
	);
	LUT2 #(
		.INIT('h2)
	) name3355 (
		_w4352_,
		_w4356_,
		_w4357_
	);
	LUT2 #(
		.INIT('h4)
	) name3356 (
		_w4352_,
		_w4356_,
		_w4358_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w4258_,
		_w4271_,
		_w4359_
	);
	LUT2 #(
		.INIT('h8)
	) name3358 (
		_w4266_,
		_w4359_,
		_w4360_
	);
	LUT2 #(
		.INIT('h1)
	) name3359 (
		_w4266_,
		_w4359_,
		_w4361_
	);
	LUT2 #(
		.INIT('h1)
	) name3360 (
		_w4360_,
		_w4361_,
		_w4362_
	);
	LUT2 #(
		.INIT('h1)
	) name3361 (
		_w4358_,
		_w4362_,
		_w4363_
	);
	LUT2 #(
		.INIT('h1)
	) name3362 (
		_w4357_,
		_w4363_,
		_w4364_
	);
	LUT2 #(
		.INIT('h1)
	) name3363 (
		_w4347_,
		_w4364_,
		_w4365_
	);
	LUT2 #(
		.INIT('h1)
	) name3364 (
		_w4346_,
		_w4365_,
		_w4366_
	);
	LUT2 #(
		.INIT('h2)
	) name3365 (
		_w4280_,
		_w4366_,
		_w4367_
	);
	LUT2 #(
		.INIT('h4)
	) name3366 (
		_w4280_,
		_w4366_,
		_w4368_
	);
	LUT2 #(
		.INIT('h1)
	) name3367 (
		_w4339_,
		_w4342_,
		_w4369_
	);
	LUT2 #(
		.INIT('h1)
	) name3368 (
		_w4338_,
		_w4369_,
		_w4370_
	);
	LUT2 #(
		.INIT('h4)
	) name3369 (
		_w4368_,
		_w4370_,
		_w4371_
	);
	LUT2 #(
		.INIT('h1)
	) name3370 (
		_w4367_,
		_w4371_,
		_w4372_
	);
	LUT2 #(
		.INIT('h1)
	) name3371 (
		_w4221_,
		_w4372_,
		_w4373_
	);
	LUT2 #(
		.INIT('h8)
	) name3372 (
		_w4221_,
		_w4372_,
		_w4374_
	);
	LUT2 #(
		.INIT('h1)
	) name3373 (
		_w4216_,
		_w4217_,
		_w4375_
	);
	LUT2 #(
		.INIT('h8)
	) name3374 (
		_w4219_,
		_w4375_,
		_w4376_
	);
	LUT2 #(
		.INIT('h1)
	) name3375 (
		_w4219_,
		_w4375_,
		_w4377_
	);
	LUT2 #(
		.INIT('h1)
	) name3376 (
		_w4376_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h1)
	) name3377 (
		_w4367_,
		_w4368_,
		_w4379_
	);
	LUT2 #(
		.INIT('h8)
	) name3378 (
		_w4370_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h1)
	) name3379 (
		_w4370_,
		_w4379_,
		_w4381_
	);
	LUT2 #(
		.INIT('h1)
	) name3380 (
		_w4380_,
		_w4381_,
		_w4382_
	);
	LUT2 #(
		.INIT('h1)
	) name3381 (
		_w4378_,
		_w4382_,
		_w4383_
	);
	LUT2 #(
		.INIT('h8)
	) name3382 (
		_w4378_,
		_w4382_,
		_w4384_
	);
	LUT2 #(
		.INIT('h1)
	) name3383 (
		_w4346_,
		_w4347_,
		_w4385_
	);
	LUT2 #(
		.INIT('h4)
	) name3384 (
		_w4364_,
		_w4385_,
		_w4386_
	);
	LUT2 #(
		.INIT('h2)
	) name3385 (
		_w4364_,
		_w4385_,
		_w4387_
	);
	LUT2 #(
		.INIT('h1)
	) name3386 (
		_w4386_,
		_w4387_,
		_w4388_
	);
	LUT2 #(
		.INIT('h1)
	) name3387 (
		_w4195_,
		_w4196_,
		_w4389_
	);
	LUT2 #(
		.INIT('h4)
	) name3388 (
		_w4213_,
		_w4389_,
		_w4390_
	);
	LUT2 #(
		.INIT('h2)
	) name3389 (
		_w4213_,
		_w4389_,
		_w4391_
	);
	LUT2 #(
		.INIT('h1)
	) name3390 (
		_w4390_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h1)
	) name3391 (
		_w4388_,
		_w4392_,
		_w4393_
	);
	LUT2 #(
		.INIT('h8)
	) name3392 (
		_w4388_,
		_w4392_,
		_w4394_
	);
	LUT2 #(
		.INIT('h1)
	) name3393 (
		_w4198_,
		_w4200_,
		_w4395_
	);
	LUT2 #(
		.INIT('h1)
	) name3394 (
		_w4201_,
		_w4395_,
		_w4396_
	);
	LUT2 #(
		.INIT('h1)
	) name3395 (
		_w4349_,
		_w4351_,
		_w4397_
	);
	LUT2 #(
		.INIT('h1)
	) name3396 (
		_w4352_,
		_w4397_,
		_w4398_
	);
	LUT2 #(
		.INIT('h8)
	) name3397 (
		_w4396_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h1)
	) name3398 (
		_w4206_,
		_w4207_,
		_w4400_
	);
	LUT2 #(
		.INIT('h4)
	) name3399 (
		_w4211_,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h2)
	) name3400 (
		_w4211_,
		_w4400_,
		_w4402_
	);
	LUT2 #(
		.INIT('h1)
	) name3401 (
		_w4401_,
		_w4402_,
		_w4403_
	);
	LUT2 #(
		.INIT('h8)
	) name3402 (
		_w4399_,
		_w4403_,
		_w4404_
	);
	LUT2 #(
		.INIT('h1)
	) name3403 (
		_w4399_,
		_w4403_,
		_w4405_
	);
	LUT2 #(
		.INIT('h1)
	) name3404 (
		_w4357_,
		_w4358_,
		_w4406_
	);
	LUT2 #(
		.INIT('h4)
	) name3405 (
		_w4362_,
		_w4406_,
		_w4407_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		_w4362_,
		_w4406_,
		_w4408_
	);
	LUT2 #(
		.INIT('h1)
	) name3407 (
		_w4407_,
		_w4408_,
		_w4409_
	);
	LUT2 #(
		.INIT('h4)
	) name3408 (
		_w4405_,
		_w4409_,
		_w4410_
	);
	LUT2 #(
		.INIT('h1)
	) name3409 (
		_w4404_,
		_w4410_,
		_w4411_
	);
	LUT2 #(
		.INIT('h4)
	) name3410 (
		_w4394_,
		_w4411_,
		_w4412_
	);
	LUT2 #(
		.INIT('h1)
	) name3411 (
		_w4393_,
		_w4412_,
		_w4413_
	);
	LUT2 #(
		.INIT('h1)
	) name3412 (
		_w4384_,
		_w4413_,
		_w4414_
	);
	LUT2 #(
		.INIT('h1)
	) name3413 (
		_w4383_,
		_w4414_,
		_w4415_
	);
	LUT2 #(
		.INIT('h4)
	) name3414 (
		_w4374_,
		_w4415_,
		_w4416_
	);
	LUT2 #(
		.INIT('h1)
	) name3415 (
		_w4373_,
		_w4416_,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name3416 (
		_w4070_,
		_w4417_,
		_w4418_
	);
	LUT2 #(
		.INIT('h8)
	) name3417 (
		_w4070_,
		_w4417_,
		_w4419_
	);
	LUT2 #(
		.INIT('h1)
	) name3418 (
		_w4026_,
		_w4027_,
		_w4420_
	);
	LUT2 #(
		.INIT('h4)
	) name3419 (
		_w4068_,
		_w4420_,
		_w4421_
	);
	LUT2 #(
		.INIT('h2)
	) name3420 (
		_w4068_,
		_w4420_,
		_w4422_
	);
	LUT2 #(
		.INIT('h1)
	) name3421 (
		_w4421_,
		_w4422_,
		_w4423_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		_w4373_,
		_w4374_,
		_w4424_
	);
	LUT2 #(
		.INIT('h4)
	) name3423 (
		_w4415_,
		_w4424_,
		_w4425_
	);
	LUT2 #(
		.INIT('h2)
	) name3424 (
		_w4415_,
		_w4424_,
		_w4426_
	);
	LUT2 #(
		.INIT('h1)
	) name3425 (
		_w4425_,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		_w4423_,
		_w4427_,
		_w4428_
	);
	LUT2 #(
		.INIT('h8)
	) name3427 (
		_w4423_,
		_w4427_,
		_w4429_
	);
	LUT2 #(
		.INIT('h1)
	) name3428 (
		_w4383_,
		_w4384_,
		_w4430_
	);
	LUT2 #(
		.INIT('h4)
	) name3429 (
		_w4413_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h2)
	) name3430 (
		_w4413_,
		_w4430_,
		_w4432_
	);
	LUT2 #(
		.INIT('h1)
	) name3431 (
		_w4431_,
		_w4432_,
		_w4433_
	);
	LUT2 #(
		.INIT('h1)
	) name3432 (
		_w4036_,
		_w4037_,
		_w4434_
	);
	LUT2 #(
		.INIT('h8)
	) name3433 (
		_w4066_,
		_w4434_,
		_w4435_
	);
	LUT2 #(
		.INIT('h1)
	) name3434 (
		_w4066_,
		_w4434_,
		_w4436_
	);
	LUT2 #(
		.INIT('h1)
	) name3435 (
		_w4435_,
		_w4436_,
		_w4437_
	);
	LUT2 #(
		.INIT('h1)
	) name3436 (
		_w4433_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h8)
	) name3437 (
		_w4433_,
		_w4437_,
		_w4439_
	);
	LUT2 #(
		.INIT('h1)
	) name3438 (
		_w4393_,
		_w4394_,
		_w4440_
	);
	LUT2 #(
		.INIT('h4)
	) name3439 (
		_w4411_,
		_w4440_,
		_w4441_
	);
	LUT2 #(
		.INIT('h2)
	) name3440 (
		_w4411_,
		_w4440_,
		_w4442_
	);
	LUT2 #(
		.INIT('h1)
	) name3441 (
		_w4441_,
		_w4442_,
		_w4443_
	);
	LUT2 #(
		.INIT('h1)
	) name3442 (
		_w4046_,
		_w4047_,
		_w4444_
	);
	LUT2 #(
		.INIT('h4)
	) name3443 (
		_w4064_,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h2)
	) name3444 (
		_w4064_,
		_w4444_,
		_w4446_
	);
	LUT2 #(
		.INIT('h1)
	) name3445 (
		_w4445_,
		_w4446_,
		_w4447_
	);
	LUT2 #(
		.INIT('h1)
	) name3446 (
		_w4443_,
		_w4447_,
		_w4448_
	);
	LUT2 #(
		.INIT('h8)
	) name3447 (
		_w4443_,
		_w4447_,
		_w4449_
	);
	LUT2 #(
		.INIT('h1)
	) name3448 (
		_w4049_,
		_w4051_,
		_w4450_
	);
	LUT2 #(
		.INIT('h1)
	) name3449 (
		_w4052_,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h1)
	) name3450 (
		_w4396_,
		_w4398_,
		_w4452_
	);
	LUT2 #(
		.INIT('h1)
	) name3451 (
		_w4399_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h8)
	) name3452 (
		_w4451_,
		_w4453_,
		_w4454_
	);
	LUT2 #(
		.INIT('h1)
	) name3453 (
		_w4057_,
		_w4058_,
		_w4455_
	);
	LUT2 #(
		.INIT('h4)
	) name3454 (
		_w4062_,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h2)
	) name3455 (
		_w4062_,
		_w4455_,
		_w4457_
	);
	LUT2 #(
		.INIT('h1)
	) name3456 (
		_w4456_,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h2)
	) name3457 (
		_w4454_,
		_w4458_,
		_w4459_
	);
	LUT2 #(
		.INIT('h4)
	) name3458 (
		_w4454_,
		_w4458_,
		_w4460_
	);
	LUT2 #(
		.INIT('h1)
	) name3459 (
		_w4404_,
		_w4405_,
		_w4461_
	);
	LUT2 #(
		.INIT('h4)
	) name3460 (
		_w4409_,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h2)
	) name3461 (
		_w4409_,
		_w4461_,
		_w4463_
	);
	LUT2 #(
		.INIT('h1)
	) name3462 (
		_w4462_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h1)
	) name3463 (
		_w4460_,
		_w4464_,
		_w4465_
	);
	LUT2 #(
		.INIT('h1)
	) name3464 (
		_w4459_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h4)
	) name3465 (
		_w4449_,
		_w4466_,
		_w4467_
	);
	LUT2 #(
		.INIT('h1)
	) name3466 (
		_w4448_,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h4)
	) name3467 (
		_w4439_,
		_w4468_,
		_w4469_
	);
	LUT2 #(
		.INIT('h1)
	) name3468 (
		_w4438_,
		_w4469_,
		_w4470_
	);
	LUT2 #(
		.INIT('h1)
	) name3469 (
		_w4429_,
		_w4470_,
		_w4471_
	);
	LUT2 #(
		.INIT('h1)
	) name3470 (
		_w4428_,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h1)
	) name3471 (
		_w4419_,
		_w4472_,
		_w4473_
	);
	LUT2 #(
		.INIT('h1)
	) name3472 (
		_w4418_,
		_w4473_,
		_w4474_
	);
	LUT2 #(
		.INIT('h1)
	) name3473 (
		_w3713_,
		_w4474_,
		_w4475_
	);
	LUT2 #(
		.INIT('h8)
	) name3474 (
		_w3713_,
		_w4474_,
		_w4476_
	);
	LUT2 #(
		.INIT('h1)
	) name3475 (
		_w3657_,
		_w3658_,
		_w4477_
	);
	LUT2 #(
		.INIT('h4)
	) name3476 (
		_w3711_,
		_w4477_,
		_w4478_
	);
	LUT2 #(
		.INIT('h2)
	) name3477 (
		_w3711_,
		_w4477_,
		_w4479_
	);
	LUT2 #(
		.INIT('h1)
	) name3478 (
		_w4478_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h1)
	) name3479 (
		_w4418_,
		_w4419_,
		_w4481_
	);
	LUT2 #(
		.INIT('h4)
	) name3480 (
		_w4472_,
		_w4481_,
		_w4482_
	);
	LUT2 #(
		.INIT('h2)
	) name3481 (
		_w4472_,
		_w4481_,
		_w4483_
	);
	LUT2 #(
		.INIT('h1)
	) name3482 (
		_w4482_,
		_w4483_,
		_w4484_
	);
	LUT2 #(
		.INIT('h2)
	) name3483 (
		_w4480_,
		_w4484_,
		_w4485_
	);
	LUT2 #(
		.INIT('h4)
	) name3484 (
		_w4480_,
		_w4484_,
		_w4486_
	);
	LUT2 #(
		.INIT('h1)
	) name3485 (
		_w4428_,
		_w4429_,
		_w4487_
	);
	LUT2 #(
		.INIT('h4)
	) name3486 (
		_w4470_,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h2)
	) name3487 (
		_w4470_,
		_w4487_,
		_w4489_
	);
	LUT2 #(
		.INIT('h1)
	) name3488 (
		_w4488_,
		_w4489_,
		_w4490_
	);
	LUT2 #(
		.INIT('h1)
	) name3489 (
		_w3667_,
		_w3668_,
		_w4491_
	);
	LUT2 #(
		.INIT('h4)
	) name3490 (
		_w3709_,
		_w4491_,
		_w4492_
	);
	LUT2 #(
		.INIT('h2)
	) name3491 (
		_w3709_,
		_w4491_,
		_w4493_
	);
	LUT2 #(
		.INIT('h1)
	) name3492 (
		_w4492_,
		_w4493_,
		_w4494_
	);
	LUT2 #(
		.INIT('h4)
	) name3493 (
		_w4490_,
		_w4494_,
		_w4495_
	);
	LUT2 #(
		.INIT('h2)
	) name3494 (
		_w4490_,
		_w4494_,
		_w4496_
	);
	LUT2 #(
		.INIT('h1)
	) name3495 (
		_w3677_,
		_w3678_,
		_w4497_
	);
	LUT2 #(
		.INIT('h4)
	) name3496 (
		_w3707_,
		_w4497_,
		_w4498_
	);
	LUT2 #(
		.INIT('h2)
	) name3497 (
		_w3707_,
		_w4497_,
		_w4499_
	);
	LUT2 #(
		.INIT('h1)
	) name3498 (
		_w4498_,
		_w4499_,
		_w4500_
	);
	LUT2 #(
		.INIT('h1)
	) name3499 (
		_w4438_,
		_w4439_,
		_w4501_
	);
	LUT2 #(
		.INIT('h8)
	) name3500 (
		_w4468_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h1)
	) name3501 (
		_w4468_,
		_w4501_,
		_w4503_
	);
	LUT2 #(
		.INIT('h1)
	) name3502 (
		_w4502_,
		_w4503_,
		_w4504_
	);
	LUT2 #(
		.INIT('h2)
	) name3503 (
		_w4500_,
		_w4504_,
		_w4505_
	);
	LUT2 #(
		.INIT('h4)
	) name3504 (
		_w4500_,
		_w4504_,
		_w4506_
	);
	LUT2 #(
		.INIT('h1)
	) name3505 (
		_w4448_,
		_w4449_,
		_w4507_
	);
	LUT2 #(
		.INIT('h4)
	) name3506 (
		_w4466_,
		_w4507_,
		_w4508_
	);
	LUT2 #(
		.INIT('h2)
	) name3507 (
		_w4466_,
		_w4507_,
		_w4509_
	);
	LUT2 #(
		.INIT('h1)
	) name3508 (
		_w4508_,
		_w4509_,
		_w4510_
	);
	LUT2 #(
		.INIT('h1)
	) name3509 (
		_w3687_,
		_w3688_,
		_w4511_
	);
	LUT2 #(
		.INIT('h4)
	) name3510 (
		_w3705_,
		_w4511_,
		_w4512_
	);
	LUT2 #(
		.INIT('h2)
	) name3511 (
		_w3705_,
		_w4511_,
		_w4513_
	);
	LUT2 #(
		.INIT('h1)
	) name3512 (
		_w4512_,
		_w4513_,
		_w4514_
	);
	LUT2 #(
		.INIT('h1)
	) name3513 (
		_w4510_,
		_w4514_,
		_w4515_
	);
	LUT2 #(
		.INIT('h8)
	) name3514 (
		_w4510_,
		_w4514_,
		_w4516_
	);
	LUT2 #(
		.INIT('h1)
	) name3515 (
		_w3690_,
		_w3692_,
		_w4517_
	);
	LUT2 #(
		.INIT('h1)
	) name3516 (
		_w3693_,
		_w4517_,
		_w4518_
	);
	LUT2 #(
		.INIT('h1)
	) name3517 (
		_w4451_,
		_w4453_,
		_w4519_
	);
	LUT2 #(
		.INIT('h1)
	) name3518 (
		_w4454_,
		_w4519_,
		_w4520_
	);
	LUT2 #(
		.INIT('h8)
	) name3519 (
		_w4518_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h1)
	) name3520 (
		_w3698_,
		_w3699_,
		_w4522_
	);
	LUT2 #(
		.INIT('h4)
	) name3521 (
		_w3703_,
		_w4522_,
		_w4523_
	);
	LUT2 #(
		.INIT('h2)
	) name3522 (
		_w3703_,
		_w4522_,
		_w4524_
	);
	LUT2 #(
		.INIT('h1)
	) name3523 (
		_w4523_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h8)
	) name3524 (
		_w4521_,
		_w4525_,
		_w4526_
	);
	LUT2 #(
		.INIT('h1)
	) name3525 (
		_w4521_,
		_w4525_,
		_w4527_
	);
	LUT2 #(
		.INIT('h1)
	) name3526 (
		_w4459_,
		_w4460_,
		_w4528_
	);
	LUT2 #(
		.INIT('h4)
	) name3527 (
		_w4464_,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h2)
	) name3528 (
		_w4464_,
		_w4528_,
		_w4530_
	);
	LUT2 #(
		.INIT('h1)
	) name3529 (
		_w4529_,
		_w4530_,
		_w4531_
	);
	LUT2 #(
		.INIT('h4)
	) name3530 (
		_w4527_,
		_w4531_,
		_w4532_
	);
	LUT2 #(
		.INIT('h1)
	) name3531 (
		_w4526_,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h4)
	) name3532 (
		_w4516_,
		_w4533_,
		_w4534_
	);
	LUT2 #(
		.INIT('h1)
	) name3533 (
		_w4515_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h1)
	) name3534 (
		_w4506_,
		_w4535_,
		_w4536_
	);
	LUT2 #(
		.INIT('h1)
	) name3535 (
		_w4505_,
		_w4536_,
		_w4537_
	);
	LUT2 #(
		.INIT('h1)
	) name3536 (
		_w4496_,
		_w4537_,
		_w4538_
	);
	LUT2 #(
		.INIT('h1)
	) name3537 (
		_w4495_,
		_w4538_,
		_w4539_
	);
	LUT2 #(
		.INIT('h1)
	) name3538 (
		_w4486_,
		_w4539_,
		_w4540_
	);
	LUT2 #(
		.INIT('h1)
	) name3539 (
		_w4485_,
		_w4540_,
		_w4541_
	);
	LUT2 #(
		.INIT('h4)
	) name3540 (
		_w4476_,
		_w4541_,
		_w4542_
	);
	LUT2 #(
		.INIT('h1)
	) name3541 (
		_w4475_,
		_w4542_,
		_w4543_
	);
	LUT2 #(
		.INIT('h8)
	) name3542 (
		\A[211] ,
		\A[212] ,
		_w4544_
	);
	LUT2 #(
		.INIT('h1)
	) name3543 (
		\A[211] ,
		\A[212] ,
		_w4545_
	);
	LUT2 #(
		.INIT('h1)
	) name3544 (
		_w4544_,
		_w4545_,
		_w4546_
	);
	LUT2 #(
		.INIT('h8)
	) name3545 (
		\A[213] ,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h1)
	) name3546 (
		_w4544_,
		_w4547_,
		_w4548_
	);
	LUT2 #(
		.INIT('h8)
	) name3547 (
		\A[214] ,
		\A[215] ,
		_w4549_
	);
	LUT2 #(
		.INIT('h1)
	) name3548 (
		\A[213] ,
		_w4546_,
		_w4550_
	);
	LUT2 #(
		.INIT('h1)
	) name3549 (
		_w4547_,
		_w4550_,
		_w4551_
	);
	LUT2 #(
		.INIT('h1)
	) name3550 (
		\A[214] ,
		\A[215] ,
		_w4552_
	);
	LUT2 #(
		.INIT('h1)
	) name3551 (
		_w4549_,
		_w4552_,
		_w4553_
	);
	LUT2 #(
		.INIT('h8)
	) name3552 (
		\A[216] ,
		_w4553_,
		_w4554_
	);
	LUT2 #(
		.INIT('h1)
	) name3553 (
		\A[216] ,
		_w4553_,
		_w4555_
	);
	LUT2 #(
		.INIT('h1)
	) name3554 (
		_w4554_,
		_w4555_,
		_w4556_
	);
	LUT2 #(
		.INIT('h8)
	) name3555 (
		_w4551_,
		_w4556_,
		_w4557_
	);
	LUT2 #(
		.INIT('h8)
	) name3556 (
		_w4549_,
		_w4557_,
		_w4558_
	);
	LUT2 #(
		.INIT('h1)
	) name3557 (
		_w4549_,
		_w4554_,
		_w4559_
	);
	LUT2 #(
		.INIT('h4)
	) name3558 (
		_w4557_,
		_w4559_,
		_w4560_
	);
	LUT2 #(
		.INIT('h1)
	) name3559 (
		_w4558_,
		_w4560_,
		_w4561_
	);
	LUT2 #(
		.INIT('h2)
	) name3560 (
		_w4548_,
		_w4561_,
		_w4562_
	);
	LUT2 #(
		.INIT('h4)
	) name3561 (
		_w4548_,
		_w4561_,
		_w4563_
	);
	LUT2 #(
		.INIT('h1)
	) name3562 (
		_w4562_,
		_w4563_,
		_w4564_
	);
	LUT2 #(
		.INIT('h8)
	) name3563 (
		\A[217] ,
		\A[218] ,
		_w4565_
	);
	LUT2 #(
		.INIT('h1)
	) name3564 (
		\A[217] ,
		\A[218] ,
		_w4566_
	);
	LUT2 #(
		.INIT('h1)
	) name3565 (
		_w4565_,
		_w4566_,
		_w4567_
	);
	LUT2 #(
		.INIT('h8)
	) name3566 (
		\A[219] ,
		_w4567_,
		_w4568_
	);
	LUT2 #(
		.INIT('h1)
	) name3567 (
		\A[219] ,
		_w4567_,
		_w4569_
	);
	LUT2 #(
		.INIT('h1)
	) name3568 (
		_w4568_,
		_w4569_,
		_w4570_
	);
	LUT2 #(
		.INIT('h8)
	) name3569 (
		\A[220] ,
		\A[221] ,
		_w4571_
	);
	LUT2 #(
		.INIT('h1)
	) name3570 (
		\A[220] ,
		\A[221] ,
		_w4572_
	);
	LUT2 #(
		.INIT('h1)
	) name3571 (
		_w4571_,
		_w4572_,
		_w4573_
	);
	LUT2 #(
		.INIT('h8)
	) name3572 (
		\A[222] ,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h1)
	) name3573 (
		\A[222] ,
		_w4573_,
		_w4575_
	);
	LUT2 #(
		.INIT('h1)
	) name3574 (
		_w4574_,
		_w4575_,
		_w4576_
	);
	LUT2 #(
		.INIT('h8)
	) name3575 (
		_w4570_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h1)
	) name3576 (
		_w4571_,
		_w4574_,
		_w4578_
	);
	LUT2 #(
		.INIT('h1)
	) name3577 (
		_w4565_,
		_w4568_,
		_w4579_
	);
	LUT2 #(
		.INIT('h1)
	) name3578 (
		_w4578_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h8)
	) name3579 (
		_w4578_,
		_w4579_,
		_w4581_
	);
	LUT2 #(
		.INIT('h1)
	) name3580 (
		_w4580_,
		_w4581_,
		_w4582_
	);
	LUT2 #(
		.INIT('h4)
	) name3581 (
		_w4577_,
		_w4582_,
		_w4583_
	);
	LUT2 #(
		.INIT('h1)
	) name3582 (
		_w4551_,
		_w4556_,
		_w4584_
	);
	LUT2 #(
		.INIT('h1)
	) name3583 (
		_w4557_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h1)
	) name3584 (
		_w4570_,
		_w4576_,
		_w4586_
	);
	LUT2 #(
		.INIT('h1)
	) name3585 (
		_w4577_,
		_w4586_,
		_w4587_
	);
	LUT2 #(
		.INIT('h8)
	) name3586 (
		_w4585_,
		_w4587_,
		_w4588_
	);
	LUT2 #(
		.INIT('h2)
	) name3587 (
		_w4577_,
		_w4582_,
		_w4589_
	);
	LUT2 #(
		.INIT('h1)
	) name3588 (
		_w4583_,
		_w4588_,
		_w4590_
	);
	LUT2 #(
		.INIT('h4)
	) name3589 (
		_w4589_,
		_w4590_,
		_w4591_
	);
	LUT2 #(
		.INIT('h2)
	) name3590 (
		_w4564_,
		_w4591_,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name3591 (
		_w4582_,
		_w4588_,
		_w4593_
	);
	LUT2 #(
		.INIT('h4)
	) name3592 (
		_w4548_,
		_w4558_,
		_w4594_
	);
	LUT2 #(
		.INIT('h2)
	) name3593 (
		_w4593_,
		_w4594_,
		_w4595_
	);
	LUT2 #(
		.INIT('h1)
	) name3594 (
		_w4592_,
		_w4595_,
		_w4596_
	);
	LUT2 #(
		.INIT('h4)
	) name3595 (
		_w4571_,
		_w4579_,
		_w4597_
	);
	LUT2 #(
		.INIT('h2)
	) name3596 (
		_w4577_,
		_w4597_,
		_w4598_
	);
	LUT2 #(
		.INIT('h1)
	) name3597 (
		_w4580_,
		_w4598_,
		_w4599_
	);
	LUT2 #(
		.INIT('h1)
	) name3598 (
		_w4596_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h1)
	) name3599 (
		_w4548_,
		_w4560_,
		_w4601_
	);
	LUT2 #(
		.INIT('h1)
	) name3600 (
		_w4558_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('h8)
	) name3601 (
		_w4596_,
		_w4599_,
		_w4603_
	);
	LUT2 #(
		.INIT('h1)
	) name3602 (
		_w4602_,
		_w4603_,
		_w4604_
	);
	LUT2 #(
		.INIT('h1)
	) name3603 (
		_w4600_,
		_w4604_,
		_w4605_
	);
	LUT2 #(
		.INIT('h8)
	) name3604 (
		\A[205] ,
		\A[206] ,
		_w4606_
	);
	LUT2 #(
		.INIT('h1)
	) name3605 (
		\A[205] ,
		\A[206] ,
		_w4607_
	);
	LUT2 #(
		.INIT('h1)
	) name3606 (
		_w4606_,
		_w4607_,
		_w4608_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		\A[207] ,
		_w4608_,
		_w4609_
	);
	LUT2 #(
		.INIT('h1)
	) name3608 (
		\A[207] ,
		_w4608_,
		_w4610_
	);
	LUT2 #(
		.INIT('h1)
	) name3609 (
		_w4609_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h8)
	) name3610 (
		\A[208] ,
		\A[209] ,
		_w4612_
	);
	LUT2 #(
		.INIT('h1)
	) name3611 (
		\A[208] ,
		\A[209] ,
		_w4613_
	);
	LUT2 #(
		.INIT('h1)
	) name3612 (
		_w4612_,
		_w4613_,
		_w4614_
	);
	LUT2 #(
		.INIT('h8)
	) name3613 (
		\A[210] ,
		_w4614_,
		_w4615_
	);
	LUT2 #(
		.INIT('h1)
	) name3614 (
		\A[210] ,
		_w4614_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name3615 (
		_w4615_,
		_w4616_,
		_w4617_
	);
	LUT2 #(
		.INIT('h8)
	) name3616 (
		_w4611_,
		_w4617_,
		_w4618_
	);
	LUT2 #(
		.INIT('h1)
	) name3617 (
		_w4611_,
		_w4617_,
		_w4619_
	);
	LUT2 #(
		.INIT('h1)
	) name3618 (
		_w4618_,
		_w4619_,
		_w4620_
	);
	LUT2 #(
		.INIT('h8)
	) name3619 (
		\A[199] ,
		\A[200] ,
		_w4621_
	);
	LUT2 #(
		.INIT('h1)
	) name3620 (
		\A[199] ,
		\A[200] ,
		_w4622_
	);
	LUT2 #(
		.INIT('h1)
	) name3621 (
		_w4621_,
		_w4622_,
		_w4623_
	);
	LUT2 #(
		.INIT('h8)
	) name3622 (
		\A[201] ,
		_w4623_,
		_w4624_
	);
	LUT2 #(
		.INIT('h1)
	) name3623 (
		\A[201] ,
		_w4623_,
		_w4625_
	);
	LUT2 #(
		.INIT('h1)
	) name3624 (
		_w4624_,
		_w4625_,
		_w4626_
	);
	LUT2 #(
		.INIT('h8)
	) name3625 (
		\A[202] ,
		\A[203] ,
		_w4627_
	);
	LUT2 #(
		.INIT('h1)
	) name3626 (
		\A[202] ,
		\A[203] ,
		_w4628_
	);
	LUT2 #(
		.INIT('h1)
	) name3627 (
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT2 #(
		.INIT('h8)
	) name3628 (
		\A[204] ,
		_w4629_,
		_w4630_
	);
	LUT2 #(
		.INIT('h1)
	) name3629 (
		\A[204] ,
		_w4629_,
		_w4631_
	);
	LUT2 #(
		.INIT('h1)
	) name3630 (
		_w4630_,
		_w4631_,
		_w4632_
	);
	LUT2 #(
		.INIT('h8)
	) name3631 (
		_w4626_,
		_w4632_,
		_w4633_
	);
	LUT2 #(
		.INIT('h1)
	) name3632 (
		_w4626_,
		_w4632_,
		_w4634_
	);
	LUT2 #(
		.INIT('h1)
	) name3633 (
		_w4633_,
		_w4634_,
		_w4635_
	);
	LUT2 #(
		.INIT('h8)
	) name3634 (
		_w4620_,
		_w4635_,
		_w4636_
	);
	LUT2 #(
		.INIT('h1)
	) name3635 (
		_w4606_,
		_w4609_,
		_w4637_
	);
	LUT2 #(
		.INIT('h1)
	) name3636 (
		_w4612_,
		_w4615_,
		_w4638_
	);
	LUT2 #(
		.INIT('h4)
	) name3637 (
		_w4618_,
		_w4638_,
		_w4639_
	);
	LUT2 #(
		.INIT('h8)
	) name3638 (
		_w4612_,
		_w4618_,
		_w4640_
	);
	LUT2 #(
		.INIT('h1)
	) name3639 (
		_w4639_,
		_w4640_,
		_w4641_
	);
	LUT2 #(
		.INIT('h2)
	) name3640 (
		_w4637_,
		_w4641_,
		_w4642_
	);
	LUT2 #(
		.INIT('h4)
	) name3641 (
		_w4637_,
		_w4641_,
		_w4643_
	);
	LUT2 #(
		.INIT('h1)
	) name3642 (
		_w4642_,
		_w4643_,
		_w4644_
	);
	LUT2 #(
		.INIT('h1)
	) name3643 (
		_w4636_,
		_w4644_,
		_w4645_
	);
	LUT2 #(
		.INIT('h1)
	) name3644 (
		_w4621_,
		_w4624_,
		_w4646_
	);
	LUT2 #(
		.INIT('h8)
	) name3645 (
		_w4627_,
		_w4633_,
		_w4647_
	);
	LUT2 #(
		.INIT('h1)
	) name3646 (
		_w4627_,
		_w4630_,
		_w4648_
	);
	LUT2 #(
		.INIT('h4)
	) name3647 (
		_w4633_,
		_w4648_,
		_w4649_
	);
	LUT2 #(
		.INIT('h1)
	) name3648 (
		_w4647_,
		_w4649_,
		_w4650_
	);
	LUT2 #(
		.INIT('h2)
	) name3649 (
		_w4646_,
		_w4650_,
		_w4651_
	);
	LUT2 #(
		.INIT('h4)
	) name3650 (
		_w4646_,
		_w4650_,
		_w4652_
	);
	LUT2 #(
		.INIT('h1)
	) name3651 (
		_w4651_,
		_w4652_,
		_w4653_
	);
	LUT2 #(
		.INIT('h4)
	) name3652 (
		_w4645_,
		_w4653_,
		_w4654_
	);
	LUT2 #(
		.INIT('h8)
	) name3653 (
		_w4636_,
		_w4644_,
		_w4655_
	);
	LUT2 #(
		.INIT('h1)
	) name3654 (
		_w4637_,
		_w4638_,
		_w4656_
	);
	LUT2 #(
		.INIT('h4)
	) name3655 (
		_w4646_,
		_w4647_,
		_w4657_
	);
	LUT2 #(
		.INIT('h1)
	) name3656 (
		_w4656_,
		_w4657_,
		_w4658_
	);
	LUT2 #(
		.INIT('h8)
	) name3657 (
		_w4655_,
		_w4658_,
		_w4659_
	);
	LUT2 #(
		.INIT('h1)
	) name3658 (
		_w4654_,
		_w4659_,
		_w4660_
	);
	LUT2 #(
		.INIT('h1)
	) name3659 (
		_w4637_,
		_w4639_,
		_w4661_
	);
	LUT2 #(
		.INIT('h1)
	) name3660 (
		_w4640_,
		_w4661_,
		_w4662_
	);
	LUT2 #(
		.INIT('h1)
	) name3661 (
		_w4660_,
		_w4662_,
		_w4663_
	);
	LUT2 #(
		.INIT('h1)
	) name3662 (
		_w4646_,
		_w4649_,
		_w4664_
	);
	LUT2 #(
		.INIT('h1)
	) name3663 (
		_w4647_,
		_w4664_,
		_w4665_
	);
	LUT2 #(
		.INIT('h8)
	) name3664 (
		_w4660_,
		_w4662_,
		_w4666_
	);
	LUT2 #(
		.INIT('h1)
	) name3665 (
		_w4665_,
		_w4666_,
		_w4667_
	);
	LUT2 #(
		.INIT('h1)
	) name3666 (
		_w4663_,
		_w4667_,
		_w4668_
	);
	LUT2 #(
		.INIT('h1)
	) name3667 (
		_w4605_,
		_w4668_,
		_w4669_
	);
	LUT2 #(
		.INIT('h8)
	) name3668 (
		_w4605_,
		_w4668_,
		_w4670_
	);
	LUT2 #(
		.INIT('h1)
	) name3669 (
		_w4663_,
		_w4666_,
		_w4671_
	);
	LUT2 #(
		.INIT('h2)
	) name3670 (
		_w4665_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h4)
	) name3671 (
		_w4665_,
		_w4671_,
		_w4673_
	);
	LUT2 #(
		.INIT('h1)
	) name3672 (
		_w4672_,
		_w4673_,
		_w4674_
	);
	LUT2 #(
		.INIT('h1)
	) name3673 (
		_w4600_,
		_w4603_,
		_w4675_
	);
	LUT2 #(
		.INIT('h2)
	) name3674 (
		_w4602_,
		_w4675_,
		_w4676_
	);
	LUT2 #(
		.INIT('h4)
	) name3675 (
		_w4602_,
		_w4675_,
		_w4677_
	);
	LUT2 #(
		.INIT('h1)
	) name3676 (
		_w4676_,
		_w4677_,
		_w4678_
	);
	LUT2 #(
		.INIT('h1)
	) name3677 (
		_w4674_,
		_w4678_,
		_w4679_
	);
	LUT2 #(
		.INIT('h1)
	) name3678 (
		_w4585_,
		_w4587_,
		_w4680_
	);
	LUT2 #(
		.INIT('h1)
	) name3679 (
		_w4588_,
		_w4680_,
		_w4681_
	);
	LUT2 #(
		.INIT('h1)
	) name3680 (
		_w4620_,
		_w4635_,
		_w4682_
	);
	LUT2 #(
		.INIT('h1)
	) name3681 (
		_w4636_,
		_w4682_,
		_w4683_
	);
	LUT2 #(
		.INIT('h8)
	) name3682 (
		_w4681_,
		_w4683_,
		_w4684_
	);
	LUT2 #(
		.INIT('h2)
	) name3683 (
		_w4592_,
		_w4595_,
		_w4685_
	);
	LUT2 #(
		.INIT('h1)
	) name3684 (
		_w4591_,
		_w4593_,
		_w4686_
	);
	LUT2 #(
		.INIT('h1)
	) name3685 (
		_w4564_,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('h1)
	) name3686 (
		_w4685_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h1)
	) name3687 (
		_w4684_,
		_w4688_,
		_w4689_
	);
	LUT2 #(
		.INIT('h2)
	) name3688 (
		_w4654_,
		_w4659_,
		_w4690_
	);
	LUT2 #(
		.INIT('h1)
	) name3689 (
		_w4645_,
		_w4655_,
		_w4691_
	);
	LUT2 #(
		.INIT('h1)
	) name3690 (
		_w4653_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h1)
	) name3691 (
		_w4690_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h8)
	) name3692 (
		_w4684_,
		_w4688_,
		_w4694_
	);
	LUT2 #(
		.INIT('h1)
	) name3693 (
		_w4693_,
		_w4694_,
		_w4695_
	);
	LUT2 #(
		.INIT('h1)
	) name3694 (
		_w4689_,
		_w4695_,
		_w4696_
	);
	LUT2 #(
		.INIT('h8)
	) name3695 (
		_w4674_,
		_w4678_,
		_w4697_
	);
	LUT2 #(
		.INIT('h1)
	) name3696 (
		_w4696_,
		_w4697_,
		_w4698_
	);
	LUT2 #(
		.INIT('h1)
	) name3697 (
		_w4679_,
		_w4698_,
		_w4699_
	);
	LUT2 #(
		.INIT('h4)
	) name3698 (
		_w4670_,
		_w4699_,
		_w4700_
	);
	LUT2 #(
		.INIT('h1)
	) name3699 (
		_w4669_,
		_w4700_,
		_w4701_
	);
	LUT2 #(
		.INIT('h8)
	) name3700 (
		\A[193] ,
		\A[194] ,
		_w4702_
	);
	LUT2 #(
		.INIT('h1)
	) name3701 (
		\A[193] ,
		\A[194] ,
		_w4703_
	);
	LUT2 #(
		.INIT('h1)
	) name3702 (
		_w4702_,
		_w4703_,
		_w4704_
	);
	LUT2 #(
		.INIT('h8)
	) name3703 (
		\A[195] ,
		_w4704_,
		_w4705_
	);
	LUT2 #(
		.INIT('h1)
	) name3704 (
		\A[195] ,
		_w4704_,
		_w4706_
	);
	LUT2 #(
		.INIT('h1)
	) name3705 (
		_w4705_,
		_w4706_,
		_w4707_
	);
	LUT2 #(
		.INIT('h8)
	) name3706 (
		\A[196] ,
		\A[197] ,
		_w4708_
	);
	LUT2 #(
		.INIT('h1)
	) name3707 (
		\A[196] ,
		\A[197] ,
		_w4709_
	);
	LUT2 #(
		.INIT('h1)
	) name3708 (
		_w4708_,
		_w4709_,
		_w4710_
	);
	LUT2 #(
		.INIT('h8)
	) name3709 (
		\A[198] ,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h1)
	) name3710 (
		\A[198] ,
		_w4710_,
		_w4712_
	);
	LUT2 #(
		.INIT('h1)
	) name3711 (
		_w4711_,
		_w4712_,
		_w4713_
	);
	LUT2 #(
		.INIT('h8)
	) name3712 (
		_w4707_,
		_w4713_,
		_w4714_
	);
	LUT2 #(
		.INIT('h1)
	) name3713 (
		_w4707_,
		_w4713_,
		_w4715_
	);
	LUT2 #(
		.INIT('h1)
	) name3714 (
		_w4714_,
		_w4715_,
		_w4716_
	);
	LUT2 #(
		.INIT('h8)
	) name3715 (
		\A[187] ,
		\A[188] ,
		_w4717_
	);
	LUT2 #(
		.INIT('h1)
	) name3716 (
		\A[187] ,
		\A[188] ,
		_w4718_
	);
	LUT2 #(
		.INIT('h1)
	) name3717 (
		_w4717_,
		_w4718_,
		_w4719_
	);
	LUT2 #(
		.INIT('h8)
	) name3718 (
		\A[189] ,
		_w4719_,
		_w4720_
	);
	LUT2 #(
		.INIT('h1)
	) name3719 (
		\A[189] ,
		_w4719_,
		_w4721_
	);
	LUT2 #(
		.INIT('h1)
	) name3720 (
		_w4720_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h8)
	) name3721 (
		\A[190] ,
		\A[191] ,
		_w4723_
	);
	LUT2 #(
		.INIT('h1)
	) name3722 (
		\A[190] ,
		\A[191] ,
		_w4724_
	);
	LUT2 #(
		.INIT('h1)
	) name3723 (
		_w4723_,
		_w4724_,
		_w4725_
	);
	LUT2 #(
		.INIT('h8)
	) name3724 (
		\A[192] ,
		_w4725_,
		_w4726_
	);
	LUT2 #(
		.INIT('h1)
	) name3725 (
		\A[192] ,
		_w4725_,
		_w4727_
	);
	LUT2 #(
		.INIT('h1)
	) name3726 (
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h8)
	) name3727 (
		_w4722_,
		_w4728_,
		_w4729_
	);
	LUT2 #(
		.INIT('h1)
	) name3728 (
		_w4722_,
		_w4728_,
		_w4730_
	);
	LUT2 #(
		.INIT('h1)
	) name3729 (
		_w4729_,
		_w4730_,
		_w4731_
	);
	LUT2 #(
		.INIT('h8)
	) name3730 (
		_w4716_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h1)
	) name3731 (
		_w4708_,
		_w4711_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name3732 (
		_w4702_,
		_w4705_,
		_w4734_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		_w4733_,
		_w4734_,
		_w4735_
	);
	LUT2 #(
		.INIT('h8)
	) name3734 (
		_w4733_,
		_w4734_,
		_w4736_
	);
	LUT2 #(
		.INIT('h1)
	) name3735 (
		_w4735_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h8)
	) name3736 (
		_w4732_,
		_w4737_,
		_w4738_
	);
	LUT2 #(
		.INIT('h1)
	) name3737 (
		_w4717_,
		_w4720_,
		_w4739_
	);
	LUT2 #(
		.INIT('h1)
	) name3738 (
		_w4723_,
		_w4726_,
		_w4740_
	);
	LUT2 #(
		.INIT('h4)
	) name3739 (
		_w4729_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h8)
	) name3740 (
		_w4723_,
		_w4729_,
		_w4742_
	);
	LUT2 #(
		.INIT('h1)
	) name3741 (
		_w4741_,
		_w4742_,
		_w4743_
	);
	LUT2 #(
		.INIT('h2)
	) name3742 (
		_w4739_,
		_w4743_,
		_w4744_
	);
	LUT2 #(
		.INIT('h4)
	) name3743 (
		_w4739_,
		_w4743_,
		_w4745_
	);
	LUT2 #(
		.INIT('h1)
	) name3744 (
		_w4744_,
		_w4745_,
		_w4746_
	);
	LUT2 #(
		.INIT('h1)
	) name3745 (
		_w4738_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h4)
	) name3746 (
		_w4714_,
		_w4737_,
		_w4748_
	);
	LUT2 #(
		.INIT('h2)
	) name3747 (
		_w4714_,
		_w4737_,
		_w4749_
	);
	LUT2 #(
		.INIT('h1)
	) name3748 (
		_w4732_,
		_w4748_,
		_w4750_
	);
	LUT2 #(
		.INIT('h4)
	) name3749 (
		_w4749_,
		_w4750_,
		_w4751_
	);
	LUT2 #(
		.INIT('h1)
	) name3750 (
		_w4747_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h1)
	) name3751 (
		_w4714_,
		_w4735_,
		_w4753_
	);
	LUT2 #(
		.INIT('h1)
	) name3752 (
		_w4736_,
		_w4753_,
		_w4754_
	);
	LUT2 #(
		.INIT('h1)
	) name3753 (
		_w4752_,
		_w4754_,
		_w4755_
	);
	LUT2 #(
		.INIT('h8)
	) name3754 (
		_w4752_,
		_w4754_,
		_w4756_
	);
	LUT2 #(
		.INIT('h1)
	) name3755 (
		_w4739_,
		_w4741_,
		_w4757_
	);
	LUT2 #(
		.INIT('h1)
	) name3756 (
		_w4742_,
		_w4757_,
		_w4758_
	);
	LUT2 #(
		.INIT('h4)
	) name3757 (
		_w4756_,
		_w4758_,
		_w4759_
	);
	LUT2 #(
		.INIT('h1)
	) name3758 (
		_w4755_,
		_w4759_,
		_w4760_
	);
	LUT2 #(
		.INIT('h1)
	) name3759 (
		_w4755_,
		_w4756_,
		_w4761_
	);
	LUT2 #(
		.INIT('h4)
	) name3760 (
		_w4758_,
		_w4761_,
		_w4762_
	);
	LUT2 #(
		.INIT('h2)
	) name3761 (
		_w4758_,
		_w4761_,
		_w4763_
	);
	LUT2 #(
		.INIT('h1)
	) name3762 (
		_w4762_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h8)
	) name3763 (
		\A[178] ,
		\A[179] ,
		_w4765_
	);
	LUT2 #(
		.INIT('h8)
	) name3764 (
		\A[175] ,
		\A[176] ,
		_w4766_
	);
	LUT2 #(
		.INIT('h1)
	) name3765 (
		\A[175] ,
		\A[176] ,
		_w4767_
	);
	LUT2 #(
		.INIT('h1)
	) name3766 (
		_w4766_,
		_w4767_,
		_w4768_
	);
	LUT2 #(
		.INIT('h8)
	) name3767 (
		\A[177] ,
		_w4768_,
		_w4769_
	);
	LUT2 #(
		.INIT('h1)
	) name3768 (
		\A[177] ,
		_w4768_,
		_w4770_
	);
	LUT2 #(
		.INIT('h1)
	) name3769 (
		_w4769_,
		_w4770_,
		_w4771_
	);
	LUT2 #(
		.INIT('h1)
	) name3770 (
		\A[178] ,
		\A[179] ,
		_w4772_
	);
	LUT2 #(
		.INIT('h1)
	) name3771 (
		_w4765_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h8)
	) name3772 (
		\A[180] ,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h1)
	) name3773 (
		\A[180] ,
		_w4773_,
		_w4775_
	);
	LUT2 #(
		.INIT('h1)
	) name3774 (
		_w4774_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h8)
	) name3775 (
		_w4771_,
		_w4776_,
		_w4777_
	);
	LUT2 #(
		.INIT('h8)
	) name3776 (
		_w4765_,
		_w4777_,
		_w4778_
	);
	LUT2 #(
		.INIT('h1)
	) name3777 (
		_w4766_,
		_w4769_,
		_w4779_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		_w4765_,
		_w4774_,
		_w4780_
	);
	LUT2 #(
		.INIT('h4)
	) name3779 (
		_w4777_,
		_w4780_,
		_w4781_
	);
	LUT2 #(
		.INIT('h1)
	) name3780 (
		_w4779_,
		_w4781_,
		_w4782_
	);
	LUT2 #(
		.INIT('h1)
	) name3781 (
		_w4778_,
		_w4782_,
		_w4783_
	);
	LUT2 #(
		.INIT('h8)
	) name3782 (
		\A[181] ,
		\A[182] ,
		_w4784_
	);
	LUT2 #(
		.INIT('h1)
	) name3783 (
		\A[181] ,
		\A[182] ,
		_w4785_
	);
	LUT2 #(
		.INIT('h1)
	) name3784 (
		_w4784_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h8)
	) name3785 (
		\A[183] ,
		_w4786_,
		_w4787_
	);
	LUT2 #(
		.INIT('h1)
	) name3786 (
		\A[183] ,
		_w4786_,
		_w4788_
	);
	LUT2 #(
		.INIT('h1)
	) name3787 (
		_w4787_,
		_w4788_,
		_w4789_
	);
	LUT2 #(
		.INIT('h8)
	) name3788 (
		\A[184] ,
		\A[185] ,
		_w4790_
	);
	LUT2 #(
		.INIT('h1)
	) name3789 (
		\A[184] ,
		\A[185] ,
		_w4791_
	);
	LUT2 #(
		.INIT('h1)
	) name3790 (
		_w4790_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h8)
	) name3791 (
		\A[186] ,
		_w4792_,
		_w4793_
	);
	LUT2 #(
		.INIT('h1)
	) name3792 (
		\A[186] ,
		_w4792_,
		_w4794_
	);
	LUT2 #(
		.INIT('h1)
	) name3793 (
		_w4793_,
		_w4794_,
		_w4795_
	);
	LUT2 #(
		.INIT('h8)
	) name3794 (
		_w4789_,
		_w4795_,
		_w4796_
	);
	LUT2 #(
		.INIT('h1)
	) name3795 (
		_w4789_,
		_w4795_,
		_w4797_
	);
	LUT2 #(
		.INIT('h1)
	) name3796 (
		_w4796_,
		_w4797_,
		_w4798_
	);
	LUT2 #(
		.INIT('h1)
	) name3797 (
		_w4771_,
		_w4776_,
		_w4799_
	);
	LUT2 #(
		.INIT('h1)
	) name3798 (
		_w4777_,
		_w4799_,
		_w4800_
	);
	LUT2 #(
		.INIT('h8)
	) name3799 (
		_w4798_,
		_w4800_,
		_w4801_
	);
	LUT2 #(
		.INIT('h1)
	) name3800 (
		_w4790_,
		_w4793_,
		_w4802_
	);
	LUT2 #(
		.INIT('h1)
	) name3801 (
		_w4784_,
		_w4787_,
		_w4803_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w4802_,
		_w4803_,
		_w4804_
	);
	LUT2 #(
		.INIT('h8)
	) name3803 (
		_w4802_,
		_w4803_,
		_w4805_
	);
	LUT2 #(
		.INIT('h1)
	) name3804 (
		_w4804_,
		_w4805_,
		_w4806_
	);
	LUT2 #(
		.INIT('h8)
	) name3805 (
		_w4801_,
		_w4806_,
		_w4807_
	);
	LUT2 #(
		.INIT('h1)
	) name3806 (
		_w4778_,
		_w4781_,
		_w4808_
	);
	LUT2 #(
		.INIT('h2)
	) name3807 (
		_w4779_,
		_w4808_,
		_w4809_
	);
	LUT2 #(
		.INIT('h4)
	) name3808 (
		_w4779_,
		_w4808_,
		_w4810_
	);
	LUT2 #(
		.INIT('h1)
	) name3809 (
		_w4809_,
		_w4810_,
		_w4811_
	);
	LUT2 #(
		.INIT('h1)
	) name3810 (
		_w4807_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('h4)
	) name3811 (
		_w4796_,
		_w4806_,
		_w4813_
	);
	LUT2 #(
		.INIT('h2)
	) name3812 (
		_w4796_,
		_w4806_,
		_w4814_
	);
	LUT2 #(
		.INIT('h1)
	) name3813 (
		_w4801_,
		_w4813_,
		_w4815_
	);
	LUT2 #(
		.INIT('h4)
	) name3814 (
		_w4814_,
		_w4815_,
		_w4816_
	);
	LUT2 #(
		.INIT('h1)
	) name3815 (
		_w4812_,
		_w4816_,
		_w4817_
	);
	LUT2 #(
		.INIT('h1)
	) name3816 (
		_w4796_,
		_w4804_,
		_w4818_
	);
	LUT2 #(
		.INIT('h1)
	) name3817 (
		_w4805_,
		_w4818_,
		_w4819_
	);
	LUT2 #(
		.INIT('h8)
	) name3818 (
		_w4817_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h1)
	) name3819 (
		_w4817_,
		_w4819_,
		_w4821_
	);
	LUT2 #(
		.INIT('h1)
	) name3820 (
		_w4820_,
		_w4821_,
		_w4822_
	);
	LUT2 #(
		.INIT('h2)
	) name3821 (
		_w4783_,
		_w4822_,
		_w4823_
	);
	LUT2 #(
		.INIT('h4)
	) name3822 (
		_w4783_,
		_w4822_,
		_w4824_
	);
	LUT2 #(
		.INIT('h1)
	) name3823 (
		_w4823_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h8)
	) name3824 (
		_w4764_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('h1)
	) name3825 (
		_w4764_,
		_w4825_,
		_w4827_
	);
	LUT2 #(
		.INIT('h1)
	) name3826 (
		_w4716_,
		_w4731_,
		_w4828_
	);
	LUT2 #(
		.INIT('h1)
	) name3827 (
		_w4732_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h1)
	) name3828 (
		_w4798_,
		_w4800_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		_w4801_,
		_w4830_,
		_w4831_
	);
	LUT2 #(
		.INIT('h8)
	) name3830 (
		_w4829_,
		_w4831_,
		_w4832_
	);
	LUT2 #(
		.INIT('h1)
	) name3831 (
		_w4738_,
		_w4751_,
		_w4833_
	);
	LUT2 #(
		.INIT('h4)
	) name3832 (
		_w4746_,
		_w4833_,
		_w4834_
	);
	LUT2 #(
		.INIT('h2)
	) name3833 (
		_w4746_,
		_w4833_,
		_w4835_
	);
	LUT2 #(
		.INIT('h1)
	) name3834 (
		_w4834_,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('h2)
	) name3835 (
		_w4832_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('h4)
	) name3836 (
		_w4832_,
		_w4836_,
		_w4838_
	);
	LUT2 #(
		.INIT('h1)
	) name3837 (
		_w4807_,
		_w4816_,
		_w4839_
	);
	LUT2 #(
		.INIT('h4)
	) name3838 (
		_w4811_,
		_w4839_,
		_w4840_
	);
	LUT2 #(
		.INIT('h2)
	) name3839 (
		_w4811_,
		_w4839_,
		_w4841_
	);
	LUT2 #(
		.INIT('h1)
	) name3840 (
		_w4840_,
		_w4841_,
		_w4842_
	);
	LUT2 #(
		.INIT('h1)
	) name3841 (
		_w4838_,
		_w4842_,
		_w4843_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		_w4837_,
		_w4843_,
		_w4844_
	);
	LUT2 #(
		.INIT('h1)
	) name3843 (
		_w4827_,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('h1)
	) name3844 (
		_w4826_,
		_w4845_,
		_w4846_
	);
	LUT2 #(
		.INIT('h2)
	) name3845 (
		_w4760_,
		_w4846_,
		_w4847_
	);
	LUT2 #(
		.INIT('h4)
	) name3846 (
		_w4760_,
		_w4846_,
		_w4848_
	);
	LUT2 #(
		.INIT('h2)
	) name3847 (
		_w4783_,
		_w4820_,
		_w4849_
	);
	LUT2 #(
		.INIT('h1)
	) name3848 (
		_w4821_,
		_w4849_,
		_w4850_
	);
	LUT2 #(
		.INIT('h4)
	) name3849 (
		_w4848_,
		_w4850_,
		_w4851_
	);
	LUT2 #(
		.INIT('h1)
	) name3850 (
		_w4847_,
		_w4851_,
		_w4852_
	);
	LUT2 #(
		.INIT('h1)
	) name3851 (
		_w4701_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h8)
	) name3852 (
		_w4701_,
		_w4852_,
		_w4854_
	);
	LUT2 #(
		.INIT('h1)
	) name3853 (
		_w4669_,
		_w4670_,
		_w4855_
	);
	LUT2 #(
		.INIT('h2)
	) name3854 (
		_w4699_,
		_w4855_,
		_w4856_
	);
	LUT2 #(
		.INIT('h4)
	) name3855 (
		_w4699_,
		_w4855_,
		_w4857_
	);
	LUT2 #(
		.INIT('h1)
	) name3856 (
		_w4856_,
		_w4857_,
		_w4858_
	);
	LUT2 #(
		.INIT('h1)
	) name3857 (
		_w4847_,
		_w4848_,
		_w4859_
	);
	LUT2 #(
		.INIT('h8)
	) name3858 (
		_w4850_,
		_w4859_,
		_w4860_
	);
	LUT2 #(
		.INIT('h1)
	) name3859 (
		_w4850_,
		_w4859_,
		_w4861_
	);
	LUT2 #(
		.INIT('h1)
	) name3860 (
		_w4860_,
		_w4861_,
		_w4862_
	);
	LUT2 #(
		.INIT('h4)
	) name3861 (
		_w4858_,
		_w4862_,
		_w4863_
	);
	LUT2 #(
		.INIT('h2)
	) name3862 (
		_w4858_,
		_w4862_,
		_w4864_
	);
	LUT2 #(
		.INIT('h1)
	) name3863 (
		_w4679_,
		_w4697_,
		_w4865_
	);
	LUT2 #(
		.INIT('h8)
	) name3864 (
		_w4696_,
		_w4865_,
		_w4866_
	);
	LUT2 #(
		.INIT('h1)
	) name3865 (
		_w4696_,
		_w4865_,
		_w4867_
	);
	LUT2 #(
		.INIT('h1)
	) name3866 (
		_w4866_,
		_w4867_,
		_w4868_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w4826_,
		_w4827_,
		_w4869_
	);
	LUT2 #(
		.INIT('h4)
	) name3868 (
		_w4844_,
		_w4869_,
		_w4870_
	);
	LUT2 #(
		.INIT('h2)
	) name3869 (
		_w4844_,
		_w4869_,
		_w4871_
	);
	LUT2 #(
		.INIT('h1)
	) name3870 (
		_w4870_,
		_w4871_,
		_w4872_
	);
	LUT2 #(
		.INIT('h8)
	) name3871 (
		_w4868_,
		_w4872_,
		_w4873_
	);
	LUT2 #(
		.INIT('h1)
	) name3872 (
		_w4868_,
		_w4872_,
		_w4874_
	);
	LUT2 #(
		.INIT('h1)
	) name3873 (
		_w4681_,
		_w4683_,
		_w4875_
	);
	LUT2 #(
		.INIT('h1)
	) name3874 (
		_w4684_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h1)
	) name3875 (
		_w4829_,
		_w4831_,
		_w4877_
	);
	LUT2 #(
		.INIT('h1)
	) name3876 (
		_w4832_,
		_w4877_,
		_w4878_
	);
	LUT2 #(
		.INIT('h8)
	) name3877 (
		_w4876_,
		_w4878_,
		_w4879_
	);
	LUT2 #(
		.INIT('h1)
	) name3878 (
		_w4689_,
		_w4694_,
		_w4880_
	);
	LUT2 #(
		.INIT('h2)
	) name3879 (
		_w4693_,
		_w4880_,
		_w4881_
	);
	LUT2 #(
		.INIT('h4)
	) name3880 (
		_w4693_,
		_w4880_,
		_w4882_
	);
	LUT2 #(
		.INIT('h1)
	) name3881 (
		_w4881_,
		_w4882_,
		_w4883_
	);
	LUT2 #(
		.INIT('h2)
	) name3882 (
		_w4879_,
		_w4883_,
		_w4884_
	);
	LUT2 #(
		.INIT('h4)
	) name3883 (
		_w4879_,
		_w4883_,
		_w4885_
	);
	LUT2 #(
		.INIT('h1)
	) name3884 (
		_w4837_,
		_w4838_,
		_w4886_
	);
	LUT2 #(
		.INIT('h4)
	) name3885 (
		_w4842_,
		_w4886_,
		_w4887_
	);
	LUT2 #(
		.INIT('h2)
	) name3886 (
		_w4842_,
		_w4886_,
		_w4888_
	);
	LUT2 #(
		.INIT('h1)
	) name3887 (
		_w4887_,
		_w4888_,
		_w4889_
	);
	LUT2 #(
		.INIT('h4)
	) name3888 (
		_w4885_,
		_w4889_,
		_w4890_
	);
	LUT2 #(
		.INIT('h1)
	) name3889 (
		_w4884_,
		_w4890_,
		_w4891_
	);
	LUT2 #(
		.INIT('h1)
	) name3890 (
		_w4874_,
		_w4891_,
		_w4892_
	);
	LUT2 #(
		.INIT('h1)
	) name3891 (
		_w4873_,
		_w4892_,
		_w4893_
	);
	LUT2 #(
		.INIT('h1)
	) name3892 (
		_w4864_,
		_w4893_,
		_w4894_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w4863_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h1)
	) name3894 (
		_w4854_,
		_w4895_,
		_w4896_
	);
	LUT2 #(
		.INIT('h1)
	) name3895 (
		_w4853_,
		_w4896_,
		_w4897_
	);
	LUT2 #(
		.INIT('h8)
	) name3896 (
		\A[259] ,
		\A[260] ,
		_w4898_
	);
	LUT2 #(
		.INIT('h1)
	) name3897 (
		\A[259] ,
		\A[260] ,
		_w4899_
	);
	LUT2 #(
		.INIT('h1)
	) name3898 (
		_w4898_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('h8)
	) name3899 (
		\A[261] ,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('h1)
	) name3900 (
		_w4898_,
		_w4901_,
		_w4902_
	);
	LUT2 #(
		.INIT('h8)
	) name3901 (
		\A[262] ,
		\A[263] ,
		_w4903_
	);
	LUT2 #(
		.INIT('h1)
	) name3902 (
		\A[261] ,
		_w4900_,
		_w4904_
	);
	LUT2 #(
		.INIT('h1)
	) name3903 (
		_w4901_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h1)
	) name3904 (
		\A[262] ,
		\A[263] ,
		_w4906_
	);
	LUT2 #(
		.INIT('h1)
	) name3905 (
		_w4903_,
		_w4906_,
		_w4907_
	);
	LUT2 #(
		.INIT('h8)
	) name3906 (
		\A[264] ,
		_w4907_,
		_w4908_
	);
	LUT2 #(
		.INIT('h1)
	) name3907 (
		\A[264] ,
		_w4907_,
		_w4909_
	);
	LUT2 #(
		.INIT('h1)
	) name3908 (
		_w4908_,
		_w4909_,
		_w4910_
	);
	LUT2 #(
		.INIT('h8)
	) name3909 (
		_w4905_,
		_w4910_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name3910 (
		_w4903_,
		_w4911_,
		_w4912_
	);
	LUT2 #(
		.INIT('h1)
	) name3911 (
		_w4903_,
		_w4908_,
		_w4913_
	);
	LUT2 #(
		.INIT('h4)
	) name3912 (
		_w4911_,
		_w4913_,
		_w4914_
	);
	LUT2 #(
		.INIT('h1)
	) name3913 (
		_w4912_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('h2)
	) name3914 (
		_w4902_,
		_w4915_,
		_w4916_
	);
	LUT2 #(
		.INIT('h4)
	) name3915 (
		_w4902_,
		_w4915_,
		_w4917_
	);
	LUT2 #(
		.INIT('h1)
	) name3916 (
		_w4916_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h8)
	) name3917 (
		\A[265] ,
		\A[266] ,
		_w4919_
	);
	LUT2 #(
		.INIT('h1)
	) name3918 (
		\A[265] ,
		\A[266] ,
		_w4920_
	);
	LUT2 #(
		.INIT('h1)
	) name3919 (
		_w4919_,
		_w4920_,
		_w4921_
	);
	LUT2 #(
		.INIT('h8)
	) name3920 (
		\A[267] ,
		_w4921_,
		_w4922_
	);
	LUT2 #(
		.INIT('h1)
	) name3921 (
		\A[267] ,
		_w4921_,
		_w4923_
	);
	LUT2 #(
		.INIT('h1)
	) name3922 (
		_w4922_,
		_w4923_,
		_w4924_
	);
	LUT2 #(
		.INIT('h8)
	) name3923 (
		\A[268] ,
		\A[269] ,
		_w4925_
	);
	LUT2 #(
		.INIT('h1)
	) name3924 (
		\A[268] ,
		\A[269] ,
		_w4926_
	);
	LUT2 #(
		.INIT('h1)
	) name3925 (
		_w4925_,
		_w4926_,
		_w4927_
	);
	LUT2 #(
		.INIT('h8)
	) name3926 (
		\A[270] ,
		_w4927_,
		_w4928_
	);
	LUT2 #(
		.INIT('h1)
	) name3927 (
		\A[270] ,
		_w4927_,
		_w4929_
	);
	LUT2 #(
		.INIT('h1)
	) name3928 (
		_w4928_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h8)
	) name3929 (
		_w4924_,
		_w4930_,
		_w4931_
	);
	LUT2 #(
		.INIT('h1)
	) name3930 (
		_w4925_,
		_w4928_,
		_w4932_
	);
	LUT2 #(
		.INIT('h1)
	) name3931 (
		_w4919_,
		_w4922_,
		_w4933_
	);
	LUT2 #(
		.INIT('h1)
	) name3932 (
		_w4932_,
		_w4933_,
		_w4934_
	);
	LUT2 #(
		.INIT('h8)
	) name3933 (
		_w4932_,
		_w4933_,
		_w4935_
	);
	LUT2 #(
		.INIT('h1)
	) name3934 (
		_w4934_,
		_w4935_,
		_w4936_
	);
	LUT2 #(
		.INIT('h4)
	) name3935 (
		_w4931_,
		_w4936_,
		_w4937_
	);
	LUT2 #(
		.INIT('h1)
	) name3936 (
		_w4905_,
		_w4910_,
		_w4938_
	);
	LUT2 #(
		.INIT('h1)
	) name3937 (
		_w4911_,
		_w4938_,
		_w4939_
	);
	LUT2 #(
		.INIT('h1)
	) name3938 (
		_w4924_,
		_w4930_,
		_w4940_
	);
	LUT2 #(
		.INIT('h1)
	) name3939 (
		_w4931_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h8)
	) name3940 (
		_w4939_,
		_w4941_,
		_w4942_
	);
	LUT2 #(
		.INIT('h2)
	) name3941 (
		_w4931_,
		_w4936_,
		_w4943_
	);
	LUT2 #(
		.INIT('h1)
	) name3942 (
		_w4937_,
		_w4942_,
		_w4944_
	);
	LUT2 #(
		.INIT('h4)
	) name3943 (
		_w4943_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('h2)
	) name3944 (
		_w4918_,
		_w4945_,
		_w4946_
	);
	LUT2 #(
		.INIT('h8)
	) name3945 (
		_w4936_,
		_w4942_,
		_w4947_
	);
	LUT2 #(
		.INIT('h4)
	) name3946 (
		_w4902_,
		_w4912_,
		_w4948_
	);
	LUT2 #(
		.INIT('h2)
	) name3947 (
		_w4947_,
		_w4948_,
		_w4949_
	);
	LUT2 #(
		.INIT('h1)
	) name3948 (
		_w4946_,
		_w4949_,
		_w4950_
	);
	LUT2 #(
		.INIT('h4)
	) name3949 (
		_w4925_,
		_w4933_,
		_w4951_
	);
	LUT2 #(
		.INIT('h2)
	) name3950 (
		_w4931_,
		_w4951_,
		_w4952_
	);
	LUT2 #(
		.INIT('h1)
	) name3951 (
		_w4934_,
		_w4952_,
		_w4953_
	);
	LUT2 #(
		.INIT('h1)
	) name3952 (
		_w4950_,
		_w4953_,
		_w4954_
	);
	LUT2 #(
		.INIT('h1)
	) name3953 (
		_w4902_,
		_w4914_,
		_w4955_
	);
	LUT2 #(
		.INIT('h1)
	) name3954 (
		_w4912_,
		_w4955_,
		_w4956_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		_w4950_,
		_w4953_,
		_w4957_
	);
	LUT2 #(
		.INIT('h1)
	) name3956 (
		_w4956_,
		_w4957_,
		_w4958_
	);
	LUT2 #(
		.INIT('h1)
	) name3957 (
		_w4954_,
		_w4958_,
		_w4959_
	);
	LUT2 #(
		.INIT('h8)
	) name3958 (
		\A[253] ,
		\A[254] ,
		_w4960_
	);
	LUT2 #(
		.INIT('h1)
	) name3959 (
		\A[253] ,
		\A[254] ,
		_w4961_
	);
	LUT2 #(
		.INIT('h1)
	) name3960 (
		_w4960_,
		_w4961_,
		_w4962_
	);
	LUT2 #(
		.INIT('h8)
	) name3961 (
		\A[255] ,
		_w4962_,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name3962 (
		\A[255] ,
		_w4962_,
		_w4964_
	);
	LUT2 #(
		.INIT('h1)
	) name3963 (
		_w4963_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h8)
	) name3964 (
		\A[256] ,
		\A[257] ,
		_w4966_
	);
	LUT2 #(
		.INIT('h1)
	) name3965 (
		\A[256] ,
		\A[257] ,
		_w4967_
	);
	LUT2 #(
		.INIT('h1)
	) name3966 (
		_w4966_,
		_w4967_,
		_w4968_
	);
	LUT2 #(
		.INIT('h8)
	) name3967 (
		\A[258] ,
		_w4968_,
		_w4969_
	);
	LUT2 #(
		.INIT('h1)
	) name3968 (
		\A[258] ,
		_w4968_,
		_w4970_
	);
	LUT2 #(
		.INIT('h1)
	) name3969 (
		_w4969_,
		_w4970_,
		_w4971_
	);
	LUT2 #(
		.INIT('h8)
	) name3970 (
		_w4965_,
		_w4971_,
		_w4972_
	);
	LUT2 #(
		.INIT('h1)
	) name3971 (
		_w4965_,
		_w4971_,
		_w4973_
	);
	LUT2 #(
		.INIT('h1)
	) name3972 (
		_w4972_,
		_w4973_,
		_w4974_
	);
	LUT2 #(
		.INIT('h8)
	) name3973 (
		\A[247] ,
		\A[248] ,
		_w4975_
	);
	LUT2 #(
		.INIT('h1)
	) name3974 (
		\A[247] ,
		\A[248] ,
		_w4976_
	);
	LUT2 #(
		.INIT('h1)
	) name3975 (
		_w4975_,
		_w4976_,
		_w4977_
	);
	LUT2 #(
		.INIT('h8)
	) name3976 (
		\A[249] ,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h1)
	) name3977 (
		\A[249] ,
		_w4977_,
		_w4979_
	);
	LUT2 #(
		.INIT('h1)
	) name3978 (
		_w4978_,
		_w4979_,
		_w4980_
	);
	LUT2 #(
		.INIT('h8)
	) name3979 (
		\A[250] ,
		\A[251] ,
		_w4981_
	);
	LUT2 #(
		.INIT('h1)
	) name3980 (
		\A[250] ,
		\A[251] ,
		_w4982_
	);
	LUT2 #(
		.INIT('h1)
	) name3981 (
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT2 #(
		.INIT('h8)
	) name3982 (
		\A[252] ,
		_w4983_,
		_w4984_
	);
	LUT2 #(
		.INIT('h1)
	) name3983 (
		\A[252] ,
		_w4983_,
		_w4985_
	);
	LUT2 #(
		.INIT('h1)
	) name3984 (
		_w4984_,
		_w4985_,
		_w4986_
	);
	LUT2 #(
		.INIT('h8)
	) name3985 (
		_w4980_,
		_w4986_,
		_w4987_
	);
	LUT2 #(
		.INIT('h1)
	) name3986 (
		_w4980_,
		_w4986_,
		_w4988_
	);
	LUT2 #(
		.INIT('h1)
	) name3987 (
		_w4987_,
		_w4988_,
		_w4989_
	);
	LUT2 #(
		.INIT('h8)
	) name3988 (
		_w4974_,
		_w4989_,
		_w4990_
	);
	LUT2 #(
		.INIT('h1)
	) name3989 (
		_w4960_,
		_w4963_,
		_w4991_
	);
	LUT2 #(
		.INIT('h1)
	) name3990 (
		_w4966_,
		_w4969_,
		_w4992_
	);
	LUT2 #(
		.INIT('h4)
	) name3991 (
		_w4972_,
		_w4992_,
		_w4993_
	);
	LUT2 #(
		.INIT('h8)
	) name3992 (
		_w4966_,
		_w4972_,
		_w4994_
	);
	LUT2 #(
		.INIT('h1)
	) name3993 (
		_w4993_,
		_w4994_,
		_w4995_
	);
	LUT2 #(
		.INIT('h2)
	) name3994 (
		_w4991_,
		_w4995_,
		_w4996_
	);
	LUT2 #(
		.INIT('h4)
	) name3995 (
		_w4991_,
		_w4995_,
		_w4997_
	);
	LUT2 #(
		.INIT('h1)
	) name3996 (
		_w4996_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h1)
	) name3997 (
		_w4990_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h1)
	) name3998 (
		_w4975_,
		_w4978_,
		_w5000_
	);
	LUT2 #(
		.INIT('h8)
	) name3999 (
		_w4981_,
		_w4987_,
		_w5001_
	);
	LUT2 #(
		.INIT('h1)
	) name4000 (
		_w4981_,
		_w4984_,
		_w5002_
	);
	LUT2 #(
		.INIT('h4)
	) name4001 (
		_w4987_,
		_w5002_,
		_w5003_
	);
	LUT2 #(
		.INIT('h1)
	) name4002 (
		_w5001_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h2)
	) name4003 (
		_w5000_,
		_w5004_,
		_w5005_
	);
	LUT2 #(
		.INIT('h4)
	) name4004 (
		_w5000_,
		_w5004_,
		_w5006_
	);
	LUT2 #(
		.INIT('h1)
	) name4005 (
		_w5005_,
		_w5006_,
		_w5007_
	);
	LUT2 #(
		.INIT('h4)
	) name4006 (
		_w4999_,
		_w5007_,
		_w5008_
	);
	LUT2 #(
		.INIT('h8)
	) name4007 (
		_w4990_,
		_w4998_,
		_w5009_
	);
	LUT2 #(
		.INIT('h1)
	) name4008 (
		_w4991_,
		_w4992_,
		_w5010_
	);
	LUT2 #(
		.INIT('h4)
	) name4009 (
		_w5000_,
		_w5001_,
		_w5011_
	);
	LUT2 #(
		.INIT('h1)
	) name4010 (
		_w5010_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h8)
	) name4011 (
		_w5009_,
		_w5012_,
		_w5013_
	);
	LUT2 #(
		.INIT('h1)
	) name4012 (
		_w5008_,
		_w5013_,
		_w5014_
	);
	LUT2 #(
		.INIT('h1)
	) name4013 (
		_w4991_,
		_w4993_,
		_w5015_
	);
	LUT2 #(
		.INIT('h1)
	) name4014 (
		_w4994_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w5014_,
		_w5016_,
		_w5017_
	);
	LUT2 #(
		.INIT('h1)
	) name4016 (
		_w5000_,
		_w5003_,
		_w5018_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		_w5001_,
		_w5018_,
		_w5019_
	);
	LUT2 #(
		.INIT('h8)
	) name4018 (
		_w5014_,
		_w5016_,
		_w5020_
	);
	LUT2 #(
		.INIT('h1)
	) name4019 (
		_w5019_,
		_w5020_,
		_w5021_
	);
	LUT2 #(
		.INIT('h1)
	) name4020 (
		_w5017_,
		_w5021_,
		_w5022_
	);
	LUT2 #(
		.INIT('h1)
	) name4021 (
		_w4959_,
		_w5022_,
		_w5023_
	);
	LUT2 #(
		.INIT('h8)
	) name4022 (
		_w4959_,
		_w5022_,
		_w5024_
	);
	LUT2 #(
		.INIT('h1)
	) name4023 (
		_w5017_,
		_w5020_,
		_w5025_
	);
	LUT2 #(
		.INIT('h2)
	) name4024 (
		_w5019_,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h4)
	) name4025 (
		_w5019_,
		_w5025_,
		_w5027_
	);
	LUT2 #(
		.INIT('h1)
	) name4026 (
		_w5026_,
		_w5027_,
		_w5028_
	);
	LUT2 #(
		.INIT('h1)
	) name4027 (
		_w4954_,
		_w4957_,
		_w5029_
	);
	LUT2 #(
		.INIT('h2)
	) name4028 (
		_w4956_,
		_w5029_,
		_w5030_
	);
	LUT2 #(
		.INIT('h4)
	) name4029 (
		_w4956_,
		_w5029_,
		_w5031_
	);
	LUT2 #(
		.INIT('h1)
	) name4030 (
		_w5030_,
		_w5031_,
		_w5032_
	);
	LUT2 #(
		.INIT('h1)
	) name4031 (
		_w5028_,
		_w5032_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name4032 (
		_w4939_,
		_w4941_,
		_w5034_
	);
	LUT2 #(
		.INIT('h1)
	) name4033 (
		_w4942_,
		_w5034_,
		_w5035_
	);
	LUT2 #(
		.INIT('h1)
	) name4034 (
		_w4974_,
		_w4989_,
		_w5036_
	);
	LUT2 #(
		.INIT('h1)
	) name4035 (
		_w4990_,
		_w5036_,
		_w5037_
	);
	LUT2 #(
		.INIT('h8)
	) name4036 (
		_w5035_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h2)
	) name4037 (
		_w4946_,
		_w4949_,
		_w5039_
	);
	LUT2 #(
		.INIT('h1)
	) name4038 (
		_w4945_,
		_w4947_,
		_w5040_
	);
	LUT2 #(
		.INIT('h1)
	) name4039 (
		_w4918_,
		_w5040_,
		_w5041_
	);
	LUT2 #(
		.INIT('h1)
	) name4040 (
		_w5039_,
		_w5041_,
		_w5042_
	);
	LUT2 #(
		.INIT('h1)
	) name4041 (
		_w5038_,
		_w5042_,
		_w5043_
	);
	LUT2 #(
		.INIT('h2)
	) name4042 (
		_w5008_,
		_w5013_,
		_w5044_
	);
	LUT2 #(
		.INIT('h1)
	) name4043 (
		_w4999_,
		_w5009_,
		_w5045_
	);
	LUT2 #(
		.INIT('h1)
	) name4044 (
		_w5007_,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h1)
	) name4045 (
		_w5044_,
		_w5046_,
		_w5047_
	);
	LUT2 #(
		.INIT('h8)
	) name4046 (
		_w5038_,
		_w5042_,
		_w5048_
	);
	LUT2 #(
		.INIT('h1)
	) name4047 (
		_w5047_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h1)
	) name4048 (
		_w5043_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h8)
	) name4049 (
		_w5028_,
		_w5032_,
		_w5051_
	);
	LUT2 #(
		.INIT('h1)
	) name4050 (
		_w5050_,
		_w5051_,
		_w5052_
	);
	LUT2 #(
		.INIT('h1)
	) name4051 (
		_w5033_,
		_w5052_,
		_w5053_
	);
	LUT2 #(
		.INIT('h4)
	) name4052 (
		_w5024_,
		_w5053_,
		_w5054_
	);
	LUT2 #(
		.INIT('h1)
	) name4053 (
		_w5023_,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('h8)
	) name4054 (
		\A[235] ,
		\A[236] ,
		_w5056_
	);
	LUT2 #(
		.INIT('h1)
	) name4055 (
		\A[235] ,
		\A[236] ,
		_w5057_
	);
	LUT2 #(
		.INIT('h1)
	) name4056 (
		_w5056_,
		_w5057_,
		_w5058_
	);
	LUT2 #(
		.INIT('h8)
	) name4057 (
		\A[237] ,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h1)
	) name4058 (
		_w5056_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h8)
	) name4059 (
		\A[238] ,
		\A[239] ,
		_w5061_
	);
	LUT2 #(
		.INIT('h1)
	) name4060 (
		\A[237] ,
		_w5058_,
		_w5062_
	);
	LUT2 #(
		.INIT('h1)
	) name4061 (
		_w5059_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h1)
	) name4062 (
		\A[238] ,
		\A[239] ,
		_w5064_
	);
	LUT2 #(
		.INIT('h1)
	) name4063 (
		_w5061_,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('h8)
	) name4064 (
		\A[240] ,
		_w5065_,
		_w5066_
	);
	LUT2 #(
		.INIT('h1)
	) name4065 (
		\A[240] ,
		_w5065_,
		_w5067_
	);
	LUT2 #(
		.INIT('h1)
	) name4066 (
		_w5066_,
		_w5067_,
		_w5068_
	);
	LUT2 #(
		.INIT('h8)
	) name4067 (
		_w5063_,
		_w5068_,
		_w5069_
	);
	LUT2 #(
		.INIT('h8)
	) name4068 (
		_w5061_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h1)
	) name4069 (
		_w5061_,
		_w5066_,
		_w5071_
	);
	LUT2 #(
		.INIT('h4)
	) name4070 (
		_w5069_,
		_w5071_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name4071 (
		_w5070_,
		_w5072_,
		_w5073_
	);
	LUT2 #(
		.INIT('h2)
	) name4072 (
		_w5060_,
		_w5073_,
		_w5074_
	);
	LUT2 #(
		.INIT('h4)
	) name4073 (
		_w5060_,
		_w5073_,
		_w5075_
	);
	LUT2 #(
		.INIT('h1)
	) name4074 (
		_w5074_,
		_w5075_,
		_w5076_
	);
	LUT2 #(
		.INIT('h8)
	) name4075 (
		\A[241] ,
		\A[242] ,
		_w5077_
	);
	LUT2 #(
		.INIT('h1)
	) name4076 (
		\A[241] ,
		\A[242] ,
		_w5078_
	);
	LUT2 #(
		.INIT('h1)
	) name4077 (
		_w5077_,
		_w5078_,
		_w5079_
	);
	LUT2 #(
		.INIT('h8)
	) name4078 (
		\A[243] ,
		_w5079_,
		_w5080_
	);
	LUT2 #(
		.INIT('h1)
	) name4079 (
		\A[243] ,
		_w5079_,
		_w5081_
	);
	LUT2 #(
		.INIT('h1)
	) name4080 (
		_w5080_,
		_w5081_,
		_w5082_
	);
	LUT2 #(
		.INIT('h8)
	) name4081 (
		\A[244] ,
		\A[245] ,
		_w5083_
	);
	LUT2 #(
		.INIT('h1)
	) name4082 (
		\A[244] ,
		\A[245] ,
		_w5084_
	);
	LUT2 #(
		.INIT('h1)
	) name4083 (
		_w5083_,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h8)
	) name4084 (
		\A[246] ,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('h1)
	) name4085 (
		\A[246] ,
		_w5085_,
		_w5087_
	);
	LUT2 #(
		.INIT('h1)
	) name4086 (
		_w5086_,
		_w5087_,
		_w5088_
	);
	LUT2 #(
		.INIT('h8)
	) name4087 (
		_w5082_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h1)
	) name4088 (
		_w5083_,
		_w5086_,
		_w5090_
	);
	LUT2 #(
		.INIT('h1)
	) name4089 (
		_w5077_,
		_w5080_,
		_w5091_
	);
	LUT2 #(
		.INIT('h1)
	) name4090 (
		_w5090_,
		_w5091_,
		_w5092_
	);
	LUT2 #(
		.INIT('h8)
	) name4091 (
		_w5090_,
		_w5091_,
		_w5093_
	);
	LUT2 #(
		.INIT('h1)
	) name4092 (
		_w5092_,
		_w5093_,
		_w5094_
	);
	LUT2 #(
		.INIT('h4)
	) name4093 (
		_w5089_,
		_w5094_,
		_w5095_
	);
	LUT2 #(
		.INIT('h1)
	) name4094 (
		_w5063_,
		_w5068_,
		_w5096_
	);
	LUT2 #(
		.INIT('h1)
	) name4095 (
		_w5069_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h1)
	) name4096 (
		_w5082_,
		_w5088_,
		_w5098_
	);
	LUT2 #(
		.INIT('h1)
	) name4097 (
		_w5089_,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h8)
	) name4098 (
		_w5097_,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('h2)
	) name4099 (
		_w5089_,
		_w5094_,
		_w5101_
	);
	LUT2 #(
		.INIT('h1)
	) name4100 (
		_w5095_,
		_w5100_,
		_w5102_
	);
	LUT2 #(
		.INIT('h4)
	) name4101 (
		_w5101_,
		_w5102_,
		_w5103_
	);
	LUT2 #(
		.INIT('h2)
	) name4102 (
		_w5076_,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h8)
	) name4103 (
		_w5094_,
		_w5100_,
		_w5105_
	);
	LUT2 #(
		.INIT('h4)
	) name4104 (
		_w5060_,
		_w5070_,
		_w5106_
	);
	LUT2 #(
		.INIT('h2)
	) name4105 (
		_w5105_,
		_w5106_,
		_w5107_
	);
	LUT2 #(
		.INIT('h1)
	) name4106 (
		_w5104_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h4)
	) name4107 (
		_w5083_,
		_w5091_,
		_w5109_
	);
	LUT2 #(
		.INIT('h2)
	) name4108 (
		_w5089_,
		_w5109_,
		_w5110_
	);
	LUT2 #(
		.INIT('h1)
	) name4109 (
		_w5092_,
		_w5110_,
		_w5111_
	);
	LUT2 #(
		.INIT('h1)
	) name4110 (
		_w5108_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h1)
	) name4111 (
		_w5060_,
		_w5072_,
		_w5113_
	);
	LUT2 #(
		.INIT('h1)
	) name4112 (
		_w5070_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h8)
	) name4113 (
		_w5108_,
		_w5111_,
		_w5115_
	);
	LUT2 #(
		.INIT('h1)
	) name4114 (
		_w5114_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('h1)
	) name4115 (
		_w5112_,
		_w5116_,
		_w5117_
	);
	LUT2 #(
		.INIT('h8)
	) name4116 (
		\A[229] ,
		\A[230] ,
		_w5118_
	);
	LUT2 #(
		.INIT('h1)
	) name4117 (
		\A[229] ,
		\A[230] ,
		_w5119_
	);
	LUT2 #(
		.INIT('h1)
	) name4118 (
		_w5118_,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('h8)
	) name4119 (
		\A[231] ,
		_w5120_,
		_w5121_
	);
	LUT2 #(
		.INIT('h1)
	) name4120 (
		\A[231] ,
		_w5120_,
		_w5122_
	);
	LUT2 #(
		.INIT('h1)
	) name4121 (
		_w5121_,
		_w5122_,
		_w5123_
	);
	LUT2 #(
		.INIT('h8)
	) name4122 (
		\A[232] ,
		\A[233] ,
		_w5124_
	);
	LUT2 #(
		.INIT('h1)
	) name4123 (
		\A[232] ,
		\A[233] ,
		_w5125_
	);
	LUT2 #(
		.INIT('h1)
	) name4124 (
		_w5124_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h8)
	) name4125 (
		\A[234] ,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h1)
	) name4126 (
		\A[234] ,
		_w5126_,
		_w5128_
	);
	LUT2 #(
		.INIT('h1)
	) name4127 (
		_w5127_,
		_w5128_,
		_w5129_
	);
	LUT2 #(
		.INIT('h8)
	) name4128 (
		_w5123_,
		_w5129_,
		_w5130_
	);
	LUT2 #(
		.INIT('h1)
	) name4129 (
		_w5123_,
		_w5129_,
		_w5131_
	);
	LUT2 #(
		.INIT('h1)
	) name4130 (
		_w5130_,
		_w5131_,
		_w5132_
	);
	LUT2 #(
		.INIT('h8)
	) name4131 (
		\A[223] ,
		\A[224] ,
		_w5133_
	);
	LUT2 #(
		.INIT('h1)
	) name4132 (
		\A[223] ,
		\A[224] ,
		_w5134_
	);
	LUT2 #(
		.INIT('h1)
	) name4133 (
		_w5133_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h8)
	) name4134 (
		\A[225] ,
		_w5135_,
		_w5136_
	);
	LUT2 #(
		.INIT('h1)
	) name4135 (
		\A[225] ,
		_w5135_,
		_w5137_
	);
	LUT2 #(
		.INIT('h1)
	) name4136 (
		_w5136_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h8)
	) name4137 (
		\A[226] ,
		\A[227] ,
		_w5139_
	);
	LUT2 #(
		.INIT('h1)
	) name4138 (
		\A[226] ,
		\A[227] ,
		_w5140_
	);
	LUT2 #(
		.INIT('h1)
	) name4139 (
		_w5139_,
		_w5140_,
		_w5141_
	);
	LUT2 #(
		.INIT('h8)
	) name4140 (
		\A[228] ,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h1)
	) name4141 (
		\A[228] ,
		_w5141_,
		_w5143_
	);
	LUT2 #(
		.INIT('h1)
	) name4142 (
		_w5142_,
		_w5143_,
		_w5144_
	);
	LUT2 #(
		.INIT('h8)
	) name4143 (
		_w5138_,
		_w5144_,
		_w5145_
	);
	LUT2 #(
		.INIT('h1)
	) name4144 (
		_w5138_,
		_w5144_,
		_w5146_
	);
	LUT2 #(
		.INIT('h1)
	) name4145 (
		_w5145_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('h8)
	) name4146 (
		_w5132_,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h1)
	) name4147 (
		_w5124_,
		_w5127_,
		_w5149_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		_w5118_,
		_w5121_,
		_w5150_
	);
	LUT2 #(
		.INIT('h1)
	) name4149 (
		_w5149_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h8)
	) name4150 (
		_w5149_,
		_w5150_,
		_w5152_
	);
	LUT2 #(
		.INIT('h1)
	) name4151 (
		_w5151_,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		_w5148_,
		_w5153_,
		_w5154_
	);
	LUT2 #(
		.INIT('h1)
	) name4153 (
		_w5139_,
		_w5142_,
		_w5155_
	);
	LUT2 #(
		.INIT('h1)
	) name4154 (
		_w5133_,
		_w5136_,
		_w5156_
	);
	LUT2 #(
		.INIT('h8)
	) name4155 (
		_w5155_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h1)
	) name4156 (
		_w5155_,
		_w5156_,
		_w5158_
	);
	LUT2 #(
		.INIT('h1)
	) name4157 (
		_w5157_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h2)
	) name4158 (
		_w5145_,
		_w5159_,
		_w5160_
	);
	LUT2 #(
		.INIT('h4)
	) name4159 (
		_w5145_,
		_w5159_,
		_w5161_
	);
	LUT2 #(
		.INIT('h1)
	) name4160 (
		_w5160_,
		_w5161_,
		_w5162_
	);
	LUT2 #(
		.INIT('h4)
	) name4161 (
		_w5154_,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h4)
	) name4162 (
		_w5130_,
		_w5153_,
		_w5164_
	);
	LUT2 #(
		.INIT('h2)
	) name4163 (
		_w5130_,
		_w5153_,
		_w5165_
	);
	LUT2 #(
		.INIT('h1)
	) name4164 (
		_w5148_,
		_w5164_,
		_w5166_
	);
	LUT2 #(
		.INIT('h4)
	) name4165 (
		_w5165_,
		_w5166_,
		_w5167_
	);
	LUT2 #(
		.INIT('h1)
	) name4166 (
		_w5163_,
		_w5167_,
		_w5168_
	);
	LUT2 #(
		.INIT('h1)
	) name4167 (
		_w5130_,
		_w5151_,
		_w5169_
	);
	LUT2 #(
		.INIT('h1)
	) name4168 (
		_w5152_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h1)
	) name4169 (
		_w5168_,
		_w5170_,
		_w5171_
	);
	LUT2 #(
		.INIT('h8)
	) name4170 (
		_w5168_,
		_w5170_,
		_w5172_
	);
	LUT2 #(
		.INIT('h1)
	) name4171 (
		_w5145_,
		_w5158_,
		_w5173_
	);
	LUT2 #(
		.INIT('h1)
	) name4172 (
		_w5157_,
		_w5173_,
		_w5174_
	);
	LUT2 #(
		.INIT('h1)
	) name4173 (
		_w5172_,
		_w5174_,
		_w5175_
	);
	LUT2 #(
		.INIT('h1)
	) name4174 (
		_w5171_,
		_w5175_,
		_w5176_
	);
	LUT2 #(
		.INIT('h4)
	) name4175 (
		_w5117_,
		_w5176_,
		_w5177_
	);
	LUT2 #(
		.INIT('h2)
	) name4176 (
		_w5117_,
		_w5176_,
		_w5178_
	);
	LUT2 #(
		.INIT('h1)
	) name4177 (
		_w5112_,
		_w5115_,
		_w5179_
	);
	LUT2 #(
		.INIT('h2)
	) name4178 (
		_w5114_,
		_w5179_,
		_w5180_
	);
	LUT2 #(
		.INIT('h4)
	) name4179 (
		_w5114_,
		_w5179_,
		_w5181_
	);
	LUT2 #(
		.INIT('h1)
	) name4180 (
		_w5180_,
		_w5181_,
		_w5182_
	);
	LUT2 #(
		.INIT('h1)
	) name4181 (
		_w5171_,
		_w5172_,
		_w5183_
	);
	LUT2 #(
		.INIT('h4)
	) name4182 (
		_w5174_,
		_w5183_,
		_w5184_
	);
	LUT2 #(
		.INIT('h2)
	) name4183 (
		_w5174_,
		_w5183_,
		_w5185_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		_w5184_,
		_w5185_,
		_w5186_
	);
	LUT2 #(
		.INIT('h2)
	) name4185 (
		_w5182_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h4)
	) name4186 (
		_w5182_,
		_w5186_,
		_w5188_
	);
	LUT2 #(
		.INIT('h1)
	) name4187 (
		_w5097_,
		_w5099_,
		_w5189_
	);
	LUT2 #(
		.INIT('h1)
	) name4188 (
		_w5100_,
		_w5189_,
		_w5190_
	);
	LUT2 #(
		.INIT('h1)
	) name4189 (
		_w5132_,
		_w5147_,
		_w5191_
	);
	LUT2 #(
		.INIT('h1)
	) name4190 (
		_w5148_,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h8)
	) name4191 (
		_w5190_,
		_w5192_,
		_w5193_
	);
	LUT2 #(
		.INIT('h2)
	) name4192 (
		_w5104_,
		_w5107_,
		_w5194_
	);
	LUT2 #(
		.INIT('h1)
	) name4193 (
		_w5103_,
		_w5105_,
		_w5195_
	);
	LUT2 #(
		.INIT('h1)
	) name4194 (
		_w5076_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h1)
	) name4195 (
		_w5194_,
		_w5196_,
		_w5197_
	);
	LUT2 #(
		.INIT('h8)
	) name4196 (
		_w5193_,
		_w5197_,
		_w5198_
	);
	LUT2 #(
		.INIT('h1)
	) name4197 (
		_w5193_,
		_w5197_,
		_w5199_
	);
	LUT2 #(
		.INIT('h1)
	) name4198 (
		_w5154_,
		_w5167_,
		_w5200_
	);
	LUT2 #(
		.INIT('h8)
	) name4199 (
		_w5162_,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h1)
	) name4200 (
		_w5162_,
		_w5200_,
		_w5202_
	);
	LUT2 #(
		.INIT('h1)
	) name4201 (
		_w5201_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h1)
	) name4202 (
		_w5199_,
		_w5203_,
		_w5204_
	);
	LUT2 #(
		.INIT('h1)
	) name4203 (
		_w5198_,
		_w5204_,
		_w5205_
	);
	LUT2 #(
		.INIT('h1)
	) name4204 (
		_w5188_,
		_w5205_,
		_w5206_
	);
	LUT2 #(
		.INIT('h1)
	) name4205 (
		_w5187_,
		_w5206_,
		_w5207_
	);
	LUT2 #(
		.INIT('h1)
	) name4206 (
		_w5178_,
		_w5207_,
		_w5208_
	);
	LUT2 #(
		.INIT('h1)
	) name4207 (
		_w5177_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		_w5055_,
		_w5209_,
		_w5210_
	);
	LUT2 #(
		.INIT('h8)
	) name4209 (
		_w5055_,
		_w5209_,
		_w5211_
	);
	LUT2 #(
		.INIT('h1)
	) name4210 (
		_w5023_,
		_w5024_,
		_w5212_
	);
	LUT2 #(
		.INIT('h2)
	) name4211 (
		_w5053_,
		_w5212_,
		_w5213_
	);
	LUT2 #(
		.INIT('h4)
	) name4212 (
		_w5053_,
		_w5212_,
		_w5214_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w5213_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h1)
	) name4214 (
		_w5177_,
		_w5178_,
		_w5216_
	);
	LUT2 #(
		.INIT('h4)
	) name4215 (
		_w5207_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h2)
	) name4216 (
		_w5207_,
		_w5216_,
		_w5218_
	);
	LUT2 #(
		.INIT('h1)
	) name4217 (
		_w5217_,
		_w5218_,
		_w5219_
	);
	LUT2 #(
		.INIT('h2)
	) name4218 (
		_w5215_,
		_w5219_,
		_w5220_
	);
	LUT2 #(
		.INIT('h4)
	) name4219 (
		_w5215_,
		_w5219_,
		_w5221_
	);
	LUT2 #(
		.INIT('h1)
	) name4220 (
		_w5033_,
		_w5051_,
		_w5222_
	);
	LUT2 #(
		.INIT('h8)
	) name4221 (
		_w5050_,
		_w5222_,
		_w5223_
	);
	LUT2 #(
		.INIT('h1)
	) name4222 (
		_w5050_,
		_w5222_,
		_w5224_
	);
	LUT2 #(
		.INIT('h1)
	) name4223 (
		_w5223_,
		_w5224_,
		_w5225_
	);
	LUT2 #(
		.INIT('h1)
	) name4224 (
		_w5187_,
		_w5188_,
		_w5226_
	);
	LUT2 #(
		.INIT('h4)
	) name4225 (
		_w5205_,
		_w5226_,
		_w5227_
	);
	LUT2 #(
		.INIT('h2)
	) name4226 (
		_w5205_,
		_w5226_,
		_w5228_
	);
	LUT2 #(
		.INIT('h1)
	) name4227 (
		_w5227_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('h8)
	) name4228 (
		_w5225_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h1)
	) name4229 (
		_w5225_,
		_w5229_,
		_w5231_
	);
	LUT2 #(
		.INIT('h1)
	) name4230 (
		_w5035_,
		_w5037_,
		_w5232_
	);
	LUT2 #(
		.INIT('h1)
	) name4231 (
		_w5038_,
		_w5232_,
		_w5233_
	);
	LUT2 #(
		.INIT('h1)
	) name4232 (
		_w5190_,
		_w5192_,
		_w5234_
	);
	LUT2 #(
		.INIT('h1)
	) name4233 (
		_w5193_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h8)
	) name4234 (
		_w5233_,
		_w5235_,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name4235 (
		_w5043_,
		_w5048_,
		_w5237_
	);
	LUT2 #(
		.INIT('h2)
	) name4236 (
		_w5047_,
		_w5237_,
		_w5238_
	);
	LUT2 #(
		.INIT('h4)
	) name4237 (
		_w5047_,
		_w5237_,
		_w5239_
	);
	LUT2 #(
		.INIT('h1)
	) name4238 (
		_w5238_,
		_w5239_,
		_w5240_
	);
	LUT2 #(
		.INIT('h2)
	) name4239 (
		_w5236_,
		_w5240_,
		_w5241_
	);
	LUT2 #(
		.INIT('h4)
	) name4240 (
		_w5236_,
		_w5240_,
		_w5242_
	);
	LUT2 #(
		.INIT('h1)
	) name4241 (
		_w5198_,
		_w5199_,
		_w5243_
	);
	LUT2 #(
		.INIT('h4)
	) name4242 (
		_w5203_,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h2)
	) name4243 (
		_w5203_,
		_w5243_,
		_w5245_
	);
	LUT2 #(
		.INIT('h1)
	) name4244 (
		_w5244_,
		_w5245_,
		_w5246_
	);
	LUT2 #(
		.INIT('h4)
	) name4245 (
		_w5242_,
		_w5246_,
		_w5247_
	);
	LUT2 #(
		.INIT('h1)
	) name4246 (
		_w5241_,
		_w5247_,
		_w5248_
	);
	LUT2 #(
		.INIT('h1)
	) name4247 (
		_w5231_,
		_w5248_,
		_w5249_
	);
	LUT2 #(
		.INIT('h1)
	) name4248 (
		_w5230_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h4)
	) name4249 (
		_w5221_,
		_w5250_,
		_w5251_
	);
	LUT2 #(
		.INIT('h1)
	) name4250 (
		_w5220_,
		_w5251_,
		_w5252_
	);
	LUT2 #(
		.INIT('h4)
	) name4251 (
		_w5211_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h1)
	) name4252 (
		_w5210_,
		_w5253_,
		_w5254_
	);
	LUT2 #(
		.INIT('h1)
	) name4253 (
		_w4897_,
		_w5254_,
		_w5255_
	);
	LUT2 #(
		.INIT('h8)
	) name4254 (
		_w4897_,
		_w5254_,
		_w5256_
	);
	LUT2 #(
		.INIT('h1)
	) name4255 (
		_w5210_,
		_w5211_,
		_w5257_
	);
	LUT2 #(
		.INIT('h4)
	) name4256 (
		_w5252_,
		_w5257_,
		_w5258_
	);
	LUT2 #(
		.INIT('h2)
	) name4257 (
		_w5252_,
		_w5257_,
		_w5259_
	);
	LUT2 #(
		.INIT('h1)
	) name4258 (
		_w5258_,
		_w5259_,
		_w5260_
	);
	LUT2 #(
		.INIT('h1)
	) name4259 (
		_w4853_,
		_w4854_,
		_w5261_
	);
	LUT2 #(
		.INIT('h4)
	) name4260 (
		_w4895_,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('h2)
	) name4261 (
		_w4895_,
		_w5261_,
		_w5263_
	);
	LUT2 #(
		.INIT('h1)
	) name4262 (
		_w5262_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h2)
	) name4263 (
		_w5260_,
		_w5264_,
		_w5265_
	);
	LUT2 #(
		.INIT('h4)
	) name4264 (
		_w5260_,
		_w5264_,
		_w5266_
	);
	LUT2 #(
		.INIT('h1)
	) name4265 (
		_w4863_,
		_w4864_,
		_w5267_
	);
	LUT2 #(
		.INIT('h4)
	) name4266 (
		_w4893_,
		_w5267_,
		_w5268_
	);
	LUT2 #(
		.INIT('h2)
	) name4267 (
		_w4893_,
		_w5267_,
		_w5269_
	);
	LUT2 #(
		.INIT('h1)
	) name4268 (
		_w5268_,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h1)
	) name4269 (
		_w5220_,
		_w5221_,
		_w5271_
	);
	LUT2 #(
		.INIT('h4)
	) name4270 (
		_w5250_,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h2)
	) name4271 (
		_w5250_,
		_w5271_,
		_w5273_
	);
	LUT2 #(
		.INIT('h1)
	) name4272 (
		_w5272_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h1)
	) name4273 (
		_w5270_,
		_w5274_,
		_w5275_
	);
	LUT2 #(
		.INIT('h8)
	) name4274 (
		_w5270_,
		_w5274_,
		_w5276_
	);
	LUT2 #(
		.INIT('h1)
	) name4275 (
		_w4873_,
		_w4874_,
		_w5277_
	);
	LUT2 #(
		.INIT('h4)
	) name4276 (
		_w4891_,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h2)
	) name4277 (
		_w4891_,
		_w5277_,
		_w5279_
	);
	LUT2 #(
		.INIT('h1)
	) name4278 (
		_w5278_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h1)
	) name4279 (
		_w5230_,
		_w5231_,
		_w5281_
	);
	LUT2 #(
		.INIT('h4)
	) name4280 (
		_w5248_,
		_w5281_,
		_w5282_
	);
	LUT2 #(
		.INIT('h2)
	) name4281 (
		_w5248_,
		_w5281_,
		_w5283_
	);
	LUT2 #(
		.INIT('h1)
	) name4282 (
		_w5282_,
		_w5283_,
		_w5284_
	);
	LUT2 #(
		.INIT('h1)
	) name4283 (
		_w5280_,
		_w5284_,
		_w5285_
	);
	LUT2 #(
		.INIT('h8)
	) name4284 (
		_w5280_,
		_w5284_,
		_w5286_
	);
	LUT2 #(
		.INIT('h1)
	) name4285 (
		_w5233_,
		_w5235_,
		_w5287_
	);
	LUT2 #(
		.INIT('h1)
	) name4286 (
		_w5236_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h1)
	) name4287 (
		_w4876_,
		_w4878_,
		_w5289_
	);
	LUT2 #(
		.INIT('h1)
	) name4288 (
		_w4879_,
		_w5289_,
		_w5290_
	);
	LUT2 #(
		.INIT('h8)
	) name4289 (
		_w5288_,
		_w5290_,
		_w5291_
	);
	LUT2 #(
		.INIT('h1)
	) name4290 (
		_w5241_,
		_w5242_,
		_w5292_
	);
	LUT2 #(
		.INIT('h4)
	) name4291 (
		_w5246_,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('h2)
	) name4292 (
		_w5246_,
		_w5292_,
		_w5294_
	);
	LUT2 #(
		.INIT('h1)
	) name4293 (
		_w5293_,
		_w5294_,
		_w5295_
	);
	LUT2 #(
		.INIT('h2)
	) name4294 (
		_w5291_,
		_w5295_,
		_w5296_
	);
	LUT2 #(
		.INIT('h4)
	) name4295 (
		_w5291_,
		_w5295_,
		_w5297_
	);
	LUT2 #(
		.INIT('h1)
	) name4296 (
		_w4884_,
		_w4885_,
		_w5298_
	);
	LUT2 #(
		.INIT('h4)
	) name4297 (
		_w4889_,
		_w5298_,
		_w5299_
	);
	LUT2 #(
		.INIT('h2)
	) name4298 (
		_w4889_,
		_w5298_,
		_w5300_
	);
	LUT2 #(
		.INIT('h1)
	) name4299 (
		_w5299_,
		_w5300_,
		_w5301_
	);
	LUT2 #(
		.INIT('h1)
	) name4300 (
		_w5297_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h1)
	) name4301 (
		_w5296_,
		_w5302_,
		_w5303_
	);
	LUT2 #(
		.INIT('h4)
	) name4302 (
		_w5286_,
		_w5303_,
		_w5304_
	);
	LUT2 #(
		.INIT('h1)
	) name4303 (
		_w5285_,
		_w5304_,
		_w5305_
	);
	LUT2 #(
		.INIT('h1)
	) name4304 (
		_w5276_,
		_w5305_,
		_w5306_
	);
	LUT2 #(
		.INIT('h1)
	) name4305 (
		_w5275_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('h1)
	) name4306 (
		_w5266_,
		_w5307_,
		_w5308_
	);
	LUT2 #(
		.INIT('h1)
	) name4307 (
		_w5265_,
		_w5308_,
		_w5309_
	);
	LUT2 #(
		.INIT('h4)
	) name4308 (
		_w5256_,
		_w5309_,
		_w5310_
	);
	LUT2 #(
		.INIT('h1)
	) name4309 (
		_w5255_,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h8)
	) name4310 (
		\A[145] ,
		\A[146] ,
		_w5312_
	);
	LUT2 #(
		.INIT('h1)
	) name4311 (
		\A[145] ,
		\A[146] ,
		_w5313_
	);
	LUT2 #(
		.INIT('h1)
	) name4312 (
		_w5312_,
		_w5313_,
		_w5314_
	);
	LUT2 #(
		.INIT('h8)
	) name4313 (
		\A[147] ,
		_w5314_,
		_w5315_
	);
	LUT2 #(
		.INIT('h1)
	) name4314 (
		\A[147] ,
		_w5314_,
		_w5316_
	);
	LUT2 #(
		.INIT('h1)
	) name4315 (
		_w5315_,
		_w5316_,
		_w5317_
	);
	LUT2 #(
		.INIT('h8)
	) name4316 (
		\A[148] ,
		\A[149] ,
		_w5318_
	);
	LUT2 #(
		.INIT('h1)
	) name4317 (
		\A[148] ,
		\A[149] ,
		_w5319_
	);
	LUT2 #(
		.INIT('h1)
	) name4318 (
		_w5318_,
		_w5319_,
		_w5320_
	);
	LUT2 #(
		.INIT('h8)
	) name4319 (
		\A[150] ,
		_w5320_,
		_w5321_
	);
	LUT2 #(
		.INIT('h1)
	) name4320 (
		\A[150] ,
		_w5320_,
		_w5322_
	);
	LUT2 #(
		.INIT('h1)
	) name4321 (
		_w5321_,
		_w5322_,
		_w5323_
	);
	LUT2 #(
		.INIT('h8)
	) name4322 (
		_w5317_,
		_w5323_,
		_w5324_
	);
	LUT2 #(
		.INIT('h1)
	) name4323 (
		_w5317_,
		_w5323_,
		_w5325_
	);
	LUT2 #(
		.INIT('h1)
	) name4324 (
		_w5324_,
		_w5325_,
		_w5326_
	);
	LUT2 #(
		.INIT('h8)
	) name4325 (
		\A[139] ,
		\A[140] ,
		_w5327_
	);
	LUT2 #(
		.INIT('h1)
	) name4326 (
		\A[139] ,
		\A[140] ,
		_w5328_
	);
	LUT2 #(
		.INIT('h1)
	) name4327 (
		_w5327_,
		_w5328_,
		_w5329_
	);
	LUT2 #(
		.INIT('h8)
	) name4328 (
		\A[141] ,
		_w5329_,
		_w5330_
	);
	LUT2 #(
		.INIT('h1)
	) name4329 (
		\A[141] ,
		_w5329_,
		_w5331_
	);
	LUT2 #(
		.INIT('h1)
	) name4330 (
		_w5330_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h8)
	) name4331 (
		\A[142] ,
		\A[143] ,
		_w5333_
	);
	LUT2 #(
		.INIT('h1)
	) name4332 (
		\A[142] ,
		\A[143] ,
		_w5334_
	);
	LUT2 #(
		.INIT('h1)
	) name4333 (
		_w5333_,
		_w5334_,
		_w5335_
	);
	LUT2 #(
		.INIT('h8)
	) name4334 (
		\A[144] ,
		_w5335_,
		_w5336_
	);
	LUT2 #(
		.INIT('h1)
	) name4335 (
		\A[144] ,
		_w5335_,
		_w5337_
	);
	LUT2 #(
		.INIT('h1)
	) name4336 (
		_w5336_,
		_w5337_,
		_w5338_
	);
	LUT2 #(
		.INIT('h8)
	) name4337 (
		_w5332_,
		_w5338_,
		_w5339_
	);
	LUT2 #(
		.INIT('h1)
	) name4338 (
		_w5332_,
		_w5338_,
		_w5340_
	);
	LUT2 #(
		.INIT('h1)
	) name4339 (
		_w5339_,
		_w5340_,
		_w5341_
	);
	LUT2 #(
		.INIT('h8)
	) name4340 (
		_w5326_,
		_w5341_,
		_w5342_
	);
	LUT2 #(
		.INIT('h1)
	) name4341 (
		_w5318_,
		_w5321_,
		_w5343_
	);
	LUT2 #(
		.INIT('h1)
	) name4342 (
		_w5312_,
		_w5315_,
		_w5344_
	);
	LUT2 #(
		.INIT('h1)
	) name4343 (
		_w5343_,
		_w5344_,
		_w5345_
	);
	LUT2 #(
		.INIT('h8)
	) name4344 (
		_w5343_,
		_w5344_,
		_w5346_
	);
	LUT2 #(
		.INIT('h1)
	) name4345 (
		_w5345_,
		_w5346_,
		_w5347_
	);
	LUT2 #(
		.INIT('h8)
	) name4346 (
		_w5342_,
		_w5347_,
		_w5348_
	);
	LUT2 #(
		.INIT('h1)
	) name4347 (
		_w5327_,
		_w5330_,
		_w5349_
	);
	LUT2 #(
		.INIT('h1)
	) name4348 (
		_w5333_,
		_w5336_,
		_w5350_
	);
	LUT2 #(
		.INIT('h4)
	) name4349 (
		_w5339_,
		_w5350_,
		_w5351_
	);
	LUT2 #(
		.INIT('h8)
	) name4350 (
		_w5333_,
		_w5339_,
		_w5352_
	);
	LUT2 #(
		.INIT('h1)
	) name4351 (
		_w5351_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h2)
	) name4352 (
		_w5349_,
		_w5353_,
		_w5354_
	);
	LUT2 #(
		.INIT('h4)
	) name4353 (
		_w5349_,
		_w5353_,
		_w5355_
	);
	LUT2 #(
		.INIT('h1)
	) name4354 (
		_w5354_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h1)
	) name4355 (
		_w5348_,
		_w5356_,
		_w5357_
	);
	LUT2 #(
		.INIT('h4)
	) name4356 (
		_w5324_,
		_w5347_,
		_w5358_
	);
	LUT2 #(
		.INIT('h2)
	) name4357 (
		_w5324_,
		_w5347_,
		_w5359_
	);
	LUT2 #(
		.INIT('h1)
	) name4358 (
		_w5342_,
		_w5358_,
		_w5360_
	);
	LUT2 #(
		.INIT('h4)
	) name4359 (
		_w5359_,
		_w5360_,
		_w5361_
	);
	LUT2 #(
		.INIT('h1)
	) name4360 (
		_w5357_,
		_w5361_,
		_w5362_
	);
	LUT2 #(
		.INIT('h1)
	) name4361 (
		_w5324_,
		_w5345_,
		_w5363_
	);
	LUT2 #(
		.INIT('h1)
	) name4362 (
		_w5346_,
		_w5363_,
		_w5364_
	);
	LUT2 #(
		.INIT('h1)
	) name4363 (
		_w5362_,
		_w5364_,
		_w5365_
	);
	LUT2 #(
		.INIT('h8)
	) name4364 (
		_w5362_,
		_w5364_,
		_w5366_
	);
	LUT2 #(
		.INIT('h1)
	) name4365 (
		_w5349_,
		_w5351_,
		_w5367_
	);
	LUT2 #(
		.INIT('h1)
	) name4366 (
		_w5352_,
		_w5367_,
		_w5368_
	);
	LUT2 #(
		.INIT('h4)
	) name4367 (
		_w5366_,
		_w5368_,
		_w5369_
	);
	LUT2 #(
		.INIT('h1)
	) name4368 (
		_w5365_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h1)
	) name4369 (
		_w5365_,
		_w5366_,
		_w5371_
	);
	LUT2 #(
		.INIT('h4)
	) name4370 (
		_w5368_,
		_w5371_,
		_w5372_
	);
	LUT2 #(
		.INIT('h2)
	) name4371 (
		_w5368_,
		_w5371_,
		_w5373_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w5372_,
		_w5373_,
		_w5374_
	);
	LUT2 #(
		.INIT('h8)
	) name4373 (
		\A[130] ,
		\A[131] ,
		_w5375_
	);
	LUT2 #(
		.INIT('h8)
	) name4374 (
		\A[127] ,
		\A[128] ,
		_w5376_
	);
	LUT2 #(
		.INIT('h1)
	) name4375 (
		\A[127] ,
		\A[128] ,
		_w5377_
	);
	LUT2 #(
		.INIT('h1)
	) name4376 (
		_w5376_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h8)
	) name4377 (
		\A[129] ,
		_w5378_,
		_w5379_
	);
	LUT2 #(
		.INIT('h1)
	) name4378 (
		\A[129] ,
		_w5378_,
		_w5380_
	);
	LUT2 #(
		.INIT('h1)
	) name4379 (
		_w5379_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h1)
	) name4380 (
		\A[130] ,
		\A[131] ,
		_w5382_
	);
	LUT2 #(
		.INIT('h1)
	) name4381 (
		_w5375_,
		_w5382_,
		_w5383_
	);
	LUT2 #(
		.INIT('h8)
	) name4382 (
		\A[132] ,
		_w5383_,
		_w5384_
	);
	LUT2 #(
		.INIT('h1)
	) name4383 (
		\A[132] ,
		_w5383_,
		_w5385_
	);
	LUT2 #(
		.INIT('h1)
	) name4384 (
		_w5384_,
		_w5385_,
		_w5386_
	);
	LUT2 #(
		.INIT('h8)
	) name4385 (
		_w5381_,
		_w5386_,
		_w5387_
	);
	LUT2 #(
		.INIT('h8)
	) name4386 (
		_w5375_,
		_w5387_,
		_w5388_
	);
	LUT2 #(
		.INIT('h1)
	) name4387 (
		_w5376_,
		_w5379_,
		_w5389_
	);
	LUT2 #(
		.INIT('h1)
	) name4388 (
		_w5375_,
		_w5384_,
		_w5390_
	);
	LUT2 #(
		.INIT('h4)
	) name4389 (
		_w5387_,
		_w5390_,
		_w5391_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		_w5389_,
		_w5391_,
		_w5392_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		_w5388_,
		_w5392_,
		_w5393_
	);
	LUT2 #(
		.INIT('h8)
	) name4392 (
		\A[133] ,
		\A[134] ,
		_w5394_
	);
	LUT2 #(
		.INIT('h1)
	) name4393 (
		\A[133] ,
		\A[134] ,
		_w5395_
	);
	LUT2 #(
		.INIT('h1)
	) name4394 (
		_w5394_,
		_w5395_,
		_w5396_
	);
	LUT2 #(
		.INIT('h8)
	) name4395 (
		\A[135] ,
		_w5396_,
		_w5397_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		\A[135] ,
		_w5396_,
		_w5398_
	);
	LUT2 #(
		.INIT('h1)
	) name4397 (
		_w5397_,
		_w5398_,
		_w5399_
	);
	LUT2 #(
		.INIT('h8)
	) name4398 (
		\A[136] ,
		\A[137] ,
		_w5400_
	);
	LUT2 #(
		.INIT('h1)
	) name4399 (
		\A[136] ,
		\A[137] ,
		_w5401_
	);
	LUT2 #(
		.INIT('h1)
	) name4400 (
		_w5400_,
		_w5401_,
		_w5402_
	);
	LUT2 #(
		.INIT('h8)
	) name4401 (
		\A[138] ,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h1)
	) name4402 (
		\A[138] ,
		_w5402_,
		_w5404_
	);
	LUT2 #(
		.INIT('h1)
	) name4403 (
		_w5403_,
		_w5404_,
		_w5405_
	);
	LUT2 #(
		.INIT('h8)
	) name4404 (
		_w5399_,
		_w5405_,
		_w5406_
	);
	LUT2 #(
		.INIT('h1)
	) name4405 (
		_w5399_,
		_w5405_,
		_w5407_
	);
	LUT2 #(
		.INIT('h1)
	) name4406 (
		_w5406_,
		_w5407_,
		_w5408_
	);
	LUT2 #(
		.INIT('h1)
	) name4407 (
		_w5381_,
		_w5386_,
		_w5409_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		_w5387_,
		_w5409_,
		_w5410_
	);
	LUT2 #(
		.INIT('h8)
	) name4409 (
		_w5408_,
		_w5410_,
		_w5411_
	);
	LUT2 #(
		.INIT('h1)
	) name4410 (
		_w5400_,
		_w5403_,
		_w5412_
	);
	LUT2 #(
		.INIT('h1)
	) name4411 (
		_w5394_,
		_w5397_,
		_w5413_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w5412_,
		_w5413_,
		_w5414_
	);
	LUT2 #(
		.INIT('h8)
	) name4413 (
		_w5412_,
		_w5413_,
		_w5415_
	);
	LUT2 #(
		.INIT('h1)
	) name4414 (
		_w5414_,
		_w5415_,
		_w5416_
	);
	LUT2 #(
		.INIT('h8)
	) name4415 (
		_w5411_,
		_w5416_,
		_w5417_
	);
	LUT2 #(
		.INIT('h1)
	) name4416 (
		_w5388_,
		_w5391_,
		_w5418_
	);
	LUT2 #(
		.INIT('h2)
	) name4417 (
		_w5389_,
		_w5418_,
		_w5419_
	);
	LUT2 #(
		.INIT('h4)
	) name4418 (
		_w5389_,
		_w5418_,
		_w5420_
	);
	LUT2 #(
		.INIT('h1)
	) name4419 (
		_w5419_,
		_w5420_,
		_w5421_
	);
	LUT2 #(
		.INIT('h1)
	) name4420 (
		_w5417_,
		_w5421_,
		_w5422_
	);
	LUT2 #(
		.INIT('h4)
	) name4421 (
		_w5406_,
		_w5416_,
		_w5423_
	);
	LUT2 #(
		.INIT('h2)
	) name4422 (
		_w5406_,
		_w5416_,
		_w5424_
	);
	LUT2 #(
		.INIT('h1)
	) name4423 (
		_w5411_,
		_w5423_,
		_w5425_
	);
	LUT2 #(
		.INIT('h4)
	) name4424 (
		_w5424_,
		_w5425_,
		_w5426_
	);
	LUT2 #(
		.INIT('h1)
	) name4425 (
		_w5422_,
		_w5426_,
		_w5427_
	);
	LUT2 #(
		.INIT('h1)
	) name4426 (
		_w5406_,
		_w5414_,
		_w5428_
	);
	LUT2 #(
		.INIT('h1)
	) name4427 (
		_w5415_,
		_w5428_,
		_w5429_
	);
	LUT2 #(
		.INIT('h1)
	) name4428 (
		_w5427_,
		_w5429_,
		_w5430_
	);
	LUT2 #(
		.INIT('h8)
	) name4429 (
		_w5427_,
		_w5429_,
		_w5431_
	);
	LUT2 #(
		.INIT('h1)
	) name4430 (
		_w5430_,
		_w5431_,
		_w5432_
	);
	LUT2 #(
		.INIT('h2)
	) name4431 (
		_w5393_,
		_w5432_,
		_w5433_
	);
	LUT2 #(
		.INIT('h4)
	) name4432 (
		_w5393_,
		_w5432_,
		_w5434_
	);
	LUT2 #(
		.INIT('h1)
	) name4433 (
		_w5433_,
		_w5434_,
		_w5435_
	);
	LUT2 #(
		.INIT('h8)
	) name4434 (
		_w5374_,
		_w5435_,
		_w5436_
	);
	LUT2 #(
		.INIT('h1)
	) name4435 (
		_w5374_,
		_w5435_,
		_w5437_
	);
	LUT2 #(
		.INIT('h1)
	) name4436 (
		_w5326_,
		_w5341_,
		_w5438_
	);
	LUT2 #(
		.INIT('h1)
	) name4437 (
		_w5342_,
		_w5438_,
		_w5439_
	);
	LUT2 #(
		.INIT('h1)
	) name4438 (
		_w5408_,
		_w5410_,
		_w5440_
	);
	LUT2 #(
		.INIT('h1)
	) name4439 (
		_w5411_,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h8)
	) name4440 (
		_w5439_,
		_w5441_,
		_w5442_
	);
	LUT2 #(
		.INIT('h1)
	) name4441 (
		_w5348_,
		_w5361_,
		_w5443_
	);
	LUT2 #(
		.INIT('h4)
	) name4442 (
		_w5356_,
		_w5443_,
		_w5444_
	);
	LUT2 #(
		.INIT('h2)
	) name4443 (
		_w5356_,
		_w5443_,
		_w5445_
	);
	LUT2 #(
		.INIT('h1)
	) name4444 (
		_w5444_,
		_w5445_,
		_w5446_
	);
	LUT2 #(
		.INIT('h2)
	) name4445 (
		_w5442_,
		_w5446_,
		_w5447_
	);
	LUT2 #(
		.INIT('h4)
	) name4446 (
		_w5442_,
		_w5446_,
		_w5448_
	);
	LUT2 #(
		.INIT('h1)
	) name4447 (
		_w5417_,
		_w5426_,
		_w5449_
	);
	LUT2 #(
		.INIT('h4)
	) name4448 (
		_w5421_,
		_w5449_,
		_w5450_
	);
	LUT2 #(
		.INIT('h2)
	) name4449 (
		_w5421_,
		_w5449_,
		_w5451_
	);
	LUT2 #(
		.INIT('h1)
	) name4450 (
		_w5450_,
		_w5451_,
		_w5452_
	);
	LUT2 #(
		.INIT('h1)
	) name4451 (
		_w5448_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h1)
	) name4452 (
		_w5447_,
		_w5453_,
		_w5454_
	);
	LUT2 #(
		.INIT('h1)
	) name4453 (
		_w5437_,
		_w5454_,
		_w5455_
	);
	LUT2 #(
		.INIT('h1)
	) name4454 (
		_w5436_,
		_w5455_,
		_w5456_
	);
	LUT2 #(
		.INIT('h4)
	) name4455 (
		_w5370_,
		_w5456_,
		_w5457_
	);
	LUT2 #(
		.INIT('h2)
	) name4456 (
		_w5370_,
		_w5456_,
		_w5458_
	);
	LUT2 #(
		.INIT('h2)
	) name4457 (
		_w5393_,
		_w5431_,
		_w5459_
	);
	LUT2 #(
		.INIT('h1)
	) name4458 (
		_w5430_,
		_w5459_,
		_w5460_
	);
	LUT2 #(
		.INIT('h1)
	) name4459 (
		_w5458_,
		_w5460_,
		_w5461_
	);
	LUT2 #(
		.INIT('h1)
	) name4460 (
		_w5457_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('h8)
	) name4461 (
		\A[169] ,
		\A[170] ,
		_w5463_
	);
	LUT2 #(
		.INIT('h1)
	) name4462 (
		\A[169] ,
		\A[170] ,
		_w5464_
	);
	LUT2 #(
		.INIT('h1)
	) name4463 (
		_w5463_,
		_w5464_,
		_w5465_
	);
	LUT2 #(
		.INIT('h8)
	) name4464 (
		\A[171] ,
		_w5465_,
		_w5466_
	);
	LUT2 #(
		.INIT('h1)
	) name4465 (
		\A[171] ,
		_w5465_,
		_w5467_
	);
	LUT2 #(
		.INIT('h1)
	) name4466 (
		_w5466_,
		_w5467_,
		_w5468_
	);
	LUT2 #(
		.INIT('h8)
	) name4467 (
		\A[172] ,
		\A[173] ,
		_w5469_
	);
	LUT2 #(
		.INIT('h1)
	) name4468 (
		\A[172] ,
		\A[173] ,
		_w5470_
	);
	LUT2 #(
		.INIT('h1)
	) name4469 (
		_w5469_,
		_w5470_,
		_w5471_
	);
	LUT2 #(
		.INIT('h8)
	) name4470 (
		\A[174] ,
		_w5471_,
		_w5472_
	);
	LUT2 #(
		.INIT('h1)
	) name4471 (
		\A[174] ,
		_w5471_,
		_w5473_
	);
	LUT2 #(
		.INIT('h1)
	) name4472 (
		_w5472_,
		_w5473_,
		_w5474_
	);
	LUT2 #(
		.INIT('h8)
	) name4473 (
		_w5468_,
		_w5474_,
		_w5475_
	);
	LUT2 #(
		.INIT('h1)
	) name4474 (
		_w5468_,
		_w5474_,
		_w5476_
	);
	LUT2 #(
		.INIT('h1)
	) name4475 (
		_w5475_,
		_w5476_,
		_w5477_
	);
	LUT2 #(
		.INIT('h8)
	) name4476 (
		\A[163] ,
		\A[164] ,
		_w5478_
	);
	LUT2 #(
		.INIT('h1)
	) name4477 (
		\A[163] ,
		\A[164] ,
		_w5479_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		_w5478_,
		_w5479_,
		_w5480_
	);
	LUT2 #(
		.INIT('h8)
	) name4479 (
		\A[165] ,
		_w5480_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name4480 (
		\A[165] ,
		_w5480_,
		_w5482_
	);
	LUT2 #(
		.INIT('h1)
	) name4481 (
		_w5481_,
		_w5482_,
		_w5483_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		\A[166] ,
		\A[167] ,
		_w5484_
	);
	LUT2 #(
		.INIT('h1)
	) name4483 (
		\A[166] ,
		\A[167] ,
		_w5485_
	);
	LUT2 #(
		.INIT('h1)
	) name4484 (
		_w5484_,
		_w5485_,
		_w5486_
	);
	LUT2 #(
		.INIT('h8)
	) name4485 (
		\A[168] ,
		_w5486_,
		_w5487_
	);
	LUT2 #(
		.INIT('h1)
	) name4486 (
		\A[168] ,
		_w5486_,
		_w5488_
	);
	LUT2 #(
		.INIT('h1)
	) name4487 (
		_w5487_,
		_w5488_,
		_w5489_
	);
	LUT2 #(
		.INIT('h8)
	) name4488 (
		_w5483_,
		_w5489_,
		_w5490_
	);
	LUT2 #(
		.INIT('h1)
	) name4489 (
		_w5483_,
		_w5489_,
		_w5491_
	);
	LUT2 #(
		.INIT('h1)
	) name4490 (
		_w5490_,
		_w5491_,
		_w5492_
	);
	LUT2 #(
		.INIT('h8)
	) name4491 (
		_w5477_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h1)
	) name4492 (
		_w5469_,
		_w5472_,
		_w5494_
	);
	LUT2 #(
		.INIT('h1)
	) name4493 (
		_w5463_,
		_w5466_,
		_w5495_
	);
	LUT2 #(
		.INIT('h1)
	) name4494 (
		_w5494_,
		_w5495_,
		_w5496_
	);
	LUT2 #(
		.INIT('h8)
	) name4495 (
		_w5494_,
		_w5495_,
		_w5497_
	);
	LUT2 #(
		.INIT('h1)
	) name4496 (
		_w5496_,
		_w5497_,
		_w5498_
	);
	LUT2 #(
		.INIT('h8)
	) name4497 (
		_w5493_,
		_w5498_,
		_w5499_
	);
	LUT2 #(
		.INIT('h1)
	) name4498 (
		_w5478_,
		_w5481_,
		_w5500_
	);
	LUT2 #(
		.INIT('h1)
	) name4499 (
		_w5484_,
		_w5487_,
		_w5501_
	);
	LUT2 #(
		.INIT('h4)
	) name4500 (
		_w5490_,
		_w5501_,
		_w5502_
	);
	LUT2 #(
		.INIT('h8)
	) name4501 (
		_w5484_,
		_w5490_,
		_w5503_
	);
	LUT2 #(
		.INIT('h1)
	) name4502 (
		_w5502_,
		_w5503_,
		_w5504_
	);
	LUT2 #(
		.INIT('h2)
	) name4503 (
		_w5500_,
		_w5504_,
		_w5505_
	);
	LUT2 #(
		.INIT('h4)
	) name4504 (
		_w5500_,
		_w5504_,
		_w5506_
	);
	LUT2 #(
		.INIT('h1)
	) name4505 (
		_w5505_,
		_w5506_,
		_w5507_
	);
	LUT2 #(
		.INIT('h1)
	) name4506 (
		_w5499_,
		_w5507_,
		_w5508_
	);
	LUT2 #(
		.INIT('h4)
	) name4507 (
		_w5475_,
		_w5498_,
		_w5509_
	);
	LUT2 #(
		.INIT('h2)
	) name4508 (
		_w5475_,
		_w5498_,
		_w5510_
	);
	LUT2 #(
		.INIT('h1)
	) name4509 (
		_w5493_,
		_w5509_,
		_w5511_
	);
	LUT2 #(
		.INIT('h4)
	) name4510 (
		_w5510_,
		_w5511_,
		_w5512_
	);
	LUT2 #(
		.INIT('h1)
	) name4511 (
		_w5508_,
		_w5512_,
		_w5513_
	);
	LUT2 #(
		.INIT('h1)
	) name4512 (
		_w5475_,
		_w5496_,
		_w5514_
	);
	LUT2 #(
		.INIT('h1)
	) name4513 (
		_w5497_,
		_w5514_,
		_w5515_
	);
	LUT2 #(
		.INIT('h1)
	) name4514 (
		_w5513_,
		_w5515_,
		_w5516_
	);
	LUT2 #(
		.INIT('h8)
	) name4515 (
		_w5513_,
		_w5515_,
		_w5517_
	);
	LUT2 #(
		.INIT('h1)
	) name4516 (
		_w5500_,
		_w5502_,
		_w5518_
	);
	LUT2 #(
		.INIT('h1)
	) name4517 (
		_w5503_,
		_w5518_,
		_w5519_
	);
	LUT2 #(
		.INIT('h4)
	) name4518 (
		_w5517_,
		_w5519_,
		_w5520_
	);
	LUT2 #(
		.INIT('h1)
	) name4519 (
		_w5516_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h1)
	) name4520 (
		_w5516_,
		_w5517_,
		_w5522_
	);
	LUT2 #(
		.INIT('h4)
	) name4521 (
		_w5519_,
		_w5522_,
		_w5523_
	);
	LUT2 #(
		.INIT('h2)
	) name4522 (
		_w5519_,
		_w5522_,
		_w5524_
	);
	LUT2 #(
		.INIT('h1)
	) name4523 (
		_w5523_,
		_w5524_,
		_w5525_
	);
	LUT2 #(
		.INIT('h8)
	) name4524 (
		\A[154] ,
		\A[155] ,
		_w5526_
	);
	LUT2 #(
		.INIT('h8)
	) name4525 (
		\A[151] ,
		\A[152] ,
		_w5527_
	);
	LUT2 #(
		.INIT('h1)
	) name4526 (
		\A[151] ,
		\A[152] ,
		_w5528_
	);
	LUT2 #(
		.INIT('h1)
	) name4527 (
		_w5527_,
		_w5528_,
		_w5529_
	);
	LUT2 #(
		.INIT('h8)
	) name4528 (
		\A[153] ,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h1)
	) name4529 (
		\A[153] ,
		_w5529_,
		_w5531_
	);
	LUT2 #(
		.INIT('h1)
	) name4530 (
		_w5530_,
		_w5531_,
		_w5532_
	);
	LUT2 #(
		.INIT('h1)
	) name4531 (
		\A[154] ,
		\A[155] ,
		_w5533_
	);
	LUT2 #(
		.INIT('h1)
	) name4532 (
		_w5526_,
		_w5533_,
		_w5534_
	);
	LUT2 #(
		.INIT('h8)
	) name4533 (
		\A[156] ,
		_w5534_,
		_w5535_
	);
	LUT2 #(
		.INIT('h1)
	) name4534 (
		\A[156] ,
		_w5534_,
		_w5536_
	);
	LUT2 #(
		.INIT('h1)
	) name4535 (
		_w5535_,
		_w5536_,
		_w5537_
	);
	LUT2 #(
		.INIT('h8)
	) name4536 (
		_w5532_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h8)
	) name4537 (
		_w5526_,
		_w5538_,
		_w5539_
	);
	LUT2 #(
		.INIT('h1)
	) name4538 (
		_w5527_,
		_w5530_,
		_w5540_
	);
	LUT2 #(
		.INIT('h1)
	) name4539 (
		_w5526_,
		_w5535_,
		_w5541_
	);
	LUT2 #(
		.INIT('h4)
	) name4540 (
		_w5538_,
		_w5541_,
		_w5542_
	);
	LUT2 #(
		.INIT('h1)
	) name4541 (
		_w5540_,
		_w5542_,
		_w5543_
	);
	LUT2 #(
		.INIT('h1)
	) name4542 (
		_w5539_,
		_w5543_,
		_w5544_
	);
	LUT2 #(
		.INIT('h8)
	) name4543 (
		\A[157] ,
		\A[158] ,
		_w5545_
	);
	LUT2 #(
		.INIT('h1)
	) name4544 (
		\A[157] ,
		\A[158] ,
		_w5546_
	);
	LUT2 #(
		.INIT('h1)
	) name4545 (
		_w5545_,
		_w5546_,
		_w5547_
	);
	LUT2 #(
		.INIT('h8)
	) name4546 (
		\A[159] ,
		_w5547_,
		_w5548_
	);
	LUT2 #(
		.INIT('h1)
	) name4547 (
		\A[159] ,
		_w5547_,
		_w5549_
	);
	LUT2 #(
		.INIT('h1)
	) name4548 (
		_w5548_,
		_w5549_,
		_w5550_
	);
	LUT2 #(
		.INIT('h8)
	) name4549 (
		\A[160] ,
		\A[161] ,
		_w5551_
	);
	LUT2 #(
		.INIT('h1)
	) name4550 (
		\A[160] ,
		\A[161] ,
		_w5552_
	);
	LUT2 #(
		.INIT('h1)
	) name4551 (
		_w5551_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h8)
	) name4552 (
		\A[162] ,
		_w5553_,
		_w5554_
	);
	LUT2 #(
		.INIT('h1)
	) name4553 (
		\A[162] ,
		_w5553_,
		_w5555_
	);
	LUT2 #(
		.INIT('h1)
	) name4554 (
		_w5554_,
		_w5555_,
		_w5556_
	);
	LUT2 #(
		.INIT('h8)
	) name4555 (
		_w5550_,
		_w5556_,
		_w5557_
	);
	LUT2 #(
		.INIT('h1)
	) name4556 (
		_w5550_,
		_w5556_,
		_w5558_
	);
	LUT2 #(
		.INIT('h1)
	) name4557 (
		_w5557_,
		_w5558_,
		_w5559_
	);
	LUT2 #(
		.INIT('h1)
	) name4558 (
		_w5532_,
		_w5537_,
		_w5560_
	);
	LUT2 #(
		.INIT('h1)
	) name4559 (
		_w5538_,
		_w5560_,
		_w5561_
	);
	LUT2 #(
		.INIT('h8)
	) name4560 (
		_w5559_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h1)
	) name4561 (
		_w5551_,
		_w5554_,
		_w5563_
	);
	LUT2 #(
		.INIT('h1)
	) name4562 (
		_w5545_,
		_w5548_,
		_w5564_
	);
	LUT2 #(
		.INIT('h1)
	) name4563 (
		_w5563_,
		_w5564_,
		_w5565_
	);
	LUT2 #(
		.INIT('h8)
	) name4564 (
		_w5563_,
		_w5564_,
		_w5566_
	);
	LUT2 #(
		.INIT('h1)
	) name4565 (
		_w5565_,
		_w5566_,
		_w5567_
	);
	LUT2 #(
		.INIT('h8)
	) name4566 (
		_w5562_,
		_w5567_,
		_w5568_
	);
	LUT2 #(
		.INIT('h1)
	) name4567 (
		_w5539_,
		_w5542_,
		_w5569_
	);
	LUT2 #(
		.INIT('h2)
	) name4568 (
		_w5540_,
		_w5569_,
		_w5570_
	);
	LUT2 #(
		.INIT('h4)
	) name4569 (
		_w5540_,
		_w5569_,
		_w5571_
	);
	LUT2 #(
		.INIT('h1)
	) name4570 (
		_w5570_,
		_w5571_,
		_w5572_
	);
	LUT2 #(
		.INIT('h1)
	) name4571 (
		_w5568_,
		_w5572_,
		_w5573_
	);
	LUT2 #(
		.INIT('h4)
	) name4572 (
		_w5557_,
		_w5567_,
		_w5574_
	);
	LUT2 #(
		.INIT('h2)
	) name4573 (
		_w5557_,
		_w5567_,
		_w5575_
	);
	LUT2 #(
		.INIT('h1)
	) name4574 (
		_w5562_,
		_w5574_,
		_w5576_
	);
	LUT2 #(
		.INIT('h4)
	) name4575 (
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('h1)
	) name4576 (
		_w5573_,
		_w5577_,
		_w5578_
	);
	LUT2 #(
		.INIT('h1)
	) name4577 (
		_w5557_,
		_w5565_,
		_w5579_
	);
	LUT2 #(
		.INIT('h1)
	) name4578 (
		_w5566_,
		_w5579_,
		_w5580_
	);
	LUT2 #(
		.INIT('h1)
	) name4579 (
		_w5578_,
		_w5580_,
		_w5581_
	);
	LUT2 #(
		.INIT('h8)
	) name4580 (
		_w5578_,
		_w5580_,
		_w5582_
	);
	LUT2 #(
		.INIT('h1)
	) name4581 (
		_w5581_,
		_w5582_,
		_w5583_
	);
	LUT2 #(
		.INIT('h2)
	) name4582 (
		_w5544_,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h4)
	) name4583 (
		_w5544_,
		_w5583_,
		_w5585_
	);
	LUT2 #(
		.INIT('h1)
	) name4584 (
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT2 #(
		.INIT('h8)
	) name4585 (
		_w5525_,
		_w5586_,
		_w5587_
	);
	LUT2 #(
		.INIT('h1)
	) name4586 (
		_w5525_,
		_w5586_,
		_w5588_
	);
	LUT2 #(
		.INIT('h1)
	) name4587 (
		_w5477_,
		_w5492_,
		_w5589_
	);
	LUT2 #(
		.INIT('h1)
	) name4588 (
		_w5493_,
		_w5589_,
		_w5590_
	);
	LUT2 #(
		.INIT('h1)
	) name4589 (
		_w5559_,
		_w5561_,
		_w5591_
	);
	LUT2 #(
		.INIT('h1)
	) name4590 (
		_w5562_,
		_w5591_,
		_w5592_
	);
	LUT2 #(
		.INIT('h8)
	) name4591 (
		_w5590_,
		_w5592_,
		_w5593_
	);
	LUT2 #(
		.INIT('h1)
	) name4592 (
		_w5499_,
		_w5512_,
		_w5594_
	);
	LUT2 #(
		.INIT('h4)
	) name4593 (
		_w5507_,
		_w5594_,
		_w5595_
	);
	LUT2 #(
		.INIT('h2)
	) name4594 (
		_w5507_,
		_w5594_,
		_w5596_
	);
	LUT2 #(
		.INIT('h1)
	) name4595 (
		_w5595_,
		_w5596_,
		_w5597_
	);
	LUT2 #(
		.INIT('h2)
	) name4596 (
		_w5593_,
		_w5597_,
		_w5598_
	);
	LUT2 #(
		.INIT('h4)
	) name4597 (
		_w5593_,
		_w5597_,
		_w5599_
	);
	LUT2 #(
		.INIT('h1)
	) name4598 (
		_w5568_,
		_w5577_,
		_w5600_
	);
	LUT2 #(
		.INIT('h4)
	) name4599 (
		_w5572_,
		_w5600_,
		_w5601_
	);
	LUT2 #(
		.INIT('h2)
	) name4600 (
		_w5572_,
		_w5600_,
		_w5602_
	);
	LUT2 #(
		.INIT('h1)
	) name4601 (
		_w5601_,
		_w5602_,
		_w5603_
	);
	LUT2 #(
		.INIT('h1)
	) name4602 (
		_w5599_,
		_w5603_,
		_w5604_
	);
	LUT2 #(
		.INIT('h1)
	) name4603 (
		_w5598_,
		_w5604_,
		_w5605_
	);
	LUT2 #(
		.INIT('h1)
	) name4604 (
		_w5588_,
		_w5605_,
		_w5606_
	);
	LUT2 #(
		.INIT('h1)
	) name4605 (
		_w5587_,
		_w5606_,
		_w5607_
	);
	LUT2 #(
		.INIT('h4)
	) name4606 (
		_w5521_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('h2)
	) name4607 (
		_w5521_,
		_w5607_,
		_w5609_
	);
	LUT2 #(
		.INIT('h2)
	) name4608 (
		_w5544_,
		_w5582_,
		_w5610_
	);
	LUT2 #(
		.INIT('h1)
	) name4609 (
		_w5581_,
		_w5610_,
		_w5611_
	);
	LUT2 #(
		.INIT('h1)
	) name4610 (
		_w5609_,
		_w5611_,
		_w5612_
	);
	LUT2 #(
		.INIT('h1)
	) name4611 (
		_w5608_,
		_w5612_,
		_w5613_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		_w5462_,
		_w5613_,
		_w5614_
	);
	LUT2 #(
		.INIT('h8)
	) name4613 (
		_w5462_,
		_w5613_,
		_w5615_
	);
	LUT2 #(
		.INIT('h1)
	) name4614 (
		_w5608_,
		_w5609_,
		_w5616_
	);
	LUT2 #(
		.INIT('h4)
	) name4615 (
		_w5611_,
		_w5616_,
		_w5617_
	);
	LUT2 #(
		.INIT('h2)
	) name4616 (
		_w5611_,
		_w5616_,
		_w5618_
	);
	LUT2 #(
		.INIT('h1)
	) name4617 (
		_w5617_,
		_w5618_,
		_w5619_
	);
	LUT2 #(
		.INIT('h1)
	) name4618 (
		_w5457_,
		_w5458_,
		_w5620_
	);
	LUT2 #(
		.INIT('h4)
	) name4619 (
		_w5460_,
		_w5620_,
		_w5621_
	);
	LUT2 #(
		.INIT('h2)
	) name4620 (
		_w5460_,
		_w5620_,
		_w5622_
	);
	LUT2 #(
		.INIT('h1)
	) name4621 (
		_w5621_,
		_w5622_,
		_w5623_
	);
	LUT2 #(
		.INIT('h8)
	) name4622 (
		_w5619_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h1)
	) name4623 (
		_w5619_,
		_w5623_,
		_w5625_
	);
	LUT2 #(
		.INIT('h1)
	) name4624 (
		_w5436_,
		_w5437_,
		_w5626_
	);
	LUT2 #(
		.INIT('h4)
	) name4625 (
		_w5454_,
		_w5626_,
		_w5627_
	);
	LUT2 #(
		.INIT('h2)
	) name4626 (
		_w5454_,
		_w5626_,
		_w5628_
	);
	LUT2 #(
		.INIT('h1)
	) name4627 (
		_w5627_,
		_w5628_,
		_w5629_
	);
	LUT2 #(
		.INIT('h1)
	) name4628 (
		_w5587_,
		_w5588_,
		_w5630_
	);
	LUT2 #(
		.INIT('h4)
	) name4629 (
		_w5605_,
		_w5630_,
		_w5631_
	);
	LUT2 #(
		.INIT('h2)
	) name4630 (
		_w5605_,
		_w5630_,
		_w5632_
	);
	LUT2 #(
		.INIT('h1)
	) name4631 (
		_w5631_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h1)
	) name4632 (
		_w5629_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h8)
	) name4633 (
		_w5629_,
		_w5633_,
		_w5635_
	);
	LUT2 #(
		.INIT('h1)
	) name4634 (
		_w5590_,
		_w5592_,
		_w5636_
	);
	LUT2 #(
		.INIT('h1)
	) name4635 (
		_w5593_,
		_w5636_,
		_w5637_
	);
	LUT2 #(
		.INIT('h1)
	) name4636 (
		_w5439_,
		_w5441_,
		_w5638_
	);
	LUT2 #(
		.INIT('h1)
	) name4637 (
		_w5442_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('h8)
	) name4638 (
		_w5637_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h1)
	) name4639 (
		_w5598_,
		_w5599_,
		_w5641_
	);
	LUT2 #(
		.INIT('h4)
	) name4640 (
		_w5603_,
		_w5641_,
		_w5642_
	);
	LUT2 #(
		.INIT('h2)
	) name4641 (
		_w5603_,
		_w5641_,
		_w5643_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w5642_,
		_w5643_,
		_w5644_
	);
	LUT2 #(
		.INIT('h8)
	) name4643 (
		_w5640_,
		_w5644_,
		_w5645_
	);
	LUT2 #(
		.INIT('h1)
	) name4644 (
		_w5640_,
		_w5644_,
		_w5646_
	);
	LUT2 #(
		.INIT('h1)
	) name4645 (
		_w5447_,
		_w5448_,
		_w5647_
	);
	LUT2 #(
		.INIT('h4)
	) name4646 (
		_w5452_,
		_w5647_,
		_w5648_
	);
	LUT2 #(
		.INIT('h2)
	) name4647 (
		_w5452_,
		_w5647_,
		_w5649_
	);
	LUT2 #(
		.INIT('h1)
	) name4648 (
		_w5648_,
		_w5649_,
		_w5650_
	);
	LUT2 #(
		.INIT('h4)
	) name4649 (
		_w5646_,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h1)
	) name4650 (
		_w5645_,
		_w5651_,
		_w5652_
	);
	LUT2 #(
		.INIT('h4)
	) name4651 (
		_w5635_,
		_w5652_,
		_w5653_
	);
	LUT2 #(
		.INIT('h1)
	) name4652 (
		_w5634_,
		_w5653_,
		_w5654_
	);
	LUT2 #(
		.INIT('h1)
	) name4653 (
		_w5625_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h1)
	) name4654 (
		_w5624_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h1)
	) name4655 (
		_w5615_,
		_w5656_,
		_w5657_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w5614_,
		_w5657_,
		_w5658_
	);
	LUT2 #(
		.INIT('h8)
	) name4657 (
		\A[97] ,
		\A[98] ,
		_w5659_
	);
	LUT2 #(
		.INIT('h1)
	) name4658 (
		\A[97] ,
		\A[98] ,
		_w5660_
	);
	LUT2 #(
		.INIT('h1)
	) name4659 (
		_w5659_,
		_w5660_,
		_w5661_
	);
	LUT2 #(
		.INIT('h8)
	) name4660 (
		\A[99] ,
		_w5661_,
		_w5662_
	);
	LUT2 #(
		.INIT('h1)
	) name4661 (
		\A[99] ,
		_w5661_,
		_w5663_
	);
	LUT2 #(
		.INIT('h1)
	) name4662 (
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT2 #(
		.INIT('h8)
	) name4663 (
		\A[100] ,
		\A[101] ,
		_w5665_
	);
	LUT2 #(
		.INIT('h1)
	) name4664 (
		\A[100] ,
		\A[101] ,
		_w5666_
	);
	LUT2 #(
		.INIT('h1)
	) name4665 (
		_w5665_,
		_w5666_,
		_w5667_
	);
	LUT2 #(
		.INIT('h8)
	) name4666 (
		\A[102] ,
		_w5667_,
		_w5668_
	);
	LUT2 #(
		.INIT('h1)
	) name4667 (
		\A[102] ,
		_w5667_,
		_w5669_
	);
	LUT2 #(
		.INIT('h1)
	) name4668 (
		_w5668_,
		_w5669_,
		_w5670_
	);
	LUT2 #(
		.INIT('h8)
	) name4669 (
		_w5664_,
		_w5670_,
		_w5671_
	);
	LUT2 #(
		.INIT('h1)
	) name4670 (
		_w5664_,
		_w5670_,
		_w5672_
	);
	LUT2 #(
		.INIT('h1)
	) name4671 (
		_w5671_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h8)
	) name4672 (
		\A[91] ,
		\A[92] ,
		_w5674_
	);
	LUT2 #(
		.INIT('h1)
	) name4673 (
		\A[91] ,
		\A[92] ,
		_w5675_
	);
	LUT2 #(
		.INIT('h1)
	) name4674 (
		_w5674_,
		_w5675_,
		_w5676_
	);
	LUT2 #(
		.INIT('h8)
	) name4675 (
		\A[93] ,
		_w5676_,
		_w5677_
	);
	LUT2 #(
		.INIT('h1)
	) name4676 (
		\A[93] ,
		_w5676_,
		_w5678_
	);
	LUT2 #(
		.INIT('h1)
	) name4677 (
		_w5677_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h8)
	) name4678 (
		\A[94] ,
		\A[95] ,
		_w5680_
	);
	LUT2 #(
		.INIT('h1)
	) name4679 (
		\A[94] ,
		\A[95] ,
		_w5681_
	);
	LUT2 #(
		.INIT('h1)
	) name4680 (
		_w5680_,
		_w5681_,
		_w5682_
	);
	LUT2 #(
		.INIT('h8)
	) name4681 (
		\A[96] ,
		_w5682_,
		_w5683_
	);
	LUT2 #(
		.INIT('h1)
	) name4682 (
		\A[96] ,
		_w5682_,
		_w5684_
	);
	LUT2 #(
		.INIT('h1)
	) name4683 (
		_w5683_,
		_w5684_,
		_w5685_
	);
	LUT2 #(
		.INIT('h8)
	) name4684 (
		_w5679_,
		_w5685_,
		_w5686_
	);
	LUT2 #(
		.INIT('h1)
	) name4685 (
		_w5679_,
		_w5685_,
		_w5687_
	);
	LUT2 #(
		.INIT('h1)
	) name4686 (
		_w5686_,
		_w5687_,
		_w5688_
	);
	LUT2 #(
		.INIT('h8)
	) name4687 (
		_w5673_,
		_w5688_,
		_w5689_
	);
	LUT2 #(
		.INIT('h1)
	) name4688 (
		_w5665_,
		_w5668_,
		_w5690_
	);
	LUT2 #(
		.INIT('h1)
	) name4689 (
		_w5659_,
		_w5662_,
		_w5691_
	);
	LUT2 #(
		.INIT('h1)
	) name4690 (
		_w5690_,
		_w5691_,
		_w5692_
	);
	LUT2 #(
		.INIT('h8)
	) name4691 (
		_w5690_,
		_w5691_,
		_w5693_
	);
	LUT2 #(
		.INIT('h1)
	) name4692 (
		_w5692_,
		_w5693_,
		_w5694_
	);
	LUT2 #(
		.INIT('h8)
	) name4693 (
		_w5689_,
		_w5694_,
		_w5695_
	);
	LUT2 #(
		.INIT('h1)
	) name4694 (
		_w5674_,
		_w5677_,
		_w5696_
	);
	LUT2 #(
		.INIT('h1)
	) name4695 (
		_w5680_,
		_w5683_,
		_w5697_
	);
	LUT2 #(
		.INIT('h4)
	) name4696 (
		_w5686_,
		_w5697_,
		_w5698_
	);
	LUT2 #(
		.INIT('h8)
	) name4697 (
		_w5680_,
		_w5686_,
		_w5699_
	);
	LUT2 #(
		.INIT('h1)
	) name4698 (
		_w5698_,
		_w5699_,
		_w5700_
	);
	LUT2 #(
		.INIT('h2)
	) name4699 (
		_w5696_,
		_w5700_,
		_w5701_
	);
	LUT2 #(
		.INIT('h4)
	) name4700 (
		_w5696_,
		_w5700_,
		_w5702_
	);
	LUT2 #(
		.INIT('h1)
	) name4701 (
		_w5701_,
		_w5702_,
		_w5703_
	);
	LUT2 #(
		.INIT('h1)
	) name4702 (
		_w5695_,
		_w5703_,
		_w5704_
	);
	LUT2 #(
		.INIT('h4)
	) name4703 (
		_w5671_,
		_w5694_,
		_w5705_
	);
	LUT2 #(
		.INIT('h2)
	) name4704 (
		_w5671_,
		_w5694_,
		_w5706_
	);
	LUT2 #(
		.INIT('h1)
	) name4705 (
		_w5689_,
		_w5705_,
		_w5707_
	);
	LUT2 #(
		.INIT('h4)
	) name4706 (
		_w5706_,
		_w5707_,
		_w5708_
	);
	LUT2 #(
		.INIT('h1)
	) name4707 (
		_w5704_,
		_w5708_,
		_w5709_
	);
	LUT2 #(
		.INIT('h1)
	) name4708 (
		_w5671_,
		_w5692_,
		_w5710_
	);
	LUT2 #(
		.INIT('h1)
	) name4709 (
		_w5693_,
		_w5710_,
		_w5711_
	);
	LUT2 #(
		.INIT('h1)
	) name4710 (
		_w5709_,
		_w5711_,
		_w5712_
	);
	LUT2 #(
		.INIT('h8)
	) name4711 (
		_w5709_,
		_w5711_,
		_w5713_
	);
	LUT2 #(
		.INIT('h1)
	) name4712 (
		_w5696_,
		_w5698_,
		_w5714_
	);
	LUT2 #(
		.INIT('h1)
	) name4713 (
		_w5699_,
		_w5714_,
		_w5715_
	);
	LUT2 #(
		.INIT('h4)
	) name4714 (
		_w5713_,
		_w5715_,
		_w5716_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w5712_,
		_w5716_,
		_w5717_
	);
	LUT2 #(
		.INIT('h1)
	) name4716 (
		_w5712_,
		_w5713_,
		_w5718_
	);
	LUT2 #(
		.INIT('h4)
	) name4717 (
		_w5715_,
		_w5718_,
		_w5719_
	);
	LUT2 #(
		.INIT('h2)
	) name4718 (
		_w5715_,
		_w5718_,
		_w5720_
	);
	LUT2 #(
		.INIT('h1)
	) name4719 (
		_w5719_,
		_w5720_,
		_w5721_
	);
	LUT2 #(
		.INIT('h8)
	) name4720 (
		\A[82] ,
		\A[83] ,
		_w5722_
	);
	LUT2 #(
		.INIT('h8)
	) name4721 (
		\A[79] ,
		\A[80] ,
		_w5723_
	);
	LUT2 #(
		.INIT('h1)
	) name4722 (
		\A[79] ,
		\A[80] ,
		_w5724_
	);
	LUT2 #(
		.INIT('h1)
	) name4723 (
		_w5723_,
		_w5724_,
		_w5725_
	);
	LUT2 #(
		.INIT('h8)
	) name4724 (
		\A[81] ,
		_w5725_,
		_w5726_
	);
	LUT2 #(
		.INIT('h1)
	) name4725 (
		\A[81] ,
		_w5725_,
		_w5727_
	);
	LUT2 #(
		.INIT('h1)
	) name4726 (
		_w5726_,
		_w5727_,
		_w5728_
	);
	LUT2 #(
		.INIT('h1)
	) name4727 (
		\A[82] ,
		\A[83] ,
		_w5729_
	);
	LUT2 #(
		.INIT('h1)
	) name4728 (
		_w5722_,
		_w5729_,
		_w5730_
	);
	LUT2 #(
		.INIT('h8)
	) name4729 (
		\A[84] ,
		_w5730_,
		_w5731_
	);
	LUT2 #(
		.INIT('h1)
	) name4730 (
		\A[84] ,
		_w5730_,
		_w5732_
	);
	LUT2 #(
		.INIT('h1)
	) name4731 (
		_w5731_,
		_w5732_,
		_w5733_
	);
	LUT2 #(
		.INIT('h8)
	) name4732 (
		_w5728_,
		_w5733_,
		_w5734_
	);
	LUT2 #(
		.INIT('h8)
	) name4733 (
		_w5722_,
		_w5734_,
		_w5735_
	);
	LUT2 #(
		.INIT('h1)
	) name4734 (
		_w5723_,
		_w5726_,
		_w5736_
	);
	LUT2 #(
		.INIT('h1)
	) name4735 (
		_w5722_,
		_w5731_,
		_w5737_
	);
	LUT2 #(
		.INIT('h4)
	) name4736 (
		_w5734_,
		_w5737_,
		_w5738_
	);
	LUT2 #(
		.INIT('h1)
	) name4737 (
		_w5736_,
		_w5738_,
		_w5739_
	);
	LUT2 #(
		.INIT('h1)
	) name4738 (
		_w5735_,
		_w5739_,
		_w5740_
	);
	LUT2 #(
		.INIT('h8)
	) name4739 (
		\A[85] ,
		\A[86] ,
		_w5741_
	);
	LUT2 #(
		.INIT('h1)
	) name4740 (
		\A[85] ,
		\A[86] ,
		_w5742_
	);
	LUT2 #(
		.INIT('h1)
	) name4741 (
		_w5741_,
		_w5742_,
		_w5743_
	);
	LUT2 #(
		.INIT('h8)
	) name4742 (
		\A[87] ,
		_w5743_,
		_w5744_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		\A[87] ,
		_w5743_,
		_w5745_
	);
	LUT2 #(
		.INIT('h1)
	) name4744 (
		_w5744_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h8)
	) name4745 (
		\A[88] ,
		\A[89] ,
		_w5747_
	);
	LUT2 #(
		.INIT('h1)
	) name4746 (
		\A[88] ,
		\A[89] ,
		_w5748_
	);
	LUT2 #(
		.INIT('h1)
	) name4747 (
		_w5747_,
		_w5748_,
		_w5749_
	);
	LUT2 #(
		.INIT('h8)
	) name4748 (
		\A[90] ,
		_w5749_,
		_w5750_
	);
	LUT2 #(
		.INIT('h1)
	) name4749 (
		\A[90] ,
		_w5749_,
		_w5751_
	);
	LUT2 #(
		.INIT('h1)
	) name4750 (
		_w5750_,
		_w5751_,
		_w5752_
	);
	LUT2 #(
		.INIT('h8)
	) name4751 (
		_w5746_,
		_w5752_,
		_w5753_
	);
	LUT2 #(
		.INIT('h1)
	) name4752 (
		_w5746_,
		_w5752_,
		_w5754_
	);
	LUT2 #(
		.INIT('h1)
	) name4753 (
		_w5753_,
		_w5754_,
		_w5755_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w5728_,
		_w5733_,
		_w5756_
	);
	LUT2 #(
		.INIT('h1)
	) name4755 (
		_w5734_,
		_w5756_,
		_w5757_
	);
	LUT2 #(
		.INIT('h8)
	) name4756 (
		_w5755_,
		_w5757_,
		_w5758_
	);
	LUT2 #(
		.INIT('h1)
	) name4757 (
		_w5747_,
		_w5750_,
		_w5759_
	);
	LUT2 #(
		.INIT('h1)
	) name4758 (
		_w5741_,
		_w5744_,
		_w5760_
	);
	LUT2 #(
		.INIT('h1)
	) name4759 (
		_w5759_,
		_w5760_,
		_w5761_
	);
	LUT2 #(
		.INIT('h8)
	) name4760 (
		_w5759_,
		_w5760_,
		_w5762_
	);
	LUT2 #(
		.INIT('h1)
	) name4761 (
		_w5761_,
		_w5762_,
		_w5763_
	);
	LUT2 #(
		.INIT('h8)
	) name4762 (
		_w5758_,
		_w5763_,
		_w5764_
	);
	LUT2 #(
		.INIT('h1)
	) name4763 (
		_w5735_,
		_w5738_,
		_w5765_
	);
	LUT2 #(
		.INIT('h2)
	) name4764 (
		_w5736_,
		_w5765_,
		_w5766_
	);
	LUT2 #(
		.INIT('h4)
	) name4765 (
		_w5736_,
		_w5765_,
		_w5767_
	);
	LUT2 #(
		.INIT('h1)
	) name4766 (
		_w5766_,
		_w5767_,
		_w5768_
	);
	LUT2 #(
		.INIT('h1)
	) name4767 (
		_w5764_,
		_w5768_,
		_w5769_
	);
	LUT2 #(
		.INIT('h4)
	) name4768 (
		_w5753_,
		_w5763_,
		_w5770_
	);
	LUT2 #(
		.INIT('h2)
	) name4769 (
		_w5753_,
		_w5763_,
		_w5771_
	);
	LUT2 #(
		.INIT('h1)
	) name4770 (
		_w5758_,
		_w5770_,
		_w5772_
	);
	LUT2 #(
		.INIT('h4)
	) name4771 (
		_w5771_,
		_w5772_,
		_w5773_
	);
	LUT2 #(
		.INIT('h1)
	) name4772 (
		_w5769_,
		_w5773_,
		_w5774_
	);
	LUT2 #(
		.INIT('h1)
	) name4773 (
		_w5753_,
		_w5761_,
		_w5775_
	);
	LUT2 #(
		.INIT('h1)
	) name4774 (
		_w5762_,
		_w5775_,
		_w5776_
	);
	LUT2 #(
		.INIT('h1)
	) name4775 (
		_w5774_,
		_w5776_,
		_w5777_
	);
	LUT2 #(
		.INIT('h8)
	) name4776 (
		_w5774_,
		_w5776_,
		_w5778_
	);
	LUT2 #(
		.INIT('h1)
	) name4777 (
		_w5777_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h2)
	) name4778 (
		_w5740_,
		_w5779_,
		_w5780_
	);
	LUT2 #(
		.INIT('h4)
	) name4779 (
		_w5740_,
		_w5779_,
		_w5781_
	);
	LUT2 #(
		.INIT('h1)
	) name4780 (
		_w5780_,
		_w5781_,
		_w5782_
	);
	LUT2 #(
		.INIT('h8)
	) name4781 (
		_w5721_,
		_w5782_,
		_w5783_
	);
	LUT2 #(
		.INIT('h1)
	) name4782 (
		_w5721_,
		_w5782_,
		_w5784_
	);
	LUT2 #(
		.INIT('h1)
	) name4783 (
		_w5673_,
		_w5688_,
		_w5785_
	);
	LUT2 #(
		.INIT('h1)
	) name4784 (
		_w5689_,
		_w5785_,
		_w5786_
	);
	LUT2 #(
		.INIT('h1)
	) name4785 (
		_w5755_,
		_w5757_,
		_w5787_
	);
	LUT2 #(
		.INIT('h1)
	) name4786 (
		_w5758_,
		_w5787_,
		_w5788_
	);
	LUT2 #(
		.INIT('h8)
	) name4787 (
		_w5786_,
		_w5788_,
		_w5789_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		_w5695_,
		_w5708_,
		_w5790_
	);
	LUT2 #(
		.INIT('h4)
	) name4789 (
		_w5703_,
		_w5790_,
		_w5791_
	);
	LUT2 #(
		.INIT('h2)
	) name4790 (
		_w5703_,
		_w5790_,
		_w5792_
	);
	LUT2 #(
		.INIT('h1)
	) name4791 (
		_w5791_,
		_w5792_,
		_w5793_
	);
	LUT2 #(
		.INIT('h2)
	) name4792 (
		_w5789_,
		_w5793_,
		_w5794_
	);
	LUT2 #(
		.INIT('h4)
	) name4793 (
		_w5789_,
		_w5793_,
		_w5795_
	);
	LUT2 #(
		.INIT('h1)
	) name4794 (
		_w5764_,
		_w5773_,
		_w5796_
	);
	LUT2 #(
		.INIT('h4)
	) name4795 (
		_w5768_,
		_w5796_,
		_w5797_
	);
	LUT2 #(
		.INIT('h2)
	) name4796 (
		_w5768_,
		_w5796_,
		_w5798_
	);
	LUT2 #(
		.INIT('h1)
	) name4797 (
		_w5797_,
		_w5798_,
		_w5799_
	);
	LUT2 #(
		.INIT('h1)
	) name4798 (
		_w5795_,
		_w5799_,
		_w5800_
	);
	LUT2 #(
		.INIT('h1)
	) name4799 (
		_w5794_,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h1)
	) name4800 (
		_w5784_,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h1)
	) name4801 (
		_w5783_,
		_w5802_,
		_w5803_
	);
	LUT2 #(
		.INIT('h4)
	) name4802 (
		_w5717_,
		_w5803_,
		_w5804_
	);
	LUT2 #(
		.INIT('h2)
	) name4803 (
		_w5717_,
		_w5803_,
		_w5805_
	);
	LUT2 #(
		.INIT('h2)
	) name4804 (
		_w5740_,
		_w5778_,
		_w5806_
	);
	LUT2 #(
		.INIT('h1)
	) name4805 (
		_w5777_,
		_w5806_,
		_w5807_
	);
	LUT2 #(
		.INIT('h1)
	) name4806 (
		_w5805_,
		_w5807_,
		_w5808_
	);
	LUT2 #(
		.INIT('h1)
	) name4807 (
		_w5804_,
		_w5808_,
		_w5809_
	);
	LUT2 #(
		.INIT('h8)
	) name4808 (
		\A[121] ,
		\A[122] ,
		_w5810_
	);
	LUT2 #(
		.INIT('h1)
	) name4809 (
		\A[121] ,
		\A[122] ,
		_w5811_
	);
	LUT2 #(
		.INIT('h1)
	) name4810 (
		_w5810_,
		_w5811_,
		_w5812_
	);
	LUT2 #(
		.INIT('h8)
	) name4811 (
		\A[123] ,
		_w5812_,
		_w5813_
	);
	LUT2 #(
		.INIT('h1)
	) name4812 (
		\A[123] ,
		_w5812_,
		_w5814_
	);
	LUT2 #(
		.INIT('h1)
	) name4813 (
		_w5813_,
		_w5814_,
		_w5815_
	);
	LUT2 #(
		.INIT('h8)
	) name4814 (
		\A[124] ,
		\A[125] ,
		_w5816_
	);
	LUT2 #(
		.INIT('h1)
	) name4815 (
		\A[124] ,
		\A[125] ,
		_w5817_
	);
	LUT2 #(
		.INIT('h1)
	) name4816 (
		_w5816_,
		_w5817_,
		_w5818_
	);
	LUT2 #(
		.INIT('h8)
	) name4817 (
		\A[126] ,
		_w5818_,
		_w5819_
	);
	LUT2 #(
		.INIT('h1)
	) name4818 (
		\A[126] ,
		_w5818_,
		_w5820_
	);
	LUT2 #(
		.INIT('h1)
	) name4819 (
		_w5819_,
		_w5820_,
		_w5821_
	);
	LUT2 #(
		.INIT('h8)
	) name4820 (
		_w5815_,
		_w5821_,
		_w5822_
	);
	LUT2 #(
		.INIT('h1)
	) name4821 (
		_w5815_,
		_w5821_,
		_w5823_
	);
	LUT2 #(
		.INIT('h1)
	) name4822 (
		_w5822_,
		_w5823_,
		_w5824_
	);
	LUT2 #(
		.INIT('h8)
	) name4823 (
		\A[115] ,
		\A[116] ,
		_w5825_
	);
	LUT2 #(
		.INIT('h1)
	) name4824 (
		\A[115] ,
		\A[116] ,
		_w5826_
	);
	LUT2 #(
		.INIT('h1)
	) name4825 (
		_w5825_,
		_w5826_,
		_w5827_
	);
	LUT2 #(
		.INIT('h8)
	) name4826 (
		\A[117] ,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h1)
	) name4827 (
		\A[117] ,
		_w5827_,
		_w5829_
	);
	LUT2 #(
		.INIT('h1)
	) name4828 (
		_w5828_,
		_w5829_,
		_w5830_
	);
	LUT2 #(
		.INIT('h8)
	) name4829 (
		\A[118] ,
		\A[119] ,
		_w5831_
	);
	LUT2 #(
		.INIT('h1)
	) name4830 (
		\A[118] ,
		\A[119] ,
		_w5832_
	);
	LUT2 #(
		.INIT('h1)
	) name4831 (
		_w5831_,
		_w5832_,
		_w5833_
	);
	LUT2 #(
		.INIT('h8)
	) name4832 (
		\A[120] ,
		_w5833_,
		_w5834_
	);
	LUT2 #(
		.INIT('h1)
	) name4833 (
		\A[120] ,
		_w5833_,
		_w5835_
	);
	LUT2 #(
		.INIT('h1)
	) name4834 (
		_w5834_,
		_w5835_,
		_w5836_
	);
	LUT2 #(
		.INIT('h8)
	) name4835 (
		_w5830_,
		_w5836_,
		_w5837_
	);
	LUT2 #(
		.INIT('h1)
	) name4836 (
		_w5830_,
		_w5836_,
		_w5838_
	);
	LUT2 #(
		.INIT('h1)
	) name4837 (
		_w5837_,
		_w5838_,
		_w5839_
	);
	LUT2 #(
		.INIT('h8)
	) name4838 (
		_w5824_,
		_w5839_,
		_w5840_
	);
	LUT2 #(
		.INIT('h1)
	) name4839 (
		_w5816_,
		_w5819_,
		_w5841_
	);
	LUT2 #(
		.INIT('h1)
	) name4840 (
		_w5810_,
		_w5813_,
		_w5842_
	);
	LUT2 #(
		.INIT('h1)
	) name4841 (
		_w5841_,
		_w5842_,
		_w5843_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		_w5841_,
		_w5842_,
		_w5844_
	);
	LUT2 #(
		.INIT('h1)
	) name4843 (
		_w5843_,
		_w5844_,
		_w5845_
	);
	LUT2 #(
		.INIT('h8)
	) name4844 (
		_w5840_,
		_w5845_,
		_w5846_
	);
	LUT2 #(
		.INIT('h1)
	) name4845 (
		_w5825_,
		_w5828_,
		_w5847_
	);
	LUT2 #(
		.INIT('h1)
	) name4846 (
		_w5831_,
		_w5834_,
		_w5848_
	);
	LUT2 #(
		.INIT('h4)
	) name4847 (
		_w5837_,
		_w5848_,
		_w5849_
	);
	LUT2 #(
		.INIT('h8)
	) name4848 (
		_w5831_,
		_w5837_,
		_w5850_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w5849_,
		_w5850_,
		_w5851_
	);
	LUT2 #(
		.INIT('h2)
	) name4850 (
		_w5847_,
		_w5851_,
		_w5852_
	);
	LUT2 #(
		.INIT('h4)
	) name4851 (
		_w5847_,
		_w5851_,
		_w5853_
	);
	LUT2 #(
		.INIT('h1)
	) name4852 (
		_w5852_,
		_w5853_,
		_w5854_
	);
	LUT2 #(
		.INIT('h1)
	) name4853 (
		_w5846_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h4)
	) name4854 (
		_w5822_,
		_w5845_,
		_w5856_
	);
	LUT2 #(
		.INIT('h2)
	) name4855 (
		_w5822_,
		_w5845_,
		_w5857_
	);
	LUT2 #(
		.INIT('h1)
	) name4856 (
		_w5840_,
		_w5856_,
		_w5858_
	);
	LUT2 #(
		.INIT('h4)
	) name4857 (
		_w5857_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('h1)
	) name4858 (
		_w5855_,
		_w5859_,
		_w5860_
	);
	LUT2 #(
		.INIT('h1)
	) name4859 (
		_w5822_,
		_w5843_,
		_w5861_
	);
	LUT2 #(
		.INIT('h1)
	) name4860 (
		_w5844_,
		_w5861_,
		_w5862_
	);
	LUT2 #(
		.INIT('h1)
	) name4861 (
		_w5860_,
		_w5862_,
		_w5863_
	);
	LUT2 #(
		.INIT('h8)
	) name4862 (
		_w5860_,
		_w5862_,
		_w5864_
	);
	LUT2 #(
		.INIT('h1)
	) name4863 (
		_w5847_,
		_w5849_,
		_w5865_
	);
	LUT2 #(
		.INIT('h1)
	) name4864 (
		_w5850_,
		_w5865_,
		_w5866_
	);
	LUT2 #(
		.INIT('h4)
	) name4865 (
		_w5864_,
		_w5866_,
		_w5867_
	);
	LUT2 #(
		.INIT('h1)
	) name4866 (
		_w5863_,
		_w5867_,
		_w5868_
	);
	LUT2 #(
		.INIT('h1)
	) name4867 (
		_w5863_,
		_w5864_,
		_w5869_
	);
	LUT2 #(
		.INIT('h4)
	) name4868 (
		_w5866_,
		_w5869_,
		_w5870_
	);
	LUT2 #(
		.INIT('h2)
	) name4869 (
		_w5866_,
		_w5869_,
		_w5871_
	);
	LUT2 #(
		.INIT('h1)
	) name4870 (
		_w5870_,
		_w5871_,
		_w5872_
	);
	LUT2 #(
		.INIT('h8)
	) name4871 (
		\A[106] ,
		\A[107] ,
		_w5873_
	);
	LUT2 #(
		.INIT('h8)
	) name4872 (
		\A[103] ,
		\A[104] ,
		_w5874_
	);
	LUT2 #(
		.INIT('h1)
	) name4873 (
		\A[103] ,
		\A[104] ,
		_w5875_
	);
	LUT2 #(
		.INIT('h1)
	) name4874 (
		_w5874_,
		_w5875_,
		_w5876_
	);
	LUT2 #(
		.INIT('h8)
	) name4875 (
		\A[105] ,
		_w5876_,
		_w5877_
	);
	LUT2 #(
		.INIT('h1)
	) name4876 (
		\A[105] ,
		_w5876_,
		_w5878_
	);
	LUT2 #(
		.INIT('h1)
	) name4877 (
		_w5877_,
		_w5878_,
		_w5879_
	);
	LUT2 #(
		.INIT('h1)
	) name4878 (
		\A[106] ,
		\A[107] ,
		_w5880_
	);
	LUT2 #(
		.INIT('h1)
	) name4879 (
		_w5873_,
		_w5880_,
		_w5881_
	);
	LUT2 #(
		.INIT('h8)
	) name4880 (
		\A[108] ,
		_w5881_,
		_w5882_
	);
	LUT2 #(
		.INIT('h1)
	) name4881 (
		\A[108] ,
		_w5881_,
		_w5883_
	);
	LUT2 #(
		.INIT('h1)
	) name4882 (
		_w5882_,
		_w5883_,
		_w5884_
	);
	LUT2 #(
		.INIT('h8)
	) name4883 (
		_w5879_,
		_w5884_,
		_w5885_
	);
	LUT2 #(
		.INIT('h8)
	) name4884 (
		_w5873_,
		_w5885_,
		_w5886_
	);
	LUT2 #(
		.INIT('h1)
	) name4885 (
		_w5874_,
		_w5877_,
		_w5887_
	);
	LUT2 #(
		.INIT('h1)
	) name4886 (
		_w5873_,
		_w5882_,
		_w5888_
	);
	LUT2 #(
		.INIT('h4)
	) name4887 (
		_w5885_,
		_w5888_,
		_w5889_
	);
	LUT2 #(
		.INIT('h1)
	) name4888 (
		_w5887_,
		_w5889_,
		_w5890_
	);
	LUT2 #(
		.INIT('h1)
	) name4889 (
		_w5886_,
		_w5890_,
		_w5891_
	);
	LUT2 #(
		.INIT('h8)
	) name4890 (
		\A[109] ,
		\A[110] ,
		_w5892_
	);
	LUT2 #(
		.INIT('h1)
	) name4891 (
		\A[109] ,
		\A[110] ,
		_w5893_
	);
	LUT2 #(
		.INIT('h1)
	) name4892 (
		_w5892_,
		_w5893_,
		_w5894_
	);
	LUT2 #(
		.INIT('h8)
	) name4893 (
		\A[111] ,
		_w5894_,
		_w5895_
	);
	LUT2 #(
		.INIT('h1)
	) name4894 (
		\A[111] ,
		_w5894_,
		_w5896_
	);
	LUT2 #(
		.INIT('h1)
	) name4895 (
		_w5895_,
		_w5896_,
		_w5897_
	);
	LUT2 #(
		.INIT('h8)
	) name4896 (
		\A[112] ,
		\A[113] ,
		_w5898_
	);
	LUT2 #(
		.INIT('h1)
	) name4897 (
		\A[112] ,
		\A[113] ,
		_w5899_
	);
	LUT2 #(
		.INIT('h1)
	) name4898 (
		_w5898_,
		_w5899_,
		_w5900_
	);
	LUT2 #(
		.INIT('h8)
	) name4899 (
		\A[114] ,
		_w5900_,
		_w5901_
	);
	LUT2 #(
		.INIT('h1)
	) name4900 (
		\A[114] ,
		_w5900_,
		_w5902_
	);
	LUT2 #(
		.INIT('h1)
	) name4901 (
		_w5901_,
		_w5902_,
		_w5903_
	);
	LUT2 #(
		.INIT('h8)
	) name4902 (
		_w5897_,
		_w5903_,
		_w5904_
	);
	LUT2 #(
		.INIT('h1)
	) name4903 (
		_w5897_,
		_w5903_,
		_w5905_
	);
	LUT2 #(
		.INIT('h1)
	) name4904 (
		_w5904_,
		_w5905_,
		_w5906_
	);
	LUT2 #(
		.INIT('h1)
	) name4905 (
		_w5879_,
		_w5884_,
		_w5907_
	);
	LUT2 #(
		.INIT('h1)
	) name4906 (
		_w5885_,
		_w5907_,
		_w5908_
	);
	LUT2 #(
		.INIT('h8)
	) name4907 (
		_w5906_,
		_w5908_,
		_w5909_
	);
	LUT2 #(
		.INIT('h1)
	) name4908 (
		_w5898_,
		_w5901_,
		_w5910_
	);
	LUT2 #(
		.INIT('h1)
	) name4909 (
		_w5892_,
		_w5895_,
		_w5911_
	);
	LUT2 #(
		.INIT('h1)
	) name4910 (
		_w5910_,
		_w5911_,
		_w5912_
	);
	LUT2 #(
		.INIT('h8)
	) name4911 (
		_w5910_,
		_w5911_,
		_w5913_
	);
	LUT2 #(
		.INIT('h1)
	) name4912 (
		_w5912_,
		_w5913_,
		_w5914_
	);
	LUT2 #(
		.INIT('h8)
	) name4913 (
		_w5909_,
		_w5914_,
		_w5915_
	);
	LUT2 #(
		.INIT('h1)
	) name4914 (
		_w5886_,
		_w5889_,
		_w5916_
	);
	LUT2 #(
		.INIT('h2)
	) name4915 (
		_w5887_,
		_w5916_,
		_w5917_
	);
	LUT2 #(
		.INIT('h4)
	) name4916 (
		_w5887_,
		_w5916_,
		_w5918_
	);
	LUT2 #(
		.INIT('h1)
	) name4917 (
		_w5917_,
		_w5918_,
		_w5919_
	);
	LUT2 #(
		.INIT('h1)
	) name4918 (
		_w5915_,
		_w5919_,
		_w5920_
	);
	LUT2 #(
		.INIT('h4)
	) name4919 (
		_w5904_,
		_w5914_,
		_w5921_
	);
	LUT2 #(
		.INIT('h2)
	) name4920 (
		_w5904_,
		_w5914_,
		_w5922_
	);
	LUT2 #(
		.INIT('h1)
	) name4921 (
		_w5909_,
		_w5921_,
		_w5923_
	);
	LUT2 #(
		.INIT('h4)
	) name4922 (
		_w5922_,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h1)
	) name4923 (
		_w5920_,
		_w5924_,
		_w5925_
	);
	LUT2 #(
		.INIT('h1)
	) name4924 (
		_w5904_,
		_w5912_,
		_w5926_
	);
	LUT2 #(
		.INIT('h1)
	) name4925 (
		_w5913_,
		_w5926_,
		_w5927_
	);
	LUT2 #(
		.INIT('h1)
	) name4926 (
		_w5925_,
		_w5927_,
		_w5928_
	);
	LUT2 #(
		.INIT('h8)
	) name4927 (
		_w5925_,
		_w5927_,
		_w5929_
	);
	LUT2 #(
		.INIT('h1)
	) name4928 (
		_w5928_,
		_w5929_,
		_w5930_
	);
	LUT2 #(
		.INIT('h2)
	) name4929 (
		_w5891_,
		_w5930_,
		_w5931_
	);
	LUT2 #(
		.INIT('h4)
	) name4930 (
		_w5891_,
		_w5930_,
		_w5932_
	);
	LUT2 #(
		.INIT('h1)
	) name4931 (
		_w5931_,
		_w5932_,
		_w5933_
	);
	LUT2 #(
		.INIT('h8)
	) name4932 (
		_w5872_,
		_w5933_,
		_w5934_
	);
	LUT2 #(
		.INIT('h1)
	) name4933 (
		_w5872_,
		_w5933_,
		_w5935_
	);
	LUT2 #(
		.INIT('h1)
	) name4934 (
		_w5824_,
		_w5839_,
		_w5936_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		_w5840_,
		_w5936_,
		_w5937_
	);
	LUT2 #(
		.INIT('h1)
	) name4936 (
		_w5906_,
		_w5908_,
		_w5938_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		_w5909_,
		_w5938_,
		_w5939_
	);
	LUT2 #(
		.INIT('h8)
	) name4938 (
		_w5937_,
		_w5939_,
		_w5940_
	);
	LUT2 #(
		.INIT('h1)
	) name4939 (
		_w5846_,
		_w5859_,
		_w5941_
	);
	LUT2 #(
		.INIT('h4)
	) name4940 (
		_w5854_,
		_w5941_,
		_w5942_
	);
	LUT2 #(
		.INIT('h2)
	) name4941 (
		_w5854_,
		_w5941_,
		_w5943_
	);
	LUT2 #(
		.INIT('h1)
	) name4942 (
		_w5942_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h2)
	) name4943 (
		_w5940_,
		_w5944_,
		_w5945_
	);
	LUT2 #(
		.INIT('h4)
	) name4944 (
		_w5940_,
		_w5944_,
		_w5946_
	);
	LUT2 #(
		.INIT('h1)
	) name4945 (
		_w5915_,
		_w5924_,
		_w5947_
	);
	LUT2 #(
		.INIT('h4)
	) name4946 (
		_w5919_,
		_w5947_,
		_w5948_
	);
	LUT2 #(
		.INIT('h2)
	) name4947 (
		_w5919_,
		_w5947_,
		_w5949_
	);
	LUT2 #(
		.INIT('h1)
	) name4948 (
		_w5948_,
		_w5949_,
		_w5950_
	);
	LUT2 #(
		.INIT('h1)
	) name4949 (
		_w5946_,
		_w5950_,
		_w5951_
	);
	LUT2 #(
		.INIT('h1)
	) name4950 (
		_w5945_,
		_w5951_,
		_w5952_
	);
	LUT2 #(
		.INIT('h1)
	) name4951 (
		_w5935_,
		_w5952_,
		_w5953_
	);
	LUT2 #(
		.INIT('h1)
	) name4952 (
		_w5934_,
		_w5953_,
		_w5954_
	);
	LUT2 #(
		.INIT('h4)
	) name4953 (
		_w5868_,
		_w5954_,
		_w5955_
	);
	LUT2 #(
		.INIT('h2)
	) name4954 (
		_w5868_,
		_w5954_,
		_w5956_
	);
	LUT2 #(
		.INIT('h2)
	) name4955 (
		_w5891_,
		_w5929_,
		_w5957_
	);
	LUT2 #(
		.INIT('h1)
	) name4956 (
		_w5928_,
		_w5957_,
		_w5958_
	);
	LUT2 #(
		.INIT('h1)
	) name4957 (
		_w5956_,
		_w5958_,
		_w5959_
	);
	LUT2 #(
		.INIT('h1)
	) name4958 (
		_w5955_,
		_w5959_,
		_w5960_
	);
	LUT2 #(
		.INIT('h1)
	) name4959 (
		_w5809_,
		_w5960_,
		_w5961_
	);
	LUT2 #(
		.INIT('h8)
	) name4960 (
		_w5809_,
		_w5960_,
		_w5962_
	);
	LUT2 #(
		.INIT('h1)
	) name4961 (
		_w5955_,
		_w5956_,
		_w5963_
	);
	LUT2 #(
		.INIT('h4)
	) name4962 (
		_w5958_,
		_w5963_,
		_w5964_
	);
	LUT2 #(
		.INIT('h2)
	) name4963 (
		_w5958_,
		_w5963_,
		_w5965_
	);
	LUT2 #(
		.INIT('h1)
	) name4964 (
		_w5964_,
		_w5965_,
		_w5966_
	);
	LUT2 #(
		.INIT('h1)
	) name4965 (
		_w5804_,
		_w5805_,
		_w5967_
	);
	LUT2 #(
		.INIT('h4)
	) name4966 (
		_w5807_,
		_w5967_,
		_w5968_
	);
	LUT2 #(
		.INIT('h2)
	) name4967 (
		_w5807_,
		_w5967_,
		_w5969_
	);
	LUT2 #(
		.INIT('h1)
	) name4968 (
		_w5968_,
		_w5969_,
		_w5970_
	);
	LUT2 #(
		.INIT('h8)
	) name4969 (
		_w5966_,
		_w5970_,
		_w5971_
	);
	LUT2 #(
		.INIT('h1)
	) name4970 (
		_w5966_,
		_w5970_,
		_w5972_
	);
	LUT2 #(
		.INIT('h1)
	) name4971 (
		_w5783_,
		_w5784_,
		_w5973_
	);
	LUT2 #(
		.INIT('h4)
	) name4972 (
		_w5801_,
		_w5973_,
		_w5974_
	);
	LUT2 #(
		.INIT('h2)
	) name4973 (
		_w5801_,
		_w5973_,
		_w5975_
	);
	LUT2 #(
		.INIT('h1)
	) name4974 (
		_w5974_,
		_w5975_,
		_w5976_
	);
	LUT2 #(
		.INIT('h1)
	) name4975 (
		_w5934_,
		_w5935_,
		_w5977_
	);
	LUT2 #(
		.INIT('h4)
	) name4976 (
		_w5952_,
		_w5977_,
		_w5978_
	);
	LUT2 #(
		.INIT('h2)
	) name4977 (
		_w5952_,
		_w5977_,
		_w5979_
	);
	LUT2 #(
		.INIT('h1)
	) name4978 (
		_w5978_,
		_w5979_,
		_w5980_
	);
	LUT2 #(
		.INIT('h1)
	) name4979 (
		_w5976_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h8)
	) name4980 (
		_w5976_,
		_w5980_,
		_w5982_
	);
	LUT2 #(
		.INIT('h1)
	) name4981 (
		_w5937_,
		_w5939_,
		_w5983_
	);
	LUT2 #(
		.INIT('h1)
	) name4982 (
		_w5940_,
		_w5983_,
		_w5984_
	);
	LUT2 #(
		.INIT('h1)
	) name4983 (
		_w5786_,
		_w5788_,
		_w5985_
	);
	LUT2 #(
		.INIT('h1)
	) name4984 (
		_w5789_,
		_w5985_,
		_w5986_
	);
	LUT2 #(
		.INIT('h8)
	) name4985 (
		_w5984_,
		_w5986_,
		_w5987_
	);
	LUT2 #(
		.INIT('h1)
	) name4986 (
		_w5945_,
		_w5946_,
		_w5988_
	);
	LUT2 #(
		.INIT('h4)
	) name4987 (
		_w5950_,
		_w5988_,
		_w5989_
	);
	LUT2 #(
		.INIT('h2)
	) name4988 (
		_w5950_,
		_w5988_,
		_w5990_
	);
	LUT2 #(
		.INIT('h1)
	) name4989 (
		_w5989_,
		_w5990_,
		_w5991_
	);
	LUT2 #(
		.INIT('h8)
	) name4990 (
		_w5987_,
		_w5991_,
		_w5992_
	);
	LUT2 #(
		.INIT('h1)
	) name4991 (
		_w5987_,
		_w5991_,
		_w5993_
	);
	LUT2 #(
		.INIT('h1)
	) name4992 (
		_w5794_,
		_w5795_,
		_w5994_
	);
	LUT2 #(
		.INIT('h4)
	) name4993 (
		_w5799_,
		_w5994_,
		_w5995_
	);
	LUT2 #(
		.INIT('h2)
	) name4994 (
		_w5799_,
		_w5994_,
		_w5996_
	);
	LUT2 #(
		.INIT('h1)
	) name4995 (
		_w5995_,
		_w5996_,
		_w5997_
	);
	LUT2 #(
		.INIT('h4)
	) name4996 (
		_w5993_,
		_w5997_,
		_w5998_
	);
	LUT2 #(
		.INIT('h1)
	) name4997 (
		_w5992_,
		_w5998_,
		_w5999_
	);
	LUT2 #(
		.INIT('h4)
	) name4998 (
		_w5982_,
		_w5999_,
		_w6000_
	);
	LUT2 #(
		.INIT('h1)
	) name4999 (
		_w5981_,
		_w6000_,
		_w6001_
	);
	LUT2 #(
		.INIT('h1)
	) name5000 (
		_w5972_,
		_w6001_,
		_w6002_
	);
	LUT2 #(
		.INIT('h1)
	) name5001 (
		_w5971_,
		_w6002_,
		_w6003_
	);
	LUT2 #(
		.INIT('h1)
	) name5002 (
		_w5962_,
		_w6003_,
		_w6004_
	);
	LUT2 #(
		.INIT('h1)
	) name5003 (
		_w5961_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h1)
	) name5004 (
		_w5658_,
		_w6005_,
		_w6006_
	);
	LUT2 #(
		.INIT('h8)
	) name5005 (
		_w5658_,
		_w6005_,
		_w6007_
	);
	LUT2 #(
		.INIT('h1)
	) name5006 (
		_w5961_,
		_w5962_,
		_w6008_
	);
	LUT2 #(
		.INIT('h4)
	) name5007 (
		_w6003_,
		_w6008_,
		_w6009_
	);
	LUT2 #(
		.INIT('h2)
	) name5008 (
		_w6003_,
		_w6008_,
		_w6010_
	);
	LUT2 #(
		.INIT('h1)
	) name5009 (
		_w6009_,
		_w6010_,
		_w6011_
	);
	LUT2 #(
		.INIT('h1)
	) name5010 (
		_w5614_,
		_w5615_,
		_w6012_
	);
	LUT2 #(
		.INIT('h4)
	) name5011 (
		_w5656_,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h2)
	) name5012 (
		_w5656_,
		_w6012_,
		_w6014_
	);
	LUT2 #(
		.INIT('h1)
	) name5013 (
		_w6013_,
		_w6014_,
		_w6015_
	);
	LUT2 #(
		.INIT('h1)
	) name5014 (
		_w6011_,
		_w6015_,
		_w6016_
	);
	LUT2 #(
		.INIT('h8)
	) name5015 (
		_w6011_,
		_w6015_,
		_w6017_
	);
	LUT2 #(
		.INIT('h1)
	) name5016 (
		_w5624_,
		_w5625_,
		_w6018_
	);
	LUT2 #(
		.INIT('h4)
	) name5017 (
		_w5654_,
		_w6018_,
		_w6019_
	);
	LUT2 #(
		.INIT('h2)
	) name5018 (
		_w5654_,
		_w6018_,
		_w6020_
	);
	LUT2 #(
		.INIT('h1)
	) name5019 (
		_w6019_,
		_w6020_,
		_w6021_
	);
	LUT2 #(
		.INIT('h1)
	) name5020 (
		_w5971_,
		_w5972_,
		_w6022_
	);
	LUT2 #(
		.INIT('h4)
	) name5021 (
		_w6001_,
		_w6022_,
		_w6023_
	);
	LUT2 #(
		.INIT('h2)
	) name5022 (
		_w6001_,
		_w6022_,
		_w6024_
	);
	LUT2 #(
		.INIT('h1)
	) name5023 (
		_w6023_,
		_w6024_,
		_w6025_
	);
	LUT2 #(
		.INIT('h1)
	) name5024 (
		_w6021_,
		_w6025_,
		_w6026_
	);
	LUT2 #(
		.INIT('h8)
	) name5025 (
		_w6021_,
		_w6025_,
		_w6027_
	);
	LUT2 #(
		.INIT('h1)
	) name5026 (
		_w5981_,
		_w5982_,
		_w6028_
	);
	LUT2 #(
		.INIT('h4)
	) name5027 (
		_w5999_,
		_w6028_,
		_w6029_
	);
	LUT2 #(
		.INIT('h2)
	) name5028 (
		_w5999_,
		_w6028_,
		_w6030_
	);
	LUT2 #(
		.INIT('h1)
	) name5029 (
		_w6029_,
		_w6030_,
		_w6031_
	);
	LUT2 #(
		.INIT('h1)
	) name5030 (
		_w5634_,
		_w5635_,
		_w6032_
	);
	LUT2 #(
		.INIT('h4)
	) name5031 (
		_w5652_,
		_w6032_,
		_w6033_
	);
	LUT2 #(
		.INIT('h2)
	) name5032 (
		_w5652_,
		_w6032_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name5033 (
		_w6033_,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h1)
	) name5034 (
		_w6031_,
		_w6035_,
		_w6036_
	);
	LUT2 #(
		.INIT('h8)
	) name5035 (
		_w6031_,
		_w6035_,
		_w6037_
	);
	LUT2 #(
		.INIT('h1)
	) name5036 (
		_w5637_,
		_w5639_,
		_w6038_
	);
	LUT2 #(
		.INIT('h1)
	) name5037 (
		_w5640_,
		_w6038_,
		_w6039_
	);
	LUT2 #(
		.INIT('h1)
	) name5038 (
		_w5984_,
		_w5986_,
		_w6040_
	);
	LUT2 #(
		.INIT('h1)
	) name5039 (
		_w5987_,
		_w6040_,
		_w6041_
	);
	LUT2 #(
		.INIT('h8)
	) name5040 (
		_w6039_,
		_w6041_,
		_w6042_
	);
	LUT2 #(
		.INIT('h1)
	) name5041 (
		_w5645_,
		_w5646_,
		_w6043_
	);
	LUT2 #(
		.INIT('h4)
	) name5042 (
		_w5650_,
		_w6043_,
		_w6044_
	);
	LUT2 #(
		.INIT('h2)
	) name5043 (
		_w5650_,
		_w6043_,
		_w6045_
	);
	LUT2 #(
		.INIT('h1)
	) name5044 (
		_w6044_,
		_w6045_,
		_w6046_
	);
	LUT2 #(
		.INIT('h2)
	) name5045 (
		_w6042_,
		_w6046_,
		_w6047_
	);
	LUT2 #(
		.INIT('h4)
	) name5046 (
		_w6042_,
		_w6046_,
		_w6048_
	);
	LUT2 #(
		.INIT('h1)
	) name5047 (
		_w5992_,
		_w5993_,
		_w6049_
	);
	LUT2 #(
		.INIT('h4)
	) name5048 (
		_w5997_,
		_w6049_,
		_w6050_
	);
	LUT2 #(
		.INIT('h2)
	) name5049 (
		_w5997_,
		_w6049_,
		_w6051_
	);
	LUT2 #(
		.INIT('h1)
	) name5050 (
		_w6050_,
		_w6051_,
		_w6052_
	);
	LUT2 #(
		.INIT('h1)
	) name5051 (
		_w6048_,
		_w6052_,
		_w6053_
	);
	LUT2 #(
		.INIT('h1)
	) name5052 (
		_w6047_,
		_w6053_,
		_w6054_
	);
	LUT2 #(
		.INIT('h4)
	) name5053 (
		_w6037_,
		_w6054_,
		_w6055_
	);
	LUT2 #(
		.INIT('h1)
	) name5054 (
		_w6036_,
		_w6055_,
		_w6056_
	);
	LUT2 #(
		.INIT('h4)
	) name5055 (
		_w6027_,
		_w6056_,
		_w6057_
	);
	LUT2 #(
		.INIT('h1)
	) name5056 (
		_w6026_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h1)
	) name5057 (
		_w6017_,
		_w6058_,
		_w6059_
	);
	LUT2 #(
		.INIT('h1)
	) name5058 (
		_w6016_,
		_w6059_,
		_w6060_
	);
	LUT2 #(
		.INIT('h4)
	) name5059 (
		_w6007_,
		_w6060_,
		_w6061_
	);
	LUT2 #(
		.INIT('h1)
	) name5060 (
		_w6006_,
		_w6061_,
		_w6062_
	);
	LUT2 #(
		.INIT('h4)
	) name5061 (
		_w5311_,
		_w6062_,
		_w6063_
	);
	LUT2 #(
		.INIT('h2)
	) name5062 (
		_w5311_,
		_w6062_,
		_w6064_
	);
	LUT2 #(
		.INIT('h1)
	) name5063 (
		_w6006_,
		_w6007_,
		_w6065_
	);
	LUT2 #(
		.INIT('h4)
	) name5064 (
		_w6060_,
		_w6065_,
		_w6066_
	);
	LUT2 #(
		.INIT('h2)
	) name5065 (
		_w6060_,
		_w6065_,
		_w6067_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		_w6066_,
		_w6067_,
		_w6068_
	);
	LUT2 #(
		.INIT('h1)
	) name5067 (
		_w5255_,
		_w5256_,
		_w6069_
	);
	LUT2 #(
		.INIT('h4)
	) name5068 (
		_w5309_,
		_w6069_,
		_w6070_
	);
	LUT2 #(
		.INIT('h2)
	) name5069 (
		_w5309_,
		_w6069_,
		_w6071_
	);
	LUT2 #(
		.INIT('h1)
	) name5070 (
		_w6070_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('h2)
	) name5071 (
		_w6068_,
		_w6072_,
		_w6073_
	);
	LUT2 #(
		.INIT('h4)
	) name5072 (
		_w6068_,
		_w6072_,
		_w6074_
	);
	LUT2 #(
		.INIT('h1)
	) name5073 (
		_w6016_,
		_w6017_,
		_w6075_
	);
	LUT2 #(
		.INIT('h4)
	) name5074 (
		_w6058_,
		_w6075_,
		_w6076_
	);
	LUT2 #(
		.INIT('h2)
	) name5075 (
		_w6058_,
		_w6075_,
		_w6077_
	);
	LUT2 #(
		.INIT('h1)
	) name5076 (
		_w6076_,
		_w6077_,
		_w6078_
	);
	LUT2 #(
		.INIT('h1)
	) name5077 (
		_w5265_,
		_w5266_,
		_w6079_
	);
	LUT2 #(
		.INIT('h4)
	) name5078 (
		_w5307_,
		_w6079_,
		_w6080_
	);
	LUT2 #(
		.INIT('h2)
	) name5079 (
		_w5307_,
		_w6079_,
		_w6081_
	);
	LUT2 #(
		.INIT('h1)
	) name5080 (
		_w6080_,
		_w6081_,
		_w6082_
	);
	LUT2 #(
		.INIT('h4)
	) name5081 (
		_w6078_,
		_w6082_,
		_w6083_
	);
	LUT2 #(
		.INIT('h2)
	) name5082 (
		_w6078_,
		_w6082_,
		_w6084_
	);
	LUT2 #(
		.INIT('h1)
	) name5083 (
		_w5275_,
		_w5276_,
		_w6085_
	);
	LUT2 #(
		.INIT('h4)
	) name5084 (
		_w5305_,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h2)
	) name5085 (
		_w5305_,
		_w6085_,
		_w6087_
	);
	LUT2 #(
		.INIT('h1)
	) name5086 (
		_w6086_,
		_w6087_,
		_w6088_
	);
	LUT2 #(
		.INIT('h1)
	) name5087 (
		_w6026_,
		_w6027_,
		_w6089_
	);
	LUT2 #(
		.INIT('h8)
	) name5088 (
		_w6056_,
		_w6089_,
		_w6090_
	);
	LUT2 #(
		.INIT('h1)
	) name5089 (
		_w6056_,
		_w6089_,
		_w6091_
	);
	LUT2 #(
		.INIT('h1)
	) name5090 (
		_w6090_,
		_w6091_,
		_w6092_
	);
	LUT2 #(
		.INIT('h2)
	) name5091 (
		_w6088_,
		_w6092_,
		_w6093_
	);
	LUT2 #(
		.INIT('h4)
	) name5092 (
		_w6088_,
		_w6092_,
		_w6094_
	);
	LUT2 #(
		.INIT('h1)
	) name5093 (
		_w6036_,
		_w6037_,
		_w6095_
	);
	LUT2 #(
		.INIT('h4)
	) name5094 (
		_w6054_,
		_w6095_,
		_w6096_
	);
	LUT2 #(
		.INIT('h2)
	) name5095 (
		_w6054_,
		_w6095_,
		_w6097_
	);
	LUT2 #(
		.INIT('h1)
	) name5096 (
		_w6096_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h1)
	) name5097 (
		_w5285_,
		_w5286_,
		_w6099_
	);
	LUT2 #(
		.INIT('h4)
	) name5098 (
		_w5303_,
		_w6099_,
		_w6100_
	);
	LUT2 #(
		.INIT('h2)
	) name5099 (
		_w5303_,
		_w6099_,
		_w6101_
	);
	LUT2 #(
		.INIT('h1)
	) name5100 (
		_w6100_,
		_w6101_,
		_w6102_
	);
	LUT2 #(
		.INIT('h1)
	) name5101 (
		_w6098_,
		_w6102_,
		_w6103_
	);
	LUT2 #(
		.INIT('h8)
	) name5102 (
		_w6098_,
		_w6102_,
		_w6104_
	);
	LUT2 #(
		.INIT('h1)
	) name5103 (
		_w5288_,
		_w5290_,
		_w6105_
	);
	LUT2 #(
		.INIT('h1)
	) name5104 (
		_w5291_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name5105 (
		_w6039_,
		_w6041_,
		_w6107_
	);
	LUT2 #(
		.INIT('h1)
	) name5106 (
		_w6042_,
		_w6107_,
		_w6108_
	);
	LUT2 #(
		.INIT('h8)
	) name5107 (
		_w6106_,
		_w6108_,
		_w6109_
	);
	LUT2 #(
		.INIT('h1)
	) name5108 (
		_w5296_,
		_w5297_,
		_w6110_
	);
	LUT2 #(
		.INIT('h4)
	) name5109 (
		_w5301_,
		_w6110_,
		_w6111_
	);
	LUT2 #(
		.INIT('h2)
	) name5110 (
		_w5301_,
		_w6110_,
		_w6112_
	);
	LUT2 #(
		.INIT('h1)
	) name5111 (
		_w6111_,
		_w6112_,
		_w6113_
	);
	LUT2 #(
		.INIT('h8)
	) name5112 (
		_w6109_,
		_w6113_,
		_w6114_
	);
	LUT2 #(
		.INIT('h1)
	) name5113 (
		_w6109_,
		_w6113_,
		_w6115_
	);
	LUT2 #(
		.INIT('h1)
	) name5114 (
		_w6047_,
		_w6048_,
		_w6116_
	);
	LUT2 #(
		.INIT('h4)
	) name5115 (
		_w6052_,
		_w6116_,
		_w6117_
	);
	LUT2 #(
		.INIT('h2)
	) name5116 (
		_w6052_,
		_w6116_,
		_w6118_
	);
	LUT2 #(
		.INIT('h1)
	) name5117 (
		_w6117_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h4)
	) name5118 (
		_w6115_,
		_w6119_,
		_w6120_
	);
	LUT2 #(
		.INIT('h1)
	) name5119 (
		_w6114_,
		_w6120_,
		_w6121_
	);
	LUT2 #(
		.INIT('h4)
	) name5120 (
		_w6104_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('h1)
	) name5121 (
		_w6103_,
		_w6122_,
		_w6123_
	);
	LUT2 #(
		.INIT('h1)
	) name5122 (
		_w6094_,
		_w6123_,
		_w6124_
	);
	LUT2 #(
		.INIT('h1)
	) name5123 (
		_w6093_,
		_w6124_,
		_w6125_
	);
	LUT2 #(
		.INIT('h1)
	) name5124 (
		_w6084_,
		_w6125_,
		_w6126_
	);
	LUT2 #(
		.INIT('h1)
	) name5125 (
		_w6083_,
		_w6126_,
		_w6127_
	);
	LUT2 #(
		.INIT('h4)
	) name5126 (
		_w6074_,
		_w6127_,
		_w6128_
	);
	LUT2 #(
		.INIT('h1)
	) name5127 (
		_w6073_,
		_w6128_,
		_w6129_
	);
	LUT2 #(
		.INIT('h1)
	) name5128 (
		_w6064_,
		_w6129_,
		_w6130_
	);
	LUT2 #(
		.INIT('h1)
	) name5129 (
		_w6063_,
		_w6130_,
		_w6131_
	);
	LUT2 #(
		.INIT('h1)
	) name5130 (
		_w4543_,
		_w6131_,
		_w6132_
	);
	LUT2 #(
		.INIT('h8)
	) name5131 (
		_w4543_,
		_w6131_,
		_w6133_
	);
	LUT2 #(
		.INIT('h1)
	) name5132 (
		_w4475_,
		_w4476_,
		_w6134_
	);
	LUT2 #(
		.INIT('h4)
	) name5133 (
		_w4541_,
		_w6134_,
		_w6135_
	);
	LUT2 #(
		.INIT('h2)
	) name5134 (
		_w4541_,
		_w6134_,
		_w6136_
	);
	LUT2 #(
		.INIT('h1)
	) name5135 (
		_w6135_,
		_w6136_,
		_w6137_
	);
	LUT2 #(
		.INIT('h1)
	) name5136 (
		_w6063_,
		_w6064_,
		_w6138_
	);
	LUT2 #(
		.INIT('h4)
	) name5137 (
		_w6129_,
		_w6138_,
		_w6139_
	);
	LUT2 #(
		.INIT('h2)
	) name5138 (
		_w6129_,
		_w6138_,
		_w6140_
	);
	LUT2 #(
		.INIT('h1)
	) name5139 (
		_w6139_,
		_w6140_,
		_w6141_
	);
	LUT2 #(
		.INIT('h2)
	) name5140 (
		_w6137_,
		_w6141_,
		_w6142_
	);
	LUT2 #(
		.INIT('h4)
	) name5141 (
		_w6137_,
		_w6141_,
		_w6143_
	);
	LUT2 #(
		.INIT('h1)
	) name5142 (
		_w6073_,
		_w6074_,
		_w6144_
	);
	LUT2 #(
		.INIT('h4)
	) name5143 (
		_w6127_,
		_w6144_,
		_w6145_
	);
	LUT2 #(
		.INIT('h2)
	) name5144 (
		_w6127_,
		_w6144_,
		_w6146_
	);
	LUT2 #(
		.INIT('h1)
	) name5145 (
		_w6145_,
		_w6146_,
		_w6147_
	);
	LUT2 #(
		.INIT('h1)
	) name5146 (
		_w4485_,
		_w4486_,
		_w6148_
	);
	LUT2 #(
		.INIT('h4)
	) name5147 (
		_w4539_,
		_w6148_,
		_w6149_
	);
	LUT2 #(
		.INIT('h2)
	) name5148 (
		_w4539_,
		_w6148_,
		_w6150_
	);
	LUT2 #(
		.INIT('h1)
	) name5149 (
		_w6149_,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h1)
	) name5150 (
		_w6147_,
		_w6151_,
		_w6152_
	);
	LUT2 #(
		.INIT('h8)
	) name5151 (
		_w6147_,
		_w6151_,
		_w6153_
	);
	LUT2 #(
		.INIT('h1)
	) name5152 (
		_w6083_,
		_w6084_,
		_w6154_
	);
	LUT2 #(
		.INIT('h4)
	) name5153 (
		_w6125_,
		_w6154_,
		_w6155_
	);
	LUT2 #(
		.INIT('h2)
	) name5154 (
		_w6125_,
		_w6154_,
		_w6156_
	);
	LUT2 #(
		.INIT('h1)
	) name5155 (
		_w6155_,
		_w6156_,
		_w6157_
	);
	LUT2 #(
		.INIT('h1)
	) name5156 (
		_w4495_,
		_w4496_,
		_w6158_
	);
	LUT2 #(
		.INIT('h4)
	) name5157 (
		_w4537_,
		_w6158_,
		_w6159_
	);
	LUT2 #(
		.INIT('h2)
	) name5158 (
		_w4537_,
		_w6158_,
		_w6160_
	);
	LUT2 #(
		.INIT('h1)
	) name5159 (
		_w6159_,
		_w6160_,
		_w6161_
	);
	LUT2 #(
		.INIT('h1)
	) name5160 (
		_w6157_,
		_w6161_,
		_w6162_
	);
	LUT2 #(
		.INIT('h8)
	) name5161 (
		_w6157_,
		_w6161_,
		_w6163_
	);
	LUT2 #(
		.INIT('h1)
	) name5162 (
		_w4505_,
		_w4506_,
		_w6164_
	);
	LUT2 #(
		.INIT('h4)
	) name5163 (
		_w4535_,
		_w6164_,
		_w6165_
	);
	LUT2 #(
		.INIT('h2)
	) name5164 (
		_w4535_,
		_w6164_,
		_w6166_
	);
	LUT2 #(
		.INIT('h1)
	) name5165 (
		_w6165_,
		_w6166_,
		_w6167_
	);
	LUT2 #(
		.INIT('h1)
	) name5166 (
		_w6093_,
		_w6094_,
		_w6168_
	);
	LUT2 #(
		.INIT('h4)
	) name5167 (
		_w6123_,
		_w6168_,
		_w6169_
	);
	LUT2 #(
		.INIT('h2)
	) name5168 (
		_w6123_,
		_w6168_,
		_w6170_
	);
	LUT2 #(
		.INIT('h1)
	) name5169 (
		_w6169_,
		_w6170_,
		_w6171_
	);
	LUT2 #(
		.INIT('h1)
	) name5170 (
		_w6167_,
		_w6171_,
		_w6172_
	);
	LUT2 #(
		.INIT('h8)
	) name5171 (
		_w6167_,
		_w6171_,
		_w6173_
	);
	LUT2 #(
		.INIT('h1)
	) name5172 (
		_w6103_,
		_w6104_,
		_w6174_
	);
	LUT2 #(
		.INIT('h4)
	) name5173 (
		_w6121_,
		_w6174_,
		_w6175_
	);
	LUT2 #(
		.INIT('h2)
	) name5174 (
		_w6121_,
		_w6174_,
		_w6176_
	);
	LUT2 #(
		.INIT('h1)
	) name5175 (
		_w6175_,
		_w6176_,
		_w6177_
	);
	LUT2 #(
		.INIT('h1)
	) name5176 (
		_w4515_,
		_w4516_,
		_w6178_
	);
	LUT2 #(
		.INIT('h4)
	) name5177 (
		_w4533_,
		_w6178_,
		_w6179_
	);
	LUT2 #(
		.INIT('h2)
	) name5178 (
		_w4533_,
		_w6178_,
		_w6180_
	);
	LUT2 #(
		.INIT('h1)
	) name5179 (
		_w6179_,
		_w6180_,
		_w6181_
	);
	LUT2 #(
		.INIT('h1)
	) name5180 (
		_w6177_,
		_w6181_,
		_w6182_
	);
	LUT2 #(
		.INIT('h8)
	) name5181 (
		_w6177_,
		_w6181_,
		_w6183_
	);
	LUT2 #(
		.INIT('h1)
	) name5182 (
		_w4518_,
		_w4520_,
		_w6184_
	);
	LUT2 #(
		.INIT('h1)
	) name5183 (
		_w4521_,
		_w6184_,
		_w6185_
	);
	LUT2 #(
		.INIT('h1)
	) name5184 (
		_w6106_,
		_w6108_,
		_w6186_
	);
	LUT2 #(
		.INIT('h1)
	) name5185 (
		_w6109_,
		_w6186_,
		_w6187_
	);
	LUT2 #(
		.INIT('h8)
	) name5186 (
		_w6185_,
		_w6187_,
		_w6188_
	);
	LUT2 #(
		.INIT('h1)
	) name5187 (
		_w4526_,
		_w4527_,
		_w6189_
	);
	LUT2 #(
		.INIT('h4)
	) name5188 (
		_w4531_,
		_w6189_,
		_w6190_
	);
	LUT2 #(
		.INIT('h2)
	) name5189 (
		_w4531_,
		_w6189_,
		_w6191_
	);
	LUT2 #(
		.INIT('h1)
	) name5190 (
		_w6190_,
		_w6191_,
		_w6192_
	);
	LUT2 #(
		.INIT('h2)
	) name5191 (
		_w6188_,
		_w6192_,
		_w6193_
	);
	LUT2 #(
		.INIT('h4)
	) name5192 (
		_w6188_,
		_w6192_,
		_w6194_
	);
	LUT2 #(
		.INIT('h1)
	) name5193 (
		_w6114_,
		_w6115_,
		_w6195_
	);
	LUT2 #(
		.INIT('h8)
	) name5194 (
		_w6119_,
		_w6195_,
		_w6196_
	);
	LUT2 #(
		.INIT('h1)
	) name5195 (
		_w6119_,
		_w6195_,
		_w6197_
	);
	LUT2 #(
		.INIT('h1)
	) name5196 (
		_w6196_,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h4)
	) name5197 (
		_w6194_,
		_w6198_,
		_w6199_
	);
	LUT2 #(
		.INIT('h1)
	) name5198 (
		_w6193_,
		_w6199_,
		_w6200_
	);
	LUT2 #(
		.INIT('h4)
	) name5199 (
		_w6183_,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h1)
	) name5200 (
		_w6182_,
		_w6201_,
		_w6202_
	);
	LUT2 #(
		.INIT('h4)
	) name5201 (
		_w6173_,
		_w6202_,
		_w6203_
	);
	LUT2 #(
		.INIT('h1)
	) name5202 (
		_w6172_,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h1)
	) name5203 (
		_w6163_,
		_w6204_,
		_w6205_
	);
	LUT2 #(
		.INIT('h1)
	) name5204 (
		_w6162_,
		_w6205_,
		_w6206_
	);
	LUT2 #(
		.INIT('h1)
	) name5205 (
		_w6153_,
		_w6206_,
		_w6207_
	);
	LUT2 #(
		.INIT('h1)
	) name5206 (
		_w6152_,
		_w6207_,
		_w6208_
	);
	LUT2 #(
		.INIT('h4)
	) name5207 (
		_w6143_,
		_w6208_,
		_w6209_
	);
	LUT2 #(
		.INIT('h1)
	) name5208 (
		_w6142_,
		_w6209_,
		_w6210_
	);
	LUT2 #(
		.INIT('h4)
	) name5209 (
		_w6133_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h1)
	) name5210 (
		_w6132_,
		_w6211_,
		_w6212_
	);
	LUT2 #(
		.INIT('h4)
	) name5211 (
		_w2945_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h2)
	) name5212 (
		_w2945_,
		_w6212_,
		_w6214_
	);
	LUT2 #(
		.INIT('h1)
	) name5213 (
		_w6213_,
		_w6214_,
		_w6215_
	);
	LUT2 #(
		.INIT('h8)
	) name5214 (
		_w2110_,
		_w2877_,
		_w6216_
	);
	LUT2 #(
		.INIT('h1)
	) name5215 (
		_w2108_,
		_w2944_,
		_w6217_
	);
	LUT2 #(
		.INIT('h1)
	) name5216 (
		_w2945_,
		_w6217_,
		_w6218_
	);
	LUT2 #(
		.INIT('h1)
	) name5217 (
		_w6216_,
		_w6218_,
		_w6219_
	);
	LUT2 #(
		.INIT('h1)
	) name5218 (
		_w6132_,
		_w6133_,
		_w6220_
	);
	LUT2 #(
		.INIT('h4)
	) name5219 (
		_w6210_,
		_w6220_,
		_w6221_
	);
	LUT2 #(
		.INIT('h2)
	) name5220 (
		_w6210_,
		_w6220_,
		_w6222_
	);
	LUT2 #(
		.INIT('h1)
	) name5221 (
		_w6221_,
		_w6222_,
		_w6223_
	);
	LUT2 #(
		.INIT('h8)
	) name5222 (
		_w6219_,
		_w6223_,
		_w6224_
	);
	LUT2 #(
		.INIT('h1)
	) name5223 (
		_w6219_,
		_w6223_,
		_w6225_
	);
	LUT2 #(
		.INIT('h1)
	) name5224 (
		_w2878_,
		_w6216_,
		_w6226_
	);
	LUT2 #(
		.INIT('h4)
	) name5225 (
		_w2943_,
		_w6226_,
		_w6227_
	);
	LUT2 #(
		.INIT('h2)
	) name5226 (
		_w2943_,
		_w6226_,
		_w6228_
	);
	LUT2 #(
		.INIT('h1)
	) name5227 (
		_w6227_,
		_w6228_,
		_w6229_
	);
	LUT2 #(
		.INIT('h1)
	) name5228 (
		_w6142_,
		_w6143_,
		_w6230_
	);
	LUT2 #(
		.INIT('h4)
	) name5229 (
		_w6208_,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h2)
	) name5230 (
		_w6208_,
		_w6230_,
		_w6232_
	);
	LUT2 #(
		.INIT('h1)
	) name5231 (
		_w6231_,
		_w6232_,
		_w6233_
	);
	LUT2 #(
		.INIT('h2)
	) name5232 (
		_w6229_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h4)
	) name5233 (
		_w6229_,
		_w6233_,
		_w6235_
	);
	LUT2 #(
		.INIT('h1)
	) name5234 (
		_w2887_,
		_w2888_,
		_w6236_
	);
	LUT2 #(
		.INIT('h4)
	) name5235 (
		_w2941_,
		_w6236_,
		_w6237_
	);
	LUT2 #(
		.INIT('h2)
	) name5236 (
		_w2941_,
		_w6236_,
		_w6238_
	);
	LUT2 #(
		.INIT('h1)
	) name5237 (
		_w6237_,
		_w6238_,
		_w6239_
	);
	LUT2 #(
		.INIT('h1)
	) name5238 (
		_w6152_,
		_w6153_,
		_w6240_
	);
	LUT2 #(
		.INIT('h4)
	) name5239 (
		_w6206_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('h2)
	) name5240 (
		_w6206_,
		_w6240_,
		_w6242_
	);
	LUT2 #(
		.INIT('h1)
	) name5241 (
		_w6241_,
		_w6242_,
		_w6243_
	);
	LUT2 #(
		.INIT('h2)
	) name5242 (
		_w6239_,
		_w6243_,
		_w6244_
	);
	LUT2 #(
		.INIT('h4)
	) name5243 (
		_w6239_,
		_w6243_,
		_w6245_
	);
	LUT2 #(
		.INIT('h1)
	) name5244 (
		_w2897_,
		_w2898_,
		_w6246_
	);
	LUT2 #(
		.INIT('h4)
	) name5245 (
		_w2939_,
		_w6246_,
		_w6247_
	);
	LUT2 #(
		.INIT('h2)
	) name5246 (
		_w2939_,
		_w6246_,
		_w6248_
	);
	LUT2 #(
		.INIT('h1)
	) name5247 (
		_w6247_,
		_w6248_,
		_w6249_
	);
	LUT2 #(
		.INIT('h1)
	) name5248 (
		_w6162_,
		_w6163_,
		_w6250_
	);
	LUT2 #(
		.INIT('h4)
	) name5249 (
		_w6204_,
		_w6250_,
		_w6251_
	);
	LUT2 #(
		.INIT('h2)
	) name5250 (
		_w6204_,
		_w6250_,
		_w6252_
	);
	LUT2 #(
		.INIT('h1)
	) name5251 (
		_w6251_,
		_w6252_,
		_w6253_
	);
	LUT2 #(
		.INIT('h2)
	) name5252 (
		_w6249_,
		_w6253_,
		_w6254_
	);
	LUT2 #(
		.INIT('h4)
	) name5253 (
		_w6249_,
		_w6253_,
		_w6255_
	);
	LUT2 #(
		.INIT('h1)
	) name5254 (
		_w6172_,
		_w6173_,
		_w6256_
	);
	LUT2 #(
		.INIT('h4)
	) name5255 (
		_w6202_,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h2)
	) name5256 (
		_w6202_,
		_w6256_,
		_w6258_
	);
	LUT2 #(
		.INIT('h1)
	) name5257 (
		_w6257_,
		_w6258_,
		_w6259_
	);
	LUT2 #(
		.INIT('h1)
	) name5258 (
		_w2907_,
		_w2908_,
		_w6260_
	);
	LUT2 #(
		.INIT('h4)
	) name5259 (
		_w2937_,
		_w6260_,
		_w6261_
	);
	LUT2 #(
		.INIT('h2)
	) name5260 (
		_w2937_,
		_w6260_,
		_w6262_
	);
	LUT2 #(
		.INIT('h1)
	) name5261 (
		_w6261_,
		_w6262_,
		_w6263_
	);
	LUT2 #(
		.INIT('h1)
	) name5262 (
		_w6259_,
		_w6263_,
		_w6264_
	);
	LUT2 #(
		.INIT('h8)
	) name5263 (
		_w6259_,
		_w6263_,
		_w6265_
	);
	LUT2 #(
		.INIT('h1)
	) name5264 (
		_w2917_,
		_w2918_,
		_w6266_
	);
	LUT2 #(
		.INIT('h4)
	) name5265 (
		_w2935_,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h2)
	) name5266 (
		_w2935_,
		_w6266_,
		_w6268_
	);
	LUT2 #(
		.INIT('h1)
	) name5267 (
		_w6267_,
		_w6268_,
		_w6269_
	);
	LUT2 #(
		.INIT('h1)
	) name5268 (
		_w6182_,
		_w6183_,
		_w6270_
	);
	LUT2 #(
		.INIT('h4)
	) name5269 (
		_w6200_,
		_w6270_,
		_w6271_
	);
	LUT2 #(
		.INIT('h2)
	) name5270 (
		_w6200_,
		_w6270_,
		_w6272_
	);
	LUT2 #(
		.INIT('h1)
	) name5271 (
		_w6271_,
		_w6272_,
		_w6273_
	);
	LUT2 #(
		.INIT('h1)
	) name5272 (
		_w6269_,
		_w6273_,
		_w6274_
	);
	LUT2 #(
		.INIT('h8)
	) name5273 (
		_w6269_,
		_w6273_,
		_w6275_
	);
	LUT2 #(
		.INIT('h1)
	) name5274 (
		_w2920_,
		_w2922_,
		_w6276_
	);
	LUT2 #(
		.INIT('h1)
	) name5275 (
		_w2923_,
		_w6276_,
		_w6277_
	);
	LUT2 #(
		.INIT('h1)
	) name5276 (
		_w6185_,
		_w6187_,
		_w6278_
	);
	LUT2 #(
		.INIT('h1)
	) name5277 (
		_w6188_,
		_w6278_,
		_w6279_
	);
	LUT2 #(
		.INIT('h8)
	) name5278 (
		_w6277_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h1)
	) name5279 (
		_w6193_,
		_w6194_,
		_w6281_
	);
	LUT2 #(
		.INIT('h4)
	) name5280 (
		_w6198_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h2)
	) name5281 (
		_w6198_,
		_w6281_,
		_w6283_
	);
	LUT2 #(
		.INIT('h1)
	) name5282 (
		_w6282_,
		_w6283_,
		_w6284_
	);
	LUT2 #(
		.INIT('h2)
	) name5283 (
		_w6280_,
		_w6284_,
		_w6285_
	);
	LUT2 #(
		.INIT('h4)
	) name5284 (
		_w6280_,
		_w6284_,
		_w6286_
	);
	LUT2 #(
		.INIT('h1)
	) name5285 (
		_w2928_,
		_w2929_,
		_w6287_
	);
	LUT2 #(
		.INIT('h4)
	) name5286 (
		_w2933_,
		_w6287_,
		_w6288_
	);
	LUT2 #(
		.INIT('h2)
	) name5287 (
		_w2933_,
		_w6287_,
		_w6289_
	);
	LUT2 #(
		.INIT('h1)
	) name5288 (
		_w6288_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h4)
	) name5289 (
		_w6286_,
		_w6290_,
		_w6291_
	);
	LUT2 #(
		.INIT('h1)
	) name5290 (
		_w6285_,
		_w6291_,
		_w6292_
	);
	LUT2 #(
		.INIT('h4)
	) name5291 (
		_w6275_,
		_w6292_,
		_w6293_
	);
	LUT2 #(
		.INIT('h1)
	) name5292 (
		_w6274_,
		_w6293_,
		_w6294_
	);
	LUT2 #(
		.INIT('h4)
	) name5293 (
		_w6265_,
		_w6294_,
		_w6295_
	);
	LUT2 #(
		.INIT('h1)
	) name5294 (
		_w6264_,
		_w6295_,
		_w6296_
	);
	LUT2 #(
		.INIT('h4)
	) name5295 (
		_w6255_,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h1)
	) name5296 (
		_w6254_,
		_w6297_,
		_w6298_
	);
	LUT2 #(
		.INIT('h1)
	) name5297 (
		_w6245_,
		_w6298_,
		_w6299_
	);
	LUT2 #(
		.INIT('h1)
	) name5298 (
		_w6244_,
		_w6299_,
		_w6300_
	);
	LUT2 #(
		.INIT('h1)
	) name5299 (
		_w6235_,
		_w6300_,
		_w6301_
	);
	LUT2 #(
		.INIT('h1)
	) name5300 (
		_w6234_,
		_w6301_,
		_w6302_
	);
	LUT2 #(
		.INIT('h1)
	) name5301 (
		_w6225_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h1)
	) name5302 (
		_w6224_,
		_w6303_,
		_w6304_
	);
	LUT2 #(
		.INIT('h2)
	) name5303 (
		_w6215_,
		_w6304_,
		_w6305_
	);
	LUT2 #(
		.INIT('h4)
	) name5304 (
		_w6215_,
		_w6304_,
		_w6306_
	);
	LUT2 #(
		.INIT('h1)
	) name5305 (
		_w6305_,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h8)
	) name5306 (
		\A[835] ,
		\A[836] ,
		_w6308_
	);
	LUT2 #(
		.INIT('h1)
	) name5307 (
		\A[835] ,
		\A[836] ,
		_w6309_
	);
	LUT2 #(
		.INIT('h1)
	) name5308 (
		_w6308_,
		_w6309_,
		_w6310_
	);
	LUT2 #(
		.INIT('h8)
	) name5309 (
		\A[837] ,
		_w6310_,
		_w6311_
	);
	LUT2 #(
		.INIT('h1)
	) name5310 (
		\A[837] ,
		_w6310_,
		_w6312_
	);
	LUT2 #(
		.INIT('h1)
	) name5311 (
		_w6311_,
		_w6312_,
		_w6313_
	);
	LUT2 #(
		.INIT('h8)
	) name5312 (
		\A[838] ,
		\A[839] ,
		_w6314_
	);
	LUT2 #(
		.INIT('h1)
	) name5313 (
		\A[838] ,
		\A[839] ,
		_w6315_
	);
	LUT2 #(
		.INIT('h1)
	) name5314 (
		_w6314_,
		_w6315_,
		_w6316_
	);
	LUT2 #(
		.INIT('h8)
	) name5315 (
		\A[840] ,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h1)
	) name5316 (
		\A[840] ,
		_w6316_,
		_w6318_
	);
	LUT2 #(
		.INIT('h1)
	) name5317 (
		_w6317_,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h8)
	) name5318 (
		_w6313_,
		_w6319_,
		_w6320_
	);
	LUT2 #(
		.INIT('h1)
	) name5319 (
		_w6313_,
		_w6319_,
		_w6321_
	);
	LUT2 #(
		.INIT('h1)
	) name5320 (
		_w6320_,
		_w6321_,
		_w6322_
	);
	LUT2 #(
		.INIT('h8)
	) name5321 (
		\A[841] ,
		\A[842] ,
		_w6323_
	);
	LUT2 #(
		.INIT('h1)
	) name5322 (
		\A[841] ,
		\A[842] ,
		_w6324_
	);
	LUT2 #(
		.INIT('h1)
	) name5323 (
		_w6323_,
		_w6324_,
		_w6325_
	);
	LUT2 #(
		.INIT('h8)
	) name5324 (
		\A[843] ,
		_w6325_,
		_w6326_
	);
	LUT2 #(
		.INIT('h1)
	) name5325 (
		\A[843] ,
		_w6325_,
		_w6327_
	);
	LUT2 #(
		.INIT('h1)
	) name5326 (
		_w6326_,
		_w6327_,
		_w6328_
	);
	LUT2 #(
		.INIT('h8)
	) name5327 (
		\A[844] ,
		\A[845] ,
		_w6329_
	);
	LUT2 #(
		.INIT('h1)
	) name5328 (
		\A[844] ,
		\A[845] ,
		_w6330_
	);
	LUT2 #(
		.INIT('h1)
	) name5329 (
		_w6329_,
		_w6330_,
		_w6331_
	);
	LUT2 #(
		.INIT('h8)
	) name5330 (
		\A[846] ,
		_w6331_,
		_w6332_
	);
	LUT2 #(
		.INIT('h1)
	) name5331 (
		\A[846] ,
		_w6331_,
		_w6333_
	);
	LUT2 #(
		.INIT('h1)
	) name5332 (
		_w6332_,
		_w6333_,
		_w6334_
	);
	LUT2 #(
		.INIT('h8)
	) name5333 (
		_w6328_,
		_w6334_,
		_w6335_
	);
	LUT2 #(
		.INIT('h1)
	) name5334 (
		_w6328_,
		_w6334_,
		_w6336_
	);
	LUT2 #(
		.INIT('h1)
	) name5335 (
		_w6335_,
		_w6336_,
		_w6337_
	);
	LUT2 #(
		.INIT('h8)
	) name5336 (
		_w6322_,
		_w6337_,
		_w6338_
	);
	LUT2 #(
		.INIT('h1)
	) name5337 (
		_w6329_,
		_w6332_,
		_w6339_
	);
	LUT2 #(
		.INIT('h1)
	) name5338 (
		_w6323_,
		_w6326_,
		_w6340_
	);
	LUT2 #(
		.INIT('h8)
	) name5339 (
		_w6339_,
		_w6340_,
		_w6341_
	);
	LUT2 #(
		.INIT('h1)
	) name5340 (
		_w6339_,
		_w6340_,
		_w6342_
	);
	LUT2 #(
		.INIT('h1)
	) name5341 (
		_w6341_,
		_w6342_,
		_w6343_
	);
	LUT2 #(
		.INIT('h8)
	) name5342 (
		_w6338_,
		_w6343_,
		_w6344_
	);
	LUT2 #(
		.INIT('h1)
	) name5343 (
		_w6308_,
		_w6311_,
		_w6345_
	);
	LUT2 #(
		.INIT('h8)
	) name5344 (
		_w6314_,
		_w6320_,
		_w6346_
	);
	LUT2 #(
		.INIT('h1)
	) name5345 (
		_w6314_,
		_w6317_,
		_w6347_
	);
	LUT2 #(
		.INIT('h4)
	) name5346 (
		_w6320_,
		_w6347_,
		_w6348_
	);
	LUT2 #(
		.INIT('h1)
	) name5347 (
		_w6346_,
		_w6348_,
		_w6349_
	);
	LUT2 #(
		.INIT('h2)
	) name5348 (
		_w6345_,
		_w6349_,
		_w6350_
	);
	LUT2 #(
		.INIT('h4)
	) name5349 (
		_w6345_,
		_w6349_,
		_w6351_
	);
	LUT2 #(
		.INIT('h1)
	) name5350 (
		_w6350_,
		_w6351_,
		_w6352_
	);
	LUT2 #(
		.INIT('h1)
	) name5351 (
		_w6344_,
		_w6352_,
		_w6353_
	);
	LUT2 #(
		.INIT('h4)
	) name5352 (
		_w6335_,
		_w6343_,
		_w6354_
	);
	LUT2 #(
		.INIT('h2)
	) name5353 (
		_w6335_,
		_w6343_,
		_w6355_
	);
	LUT2 #(
		.INIT('h1)
	) name5354 (
		_w6338_,
		_w6354_,
		_w6356_
	);
	LUT2 #(
		.INIT('h4)
	) name5355 (
		_w6355_,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h1)
	) name5356 (
		_w6353_,
		_w6357_,
		_w6358_
	);
	LUT2 #(
		.INIT('h2)
	) name5357 (
		_w6335_,
		_w6341_,
		_w6359_
	);
	LUT2 #(
		.INIT('h1)
	) name5358 (
		_w6342_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h2)
	) name5359 (
		_w6358_,
		_w6360_,
		_w6361_
	);
	LUT2 #(
		.INIT('h4)
	) name5360 (
		_w6358_,
		_w6360_,
		_w6362_
	);
	LUT2 #(
		.INIT('h1)
	) name5361 (
		_w6345_,
		_w6348_,
		_w6363_
	);
	LUT2 #(
		.INIT('h1)
	) name5362 (
		_w6346_,
		_w6363_,
		_w6364_
	);
	LUT2 #(
		.INIT('h1)
	) name5363 (
		_w6362_,
		_w6364_,
		_w6365_
	);
	LUT2 #(
		.INIT('h1)
	) name5364 (
		_w6361_,
		_w6365_,
		_w6366_
	);
	LUT2 #(
		.INIT('h8)
	) name5365 (
		\A[823] ,
		\A[824] ,
		_w6367_
	);
	LUT2 #(
		.INIT('h1)
	) name5366 (
		\A[823] ,
		\A[824] ,
		_w6368_
	);
	LUT2 #(
		.INIT('h1)
	) name5367 (
		_w6367_,
		_w6368_,
		_w6369_
	);
	LUT2 #(
		.INIT('h8)
	) name5368 (
		\A[825] ,
		_w6369_,
		_w6370_
	);
	LUT2 #(
		.INIT('h1)
	) name5369 (
		\A[825] ,
		_w6369_,
		_w6371_
	);
	LUT2 #(
		.INIT('h1)
	) name5370 (
		_w6370_,
		_w6371_,
		_w6372_
	);
	LUT2 #(
		.INIT('h8)
	) name5371 (
		\A[826] ,
		\A[827] ,
		_w6373_
	);
	LUT2 #(
		.INIT('h1)
	) name5372 (
		\A[826] ,
		\A[827] ,
		_w6374_
	);
	LUT2 #(
		.INIT('h1)
	) name5373 (
		_w6373_,
		_w6374_,
		_w6375_
	);
	LUT2 #(
		.INIT('h8)
	) name5374 (
		\A[828] ,
		_w6375_,
		_w6376_
	);
	LUT2 #(
		.INIT('h1)
	) name5375 (
		\A[828] ,
		_w6375_,
		_w6377_
	);
	LUT2 #(
		.INIT('h1)
	) name5376 (
		_w6376_,
		_w6377_,
		_w6378_
	);
	LUT2 #(
		.INIT('h8)
	) name5377 (
		_w6372_,
		_w6378_,
		_w6379_
	);
	LUT2 #(
		.INIT('h1)
	) name5378 (
		_w6372_,
		_w6378_,
		_w6380_
	);
	LUT2 #(
		.INIT('h1)
	) name5379 (
		_w6379_,
		_w6380_,
		_w6381_
	);
	LUT2 #(
		.INIT('h8)
	) name5380 (
		\A[829] ,
		\A[830] ,
		_w6382_
	);
	LUT2 #(
		.INIT('h1)
	) name5381 (
		\A[829] ,
		\A[830] ,
		_w6383_
	);
	LUT2 #(
		.INIT('h1)
	) name5382 (
		_w6382_,
		_w6383_,
		_w6384_
	);
	LUT2 #(
		.INIT('h8)
	) name5383 (
		\A[831] ,
		_w6384_,
		_w6385_
	);
	LUT2 #(
		.INIT('h1)
	) name5384 (
		\A[831] ,
		_w6384_,
		_w6386_
	);
	LUT2 #(
		.INIT('h1)
	) name5385 (
		_w6385_,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h8)
	) name5386 (
		\A[832] ,
		\A[833] ,
		_w6388_
	);
	LUT2 #(
		.INIT('h1)
	) name5387 (
		\A[832] ,
		\A[833] ,
		_w6389_
	);
	LUT2 #(
		.INIT('h1)
	) name5388 (
		_w6388_,
		_w6389_,
		_w6390_
	);
	LUT2 #(
		.INIT('h8)
	) name5389 (
		\A[834] ,
		_w6390_,
		_w6391_
	);
	LUT2 #(
		.INIT('h1)
	) name5390 (
		\A[834] ,
		_w6390_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name5391 (
		_w6391_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h8)
	) name5392 (
		_w6387_,
		_w6393_,
		_w6394_
	);
	LUT2 #(
		.INIT('h1)
	) name5393 (
		_w6387_,
		_w6393_,
		_w6395_
	);
	LUT2 #(
		.INIT('h1)
	) name5394 (
		_w6394_,
		_w6395_,
		_w6396_
	);
	LUT2 #(
		.INIT('h8)
	) name5395 (
		_w6381_,
		_w6396_,
		_w6397_
	);
	LUT2 #(
		.INIT('h1)
	) name5396 (
		_w6388_,
		_w6391_,
		_w6398_
	);
	LUT2 #(
		.INIT('h1)
	) name5397 (
		_w6382_,
		_w6385_,
		_w6399_
	);
	LUT2 #(
		.INIT('h8)
	) name5398 (
		_w6398_,
		_w6399_,
		_w6400_
	);
	LUT2 #(
		.INIT('h1)
	) name5399 (
		_w6398_,
		_w6399_,
		_w6401_
	);
	LUT2 #(
		.INIT('h1)
	) name5400 (
		_w6400_,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h8)
	) name5401 (
		_w6397_,
		_w6402_,
		_w6403_
	);
	LUT2 #(
		.INIT('h1)
	) name5402 (
		_w6367_,
		_w6370_,
		_w6404_
	);
	LUT2 #(
		.INIT('h8)
	) name5403 (
		_w6373_,
		_w6379_,
		_w6405_
	);
	LUT2 #(
		.INIT('h1)
	) name5404 (
		_w6373_,
		_w6376_,
		_w6406_
	);
	LUT2 #(
		.INIT('h4)
	) name5405 (
		_w6379_,
		_w6406_,
		_w6407_
	);
	LUT2 #(
		.INIT('h1)
	) name5406 (
		_w6405_,
		_w6407_,
		_w6408_
	);
	LUT2 #(
		.INIT('h2)
	) name5407 (
		_w6404_,
		_w6408_,
		_w6409_
	);
	LUT2 #(
		.INIT('h4)
	) name5408 (
		_w6404_,
		_w6408_,
		_w6410_
	);
	LUT2 #(
		.INIT('h1)
	) name5409 (
		_w6409_,
		_w6410_,
		_w6411_
	);
	LUT2 #(
		.INIT('h1)
	) name5410 (
		_w6403_,
		_w6411_,
		_w6412_
	);
	LUT2 #(
		.INIT('h4)
	) name5411 (
		_w6394_,
		_w6402_,
		_w6413_
	);
	LUT2 #(
		.INIT('h2)
	) name5412 (
		_w6394_,
		_w6402_,
		_w6414_
	);
	LUT2 #(
		.INIT('h1)
	) name5413 (
		_w6397_,
		_w6413_,
		_w6415_
	);
	LUT2 #(
		.INIT('h4)
	) name5414 (
		_w6414_,
		_w6415_,
		_w6416_
	);
	LUT2 #(
		.INIT('h1)
	) name5415 (
		_w6412_,
		_w6416_,
		_w6417_
	);
	LUT2 #(
		.INIT('h2)
	) name5416 (
		_w6394_,
		_w6400_,
		_w6418_
	);
	LUT2 #(
		.INIT('h1)
	) name5417 (
		_w6401_,
		_w6418_,
		_w6419_
	);
	LUT2 #(
		.INIT('h2)
	) name5418 (
		_w6417_,
		_w6419_,
		_w6420_
	);
	LUT2 #(
		.INIT('h4)
	) name5419 (
		_w6417_,
		_w6419_,
		_w6421_
	);
	LUT2 #(
		.INIT('h1)
	) name5420 (
		_w6404_,
		_w6407_,
		_w6422_
	);
	LUT2 #(
		.INIT('h1)
	) name5421 (
		_w6405_,
		_w6422_,
		_w6423_
	);
	LUT2 #(
		.INIT('h1)
	) name5422 (
		_w6421_,
		_w6423_,
		_w6424_
	);
	LUT2 #(
		.INIT('h1)
	) name5423 (
		_w6420_,
		_w6424_,
		_w6425_
	);
	LUT2 #(
		.INIT('h1)
	) name5424 (
		_w6366_,
		_w6425_,
		_w6426_
	);
	LUT2 #(
		.INIT('h8)
	) name5425 (
		_w6366_,
		_w6425_,
		_w6427_
	);
	LUT2 #(
		.INIT('h1)
	) name5426 (
		_w6426_,
		_w6427_,
		_w6428_
	);
	LUT2 #(
		.INIT('h1)
	) name5427 (
		_w6420_,
		_w6421_,
		_w6429_
	);
	LUT2 #(
		.INIT('h4)
	) name5428 (
		_w6423_,
		_w6429_,
		_w6430_
	);
	LUT2 #(
		.INIT('h2)
	) name5429 (
		_w6423_,
		_w6429_,
		_w6431_
	);
	LUT2 #(
		.INIT('h1)
	) name5430 (
		_w6430_,
		_w6431_,
		_w6432_
	);
	LUT2 #(
		.INIT('h1)
	) name5431 (
		_w6361_,
		_w6362_,
		_w6433_
	);
	LUT2 #(
		.INIT('h4)
	) name5432 (
		_w6364_,
		_w6433_,
		_w6434_
	);
	LUT2 #(
		.INIT('h2)
	) name5433 (
		_w6364_,
		_w6433_,
		_w6435_
	);
	LUT2 #(
		.INIT('h1)
	) name5434 (
		_w6434_,
		_w6435_,
		_w6436_
	);
	LUT2 #(
		.INIT('h1)
	) name5435 (
		_w6432_,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('h8)
	) name5436 (
		_w6432_,
		_w6436_,
		_w6438_
	);
	LUT2 #(
		.INIT('h1)
	) name5437 (
		_w6322_,
		_w6337_,
		_w6439_
	);
	LUT2 #(
		.INIT('h1)
	) name5438 (
		_w6338_,
		_w6439_,
		_w6440_
	);
	LUT2 #(
		.INIT('h1)
	) name5439 (
		_w6381_,
		_w6396_,
		_w6441_
	);
	LUT2 #(
		.INIT('h1)
	) name5440 (
		_w6397_,
		_w6441_,
		_w6442_
	);
	LUT2 #(
		.INIT('h8)
	) name5441 (
		_w6440_,
		_w6442_,
		_w6443_
	);
	LUT2 #(
		.INIT('h1)
	) name5442 (
		_w6344_,
		_w6357_,
		_w6444_
	);
	LUT2 #(
		.INIT('h4)
	) name5443 (
		_w6352_,
		_w6444_,
		_w6445_
	);
	LUT2 #(
		.INIT('h2)
	) name5444 (
		_w6352_,
		_w6444_,
		_w6446_
	);
	LUT2 #(
		.INIT('h1)
	) name5445 (
		_w6445_,
		_w6446_,
		_w6447_
	);
	LUT2 #(
		.INIT('h2)
	) name5446 (
		_w6443_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h4)
	) name5447 (
		_w6443_,
		_w6447_,
		_w6449_
	);
	LUT2 #(
		.INIT('h1)
	) name5448 (
		_w6403_,
		_w6416_,
		_w6450_
	);
	LUT2 #(
		.INIT('h4)
	) name5449 (
		_w6411_,
		_w6450_,
		_w6451_
	);
	LUT2 #(
		.INIT('h2)
	) name5450 (
		_w6411_,
		_w6450_,
		_w6452_
	);
	LUT2 #(
		.INIT('h1)
	) name5451 (
		_w6451_,
		_w6452_,
		_w6453_
	);
	LUT2 #(
		.INIT('h1)
	) name5452 (
		_w6449_,
		_w6453_,
		_w6454_
	);
	LUT2 #(
		.INIT('h1)
	) name5453 (
		_w6448_,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('h4)
	) name5454 (
		_w6438_,
		_w6455_,
		_w6456_
	);
	LUT2 #(
		.INIT('h1)
	) name5455 (
		_w6437_,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h2)
	) name5456 (
		_w6428_,
		_w6457_,
		_w6458_
	);
	LUT2 #(
		.INIT('h4)
	) name5457 (
		_w6428_,
		_w6457_,
		_w6459_
	);
	LUT2 #(
		.INIT('h1)
	) name5458 (
		_w6458_,
		_w6459_,
		_w6460_
	);
	LUT2 #(
		.INIT('h8)
	) name5459 (
		\A[811] ,
		\A[812] ,
		_w6461_
	);
	LUT2 #(
		.INIT('h1)
	) name5460 (
		\A[811] ,
		\A[812] ,
		_w6462_
	);
	LUT2 #(
		.INIT('h1)
	) name5461 (
		_w6461_,
		_w6462_,
		_w6463_
	);
	LUT2 #(
		.INIT('h8)
	) name5462 (
		\A[813] ,
		_w6463_,
		_w6464_
	);
	LUT2 #(
		.INIT('h1)
	) name5463 (
		\A[813] ,
		_w6463_,
		_w6465_
	);
	LUT2 #(
		.INIT('h1)
	) name5464 (
		_w6464_,
		_w6465_,
		_w6466_
	);
	LUT2 #(
		.INIT('h8)
	) name5465 (
		\A[814] ,
		\A[815] ,
		_w6467_
	);
	LUT2 #(
		.INIT('h1)
	) name5466 (
		\A[814] ,
		\A[815] ,
		_w6468_
	);
	LUT2 #(
		.INIT('h1)
	) name5467 (
		_w6467_,
		_w6468_,
		_w6469_
	);
	LUT2 #(
		.INIT('h8)
	) name5468 (
		\A[816] ,
		_w6469_,
		_w6470_
	);
	LUT2 #(
		.INIT('h1)
	) name5469 (
		\A[816] ,
		_w6469_,
		_w6471_
	);
	LUT2 #(
		.INIT('h1)
	) name5470 (
		_w6470_,
		_w6471_,
		_w6472_
	);
	LUT2 #(
		.INIT('h8)
	) name5471 (
		_w6466_,
		_w6472_,
		_w6473_
	);
	LUT2 #(
		.INIT('h1)
	) name5472 (
		_w6466_,
		_w6472_,
		_w6474_
	);
	LUT2 #(
		.INIT('h1)
	) name5473 (
		_w6473_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h8)
	) name5474 (
		\A[817] ,
		\A[818] ,
		_w6476_
	);
	LUT2 #(
		.INIT('h1)
	) name5475 (
		\A[817] ,
		\A[818] ,
		_w6477_
	);
	LUT2 #(
		.INIT('h1)
	) name5476 (
		_w6476_,
		_w6477_,
		_w6478_
	);
	LUT2 #(
		.INIT('h8)
	) name5477 (
		\A[819] ,
		_w6478_,
		_w6479_
	);
	LUT2 #(
		.INIT('h1)
	) name5478 (
		\A[819] ,
		_w6478_,
		_w6480_
	);
	LUT2 #(
		.INIT('h1)
	) name5479 (
		_w6479_,
		_w6480_,
		_w6481_
	);
	LUT2 #(
		.INIT('h8)
	) name5480 (
		\A[820] ,
		\A[821] ,
		_w6482_
	);
	LUT2 #(
		.INIT('h1)
	) name5481 (
		\A[820] ,
		\A[821] ,
		_w6483_
	);
	LUT2 #(
		.INIT('h1)
	) name5482 (
		_w6482_,
		_w6483_,
		_w6484_
	);
	LUT2 #(
		.INIT('h8)
	) name5483 (
		\A[822] ,
		_w6484_,
		_w6485_
	);
	LUT2 #(
		.INIT('h1)
	) name5484 (
		\A[822] ,
		_w6484_,
		_w6486_
	);
	LUT2 #(
		.INIT('h1)
	) name5485 (
		_w6485_,
		_w6486_,
		_w6487_
	);
	LUT2 #(
		.INIT('h8)
	) name5486 (
		_w6481_,
		_w6487_,
		_w6488_
	);
	LUT2 #(
		.INIT('h1)
	) name5487 (
		_w6481_,
		_w6487_,
		_w6489_
	);
	LUT2 #(
		.INIT('h1)
	) name5488 (
		_w6488_,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('h8)
	) name5489 (
		_w6475_,
		_w6490_,
		_w6491_
	);
	LUT2 #(
		.INIT('h1)
	) name5490 (
		_w6482_,
		_w6485_,
		_w6492_
	);
	LUT2 #(
		.INIT('h1)
	) name5491 (
		_w6476_,
		_w6479_,
		_w6493_
	);
	LUT2 #(
		.INIT('h8)
	) name5492 (
		_w6492_,
		_w6493_,
		_w6494_
	);
	LUT2 #(
		.INIT('h1)
	) name5493 (
		_w6492_,
		_w6493_,
		_w6495_
	);
	LUT2 #(
		.INIT('h1)
	) name5494 (
		_w6494_,
		_w6495_,
		_w6496_
	);
	LUT2 #(
		.INIT('h8)
	) name5495 (
		_w6491_,
		_w6496_,
		_w6497_
	);
	LUT2 #(
		.INIT('h1)
	) name5496 (
		_w6461_,
		_w6464_,
		_w6498_
	);
	LUT2 #(
		.INIT('h8)
	) name5497 (
		_w6467_,
		_w6473_,
		_w6499_
	);
	LUT2 #(
		.INIT('h1)
	) name5498 (
		_w6467_,
		_w6470_,
		_w6500_
	);
	LUT2 #(
		.INIT('h4)
	) name5499 (
		_w6473_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h1)
	) name5500 (
		_w6499_,
		_w6501_,
		_w6502_
	);
	LUT2 #(
		.INIT('h2)
	) name5501 (
		_w6498_,
		_w6502_,
		_w6503_
	);
	LUT2 #(
		.INIT('h4)
	) name5502 (
		_w6498_,
		_w6502_,
		_w6504_
	);
	LUT2 #(
		.INIT('h1)
	) name5503 (
		_w6503_,
		_w6504_,
		_w6505_
	);
	LUT2 #(
		.INIT('h1)
	) name5504 (
		_w6497_,
		_w6505_,
		_w6506_
	);
	LUT2 #(
		.INIT('h4)
	) name5505 (
		_w6488_,
		_w6496_,
		_w6507_
	);
	LUT2 #(
		.INIT('h2)
	) name5506 (
		_w6488_,
		_w6496_,
		_w6508_
	);
	LUT2 #(
		.INIT('h1)
	) name5507 (
		_w6491_,
		_w6507_,
		_w6509_
	);
	LUT2 #(
		.INIT('h4)
	) name5508 (
		_w6508_,
		_w6509_,
		_w6510_
	);
	LUT2 #(
		.INIT('h1)
	) name5509 (
		_w6506_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('h2)
	) name5510 (
		_w6488_,
		_w6494_,
		_w6512_
	);
	LUT2 #(
		.INIT('h1)
	) name5511 (
		_w6495_,
		_w6512_,
		_w6513_
	);
	LUT2 #(
		.INIT('h2)
	) name5512 (
		_w6511_,
		_w6513_,
		_w6514_
	);
	LUT2 #(
		.INIT('h4)
	) name5513 (
		_w6511_,
		_w6513_,
		_w6515_
	);
	LUT2 #(
		.INIT('h1)
	) name5514 (
		_w6498_,
		_w6501_,
		_w6516_
	);
	LUT2 #(
		.INIT('h1)
	) name5515 (
		_w6499_,
		_w6516_,
		_w6517_
	);
	LUT2 #(
		.INIT('h1)
	) name5516 (
		_w6515_,
		_w6517_,
		_w6518_
	);
	LUT2 #(
		.INIT('h1)
	) name5517 (
		_w6514_,
		_w6518_,
		_w6519_
	);
	LUT2 #(
		.INIT('h8)
	) name5518 (
		\A[805] ,
		\A[806] ,
		_w6520_
	);
	LUT2 #(
		.INIT('h1)
	) name5519 (
		\A[805] ,
		\A[806] ,
		_w6521_
	);
	LUT2 #(
		.INIT('h1)
	) name5520 (
		_w6520_,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h8)
	) name5521 (
		\A[807] ,
		_w6522_,
		_w6523_
	);
	LUT2 #(
		.INIT('h1)
	) name5522 (
		\A[807] ,
		_w6522_,
		_w6524_
	);
	LUT2 #(
		.INIT('h1)
	) name5523 (
		_w6523_,
		_w6524_,
		_w6525_
	);
	LUT2 #(
		.INIT('h8)
	) name5524 (
		\A[808] ,
		\A[809] ,
		_w6526_
	);
	LUT2 #(
		.INIT('h1)
	) name5525 (
		\A[808] ,
		\A[809] ,
		_w6527_
	);
	LUT2 #(
		.INIT('h1)
	) name5526 (
		_w6526_,
		_w6527_,
		_w6528_
	);
	LUT2 #(
		.INIT('h8)
	) name5527 (
		\A[810] ,
		_w6528_,
		_w6529_
	);
	LUT2 #(
		.INIT('h1)
	) name5528 (
		\A[810] ,
		_w6528_,
		_w6530_
	);
	LUT2 #(
		.INIT('h1)
	) name5529 (
		_w6529_,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h8)
	) name5530 (
		_w6525_,
		_w6531_,
		_w6532_
	);
	LUT2 #(
		.INIT('h1)
	) name5531 (
		_w6525_,
		_w6531_,
		_w6533_
	);
	LUT2 #(
		.INIT('h1)
	) name5532 (
		_w6532_,
		_w6533_,
		_w6534_
	);
	LUT2 #(
		.INIT('h8)
	) name5533 (
		\A[799] ,
		\A[800] ,
		_w6535_
	);
	LUT2 #(
		.INIT('h1)
	) name5534 (
		\A[799] ,
		\A[800] ,
		_w6536_
	);
	LUT2 #(
		.INIT('h1)
	) name5535 (
		_w6535_,
		_w6536_,
		_w6537_
	);
	LUT2 #(
		.INIT('h8)
	) name5536 (
		\A[801] ,
		_w6537_,
		_w6538_
	);
	LUT2 #(
		.INIT('h1)
	) name5537 (
		\A[801] ,
		_w6537_,
		_w6539_
	);
	LUT2 #(
		.INIT('h1)
	) name5538 (
		_w6538_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h8)
	) name5539 (
		\A[802] ,
		\A[803] ,
		_w6541_
	);
	LUT2 #(
		.INIT('h1)
	) name5540 (
		\A[802] ,
		\A[803] ,
		_w6542_
	);
	LUT2 #(
		.INIT('h1)
	) name5541 (
		_w6541_,
		_w6542_,
		_w6543_
	);
	LUT2 #(
		.INIT('h8)
	) name5542 (
		\A[804] ,
		_w6543_,
		_w6544_
	);
	LUT2 #(
		.INIT('h1)
	) name5543 (
		\A[804] ,
		_w6543_,
		_w6545_
	);
	LUT2 #(
		.INIT('h1)
	) name5544 (
		_w6544_,
		_w6545_,
		_w6546_
	);
	LUT2 #(
		.INIT('h8)
	) name5545 (
		_w6540_,
		_w6546_,
		_w6547_
	);
	LUT2 #(
		.INIT('h1)
	) name5546 (
		_w6540_,
		_w6546_,
		_w6548_
	);
	LUT2 #(
		.INIT('h1)
	) name5547 (
		_w6547_,
		_w6548_,
		_w6549_
	);
	LUT2 #(
		.INIT('h8)
	) name5548 (
		_w6534_,
		_w6549_,
		_w6550_
	);
	LUT2 #(
		.INIT('h1)
	) name5549 (
		_w6526_,
		_w6529_,
		_w6551_
	);
	LUT2 #(
		.INIT('h1)
	) name5550 (
		_w6520_,
		_w6523_,
		_w6552_
	);
	LUT2 #(
		.INIT('h1)
	) name5551 (
		_w6551_,
		_w6552_,
		_w6553_
	);
	LUT2 #(
		.INIT('h8)
	) name5552 (
		_w6551_,
		_w6552_,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name5553 (
		_w6553_,
		_w6554_,
		_w6555_
	);
	LUT2 #(
		.INIT('h8)
	) name5554 (
		_w6550_,
		_w6555_,
		_w6556_
	);
	LUT2 #(
		.INIT('h1)
	) name5555 (
		_w6541_,
		_w6544_,
		_w6557_
	);
	LUT2 #(
		.INIT('h1)
	) name5556 (
		_w6535_,
		_w6538_,
		_w6558_
	);
	LUT2 #(
		.INIT('h1)
	) name5557 (
		_w6557_,
		_w6558_,
		_w6559_
	);
	LUT2 #(
		.INIT('h8)
	) name5558 (
		_w6557_,
		_w6558_,
		_w6560_
	);
	LUT2 #(
		.INIT('h1)
	) name5559 (
		_w6559_,
		_w6560_,
		_w6561_
	);
	LUT2 #(
		.INIT('h2)
	) name5560 (
		_w6547_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h4)
	) name5561 (
		_w6547_,
		_w6561_,
		_w6563_
	);
	LUT2 #(
		.INIT('h1)
	) name5562 (
		_w6562_,
		_w6563_,
		_w6564_
	);
	LUT2 #(
		.INIT('h4)
	) name5563 (
		_w6556_,
		_w6564_,
		_w6565_
	);
	LUT2 #(
		.INIT('h4)
	) name5564 (
		_w6532_,
		_w6555_,
		_w6566_
	);
	LUT2 #(
		.INIT('h2)
	) name5565 (
		_w6532_,
		_w6555_,
		_w6567_
	);
	LUT2 #(
		.INIT('h1)
	) name5566 (
		_w6550_,
		_w6566_,
		_w6568_
	);
	LUT2 #(
		.INIT('h4)
	) name5567 (
		_w6567_,
		_w6568_,
		_w6569_
	);
	LUT2 #(
		.INIT('h1)
	) name5568 (
		_w6565_,
		_w6569_,
		_w6570_
	);
	LUT2 #(
		.INIT('h1)
	) name5569 (
		_w6532_,
		_w6553_,
		_w6571_
	);
	LUT2 #(
		.INIT('h1)
	) name5570 (
		_w6554_,
		_w6571_,
		_w6572_
	);
	LUT2 #(
		.INIT('h1)
	) name5571 (
		_w6570_,
		_w6572_,
		_w6573_
	);
	LUT2 #(
		.INIT('h8)
	) name5572 (
		_w6570_,
		_w6572_,
		_w6574_
	);
	LUT2 #(
		.INIT('h1)
	) name5573 (
		_w6547_,
		_w6559_,
		_w6575_
	);
	LUT2 #(
		.INIT('h1)
	) name5574 (
		_w6560_,
		_w6575_,
		_w6576_
	);
	LUT2 #(
		.INIT('h1)
	) name5575 (
		_w6574_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h1)
	) name5576 (
		_w6573_,
		_w6577_,
		_w6578_
	);
	LUT2 #(
		.INIT('h4)
	) name5577 (
		_w6519_,
		_w6578_,
		_w6579_
	);
	LUT2 #(
		.INIT('h2)
	) name5578 (
		_w6519_,
		_w6578_,
		_w6580_
	);
	LUT2 #(
		.INIT('h1)
	) name5579 (
		_w6579_,
		_w6580_,
		_w6581_
	);
	LUT2 #(
		.INIT('h1)
	) name5580 (
		_w6573_,
		_w6574_,
		_w6582_
	);
	LUT2 #(
		.INIT('h4)
	) name5581 (
		_w6576_,
		_w6582_,
		_w6583_
	);
	LUT2 #(
		.INIT('h2)
	) name5582 (
		_w6576_,
		_w6582_,
		_w6584_
	);
	LUT2 #(
		.INIT('h1)
	) name5583 (
		_w6583_,
		_w6584_,
		_w6585_
	);
	LUT2 #(
		.INIT('h1)
	) name5584 (
		_w6514_,
		_w6515_,
		_w6586_
	);
	LUT2 #(
		.INIT('h4)
	) name5585 (
		_w6517_,
		_w6586_,
		_w6587_
	);
	LUT2 #(
		.INIT('h2)
	) name5586 (
		_w6517_,
		_w6586_,
		_w6588_
	);
	LUT2 #(
		.INIT('h1)
	) name5587 (
		_w6587_,
		_w6588_,
		_w6589_
	);
	LUT2 #(
		.INIT('h4)
	) name5588 (
		_w6585_,
		_w6589_,
		_w6590_
	);
	LUT2 #(
		.INIT('h2)
	) name5589 (
		_w6585_,
		_w6589_,
		_w6591_
	);
	LUT2 #(
		.INIT('h1)
	) name5590 (
		_w6475_,
		_w6490_,
		_w6592_
	);
	LUT2 #(
		.INIT('h1)
	) name5591 (
		_w6491_,
		_w6592_,
		_w6593_
	);
	LUT2 #(
		.INIT('h1)
	) name5592 (
		_w6534_,
		_w6549_,
		_w6594_
	);
	LUT2 #(
		.INIT('h1)
	) name5593 (
		_w6550_,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h8)
	) name5594 (
		_w6593_,
		_w6595_,
		_w6596_
	);
	LUT2 #(
		.INIT('h1)
	) name5595 (
		_w6497_,
		_w6510_,
		_w6597_
	);
	LUT2 #(
		.INIT('h4)
	) name5596 (
		_w6505_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h2)
	) name5597 (
		_w6505_,
		_w6597_,
		_w6599_
	);
	LUT2 #(
		.INIT('h1)
	) name5598 (
		_w6598_,
		_w6599_,
		_w6600_
	);
	LUT2 #(
		.INIT('h2)
	) name5599 (
		_w6596_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h4)
	) name5600 (
		_w6596_,
		_w6600_,
		_w6602_
	);
	LUT2 #(
		.INIT('h1)
	) name5601 (
		_w6556_,
		_w6569_,
		_w6603_
	);
	LUT2 #(
		.INIT('h8)
	) name5602 (
		_w6564_,
		_w6603_,
		_w6604_
	);
	LUT2 #(
		.INIT('h1)
	) name5603 (
		_w6564_,
		_w6603_,
		_w6605_
	);
	LUT2 #(
		.INIT('h1)
	) name5604 (
		_w6604_,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h1)
	) name5605 (
		_w6602_,
		_w6606_,
		_w6607_
	);
	LUT2 #(
		.INIT('h1)
	) name5606 (
		_w6601_,
		_w6607_,
		_w6608_
	);
	LUT2 #(
		.INIT('h1)
	) name5607 (
		_w6591_,
		_w6608_,
		_w6609_
	);
	LUT2 #(
		.INIT('h1)
	) name5608 (
		_w6590_,
		_w6609_,
		_w6610_
	);
	LUT2 #(
		.INIT('h2)
	) name5609 (
		_w6581_,
		_w6610_,
		_w6611_
	);
	LUT2 #(
		.INIT('h4)
	) name5610 (
		_w6581_,
		_w6610_,
		_w6612_
	);
	LUT2 #(
		.INIT('h1)
	) name5611 (
		_w6611_,
		_w6612_,
		_w6613_
	);
	LUT2 #(
		.INIT('h2)
	) name5612 (
		_w6460_,
		_w6613_,
		_w6614_
	);
	LUT2 #(
		.INIT('h4)
	) name5613 (
		_w6460_,
		_w6613_,
		_w6615_
	);
	LUT2 #(
		.INIT('h1)
	) name5614 (
		_w6590_,
		_w6591_,
		_w6616_
	);
	LUT2 #(
		.INIT('h4)
	) name5615 (
		_w6608_,
		_w6616_,
		_w6617_
	);
	LUT2 #(
		.INIT('h2)
	) name5616 (
		_w6608_,
		_w6616_,
		_w6618_
	);
	LUT2 #(
		.INIT('h1)
	) name5617 (
		_w6617_,
		_w6618_,
		_w6619_
	);
	LUT2 #(
		.INIT('h1)
	) name5618 (
		_w6437_,
		_w6438_,
		_w6620_
	);
	LUT2 #(
		.INIT('h4)
	) name5619 (
		_w6455_,
		_w6620_,
		_w6621_
	);
	LUT2 #(
		.INIT('h2)
	) name5620 (
		_w6455_,
		_w6620_,
		_w6622_
	);
	LUT2 #(
		.INIT('h1)
	) name5621 (
		_w6621_,
		_w6622_,
		_w6623_
	);
	LUT2 #(
		.INIT('h1)
	) name5622 (
		_w6619_,
		_w6623_,
		_w6624_
	);
	LUT2 #(
		.INIT('h8)
	) name5623 (
		_w6619_,
		_w6623_,
		_w6625_
	);
	LUT2 #(
		.INIT('h1)
	) name5624 (
		_w6440_,
		_w6442_,
		_w6626_
	);
	LUT2 #(
		.INIT('h1)
	) name5625 (
		_w6443_,
		_w6626_,
		_w6627_
	);
	LUT2 #(
		.INIT('h1)
	) name5626 (
		_w6593_,
		_w6595_,
		_w6628_
	);
	LUT2 #(
		.INIT('h1)
	) name5627 (
		_w6596_,
		_w6628_,
		_w6629_
	);
	LUT2 #(
		.INIT('h8)
	) name5628 (
		_w6627_,
		_w6629_,
		_w6630_
	);
	LUT2 #(
		.INIT('h1)
	) name5629 (
		_w6448_,
		_w6449_,
		_w6631_
	);
	LUT2 #(
		.INIT('h4)
	) name5630 (
		_w6453_,
		_w6631_,
		_w6632_
	);
	LUT2 #(
		.INIT('h2)
	) name5631 (
		_w6453_,
		_w6631_,
		_w6633_
	);
	LUT2 #(
		.INIT('h1)
	) name5632 (
		_w6632_,
		_w6633_,
		_w6634_
	);
	LUT2 #(
		.INIT('h8)
	) name5633 (
		_w6630_,
		_w6634_,
		_w6635_
	);
	LUT2 #(
		.INIT('h1)
	) name5634 (
		_w6630_,
		_w6634_,
		_w6636_
	);
	LUT2 #(
		.INIT('h1)
	) name5635 (
		_w6601_,
		_w6602_,
		_w6637_
	);
	LUT2 #(
		.INIT('h4)
	) name5636 (
		_w6606_,
		_w6637_,
		_w6638_
	);
	LUT2 #(
		.INIT('h2)
	) name5637 (
		_w6606_,
		_w6637_,
		_w6639_
	);
	LUT2 #(
		.INIT('h1)
	) name5638 (
		_w6638_,
		_w6639_,
		_w6640_
	);
	LUT2 #(
		.INIT('h4)
	) name5639 (
		_w6636_,
		_w6640_,
		_w6641_
	);
	LUT2 #(
		.INIT('h1)
	) name5640 (
		_w6635_,
		_w6641_,
		_w6642_
	);
	LUT2 #(
		.INIT('h4)
	) name5641 (
		_w6625_,
		_w6642_,
		_w6643_
	);
	LUT2 #(
		.INIT('h1)
	) name5642 (
		_w6624_,
		_w6643_,
		_w6644_
	);
	LUT2 #(
		.INIT('h1)
	) name5643 (
		_w6615_,
		_w6644_,
		_w6645_
	);
	LUT2 #(
		.INIT('h1)
	) name5644 (
		_w6614_,
		_w6645_,
		_w6646_
	);
	LUT2 #(
		.INIT('h4)
	) name5645 (
		_w6427_,
		_w6457_,
		_w6647_
	);
	LUT2 #(
		.INIT('h1)
	) name5646 (
		_w6426_,
		_w6647_,
		_w6648_
	);
	LUT2 #(
		.INIT('h2)
	) name5647 (
		_w6646_,
		_w6648_,
		_w6649_
	);
	LUT2 #(
		.INIT('h4)
	) name5648 (
		_w6646_,
		_w6648_,
		_w6650_
	);
	LUT2 #(
		.INIT('h1)
	) name5649 (
		_w6580_,
		_w6610_,
		_w6651_
	);
	LUT2 #(
		.INIT('h1)
	) name5650 (
		_w6579_,
		_w6651_,
		_w6652_
	);
	LUT2 #(
		.INIT('h1)
	) name5651 (
		_w6650_,
		_w6652_,
		_w6653_
	);
	LUT2 #(
		.INIT('h1)
	) name5652 (
		_w6649_,
		_w6653_,
		_w6654_
	);
	LUT2 #(
		.INIT('h8)
	) name5653 (
		\A[787] ,
		\A[788] ,
		_w6655_
	);
	LUT2 #(
		.INIT('h1)
	) name5654 (
		\A[787] ,
		\A[788] ,
		_w6656_
	);
	LUT2 #(
		.INIT('h1)
	) name5655 (
		_w6655_,
		_w6656_,
		_w6657_
	);
	LUT2 #(
		.INIT('h8)
	) name5656 (
		\A[789] ,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h1)
	) name5657 (
		\A[789] ,
		_w6657_,
		_w6659_
	);
	LUT2 #(
		.INIT('h1)
	) name5658 (
		_w6658_,
		_w6659_,
		_w6660_
	);
	LUT2 #(
		.INIT('h8)
	) name5659 (
		\A[790] ,
		\A[791] ,
		_w6661_
	);
	LUT2 #(
		.INIT('h1)
	) name5660 (
		\A[790] ,
		\A[791] ,
		_w6662_
	);
	LUT2 #(
		.INIT('h1)
	) name5661 (
		_w6661_,
		_w6662_,
		_w6663_
	);
	LUT2 #(
		.INIT('h8)
	) name5662 (
		\A[792] ,
		_w6663_,
		_w6664_
	);
	LUT2 #(
		.INIT('h1)
	) name5663 (
		\A[792] ,
		_w6663_,
		_w6665_
	);
	LUT2 #(
		.INIT('h1)
	) name5664 (
		_w6664_,
		_w6665_,
		_w6666_
	);
	LUT2 #(
		.INIT('h8)
	) name5665 (
		_w6660_,
		_w6666_,
		_w6667_
	);
	LUT2 #(
		.INIT('h1)
	) name5666 (
		_w6660_,
		_w6666_,
		_w6668_
	);
	LUT2 #(
		.INIT('h1)
	) name5667 (
		_w6667_,
		_w6668_,
		_w6669_
	);
	LUT2 #(
		.INIT('h8)
	) name5668 (
		\A[793] ,
		\A[794] ,
		_w6670_
	);
	LUT2 #(
		.INIT('h1)
	) name5669 (
		\A[793] ,
		\A[794] ,
		_w6671_
	);
	LUT2 #(
		.INIT('h1)
	) name5670 (
		_w6670_,
		_w6671_,
		_w6672_
	);
	LUT2 #(
		.INIT('h8)
	) name5671 (
		\A[795] ,
		_w6672_,
		_w6673_
	);
	LUT2 #(
		.INIT('h1)
	) name5672 (
		\A[795] ,
		_w6672_,
		_w6674_
	);
	LUT2 #(
		.INIT('h1)
	) name5673 (
		_w6673_,
		_w6674_,
		_w6675_
	);
	LUT2 #(
		.INIT('h8)
	) name5674 (
		\A[796] ,
		\A[797] ,
		_w6676_
	);
	LUT2 #(
		.INIT('h1)
	) name5675 (
		\A[796] ,
		\A[797] ,
		_w6677_
	);
	LUT2 #(
		.INIT('h1)
	) name5676 (
		_w6676_,
		_w6677_,
		_w6678_
	);
	LUT2 #(
		.INIT('h8)
	) name5677 (
		\A[798] ,
		_w6678_,
		_w6679_
	);
	LUT2 #(
		.INIT('h1)
	) name5678 (
		\A[798] ,
		_w6678_,
		_w6680_
	);
	LUT2 #(
		.INIT('h1)
	) name5679 (
		_w6679_,
		_w6680_,
		_w6681_
	);
	LUT2 #(
		.INIT('h8)
	) name5680 (
		_w6675_,
		_w6681_,
		_w6682_
	);
	LUT2 #(
		.INIT('h1)
	) name5681 (
		_w6675_,
		_w6681_,
		_w6683_
	);
	LUT2 #(
		.INIT('h1)
	) name5682 (
		_w6682_,
		_w6683_,
		_w6684_
	);
	LUT2 #(
		.INIT('h8)
	) name5683 (
		_w6669_,
		_w6684_,
		_w6685_
	);
	LUT2 #(
		.INIT('h1)
	) name5684 (
		_w6676_,
		_w6679_,
		_w6686_
	);
	LUT2 #(
		.INIT('h1)
	) name5685 (
		_w6670_,
		_w6673_,
		_w6687_
	);
	LUT2 #(
		.INIT('h8)
	) name5686 (
		_w6686_,
		_w6687_,
		_w6688_
	);
	LUT2 #(
		.INIT('h1)
	) name5687 (
		_w6686_,
		_w6687_,
		_w6689_
	);
	LUT2 #(
		.INIT('h1)
	) name5688 (
		_w6688_,
		_w6689_,
		_w6690_
	);
	LUT2 #(
		.INIT('h8)
	) name5689 (
		_w6685_,
		_w6690_,
		_w6691_
	);
	LUT2 #(
		.INIT('h1)
	) name5690 (
		_w6655_,
		_w6658_,
		_w6692_
	);
	LUT2 #(
		.INIT('h8)
	) name5691 (
		_w6661_,
		_w6667_,
		_w6693_
	);
	LUT2 #(
		.INIT('h1)
	) name5692 (
		_w6661_,
		_w6664_,
		_w6694_
	);
	LUT2 #(
		.INIT('h4)
	) name5693 (
		_w6667_,
		_w6694_,
		_w6695_
	);
	LUT2 #(
		.INIT('h1)
	) name5694 (
		_w6693_,
		_w6695_,
		_w6696_
	);
	LUT2 #(
		.INIT('h2)
	) name5695 (
		_w6692_,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h4)
	) name5696 (
		_w6692_,
		_w6696_,
		_w6698_
	);
	LUT2 #(
		.INIT('h1)
	) name5697 (
		_w6697_,
		_w6698_,
		_w6699_
	);
	LUT2 #(
		.INIT('h1)
	) name5698 (
		_w6691_,
		_w6699_,
		_w6700_
	);
	LUT2 #(
		.INIT('h4)
	) name5699 (
		_w6682_,
		_w6690_,
		_w6701_
	);
	LUT2 #(
		.INIT('h2)
	) name5700 (
		_w6682_,
		_w6690_,
		_w6702_
	);
	LUT2 #(
		.INIT('h1)
	) name5701 (
		_w6685_,
		_w6701_,
		_w6703_
	);
	LUT2 #(
		.INIT('h4)
	) name5702 (
		_w6702_,
		_w6703_,
		_w6704_
	);
	LUT2 #(
		.INIT('h1)
	) name5703 (
		_w6700_,
		_w6704_,
		_w6705_
	);
	LUT2 #(
		.INIT('h2)
	) name5704 (
		_w6682_,
		_w6688_,
		_w6706_
	);
	LUT2 #(
		.INIT('h1)
	) name5705 (
		_w6689_,
		_w6706_,
		_w6707_
	);
	LUT2 #(
		.INIT('h2)
	) name5706 (
		_w6705_,
		_w6707_,
		_w6708_
	);
	LUT2 #(
		.INIT('h4)
	) name5707 (
		_w6705_,
		_w6707_,
		_w6709_
	);
	LUT2 #(
		.INIT('h1)
	) name5708 (
		_w6692_,
		_w6695_,
		_w6710_
	);
	LUT2 #(
		.INIT('h1)
	) name5709 (
		_w6693_,
		_w6710_,
		_w6711_
	);
	LUT2 #(
		.INIT('h1)
	) name5710 (
		_w6709_,
		_w6711_,
		_w6712_
	);
	LUT2 #(
		.INIT('h1)
	) name5711 (
		_w6708_,
		_w6712_,
		_w6713_
	);
	LUT2 #(
		.INIT('h8)
	) name5712 (
		\A[775] ,
		\A[776] ,
		_w6714_
	);
	LUT2 #(
		.INIT('h1)
	) name5713 (
		\A[775] ,
		\A[776] ,
		_w6715_
	);
	LUT2 #(
		.INIT('h1)
	) name5714 (
		_w6714_,
		_w6715_,
		_w6716_
	);
	LUT2 #(
		.INIT('h8)
	) name5715 (
		\A[777] ,
		_w6716_,
		_w6717_
	);
	LUT2 #(
		.INIT('h1)
	) name5716 (
		\A[777] ,
		_w6716_,
		_w6718_
	);
	LUT2 #(
		.INIT('h1)
	) name5717 (
		_w6717_,
		_w6718_,
		_w6719_
	);
	LUT2 #(
		.INIT('h8)
	) name5718 (
		\A[778] ,
		\A[779] ,
		_w6720_
	);
	LUT2 #(
		.INIT('h1)
	) name5719 (
		\A[778] ,
		\A[779] ,
		_w6721_
	);
	LUT2 #(
		.INIT('h1)
	) name5720 (
		_w6720_,
		_w6721_,
		_w6722_
	);
	LUT2 #(
		.INIT('h8)
	) name5721 (
		\A[780] ,
		_w6722_,
		_w6723_
	);
	LUT2 #(
		.INIT('h1)
	) name5722 (
		\A[780] ,
		_w6722_,
		_w6724_
	);
	LUT2 #(
		.INIT('h1)
	) name5723 (
		_w6723_,
		_w6724_,
		_w6725_
	);
	LUT2 #(
		.INIT('h8)
	) name5724 (
		_w6719_,
		_w6725_,
		_w6726_
	);
	LUT2 #(
		.INIT('h1)
	) name5725 (
		_w6719_,
		_w6725_,
		_w6727_
	);
	LUT2 #(
		.INIT('h1)
	) name5726 (
		_w6726_,
		_w6727_,
		_w6728_
	);
	LUT2 #(
		.INIT('h8)
	) name5727 (
		\A[781] ,
		\A[782] ,
		_w6729_
	);
	LUT2 #(
		.INIT('h1)
	) name5728 (
		\A[781] ,
		\A[782] ,
		_w6730_
	);
	LUT2 #(
		.INIT('h1)
	) name5729 (
		_w6729_,
		_w6730_,
		_w6731_
	);
	LUT2 #(
		.INIT('h8)
	) name5730 (
		\A[783] ,
		_w6731_,
		_w6732_
	);
	LUT2 #(
		.INIT('h1)
	) name5731 (
		\A[783] ,
		_w6731_,
		_w6733_
	);
	LUT2 #(
		.INIT('h1)
	) name5732 (
		_w6732_,
		_w6733_,
		_w6734_
	);
	LUT2 #(
		.INIT('h8)
	) name5733 (
		\A[784] ,
		\A[785] ,
		_w6735_
	);
	LUT2 #(
		.INIT('h1)
	) name5734 (
		\A[784] ,
		\A[785] ,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name5735 (
		_w6735_,
		_w6736_,
		_w6737_
	);
	LUT2 #(
		.INIT('h8)
	) name5736 (
		\A[786] ,
		_w6737_,
		_w6738_
	);
	LUT2 #(
		.INIT('h1)
	) name5737 (
		\A[786] ,
		_w6737_,
		_w6739_
	);
	LUT2 #(
		.INIT('h1)
	) name5738 (
		_w6738_,
		_w6739_,
		_w6740_
	);
	LUT2 #(
		.INIT('h8)
	) name5739 (
		_w6734_,
		_w6740_,
		_w6741_
	);
	LUT2 #(
		.INIT('h1)
	) name5740 (
		_w6734_,
		_w6740_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name5741 (
		_w6741_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h8)
	) name5742 (
		_w6728_,
		_w6743_,
		_w6744_
	);
	LUT2 #(
		.INIT('h1)
	) name5743 (
		_w6735_,
		_w6738_,
		_w6745_
	);
	LUT2 #(
		.INIT('h1)
	) name5744 (
		_w6729_,
		_w6732_,
		_w6746_
	);
	LUT2 #(
		.INIT('h8)
	) name5745 (
		_w6745_,
		_w6746_,
		_w6747_
	);
	LUT2 #(
		.INIT('h1)
	) name5746 (
		_w6745_,
		_w6746_,
		_w6748_
	);
	LUT2 #(
		.INIT('h1)
	) name5747 (
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h8)
	) name5748 (
		_w6744_,
		_w6749_,
		_w6750_
	);
	LUT2 #(
		.INIT('h1)
	) name5749 (
		_w6714_,
		_w6717_,
		_w6751_
	);
	LUT2 #(
		.INIT('h8)
	) name5750 (
		_w6720_,
		_w6726_,
		_w6752_
	);
	LUT2 #(
		.INIT('h1)
	) name5751 (
		_w6720_,
		_w6723_,
		_w6753_
	);
	LUT2 #(
		.INIT('h4)
	) name5752 (
		_w6726_,
		_w6753_,
		_w6754_
	);
	LUT2 #(
		.INIT('h1)
	) name5753 (
		_w6752_,
		_w6754_,
		_w6755_
	);
	LUT2 #(
		.INIT('h2)
	) name5754 (
		_w6751_,
		_w6755_,
		_w6756_
	);
	LUT2 #(
		.INIT('h4)
	) name5755 (
		_w6751_,
		_w6755_,
		_w6757_
	);
	LUT2 #(
		.INIT('h1)
	) name5756 (
		_w6756_,
		_w6757_,
		_w6758_
	);
	LUT2 #(
		.INIT('h1)
	) name5757 (
		_w6750_,
		_w6758_,
		_w6759_
	);
	LUT2 #(
		.INIT('h4)
	) name5758 (
		_w6741_,
		_w6749_,
		_w6760_
	);
	LUT2 #(
		.INIT('h2)
	) name5759 (
		_w6741_,
		_w6749_,
		_w6761_
	);
	LUT2 #(
		.INIT('h1)
	) name5760 (
		_w6744_,
		_w6760_,
		_w6762_
	);
	LUT2 #(
		.INIT('h4)
	) name5761 (
		_w6761_,
		_w6762_,
		_w6763_
	);
	LUT2 #(
		.INIT('h1)
	) name5762 (
		_w6759_,
		_w6763_,
		_w6764_
	);
	LUT2 #(
		.INIT('h2)
	) name5763 (
		_w6741_,
		_w6747_,
		_w6765_
	);
	LUT2 #(
		.INIT('h1)
	) name5764 (
		_w6748_,
		_w6765_,
		_w6766_
	);
	LUT2 #(
		.INIT('h2)
	) name5765 (
		_w6764_,
		_w6766_,
		_w6767_
	);
	LUT2 #(
		.INIT('h4)
	) name5766 (
		_w6764_,
		_w6766_,
		_w6768_
	);
	LUT2 #(
		.INIT('h1)
	) name5767 (
		_w6751_,
		_w6754_,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name5768 (
		_w6752_,
		_w6769_,
		_w6770_
	);
	LUT2 #(
		.INIT('h1)
	) name5769 (
		_w6768_,
		_w6770_,
		_w6771_
	);
	LUT2 #(
		.INIT('h1)
	) name5770 (
		_w6767_,
		_w6771_,
		_w6772_
	);
	LUT2 #(
		.INIT('h1)
	) name5771 (
		_w6713_,
		_w6772_,
		_w6773_
	);
	LUT2 #(
		.INIT('h8)
	) name5772 (
		_w6713_,
		_w6772_,
		_w6774_
	);
	LUT2 #(
		.INIT('h1)
	) name5773 (
		_w6767_,
		_w6768_,
		_w6775_
	);
	LUT2 #(
		.INIT('h4)
	) name5774 (
		_w6770_,
		_w6775_,
		_w6776_
	);
	LUT2 #(
		.INIT('h2)
	) name5775 (
		_w6770_,
		_w6775_,
		_w6777_
	);
	LUT2 #(
		.INIT('h1)
	) name5776 (
		_w6776_,
		_w6777_,
		_w6778_
	);
	LUT2 #(
		.INIT('h1)
	) name5777 (
		_w6708_,
		_w6709_,
		_w6779_
	);
	LUT2 #(
		.INIT('h4)
	) name5778 (
		_w6711_,
		_w6779_,
		_w6780_
	);
	LUT2 #(
		.INIT('h2)
	) name5779 (
		_w6711_,
		_w6779_,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name5780 (
		_w6780_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h1)
	) name5781 (
		_w6778_,
		_w6782_,
		_w6783_
	);
	LUT2 #(
		.INIT('h8)
	) name5782 (
		_w6778_,
		_w6782_,
		_w6784_
	);
	LUT2 #(
		.INIT('h1)
	) name5783 (
		_w6669_,
		_w6684_,
		_w6785_
	);
	LUT2 #(
		.INIT('h1)
	) name5784 (
		_w6685_,
		_w6785_,
		_w6786_
	);
	LUT2 #(
		.INIT('h1)
	) name5785 (
		_w6728_,
		_w6743_,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name5786 (
		_w6744_,
		_w6787_,
		_w6788_
	);
	LUT2 #(
		.INIT('h8)
	) name5787 (
		_w6786_,
		_w6788_,
		_w6789_
	);
	LUT2 #(
		.INIT('h1)
	) name5788 (
		_w6691_,
		_w6704_,
		_w6790_
	);
	LUT2 #(
		.INIT('h4)
	) name5789 (
		_w6699_,
		_w6790_,
		_w6791_
	);
	LUT2 #(
		.INIT('h2)
	) name5790 (
		_w6699_,
		_w6790_,
		_w6792_
	);
	LUT2 #(
		.INIT('h1)
	) name5791 (
		_w6791_,
		_w6792_,
		_w6793_
	);
	LUT2 #(
		.INIT('h2)
	) name5792 (
		_w6789_,
		_w6793_,
		_w6794_
	);
	LUT2 #(
		.INIT('h4)
	) name5793 (
		_w6789_,
		_w6793_,
		_w6795_
	);
	LUT2 #(
		.INIT('h1)
	) name5794 (
		_w6750_,
		_w6763_,
		_w6796_
	);
	LUT2 #(
		.INIT('h4)
	) name5795 (
		_w6758_,
		_w6796_,
		_w6797_
	);
	LUT2 #(
		.INIT('h2)
	) name5796 (
		_w6758_,
		_w6796_,
		_w6798_
	);
	LUT2 #(
		.INIT('h1)
	) name5797 (
		_w6797_,
		_w6798_,
		_w6799_
	);
	LUT2 #(
		.INIT('h1)
	) name5798 (
		_w6795_,
		_w6799_,
		_w6800_
	);
	LUT2 #(
		.INIT('h1)
	) name5799 (
		_w6794_,
		_w6800_,
		_w6801_
	);
	LUT2 #(
		.INIT('h4)
	) name5800 (
		_w6784_,
		_w6801_,
		_w6802_
	);
	LUT2 #(
		.INIT('h1)
	) name5801 (
		_w6783_,
		_w6802_,
		_w6803_
	);
	LUT2 #(
		.INIT('h4)
	) name5802 (
		_w6774_,
		_w6803_,
		_w6804_
	);
	LUT2 #(
		.INIT('h1)
	) name5803 (
		_w6773_,
		_w6804_,
		_w6805_
	);
	LUT2 #(
		.INIT('h8)
	) name5804 (
		\A[757] ,
		\A[758] ,
		_w6806_
	);
	LUT2 #(
		.INIT('h1)
	) name5805 (
		\A[757] ,
		\A[758] ,
		_w6807_
	);
	LUT2 #(
		.INIT('h1)
	) name5806 (
		_w6806_,
		_w6807_,
		_w6808_
	);
	LUT2 #(
		.INIT('h8)
	) name5807 (
		\A[759] ,
		_w6808_,
		_w6809_
	);
	LUT2 #(
		.INIT('h1)
	) name5808 (
		\A[759] ,
		_w6808_,
		_w6810_
	);
	LUT2 #(
		.INIT('h1)
	) name5809 (
		_w6809_,
		_w6810_,
		_w6811_
	);
	LUT2 #(
		.INIT('h8)
	) name5810 (
		\A[760] ,
		\A[761] ,
		_w6812_
	);
	LUT2 #(
		.INIT('h1)
	) name5811 (
		\A[760] ,
		\A[761] ,
		_w6813_
	);
	LUT2 #(
		.INIT('h1)
	) name5812 (
		_w6812_,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h8)
	) name5813 (
		\A[762] ,
		_w6814_,
		_w6815_
	);
	LUT2 #(
		.INIT('h1)
	) name5814 (
		\A[762] ,
		_w6814_,
		_w6816_
	);
	LUT2 #(
		.INIT('h1)
	) name5815 (
		_w6815_,
		_w6816_,
		_w6817_
	);
	LUT2 #(
		.INIT('h8)
	) name5816 (
		_w6811_,
		_w6817_,
		_w6818_
	);
	LUT2 #(
		.INIT('h1)
	) name5817 (
		_w6811_,
		_w6817_,
		_w6819_
	);
	LUT2 #(
		.INIT('h1)
	) name5818 (
		_w6818_,
		_w6819_,
		_w6820_
	);
	LUT2 #(
		.INIT('h8)
	) name5819 (
		\A[751] ,
		\A[752] ,
		_w6821_
	);
	LUT2 #(
		.INIT('h1)
	) name5820 (
		\A[751] ,
		\A[752] ,
		_w6822_
	);
	LUT2 #(
		.INIT('h1)
	) name5821 (
		_w6821_,
		_w6822_,
		_w6823_
	);
	LUT2 #(
		.INIT('h8)
	) name5822 (
		\A[753] ,
		_w6823_,
		_w6824_
	);
	LUT2 #(
		.INIT('h1)
	) name5823 (
		\A[753] ,
		_w6823_,
		_w6825_
	);
	LUT2 #(
		.INIT('h1)
	) name5824 (
		_w6824_,
		_w6825_,
		_w6826_
	);
	LUT2 #(
		.INIT('h8)
	) name5825 (
		\A[754] ,
		\A[755] ,
		_w6827_
	);
	LUT2 #(
		.INIT('h1)
	) name5826 (
		\A[754] ,
		\A[755] ,
		_w6828_
	);
	LUT2 #(
		.INIT('h1)
	) name5827 (
		_w6827_,
		_w6828_,
		_w6829_
	);
	LUT2 #(
		.INIT('h8)
	) name5828 (
		\A[756] ,
		_w6829_,
		_w6830_
	);
	LUT2 #(
		.INIT('h1)
	) name5829 (
		\A[756] ,
		_w6829_,
		_w6831_
	);
	LUT2 #(
		.INIT('h1)
	) name5830 (
		_w6830_,
		_w6831_,
		_w6832_
	);
	LUT2 #(
		.INIT('h8)
	) name5831 (
		_w6826_,
		_w6832_,
		_w6833_
	);
	LUT2 #(
		.INIT('h1)
	) name5832 (
		_w6826_,
		_w6832_,
		_w6834_
	);
	LUT2 #(
		.INIT('h1)
	) name5833 (
		_w6833_,
		_w6834_,
		_w6835_
	);
	LUT2 #(
		.INIT('h8)
	) name5834 (
		_w6820_,
		_w6835_,
		_w6836_
	);
	LUT2 #(
		.INIT('h1)
	) name5835 (
		_w6812_,
		_w6815_,
		_w6837_
	);
	LUT2 #(
		.INIT('h1)
	) name5836 (
		_w6806_,
		_w6809_,
		_w6838_
	);
	LUT2 #(
		.INIT('h8)
	) name5837 (
		_w6837_,
		_w6838_,
		_w6839_
	);
	LUT2 #(
		.INIT('h1)
	) name5838 (
		_w6837_,
		_w6838_,
		_w6840_
	);
	LUT2 #(
		.INIT('h1)
	) name5839 (
		_w6839_,
		_w6840_,
		_w6841_
	);
	LUT2 #(
		.INIT('h8)
	) name5840 (
		_w6836_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h1)
	) name5841 (
		_w6827_,
		_w6830_,
		_w6843_
	);
	LUT2 #(
		.INIT('h1)
	) name5842 (
		_w6821_,
		_w6824_,
		_w6844_
	);
	LUT2 #(
		.INIT('h1)
	) name5843 (
		_w6843_,
		_w6844_,
		_w6845_
	);
	LUT2 #(
		.INIT('h8)
	) name5844 (
		_w6843_,
		_w6844_,
		_w6846_
	);
	LUT2 #(
		.INIT('h1)
	) name5845 (
		_w6845_,
		_w6846_,
		_w6847_
	);
	LUT2 #(
		.INIT('h2)
	) name5846 (
		_w6833_,
		_w6847_,
		_w6848_
	);
	LUT2 #(
		.INIT('h4)
	) name5847 (
		_w6833_,
		_w6847_,
		_w6849_
	);
	LUT2 #(
		.INIT('h1)
	) name5848 (
		_w6848_,
		_w6849_,
		_w6850_
	);
	LUT2 #(
		.INIT('h4)
	) name5849 (
		_w6842_,
		_w6850_,
		_w6851_
	);
	LUT2 #(
		.INIT('h4)
	) name5850 (
		_w6818_,
		_w6841_,
		_w6852_
	);
	LUT2 #(
		.INIT('h2)
	) name5851 (
		_w6818_,
		_w6841_,
		_w6853_
	);
	LUT2 #(
		.INIT('h1)
	) name5852 (
		_w6836_,
		_w6852_,
		_w6854_
	);
	LUT2 #(
		.INIT('h4)
	) name5853 (
		_w6853_,
		_w6854_,
		_w6855_
	);
	LUT2 #(
		.INIT('h1)
	) name5854 (
		_w6851_,
		_w6855_,
		_w6856_
	);
	LUT2 #(
		.INIT('h1)
	) name5855 (
		_w6833_,
		_w6845_,
		_w6857_
	);
	LUT2 #(
		.INIT('h1)
	) name5856 (
		_w6846_,
		_w6857_,
		_w6858_
	);
	LUT2 #(
		.INIT('h8)
	) name5857 (
		_w6856_,
		_w6858_,
		_w6859_
	);
	LUT2 #(
		.INIT('h1)
	) name5858 (
		_w6856_,
		_w6858_,
		_w6860_
	);
	LUT2 #(
		.INIT('h1)
	) name5859 (
		_w6859_,
		_w6860_,
		_w6861_
	);
	LUT2 #(
		.INIT('h1)
	) name5860 (
		_w6818_,
		_w6840_,
		_w6862_
	);
	LUT2 #(
		.INIT('h1)
	) name5861 (
		_w6839_,
		_w6862_,
		_w6863_
	);
	LUT2 #(
		.INIT('h2)
	) name5862 (
		_w6861_,
		_w6863_,
		_w6864_
	);
	LUT2 #(
		.INIT('h4)
	) name5863 (
		_w6861_,
		_w6863_,
		_w6865_
	);
	LUT2 #(
		.INIT('h1)
	) name5864 (
		_w6864_,
		_w6865_,
		_w6866_
	);
	LUT2 #(
		.INIT('h8)
	) name5865 (
		\A[766] ,
		\A[767] ,
		_w6867_
	);
	LUT2 #(
		.INIT('h8)
	) name5866 (
		\A[763] ,
		\A[764] ,
		_w6868_
	);
	LUT2 #(
		.INIT('h1)
	) name5867 (
		\A[763] ,
		\A[764] ,
		_w6869_
	);
	LUT2 #(
		.INIT('h1)
	) name5868 (
		_w6868_,
		_w6869_,
		_w6870_
	);
	LUT2 #(
		.INIT('h8)
	) name5869 (
		\A[765] ,
		_w6870_,
		_w6871_
	);
	LUT2 #(
		.INIT('h1)
	) name5870 (
		\A[765] ,
		_w6870_,
		_w6872_
	);
	LUT2 #(
		.INIT('h1)
	) name5871 (
		_w6871_,
		_w6872_,
		_w6873_
	);
	LUT2 #(
		.INIT('h1)
	) name5872 (
		\A[766] ,
		\A[767] ,
		_w6874_
	);
	LUT2 #(
		.INIT('h1)
	) name5873 (
		_w6867_,
		_w6874_,
		_w6875_
	);
	LUT2 #(
		.INIT('h8)
	) name5874 (
		\A[768] ,
		_w6875_,
		_w6876_
	);
	LUT2 #(
		.INIT('h1)
	) name5875 (
		\A[768] ,
		_w6875_,
		_w6877_
	);
	LUT2 #(
		.INIT('h1)
	) name5876 (
		_w6876_,
		_w6877_,
		_w6878_
	);
	LUT2 #(
		.INIT('h8)
	) name5877 (
		_w6873_,
		_w6878_,
		_w6879_
	);
	LUT2 #(
		.INIT('h8)
	) name5878 (
		_w6867_,
		_w6879_,
		_w6880_
	);
	LUT2 #(
		.INIT('h1)
	) name5879 (
		_w6868_,
		_w6871_,
		_w6881_
	);
	LUT2 #(
		.INIT('h1)
	) name5880 (
		_w6867_,
		_w6876_,
		_w6882_
	);
	LUT2 #(
		.INIT('h4)
	) name5881 (
		_w6879_,
		_w6882_,
		_w6883_
	);
	LUT2 #(
		.INIT('h1)
	) name5882 (
		_w6881_,
		_w6883_,
		_w6884_
	);
	LUT2 #(
		.INIT('h1)
	) name5883 (
		_w6880_,
		_w6884_,
		_w6885_
	);
	LUT2 #(
		.INIT('h8)
	) name5884 (
		\A[772] ,
		\A[773] ,
		_w6886_
	);
	LUT2 #(
		.INIT('h1)
	) name5885 (
		\A[772] ,
		\A[773] ,
		_w6887_
	);
	LUT2 #(
		.INIT('h1)
	) name5886 (
		_w6886_,
		_w6887_,
		_w6888_
	);
	LUT2 #(
		.INIT('h8)
	) name5887 (
		\A[774] ,
		_w6888_,
		_w6889_
	);
	LUT2 #(
		.INIT('h1)
	) name5888 (
		_w6886_,
		_w6889_,
		_w6890_
	);
	LUT2 #(
		.INIT('h8)
	) name5889 (
		\A[769] ,
		\A[770] ,
		_w6891_
	);
	LUT2 #(
		.INIT('h1)
	) name5890 (
		\A[769] ,
		\A[770] ,
		_w6892_
	);
	LUT2 #(
		.INIT('h1)
	) name5891 (
		_w6891_,
		_w6892_,
		_w6893_
	);
	LUT2 #(
		.INIT('h8)
	) name5892 (
		\A[771] ,
		_w6893_,
		_w6894_
	);
	LUT2 #(
		.INIT('h1)
	) name5893 (
		_w6891_,
		_w6894_,
		_w6895_
	);
	LUT2 #(
		.INIT('h8)
	) name5894 (
		_w6890_,
		_w6895_,
		_w6896_
	);
	LUT2 #(
		.INIT('h1)
	) name5895 (
		_w6890_,
		_w6895_,
		_w6897_
	);
	LUT2 #(
		.INIT('h1)
	) name5896 (
		\A[771] ,
		_w6893_,
		_w6898_
	);
	LUT2 #(
		.INIT('h1)
	) name5897 (
		_w6894_,
		_w6898_,
		_w6899_
	);
	LUT2 #(
		.INIT('h1)
	) name5898 (
		\A[774] ,
		_w6888_,
		_w6900_
	);
	LUT2 #(
		.INIT('h1)
	) name5899 (
		_w6889_,
		_w6900_,
		_w6901_
	);
	LUT2 #(
		.INIT('h8)
	) name5900 (
		_w6899_,
		_w6901_,
		_w6902_
	);
	LUT2 #(
		.INIT('h1)
	) name5901 (
		_w6897_,
		_w6902_,
		_w6903_
	);
	LUT2 #(
		.INIT('h1)
	) name5902 (
		_w6896_,
		_w6903_,
		_w6904_
	);
	LUT2 #(
		.INIT('h1)
	) name5903 (
		_w6899_,
		_w6901_,
		_w6905_
	);
	LUT2 #(
		.INIT('h1)
	) name5904 (
		_w6902_,
		_w6905_,
		_w6906_
	);
	LUT2 #(
		.INIT('h1)
	) name5905 (
		_w6873_,
		_w6878_,
		_w6907_
	);
	LUT2 #(
		.INIT('h1)
	) name5906 (
		_w6879_,
		_w6907_,
		_w6908_
	);
	LUT2 #(
		.INIT('h8)
	) name5907 (
		_w6906_,
		_w6908_,
		_w6909_
	);
	LUT2 #(
		.INIT('h2)
	) name5908 (
		_w6880_,
		_w6881_,
		_w6910_
	);
	LUT2 #(
		.INIT('h2)
	) name5909 (
		_w6909_,
		_w6910_,
		_w6911_
	);
	LUT2 #(
		.INIT('h1)
	) name5910 (
		_w6896_,
		_w6897_,
		_w6912_
	);
	LUT2 #(
		.INIT('h2)
	) name5911 (
		_w6902_,
		_w6912_,
		_w6913_
	);
	LUT2 #(
		.INIT('h4)
	) name5912 (
		_w6902_,
		_w6912_,
		_w6914_
	);
	LUT2 #(
		.INIT('h1)
	) name5913 (
		_w6913_,
		_w6914_,
		_w6915_
	);
	LUT2 #(
		.INIT('h2)
	) name5914 (
		_w6911_,
		_w6915_,
		_w6916_
	);
	LUT2 #(
		.INIT('h4)
	) name5915 (
		_w6911_,
		_w6915_,
		_w6917_
	);
	LUT2 #(
		.INIT('h1)
	) name5916 (
		_w6880_,
		_w6883_,
		_w6918_
	);
	LUT2 #(
		.INIT('h2)
	) name5917 (
		_w6881_,
		_w6918_,
		_w6919_
	);
	LUT2 #(
		.INIT('h4)
	) name5918 (
		_w6881_,
		_w6918_,
		_w6920_
	);
	LUT2 #(
		.INIT('h1)
	) name5919 (
		_w6919_,
		_w6920_,
		_w6921_
	);
	LUT2 #(
		.INIT('h4)
	) name5920 (
		_w6917_,
		_w6921_,
		_w6922_
	);
	LUT2 #(
		.INIT('h1)
	) name5921 (
		_w6916_,
		_w6922_,
		_w6923_
	);
	LUT2 #(
		.INIT('h2)
	) name5922 (
		_w6904_,
		_w6923_,
		_w6924_
	);
	LUT2 #(
		.INIT('h4)
	) name5923 (
		_w6904_,
		_w6923_,
		_w6925_
	);
	LUT2 #(
		.INIT('h1)
	) name5924 (
		_w6924_,
		_w6925_,
		_w6926_
	);
	LUT2 #(
		.INIT('h8)
	) name5925 (
		_w6885_,
		_w6926_,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name5926 (
		_w6885_,
		_w6926_,
		_w6928_
	);
	LUT2 #(
		.INIT('h1)
	) name5927 (
		_w6927_,
		_w6928_,
		_w6929_
	);
	LUT2 #(
		.INIT('h1)
	) name5928 (
		_w6866_,
		_w6929_,
		_w6930_
	);
	LUT2 #(
		.INIT('h8)
	) name5929 (
		_w6866_,
		_w6929_,
		_w6931_
	);
	LUT2 #(
		.INIT('h1)
	) name5930 (
		_w6906_,
		_w6908_,
		_w6932_
	);
	LUT2 #(
		.INIT('h1)
	) name5931 (
		_w6909_,
		_w6932_,
		_w6933_
	);
	LUT2 #(
		.INIT('h1)
	) name5932 (
		_w6820_,
		_w6835_,
		_w6934_
	);
	LUT2 #(
		.INIT('h1)
	) name5933 (
		_w6836_,
		_w6934_,
		_w6935_
	);
	LUT2 #(
		.INIT('h8)
	) name5934 (
		_w6933_,
		_w6935_,
		_w6936_
	);
	LUT2 #(
		.INIT('h1)
	) name5935 (
		_w6916_,
		_w6917_,
		_w6937_
	);
	LUT2 #(
		.INIT('h8)
	) name5936 (
		_w6921_,
		_w6937_,
		_w6938_
	);
	LUT2 #(
		.INIT('h1)
	) name5937 (
		_w6921_,
		_w6937_,
		_w6939_
	);
	LUT2 #(
		.INIT('h1)
	) name5938 (
		_w6938_,
		_w6939_,
		_w6940_
	);
	LUT2 #(
		.INIT('h8)
	) name5939 (
		_w6936_,
		_w6940_,
		_w6941_
	);
	LUT2 #(
		.INIT('h1)
	) name5940 (
		_w6936_,
		_w6940_,
		_w6942_
	);
	LUT2 #(
		.INIT('h1)
	) name5941 (
		_w6842_,
		_w6855_,
		_w6943_
	);
	LUT2 #(
		.INIT('h8)
	) name5942 (
		_w6850_,
		_w6943_,
		_w6944_
	);
	LUT2 #(
		.INIT('h1)
	) name5943 (
		_w6850_,
		_w6943_,
		_w6945_
	);
	LUT2 #(
		.INIT('h1)
	) name5944 (
		_w6944_,
		_w6945_,
		_w6946_
	);
	LUT2 #(
		.INIT('h1)
	) name5945 (
		_w6942_,
		_w6946_,
		_w6947_
	);
	LUT2 #(
		.INIT('h1)
	) name5946 (
		_w6941_,
		_w6947_,
		_w6948_
	);
	LUT2 #(
		.INIT('h1)
	) name5947 (
		_w6931_,
		_w6948_,
		_w6949_
	);
	LUT2 #(
		.INIT('h1)
	) name5948 (
		_w6930_,
		_w6949_,
		_w6950_
	);
	LUT2 #(
		.INIT('h1)
	) name5949 (
		_w6885_,
		_w6925_,
		_w6951_
	);
	LUT2 #(
		.INIT('h1)
	) name5950 (
		_w6924_,
		_w6951_,
		_w6952_
	);
	LUT2 #(
		.INIT('h8)
	) name5951 (
		_w6950_,
		_w6952_,
		_w6953_
	);
	LUT2 #(
		.INIT('h1)
	) name5952 (
		_w6950_,
		_w6952_,
		_w6954_
	);
	LUT2 #(
		.INIT('h1)
	) name5953 (
		_w6859_,
		_w6863_,
		_w6955_
	);
	LUT2 #(
		.INIT('h1)
	) name5954 (
		_w6860_,
		_w6955_,
		_w6956_
	);
	LUT2 #(
		.INIT('h1)
	) name5955 (
		_w6954_,
		_w6956_,
		_w6957_
	);
	LUT2 #(
		.INIT('h1)
	) name5956 (
		_w6953_,
		_w6957_,
		_w6958_
	);
	LUT2 #(
		.INIT('h4)
	) name5957 (
		_w6805_,
		_w6958_,
		_w6959_
	);
	LUT2 #(
		.INIT('h2)
	) name5958 (
		_w6805_,
		_w6958_,
		_w6960_
	);
	LUT2 #(
		.INIT('h1)
	) name5959 (
		_w6773_,
		_w6774_,
		_w6961_
	);
	LUT2 #(
		.INIT('h4)
	) name5960 (
		_w6803_,
		_w6961_,
		_w6962_
	);
	LUT2 #(
		.INIT('h2)
	) name5961 (
		_w6803_,
		_w6961_,
		_w6963_
	);
	LUT2 #(
		.INIT('h1)
	) name5962 (
		_w6962_,
		_w6963_,
		_w6964_
	);
	LUT2 #(
		.INIT('h1)
	) name5963 (
		_w6953_,
		_w6954_,
		_w6965_
	);
	LUT2 #(
		.INIT('h4)
	) name5964 (
		_w6956_,
		_w6965_,
		_w6966_
	);
	LUT2 #(
		.INIT('h2)
	) name5965 (
		_w6956_,
		_w6965_,
		_w6967_
	);
	LUT2 #(
		.INIT('h1)
	) name5966 (
		_w6966_,
		_w6967_,
		_w6968_
	);
	LUT2 #(
		.INIT('h1)
	) name5967 (
		_w6964_,
		_w6968_,
		_w6969_
	);
	LUT2 #(
		.INIT('h8)
	) name5968 (
		_w6964_,
		_w6968_,
		_w6970_
	);
	LUT2 #(
		.INIT('h1)
	) name5969 (
		_w6930_,
		_w6931_,
		_w6971_
	);
	LUT2 #(
		.INIT('h4)
	) name5970 (
		_w6948_,
		_w6971_,
		_w6972_
	);
	LUT2 #(
		.INIT('h2)
	) name5971 (
		_w6948_,
		_w6971_,
		_w6973_
	);
	LUT2 #(
		.INIT('h1)
	) name5972 (
		_w6972_,
		_w6973_,
		_w6974_
	);
	LUT2 #(
		.INIT('h1)
	) name5973 (
		_w6783_,
		_w6784_,
		_w6975_
	);
	LUT2 #(
		.INIT('h4)
	) name5974 (
		_w6801_,
		_w6975_,
		_w6976_
	);
	LUT2 #(
		.INIT('h2)
	) name5975 (
		_w6801_,
		_w6975_,
		_w6977_
	);
	LUT2 #(
		.INIT('h1)
	) name5976 (
		_w6976_,
		_w6977_,
		_w6978_
	);
	LUT2 #(
		.INIT('h1)
	) name5977 (
		_w6974_,
		_w6978_,
		_w6979_
	);
	LUT2 #(
		.INIT('h8)
	) name5978 (
		_w6974_,
		_w6978_,
		_w6980_
	);
	LUT2 #(
		.INIT('h1)
	) name5979 (
		_w6786_,
		_w6788_,
		_w6981_
	);
	LUT2 #(
		.INIT('h1)
	) name5980 (
		_w6789_,
		_w6981_,
		_w6982_
	);
	LUT2 #(
		.INIT('h1)
	) name5981 (
		_w6933_,
		_w6935_,
		_w6983_
	);
	LUT2 #(
		.INIT('h1)
	) name5982 (
		_w6936_,
		_w6983_,
		_w6984_
	);
	LUT2 #(
		.INIT('h8)
	) name5983 (
		_w6982_,
		_w6984_,
		_w6985_
	);
	LUT2 #(
		.INIT('h1)
	) name5984 (
		_w6794_,
		_w6795_,
		_w6986_
	);
	LUT2 #(
		.INIT('h4)
	) name5985 (
		_w6799_,
		_w6986_,
		_w6987_
	);
	LUT2 #(
		.INIT('h2)
	) name5986 (
		_w6799_,
		_w6986_,
		_w6988_
	);
	LUT2 #(
		.INIT('h1)
	) name5987 (
		_w6987_,
		_w6988_,
		_w6989_
	);
	LUT2 #(
		.INIT('h8)
	) name5988 (
		_w6985_,
		_w6989_,
		_w6990_
	);
	LUT2 #(
		.INIT('h1)
	) name5989 (
		_w6985_,
		_w6989_,
		_w6991_
	);
	LUT2 #(
		.INIT('h1)
	) name5990 (
		_w6941_,
		_w6942_,
		_w6992_
	);
	LUT2 #(
		.INIT('h4)
	) name5991 (
		_w6946_,
		_w6992_,
		_w6993_
	);
	LUT2 #(
		.INIT('h2)
	) name5992 (
		_w6946_,
		_w6992_,
		_w6994_
	);
	LUT2 #(
		.INIT('h1)
	) name5993 (
		_w6993_,
		_w6994_,
		_w6995_
	);
	LUT2 #(
		.INIT('h4)
	) name5994 (
		_w6991_,
		_w6995_,
		_w6996_
	);
	LUT2 #(
		.INIT('h1)
	) name5995 (
		_w6990_,
		_w6996_,
		_w6997_
	);
	LUT2 #(
		.INIT('h4)
	) name5996 (
		_w6980_,
		_w6997_,
		_w6998_
	);
	LUT2 #(
		.INIT('h1)
	) name5997 (
		_w6979_,
		_w6998_,
		_w6999_
	);
	LUT2 #(
		.INIT('h4)
	) name5998 (
		_w6970_,
		_w6999_,
		_w7000_
	);
	LUT2 #(
		.INIT('h1)
	) name5999 (
		_w6969_,
		_w7000_,
		_w7001_
	);
	LUT2 #(
		.INIT('h1)
	) name6000 (
		_w6960_,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('h1)
	) name6001 (
		_w6959_,
		_w7002_,
		_w7003_
	);
	LUT2 #(
		.INIT('h1)
	) name6002 (
		_w6654_,
		_w7003_,
		_w7004_
	);
	LUT2 #(
		.INIT('h8)
	) name6003 (
		_w6654_,
		_w7003_,
		_w7005_
	);
	LUT2 #(
		.INIT('h1)
	) name6004 (
		_w6959_,
		_w6960_,
		_w7006_
	);
	LUT2 #(
		.INIT('h4)
	) name6005 (
		_w7001_,
		_w7006_,
		_w7007_
	);
	LUT2 #(
		.INIT('h2)
	) name6006 (
		_w7001_,
		_w7006_,
		_w7008_
	);
	LUT2 #(
		.INIT('h1)
	) name6007 (
		_w7007_,
		_w7008_,
		_w7009_
	);
	LUT2 #(
		.INIT('h1)
	) name6008 (
		_w6649_,
		_w6650_,
		_w7010_
	);
	LUT2 #(
		.INIT('h8)
	) name6009 (
		_w6652_,
		_w7010_,
		_w7011_
	);
	LUT2 #(
		.INIT('h1)
	) name6010 (
		_w6652_,
		_w7010_,
		_w7012_
	);
	LUT2 #(
		.INIT('h1)
	) name6011 (
		_w7011_,
		_w7012_,
		_w7013_
	);
	LUT2 #(
		.INIT('h2)
	) name6012 (
		_w7009_,
		_w7013_,
		_w7014_
	);
	LUT2 #(
		.INIT('h4)
	) name6013 (
		_w7009_,
		_w7013_,
		_w7015_
	);
	LUT2 #(
		.INIT('h1)
	) name6014 (
		_w6614_,
		_w6615_,
		_w7016_
	);
	LUT2 #(
		.INIT('h4)
	) name6015 (
		_w6644_,
		_w7016_,
		_w7017_
	);
	LUT2 #(
		.INIT('h2)
	) name6016 (
		_w6644_,
		_w7016_,
		_w7018_
	);
	LUT2 #(
		.INIT('h1)
	) name6017 (
		_w7017_,
		_w7018_,
		_w7019_
	);
	LUT2 #(
		.INIT('h1)
	) name6018 (
		_w6969_,
		_w6970_,
		_w7020_
	);
	LUT2 #(
		.INIT('h8)
	) name6019 (
		_w6999_,
		_w7020_,
		_w7021_
	);
	LUT2 #(
		.INIT('h1)
	) name6020 (
		_w6999_,
		_w7020_,
		_w7022_
	);
	LUT2 #(
		.INIT('h1)
	) name6021 (
		_w7021_,
		_w7022_,
		_w7023_
	);
	LUT2 #(
		.INIT('h2)
	) name6022 (
		_w7019_,
		_w7023_,
		_w7024_
	);
	LUT2 #(
		.INIT('h4)
	) name6023 (
		_w7019_,
		_w7023_,
		_w7025_
	);
	LUT2 #(
		.INIT('h1)
	) name6024 (
		_w6979_,
		_w6980_,
		_w7026_
	);
	LUT2 #(
		.INIT('h4)
	) name6025 (
		_w6997_,
		_w7026_,
		_w7027_
	);
	LUT2 #(
		.INIT('h2)
	) name6026 (
		_w6997_,
		_w7026_,
		_w7028_
	);
	LUT2 #(
		.INIT('h1)
	) name6027 (
		_w7027_,
		_w7028_,
		_w7029_
	);
	LUT2 #(
		.INIT('h1)
	) name6028 (
		_w6624_,
		_w6625_,
		_w7030_
	);
	LUT2 #(
		.INIT('h4)
	) name6029 (
		_w6642_,
		_w7030_,
		_w7031_
	);
	LUT2 #(
		.INIT('h2)
	) name6030 (
		_w6642_,
		_w7030_,
		_w7032_
	);
	LUT2 #(
		.INIT('h1)
	) name6031 (
		_w7031_,
		_w7032_,
		_w7033_
	);
	LUT2 #(
		.INIT('h1)
	) name6032 (
		_w7029_,
		_w7033_,
		_w7034_
	);
	LUT2 #(
		.INIT('h8)
	) name6033 (
		_w7029_,
		_w7033_,
		_w7035_
	);
	LUT2 #(
		.INIT('h1)
	) name6034 (
		_w6627_,
		_w6629_,
		_w7036_
	);
	LUT2 #(
		.INIT('h1)
	) name6035 (
		_w6630_,
		_w7036_,
		_w7037_
	);
	LUT2 #(
		.INIT('h1)
	) name6036 (
		_w6982_,
		_w6984_,
		_w7038_
	);
	LUT2 #(
		.INIT('h1)
	) name6037 (
		_w6985_,
		_w7038_,
		_w7039_
	);
	LUT2 #(
		.INIT('h8)
	) name6038 (
		_w7037_,
		_w7039_,
		_w7040_
	);
	LUT2 #(
		.INIT('h1)
	) name6039 (
		_w6635_,
		_w6636_,
		_w7041_
	);
	LUT2 #(
		.INIT('h4)
	) name6040 (
		_w6640_,
		_w7041_,
		_w7042_
	);
	LUT2 #(
		.INIT('h2)
	) name6041 (
		_w6640_,
		_w7041_,
		_w7043_
	);
	LUT2 #(
		.INIT('h1)
	) name6042 (
		_w7042_,
		_w7043_,
		_w7044_
	);
	LUT2 #(
		.INIT('h2)
	) name6043 (
		_w7040_,
		_w7044_,
		_w7045_
	);
	LUT2 #(
		.INIT('h4)
	) name6044 (
		_w7040_,
		_w7044_,
		_w7046_
	);
	LUT2 #(
		.INIT('h1)
	) name6045 (
		_w6990_,
		_w6991_,
		_w7047_
	);
	LUT2 #(
		.INIT('h4)
	) name6046 (
		_w6995_,
		_w7047_,
		_w7048_
	);
	LUT2 #(
		.INIT('h2)
	) name6047 (
		_w6995_,
		_w7047_,
		_w7049_
	);
	LUT2 #(
		.INIT('h1)
	) name6048 (
		_w7048_,
		_w7049_,
		_w7050_
	);
	LUT2 #(
		.INIT('h1)
	) name6049 (
		_w7046_,
		_w7050_,
		_w7051_
	);
	LUT2 #(
		.INIT('h1)
	) name6050 (
		_w7045_,
		_w7051_,
		_w7052_
	);
	LUT2 #(
		.INIT('h4)
	) name6051 (
		_w7035_,
		_w7052_,
		_w7053_
	);
	LUT2 #(
		.INIT('h1)
	) name6052 (
		_w7034_,
		_w7053_,
		_w7054_
	);
	LUT2 #(
		.INIT('h1)
	) name6053 (
		_w7025_,
		_w7054_,
		_w7055_
	);
	LUT2 #(
		.INIT('h1)
	) name6054 (
		_w7024_,
		_w7055_,
		_w7056_
	);
	LUT2 #(
		.INIT('h4)
	) name6055 (
		_w7015_,
		_w7056_,
		_w7057_
	);
	LUT2 #(
		.INIT('h1)
	) name6056 (
		_w7014_,
		_w7057_,
		_w7058_
	);
	LUT2 #(
		.INIT('h1)
	) name6057 (
		_w7005_,
		_w7058_,
		_w7059_
	);
	LUT2 #(
		.INIT('h1)
	) name6058 (
		_w7004_,
		_w7059_,
		_w7060_
	);
	LUT2 #(
		.INIT('h8)
	) name6059 (
		\A[739] ,
		\A[740] ,
		_w7061_
	);
	LUT2 #(
		.INIT('h1)
	) name6060 (
		\A[739] ,
		\A[740] ,
		_w7062_
	);
	LUT2 #(
		.INIT('h1)
	) name6061 (
		_w7061_,
		_w7062_,
		_w7063_
	);
	LUT2 #(
		.INIT('h8)
	) name6062 (
		\A[741] ,
		_w7063_,
		_w7064_
	);
	LUT2 #(
		.INIT('h1)
	) name6063 (
		\A[741] ,
		_w7063_,
		_w7065_
	);
	LUT2 #(
		.INIT('h1)
	) name6064 (
		_w7064_,
		_w7065_,
		_w7066_
	);
	LUT2 #(
		.INIT('h8)
	) name6065 (
		\A[742] ,
		\A[743] ,
		_w7067_
	);
	LUT2 #(
		.INIT('h1)
	) name6066 (
		\A[742] ,
		\A[743] ,
		_w7068_
	);
	LUT2 #(
		.INIT('h1)
	) name6067 (
		_w7067_,
		_w7068_,
		_w7069_
	);
	LUT2 #(
		.INIT('h8)
	) name6068 (
		\A[744] ,
		_w7069_,
		_w7070_
	);
	LUT2 #(
		.INIT('h1)
	) name6069 (
		\A[744] ,
		_w7069_,
		_w7071_
	);
	LUT2 #(
		.INIT('h1)
	) name6070 (
		_w7070_,
		_w7071_,
		_w7072_
	);
	LUT2 #(
		.INIT('h8)
	) name6071 (
		_w7066_,
		_w7072_,
		_w7073_
	);
	LUT2 #(
		.INIT('h1)
	) name6072 (
		_w7066_,
		_w7072_,
		_w7074_
	);
	LUT2 #(
		.INIT('h1)
	) name6073 (
		_w7073_,
		_w7074_,
		_w7075_
	);
	LUT2 #(
		.INIT('h8)
	) name6074 (
		\A[745] ,
		\A[746] ,
		_w7076_
	);
	LUT2 #(
		.INIT('h1)
	) name6075 (
		\A[745] ,
		\A[746] ,
		_w7077_
	);
	LUT2 #(
		.INIT('h1)
	) name6076 (
		_w7076_,
		_w7077_,
		_w7078_
	);
	LUT2 #(
		.INIT('h8)
	) name6077 (
		\A[747] ,
		_w7078_,
		_w7079_
	);
	LUT2 #(
		.INIT('h1)
	) name6078 (
		\A[747] ,
		_w7078_,
		_w7080_
	);
	LUT2 #(
		.INIT('h1)
	) name6079 (
		_w7079_,
		_w7080_,
		_w7081_
	);
	LUT2 #(
		.INIT('h8)
	) name6080 (
		\A[748] ,
		\A[749] ,
		_w7082_
	);
	LUT2 #(
		.INIT('h1)
	) name6081 (
		\A[748] ,
		\A[749] ,
		_w7083_
	);
	LUT2 #(
		.INIT('h1)
	) name6082 (
		_w7082_,
		_w7083_,
		_w7084_
	);
	LUT2 #(
		.INIT('h8)
	) name6083 (
		\A[750] ,
		_w7084_,
		_w7085_
	);
	LUT2 #(
		.INIT('h1)
	) name6084 (
		\A[750] ,
		_w7084_,
		_w7086_
	);
	LUT2 #(
		.INIT('h1)
	) name6085 (
		_w7085_,
		_w7086_,
		_w7087_
	);
	LUT2 #(
		.INIT('h8)
	) name6086 (
		_w7081_,
		_w7087_,
		_w7088_
	);
	LUT2 #(
		.INIT('h1)
	) name6087 (
		_w7081_,
		_w7087_,
		_w7089_
	);
	LUT2 #(
		.INIT('h1)
	) name6088 (
		_w7088_,
		_w7089_,
		_w7090_
	);
	LUT2 #(
		.INIT('h8)
	) name6089 (
		_w7075_,
		_w7090_,
		_w7091_
	);
	LUT2 #(
		.INIT('h1)
	) name6090 (
		_w7082_,
		_w7085_,
		_w7092_
	);
	LUT2 #(
		.INIT('h1)
	) name6091 (
		_w7076_,
		_w7079_,
		_w7093_
	);
	LUT2 #(
		.INIT('h8)
	) name6092 (
		_w7092_,
		_w7093_,
		_w7094_
	);
	LUT2 #(
		.INIT('h1)
	) name6093 (
		_w7092_,
		_w7093_,
		_w7095_
	);
	LUT2 #(
		.INIT('h1)
	) name6094 (
		_w7094_,
		_w7095_,
		_w7096_
	);
	LUT2 #(
		.INIT('h8)
	) name6095 (
		_w7091_,
		_w7096_,
		_w7097_
	);
	LUT2 #(
		.INIT('h1)
	) name6096 (
		_w7061_,
		_w7064_,
		_w7098_
	);
	LUT2 #(
		.INIT('h8)
	) name6097 (
		_w7067_,
		_w7073_,
		_w7099_
	);
	LUT2 #(
		.INIT('h1)
	) name6098 (
		_w7067_,
		_w7070_,
		_w7100_
	);
	LUT2 #(
		.INIT('h4)
	) name6099 (
		_w7073_,
		_w7100_,
		_w7101_
	);
	LUT2 #(
		.INIT('h1)
	) name6100 (
		_w7099_,
		_w7101_,
		_w7102_
	);
	LUT2 #(
		.INIT('h2)
	) name6101 (
		_w7098_,
		_w7102_,
		_w7103_
	);
	LUT2 #(
		.INIT('h4)
	) name6102 (
		_w7098_,
		_w7102_,
		_w7104_
	);
	LUT2 #(
		.INIT('h1)
	) name6103 (
		_w7103_,
		_w7104_,
		_w7105_
	);
	LUT2 #(
		.INIT('h1)
	) name6104 (
		_w7097_,
		_w7105_,
		_w7106_
	);
	LUT2 #(
		.INIT('h4)
	) name6105 (
		_w7088_,
		_w7096_,
		_w7107_
	);
	LUT2 #(
		.INIT('h2)
	) name6106 (
		_w7088_,
		_w7096_,
		_w7108_
	);
	LUT2 #(
		.INIT('h1)
	) name6107 (
		_w7091_,
		_w7107_,
		_w7109_
	);
	LUT2 #(
		.INIT('h4)
	) name6108 (
		_w7108_,
		_w7109_,
		_w7110_
	);
	LUT2 #(
		.INIT('h1)
	) name6109 (
		_w7106_,
		_w7110_,
		_w7111_
	);
	LUT2 #(
		.INIT('h2)
	) name6110 (
		_w7088_,
		_w7094_,
		_w7112_
	);
	LUT2 #(
		.INIT('h1)
	) name6111 (
		_w7095_,
		_w7112_,
		_w7113_
	);
	LUT2 #(
		.INIT('h2)
	) name6112 (
		_w7111_,
		_w7113_,
		_w7114_
	);
	LUT2 #(
		.INIT('h4)
	) name6113 (
		_w7111_,
		_w7113_,
		_w7115_
	);
	LUT2 #(
		.INIT('h1)
	) name6114 (
		_w7098_,
		_w7101_,
		_w7116_
	);
	LUT2 #(
		.INIT('h1)
	) name6115 (
		_w7099_,
		_w7116_,
		_w7117_
	);
	LUT2 #(
		.INIT('h1)
	) name6116 (
		_w7115_,
		_w7117_,
		_w7118_
	);
	LUT2 #(
		.INIT('h1)
	) name6117 (
		_w7114_,
		_w7118_,
		_w7119_
	);
	LUT2 #(
		.INIT('h8)
	) name6118 (
		\A[727] ,
		\A[728] ,
		_w7120_
	);
	LUT2 #(
		.INIT('h1)
	) name6119 (
		\A[727] ,
		\A[728] ,
		_w7121_
	);
	LUT2 #(
		.INIT('h1)
	) name6120 (
		_w7120_,
		_w7121_,
		_w7122_
	);
	LUT2 #(
		.INIT('h8)
	) name6121 (
		\A[729] ,
		_w7122_,
		_w7123_
	);
	LUT2 #(
		.INIT('h1)
	) name6122 (
		\A[729] ,
		_w7122_,
		_w7124_
	);
	LUT2 #(
		.INIT('h1)
	) name6123 (
		_w7123_,
		_w7124_,
		_w7125_
	);
	LUT2 #(
		.INIT('h8)
	) name6124 (
		\A[730] ,
		\A[731] ,
		_w7126_
	);
	LUT2 #(
		.INIT('h1)
	) name6125 (
		\A[730] ,
		\A[731] ,
		_w7127_
	);
	LUT2 #(
		.INIT('h1)
	) name6126 (
		_w7126_,
		_w7127_,
		_w7128_
	);
	LUT2 #(
		.INIT('h8)
	) name6127 (
		\A[732] ,
		_w7128_,
		_w7129_
	);
	LUT2 #(
		.INIT('h1)
	) name6128 (
		\A[732] ,
		_w7128_,
		_w7130_
	);
	LUT2 #(
		.INIT('h1)
	) name6129 (
		_w7129_,
		_w7130_,
		_w7131_
	);
	LUT2 #(
		.INIT('h8)
	) name6130 (
		_w7125_,
		_w7131_,
		_w7132_
	);
	LUT2 #(
		.INIT('h1)
	) name6131 (
		_w7125_,
		_w7131_,
		_w7133_
	);
	LUT2 #(
		.INIT('h1)
	) name6132 (
		_w7132_,
		_w7133_,
		_w7134_
	);
	LUT2 #(
		.INIT('h8)
	) name6133 (
		\A[733] ,
		\A[734] ,
		_w7135_
	);
	LUT2 #(
		.INIT('h1)
	) name6134 (
		\A[733] ,
		\A[734] ,
		_w7136_
	);
	LUT2 #(
		.INIT('h1)
	) name6135 (
		_w7135_,
		_w7136_,
		_w7137_
	);
	LUT2 #(
		.INIT('h8)
	) name6136 (
		\A[735] ,
		_w7137_,
		_w7138_
	);
	LUT2 #(
		.INIT('h1)
	) name6137 (
		\A[735] ,
		_w7137_,
		_w7139_
	);
	LUT2 #(
		.INIT('h1)
	) name6138 (
		_w7138_,
		_w7139_,
		_w7140_
	);
	LUT2 #(
		.INIT('h8)
	) name6139 (
		\A[736] ,
		\A[737] ,
		_w7141_
	);
	LUT2 #(
		.INIT('h1)
	) name6140 (
		\A[736] ,
		\A[737] ,
		_w7142_
	);
	LUT2 #(
		.INIT('h1)
	) name6141 (
		_w7141_,
		_w7142_,
		_w7143_
	);
	LUT2 #(
		.INIT('h8)
	) name6142 (
		\A[738] ,
		_w7143_,
		_w7144_
	);
	LUT2 #(
		.INIT('h1)
	) name6143 (
		\A[738] ,
		_w7143_,
		_w7145_
	);
	LUT2 #(
		.INIT('h1)
	) name6144 (
		_w7144_,
		_w7145_,
		_w7146_
	);
	LUT2 #(
		.INIT('h8)
	) name6145 (
		_w7140_,
		_w7146_,
		_w7147_
	);
	LUT2 #(
		.INIT('h1)
	) name6146 (
		_w7140_,
		_w7146_,
		_w7148_
	);
	LUT2 #(
		.INIT('h1)
	) name6147 (
		_w7147_,
		_w7148_,
		_w7149_
	);
	LUT2 #(
		.INIT('h8)
	) name6148 (
		_w7134_,
		_w7149_,
		_w7150_
	);
	LUT2 #(
		.INIT('h1)
	) name6149 (
		_w7141_,
		_w7144_,
		_w7151_
	);
	LUT2 #(
		.INIT('h1)
	) name6150 (
		_w7135_,
		_w7138_,
		_w7152_
	);
	LUT2 #(
		.INIT('h8)
	) name6151 (
		_w7151_,
		_w7152_,
		_w7153_
	);
	LUT2 #(
		.INIT('h1)
	) name6152 (
		_w7151_,
		_w7152_,
		_w7154_
	);
	LUT2 #(
		.INIT('h1)
	) name6153 (
		_w7153_,
		_w7154_,
		_w7155_
	);
	LUT2 #(
		.INIT('h8)
	) name6154 (
		_w7150_,
		_w7155_,
		_w7156_
	);
	LUT2 #(
		.INIT('h1)
	) name6155 (
		_w7120_,
		_w7123_,
		_w7157_
	);
	LUT2 #(
		.INIT('h8)
	) name6156 (
		_w7126_,
		_w7132_,
		_w7158_
	);
	LUT2 #(
		.INIT('h1)
	) name6157 (
		_w7126_,
		_w7129_,
		_w7159_
	);
	LUT2 #(
		.INIT('h4)
	) name6158 (
		_w7132_,
		_w7159_,
		_w7160_
	);
	LUT2 #(
		.INIT('h1)
	) name6159 (
		_w7158_,
		_w7160_,
		_w7161_
	);
	LUT2 #(
		.INIT('h2)
	) name6160 (
		_w7157_,
		_w7161_,
		_w7162_
	);
	LUT2 #(
		.INIT('h4)
	) name6161 (
		_w7157_,
		_w7161_,
		_w7163_
	);
	LUT2 #(
		.INIT('h1)
	) name6162 (
		_w7162_,
		_w7163_,
		_w7164_
	);
	LUT2 #(
		.INIT('h1)
	) name6163 (
		_w7156_,
		_w7164_,
		_w7165_
	);
	LUT2 #(
		.INIT('h4)
	) name6164 (
		_w7147_,
		_w7155_,
		_w7166_
	);
	LUT2 #(
		.INIT('h2)
	) name6165 (
		_w7147_,
		_w7155_,
		_w7167_
	);
	LUT2 #(
		.INIT('h1)
	) name6166 (
		_w7150_,
		_w7166_,
		_w7168_
	);
	LUT2 #(
		.INIT('h4)
	) name6167 (
		_w7167_,
		_w7168_,
		_w7169_
	);
	LUT2 #(
		.INIT('h1)
	) name6168 (
		_w7165_,
		_w7169_,
		_w7170_
	);
	LUT2 #(
		.INIT('h2)
	) name6169 (
		_w7147_,
		_w7153_,
		_w7171_
	);
	LUT2 #(
		.INIT('h1)
	) name6170 (
		_w7154_,
		_w7171_,
		_w7172_
	);
	LUT2 #(
		.INIT('h2)
	) name6171 (
		_w7170_,
		_w7172_,
		_w7173_
	);
	LUT2 #(
		.INIT('h4)
	) name6172 (
		_w7170_,
		_w7172_,
		_w7174_
	);
	LUT2 #(
		.INIT('h1)
	) name6173 (
		_w7157_,
		_w7160_,
		_w7175_
	);
	LUT2 #(
		.INIT('h1)
	) name6174 (
		_w7158_,
		_w7175_,
		_w7176_
	);
	LUT2 #(
		.INIT('h1)
	) name6175 (
		_w7174_,
		_w7176_,
		_w7177_
	);
	LUT2 #(
		.INIT('h1)
	) name6176 (
		_w7173_,
		_w7177_,
		_w7178_
	);
	LUT2 #(
		.INIT('h1)
	) name6177 (
		_w7119_,
		_w7178_,
		_w7179_
	);
	LUT2 #(
		.INIT('h8)
	) name6178 (
		_w7119_,
		_w7178_,
		_w7180_
	);
	LUT2 #(
		.INIT('h1)
	) name6179 (
		_w7179_,
		_w7180_,
		_w7181_
	);
	LUT2 #(
		.INIT('h1)
	) name6180 (
		_w7173_,
		_w7174_,
		_w7182_
	);
	LUT2 #(
		.INIT('h4)
	) name6181 (
		_w7176_,
		_w7182_,
		_w7183_
	);
	LUT2 #(
		.INIT('h2)
	) name6182 (
		_w7176_,
		_w7182_,
		_w7184_
	);
	LUT2 #(
		.INIT('h1)
	) name6183 (
		_w7183_,
		_w7184_,
		_w7185_
	);
	LUT2 #(
		.INIT('h1)
	) name6184 (
		_w7114_,
		_w7115_,
		_w7186_
	);
	LUT2 #(
		.INIT('h4)
	) name6185 (
		_w7117_,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h2)
	) name6186 (
		_w7117_,
		_w7186_,
		_w7188_
	);
	LUT2 #(
		.INIT('h1)
	) name6187 (
		_w7187_,
		_w7188_,
		_w7189_
	);
	LUT2 #(
		.INIT('h1)
	) name6188 (
		_w7185_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h8)
	) name6189 (
		_w7185_,
		_w7189_,
		_w7191_
	);
	LUT2 #(
		.INIT('h1)
	) name6190 (
		_w7075_,
		_w7090_,
		_w7192_
	);
	LUT2 #(
		.INIT('h1)
	) name6191 (
		_w7091_,
		_w7192_,
		_w7193_
	);
	LUT2 #(
		.INIT('h1)
	) name6192 (
		_w7134_,
		_w7149_,
		_w7194_
	);
	LUT2 #(
		.INIT('h1)
	) name6193 (
		_w7150_,
		_w7194_,
		_w7195_
	);
	LUT2 #(
		.INIT('h8)
	) name6194 (
		_w7193_,
		_w7195_,
		_w7196_
	);
	LUT2 #(
		.INIT('h1)
	) name6195 (
		_w7097_,
		_w7110_,
		_w7197_
	);
	LUT2 #(
		.INIT('h4)
	) name6196 (
		_w7105_,
		_w7197_,
		_w7198_
	);
	LUT2 #(
		.INIT('h2)
	) name6197 (
		_w7105_,
		_w7197_,
		_w7199_
	);
	LUT2 #(
		.INIT('h1)
	) name6198 (
		_w7198_,
		_w7199_,
		_w7200_
	);
	LUT2 #(
		.INIT('h2)
	) name6199 (
		_w7196_,
		_w7200_,
		_w7201_
	);
	LUT2 #(
		.INIT('h4)
	) name6200 (
		_w7196_,
		_w7200_,
		_w7202_
	);
	LUT2 #(
		.INIT('h1)
	) name6201 (
		_w7156_,
		_w7169_,
		_w7203_
	);
	LUT2 #(
		.INIT('h4)
	) name6202 (
		_w7164_,
		_w7203_,
		_w7204_
	);
	LUT2 #(
		.INIT('h2)
	) name6203 (
		_w7164_,
		_w7203_,
		_w7205_
	);
	LUT2 #(
		.INIT('h1)
	) name6204 (
		_w7204_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('h1)
	) name6205 (
		_w7202_,
		_w7206_,
		_w7207_
	);
	LUT2 #(
		.INIT('h1)
	) name6206 (
		_w7201_,
		_w7207_,
		_w7208_
	);
	LUT2 #(
		.INIT('h4)
	) name6207 (
		_w7191_,
		_w7208_,
		_w7209_
	);
	LUT2 #(
		.INIT('h1)
	) name6208 (
		_w7190_,
		_w7209_,
		_w7210_
	);
	LUT2 #(
		.INIT('h2)
	) name6209 (
		_w7181_,
		_w7210_,
		_w7211_
	);
	LUT2 #(
		.INIT('h4)
	) name6210 (
		_w7181_,
		_w7210_,
		_w7212_
	);
	LUT2 #(
		.INIT('h1)
	) name6211 (
		_w7211_,
		_w7212_,
		_w7213_
	);
	LUT2 #(
		.INIT('h8)
	) name6212 (
		\A[715] ,
		\A[716] ,
		_w7214_
	);
	LUT2 #(
		.INIT('h1)
	) name6213 (
		\A[715] ,
		\A[716] ,
		_w7215_
	);
	LUT2 #(
		.INIT('h1)
	) name6214 (
		_w7214_,
		_w7215_,
		_w7216_
	);
	LUT2 #(
		.INIT('h8)
	) name6215 (
		\A[717] ,
		_w7216_,
		_w7217_
	);
	LUT2 #(
		.INIT('h1)
	) name6216 (
		\A[717] ,
		_w7216_,
		_w7218_
	);
	LUT2 #(
		.INIT('h1)
	) name6217 (
		_w7217_,
		_w7218_,
		_w7219_
	);
	LUT2 #(
		.INIT('h8)
	) name6218 (
		\A[718] ,
		\A[719] ,
		_w7220_
	);
	LUT2 #(
		.INIT('h1)
	) name6219 (
		\A[718] ,
		\A[719] ,
		_w7221_
	);
	LUT2 #(
		.INIT('h1)
	) name6220 (
		_w7220_,
		_w7221_,
		_w7222_
	);
	LUT2 #(
		.INIT('h8)
	) name6221 (
		\A[720] ,
		_w7222_,
		_w7223_
	);
	LUT2 #(
		.INIT('h1)
	) name6222 (
		\A[720] ,
		_w7222_,
		_w7224_
	);
	LUT2 #(
		.INIT('h1)
	) name6223 (
		_w7223_,
		_w7224_,
		_w7225_
	);
	LUT2 #(
		.INIT('h8)
	) name6224 (
		_w7219_,
		_w7225_,
		_w7226_
	);
	LUT2 #(
		.INIT('h1)
	) name6225 (
		_w7219_,
		_w7225_,
		_w7227_
	);
	LUT2 #(
		.INIT('h1)
	) name6226 (
		_w7226_,
		_w7227_,
		_w7228_
	);
	LUT2 #(
		.INIT('h8)
	) name6227 (
		\A[721] ,
		\A[722] ,
		_w7229_
	);
	LUT2 #(
		.INIT('h1)
	) name6228 (
		\A[721] ,
		\A[722] ,
		_w7230_
	);
	LUT2 #(
		.INIT('h1)
	) name6229 (
		_w7229_,
		_w7230_,
		_w7231_
	);
	LUT2 #(
		.INIT('h8)
	) name6230 (
		\A[723] ,
		_w7231_,
		_w7232_
	);
	LUT2 #(
		.INIT('h1)
	) name6231 (
		\A[723] ,
		_w7231_,
		_w7233_
	);
	LUT2 #(
		.INIT('h1)
	) name6232 (
		_w7232_,
		_w7233_,
		_w7234_
	);
	LUT2 #(
		.INIT('h8)
	) name6233 (
		\A[724] ,
		\A[725] ,
		_w7235_
	);
	LUT2 #(
		.INIT('h1)
	) name6234 (
		\A[724] ,
		\A[725] ,
		_w7236_
	);
	LUT2 #(
		.INIT('h1)
	) name6235 (
		_w7235_,
		_w7236_,
		_w7237_
	);
	LUT2 #(
		.INIT('h8)
	) name6236 (
		\A[726] ,
		_w7237_,
		_w7238_
	);
	LUT2 #(
		.INIT('h1)
	) name6237 (
		\A[726] ,
		_w7237_,
		_w7239_
	);
	LUT2 #(
		.INIT('h1)
	) name6238 (
		_w7238_,
		_w7239_,
		_w7240_
	);
	LUT2 #(
		.INIT('h8)
	) name6239 (
		_w7234_,
		_w7240_,
		_w7241_
	);
	LUT2 #(
		.INIT('h1)
	) name6240 (
		_w7234_,
		_w7240_,
		_w7242_
	);
	LUT2 #(
		.INIT('h1)
	) name6241 (
		_w7241_,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h8)
	) name6242 (
		_w7228_,
		_w7243_,
		_w7244_
	);
	LUT2 #(
		.INIT('h1)
	) name6243 (
		_w7235_,
		_w7238_,
		_w7245_
	);
	LUT2 #(
		.INIT('h1)
	) name6244 (
		_w7229_,
		_w7232_,
		_w7246_
	);
	LUT2 #(
		.INIT('h8)
	) name6245 (
		_w7245_,
		_w7246_,
		_w7247_
	);
	LUT2 #(
		.INIT('h1)
	) name6246 (
		_w7245_,
		_w7246_,
		_w7248_
	);
	LUT2 #(
		.INIT('h1)
	) name6247 (
		_w7247_,
		_w7248_,
		_w7249_
	);
	LUT2 #(
		.INIT('h8)
	) name6248 (
		_w7244_,
		_w7249_,
		_w7250_
	);
	LUT2 #(
		.INIT('h1)
	) name6249 (
		_w7214_,
		_w7217_,
		_w7251_
	);
	LUT2 #(
		.INIT('h8)
	) name6250 (
		_w7220_,
		_w7226_,
		_w7252_
	);
	LUT2 #(
		.INIT('h1)
	) name6251 (
		_w7220_,
		_w7223_,
		_w7253_
	);
	LUT2 #(
		.INIT('h4)
	) name6252 (
		_w7226_,
		_w7253_,
		_w7254_
	);
	LUT2 #(
		.INIT('h1)
	) name6253 (
		_w7252_,
		_w7254_,
		_w7255_
	);
	LUT2 #(
		.INIT('h2)
	) name6254 (
		_w7251_,
		_w7255_,
		_w7256_
	);
	LUT2 #(
		.INIT('h4)
	) name6255 (
		_w7251_,
		_w7255_,
		_w7257_
	);
	LUT2 #(
		.INIT('h1)
	) name6256 (
		_w7256_,
		_w7257_,
		_w7258_
	);
	LUT2 #(
		.INIT('h1)
	) name6257 (
		_w7250_,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('h4)
	) name6258 (
		_w7241_,
		_w7249_,
		_w7260_
	);
	LUT2 #(
		.INIT('h2)
	) name6259 (
		_w7241_,
		_w7249_,
		_w7261_
	);
	LUT2 #(
		.INIT('h1)
	) name6260 (
		_w7244_,
		_w7260_,
		_w7262_
	);
	LUT2 #(
		.INIT('h4)
	) name6261 (
		_w7261_,
		_w7262_,
		_w7263_
	);
	LUT2 #(
		.INIT('h1)
	) name6262 (
		_w7259_,
		_w7263_,
		_w7264_
	);
	LUT2 #(
		.INIT('h2)
	) name6263 (
		_w7241_,
		_w7247_,
		_w7265_
	);
	LUT2 #(
		.INIT('h1)
	) name6264 (
		_w7248_,
		_w7265_,
		_w7266_
	);
	LUT2 #(
		.INIT('h2)
	) name6265 (
		_w7264_,
		_w7266_,
		_w7267_
	);
	LUT2 #(
		.INIT('h4)
	) name6266 (
		_w7264_,
		_w7266_,
		_w7268_
	);
	LUT2 #(
		.INIT('h1)
	) name6267 (
		_w7251_,
		_w7254_,
		_w7269_
	);
	LUT2 #(
		.INIT('h1)
	) name6268 (
		_w7252_,
		_w7269_,
		_w7270_
	);
	LUT2 #(
		.INIT('h1)
	) name6269 (
		_w7268_,
		_w7270_,
		_w7271_
	);
	LUT2 #(
		.INIT('h1)
	) name6270 (
		_w7267_,
		_w7271_,
		_w7272_
	);
	LUT2 #(
		.INIT('h8)
	) name6271 (
		\A[709] ,
		\A[710] ,
		_w7273_
	);
	LUT2 #(
		.INIT('h1)
	) name6272 (
		\A[709] ,
		\A[710] ,
		_w7274_
	);
	LUT2 #(
		.INIT('h1)
	) name6273 (
		_w7273_,
		_w7274_,
		_w7275_
	);
	LUT2 #(
		.INIT('h8)
	) name6274 (
		\A[711] ,
		_w7275_,
		_w7276_
	);
	LUT2 #(
		.INIT('h1)
	) name6275 (
		\A[711] ,
		_w7275_,
		_w7277_
	);
	LUT2 #(
		.INIT('h1)
	) name6276 (
		_w7276_,
		_w7277_,
		_w7278_
	);
	LUT2 #(
		.INIT('h8)
	) name6277 (
		\A[712] ,
		\A[713] ,
		_w7279_
	);
	LUT2 #(
		.INIT('h1)
	) name6278 (
		\A[712] ,
		\A[713] ,
		_w7280_
	);
	LUT2 #(
		.INIT('h1)
	) name6279 (
		_w7279_,
		_w7280_,
		_w7281_
	);
	LUT2 #(
		.INIT('h8)
	) name6280 (
		\A[714] ,
		_w7281_,
		_w7282_
	);
	LUT2 #(
		.INIT('h1)
	) name6281 (
		\A[714] ,
		_w7281_,
		_w7283_
	);
	LUT2 #(
		.INIT('h1)
	) name6282 (
		_w7282_,
		_w7283_,
		_w7284_
	);
	LUT2 #(
		.INIT('h8)
	) name6283 (
		_w7278_,
		_w7284_,
		_w7285_
	);
	LUT2 #(
		.INIT('h1)
	) name6284 (
		_w7278_,
		_w7284_,
		_w7286_
	);
	LUT2 #(
		.INIT('h1)
	) name6285 (
		_w7285_,
		_w7286_,
		_w7287_
	);
	LUT2 #(
		.INIT('h8)
	) name6286 (
		\A[703] ,
		\A[704] ,
		_w7288_
	);
	LUT2 #(
		.INIT('h1)
	) name6287 (
		\A[703] ,
		\A[704] ,
		_w7289_
	);
	LUT2 #(
		.INIT('h1)
	) name6288 (
		_w7288_,
		_w7289_,
		_w7290_
	);
	LUT2 #(
		.INIT('h8)
	) name6289 (
		\A[705] ,
		_w7290_,
		_w7291_
	);
	LUT2 #(
		.INIT('h1)
	) name6290 (
		\A[705] ,
		_w7290_,
		_w7292_
	);
	LUT2 #(
		.INIT('h1)
	) name6291 (
		_w7291_,
		_w7292_,
		_w7293_
	);
	LUT2 #(
		.INIT('h8)
	) name6292 (
		\A[706] ,
		\A[707] ,
		_w7294_
	);
	LUT2 #(
		.INIT('h1)
	) name6293 (
		\A[706] ,
		\A[707] ,
		_w7295_
	);
	LUT2 #(
		.INIT('h1)
	) name6294 (
		_w7294_,
		_w7295_,
		_w7296_
	);
	LUT2 #(
		.INIT('h8)
	) name6295 (
		\A[708] ,
		_w7296_,
		_w7297_
	);
	LUT2 #(
		.INIT('h1)
	) name6296 (
		\A[708] ,
		_w7296_,
		_w7298_
	);
	LUT2 #(
		.INIT('h1)
	) name6297 (
		_w7297_,
		_w7298_,
		_w7299_
	);
	LUT2 #(
		.INIT('h8)
	) name6298 (
		_w7293_,
		_w7299_,
		_w7300_
	);
	LUT2 #(
		.INIT('h1)
	) name6299 (
		_w7293_,
		_w7299_,
		_w7301_
	);
	LUT2 #(
		.INIT('h1)
	) name6300 (
		_w7300_,
		_w7301_,
		_w7302_
	);
	LUT2 #(
		.INIT('h8)
	) name6301 (
		_w7287_,
		_w7302_,
		_w7303_
	);
	LUT2 #(
		.INIT('h1)
	) name6302 (
		_w7279_,
		_w7282_,
		_w7304_
	);
	LUT2 #(
		.INIT('h1)
	) name6303 (
		_w7273_,
		_w7276_,
		_w7305_
	);
	LUT2 #(
		.INIT('h1)
	) name6304 (
		_w7304_,
		_w7305_,
		_w7306_
	);
	LUT2 #(
		.INIT('h8)
	) name6305 (
		_w7304_,
		_w7305_,
		_w7307_
	);
	LUT2 #(
		.INIT('h1)
	) name6306 (
		_w7306_,
		_w7307_,
		_w7308_
	);
	LUT2 #(
		.INIT('h8)
	) name6307 (
		_w7303_,
		_w7308_,
		_w7309_
	);
	LUT2 #(
		.INIT('h1)
	) name6308 (
		_w7294_,
		_w7297_,
		_w7310_
	);
	LUT2 #(
		.INIT('h1)
	) name6309 (
		_w7288_,
		_w7291_,
		_w7311_
	);
	LUT2 #(
		.INIT('h1)
	) name6310 (
		_w7310_,
		_w7311_,
		_w7312_
	);
	LUT2 #(
		.INIT('h8)
	) name6311 (
		_w7310_,
		_w7311_,
		_w7313_
	);
	LUT2 #(
		.INIT('h1)
	) name6312 (
		_w7312_,
		_w7313_,
		_w7314_
	);
	LUT2 #(
		.INIT('h2)
	) name6313 (
		_w7300_,
		_w7314_,
		_w7315_
	);
	LUT2 #(
		.INIT('h4)
	) name6314 (
		_w7300_,
		_w7314_,
		_w7316_
	);
	LUT2 #(
		.INIT('h1)
	) name6315 (
		_w7315_,
		_w7316_,
		_w7317_
	);
	LUT2 #(
		.INIT('h4)
	) name6316 (
		_w7309_,
		_w7317_,
		_w7318_
	);
	LUT2 #(
		.INIT('h4)
	) name6317 (
		_w7285_,
		_w7308_,
		_w7319_
	);
	LUT2 #(
		.INIT('h2)
	) name6318 (
		_w7285_,
		_w7308_,
		_w7320_
	);
	LUT2 #(
		.INIT('h1)
	) name6319 (
		_w7303_,
		_w7319_,
		_w7321_
	);
	LUT2 #(
		.INIT('h4)
	) name6320 (
		_w7320_,
		_w7321_,
		_w7322_
	);
	LUT2 #(
		.INIT('h1)
	) name6321 (
		_w7318_,
		_w7322_,
		_w7323_
	);
	LUT2 #(
		.INIT('h1)
	) name6322 (
		_w7285_,
		_w7306_,
		_w7324_
	);
	LUT2 #(
		.INIT('h1)
	) name6323 (
		_w7307_,
		_w7324_,
		_w7325_
	);
	LUT2 #(
		.INIT('h1)
	) name6324 (
		_w7323_,
		_w7325_,
		_w7326_
	);
	LUT2 #(
		.INIT('h8)
	) name6325 (
		_w7323_,
		_w7325_,
		_w7327_
	);
	LUT2 #(
		.INIT('h1)
	) name6326 (
		_w7300_,
		_w7312_,
		_w7328_
	);
	LUT2 #(
		.INIT('h1)
	) name6327 (
		_w7313_,
		_w7328_,
		_w7329_
	);
	LUT2 #(
		.INIT('h1)
	) name6328 (
		_w7327_,
		_w7329_,
		_w7330_
	);
	LUT2 #(
		.INIT('h1)
	) name6329 (
		_w7326_,
		_w7330_,
		_w7331_
	);
	LUT2 #(
		.INIT('h4)
	) name6330 (
		_w7272_,
		_w7331_,
		_w7332_
	);
	LUT2 #(
		.INIT('h2)
	) name6331 (
		_w7272_,
		_w7331_,
		_w7333_
	);
	LUT2 #(
		.INIT('h1)
	) name6332 (
		_w7332_,
		_w7333_,
		_w7334_
	);
	LUT2 #(
		.INIT('h1)
	) name6333 (
		_w7326_,
		_w7327_,
		_w7335_
	);
	LUT2 #(
		.INIT('h4)
	) name6334 (
		_w7329_,
		_w7335_,
		_w7336_
	);
	LUT2 #(
		.INIT('h2)
	) name6335 (
		_w7329_,
		_w7335_,
		_w7337_
	);
	LUT2 #(
		.INIT('h1)
	) name6336 (
		_w7336_,
		_w7337_,
		_w7338_
	);
	LUT2 #(
		.INIT('h1)
	) name6337 (
		_w7267_,
		_w7268_,
		_w7339_
	);
	LUT2 #(
		.INIT('h4)
	) name6338 (
		_w7270_,
		_w7339_,
		_w7340_
	);
	LUT2 #(
		.INIT('h2)
	) name6339 (
		_w7270_,
		_w7339_,
		_w7341_
	);
	LUT2 #(
		.INIT('h1)
	) name6340 (
		_w7340_,
		_w7341_,
		_w7342_
	);
	LUT2 #(
		.INIT('h4)
	) name6341 (
		_w7338_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h2)
	) name6342 (
		_w7338_,
		_w7342_,
		_w7344_
	);
	LUT2 #(
		.INIT('h1)
	) name6343 (
		_w7228_,
		_w7243_,
		_w7345_
	);
	LUT2 #(
		.INIT('h1)
	) name6344 (
		_w7244_,
		_w7345_,
		_w7346_
	);
	LUT2 #(
		.INIT('h1)
	) name6345 (
		_w7287_,
		_w7302_,
		_w7347_
	);
	LUT2 #(
		.INIT('h1)
	) name6346 (
		_w7303_,
		_w7347_,
		_w7348_
	);
	LUT2 #(
		.INIT('h8)
	) name6347 (
		_w7346_,
		_w7348_,
		_w7349_
	);
	LUT2 #(
		.INIT('h1)
	) name6348 (
		_w7250_,
		_w7263_,
		_w7350_
	);
	LUT2 #(
		.INIT('h4)
	) name6349 (
		_w7258_,
		_w7350_,
		_w7351_
	);
	LUT2 #(
		.INIT('h2)
	) name6350 (
		_w7258_,
		_w7350_,
		_w7352_
	);
	LUT2 #(
		.INIT('h1)
	) name6351 (
		_w7351_,
		_w7352_,
		_w7353_
	);
	LUT2 #(
		.INIT('h2)
	) name6352 (
		_w7349_,
		_w7353_,
		_w7354_
	);
	LUT2 #(
		.INIT('h4)
	) name6353 (
		_w7349_,
		_w7353_,
		_w7355_
	);
	LUT2 #(
		.INIT('h1)
	) name6354 (
		_w7309_,
		_w7322_,
		_w7356_
	);
	LUT2 #(
		.INIT('h8)
	) name6355 (
		_w7317_,
		_w7356_,
		_w7357_
	);
	LUT2 #(
		.INIT('h1)
	) name6356 (
		_w7317_,
		_w7356_,
		_w7358_
	);
	LUT2 #(
		.INIT('h1)
	) name6357 (
		_w7357_,
		_w7358_,
		_w7359_
	);
	LUT2 #(
		.INIT('h1)
	) name6358 (
		_w7355_,
		_w7359_,
		_w7360_
	);
	LUT2 #(
		.INIT('h1)
	) name6359 (
		_w7354_,
		_w7360_,
		_w7361_
	);
	LUT2 #(
		.INIT('h1)
	) name6360 (
		_w7344_,
		_w7361_,
		_w7362_
	);
	LUT2 #(
		.INIT('h1)
	) name6361 (
		_w7343_,
		_w7362_,
		_w7363_
	);
	LUT2 #(
		.INIT('h2)
	) name6362 (
		_w7334_,
		_w7363_,
		_w7364_
	);
	LUT2 #(
		.INIT('h4)
	) name6363 (
		_w7334_,
		_w7363_,
		_w7365_
	);
	LUT2 #(
		.INIT('h1)
	) name6364 (
		_w7364_,
		_w7365_,
		_w7366_
	);
	LUT2 #(
		.INIT('h2)
	) name6365 (
		_w7213_,
		_w7366_,
		_w7367_
	);
	LUT2 #(
		.INIT('h4)
	) name6366 (
		_w7213_,
		_w7366_,
		_w7368_
	);
	LUT2 #(
		.INIT('h1)
	) name6367 (
		_w7343_,
		_w7344_,
		_w7369_
	);
	LUT2 #(
		.INIT('h4)
	) name6368 (
		_w7361_,
		_w7369_,
		_w7370_
	);
	LUT2 #(
		.INIT('h2)
	) name6369 (
		_w7361_,
		_w7369_,
		_w7371_
	);
	LUT2 #(
		.INIT('h1)
	) name6370 (
		_w7370_,
		_w7371_,
		_w7372_
	);
	LUT2 #(
		.INIT('h1)
	) name6371 (
		_w7190_,
		_w7191_,
		_w7373_
	);
	LUT2 #(
		.INIT('h4)
	) name6372 (
		_w7208_,
		_w7373_,
		_w7374_
	);
	LUT2 #(
		.INIT('h2)
	) name6373 (
		_w7208_,
		_w7373_,
		_w7375_
	);
	LUT2 #(
		.INIT('h1)
	) name6374 (
		_w7374_,
		_w7375_,
		_w7376_
	);
	LUT2 #(
		.INIT('h1)
	) name6375 (
		_w7372_,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('h8)
	) name6376 (
		_w7372_,
		_w7376_,
		_w7378_
	);
	LUT2 #(
		.INIT('h1)
	) name6377 (
		_w7193_,
		_w7195_,
		_w7379_
	);
	LUT2 #(
		.INIT('h1)
	) name6378 (
		_w7196_,
		_w7379_,
		_w7380_
	);
	LUT2 #(
		.INIT('h1)
	) name6379 (
		_w7346_,
		_w7348_,
		_w7381_
	);
	LUT2 #(
		.INIT('h1)
	) name6380 (
		_w7349_,
		_w7381_,
		_w7382_
	);
	LUT2 #(
		.INIT('h8)
	) name6381 (
		_w7380_,
		_w7382_,
		_w7383_
	);
	LUT2 #(
		.INIT('h1)
	) name6382 (
		_w7201_,
		_w7202_,
		_w7384_
	);
	LUT2 #(
		.INIT('h4)
	) name6383 (
		_w7206_,
		_w7384_,
		_w7385_
	);
	LUT2 #(
		.INIT('h2)
	) name6384 (
		_w7206_,
		_w7384_,
		_w7386_
	);
	LUT2 #(
		.INIT('h1)
	) name6385 (
		_w7385_,
		_w7386_,
		_w7387_
	);
	LUT2 #(
		.INIT('h8)
	) name6386 (
		_w7383_,
		_w7387_,
		_w7388_
	);
	LUT2 #(
		.INIT('h1)
	) name6387 (
		_w7383_,
		_w7387_,
		_w7389_
	);
	LUT2 #(
		.INIT('h1)
	) name6388 (
		_w7354_,
		_w7355_,
		_w7390_
	);
	LUT2 #(
		.INIT('h4)
	) name6389 (
		_w7359_,
		_w7390_,
		_w7391_
	);
	LUT2 #(
		.INIT('h2)
	) name6390 (
		_w7359_,
		_w7390_,
		_w7392_
	);
	LUT2 #(
		.INIT('h1)
	) name6391 (
		_w7391_,
		_w7392_,
		_w7393_
	);
	LUT2 #(
		.INIT('h4)
	) name6392 (
		_w7389_,
		_w7393_,
		_w7394_
	);
	LUT2 #(
		.INIT('h1)
	) name6393 (
		_w7388_,
		_w7394_,
		_w7395_
	);
	LUT2 #(
		.INIT('h4)
	) name6394 (
		_w7378_,
		_w7395_,
		_w7396_
	);
	LUT2 #(
		.INIT('h1)
	) name6395 (
		_w7377_,
		_w7396_,
		_w7397_
	);
	LUT2 #(
		.INIT('h1)
	) name6396 (
		_w7368_,
		_w7397_,
		_w7398_
	);
	LUT2 #(
		.INIT('h1)
	) name6397 (
		_w7367_,
		_w7398_,
		_w7399_
	);
	LUT2 #(
		.INIT('h4)
	) name6398 (
		_w7180_,
		_w7210_,
		_w7400_
	);
	LUT2 #(
		.INIT('h1)
	) name6399 (
		_w7179_,
		_w7400_,
		_w7401_
	);
	LUT2 #(
		.INIT('h2)
	) name6400 (
		_w7399_,
		_w7401_,
		_w7402_
	);
	LUT2 #(
		.INIT('h4)
	) name6401 (
		_w7399_,
		_w7401_,
		_w7403_
	);
	LUT2 #(
		.INIT('h1)
	) name6402 (
		_w7333_,
		_w7363_,
		_w7404_
	);
	LUT2 #(
		.INIT('h1)
	) name6403 (
		_w7332_,
		_w7404_,
		_w7405_
	);
	LUT2 #(
		.INIT('h1)
	) name6404 (
		_w7403_,
		_w7405_,
		_w7406_
	);
	LUT2 #(
		.INIT('h1)
	) name6405 (
		_w7402_,
		_w7406_,
		_w7407_
	);
	LUT2 #(
		.INIT('h8)
	) name6406 (
		\A[658] ,
		\A[659] ,
		_w7408_
	);
	LUT2 #(
		.INIT('h8)
	) name6407 (
		\A[655] ,
		\A[656] ,
		_w7409_
	);
	LUT2 #(
		.INIT('h1)
	) name6408 (
		\A[655] ,
		\A[656] ,
		_w7410_
	);
	LUT2 #(
		.INIT('h1)
	) name6409 (
		_w7409_,
		_w7410_,
		_w7411_
	);
	LUT2 #(
		.INIT('h8)
	) name6410 (
		\A[657] ,
		_w7411_,
		_w7412_
	);
	LUT2 #(
		.INIT('h1)
	) name6411 (
		\A[657] ,
		_w7411_,
		_w7413_
	);
	LUT2 #(
		.INIT('h1)
	) name6412 (
		_w7412_,
		_w7413_,
		_w7414_
	);
	LUT2 #(
		.INIT('h1)
	) name6413 (
		\A[658] ,
		\A[659] ,
		_w7415_
	);
	LUT2 #(
		.INIT('h1)
	) name6414 (
		_w7408_,
		_w7415_,
		_w7416_
	);
	LUT2 #(
		.INIT('h8)
	) name6415 (
		\A[660] ,
		_w7416_,
		_w7417_
	);
	LUT2 #(
		.INIT('h1)
	) name6416 (
		\A[660] ,
		_w7416_,
		_w7418_
	);
	LUT2 #(
		.INIT('h1)
	) name6417 (
		_w7417_,
		_w7418_,
		_w7419_
	);
	LUT2 #(
		.INIT('h8)
	) name6418 (
		_w7414_,
		_w7419_,
		_w7420_
	);
	LUT2 #(
		.INIT('h8)
	) name6419 (
		_w7408_,
		_w7420_,
		_w7421_
	);
	LUT2 #(
		.INIT('h1)
	) name6420 (
		_w7409_,
		_w7412_,
		_w7422_
	);
	LUT2 #(
		.INIT('h1)
	) name6421 (
		_w7408_,
		_w7417_,
		_w7423_
	);
	LUT2 #(
		.INIT('h4)
	) name6422 (
		_w7420_,
		_w7423_,
		_w7424_
	);
	LUT2 #(
		.INIT('h1)
	) name6423 (
		_w7422_,
		_w7424_,
		_w7425_
	);
	LUT2 #(
		.INIT('h1)
	) name6424 (
		_w7421_,
		_w7425_,
		_w7426_
	);
	LUT2 #(
		.INIT('h8)
	) name6425 (
		\A[664] ,
		\A[665] ,
		_w7427_
	);
	LUT2 #(
		.INIT('h1)
	) name6426 (
		\A[664] ,
		\A[665] ,
		_w7428_
	);
	LUT2 #(
		.INIT('h1)
	) name6427 (
		_w7427_,
		_w7428_,
		_w7429_
	);
	LUT2 #(
		.INIT('h8)
	) name6428 (
		\A[666] ,
		_w7429_,
		_w7430_
	);
	LUT2 #(
		.INIT('h1)
	) name6429 (
		_w7427_,
		_w7430_,
		_w7431_
	);
	LUT2 #(
		.INIT('h8)
	) name6430 (
		\A[661] ,
		\A[662] ,
		_w7432_
	);
	LUT2 #(
		.INIT('h1)
	) name6431 (
		\A[661] ,
		\A[662] ,
		_w7433_
	);
	LUT2 #(
		.INIT('h1)
	) name6432 (
		_w7432_,
		_w7433_,
		_w7434_
	);
	LUT2 #(
		.INIT('h8)
	) name6433 (
		\A[663] ,
		_w7434_,
		_w7435_
	);
	LUT2 #(
		.INIT('h1)
	) name6434 (
		_w7432_,
		_w7435_,
		_w7436_
	);
	LUT2 #(
		.INIT('h8)
	) name6435 (
		_w7431_,
		_w7436_,
		_w7437_
	);
	LUT2 #(
		.INIT('h1)
	) name6436 (
		_w7431_,
		_w7436_,
		_w7438_
	);
	LUT2 #(
		.INIT('h1)
	) name6437 (
		\A[663] ,
		_w7434_,
		_w7439_
	);
	LUT2 #(
		.INIT('h1)
	) name6438 (
		_w7435_,
		_w7439_,
		_w7440_
	);
	LUT2 #(
		.INIT('h1)
	) name6439 (
		\A[666] ,
		_w7429_,
		_w7441_
	);
	LUT2 #(
		.INIT('h1)
	) name6440 (
		_w7430_,
		_w7441_,
		_w7442_
	);
	LUT2 #(
		.INIT('h8)
	) name6441 (
		_w7440_,
		_w7442_,
		_w7443_
	);
	LUT2 #(
		.INIT('h1)
	) name6442 (
		_w7438_,
		_w7443_,
		_w7444_
	);
	LUT2 #(
		.INIT('h1)
	) name6443 (
		_w7437_,
		_w7444_,
		_w7445_
	);
	LUT2 #(
		.INIT('h1)
	) name6444 (
		_w7440_,
		_w7442_,
		_w7446_
	);
	LUT2 #(
		.INIT('h1)
	) name6445 (
		_w7443_,
		_w7446_,
		_w7447_
	);
	LUT2 #(
		.INIT('h1)
	) name6446 (
		_w7414_,
		_w7419_,
		_w7448_
	);
	LUT2 #(
		.INIT('h1)
	) name6447 (
		_w7420_,
		_w7448_,
		_w7449_
	);
	LUT2 #(
		.INIT('h8)
	) name6448 (
		_w7447_,
		_w7449_,
		_w7450_
	);
	LUT2 #(
		.INIT('h2)
	) name6449 (
		_w7421_,
		_w7422_,
		_w7451_
	);
	LUT2 #(
		.INIT('h2)
	) name6450 (
		_w7450_,
		_w7451_,
		_w7452_
	);
	LUT2 #(
		.INIT('h1)
	) name6451 (
		_w7437_,
		_w7438_,
		_w7453_
	);
	LUT2 #(
		.INIT('h2)
	) name6452 (
		_w7443_,
		_w7453_,
		_w7454_
	);
	LUT2 #(
		.INIT('h4)
	) name6453 (
		_w7443_,
		_w7453_,
		_w7455_
	);
	LUT2 #(
		.INIT('h1)
	) name6454 (
		_w7454_,
		_w7455_,
		_w7456_
	);
	LUT2 #(
		.INIT('h2)
	) name6455 (
		_w7452_,
		_w7456_,
		_w7457_
	);
	LUT2 #(
		.INIT('h4)
	) name6456 (
		_w7452_,
		_w7456_,
		_w7458_
	);
	LUT2 #(
		.INIT('h1)
	) name6457 (
		_w7421_,
		_w7424_,
		_w7459_
	);
	LUT2 #(
		.INIT('h2)
	) name6458 (
		_w7422_,
		_w7459_,
		_w7460_
	);
	LUT2 #(
		.INIT('h4)
	) name6459 (
		_w7422_,
		_w7459_,
		_w7461_
	);
	LUT2 #(
		.INIT('h1)
	) name6460 (
		_w7460_,
		_w7461_,
		_w7462_
	);
	LUT2 #(
		.INIT('h4)
	) name6461 (
		_w7458_,
		_w7462_,
		_w7463_
	);
	LUT2 #(
		.INIT('h1)
	) name6462 (
		_w7457_,
		_w7463_,
		_w7464_
	);
	LUT2 #(
		.INIT('h2)
	) name6463 (
		_w7445_,
		_w7464_,
		_w7465_
	);
	LUT2 #(
		.INIT('h4)
	) name6464 (
		_w7445_,
		_w7464_,
		_w7466_
	);
	LUT2 #(
		.INIT('h1)
	) name6465 (
		_w7465_,
		_w7466_,
		_w7467_
	);
	LUT2 #(
		.INIT('h8)
	) name6466 (
		_w7426_,
		_w7467_,
		_w7468_
	);
	LUT2 #(
		.INIT('h1)
	) name6467 (
		_w7426_,
		_w7467_,
		_w7469_
	);
	LUT2 #(
		.INIT('h1)
	) name6468 (
		_w7468_,
		_w7469_,
		_w7470_
	);
	LUT2 #(
		.INIT('h8)
	) name6469 (
		\A[670] ,
		\A[671] ,
		_w7471_
	);
	LUT2 #(
		.INIT('h8)
	) name6470 (
		\A[667] ,
		\A[668] ,
		_w7472_
	);
	LUT2 #(
		.INIT('h1)
	) name6471 (
		\A[667] ,
		\A[668] ,
		_w7473_
	);
	LUT2 #(
		.INIT('h1)
	) name6472 (
		_w7472_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h8)
	) name6473 (
		\A[669] ,
		_w7474_,
		_w7475_
	);
	LUT2 #(
		.INIT('h1)
	) name6474 (
		\A[669] ,
		_w7474_,
		_w7476_
	);
	LUT2 #(
		.INIT('h1)
	) name6475 (
		_w7475_,
		_w7476_,
		_w7477_
	);
	LUT2 #(
		.INIT('h1)
	) name6476 (
		\A[670] ,
		\A[671] ,
		_w7478_
	);
	LUT2 #(
		.INIT('h1)
	) name6477 (
		_w7471_,
		_w7478_,
		_w7479_
	);
	LUT2 #(
		.INIT('h8)
	) name6478 (
		\A[672] ,
		_w7479_,
		_w7480_
	);
	LUT2 #(
		.INIT('h1)
	) name6479 (
		\A[672] ,
		_w7479_,
		_w7481_
	);
	LUT2 #(
		.INIT('h1)
	) name6480 (
		_w7480_,
		_w7481_,
		_w7482_
	);
	LUT2 #(
		.INIT('h8)
	) name6481 (
		_w7477_,
		_w7482_,
		_w7483_
	);
	LUT2 #(
		.INIT('h8)
	) name6482 (
		_w7471_,
		_w7483_,
		_w7484_
	);
	LUT2 #(
		.INIT('h1)
	) name6483 (
		_w7472_,
		_w7475_,
		_w7485_
	);
	LUT2 #(
		.INIT('h1)
	) name6484 (
		_w7471_,
		_w7480_,
		_w7486_
	);
	LUT2 #(
		.INIT('h4)
	) name6485 (
		_w7483_,
		_w7486_,
		_w7487_
	);
	LUT2 #(
		.INIT('h1)
	) name6486 (
		_w7485_,
		_w7487_,
		_w7488_
	);
	LUT2 #(
		.INIT('h1)
	) name6487 (
		_w7484_,
		_w7488_,
		_w7489_
	);
	LUT2 #(
		.INIT('h8)
	) name6488 (
		\A[676] ,
		\A[677] ,
		_w7490_
	);
	LUT2 #(
		.INIT('h1)
	) name6489 (
		\A[676] ,
		\A[677] ,
		_w7491_
	);
	LUT2 #(
		.INIT('h1)
	) name6490 (
		_w7490_,
		_w7491_,
		_w7492_
	);
	LUT2 #(
		.INIT('h8)
	) name6491 (
		\A[678] ,
		_w7492_,
		_w7493_
	);
	LUT2 #(
		.INIT('h1)
	) name6492 (
		_w7490_,
		_w7493_,
		_w7494_
	);
	LUT2 #(
		.INIT('h8)
	) name6493 (
		\A[673] ,
		\A[674] ,
		_w7495_
	);
	LUT2 #(
		.INIT('h1)
	) name6494 (
		\A[673] ,
		\A[674] ,
		_w7496_
	);
	LUT2 #(
		.INIT('h1)
	) name6495 (
		_w7495_,
		_w7496_,
		_w7497_
	);
	LUT2 #(
		.INIT('h8)
	) name6496 (
		\A[675] ,
		_w7497_,
		_w7498_
	);
	LUT2 #(
		.INIT('h1)
	) name6497 (
		_w7495_,
		_w7498_,
		_w7499_
	);
	LUT2 #(
		.INIT('h8)
	) name6498 (
		_w7494_,
		_w7499_,
		_w7500_
	);
	LUT2 #(
		.INIT('h1)
	) name6499 (
		_w7494_,
		_w7499_,
		_w7501_
	);
	LUT2 #(
		.INIT('h1)
	) name6500 (
		\A[675] ,
		_w7497_,
		_w7502_
	);
	LUT2 #(
		.INIT('h1)
	) name6501 (
		_w7498_,
		_w7502_,
		_w7503_
	);
	LUT2 #(
		.INIT('h1)
	) name6502 (
		\A[678] ,
		_w7492_,
		_w7504_
	);
	LUT2 #(
		.INIT('h1)
	) name6503 (
		_w7493_,
		_w7504_,
		_w7505_
	);
	LUT2 #(
		.INIT('h8)
	) name6504 (
		_w7503_,
		_w7505_,
		_w7506_
	);
	LUT2 #(
		.INIT('h1)
	) name6505 (
		_w7501_,
		_w7506_,
		_w7507_
	);
	LUT2 #(
		.INIT('h1)
	) name6506 (
		_w7500_,
		_w7507_,
		_w7508_
	);
	LUT2 #(
		.INIT('h1)
	) name6507 (
		_w7503_,
		_w7505_,
		_w7509_
	);
	LUT2 #(
		.INIT('h1)
	) name6508 (
		_w7506_,
		_w7509_,
		_w7510_
	);
	LUT2 #(
		.INIT('h1)
	) name6509 (
		_w7477_,
		_w7482_,
		_w7511_
	);
	LUT2 #(
		.INIT('h1)
	) name6510 (
		_w7483_,
		_w7511_,
		_w7512_
	);
	LUT2 #(
		.INIT('h8)
	) name6511 (
		_w7510_,
		_w7512_,
		_w7513_
	);
	LUT2 #(
		.INIT('h2)
	) name6512 (
		_w7484_,
		_w7485_,
		_w7514_
	);
	LUT2 #(
		.INIT('h2)
	) name6513 (
		_w7513_,
		_w7514_,
		_w7515_
	);
	LUT2 #(
		.INIT('h1)
	) name6514 (
		_w7500_,
		_w7501_,
		_w7516_
	);
	LUT2 #(
		.INIT('h2)
	) name6515 (
		_w7506_,
		_w7516_,
		_w7517_
	);
	LUT2 #(
		.INIT('h4)
	) name6516 (
		_w7506_,
		_w7516_,
		_w7518_
	);
	LUT2 #(
		.INIT('h1)
	) name6517 (
		_w7517_,
		_w7518_,
		_w7519_
	);
	LUT2 #(
		.INIT('h2)
	) name6518 (
		_w7515_,
		_w7519_,
		_w7520_
	);
	LUT2 #(
		.INIT('h4)
	) name6519 (
		_w7515_,
		_w7519_,
		_w7521_
	);
	LUT2 #(
		.INIT('h1)
	) name6520 (
		_w7484_,
		_w7487_,
		_w7522_
	);
	LUT2 #(
		.INIT('h2)
	) name6521 (
		_w7485_,
		_w7522_,
		_w7523_
	);
	LUT2 #(
		.INIT('h4)
	) name6522 (
		_w7485_,
		_w7522_,
		_w7524_
	);
	LUT2 #(
		.INIT('h1)
	) name6523 (
		_w7523_,
		_w7524_,
		_w7525_
	);
	LUT2 #(
		.INIT('h4)
	) name6524 (
		_w7521_,
		_w7525_,
		_w7526_
	);
	LUT2 #(
		.INIT('h1)
	) name6525 (
		_w7520_,
		_w7526_,
		_w7527_
	);
	LUT2 #(
		.INIT('h2)
	) name6526 (
		_w7508_,
		_w7527_,
		_w7528_
	);
	LUT2 #(
		.INIT('h4)
	) name6527 (
		_w7508_,
		_w7527_,
		_w7529_
	);
	LUT2 #(
		.INIT('h1)
	) name6528 (
		_w7528_,
		_w7529_,
		_w7530_
	);
	LUT2 #(
		.INIT('h8)
	) name6529 (
		_w7489_,
		_w7530_,
		_w7531_
	);
	LUT2 #(
		.INIT('h1)
	) name6530 (
		_w7489_,
		_w7530_,
		_w7532_
	);
	LUT2 #(
		.INIT('h1)
	) name6531 (
		_w7531_,
		_w7532_,
		_w7533_
	);
	LUT2 #(
		.INIT('h1)
	) name6532 (
		_w7470_,
		_w7533_,
		_w7534_
	);
	LUT2 #(
		.INIT('h8)
	) name6533 (
		_w7470_,
		_w7533_,
		_w7535_
	);
	LUT2 #(
		.INIT('h1)
	) name6534 (
		_w7510_,
		_w7512_,
		_w7536_
	);
	LUT2 #(
		.INIT('h1)
	) name6535 (
		_w7513_,
		_w7536_,
		_w7537_
	);
	LUT2 #(
		.INIT('h1)
	) name6536 (
		_w7447_,
		_w7449_,
		_w7538_
	);
	LUT2 #(
		.INIT('h1)
	) name6537 (
		_w7450_,
		_w7538_,
		_w7539_
	);
	LUT2 #(
		.INIT('h8)
	) name6538 (
		_w7537_,
		_w7539_,
		_w7540_
	);
	LUT2 #(
		.INIT('h1)
	) name6539 (
		_w7520_,
		_w7521_,
		_w7541_
	);
	LUT2 #(
		.INIT('h8)
	) name6540 (
		_w7525_,
		_w7541_,
		_w7542_
	);
	LUT2 #(
		.INIT('h1)
	) name6541 (
		_w7525_,
		_w7541_,
		_w7543_
	);
	LUT2 #(
		.INIT('h1)
	) name6542 (
		_w7542_,
		_w7543_,
		_w7544_
	);
	LUT2 #(
		.INIT('h8)
	) name6543 (
		_w7540_,
		_w7544_,
		_w7545_
	);
	LUT2 #(
		.INIT('h1)
	) name6544 (
		_w7540_,
		_w7544_,
		_w7546_
	);
	LUT2 #(
		.INIT('h1)
	) name6545 (
		_w7457_,
		_w7458_,
		_w7547_
	);
	LUT2 #(
		.INIT('h8)
	) name6546 (
		_w7462_,
		_w7547_,
		_w7548_
	);
	LUT2 #(
		.INIT('h1)
	) name6547 (
		_w7462_,
		_w7547_,
		_w7549_
	);
	LUT2 #(
		.INIT('h1)
	) name6548 (
		_w7548_,
		_w7549_,
		_w7550_
	);
	LUT2 #(
		.INIT('h4)
	) name6549 (
		_w7546_,
		_w7550_,
		_w7551_
	);
	LUT2 #(
		.INIT('h1)
	) name6550 (
		_w7545_,
		_w7551_,
		_w7552_
	);
	LUT2 #(
		.INIT('h1)
	) name6551 (
		_w7535_,
		_w7552_,
		_w7553_
	);
	LUT2 #(
		.INIT('h1)
	) name6552 (
		_w7534_,
		_w7553_,
		_w7554_
	);
	LUT2 #(
		.INIT('h1)
	) name6553 (
		_w7489_,
		_w7529_,
		_w7555_
	);
	LUT2 #(
		.INIT('h1)
	) name6554 (
		_w7528_,
		_w7555_,
		_w7556_
	);
	LUT2 #(
		.INIT('h1)
	) name6555 (
		_w7554_,
		_w7556_,
		_w7557_
	);
	LUT2 #(
		.INIT('h8)
	) name6556 (
		_w7554_,
		_w7556_,
		_w7558_
	);
	LUT2 #(
		.INIT('h1)
	) name6557 (
		_w7426_,
		_w7466_,
		_w7559_
	);
	LUT2 #(
		.INIT('h1)
	) name6558 (
		_w7465_,
		_w7559_,
		_w7560_
	);
	LUT2 #(
		.INIT('h1)
	) name6559 (
		_w7558_,
		_w7560_,
		_w7561_
	);
	LUT2 #(
		.INIT('h1)
	) name6560 (
		_w7557_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('h8)
	) name6561 (
		\A[682] ,
		\A[683] ,
		_w7563_
	);
	LUT2 #(
		.INIT('h8)
	) name6562 (
		\A[679] ,
		\A[680] ,
		_w7564_
	);
	LUT2 #(
		.INIT('h1)
	) name6563 (
		\A[679] ,
		\A[680] ,
		_w7565_
	);
	LUT2 #(
		.INIT('h1)
	) name6564 (
		_w7564_,
		_w7565_,
		_w7566_
	);
	LUT2 #(
		.INIT('h8)
	) name6565 (
		\A[681] ,
		_w7566_,
		_w7567_
	);
	LUT2 #(
		.INIT('h1)
	) name6566 (
		\A[681] ,
		_w7566_,
		_w7568_
	);
	LUT2 #(
		.INIT('h1)
	) name6567 (
		_w7567_,
		_w7568_,
		_w7569_
	);
	LUT2 #(
		.INIT('h1)
	) name6568 (
		\A[682] ,
		\A[683] ,
		_w7570_
	);
	LUT2 #(
		.INIT('h1)
	) name6569 (
		_w7563_,
		_w7570_,
		_w7571_
	);
	LUT2 #(
		.INIT('h8)
	) name6570 (
		\A[684] ,
		_w7571_,
		_w7572_
	);
	LUT2 #(
		.INIT('h1)
	) name6571 (
		\A[684] ,
		_w7571_,
		_w7573_
	);
	LUT2 #(
		.INIT('h1)
	) name6572 (
		_w7572_,
		_w7573_,
		_w7574_
	);
	LUT2 #(
		.INIT('h8)
	) name6573 (
		_w7569_,
		_w7574_,
		_w7575_
	);
	LUT2 #(
		.INIT('h8)
	) name6574 (
		_w7563_,
		_w7575_,
		_w7576_
	);
	LUT2 #(
		.INIT('h1)
	) name6575 (
		_w7564_,
		_w7567_,
		_w7577_
	);
	LUT2 #(
		.INIT('h1)
	) name6576 (
		_w7563_,
		_w7572_,
		_w7578_
	);
	LUT2 #(
		.INIT('h4)
	) name6577 (
		_w7575_,
		_w7578_,
		_w7579_
	);
	LUT2 #(
		.INIT('h1)
	) name6578 (
		_w7577_,
		_w7579_,
		_w7580_
	);
	LUT2 #(
		.INIT('h1)
	) name6579 (
		_w7576_,
		_w7580_,
		_w7581_
	);
	LUT2 #(
		.INIT('h8)
	) name6580 (
		\A[688] ,
		\A[689] ,
		_w7582_
	);
	LUT2 #(
		.INIT('h1)
	) name6581 (
		\A[688] ,
		\A[689] ,
		_w7583_
	);
	LUT2 #(
		.INIT('h1)
	) name6582 (
		_w7582_,
		_w7583_,
		_w7584_
	);
	LUT2 #(
		.INIT('h8)
	) name6583 (
		\A[690] ,
		_w7584_,
		_w7585_
	);
	LUT2 #(
		.INIT('h1)
	) name6584 (
		_w7582_,
		_w7585_,
		_w7586_
	);
	LUT2 #(
		.INIT('h8)
	) name6585 (
		\A[685] ,
		\A[686] ,
		_w7587_
	);
	LUT2 #(
		.INIT('h1)
	) name6586 (
		\A[685] ,
		\A[686] ,
		_w7588_
	);
	LUT2 #(
		.INIT('h1)
	) name6587 (
		_w7587_,
		_w7588_,
		_w7589_
	);
	LUT2 #(
		.INIT('h8)
	) name6588 (
		\A[687] ,
		_w7589_,
		_w7590_
	);
	LUT2 #(
		.INIT('h1)
	) name6589 (
		_w7587_,
		_w7590_,
		_w7591_
	);
	LUT2 #(
		.INIT('h8)
	) name6590 (
		_w7586_,
		_w7591_,
		_w7592_
	);
	LUT2 #(
		.INIT('h1)
	) name6591 (
		_w7586_,
		_w7591_,
		_w7593_
	);
	LUT2 #(
		.INIT('h1)
	) name6592 (
		\A[687] ,
		_w7589_,
		_w7594_
	);
	LUT2 #(
		.INIT('h1)
	) name6593 (
		_w7590_,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('h1)
	) name6594 (
		\A[690] ,
		_w7584_,
		_w7596_
	);
	LUT2 #(
		.INIT('h1)
	) name6595 (
		_w7585_,
		_w7596_,
		_w7597_
	);
	LUT2 #(
		.INIT('h8)
	) name6596 (
		_w7595_,
		_w7597_,
		_w7598_
	);
	LUT2 #(
		.INIT('h1)
	) name6597 (
		_w7593_,
		_w7598_,
		_w7599_
	);
	LUT2 #(
		.INIT('h1)
	) name6598 (
		_w7592_,
		_w7599_,
		_w7600_
	);
	LUT2 #(
		.INIT('h1)
	) name6599 (
		_w7595_,
		_w7597_,
		_w7601_
	);
	LUT2 #(
		.INIT('h1)
	) name6600 (
		_w7598_,
		_w7601_,
		_w7602_
	);
	LUT2 #(
		.INIT('h1)
	) name6601 (
		_w7569_,
		_w7574_,
		_w7603_
	);
	LUT2 #(
		.INIT('h1)
	) name6602 (
		_w7575_,
		_w7603_,
		_w7604_
	);
	LUT2 #(
		.INIT('h8)
	) name6603 (
		_w7602_,
		_w7604_,
		_w7605_
	);
	LUT2 #(
		.INIT('h2)
	) name6604 (
		_w7576_,
		_w7577_,
		_w7606_
	);
	LUT2 #(
		.INIT('h2)
	) name6605 (
		_w7605_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h1)
	) name6606 (
		_w7592_,
		_w7593_,
		_w7608_
	);
	LUT2 #(
		.INIT('h2)
	) name6607 (
		_w7598_,
		_w7608_,
		_w7609_
	);
	LUT2 #(
		.INIT('h4)
	) name6608 (
		_w7598_,
		_w7608_,
		_w7610_
	);
	LUT2 #(
		.INIT('h1)
	) name6609 (
		_w7609_,
		_w7610_,
		_w7611_
	);
	LUT2 #(
		.INIT('h2)
	) name6610 (
		_w7607_,
		_w7611_,
		_w7612_
	);
	LUT2 #(
		.INIT('h4)
	) name6611 (
		_w7607_,
		_w7611_,
		_w7613_
	);
	LUT2 #(
		.INIT('h1)
	) name6612 (
		_w7576_,
		_w7579_,
		_w7614_
	);
	LUT2 #(
		.INIT('h2)
	) name6613 (
		_w7577_,
		_w7614_,
		_w7615_
	);
	LUT2 #(
		.INIT('h4)
	) name6614 (
		_w7577_,
		_w7614_,
		_w7616_
	);
	LUT2 #(
		.INIT('h1)
	) name6615 (
		_w7615_,
		_w7616_,
		_w7617_
	);
	LUT2 #(
		.INIT('h4)
	) name6616 (
		_w7613_,
		_w7617_,
		_w7618_
	);
	LUT2 #(
		.INIT('h1)
	) name6617 (
		_w7612_,
		_w7618_,
		_w7619_
	);
	LUT2 #(
		.INIT('h2)
	) name6618 (
		_w7600_,
		_w7619_,
		_w7620_
	);
	LUT2 #(
		.INIT('h4)
	) name6619 (
		_w7600_,
		_w7619_,
		_w7621_
	);
	LUT2 #(
		.INIT('h1)
	) name6620 (
		_w7620_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('h8)
	) name6621 (
		_w7581_,
		_w7622_,
		_w7623_
	);
	LUT2 #(
		.INIT('h1)
	) name6622 (
		_w7581_,
		_w7622_,
		_w7624_
	);
	LUT2 #(
		.INIT('h1)
	) name6623 (
		_w7623_,
		_w7624_,
		_w7625_
	);
	LUT2 #(
		.INIT('h8)
	) name6624 (
		\A[694] ,
		\A[695] ,
		_w7626_
	);
	LUT2 #(
		.INIT('h8)
	) name6625 (
		\A[691] ,
		\A[692] ,
		_w7627_
	);
	LUT2 #(
		.INIT('h1)
	) name6626 (
		\A[691] ,
		\A[692] ,
		_w7628_
	);
	LUT2 #(
		.INIT('h1)
	) name6627 (
		_w7627_,
		_w7628_,
		_w7629_
	);
	LUT2 #(
		.INIT('h8)
	) name6628 (
		\A[693] ,
		_w7629_,
		_w7630_
	);
	LUT2 #(
		.INIT('h1)
	) name6629 (
		\A[693] ,
		_w7629_,
		_w7631_
	);
	LUT2 #(
		.INIT('h1)
	) name6630 (
		_w7630_,
		_w7631_,
		_w7632_
	);
	LUT2 #(
		.INIT('h1)
	) name6631 (
		\A[694] ,
		\A[695] ,
		_w7633_
	);
	LUT2 #(
		.INIT('h1)
	) name6632 (
		_w7626_,
		_w7633_,
		_w7634_
	);
	LUT2 #(
		.INIT('h8)
	) name6633 (
		\A[696] ,
		_w7634_,
		_w7635_
	);
	LUT2 #(
		.INIT('h1)
	) name6634 (
		\A[696] ,
		_w7634_,
		_w7636_
	);
	LUT2 #(
		.INIT('h1)
	) name6635 (
		_w7635_,
		_w7636_,
		_w7637_
	);
	LUT2 #(
		.INIT('h8)
	) name6636 (
		_w7632_,
		_w7637_,
		_w7638_
	);
	LUT2 #(
		.INIT('h8)
	) name6637 (
		_w7626_,
		_w7638_,
		_w7639_
	);
	LUT2 #(
		.INIT('h1)
	) name6638 (
		_w7627_,
		_w7630_,
		_w7640_
	);
	LUT2 #(
		.INIT('h1)
	) name6639 (
		_w7626_,
		_w7635_,
		_w7641_
	);
	LUT2 #(
		.INIT('h4)
	) name6640 (
		_w7638_,
		_w7641_,
		_w7642_
	);
	LUT2 #(
		.INIT('h1)
	) name6641 (
		_w7640_,
		_w7642_,
		_w7643_
	);
	LUT2 #(
		.INIT('h1)
	) name6642 (
		_w7639_,
		_w7643_,
		_w7644_
	);
	LUT2 #(
		.INIT('h8)
	) name6643 (
		\A[700] ,
		\A[701] ,
		_w7645_
	);
	LUT2 #(
		.INIT('h1)
	) name6644 (
		\A[700] ,
		\A[701] ,
		_w7646_
	);
	LUT2 #(
		.INIT('h1)
	) name6645 (
		_w7645_,
		_w7646_,
		_w7647_
	);
	LUT2 #(
		.INIT('h8)
	) name6646 (
		\A[702] ,
		_w7647_,
		_w7648_
	);
	LUT2 #(
		.INIT('h1)
	) name6647 (
		_w7645_,
		_w7648_,
		_w7649_
	);
	LUT2 #(
		.INIT('h8)
	) name6648 (
		\A[697] ,
		\A[698] ,
		_w7650_
	);
	LUT2 #(
		.INIT('h1)
	) name6649 (
		\A[697] ,
		\A[698] ,
		_w7651_
	);
	LUT2 #(
		.INIT('h1)
	) name6650 (
		_w7650_,
		_w7651_,
		_w7652_
	);
	LUT2 #(
		.INIT('h8)
	) name6651 (
		\A[699] ,
		_w7652_,
		_w7653_
	);
	LUT2 #(
		.INIT('h1)
	) name6652 (
		_w7650_,
		_w7653_,
		_w7654_
	);
	LUT2 #(
		.INIT('h8)
	) name6653 (
		_w7649_,
		_w7654_,
		_w7655_
	);
	LUT2 #(
		.INIT('h1)
	) name6654 (
		_w7649_,
		_w7654_,
		_w7656_
	);
	LUT2 #(
		.INIT('h1)
	) name6655 (
		\A[699] ,
		_w7652_,
		_w7657_
	);
	LUT2 #(
		.INIT('h1)
	) name6656 (
		_w7653_,
		_w7657_,
		_w7658_
	);
	LUT2 #(
		.INIT('h1)
	) name6657 (
		\A[702] ,
		_w7647_,
		_w7659_
	);
	LUT2 #(
		.INIT('h1)
	) name6658 (
		_w7648_,
		_w7659_,
		_w7660_
	);
	LUT2 #(
		.INIT('h8)
	) name6659 (
		_w7658_,
		_w7660_,
		_w7661_
	);
	LUT2 #(
		.INIT('h1)
	) name6660 (
		_w7656_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h1)
	) name6661 (
		_w7655_,
		_w7662_,
		_w7663_
	);
	LUT2 #(
		.INIT('h1)
	) name6662 (
		_w7658_,
		_w7660_,
		_w7664_
	);
	LUT2 #(
		.INIT('h1)
	) name6663 (
		_w7661_,
		_w7664_,
		_w7665_
	);
	LUT2 #(
		.INIT('h1)
	) name6664 (
		_w7632_,
		_w7637_,
		_w7666_
	);
	LUT2 #(
		.INIT('h1)
	) name6665 (
		_w7638_,
		_w7666_,
		_w7667_
	);
	LUT2 #(
		.INIT('h8)
	) name6666 (
		_w7665_,
		_w7667_,
		_w7668_
	);
	LUT2 #(
		.INIT('h2)
	) name6667 (
		_w7639_,
		_w7640_,
		_w7669_
	);
	LUT2 #(
		.INIT('h2)
	) name6668 (
		_w7668_,
		_w7669_,
		_w7670_
	);
	LUT2 #(
		.INIT('h1)
	) name6669 (
		_w7655_,
		_w7656_,
		_w7671_
	);
	LUT2 #(
		.INIT('h2)
	) name6670 (
		_w7661_,
		_w7671_,
		_w7672_
	);
	LUT2 #(
		.INIT('h4)
	) name6671 (
		_w7661_,
		_w7671_,
		_w7673_
	);
	LUT2 #(
		.INIT('h1)
	) name6672 (
		_w7672_,
		_w7673_,
		_w7674_
	);
	LUT2 #(
		.INIT('h2)
	) name6673 (
		_w7670_,
		_w7674_,
		_w7675_
	);
	LUT2 #(
		.INIT('h4)
	) name6674 (
		_w7670_,
		_w7674_,
		_w7676_
	);
	LUT2 #(
		.INIT('h1)
	) name6675 (
		_w7639_,
		_w7642_,
		_w7677_
	);
	LUT2 #(
		.INIT('h2)
	) name6676 (
		_w7640_,
		_w7677_,
		_w7678_
	);
	LUT2 #(
		.INIT('h4)
	) name6677 (
		_w7640_,
		_w7677_,
		_w7679_
	);
	LUT2 #(
		.INIT('h1)
	) name6678 (
		_w7678_,
		_w7679_,
		_w7680_
	);
	LUT2 #(
		.INIT('h4)
	) name6679 (
		_w7676_,
		_w7680_,
		_w7681_
	);
	LUT2 #(
		.INIT('h1)
	) name6680 (
		_w7675_,
		_w7681_,
		_w7682_
	);
	LUT2 #(
		.INIT('h2)
	) name6681 (
		_w7663_,
		_w7682_,
		_w7683_
	);
	LUT2 #(
		.INIT('h4)
	) name6682 (
		_w7663_,
		_w7682_,
		_w7684_
	);
	LUT2 #(
		.INIT('h1)
	) name6683 (
		_w7683_,
		_w7684_,
		_w7685_
	);
	LUT2 #(
		.INIT('h8)
	) name6684 (
		_w7644_,
		_w7685_,
		_w7686_
	);
	LUT2 #(
		.INIT('h1)
	) name6685 (
		_w7644_,
		_w7685_,
		_w7687_
	);
	LUT2 #(
		.INIT('h1)
	) name6686 (
		_w7686_,
		_w7687_,
		_w7688_
	);
	LUT2 #(
		.INIT('h1)
	) name6687 (
		_w7625_,
		_w7688_,
		_w7689_
	);
	LUT2 #(
		.INIT('h8)
	) name6688 (
		_w7625_,
		_w7688_,
		_w7690_
	);
	LUT2 #(
		.INIT('h1)
	) name6689 (
		_w7665_,
		_w7667_,
		_w7691_
	);
	LUT2 #(
		.INIT('h1)
	) name6690 (
		_w7668_,
		_w7691_,
		_w7692_
	);
	LUT2 #(
		.INIT('h1)
	) name6691 (
		_w7602_,
		_w7604_,
		_w7693_
	);
	LUT2 #(
		.INIT('h1)
	) name6692 (
		_w7605_,
		_w7693_,
		_w7694_
	);
	LUT2 #(
		.INIT('h8)
	) name6693 (
		_w7692_,
		_w7694_,
		_w7695_
	);
	LUT2 #(
		.INIT('h1)
	) name6694 (
		_w7675_,
		_w7676_,
		_w7696_
	);
	LUT2 #(
		.INIT('h8)
	) name6695 (
		_w7680_,
		_w7696_,
		_w7697_
	);
	LUT2 #(
		.INIT('h1)
	) name6696 (
		_w7680_,
		_w7696_,
		_w7698_
	);
	LUT2 #(
		.INIT('h1)
	) name6697 (
		_w7697_,
		_w7698_,
		_w7699_
	);
	LUT2 #(
		.INIT('h8)
	) name6698 (
		_w7695_,
		_w7699_,
		_w7700_
	);
	LUT2 #(
		.INIT('h1)
	) name6699 (
		_w7695_,
		_w7699_,
		_w7701_
	);
	LUT2 #(
		.INIT('h1)
	) name6700 (
		_w7612_,
		_w7613_,
		_w7702_
	);
	LUT2 #(
		.INIT('h8)
	) name6701 (
		_w7617_,
		_w7702_,
		_w7703_
	);
	LUT2 #(
		.INIT('h1)
	) name6702 (
		_w7617_,
		_w7702_,
		_w7704_
	);
	LUT2 #(
		.INIT('h1)
	) name6703 (
		_w7703_,
		_w7704_,
		_w7705_
	);
	LUT2 #(
		.INIT('h4)
	) name6704 (
		_w7701_,
		_w7705_,
		_w7706_
	);
	LUT2 #(
		.INIT('h1)
	) name6705 (
		_w7700_,
		_w7706_,
		_w7707_
	);
	LUT2 #(
		.INIT('h1)
	) name6706 (
		_w7690_,
		_w7707_,
		_w7708_
	);
	LUT2 #(
		.INIT('h1)
	) name6707 (
		_w7689_,
		_w7708_,
		_w7709_
	);
	LUT2 #(
		.INIT('h1)
	) name6708 (
		_w7644_,
		_w7684_,
		_w7710_
	);
	LUT2 #(
		.INIT('h1)
	) name6709 (
		_w7683_,
		_w7710_,
		_w7711_
	);
	LUT2 #(
		.INIT('h1)
	) name6710 (
		_w7709_,
		_w7711_,
		_w7712_
	);
	LUT2 #(
		.INIT('h8)
	) name6711 (
		_w7709_,
		_w7711_,
		_w7713_
	);
	LUT2 #(
		.INIT('h1)
	) name6712 (
		_w7712_,
		_w7713_,
		_w7714_
	);
	LUT2 #(
		.INIT('h1)
	) name6713 (
		_w7581_,
		_w7621_,
		_w7715_
	);
	LUT2 #(
		.INIT('h1)
	) name6714 (
		_w7620_,
		_w7715_,
		_w7716_
	);
	LUT2 #(
		.INIT('h2)
	) name6715 (
		_w7714_,
		_w7716_,
		_w7717_
	);
	LUT2 #(
		.INIT('h4)
	) name6716 (
		_w7714_,
		_w7716_,
		_w7718_
	);
	LUT2 #(
		.INIT('h1)
	) name6717 (
		_w7717_,
		_w7718_,
		_w7719_
	);
	LUT2 #(
		.INIT('h1)
	) name6718 (
		_w7557_,
		_w7558_,
		_w7720_
	);
	LUT2 #(
		.INIT('h4)
	) name6719 (
		_w7560_,
		_w7720_,
		_w7721_
	);
	LUT2 #(
		.INIT('h2)
	) name6720 (
		_w7560_,
		_w7720_,
		_w7722_
	);
	LUT2 #(
		.INIT('h1)
	) name6721 (
		_w7721_,
		_w7722_,
		_w7723_
	);
	LUT2 #(
		.INIT('h1)
	) name6722 (
		_w7719_,
		_w7723_,
		_w7724_
	);
	LUT2 #(
		.INIT('h8)
	) name6723 (
		_w7719_,
		_w7723_,
		_w7725_
	);
	LUT2 #(
		.INIT('h1)
	) name6724 (
		_w7534_,
		_w7535_,
		_w7726_
	);
	LUT2 #(
		.INIT('h4)
	) name6725 (
		_w7552_,
		_w7726_,
		_w7727_
	);
	LUT2 #(
		.INIT('h2)
	) name6726 (
		_w7552_,
		_w7726_,
		_w7728_
	);
	LUT2 #(
		.INIT('h1)
	) name6727 (
		_w7727_,
		_w7728_,
		_w7729_
	);
	LUT2 #(
		.INIT('h1)
	) name6728 (
		_w7689_,
		_w7690_,
		_w7730_
	);
	LUT2 #(
		.INIT('h4)
	) name6729 (
		_w7707_,
		_w7730_,
		_w7731_
	);
	LUT2 #(
		.INIT('h2)
	) name6730 (
		_w7707_,
		_w7730_,
		_w7732_
	);
	LUT2 #(
		.INIT('h1)
	) name6731 (
		_w7731_,
		_w7732_,
		_w7733_
	);
	LUT2 #(
		.INIT('h1)
	) name6732 (
		_w7729_,
		_w7733_,
		_w7734_
	);
	LUT2 #(
		.INIT('h8)
	) name6733 (
		_w7729_,
		_w7733_,
		_w7735_
	);
	LUT2 #(
		.INIT('h1)
	) name6734 (
		_w7692_,
		_w7694_,
		_w7736_
	);
	LUT2 #(
		.INIT('h1)
	) name6735 (
		_w7695_,
		_w7736_,
		_w7737_
	);
	LUT2 #(
		.INIT('h1)
	) name6736 (
		_w7537_,
		_w7539_,
		_w7738_
	);
	LUT2 #(
		.INIT('h1)
	) name6737 (
		_w7540_,
		_w7738_,
		_w7739_
	);
	LUT2 #(
		.INIT('h8)
	) name6738 (
		_w7737_,
		_w7739_,
		_w7740_
	);
	LUT2 #(
		.INIT('h1)
	) name6739 (
		_w7700_,
		_w7701_,
		_w7741_
	);
	LUT2 #(
		.INIT('h4)
	) name6740 (
		_w7705_,
		_w7741_,
		_w7742_
	);
	LUT2 #(
		.INIT('h2)
	) name6741 (
		_w7705_,
		_w7741_,
		_w7743_
	);
	LUT2 #(
		.INIT('h1)
	) name6742 (
		_w7742_,
		_w7743_,
		_w7744_
	);
	LUT2 #(
		.INIT('h2)
	) name6743 (
		_w7740_,
		_w7744_,
		_w7745_
	);
	LUT2 #(
		.INIT('h4)
	) name6744 (
		_w7740_,
		_w7744_,
		_w7746_
	);
	LUT2 #(
		.INIT('h1)
	) name6745 (
		_w7545_,
		_w7546_,
		_w7747_
	);
	LUT2 #(
		.INIT('h4)
	) name6746 (
		_w7550_,
		_w7747_,
		_w7748_
	);
	LUT2 #(
		.INIT('h2)
	) name6747 (
		_w7550_,
		_w7747_,
		_w7749_
	);
	LUT2 #(
		.INIT('h1)
	) name6748 (
		_w7748_,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('h1)
	) name6749 (
		_w7746_,
		_w7750_,
		_w7751_
	);
	LUT2 #(
		.INIT('h1)
	) name6750 (
		_w7745_,
		_w7751_,
		_w7752_
	);
	LUT2 #(
		.INIT('h4)
	) name6751 (
		_w7735_,
		_w7752_,
		_w7753_
	);
	LUT2 #(
		.INIT('h1)
	) name6752 (
		_w7734_,
		_w7753_,
		_w7754_
	);
	LUT2 #(
		.INIT('h1)
	) name6753 (
		_w7725_,
		_w7754_,
		_w7755_
	);
	LUT2 #(
		.INIT('h1)
	) name6754 (
		_w7724_,
		_w7755_,
		_w7756_
	);
	LUT2 #(
		.INIT('h2)
	) name6755 (
		_w7562_,
		_w7756_,
		_w7757_
	);
	LUT2 #(
		.INIT('h4)
	) name6756 (
		_w7562_,
		_w7756_,
		_w7758_
	);
	LUT2 #(
		.INIT('h1)
	) name6757 (
		_w7713_,
		_w7716_,
		_w7759_
	);
	LUT2 #(
		.INIT('h1)
	) name6758 (
		_w7712_,
		_w7759_,
		_w7760_
	);
	LUT2 #(
		.INIT('h4)
	) name6759 (
		_w7758_,
		_w7760_,
		_w7761_
	);
	LUT2 #(
		.INIT('h1)
	) name6760 (
		_w7757_,
		_w7761_,
		_w7762_
	);
	LUT2 #(
		.INIT('h4)
	) name6761 (
		_w7407_,
		_w7762_,
		_w7763_
	);
	LUT2 #(
		.INIT('h2)
	) name6762 (
		_w7407_,
		_w7762_,
		_w7764_
	);
	LUT2 #(
		.INIT('h1)
	) name6763 (
		_w7757_,
		_w7758_,
		_w7765_
	);
	LUT2 #(
		.INIT('h8)
	) name6764 (
		_w7760_,
		_w7765_,
		_w7766_
	);
	LUT2 #(
		.INIT('h1)
	) name6765 (
		_w7760_,
		_w7765_,
		_w7767_
	);
	LUT2 #(
		.INIT('h1)
	) name6766 (
		_w7766_,
		_w7767_,
		_w7768_
	);
	LUT2 #(
		.INIT('h1)
	) name6767 (
		_w7402_,
		_w7403_,
		_w7769_
	);
	LUT2 #(
		.INIT('h4)
	) name6768 (
		_w7405_,
		_w7769_,
		_w7770_
	);
	LUT2 #(
		.INIT('h2)
	) name6769 (
		_w7405_,
		_w7769_,
		_w7771_
	);
	LUT2 #(
		.INIT('h1)
	) name6770 (
		_w7770_,
		_w7771_,
		_w7772_
	);
	LUT2 #(
		.INIT('h4)
	) name6771 (
		_w7768_,
		_w7772_,
		_w7773_
	);
	LUT2 #(
		.INIT('h2)
	) name6772 (
		_w7768_,
		_w7772_,
		_w7774_
	);
	LUT2 #(
		.INIT('h1)
	) name6773 (
		_w7367_,
		_w7368_,
		_w7775_
	);
	LUT2 #(
		.INIT('h4)
	) name6774 (
		_w7397_,
		_w7775_,
		_w7776_
	);
	LUT2 #(
		.INIT('h2)
	) name6775 (
		_w7397_,
		_w7775_,
		_w7777_
	);
	LUT2 #(
		.INIT('h1)
	) name6776 (
		_w7776_,
		_w7777_,
		_w7778_
	);
	LUT2 #(
		.INIT('h1)
	) name6777 (
		_w7724_,
		_w7725_,
		_w7779_
	);
	LUT2 #(
		.INIT('h4)
	) name6778 (
		_w7754_,
		_w7779_,
		_w7780_
	);
	LUT2 #(
		.INIT('h2)
	) name6779 (
		_w7754_,
		_w7779_,
		_w7781_
	);
	LUT2 #(
		.INIT('h1)
	) name6780 (
		_w7780_,
		_w7781_,
		_w7782_
	);
	LUT2 #(
		.INIT('h1)
	) name6781 (
		_w7778_,
		_w7782_,
		_w7783_
	);
	LUT2 #(
		.INIT('h8)
	) name6782 (
		_w7778_,
		_w7782_,
		_w7784_
	);
	LUT2 #(
		.INIT('h1)
	) name6783 (
		_w7734_,
		_w7735_,
		_w7785_
	);
	LUT2 #(
		.INIT('h4)
	) name6784 (
		_w7752_,
		_w7785_,
		_w7786_
	);
	LUT2 #(
		.INIT('h2)
	) name6785 (
		_w7752_,
		_w7785_,
		_w7787_
	);
	LUT2 #(
		.INIT('h1)
	) name6786 (
		_w7786_,
		_w7787_,
		_w7788_
	);
	LUT2 #(
		.INIT('h1)
	) name6787 (
		_w7377_,
		_w7378_,
		_w7789_
	);
	LUT2 #(
		.INIT('h4)
	) name6788 (
		_w7395_,
		_w7789_,
		_w7790_
	);
	LUT2 #(
		.INIT('h2)
	) name6789 (
		_w7395_,
		_w7789_,
		_w7791_
	);
	LUT2 #(
		.INIT('h1)
	) name6790 (
		_w7790_,
		_w7791_,
		_w7792_
	);
	LUT2 #(
		.INIT('h1)
	) name6791 (
		_w7788_,
		_w7792_,
		_w7793_
	);
	LUT2 #(
		.INIT('h8)
	) name6792 (
		_w7788_,
		_w7792_,
		_w7794_
	);
	LUT2 #(
		.INIT('h1)
	) name6793 (
		_w7380_,
		_w7382_,
		_w7795_
	);
	LUT2 #(
		.INIT('h1)
	) name6794 (
		_w7383_,
		_w7795_,
		_w7796_
	);
	LUT2 #(
		.INIT('h1)
	) name6795 (
		_w7737_,
		_w7739_,
		_w7797_
	);
	LUT2 #(
		.INIT('h1)
	) name6796 (
		_w7740_,
		_w7797_,
		_w7798_
	);
	LUT2 #(
		.INIT('h8)
	) name6797 (
		_w7796_,
		_w7798_,
		_w7799_
	);
	LUT2 #(
		.INIT('h1)
	) name6798 (
		_w7388_,
		_w7389_,
		_w7800_
	);
	LUT2 #(
		.INIT('h4)
	) name6799 (
		_w7393_,
		_w7800_,
		_w7801_
	);
	LUT2 #(
		.INIT('h2)
	) name6800 (
		_w7393_,
		_w7800_,
		_w7802_
	);
	LUT2 #(
		.INIT('h1)
	) name6801 (
		_w7801_,
		_w7802_,
		_w7803_
	);
	LUT2 #(
		.INIT('h2)
	) name6802 (
		_w7799_,
		_w7803_,
		_w7804_
	);
	LUT2 #(
		.INIT('h4)
	) name6803 (
		_w7799_,
		_w7803_,
		_w7805_
	);
	LUT2 #(
		.INIT('h1)
	) name6804 (
		_w7745_,
		_w7746_,
		_w7806_
	);
	LUT2 #(
		.INIT('h4)
	) name6805 (
		_w7750_,
		_w7806_,
		_w7807_
	);
	LUT2 #(
		.INIT('h2)
	) name6806 (
		_w7750_,
		_w7806_,
		_w7808_
	);
	LUT2 #(
		.INIT('h1)
	) name6807 (
		_w7807_,
		_w7808_,
		_w7809_
	);
	LUT2 #(
		.INIT('h4)
	) name6808 (
		_w7805_,
		_w7809_,
		_w7810_
	);
	LUT2 #(
		.INIT('h1)
	) name6809 (
		_w7804_,
		_w7810_,
		_w7811_
	);
	LUT2 #(
		.INIT('h4)
	) name6810 (
		_w7794_,
		_w7811_,
		_w7812_
	);
	LUT2 #(
		.INIT('h1)
	) name6811 (
		_w7793_,
		_w7812_,
		_w7813_
	);
	LUT2 #(
		.INIT('h4)
	) name6812 (
		_w7784_,
		_w7813_,
		_w7814_
	);
	LUT2 #(
		.INIT('h1)
	) name6813 (
		_w7783_,
		_w7814_,
		_w7815_
	);
	LUT2 #(
		.INIT('h1)
	) name6814 (
		_w7774_,
		_w7815_,
		_w7816_
	);
	LUT2 #(
		.INIT('h1)
	) name6815 (
		_w7773_,
		_w7816_,
		_w7817_
	);
	LUT2 #(
		.INIT('h1)
	) name6816 (
		_w7764_,
		_w7817_,
		_w7818_
	);
	LUT2 #(
		.INIT('h1)
	) name6817 (
		_w7763_,
		_w7818_,
		_w7819_
	);
	LUT2 #(
		.INIT('h1)
	) name6818 (
		_w7060_,
		_w7819_,
		_w7820_
	);
	LUT2 #(
		.INIT('h8)
	) name6819 (
		_w7060_,
		_w7819_,
		_w7821_
	);
	LUT2 #(
		.INIT('h1)
	) name6820 (
		_w7004_,
		_w7005_,
		_w7822_
	);
	LUT2 #(
		.INIT('h4)
	) name6821 (
		_w7058_,
		_w7822_,
		_w7823_
	);
	LUT2 #(
		.INIT('h2)
	) name6822 (
		_w7058_,
		_w7822_,
		_w7824_
	);
	LUT2 #(
		.INIT('h1)
	) name6823 (
		_w7823_,
		_w7824_,
		_w7825_
	);
	LUT2 #(
		.INIT('h1)
	) name6824 (
		_w7763_,
		_w7764_,
		_w7826_
	);
	LUT2 #(
		.INIT('h4)
	) name6825 (
		_w7817_,
		_w7826_,
		_w7827_
	);
	LUT2 #(
		.INIT('h2)
	) name6826 (
		_w7817_,
		_w7826_,
		_w7828_
	);
	LUT2 #(
		.INIT('h1)
	) name6827 (
		_w7827_,
		_w7828_,
		_w7829_
	);
	LUT2 #(
		.INIT('h1)
	) name6828 (
		_w7825_,
		_w7829_,
		_w7830_
	);
	LUT2 #(
		.INIT('h8)
	) name6829 (
		_w7825_,
		_w7829_,
		_w7831_
	);
	LUT2 #(
		.INIT('h1)
	) name6830 (
		_w7014_,
		_w7015_,
		_w7832_
	);
	LUT2 #(
		.INIT('h4)
	) name6831 (
		_w7056_,
		_w7832_,
		_w7833_
	);
	LUT2 #(
		.INIT('h2)
	) name6832 (
		_w7056_,
		_w7832_,
		_w7834_
	);
	LUT2 #(
		.INIT('h1)
	) name6833 (
		_w7833_,
		_w7834_,
		_w7835_
	);
	LUT2 #(
		.INIT('h1)
	) name6834 (
		_w7773_,
		_w7774_,
		_w7836_
	);
	LUT2 #(
		.INIT('h4)
	) name6835 (
		_w7815_,
		_w7836_,
		_w7837_
	);
	LUT2 #(
		.INIT('h2)
	) name6836 (
		_w7815_,
		_w7836_,
		_w7838_
	);
	LUT2 #(
		.INIT('h1)
	) name6837 (
		_w7837_,
		_w7838_,
		_w7839_
	);
	LUT2 #(
		.INIT('h2)
	) name6838 (
		_w7835_,
		_w7839_,
		_w7840_
	);
	LUT2 #(
		.INIT('h4)
	) name6839 (
		_w7835_,
		_w7839_,
		_w7841_
	);
	LUT2 #(
		.INIT('h1)
	) name6840 (
		_w7024_,
		_w7025_,
		_w7842_
	);
	LUT2 #(
		.INIT('h4)
	) name6841 (
		_w7054_,
		_w7842_,
		_w7843_
	);
	LUT2 #(
		.INIT('h2)
	) name6842 (
		_w7054_,
		_w7842_,
		_w7844_
	);
	LUT2 #(
		.INIT('h1)
	) name6843 (
		_w7843_,
		_w7844_,
		_w7845_
	);
	LUT2 #(
		.INIT('h1)
	) name6844 (
		_w7783_,
		_w7784_,
		_w7846_
	);
	LUT2 #(
		.INIT('h8)
	) name6845 (
		_w7813_,
		_w7846_,
		_w7847_
	);
	LUT2 #(
		.INIT('h1)
	) name6846 (
		_w7813_,
		_w7846_,
		_w7848_
	);
	LUT2 #(
		.INIT('h1)
	) name6847 (
		_w7847_,
		_w7848_,
		_w7849_
	);
	LUT2 #(
		.INIT('h2)
	) name6848 (
		_w7845_,
		_w7849_,
		_w7850_
	);
	LUT2 #(
		.INIT('h4)
	) name6849 (
		_w7845_,
		_w7849_,
		_w7851_
	);
	LUT2 #(
		.INIT('h1)
	) name6850 (
		_w7793_,
		_w7794_,
		_w7852_
	);
	LUT2 #(
		.INIT('h4)
	) name6851 (
		_w7811_,
		_w7852_,
		_w7853_
	);
	LUT2 #(
		.INIT('h2)
	) name6852 (
		_w7811_,
		_w7852_,
		_w7854_
	);
	LUT2 #(
		.INIT('h1)
	) name6853 (
		_w7853_,
		_w7854_,
		_w7855_
	);
	LUT2 #(
		.INIT('h1)
	) name6854 (
		_w7034_,
		_w7035_,
		_w7856_
	);
	LUT2 #(
		.INIT('h4)
	) name6855 (
		_w7052_,
		_w7856_,
		_w7857_
	);
	LUT2 #(
		.INIT('h2)
	) name6856 (
		_w7052_,
		_w7856_,
		_w7858_
	);
	LUT2 #(
		.INIT('h1)
	) name6857 (
		_w7857_,
		_w7858_,
		_w7859_
	);
	LUT2 #(
		.INIT('h1)
	) name6858 (
		_w7855_,
		_w7859_,
		_w7860_
	);
	LUT2 #(
		.INIT('h8)
	) name6859 (
		_w7855_,
		_w7859_,
		_w7861_
	);
	LUT2 #(
		.INIT('h1)
	) name6860 (
		_w7037_,
		_w7039_,
		_w7862_
	);
	LUT2 #(
		.INIT('h1)
	) name6861 (
		_w7040_,
		_w7862_,
		_w7863_
	);
	LUT2 #(
		.INIT('h1)
	) name6862 (
		_w7796_,
		_w7798_,
		_w7864_
	);
	LUT2 #(
		.INIT('h1)
	) name6863 (
		_w7799_,
		_w7864_,
		_w7865_
	);
	LUT2 #(
		.INIT('h8)
	) name6864 (
		_w7863_,
		_w7865_,
		_w7866_
	);
	LUT2 #(
		.INIT('h1)
	) name6865 (
		_w7045_,
		_w7046_,
		_w7867_
	);
	LUT2 #(
		.INIT('h4)
	) name6866 (
		_w7050_,
		_w7867_,
		_w7868_
	);
	LUT2 #(
		.INIT('h2)
	) name6867 (
		_w7050_,
		_w7867_,
		_w7869_
	);
	LUT2 #(
		.INIT('h1)
	) name6868 (
		_w7868_,
		_w7869_,
		_w7870_
	);
	LUT2 #(
		.INIT('h8)
	) name6869 (
		_w7866_,
		_w7870_,
		_w7871_
	);
	LUT2 #(
		.INIT('h1)
	) name6870 (
		_w7866_,
		_w7870_,
		_w7872_
	);
	LUT2 #(
		.INIT('h1)
	) name6871 (
		_w7804_,
		_w7805_,
		_w7873_
	);
	LUT2 #(
		.INIT('h4)
	) name6872 (
		_w7809_,
		_w7873_,
		_w7874_
	);
	LUT2 #(
		.INIT('h2)
	) name6873 (
		_w7809_,
		_w7873_,
		_w7875_
	);
	LUT2 #(
		.INIT('h1)
	) name6874 (
		_w7874_,
		_w7875_,
		_w7876_
	);
	LUT2 #(
		.INIT('h1)
	) name6875 (
		_w7872_,
		_w7876_,
		_w7877_
	);
	LUT2 #(
		.INIT('h1)
	) name6876 (
		_w7871_,
		_w7877_,
		_w7878_
	);
	LUT2 #(
		.INIT('h4)
	) name6877 (
		_w7861_,
		_w7878_,
		_w7879_
	);
	LUT2 #(
		.INIT('h1)
	) name6878 (
		_w7860_,
		_w7879_,
		_w7880_
	);
	LUT2 #(
		.INIT('h1)
	) name6879 (
		_w7851_,
		_w7880_,
		_w7881_
	);
	LUT2 #(
		.INIT('h1)
	) name6880 (
		_w7850_,
		_w7881_,
		_w7882_
	);
	LUT2 #(
		.INIT('h1)
	) name6881 (
		_w7841_,
		_w7882_,
		_w7883_
	);
	LUT2 #(
		.INIT('h1)
	) name6882 (
		_w7840_,
		_w7883_,
		_w7884_
	);
	LUT2 #(
		.INIT('h1)
	) name6883 (
		_w7831_,
		_w7884_,
		_w7885_
	);
	LUT2 #(
		.INIT('h1)
	) name6884 (
		_w7830_,
		_w7885_,
		_w7886_
	);
	LUT2 #(
		.INIT('h4)
	) name6885 (
		_w7821_,
		_w7886_,
		_w7887_
	);
	LUT2 #(
		.INIT('h1)
	) name6886 (
		_w7820_,
		_w7887_,
		_w7888_
	);
	LUT2 #(
		.INIT('h8)
	) name6887 (
		\A[562] ,
		\A[563] ,
		_w7889_
	);
	LUT2 #(
		.INIT('h8)
	) name6888 (
		\A[559] ,
		\A[560] ,
		_w7890_
	);
	LUT2 #(
		.INIT('h1)
	) name6889 (
		\A[559] ,
		\A[560] ,
		_w7891_
	);
	LUT2 #(
		.INIT('h1)
	) name6890 (
		_w7890_,
		_w7891_,
		_w7892_
	);
	LUT2 #(
		.INIT('h8)
	) name6891 (
		\A[561] ,
		_w7892_,
		_w7893_
	);
	LUT2 #(
		.INIT('h1)
	) name6892 (
		\A[561] ,
		_w7892_,
		_w7894_
	);
	LUT2 #(
		.INIT('h1)
	) name6893 (
		_w7893_,
		_w7894_,
		_w7895_
	);
	LUT2 #(
		.INIT('h1)
	) name6894 (
		\A[562] ,
		\A[563] ,
		_w7896_
	);
	LUT2 #(
		.INIT('h1)
	) name6895 (
		_w7889_,
		_w7896_,
		_w7897_
	);
	LUT2 #(
		.INIT('h8)
	) name6896 (
		\A[564] ,
		_w7897_,
		_w7898_
	);
	LUT2 #(
		.INIT('h1)
	) name6897 (
		\A[564] ,
		_w7897_,
		_w7899_
	);
	LUT2 #(
		.INIT('h1)
	) name6898 (
		_w7898_,
		_w7899_,
		_w7900_
	);
	LUT2 #(
		.INIT('h8)
	) name6899 (
		_w7895_,
		_w7900_,
		_w7901_
	);
	LUT2 #(
		.INIT('h8)
	) name6900 (
		_w7889_,
		_w7901_,
		_w7902_
	);
	LUT2 #(
		.INIT('h1)
	) name6901 (
		_w7890_,
		_w7893_,
		_w7903_
	);
	LUT2 #(
		.INIT('h1)
	) name6902 (
		_w7889_,
		_w7898_,
		_w7904_
	);
	LUT2 #(
		.INIT('h4)
	) name6903 (
		_w7901_,
		_w7904_,
		_w7905_
	);
	LUT2 #(
		.INIT('h1)
	) name6904 (
		_w7903_,
		_w7905_,
		_w7906_
	);
	LUT2 #(
		.INIT('h1)
	) name6905 (
		_w7902_,
		_w7906_,
		_w7907_
	);
	LUT2 #(
		.INIT('h8)
	) name6906 (
		\A[568] ,
		\A[569] ,
		_w7908_
	);
	LUT2 #(
		.INIT('h1)
	) name6907 (
		\A[568] ,
		\A[569] ,
		_w7909_
	);
	LUT2 #(
		.INIT('h1)
	) name6908 (
		_w7908_,
		_w7909_,
		_w7910_
	);
	LUT2 #(
		.INIT('h8)
	) name6909 (
		\A[570] ,
		_w7910_,
		_w7911_
	);
	LUT2 #(
		.INIT('h1)
	) name6910 (
		_w7908_,
		_w7911_,
		_w7912_
	);
	LUT2 #(
		.INIT('h8)
	) name6911 (
		\A[565] ,
		\A[566] ,
		_w7913_
	);
	LUT2 #(
		.INIT('h1)
	) name6912 (
		\A[565] ,
		\A[566] ,
		_w7914_
	);
	LUT2 #(
		.INIT('h1)
	) name6913 (
		_w7913_,
		_w7914_,
		_w7915_
	);
	LUT2 #(
		.INIT('h8)
	) name6914 (
		\A[567] ,
		_w7915_,
		_w7916_
	);
	LUT2 #(
		.INIT('h1)
	) name6915 (
		_w7913_,
		_w7916_,
		_w7917_
	);
	LUT2 #(
		.INIT('h8)
	) name6916 (
		_w7912_,
		_w7917_,
		_w7918_
	);
	LUT2 #(
		.INIT('h1)
	) name6917 (
		_w7912_,
		_w7917_,
		_w7919_
	);
	LUT2 #(
		.INIT('h1)
	) name6918 (
		\A[567] ,
		_w7915_,
		_w7920_
	);
	LUT2 #(
		.INIT('h1)
	) name6919 (
		_w7916_,
		_w7920_,
		_w7921_
	);
	LUT2 #(
		.INIT('h1)
	) name6920 (
		\A[570] ,
		_w7910_,
		_w7922_
	);
	LUT2 #(
		.INIT('h1)
	) name6921 (
		_w7911_,
		_w7922_,
		_w7923_
	);
	LUT2 #(
		.INIT('h8)
	) name6922 (
		_w7921_,
		_w7923_,
		_w7924_
	);
	LUT2 #(
		.INIT('h1)
	) name6923 (
		_w7919_,
		_w7924_,
		_w7925_
	);
	LUT2 #(
		.INIT('h1)
	) name6924 (
		_w7918_,
		_w7925_,
		_w7926_
	);
	LUT2 #(
		.INIT('h1)
	) name6925 (
		_w7921_,
		_w7923_,
		_w7927_
	);
	LUT2 #(
		.INIT('h1)
	) name6926 (
		_w7924_,
		_w7927_,
		_w7928_
	);
	LUT2 #(
		.INIT('h1)
	) name6927 (
		_w7895_,
		_w7900_,
		_w7929_
	);
	LUT2 #(
		.INIT('h1)
	) name6928 (
		_w7901_,
		_w7929_,
		_w7930_
	);
	LUT2 #(
		.INIT('h8)
	) name6929 (
		_w7928_,
		_w7930_,
		_w7931_
	);
	LUT2 #(
		.INIT('h2)
	) name6930 (
		_w7902_,
		_w7903_,
		_w7932_
	);
	LUT2 #(
		.INIT('h2)
	) name6931 (
		_w7931_,
		_w7932_,
		_w7933_
	);
	LUT2 #(
		.INIT('h1)
	) name6932 (
		_w7918_,
		_w7919_,
		_w7934_
	);
	LUT2 #(
		.INIT('h2)
	) name6933 (
		_w7924_,
		_w7934_,
		_w7935_
	);
	LUT2 #(
		.INIT('h4)
	) name6934 (
		_w7924_,
		_w7934_,
		_w7936_
	);
	LUT2 #(
		.INIT('h1)
	) name6935 (
		_w7935_,
		_w7936_,
		_w7937_
	);
	LUT2 #(
		.INIT('h2)
	) name6936 (
		_w7933_,
		_w7937_,
		_w7938_
	);
	LUT2 #(
		.INIT('h4)
	) name6937 (
		_w7933_,
		_w7937_,
		_w7939_
	);
	LUT2 #(
		.INIT('h1)
	) name6938 (
		_w7902_,
		_w7905_,
		_w7940_
	);
	LUT2 #(
		.INIT('h2)
	) name6939 (
		_w7903_,
		_w7940_,
		_w7941_
	);
	LUT2 #(
		.INIT('h4)
	) name6940 (
		_w7903_,
		_w7940_,
		_w7942_
	);
	LUT2 #(
		.INIT('h1)
	) name6941 (
		_w7941_,
		_w7942_,
		_w7943_
	);
	LUT2 #(
		.INIT('h4)
	) name6942 (
		_w7939_,
		_w7943_,
		_w7944_
	);
	LUT2 #(
		.INIT('h1)
	) name6943 (
		_w7938_,
		_w7944_,
		_w7945_
	);
	LUT2 #(
		.INIT('h2)
	) name6944 (
		_w7926_,
		_w7945_,
		_w7946_
	);
	LUT2 #(
		.INIT('h4)
	) name6945 (
		_w7926_,
		_w7945_,
		_w7947_
	);
	LUT2 #(
		.INIT('h1)
	) name6946 (
		_w7946_,
		_w7947_,
		_w7948_
	);
	LUT2 #(
		.INIT('h8)
	) name6947 (
		_w7907_,
		_w7948_,
		_w7949_
	);
	LUT2 #(
		.INIT('h1)
	) name6948 (
		_w7907_,
		_w7948_,
		_w7950_
	);
	LUT2 #(
		.INIT('h1)
	) name6949 (
		_w7949_,
		_w7950_,
		_w7951_
	);
	LUT2 #(
		.INIT('h8)
	) name6950 (
		\A[574] ,
		\A[575] ,
		_w7952_
	);
	LUT2 #(
		.INIT('h8)
	) name6951 (
		\A[571] ,
		\A[572] ,
		_w7953_
	);
	LUT2 #(
		.INIT('h1)
	) name6952 (
		\A[571] ,
		\A[572] ,
		_w7954_
	);
	LUT2 #(
		.INIT('h1)
	) name6953 (
		_w7953_,
		_w7954_,
		_w7955_
	);
	LUT2 #(
		.INIT('h8)
	) name6954 (
		\A[573] ,
		_w7955_,
		_w7956_
	);
	LUT2 #(
		.INIT('h1)
	) name6955 (
		\A[573] ,
		_w7955_,
		_w7957_
	);
	LUT2 #(
		.INIT('h1)
	) name6956 (
		_w7956_,
		_w7957_,
		_w7958_
	);
	LUT2 #(
		.INIT('h1)
	) name6957 (
		\A[574] ,
		\A[575] ,
		_w7959_
	);
	LUT2 #(
		.INIT('h1)
	) name6958 (
		_w7952_,
		_w7959_,
		_w7960_
	);
	LUT2 #(
		.INIT('h8)
	) name6959 (
		\A[576] ,
		_w7960_,
		_w7961_
	);
	LUT2 #(
		.INIT('h1)
	) name6960 (
		\A[576] ,
		_w7960_,
		_w7962_
	);
	LUT2 #(
		.INIT('h1)
	) name6961 (
		_w7961_,
		_w7962_,
		_w7963_
	);
	LUT2 #(
		.INIT('h8)
	) name6962 (
		_w7958_,
		_w7963_,
		_w7964_
	);
	LUT2 #(
		.INIT('h8)
	) name6963 (
		_w7952_,
		_w7964_,
		_w7965_
	);
	LUT2 #(
		.INIT('h1)
	) name6964 (
		_w7953_,
		_w7956_,
		_w7966_
	);
	LUT2 #(
		.INIT('h1)
	) name6965 (
		_w7952_,
		_w7961_,
		_w7967_
	);
	LUT2 #(
		.INIT('h4)
	) name6966 (
		_w7964_,
		_w7967_,
		_w7968_
	);
	LUT2 #(
		.INIT('h1)
	) name6967 (
		_w7966_,
		_w7968_,
		_w7969_
	);
	LUT2 #(
		.INIT('h1)
	) name6968 (
		_w7965_,
		_w7969_,
		_w7970_
	);
	LUT2 #(
		.INIT('h8)
	) name6969 (
		\A[580] ,
		\A[581] ,
		_w7971_
	);
	LUT2 #(
		.INIT('h1)
	) name6970 (
		\A[580] ,
		\A[581] ,
		_w7972_
	);
	LUT2 #(
		.INIT('h1)
	) name6971 (
		_w7971_,
		_w7972_,
		_w7973_
	);
	LUT2 #(
		.INIT('h8)
	) name6972 (
		\A[582] ,
		_w7973_,
		_w7974_
	);
	LUT2 #(
		.INIT('h1)
	) name6973 (
		_w7971_,
		_w7974_,
		_w7975_
	);
	LUT2 #(
		.INIT('h8)
	) name6974 (
		\A[577] ,
		\A[578] ,
		_w7976_
	);
	LUT2 #(
		.INIT('h1)
	) name6975 (
		\A[577] ,
		\A[578] ,
		_w7977_
	);
	LUT2 #(
		.INIT('h1)
	) name6976 (
		_w7976_,
		_w7977_,
		_w7978_
	);
	LUT2 #(
		.INIT('h8)
	) name6977 (
		\A[579] ,
		_w7978_,
		_w7979_
	);
	LUT2 #(
		.INIT('h1)
	) name6978 (
		_w7976_,
		_w7979_,
		_w7980_
	);
	LUT2 #(
		.INIT('h8)
	) name6979 (
		_w7975_,
		_w7980_,
		_w7981_
	);
	LUT2 #(
		.INIT('h1)
	) name6980 (
		_w7975_,
		_w7980_,
		_w7982_
	);
	LUT2 #(
		.INIT('h1)
	) name6981 (
		\A[579] ,
		_w7978_,
		_w7983_
	);
	LUT2 #(
		.INIT('h1)
	) name6982 (
		_w7979_,
		_w7983_,
		_w7984_
	);
	LUT2 #(
		.INIT('h1)
	) name6983 (
		\A[582] ,
		_w7973_,
		_w7985_
	);
	LUT2 #(
		.INIT('h1)
	) name6984 (
		_w7974_,
		_w7985_,
		_w7986_
	);
	LUT2 #(
		.INIT('h8)
	) name6985 (
		_w7984_,
		_w7986_,
		_w7987_
	);
	LUT2 #(
		.INIT('h1)
	) name6986 (
		_w7982_,
		_w7987_,
		_w7988_
	);
	LUT2 #(
		.INIT('h1)
	) name6987 (
		_w7981_,
		_w7988_,
		_w7989_
	);
	LUT2 #(
		.INIT('h1)
	) name6988 (
		_w7984_,
		_w7986_,
		_w7990_
	);
	LUT2 #(
		.INIT('h1)
	) name6989 (
		_w7987_,
		_w7990_,
		_w7991_
	);
	LUT2 #(
		.INIT('h1)
	) name6990 (
		_w7958_,
		_w7963_,
		_w7992_
	);
	LUT2 #(
		.INIT('h1)
	) name6991 (
		_w7964_,
		_w7992_,
		_w7993_
	);
	LUT2 #(
		.INIT('h8)
	) name6992 (
		_w7991_,
		_w7993_,
		_w7994_
	);
	LUT2 #(
		.INIT('h2)
	) name6993 (
		_w7965_,
		_w7966_,
		_w7995_
	);
	LUT2 #(
		.INIT('h2)
	) name6994 (
		_w7994_,
		_w7995_,
		_w7996_
	);
	LUT2 #(
		.INIT('h1)
	) name6995 (
		_w7981_,
		_w7982_,
		_w7997_
	);
	LUT2 #(
		.INIT('h2)
	) name6996 (
		_w7987_,
		_w7997_,
		_w7998_
	);
	LUT2 #(
		.INIT('h4)
	) name6997 (
		_w7987_,
		_w7997_,
		_w7999_
	);
	LUT2 #(
		.INIT('h1)
	) name6998 (
		_w7998_,
		_w7999_,
		_w8000_
	);
	LUT2 #(
		.INIT('h2)
	) name6999 (
		_w7996_,
		_w8000_,
		_w8001_
	);
	LUT2 #(
		.INIT('h4)
	) name7000 (
		_w7996_,
		_w8000_,
		_w8002_
	);
	LUT2 #(
		.INIT('h1)
	) name7001 (
		_w7965_,
		_w7968_,
		_w8003_
	);
	LUT2 #(
		.INIT('h2)
	) name7002 (
		_w7966_,
		_w8003_,
		_w8004_
	);
	LUT2 #(
		.INIT('h4)
	) name7003 (
		_w7966_,
		_w8003_,
		_w8005_
	);
	LUT2 #(
		.INIT('h1)
	) name7004 (
		_w8004_,
		_w8005_,
		_w8006_
	);
	LUT2 #(
		.INIT('h4)
	) name7005 (
		_w8002_,
		_w8006_,
		_w8007_
	);
	LUT2 #(
		.INIT('h1)
	) name7006 (
		_w8001_,
		_w8007_,
		_w8008_
	);
	LUT2 #(
		.INIT('h2)
	) name7007 (
		_w7989_,
		_w8008_,
		_w8009_
	);
	LUT2 #(
		.INIT('h4)
	) name7008 (
		_w7989_,
		_w8008_,
		_w8010_
	);
	LUT2 #(
		.INIT('h1)
	) name7009 (
		_w8009_,
		_w8010_,
		_w8011_
	);
	LUT2 #(
		.INIT('h8)
	) name7010 (
		_w7970_,
		_w8011_,
		_w8012_
	);
	LUT2 #(
		.INIT('h1)
	) name7011 (
		_w7970_,
		_w8011_,
		_w8013_
	);
	LUT2 #(
		.INIT('h1)
	) name7012 (
		_w8012_,
		_w8013_,
		_w8014_
	);
	LUT2 #(
		.INIT('h1)
	) name7013 (
		_w7951_,
		_w8014_,
		_w8015_
	);
	LUT2 #(
		.INIT('h8)
	) name7014 (
		_w7951_,
		_w8014_,
		_w8016_
	);
	LUT2 #(
		.INIT('h1)
	) name7015 (
		_w7991_,
		_w7993_,
		_w8017_
	);
	LUT2 #(
		.INIT('h1)
	) name7016 (
		_w7994_,
		_w8017_,
		_w8018_
	);
	LUT2 #(
		.INIT('h1)
	) name7017 (
		_w7928_,
		_w7930_,
		_w8019_
	);
	LUT2 #(
		.INIT('h1)
	) name7018 (
		_w7931_,
		_w8019_,
		_w8020_
	);
	LUT2 #(
		.INIT('h8)
	) name7019 (
		_w8018_,
		_w8020_,
		_w8021_
	);
	LUT2 #(
		.INIT('h1)
	) name7020 (
		_w8001_,
		_w8002_,
		_w8022_
	);
	LUT2 #(
		.INIT('h8)
	) name7021 (
		_w8006_,
		_w8022_,
		_w8023_
	);
	LUT2 #(
		.INIT('h1)
	) name7022 (
		_w8006_,
		_w8022_,
		_w8024_
	);
	LUT2 #(
		.INIT('h1)
	) name7023 (
		_w8023_,
		_w8024_,
		_w8025_
	);
	LUT2 #(
		.INIT('h8)
	) name7024 (
		_w8021_,
		_w8025_,
		_w8026_
	);
	LUT2 #(
		.INIT('h1)
	) name7025 (
		_w8021_,
		_w8025_,
		_w8027_
	);
	LUT2 #(
		.INIT('h1)
	) name7026 (
		_w7938_,
		_w7939_,
		_w8028_
	);
	LUT2 #(
		.INIT('h8)
	) name7027 (
		_w7943_,
		_w8028_,
		_w8029_
	);
	LUT2 #(
		.INIT('h1)
	) name7028 (
		_w7943_,
		_w8028_,
		_w8030_
	);
	LUT2 #(
		.INIT('h1)
	) name7029 (
		_w8029_,
		_w8030_,
		_w8031_
	);
	LUT2 #(
		.INIT('h4)
	) name7030 (
		_w8027_,
		_w8031_,
		_w8032_
	);
	LUT2 #(
		.INIT('h1)
	) name7031 (
		_w8026_,
		_w8032_,
		_w8033_
	);
	LUT2 #(
		.INIT('h1)
	) name7032 (
		_w8016_,
		_w8033_,
		_w8034_
	);
	LUT2 #(
		.INIT('h1)
	) name7033 (
		_w8015_,
		_w8034_,
		_w8035_
	);
	LUT2 #(
		.INIT('h1)
	) name7034 (
		_w7970_,
		_w8010_,
		_w8036_
	);
	LUT2 #(
		.INIT('h1)
	) name7035 (
		_w8009_,
		_w8036_,
		_w8037_
	);
	LUT2 #(
		.INIT('h1)
	) name7036 (
		_w8035_,
		_w8037_,
		_w8038_
	);
	LUT2 #(
		.INIT('h8)
	) name7037 (
		_w8035_,
		_w8037_,
		_w8039_
	);
	LUT2 #(
		.INIT('h1)
	) name7038 (
		_w7907_,
		_w7947_,
		_w8040_
	);
	LUT2 #(
		.INIT('h1)
	) name7039 (
		_w7946_,
		_w8040_,
		_w8041_
	);
	LUT2 #(
		.INIT('h1)
	) name7040 (
		_w8039_,
		_w8041_,
		_w8042_
	);
	LUT2 #(
		.INIT('h1)
	) name7041 (
		_w8038_,
		_w8042_,
		_w8043_
	);
	LUT2 #(
		.INIT('h8)
	) name7042 (
		\A[586] ,
		\A[587] ,
		_w8044_
	);
	LUT2 #(
		.INIT('h8)
	) name7043 (
		\A[583] ,
		\A[584] ,
		_w8045_
	);
	LUT2 #(
		.INIT('h1)
	) name7044 (
		\A[583] ,
		\A[584] ,
		_w8046_
	);
	LUT2 #(
		.INIT('h1)
	) name7045 (
		_w8045_,
		_w8046_,
		_w8047_
	);
	LUT2 #(
		.INIT('h8)
	) name7046 (
		\A[585] ,
		_w8047_,
		_w8048_
	);
	LUT2 #(
		.INIT('h1)
	) name7047 (
		\A[585] ,
		_w8047_,
		_w8049_
	);
	LUT2 #(
		.INIT('h1)
	) name7048 (
		_w8048_,
		_w8049_,
		_w8050_
	);
	LUT2 #(
		.INIT('h1)
	) name7049 (
		\A[586] ,
		\A[587] ,
		_w8051_
	);
	LUT2 #(
		.INIT('h1)
	) name7050 (
		_w8044_,
		_w8051_,
		_w8052_
	);
	LUT2 #(
		.INIT('h8)
	) name7051 (
		\A[588] ,
		_w8052_,
		_w8053_
	);
	LUT2 #(
		.INIT('h1)
	) name7052 (
		\A[588] ,
		_w8052_,
		_w8054_
	);
	LUT2 #(
		.INIT('h1)
	) name7053 (
		_w8053_,
		_w8054_,
		_w8055_
	);
	LUT2 #(
		.INIT('h8)
	) name7054 (
		_w8050_,
		_w8055_,
		_w8056_
	);
	LUT2 #(
		.INIT('h8)
	) name7055 (
		_w8044_,
		_w8056_,
		_w8057_
	);
	LUT2 #(
		.INIT('h1)
	) name7056 (
		_w8045_,
		_w8048_,
		_w8058_
	);
	LUT2 #(
		.INIT('h1)
	) name7057 (
		_w8044_,
		_w8053_,
		_w8059_
	);
	LUT2 #(
		.INIT('h4)
	) name7058 (
		_w8056_,
		_w8059_,
		_w8060_
	);
	LUT2 #(
		.INIT('h1)
	) name7059 (
		_w8058_,
		_w8060_,
		_w8061_
	);
	LUT2 #(
		.INIT('h1)
	) name7060 (
		_w8057_,
		_w8061_,
		_w8062_
	);
	LUT2 #(
		.INIT('h8)
	) name7061 (
		\A[592] ,
		\A[593] ,
		_w8063_
	);
	LUT2 #(
		.INIT('h1)
	) name7062 (
		\A[592] ,
		\A[593] ,
		_w8064_
	);
	LUT2 #(
		.INIT('h1)
	) name7063 (
		_w8063_,
		_w8064_,
		_w8065_
	);
	LUT2 #(
		.INIT('h8)
	) name7064 (
		\A[594] ,
		_w8065_,
		_w8066_
	);
	LUT2 #(
		.INIT('h1)
	) name7065 (
		_w8063_,
		_w8066_,
		_w8067_
	);
	LUT2 #(
		.INIT('h8)
	) name7066 (
		\A[589] ,
		\A[590] ,
		_w8068_
	);
	LUT2 #(
		.INIT('h1)
	) name7067 (
		\A[589] ,
		\A[590] ,
		_w8069_
	);
	LUT2 #(
		.INIT('h1)
	) name7068 (
		_w8068_,
		_w8069_,
		_w8070_
	);
	LUT2 #(
		.INIT('h8)
	) name7069 (
		\A[591] ,
		_w8070_,
		_w8071_
	);
	LUT2 #(
		.INIT('h1)
	) name7070 (
		_w8068_,
		_w8071_,
		_w8072_
	);
	LUT2 #(
		.INIT('h8)
	) name7071 (
		_w8067_,
		_w8072_,
		_w8073_
	);
	LUT2 #(
		.INIT('h1)
	) name7072 (
		_w8067_,
		_w8072_,
		_w8074_
	);
	LUT2 #(
		.INIT('h1)
	) name7073 (
		\A[591] ,
		_w8070_,
		_w8075_
	);
	LUT2 #(
		.INIT('h1)
	) name7074 (
		_w8071_,
		_w8075_,
		_w8076_
	);
	LUT2 #(
		.INIT('h1)
	) name7075 (
		\A[594] ,
		_w8065_,
		_w8077_
	);
	LUT2 #(
		.INIT('h1)
	) name7076 (
		_w8066_,
		_w8077_,
		_w8078_
	);
	LUT2 #(
		.INIT('h8)
	) name7077 (
		_w8076_,
		_w8078_,
		_w8079_
	);
	LUT2 #(
		.INIT('h1)
	) name7078 (
		_w8074_,
		_w8079_,
		_w8080_
	);
	LUT2 #(
		.INIT('h1)
	) name7079 (
		_w8073_,
		_w8080_,
		_w8081_
	);
	LUT2 #(
		.INIT('h1)
	) name7080 (
		_w8076_,
		_w8078_,
		_w8082_
	);
	LUT2 #(
		.INIT('h1)
	) name7081 (
		_w8079_,
		_w8082_,
		_w8083_
	);
	LUT2 #(
		.INIT('h1)
	) name7082 (
		_w8050_,
		_w8055_,
		_w8084_
	);
	LUT2 #(
		.INIT('h1)
	) name7083 (
		_w8056_,
		_w8084_,
		_w8085_
	);
	LUT2 #(
		.INIT('h8)
	) name7084 (
		_w8083_,
		_w8085_,
		_w8086_
	);
	LUT2 #(
		.INIT('h2)
	) name7085 (
		_w8057_,
		_w8058_,
		_w8087_
	);
	LUT2 #(
		.INIT('h2)
	) name7086 (
		_w8086_,
		_w8087_,
		_w8088_
	);
	LUT2 #(
		.INIT('h1)
	) name7087 (
		_w8073_,
		_w8074_,
		_w8089_
	);
	LUT2 #(
		.INIT('h2)
	) name7088 (
		_w8079_,
		_w8089_,
		_w8090_
	);
	LUT2 #(
		.INIT('h4)
	) name7089 (
		_w8079_,
		_w8089_,
		_w8091_
	);
	LUT2 #(
		.INIT('h1)
	) name7090 (
		_w8090_,
		_w8091_,
		_w8092_
	);
	LUT2 #(
		.INIT('h2)
	) name7091 (
		_w8088_,
		_w8092_,
		_w8093_
	);
	LUT2 #(
		.INIT('h4)
	) name7092 (
		_w8088_,
		_w8092_,
		_w8094_
	);
	LUT2 #(
		.INIT('h1)
	) name7093 (
		_w8057_,
		_w8060_,
		_w8095_
	);
	LUT2 #(
		.INIT('h2)
	) name7094 (
		_w8058_,
		_w8095_,
		_w8096_
	);
	LUT2 #(
		.INIT('h4)
	) name7095 (
		_w8058_,
		_w8095_,
		_w8097_
	);
	LUT2 #(
		.INIT('h1)
	) name7096 (
		_w8096_,
		_w8097_,
		_w8098_
	);
	LUT2 #(
		.INIT('h4)
	) name7097 (
		_w8094_,
		_w8098_,
		_w8099_
	);
	LUT2 #(
		.INIT('h1)
	) name7098 (
		_w8093_,
		_w8099_,
		_w8100_
	);
	LUT2 #(
		.INIT('h2)
	) name7099 (
		_w8081_,
		_w8100_,
		_w8101_
	);
	LUT2 #(
		.INIT('h4)
	) name7100 (
		_w8081_,
		_w8100_,
		_w8102_
	);
	LUT2 #(
		.INIT('h1)
	) name7101 (
		_w8101_,
		_w8102_,
		_w8103_
	);
	LUT2 #(
		.INIT('h8)
	) name7102 (
		_w8062_,
		_w8103_,
		_w8104_
	);
	LUT2 #(
		.INIT('h1)
	) name7103 (
		_w8062_,
		_w8103_,
		_w8105_
	);
	LUT2 #(
		.INIT('h1)
	) name7104 (
		_w8104_,
		_w8105_,
		_w8106_
	);
	LUT2 #(
		.INIT('h8)
	) name7105 (
		\A[598] ,
		\A[599] ,
		_w8107_
	);
	LUT2 #(
		.INIT('h8)
	) name7106 (
		\A[595] ,
		\A[596] ,
		_w8108_
	);
	LUT2 #(
		.INIT('h1)
	) name7107 (
		\A[595] ,
		\A[596] ,
		_w8109_
	);
	LUT2 #(
		.INIT('h1)
	) name7108 (
		_w8108_,
		_w8109_,
		_w8110_
	);
	LUT2 #(
		.INIT('h8)
	) name7109 (
		\A[597] ,
		_w8110_,
		_w8111_
	);
	LUT2 #(
		.INIT('h1)
	) name7110 (
		\A[597] ,
		_w8110_,
		_w8112_
	);
	LUT2 #(
		.INIT('h1)
	) name7111 (
		_w8111_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h1)
	) name7112 (
		\A[598] ,
		\A[599] ,
		_w8114_
	);
	LUT2 #(
		.INIT('h1)
	) name7113 (
		_w8107_,
		_w8114_,
		_w8115_
	);
	LUT2 #(
		.INIT('h8)
	) name7114 (
		\A[600] ,
		_w8115_,
		_w8116_
	);
	LUT2 #(
		.INIT('h1)
	) name7115 (
		\A[600] ,
		_w8115_,
		_w8117_
	);
	LUT2 #(
		.INIT('h1)
	) name7116 (
		_w8116_,
		_w8117_,
		_w8118_
	);
	LUT2 #(
		.INIT('h8)
	) name7117 (
		_w8113_,
		_w8118_,
		_w8119_
	);
	LUT2 #(
		.INIT('h8)
	) name7118 (
		_w8107_,
		_w8119_,
		_w8120_
	);
	LUT2 #(
		.INIT('h1)
	) name7119 (
		_w8108_,
		_w8111_,
		_w8121_
	);
	LUT2 #(
		.INIT('h1)
	) name7120 (
		_w8107_,
		_w8116_,
		_w8122_
	);
	LUT2 #(
		.INIT('h4)
	) name7121 (
		_w8119_,
		_w8122_,
		_w8123_
	);
	LUT2 #(
		.INIT('h1)
	) name7122 (
		_w8121_,
		_w8123_,
		_w8124_
	);
	LUT2 #(
		.INIT('h1)
	) name7123 (
		_w8120_,
		_w8124_,
		_w8125_
	);
	LUT2 #(
		.INIT('h8)
	) name7124 (
		\A[604] ,
		\A[605] ,
		_w8126_
	);
	LUT2 #(
		.INIT('h1)
	) name7125 (
		\A[604] ,
		\A[605] ,
		_w8127_
	);
	LUT2 #(
		.INIT('h1)
	) name7126 (
		_w8126_,
		_w8127_,
		_w8128_
	);
	LUT2 #(
		.INIT('h8)
	) name7127 (
		\A[606] ,
		_w8128_,
		_w8129_
	);
	LUT2 #(
		.INIT('h1)
	) name7128 (
		_w8126_,
		_w8129_,
		_w8130_
	);
	LUT2 #(
		.INIT('h8)
	) name7129 (
		\A[601] ,
		\A[602] ,
		_w8131_
	);
	LUT2 #(
		.INIT('h1)
	) name7130 (
		\A[601] ,
		\A[602] ,
		_w8132_
	);
	LUT2 #(
		.INIT('h1)
	) name7131 (
		_w8131_,
		_w8132_,
		_w8133_
	);
	LUT2 #(
		.INIT('h8)
	) name7132 (
		\A[603] ,
		_w8133_,
		_w8134_
	);
	LUT2 #(
		.INIT('h1)
	) name7133 (
		_w8131_,
		_w8134_,
		_w8135_
	);
	LUT2 #(
		.INIT('h8)
	) name7134 (
		_w8130_,
		_w8135_,
		_w8136_
	);
	LUT2 #(
		.INIT('h1)
	) name7135 (
		_w8130_,
		_w8135_,
		_w8137_
	);
	LUT2 #(
		.INIT('h1)
	) name7136 (
		\A[603] ,
		_w8133_,
		_w8138_
	);
	LUT2 #(
		.INIT('h1)
	) name7137 (
		_w8134_,
		_w8138_,
		_w8139_
	);
	LUT2 #(
		.INIT('h1)
	) name7138 (
		\A[606] ,
		_w8128_,
		_w8140_
	);
	LUT2 #(
		.INIT('h1)
	) name7139 (
		_w8129_,
		_w8140_,
		_w8141_
	);
	LUT2 #(
		.INIT('h8)
	) name7140 (
		_w8139_,
		_w8141_,
		_w8142_
	);
	LUT2 #(
		.INIT('h1)
	) name7141 (
		_w8137_,
		_w8142_,
		_w8143_
	);
	LUT2 #(
		.INIT('h1)
	) name7142 (
		_w8136_,
		_w8143_,
		_w8144_
	);
	LUT2 #(
		.INIT('h1)
	) name7143 (
		_w8139_,
		_w8141_,
		_w8145_
	);
	LUT2 #(
		.INIT('h1)
	) name7144 (
		_w8142_,
		_w8145_,
		_w8146_
	);
	LUT2 #(
		.INIT('h1)
	) name7145 (
		_w8113_,
		_w8118_,
		_w8147_
	);
	LUT2 #(
		.INIT('h1)
	) name7146 (
		_w8119_,
		_w8147_,
		_w8148_
	);
	LUT2 #(
		.INIT('h8)
	) name7147 (
		_w8146_,
		_w8148_,
		_w8149_
	);
	LUT2 #(
		.INIT('h2)
	) name7148 (
		_w8120_,
		_w8121_,
		_w8150_
	);
	LUT2 #(
		.INIT('h2)
	) name7149 (
		_w8149_,
		_w8150_,
		_w8151_
	);
	LUT2 #(
		.INIT('h1)
	) name7150 (
		_w8136_,
		_w8137_,
		_w8152_
	);
	LUT2 #(
		.INIT('h2)
	) name7151 (
		_w8142_,
		_w8152_,
		_w8153_
	);
	LUT2 #(
		.INIT('h4)
	) name7152 (
		_w8142_,
		_w8152_,
		_w8154_
	);
	LUT2 #(
		.INIT('h1)
	) name7153 (
		_w8153_,
		_w8154_,
		_w8155_
	);
	LUT2 #(
		.INIT('h2)
	) name7154 (
		_w8151_,
		_w8155_,
		_w8156_
	);
	LUT2 #(
		.INIT('h4)
	) name7155 (
		_w8151_,
		_w8155_,
		_w8157_
	);
	LUT2 #(
		.INIT('h1)
	) name7156 (
		_w8120_,
		_w8123_,
		_w8158_
	);
	LUT2 #(
		.INIT('h2)
	) name7157 (
		_w8121_,
		_w8158_,
		_w8159_
	);
	LUT2 #(
		.INIT('h4)
	) name7158 (
		_w8121_,
		_w8158_,
		_w8160_
	);
	LUT2 #(
		.INIT('h1)
	) name7159 (
		_w8159_,
		_w8160_,
		_w8161_
	);
	LUT2 #(
		.INIT('h4)
	) name7160 (
		_w8157_,
		_w8161_,
		_w8162_
	);
	LUT2 #(
		.INIT('h1)
	) name7161 (
		_w8156_,
		_w8162_,
		_w8163_
	);
	LUT2 #(
		.INIT('h2)
	) name7162 (
		_w8144_,
		_w8163_,
		_w8164_
	);
	LUT2 #(
		.INIT('h4)
	) name7163 (
		_w8144_,
		_w8163_,
		_w8165_
	);
	LUT2 #(
		.INIT('h1)
	) name7164 (
		_w8164_,
		_w8165_,
		_w8166_
	);
	LUT2 #(
		.INIT('h8)
	) name7165 (
		_w8125_,
		_w8166_,
		_w8167_
	);
	LUT2 #(
		.INIT('h1)
	) name7166 (
		_w8125_,
		_w8166_,
		_w8168_
	);
	LUT2 #(
		.INIT('h1)
	) name7167 (
		_w8167_,
		_w8168_,
		_w8169_
	);
	LUT2 #(
		.INIT('h1)
	) name7168 (
		_w8106_,
		_w8169_,
		_w8170_
	);
	LUT2 #(
		.INIT('h8)
	) name7169 (
		_w8106_,
		_w8169_,
		_w8171_
	);
	LUT2 #(
		.INIT('h1)
	) name7170 (
		_w8146_,
		_w8148_,
		_w8172_
	);
	LUT2 #(
		.INIT('h1)
	) name7171 (
		_w8149_,
		_w8172_,
		_w8173_
	);
	LUT2 #(
		.INIT('h1)
	) name7172 (
		_w8083_,
		_w8085_,
		_w8174_
	);
	LUT2 #(
		.INIT('h1)
	) name7173 (
		_w8086_,
		_w8174_,
		_w8175_
	);
	LUT2 #(
		.INIT('h8)
	) name7174 (
		_w8173_,
		_w8175_,
		_w8176_
	);
	LUT2 #(
		.INIT('h1)
	) name7175 (
		_w8156_,
		_w8157_,
		_w8177_
	);
	LUT2 #(
		.INIT('h8)
	) name7176 (
		_w8161_,
		_w8177_,
		_w8178_
	);
	LUT2 #(
		.INIT('h1)
	) name7177 (
		_w8161_,
		_w8177_,
		_w8179_
	);
	LUT2 #(
		.INIT('h1)
	) name7178 (
		_w8178_,
		_w8179_,
		_w8180_
	);
	LUT2 #(
		.INIT('h8)
	) name7179 (
		_w8176_,
		_w8180_,
		_w8181_
	);
	LUT2 #(
		.INIT('h1)
	) name7180 (
		_w8176_,
		_w8180_,
		_w8182_
	);
	LUT2 #(
		.INIT('h1)
	) name7181 (
		_w8093_,
		_w8094_,
		_w8183_
	);
	LUT2 #(
		.INIT('h8)
	) name7182 (
		_w8098_,
		_w8183_,
		_w8184_
	);
	LUT2 #(
		.INIT('h1)
	) name7183 (
		_w8098_,
		_w8183_,
		_w8185_
	);
	LUT2 #(
		.INIT('h1)
	) name7184 (
		_w8184_,
		_w8185_,
		_w8186_
	);
	LUT2 #(
		.INIT('h4)
	) name7185 (
		_w8182_,
		_w8186_,
		_w8187_
	);
	LUT2 #(
		.INIT('h1)
	) name7186 (
		_w8181_,
		_w8187_,
		_w8188_
	);
	LUT2 #(
		.INIT('h1)
	) name7187 (
		_w8171_,
		_w8188_,
		_w8189_
	);
	LUT2 #(
		.INIT('h1)
	) name7188 (
		_w8170_,
		_w8189_,
		_w8190_
	);
	LUT2 #(
		.INIT('h1)
	) name7189 (
		_w8125_,
		_w8165_,
		_w8191_
	);
	LUT2 #(
		.INIT('h1)
	) name7190 (
		_w8164_,
		_w8191_,
		_w8192_
	);
	LUT2 #(
		.INIT('h1)
	) name7191 (
		_w8190_,
		_w8192_,
		_w8193_
	);
	LUT2 #(
		.INIT('h8)
	) name7192 (
		_w8190_,
		_w8192_,
		_w8194_
	);
	LUT2 #(
		.INIT('h1)
	) name7193 (
		_w8193_,
		_w8194_,
		_w8195_
	);
	LUT2 #(
		.INIT('h1)
	) name7194 (
		_w8062_,
		_w8102_,
		_w8196_
	);
	LUT2 #(
		.INIT('h1)
	) name7195 (
		_w8101_,
		_w8196_,
		_w8197_
	);
	LUT2 #(
		.INIT('h2)
	) name7196 (
		_w8195_,
		_w8197_,
		_w8198_
	);
	LUT2 #(
		.INIT('h4)
	) name7197 (
		_w8195_,
		_w8197_,
		_w8199_
	);
	LUT2 #(
		.INIT('h1)
	) name7198 (
		_w8198_,
		_w8199_,
		_w8200_
	);
	LUT2 #(
		.INIT('h1)
	) name7199 (
		_w8038_,
		_w8039_,
		_w8201_
	);
	LUT2 #(
		.INIT('h4)
	) name7200 (
		_w8041_,
		_w8201_,
		_w8202_
	);
	LUT2 #(
		.INIT('h2)
	) name7201 (
		_w8041_,
		_w8201_,
		_w8203_
	);
	LUT2 #(
		.INIT('h1)
	) name7202 (
		_w8202_,
		_w8203_,
		_w8204_
	);
	LUT2 #(
		.INIT('h1)
	) name7203 (
		_w8200_,
		_w8204_,
		_w8205_
	);
	LUT2 #(
		.INIT('h8)
	) name7204 (
		_w8200_,
		_w8204_,
		_w8206_
	);
	LUT2 #(
		.INIT('h1)
	) name7205 (
		_w8015_,
		_w8016_,
		_w8207_
	);
	LUT2 #(
		.INIT('h4)
	) name7206 (
		_w8033_,
		_w8207_,
		_w8208_
	);
	LUT2 #(
		.INIT('h2)
	) name7207 (
		_w8033_,
		_w8207_,
		_w8209_
	);
	LUT2 #(
		.INIT('h1)
	) name7208 (
		_w8208_,
		_w8209_,
		_w8210_
	);
	LUT2 #(
		.INIT('h1)
	) name7209 (
		_w8170_,
		_w8171_,
		_w8211_
	);
	LUT2 #(
		.INIT('h4)
	) name7210 (
		_w8188_,
		_w8211_,
		_w8212_
	);
	LUT2 #(
		.INIT('h2)
	) name7211 (
		_w8188_,
		_w8211_,
		_w8213_
	);
	LUT2 #(
		.INIT('h1)
	) name7212 (
		_w8212_,
		_w8213_,
		_w8214_
	);
	LUT2 #(
		.INIT('h1)
	) name7213 (
		_w8210_,
		_w8214_,
		_w8215_
	);
	LUT2 #(
		.INIT('h8)
	) name7214 (
		_w8210_,
		_w8214_,
		_w8216_
	);
	LUT2 #(
		.INIT('h1)
	) name7215 (
		_w8173_,
		_w8175_,
		_w8217_
	);
	LUT2 #(
		.INIT('h1)
	) name7216 (
		_w8176_,
		_w8217_,
		_w8218_
	);
	LUT2 #(
		.INIT('h1)
	) name7217 (
		_w8018_,
		_w8020_,
		_w8219_
	);
	LUT2 #(
		.INIT('h1)
	) name7218 (
		_w8021_,
		_w8219_,
		_w8220_
	);
	LUT2 #(
		.INIT('h8)
	) name7219 (
		_w8218_,
		_w8220_,
		_w8221_
	);
	LUT2 #(
		.INIT('h1)
	) name7220 (
		_w8181_,
		_w8182_,
		_w8222_
	);
	LUT2 #(
		.INIT('h4)
	) name7221 (
		_w8186_,
		_w8222_,
		_w8223_
	);
	LUT2 #(
		.INIT('h2)
	) name7222 (
		_w8186_,
		_w8222_,
		_w8224_
	);
	LUT2 #(
		.INIT('h1)
	) name7223 (
		_w8223_,
		_w8224_,
		_w8225_
	);
	LUT2 #(
		.INIT('h2)
	) name7224 (
		_w8221_,
		_w8225_,
		_w8226_
	);
	LUT2 #(
		.INIT('h4)
	) name7225 (
		_w8221_,
		_w8225_,
		_w8227_
	);
	LUT2 #(
		.INIT('h1)
	) name7226 (
		_w8026_,
		_w8027_,
		_w8228_
	);
	LUT2 #(
		.INIT('h4)
	) name7227 (
		_w8031_,
		_w8228_,
		_w8229_
	);
	LUT2 #(
		.INIT('h2)
	) name7228 (
		_w8031_,
		_w8228_,
		_w8230_
	);
	LUT2 #(
		.INIT('h1)
	) name7229 (
		_w8229_,
		_w8230_,
		_w8231_
	);
	LUT2 #(
		.INIT('h1)
	) name7230 (
		_w8227_,
		_w8231_,
		_w8232_
	);
	LUT2 #(
		.INIT('h1)
	) name7231 (
		_w8226_,
		_w8232_,
		_w8233_
	);
	LUT2 #(
		.INIT('h4)
	) name7232 (
		_w8216_,
		_w8233_,
		_w8234_
	);
	LUT2 #(
		.INIT('h1)
	) name7233 (
		_w8215_,
		_w8234_,
		_w8235_
	);
	LUT2 #(
		.INIT('h1)
	) name7234 (
		_w8206_,
		_w8235_,
		_w8236_
	);
	LUT2 #(
		.INIT('h1)
	) name7235 (
		_w8205_,
		_w8236_,
		_w8237_
	);
	LUT2 #(
		.INIT('h2)
	) name7236 (
		_w8043_,
		_w8237_,
		_w8238_
	);
	LUT2 #(
		.INIT('h4)
	) name7237 (
		_w8043_,
		_w8237_,
		_w8239_
	);
	LUT2 #(
		.INIT('h1)
	) name7238 (
		_w8238_,
		_w8239_,
		_w8240_
	);
	LUT2 #(
		.INIT('h1)
	) name7239 (
		_w8194_,
		_w8197_,
		_w8241_
	);
	LUT2 #(
		.INIT('h1)
	) name7240 (
		_w8193_,
		_w8241_,
		_w8242_
	);
	LUT2 #(
		.INIT('h8)
	) name7241 (
		_w8240_,
		_w8242_,
		_w8243_
	);
	LUT2 #(
		.INIT('h1)
	) name7242 (
		_w8240_,
		_w8242_,
		_w8244_
	);
	LUT2 #(
		.INIT('h1)
	) name7243 (
		_w8243_,
		_w8244_,
		_w8245_
	);
	LUT2 #(
		.INIT('h8)
	) name7244 (
		\A[634] ,
		\A[635] ,
		_w8246_
	);
	LUT2 #(
		.INIT('h8)
	) name7245 (
		\A[631] ,
		\A[632] ,
		_w8247_
	);
	LUT2 #(
		.INIT('h1)
	) name7246 (
		\A[631] ,
		\A[632] ,
		_w8248_
	);
	LUT2 #(
		.INIT('h1)
	) name7247 (
		_w8247_,
		_w8248_,
		_w8249_
	);
	LUT2 #(
		.INIT('h8)
	) name7248 (
		\A[633] ,
		_w8249_,
		_w8250_
	);
	LUT2 #(
		.INIT('h1)
	) name7249 (
		\A[633] ,
		_w8249_,
		_w8251_
	);
	LUT2 #(
		.INIT('h1)
	) name7250 (
		_w8250_,
		_w8251_,
		_w8252_
	);
	LUT2 #(
		.INIT('h1)
	) name7251 (
		\A[634] ,
		\A[635] ,
		_w8253_
	);
	LUT2 #(
		.INIT('h1)
	) name7252 (
		_w8246_,
		_w8253_,
		_w8254_
	);
	LUT2 #(
		.INIT('h8)
	) name7253 (
		\A[636] ,
		_w8254_,
		_w8255_
	);
	LUT2 #(
		.INIT('h1)
	) name7254 (
		\A[636] ,
		_w8254_,
		_w8256_
	);
	LUT2 #(
		.INIT('h1)
	) name7255 (
		_w8255_,
		_w8256_,
		_w8257_
	);
	LUT2 #(
		.INIT('h8)
	) name7256 (
		_w8252_,
		_w8257_,
		_w8258_
	);
	LUT2 #(
		.INIT('h8)
	) name7257 (
		_w8246_,
		_w8258_,
		_w8259_
	);
	LUT2 #(
		.INIT('h1)
	) name7258 (
		_w8247_,
		_w8250_,
		_w8260_
	);
	LUT2 #(
		.INIT('h1)
	) name7259 (
		_w8246_,
		_w8255_,
		_w8261_
	);
	LUT2 #(
		.INIT('h4)
	) name7260 (
		_w8258_,
		_w8261_,
		_w8262_
	);
	LUT2 #(
		.INIT('h1)
	) name7261 (
		_w8260_,
		_w8262_,
		_w8263_
	);
	LUT2 #(
		.INIT('h1)
	) name7262 (
		_w8259_,
		_w8263_,
		_w8264_
	);
	LUT2 #(
		.INIT('h8)
	) name7263 (
		\A[640] ,
		\A[641] ,
		_w8265_
	);
	LUT2 #(
		.INIT('h1)
	) name7264 (
		\A[640] ,
		\A[641] ,
		_w8266_
	);
	LUT2 #(
		.INIT('h1)
	) name7265 (
		_w8265_,
		_w8266_,
		_w8267_
	);
	LUT2 #(
		.INIT('h8)
	) name7266 (
		\A[642] ,
		_w8267_,
		_w8268_
	);
	LUT2 #(
		.INIT('h1)
	) name7267 (
		_w8265_,
		_w8268_,
		_w8269_
	);
	LUT2 #(
		.INIT('h8)
	) name7268 (
		\A[637] ,
		\A[638] ,
		_w8270_
	);
	LUT2 #(
		.INIT('h1)
	) name7269 (
		\A[637] ,
		\A[638] ,
		_w8271_
	);
	LUT2 #(
		.INIT('h1)
	) name7270 (
		_w8270_,
		_w8271_,
		_w8272_
	);
	LUT2 #(
		.INIT('h8)
	) name7271 (
		\A[639] ,
		_w8272_,
		_w8273_
	);
	LUT2 #(
		.INIT('h1)
	) name7272 (
		_w8270_,
		_w8273_,
		_w8274_
	);
	LUT2 #(
		.INIT('h8)
	) name7273 (
		_w8269_,
		_w8274_,
		_w8275_
	);
	LUT2 #(
		.INIT('h1)
	) name7274 (
		_w8269_,
		_w8274_,
		_w8276_
	);
	LUT2 #(
		.INIT('h1)
	) name7275 (
		\A[639] ,
		_w8272_,
		_w8277_
	);
	LUT2 #(
		.INIT('h1)
	) name7276 (
		_w8273_,
		_w8277_,
		_w8278_
	);
	LUT2 #(
		.INIT('h1)
	) name7277 (
		\A[642] ,
		_w8267_,
		_w8279_
	);
	LUT2 #(
		.INIT('h1)
	) name7278 (
		_w8268_,
		_w8279_,
		_w8280_
	);
	LUT2 #(
		.INIT('h8)
	) name7279 (
		_w8278_,
		_w8280_,
		_w8281_
	);
	LUT2 #(
		.INIT('h1)
	) name7280 (
		_w8276_,
		_w8281_,
		_w8282_
	);
	LUT2 #(
		.INIT('h1)
	) name7281 (
		_w8275_,
		_w8282_,
		_w8283_
	);
	LUT2 #(
		.INIT('h1)
	) name7282 (
		_w8278_,
		_w8280_,
		_w8284_
	);
	LUT2 #(
		.INIT('h1)
	) name7283 (
		_w8281_,
		_w8284_,
		_w8285_
	);
	LUT2 #(
		.INIT('h1)
	) name7284 (
		_w8252_,
		_w8257_,
		_w8286_
	);
	LUT2 #(
		.INIT('h1)
	) name7285 (
		_w8258_,
		_w8286_,
		_w8287_
	);
	LUT2 #(
		.INIT('h8)
	) name7286 (
		_w8285_,
		_w8287_,
		_w8288_
	);
	LUT2 #(
		.INIT('h2)
	) name7287 (
		_w8259_,
		_w8260_,
		_w8289_
	);
	LUT2 #(
		.INIT('h2)
	) name7288 (
		_w8288_,
		_w8289_,
		_w8290_
	);
	LUT2 #(
		.INIT('h1)
	) name7289 (
		_w8275_,
		_w8276_,
		_w8291_
	);
	LUT2 #(
		.INIT('h2)
	) name7290 (
		_w8281_,
		_w8291_,
		_w8292_
	);
	LUT2 #(
		.INIT('h4)
	) name7291 (
		_w8281_,
		_w8291_,
		_w8293_
	);
	LUT2 #(
		.INIT('h1)
	) name7292 (
		_w8292_,
		_w8293_,
		_w8294_
	);
	LUT2 #(
		.INIT('h2)
	) name7293 (
		_w8290_,
		_w8294_,
		_w8295_
	);
	LUT2 #(
		.INIT('h4)
	) name7294 (
		_w8290_,
		_w8294_,
		_w8296_
	);
	LUT2 #(
		.INIT('h1)
	) name7295 (
		_w8259_,
		_w8262_,
		_w8297_
	);
	LUT2 #(
		.INIT('h2)
	) name7296 (
		_w8260_,
		_w8297_,
		_w8298_
	);
	LUT2 #(
		.INIT('h4)
	) name7297 (
		_w8260_,
		_w8297_,
		_w8299_
	);
	LUT2 #(
		.INIT('h1)
	) name7298 (
		_w8298_,
		_w8299_,
		_w8300_
	);
	LUT2 #(
		.INIT('h4)
	) name7299 (
		_w8296_,
		_w8300_,
		_w8301_
	);
	LUT2 #(
		.INIT('h1)
	) name7300 (
		_w8295_,
		_w8301_,
		_w8302_
	);
	LUT2 #(
		.INIT('h2)
	) name7301 (
		_w8283_,
		_w8302_,
		_w8303_
	);
	LUT2 #(
		.INIT('h4)
	) name7302 (
		_w8283_,
		_w8302_,
		_w8304_
	);
	LUT2 #(
		.INIT('h1)
	) name7303 (
		_w8303_,
		_w8304_,
		_w8305_
	);
	LUT2 #(
		.INIT('h8)
	) name7304 (
		_w8264_,
		_w8305_,
		_w8306_
	);
	LUT2 #(
		.INIT('h1)
	) name7305 (
		_w8264_,
		_w8305_,
		_w8307_
	);
	LUT2 #(
		.INIT('h1)
	) name7306 (
		_w8306_,
		_w8307_,
		_w8308_
	);
	LUT2 #(
		.INIT('h8)
	) name7307 (
		\A[646] ,
		\A[647] ,
		_w8309_
	);
	LUT2 #(
		.INIT('h8)
	) name7308 (
		\A[643] ,
		\A[644] ,
		_w8310_
	);
	LUT2 #(
		.INIT('h1)
	) name7309 (
		\A[643] ,
		\A[644] ,
		_w8311_
	);
	LUT2 #(
		.INIT('h1)
	) name7310 (
		_w8310_,
		_w8311_,
		_w8312_
	);
	LUT2 #(
		.INIT('h8)
	) name7311 (
		\A[645] ,
		_w8312_,
		_w8313_
	);
	LUT2 #(
		.INIT('h1)
	) name7312 (
		\A[645] ,
		_w8312_,
		_w8314_
	);
	LUT2 #(
		.INIT('h1)
	) name7313 (
		_w8313_,
		_w8314_,
		_w8315_
	);
	LUT2 #(
		.INIT('h1)
	) name7314 (
		\A[646] ,
		\A[647] ,
		_w8316_
	);
	LUT2 #(
		.INIT('h1)
	) name7315 (
		_w8309_,
		_w8316_,
		_w8317_
	);
	LUT2 #(
		.INIT('h8)
	) name7316 (
		\A[648] ,
		_w8317_,
		_w8318_
	);
	LUT2 #(
		.INIT('h1)
	) name7317 (
		\A[648] ,
		_w8317_,
		_w8319_
	);
	LUT2 #(
		.INIT('h1)
	) name7318 (
		_w8318_,
		_w8319_,
		_w8320_
	);
	LUT2 #(
		.INIT('h8)
	) name7319 (
		_w8315_,
		_w8320_,
		_w8321_
	);
	LUT2 #(
		.INIT('h8)
	) name7320 (
		_w8309_,
		_w8321_,
		_w8322_
	);
	LUT2 #(
		.INIT('h1)
	) name7321 (
		_w8310_,
		_w8313_,
		_w8323_
	);
	LUT2 #(
		.INIT('h1)
	) name7322 (
		_w8309_,
		_w8318_,
		_w8324_
	);
	LUT2 #(
		.INIT('h4)
	) name7323 (
		_w8321_,
		_w8324_,
		_w8325_
	);
	LUT2 #(
		.INIT('h1)
	) name7324 (
		_w8323_,
		_w8325_,
		_w8326_
	);
	LUT2 #(
		.INIT('h1)
	) name7325 (
		_w8322_,
		_w8326_,
		_w8327_
	);
	LUT2 #(
		.INIT('h8)
	) name7326 (
		\A[652] ,
		\A[653] ,
		_w8328_
	);
	LUT2 #(
		.INIT('h1)
	) name7327 (
		\A[652] ,
		\A[653] ,
		_w8329_
	);
	LUT2 #(
		.INIT('h1)
	) name7328 (
		_w8328_,
		_w8329_,
		_w8330_
	);
	LUT2 #(
		.INIT('h8)
	) name7329 (
		\A[654] ,
		_w8330_,
		_w8331_
	);
	LUT2 #(
		.INIT('h1)
	) name7330 (
		_w8328_,
		_w8331_,
		_w8332_
	);
	LUT2 #(
		.INIT('h8)
	) name7331 (
		\A[649] ,
		\A[650] ,
		_w8333_
	);
	LUT2 #(
		.INIT('h1)
	) name7332 (
		\A[649] ,
		\A[650] ,
		_w8334_
	);
	LUT2 #(
		.INIT('h1)
	) name7333 (
		_w8333_,
		_w8334_,
		_w8335_
	);
	LUT2 #(
		.INIT('h8)
	) name7334 (
		\A[651] ,
		_w8335_,
		_w8336_
	);
	LUT2 #(
		.INIT('h1)
	) name7335 (
		_w8333_,
		_w8336_,
		_w8337_
	);
	LUT2 #(
		.INIT('h8)
	) name7336 (
		_w8332_,
		_w8337_,
		_w8338_
	);
	LUT2 #(
		.INIT('h1)
	) name7337 (
		_w8332_,
		_w8337_,
		_w8339_
	);
	LUT2 #(
		.INIT('h1)
	) name7338 (
		\A[651] ,
		_w8335_,
		_w8340_
	);
	LUT2 #(
		.INIT('h1)
	) name7339 (
		_w8336_,
		_w8340_,
		_w8341_
	);
	LUT2 #(
		.INIT('h1)
	) name7340 (
		\A[654] ,
		_w8330_,
		_w8342_
	);
	LUT2 #(
		.INIT('h1)
	) name7341 (
		_w8331_,
		_w8342_,
		_w8343_
	);
	LUT2 #(
		.INIT('h8)
	) name7342 (
		_w8341_,
		_w8343_,
		_w8344_
	);
	LUT2 #(
		.INIT('h1)
	) name7343 (
		_w8339_,
		_w8344_,
		_w8345_
	);
	LUT2 #(
		.INIT('h1)
	) name7344 (
		_w8338_,
		_w8345_,
		_w8346_
	);
	LUT2 #(
		.INIT('h1)
	) name7345 (
		_w8341_,
		_w8343_,
		_w8347_
	);
	LUT2 #(
		.INIT('h1)
	) name7346 (
		_w8344_,
		_w8347_,
		_w8348_
	);
	LUT2 #(
		.INIT('h1)
	) name7347 (
		_w8315_,
		_w8320_,
		_w8349_
	);
	LUT2 #(
		.INIT('h1)
	) name7348 (
		_w8321_,
		_w8349_,
		_w8350_
	);
	LUT2 #(
		.INIT('h8)
	) name7349 (
		_w8348_,
		_w8350_,
		_w8351_
	);
	LUT2 #(
		.INIT('h2)
	) name7350 (
		_w8322_,
		_w8323_,
		_w8352_
	);
	LUT2 #(
		.INIT('h2)
	) name7351 (
		_w8351_,
		_w8352_,
		_w8353_
	);
	LUT2 #(
		.INIT('h1)
	) name7352 (
		_w8338_,
		_w8339_,
		_w8354_
	);
	LUT2 #(
		.INIT('h2)
	) name7353 (
		_w8344_,
		_w8354_,
		_w8355_
	);
	LUT2 #(
		.INIT('h4)
	) name7354 (
		_w8344_,
		_w8354_,
		_w8356_
	);
	LUT2 #(
		.INIT('h1)
	) name7355 (
		_w8355_,
		_w8356_,
		_w8357_
	);
	LUT2 #(
		.INIT('h2)
	) name7356 (
		_w8353_,
		_w8357_,
		_w8358_
	);
	LUT2 #(
		.INIT('h4)
	) name7357 (
		_w8353_,
		_w8357_,
		_w8359_
	);
	LUT2 #(
		.INIT('h1)
	) name7358 (
		_w8322_,
		_w8325_,
		_w8360_
	);
	LUT2 #(
		.INIT('h2)
	) name7359 (
		_w8323_,
		_w8360_,
		_w8361_
	);
	LUT2 #(
		.INIT('h4)
	) name7360 (
		_w8323_,
		_w8360_,
		_w8362_
	);
	LUT2 #(
		.INIT('h1)
	) name7361 (
		_w8361_,
		_w8362_,
		_w8363_
	);
	LUT2 #(
		.INIT('h4)
	) name7362 (
		_w8359_,
		_w8363_,
		_w8364_
	);
	LUT2 #(
		.INIT('h1)
	) name7363 (
		_w8358_,
		_w8364_,
		_w8365_
	);
	LUT2 #(
		.INIT('h2)
	) name7364 (
		_w8346_,
		_w8365_,
		_w8366_
	);
	LUT2 #(
		.INIT('h4)
	) name7365 (
		_w8346_,
		_w8365_,
		_w8367_
	);
	LUT2 #(
		.INIT('h1)
	) name7366 (
		_w8366_,
		_w8367_,
		_w8368_
	);
	LUT2 #(
		.INIT('h8)
	) name7367 (
		_w8327_,
		_w8368_,
		_w8369_
	);
	LUT2 #(
		.INIT('h1)
	) name7368 (
		_w8327_,
		_w8368_,
		_w8370_
	);
	LUT2 #(
		.INIT('h1)
	) name7369 (
		_w8369_,
		_w8370_,
		_w8371_
	);
	LUT2 #(
		.INIT('h1)
	) name7370 (
		_w8308_,
		_w8371_,
		_w8372_
	);
	LUT2 #(
		.INIT('h8)
	) name7371 (
		_w8308_,
		_w8371_,
		_w8373_
	);
	LUT2 #(
		.INIT('h1)
	) name7372 (
		_w8348_,
		_w8350_,
		_w8374_
	);
	LUT2 #(
		.INIT('h1)
	) name7373 (
		_w8351_,
		_w8374_,
		_w8375_
	);
	LUT2 #(
		.INIT('h1)
	) name7374 (
		_w8285_,
		_w8287_,
		_w8376_
	);
	LUT2 #(
		.INIT('h1)
	) name7375 (
		_w8288_,
		_w8376_,
		_w8377_
	);
	LUT2 #(
		.INIT('h8)
	) name7376 (
		_w8375_,
		_w8377_,
		_w8378_
	);
	LUT2 #(
		.INIT('h1)
	) name7377 (
		_w8358_,
		_w8359_,
		_w8379_
	);
	LUT2 #(
		.INIT('h8)
	) name7378 (
		_w8363_,
		_w8379_,
		_w8380_
	);
	LUT2 #(
		.INIT('h1)
	) name7379 (
		_w8363_,
		_w8379_,
		_w8381_
	);
	LUT2 #(
		.INIT('h1)
	) name7380 (
		_w8380_,
		_w8381_,
		_w8382_
	);
	LUT2 #(
		.INIT('h8)
	) name7381 (
		_w8378_,
		_w8382_,
		_w8383_
	);
	LUT2 #(
		.INIT('h1)
	) name7382 (
		_w8378_,
		_w8382_,
		_w8384_
	);
	LUT2 #(
		.INIT('h1)
	) name7383 (
		_w8295_,
		_w8296_,
		_w8385_
	);
	LUT2 #(
		.INIT('h8)
	) name7384 (
		_w8300_,
		_w8385_,
		_w8386_
	);
	LUT2 #(
		.INIT('h1)
	) name7385 (
		_w8300_,
		_w8385_,
		_w8387_
	);
	LUT2 #(
		.INIT('h1)
	) name7386 (
		_w8386_,
		_w8387_,
		_w8388_
	);
	LUT2 #(
		.INIT('h4)
	) name7387 (
		_w8384_,
		_w8388_,
		_w8389_
	);
	LUT2 #(
		.INIT('h1)
	) name7388 (
		_w8383_,
		_w8389_,
		_w8390_
	);
	LUT2 #(
		.INIT('h1)
	) name7389 (
		_w8373_,
		_w8390_,
		_w8391_
	);
	LUT2 #(
		.INIT('h1)
	) name7390 (
		_w8372_,
		_w8391_,
		_w8392_
	);
	LUT2 #(
		.INIT('h1)
	) name7391 (
		_w8327_,
		_w8367_,
		_w8393_
	);
	LUT2 #(
		.INIT('h1)
	) name7392 (
		_w8366_,
		_w8393_,
		_w8394_
	);
	LUT2 #(
		.INIT('h1)
	) name7393 (
		_w8392_,
		_w8394_,
		_w8395_
	);
	LUT2 #(
		.INIT('h8)
	) name7394 (
		_w8392_,
		_w8394_,
		_w8396_
	);
	LUT2 #(
		.INIT('h1)
	) name7395 (
		_w8264_,
		_w8304_,
		_w8397_
	);
	LUT2 #(
		.INIT('h1)
	) name7396 (
		_w8303_,
		_w8397_,
		_w8398_
	);
	LUT2 #(
		.INIT('h1)
	) name7397 (
		_w8396_,
		_w8398_,
		_w8399_
	);
	LUT2 #(
		.INIT('h1)
	) name7398 (
		_w8395_,
		_w8399_,
		_w8400_
	);
	LUT2 #(
		.INIT('h1)
	) name7399 (
		_w8395_,
		_w8396_,
		_w8401_
	);
	LUT2 #(
		.INIT('h4)
	) name7400 (
		_w8398_,
		_w8401_,
		_w8402_
	);
	LUT2 #(
		.INIT('h2)
	) name7401 (
		_w8398_,
		_w8401_,
		_w8403_
	);
	LUT2 #(
		.INIT('h1)
	) name7402 (
		_w8402_,
		_w8403_,
		_w8404_
	);
	LUT2 #(
		.INIT('h8)
	) name7403 (
		\A[610] ,
		\A[611] ,
		_w8405_
	);
	LUT2 #(
		.INIT('h8)
	) name7404 (
		\A[607] ,
		\A[608] ,
		_w8406_
	);
	LUT2 #(
		.INIT('h1)
	) name7405 (
		\A[607] ,
		\A[608] ,
		_w8407_
	);
	LUT2 #(
		.INIT('h1)
	) name7406 (
		_w8406_,
		_w8407_,
		_w8408_
	);
	LUT2 #(
		.INIT('h8)
	) name7407 (
		\A[609] ,
		_w8408_,
		_w8409_
	);
	LUT2 #(
		.INIT('h1)
	) name7408 (
		\A[609] ,
		_w8408_,
		_w8410_
	);
	LUT2 #(
		.INIT('h1)
	) name7409 (
		_w8409_,
		_w8410_,
		_w8411_
	);
	LUT2 #(
		.INIT('h1)
	) name7410 (
		\A[610] ,
		\A[611] ,
		_w8412_
	);
	LUT2 #(
		.INIT('h1)
	) name7411 (
		_w8405_,
		_w8412_,
		_w8413_
	);
	LUT2 #(
		.INIT('h8)
	) name7412 (
		\A[612] ,
		_w8413_,
		_w8414_
	);
	LUT2 #(
		.INIT('h1)
	) name7413 (
		\A[612] ,
		_w8413_,
		_w8415_
	);
	LUT2 #(
		.INIT('h1)
	) name7414 (
		_w8414_,
		_w8415_,
		_w8416_
	);
	LUT2 #(
		.INIT('h8)
	) name7415 (
		_w8411_,
		_w8416_,
		_w8417_
	);
	LUT2 #(
		.INIT('h8)
	) name7416 (
		_w8405_,
		_w8417_,
		_w8418_
	);
	LUT2 #(
		.INIT('h1)
	) name7417 (
		_w8406_,
		_w8409_,
		_w8419_
	);
	LUT2 #(
		.INIT('h1)
	) name7418 (
		_w8405_,
		_w8414_,
		_w8420_
	);
	LUT2 #(
		.INIT('h4)
	) name7419 (
		_w8417_,
		_w8420_,
		_w8421_
	);
	LUT2 #(
		.INIT('h1)
	) name7420 (
		_w8419_,
		_w8421_,
		_w8422_
	);
	LUT2 #(
		.INIT('h1)
	) name7421 (
		_w8418_,
		_w8422_,
		_w8423_
	);
	LUT2 #(
		.INIT('h8)
	) name7422 (
		\A[616] ,
		\A[617] ,
		_w8424_
	);
	LUT2 #(
		.INIT('h1)
	) name7423 (
		\A[616] ,
		\A[617] ,
		_w8425_
	);
	LUT2 #(
		.INIT('h1)
	) name7424 (
		_w8424_,
		_w8425_,
		_w8426_
	);
	LUT2 #(
		.INIT('h8)
	) name7425 (
		\A[618] ,
		_w8426_,
		_w8427_
	);
	LUT2 #(
		.INIT('h1)
	) name7426 (
		_w8424_,
		_w8427_,
		_w8428_
	);
	LUT2 #(
		.INIT('h8)
	) name7427 (
		\A[613] ,
		\A[614] ,
		_w8429_
	);
	LUT2 #(
		.INIT('h1)
	) name7428 (
		\A[613] ,
		\A[614] ,
		_w8430_
	);
	LUT2 #(
		.INIT('h1)
	) name7429 (
		_w8429_,
		_w8430_,
		_w8431_
	);
	LUT2 #(
		.INIT('h8)
	) name7430 (
		\A[615] ,
		_w8431_,
		_w8432_
	);
	LUT2 #(
		.INIT('h1)
	) name7431 (
		_w8429_,
		_w8432_,
		_w8433_
	);
	LUT2 #(
		.INIT('h8)
	) name7432 (
		_w8428_,
		_w8433_,
		_w8434_
	);
	LUT2 #(
		.INIT('h1)
	) name7433 (
		_w8428_,
		_w8433_,
		_w8435_
	);
	LUT2 #(
		.INIT('h1)
	) name7434 (
		\A[615] ,
		_w8431_,
		_w8436_
	);
	LUT2 #(
		.INIT('h1)
	) name7435 (
		_w8432_,
		_w8436_,
		_w8437_
	);
	LUT2 #(
		.INIT('h1)
	) name7436 (
		\A[618] ,
		_w8426_,
		_w8438_
	);
	LUT2 #(
		.INIT('h1)
	) name7437 (
		_w8427_,
		_w8438_,
		_w8439_
	);
	LUT2 #(
		.INIT('h8)
	) name7438 (
		_w8437_,
		_w8439_,
		_w8440_
	);
	LUT2 #(
		.INIT('h1)
	) name7439 (
		_w8435_,
		_w8440_,
		_w8441_
	);
	LUT2 #(
		.INIT('h1)
	) name7440 (
		_w8434_,
		_w8441_,
		_w8442_
	);
	LUT2 #(
		.INIT('h1)
	) name7441 (
		_w8437_,
		_w8439_,
		_w8443_
	);
	LUT2 #(
		.INIT('h1)
	) name7442 (
		_w8440_,
		_w8443_,
		_w8444_
	);
	LUT2 #(
		.INIT('h1)
	) name7443 (
		_w8411_,
		_w8416_,
		_w8445_
	);
	LUT2 #(
		.INIT('h1)
	) name7444 (
		_w8417_,
		_w8445_,
		_w8446_
	);
	LUT2 #(
		.INIT('h8)
	) name7445 (
		_w8444_,
		_w8446_,
		_w8447_
	);
	LUT2 #(
		.INIT('h2)
	) name7446 (
		_w8418_,
		_w8419_,
		_w8448_
	);
	LUT2 #(
		.INIT('h2)
	) name7447 (
		_w8447_,
		_w8448_,
		_w8449_
	);
	LUT2 #(
		.INIT('h1)
	) name7448 (
		_w8434_,
		_w8435_,
		_w8450_
	);
	LUT2 #(
		.INIT('h2)
	) name7449 (
		_w8440_,
		_w8450_,
		_w8451_
	);
	LUT2 #(
		.INIT('h4)
	) name7450 (
		_w8440_,
		_w8450_,
		_w8452_
	);
	LUT2 #(
		.INIT('h1)
	) name7451 (
		_w8451_,
		_w8452_,
		_w8453_
	);
	LUT2 #(
		.INIT('h2)
	) name7452 (
		_w8449_,
		_w8453_,
		_w8454_
	);
	LUT2 #(
		.INIT('h4)
	) name7453 (
		_w8449_,
		_w8453_,
		_w8455_
	);
	LUT2 #(
		.INIT('h1)
	) name7454 (
		_w8418_,
		_w8421_,
		_w8456_
	);
	LUT2 #(
		.INIT('h2)
	) name7455 (
		_w8419_,
		_w8456_,
		_w8457_
	);
	LUT2 #(
		.INIT('h4)
	) name7456 (
		_w8419_,
		_w8456_,
		_w8458_
	);
	LUT2 #(
		.INIT('h1)
	) name7457 (
		_w8457_,
		_w8458_,
		_w8459_
	);
	LUT2 #(
		.INIT('h4)
	) name7458 (
		_w8455_,
		_w8459_,
		_w8460_
	);
	LUT2 #(
		.INIT('h1)
	) name7459 (
		_w8454_,
		_w8460_,
		_w8461_
	);
	LUT2 #(
		.INIT('h2)
	) name7460 (
		_w8442_,
		_w8461_,
		_w8462_
	);
	LUT2 #(
		.INIT('h4)
	) name7461 (
		_w8442_,
		_w8461_,
		_w8463_
	);
	LUT2 #(
		.INIT('h1)
	) name7462 (
		_w8462_,
		_w8463_,
		_w8464_
	);
	LUT2 #(
		.INIT('h8)
	) name7463 (
		_w8423_,
		_w8464_,
		_w8465_
	);
	LUT2 #(
		.INIT('h1)
	) name7464 (
		_w8423_,
		_w8464_,
		_w8466_
	);
	LUT2 #(
		.INIT('h1)
	) name7465 (
		_w8465_,
		_w8466_,
		_w8467_
	);
	LUT2 #(
		.INIT('h8)
	) name7466 (
		\A[622] ,
		\A[623] ,
		_w8468_
	);
	LUT2 #(
		.INIT('h8)
	) name7467 (
		\A[619] ,
		\A[620] ,
		_w8469_
	);
	LUT2 #(
		.INIT('h1)
	) name7468 (
		\A[619] ,
		\A[620] ,
		_w8470_
	);
	LUT2 #(
		.INIT('h1)
	) name7469 (
		_w8469_,
		_w8470_,
		_w8471_
	);
	LUT2 #(
		.INIT('h8)
	) name7470 (
		\A[621] ,
		_w8471_,
		_w8472_
	);
	LUT2 #(
		.INIT('h1)
	) name7471 (
		\A[621] ,
		_w8471_,
		_w8473_
	);
	LUT2 #(
		.INIT('h1)
	) name7472 (
		_w8472_,
		_w8473_,
		_w8474_
	);
	LUT2 #(
		.INIT('h1)
	) name7473 (
		\A[622] ,
		\A[623] ,
		_w8475_
	);
	LUT2 #(
		.INIT('h1)
	) name7474 (
		_w8468_,
		_w8475_,
		_w8476_
	);
	LUT2 #(
		.INIT('h8)
	) name7475 (
		\A[624] ,
		_w8476_,
		_w8477_
	);
	LUT2 #(
		.INIT('h1)
	) name7476 (
		\A[624] ,
		_w8476_,
		_w8478_
	);
	LUT2 #(
		.INIT('h1)
	) name7477 (
		_w8477_,
		_w8478_,
		_w8479_
	);
	LUT2 #(
		.INIT('h8)
	) name7478 (
		_w8474_,
		_w8479_,
		_w8480_
	);
	LUT2 #(
		.INIT('h8)
	) name7479 (
		_w8468_,
		_w8480_,
		_w8481_
	);
	LUT2 #(
		.INIT('h1)
	) name7480 (
		_w8469_,
		_w8472_,
		_w8482_
	);
	LUT2 #(
		.INIT('h1)
	) name7481 (
		_w8468_,
		_w8477_,
		_w8483_
	);
	LUT2 #(
		.INIT('h4)
	) name7482 (
		_w8480_,
		_w8483_,
		_w8484_
	);
	LUT2 #(
		.INIT('h1)
	) name7483 (
		_w8482_,
		_w8484_,
		_w8485_
	);
	LUT2 #(
		.INIT('h1)
	) name7484 (
		_w8481_,
		_w8485_,
		_w8486_
	);
	LUT2 #(
		.INIT('h8)
	) name7485 (
		\A[628] ,
		\A[629] ,
		_w8487_
	);
	LUT2 #(
		.INIT('h1)
	) name7486 (
		\A[628] ,
		\A[629] ,
		_w8488_
	);
	LUT2 #(
		.INIT('h1)
	) name7487 (
		_w8487_,
		_w8488_,
		_w8489_
	);
	LUT2 #(
		.INIT('h8)
	) name7488 (
		\A[630] ,
		_w8489_,
		_w8490_
	);
	LUT2 #(
		.INIT('h1)
	) name7489 (
		_w8487_,
		_w8490_,
		_w8491_
	);
	LUT2 #(
		.INIT('h8)
	) name7490 (
		\A[625] ,
		\A[626] ,
		_w8492_
	);
	LUT2 #(
		.INIT('h1)
	) name7491 (
		\A[625] ,
		\A[626] ,
		_w8493_
	);
	LUT2 #(
		.INIT('h1)
	) name7492 (
		_w8492_,
		_w8493_,
		_w8494_
	);
	LUT2 #(
		.INIT('h8)
	) name7493 (
		\A[627] ,
		_w8494_,
		_w8495_
	);
	LUT2 #(
		.INIT('h1)
	) name7494 (
		_w8492_,
		_w8495_,
		_w8496_
	);
	LUT2 #(
		.INIT('h8)
	) name7495 (
		_w8491_,
		_w8496_,
		_w8497_
	);
	LUT2 #(
		.INIT('h1)
	) name7496 (
		_w8491_,
		_w8496_,
		_w8498_
	);
	LUT2 #(
		.INIT('h1)
	) name7497 (
		\A[627] ,
		_w8494_,
		_w8499_
	);
	LUT2 #(
		.INIT('h1)
	) name7498 (
		_w8495_,
		_w8499_,
		_w8500_
	);
	LUT2 #(
		.INIT('h1)
	) name7499 (
		\A[630] ,
		_w8489_,
		_w8501_
	);
	LUT2 #(
		.INIT('h1)
	) name7500 (
		_w8490_,
		_w8501_,
		_w8502_
	);
	LUT2 #(
		.INIT('h8)
	) name7501 (
		_w8500_,
		_w8502_,
		_w8503_
	);
	LUT2 #(
		.INIT('h1)
	) name7502 (
		_w8498_,
		_w8503_,
		_w8504_
	);
	LUT2 #(
		.INIT('h1)
	) name7503 (
		_w8497_,
		_w8504_,
		_w8505_
	);
	LUT2 #(
		.INIT('h1)
	) name7504 (
		_w8500_,
		_w8502_,
		_w8506_
	);
	LUT2 #(
		.INIT('h1)
	) name7505 (
		_w8503_,
		_w8506_,
		_w8507_
	);
	LUT2 #(
		.INIT('h1)
	) name7506 (
		_w8474_,
		_w8479_,
		_w8508_
	);
	LUT2 #(
		.INIT('h1)
	) name7507 (
		_w8480_,
		_w8508_,
		_w8509_
	);
	LUT2 #(
		.INIT('h8)
	) name7508 (
		_w8507_,
		_w8509_,
		_w8510_
	);
	LUT2 #(
		.INIT('h2)
	) name7509 (
		_w8481_,
		_w8482_,
		_w8511_
	);
	LUT2 #(
		.INIT('h2)
	) name7510 (
		_w8510_,
		_w8511_,
		_w8512_
	);
	LUT2 #(
		.INIT('h1)
	) name7511 (
		_w8497_,
		_w8498_,
		_w8513_
	);
	LUT2 #(
		.INIT('h2)
	) name7512 (
		_w8503_,
		_w8513_,
		_w8514_
	);
	LUT2 #(
		.INIT('h4)
	) name7513 (
		_w8503_,
		_w8513_,
		_w8515_
	);
	LUT2 #(
		.INIT('h1)
	) name7514 (
		_w8514_,
		_w8515_,
		_w8516_
	);
	LUT2 #(
		.INIT('h2)
	) name7515 (
		_w8512_,
		_w8516_,
		_w8517_
	);
	LUT2 #(
		.INIT('h4)
	) name7516 (
		_w8512_,
		_w8516_,
		_w8518_
	);
	LUT2 #(
		.INIT('h1)
	) name7517 (
		_w8481_,
		_w8484_,
		_w8519_
	);
	LUT2 #(
		.INIT('h2)
	) name7518 (
		_w8482_,
		_w8519_,
		_w8520_
	);
	LUT2 #(
		.INIT('h4)
	) name7519 (
		_w8482_,
		_w8519_,
		_w8521_
	);
	LUT2 #(
		.INIT('h1)
	) name7520 (
		_w8520_,
		_w8521_,
		_w8522_
	);
	LUT2 #(
		.INIT('h4)
	) name7521 (
		_w8518_,
		_w8522_,
		_w8523_
	);
	LUT2 #(
		.INIT('h1)
	) name7522 (
		_w8517_,
		_w8523_,
		_w8524_
	);
	LUT2 #(
		.INIT('h2)
	) name7523 (
		_w8505_,
		_w8524_,
		_w8525_
	);
	LUT2 #(
		.INIT('h4)
	) name7524 (
		_w8505_,
		_w8524_,
		_w8526_
	);
	LUT2 #(
		.INIT('h1)
	) name7525 (
		_w8525_,
		_w8526_,
		_w8527_
	);
	LUT2 #(
		.INIT('h8)
	) name7526 (
		_w8486_,
		_w8527_,
		_w8528_
	);
	LUT2 #(
		.INIT('h1)
	) name7527 (
		_w8486_,
		_w8527_,
		_w8529_
	);
	LUT2 #(
		.INIT('h1)
	) name7528 (
		_w8528_,
		_w8529_,
		_w8530_
	);
	LUT2 #(
		.INIT('h1)
	) name7529 (
		_w8467_,
		_w8530_,
		_w8531_
	);
	LUT2 #(
		.INIT('h8)
	) name7530 (
		_w8467_,
		_w8530_,
		_w8532_
	);
	LUT2 #(
		.INIT('h1)
	) name7531 (
		_w8507_,
		_w8509_,
		_w8533_
	);
	LUT2 #(
		.INIT('h1)
	) name7532 (
		_w8510_,
		_w8533_,
		_w8534_
	);
	LUT2 #(
		.INIT('h1)
	) name7533 (
		_w8444_,
		_w8446_,
		_w8535_
	);
	LUT2 #(
		.INIT('h1)
	) name7534 (
		_w8447_,
		_w8535_,
		_w8536_
	);
	LUT2 #(
		.INIT('h8)
	) name7535 (
		_w8534_,
		_w8536_,
		_w8537_
	);
	LUT2 #(
		.INIT('h1)
	) name7536 (
		_w8517_,
		_w8518_,
		_w8538_
	);
	LUT2 #(
		.INIT('h8)
	) name7537 (
		_w8522_,
		_w8538_,
		_w8539_
	);
	LUT2 #(
		.INIT('h1)
	) name7538 (
		_w8522_,
		_w8538_,
		_w8540_
	);
	LUT2 #(
		.INIT('h1)
	) name7539 (
		_w8539_,
		_w8540_,
		_w8541_
	);
	LUT2 #(
		.INIT('h8)
	) name7540 (
		_w8537_,
		_w8541_,
		_w8542_
	);
	LUT2 #(
		.INIT('h1)
	) name7541 (
		_w8537_,
		_w8541_,
		_w8543_
	);
	LUT2 #(
		.INIT('h1)
	) name7542 (
		_w8454_,
		_w8455_,
		_w8544_
	);
	LUT2 #(
		.INIT('h8)
	) name7543 (
		_w8459_,
		_w8544_,
		_w8545_
	);
	LUT2 #(
		.INIT('h1)
	) name7544 (
		_w8459_,
		_w8544_,
		_w8546_
	);
	LUT2 #(
		.INIT('h1)
	) name7545 (
		_w8545_,
		_w8546_,
		_w8547_
	);
	LUT2 #(
		.INIT('h4)
	) name7546 (
		_w8543_,
		_w8547_,
		_w8548_
	);
	LUT2 #(
		.INIT('h1)
	) name7547 (
		_w8542_,
		_w8548_,
		_w8549_
	);
	LUT2 #(
		.INIT('h1)
	) name7548 (
		_w8532_,
		_w8549_,
		_w8550_
	);
	LUT2 #(
		.INIT('h1)
	) name7549 (
		_w8531_,
		_w8550_,
		_w8551_
	);
	LUT2 #(
		.INIT('h1)
	) name7550 (
		_w8486_,
		_w8526_,
		_w8552_
	);
	LUT2 #(
		.INIT('h1)
	) name7551 (
		_w8525_,
		_w8552_,
		_w8553_
	);
	LUT2 #(
		.INIT('h1)
	) name7552 (
		_w8551_,
		_w8553_,
		_w8554_
	);
	LUT2 #(
		.INIT('h8)
	) name7553 (
		_w8551_,
		_w8553_,
		_w8555_
	);
	LUT2 #(
		.INIT('h1)
	) name7554 (
		_w8554_,
		_w8555_,
		_w8556_
	);
	LUT2 #(
		.INIT('h1)
	) name7555 (
		_w8423_,
		_w8463_,
		_w8557_
	);
	LUT2 #(
		.INIT('h1)
	) name7556 (
		_w8462_,
		_w8557_,
		_w8558_
	);
	LUT2 #(
		.INIT('h2)
	) name7557 (
		_w8556_,
		_w8558_,
		_w8559_
	);
	LUT2 #(
		.INIT('h4)
	) name7558 (
		_w8556_,
		_w8558_,
		_w8560_
	);
	LUT2 #(
		.INIT('h1)
	) name7559 (
		_w8559_,
		_w8560_,
		_w8561_
	);
	LUT2 #(
		.INIT('h1)
	) name7560 (
		_w8404_,
		_w8561_,
		_w8562_
	);
	LUT2 #(
		.INIT('h8)
	) name7561 (
		_w8404_,
		_w8561_,
		_w8563_
	);
	LUT2 #(
		.INIT('h1)
	) name7562 (
		_w8531_,
		_w8532_,
		_w8564_
	);
	LUT2 #(
		.INIT('h4)
	) name7563 (
		_w8549_,
		_w8564_,
		_w8565_
	);
	LUT2 #(
		.INIT('h2)
	) name7564 (
		_w8549_,
		_w8564_,
		_w8566_
	);
	LUT2 #(
		.INIT('h1)
	) name7565 (
		_w8565_,
		_w8566_,
		_w8567_
	);
	LUT2 #(
		.INIT('h1)
	) name7566 (
		_w8372_,
		_w8373_,
		_w8568_
	);
	LUT2 #(
		.INIT('h4)
	) name7567 (
		_w8390_,
		_w8568_,
		_w8569_
	);
	LUT2 #(
		.INIT('h2)
	) name7568 (
		_w8390_,
		_w8568_,
		_w8570_
	);
	LUT2 #(
		.INIT('h1)
	) name7569 (
		_w8569_,
		_w8570_,
		_w8571_
	);
	LUT2 #(
		.INIT('h1)
	) name7570 (
		_w8567_,
		_w8571_,
		_w8572_
	);
	LUT2 #(
		.INIT('h8)
	) name7571 (
		_w8567_,
		_w8571_,
		_w8573_
	);
	LUT2 #(
		.INIT('h1)
	) name7572 (
		_w8375_,
		_w8377_,
		_w8574_
	);
	LUT2 #(
		.INIT('h1)
	) name7573 (
		_w8378_,
		_w8574_,
		_w8575_
	);
	LUT2 #(
		.INIT('h1)
	) name7574 (
		_w8534_,
		_w8536_,
		_w8576_
	);
	LUT2 #(
		.INIT('h1)
	) name7575 (
		_w8537_,
		_w8576_,
		_w8577_
	);
	LUT2 #(
		.INIT('h8)
	) name7576 (
		_w8575_,
		_w8577_,
		_w8578_
	);
	LUT2 #(
		.INIT('h1)
	) name7577 (
		_w8383_,
		_w8384_,
		_w8579_
	);
	LUT2 #(
		.INIT('h4)
	) name7578 (
		_w8388_,
		_w8579_,
		_w8580_
	);
	LUT2 #(
		.INIT('h2)
	) name7579 (
		_w8388_,
		_w8579_,
		_w8581_
	);
	LUT2 #(
		.INIT('h1)
	) name7580 (
		_w8580_,
		_w8581_,
		_w8582_
	);
	LUT2 #(
		.INIT('h2)
	) name7581 (
		_w8578_,
		_w8582_,
		_w8583_
	);
	LUT2 #(
		.INIT('h4)
	) name7582 (
		_w8578_,
		_w8582_,
		_w8584_
	);
	LUT2 #(
		.INIT('h1)
	) name7583 (
		_w8542_,
		_w8543_,
		_w8585_
	);
	LUT2 #(
		.INIT('h4)
	) name7584 (
		_w8547_,
		_w8585_,
		_w8586_
	);
	LUT2 #(
		.INIT('h2)
	) name7585 (
		_w8547_,
		_w8585_,
		_w8587_
	);
	LUT2 #(
		.INIT('h1)
	) name7586 (
		_w8586_,
		_w8587_,
		_w8588_
	);
	LUT2 #(
		.INIT('h1)
	) name7587 (
		_w8584_,
		_w8588_,
		_w8589_
	);
	LUT2 #(
		.INIT('h1)
	) name7588 (
		_w8583_,
		_w8589_,
		_w8590_
	);
	LUT2 #(
		.INIT('h4)
	) name7589 (
		_w8573_,
		_w8590_,
		_w8591_
	);
	LUT2 #(
		.INIT('h1)
	) name7590 (
		_w8572_,
		_w8591_,
		_w8592_
	);
	LUT2 #(
		.INIT('h1)
	) name7591 (
		_w8563_,
		_w8592_,
		_w8593_
	);
	LUT2 #(
		.INIT('h1)
	) name7592 (
		_w8562_,
		_w8593_,
		_w8594_
	);
	LUT2 #(
		.INIT('h2)
	) name7593 (
		_w8400_,
		_w8594_,
		_w8595_
	);
	LUT2 #(
		.INIT('h4)
	) name7594 (
		_w8400_,
		_w8594_,
		_w8596_
	);
	LUT2 #(
		.INIT('h1)
	) name7595 (
		_w8595_,
		_w8596_,
		_w8597_
	);
	LUT2 #(
		.INIT('h1)
	) name7596 (
		_w8555_,
		_w8558_,
		_w8598_
	);
	LUT2 #(
		.INIT('h1)
	) name7597 (
		_w8554_,
		_w8598_,
		_w8599_
	);
	LUT2 #(
		.INIT('h8)
	) name7598 (
		_w8597_,
		_w8599_,
		_w8600_
	);
	LUT2 #(
		.INIT('h1)
	) name7599 (
		_w8597_,
		_w8599_,
		_w8601_
	);
	LUT2 #(
		.INIT('h1)
	) name7600 (
		_w8600_,
		_w8601_,
		_w8602_
	);
	LUT2 #(
		.INIT('h1)
	) name7601 (
		_w8245_,
		_w8602_,
		_w8603_
	);
	LUT2 #(
		.INIT('h8)
	) name7602 (
		_w8245_,
		_w8602_,
		_w8604_
	);
	LUT2 #(
		.INIT('h1)
	) name7603 (
		_w8562_,
		_w8563_,
		_w8605_
	);
	LUT2 #(
		.INIT('h4)
	) name7604 (
		_w8592_,
		_w8605_,
		_w8606_
	);
	LUT2 #(
		.INIT('h2)
	) name7605 (
		_w8592_,
		_w8605_,
		_w8607_
	);
	LUT2 #(
		.INIT('h1)
	) name7606 (
		_w8606_,
		_w8607_,
		_w8608_
	);
	LUT2 #(
		.INIT('h1)
	) name7607 (
		_w8205_,
		_w8206_,
		_w8609_
	);
	LUT2 #(
		.INIT('h4)
	) name7608 (
		_w8235_,
		_w8609_,
		_w8610_
	);
	LUT2 #(
		.INIT('h2)
	) name7609 (
		_w8235_,
		_w8609_,
		_w8611_
	);
	LUT2 #(
		.INIT('h1)
	) name7610 (
		_w8610_,
		_w8611_,
		_w8612_
	);
	LUT2 #(
		.INIT('h1)
	) name7611 (
		_w8608_,
		_w8612_,
		_w8613_
	);
	LUT2 #(
		.INIT('h8)
	) name7612 (
		_w8608_,
		_w8612_,
		_w8614_
	);
	LUT2 #(
		.INIT('h1)
	) name7613 (
		_w8215_,
		_w8216_,
		_w8615_
	);
	LUT2 #(
		.INIT('h4)
	) name7614 (
		_w8233_,
		_w8615_,
		_w8616_
	);
	LUT2 #(
		.INIT('h2)
	) name7615 (
		_w8233_,
		_w8615_,
		_w8617_
	);
	LUT2 #(
		.INIT('h1)
	) name7616 (
		_w8616_,
		_w8617_,
		_w8618_
	);
	LUT2 #(
		.INIT('h1)
	) name7617 (
		_w8572_,
		_w8573_,
		_w8619_
	);
	LUT2 #(
		.INIT('h4)
	) name7618 (
		_w8590_,
		_w8619_,
		_w8620_
	);
	LUT2 #(
		.INIT('h2)
	) name7619 (
		_w8590_,
		_w8619_,
		_w8621_
	);
	LUT2 #(
		.INIT('h1)
	) name7620 (
		_w8620_,
		_w8621_,
		_w8622_
	);
	LUT2 #(
		.INIT('h1)
	) name7621 (
		_w8618_,
		_w8622_,
		_w8623_
	);
	LUT2 #(
		.INIT('h8)
	) name7622 (
		_w8618_,
		_w8622_,
		_w8624_
	);
	LUT2 #(
		.INIT('h1)
	) name7623 (
		_w8575_,
		_w8577_,
		_w8625_
	);
	LUT2 #(
		.INIT('h1)
	) name7624 (
		_w8578_,
		_w8625_,
		_w8626_
	);
	LUT2 #(
		.INIT('h1)
	) name7625 (
		_w8218_,
		_w8220_,
		_w8627_
	);
	LUT2 #(
		.INIT('h1)
	) name7626 (
		_w8221_,
		_w8627_,
		_w8628_
	);
	LUT2 #(
		.INIT('h8)
	) name7627 (
		_w8626_,
		_w8628_,
		_w8629_
	);
	LUT2 #(
		.INIT('h1)
	) name7628 (
		_w8583_,
		_w8584_,
		_w8630_
	);
	LUT2 #(
		.INIT('h4)
	) name7629 (
		_w8588_,
		_w8630_,
		_w8631_
	);
	LUT2 #(
		.INIT('h2)
	) name7630 (
		_w8588_,
		_w8630_,
		_w8632_
	);
	LUT2 #(
		.INIT('h1)
	) name7631 (
		_w8631_,
		_w8632_,
		_w8633_
	);
	LUT2 #(
		.INIT('h8)
	) name7632 (
		_w8629_,
		_w8633_,
		_w8634_
	);
	LUT2 #(
		.INIT('h1)
	) name7633 (
		_w8629_,
		_w8633_,
		_w8635_
	);
	LUT2 #(
		.INIT('h1)
	) name7634 (
		_w8226_,
		_w8227_,
		_w8636_
	);
	LUT2 #(
		.INIT('h4)
	) name7635 (
		_w8231_,
		_w8636_,
		_w8637_
	);
	LUT2 #(
		.INIT('h2)
	) name7636 (
		_w8231_,
		_w8636_,
		_w8638_
	);
	LUT2 #(
		.INIT('h1)
	) name7637 (
		_w8637_,
		_w8638_,
		_w8639_
	);
	LUT2 #(
		.INIT('h4)
	) name7638 (
		_w8635_,
		_w8639_,
		_w8640_
	);
	LUT2 #(
		.INIT('h1)
	) name7639 (
		_w8634_,
		_w8640_,
		_w8641_
	);
	LUT2 #(
		.INIT('h4)
	) name7640 (
		_w8624_,
		_w8641_,
		_w8642_
	);
	LUT2 #(
		.INIT('h1)
	) name7641 (
		_w8623_,
		_w8642_,
		_w8643_
	);
	LUT2 #(
		.INIT('h4)
	) name7642 (
		_w8614_,
		_w8643_,
		_w8644_
	);
	LUT2 #(
		.INIT('h1)
	) name7643 (
		_w8613_,
		_w8644_,
		_w8645_
	);
	LUT2 #(
		.INIT('h1)
	) name7644 (
		_w8604_,
		_w8645_,
		_w8646_
	);
	LUT2 #(
		.INIT('h1)
	) name7645 (
		_w8603_,
		_w8646_,
		_w8647_
	);
	LUT2 #(
		.INIT('h4)
	) name7646 (
		_w8239_,
		_w8242_,
		_w8648_
	);
	LUT2 #(
		.INIT('h1)
	) name7647 (
		_w8238_,
		_w8648_,
		_w8649_
	);
	LUT2 #(
		.INIT('h2)
	) name7648 (
		_w8647_,
		_w8649_,
		_w8650_
	);
	LUT2 #(
		.INIT('h4)
	) name7649 (
		_w8647_,
		_w8649_,
		_w8651_
	);
	LUT2 #(
		.INIT('h4)
	) name7650 (
		_w8596_,
		_w8599_,
		_w8652_
	);
	LUT2 #(
		.INIT('h1)
	) name7651 (
		_w8595_,
		_w8652_,
		_w8653_
	);
	LUT2 #(
		.INIT('h1)
	) name7652 (
		_w8651_,
		_w8653_,
		_w8654_
	);
	LUT2 #(
		.INIT('h1)
	) name7653 (
		_w8650_,
		_w8654_,
		_w8655_
	);
	LUT2 #(
		.INIT('h8)
	) name7654 (
		\A[466] ,
		\A[467] ,
		_w8656_
	);
	LUT2 #(
		.INIT('h1)
	) name7655 (
		\A[466] ,
		\A[467] ,
		_w8657_
	);
	LUT2 #(
		.INIT('h1)
	) name7656 (
		_w8656_,
		_w8657_,
		_w8658_
	);
	LUT2 #(
		.INIT('h8)
	) name7657 (
		\A[468] ,
		_w8658_,
		_w8659_
	);
	LUT2 #(
		.INIT('h1)
	) name7658 (
		\A[468] ,
		_w8658_,
		_w8660_
	);
	LUT2 #(
		.INIT('h1)
	) name7659 (
		_w8659_,
		_w8660_,
		_w8661_
	);
	LUT2 #(
		.INIT('h8)
	) name7660 (
		\A[463] ,
		\A[464] ,
		_w8662_
	);
	LUT2 #(
		.INIT('h1)
	) name7661 (
		\A[463] ,
		\A[464] ,
		_w8663_
	);
	LUT2 #(
		.INIT('h1)
	) name7662 (
		_w8662_,
		_w8663_,
		_w8664_
	);
	LUT2 #(
		.INIT('h8)
	) name7663 (
		\A[465] ,
		_w8664_,
		_w8665_
	);
	LUT2 #(
		.INIT('h1)
	) name7664 (
		\A[465] ,
		_w8664_,
		_w8666_
	);
	LUT2 #(
		.INIT('h1)
	) name7665 (
		_w8665_,
		_w8666_,
		_w8667_
	);
	LUT2 #(
		.INIT('h8)
	) name7666 (
		_w8661_,
		_w8667_,
		_w8668_
	);
	LUT2 #(
		.INIT('h8)
	) name7667 (
		_w8656_,
		_w8668_,
		_w8669_
	);
	LUT2 #(
		.INIT('h1)
	) name7668 (
		_w8662_,
		_w8665_,
		_w8670_
	);
	LUT2 #(
		.INIT('h1)
	) name7669 (
		_w8656_,
		_w8659_,
		_w8671_
	);
	LUT2 #(
		.INIT('h4)
	) name7670 (
		_w8668_,
		_w8671_,
		_w8672_
	);
	LUT2 #(
		.INIT('h1)
	) name7671 (
		_w8670_,
		_w8672_,
		_w8673_
	);
	LUT2 #(
		.INIT('h1)
	) name7672 (
		_w8669_,
		_w8673_,
		_w8674_
	);
	LUT2 #(
		.INIT('h8)
	) name7673 (
		\A[472] ,
		\A[473] ,
		_w8675_
	);
	LUT2 #(
		.INIT('h1)
	) name7674 (
		\A[472] ,
		\A[473] ,
		_w8676_
	);
	LUT2 #(
		.INIT('h1)
	) name7675 (
		_w8675_,
		_w8676_,
		_w8677_
	);
	LUT2 #(
		.INIT('h8)
	) name7676 (
		\A[474] ,
		_w8677_,
		_w8678_
	);
	LUT2 #(
		.INIT('h1)
	) name7677 (
		_w8675_,
		_w8678_,
		_w8679_
	);
	LUT2 #(
		.INIT('h8)
	) name7678 (
		\A[469] ,
		\A[470] ,
		_w8680_
	);
	LUT2 #(
		.INIT('h1)
	) name7679 (
		\A[469] ,
		\A[470] ,
		_w8681_
	);
	LUT2 #(
		.INIT('h1)
	) name7680 (
		_w8680_,
		_w8681_,
		_w8682_
	);
	LUT2 #(
		.INIT('h8)
	) name7681 (
		\A[471] ,
		_w8682_,
		_w8683_
	);
	LUT2 #(
		.INIT('h1)
	) name7682 (
		_w8680_,
		_w8683_,
		_w8684_
	);
	LUT2 #(
		.INIT('h8)
	) name7683 (
		_w8679_,
		_w8684_,
		_w8685_
	);
	LUT2 #(
		.INIT('h1)
	) name7684 (
		_w8679_,
		_w8684_,
		_w8686_
	);
	LUT2 #(
		.INIT('h1)
	) name7685 (
		\A[471] ,
		_w8682_,
		_w8687_
	);
	LUT2 #(
		.INIT('h1)
	) name7686 (
		_w8683_,
		_w8687_,
		_w8688_
	);
	LUT2 #(
		.INIT('h1)
	) name7687 (
		\A[474] ,
		_w8677_,
		_w8689_
	);
	LUT2 #(
		.INIT('h1)
	) name7688 (
		_w8678_,
		_w8689_,
		_w8690_
	);
	LUT2 #(
		.INIT('h8)
	) name7689 (
		_w8688_,
		_w8690_,
		_w8691_
	);
	LUT2 #(
		.INIT('h1)
	) name7690 (
		_w8686_,
		_w8691_,
		_w8692_
	);
	LUT2 #(
		.INIT('h1)
	) name7691 (
		_w8685_,
		_w8692_,
		_w8693_
	);
	LUT2 #(
		.INIT('h1)
	) name7692 (
		_w8688_,
		_w8690_,
		_w8694_
	);
	LUT2 #(
		.INIT('h1)
	) name7693 (
		_w8691_,
		_w8694_,
		_w8695_
	);
	LUT2 #(
		.INIT('h1)
	) name7694 (
		_w8661_,
		_w8667_,
		_w8696_
	);
	LUT2 #(
		.INIT('h1)
	) name7695 (
		_w8668_,
		_w8696_,
		_w8697_
	);
	LUT2 #(
		.INIT('h8)
	) name7696 (
		_w8695_,
		_w8697_,
		_w8698_
	);
	LUT2 #(
		.INIT('h2)
	) name7697 (
		_w8669_,
		_w8670_,
		_w8699_
	);
	LUT2 #(
		.INIT('h2)
	) name7698 (
		_w8698_,
		_w8699_,
		_w8700_
	);
	LUT2 #(
		.INIT('h1)
	) name7699 (
		_w8685_,
		_w8686_,
		_w8701_
	);
	LUT2 #(
		.INIT('h2)
	) name7700 (
		_w8691_,
		_w8701_,
		_w8702_
	);
	LUT2 #(
		.INIT('h4)
	) name7701 (
		_w8691_,
		_w8701_,
		_w8703_
	);
	LUT2 #(
		.INIT('h1)
	) name7702 (
		_w8702_,
		_w8703_,
		_w8704_
	);
	LUT2 #(
		.INIT('h2)
	) name7703 (
		_w8700_,
		_w8704_,
		_w8705_
	);
	LUT2 #(
		.INIT('h4)
	) name7704 (
		_w8700_,
		_w8704_,
		_w8706_
	);
	LUT2 #(
		.INIT('h1)
	) name7705 (
		_w8669_,
		_w8672_,
		_w8707_
	);
	LUT2 #(
		.INIT('h2)
	) name7706 (
		_w8670_,
		_w8707_,
		_w8708_
	);
	LUT2 #(
		.INIT('h4)
	) name7707 (
		_w8670_,
		_w8707_,
		_w8709_
	);
	LUT2 #(
		.INIT('h1)
	) name7708 (
		_w8708_,
		_w8709_,
		_w8710_
	);
	LUT2 #(
		.INIT('h4)
	) name7709 (
		_w8706_,
		_w8710_,
		_w8711_
	);
	LUT2 #(
		.INIT('h1)
	) name7710 (
		_w8705_,
		_w8711_,
		_w8712_
	);
	LUT2 #(
		.INIT('h2)
	) name7711 (
		_w8693_,
		_w8712_,
		_w8713_
	);
	LUT2 #(
		.INIT('h4)
	) name7712 (
		_w8693_,
		_w8712_,
		_w8714_
	);
	LUT2 #(
		.INIT('h1)
	) name7713 (
		_w8713_,
		_w8714_,
		_w8715_
	);
	LUT2 #(
		.INIT('h8)
	) name7714 (
		_w8674_,
		_w8715_,
		_w8716_
	);
	LUT2 #(
		.INIT('h1)
	) name7715 (
		_w8674_,
		_w8715_,
		_w8717_
	);
	LUT2 #(
		.INIT('h1)
	) name7716 (
		_w8716_,
		_w8717_,
		_w8718_
	);
	LUT2 #(
		.INIT('h8)
	) name7717 (
		\A[478] ,
		\A[479] ,
		_w8719_
	);
	LUT2 #(
		.INIT('h8)
	) name7718 (
		\A[475] ,
		\A[476] ,
		_w8720_
	);
	LUT2 #(
		.INIT('h1)
	) name7719 (
		\A[475] ,
		\A[476] ,
		_w8721_
	);
	LUT2 #(
		.INIT('h1)
	) name7720 (
		_w8720_,
		_w8721_,
		_w8722_
	);
	LUT2 #(
		.INIT('h8)
	) name7721 (
		\A[477] ,
		_w8722_,
		_w8723_
	);
	LUT2 #(
		.INIT('h1)
	) name7722 (
		\A[477] ,
		_w8722_,
		_w8724_
	);
	LUT2 #(
		.INIT('h1)
	) name7723 (
		_w8723_,
		_w8724_,
		_w8725_
	);
	LUT2 #(
		.INIT('h1)
	) name7724 (
		\A[478] ,
		\A[479] ,
		_w8726_
	);
	LUT2 #(
		.INIT('h1)
	) name7725 (
		_w8719_,
		_w8726_,
		_w8727_
	);
	LUT2 #(
		.INIT('h8)
	) name7726 (
		\A[480] ,
		_w8727_,
		_w8728_
	);
	LUT2 #(
		.INIT('h1)
	) name7727 (
		\A[480] ,
		_w8727_,
		_w8729_
	);
	LUT2 #(
		.INIT('h1)
	) name7728 (
		_w8728_,
		_w8729_,
		_w8730_
	);
	LUT2 #(
		.INIT('h8)
	) name7729 (
		_w8725_,
		_w8730_,
		_w8731_
	);
	LUT2 #(
		.INIT('h8)
	) name7730 (
		_w8719_,
		_w8731_,
		_w8732_
	);
	LUT2 #(
		.INIT('h1)
	) name7731 (
		_w8720_,
		_w8723_,
		_w8733_
	);
	LUT2 #(
		.INIT('h1)
	) name7732 (
		_w8719_,
		_w8728_,
		_w8734_
	);
	LUT2 #(
		.INIT('h4)
	) name7733 (
		_w8731_,
		_w8734_,
		_w8735_
	);
	LUT2 #(
		.INIT('h1)
	) name7734 (
		_w8733_,
		_w8735_,
		_w8736_
	);
	LUT2 #(
		.INIT('h1)
	) name7735 (
		_w8732_,
		_w8736_,
		_w8737_
	);
	LUT2 #(
		.INIT('h8)
	) name7736 (
		\A[484] ,
		\A[485] ,
		_w8738_
	);
	LUT2 #(
		.INIT('h1)
	) name7737 (
		\A[484] ,
		\A[485] ,
		_w8739_
	);
	LUT2 #(
		.INIT('h1)
	) name7738 (
		_w8738_,
		_w8739_,
		_w8740_
	);
	LUT2 #(
		.INIT('h8)
	) name7739 (
		\A[486] ,
		_w8740_,
		_w8741_
	);
	LUT2 #(
		.INIT('h1)
	) name7740 (
		_w8738_,
		_w8741_,
		_w8742_
	);
	LUT2 #(
		.INIT('h8)
	) name7741 (
		\A[481] ,
		\A[482] ,
		_w8743_
	);
	LUT2 #(
		.INIT('h1)
	) name7742 (
		\A[481] ,
		\A[482] ,
		_w8744_
	);
	LUT2 #(
		.INIT('h1)
	) name7743 (
		_w8743_,
		_w8744_,
		_w8745_
	);
	LUT2 #(
		.INIT('h8)
	) name7744 (
		\A[483] ,
		_w8745_,
		_w8746_
	);
	LUT2 #(
		.INIT('h1)
	) name7745 (
		_w8743_,
		_w8746_,
		_w8747_
	);
	LUT2 #(
		.INIT('h8)
	) name7746 (
		_w8742_,
		_w8747_,
		_w8748_
	);
	LUT2 #(
		.INIT('h1)
	) name7747 (
		_w8742_,
		_w8747_,
		_w8749_
	);
	LUT2 #(
		.INIT('h1)
	) name7748 (
		\A[483] ,
		_w8745_,
		_w8750_
	);
	LUT2 #(
		.INIT('h1)
	) name7749 (
		_w8746_,
		_w8750_,
		_w8751_
	);
	LUT2 #(
		.INIT('h1)
	) name7750 (
		\A[486] ,
		_w8740_,
		_w8752_
	);
	LUT2 #(
		.INIT('h1)
	) name7751 (
		_w8741_,
		_w8752_,
		_w8753_
	);
	LUT2 #(
		.INIT('h8)
	) name7752 (
		_w8751_,
		_w8753_,
		_w8754_
	);
	LUT2 #(
		.INIT('h1)
	) name7753 (
		_w8749_,
		_w8754_,
		_w8755_
	);
	LUT2 #(
		.INIT('h1)
	) name7754 (
		_w8748_,
		_w8755_,
		_w8756_
	);
	LUT2 #(
		.INIT('h1)
	) name7755 (
		_w8751_,
		_w8753_,
		_w8757_
	);
	LUT2 #(
		.INIT('h1)
	) name7756 (
		_w8754_,
		_w8757_,
		_w8758_
	);
	LUT2 #(
		.INIT('h1)
	) name7757 (
		_w8725_,
		_w8730_,
		_w8759_
	);
	LUT2 #(
		.INIT('h1)
	) name7758 (
		_w8731_,
		_w8759_,
		_w8760_
	);
	LUT2 #(
		.INIT('h8)
	) name7759 (
		_w8758_,
		_w8760_,
		_w8761_
	);
	LUT2 #(
		.INIT('h2)
	) name7760 (
		_w8732_,
		_w8733_,
		_w8762_
	);
	LUT2 #(
		.INIT('h2)
	) name7761 (
		_w8761_,
		_w8762_,
		_w8763_
	);
	LUT2 #(
		.INIT('h1)
	) name7762 (
		_w8748_,
		_w8749_,
		_w8764_
	);
	LUT2 #(
		.INIT('h2)
	) name7763 (
		_w8754_,
		_w8764_,
		_w8765_
	);
	LUT2 #(
		.INIT('h4)
	) name7764 (
		_w8754_,
		_w8764_,
		_w8766_
	);
	LUT2 #(
		.INIT('h1)
	) name7765 (
		_w8765_,
		_w8766_,
		_w8767_
	);
	LUT2 #(
		.INIT('h2)
	) name7766 (
		_w8763_,
		_w8767_,
		_w8768_
	);
	LUT2 #(
		.INIT('h4)
	) name7767 (
		_w8763_,
		_w8767_,
		_w8769_
	);
	LUT2 #(
		.INIT('h1)
	) name7768 (
		_w8732_,
		_w8735_,
		_w8770_
	);
	LUT2 #(
		.INIT('h2)
	) name7769 (
		_w8733_,
		_w8770_,
		_w8771_
	);
	LUT2 #(
		.INIT('h4)
	) name7770 (
		_w8733_,
		_w8770_,
		_w8772_
	);
	LUT2 #(
		.INIT('h1)
	) name7771 (
		_w8771_,
		_w8772_,
		_w8773_
	);
	LUT2 #(
		.INIT('h4)
	) name7772 (
		_w8769_,
		_w8773_,
		_w8774_
	);
	LUT2 #(
		.INIT('h1)
	) name7773 (
		_w8768_,
		_w8774_,
		_w8775_
	);
	LUT2 #(
		.INIT('h2)
	) name7774 (
		_w8756_,
		_w8775_,
		_w8776_
	);
	LUT2 #(
		.INIT('h4)
	) name7775 (
		_w8756_,
		_w8775_,
		_w8777_
	);
	LUT2 #(
		.INIT('h1)
	) name7776 (
		_w8776_,
		_w8777_,
		_w8778_
	);
	LUT2 #(
		.INIT('h8)
	) name7777 (
		_w8737_,
		_w8778_,
		_w8779_
	);
	LUT2 #(
		.INIT('h1)
	) name7778 (
		_w8737_,
		_w8778_,
		_w8780_
	);
	LUT2 #(
		.INIT('h1)
	) name7779 (
		_w8779_,
		_w8780_,
		_w8781_
	);
	LUT2 #(
		.INIT('h1)
	) name7780 (
		_w8718_,
		_w8781_,
		_w8782_
	);
	LUT2 #(
		.INIT('h8)
	) name7781 (
		_w8718_,
		_w8781_,
		_w8783_
	);
	LUT2 #(
		.INIT('h1)
	) name7782 (
		_w8695_,
		_w8697_,
		_w8784_
	);
	LUT2 #(
		.INIT('h1)
	) name7783 (
		_w8698_,
		_w8784_,
		_w8785_
	);
	LUT2 #(
		.INIT('h1)
	) name7784 (
		_w8758_,
		_w8760_,
		_w8786_
	);
	LUT2 #(
		.INIT('h1)
	) name7785 (
		_w8761_,
		_w8786_,
		_w8787_
	);
	LUT2 #(
		.INIT('h8)
	) name7786 (
		_w8785_,
		_w8787_,
		_w8788_
	);
	LUT2 #(
		.INIT('h1)
	) name7787 (
		_w8768_,
		_w8769_,
		_w8789_
	);
	LUT2 #(
		.INIT('h8)
	) name7788 (
		_w8773_,
		_w8789_,
		_w8790_
	);
	LUT2 #(
		.INIT('h1)
	) name7789 (
		_w8773_,
		_w8789_,
		_w8791_
	);
	LUT2 #(
		.INIT('h1)
	) name7790 (
		_w8790_,
		_w8791_,
		_w8792_
	);
	LUT2 #(
		.INIT('h8)
	) name7791 (
		_w8788_,
		_w8792_,
		_w8793_
	);
	LUT2 #(
		.INIT('h1)
	) name7792 (
		_w8788_,
		_w8792_,
		_w8794_
	);
	LUT2 #(
		.INIT('h1)
	) name7793 (
		_w8705_,
		_w8706_,
		_w8795_
	);
	LUT2 #(
		.INIT('h8)
	) name7794 (
		_w8710_,
		_w8795_,
		_w8796_
	);
	LUT2 #(
		.INIT('h1)
	) name7795 (
		_w8710_,
		_w8795_,
		_w8797_
	);
	LUT2 #(
		.INIT('h1)
	) name7796 (
		_w8796_,
		_w8797_,
		_w8798_
	);
	LUT2 #(
		.INIT('h4)
	) name7797 (
		_w8794_,
		_w8798_,
		_w8799_
	);
	LUT2 #(
		.INIT('h1)
	) name7798 (
		_w8793_,
		_w8799_,
		_w8800_
	);
	LUT2 #(
		.INIT('h1)
	) name7799 (
		_w8783_,
		_w8800_,
		_w8801_
	);
	LUT2 #(
		.INIT('h1)
	) name7800 (
		_w8782_,
		_w8801_,
		_w8802_
	);
	LUT2 #(
		.INIT('h1)
	) name7801 (
		_w8737_,
		_w8777_,
		_w8803_
	);
	LUT2 #(
		.INIT('h1)
	) name7802 (
		_w8776_,
		_w8803_,
		_w8804_
	);
	LUT2 #(
		.INIT('h1)
	) name7803 (
		_w8802_,
		_w8804_,
		_w8805_
	);
	LUT2 #(
		.INIT('h8)
	) name7804 (
		_w8802_,
		_w8804_,
		_w8806_
	);
	LUT2 #(
		.INIT('h1)
	) name7805 (
		_w8674_,
		_w8714_,
		_w8807_
	);
	LUT2 #(
		.INIT('h1)
	) name7806 (
		_w8713_,
		_w8807_,
		_w8808_
	);
	LUT2 #(
		.INIT('h1)
	) name7807 (
		_w8806_,
		_w8808_,
		_w8809_
	);
	LUT2 #(
		.INIT('h1)
	) name7808 (
		_w8805_,
		_w8809_,
		_w8810_
	);
	LUT2 #(
		.INIT('h8)
	) name7809 (
		\A[490] ,
		\A[491] ,
		_w8811_
	);
	LUT2 #(
		.INIT('h8)
	) name7810 (
		\A[487] ,
		\A[488] ,
		_w8812_
	);
	LUT2 #(
		.INIT('h1)
	) name7811 (
		\A[487] ,
		\A[488] ,
		_w8813_
	);
	LUT2 #(
		.INIT('h1)
	) name7812 (
		_w8812_,
		_w8813_,
		_w8814_
	);
	LUT2 #(
		.INIT('h8)
	) name7813 (
		\A[489] ,
		_w8814_,
		_w8815_
	);
	LUT2 #(
		.INIT('h1)
	) name7814 (
		\A[489] ,
		_w8814_,
		_w8816_
	);
	LUT2 #(
		.INIT('h1)
	) name7815 (
		_w8815_,
		_w8816_,
		_w8817_
	);
	LUT2 #(
		.INIT('h1)
	) name7816 (
		\A[490] ,
		\A[491] ,
		_w8818_
	);
	LUT2 #(
		.INIT('h1)
	) name7817 (
		_w8811_,
		_w8818_,
		_w8819_
	);
	LUT2 #(
		.INIT('h8)
	) name7818 (
		\A[492] ,
		_w8819_,
		_w8820_
	);
	LUT2 #(
		.INIT('h1)
	) name7819 (
		\A[492] ,
		_w8819_,
		_w8821_
	);
	LUT2 #(
		.INIT('h1)
	) name7820 (
		_w8820_,
		_w8821_,
		_w8822_
	);
	LUT2 #(
		.INIT('h8)
	) name7821 (
		_w8817_,
		_w8822_,
		_w8823_
	);
	LUT2 #(
		.INIT('h8)
	) name7822 (
		_w8811_,
		_w8823_,
		_w8824_
	);
	LUT2 #(
		.INIT('h1)
	) name7823 (
		_w8812_,
		_w8815_,
		_w8825_
	);
	LUT2 #(
		.INIT('h1)
	) name7824 (
		_w8811_,
		_w8820_,
		_w8826_
	);
	LUT2 #(
		.INIT('h4)
	) name7825 (
		_w8823_,
		_w8826_,
		_w8827_
	);
	LUT2 #(
		.INIT('h1)
	) name7826 (
		_w8825_,
		_w8827_,
		_w8828_
	);
	LUT2 #(
		.INIT('h1)
	) name7827 (
		_w8824_,
		_w8828_,
		_w8829_
	);
	LUT2 #(
		.INIT('h8)
	) name7828 (
		\A[496] ,
		\A[497] ,
		_w8830_
	);
	LUT2 #(
		.INIT('h1)
	) name7829 (
		\A[496] ,
		\A[497] ,
		_w8831_
	);
	LUT2 #(
		.INIT('h1)
	) name7830 (
		_w8830_,
		_w8831_,
		_w8832_
	);
	LUT2 #(
		.INIT('h8)
	) name7831 (
		\A[498] ,
		_w8832_,
		_w8833_
	);
	LUT2 #(
		.INIT('h1)
	) name7832 (
		_w8830_,
		_w8833_,
		_w8834_
	);
	LUT2 #(
		.INIT('h8)
	) name7833 (
		\A[493] ,
		\A[494] ,
		_w8835_
	);
	LUT2 #(
		.INIT('h1)
	) name7834 (
		\A[493] ,
		\A[494] ,
		_w8836_
	);
	LUT2 #(
		.INIT('h1)
	) name7835 (
		_w8835_,
		_w8836_,
		_w8837_
	);
	LUT2 #(
		.INIT('h8)
	) name7836 (
		\A[495] ,
		_w8837_,
		_w8838_
	);
	LUT2 #(
		.INIT('h1)
	) name7837 (
		_w8835_,
		_w8838_,
		_w8839_
	);
	LUT2 #(
		.INIT('h8)
	) name7838 (
		_w8834_,
		_w8839_,
		_w8840_
	);
	LUT2 #(
		.INIT('h1)
	) name7839 (
		_w8834_,
		_w8839_,
		_w8841_
	);
	LUT2 #(
		.INIT('h1)
	) name7840 (
		\A[495] ,
		_w8837_,
		_w8842_
	);
	LUT2 #(
		.INIT('h1)
	) name7841 (
		_w8838_,
		_w8842_,
		_w8843_
	);
	LUT2 #(
		.INIT('h1)
	) name7842 (
		\A[498] ,
		_w8832_,
		_w8844_
	);
	LUT2 #(
		.INIT('h1)
	) name7843 (
		_w8833_,
		_w8844_,
		_w8845_
	);
	LUT2 #(
		.INIT('h8)
	) name7844 (
		_w8843_,
		_w8845_,
		_w8846_
	);
	LUT2 #(
		.INIT('h1)
	) name7845 (
		_w8841_,
		_w8846_,
		_w8847_
	);
	LUT2 #(
		.INIT('h1)
	) name7846 (
		_w8840_,
		_w8847_,
		_w8848_
	);
	LUT2 #(
		.INIT('h1)
	) name7847 (
		_w8843_,
		_w8845_,
		_w8849_
	);
	LUT2 #(
		.INIT('h1)
	) name7848 (
		_w8846_,
		_w8849_,
		_w8850_
	);
	LUT2 #(
		.INIT('h1)
	) name7849 (
		_w8817_,
		_w8822_,
		_w8851_
	);
	LUT2 #(
		.INIT('h1)
	) name7850 (
		_w8823_,
		_w8851_,
		_w8852_
	);
	LUT2 #(
		.INIT('h8)
	) name7851 (
		_w8850_,
		_w8852_,
		_w8853_
	);
	LUT2 #(
		.INIT('h2)
	) name7852 (
		_w8824_,
		_w8825_,
		_w8854_
	);
	LUT2 #(
		.INIT('h2)
	) name7853 (
		_w8853_,
		_w8854_,
		_w8855_
	);
	LUT2 #(
		.INIT('h1)
	) name7854 (
		_w8840_,
		_w8841_,
		_w8856_
	);
	LUT2 #(
		.INIT('h2)
	) name7855 (
		_w8846_,
		_w8856_,
		_w8857_
	);
	LUT2 #(
		.INIT('h4)
	) name7856 (
		_w8846_,
		_w8856_,
		_w8858_
	);
	LUT2 #(
		.INIT('h1)
	) name7857 (
		_w8857_,
		_w8858_,
		_w8859_
	);
	LUT2 #(
		.INIT('h2)
	) name7858 (
		_w8855_,
		_w8859_,
		_w8860_
	);
	LUT2 #(
		.INIT('h4)
	) name7859 (
		_w8855_,
		_w8859_,
		_w8861_
	);
	LUT2 #(
		.INIT('h1)
	) name7860 (
		_w8824_,
		_w8827_,
		_w8862_
	);
	LUT2 #(
		.INIT('h2)
	) name7861 (
		_w8825_,
		_w8862_,
		_w8863_
	);
	LUT2 #(
		.INIT('h4)
	) name7862 (
		_w8825_,
		_w8862_,
		_w8864_
	);
	LUT2 #(
		.INIT('h1)
	) name7863 (
		_w8863_,
		_w8864_,
		_w8865_
	);
	LUT2 #(
		.INIT('h4)
	) name7864 (
		_w8861_,
		_w8865_,
		_w8866_
	);
	LUT2 #(
		.INIT('h1)
	) name7865 (
		_w8860_,
		_w8866_,
		_w8867_
	);
	LUT2 #(
		.INIT('h2)
	) name7866 (
		_w8848_,
		_w8867_,
		_w8868_
	);
	LUT2 #(
		.INIT('h4)
	) name7867 (
		_w8848_,
		_w8867_,
		_w8869_
	);
	LUT2 #(
		.INIT('h1)
	) name7868 (
		_w8868_,
		_w8869_,
		_w8870_
	);
	LUT2 #(
		.INIT('h8)
	) name7869 (
		_w8829_,
		_w8870_,
		_w8871_
	);
	LUT2 #(
		.INIT('h1)
	) name7870 (
		_w8829_,
		_w8870_,
		_w8872_
	);
	LUT2 #(
		.INIT('h1)
	) name7871 (
		_w8871_,
		_w8872_,
		_w8873_
	);
	LUT2 #(
		.INIT('h8)
	) name7872 (
		\A[502] ,
		\A[503] ,
		_w8874_
	);
	LUT2 #(
		.INIT('h8)
	) name7873 (
		\A[499] ,
		\A[500] ,
		_w8875_
	);
	LUT2 #(
		.INIT('h1)
	) name7874 (
		\A[499] ,
		\A[500] ,
		_w8876_
	);
	LUT2 #(
		.INIT('h1)
	) name7875 (
		_w8875_,
		_w8876_,
		_w8877_
	);
	LUT2 #(
		.INIT('h8)
	) name7876 (
		\A[501] ,
		_w8877_,
		_w8878_
	);
	LUT2 #(
		.INIT('h1)
	) name7877 (
		\A[501] ,
		_w8877_,
		_w8879_
	);
	LUT2 #(
		.INIT('h1)
	) name7878 (
		_w8878_,
		_w8879_,
		_w8880_
	);
	LUT2 #(
		.INIT('h1)
	) name7879 (
		\A[502] ,
		\A[503] ,
		_w8881_
	);
	LUT2 #(
		.INIT('h1)
	) name7880 (
		_w8874_,
		_w8881_,
		_w8882_
	);
	LUT2 #(
		.INIT('h8)
	) name7881 (
		\A[504] ,
		_w8882_,
		_w8883_
	);
	LUT2 #(
		.INIT('h1)
	) name7882 (
		\A[504] ,
		_w8882_,
		_w8884_
	);
	LUT2 #(
		.INIT('h1)
	) name7883 (
		_w8883_,
		_w8884_,
		_w8885_
	);
	LUT2 #(
		.INIT('h8)
	) name7884 (
		_w8880_,
		_w8885_,
		_w8886_
	);
	LUT2 #(
		.INIT('h8)
	) name7885 (
		_w8874_,
		_w8886_,
		_w8887_
	);
	LUT2 #(
		.INIT('h1)
	) name7886 (
		_w8875_,
		_w8878_,
		_w8888_
	);
	LUT2 #(
		.INIT('h1)
	) name7887 (
		_w8874_,
		_w8883_,
		_w8889_
	);
	LUT2 #(
		.INIT('h4)
	) name7888 (
		_w8886_,
		_w8889_,
		_w8890_
	);
	LUT2 #(
		.INIT('h1)
	) name7889 (
		_w8888_,
		_w8890_,
		_w8891_
	);
	LUT2 #(
		.INIT('h1)
	) name7890 (
		_w8887_,
		_w8891_,
		_w8892_
	);
	LUT2 #(
		.INIT('h8)
	) name7891 (
		\A[508] ,
		\A[509] ,
		_w8893_
	);
	LUT2 #(
		.INIT('h1)
	) name7892 (
		\A[508] ,
		\A[509] ,
		_w8894_
	);
	LUT2 #(
		.INIT('h1)
	) name7893 (
		_w8893_,
		_w8894_,
		_w8895_
	);
	LUT2 #(
		.INIT('h8)
	) name7894 (
		\A[510] ,
		_w8895_,
		_w8896_
	);
	LUT2 #(
		.INIT('h1)
	) name7895 (
		_w8893_,
		_w8896_,
		_w8897_
	);
	LUT2 #(
		.INIT('h8)
	) name7896 (
		\A[505] ,
		\A[506] ,
		_w8898_
	);
	LUT2 #(
		.INIT('h1)
	) name7897 (
		\A[505] ,
		\A[506] ,
		_w8899_
	);
	LUT2 #(
		.INIT('h1)
	) name7898 (
		_w8898_,
		_w8899_,
		_w8900_
	);
	LUT2 #(
		.INIT('h8)
	) name7899 (
		\A[507] ,
		_w8900_,
		_w8901_
	);
	LUT2 #(
		.INIT('h1)
	) name7900 (
		_w8898_,
		_w8901_,
		_w8902_
	);
	LUT2 #(
		.INIT('h8)
	) name7901 (
		_w8897_,
		_w8902_,
		_w8903_
	);
	LUT2 #(
		.INIT('h1)
	) name7902 (
		_w8897_,
		_w8902_,
		_w8904_
	);
	LUT2 #(
		.INIT('h1)
	) name7903 (
		\A[507] ,
		_w8900_,
		_w8905_
	);
	LUT2 #(
		.INIT('h1)
	) name7904 (
		_w8901_,
		_w8905_,
		_w8906_
	);
	LUT2 #(
		.INIT('h1)
	) name7905 (
		\A[510] ,
		_w8895_,
		_w8907_
	);
	LUT2 #(
		.INIT('h1)
	) name7906 (
		_w8896_,
		_w8907_,
		_w8908_
	);
	LUT2 #(
		.INIT('h8)
	) name7907 (
		_w8906_,
		_w8908_,
		_w8909_
	);
	LUT2 #(
		.INIT('h1)
	) name7908 (
		_w8904_,
		_w8909_,
		_w8910_
	);
	LUT2 #(
		.INIT('h1)
	) name7909 (
		_w8903_,
		_w8910_,
		_w8911_
	);
	LUT2 #(
		.INIT('h1)
	) name7910 (
		_w8906_,
		_w8908_,
		_w8912_
	);
	LUT2 #(
		.INIT('h1)
	) name7911 (
		_w8909_,
		_w8912_,
		_w8913_
	);
	LUT2 #(
		.INIT('h1)
	) name7912 (
		_w8880_,
		_w8885_,
		_w8914_
	);
	LUT2 #(
		.INIT('h1)
	) name7913 (
		_w8886_,
		_w8914_,
		_w8915_
	);
	LUT2 #(
		.INIT('h8)
	) name7914 (
		_w8913_,
		_w8915_,
		_w8916_
	);
	LUT2 #(
		.INIT('h2)
	) name7915 (
		_w8887_,
		_w8888_,
		_w8917_
	);
	LUT2 #(
		.INIT('h2)
	) name7916 (
		_w8916_,
		_w8917_,
		_w8918_
	);
	LUT2 #(
		.INIT('h1)
	) name7917 (
		_w8903_,
		_w8904_,
		_w8919_
	);
	LUT2 #(
		.INIT('h2)
	) name7918 (
		_w8909_,
		_w8919_,
		_w8920_
	);
	LUT2 #(
		.INIT('h4)
	) name7919 (
		_w8909_,
		_w8919_,
		_w8921_
	);
	LUT2 #(
		.INIT('h1)
	) name7920 (
		_w8920_,
		_w8921_,
		_w8922_
	);
	LUT2 #(
		.INIT('h2)
	) name7921 (
		_w8918_,
		_w8922_,
		_w8923_
	);
	LUT2 #(
		.INIT('h4)
	) name7922 (
		_w8918_,
		_w8922_,
		_w8924_
	);
	LUT2 #(
		.INIT('h1)
	) name7923 (
		_w8887_,
		_w8890_,
		_w8925_
	);
	LUT2 #(
		.INIT('h2)
	) name7924 (
		_w8888_,
		_w8925_,
		_w8926_
	);
	LUT2 #(
		.INIT('h4)
	) name7925 (
		_w8888_,
		_w8925_,
		_w8927_
	);
	LUT2 #(
		.INIT('h1)
	) name7926 (
		_w8926_,
		_w8927_,
		_w8928_
	);
	LUT2 #(
		.INIT('h4)
	) name7927 (
		_w8924_,
		_w8928_,
		_w8929_
	);
	LUT2 #(
		.INIT('h1)
	) name7928 (
		_w8923_,
		_w8929_,
		_w8930_
	);
	LUT2 #(
		.INIT('h2)
	) name7929 (
		_w8911_,
		_w8930_,
		_w8931_
	);
	LUT2 #(
		.INIT('h4)
	) name7930 (
		_w8911_,
		_w8930_,
		_w8932_
	);
	LUT2 #(
		.INIT('h1)
	) name7931 (
		_w8931_,
		_w8932_,
		_w8933_
	);
	LUT2 #(
		.INIT('h8)
	) name7932 (
		_w8892_,
		_w8933_,
		_w8934_
	);
	LUT2 #(
		.INIT('h1)
	) name7933 (
		_w8892_,
		_w8933_,
		_w8935_
	);
	LUT2 #(
		.INIT('h1)
	) name7934 (
		_w8934_,
		_w8935_,
		_w8936_
	);
	LUT2 #(
		.INIT('h1)
	) name7935 (
		_w8873_,
		_w8936_,
		_w8937_
	);
	LUT2 #(
		.INIT('h8)
	) name7936 (
		_w8873_,
		_w8936_,
		_w8938_
	);
	LUT2 #(
		.INIT('h1)
	) name7937 (
		_w8913_,
		_w8915_,
		_w8939_
	);
	LUT2 #(
		.INIT('h1)
	) name7938 (
		_w8916_,
		_w8939_,
		_w8940_
	);
	LUT2 #(
		.INIT('h1)
	) name7939 (
		_w8850_,
		_w8852_,
		_w8941_
	);
	LUT2 #(
		.INIT('h1)
	) name7940 (
		_w8853_,
		_w8941_,
		_w8942_
	);
	LUT2 #(
		.INIT('h8)
	) name7941 (
		_w8940_,
		_w8942_,
		_w8943_
	);
	LUT2 #(
		.INIT('h1)
	) name7942 (
		_w8923_,
		_w8924_,
		_w8944_
	);
	LUT2 #(
		.INIT('h8)
	) name7943 (
		_w8928_,
		_w8944_,
		_w8945_
	);
	LUT2 #(
		.INIT('h1)
	) name7944 (
		_w8928_,
		_w8944_,
		_w8946_
	);
	LUT2 #(
		.INIT('h1)
	) name7945 (
		_w8945_,
		_w8946_,
		_w8947_
	);
	LUT2 #(
		.INIT('h8)
	) name7946 (
		_w8943_,
		_w8947_,
		_w8948_
	);
	LUT2 #(
		.INIT('h1)
	) name7947 (
		_w8943_,
		_w8947_,
		_w8949_
	);
	LUT2 #(
		.INIT('h1)
	) name7948 (
		_w8860_,
		_w8861_,
		_w8950_
	);
	LUT2 #(
		.INIT('h8)
	) name7949 (
		_w8865_,
		_w8950_,
		_w8951_
	);
	LUT2 #(
		.INIT('h1)
	) name7950 (
		_w8865_,
		_w8950_,
		_w8952_
	);
	LUT2 #(
		.INIT('h1)
	) name7951 (
		_w8951_,
		_w8952_,
		_w8953_
	);
	LUT2 #(
		.INIT('h4)
	) name7952 (
		_w8949_,
		_w8953_,
		_w8954_
	);
	LUT2 #(
		.INIT('h1)
	) name7953 (
		_w8948_,
		_w8954_,
		_w8955_
	);
	LUT2 #(
		.INIT('h1)
	) name7954 (
		_w8938_,
		_w8955_,
		_w8956_
	);
	LUT2 #(
		.INIT('h1)
	) name7955 (
		_w8937_,
		_w8956_,
		_w8957_
	);
	LUT2 #(
		.INIT('h1)
	) name7956 (
		_w8892_,
		_w8932_,
		_w8958_
	);
	LUT2 #(
		.INIT('h1)
	) name7957 (
		_w8931_,
		_w8958_,
		_w8959_
	);
	LUT2 #(
		.INIT('h1)
	) name7958 (
		_w8957_,
		_w8959_,
		_w8960_
	);
	LUT2 #(
		.INIT('h8)
	) name7959 (
		_w8957_,
		_w8959_,
		_w8961_
	);
	LUT2 #(
		.INIT('h1)
	) name7960 (
		_w8960_,
		_w8961_,
		_w8962_
	);
	LUT2 #(
		.INIT('h1)
	) name7961 (
		_w8829_,
		_w8869_,
		_w8963_
	);
	LUT2 #(
		.INIT('h1)
	) name7962 (
		_w8868_,
		_w8963_,
		_w8964_
	);
	LUT2 #(
		.INIT('h2)
	) name7963 (
		_w8962_,
		_w8964_,
		_w8965_
	);
	LUT2 #(
		.INIT('h4)
	) name7964 (
		_w8962_,
		_w8964_,
		_w8966_
	);
	LUT2 #(
		.INIT('h1)
	) name7965 (
		_w8965_,
		_w8966_,
		_w8967_
	);
	LUT2 #(
		.INIT('h1)
	) name7966 (
		_w8805_,
		_w8806_,
		_w8968_
	);
	LUT2 #(
		.INIT('h4)
	) name7967 (
		_w8808_,
		_w8968_,
		_w8969_
	);
	LUT2 #(
		.INIT('h2)
	) name7968 (
		_w8808_,
		_w8968_,
		_w8970_
	);
	LUT2 #(
		.INIT('h1)
	) name7969 (
		_w8969_,
		_w8970_,
		_w8971_
	);
	LUT2 #(
		.INIT('h1)
	) name7970 (
		_w8967_,
		_w8971_,
		_w8972_
	);
	LUT2 #(
		.INIT('h8)
	) name7971 (
		_w8967_,
		_w8971_,
		_w8973_
	);
	LUT2 #(
		.INIT('h1)
	) name7972 (
		_w8782_,
		_w8783_,
		_w8974_
	);
	LUT2 #(
		.INIT('h4)
	) name7973 (
		_w8800_,
		_w8974_,
		_w8975_
	);
	LUT2 #(
		.INIT('h2)
	) name7974 (
		_w8800_,
		_w8974_,
		_w8976_
	);
	LUT2 #(
		.INIT('h1)
	) name7975 (
		_w8975_,
		_w8976_,
		_w8977_
	);
	LUT2 #(
		.INIT('h1)
	) name7976 (
		_w8937_,
		_w8938_,
		_w8978_
	);
	LUT2 #(
		.INIT('h4)
	) name7977 (
		_w8955_,
		_w8978_,
		_w8979_
	);
	LUT2 #(
		.INIT('h2)
	) name7978 (
		_w8955_,
		_w8978_,
		_w8980_
	);
	LUT2 #(
		.INIT('h1)
	) name7979 (
		_w8979_,
		_w8980_,
		_w8981_
	);
	LUT2 #(
		.INIT('h1)
	) name7980 (
		_w8977_,
		_w8981_,
		_w8982_
	);
	LUT2 #(
		.INIT('h8)
	) name7981 (
		_w8977_,
		_w8981_,
		_w8983_
	);
	LUT2 #(
		.INIT('h1)
	) name7982 (
		_w8785_,
		_w8787_,
		_w8984_
	);
	LUT2 #(
		.INIT('h1)
	) name7983 (
		_w8788_,
		_w8984_,
		_w8985_
	);
	LUT2 #(
		.INIT('h1)
	) name7984 (
		_w8940_,
		_w8942_,
		_w8986_
	);
	LUT2 #(
		.INIT('h1)
	) name7985 (
		_w8943_,
		_w8986_,
		_w8987_
	);
	LUT2 #(
		.INIT('h8)
	) name7986 (
		_w8985_,
		_w8987_,
		_w8988_
	);
	LUT2 #(
		.INIT('h1)
	) name7987 (
		_w8948_,
		_w8949_,
		_w8989_
	);
	LUT2 #(
		.INIT('h4)
	) name7988 (
		_w8953_,
		_w8989_,
		_w8990_
	);
	LUT2 #(
		.INIT('h2)
	) name7989 (
		_w8953_,
		_w8989_,
		_w8991_
	);
	LUT2 #(
		.INIT('h1)
	) name7990 (
		_w8990_,
		_w8991_,
		_w8992_
	);
	LUT2 #(
		.INIT('h2)
	) name7991 (
		_w8988_,
		_w8992_,
		_w8993_
	);
	LUT2 #(
		.INIT('h4)
	) name7992 (
		_w8988_,
		_w8992_,
		_w8994_
	);
	LUT2 #(
		.INIT('h1)
	) name7993 (
		_w8793_,
		_w8794_,
		_w8995_
	);
	LUT2 #(
		.INIT('h4)
	) name7994 (
		_w8798_,
		_w8995_,
		_w8996_
	);
	LUT2 #(
		.INIT('h2)
	) name7995 (
		_w8798_,
		_w8995_,
		_w8997_
	);
	LUT2 #(
		.INIT('h1)
	) name7996 (
		_w8996_,
		_w8997_,
		_w8998_
	);
	LUT2 #(
		.INIT('h1)
	) name7997 (
		_w8994_,
		_w8998_,
		_w8999_
	);
	LUT2 #(
		.INIT('h1)
	) name7998 (
		_w8993_,
		_w8999_,
		_w9000_
	);
	LUT2 #(
		.INIT('h4)
	) name7999 (
		_w8983_,
		_w9000_,
		_w9001_
	);
	LUT2 #(
		.INIT('h1)
	) name8000 (
		_w8982_,
		_w9001_,
		_w9002_
	);
	LUT2 #(
		.INIT('h1)
	) name8001 (
		_w8973_,
		_w9002_,
		_w9003_
	);
	LUT2 #(
		.INIT('h1)
	) name8002 (
		_w8972_,
		_w9003_,
		_w9004_
	);
	LUT2 #(
		.INIT('h2)
	) name8003 (
		_w8810_,
		_w9004_,
		_w9005_
	);
	LUT2 #(
		.INIT('h4)
	) name8004 (
		_w8810_,
		_w9004_,
		_w9006_
	);
	LUT2 #(
		.INIT('h1)
	) name8005 (
		_w9005_,
		_w9006_,
		_w9007_
	);
	LUT2 #(
		.INIT('h1)
	) name8006 (
		_w8961_,
		_w8964_,
		_w9008_
	);
	LUT2 #(
		.INIT('h1)
	) name8007 (
		_w8960_,
		_w9008_,
		_w9009_
	);
	LUT2 #(
		.INIT('h8)
	) name8008 (
		_w9007_,
		_w9009_,
		_w9010_
	);
	LUT2 #(
		.INIT('h1)
	) name8009 (
		_w9007_,
		_w9009_,
		_w9011_
	);
	LUT2 #(
		.INIT('h1)
	) name8010 (
		_w9010_,
		_w9011_,
		_w9012_
	);
	LUT2 #(
		.INIT('h8)
	) name8011 (
		\A[538] ,
		\A[539] ,
		_w9013_
	);
	LUT2 #(
		.INIT('h8)
	) name8012 (
		\A[535] ,
		\A[536] ,
		_w9014_
	);
	LUT2 #(
		.INIT('h1)
	) name8013 (
		\A[535] ,
		\A[536] ,
		_w9015_
	);
	LUT2 #(
		.INIT('h1)
	) name8014 (
		_w9014_,
		_w9015_,
		_w9016_
	);
	LUT2 #(
		.INIT('h8)
	) name8015 (
		\A[537] ,
		_w9016_,
		_w9017_
	);
	LUT2 #(
		.INIT('h1)
	) name8016 (
		\A[537] ,
		_w9016_,
		_w9018_
	);
	LUT2 #(
		.INIT('h1)
	) name8017 (
		_w9017_,
		_w9018_,
		_w9019_
	);
	LUT2 #(
		.INIT('h1)
	) name8018 (
		\A[538] ,
		\A[539] ,
		_w9020_
	);
	LUT2 #(
		.INIT('h1)
	) name8019 (
		_w9013_,
		_w9020_,
		_w9021_
	);
	LUT2 #(
		.INIT('h8)
	) name8020 (
		\A[540] ,
		_w9021_,
		_w9022_
	);
	LUT2 #(
		.INIT('h1)
	) name8021 (
		\A[540] ,
		_w9021_,
		_w9023_
	);
	LUT2 #(
		.INIT('h1)
	) name8022 (
		_w9022_,
		_w9023_,
		_w9024_
	);
	LUT2 #(
		.INIT('h8)
	) name8023 (
		_w9019_,
		_w9024_,
		_w9025_
	);
	LUT2 #(
		.INIT('h8)
	) name8024 (
		_w9013_,
		_w9025_,
		_w9026_
	);
	LUT2 #(
		.INIT('h1)
	) name8025 (
		_w9014_,
		_w9017_,
		_w9027_
	);
	LUT2 #(
		.INIT('h1)
	) name8026 (
		_w9013_,
		_w9022_,
		_w9028_
	);
	LUT2 #(
		.INIT('h4)
	) name8027 (
		_w9025_,
		_w9028_,
		_w9029_
	);
	LUT2 #(
		.INIT('h1)
	) name8028 (
		_w9027_,
		_w9029_,
		_w9030_
	);
	LUT2 #(
		.INIT('h1)
	) name8029 (
		_w9026_,
		_w9030_,
		_w9031_
	);
	LUT2 #(
		.INIT('h8)
	) name8030 (
		\A[544] ,
		\A[545] ,
		_w9032_
	);
	LUT2 #(
		.INIT('h1)
	) name8031 (
		\A[544] ,
		\A[545] ,
		_w9033_
	);
	LUT2 #(
		.INIT('h1)
	) name8032 (
		_w9032_,
		_w9033_,
		_w9034_
	);
	LUT2 #(
		.INIT('h8)
	) name8033 (
		\A[546] ,
		_w9034_,
		_w9035_
	);
	LUT2 #(
		.INIT('h1)
	) name8034 (
		_w9032_,
		_w9035_,
		_w9036_
	);
	LUT2 #(
		.INIT('h8)
	) name8035 (
		\A[541] ,
		\A[542] ,
		_w9037_
	);
	LUT2 #(
		.INIT('h1)
	) name8036 (
		\A[541] ,
		\A[542] ,
		_w9038_
	);
	LUT2 #(
		.INIT('h1)
	) name8037 (
		_w9037_,
		_w9038_,
		_w9039_
	);
	LUT2 #(
		.INIT('h8)
	) name8038 (
		\A[543] ,
		_w9039_,
		_w9040_
	);
	LUT2 #(
		.INIT('h1)
	) name8039 (
		_w9037_,
		_w9040_,
		_w9041_
	);
	LUT2 #(
		.INIT('h8)
	) name8040 (
		_w9036_,
		_w9041_,
		_w9042_
	);
	LUT2 #(
		.INIT('h1)
	) name8041 (
		_w9036_,
		_w9041_,
		_w9043_
	);
	LUT2 #(
		.INIT('h1)
	) name8042 (
		\A[543] ,
		_w9039_,
		_w9044_
	);
	LUT2 #(
		.INIT('h1)
	) name8043 (
		_w9040_,
		_w9044_,
		_w9045_
	);
	LUT2 #(
		.INIT('h1)
	) name8044 (
		\A[546] ,
		_w9034_,
		_w9046_
	);
	LUT2 #(
		.INIT('h1)
	) name8045 (
		_w9035_,
		_w9046_,
		_w9047_
	);
	LUT2 #(
		.INIT('h8)
	) name8046 (
		_w9045_,
		_w9047_,
		_w9048_
	);
	LUT2 #(
		.INIT('h1)
	) name8047 (
		_w9043_,
		_w9048_,
		_w9049_
	);
	LUT2 #(
		.INIT('h1)
	) name8048 (
		_w9042_,
		_w9049_,
		_w9050_
	);
	LUT2 #(
		.INIT('h1)
	) name8049 (
		_w9045_,
		_w9047_,
		_w9051_
	);
	LUT2 #(
		.INIT('h1)
	) name8050 (
		_w9048_,
		_w9051_,
		_w9052_
	);
	LUT2 #(
		.INIT('h1)
	) name8051 (
		_w9019_,
		_w9024_,
		_w9053_
	);
	LUT2 #(
		.INIT('h1)
	) name8052 (
		_w9025_,
		_w9053_,
		_w9054_
	);
	LUT2 #(
		.INIT('h8)
	) name8053 (
		_w9052_,
		_w9054_,
		_w9055_
	);
	LUT2 #(
		.INIT('h2)
	) name8054 (
		_w9026_,
		_w9027_,
		_w9056_
	);
	LUT2 #(
		.INIT('h2)
	) name8055 (
		_w9055_,
		_w9056_,
		_w9057_
	);
	LUT2 #(
		.INIT('h1)
	) name8056 (
		_w9042_,
		_w9043_,
		_w9058_
	);
	LUT2 #(
		.INIT('h2)
	) name8057 (
		_w9048_,
		_w9058_,
		_w9059_
	);
	LUT2 #(
		.INIT('h4)
	) name8058 (
		_w9048_,
		_w9058_,
		_w9060_
	);
	LUT2 #(
		.INIT('h1)
	) name8059 (
		_w9059_,
		_w9060_,
		_w9061_
	);
	LUT2 #(
		.INIT('h2)
	) name8060 (
		_w9057_,
		_w9061_,
		_w9062_
	);
	LUT2 #(
		.INIT('h4)
	) name8061 (
		_w9057_,
		_w9061_,
		_w9063_
	);
	LUT2 #(
		.INIT('h1)
	) name8062 (
		_w9026_,
		_w9029_,
		_w9064_
	);
	LUT2 #(
		.INIT('h2)
	) name8063 (
		_w9027_,
		_w9064_,
		_w9065_
	);
	LUT2 #(
		.INIT('h4)
	) name8064 (
		_w9027_,
		_w9064_,
		_w9066_
	);
	LUT2 #(
		.INIT('h1)
	) name8065 (
		_w9065_,
		_w9066_,
		_w9067_
	);
	LUT2 #(
		.INIT('h4)
	) name8066 (
		_w9063_,
		_w9067_,
		_w9068_
	);
	LUT2 #(
		.INIT('h1)
	) name8067 (
		_w9062_,
		_w9068_,
		_w9069_
	);
	LUT2 #(
		.INIT('h2)
	) name8068 (
		_w9050_,
		_w9069_,
		_w9070_
	);
	LUT2 #(
		.INIT('h4)
	) name8069 (
		_w9050_,
		_w9069_,
		_w9071_
	);
	LUT2 #(
		.INIT('h1)
	) name8070 (
		_w9070_,
		_w9071_,
		_w9072_
	);
	LUT2 #(
		.INIT('h8)
	) name8071 (
		_w9031_,
		_w9072_,
		_w9073_
	);
	LUT2 #(
		.INIT('h1)
	) name8072 (
		_w9031_,
		_w9072_,
		_w9074_
	);
	LUT2 #(
		.INIT('h1)
	) name8073 (
		_w9073_,
		_w9074_,
		_w9075_
	);
	LUT2 #(
		.INIT('h8)
	) name8074 (
		\A[550] ,
		\A[551] ,
		_w9076_
	);
	LUT2 #(
		.INIT('h8)
	) name8075 (
		\A[547] ,
		\A[548] ,
		_w9077_
	);
	LUT2 #(
		.INIT('h1)
	) name8076 (
		\A[547] ,
		\A[548] ,
		_w9078_
	);
	LUT2 #(
		.INIT('h1)
	) name8077 (
		_w9077_,
		_w9078_,
		_w9079_
	);
	LUT2 #(
		.INIT('h8)
	) name8078 (
		\A[549] ,
		_w9079_,
		_w9080_
	);
	LUT2 #(
		.INIT('h1)
	) name8079 (
		\A[549] ,
		_w9079_,
		_w9081_
	);
	LUT2 #(
		.INIT('h1)
	) name8080 (
		_w9080_,
		_w9081_,
		_w9082_
	);
	LUT2 #(
		.INIT('h1)
	) name8081 (
		\A[550] ,
		\A[551] ,
		_w9083_
	);
	LUT2 #(
		.INIT('h1)
	) name8082 (
		_w9076_,
		_w9083_,
		_w9084_
	);
	LUT2 #(
		.INIT('h8)
	) name8083 (
		\A[552] ,
		_w9084_,
		_w9085_
	);
	LUT2 #(
		.INIT('h1)
	) name8084 (
		\A[552] ,
		_w9084_,
		_w9086_
	);
	LUT2 #(
		.INIT('h1)
	) name8085 (
		_w9085_,
		_w9086_,
		_w9087_
	);
	LUT2 #(
		.INIT('h8)
	) name8086 (
		_w9082_,
		_w9087_,
		_w9088_
	);
	LUT2 #(
		.INIT('h8)
	) name8087 (
		_w9076_,
		_w9088_,
		_w9089_
	);
	LUT2 #(
		.INIT('h1)
	) name8088 (
		_w9077_,
		_w9080_,
		_w9090_
	);
	LUT2 #(
		.INIT('h1)
	) name8089 (
		_w9076_,
		_w9085_,
		_w9091_
	);
	LUT2 #(
		.INIT('h4)
	) name8090 (
		_w9088_,
		_w9091_,
		_w9092_
	);
	LUT2 #(
		.INIT('h1)
	) name8091 (
		_w9090_,
		_w9092_,
		_w9093_
	);
	LUT2 #(
		.INIT('h1)
	) name8092 (
		_w9089_,
		_w9093_,
		_w9094_
	);
	LUT2 #(
		.INIT('h8)
	) name8093 (
		\A[556] ,
		\A[557] ,
		_w9095_
	);
	LUT2 #(
		.INIT('h1)
	) name8094 (
		\A[556] ,
		\A[557] ,
		_w9096_
	);
	LUT2 #(
		.INIT('h1)
	) name8095 (
		_w9095_,
		_w9096_,
		_w9097_
	);
	LUT2 #(
		.INIT('h8)
	) name8096 (
		\A[558] ,
		_w9097_,
		_w9098_
	);
	LUT2 #(
		.INIT('h1)
	) name8097 (
		_w9095_,
		_w9098_,
		_w9099_
	);
	LUT2 #(
		.INIT('h8)
	) name8098 (
		\A[553] ,
		\A[554] ,
		_w9100_
	);
	LUT2 #(
		.INIT('h1)
	) name8099 (
		\A[553] ,
		\A[554] ,
		_w9101_
	);
	LUT2 #(
		.INIT('h1)
	) name8100 (
		_w9100_,
		_w9101_,
		_w9102_
	);
	LUT2 #(
		.INIT('h8)
	) name8101 (
		\A[555] ,
		_w9102_,
		_w9103_
	);
	LUT2 #(
		.INIT('h1)
	) name8102 (
		_w9100_,
		_w9103_,
		_w9104_
	);
	LUT2 #(
		.INIT('h8)
	) name8103 (
		_w9099_,
		_w9104_,
		_w9105_
	);
	LUT2 #(
		.INIT('h1)
	) name8104 (
		_w9099_,
		_w9104_,
		_w9106_
	);
	LUT2 #(
		.INIT('h1)
	) name8105 (
		\A[555] ,
		_w9102_,
		_w9107_
	);
	LUT2 #(
		.INIT('h1)
	) name8106 (
		_w9103_,
		_w9107_,
		_w9108_
	);
	LUT2 #(
		.INIT('h1)
	) name8107 (
		\A[558] ,
		_w9097_,
		_w9109_
	);
	LUT2 #(
		.INIT('h1)
	) name8108 (
		_w9098_,
		_w9109_,
		_w9110_
	);
	LUT2 #(
		.INIT('h8)
	) name8109 (
		_w9108_,
		_w9110_,
		_w9111_
	);
	LUT2 #(
		.INIT('h1)
	) name8110 (
		_w9106_,
		_w9111_,
		_w9112_
	);
	LUT2 #(
		.INIT('h1)
	) name8111 (
		_w9105_,
		_w9112_,
		_w9113_
	);
	LUT2 #(
		.INIT('h1)
	) name8112 (
		_w9108_,
		_w9110_,
		_w9114_
	);
	LUT2 #(
		.INIT('h1)
	) name8113 (
		_w9111_,
		_w9114_,
		_w9115_
	);
	LUT2 #(
		.INIT('h1)
	) name8114 (
		_w9082_,
		_w9087_,
		_w9116_
	);
	LUT2 #(
		.INIT('h1)
	) name8115 (
		_w9088_,
		_w9116_,
		_w9117_
	);
	LUT2 #(
		.INIT('h8)
	) name8116 (
		_w9115_,
		_w9117_,
		_w9118_
	);
	LUT2 #(
		.INIT('h2)
	) name8117 (
		_w9089_,
		_w9090_,
		_w9119_
	);
	LUT2 #(
		.INIT('h2)
	) name8118 (
		_w9118_,
		_w9119_,
		_w9120_
	);
	LUT2 #(
		.INIT('h1)
	) name8119 (
		_w9105_,
		_w9106_,
		_w9121_
	);
	LUT2 #(
		.INIT('h2)
	) name8120 (
		_w9111_,
		_w9121_,
		_w9122_
	);
	LUT2 #(
		.INIT('h4)
	) name8121 (
		_w9111_,
		_w9121_,
		_w9123_
	);
	LUT2 #(
		.INIT('h1)
	) name8122 (
		_w9122_,
		_w9123_,
		_w9124_
	);
	LUT2 #(
		.INIT('h2)
	) name8123 (
		_w9120_,
		_w9124_,
		_w9125_
	);
	LUT2 #(
		.INIT('h4)
	) name8124 (
		_w9120_,
		_w9124_,
		_w9126_
	);
	LUT2 #(
		.INIT('h1)
	) name8125 (
		_w9089_,
		_w9092_,
		_w9127_
	);
	LUT2 #(
		.INIT('h2)
	) name8126 (
		_w9090_,
		_w9127_,
		_w9128_
	);
	LUT2 #(
		.INIT('h4)
	) name8127 (
		_w9090_,
		_w9127_,
		_w9129_
	);
	LUT2 #(
		.INIT('h1)
	) name8128 (
		_w9128_,
		_w9129_,
		_w9130_
	);
	LUT2 #(
		.INIT('h4)
	) name8129 (
		_w9126_,
		_w9130_,
		_w9131_
	);
	LUT2 #(
		.INIT('h1)
	) name8130 (
		_w9125_,
		_w9131_,
		_w9132_
	);
	LUT2 #(
		.INIT('h2)
	) name8131 (
		_w9113_,
		_w9132_,
		_w9133_
	);
	LUT2 #(
		.INIT('h4)
	) name8132 (
		_w9113_,
		_w9132_,
		_w9134_
	);
	LUT2 #(
		.INIT('h1)
	) name8133 (
		_w9133_,
		_w9134_,
		_w9135_
	);
	LUT2 #(
		.INIT('h8)
	) name8134 (
		_w9094_,
		_w9135_,
		_w9136_
	);
	LUT2 #(
		.INIT('h1)
	) name8135 (
		_w9094_,
		_w9135_,
		_w9137_
	);
	LUT2 #(
		.INIT('h1)
	) name8136 (
		_w9136_,
		_w9137_,
		_w9138_
	);
	LUT2 #(
		.INIT('h1)
	) name8137 (
		_w9075_,
		_w9138_,
		_w9139_
	);
	LUT2 #(
		.INIT('h8)
	) name8138 (
		_w9075_,
		_w9138_,
		_w9140_
	);
	LUT2 #(
		.INIT('h1)
	) name8139 (
		_w9115_,
		_w9117_,
		_w9141_
	);
	LUT2 #(
		.INIT('h1)
	) name8140 (
		_w9118_,
		_w9141_,
		_w9142_
	);
	LUT2 #(
		.INIT('h1)
	) name8141 (
		_w9052_,
		_w9054_,
		_w9143_
	);
	LUT2 #(
		.INIT('h1)
	) name8142 (
		_w9055_,
		_w9143_,
		_w9144_
	);
	LUT2 #(
		.INIT('h8)
	) name8143 (
		_w9142_,
		_w9144_,
		_w9145_
	);
	LUT2 #(
		.INIT('h1)
	) name8144 (
		_w9125_,
		_w9126_,
		_w9146_
	);
	LUT2 #(
		.INIT('h8)
	) name8145 (
		_w9130_,
		_w9146_,
		_w9147_
	);
	LUT2 #(
		.INIT('h1)
	) name8146 (
		_w9130_,
		_w9146_,
		_w9148_
	);
	LUT2 #(
		.INIT('h1)
	) name8147 (
		_w9147_,
		_w9148_,
		_w9149_
	);
	LUT2 #(
		.INIT('h8)
	) name8148 (
		_w9145_,
		_w9149_,
		_w9150_
	);
	LUT2 #(
		.INIT('h1)
	) name8149 (
		_w9145_,
		_w9149_,
		_w9151_
	);
	LUT2 #(
		.INIT('h1)
	) name8150 (
		_w9062_,
		_w9063_,
		_w9152_
	);
	LUT2 #(
		.INIT('h8)
	) name8151 (
		_w9067_,
		_w9152_,
		_w9153_
	);
	LUT2 #(
		.INIT('h1)
	) name8152 (
		_w9067_,
		_w9152_,
		_w9154_
	);
	LUT2 #(
		.INIT('h1)
	) name8153 (
		_w9153_,
		_w9154_,
		_w9155_
	);
	LUT2 #(
		.INIT('h4)
	) name8154 (
		_w9151_,
		_w9155_,
		_w9156_
	);
	LUT2 #(
		.INIT('h1)
	) name8155 (
		_w9150_,
		_w9156_,
		_w9157_
	);
	LUT2 #(
		.INIT('h1)
	) name8156 (
		_w9140_,
		_w9157_,
		_w9158_
	);
	LUT2 #(
		.INIT('h1)
	) name8157 (
		_w9139_,
		_w9158_,
		_w9159_
	);
	LUT2 #(
		.INIT('h1)
	) name8158 (
		_w9094_,
		_w9134_,
		_w9160_
	);
	LUT2 #(
		.INIT('h1)
	) name8159 (
		_w9133_,
		_w9160_,
		_w9161_
	);
	LUT2 #(
		.INIT('h1)
	) name8160 (
		_w9159_,
		_w9161_,
		_w9162_
	);
	LUT2 #(
		.INIT('h8)
	) name8161 (
		_w9159_,
		_w9161_,
		_w9163_
	);
	LUT2 #(
		.INIT('h1)
	) name8162 (
		_w9031_,
		_w9071_,
		_w9164_
	);
	LUT2 #(
		.INIT('h1)
	) name8163 (
		_w9070_,
		_w9164_,
		_w9165_
	);
	LUT2 #(
		.INIT('h1)
	) name8164 (
		_w9163_,
		_w9165_,
		_w9166_
	);
	LUT2 #(
		.INIT('h1)
	) name8165 (
		_w9162_,
		_w9166_,
		_w9167_
	);
	LUT2 #(
		.INIT('h1)
	) name8166 (
		_w9162_,
		_w9163_,
		_w9168_
	);
	LUT2 #(
		.INIT('h4)
	) name8167 (
		_w9165_,
		_w9168_,
		_w9169_
	);
	LUT2 #(
		.INIT('h2)
	) name8168 (
		_w9165_,
		_w9168_,
		_w9170_
	);
	LUT2 #(
		.INIT('h1)
	) name8169 (
		_w9169_,
		_w9170_,
		_w9171_
	);
	LUT2 #(
		.INIT('h8)
	) name8170 (
		\A[514] ,
		\A[515] ,
		_w9172_
	);
	LUT2 #(
		.INIT('h8)
	) name8171 (
		\A[511] ,
		\A[512] ,
		_w9173_
	);
	LUT2 #(
		.INIT('h1)
	) name8172 (
		\A[511] ,
		\A[512] ,
		_w9174_
	);
	LUT2 #(
		.INIT('h1)
	) name8173 (
		_w9173_,
		_w9174_,
		_w9175_
	);
	LUT2 #(
		.INIT('h8)
	) name8174 (
		\A[513] ,
		_w9175_,
		_w9176_
	);
	LUT2 #(
		.INIT('h1)
	) name8175 (
		\A[513] ,
		_w9175_,
		_w9177_
	);
	LUT2 #(
		.INIT('h1)
	) name8176 (
		_w9176_,
		_w9177_,
		_w9178_
	);
	LUT2 #(
		.INIT('h1)
	) name8177 (
		\A[514] ,
		\A[515] ,
		_w9179_
	);
	LUT2 #(
		.INIT('h1)
	) name8178 (
		_w9172_,
		_w9179_,
		_w9180_
	);
	LUT2 #(
		.INIT('h8)
	) name8179 (
		\A[516] ,
		_w9180_,
		_w9181_
	);
	LUT2 #(
		.INIT('h1)
	) name8180 (
		\A[516] ,
		_w9180_,
		_w9182_
	);
	LUT2 #(
		.INIT('h1)
	) name8181 (
		_w9181_,
		_w9182_,
		_w9183_
	);
	LUT2 #(
		.INIT('h8)
	) name8182 (
		_w9178_,
		_w9183_,
		_w9184_
	);
	LUT2 #(
		.INIT('h8)
	) name8183 (
		_w9172_,
		_w9184_,
		_w9185_
	);
	LUT2 #(
		.INIT('h1)
	) name8184 (
		_w9173_,
		_w9176_,
		_w9186_
	);
	LUT2 #(
		.INIT('h1)
	) name8185 (
		_w9172_,
		_w9181_,
		_w9187_
	);
	LUT2 #(
		.INIT('h4)
	) name8186 (
		_w9184_,
		_w9187_,
		_w9188_
	);
	LUT2 #(
		.INIT('h1)
	) name8187 (
		_w9186_,
		_w9188_,
		_w9189_
	);
	LUT2 #(
		.INIT('h1)
	) name8188 (
		_w9185_,
		_w9189_,
		_w9190_
	);
	LUT2 #(
		.INIT('h8)
	) name8189 (
		\A[520] ,
		\A[521] ,
		_w9191_
	);
	LUT2 #(
		.INIT('h1)
	) name8190 (
		\A[520] ,
		\A[521] ,
		_w9192_
	);
	LUT2 #(
		.INIT('h1)
	) name8191 (
		_w9191_,
		_w9192_,
		_w9193_
	);
	LUT2 #(
		.INIT('h8)
	) name8192 (
		\A[522] ,
		_w9193_,
		_w9194_
	);
	LUT2 #(
		.INIT('h1)
	) name8193 (
		_w9191_,
		_w9194_,
		_w9195_
	);
	LUT2 #(
		.INIT('h8)
	) name8194 (
		\A[517] ,
		\A[518] ,
		_w9196_
	);
	LUT2 #(
		.INIT('h1)
	) name8195 (
		\A[517] ,
		\A[518] ,
		_w9197_
	);
	LUT2 #(
		.INIT('h1)
	) name8196 (
		_w9196_,
		_w9197_,
		_w9198_
	);
	LUT2 #(
		.INIT('h8)
	) name8197 (
		\A[519] ,
		_w9198_,
		_w9199_
	);
	LUT2 #(
		.INIT('h1)
	) name8198 (
		_w9196_,
		_w9199_,
		_w9200_
	);
	LUT2 #(
		.INIT('h8)
	) name8199 (
		_w9195_,
		_w9200_,
		_w9201_
	);
	LUT2 #(
		.INIT('h1)
	) name8200 (
		_w9195_,
		_w9200_,
		_w9202_
	);
	LUT2 #(
		.INIT('h1)
	) name8201 (
		\A[519] ,
		_w9198_,
		_w9203_
	);
	LUT2 #(
		.INIT('h1)
	) name8202 (
		_w9199_,
		_w9203_,
		_w9204_
	);
	LUT2 #(
		.INIT('h1)
	) name8203 (
		\A[522] ,
		_w9193_,
		_w9205_
	);
	LUT2 #(
		.INIT('h1)
	) name8204 (
		_w9194_,
		_w9205_,
		_w9206_
	);
	LUT2 #(
		.INIT('h8)
	) name8205 (
		_w9204_,
		_w9206_,
		_w9207_
	);
	LUT2 #(
		.INIT('h1)
	) name8206 (
		_w9202_,
		_w9207_,
		_w9208_
	);
	LUT2 #(
		.INIT('h1)
	) name8207 (
		_w9201_,
		_w9208_,
		_w9209_
	);
	LUT2 #(
		.INIT('h1)
	) name8208 (
		_w9204_,
		_w9206_,
		_w9210_
	);
	LUT2 #(
		.INIT('h1)
	) name8209 (
		_w9207_,
		_w9210_,
		_w9211_
	);
	LUT2 #(
		.INIT('h1)
	) name8210 (
		_w9178_,
		_w9183_,
		_w9212_
	);
	LUT2 #(
		.INIT('h1)
	) name8211 (
		_w9184_,
		_w9212_,
		_w9213_
	);
	LUT2 #(
		.INIT('h8)
	) name8212 (
		_w9211_,
		_w9213_,
		_w9214_
	);
	LUT2 #(
		.INIT('h2)
	) name8213 (
		_w9185_,
		_w9186_,
		_w9215_
	);
	LUT2 #(
		.INIT('h2)
	) name8214 (
		_w9214_,
		_w9215_,
		_w9216_
	);
	LUT2 #(
		.INIT('h1)
	) name8215 (
		_w9201_,
		_w9202_,
		_w9217_
	);
	LUT2 #(
		.INIT('h2)
	) name8216 (
		_w9207_,
		_w9217_,
		_w9218_
	);
	LUT2 #(
		.INIT('h4)
	) name8217 (
		_w9207_,
		_w9217_,
		_w9219_
	);
	LUT2 #(
		.INIT('h1)
	) name8218 (
		_w9218_,
		_w9219_,
		_w9220_
	);
	LUT2 #(
		.INIT('h2)
	) name8219 (
		_w9216_,
		_w9220_,
		_w9221_
	);
	LUT2 #(
		.INIT('h4)
	) name8220 (
		_w9216_,
		_w9220_,
		_w9222_
	);
	LUT2 #(
		.INIT('h1)
	) name8221 (
		_w9185_,
		_w9188_,
		_w9223_
	);
	LUT2 #(
		.INIT('h2)
	) name8222 (
		_w9186_,
		_w9223_,
		_w9224_
	);
	LUT2 #(
		.INIT('h4)
	) name8223 (
		_w9186_,
		_w9223_,
		_w9225_
	);
	LUT2 #(
		.INIT('h1)
	) name8224 (
		_w9224_,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('h4)
	) name8225 (
		_w9222_,
		_w9226_,
		_w9227_
	);
	LUT2 #(
		.INIT('h1)
	) name8226 (
		_w9221_,
		_w9227_,
		_w9228_
	);
	LUT2 #(
		.INIT('h2)
	) name8227 (
		_w9209_,
		_w9228_,
		_w9229_
	);
	LUT2 #(
		.INIT('h4)
	) name8228 (
		_w9209_,
		_w9228_,
		_w9230_
	);
	LUT2 #(
		.INIT('h1)
	) name8229 (
		_w9229_,
		_w9230_,
		_w9231_
	);
	LUT2 #(
		.INIT('h8)
	) name8230 (
		_w9190_,
		_w9231_,
		_w9232_
	);
	LUT2 #(
		.INIT('h1)
	) name8231 (
		_w9190_,
		_w9231_,
		_w9233_
	);
	LUT2 #(
		.INIT('h1)
	) name8232 (
		_w9232_,
		_w9233_,
		_w9234_
	);
	LUT2 #(
		.INIT('h8)
	) name8233 (
		\A[526] ,
		\A[527] ,
		_w9235_
	);
	LUT2 #(
		.INIT('h8)
	) name8234 (
		\A[523] ,
		\A[524] ,
		_w9236_
	);
	LUT2 #(
		.INIT('h1)
	) name8235 (
		\A[523] ,
		\A[524] ,
		_w9237_
	);
	LUT2 #(
		.INIT('h1)
	) name8236 (
		_w9236_,
		_w9237_,
		_w9238_
	);
	LUT2 #(
		.INIT('h8)
	) name8237 (
		\A[525] ,
		_w9238_,
		_w9239_
	);
	LUT2 #(
		.INIT('h1)
	) name8238 (
		\A[525] ,
		_w9238_,
		_w9240_
	);
	LUT2 #(
		.INIT('h1)
	) name8239 (
		_w9239_,
		_w9240_,
		_w9241_
	);
	LUT2 #(
		.INIT('h1)
	) name8240 (
		\A[526] ,
		\A[527] ,
		_w9242_
	);
	LUT2 #(
		.INIT('h1)
	) name8241 (
		_w9235_,
		_w9242_,
		_w9243_
	);
	LUT2 #(
		.INIT('h8)
	) name8242 (
		\A[528] ,
		_w9243_,
		_w9244_
	);
	LUT2 #(
		.INIT('h1)
	) name8243 (
		\A[528] ,
		_w9243_,
		_w9245_
	);
	LUT2 #(
		.INIT('h1)
	) name8244 (
		_w9244_,
		_w9245_,
		_w9246_
	);
	LUT2 #(
		.INIT('h8)
	) name8245 (
		_w9241_,
		_w9246_,
		_w9247_
	);
	LUT2 #(
		.INIT('h8)
	) name8246 (
		_w9235_,
		_w9247_,
		_w9248_
	);
	LUT2 #(
		.INIT('h1)
	) name8247 (
		_w9236_,
		_w9239_,
		_w9249_
	);
	LUT2 #(
		.INIT('h1)
	) name8248 (
		_w9235_,
		_w9244_,
		_w9250_
	);
	LUT2 #(
		.INIT('h4)
	) name8249 (
		_w9247_,
		_w9250_,
		_w9251_
	);
	LUT2 #(
		.INIT('h1)
	) name8250 (
		_w9249_,
		_w9251_,
		_w9252_
	);
	LUT2 #(
		.INIT('h1)
	) name8251 (
		_w9248_,
		_w9252_,
		_w9253_
	);
	LUT2 #(
		.INIT('h8)
	) name8252 (
		\A[532] ,
		\A[533] ,
		_w9254_
	);
	LUT2 #(
		.INIT('h1)
	) name8253 (
		\A[532] ,
		\A[533] ,
		_w9255_
	);
	LUT2 #(
		.INIT('h1)
	) name8254 (
		_w9254_,
		_w9255_,
		_w9256_
	);
	LUT2 #(
		.INIT('h8)
	) name8255 (
		\A[534] ,
		_w9256_,
		_w9257_
	);
	LUT2 #(
		.INIT('h1)
	) name8256 (
		_w9254_,
		_w9257_,
		_w9258_
	);
	LUT2 #(
		.INIT('h8)
	) name8257 (
		\A[529] ,
		\A[530] ,
		_w9259_
	);
	LUT2 #(
		.INIT('h1)
	) name8258 (
		\A[529] ,
		\A[530] ,
		_w9260_
	);
	LUT2 #(
		.INIT('h1)
	) name8259 (
		_w9259_,
		_w9260_,
		_w9261_
	);
	LUT2 #(
		.INIT('h8)
	) name8260 (
		\A[531] ,
		_w9261_,
		_w9262_
	);
	LUT2 #(
		.INIT('h1)
	) name8261 (
		_w9259_,
		_w9262_,
		_w9263_
	);
	LUT2 #(
		.INIT('h8)
	) name8262 (
		_w9258_,
		_w9263_,
		_w9264_
	);
	LUT2 #(
		.INIT('h1)
	) name8263 (
		_w9258_,
		_w9263_,
		_w9265_
	);
	LUT2 #(
		.INIT('h1)
	) name8264 (
		\A[531] ,
		_w9261_,
		_w9266_
	);
	LUT2 #(
		.INIT('h1)
	) name8265 (
		_w9262_,
		_w9266_,
		_w9267_
	);
	LUT2 #(
		.INIT('h1)
	) name8266 (
		\A[534] ,
		_w9256_,
		_w9268_
	);
	LUT2 #(
		.INIT('h1)
	) name8267 (
		_w9257_,
		_w9268_,
		_w9269_
	);
	LUT2 #(
		.INIT('h8)
	) name8268 (
		_w9267_,
		_w9269_,
		_w9270_
	);
	LUT2 #(
		.INIT('h1)
	) name8269 (
		_w9265_,
		_w9270_,
		_w9271_
	);
	LUT2 #(
		.INIT('h1)
	) name8270 (
		_w9264_,
		_w9271_,
		_w9272_
	);
	LUT2 #(
		.INIT('h1)
	) name8271 (
		_w9267_,
		_w9269_,
		_w9273_
	);
	LUT2 #(
		.INIT('h1)
	) name8272 (
		_w9270_,
		_w9273_,
		_w9274_
	);
	LUT2 #(
		.INIT('h1)
	) name8273 (
		_w9241_,
		_w9246_,
		_w9275_
	);
	LUT2 #(
		.INIT('h1)
	) name8274 (
		_w9247_,
		_w9275_,
		_w9276_
	);
	LUT2 #(
		.INIT('h8)
	) name8275 (
		_w9274_,
		_w9276_,
		_w9277_
	);
	LUT2 #(
		.INIT('h2)
	) name8276 (
		_w9248_,
		_w9249_,
		_w9278_
	);
	LUT2 #(
		.INIT('h2)
	) name8277 (
		_w9277_,
		_w9278_,
		_w9279_
	);
	LUT2 #(
		.INIT('h1)
	) name8278 (
		_w9264_,
		_w9265_,
		_w9280_
	);
	LUT2 #(
		.INIT('h2)
	) name8279 (
		_w9270_,
		_w9280_,
		_w9281_
	);
	LUT2 #(
		.INIT('h4)
	) name8280 (
		_w9270_,
		_w9280_,
		_w9282_
	);
	LUT2 #(
		.INIT('h1)
	) name8281 (
		_w9281_,
		_w9282_,
		_w9283_
	);
	LUT2 #(
		.INIT('h2)
	) name8282 (
		_w9279_,
		_w9283_,
		_w9284_
	);
	LUT2 #(
		.INIT('h4)
	) name8283 (
		_w9279_,
		_w9283_,
		_w9285_
	);
	LUT2 #(
		.INIT('h1)
	) name8284 (
		_w9248_,
		_w9251_,
		_w9286_
	);
	LUT2 #(
		.INIT('h2)
	) name8285 (
		_w9249_,
		_w9286_,
		_w9287_
	);
	LUT2 #(
		.INIT('h4)
	) name8286 (
		_w9249_,
		_w9286_,
		_w9288_
	);
	LUT2 #(
		.INIT('h1)
	) name8287 (
		_w9287_,
		_w9288_,
		_w9289_
	);
	LUT2 #(
		.INIT('h4)
	) name8288 (
		_w9285_,
		_w9289_,
		_w9290_
	);
	LUT2 #(
		.INIT('h1)
	) name8289 (
		_w9284_,
		_w9290_,
		_w9291_
	);
	LUT2 #(
		.INIT('h2)
	) name8290 (
		_w9272_,
		_w9291_,
		_w9292_
	);
	LUT2 #(
		.INIT('h4)
	) name8291 (
		_w9272_,
		_w9291_,
		_w9293_
	);
	LUT2 #(
		.INIT('h1)
	) name8292 (
		_w9292_,
		_w9293_,
		_w9294_
	);
	LUT2 #(
		.INIT('h8)
	) name8293 (
		_w9253_,
		_w9294_,
		_w9295_
	);
	LUT2 #(
		.INIT('h1)
	) name8294 (
		_w9253_,
		_w9294_,
		_w9296_
	);
	LUT2 #(
		.INIT('h1)
	) name8295 (
		_w9295_,
		_w9296_,
		_w9297_
	);
	LUT2 #(
		.INIT('h1)
	) name8296 (
		_w9234_,
		_w9297_,
		_w9298_
	);
	LUT2 #(
		.INIT('h8)
	) name8297 (
		_w9234_,
		_w9297_,
		_w9299_
	);
	LUT2 #(
		.INIT('h1)
	) name8298 (
		_w9274_,
		_w9276_,
		_w9300_
	);
	LUT2 #(
		.INIT('h1)
	) name8299 (
		_w9277_,
		_w9300_,
		_w9301_
	);
	LUT2 #(
		.INIT('h1)
	) name8300 (
		_w9211_,
		_w9213_,
		_w9302_
	);
	LUT2 #(
		.INIT('h1)
	) name8301 (
		_w9214_,
		_w9302_,
		_w9303_
	);
	LUT2 #(
		.INIT('h8)
	) name8302 (
		_w9301_,
		_w9303_,
		_w9304_
	);
	LUT2 #(
		.INIT('h1)
	) name8303 (
		_w9284_,
		_w9285_,
		_w9305_
	);
	LUT2 #(
		.INIT('h8)
	) name8304 (
		_w9289_,
		_w9305_,
		_w9306_
	);
	LUT2 #(
		.INIT('h1)
	) name8305 (
		_w9289_,
		_w9305_,
		_w9307_
	);
	LUT2 #(
		.INIT('h1)
	) name8306 (
		_w9306_,
		_w9307_,
		_w9308_
	);
	LUT2 #(
		.INIT('h8)
	) name8307 (
		_w9304_,
		_w9308_,
		_w9309_
	);
	LUT2 #(
		.INIT('h1)
	) name8308 (
		_w9304_,
		_w9308_,
		_w9310_
	);
	LUT2 #(
		.INIT('h1)
	) name8309 (
		_w9221_,
		_w9222_,
		_w9311_
	);
	LUT2 #(
		.INIT('h8)
	) name8310 (
		_w9226_,
		_w9311_,
		_w9312_
	);
	LUT2 #(
		.INIT('h1)
	) name8311 (
		_w9226_,
		_w9311_,
		_w9313_
	);
	LUT2 #(
		.INIT('h1)
	) name8312 (
		_w9312_,
		_w9313_,
		_w9314_
	);
	LUT2 #(
		.INIT('h4)
	) name8313 (
		_w9310_,
		_w9314_,
		_w9315_
	);
	LUT2 #(
		.INIT('h1)
	) name8314 (
		_w9309_,
		_w9315_,
		_w9316_
	);
	LUT2 #(
		.INIT('h1)
	) name8315 (
		_w9299_,
		_w9316_,
		_w9317_
	);
	LUT2 #(
		.INIT('h1)
	) name8316 (
		_w9298_,
		_w9317_,
		_w9318_
	);
	LUT2 #(
		.INIT('h1)
	) name8317 (
		_w9253_,
		_w9293_,
		_w9319_
	);
	LUT2 #(
		.INIT('h1)
	) name8318 (
		_w9292_,
		_w9319_,
		_w9320_
	);
	LUT2 #(
		.INIT('h1)
	) name8319 (
		_w9318_,
		_w9320_,
		_w9321_
	);
	LUT2 #(
		.INIT('h8)
	) name8320 (
		_w9318_,
		_w9320_,
		_w9322_
	);
	LUT2 #(
		.INIT('h1)
	) name8321 (
		_w9321_,
		_w9322_,
		_w9323_
	);
	LUT2 #(
		.INIT('h1)
	) name8322 (
		_w9190_,
		_w9230_,
		_w9324_
	);
	LUT2 #(
		.INIT('h1)
	) name8323 (
		_w9229_,
		_w9324_,
		_w9325_
	);
	LUT2 #(
		.INIT('h2)
	) name8324 (
		_w9323_,
		_w9325_,
		_w9326_
	);
	LUT2 #(
		.INIT('h4)
	) name8325 (
		_w9323_,
		_w9325_,
		_w9327_
	);
	LUT2 #(
		.INIT('h1)
	) name8326 (
		_w9326_,
		_w9327_,
		_w9328_
	);
	LUT2 #(
		.INIT('h1)
	) name8327 (
		_w9171_,
		_w9328_,
		_w9329_
	);
	LUT2 #(
		.INIT('h8)
	) name8328 (
		_w9171_,
		_w9328_,
		_w9330_
	);
	LUT2 #(
		.INIT('h1)
	) name8329 (
		_w9298_,
		_w9299_,
		_w9331_
	);
	LUT2 #(
		.INIT('h4)
	) name8330 (
		_w9316_,
		_w9331_,
		_w9332_
	);
	LUT2 #(
		.INIT('h2)
	) name8331 (
		_w9316_,
		_w9331_,
		_w9333_
	);
	LUT2 #(
		.INIT('h1)
	) name8332 (
		_w9332_,
		_w9333_,
		_w9334_
	);
	LUT2 #(
		.INIT('h1)
	) name8333 (
		_w9139_,
		_w9140_,
		_w9335_
	);
	LUT2 #(
		.INIT('h4)
	) name8334 (
		_w9157_,
		_w9335_,
		_w9336_
	);
	LUT2 #(
		.INIT('h2)
	) name8335 (
		_w9157_,
		_w9335_,
		_w9337_
	);
	LUT2 #(
		.INIT('h1)
	) name8336 (
		_w9336_,
		_w9337_,
		_w9338_
	);
	LUT2 #(
		.INIT('h1)
	) name8337 (
		_w9334_,
		_w9338_,
		_w9339_
	);
	LUT2 #(
		.INIT('h8)
	) name8338 (
		_w9334_,
		_w9338_,
		_w9340_
	);
	LUT2 #(
		.INIT('h1)
	) name8339 (
		_w9142_,
		_w9144_,
		_w9341_
	);
	LUT2 #(
		.INIT('h1)
	) name8340 (
		_w9145_,
		_w9341_,
		_w9342_
	);
	LUT2 #(
		.INIT('h1)
	) name8341 (
		_w9301_,
		_w9303_,
		_w9343_
	);
	LUT2 #(
		.INIT('h1)
	) name8342 (
		_w9304_,
		_w9343_,
		_w9344_
	);
	LUT2 #(
		.INIT('h8)
	) name8343 (
		_w9342_,
		_w9344_,
		_w9345_
	);
	LUT2 #(
		.INIT('h1)
	) name8344 (
		_w9150_,
		_w9151_,
		_w9346_
	);
	LUT2 #(
		.INIT('h4)
	) name8345 (
		_w9155_,
		_w9346_,
		_w9347_
	);
	LUT2 #(
		.INIT('h2)
	) name8346 (
		_w9155_,
		_w9346_,
		_w9348_
	);
	LUT2 #(
		.INIT('h1)
	) name8347 (
		_w9347_,
		_w9348_,
		_w9349_
	);
	LUT2 #(
		.INIT('h2)
	) name8348 (
		_w9345_,
		_w9349_,
		_w9350_
	);
	LUT2 #(
		.INIT('h4)
	) name8349 (
		_w9345_,
		_w9349_,
		_w9351_
	);
	LUT2 #(
		.INIT('h1)
	) name8350 (
		_w9309_,
		_w9310_,
		_w9352_
	);
	LUT2 #(
		.INIT('h4)
	) name8351 (
		_w9314_,
		_w9352_,
		_w9353_
	);
	LUT2 #(
		.INIT('h2)
	) name8352 (
		_w9314_,
		_w9352_,
		_w9354_
	);
	LUT2 #(
		.INIT('h1)
	) name8353 (
		_w9353_,
		_w9354_,
		_w9355_
	);
	LUT2 #(
		.INIT('h1)
	) name8354 (
		_w9351_,
		_w9355_,
		_w9356_
	);
	LUT2 #(
		.INIT('h1)
	) name8355 (
		_w9350_,
		_w9356_,
		_w9357_
	);
	LUT2 #(
		.INIT('h4)
	) name8356 (
		_w9340_,
		_w9357_,
		_w9358_
	);
	LUT2 #(
		.INIT('h1)
	) name8357 (
		_w9339_,
		_w9358_,
		_w9359_
	);
	LUT2 #(
		.INIT('h1)
	) name8358 (
		_w9330_,
		_w9359_,
		_w9360_
	);
	LUT2 #(
		.INIT('h1)
	) name8359 (
		_w9329_,
		_w9360_,
		_w9361_
	);
	LUT2 #(
		.INIT('h2)
	) name8360 (
		_w9167_,
		_w9361_,
		_w9362_
	);
	LUT2 #(
		.INIT('h4)
	) name8361 (
		_w9167_,
		_w9361_,
		_w9363_
	);
	LUT2 #(
		.INIT('h1)
	) name8362 (
		_w9362_,
		_w9363_,
		_w9364_
	);
	LUT2 #(
		.INIT('h1)
	) name8363 (
		_w9322_,
		_w9325_,
		_w9365_
	);
	LUT2 #(
		.INIT('h1)
	) name8364 (
		_w9321_,
		_w9365_,
		_w9366_
	);
	LUT2 #(
		.INIT('h8)
	) name8365 (
		_w9364_,
		_w9366_,
		_w9367_
	);
	LUT2 #(
		.INIT('h1)
	) name8366 (
		_w9364_,
		_w9366_,
		_w9368_
	);
	LUT2 #(
		.INIT('h1)
	) name8367 (
		_w9367_,
		_w9368_,
		_w9369_
	);
	LUT2 #(
		.INIT('h1)
	) name8368 (
		_w9012_,
		_w9369_,
		_w9370_
	);
	LUT2 #(
		.INIT('h8)
	) name8369 (
		_w9012_,
		_w9369_,
		_w9371_
	);
	LUT2 #(
		.INIT('h1)
	) name8370 (
		_w9329_,
		_w9330_,
		_w9372_
	);
	LUT2 #(
		.INIT('h4)
	) name8371 (
		_w9359_,
		_w9372_,
		_w9373_
	);
	LUT2 #(
		.INIT('h2)
	) name8372 (
		_w9359_,
		_w9372_,
		_w9374_
	);
	LUT2 #(
		.INIT('h1)
	) name8373 (
		_w9373_,
		_w9374_,
		_w9375_
	);
	LUT2 #(
		.INIT('h1)
	) name8374 (
		_w8972_,
		_w8973_,
		_w9376_
	);
	LUT2 #(
		.INIT('h4)
	) name8375 (
		_w9002_,
		_w9376_,
		_w9377_
	);
	LUT2 #(
		.INIT('h2)
	) name8376 (
		_w9002_,
		_w9376_,
		_w9378_
	);
	LUT2 #(
		.INIT('h1)
	) name8377 (
		_w9377_,
		_w9378_,
		_w9379_
	);
	LUT2 #(
		.INIT('h1)
	) name8378 (
		_w9375_,
		_w9379_,
		_w9380_
	);
	LUT2 #(
		.INIT('h8)
	) name8379 (
		_w9375_,
		_w9379_,
		_w9381_
	);
	LUT2 #(
		.INIT('h1)
	) name8380 (
		_w8982_,
		_w8983_,
		_w9382_
	);
	LUT2 #(
		.INIT('h4)
	) name8381 (
		_w9000_,
		_w9382_,
		_w9383_
	);
	LUT2 #(
		.INIT('h2)
	) name8382 (
		_w9000_,
		_w9382_,
		_w9384_
	);
	LUT2 #(
		.INIT('h1)
	) name8383 (
		_w9383_,
		_w9384_,
		_w9385_
	);
	LUT2 #(
		.INIT('h1)
	) name8384 (
		_w9339_,
		_w9340_,
		_w9386_
	);
	LUT2 #(
		.INIT('h4)
	) name8385 (
		_w9357_,
		_w9386_,
		_w9387_
	);
	LUT2 #(
		.INIT('h2)
	) name8386 (
		_w9357_,
		_w9386_,
		_w9388_
	);
	LUT2 #(
		.INIT('h1)
	) name8387 (
		_w9387_,
		_w9388_,
		_w9389_
	);
	LUT2 #(
		.INIT('h1)
	) name8388 (
		_w9385_,
		_w9389_,
		_w9390_
	);
	LUT2 #(
		.INIT('h8)
	) name8389 (
		_w9385_,
		_w9389_,
		_w9391_
	);
	LUT2 #(
		.INIT('h1)
	) name8390 (
		_w8985_,
		_w8987_,
		_w9392_
	);
	LUT2 #(
		.INIT('h1)
	) name8391 (
		_w8988_,
		_w9392_,
		_w9393_
	);
	LUT2 #(
		.INIT('h1)
	) name8392 (
		_w9342_,
		_w9344_,
		_w9394_
	);
	LUT2 #(
		.INIT('h1)
	) name8393 (
		_w9345_,
		_w9394_,
		_w9395_
	);
	LUT2 #(
		.INIT('h8)
	) name8394 (
		_w9393_,
		_w9395_,
		_w9396_
	);
	LUT2 #(
		.INIT('h1)
	) name8395 (
		_w9350_,
		_w9351_,
		_w9397_
	);
	LUT2 #(
		.INIT('h4)
	) name8396 (
		_w9355_,
		_w9397_,
		_w9398_
	);
	LUT2 #(
		.INIT('h2)
	) name8397 (
		_w9355_,
		_w9397_,
		_w9399_
	);
	LUT2 #(
		.INIT('h1)
	) name8398 (
		_w9398_,
		_w9399_,
		_w9400_
	);
	LUT2 #(
		.INIT('h8)
	) name8399 (
		_w9396_,
		_w9400_,
		_w9401_
	);
	LUT2 #(
		.INIT('h1)
	) name8400 (
		_w9396_,
		_w9400_,
		_w9402_
	);
	LUT2 #(
		.INIT('h1)
	) name8401 (
		_w8993_,
		_w8994_,
		_w9403_
	);
	LUT2 #(
		.INIT('h4)
	) name8402 (
		_w8998_,
		_w9403_,
		_w9404_
	);
	LUT2 #(
		.INIT('h2)
	) name8403 (
		_w8998_,
		_w9403_,
		_w9405_
	);
	LUT2 #(
		.INIT('h1)
	) name8404 (
		_w9404_,
		_w9405_,
		_w9406_
	);
	LUT2 #(
		.INIT('h4)
	) name8405 (
		_w9402_,
		_w9406_,
		_w9407_
	);
	LUT2 #(
		.INIT('h1)
	) name8406 (
		_w9401_,
		_w9407_,
		_w9408_
	);
	LUT2 #(
		.INIT('h4)
	) name8407 (
		_w9391_,
		_w9408_,
		_w9409_
	);
	LUT2 #(
		.INIT('h1)
	) name8408 (
		_w9390_,
		_w9409_,
		_w9410_
	);
	LUT2 #(
		.INIT('h4)
	) name8409 (
		_w9381_,
		_w9410_,
		_w9411_
	);
	LUT2 #(
		.INIT('h1)
	) name8410 (
		_w9380_,
		_w9411_,
		_w9412_
	);
	LUT2 #(
		.INIT('h1)
	) name8411 (
		_w9371_,
		_w9412_,
		_w9413_
	);
	LUT2 #(
		.INIT('h1)
	) name8412 (
		_w9370_,
		_w9413_,
		_w9414_
	);
	LUT2 #(
		.INIT('h4)
	) name8413 (
		_w9006_,
		_w9009_,
		_w9415_
	);
	LUT2 #(
		.INIT('h1)
	) name8414 (
		_w9005_,
		_w9415_,
		_w9416_
	);
	LUT2 #(
		.INIT('h2)
	) name8415 (
		_w9414_,
		_w9416_,
		_w9417_
	);
	LUT2 #(
		.INIT('h4)
	) name8416 (
		_w9414_,
		_w9416_,
		_w9418_
	);
	LUT2 #(
		.INIT('h4)
	) name8417 (
		_w9363_,
		_w9366_,
		_w9419_
	);
	LUT2 #(
		.INIT('h1)
	) name8418 (
		_w9362_,
		_w9419_,
		_w9420_
	);
	LUT2 #(
		.INIT('h1)
	) name8419 (
		_w9418_,
		_w9420_,
		_w9421_
	);
	LUT2 #(
		.INIT('h1)
	) name8420 (
		_w9417_,
		_w9421_,
		_w9422_
	);
	LUT2 #(
		.INIT('h8)
	) name8421 (
		_w8655_,
		_w9422_,
		_w9423_
	);
	LUT2 #(
		.INIT('h1)
	) name8422 (
		_w8655_,
		_w9422_,
		_w9424_
	);
	LUT2 #(
		.INIT('h1)
	) name8423 (
		_w8650_,
		_w8651_,
		_w9425_
	);
	LUT2 #(
		.INIT('h4)
	) name8424 (
		_w8653_,
		_w9425_,
		_w9426_
	);
	LUT2 #(
		.INIT('h2)
	) name8425 (
		_w8653_,
		_w9425_,
		_w9427_
	);
	LUT2 #(
		.INIT('h1)
	) name8426 (
		_w9426_,
		_w9427_,
		_w9428_
	);
	LUT2 #(
		.INIT('h1)
	) name8427 (
		_w9417_,
		_w9418_,
		_w9429_
	);
	LUT2 #(
		.INIT('h4)
	) name8428 (
		_w9420_,
		_w9429_,
		_w9430_
	);
	LUT2 #(
		.INIT('h2)
	) name8429 (
		_w9420_,
		_w9429_,
		_w9431_
	);
	LUT2 #(
		.INIT('h1)
	) name8430 (
		_w9430_,
		_w9431_,
		_w9432_
	);
	LUT2 #(
		.INIT('h1)
	) name8431 (
		_w9428_,
		_w9432_,
		_w9433_
	);
	LUT2 #(
		.INIT('h8)
	) name8432 (
		_w9428_,
		_w9432_,
		_w9434_
	);
	LUT2 #(
		.INIT('h1)
	) name8433 (
		_w9370_,
		_w9371_,
		_w9435_
	);
	LUT2 #(
		.INIT('h4)
	) name8434 (
		_w9412_,
		_w9435_,
		_w9436_
	);
	LUT2 #(
		.INIT('h2)
	) name8435 (
		_w9412_,
		_w9435_,
		_w9437_
	);
	LUT2 #(
		.INIT('h1)
	) name8436 (
		_w9436_,
		_w9437_,
		_w9438_
	);
	LUT2 #(
		.INIT('h1)
	) name8437 (
		_w8603_,
		_w8604_,
		_w9439_
	);
	LUT2 #(
		.INIT('h4)
	) name8438 (
		_w8645_,
		_w9439_,
		_w9440_
	);
	LUT2 #(
		.INIT('h2)
	) name8439 (
		_w8645_,
		_w9439_,
		_w9441_
	);
	LUT2 #(
		.INIT('h1)
	) name8440 (
		_w9440_,
		_w9441_,
		_w9442_
	);
	LUT2 #(
		.INIT('h1)
	) name8441 (
		_w9438_,
		_w9442_,
		_w9443_
	);
	LUT2 #(
		.INIT('h8)
	) name8442 (
		_w9438_,
		_w9442_,
		_w9444_
	);
	LUT2 #(
		.INIT('h1)
	) name8443 (
		_w8613_,
		_w8614_,
		_w9445_
	);
	LUT2 #(
		.INIT('h8)
	) name8444 (
		_w8643_,
		_w9445_,
		_w9446_
	);
	LUT2 #(
		.INIT('h1)
	) name8445 (
		_w8643_,
		_w9445_,
		_w9447_
	);
	LUT2 #(
		.INIT('h1)
	) name8446 (
		_w9446_,
		_w9447_,
		_w9448_
	);
	LUT2 #(
		.INIT('h1)
	) name8447 (
		_w9380_,
		_w9381_,
		_w9449_
	);
	LUT2 #(
		.INIT('h8)
	) name8448 (
		_w9410_,
		_w9449_,
		_w9450_
	);
	LUT2 #(
		.INIT('h1)
	) name8449 (
		_w9410_,
		_w9449_,
		_w9451_
	);
	LUT2 #(
		.INIT('h1)
	) name8450 (
		_w9450_,
		_w9451_,
		_w9452_
	);
	LUT2 #(
		.INIT('h1)
	) name8451 (
		_w9448_,
		_w9452_,
		_w9453_
	);
	LUT2 #(
		.INIT('h8)
	) name8452 (
		_w9448_,
		_w9452_,
		_w9454_
	);
	LUT2 #(
		.INIT('h1)
	) name8453 (
		_w9390_,
		_w9391_,
		_w9455_
	);
	LUT2 #(
		.INIT('h4)
	) name8454 (
		_w9408_,
		_w9455_,
		_w9456_
	);
	LUT2 #(
		.INIT('h2)
	) name8455 (
		_w9408_,
		_w9455_,
		_w9457_
	);
	LUT2 #(
		.INIT('h1)
	) name8456 (
		_w9456_,
		_w9457_,
		_w9458_
	);
	LUT2 #(
		.INIT('h1)
	) name8457 (
		_w8623_,
		_w8624_,
		_w9459_
	);
	LUT2 #(
		.INIT('h4)
	) name8458 (
		_w8641_,
		_w9459_,
		_w9460_
	);
	LUT2 #(
		.INIT('h2)
	) name8459 (
		_w8641_,
		_w9459_,
		_w9461_
	);
	LUT2 #(
		.INIT('h1)
	) name8460 (
		_w9460_,
		_w9461_,
		_w9462_
	);
	LUT2 #(
		.INIT('h1)
	) name8461 (
		_w9458_,
		_w9462_,
		_w9463_
	);
	LUT2 #(
		.INIT('h8)
	) name8462 (
		_w9458_,
		_w9462_,
		_w9464_
	);
	LUT2 #(
		.INIT('h1)
	) name8463 (
		_w9393_,
		_w9395_,
		_w9465_
	);
	LUT2 #(
		.INIT('h1)
	) name8464 (
		_w9396_,
		_w9465_,
		_w9466_
	);
	LUT2 #(
		.INIT('h1)
	) name8465 (
		_w8626_,
		_w8628_,
		_w9467_
	);
	LUT2 #(
		.INIT('h1)
	) name8466 (
		_w8629_,
		_w9467_,
		_w9468_
	);
	LUT2 #(
		.INIT('h8)
	) name8467 (
		_w9466_,
		_w9468_,
		_w9469_
	);
	LUT2 #(
		.INIT('h1)
	) name8468 (
		_w8634_,
		_w8635_,
		_w9470_
	);
	LUT2 #(
		.INIT('h4)
	) name8469 (
		_w8639_,
		_w9470_,
		_w9471_
	);
	LUT2 #(
		.INIT('h2)
	) name8470 (
		_w8639_,
		_w9470_,
		_w9472_
	);
	LUT2 #(
		.INIT('h1)
	) name8471 (
		_w9471_,
		_w9472_,
		_w9473_
	);
	LUT2 #(
		.INIT('h2)
	) name8472 (
		_w9469_,
		_w9473_,
		_w9474_
	);
	LUT2 #(
		.INIT('h4)
	) name8473 (
		_w9469_,
		_w9473_,
		_w9475_
	);
	LUT2 #(
		.INIT('h1)
	) name8474 (
		_w9401_,
		_w9402_,
		_w9476_
	);
	LUT2 #(
		.INIT('h4)
	) name8475 (
		_w9406_,
		_w9476_,
		_w9477_
	);
	LUT2 #(
		.INIT('h2)
	) name8476 (
		_w9406_,
		_w9476_,
		_w9478_
	);
	LUT2 #(
		.INIT('h1)
	) name8477 (
		_w9477_,
		_w9478_,
		_w9479_
	);
	LUT2 #(
		.INIT('h1)
	) name8478 (
		_w9475_,
		_w9479_,
		_w9480_
	);
	LUT2 #(
		.INIT('h1)
	) name8479 (
		_w9474_,
		_w9480_,
		_w9481_
	);
	LUT2 #(
		.INIT('h4)
	) name8480 (
		_w9464_,
		_w9481_,
		_w9482_
	);
	LUT2 #(
		.INIT('h1)
	) name8481 (
		_w9463_,
		_w9482_,
		_w9483_
	);
	LUT2 #(
		.INIT('h1)
	) name8482 (
		_w9454_,
		_w9483_,
		_w9484_
	);
	LUT2 #(
		.INIT('h1)
	) name8483 (
		_w9453_,
		_w9484_,
		_w9485_
	);
	LUT2 #(
		.INIT('h1)
	) name8484 (
		_w9444_,
		_w9485_,
		_w9486_
	);
	LUT2 #(
		.INIT('h1)
	) name8485 (
		_w9443_,
		_w9486_,
		_w9487_
	);
	LUT2 #(
		.INIT('h4)
	) name8486 (
		_w9434_,
		_w9487_,
		_w9488_
	);
	LUT2 #(
		.INIT('h1)
	) name8487 (
		_w9433_,
		_w9488_,
		_w9489_
	);
	LUT2 #(
		.INIT('h1)
	) name8488 (
		_w9424_,
		_w9489_,
		_w9490_
	);
	LUT2 #(
		.INIT('h1)
	) name8489 (
		_w9423_,
		_w9490_,
		_w9491_
	);
	LUT2 #(
		.INIT('h1)
	) name8490 (
		_w7888_,
		_w9491_,
		_w9492_
	);
	LUT2 #(
		.INIT('h8)
	) name8491 (
		_w7888_,
		_w9491_,
		_w9493_
	);
	LUT2 #(
		.INIT('h1)
	) name8492 (
		_w9423_,
		_w9424_,
		_w9494_
	);
	LUT2 #(
		.INIT('h4)
	) name8493 (
		_w9489_,
		_w9494_,
		_w9495_
	);
	LUT2 #(
		.INIT('h2)
	) name8494 (
		_w9489_,
		_w9494_,
		_w9496_
	);
	LUT2 #(
		.INIT('h1)
	) name8495 (
		_w9495_,
		_w9496_,
		_w9497_
	);
	LUT2 #(
		.INIT('h1)
	) name8496 (
		_w7820_,
		_w7821_,
		_w9498_
	);
	LUT2 #(
		.INIT('h4)
	) name8497 (
		_w7886_,
		_w9498_,
		_w9499_
	);
	LUT2 #(
		.INIT('h2)
	) name8498 (
		_w7886_,
		_w9498_,
		_w9500_
	);
	LUT2 #(
		.INIT('h1)
	) name8499 (
		_w9499_,
		_w9500_,
		_w9501_
	);
	LUT2 #(
		.INIT('h2)
	) name8500 (
		_w9497_,
		_w9501_,
		_w9502_
	);
	LUT2 #(
		.INIT('h4)
	) name8501 (
		_w9497_,
		_w9501_,
		_w9503_
	);
	LUT2 #(
		.INIT('h1)
	) name8502 (
		_w7830_,
		_w7831_,
		_w9504_
	);
	LUT2 #(
		.INIT('h4)
	) name8503 (
		_w7884_,
		_w9504_,
		_w9505_
	);
	LUT2 #(
		.INIT('h2)
	) name8504 (
		_w7884_,
		_w9504_,
		_w9506_
	);
	LUT2 #(
		.INIT('h1)
	) name8505 (
		_w9505_,
		_w9506_,
		_w9507_
	);
	LUT2 #(
		.INIT('h1)
	) name8506 (
		_w9433_,
		_w9434_,
		_w9508_
	);
	LUT2 #(
		.INIT('h4)
	) name8507 (
		_w9487_,
		_w9508_,
		_w9509_
	);
	LUT2 #(
		.INIT('h2)
	) name8508 (
		_w9487_,
		_w9508_,
		_w9510_
	);
	LUT2 #(
		.INIT('h1)
	) name8509 (
		_w9509_,
		_w9510_,
		_w9511_
	);
	LUT2 #(
		.INIT('h1)
	) name8510 (
		_w9507_,
		_w9511_,
		_w9512_
	);
	LUT2 #(
		.INIT('h8)
	) name8511 (
		_w9507_,
		_w9511_,
		_w9513_
	);
	LUT2 #(
		.INIT('h1)
	) name8512 (
		_w9443_,
		_w9444_,
		_w9514_
	);
	LUT2 #(
		.INIT('h4)
	) name8513 (
		_w9485_,
		_w9514_,
		_w9515_
	);
	LUT2 #(
		.INIT('h2)
	) name8514 (
		_w9485_,
		_w9514_,
		_w9516_
	);
	LUT2 #(
		.INIT('h1)
	) name8515 (
		_w9515_,
		_w9516_,
		_w9517_
	);
	LUT2 #(
		.INIT('h1)
	) name8516 (
		_w7840_,
		_w7841_,
		_w9518_
	);
	LUT2 #(
		.INIT('h4)
	) name8517 (
		_w7882_,
		_w9518_,
		_w9519_
	);
	LUT2 #(
		.INIT('h2)
	) name8518 (
		_w7882_,
		_w9518_,
		_w9520_
	);
	LUT2 #(
		.INIT('h1)
	) name8519 (
		_w9519_,
		_w9520_,
		_w9521_
	);
	LUT2 #(
		.INIT('h1)
	) name8520 (
		_w9517_,
		_w9521_,
		_w9522_
	);
	LUT2 #(
		.INIT('h8)
	) name8521 (
		_w9517_,
		_w9521_,
		_w9523_
	);
	LUT2 #(
		.INIT('h1)
	) name8522 (
		_w7850_,
		_w7851_,
		_w9524_
	);
	LUT2 #(
		.INIT('h4)
	) name8523 (
		_w7880_,
		_w9524_,
		_w9525_
	);
	LUT2 #(
		.INIT('h2)
	) name8524 (
		_w7880_,
		_w9524_,
		_w9526_
	);
	LUT2 #(
		.INIT('h1)
	) name8525 (
		_w9525_,
		_w9526_,
		_w9527_
	);
	LUT2 #(
		.INIT('h1)
	) name8526 (
		_w9453_,
		_w9454_,
		_w9528_
	);
	LUT2 #(
		.INIT('h4)
	) name8527 (
		_w9483_,
		_w9528_,
		_w9529_
	);
	LUT2 #(
		.INIT('h2)
	) name8528 (
		_w9483_,
		_w9528_,
		_w9530_
	);
	LUT2 #(
		.INIT('h1)
	) name8529 (
		_w9529_,
		_w9530_,
		_w9531_
	);
	LUT2 #(
		.INIT('h1)
	) name8530 (
		_w9527_,
		_w9531_,
		_w9532_
	);
	LUT2 #(
		.INIT('h8)
	) name8531 (
		_w9527_,
		_w9531_,
		_w9533_
	);
	LUT2 #(
		.INIT('h1)
	) name8532 (
		_w9463_,
		_w9464_,
		_w9534_
	);
	LUT2 #(
		.INIT('h4)
	) name8533 (
		_w9481_,
		_w9534_,
		_w9535_
	);
	LUT2 #(
		.INIT('h2)
	) name8534 (
		_w9481_,
		_w9534_,
		_w9536_
	);
	LUT2 #(
		.INIT('h1)
	) name8535 (
		_w9535_,
		_w9536_,
		_w9537_
	);
	LUT2 #(
		.INIT('h1)
	) name8536 (
		_w7860_,
		_w7861_,
		_w9538_
	);
	LUT2 #(
		.INIT('h4)
	) name8537 (
		_w7878_,
		_w9538_,
		_w9539_
	);
	LUT2 #(
		.INIT('h2)
	) name8538 (
		_w7878_,
		_w9538_,
		_w9540_
	);
	LUT2 #(
		.INIT('h1)
	) name8539 (
		_w9539_,
		_w9540_,
		_w9541_
	);
	LUT2 #(
		.INIT('h1)
	) name8540 (
		_w9537_,
		_w9541_,
		_w9542_
	);
	LUT2 #(
		.INIT('h8)
	) name8541 (
		_w9537_,
		_w9541_,
		_w9543_
	);
	LUT2 #(
		.INIT('h1)
	) name8542 (
		_w9466_,
		_w9468_,
		_w9544_
	);
	LUT2 #(
		.INIT('h1)
	) name8543 (
		_w9469_,
		_w9544_,
		_w9545_
	);
	LUT2 #(
		.INIT('h1)
	) name8544 (
		_w7863_,
		_w7865_,
		_w9546_
	);
	LUT2 #(
		.INIT('h1)
	) name8545 (
		_w7866_,
		_w9546_,
		_w9547_
	);
	LUT2 #(
		.INIT('h8)
	) name8546 (
		_w9545_,
		_w9547_,
		_w9548_
	);
	LUT2 #(
		.INIT('h1)
	) name8547 (
		_w7871_,
		_w7872_,
		_w9549_
	);
	LUT2 #(
		.INIT('h4)
	) name8548 (
		_w7876_,
		_w9549_,
		_w9550_
	);
	LUT2 #(
		.INIT('h2)
	) name8549 (
		_w7876_,
		_w9549_,
		_w9551_
	);
	LUT2 #(
		.INIT('h1)
	) name8550 (
		_w9550_,
		_w9551_,
		_w9552_
	);
	LUT2 #(
		.INIT('h8)
	) name8551 (
		_w9548_,
		_w9552_,
		_w9553_
	);
	LUT2 #(
		.INIT('h1)
	) name8552 (
		_w9548_,
		_w9552_,
		_w9554_
	);
	LUT2 #(
		.INIT('h1)
	) name8553 (
		_w9474_,
		_w9475_,
		_w9555_
	);
	LUT2 #(
		.INIT('h4)
	) name8554 (
		_w9479_,
		_w9555_,
		_w9556_
	);
	LUT2 #(
		.INIT('h2)
	) name8555 (
		_w9479_,
		_w9555_,
		_w9557_
	);
	LUT2 #(
		.INIT('h1)
	) name8556 (
		_w9556_,
		_w9557_,
		_w9558_
	);
	LUT2 #(
		.INIT('h4)
	) name8557 (
		_w9554_,
		_w9558_,
		_w9559_
	);
	LUT2 #(
		.INIT('h1)
	) name8558 (
		_w9553_,
		_w9559_,
		_w9560_
	);
	LUT2 #(
		.INIT('h4)
	) name8559 (
		_w9543_,
		_w9560_,
		_w9561_
	);
	LUT2 #(
		.INIT('h1)
	) name8560 (
		_w9542_,
		_w9561_,
		_w9562_
	);
	LUT2 #(
		.INIT('h4)
	) name8561 (
		_w9533_,
		_w9562_,
		_w9563_
	);
	LUT2 #(
		.INIT('h1)
	) name8562 (
		_w9532_,
		_w9563_,
		_w9564_
	);
	LUT2 #(
		.INIT('h1)
	) name8563 (
		_w9523_,
		_w9564_,
		_w9565_
	);
	LUT2 #(
		.INIT('h1)
	) name8564 (
		_w9522_,
		_w9565_,
		_w9566_
	);
	LUT2 #(
		.INIT('h1)
	) name8565 (
		_w9513_,
		_w9566_,
		_w9567_
	);
	LUT2 #(
		.INIT('h1)
	) name8566 (
		_w9512_,
		_w9567_,
		_w9568_
	);
	LUT2 #(
		.INIT('h1)
	) name8567 (
		_w9503_,
		_w9568_,
		_w9569_
	);
	LUT2 #(
		.INIT('h1)
	) name8568 (
		_w9502_,
		_w9569_,
		_w9570_
	);
	LUT2 #(
		.INIT('h1)
	) name8569 (
		_w9493_,
		_w9570_,
		_w9571_
	);
	LUT2 #(
		.INIT('h1)
	) name8570 (
		_w9492_,
		_w9571_,
		_w9572_
	);
	LUT2 #(
		.INIT('h8)
	) name8571 (
		_w6307_,
		_w9572_,
		_w9573_
	);
	LUT2 #(
		.INIT('h1)
	) name8572 (
		_w6224_,
		_w6225_,
		_w9574_
	);
	LUT2 #(
		.INIT('h4)
	) name8573 (
		_w6302_,
		_w9574_,
		_w9575_
	);
	LUT2 #(
		.INIT('h2)
	) name8574 (
		_w6302_,
		_w9574_,
		_w9576_
	);
	LUT2 #(
		.INIT('h1)
	) name8575 (
		_w9575_,
		_w9576_,
		_w9577_
	);
	LUT2 #(
		.INIT('h1)
	) name8576 (
		_w9492_,
		_w9493_,
		_w9578_
	);
	LUT2 #(
		.INIT('h4)
	) name8577 (
		_w9570_,
		_w9578_,
		_w9579_
	);
	LUT2 #(
		.INIT('h2)
	) name8578 (
		_w9570_,
		_w9578_,
		_w9580_
	);
	LUT2 #(
		.INIT('h1)
	) name8579 (
		_w9579_,
		_w9580_,
		_w9581_
	);
	LUT2 #(
		.INIT('h2)
	) name8580 (
		_w9577_,
		_w9581_,
		_w9582_
	);
	LUT2 #(
		.INIT('h4)
	) name8581 (
		_w9577_,
		_w9581_,
		_w9583_
	);
	LUT2 #(
		.INIT('h1)
	) name8582 (
		_w6234_,
		_w6235_,
		_w9584_
	);
	LUT2 #(
		.INIT('h4)
	) name8583 (
		_w6300_,
		_w9584_,
		_w9585_
	);
	LUT2 #(
		.INIT('h2)
	) name8584 (
		_w6300_,
		_w9584_,
		_w9586_
	);
	LUT2 #(
		.INIT('h1)
	) name8585 (
		_w9585_,
		_w9586_,
		_w9587_
	);
	LUT2 #(
		.INIT('h1)
	) name8586 (
		_w9502_,
		_w9503_,
		_w9588_
	);
	LUT2 #(
		.INIT('h4)
	) name8587 (
		_w9568_,
		_w9588_,
		_w9589_
	);
	LUT2 #(
		.INIT('h2)
	) name8588 (
		_w9568_,
		_w9588_,
		_w9590_
	);
	LUT2 #(
		.INIT('h1)
	) name8589 (
		_w9589_,
		_w9590_,
		_w9591_
	);
	LUT2 #(
		.INIT('h2)
	) name8590 (
		_w9587_,
		_w9591_,
		_w9592_
	);
	LUT2 #(
		.INIT('h4)
	) name8591 (
		_w9587_,
		_w9591_,
		_w9593_
	);
	LUT2 #(
		.INIT('h1)
	) name8592 (
		_w6244_,
		_w6245_,
		_w9594_
	);
	LUT2 #(
		.INIT('h4)
	) name8593 (
		_w6298_,
		_w9594_,
		_w9595_
	);
	LUT2 #(
		.INIT('h2)
	) name8594 (
		_w6298_,
		_w9594_,
		_w9596_
	);
	LUT2 #(
		.INIT('h1)
	) name8595 (
		_w9595_,
		_w9596_,
		_w9597_
	);
	LUT2 #(
		.INIT('h1)
	) name8596 (
		_w9512_,
		_w9513_,
		_w9598_
	);
	LUT2 #(
		.INIT('h4)
	) name8597 (
		_w9566_,
		_w9598_,
		_w9599_
	);
	LUT2 #(
		.INIT('h2)
	) name8598 (
		_w9566_,
		_w9598_,
		_w9600_
	);
	LUT2 #(
		.INIT('h1)
	) name8599 (
		_w9599_,
		_w9600_,
		_w9601_
	);
	LUT2 #(
		.INIT('h4)
	) name8600 (
		_w9597_,
		_w9601_,
		_w9602_
	);
	LUT2 #(
		.INIT('h2)
	) name8601 (
		_w9597_,
		_w9601_,
		_w9603_
	);
	LUT2 #(
		.INIT('h1)
	) name8602 (
		_w6254_,
		_w6255_,
		_w9604_
	);
	LUT2 #(
		.INIT('h4)
	) name8603 (
		_w6296_,
		_w9604_,
		_w9605_
	);
	LUT2 #(
		.INIT('h2)
	) name8604 (
		_w6296_,
		_w9604_,
		_w9606_
	);
	LUT2 #(
		.INIT('h1)
	) name8605 (
		_w9605_,
		_w9606_,
		_w9607_
	);
	LUT2 #(
		.INIT('h1)
	) name8606 (
		_w9522_,
		_w9523_,
		_w9608_
	);
	LUT2 #(
		.INIT('h4)
	) name8607 (
		_w9564_,
		_w9608_,
		_w9609_
	);
	LUT2 #(
		.INIT('h2)
	) name8608 (
		_w9564_,
		_w9608_,
		_w9610_
	);
	LUT2 #(
		.INIT('h1)
	) name8609 (
		_w9609_,
		_w9610_,
		_w9611_
	);
	LUT2 #(
		.INIT('h1)
	) name8610 (
		_w9607_,
		_w9611_,
		_w9612_
	);
	LUT2 #(
		.INIT('h8)
	) name8611 (
		_w9607_,
		_w9611_,
		_w9613_
	);
	LUT2 #(
		.INIT('h1)
	) name8612 (
		_w6264_,
		_w6265_,
		_w9614_
	);
	LUT2 #(
		.INIT('h8)
	) name8613 (
		_w6294_,
		_w9614_,
		_w9615_
	);
	LUT2 #(
		.INIT('h1)
	) name8614 (
		_w6294_,
		_w9614_,
		_w9616_
	);
	LUT2 #(
		.INIT('h1)
	) name8615 (
		_w9615_,
		_w9616_,
		_w9617_
	);
	LUT2 #(
		.INIT('h1)
	) name8616 (
		_w9532_,
		_w9533_,
		_w9618_
	);
	LUT2 #(
		.INIT('h8)
	) name8617 (
		_w9562_,
		_w9618_,
		_w9619_
	);
	LUT2 #(
		.INIT('h1)
	) name8618 (
		_w9562_,
		_w9618_,
		_w9620_
	);
	LUT2 #(
		.INIT('h1)
	) name8619 (
		_w9619_,
		_w9620_,
		_w9621_
	);
	LUT2 #(
		.INIT('h1)
	) name8620 (
		_w9617_,
		_w9621_,
		_w9622_
	);
	LUT2 #(
		.INIT('h8)
	) name8621 (
		_w9617_,
		_w9621_,
		_w9623_
	);
	LUT2 #(
		.INIT('h1)
	) name8622 (
		_w6274_,
		_w6275_,
		_w9624_
	);
	LUT2 #(
		.INIT('h4)
	) name8623 (
		_w6292_,
		_w9624_,
		_w9625_
	);
	LUT2 #(
		.INIT('h2)
	) name8624 (
		_w6292_,
		_w9624_,
		_w9626_
	);
	LUT2 #(
		.INIT('h1)
	) name8625 (
		_w9625_,
		_w9626_,
		_w9627_
	);
	LUT2 #(
		.INIT('h1)
	) name8626 (
		_w9542_,
		_w9543_,
		_w9628_
	);
	LUT2 #(
		.INIT('h4)
	) name8627 (
		_w9560_,
		_w9628_,
		_w9629_
	);
	LUT2 #(
		.INIT('h2)
	) name8628 (
		_w9560_,
		_w9628_,
		_w9630_
	);
	LUT2 #(
		.INIT('h1)
	) name8629 (
		_w9629_,
		_w9630_,
		_w9631_
	);
	LUT2 #(
		.INIT('h8)
	) name8630 (
		_w9627_,
		_w9631_,
		_w9632_
	);
	LUT2 #(
		.INIT('h1)
	) name8631 (
		_w9627_,
		_w9631_,
		_w9633_
	);
	LUT2 #(
		.INIT('h1)
	) name8632 (
		_w9545_,
		_w9547_,
		_w9634_
	);
	LUT2 #(
		.INIT('h1)
	) name8633 (
		_w9548_,
		_w9634_,
		_w9635_
	);
	LUT2 #(
		.INIT('h1)
	) name8634 (
		_w6277_,
		_w6279_,
		_w9636_
	);
	LUT2 #(
		.INIT('h1)
	) name8635 (
		_w6280_,
		_w9636_,
		_w9637_
	);
	LUT2 #(
		.INIT('h8)
	) name8636 (
		_w9635_,
		_w9637_,
		_w9638_
	);
	LUT2 #(
		.INIT('h1)
	) name8637 (
		_w6285_,
		_w6286_,
		_w9639_
	);
	LUT2 #(
		.INIT('h4)
	) name8638 (
		_w6290_,
		_w9639_,
		_w9640_
	);
	LUT2 #(
		.INIT('h2)
	) name8639 (
		_w6290_,
		_w9639_,
		_w9641_
	);
	LUT2 #(
		.INIT('h1)
	) name8640 (
		_w9640_,
		_w9641_,
		_w9642_
	);
	LUT2 #(
		.INIT('h4)
	) name8641 (
		_w9638_,
		_w9642_,
		_w9643_
	);
	LUT2 #(
		.INIT('h2)
	) name8642 (
		_w9638_,
		_w9642_,
		_w9644_
	);
	LUT2 #(
		.INIT('h1)
	) name8643 (
		_w9553_,
		_w9554_,
		_w9645_
	);
	LUT2 #(
		.INIT('h4)
	) name8644 (
		_w9558_,
		_w9645_,
		_w9646_
	);
	LUT2 #(
		.INIT('h2)
	) name8645 (
		_w9558_,
		_w9645_,
		_w9647_
	);
	LUT2 #(
		.INIT('h1)
	) name8646 (
		_w9646_,
		_w9647_,
		_w9648_
	);
	LUT2 #(
		.INIT('h4)
	) name8647 (
		_w9644_,
		_w9648_,
		_w9649_
	);
	LUT2 #(
		.INIT('h1)
	) name8648 (
		_w9643_,
		_w9649_,
		_w9650_
	);
	LUT2 #(
		.INIT('h4)
	) name8649 (
		_w9633_,
		_w9650_,
		_w9651_
	);
	LUT2 #(
		.INIT('h1)
	) name8650 (
		_w9632_,
		_w9651_,
		_w9652_
	);
	LUT2 #(
		.INIT('h4)
	) name8651 (
		_w9623_,
		_w9652_,
		_w9653_
	);
	LUT2 #(
		.INIT('h1)
	) name8652 (
		_w9622_,
		_w9653_,
		_w9654_
	);
	LUT2 #(
		.INIT('h1)
	) name8653 (
		_w9613_,
		_w9654_,
		_w9655_
	);
	LUT2 #(
		.INIT('h1)
	) name8654 (
		_w9612_,
		_w9655_,
		_w9656_
	);
	LUT2 #(
		.INIT('h4)
	) name8655 (
		_w9603_,
		_w9656_,
		_w9657_
	);
	LUT2 #(
		.INIT('h1)
	) name8656 (
		_w9602_,
		_w9657_,
		_w9658_
	);
	LUT2 #(
		.INIT('h4)
	) name8657 (
		_w9593_,
		_w9658_,
		_w9659_
	);
	LUT2 #(
		.INIT('h1)
	) name8658 (
		_w9592_,
		_w9659_,
		_w9660_
	);
	LUT2 #(
		.INIT('h1)
	) name8659 (
		_w9583_,
		_w9660_,
		_w9661_
	);
	LUT2 #(
		.INIT('h1)
	) name8660 (
		_w9582_,
		_w9661_,
		_w9662_
	);
	LUT2 #(
		.INIT('h2)
	) name8661 (
		_w9573_,
		_w9662_,
		_w9663_
	);
	LUT2 #(
		.INIT('h1)
	) name8662 (
		_w9612_,
		_w9613_,
		_w9664_
	);
	LUT2 #(
		.INIT('h2)
	) name8663 (
		_w9654_,
		_w9664_,
		_w9665_
	);
	LUT2 #(
		.INIT('h4)
	) name8664 (
		_w9654_,
		_w9664_,
		_w9666_
	);
	LUT2 #(
		.INIT('h1)
	) name8665 (
		_w9665_,
		_w9666_,
		_w9667_
	);
	LUT2 #(
		.INIT('h1)
	) name8666 (
		_w9592_,
		_w9593_,
		_w9668_
	);
	LUT2 #(
		.INIT('h2)
	) name8667 (
		_w9658_,
		_w9668_,
		_w9669_
	);
	LUT2 #(
		.INIT('h4)
	) name8668 (
		_w9658_,
		_w9668_,
		_w9670_
	);
	LUT2 #(
		.INIT('h1)
	) name8669 (
		_w9602_,
		_w9603_,
		_w9671_
	);
	LUT2 #(
		.INIT('h8)
	) name8670 (
		_w9656_,
		_w9671_,
		_w9672_
	);
	LUT2 #(
		.INIT('h1)
	) name8671 (
		_w9656_,
		_w9671_,
		_w9673_
	);
	LUT2 #(
		.INIT('h1)
	) name8672 (
		_w9632_,
		_w9633_,
		_w9674_
	);
	LUT2 #(
		.INIT('h1)
	) name8673 (
		_w9650_,
		_w9674_,
		_w9675_
	);
	LUT2 #(
		.INIT('h4)
	) name8674 (
		_w9643_,
		_w9649_,
		_w9676_
	);
	LUT2 #(
		.INIT('h1)
	) name8675 (
		_w9643_,
		_w9644_,
		_w9677_
	);
	LUT2 #(
		.INIT('h1)
	) name8676 (
		_w9648_,
		_w9677_,
		_w9678_
	);
	LUT2 #(
		.INIT('h1)
	) name8677 (
		_w9635_,
		_w9637_,
		_w9679_
	);
	LUT2 #(
		.INIT('h1)
	) name8678 (
		_w9638_,
		_w9679_,
		_w9680_
	);
	LUT2 #(
		.INIT('h1)
	) name8679 (
		\A[1000] ,
		_w9680_,
		_w9681_
	);
	LUT2 #(
		.INIT('h4)
	) name8680 (
		_w9676_,
		_w9681_,
		_w9682_
	);
	LUT2 #(
		.INIT('h4)
	) name8681 (
		_w9678_,
		_w9682_,
		_w9683_
	);
	LUT2 #(
		.INIT('h4)
	) name8682 (
		_w9632_,
		_w9651_,
		_w9684_
	);
	LUT2 #(
		.INIT('h1)
	) name8683 (
		_w9675_,
		_w9683_,
		_w9685_
	);
	LUT2 #(
		.INIT('h4)
	) name8684 (
		_w9684_,
		_w9685_,
		_w9686_
	);
	LUT2 #(
		.INIT('h1)
	) name8685 (
		_w9622_,
		_w9623_,
		_w9687_
	);
	LUT2 #(
		.INIT('h1)
	) name8686 (
		_w9652_,
		_w9687_,
		_w9688_
	);
	LUT2 #(
		.INIT('h8)
	) name8687 (
		_w9652_,
		_w9687_,
		_w9689_
	);
	LUT2 #(
		.INIT('h1)
	) name8688 (
		_w9686_,
		_w9688_,
		_w9690_
	);
	LUT2 #(
		.INIT('h4)
	) name8689 (
		_w9689_,
		_w9690_,
		_w9691_
	);
	LUT2 #(
		.INIT('h1)
	) name8690 (
		_w9582_,
		_w9583_,
		_w9692_
	);
	LUT2 #(
		.INIT('h4)
	) name8691 (
		_w9660_,
		_w9692_,
		_w9693_
	);
	LUT2 #(
		.INIT('h2)
	) name8692 (
		_w9660_,
		_w9692_,
		_w9694_
	);
	LUT2 #(
		.INIT('h1)
	) name8693 (
		_w9693_,
		_w9694_,
		_w9695_
	);
	LUT2 #(
		.INIT('h1)
	) name8694 (
		_w9667_,
		_w9691_,
		_w9696_
	);
	LUT2 #(
		.INIT('h4)
	) name8695 (
		_w9672_,
		_w9696_,
		_w9697_
	);
	LUT2 #(
		.INIT('h4)
	) name8696 (
		_w9673_,
		_w9697_,
		_w9698_
	);
	LUT2 #(
		.INIT('h4)
	) name8697 (
		_w9669_,
		_w9698_,
		_w9699_
	);
	LUT2 #(
		.INIT('h4)
	) name8698 (
		_w9670_,
		_w9699_,
		_w9700_
	);
	LUT2 #(
		.INIT('h4)
	) name8699 (
		_w9695_,
		_w9700_,
		_w9701_
	);
	LUT2 #(
		.INIT('h4)
	) name8700 (
		_w9663_,
		_w9701_,
		_w9702_
	);
	LUT2 #(
		.INIT('h4)
	) name8701 (
		_w9573_,
		_w9662_,
		_w9703_
	);
	LUT2 #(
		.INIT('h4)
	) name8702 (
		_w6213_,
		_w6304_,
		_w9704_
	);
	LUT2 #(
		.INIT('h1)
	) name8703 (
		_w6307_,
		_w9572_,
		_w9705_
	);
	LUT2 #(
		.INIT('h1)
	) name8704 (
		_w6214_,
		_w9704_,
		_w9706_
	);
	LUT2 #(
		.INIT('h4)
	) name8705 (
		_w9705_,
		_w9706_,
		_w9707_
	);
	LUT2 #(
		.INIT('h4)
	) name8706 (
		_w9703_,
		_w9707_,
		_w9708_
	);
	LUT2 #(
		.INIT('h4)
	) name8707 (
		_w9702_,
		_w9708_,
		_w9709_
	);
	assign maj = _w9709_ ;
endmodule;