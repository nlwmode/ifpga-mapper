module top( \addroundkey_ready_o_reg/NET0131  , \addroundkey_round_reg[0]/NET0131  , \addroundkey_round_reg[1]/NET0131  , \addroundkey_round_reg[2]/NET0131  , \addroundkey_round_reg[3]/NET0131  , \addroundkey_start_i_reg/NET0131  , \data_i[0]_pad  , \data_i[100]_pad  , \data_i[101]_pad  , \data_i[102]_pad  , \data_i[103]_pad  , \data_i[104]_pad  , \data_i[105]_pad  , \data_i[106]_pad  , \data_i[107]_pad  , \data_i[108]_pad  , \data_i[109]_pad  , \data_i[10]_pad  , \data_i[110]_pad  , \data_i[111]_pad  , \data_i[112]_pad  , \data_i[113]_pad  , \data_i[114]_pad  , \data_i[115]_pad  , \data_i[116]_pad  , \data_i[117]_pad  , \data_i[118]_pad  , \data_i[119]_pad  , \data_i[11]_pad  , \data_i[120]_pad  , \data_i[121]_pad  , \data_i[122]_pad  , \data_i[123]_pad  , \data_i[124]_pad  , \data_i[125]_pad  , \data_i[126]_pad  , \data_i[127]_pad  , \data_i[12]_pad  , \data_i[13]_pad  , \data_i[14]_pad  , \data_i[15]_pad  , \data_i[16]_pad  , \data_i[17]_pad  , \data_i[18]_pad  , \data_i[19]_pad  , \data_i[1]_pad  , \data_i[20]_pad  , \data_i[21]_pad  , \data_i[22]_pad  , \data_i[23]_pad  , \data_i[24]_pad  , \data_i[25]_pad  , \data_i[26]_pad  , \data_i[27]_pad  , \data_i[28]_pad  , \data_i[29]_pad  , \data_i[2]_pad  , \data_i[30]_pad  , \data_i[31]_pad  , \data_i[32]_pad  , \data_i[33]_pad  , \data_i[34]_pad  , \data_i[35]_pad  , \data_i[36]_pad  , \data_i[37]_pad  , \data_i[38]_pad  , \data_i[39]_pad  , \data_i[3]_pad  , \data_i[40]_pad  , \data_i[41]_pad  , \data_i[42]_pad  , \data_i[43]_pad  , \data_i[44]_pad  , \data_i[45]_pad  , \data_i[46]_pad  , \data_i[47]_pad  , \data_i[48]_pad  , \data_i[49]_pad  , \data_i[4]_pad  , \data_i[50]_pad  , \data_i[51]_pad  , \data_i[52]_pad  , \data_i[53]_pad  , \data_i[54]_pad  , \data_i[55]_pad  , \data_i[56]_pad  , \data_i[57]_pad  , \data_i[58]_pad  , \data_i[59]_pad  , \data_i[5]_pad  , \data_i[60]_pad  , \data_i[61]_pad  , \data_i[62]_pad  , \data_i[63]_pad  , \data_i[64]_pad  , \data_i[65]_pad  , \data_i[66]_pad  , \data_i[67]_pad  , \data_i[68]_pad  , \data_i[69]_pad  , \data_i[6]_pad  , \data_i[70]_pad  , \data_i[71]_pad  , \data_i[72]_pad  , \data_i[73]_pad  , \data_i[74]_pad  , \data_i[75]_pad  , \data_i[76]_pad  , \data_i[77]_pad  , \data_i[78]_pad  , \data_i[79]_pad  , \data_i[7]_pad  , \data_i[80]_pad  , \data_i[81]_pad  , \data_i[82]_pad  , \data_i[83]_pad  , \data_i[84]_pad  , \data_i[85]_pad  , \data_i[86]_pad  , \data_i[87]_pad  , \data_i[88]_pad  , \data_i[89]_pad  , \data_i[8]_pad  , \data_i[90]_pad  , \data_i[91]_pad  , \data_i[92]_pad  , \data_i[93]_pad  , \data_i[94]_pad  , \data_i[95]_pad  , \data_i[96]_pad  , \data_i[97]_pad  , \data_i[98]_pad  , \data_i[99]_pad  , \data_i[9]_pad  , \data_o[0]_pad  , \data_o[100]_pad  , \data_o[101]_pad  , \data_o[102]_pad  , \data_o[103]_pad  , \data_o[104]_pad  , \data_o[105]_pad  , \data_o[106]_pad  , \data_o[107]_pad  , \data_o[108]_pad  , \data_o[109]_pad  , \data_o[10]_pad  , \data_o[110]_pad  , \data_o[111]_pad  , \data_o[112]_pad  , \data_o[113]_pad  , \data_o[114]_pad  , \data_o[115]_pad  , \data_o[116]_pad  , \data_o[117]_pad  , \data_o[118]_pad  , \data_o[119]_pad  , \data_o[11]_pad  , \data_o[120]_pad  , \data_o[121]_pad  , \data_o[122]_pad  , \data_o[123]_pad  , \data_o[124]_pad  , \data_o[125]_pad  , \data_o[126]_pad  , \data_o[127]_pad  , \data_o[12]_pad  , \data_o[13]_pad  , \data_o[14]_pad  , \data_o[15]_pad  , \data_o[16]_pad  , \data_o[17]_pad  , \data_o[18]_pad  , \data_o[19]_pad  , \data_o[1]_pad  , \data_o[20]_pad  , \data_o[21]_pad  , \data_o[22]_pad  , \data_o[23]_pad  , \data_o[24]_pad  , \data_o[25]_pad  , \data_o[26]_pad  , \data_o[27]_pad  , \data_o[28]_pad  , \data_o[29]_pad  , \data_o[2]_pad  , \data_o[30]_pad  , \data_o[31]_pad  , \data_o[32]_pad  , \data_o[33]_pad  , \data_o[34]_pad  , \data_o[35]_pad  , \data_o[36]_pad  , \data_o[37]_pad  , \data_o[38]_pad  , \data_o[39]_pad  , \data_o[3]_pad  , \data_o[40]_pad  , \data_o[41]_pad  , \data_o[42]_pad  , \data_o[43]_pad  , \data_o[44]_pad  , \data_o[45]_pad  , \data_o[46]_pad  , \data_o[47]_pad  , \data_o[48]_pad  , \data_o[49]_pad  , \data_o[4]_pad  , \data_o[50]_pad  , \data_o[51]_pad  , \data_o[52]_pad  , \data_o[53]_pad  , \data_o[54]_pad  , \data_o[55]_pad  , \data_o[56]_pad  , \data_o[57]_pad  , \data_o[58]_pad  , \data_o[59]_pad  , \data_o[5]_pad  , \data_o[60]_pad  , \data_o[61]_pad  , \data_o[62]_pad  , \data_o[63]_pad  , \data_o[64]_pad  , \data_o[65]_pad  , \data_o[66]_pad  , \data_o[67]_pad  , \data_o[68]_pad  , \data_o[69]_pad  , \data_o[6]_pad  , \data_o[70]_pad  , \data_o[71]_pad  , \data_o[72]_pad  , \data_o[73]_pad  , \data_o[74]_pad  , \data_o[75]_pad  , \data_o[76]_pad  , \data_o[77]_pad  , \data_o[78]_pad  , \data_o[79]_pad  , \data_o[7]_pad  , \data_o[80]_pad  , \data_o[81]_pad  , \data_o[82]_pad  , \data_o[83]_pad  , \data_o[84]_pad  , \data_o[85]_pad  , \data_o[86]_pad  , \data_o[87]_pad  , \data_o[88]_pad  , \data_o[89]_pad  , \data_o[8]_pad  , \data_o[90]_pad  , \data_o[91]_pad  , \data_o[92]_pad  , \data_o[93]_pad  , \data_o[94]_pad  , \data_o[95]_pad  , \data_o[96]_pad  , \data_o[97]_pad  , \data_o[98]_pad  , \data_o[99]_pad  , \data_o[9]_pad  , decrypt_i_pad , \first_round_reg_reg/NET0131  , \key_i[0]_pad  , \key_i[100]_pad  , \key_i[101]_pad  , \key_i[102]_pad  , \key_i[103]_pad  , \key_i[104]_pad  , \key_i[105]_pad  , \key_i[106]_pad  , \key_i[107]_pad  , \key_i[108]_pad  , \key_i[109]_pad  , \key_i[10]_pad  , \key_i[110]_pad  , \key_i[111]_pad  , \key_i[112]_pad  , \key_i[113]_pad  , \key_i[114]_pad  , \key_i[115]_pad  , \key_i[116]_pad  , \key_i[117]_pad  , \key_i[118]_pad  , \key_i[119]_pad  , \key_i[11]_pad  , \key_i[120]_pad  , \key_i[121]_pad  , \key_i[122]_pad  , \key_i[123]_pad  , \key_i[124]_pad  , \key_i[125]_pad  , \key_i[126]_pad  , \key_i[127]_pad  , \key_i[12]_pad  , \key_i[13]_pad  , \key_i[14]_pad  , \key_i[15]_pad  , \key_i[16]_pad  , \key_i[17]_pad  , \key_i[18]_pad  , \key_i[19]_pad  , \key_i[1]_pad  , \key_i[20]_pad  , \key_i[21]_pad  , \key_i[22]_pad  , \key_i[23]_pad  , \key_i[24]_pad  , \key_i[25]_pad  , \key_i[26]_pad  , \key_i[27]_pad  , \key_i[28]_pad  , \key_i[29]_pad  , \key_i[2]_pad  , \key_i[30]_pad  , \key_i[31]_pad  , \key_i[32]_pad  , \key_i[33]_pad  , \key_i[34]_pad  , \key_i[35]_pad  , \key_i[36]_pad  , \key_i[37]_pad  , \key_i[38]_pad  , \key_i[39]_pad  , \key_i[3]_pad  , \key_i[40]_pad  , \key_i[41]_pad  , \key_i[42]_pad  , \key_i[43]_pad  , \key_i[44]_pad  , \key_i[45]_pad  , \key_i[46]_pad  , \key_i[47]_pad  , \key_i[48]_pad  , \key_i[49]_pad  , \key_i[4]_pad  , \key_i[50]_pad  , \key_i[51]_pad  , \key_i[52]_pad  , \key_i[53]_pad  , \key_i[54]_pad  , \key_i[55]_pad  , \key_i[56]_pad  , \key_i[57]_pad  , \key_i[58]_pad  , \key_i[59]_pad  , \key_i[5]_pad  , \key_i[60]_pad  , \key_i[61]_pad  , \key_i[62]_pad  , \key_i[63]_pad  , \key_i[64]_pad  , \key_i[65]_pad  , \key_i[66]_pad  , \key_i[67]_pad  , \key_i[68]_pad  , \key_i[69]_pad  , \key_i[6]_pad  , \key_i[70]_pad  , \key_i[71]_pad  , \key_i[72]_pad  , \key_i[73]_pad  , \key_i[74]_pad  , \key_i[75]_pad  , \key_i[76]_pad  , \key_i[77]_pad  , \key_i[78]_pad  , \key_i[79]_pad  , \key_i[7]_pad  , \key_i[80]_pad  , \key_i[81]_pad  , \key_i[82]_pad  , \key_i[83]_pad  , \key_i[84]_pad  , \key_i[85]_pad  , \key_i[86]_pad  , \key_i[87]_pad  , \key_i[88]_pad  , \key_i[89]_pad  , \key_i[8]_pad  , \key_i[90]_pad  , \key_i[91]_pad  , \key_i[92]_pad  , \key_i[93]_pad  , \key_i[94]_pad  , \key_i[95]_pad  , \key_i[96]_pad  , \key_i[97]_pad  , \key_i[98]_pad  , \key_i[99]_pad  , \key_i[9]_pad  , \ks1_col_reg[0]/NET0131  , \ks1_col_reg[16]/NET0131  , \ks1_col_reg[17]/NET0131  , \ks1_col_reg[18]/NET0131  , \ks1_col_reg[19]/NET0131  , \ks1_col_reg[1]/NET0131  , \ks1_col_reg[20]/NET0131  , \ks1_col_reg[21]/NET0131  , \ks1_col_reg[22]/NET0131  , \ks1_col_reg[23]/NET0131  , \ks1_col_reg[24]/NET0131  , \ks1_col_reg[25]/NET0131  , \ks1_col_reg[26]/NET0131  , \ks1_col_reg[27]/NET0131  , \ks1_col_reg[28]/NET0131  , \ks1_col_reg[29]/NET0131  , \ks1_col_reg[2]/NET0131  , \ks1_col_reg[30]/NET0131  , \ks1_col_reg[31]/NET0131  , \ks1_col_reg[3]/NET0131  , \ks1_col_reg[4]/NET0131  , \ks1_col_reg[5]/NET0131  , \ks1_col_reg[6]/NET0131  , \ks1_col_reg[7]/NET0131  , \ks1_key_reg_reg[0]/NET0131  , \ks1_key_reg_reg[100]/NET0131  , \ks1_key_reg_reg[101]/NET0131  , \ks1_key_reg_reg[102]/NET0131  , \ks1_key_reg_reg[103]/NET0131  , \ks1_key_reg_reg[104]/NET0131  , \ks1_key_reg_reg[105]/NET0131  , \ks1_key_reg_reg[106]/NET0131  , \ks1_key_reg_reg[107]/NET0131  , \ks1_key_reg_reg[108]/NET0131  , \ks1_key_reg_reg[109]/P0002  , \ks1_key_reg_reg[10]/NET0131  , \ks1_key_reg_reg[110]/P0002  , \ks1_key_reg_reg[111]/NET0131  , \ks1_key_reg_reg[112]/NET0131  , \ks1_key_reg_reg[113]/NET0131  , \ks1_key_reg_reg[114]/NET0131  , \ks1_key_reg_reg[115]/NET0131  , \ks1_key_reg_reg[116]/NET0131  , \ks1_key_reg_reg[117]/NET0131  , \ks1_key_reg_reg[118]/NET0131  , \ks1_key_reg_reg[119]/NET0131  , \ks1_key_reg_reg[11]/NET0131  , \ks1_key_reg_reg[120]/NET0131  , \ks1_key_reg_reg[121]/NET0131  , \ks1_key_reg_reg[122]/NET0131  , \ks1_key_reg_reg[123]/NET0131  , \ks1_key_reg_reg[124]/NET0131  , \ks1_key_reg_reg[125]/NET0131  , \ks1_key_reg_reg[126]/NET0131  , \ks1_key_reg_reg[127]/NET0131  , \ks1_key_reg_reg[12]/NET0131  , \ks1_key_reg_reg[13]/NET0131  , \ks1_key_reg_reg[14]/NET0131  , \ks1_key_reg_reg[15]/NET0131  , \ks1_key_reg_reg[16]/NET0131  , \ks1_key_reg_reg[17]/NET0131  , \ks1_key_reg_reg[18]/NET0131  , \ks1_key_reg_reg[19]/NET0131  , \ks1_key_reg_reg[1]/NET0131  , \ks1_key_reg_reg[20]/NET0131  , \ks1_key_reg_reg[21]/NET0131  , \ks1_key_reg_reg[22]/NET0131  , \ks1_key_reg_reg[23]/NET0131  , \ks1_key_reg_reg[24]/NET0131  , \ks1_key_reg_reg[25]/NET0131  , \ks1_key_reg_reg[26]/NET0131  , \ks1_key_reg_reg[27]/NET0131  , \ks1_key_reg_reg[28]/NET0131  , \ks1_key_reg_reg[29]/NET0131  , \ks1_key_reg_reg[2]/NET0131  , \ks1_key_reg_reg[30]/NET0131  , \ks1_key_reg_reg[31]/NET0131  , \ks1_key_reg_reg[32]/NET0131  , \ks1_key_reg_reg[33]/NET0131  , \ks1_key_reg_reg[34]/NET0131  , \ks1_key_reg_reg[35]/NET0131  , \ks1_key_reg_reg[36]/NET0131  , \ks1_key_reg_reg[37]/NET0131  , \ks1_key_reg_reg[38]/NET0131  , \ks1_key_reg_reg[39]/NET0131  , \ks1_key_reg_reg[3]/NET0131  , \ks1_key_reg_reg[40]/P0002  , \ks1_key_reg_reg[41]/P0002  , \ks1_key_reg_reg[42]/P0002  , \ks1_key_reg_reg[43]/P0002  , \ks1_key_reg_reg[44]/P0002  , \ks1_key_reg_reg[45]/P0002  , \ks1_key_reg_reg[46]/P0002  , \ks1_key_reg_reg[47]/P0002  , \ks1_key_reg_reg[48]/NET0131  , \ks1_key_reg_reg[49]/NET0131  , \ks1_key_reg_reg[4]/NET0131  , \ks1_key_reg_reg[50]/NET0131  , \ks1_key_reg_reg[51]/NET0131  , \ks1_key_reg_reg[52]/NET0131  , \ks1_key_reg_reg[53]/NET0131  , \ks1_key_reg_reg[54]/NET0131  , \ks1_key_reg_reg[55]/NET0131  , \ks1_key_reg_reg[56]/NET0131  , \ks1_key_reg_reg[57]/NET0131  , \ks1_key_reg_reg[58]/NET0131  , \ks1_key_reg_reg[59]/NET0131  , \ks1_key_reg_reg[5]/NET0131  , \ks1_key_reg_reg[60]/NET0131  , \ks1_key_reg_reg[61]/NET0131  , \ks1_key_reg_reg[62]/NET0131  , \ks1_key_reg_reg[63]/NET0131  , \ks1_key_reg_reg[64]/NET0131  , \ks1_key_reg_reg[65]/NET0131  , \ks1_key_reg_reg[66]/NET0131  , \ks1_key_reg_reg[67]/NET0131  , \ks1_key_reg_reg[68]/NET0131  , \ks1_key_reg_reg[69]/NET0131  , \ks1_key_reg_reg[6]/NET0131  , \ks1_key_reg_reg[70]/NET0131  , \ks1_key_reg_reg[71]/NET0131  , \ks1_key_reg_reg[72]/P0002  , \ks1_key_reg_reg[73]/NET0131  , \ks1_key_reg_reg[74]/NET0131  , \ks1_key_reg_reg[75]/P0002  , \ks1_key_reg_reg[76]/P0002  , \ks1_key_reg_reg[77]/P0002  , \ks1_key_reg_reg[78]/P0002  , \ks1_key_reg_reg[79]/P0002  , \ks1_key_reg_reg[7]/NET0131  , \ks1_key_reg_reg[80]/NET0131  , \ks1_key_reg_reg[81]/NET0131  , \ks1_key_reg_reg[82]/NET0131  , \ks1_key_reg_reg[83]/NET0131  , \ks1_key_reg_reg[84]/NET0131  , \ks1_key_reg_reg[85]/NET0131  , \ks1_key_reg_reg[86]/NET0131  , \ks1_key_reg_reg[87]/NET0131  , \ks1_key_reg_reg[88]/NET0131  , \ks1_key_reg_reg[89]/NET0131  , \ks1_key_reg_reg[8]/NET0131  , \ks1_key_reg_reg[90]/NET0131  , \ks1_key_reg_reg[91]/NET0131  , \ks1_key_reg_reg[92]/NET0131  , \ks1_key_reg_reg[93]/NET0131  , \ks1_key_reg_reg[94]/NET0131  , \ks1_key_reg_reg[95]/NET0131  , \ks1_key_reg_reg[96]/NET0131  , \ks1_key_reg_reg[97]/NET0131  , \ks1_key_reg_reg[98]/NET0131  , \ks1_key_reg_reg[99]/NET0131  , \ks1_key_reg_reg[9]/NET0131  , \ks1_ready_o_reg/NET0131  , \ks1_state_reg[0]/NET0131  , \ks1_state_reg[1]/NET0131  , \ks1_state_reg[2]/NET0131  , load_i_pad , \mix1_data_o_reg_reg[0]/NET0131  , \mix1_data_o_reg_reg[100]/NET0131  , \mix1_data_o_reg_reg[101]/NET0131  , \mix1_data_o_reg_reg[102]/NET0131  , \mix1_data_o_reg_reg[103]/NET0131  , \mix1_data_o_reg_reg[104]/NET0131  , \mix1_data_o_reg_reg[105]/NET0131  , \mix1_data_o_reg_reg[106]/NET0131  , \mix1_data_o_reg_reg[107]/NET0131  , \mix1_data_o_reg_reg[108]/NET0131  , \mix1_data_o_reg_reg[109]/NET0131  , \mix1_data_o_reg_reg[10]/NET0131  , \mix1_data_o_reg_reg[110]/NET0131  , \mix1_data_o_reg_reg[111]/NET0131  , \mix1_data_o_reg_reg[112]/NET0131  , \mix1_data_o_reg_reg[113]/NET0131  , \mix1_data_o_reg_reg[114]/NET0131  , \mix1_data_o_reg_reg[115]/NET0131  , \mix1_data_o_reg_reg[116]/NET0131  , \mix1_data_o_reg_reg[117]/NET0131  , \mix1_data_o_reg_reg[118]/NET0131  , \mix1_data_o_reg_reg[119]/NET0131  , \mix1_data_o_reg_reg[11]/NET0131  , \mix1_data_o_reg_reg[120]/NET0131  , \mix1_data_o_reg_reg[121]/NET0131  , \mix1_data_o_reg_reg[122]/NET0131  , \mix1_data_o_reg_reg[123]/NET0131  , \mix1_data_o_reg_reg[124]/NET0131  , \mix1_data_o_reg_reg[125]/NET0131  , \mix1_data_o_reg_reg[126]/NET0131  , \mix1_data_o_reg_reg[127]/NET0131  , \mix1_data_o_reg_reg[12]/NET0131  , \mix1_data_o_reg_reg[13]/NET0131  , \mix1_data_o_reg_reg[14]/NET0131  , \mix1_data_o_reg_reg[15]/NET0131  , \mix1_data_o_reg_reg[16]/NET0131  , \mix1_data_o_reg_reg[17]/NET0131  , \mix1_data_o_reg_reg[18]/NET0131  , \mix1_data_o_reg_reg[19]/NET0131  , \mix1_data_o_reg_reg[1]/NET0131  , \mix1_data_o_reg_reg[20]/NET0131  , \mix1_data_o_reg_reg[21]/NET0131  , \mix1_data_o_reg_reg[22]/NET0131  , \mix1_data_o_reg_reg[23]/NET0131  , \mix1_data_o_reg_reg[24]/NET0131  , \mix1_data_o_reg_reg[25]/NET0131  , \mix1_data_o_reg_reg[26]/NET0131  , \mix1_data_o_reg_reg[27]/NET0131  , \mix1_data_o_reg_reg[28]/NET0131  , \mix1_data_o_reg_reg[29]/NET0131  , \mix1_data_o_reg_reg[2]/NET0131  , \mix1_data_o_reg_reg[30]/NET0131  , \mix1_data_o_reg_reg[31]/NET0131  , \mix1_data_o_reg_reg[32]/NET0131  , \mix1_data_o_reg_reg[33]/NET0131  , \mix1_data_o_reg_reg[34]/NET0131  , \mix1_data_o_reg_reg[35]/NET0131  , \mix1_data_o_reg_reg[36]/NET0131  , \mix1_data_o_reg_reg[37]/NET0131  , \mix1_data_o_reg_reg[38]/NET0131  , \mix1_data_o_reg_reg[39]/NET0131  , \mix1_data_o_reg_reg[3]/NET0131  , \mix1_data_o_reg_reg[40]/NET0131  , \mix1_data_o_reg_reg[41]/NET0131  , \mix1_data_o_reg_reg[42]/NET0131  , \mix1_data_o_reg_reg[43]/NET0131  , \mix1_data_o_reg_reg[44]/NET0131  , \mix1_data_o_reg_reg[45]/NET0131  , \mix1_data_o_reg_reg[46]/NET0131  , \mix1_data_o_reg_reg[47]/NET0131  , \mix1_data_o_reg_reg[48]/NET0131  , \mix1_data_o_reg_reg[49]/NET0131  , \mix1_data_o_reg_reg[4]/NET0131  , \mix1_data_o_reg_reg[50]/NET0131  , \mix1_data_o_reg_reg[51]/NET0131  , \mix1_data_o_reg_reg[52]/NET0131  , \mix1_data_o_reg_reg[53]/NET0131  , \mix1_data_o_reg_reg[54]/NET0131  , \mix1_data_o_reg_reg[55]/NET0131  , \mix1_data_o_reg_reg[56]/NET0131  , \mix1_data_o_reg_reg[57]/NET0131  , \mix1_data_o_reg_reg[58]/NET0131  , \mix1_data_o_reg_reg[59]/NET0131  , \mix1_data_o_reg_reg[5]/NET0131  , \mix1_data_o_reg_reg[60]/NET0131  , \mix1_data_o_reg_reg[61]/NET0131  , \mix1_data_o_reg_reg[62]/NET0131  , \mix1_data_o_reg_reg[63]/NET0131  , \mix1_data_o_reg_reg[64]/NET0131  , \mix1_data_o_reg_reg[65]/NET0131  , \mix1_data_o_reg_reg[66]/NET0131  , \mix1_data_o_reg_reg[67]/NET0131  , \mix1_data_o_reg_reg[68]/NET0131  , \mix1_data_o_reg_reg[69]/NET0131  , \mix1_data_o_reg_reg[6]/NET0131  , \mix1_data_o_reg_reg[70]/NET0131  , \mix1_data_o_reg_reg[71]/NET0131  , \mix1_data_o_reg_reg[72]/NET0131  , \mix1_data_o_reg_reg[73]/NET0131  , \mix1_data_o_reg_reg[74]/NET0131  , \mix1_data_o_reg_reg[75]/NET0131  , \mix1_data_o_reg_reg[76]/NET0131  , \mix1_data_o_reg_reg[77]/NET0131  , \mix1_data_o_reg_reg[78]/NET0131  , \mix1_data_o_reg_reg[79]/NET0131  , \mix1_data_o_reg_reg[7]/NET0131  , \mix1_data_o_reg_reg[80]/NET0131  , \mix1_data_o_reg_reg[81]/NET0131  , \mix1_data_o_reg_reg[82]/NET0131  , \mix1_data_o_reg_reg[83]/NET0131  , \mix1_data_o_reg_reg[84]/NET0131  , \mix1_data_o_reg_reg[85]/NET0131  , \mix1_data_o_reg_reg[86]/NET0131  , \mix1_data_o_reg_reg[87]/NET0131  , \mix1_data_o_reg_reg[88]/NET0131  , \mix1_data_o_reg_reg[89]/NET0131  , \mix1_data_o_reg_reg[8]/NET0131  , \mix1_data_o_reg_reg[90]/NET0131  , \mix1_data_o_reg_reg[91]/NET0131  , \mix1_data_o_reg_reg[92]/NET0131  , \mix1_data_o_reg_reg[93]/NET0131  , \mix1_data_o_reg_reg[94]/NET0131  , \mix1_data_o_reg_reg[95]/NET0131  , \mix1_data_o_reg_reg[96]/NET0131  , \mix1_data_o_reg_reg[97]/NET0131  , \mix1_data_o_reg_reg[98]/NET0131  , \mix1_data_o_reg_reg[99]/NET0131  , \mix1_data_o_reg_reg[9]/NET0131  , \mix1_data_reg_reg[100]/NET0131  , \mix1_data_reg_reg[101]/NET0131  , \mix1_data_reg_reg[102]/NET0131  , \mix1_data_reg_reg[103]/NET0131  , \mix1_data_reg_reg[104]/NET0131  , \mix1_data_reg_reg[105]/NET0131  , \mix1_data_reg_reg[106]/NET0131  , \mix1_data_reg_reg[107]/NET0131  , \mix1_data_reg_reg[108]/NET0131  , \mix1_data_reg_reg[109]/NET0131  , \mix1_data_reg_reg[110]/NET0131  , \mix1_data_reg_reg[111]/NET0131  , \mix1_data_reg_reg[112]/NET0131  , \mix1_data_reg_reg[113]/NET0131  , \mix1_data_reg_reg[114]/NET0131  , \mix1_data_reg_reg[115]/NET0131  , \mix1_data_reg_reg[116]/NET0131  , \mix1_data_reg_reg[117]/NET0131  , \mix1_data_reg_reg[118]/NET0131  , \mix1_data_reg_reg[119]/NET0131  , \mix1_data_reg_reg[120]/NET0131  , \mix1_data_reg_reg[121]/NET0131  , \mix1_data_reg_reg[122]/NET0131  , \mix1_data_reg_reg[123]/NET0131  , \mix1_data_reg_reg[124]/NET0131  , \mix1_data_reg_reg[125]/NET0131  , \mix1_data_reg_reg[126]/NET0131  , \mix1_data_reg_reg[127]/NET0131  , \mix1_data_reg_reg[32]/NET0131  , \mix1_data_reg_reg[33]/NET0131  , \mix1_data_reg_reg[34]/NET0131  , \mix1_data_reg_reg[35]/NET0131  , \mix1_data_reg_reg[36]/NET0131  , \mix1_data_reg_reg[37]/NET0131  , \mix1_data_reg_reg[38]/NET0131  , \mix1_data_reg_reg[39]/NET0131  , \mix1_data_reg_reg[40]/NET0131  , \mix1_data_reg_reg[41]/NET0131  , \mix1_data_reg_reg[42]/NET0131  , \mix1_data_reg_reg[43]/NET0131  , \mix1_data_reg_reg[44]/NET0131  , \mix1_data_reg_reg[45]/NET0131  , \mix1_data_reg_reg[46]/NET0131  , \mix1_data_reg_reg[47]/NET0131  , \mix1_data_reg_reg[48]/NET0131  , \mix1_data_reg_reg[49]/NET0131  , \mix1_data_reg_reg[50]/NET0131  , \mix1_data_reg_reg[51]/NET0131  , \mix1_data_reg_reg[52]/NET0131  , \mix1_data_reg_reg[53]/NET0131  , \mix1_data_reg_reg[54]/NET0131  , \mix1_data_reg_reg[55]/NET0131  , \mix1_data_reg_reg[56]/NET0131  , \mix1_data_reg_reg[57]/NET0131  , \mix1_data_reg_reg[58]/NET0131  , \mix1_data_reg_reg[59]/NET0131  , \mix1_data_reg_reg[60]/NET0131  , \mix1_data_reg_reg[61]/NET0131  , \mix1_data_reg_reg[62]/NET0131  , \mix1_data_reg_reg[63]/NET0131  , \mix1_data_reg_reg[64]/NET0131  , \mix1_data_reg_reg[65]/NET0131  , \mix1_data_reg_reg[66]/NET0131  , \mix1_data_reg_reg[67]/NET0131  , \mix1_data_reg_reg[68]/NET0131  , \mix1_data_reg_reg[69]/NET0131  , \mix1_data_reg_reg[70]/NET0131  , \mix1_data_reg_reg[71]/NET0131  , \mix1_data_reg_reg[72]/NET0131  , \mix1_data_reg_reg[73]/NET0131  , \mix1_data_reg_reg[74]/NET0131  , \mix1_data_reg_reg[75]/NET0131  , \mix1_data_reg_reg[76]/NET0131  , \mix1_data_reg_reg[77]/NET0131  , \mix1_data_reg_reg[78]/NET0131  , \mix1_data_reg_reg[79]/NET0131  , \mix1_data_reg_reg[80]/NET0131  , \mix1_data_reg_reg[81]/NET0131  , \mix1_data_reg_reg[82]/NET0131  , \mix1_data_reg_reg[83]/NET0131  , \mix1_data_reg_reg[84]/NET0131  , \mix1_data_reg_reg[85]/NET0131  , \mix1_data_reg_reg[86]/NET0131  , \mix1_data_reg_reg[87]/NET0131  , \mix1_data_reg_reg[88]/NET0131  , \mix1_data_reg_reg[89]/NET0131  , \mix1_data_reg_reg[90]/NET0131  , \mix1_data_reg_reg[91]/NET0131  , \mix1_data_reg_reg[92]/NET0131  , \mix1_data_reg_reg[93]/NET0131  , \mix1_data_reg_reg[94]/NET0131  , \mix1_data_reg_reg[95]/NET0131  , \mix1_data_reg_reg[96]/NET0131  , \mix1_data_reg_reg[97]/NET0131  , \mix1_data_reg_reg[98]/NET0131  , \mix1_data_reg_reg[99]/NET0131  , \mix1_ready_o_reg/NET0131  , \mix1_state_reg[0]/NET0131  , \mix1_state_reg[1]/NET0131  , \round_reg[0]/NET0131  , \round_reg[1]/NET0131  , \round_reg[2]/NET0131  , \round_reg[3]/NET0131  , \sbox1_ah_reg_reg[0]/NET0131  , \sbox1_ah_reg_reg[1]/NET0131  , \sbox1_ah_reg_reg[2]/NET0131  , \sbox1_ah_reg_reg[3]/NET0131  , \sbox1_alph_reg[0]/NET0131  , \sbox1_alph_reg[1]/NET0131  , \sbox1_alph_reg[2]/NET0131  , \sbox1_alph_reg[3]/NET0131  , \sbox1_to_invert_reg[0]/NET0131  , \sbox1_to_invert_reg[1]/NET0131  , \sbox1_to_invert_reg[2]/NET0131  , \sbox1_to_invert_reg[3]/NET0131  , \state_reg/NET0131  , \sub1_data_reg_reg[0]/NET0131  , \sub1_data_reg_reg[100]/NET0131  , \sub1_data_reg_reg[101]/NET0131  , \sub1_data_reg_reg[102]/NET0131  , \sub1_data_reg_reg[103]/NET0131  , \sub1_data_reg_reg[104]/NET0131  , \sub1_data_reg_reg[105]/NET0131  , \sub1_data_reg_reg[106]/NET0131  , \sub1_data_reg_reg[107]/NET0131  , \sub1_data_reg_reg[108]/NET0131  , \sub1_data_reg_reg[109]/NET0131  , \sub1_data_reg_reg[10]/NET0131  , \sub1_data_reg_reg[110]/NET0131  , \sub1_data_reg_reg[111]/NET0131  , \sub1_data_reg_reg[112]/NET0131  , \sub1_data_reg_reg[113]/NET0131  , \sub1_data_reg_reg[114]/NET0131  , \sub1_data_reg_reg[115]/NET0131  , \sub1_data_reg_reg[116]/NET0131  , \sub1_data_reg_reg[117]/NET0131  , \sub1_data_reg_reg[118]/NET0131  , \sub1_data_reg_reg[119]/NET0131  , \sub1_data_reg_reg[11]/NET0131  , \sub1_data_reg_reg[120]/NET0131  , \sub1_data_reg_reg[121]/NET0131  , \sub1_data_reg_reg[122]/NET0131  , \sub1_data_reg_reg[123]/NET0131  , \sub1_data_reg_reg[124]/NET0131  , \sub1_data_reg_reg[125]/NET0131  , \sub1_data_reg_reg[126]/NET0131  , \sub1_data_reg_reg[127]/NET0131  , \sub1_data_reg_reg[12]/NET0131  , \sub1_data_reg_reg[13]/NET0131  , \sub1_data_reg_reg[14]/NET0131  , \sub1_data_reg_reg[15]/NET0131  , \sub1_data_reg_reg[16]/NET0131  , \sub1_data_reg_reg[17]/NET0131  , \sub1_data_reg_reg[18]/NET0131  , \sub1_data_reg_reg[19]/NET0131  , \sub1_data_reg_reg[1]/NET0131  , \sub1_data_reg_reg[20]/NET0131  , \sub1_data_reg_reg[21]/NET0131  , \sub1_data_reg_reg[22]/NET0131  , \sub1_data_reg_reg[23]/NET0131  , \sub1_data_reg_reg[24]/NET0131  , \sub1_data_reg_reg[25]/NET0131  , \sub1_data_reg_reg[26]/NET0131  , \sub1_data_reg_reg[27]/NET0131  , \sub1_data_reg_reg[28]/NET0131  , \sub1_data_reg_reg[29]/NET0131  , \sub1_data_reg_reg[2]/NET0131  , \sub1_data_reg_reg[30]/NET0131  , \sub1_data_reg_reg[31]/NET0131  , \sub1_data_reg_reg[32]/NET0131  , \sub1_data_reg_reg[33]/NET0131  , \sub1_data_reg_reg[34]/NET0131  , \sub1_data_reg_reg[35]/NET0131  , \sub1_data_reg_reg[36]/NET0131  , \sub1_data_reg_reg[37]/NET0131  , \sub1_data_reg_reg[38]/NET0131  , \sub1_data_reg_reg[39]/NET0131  , \sub1_data_reg_reg[3]/NET0131  , \sub1_data_reg_reg[40]/NET0131  , \sub1_data_reg_reg[41]/NET0131  , \sub1_data_reg_reg[42]/NET0131  , \sub1_data_reg_reg[43]/NET0131  , \sub1_data_reg_reg[44]/NET0131  , \sub1_data_reg_reg[45]/NET0131  , \sub1_data_reg_reg[46]/NET0131  , \sub1_data_reg_reg[47]/NET0131  , \sub1_data_reg_reg[48]/NET0131  , \sub1_data_reg_reg[49]/NET0131  , \sub1_data_reg_reg[4]/NET0131  , \sub1_data_reg_reg[50]/NET0131  , \sub1_data_reg_reg[51]/NET0131  , \sub1_data_reg_reg[52]/NET0131  , \sub1_data_reg_reg[53]/NET0131  , \sub1_data_reg_reg[54]/NET0131  , \sub1_data_reg_reg[55]/NET0131  , \sub1_data_reg_reg[56]/NET0131  , \sub1_data_reg_reg[57]/NET0131  , \sub1_data_reg_reg[58]/NET0131  , \sub1_data_reg_reg[59]/NET0131  , \sub1_data_reg_reg[5]/NET0131  , \sub1_data_reg_reg[60]/NET0131  , \sub1_data_reg_reg[61]/NET0131  , \sub1_data_reg_reg[62]/NET0131  , \sub1_data_reg_reg[63]/NET0131  , \sub1_data_reg_reg[64]/NET0131  , \sub1_data_reg_reg[65]/NET0131  , \sub1_data_reg_reg[66]/NET0131  , \sub1_data_reg_reg[67]/NET0131  , \sub1_data_reg_reg[68]/NET0131  , \sub1_data_reg_reg[69]/NET0131  , \sub1_data_reg_reg[6]/NET0131  , \sub1_data_reg_reg[70]/NET0131  , \sub1_data_reg_reg[71]/NET0131  , \sub1_data_reg_reg[72]/NET0131  , \sub1_data_reg_reg[73]/NET0131  , \sub1_data_reg_reg[74]/NET0131  , \sub1_data_reg_reg[75]/NET0131  , \sub1_data_reg_reg[76]/NET0131  , \sub1_data_reg_reg[77]/NET0131  , \sub1_data_reg_reg[78]/NET0131  , \sub1_data_reg_reg[79]/NET0131  , \sub1_data_reg_reg[7]/NET0131  , \sub1_data_reg_reg[80]/NET0131  , \sub1_data_reg_reg[81]/NET0131  , \sub1_data_reg_reg[82]/NET0131  , \sub1_data_reg_reg[83]/NET0131  , \sub1_data_reg_reg[84]/NET0131  , \sub1_data_reg_reg[85]/NET0131  , \sub1_data_reg_reg[86]/NET0131  , \sub1_data_reg_reg[87]/NET0131  , \sub1_data_reg_reg[88]/NET0131  , \sub1_data_reg_reg[89]/NET0131  , \sub1_data_reg_reg[8]/NET0131  , \sub1_data_reg_reg[90]/NET0131  , \sub1_data_reg_reg[91]/NET0131  , \sub1_data_reg_reg[92]/NET0131  , \sub1_data_reg_reg[93]/NET0131  , \sub1_data_reg_reg[94]/NET0131  , \sub1_data_reg_reg[95]/NET0131  , \sub1_data_reg_reg[96]/NET0131  , \sub1_data_reg_reg[97]/NET0131  , \sub1_data_reg_reg[98]/NET0131  , \sub1_data_reg_reg[99]/NET0131  , \sub1_data_reg_reg[9]/NET0131  , \sub1_ready_o_reg/NET0131  , \sub1_state_reg[0]/NET0131  , \sub1_state_reg[1]/NET0131  , \sub1_state_reg[2]/NET0131  , \sub1_state_reg[3]/NET0131  , \sub1_state_reg[4]/NET0131  , \_al_n0  , \_al_n1  , \g27929/_0_  , \g27942/_3_  , \g27943/_3_  , \g27944/_3_  , \g27945/_0_  , \g27995/_0_  , \g27998/_0_  , \g28019/_0_  , \g28020/_0_  , \g28021/_0_  , \g28022/_0_  , \g28023/_0_  , \g28024/_0_  , \g28025/_0_  , \g28026/_0_  , \g28027/_0_  , \g28028/_0_  , \g28029/_0_  , \g28030/_0_  , \g28031/_0_  , \g28032/_0_  , \g28033/_0_  , \g28034/_0_  , \g28044/_0_  , \g28045/_0_  , \g28046/_0_  , \g28047/_0_  , \g28048/_0_  , \g28049/_0_  , \g28050/_0_  , \g28051/_0_  , \g28151/_0_  , \g28177/_0_  , \g28178/_0_  , \g28179/_0_  , \g28180/_0_  , \g28181/_0_  , \g28182/_0_  , \g28183/_0_  , \g28184/_0_  , \g28185/_0_  , \g28186/_0_  , \g28187/_0_  , \g28188/_0_  , \g28189/_0_  , \g28190/_0_  , \g28191/_0_  , \g28192/_0_  , \g28193/_0_  , \g28194/_0_  , \g28195/_0_  , \g28196/_0_  , \g28197/_0_  , \g28198/_0_  , \g28199/_0_  , \g28200/_0_  , \g28201/_0_  , \g28202/_0_  , \g28203/_0_  , \g28253/_0_  , \g28254/_0_  , \g28255/_0_  , \g28256/_0_  , \g28257/_0_  , \g28258/_0_  , \g28259/_0_  , \g28260/_0_  , \g28261/_0_  , \g28262/_0_  , \g28263/_0_  , \g28264/_0_  , \g28265/_0_  , \g28266/_0_  , \g28267/_0_  , \g28268/_0_  , \g28269/_0_  , \g28270/_0_  , \g28271/_0_  , \g28272/_0_  , \g28273/_0_  , \g28274/_0_  , \g28275/_0_  , \g28276/_0_  , \g28277/_0_  , \g28278/_0_  , \g28279/_0_  , \g28384/_2_  , \g28385/_2_  , \g28388/_2_  , \g28389/_2_  , \g28394/_2_  , \g28395/_2_  , \g28401/_2_  , \g28402/_2_  , \g28403/_0_  , \g28404/_0_  , \g28408/_0_  , \g28410/_0_  , \g28440/_0_  , \g28441/_0_  , \g28442/_0_  , \g28443/_0_  , \g28444/_0_  , \g28445/_0_  , \g28446/_0_  , \g28447/_0_  , \g28448/_0_  , \g28449/_0_  , \g28450/_0_  , \g28451/_0_  , \g28452/_0_  , \g28453/_0_  , \g28538/_0_  , \g28539/_0_  , \g28540/_0_  , \g28541/_0_  , \g28542/_0_  , \g28543/_0_  , \g28544/_0_  , \g28545/_0_  , \g28546/_0_  , \g28547/_0_  , \g28548/_0_  , \g28549/_0_  , \g28550/_0_  , \g28551/_0_  , \g28552/_0_  , \g28557/_0_  , \g28558/_0_  , \g28563/_0_  , \g28564/_0_  , \g28565/_0_  , \g28566/_0_  , \g28567/_0_  , \g28625/_2_  , \g28626/_2_  , \g28633/_2_  , \g28639/_2_  , \g28655/_2_  , \g28656/_2_  , \g28657/_2_  , \g28660/_2_  , \g28661/_2_  , \g28662/_2_  , \g28666/_2_  , \g28667/_2_  , \g28668/_2_  , \g28678/_2_  , \g28679/_2_  , \g28680/_2_  , \g28690/_0_  , \g28710/_0_  , \g28716/_0_  , \g28795/_0_  , \g28796/_0_  , \g28798/_0_  , \g28799/_0_  , \g28800/_0_  , \g28801/_0_  , \g28804/_0_  , \g28825/_2_  , \g28826/_2_  , \g28830/_2_  , \g28834/_2_  , \g28842/_2_  , \g28843/_2_  , \g28845/_2_  , \g28848/_2_  , \g28890/_0_  , \g28936/_0_  , \g28982/_0_  , \g29050/_0_  , \g29051/_0_  , \g29052/_0_  , \g29053/_0_  , \g29054/_0_  , \g29055/_0_  , \g29056/_0_  , \g29057/_0_  , \g29058/_0_  , \g29059/_0_  , \g29060/_0_  , \g29061/_0_  , \g29328/_0_  , \g29329/_0_  , \g29330/_0_  , \g29331/_0_  , \g29332/_0_  , \g29333/_0_  , \g29334/_0_  , \g29335/_0_  , \g29336/_0_  , \g29337/_0_  , \g29338/_0_  , \g29339/_0_  , \g29340/_0_  , \g29341/_0_  , \g29342/_0_  , \g29343/_0_  , \g29344/_0_  , \g29345/_0_  , \g29346/_0_  , \g29347/_0_  , \g29348/_0_  , \g29349/_0_  , \g29350/_0_  , \g29351/_0_  , \g29352/_0_  , \g29353/_0_  , \g29354/_0_  , \g29355/_0_  , \g29356/_0_  , \g29357/_0_  , \g29358/_0_  , \g29359/_0_  , \g29360/_0_  , \g29361/_0_  , \g29362/_0_  , \g29363/_0_  , \g29364/_0_  , \g29365/_0_  , \g29366/_0_  , \g29367/_0_  , \g29395/_0_  , \g29396/_0_  , \g29453/_0_  , \g29454/_0_  , \g29455/_0_  , \g29456/_0_  , \g29457/_0_  , \g29458/_0_  , \g29459/_0_  , \g29460/_0_  , \g29461/_0_  , \g29462/_0_  , \g29463/_0_  , \g29464/_0_  , \g29465/_0_  , \g29466/_0_  , \g29467/_0_  , \g29468/_0_  , \g29469/_0_  , \g29470/_0_  , \g29471/_0_  , \g29472/_0_  , \g29473/_0_  , \g29474/_0_  , \g29475/_0_  , \g29476/_0_  , \g29477/_0_  , \g29478/_0_  , \g29479/_0_  , \g29480/_0_  , \g29481/_0_  , \g29482/_0_  , \g29483/_0_  , \g29484/_0_  , \g29485/_0_  , \g29486/_0_  , \g29487/_0_  , \g29488/_0_  , \g29489/_0_  , \g29490/_0_  , \g29491/_0_  , \g29492/_0_  , \g29493/_0_  , \g29494/_0_  , \g29495/_0_  , \g29496/_0_  , \g29497/_0_  , \g29498/_0_  , \g29499/_0_  , \g29500/_0_  , \g29501/_0_  , \g29502/_0_  , \g29503/_0_  , \g29504/_0_  , \g29505/_0_  , \g29506/_0_  , \g29507/_0_  , \g29508/_0_  , \g29509/_0_  , \g29510/_0_  , \g29511/_0_  , \g29512/_0_  , \g29513/_0_  , \g29514/_0_  , \g29515/_0_  , \g29516/_0_  , \g29517/_0_  , \g29518/_0_  , \g29519/_0_  , \g29520/_0_  , \g29521/_0_  , \g29522/_0_  , \g29523/_0_  , \g29524/_0_  , \g29525/_0_  , \g29526/_0_  , \g29527/_0_  , \g29528/_0_  , \g29529/_0_  , \g29530/_0_  , \g29531/_0_  , \g29532/_0_  , \g29533/_0_  , \g29534/_0_  , \g29535/_0_  , \g29536/_0_  , \g29537/_0_  , \g29538/_0_  , \g29539/_0_  , \g29540/_0_  , \g29541/_0_  , \g29542/_0_  , \g29543/_0_  , \g29544/_0_  , \g29545/_0_  , \g29546/_0_  , \g29547/_0_  , \g29548/_0_  , \g29549/_0_  , \g29550/_0_  , \g29551/_0_  , \g29552/_0_  , \g29553/_0_  , \g29554/_0_  , \g29555/_0_  , \g29556/_0_  , \g29557/_0_  , \g29558/_0_  , \g29559/_0_  , \g29560/_0_  , \g29561/_0_  , \g29562/_0_  , \g29563/_0_  , \g29564/_0_  , \g29565/_0_  , \g29566/_0_  , \g29567/_0_  , \g29568/_0_  , \g29569/_0_  , \g29570/_0_  , \g29571/_0_  , \g29572/_0_  , \g29573/_0_  , \g29574/_0_  , \g29575/_0_  , \g29576/_0_  , \g29577/_0_  , \g29578/_0_  , \g29579/_0_  , \g29580/_0_  , \g29582/_0_  , \g29583/_0_  , \g29584/_0_  , \g29585/_0_  , \g29586/_0_  , \g29587/_0_  , \g29588/_0_  , \g29589/_0_  , \g29590/_0_  , \g29591/_0_  , \g29592/_0_  , \g29593/_0_  , \g29634/_0_  , \g29635/_0_  , \g29636/_0_  , \g29637/_0_  , \g29645/_0_  , \g29646/_0_  , \g29647/_0_  , \g29824/_0_  , \g29828/_0_  , \g29832/_0_  , \g29836/_0_  , \g29837/_0_  , \g29838/_0_  , \g29839/_0_  , \g29840/_0_  , \g29841/_0_  , \g29842/_0_  , \g29843/_0_  , \g29844/_0_  , \g29845/_0_  , \g29846/_0_  , \g29847/_0_  , \g29848/_0_  , \g29849/_0_  , \g29850/_0_  , \g29851/_0_  , \g29852/_0_  , \g29853/_0_  , \g29854/_0_  , \g29855/_0_  , \g29856/_0_  , \g29857/_0_  , \g29858/_0_  , \g29859/_0_  , \g29860/_0_  , \g29861/_0_  , \g29862/_0_  , \g29863/_0_  , \g29864/_0_  , \g29865/_0_  , \g29866/_0_  , \g29867/_0_  , \g29868/_0_  , \g30081/_0_  , \g30082/_0_  , \g30083/_0_  , \g30084/_0_  , \g30085/_0_  , \g30086/_0_  , \g30087/_0_  , \g30088/_0_  , \g30089/_0_  , \g30090/_0_  , \g30091/_0_  , \g30092/_0_  , \g30093/_0_  , \g30094/_0_  , \g30095/_0_  , \g30096/_0_  , \g30135/_0_  , \g30137/_0_  , \g30164/_0_  , \g30165/_0_  , \g30166/_0_  , \g30167/_0_  , \g30168/_0_  , \g30169/_0_  , \g30170/_0_  , \g30231/_0_  , \g30232/_0_  , \g30233/_0_  , \g30234/_0_  , \g30235/_0_  , \g30236/_0_  , \g30237/_0_  , \g30238/_0_  , \g30286/_0_  , \g30287/_0_  , \g30288/_0_  , \g30289/_0_  , \g30290/_0_  , \g30291/_0_  , \g30292/_0_  , \g30293/_0_  , \g30294/_0_  , \g30295/_0_  , \g30296/_0_  , \g30297/_0_  , \g30298/_0_  , \g30299/_0_  , \g30300/_0_  , \g30301/_0_  , \g30303/_0_  , \g30304/_0_  , \g30305/_0_  , \g30306/_0_  , \g30307/_0_  , \g30308/_0_  , \g30309/_0_  , \g30310/_0_  , \g30311/_0_  , \g30312/_0_  , \g30313/_0_  , \g30314/_0_  , \g30315/_0_  , \g30316/_0_  , \g30317/_0_  , \g30318/_0_  , \g30319/_0_  , \g30481/_0_  , \g30482/_0_  , \g30483/_0_  , \g30484/_0_  , \g30493/_0_  , \g30495/_0_  , \g30536/_0_  , \g30537/_0_  , \g30538/_0_  , \g30735/_0_  , \g30927/_0_  , \g30928/_0_  , \g30929/_0_  , \g30971/_0_  , \g30972/_0_  , \g30973/_0_  , \g30974/_0_  , \g31129/_0_  , \g31130/_0_  , \g31131/_0_  , \g31132/_0_  , \g31133/_0_  , \g31134/_0_  , \g31135/_0_  , \g31136/_0_  , \g31137/_0_  , \g31138/_0_  , \g31139/_0_  , \g31140/_0_  , \g31141/_0_  , \g31142/_0_  , \g31143/_0_  , \g31144/_0_  , \g31352/_0_  , \g31353/_0_  , \g31354/_0_  , \g31355/_0_  , \g31356/_0_  , \g31357/_0_  , \g31358/_0_  , \g31359/_0_  , \g31360/_0_  , \g31361/_0_  , \g31362/_0_  , \g31363/_0_  , \g31364/_0_  , \g31365/_0_  , \g31366/_0_  , \g31367/_0_  , \g31706/_0_  , \g32001/_0_  , \g32008/_0_  , \g32009/_0_  , \g32010/_0_  , \g32011/_0_  , \g32118/_0_  , \g33261/_0_  , \g33262/_0_  , \g33263/_0_  , \g33264/_0_  , \g33265/_0_  , \g33266/_0_  , \g33450/_0_  , \g33451/_0_  , \g33453/_0_  , \g33485/_0_  , \g33679/_2_  , \g34838/_2_  , \g34971/_0_  , \g34972/_0_  , \g34973/_0_  , \g34974/_0_  , \g34975/_0_  , \g34976/_0_  , \g34977/_0_  , \g34978/_0_  , \g34979/_0_  , \g34980/_0_  , \g34981/_0_  , \g34982/_0_  , \g34983/_0_  , \g34984/_0_  , \g34985/_0_  , \g34986/_0_  , \g34987/_0_  , \g34988/_0_  , \g34989/_0_  , \g34990/_0_  , \g34991/_0_  , \g34992/_0_  , \g34993/_0_  , \g34994/_0_  , \g34995/_0_  , \g34996/_0_  , \g34997/_0_  , \g34998/_0_  , \g34999/_0_  , \g35000/_0_  , \g35001/_0_  , \g35002/_0_  , \g35003/_0_  , \g35004/_0_  , \g35005/_0_  , \g35006/_0_  , \g35007/_0_  , \g35008/_0_  , \g35009/_0_  , \g35010/_0_  , \g35011/_0_  , \g35012/_0_  , \g35013/_0_  , \g35014/_0_  , \g35015/_0_  , \g35016/_0_  , \g35017/_0_  , \g35018/_0_  , \g35019/_0_  , \g35020/_0_  , \g35021/_0_  , \g35022/_0_  , \g35023/_0_  , \g35024/_0_  , \g35025/_0_  , \g35026/_0_  , \g35027/_0_  , \g35028/_0_  , \g35029/_0_  , \g35030/_0_  , \g35031/_0_  , \g35032/_0_  , \g35033/_0_  , \g35034/_0_  , \g35035/_0_  , \g35036/_0_  , \g35037/_0_  , \g35038/_0_  , \g35039/_0_  , \g35040/_0_  , \g35041/_0_  , \g35042/_0_  , \g35043/_0_  , \g35044/_0_  , \g35045/_0_  , \g35046/_0_  , \g35047/_0_  , \g35048/_0_  , \g35049/_0_  , \g35050/_0_  , \g35051/_0_  , \g35052/_0_  , \g35053/_0_  , \g35054/_0_  , \g35055/_0_  , \g35056/_0_  , \g35057/_0_  , \g35058/_0_  , \g35059/_0_  , \g35060/_0_  , \g35061/_0_  , \g35062/_0_  , \g35063/_0_  , \g35064/_0_  , \g35065/_0_  , \g35066/_0_  , \g35538/_0_  , \g35956/_0_  , \g36298/_1_  , \g36324/_0_  , \g36375/_0_  , \g38269/_0_  , \g38473/_0_  , \g38501/_0_  , \g38569/_0_  , \g38629/_0_  , \g38721_dup/_3_  , \g38735/_0_  , \g38753/_0_  , \g38849/_3_  , \g39071/_0_  , \g39073/_0_  , \g39077/_0_  , \g39080/_0_  , \g39135/_0_  , \g39138/_0_  , \g39182/_0_  , \g39197/_3_  , \g39207/_3_  , \g39241/_0_  , \g39272/_0_  , \g39307/_0_  , \g39308/_0_  , \g39361/_0_  , \g39494/_0_  , \g39558/_0_  , \g39575/_0_  , \g39583/_0_  );
  input \addroundkey_ready_o_reg/NET0131  ;
  input \addroundkey_round_reg[0]/NET0131  ;
  input \addroundkey_round_reg[1]/NET0131  ;
  input \addroundkey_round_reg[2]/NET0131  ;
  input \addroundkey_round_reg[3]/NET0131  ;
  input \addroundkey_start_i_reg/NET0131  ;
  input \data_i[0]_pad  ;
  input \data_i[100]_pad  ;
  input \data_i[101]_pad  ;
  input \data_i[102]_pad  ;
  input \data_i[103]_pad  ;
  input \data_i[104]_pad  ;
  input \data_i[105]_pad  ;
  input \data_i[106]_pad  ;
  input \data_i[107]_pad  ;
  input \data_i[108]_pad  ;
  input \data_i[109]_pad  ;
  input \data_i[10]_pad  ;
  input \data_i[110]_pad  ;
  input \data_i[111]_pad  ;
  input \data_i[112]_pad  ;
  input \data_i[113]_pad  ;
  input \data_i[114]_pad  ;
  input \data_i[115]_pad  ;
  input \data_i[116]_pad  ;
  input \data_i[117]_pad  ;
  input \data_i[118]_pad  ;
  input \data_i[119]_pad  ;
  input \data_i[11]_pad  ;
  input \data_i[120]_pad  ;
  input \data_i[121]_pad  ;
  input \data_i[122]_pad  ;
  input \data_i[123]_pad  ;
  input \data_i[124]_pad  ;
  input \data_i[125]_pad  ;
  input \data_i[126]_pad  ;
  input \data_i[127]_pad  ;
  input \data_i[12]_pad  ;
  input \data_i[13]_pad  ;
  input \data_i[14]_pad  ;
  input \data_i[15]_pad  ;
  input \data_i[16]_pad  ;
  input \data_i[17]_pad  ;
  input \data_i[18]_pad  ;
  input \data_i[19]_pad  ;
  input \data_i[1]_pad  ;
  input \data_i[20]_pad  ;
  input \data_i[21]_pad  ;
  input \data_i[22]_pad  ;
  input \data_i[23]_pad  ;
  input \data_i[24]_pad  ;
  input \data_i[25]_pad  ;
  input \data_i[26]_pad  ;
  input \data_i[27]_pad  ;
  input \data_i[28]_pad  ;
  input \data_i[29]_pad  ;
  input \data_i[2]_pad  ;
  input \data_i[30]_pad  ;
  input \data_i[31]_pad  ;
  input \data_i[32]_pad  ;
  input \data_i[33]_pad  ;
  input \data_i[34]_pad  ;
  input \data_i[35]_pad  ;
  input \data_i[36]_pad  ;
  input \data_i[37]_pad  ;
  input \data_i[38]_pad  ;
  input \data_i[39]_pad  ;
  input \data_i[3]_pad  ;
  input \data_i[40]_pad  ;
  input \data_i[41]_pad  ;
  input \data_i[42]_pad  ;
  input \data_i[43]_pad  ;
  input \data_i[44]_pad  ;
  input \data_i[45]_pad  ;
  input \data_i[46]_pad  ;
  input \data_i[47]_pad  ;
  input \data_i[48]_pad  ;
  input \data_i[49]_pad  ;
  input \data_i[4]_pad  ;
  input \data_i[50]_pad  ;
  input \data_i[51]_pad  ;
  input \data_i[52]_pad  ;
  input \data_i[53]_pad  ;
  input \data_i[54]_pad  ;
  input \data_i[55]_pad  ;
  input \data_i[56]_pad  ;
  input \data_i[57]_pad  ;
  input \data_i[58]_pad  ;
  input \data_i[59]_pad  ;
  input \data_i[5]_pad  ;
  input \data_i[60]_pad  ;
  input \data_i[61]_pad  ;
  input \data_i[62]_pad  ;
  input \data_i[63]_pad  ;
  input \data_i[64]_pad  ;
  input \data_i[65]_pad  ;
  input \data_i[66]_pad  ;
  input \data_i[67]_pad  ;
  input \data_i[68]_pad  ;
  input \data_i[69]_pad  ;
  input \data_i[6]_pad  ;
  input \data_i[70]_pad  ;
  input \data_i[71]_pad  ;
  input \data_i[72]_pad  ;
  input \data_i[73]_pad  ;
  input \data_i[74]_pad  ;
  input \data_i[75]_pad  ;
  input \data_i[76]_pad  ;
  input \data_i[77]_pad  ;
  input \data_i[78]_pad  ;
  input \data_i[79]_pad  ;
  input \data_i[7]_pad  ;
  input \data_i[80]_pad  ;
  input \data_i[81]_pad  ;
  input \data_i[82]_pad  ;
  input \data_i[83]_pad  ;
  input \data_i[84]_pad  ;
  input \data_i[85]_pad  ;
  input \data_i[86]_pad  ;
  input \data_i[87]_pad  ;
  input \data_i[88]_pad  ;
  input \data_i[89]_pad  ;
  input \data_i[8]_pad  ;
  input \data_i[90]_pad  ;
  input \data_i[91]_pad  ;
  input \data_i[92]_pad  ;
  input \data_i[93]_pad  ;
  input \data_i[94]_pad  ;
  input \data_i[95]_pad  ;
  input \data_i[96]_pad  ;
  input \data_i[97]_pad  ;
  input \data_i[98]_pad  ;
  input \data_i[99]_pad  ;
  input \data_i[9]_pad  ;
  input \data_o[0]_pad  ;
  input \data_o[100]_pad  ;
  input \data_o[101]_pad  ;
  input \data_o[102]_pad  ;
  input \data_o[103]_pad  ;
  input \data_o[104]_pad  ;
  input \data_o[105]_pad  ;
  input \data_o[106]_pad  ;
  input \data_o[107]_pad  ;
  input \data_o[108]_pad  ;
  input \data_o[109]_pad  ;
  input \data_o[10]_pad  ;
  input \data_o[110]_pad  ;
  input \data_o[111]_pad  ;
  input \data_o[112]_pad  ;
  input \data_o[113]_pad  ;
  input \data_o[114]_pad  ;
  input \data_o[115]_pad  ;
  input \data_o[116]_pad  ;
  input \data_o[117]_pad  ;
  input \data_o[118]_pad  ;
  input \data_o[119]_pad  ;
  input \data_o[11]_pad  ;
  input \data_o[120]_pad  ;
  input \data_o[121]_pad  ;
  input \data_o[122]_pad  ;
  input \data_o[123]_pad  ;
  input \data_o[124]_pad  ;
  input \data_o[125]_pad  ;
  input \data_o[126]_pad  ;
  input \data_o[127]_pad  ;
  input \data_o[12]_pad  ;
  input \data_o[13]_pad  ;
  input \data_o[14]_pad  ;
  input \data_o[15]_pad  ;
  input \data_o[16]_pad  ;
  input \data_o[17]_pad  ;
  input \data_o[18]_pad  ;
  input \data_o[19]_pad  ;
  input \data_o[1]_pad  ;
  input \data_o[20]_pad  ;
  input \data_o[21]_pad  ;
  input \data_o[22]_pad  ;
  input \data_o[23]_pad  ;
  input \data_o[24]_pad  ;
  input \data_o[25]_pad  ;
  input \data_o[26]_pad  ;
  input \data_o[27]_pad  ;
  input \data_o[28]_pad  ;
  input \data_o[29]_pad  ;
  input \data_o[2]_pad  ;
  input \data_o[30]_pad  ;
  input \data_o[31]_pad  ;
  input \data_o[32]_pad  ;
  input \data_o[33]_pad  ;
  input \data_o[34]_pad  ;
  input \data_o[35]_pad  ;
  input \data_o[36]_pad  ;
  input \data_o[37]_pad  ;
  input \data_o[38]_pad  ;
  input \data_o[39]_pad  ;
  input \data_o[3]_pad  ;
  input \data_o[40]_pad  ;
  input \data_o[41]_pad  ;
  input \data_o[42]_pad  ;
  input \data_o[43]_pad  ;
  input \data_o[44]_pad  ;
  input \data_o[45]_pad  ;
  input \data_o[46]_pad  ;
  input \data_o[47]_pad  ;
  input \data_o[48]_pad  ;
  input \data_o[49]_pad  ;
  input \data_o[4]_pad  ;
  input \data_o[50]_pad  ;
  input \data_o[51]_pad  ;
  input \data_o[52]_pad  ;
  input \data_o[53]_pad  ;
  input \data_o[54]_pad  ;
  input \data_o[55]_pad  ;
  input \data_o[56]_pad  ;
  input \data_o[57]_pad  ;
  input \data_o[58]_pad  ;
  input \data_o[59]_pad  ;
  input \data_o[5]_pad  ;
  input \data_o[60]_pad  ;
  input \data_o[61]_pad  ;
  input \data_o[62]_pad  ;
  input \data_o[63]_pad  ;
  input \data_o[64]_pad  ;
  input \data_o[65]_pad  ;
  input \data_o[66]_pad  ;
  input \data_o[67]_pad  ;
  input \data_o[68]_pad  ;
  input \data_o[69]_pad  ;
  input \data_o[6]_pad  ;
  input \data_o[70]_pad  ;
  input \data_o[71]_pad  ;
  input \data_o[72]_pad  ;
  input \data_o[73]_pad  ;
  input \data_o[74]_pad  ;
  input \data_o[75]_pad  ;
  input \data_o[76]_pad  ;
  input \data_o[77]_pad  ;
  input \data_o[78]_pad  ;
  input \data_o[79]_pad  ;
  input \data_o[7]_pad  ;
  input \data_o[80]_pad  ;
  input \data_o[81]_pad  ;
  input \data_o[82]_pad  ;
  input \data_o[83]_pad  ;
  input \data_o[84]_pad  ;
  input \data_o[85]_pad  ;
  input \data_o[86]_pad  ;
  input \data_o[87]_pad  ;
  input \data_o[88]_pad  ;
  input \data_o[89]_pad  ;
  input \data_o[8]_pad  ;
  input \data_o[90]_pad  ;
  input \data_o[91]_pad  ;
  input \data_o[92]_pad  ;
  input \data_o[93]_pad  ;
  input \data_o[94]_pad  ;
  input \data_o[95]_pad  ;
  input \data_o[96]_pad  ;
  input \data_o[97]_pad  ;
  input \data_o[98]_pad  ;
  input \data_o[99]_pad  ;
  input \data_o[9]_pad  ;
  input decrypt_i_pad ;
  input \first_round_reg_reg/NET0131  ;
  input \key_i[0]_pad  ;
  input \key_i[100]_pad  ;
  input \key_i[101]_pad  ;
  input \key_i[102]_pad  ;
  input \key_i[103]_pad  ;
  input \key_i[104]_pad  ;
  input \key_i[105]_pad  ;
  input \key_i[106]_pad  ;
  input \key_i[107]_pad  ;
  input \key_i[108]_pad  ;
  input \key_i[109]_pad  ;
  input \key_i[10]_pad  ;
  input \key_i[110]_pad  ;
  input \key_i[111]_pad  ;
  input \key_i[112]_pad  ;
  input \key_i[113]_pad  ;
  input \key_i[114]_pad  ;
  input \key_i[115]_pad  ;
  input \key_i[116]_pad  ;
  input \key_i[117]_pad  ;
  input \key_i[118]_pad  ;
  input \key_i[119]_pad  ;
  input \key_i[11]_pad  ;
  input \key_i[120]_pad  ;
  input \key_i[121]_pad  ;
  input \key_i[122]_pad  ;
  input \key_i[123]_pad  ;
  input \key_i[124]_pad  ;
  input \key_i[125]_pad  ;
  input \key_i[126]_pad  ;
  input \key_i[127]_pad  ;
  input \key_i[12]_pad  ;
  input \key_i[13]_pad  ;
  input \key_i[14]_pad  ;
  input \key_i[15]_pad  ;
  input \key_i[16]_pad  ;
  input \key_i[17]_pad  ;
  input \key_i[18]_pad  ;
  input \key_i[19]_pad  ;
  input \key_i[1]_pad  ;
  input \key_i[20]_pad  ;
  input \key_i[21]_pad  ;
  input \key_i[22]_pad  ;
  input \key_i[23]_pad  ;
  input \key_i[24]_pad  ;
  input \key_i[25]_pad  ;
  input \key_i[26]_pad  ;
  input \key_i[27]_pad  ;
  input \key_i[28]_pad  ;
  input \key_i[29]_pad  ;
  input \key_i[2]_pad  ;
  input \key_i[30]_pad  ;
  input \key_i[31]_pad  ;
  input \key_i[32]_pad  ;
  input \key_i[33]_pad  ;
  input \key_i[34]_pad  ;
  input \key_i[35]_pad  ;
  input \key_i[36]_pad  ;
  input \key_i[37]_pad  ;
  input \key_i[38]_pad  ;
  input \key_i[39]_pad  ;
  input \key_i[3]_pad  ;
  input \key_i[40]_pad  ;
  input \key_i[41]_pad  ;
  input \key_i[42]_pad  ;
  input \key_i[43]_pad  ;
  input \key_i[44]_pad  ;
  input \key_i[45]_pad  ;
  input \key_i[46]_pad  ;
  input \key_i[47]_pad  ;
  input \key_i[48]_pad  ;
  input \key_i[49]_pad  ;
  input \key_i[4]_pad  ;
  input \key_i[50]_pad  ;
  input \key_i[51]_pad  ;
  input \key_i[52]_pad  ;
  input \key_i[53]_pad  ;
  input \key_i[54]_pad  ;
  input \key_i[55]_pad  ;
  input \key_i[56]_pad  ;
  input \key_i[57]_pad  ;
  input \key_i[58]_pad  ;
  input \key_i[59]_pad  ;
  input \key_i[5]_pad  ;
  input \key_i[60]_pad  ;
  input \key_i[61]_pad  ;
  input \key_i[62]_pad  ;
  input \key_i[63]_pad  ;
  input \key_i[64]_pad  ;
  input \key_i[65]_pad  ;
  input \key_i[66]_pad  ;
  input \key_i[67]_pad  ;
  input \key_i[68]_pad  ;
  input \key_i[69]_pad  ;
  input \key_i[6]_pad  ;
  input \key_i[70]_pad  ;
  input \key_i[71]_pad  ;
  input \key_i[72]_pad  ;
  input \key_i[73]_pad  ;
  input \key_i[74]_pad  ;
  input \key_i[75]_pad  ;
  input \key_i[76]_pad  ;
  input \key_i[77]_pad  ;
  input \key_i[78]_pad  ;
  input \key_i[79]_pad  ;
  input \key_i[7]_pad  ;
  input \key_i[80]_pad  ;
  input \key_i[81]_pad  ;
  input \key_i[82]_pad  ;
  input \key_i[83]_pad  ;
  input \key_i[84]_pad  ;
  input \key_i[85]_pad  ;
  input \key_i[86]_pad  ;
  input \key_i[87]_pad  ;
  input \key_i[88]_pad  ;
  input \key_i[89]_pad  ;
  input \key_i[8]_pad  ;
  input \key_i[90]_pad  ;
  input \key_i[91]_pad  ;
  input \key_i[92]_pad  ;
  input \key_i[93]_pad  ;
  input \key_i[94]_pad  ;
  input \key_i[95]_pad  ;
  input \key_i[96]_pad  ;
  input \key_i[97]_pad  ;
  input \key_i[98]_pad  ;
  input \key_i[99]_pad  ;
  input \key_i[9]_pad  ;
  input \ks1_col_reg[0]/NET0131  ;
  input \ks1_col_reg[16]/NET0131  ;
  input \ks1_col_reg[17]/NET0131  ;
  input \ks1_col_reg[18]/NET0131  ;
  input \ks1_col_reg[19]/NET0131  ;
  input \ks1_col_reg[1]/NET0131  ;
  input \ks1_col_reg[20]/NET0131  ;
  input \ks1_col_reg[21]/NET0131  ;
  input \ks1_col_reg[22]/NET0131  ;
  input \ks1_col_reg[23]/NET0131  ;
  input \ks1_col_reg[24]/NET0131  ;
  input \ks1_col_reg[25]/NET0131  ;
  input \ks1_col_reg[26]/NET0131  ;
  input \ks1_col_reg[27]/NET0131  ;
  input \ks1_col_reg[28]/NET0131  ;
  input \ks1_col_reg[29]/NET0131  ;
  input \ks1_col_reg[2]/NET0131  ;
  input \ks1_col_reg[30]/NET0131  ;
  input \ks1_col_reg[31]/NET0131  ;
  input \ks1_col_reg[3]/NET0131  ;
  input \ks1_col_reg[4]/NET0131  ;
  input \ks1_col_reg[5]/NET0131  ;
  input \ks1_col_reg[6]/NET0131  ;
  input \ks1_col_reg[7]/NET0131  ;
  input \ks1_key_reg_reg[0]/NET0131  ;
  input \ks1_key_reg_reg[100]/NET0131  ;
  input \ks1_key_reg_reg[101]/NET0131  ;
  input \ks1_key_reg_reg[102]/NET0131  ;
  input \ks1_key_reg_reg[103]/NET0131  ;
  input \ks1_key_reg_reg[104]/NET0131  ;
  input \ks1_key_reg_reg[105]/NET0131  ;
  input \ks1_key_reg_reg[106]/NET0131  ;
  input \ks1_key_reg_reg[107]/NET0131  ;
  input \ks1_key_reg_reg[108]/NET0131  ;
  input \ks1_key_reg_reg[109]/P0002  ;
  input \ks1_key_reg_reg[10]/NET0131  ;
  input \ks1_key_reg_reg[110]/P0002  ;
  input \ks1_key_reg_reg[111]/NET0131  ;
  input \ks1_key_reg_reg[112]/NET0131  ;
  input \ks1_key_reg_reg[113]/NET0131  ;
  input \ks1_key_reg_reg[114]/NET0131  ;
  input \ks1_key_reg_reg[115]/NET0131  ;
  input \ks1_key_reg_reg[116]/NET0131  ;
  input \ks1_key_reg_reg[117]/NET0131  ;
  input \ks1_key_reg_reg[118]/NET0131  ;
  input \ks1_key_reg_reg[119]/NET0131  ;
  input \ks1_key_reg_reg[11]/NET0131  ;
  input \ks1_key_reg_reg[120]/NET0131  ;
  input \ks1_key_reg_reg[121]/NET0131  ;
  input \ks1_key_reg_reg[122]/NET0131  ;
  input \ks1_key_reg_reg[123]/NET0131  ;
  input \ks1_key_reg_reg[124]/NET0131  ;
  input \ks1_key_reg_reg[125]/NET0131  ;
  input \ks1_key_reg_reg[126]/NET0131  ;
  input \ks1_key_reg_reg[127]/NET0131  ;
  input \ks1_key_reg_reg[12]/NET0131  ;
  input \ks1_key_reg_reg[13]/NET0131  ;
  input \ks1_key_reg_reg[14]/NET0131  ;
  input \ks1_key_reg_reg[15]/NET0131  ;
  input \ks1_key_reg_reg[16]/NET0131  ;
  input \ks1_key_reg_reg[17]/NET0131  ;
  input \ks1_key_reg_reg[18]/NET0131  ;
  input \ks1_key_reg_reg[19]/NET0131  ;
  input \ks1_key_reg_reg[1]/NET0131  ;
  input \ks1_key_reg_reg[20]/NET0131  ;
  input \ks1_key_reg_reg[21]/NET0131  ;
  input \ks1_key_reg_reg[22]/NET0131  ;
  input \ks1_key_reg_reg[23]/NET0131  ;
  input \ks1_key_reg_reg[24]/NET0131  ;
  input \ks1_key_reg_reg[25]/NET0131  ;
  input \ks1_key_reg_reg[26]/NET0131  ;
  input \ks1_key_reg_reg[27]/NET0131  ;
  input \ks1_key_reg_reg[28]/NET0131  ;
  input \ks1_key_reg_reg[29]/NET0131  ;
  input \ks1_key_reg_reg[2]/NET0131  ;
  input \ks1_key_reg_reg[30]/NET0131  ;
  input \ks1_key_reg_reg[31]/NET0131  ;
  input \ks1_key_reg_reg[32]/NET0131  ;
  input \ks1_key_reg_reg[33]/NET0131  ;
  input \ks1_key_reg_reg[34]/NET0131  ;
  input \ks1_key_reg_reg[35]/NET0131  ;
  input \ks1_key_reg_reg[36]/NET0131  ;
  input \ks1_key_reg_reg[37]/NET0131  ;
  input \ks1_key_reg_reg[38]/NET0131  ;
  input \ks1_key_reg_reg[39]/NET0131  ;
  input \ks1_key_reg_reg[3]/NET0131  ;
  input \ks1_key_reg_reg[40]/P0002  ;
  input \ks1_key_reg_reg[41]/P0002  ;
  input \ks1_key_reg_reg[42]/P0002  ;
  input \ks1_key_reg_reg[43]/P0002  ;
  input \ks1_key_reg_reg[44]/P0002  ;
  input \ks1_key_reg_reg[45]/P0002  ;
  input \ks1_key_reg_reg[46]/P0002  ;
  input \ks1_key_reg_reg[47]/P0002  ;
  input \ks1_key_reg_reg[48]/NET0131  ;
  input \ks1_key_reg_reg[49]/NET0131  ;
  input \ks1_key_reg_reg[4]/NET0131  ;
  input \ks1_key_reg_reg[50]/NET0131  ;
  input \ks1_key_reg_reg[51]/NET0131  ;
  input \ks1_key_reg_reg[52]/NET0131  ;
  input \ks1_key_reg_reg[53]/NET0131  ;
  input \ks1_key_reg_reg[54]/NET0131  ;
  input \ks1_key_reg_reg[55]/NET0131  ;
  input \ks1_key_reg_reg[56]/NET0131  ;
  input \ks1_key_reg_reg[57]/NET0131  ;
  input \ks1_key_reg_reg[58]/NET0131  ;
  input \ks1_key_reg_reg[59]/NET0131  ;
  input \ks1_key_reg_reg[5]/NET0131  ;
  input \ks1_key_reg_reg[60]/NET0131  ;
  input \ks1_key_reg_reg[61]/NET0131  ;
  input \ks1_key_reg_reg[62]/NET0131  ;
  input \ks1_key_reg_reg[63]/NET0131  ;
  input \ks1_key_reg_reg[64]/NET0131  ;
  input \ks1_key_reg_reg[65]/NET0131  ;
  input \ks1_key_reg_reg[66]/NET0131  ;
  input \ks1_key_reg_reg[67]/NET0131  ;
  input \ks1_key_reg_reg[68]/NET0131  ;
  input \ks1_key_reg_reg[69]/NET0131  ;
  input \ks1_key_reg_reg[6]/NET0131  ;
  input \ks1_key_reg_reg[70]/NET0131  ;
  input \ks1_key_reg_reg[71]/NET0131  ;
  input \ks1_key_reg_reg[72]/P0002  ;
  input \ks1_key_reg_reg[73]/NET0131  ;
  input \ks1_key_reg_reg[74]/NET0131  ;
  input \ks1_key_reg_reg[75]/P0002  ;
  input \ks1_key_reg_reg[76]/P0002  ;
  input \ks1_key_reg_reg[77]/P0002  ;
  input \ks1_key_reg_reg[78]/P0002  ;
  input \ks1_key_reg_reg[79]/P0002  ;
  input \ks1_key_reg_reg[7]/NET0131  ;
  input \ks1_key_reg_reg[80]/NET0131  ;
  input \ks1_key_reg_reg[81]/NET0131  ;
  input \ks1_key_reg_reg[82]/NET0131  ;
  input \ks1_key_reg_reg[83]/NET0131  ;
  input \ks1_key_reg_reg[84]/NET0131  ;
  input \ks1_key_reg_reg[85]/NET0131  ;
  input \ks1_key_reg_reg[86]/NET0131  ;
  input \ks1_key_reg_reg[87]/NET0131  ;
  input \ks1_key_reg_reg[88]/NET0131  ;
  input \ks1_key_reg_reg[89]/NET0131  ;
  input \ks1_key_reg_reg[8]/NET0131  ;
  input \ks1_key_reg_reg[90]/NET0131  ;
  input \ks1_key_reg_reg[91]/NET0131  ;
  input \ks1_key_reg_reg[92]/NET0131  ;
  input \ks1_key_reg_reg[93]/NET0131  ;
  input \ks1_key_reg_reg[94]/NET0131  ;
  input \ks1_key_reg_reg[95]/NET0131  ;
  input \ks1_key_reg_reg[96]/NET0131  ;
  input \ks1_key_reg_reg[97]/NET0131  ;
  input \ks1_key_reg_reg[98]/NET0131  ;
  input \ks1_key_reg_reg[99]/NET0131  ;
  input \ks1_key_reg_reg[9]/NET0131  ;
  input \ks1_ready_o_reg/NET0131  ;
  input \ks1_state_reg[0]/NET0131  ;
  input \ks1_state_reg[1]/NET0131  ;
  input \ks1_state_reg[2]/NET0131  ;
  input load_i_pad ;
  input \mix1_data_o_reg_reg[0]/NET0131  ;
  input \mix1_data_o_reg_reg[100]/NET0131  ;
  input \mix1_data_o_reg_reg[101]/NET0131  ;
  input \mix1_data_o_reg_reg[102]/NET0131  ;
  input \mix1_data_o_reg_reg[103]/NET0131  ;
  input \mix1_data_o_reg_reg[104]/NET0131  ;
  input \mix1_data_o_reg_reg[105]/NET0131  ;
  input \mix1_data_o_reg_reg[106]/NET0131  ;
  input \mix1_data_o_reg_reg[107]/NET0131  ;
  input \mix1_data_o_reg_reg[108]/NET0131  ;
  input \mix1_data_o_reg_reg[109]/NET0131  ;
  input \mix1_data_o_reg_reg[10]/NET0131  ;
  input \mix1_data_o_reg_reg[110]/NET0131  ;
  input \mix1_data_o_reg_reg[111]/NET0131  ;
  input \mix1_data_o_reg_reg[112]/NET0131  ;
  input \mix1_data_o_reg_reg[113]/NET0131  ;
  input \mix1_data_o_reg_reg[114]/NET0131  ;
  input \mix1_data_o_reg_reg[115]/NET0131  ;
  input \mix1_data_o_reg_reg[116]/NET0131  ;
  input \mix1_data_o_reg_reg[117]/NET0131  ;
  input \mix1_data_o_reg_reg[118]/NET0131  ;
  input \mix1_data_o_reg_reg[119]/NET0131  ;
  input \mix1_data_o_reg_reg[11]/NET0131  ;
  input \mix1_data_o_reg_reg[120]/NET0131  ;
  input \mix1_data_o_reg_reg[121]/NET0131  ;
  input \mix1_data_o_reg_reg[122]/NET0131  ;
  input \mix1_data_o_reg_reg[123]/NET0131  ;
  input \mix1_data_o_reg_reg[124]/NET0131  ;
  input \mix1_data_o_reg_reg[125]/NET0131  ;
  input \mix1_data_o_reg_reg[126]/NET0131  ;
  input \mix1_data_o_reg_reg[127]/NET0131  ;
  input \mix1_data_o_reg_reg[12]/NET0131  ;
  input \mix1_data_o_reg_reg[13]/NET0131  ;
  input \mix1_data_o_reg_reg[14]/NET0131  ;
  input \mix1_data_o_reg_reg[15]/NET0131  ;
  input \mix1_data_o_reg_reg[16]/NET0131  ;
  input \mix1_data_o_reg_reg[17]/NET0131  ;
  input \mix1_data_o_reg_reg[18]/NET0131  ;
  input \mix1_data_o_reg_reg[19]/NET0131  ;
  input \mix1_data_o_reg_reg[1]/NET0131  ;
  input \mix1_data_o_reg_reg[20]/NET0131  ;
  input \mix1_data_o_reg_reg[21]/NET0131  ;
  input \mix1_data_o_reg_reg[22]/NET0131  ;
  input \mix1_data_o_reg_reg[23]/NET0131  ;
  input \mix1_data_o_reg_reg[24]/NET0131  ;
  input \mix1_data_o_reg_reg[25]/NET0131  ;
  input \mix1_data_o_reg_reg[26]/NET0131  ;
  input \mix1_data_o_reg_reg[27]/NET0131  ;
  input \mix1_data_o_reg_reg[28]/NET0131  ;
  input \mix1_data_o_reg_reg[29]/NET0131  ;
  input \mix1_data_o_reg_reg[2]/NET0131  ;
  input \mix1_data_o_reg_reg[30]/NET0131  ;
  input \mix1_data_o_reg_reg[31]/NET0131  ;
  input \mix1_data_o_reg_reg[32]/NET0131  ;
  input \mix1_data_o_reg_reg[33]/NET0131  ;
  input \mix1_data_o_reg_reg[34]/NET0131  ;
  input \mix1_data_o_reg_reg[35]/NET0131  ;
  input \mix1_data_o_reg_reg[36]/NET0131  ;
  input \mix1_data_o_reg_reg[37]/NET0131  ;
  input \mix1_data_o_reg_reg[38]/NET0131  ;
  input \mix1_data_o_reg_reg[39]/NET0131  ;
  input \mix1_data_o_reg_reg[3]/NET0131  ;
  input \mix1_data_o_reg_reg[40]/NET0131  ;
  input \mix1_data_o_reg_reg[41]/NET0131  ;
  input \mix1_data_o_reg_reg[42]/NET0131  ;
  input \mix1_data_o_reg_reg[43]/NET0131  ;
  input \mix1_data_o_reg_reg[44]/NET0131  ;
  input \mix1_data_o_reg_reg[45]/NET0131  ;
  input \mix1_data_o_reg_reg[46]/NET0131  ;
  input \mix1_data_o_reg_reg[47]/NET0131  ;
  input \mix1_data_o_reg_reg[48]/NET0131  ;
  input \mix1_data_o_reg_reg[49]/NET0131  ;
  input \mix1_data_o_reg_reg[4]/NET0131  ;
  input \mix1_data_o_reg_reg[50]/NET0131  ;
  input \mix1_data_o_reg_reg[51]/NET0131  ;
  input \mix1_data_o_reg_reg[52]/NET0131  ;
  input \mix1_data_o_reg_reg[53]/NET0131  ;
  input \mix1_data_o_reg_reg[54]/NET0131  ;
  input \mix1_data_o_reg_reg[55]/NET0131  ;
  input \mix1_data_o_reg_reg[56]/NET0131  ;
  input \mix1_data_o_reg_reg[57]/NET0131  ;
  input \mix1_data_o_reg_reg[58]/NET0131  ;
  input \mix1_data_o_reg_reg[59]/NET0131  ;
  input \mix1_data_o_reg_reg[5]/NET0131  ;
  input \mix1_data_o_reg_reg[60]/NET0131  ;
  input \mix1_data_o_reg_reg[61]/NET0131  ;
  input \mix1_data_o_reg_reg[62]/NET0131  ;
  input \mix1_data_o_reg_reg[63]/NET0131  ;
  input \mix1_data_o_reg_reg[64]/NET0131  ;
  input \mix1_data_o_reg_reg[65]/NET0131  ;
  input \mix1_data_o_reg_reg[66]/NET0131  ;
  input \mix1_data_o_reg_reg[67]/NET0131  ;
  input \mix1_data_o_reg_reg[68]/NET0131  ;
  input \mix1_data_o_reg_reg[69]/NET0131  ;
  input \mix1_data_o_reg_reg[6]/NET0131  ;
  input \mix1_data_o_reg_reg[70]/NET0131  ;
  input \mix1_data_o_reg_reg[71]/NET0131  ;
  input \mix1_data_o_reg_reg[72]/NET0131  ;
  input \mix1_data_o_reg_reg[73]/NET0131  ;
  input \mix1_data_o_reg_reg[74]/NET0131  ;
  input \mix1_data_o_reg_reg[75]/NET0131  ;
  input \mix1_data_o_reg_reg[76]/NET0131  ;
  input \mix1_data_o_reg_reg[77]/NET0131  ;
  input \mix1_data_o_reg_reg[78]/NET0131  ;
  input \mix1_data_o_reg_reg[79]/NET0131  ;
  input \mix1_data_o_reg_reg[7]/NET0131  ;
  input \mix1_data_o_reg_reg[80]/NET0131  ;
  input \mix1_data_o_reg_reg[81]/NET0131  ;
  input \mix1_data_o_reg_reg[82]/NET0131  ;
  input \mix1_data_o_reg_reg[83]/NET0131  ;
  input \mix1_data_o_reg_reg[84]/NET0131  ;
  input \mix1_data_o_reg_reg[85]/NET0131  ;
  input \mix1_data_o_reg_reg[86]/NET0131  ;
  input \mix1_data_o_reg_reg[87]/NET0131  ;
  input \mix1_data_o_reg_reg[88]/NET0131  ;
  input \mix1_data_o_reg_reg[89]/NET0131  ;
  input \mix1_data_o_reg_reg[8]/NET0131  ;
  input \mix1_data_o_reg_reg[90]/NET0131  ;
  input \mix1_data_o_reg_reg[91]/NET0131  ;
  input \mix1_data_o_reg_reg[92]/NET0131  ;
  input \mix1_data_o_reg_reg[93]/NET0131  ;
  input \mix1_data_o_reg_reg[94]/NET0131  ;
  input \mix1_data_o_reg_reg[95]/NET0131  ;
  input \mix1_data_o_reg_reg[96]/NET0131  ;
  input \mix1_data_o_reg_reg[97]/NET0131  ;
  input \mix1_data_o_reg_reg[98]/NET0131  ;
  input \mix1_data_o_reg_reg[99]/NET0131  ;
  input \mix1_data_o_reg_reg[9]/NET0131  ;
  input \mix1_data_reg_reg[100]/NET0131  ;
  input \mix1_data_reg_reg[101]/NET0131  ;
  input \mix1_data_reg_reg[102]/NET0131  ;
  input \mix1_data_reg_reg[103]/NET0131  ;
  input \mix1_data_reg_reg[104]/NET0131  ;
  input \mix1_data_reg_reg[105]/NET0131  ;
  input \mix1_data_reg_reg[106]/NET0131  ;
  input \mix1_data_reg_reg[107]/NET0131  ;
  input \mix1_data_reg_reg[108]/NET0131  ;
  input \mix1_data_reg_reg[109]/NET0131  ;
  input \mix1_data_reg_reg[110]/NET0131  ;
  input \mix1_data_reg_reg[111]/NET0131  ;
  input \mix1_data_reg_reg[112]/NET0131  ;
  input \mix1_data_reg_reg[113]/NET0131  ;
  input \mix1_data_reg_reg[114]/NET0131  ;
  input \mix1_data_reg_reg[115]/NET0131  ;
  input \mix1_data_reg_reg[116]/NET0131  ;
  input \mix1_data_reg_reg[117]/NET0131  ;
  input \mix1_data_reg_reg[118]/NET0131  ;
  input \mix1_data_reg_reg[119]/NET0131  ;
  input \mix1_data_reg_reg[120]/NET0131  ;
  input \mix1_data_reg_reg[121]/NET0131  ;
  input \mix1_data_reg_reg[122]/NET0131  ;
  input \mix1_data_reg_reg[123]/NET0131  ;
  input \mix1_data_reg_reg[124]/NET0131  ;
  input \mix1_data_reg_reg[125]/NET0131  ;
  input \mix1_data_reg_reg[126]/NET0131  ;
  input \mix1_data_reg_reg[127]/NET0131  ;
  input \mix1_data_reg_reg[32]/NET0131  ;
  input \mix1_data_reg_reg[33]/NET0131  ;
  input \mix1_data_reg_reg[34]/NET0131  ;
  input \mix1_data_reg_reg[35]/NET0131  ;
  input \mix1_data_reg_reg[36]/NET0131  ;
  input \mix1_data_reg_reg[37]/NET0131  ;
  input \mix1_data_reg_reg[38]/NET0131  ;
  input \mix1_data_reg_reg[39]/NET0131  ;
  input \mix1_data_reg_reg[40]/NET0131  ;
  input \mix1_data_reg_reg[41]/NET0131  ;
  input \mix1_data_reg_reg[42]/NET0131  ;
  input \mix1_data_reg_reg[43]/NET0131  ;
  input \mix1_data_reg_reg[44]/NET0131  ;
  input \mix1_data_reg_reg[45]/NET0131  ;
  input \mix1_data_reg_reg[46]/NET0131  ;
  input \mix1_data_reg_reg[47]/NET0131  ;
  input \mix1_data_reg_reg[48]/NET0131  ;
  input \mix1_data_reg_reg[49]/NET0131  ;
  input \mix1_data_reg_reg[50]/NET0131  ;
  input \mix1_data_reg_reg[51]/NET0131  ;
  input \mix1_data_reg_reg[52]/NET0131  ;
  input \mix1_data_reg_reg[53]/NET0131  ;
  input \mix1_data_reg_reg[54]/NET0131  ;
  input \mix1_data_reg_reg[55]/NET0131  ;
  input \mix1_data_reg_reg[56]/NET0131  ;
  input \mix1_data_reg_reg[57]/NET0131  ;
  input \mix1_data_reg_reg[58]/NET0131  ;
  input \mix1_data_reg_reg[59]/NET0131  ;
  input \mix1_data_reg_reg[60]/NET0131  ;
  input \mix1_data_reg_reg[61]/NET0131  ;
  input \mix1_data_reg_reg[62]/NET0131  ;
  input \mix1_data_reg_reg[63]/NET0131  ;
  input \mix1_data_reg_reg[64]/NET0131  ;
  input \mix1_data_reg_reg[65]/NET0131  ;
  input \mix1_data_reg_reg[66]/NET0131  ;
  input \mix1_data_reg_reg[67]/NET0131  ;
  input \mix1_data_reg_reg[68]/NET0131  ;
  input \mix1_data_reg_reg[69]/NET0131  ;
  input \mix1_data_reg_reg[70]/NET0131  ;
  input \mix1_data_reg_reg[71]/NET0131  ;
  input \mix1_data_reg_reg[72]/NET0131  ;
  input \mix1_data_reg_reg[73]/NET0131  ;
  input \mix1_data_reg_reg[74]/NET0131  ;
  input \mix1_data_reg_reg[75]/NET0131  ;
  input \mix1_data_reg_reg[76]/NET0131  ;
  input \mix1_data_reg_reg[77]/NET0131  ;
  input \mix1_data_reg_reg[78]/NET0131  ;
  input \mix1_data_reg_reg[79]/NET0131  ;
  input \mix1_data_reg_reg[80]/NET0131  ;
  input \mix1_data_reg_reg[81]/NET0131  ;
  input \mix1_data_reg_reg[82]/NET0131  ;
  input \mix1_data_reg_reg[83]/NET0131  ;
  input \mix1_data_reg_reg[84]/NET0131  ;
  input \mix1_data_reg_reg[85]/NET0131  ;
  input \mix1_data_reg_reg[86]/NET0131  ;
  input \mix1_data_reg_reg[87]/NET0131  ;
  input \mix1_data_reg_reg[88]/NET0131  ;
  input \mix1_data_reg_reg[89]/NET0131  ;
  input \mix1_data_reg_reg[90]/NET0131  ;
  input \mix1_data_reg_reg[91]/NET0131  ;
  input \mix1_data_reg_reg[92]/NET0131  ;
  input \mix1_data_reg_reg[93]/NET0131  ;
  input \mix1_data_reg_reg[94]/NET0131  ;
  input \mix1_data_reg_reg[95]/NET0131  ;
  input \mix1_data_reg_reg[96]/NET0131  ;
  input \mix1_data_reg_reg[97]/NET0131  ;
  input \mix1_data_reg_reg[98]/NET0131  ;
  input \mix1_data_reg_reg[99]/NET0131  ;
  input \mix1_ready_o_reg/NET0131  ;
  input \mix1_state_reg[0]/NET0131  ;
  input \mix1_state_reg[1]/NET0131  ;
  input \round_reg[0]/NET0131  ;
  input \round_reg[1]/NET0131  ;
  input \round_reg[2]/NET0131  ;
  input \round_reg[3]/NET0131  ;
  input \sbox1_ah_reg_reg[0]/NET0131  ;
  input \sbox1_ah_reg_reg[1]/NET0131  ;
  input \sbox1_ah_reg_reg[2]/NET0131  ;
  input \sbox1_ah_reg_reg[3]/NET0131  ;
  input \sbox1_alph_reg[0]/NET0131  ;
  input \sbox1_alph_reg[1]/NET0131  ;
  input \sbox1_alph_reg[2]/NET0131  ;
  input \sbox1_alph_reg[3]/NET0131  ;
  input \sbox1_to_invert_reg[0]/NET0131  ;
  input \sbox1_to_invert_reg[1]/NET0131  ;
  input \sbox1_to_invert_reg[2]/NET0131  ;
  input \sbox1_to_invert_reg[3]/NET0131  ;
  input \state_reg/NET0131  ;
  input \sub1_data_reg_reg[0]/NET0131  ;
  input \sub1_data_reg_reg[100]/NET0131  ;
  input \sub1_data_reg_reg[101]/NET0131  ;
  input \sub1_data_reg_reg[102]/NET0131  ;
  input \sub1_data_reg_reg[103]/NET0131  ;
  input \sub1_data_reg_reg[104]/NET0131  ;
  input \sub1_data_reg_reg[105]/NET0131  ;
  input \sub1_data_reg_reg[106]/NET0131  ;
  input \sub1_data_reg_reg[107]/NET0131  ;
  input \sub1_data_reg_reg[108]/NET0131  ;
  input \sub1_data_reg_reg[109]/NET0131  ;
  input \sub1_data_reg_reg[10]/NET0131  ;
  input \sub1_data_reg_reg[110]/NET0131  ;
  input \sub1_data_reg_reg[111]/NET0131  ;
  input \sub1_data_reg_reg[112]/NET0131  ;
  input \sub1_data_reg_reg[113]/NET0131  ;
  input \sub1_data_reg_reg[114]/NET0131  ;
  input \sub1_data_reg_reg[115]/NET0131  ;
  input \sub1_data_reg_reg[116]/NET0131  ;
  input \sub1_data_reg_reg[117]/NET0131  ;
  input \sub1_data_reg_reg[118]/NET0131  ;
  input \sub1_data_reg_reg[119]/NET0131  ;
  input \sub1_data_reg_reg[11]/NET0131  ;
  input \sub1_data_reg_reg[120]/NET0131  ;
  input \sub1_data_reg_reg[121]/NET0131  ;
  input \sub1_data_reg_reg[122]/NET0131  ;
  input \sub1_data_reg_reg[123]/NET0131  ;
  input \sub1_data_reg_reg[124]/NET0131  ;
  input \sub1_data_reg_reg[125]/NET0131  ;
  input \sub1_data_reg_reg[126]/NET0131  ;
  input \sub1_data_reg_reg[127]/NET0131  ;
  input \sub1_data_reg_reg[12]/NET0131  ;
  input \sub1_data_reg_reg[13]/NET0131  ;
  input \sub1_data_reg_reg[14]/NET0131  ;
  input \sub1_data_reg_reg[15]/NET0131  ;
  input \sub1_data_reg_reg[16]/NET0131  ;
  input \sub1_data_reg_reg[17]/NET0131  ;
  input \sub1_data_reg_reg[18]/NET0131  ;
  input \sub1_data_reg_reg[19]/NET0131  ;
  input \sub1_data_reg_reg[1]/NET0131  ;
  input \sub1_data_reg_reg[20]/NET0131  ;
  input \sub1_data_reg_reg[21]/NET0131  ;
  input \sub1_data_reg_reg[22]/NET0131  ;
  input \sub1_data_reg_reg[23]/NET0131  ;
  input \sub1_data_reg_reg[24]/NET0131  ;
  input \sub1_data_reg_reg[25]/NET0131  ;
  input \sub1_data_reg_reg[26]/NET0131  ;
  input \sub1_data_reg_reg[27]/NET0131  ;
  input \sub1_data_reg_reg[28]/NET0131  ;
  input \sub1_data_reg_reg[29]/NET0131  ;
  input \sub1_data_reg_reg[2]/NET0131  ;
  input \sub1_data_reg_reg[30]/NET0131  ;
  input \sub1_data_reg_reg[31]/NET0131  ;
  input \sub1_data_reg_reg[32]/NET0131  ;
  input \sub1_data_reg_reg[33]/NET0131  ;
  input \sub1_data_reg_reg[34]/NET0131  ;
  input \sub1_data_reg_reg[35]/NET0131  ;
  input \sub1_data_reg_reg[36]/NET0131  ;
  input \sub1_data_reg_reg[37]/NET0131  ;
  input \sub1_data_reg_reg[38]/NET0131  ;
  input \sub1_data_reg_reg[39]/NET0131  ;
  input \sub1_data_reg_reg[3]/NET0131  ;
  input \sub1_data_reg_reg[40]/NET0131  ;
  input \sub1_data_reg_reg[41]/NET0131  ;
  input \sub1_data_reg_reg[42]/NET0131  ;
  input \sub1_data_reg_reg[43]/NET0131  ;
  input \sub1_data_reg_reg[44]/NET0131  ;
  input \sub1_data_reg_reg[45]/NET0131  ;
  input \sub1_data_reg_reg[46]/NET0131  ;
  input \sub1_data_reg_reg[47]/NET0131  ;
  input \sub1_data_reg_reg[48]/NET0131  ;
  input \sub1_data_reg_reg[49]/NET0131  ;
  input \sub1_data_reg_reg[4]/NET0131  ;
  input \sub1_data_reg_reg[50]/NET0131  ;
  input \sub1_data_reg_reg[51]/NET0131  ;
  input \sub1_data_reg_reg[52]/NET0131  ;
  input \sub1_data_reg_reg[53]/NET0131  ;
  input \sub1_data_reg_reg[54]/NET0131  ;
  input \sub1_data_reg_reg[55]/NET0131  ;
  input \sub1_data_reg_reg[56]/NET0131  ;
  input \sub1_data_reg_reg[57]/NET0131  ;
  input \sub1_data_reg_reg[58]/NET0131  ;
  input \sub1_data_reg_reg[59]/NET0131  ;
  input \sub1_data_reg_reg[5]/NET0131  ;
  input \sub1_data_reg_reg[60]/NET0131  ;
  input \sub1_data_reg_reg[61]/NET0131  ;
  input \sub1_data_reg_reg[62]/NET0131  ;
  input \sub1_data_reg_reg[63]/NET0131  ;
  input \sub1_data_reg_reg[64]/NET0131  ;
  input \sub1_data_reg_reg[65]/NET0131  ;
  input \sub1_data_reg_reg[66]/NET0131  ;
  input \sub1_data_reg_reg[67]/NET0131  ;
  input \sub1_data_reg_reg[68]/NET0131  ;
  input \sub1_data_reg_reg[69]/NET0131  ;
  input \sub1_data_reg_reg[6]/NET0131  ;
  input \sub1_data_reg_reg[70]/NET0131  ;
  input \sub1_data_reg_reg[71]/NET0131  ;
  input \sub1_data_reg_reg[72]/NET0131  ;
  input \sub1_data_reg_reg[73]/NET0131  ;
  input \sub1_data_reg_reg[74]/NET0131  ;
  input \sub1_data_reg_reg[75]/NET0131  ;
  input \sub1_data_reg_reg[76]/NET0131  ;
  input \sub1_data_reg_reg[77]/NET0131  ;
  input \sub1_data_reg_reg[78]/NET0131  ;
  input \sub1_data_reg_reg[79]/NET0131  ;
  input \sub1_data_reg_reg[7]/NET0131  ;
  input \sub1_data_reg_reg[80]/NET0131  ;
  input \sub1_data_reg_reg[81]/NET0131  ;
  input \sub1_data_reg_reg[82]/NET0131  ;
  input \sub1_data_reg_reg[83]/NET0131  ;
  input \sub1_data_reg_reg[84]/NET0131  ;
  input \sub1_data_reg_reg[85]/NET0131  ;
  input \sub1_data_reg_reg[86]/NET0131  ;
  input \sub1_data_reg_reg[87]/NET0131  ;
  input \sub1_data_reg_reg[88]/NET0131  ;
  input \sub1_data_reg_reg[89]/NET0131  ;
  input \sub1_data_reg_reg[8]/NET0131  ;
  input \sub1_data_reg_reg[90]/NET0131  ;
  input \sub1_data_reg_reg[91]/NET0131  ;
  input \sub1_data_reg_reg[92]/NET0131  ;
  input \sub1_data_reg_reg[93]/NET0131  ;
  input \sub1_data_reg_reg[94]/NET0131  ;
  input \sub1_data_reg_reg[95]/NET0131  ;
  input \sub1_data_reg_reg[96]/NET0131  ;
  input \sub1_data_reg_reg[97]/NET0131  ;
  input \sub1_data_reg_reg[98]/NET0131  ;
  input \sub1_data_reg_reg[99]/NET0131  ;
  input \sub1_data_reg_reg[9]/NET0131  ;
  input \sub1_ready_o_reg/NET0131  ;
  input \sub1_state_reg[0]/NET0131  ;
  input \sub1_state_reg[1]/NET0131  ;
  input \sub1_state_reg[2]/NET0131  ;
  input \sub1_state_reg[3]/NET0131  ;
  input \sub1_state_reg[4]/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g27929/_0_  ;
  output \g27942/_3_  ;
  output \g27943/_3_  ;
  output \g27944/_3_  ;
  output \g27945/_0_  ;
  output \g27995/_0_  ;
  output \g27998/_0_  ;
  output \g28019/_0_  ;
  output \g28020/_0_  ;
  output \g28021/_0_  ;
  output \g28022/_0_  ;
  output \g28023/_0_  ;
  output \g28024/_0_  ;
  output \g28025/_0_  ;
  output \g28026/_0_  ;
  output \g28027/_0_  ;
  output \g28028/_0_  ;
  output \g28029/_0_  ;
  output \g28030/_0_  ;
  output \g28031/_0_  ;
  output \g28032/_0_  ;
  output \g28033/_0_  ;
  output \g28034/_0_  ;
  output \g28044/_0_  ;
  output \g28045/_0_  ;
  output \g28046/_0_  ;
  output \g28047/_0_  ;
  output \g28048/_0_  ;
  output \g28049/_0_  ;
  output \g28050/_0_  ;
  output \g28051/_0_  ;
  output \g28151/_0_  ;
  output \g28177/_0_  ;
  output \g28178/_0_  ;
  output \g28179/_0_  ;
  output \g28180/_0_  ;
  output \g28181/_0_  ;
  output \g28182/_0_  ;
  output \g28183/_0_  ;
  output \g28184/_0_  ;
  output \g28185/_0_  ;
  output \g28186/_0_  ;
  output \g28187/_0_  ;
  output \g28188/_0_  ;
  output \g28189/_0_  ;
  output \g28190/_0_  ;
  output \g28191/_0_  ;
  output \g28192/_0_  ;
  output \g28193/_0_  ;
  output \g28194/_0_  ;
  output \g28195/_0_  ;
  output \g28196/_0_  ;
  output \g28197/_0_  ;
  output \g28198/_0_  ;
  output \g28199/_0_  ;
  output \g28200/_0_  ;
  output \g28201/_0_  ;
  output \g28202/_0_  ;
  output \g28203/_0_  ;
  output \g28253/_0_  ;
  output \g28254/_0_  ;
  output \g28255/_0_  ;
  output \g28256/_0_  ;
  output \g28257/_0_  ;
  output \g28258/_0_  ;
  output \g28259/_0_  ;
  output \g28260/_0_  ;
  output \g28261/_0_  ;
  output \g28262/_0_  ;
  output \g28263/_0_  ;
  output \g28264/_0_  ;
  output \g28265/_0_  ;
  output \g28266/_0_  ;
  output \g28267/_0_  ;
  output \g28268/_0_  ;
  output \g28269/_0_  ;
  output \g28270/_0_  ;
  output \g28271/_0_  ;
  output \g28272/_0_  ;
  output \g28273/_0_  ;
  output \g28274/_0_  ;
  output \g28275/_0_  ;
  output \g28276/_0_  ;
  output \g28277/_0_  ;
  output \g28278/_0_  ;
  output \g28279/_0_  ;
  output \g28384/_2_  ;
  output \g28385/_2_  ;
  output \g28388/_2_  ;
  output \g28389/_2_  ;
  output \g28394/_2_  ;
  output \g28395/_2_  ;
  output \g28401/_2_  ;
  output \g28402/_2_  ;
  output \g28403/_0_  ;
  output \g28404/_0_  ;
  output \g28408/_0_  ;
  output \g28410/_0_  ;
  output \g28440/_0_  ;
  output \g28441/_0_  ;
  output \g28442/_0_  ;
  output \g28443/_0_  ;
  output \g28444/_0_  ;
  output \g28445/_0_  ;
  output \g28446/_0_  ;
  output \g28447/_0_  ;
  output \g28448/_0_  ;
  output \g28449/_0_  ;
  output \g28450/_0_  ;
  output \g28451/_0_  ;
  output \g28452/_0_  ;
  output \g28453/_0_  ;
  output \g28538/_0_  ;
  output \g28539/_0_  ;
  output \g28540/_0_  ;
  output \g28541/_0_  ;
  output \g28542/_0_  ;
  output \g28543/_0_  ;
  output \g28544/_0_  ;
  output \g28545/_0_  ;
  output \g28546/_0_  ;
  output \g28547/_0_  ;
  output \g28548/_0_  ;
  output \g28549/_0_  ;
  output \g28550/_0_  ;
  output \g28551/_0_  ;
  output \g28552/_0_  ;
  output \g28557/_0_  ;
  output \g28558/_0_  ;
  output \g28563/_0_  ;
  output \g28564/_0_  ;
  output \g28565/_0_  ;
  output \g28566/_0_  ;
  output \g28567/_0_  ;
  output \g28625/_2_  ;
  output \g28626/_2_  ;
  output \g28633/_2_  ;
  output \g28639/_2_  ;
  output \g28655/_2_  ;
  output \g28656/_2_  ;
  output \g28657/_2_  ;
  output \g28660/_2_  ;
  output \g28661/_2_  ;
  output \g28662/_2_  ;
  output \g28666/_2_  ;
  output \g28667/_2_  ;
  output \g28668/_2_  ;
  output \g28678/_2_  ;
  output \g28679/_2_  ;
  output \g28680/_2_  ;
  output \g28690/_0_  ;
  output \g28710/_0_  ;
  output \g28716/_0_  ;
  output \g28795/_0_  ;
  output \g28796/_0_  ;
  output \g28798/_0_  ;
  output \g28799/_0_  ;
  output \g28800/_0_  ;
  output \g28801/_0_  ;
  output \g28804/_0_  ;
  output \g28825/_2_  ;
  output \g28826/_2_  ;
  output \g28830/_2_  ;
  output \g28834/_2_  ;
  output \g28842/_2_  ;
  output \g28843/_2_  ;
  output \g28845/_2_  ;
  output \g28848/_2_  ;
  output \g28890/_0_  ;
  output \g28936/_0_  ;
  output \g28982/_0_  ;
  output \g29050/_0_  ;
  output \g29051/_0_  ;
  output \g29052/_0_  ;
  output \g29053/_0_  ;
  output \g29054/_0_  ;
  output \g29055/_0_  ;
  output \g29056/_0_  ;
  output \g29057/_0_  ;
  output \g29058/_0_  ;
  output \g29059/_0_  ;
  output \g29060/_0_  ;
  output \g29061/_0_  ;
  output \g29328/_0_  ;
  output \g29329/_0_  ;
  output \g29330/_0_  ;
  output \g29331/_0_  ;
  output \g29332/_0_  ;
  output \g29333/_0_  ;
  output \g29334/_0_  ;
  output \g29335/_0_  ;
  output \g29336/_0_  ;
  output \g29337/_0_  ;
  output \g29338/_0_  ;
  output \g29339/_0_  ;
  output \g29340/_0_  ;
  output \g29341/_0_  ;
  output \g29342/_0_  ;
  output \g29343/_0_  ;
  output \g29344/_0_  ;
  output \g29345/_0_  ;
  output \g29346/_0_  ;
  output \g29347/_0_  ;
  output \g29348/_0_  ;
  output \g29349/_0_  ;
  output \g29350/_0_  ;
  output \g29351/_0_  ;
  output \g29352/_0_  ;
  output \g29353/_0_  ;
  output \g29354/_0_  ;
  output \g29355/_0_  ;
  output \g29356/_0_  ;
  output \g29357/_0_  ;
  output \g29358/_0_  ;
  output \g29359/_0_  ;
  output \g29360/_0_  ;
  output \g29361/_0_  ;
  output \g29362/_0_  ;
  output \g29363/_0_  ;
  output \g29364/_0_  ;
  output \g29365/_0_  ;
  output \g29366/_0_  ;
  output \g29367/_0_  ;
  output \g29395/_0_  ;
  output \g29396/_0_  ;
  output \g29453/_0_  ;
  output \g29454/_0_  ;
  output \g29455/_0_  ;
  output \g29456/_0_  ;
  output \g29457/_0_  ;
  output \g29458/_0_  ;
  output \g29459/_0_  ;
  output \g29460/_0_  ;
  output \g29461/_0_  ;
  output \g29462/_0_  ;
  output \g29463/_0_  ;
  output \g29464/_0_  ;
  output \g29465/_0_  ;
  output \g29466/_0_  ;
  output \g29467/_0_  ;
  output \g29468/_0_  ;
  output \g29469/_0_  ;
  output \g29470/_0_  ;
  output \g29471/_0_  ;
  output \g29472/_0_  ;
  output \g29473/_0_  ;
  output \g29474/_0_  ;
  output \g29475/_0_  ;
  output \g29476/_0_  ;
  output \g29477/_0_  ;
  output \g29478/_0_  ;
  output \g29479/_0_  ;
  output \g29480/_0_  ;
  output \g29481/_0_  ;
  output \g29482/_0_  ;
  output \g29483/_0_  ;
  output \g29484/_0_  ;
  output \g29485/_0_  ;
  output \g29486/_0_  ;
  output \g29487/_0_  ;
  output \g29488/_0_  ;
  output \g29489/_0_  ;
  output \g29490/_0_  ;
  output \g29491/_0_  ;
  output \g29492/_0_  ;
  output \g29493/_0_  ;
  output \g29494/_0_  ;
  output \g29495/_0_  ;
  output \g29496/_0_  ;
  output \g29497/_0_  ;
  output \g29498/_0_  ;
  output \g29499/_0_  ;
  output \g29500/_0_  ;
  output \g29501/_0_  ;
  output \g29502/_0_  ;
  output \g29503/_0_  ;
  output \g29504/_0_  ;
  output \g29505/_0_  ;
  output \g29506/_0_  ;
  output \g29507/_0_  ;
  output \g29508/_0_  ;
  output \g29509/_0_  ;
  output \g29510/_0_  ;
  output \g29511/_0_  ;
  output \g29512/_0_  ;
  output \g29513/_0_  ;
  output \g29514/_0_  ;
  output \g29515/_0_  ;
  output \g29516/_0_  ;
  output \g29517/_0_  ;
  output \g29518/_0_  ;
  output \g29519/_0_  ;
  output \g29520/_0_  ;
  output \g29521/_0_  ;
  output \g29522/_0_  ;
  output \g29523/_0_  ;
  output \g29524/_0_  ;
  output \g29525/_0_  ;
  output \g29526/_0_  ;
  output \g29527/_0_  ;
  output \g29528/_0_  ;
  output \g29529/_0_  ;
  output \g29530/_0_  ;
  output \g29531/_0_  ;
  output \g29532/_0_  ;
  output \g29533/_0_  ;
  output \g29534/_0_  ;
  output \g29535/_0_  ;
  output \g29536/_0_  ;
  output \g29537/_0_  ;
  output \g29538/_0_  ;
  output \g29539/_0_  ;
  output \g29540/_0_  ;
  output \g29541/_0_  ;
  output \g29542/_0_  ;
  output \g29543/_0_  ;
  output \g29544/_0_  ;
  output \g29545/_0_  ;
  output \g29546/_0_  ;
  output \g29547/_0_  ;
  output \g29548/_0_  ;
  output \g29549/_0_  ;
  output \g29550/_0_  ;
  output \g29551/_0_  ;
  output \g29552/_0_  ;
  output \g29553/_0_  ;
  output \g29554/_0_  ;
  output \g29555/_0_  ;
  output \g29556/_0_  ;
  output \g29557/_0_  ;
  output \g29558/_0_  ;
  output \g29559/_0_  ;
  output \g29560/_0_  ;
  output \g29561/_0_  ;
  output \g29562/_0_  ;
  output \g29563/_0_  ;
  output \g29564/_0_  ;
  output \g29565/_0_  ;
  output \g29566/_0_  ;
  output \g29567/_0_  ;
  output \g29568/_0_  ;
  output \g29569/_0_  ;
  output \g29570/_0_  ;
  output \g29571/_0_  ;
  output \g29572/_0_  ;
  output \g29573/_0_  ;
  output \g29574/_0_  ;
  output \g29575/_0_  ;
  output \g29576/_0_  ;
  output \g29577/_0_  ;
  output \g29578/_0_  ;
  output \g29579/_0_  ;
  output \g29580/_0_  ;
  output \g29582/_0_  ;
  output \g29583/_0_  ;
  output \g29584/_0_  ;
  output \g29585/_0_  ;
  output \g29586/_0_  ;
  output \g29587/_0_  ;
  output \g29588/_0_  ;
  output \g29589/_0_  ;
  output \g29590/_0_  ;
  output \g29591/_0_  ;
  output \g29592/_0_  ;
  output \g29593/_0_  ;
  output \g29634/_0_  ;
  output \g29635/_0_  ;
  output \g29636/_0_  ;
  output \g29637/_0_  ;
  output \g29645/_0_  ;
  output \g29646/_0_  ;
  output \g29647/_0_  ;
  output \g29824/_0_  ;
  output \g29828/_0_  ;
  output \g29832/_0_  ;
  output \g29836/_0_  ;
  output \g29837/_0_  ;
  output \g29838/_0_  ;
  output \g29839/_0_  ;
  output \g29840/_0_  ;
  output \g29841/_0_  ;
  output \g29842/_0_  ;
  output \g29843/_0_  ;
  output \g29844/_0_  ;
  output \g29845/_0_  ;
  output \g29846/_0_  ;
  output \g29847/_0_  ;
  output \g29848/_0_  ;
  output \g29849/_0_  ;
  output \g29850/_0_  ;
  output \g29851/_0_  ;
  output \g29852/_0_  ;
  output \g29853/_0_  ;
  output \g29854/_0_  ;
  output \g29855/_0_  ;
  output \g29856/_0_  ;
  output \g29857/_0_  ;
  output \g29858/_0_  ;
  output \g29859/_0_  ;
  output \g29860/_0_  ;
  output \g29861/_0_  ;
  output \g29862/_0_  ;
  output \g29863/_0_  ;
  output \g29864/_0_  ;
  output \g29865/_0_  ;
  output \g29866/_0_  ;
  output \g29867/_0_  ;
  output \g29868/_0_  ;
  output \g30081/_0_  ;
  output \g30082/_0_  ;
  output \g30083/_0_  ;
  output \g30084/_0_  ;
  output \g30085/_0_  ;
  output \g30086/_0_  ;
  output \g30087/_0_  ;
  output \g30088/_0_  ;
  output \g30089/_0_  ;
  output \g30090/_0_  ;
  output \g30091/_0_  ;
  output \g30092/_0_  ;
  output \g30093/_0_  ;
  output \g30094/_0_  ;
  output \g30095/_0_  ;
  output \g30096/_0_  ;
  output \g30135/_0_  ;
  output \g30137/_0_  ;
  output \g30164/_0_  ;
  output \g30165/_0_  ;
  output \g30166/_0_  ;
  output \g30167/_0_  ;
  output \g30168/_0_  ;
  output \g30169/_0_  ;
  output \g30170/_0_  ;
  output \g30231/_0_  ;
  output \g30232/_0_  ;
  output \g30233/_0_  ;
  output \g30234/_0_  ;
  output \g30235/_0_  ;
  output \g30236/_0_  ;
  output \g30237/_0_  ;
  output \g30238/_0_  ;
  output \g30286/_0_  ;
  output \g30287/_0_  ;
  output \g30288/_0_  ;
  output \g30289/_0_  ;
  output \g30290/_0_  ;
  output \g30291/_0_  ;
  output \g30292/_0_  ;
  output \g30293/_0_  ;
  output \g30294/_0_  ;
  output \g30295/_0_  ;
  output \g30296/_0_  ;
  output \g30297/_0_  ;
  output \g30298/_0_  ;
  output \g30299/_0_  ;
  output \g30300/_0_  ;
  output \g30301/_0_  ;
  output \g30303/_0_  ;
  output \g30304/_0_  ;
  output \g30305/_0_  ;
  output \g30306/_0_  ;
  output \g30307/_0_  ;
  output \g30308/_0_  ;
  output \g30309/_0_  ;
  output \g30310/_0_  ;
  output \g30311/_0_  ;
  output \g30312/_0_  ;
  output \g30313/_0_  ;
  output \g30314/_0_  ;
  output \g30315/_0_  ;
  output \g30316/_0_  ;
  output \g30317/_0_  ;
  output \g30318/_0_  ;
  output \g30319/_0_  ;
  output \g30481/_0_  ;
  output \g30482/_0_  ;
  output \g30483/_0_  ;
  output \g30484/_0_  ;
  output \g30493/_0_  ;
  output \g30495/_0_  ;
  output \g30536/_0_  ;
  output \g30537/_0_  ;
  output \g30538/_0_  ;
  output \g30735/_0_  ;
  output \g30927/_0_  ;
  output \g30928/_0_  ;
  output \g30929/_0_  ;
  output \g30971/_0_  ;
  output \g30972/_0_  ;
  output \g30973/_0_  ;
  output \g30974/_0_  ;
  output \g31129/_0_  ;
  output \g31130/_0_  ;
  output \g31131/_0_  ;
  output \g31132/_0_  ;
  output \g31133/_0_  ;
  output \g31134/_0_  ;
  output \g31135/_0_  ;
  output \g31136/_0_  ;
  output \g31137/_0_  ;
  output \g31138/_0_  ;
  output \g31139/_0_  ;
  output \g31140/_0_  ;
  output \g31141/_0_  ;
  output \g31142/_0_  ;
  output \g31143/_0_  ;
  output \g31144/_0_  ;
  output \g31352/_0_  ;
  output \g31353/_0_  ;
  output \g31354/_0_  ;
  output \g31355/_0_  ;
  output \g31356/_0_  ;
  output \g31357/_0_  ;
  output \g31358/_0_  ;
  output \g31359/_0_  ;
  output \g31360/_0_  ;
  output \g31361/_0_  ;
  output \g31362/_0_  ;
  output \g31363/_0_  ;
  output \g31364/_0_  ;
  output \g31365/_0_  ;
  output \g31366/_0_  ;
  output \g31367/_0_  ;
  output \g31706/_0_  ;
  output \g32001/_0_  ;
  output \g32008/_0_  ;
  output \g32009/_0_  ;
  output \g32010/_0_  ;
  output \g32011/_0_  ;
  output \g32118/_0_  ;
  output \g33261/_0_  ;
  output \g33262/_0_  ;
  output \g33263/_0_  ;
  output \g33264/_0_  ;
  output \g33265/_0_  ;
  output \g33266/_0_  ;
  output \g33450/_0_  ;
  output \g33451/_0_  ;
  output \g33453/_0_  ;
  output \g33485/_0_  ;
  output \g33679/_2_  ;
  output \g34838/_2_  ;
  output \g34971/_0_  ;
  output \g34972/_0_  ;
  output \g34973/_0_  ;
  output \g34974/_0_  ;
  output \g34975/_0_  ;
  output \g34976/_0_  ;
  output \g34977/_0_  ;
  output \g34978/_0_  ;
  output \g34979/_0_  ;
  output \g34980/_0_  ;
  output \g34981/_0_  ;
  output \g34982/_0_  ;
  output \g34983/_0_  ;
  output \g34984/_0_  ;
  output \g34985/_0_  ;
  output \g34986/_0_  ;
  output \g34987/_0_  ;
  output \g34988/_0_  ;
  output \g34989/_0_  ;
  output \g34990/_0_  ;
  output \g34991/_0_  ;
  output \g34992/_0_  ;
  output \g34993/_0_  ;
  output \g34994/_0_  ;
  output \g34995/_0_  ;
  output \g34996/_0_  ;
  output \g34997/_0_  ;
  output \g34998/_0_  ;
  output \g34999/_0_  ;
  output \g35000/_0_  ;
  output \g35001/_0_  ;
  output \g35002/_0_  ;
  output \g35003/_0_  ;
  output \g35004/_0_  ;
  output \g35005/_0_  ;
  output \g35006/_0_  ;
  output \g35007/_0_  ;
  output \g35008/_0_  ;
  output \g35009/_0_  ;
  output \g35010/_0_  ;
  output \g35011/_0_  ;
  output \g35012/_0_  ;
  output \g35013/_0_  ;
  output \g35014/_0_  ;
  output \g35015/_0_  ;
  output \g35016/_0_  ;
  output \g35017/_0_  ;
  output \g35018/_0_  ;
  output \g35019/_0_  ;
  output \g35020/_0_  ;
  output \g35021/_0_  ;
  output \g35022/_0_  ;
  output \g35023/_0_  ;
  output \g35024/_0_  ;
  output \g35025/_0_  ;
  output \g35026/_0_  ;
  output \g35027/_0_  ;
  output \g35028/_0_  ;
  output \g35029/_0_  ;
  output \g35030/_0_  ;
  output \g35031/_0_  ;
  output \g35032/_0_  ;
  output \g35033/_0_  ;
  output \g35034/_0_  ;
  output \g35035/_0_  ;
  output \g35036/_0_  ;
  output \g35037/_0_  ;
  output \g35038/_0_  ;
  output \g35039/_0_  ;
  output \g35040/_0_  ;
  output \g35041/_0_  ;
  output \g35042/_0_  ;
  output \g35043/_0_  ;
  output \g35044/_0_  ;
  output \g35045/_0_  ;
  output \g35046/_0_  ;
  output \g35047/_0_  ;
  output \g35048/_0_  ;
  output \g35049/_0_  ;
  output \g35050/_0_  ;
  output \g35051/_0_  ;
  output \g35052/_0_  ;
  output \g35053/_0_  ;
  output \g35054/_0_  ;
  output \g35055/_0_  ;
  output \g35056/_0_  ;
  output \g35057/_0_  ;
  output \g35058/_0_  ;
  output \g35059/_0_  ;
  output \g35060/_0_  ;
  output \g35061/_0_  ;
  output \g35062/_0_  ;
  output \g35063/_0_  ;
  output \g35064/_0_  ;
  output \g35065/_0_  ;
  output \g35066/_0_  ;
  output \g35538/_0_  ;
  output \g35956/_0_  ;
  output \g36298/_1_  ;
  output \g36324/_0_  ;
  output \g36375/_0_  ;
  output \g38269/_0_  ;
  output \g38473/_0_  ;
  output \g38501/_0_  ;
  output \g38569/_0_  ;
  output \g38629/_0_  ;
  output \g38721_dup/_3_  ;
  output \g38735/_0_  ;
  output \g38753/_0_  ;
  output \g38849/_3_  ;
  output \g39071/_0_  ;
  output \g39073/_0_  ;
  output \g39077/_0_  ;
  output \g39080/_0_  ;
  output \g39135/_0_  ;
  output \g39138/_0_  ;
  output \g39182/_0_  ;
  output \g39197/_3_  ;
  output \g39207/_3_  ;
  output \g39241/_0_  ;
  output \g39272/_0_  ;
  output \g39307/_0_  ;
  output \g39308/_0_  ;
  output \g39361/_0_  ;
  output \g39494/_0_  ;
  output \g39558/_0_  ;
  output \g39575/_0_  ;
  output \g39583/_0_  ;
  wire n928 , n929 , n930 , n931 , n932 , n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 , n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 , n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 , n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 , n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 , n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 , n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 , n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 , n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 , n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 , n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 , n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 , n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 , n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 , n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 , n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 , n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 , n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 , n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 , n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 , n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 , n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 , n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 , n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 , n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 , n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 , n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 , n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 , n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 , n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 , n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 , n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 , n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 , n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 , n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 , n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 , n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 , n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 , n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 , n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 , n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 , n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 , n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 , n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 , n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 , n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 , n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 , n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 , n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 , n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 , n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 , n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 , n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 , n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 , n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 , n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 , n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 , n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 , n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 , n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 , n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 , n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 , n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 , n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 , n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 , n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 , n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 , n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 , n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 , n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 , n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 , n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 , n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 , n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 , n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 , n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 , n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 , n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 , n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 , n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 , n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 , n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 , n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 , n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 , n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 , n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 , n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 , n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 , n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 , n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 , n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 , n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 , n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 , n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 , n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 , n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 , n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 , n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 , n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 , n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 , n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 , n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 , n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 , n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 , n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 , n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 , n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 , n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 , n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 , n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 , n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 , n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 , n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 , n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 , n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 , n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 , n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 , n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 , n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 , n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 , n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 , n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 , n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 , n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 , n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 , n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 , n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 , n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 , n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 , n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 , n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 , n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 , n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 , n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 , n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 , n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 , n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 , n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 , n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 , n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 , n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 , n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 , n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 , n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 , n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 , n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 , n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 , n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 , n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 , n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 , n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 , n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 , n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 , n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 , n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 , n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 , n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 , n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 , n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 , n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 , n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 , n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 , n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 , n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 , n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 , n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 , n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 , n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 , n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 , n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 , n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 , n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 , n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 , n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 , n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 , n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 , n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 , n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 , n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 , n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 , n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 , n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 , n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 , n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 , n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 , n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 , n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 , n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 , n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 , n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 , n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 , n10273 , n10274 , n10275 ;
  assign n928 = ~\ks1_state_reg[0]/NET0131  & ~\ks1_state_reg[1]/NET0131  ;
  assign n929 = \ks1_state_reg[2]/NET0131  & n928 ;
  assign n930 = ~\round_reg[0]/NET0131  & ~\round_reg[1]/NET0131  ;
  assign n931 = ~\round_reg[2]/NET0131  & ~\round_reg[3]/NET0131  ;
  assign n932 = n930 & n931 ;
  assign n933 = \addroundkey_start_i_reg/NET0131  & n932 ;
  assign n936 = ~\addroundkey_round_reg[0]/NET0131  & ~\round_reg[0]/NET0131  ;
  assign n937 = \addroundkey_round_reg[0]/NET0131  & \round_reg[0]/NET0131  ;
  assign n938 = ~n936 & ~n937 ;
  assign n934 = \addroundkey_round_reg[2]/NET0131  & ~\round_reg[2]/NET0131  ;
  assign n935 = ~\addroundkey_round_reg[2]/NET0131  & \round_reg[2]/NET0131  ;
  assign n945 = ~n934 & ~n935 ;
  assign n946 = ~n938 & n945 ;
  assign n939 = ~\addroundkey_round_reg[1]/NET0131  & ~\round_reg[1]/NET0131  ;
  assign n940 = \addroundkey_round_reg[1]/NET0131  & \round_reg[1]/NET0131  ;
  assign n941 = ~n939 & ~n940 ;
  assign n942 = ~\addroundkey_round_reg[3]/NET0131  & ~\round_reg[3]/NET0131  ;
  assign n943 = \addroundkey_round_reg[3]/NET0131  & \round_reg[3]/NET0131  ;
  assign n944 = ~n942 & ~n943 ;
  assign n947 = ~n941 & ~n944 ;
  assign n948 = n946 & n947 ;
  assign n949 = \ks1_ready_o_reg/NET0131  & ~n948 ;
  assign n950 = ~\addroundkey_round_reg[1]/NET0131  & ~\addroundkey_round_reg[2]/NET0131  ;
  assign n951 = ~\addroundkey_round_reg[3]/NET0131  & n950 ;
  assign n952 = ~n949 & n951 ;
  assign n953 = ~\addroundkey_start_i_reg/NET0131  & ~n952 ;
  assign n954 = \key_i[14]_pad  & ~n953 ;
  assign n955 = \addroundkey_start_i_reg/NET0131  & ~n932 ;
  assign n956 = ~n952 & ~n955 ;
  assign n957 = \ks1_key_reg_reg[14]/NET0131  & n956 ;
  assign n958 = ~n954 & ~n957 ;
  assign n959 = ~n933 & ~n958 ;
  assign n961 = ~\key_i[14]_pad  & n951 ;
  assign n960 = ~\ks1_key_reg_reg[14]/NET0131  & ~n951 ;
  assign n962 = n933 & ~n960 ;
  assign n963 = ~n961 & n962 ;
  assign n964 = ~n959 & ~n963 ;
  assign n967 = ~\addroundkey_start_i_reg/NET0131  & \ks1_ready_o_reg/NET0131  ;
  assign n968 = ~n948 & n967 ;
  assign n969 = ~n955 & ~n968 ;
  assign n966 = ~\ks1_state_reg[0]/NET0131  & ~\ks1_state_reg[2]/NET0131  ;
  assign n970 = ~\ks1_state_reg[1]/NET0131  & n966 ;
  assign n971 = ~n969 & n970 ;
  assign n965 = ~\ks1_state_reg[2]/NET0131  & ~n928 ;
  assign n972 = ~n929 & ~n965 ;
  assign n973 = ~n971 & n972 ;
  assign n974 = decrypt_i_pad & n973 ;
  assign n975 = \sbox1_to_invert_reg[1]/NET0131  & \sbox1_to_invert_reg[2]/NET0131  ;
  assign n976 = \sbox1_to_invert_reg[0]/NET0131  & \sbox1_to_invert_reg[3]/NET0131  ;
  assign n977 = ~n975 & n976 ;
  assign n978 = ~\sbox1_to_invert_reg[1]/NET0131  & ~\sbox1_to_invert_reg[2]/NET0131  ;
  assign n979 = ~\sbox1_to_invert_reg[3]/NET0131  & n978 ;
  assign n980 = ~n975 & ~n979 ;
  assign n981 = ~n976 & ~n980 ;
  assign n982 = ~n977 & ~n981 ;
  assign n983 = \sbox1_ah_reg_reg[1]/NET0131  & n982 ;
  assign n984 = \sbox1_to_invert_reg[3]/NET0131  & ~n978 ;
  assign n985 = ~n979 & ~n984 ;
  assign n986 = ~n975 & ~n985 ;
  assign n987 = ~\sbox1_to_invert_reg[1]/NET0131  & \sbox1_to_invert_reg[2]/NET0131  ;
  assign n988 = \sbox1_to_invert_reg[0]/NET0131  & ~n987 ;
  assign n989 = ~n986 & ~n988 ;
  assign n990 = \sbox1_to_invert_reg[0]/NET0131  & ~\sbox1_to_invert_reg[2]/NET0131  ;
  assign n991 = n986 & n990 ;
  assign n992 = ~n989 & ~n991 ;
  assign n993 = \sbox1_ah_reg_reg[0]/NET0131  & ~n992 ;
  assign n994 = ~\sbox1_to_invert_reg[1]/NET0131  & \sbox1_to_invert_reg[3]/NET0131  ;
  assign n995 = ~\sbox1_to_invert_reg[0]/NET0131  & ~n975 ;
  assign n996 = ~n994 & n995 ;
  assign n997 = n976 & ~n978 ;
  assign n998 = ~n979 & ~n997 ;
  assign n999 = ~n996 & n998 ;
  assign n1000 = \sbox1_ah_reg_reg[3]/NET0131  & n999 ;
  assign n1001 = \sbox1_to_invert_reg[3]/NET0131  & ~n990 ;
  assign n1002 = \sbox1_to_invert_reg[0]/NET0131  & ~\sbox1_to_invert_reg[1]/NET0131  ;
  assign n1003 = ~\sbox1_to_invert_reg[0]/NET0131  & ~\sbox1_to_invert_reg[2]/NET0131  ;
  assign n1004 = ~n1002 & ~n1003 ;
  assign n1005 = n1001 & ~n1004 ;
  assign n1006 = ~n1001 & n1004 ;
  assign n1007 = ~n1005 & ~n1006 ;
  assign n1008 = \sbox1_ah_reg_reg[2]/NET0131  & ~n1007 ;
  assign n1009 = n1000 & ~n1008 ;
  assign n1010 = ~n1000 & n1008 ;
  assign n1011 = ~n1009 & ~n1010 ;
  assign n1012 = n993 & n1011 ;
  assign n1013 = ~n993 & ~n1011 ;
  assign n1014 = ~n1012 & ~n1013 ;
  assign n1015 = n983 & ~n1014 ;
  assign n1016 = ~n983 & n1014 ;
  assign n1017 = ~n1015 & ~n1016 ;
  assign n1018 = \sbox1_ah_reg_reg[2]/NET0131  & n999 ;
  assign n1019 = \sbox1_ah_reg_reg[1]/NET0131  & ~n1007 ;
  assign n1020 = \sbox1_ah_reg_reg[3]/NET0131  & ~n992 ;
  assign n1021 = n1019 & ~n1020 ;
  assign n1022 = ~n1019 & n1020 ;
  assign n1023 = ~n1021 & ~n1022 ;
  assign n1024 = \sbox1_ah_reg_reg[0]/NET0131  & ~\sbox1_ah_reg_reg[3]/NET0131  ;
  assign n1025 = ~\sbox1_ah_reg_reg[0]/NET0131  & \sbox1_ah_reg_reg[3]/NET0131  ;
  assign n1026 = ~n1024 & ~n1025 ;
  assign n1027 = n982 & ~n1026 ;
  assign n1028 = n1023 & ~n1027 ;
  assign n1029 = ~n1023 & n1027 ;
  assign n1030 = ~n1028 & ~n1029 ;
  assign n1031 = n1018 & n1030 ;
  assign n1032 = ~n1018 & ~n1030 ;
  assign n1033 = ~n1031 & ~n1032 ;
  assign n1034 = ~n982 & n1007 ;
  assign n1035 = n982 & ~n1007 ;
  assign n1036 = ~n1034 & ~n1035 ;
  assign n1037 = \sbox1_ah_reg_reg[3]/NET0131  & n1036 ;
  assign n1038 = n982 & ~n992 ;
  assign n1039 = ~n982 & n992 ;
  assign n1040 = ~n1038 & ~n1039 ;
  assign n1041 = \sbox1_ah_reg_reg[2]/NET0131  & n1040 ;
  assign n1042 = \sbox1_ah_reg_reg[0]/NET0131  & ~n1007 ;
  assign n1043 = \sbox1_ah_reg_reg[1]/NET0131  & n999 ;
  assign n1044 = n1042 & ~n1043 ;
  assign n1045 = ~n1042 & n1043 ;
  assign n1046 = ~n1044 & ~n1045 ;
  assign n1047 = n1041 & ~n1046 ;
  assign n1048 = ~n1041 & n1046 ;
  assign n1049 = ~n1047 & ~n1048 ;
  assign n1050 = n1037 & n1049 ;
  assign n1051 = ~n1037 & ~n1049 ;
  assign n1052 = ~n1050 & ~n1051 ;
  assign n1053 = n1033 & ~n1052 ;
  assign n1054 = ~n1033 & n1052 ;
  assign n1055 = ~n1053 & ~n1054 ;
  assign n1056 = n1017 & n1055 ;
  assign n1057 = ~n1017 & ~n1055 ;
  assign n1058 = ~n1056 & ~n1057 ;
  assign n1059 = ~n974 & n1058 ;
  assign n1060 = \sbox1_alph_reg[2]/NET0131  & n1040 ;
  assign n1061 = \sbox1_alph_reg[1]/NET0131  & n999 ;
  assign n1062 = \sbox1_alph_reg[3]/NET0131  & n1036 ;
  assign n1063 = \sbox1_alph_reg[0]/NET0131  & ~n1007 ;
  assign n1064 = n1062 & ~n1063 ;
  assign n1065 = ~n1062 & n1063 ;
  assign n1066 = ~n1064 & ~n1065 ;
  assign n1067 = n1061 & ~n1066 ;
  assign n1068 = ~n1061 & n1066 ;
  assign n1069 = ~n1067 & ~n1068 ;
  assign n1070 = n1060 & n1069 ;
  assign n1071 = ~n1060 & ~n1069 ;
  assign n1072 = ~n1070 & ~n1071 ;
  assign n1073 = n1033 & n1072 ;
  assign n1074 = ~n1033 & ~n1072 ;
  assign n1075 = ~n1073 & ~n1074 ;
  assign n1076 = \sbox1_alph_reg[2]/NET0131  & n1036 ;
  assign n1077 = \sbox1_alph_reg[1]/NET0131  & n1040 ;
  assign n1078 = n1076 & ~n1077 ;
  assign n1079 = ~n1076 & n1077 ;
  assign n1080 = ~n1078 & ~n1079 ;
  assign n1081 = ~\sbox1_alph_reg[0]/NET0131  & n999 ;
  assign n1082 = \sbox1_alph_reg[3]/NET0131  & n1007 ;
  assign n1083 = ~n1081 & n1082 ;
  assign n1084 = ~\sbox1_alph_reg[3]/NET0131  & ~n999 ;
  assign n1085 = ~n1081 & ~n1084 ;
  assign n1086 = ~n1082 & ~n1085 ;
  assign n1087 = ~n1083 & ~n1086 ;
  assign n1088 = n1080 & ~n1087 ;
  assign n1089 = ~n1080 & n1087 ;
  assign n1090 = ~n1088 & ~n1089 ;
  assign n1091 = \sbox1_alph_reg[0]/NET0131  & n982 ;
  assign n1092 = \sbox1_alph_reg[3]/NET0131  & n1040 ;
  assign n1093 = \sbox1_alph_reg[2]/NET0131  & n999 ;
  assign n1094 = \sbox1_alph_reg[1]/NET0131  & ~n1007 ;
  assign n1095 = n1093 & ~n1094 ;
  assign n1096 = ~n1093 & n1094 ;
  assign n1097 = ~n1095 & ~n1096 ;
  assign n1098 = n1092 & ~n1097 ;
  assign n1099 = ~n1092 & n1097 ;
  assign n1100 = ~n1098 & ~n1099 ;
  assign n1101 = n1091 & ~n1100 ;
  assign n1102 = ~n1091 & n1100 ;
  assign n1103 = ~n1101 & ~n1102 ;
  assign n1104 = n1090 & n1103 ;
  assign n1105 = ~n1090 & ~n1103 ;
  assign n1106 = ~n1104 & ~n1105 ;
  assign n1107 = n1075 & n1106 ;
  assign n1108 = ~n1075 & ~n1106 ;
  assign n1109 = ~n1107 & ~n1108 ;
  assign n1111 = n1017 & ~n1109 ;
  assign n1110 = ~n1017 & n1109 ;
  assign n1112 = n974 & ~n1110 ;
  assign n1113 = ~n1111 & n1112 ;
  assign n1114 = ~n1059 & ~n1113 ;
  assign n1115 = n951 & ~n968 ;
  assign n1116 = ~n955 & ~n1115 ;
  assign n1117 = ~\ks1_key_reg_reg[110]/P0002  & n1116 ;
  assign n1118 = ~\key_i[110]_pad  & ~n1116 ;
  assign n1119 = ~n1117 & ~n1118 ;
  assign n1120 = n1114 & ~n1119 ;
  assign n1121 = ~n1114 & n1119 ;
  assign n1122 = ~n1120 & ~n1121 ;
  assign n1123 = ~\ks1_key_reg_reg[78]/P0002  & n1116 ;
  assign n1124 = ~\key_i[78]_pad  & ~n1116 ;
  assign n1125 = ~n1123 & ~n1124 ;
  assign n1126 = n1122 & ~n1125 ;
  assign n1127 = ~n1122 & n1125 ;
  assign n1128 = ~n1126 & ~n1127 ;
  assign n1129 = ~\ks1_key_reg_reg[46]/P0002  & n1116 ;
  assign n1130 = ~\key_i[46]_pad  & ~n1116 ;
  assign n1131 = ~n1129 & ~n1130 ;
  assign n1132 = n1128 & ~n1131 ;
  assign n1133 = ~n1128 & n1131 ;
  assign n1134 = ~n1132 & ~n1133 ;
  assign n1135 = n964 & ~n1134 ;
  assign n1136 = ~n964 & n1134 ;
  assign n1137 = ~n1135 & ~n1136 ;
  assign n1138 = n929 & ~n1137 ;
  assign n1139 = ~\ks1_key_reg_reg[14]/NET0131  & ~n929 ;
  assign n1140 = ~n1138 & ~n1139 ;
  assign n1156 = ~\round_reg[2]/NET0131  & \round_reg[3]/NET0131  ;
  assign n1157 = ~\round_reg[0]/NET0131  & \round_reg[1]/NET0131  ;
  assign n1158 = n1156 & n1157 ;
  assign n1159 = decrypt_i_pad & ~n1158 ;
  assign n1186 = ~\mix1_data_o_reg_reg[60]/NET0131  & n1159 ;
  assign n1171 = ~\sub1_state_reg[0]/NET0131  & ~\sub1_state_reg[1]/NET0131  ;
  assign n1183 = ~\sub1_state_reg[2]/NET0131  & n1171 ;
  assign n1184 = \sub1_state_reg[3]/NET0131  & n1183 ;
  assign n1185 = ~\data_o[60]_pad  & ~n1159 ;
  assign n1187 = n1184 & ~n1185 ;
  assign n1188 = ~n1186 & n1187 ;
  assign n1191 = ~\mix1_data_o_reg_reg[116]/NET0131  & n1159 ;
  assign n1164 = ~\sub1_state_reg[2]/NET0131  & ~\sub1_state_reg[3]/NET0131  ;
  assign n1177 = \sub1_state_reg[0]/NET0131  & ~\sub1_state_reg[1]/NET0131  ;
  assign n1189 = n1164 & n1177 ;
  assign n1190 = ~\data_o[116]_pad  & ~n1159 ;
  assign n1192 = n1189 & ~n1190 ;
  assign n1193 = ~n1191 & n1192 ;
  assign n1244 = ~n1188 & ~n1193 ;
  assign n1197 = ~\mix1_data_o_reg_reg[44]/NET0131  & n1159 ;
  assign n1153 = ~\sub1_state_reg[0]/NET0131  & \sub1_state_reg[1]/NET0131  ;
  assign n1194 = ~\sub1_state_reg[2]/NET0131  & \sub1_state_reg[3]/NET0131  ;
  assign n1195 = n1153 & n1194 ;
  assign n1196 = ~\data_o[44]_pad  & ~n1159 ;
  assign n1198 = n1195 & ~n1196 ;
  assign n1199 = ~n1197 & n1198 ;
  assign n1203 = ~\mix1_data_o_reg_reg[4]/NET0131  & n1159 ;
  assign n1165 = \sub1_state_reg[0]/NET0131  & \sub1_state_reg[1]/NET0131  ;
  assign n1200 = \sub1_state_reg[2]/NET0131  & n1165 ;
  assign n1201 = \sub1_state_reg[3]/NET0131  & n1200 ;
  assign n1202 = ~\data_o[4]_pad  & ~n1159 ;
  assign n1204 = n1201 & ~n1202 ;
  assign n1205 = ~n1203 & n1204 ;
  assign n1245 = ~n1199 & ~n1205 ;
  assign n1251 = n1244 & n1245 ;
  assign n1161 = ~\mix1_data_o_reg_reg[12]/NET0131  & n1159 ;
  assign n1154 = \sub1_state_reg[2]/NET0131  & \sub1_state_reg[3]/NET0131  ;
  assign n1155 = n1153 & n1154 ;
  assign n1160 = ~\data_o[12]_pad  & ~n1159 ;
  assign n1162 = n1155 & ~n1160 ;
  assign n1163 = ~n1161 & n1162 ;
  assign n1168 = ~\mix1_data_o_reg_reg[100]/NET0131  & n1159 ;
  assign n1166 = n1164 & n1165 ;
  assign n1167 = ~\data_o[100]_pad  & ~n1159 ;
  assign n1169 = n1166 & ~n1167 ;
  assign n1170 = ~n1168 & n1169 ;
  assign n1242 = ~n1163 & ~n1170 ;
  assign n1174 = ~\mix1_data_o_reg_reg[28]/NET0131  & n1159 ;
  assign n1172 = n1154 & n1171 ;
  assign n1173 = ~\data_o[28]_pad  & ~n1159 ;
  assign n1175 = n1172 & ~n1173 ;
  assign n1176 = ~n1174 & n1175 ;
  assign n1180 = ~\mix1_data_o_reg_reg[20]/NET0131  & n1159 ;
  assign n1178 = n1154 & n1177 ;
  assign n1179 = ~\data_o[20]_pad  & ~n1159 ;
  assign n1181 = n1178 & ~n1179 ;
  assign n1182 = ~n1180 & n1181 ;
  assign n1243 = ~n1176 & ~n1182 ;
  assign n1252 = n1242 & n1243 ;
  assign n1253 = n1251 & n1252 ;
  assign n1239 = ~\mix1_data_o_reg_reg[108]/NET0131  & n1159 ;
  assign n1237 = n1153 & n1164 ;
  assign n1238 = ~\data_o[108]_pad  & ~n1159 ;
  assign n1240 = n1237 & ~n1238 ;
  assign n1241 = ~n1239 & n1240 ;
  assign n1229 = ~\mix1_data_o_reg_reg[92]/NET0131  & n1159 ;
  assign n1221 = \sub1_state_reg[2]/NET0131  & ~\sub1_state_reg[3]/NET0131  ;
  assign n1227 = n1171 & n1221 ;
  assign n1228 = ~\data_o[92]_pad  & ~n1159 ;
  assign n1230 = n1227 & ~n1228 ;
  assign n1231 = ~n1229 & n1230 ;
  assign n1234 = ~\mix1_data_o_reg_reg[76]/NET0131  & n1159 ;
  assign n1232 = n1153 & n1221 ;
  assign n1233 = ~\data_o[76]_pad  & ~n1159 ;
  assign n1235 = n1232 & ~n1233 ;
  assign n1236 = ~n1234 & n1235 ;
  assign n1248 = ~n1231 & ~n1236 ;
  assign n1249 = ~n1241 & n1248 ;
  assign n1208 = ~\mix1_data_o_reg_reg[68]/NET0131  & n1159 ;
  assign n1206 = ~\sub1_state_reg[3]/NET0131  & n1200 ;
  assign n1207 = ~\data_o[68]_pad  & ~n1159 ;
  assign n1209 = n1206 & ~n1207 ;
  assign n1210 = ~n1208 & n1209 ;
  assign n1213 = ~\mix1_data_o_reg_reg[36]/NET0131  & n1159 ;
  assign n1211 = n1165 & n1194 ;
  assign n1212 = ~\data_o[36]_pad  & ~n1159 ;
  assign n1214 = n1211 & ~n1212 ;
  assign n1215 = ~n1213 & n1214 ;
  assign n1246 = ~n1210 & ~n1215 ;
  assign n1218 = ~\mix1_data_o_reg_reg[52]/NET0131  & n1159 ;
  assign n1216 = n1177 & n1194 ;
  assign n1217 = ~\data_o[52]_pad  & ~n1159 ;
  assign n1219 = n1216 & ~n1217 ;
  assign n1220 = ~n1218 & n1219 ;
  assign n1224 = ~\mix1_data_o_reg_reg[84]/NET0131  & n1159 ;
  assign n1222 = n1177 & n1221 ;
  assign n1223 = ~\data_o[84]_pad  & ~n1159 ;
  assign n1225 = n1222 & ~n1223 ;
  assign n1226 = ~n1224 & n1225 ;
  assign n1247 = ~n1220 & ~n1226 ;
  assign n1250 = n1246 & n1247 ;
  assign n1254 = n1249 & n1250 ;
  assign n1255 = n1253 & n1254 ;
  assign n1256 = ~\sub1_state_reg[3]/NET0131  & n1183 ;
  assign n1257 = ~n1255 & ~n1256 ;
  assign n1259 = ~decrypt_i_pad & n1158 ;
  assign n1260 = decrypt_i_pad & n932 ;
  assign n1261 = ~n1259 & ~n1260 ;
  assign n1262 = \state_reg/NET0131  & ~n1261 ;
  assign n1263 = \addroundkey_ready_o_reg/NET0131  & ~n1159 ;
  assign n1264 = decrypt_i_pad & \mix1_ready_o_reg/NET0131  ;
  assign n1265 = ~n1263 & ~n1264 ;
  assign n1266 = ~n1262 & ~n1265 ;
  assign n1268 = ~\data_o[124]_pad  & ~n1159 ;
  assign n1258 = ~\mix1_data_o_reg_reg[124]/NET0131  & n1159 ;
  assign n1267 = ~\sub1_state_reg[4]/NET0131  & n1256 ;
  assign n1269 = ~n1258 & n1267 ;
  assign n1270 = ~n1268 & n1269 ;
  assign n1271 = n1266 & n1270 ;
  assign n1272 = ~n1257 & ~n1271 ;
  assign n1273 = n973 & ~n1272 ;
  assign n1141 = \ks1_state_reg[0]/NET0131  & \ks1_state_reg[1]/NET0131  ;
  assign n1142 = ~\ks1_state_reg[2]/NET0131  & n1141 ;
  assign n1143 = \key_i[4]_pad  & ~n953 ;
  assign n1144 = \ks1_key_reg_reg[4]/NET0131  & n956 ;
  assign n1145 = ~n1143 & ~n1144 ;
  assign n1146 = ~n933 & ~n1145 ;
  assign n1148 = ~\key_i[4]_pad  & n951 ;
  assign n1147 = ~\ks1_key_reg_reg[4]/NET0131  & ~n951 ;
  assign n1149 = n933 & ~n1147 ;
  assign n1150 = ~n1148 & n1149 ;
  assign n1151 = ~n1146 & ~n1150 ;
  assign n1152 = n1142 & ~n1151 ;
  assign n1274 = \ks1_state_reg[1]/NET0131  & n966 ;
  assign n1275 = \key_i[12]_pad  & ~n953 ;
  assign n1276 = \ks1_key_reg_reg[12]/NET0131  & n956 ;
  assign n1277 = ~n1275 & ~n1276 ;
  assign n1278 = ~n933 & ~n1277 ;
  assign n1280 = ~\key_i[12]_pad  & n951 ;
  assign n1279 = ~\ks1_key_reg_reg[12]/NET0131  & ~n951 ;
  assign n1281 = n933 & ~n1279 ;
  assign n1282 = ~n1280 & n1281 ;
  assign n1283 = ~n1278 & ~n1282 ;
  assign n1284 = n1274 & ~n1283 ;
  assign n1307 = ~n1152 & ~n1284 ;
  assign n1285 = \ks1_state_reg[0]/NET0131  & ~\ks1_state_reg[1]/NET0131  ;
  assign n1286 = ~\ks1_state_reg[2]/NET0131  & n1285 ;
  assign n1287 = \key_i[20]_pad  & ~n953 ;
  assign n1288 = \ks1_key_reg_reg[20]/NET0131  & n956 ;
  assign n1289 = ~n1287 & ~n1288 ;
  assign n1290 = ~n933 & ~n1289 ;
  assign n1292 = ~\key_i[20]_pad  & n951 ;
  assign n1291 = ~\ks1_key_reg_reg[20]/NET0131  & ~n951 ;
  assign n1293 = n933 & ~n1291 ;
  assign n1294 = ~n1292 & n1293 ;
  assign n1295 = ~n1290 & ~n1294 ;
  assign n1296 = n1286 & ~n1295 ;
  assign n1297 = \key_i[28]_pad  & ~n953 ;
  assign n1298 = \ks1_key_reg_reg[28]/NET0131  & n956 ;
  assign n1299 = ~n1297 & ~n1298 ;
  assign n1300 = ~n933 & ~n1299 ;
  assign n1302 = ~\key_i[28]_pad  & n951 ;
  assign n1301 = ~\ks1_key_reg_reg[28]/NET0131  & ~n951 ;
  assign n1303 = n933 & ~n1301 ;
  assign n1304 = ~n1302 & n1303 ;
  assign n1305 = ~n1300 & ~n1304 ;
  assign n1306 = n971 & ~n1305 ;
  assign n1308 = ~n1296 & ~n1306 ;
  assign n1309 = n1307 & n1308 ;
  assign n1310 = ~n1273 & n1309 ;
  assign n1311 = ~n974 & ~n1310 ;
  assign n1329 = ~\mix1_data_o_reg_reg[70]/NET0131  & n1159 ;
  assign n1328 = ~\data_o[70]_pad  & ~n1159 ;
  assign n1330 = n1206 & ~n1328 ;
  assign n1331 = ~n1329 & n1330 ;
  assign n1333 = ~\mix1_data_o_reg_reg[30]/NET0131  & n1159 ;
  assign n1332 = ~\data_o[30]_pad  & ~n1159 ;
  assign n1334 = n1172 & ~n1332 ;
  assign n1335 = ~n1333 & n1334 ;
  assign n1374 = ~n1331 & ~n1335 ;
  assign n1337 = ~\mix1_data_o_reg_reg[54]/NET0131  & n1159 ;
  assign n1336 = ~\data_o[54]_pad  & ~n1159 ;
  assign n1338 = n1216 & ~n1336 ;
  assign n1339 = ~n1337 & n1338 ;
  assign n1341 = ~\mix1_data_o_reg_reg[22]/NET0131  & n1159 ;
  assign n1340 = ~\data_o[22]_pad  & ~n1159 ;
  assign n1342 = n1178 & ~n1340 ;
  assign n1343 = ~n1341 & n1342 ;
  assign n1375 = ~n1339 & ~n1343 ;
  assign n1381 = n1374 & n1375 ;
  assign n1313 = ~\mix1_data_o_reg_reg[118]/NET0131  & n1159 ;
  assign n1312 = ~\data_o[118]_pad  & ~n1159 ;
  assign n1314 = n1189 & ~n1312 ;
  assign n1315 = ~n1313 & n1314 ;
  assign n1317 = ~\mix1_data_o_reg_reg[110]/NET0131  & n1159 ;
  assign n1316 = ~\data_o[110]_pad  & ~n1159 ;
  assign n1318 = n1237 & ~n1316 ;
  assign n1319 = ~n1317 & n1318 ;
  assign n1372 = ~n1315 & ~n1319 ;
  assign n1321 = ~\mix1_data_o_reg_reg[102]/NET0131  & n1159 ;
  assign n1320 = ~\data_o[102]_pad  & ~n1159 ;
  assign n1322 = n1166 & ~n1320 ;
  assign n1323 = ~n1321 & n1322 ;
  assign n1325 = ~\mix1_data_o_reg_reg[46]/NET0131  & n1159 ;
  assign n1324 = ~\data_o[46]_pad  & ~n1159 ;
  assign n1326 = n1195 & ~n1324 ;
  assign n1327 = ~n1325 & n1326 ;
  assign n1373 = ~n1323 & ~n1327 ;
  assign n1382 = n1372 & n1373 ;
  assign n1383 = n1381 & n1382 ;
  assign n1369 = ~\mix1_data_o_reg_reg[14]/NET0131  & n1159 ;
  assign n1368 = ~\data_o[14]_pad  & ~n1159 ;
  assign n1370 = n1155 & ~n1368 ;
  assign n1371 = ~n1369 & n1370 ;
  assign n1361 = ~\mix1_data_o_reg_reg[62]/NET0131  & n1159 ;
  assign n1360 = ~\data_o[62]_pad  & ~n1159 ;
  assign n1362 = n1184 & ~n1360 ;
  assign n1363 = ~n1361 & n1362 ;
  assign n1365 = ~\mix1_data_o_reg_reg[86]/NET0131  & n1159 ;
  assign n1364 = ~\data_o[86]_pad  & ~n1159 ;
  assign n1366 = n1222 & ~n1364 ;
  assign n1367 = ~n1365 & n1366 ;
  assign n1378 = ~n1363 & ~n1367 ;
  assign n1379 = ~n1371 & n1378 ;
  assign n1345 = ~\mix1_data_o_reg_reg[6]/NET0131  & n1159 ;
  assign n1344 = ~\data_o[6]_pad  & ~n1159 ;
  assign n1346 = n1201 & ~n1344 ;
  assign n1347 = ~n1345 & n1346 ;
  assign n1349 = ~\mix1_data_o_reg_reg[94]/NET0131  & n1159 ;
  assign n1348 = ~\data_o[94]_pad  & ~n1159 ;
  assign n1350 = n1227 & ~n1348 ;
  assign n1351 = ~n1349 & n1350 ;
  assign n1376 = ~n1347 & ~n1351 ;
  assign n1353 = ~\mix1_data_o_reg_reg[78]/NET0131  & n1159 ;
  assign n1352 = ~\data_o[78]_pad  & ~n1159 ;
  assign n1354 = n1232 & ~n1352 ;
  assign n1355 = ~n1353 & n1354 ;
  assign n1357 = ~\mix1_data_o_reg_reg[38]/NET0131  & n1159 ;
  assign n1356 = ~\data_o[38]_pad  & ~n1159 ;
  assign n1358 = n1211 & ~n1356 ;
  assign n1359 = ~n1357 & n1358 ;
  assign n1377 = ~n1355 & ~n1359 ;
  assign n1380 = n1376 & n1377 ;
  assign n1384 = n1379 & n1380 ;
  assign n1385 = n1383 & n1384 ;
  assign n1386 = ~n1256 & ~n1385 ;
  assign n1388 = ~\data_o[126]_pad  & ~n1159 ;
  assign n1387 = ~\mix1_data_o_reg_reg[126]/NET0131  & n1159 ;
  assign n1389 = n1267 & ~n1387 ;
  assign n1390 = ~n1388 & n1389 ;
  assign n1391 = n1266 & n1390 ;
  assign n1392 = ~n1386 & ~n1391 ;
  assign n1393 = n973 & ~n1392 ;
  assign n1412 = ~n964 & n1274 ;
  assign n1394 = \key_i[30]_pad  & ~n953 ;
  assign n1395 = \ks1_key_reg_reg[30]/NET0131  & n956 ;
  assign n1396 = ~n1394 & ~n1395 ;
  assign n1397 = ~n933 & ~n1396 ;
  assign n1399 = ~\key_i[30]_pad  & n951 ;
  assign n1398 = ~\ks1_key_reg_reg[30]/NET0131  & ~n951 ;
  assign n1400 = n933 & ~n1398 ;
  assign n1401 = ~n1399 & n1400 ;
  assign n1402 = ~n1397 & ~n1401 ;
  assign n1403 = n971 & ~n1402 ;
  assign n1404 = \key_i[6]_pad  & ~n1116 ;
  assign n1405 = \ks1_key_reg_reg[6]/NET0131  & n1116 ;
  assign n1406 = ~n1404 & ~n1405 ;
  assign n1407 = n1142 & ~n1406 ;
  assign n1408 = \key_i[22]_pad  & ~n1116 ;
  assign n1409 = \ks1_key_reg_reg[22]/NET0131  & n1116 ;
  assign n1410 = ~n1408 & ~n1409 ;
  assign n1411 = n1286 & ~n1410 ;
  assign n1413 = ~n1407 & ~n1411 ;
  assign n1414 = ~n1403 & n1413 ;
  assign n1415 = ~n1412 & n1414 ;
  assign n1416 = ~n1393 & n1415 ;
  assign n1434 = ~\mix1_data_o_reg_reg[67]/NET0131  & n1159 ;
  assign n1433 = ~\data_o[67]_pad  & ~n1159 ;
  assign n1435 = n1206 & ~n1433 ;
  assign n1436 = ~n1434 & n1435 ;
  assign n1438 = ~\mix1_data_o_reg_reg[115]/NET0131  & n1159 ;
  assign n1437 = ~\data_o[115]_pad  & ~n1159 ;
  assign n1439 = n1189 & ~n1437 ;
  assign n1440 = ~n1438 & n1439 ;
  assign n1479 = ~n1436 & ~n1440 ;
  assign n1442 = ~\mix1_data_o_reg_reg[43]/NET0131  & n1159 ;
  assign n1441 = ~\data_o[43]_pad  & ~n1159 ;
  assign n1443 = n1195 & ~n1441 ;
  assign n1444 = ~n1442 & n1443 ;
  assign n1446 = ~\mix1_data_o_reg_reg[51]/NET0131  & n1159 ;
  assign n1445 = ~\data_o[51]_pad  & ~n1159 ;
  assign n1447 = n1216 & ~n1445 ;
  assign n1448 = ~n1446 & n1447 ;
  assign n1480 = ~n1444 & ~n1448 ;
  assign n1486 = n1479 & n1480 ;
  assign n1418 = ~\mix1_data_o_reg_reg[99]/NET0131  & n1159 ;
  assign n1417 = ~\data_o[99]_pad  & ~n1159 ;
  assign n1419 = n1166 & ~n1417 ;
  assign n1420 = ~n1418 & n1419 ;
  assign n1422 = ~\mix1_data_o_reg_reg[83]/NET0131  & n1159 ;
  assign n1421 = ~\data_o[83]_pad  & ~n1159 ;
  assign n1423 = n1222 & ~n1421 ;
  assign n1424 = ~n1422 & n1423 ;
  assign n1477 = ~n1420 & ~n1424 ;
  assign n1426 = ~\mix1_data_o_reg_reg[35]/NET0131  & n1159 ;
  assign n1425 = ~\data_o[35]_pad  & ~n1159 ;
  assign n1427 = n1211 & ~n1425 ;
  assign n1428 = ~n1426 & n1427 ;
  assign n1430 = ~\mix1_data_o_reg_reg[91]/NET0131  & n1159 ;
  assign n1429 = ~\data_o[91]_pad  & ~n1159 ;
  assign n1431 = n1227 & ~n1429 ;
  assign n1432 = ~n1430 & n1431 ;
  assign n1478 = ~n1428 & ~n1432 ;
  assign n1487 = n1477 & n1478 ;
  assign n1488 = n1486 & n1487 ;
  assign n1474 = ~\mix1_data_o_reg_reg[27]/NET0131  & n1159 ;
  assign n1473 = ~\data_o[27]_pad  & ~n1159 ;
  assign n1475 = n1172 & ~n1473 ;
  assign n1476 = ~n1474 & n1475 ;
  assign n1466 = ~\mix1_data_o_reg_reg[59]/NET0131  & n1159 ;
  assign n1465 = ~\data_o[59]_pad  & ~n1159 ;
  assign n1467 = n1184 & ~n1465 ;
  assign n1468 = ~n1466 & n1467 ;
  assign n1470 = ~\mix1_data_o_reg_reg[107]/NET0131  & n1159 ;
  assign n1469 = ~\data_o[107]_pad  & ~n1159 ;
  assign n1471 = n1237 & ~n1469 ;
  assign n1472 = ~n1470 & n1471 ;
  assign n1483 = ~n1468 & ~n1472 ;
  assign n1484 = ~n1476 & n1483 ;
  assign n1450 = ~\mix1_data_o_reg_reg[3]/NET0131  & n1159 ;
  assign n1449 = ~\data_o[3]_pad  & ~n1159 ;
  assign n1451 = n1201 & ~n1449 ;
  assign n1452 = ~n1450 & n1451 ;
  assign n1454 = ~\mix1_data_o_reg_reg[75]/NET0131  & n1159 ;
  assign n1453 = ~\data_o[75]_pad  & ~n1159 ;
  assign n1455 = n1232 & ~n1453 ;
  assign n1456 = ~n1454 & n1455 ;
  assign n1481 = ~n1452 & ~n1456 ;
  assign n1458 = ~\mix1_data_o_reg_reg[19]/NET0131  & n1159 ;
  assign n1457 = ~\data_o[19]_pad  & ~n1159 ;
  assign n1459 = n1178 & ~n1457 ;
  assign n1460 = ~n1458 & n1459 ;
  assign n1462 = ~\mix1_data_o_reg_reg[11]/NET0131  & n1159 ;
  assign n1461 = ~\data_o[11]_pad  & ~n1159 ;
  assign n1463 = n1155 & ~n1461 ;
  assign n1464 = ~n1462 & n1463 ;
  assign n1482 = ~n1460 & ~n1464 ;
  assign n1485 = n1481 & n1482 ;
  assign n1489 = n1484 & n1485 ;
  assign n1490 = n1488 & n1489 ;
  assign n1491 = ~n1256 & ~n1490 ;
  assign n1493 = ~\data_o[123]_pad  & ~n1159 ;
  assign n1492 = ~\mix1_data_o_reg_reg[123]/NET0131  & n1159 ;
  assign n1494 = n1267 & ~n1492 ;
  assign n1495 = ~n1493 & n1494 ;
  assign n1496 = n1266 & n1495 ;
  assign n1497 = ~n1491 & ~n1496 ;
  assign n1498 = n973 & ~n1497 ;
  assign n1499 = \key_i[3]_pad  & ~n953 ;
  assign n1500 = \ks1_key_reg_reg[3]/NET0131  & n956 ;
  assign n1501 = ~n1499 & ~n1500 ;
  assign n1502 = ~n933 & ~n1501 ;
  assign n1504 = ~\key_i[3]_pad  & n951 ;
  assign n1503 = ~\ks1_key_reg_reg[3]/NET0131  & ~n951 ;
  assign n1505 = n933 & ~n1503 ;
  assign n1506 = ~n1504 & n1505 ;
  assign n1507 = ~n1502 & ~n1506 ;
  assign n1508 = n1142 & ~n1507 ;
  assign n1509 = \key_i[19]_pad  & ~n953 ;
  assign n1510 = \ks1_key_reg_reg[19]/NET0131  & n956 ;
  assign n1511 = ~n1509 & ~n1510 ;
  assign n1512 = ~n933 & ~n1511 ;
  assign n1514 = ~\key_i[19]_pad  & n951 ;
  assign n1513 = ~\ks1_key_reg_reg[19]/NET0131  & ~n951 ;
  assign n1515 = n933 & ~n1513 ;
  assign n1516 = ~n1514 & n1515 ;
  assign n1517 = ~n1512 & ~n1516 ;
  assign n1518 = n1286 & ~n1517 ;
  assign n1539 = ~n1508 & ~n1518 ;
  assign n1519 = \key_i[11]_pad  & ~n953 ;
  assign n1520 = \ks1_key_reg_reg[11]/NET0131  & n956 ;
  assign n1521 = ~n1519 & ~n1520 ;
  assign n1522 = ~n933 & ~n1521 ;
  assign n1524 = ~\key_i[11]_pad  & n951 ;
  assign n1523 = ~\ks1_key_reg_reg[11]/NET0131  & ~n951 ;
  assign n1525 = n933 & ~n1523 ;
  assign n1526 = ~n1524 & n1525 ;
  assign n1527 = ~n1522 & ~n1526 ;
  assign n1528 = n1274 & ~n1527 ;
  assign n1529 = \key_i[27]_pad  & ~n953 ;
  assign n1530 = \ks1_key_reg_reg[27]/NET0131  & n956 ;
  assign n1531 = ~n1529 & ~n1530 ;
  assign n1532 = ~n933 & ~n1531 ;
  assign n1534 = ~\key_i[27]_pad  & n951 ;
  assign n1533 = ~\ks1_key_reg_reg[27]/NET0131  & ~n951 ;
  assign n1535 = n933 & ~n1533 ;
  assign n1536 = ~n1534 & n1535 ;
  assign n1537 = ~n1532 & ~n1536 ;
  assign n1538 = n971 & ~n1537 ;
  assign n1540 = ~n1528 & ~n1538 ;
  assign n1541 = n1539 & n1540 ;
  assign n1542 = ~n1498 & n1541 ;
  assign n1543 = n1416 & ~n1542 ;
  assign n1544 = ~n1416 & n1542 ;
  assign n1545 = ~n1543 & ~n1544 ;
  assign n1573 = ~\mix1_data_o_reg_reg[9]/NET0131  & n1159 ;
  assign n1572 = ~\data_o[9]_pad  & ~n1159 ;
  assign n1574 = n1155 & ~n1572 ;
  assign n1575 = ~n1573 & n1574 ;
  assign n1577 = ~\mix1_data_o_reg_reg[57]/NET0131  & n1159 ;
  assign n1576 = ~\data_o[57]_pad  & ~n1159 ;
  assign n1578 = n1184 & ~n1576 ;
  assign n1579 = ~n1577 & n1578 ;
  assign n1618 = ~n1575 & ~n1579 ;
  assign n1581 = ~\mix1_data_o_reg_reg[49]/NET0131  & n1159 ;
  assign n1580 = ~\data_o[49]_pad  & ~n1159 ;
  assign n1582 = n1216 & ~n1580 ;
  assign n1583 = ~n1581 & n1582 ;
  assign n1585 = ~\mix1_data_o_reg_reg[89]/NET0131  & n1159 ;
  assign n1584 = ~\data_o[89]_pad  & ~n1159 ;
  assign n1586 = n1227 & ~n1584 ;
  assign n1587 = ~n1585 & n1586 ;
  assign n1619 = ~n1583 & ~n1587 ;
  assign n1625 = n1618 & n1619 ;
  assign n1557 = ~\mix1_data_o_reg_reg[105]/NET0131  & n1159 ;
  assign n1556 = ~\data_o[105]_pad  & ~n1159 ;
  assign n1558 = n1237 & ~n1556 ;
  assign n1559 = ~n1557 & n1558 ;
  assign n1561 = ~\mix1_data_o_reg_reg[81]/NET0131  & n1159 ;
  assign n1560 = ~\data_o[81]_pad  & ~n1159 ;
  assign n1562 = n1222 & ~n1560 ;
  assign n1563 = ~n1561 & n1562 ;
  assign n1616 = ~n1559 & ~n1563 ;
  assign n1565 = ~\mix1_data_o_reg_reg[113]/NET0131  & n1159 ;
  assign n1564 = ~\data_o[113]_pad  & ~n1159 ;
  assign n1566 = n1189 & ~n1564 ;
  assign n1567 = ~n1565 & n1566 ;
  assign n1569 = ~\mix1_data_o_reg_reg[17]/NET0131  & n1159 ;
  assign n1568 = ~\data_o[17]_pad  & ~n1159 ;
  assign n1570 = n1178 & ~n1568 ;
  assign n1571 = ~n1569 & n1570 ;
  assign n1617 = ~n1567 & ~n1571 ;
  assign n1626 = n1616 & n1617 ;
  assign n1627 = n1625 & n1626 ;
  assign n1613 = ~\mix1_data_o_reg_reg[97]/NET0131  & n1159 ;
  assign n1612 = ~\data_o[97]_pad  & ~n1159 ;
  assign n1614 = n1166 & ~n1612 ;
  assign n1615 = ~n1613 & n1614 ;
  assign n1605 = ~\mix1_data_o_reg_reg[73]/NET0131  & n1159 ;
  assign n1604 = ~\data_o[73]_pad  & ~n1159 ;
  assign n1606 = n1232 & ~n1604 ;
  assign n1607 = ~n1605 & n1606 ;
  assign n1609 = ~\mix1_data_o_reg_reg[1]/NET0131  & n1159 ;
  assign n1608 = ~\data_o[1]_pad  & ~n1159 ;
  assign n1610 = n1201 & ~n1608 ;
  assign n1611 = ~n1609 & n1610 ;
  assign n1622 = ~n1607 & ~n1611 ;
  assign n1623 = ~n1615 & n1622 ;
  assign n1589 = ~\mix1_data_o_reg_reg[41]/NET0131  & n1159 ;
  assign n1588 = ~\data_o[41]_pad  & ~n1159 ;
  assign n1590 = n1195 & ~n1588 ;
  assign n1591 = ~n1589 & n1590 ;
  assign n1593 = ~\mix1_data_o_reg_reg[25]/NET0131  & n1159 ;
  assign n1592 = ~\data_o[25]_pad  & ~n1159 ;
  assign n1594 = n1172 & ~n1592 ;
  assign n1595 = ~n1593 & n1594 ;
  assign n1620 = ~n1591 & ~n1595 ;
  assign n1597 = ~\mix1_data_o_reg_reg[65]/NET0131  & n1159 ;
  assign n1596 = ~\data_o[65]_pad  & ~n1159 ;
  assign n1598 = n1206 & ~n1596 ;
  assign n1599 = ~n1597 & n1598 ;
  assign n1601 = ~\mix1_data_o_reg_reg[33]/NET0131  & n1159 ;
  assign n1600 = ~\data_o[33]_pad  & ~n1159 ;
  assign n1602 = n1211 & ~n1600 ;
  assign n1603 = ~n1601 & n1602 ;
  assign n1621 = ~n1599 & ~n1603 ;
  assign n1624 = n1620 & n1621 ;
  assign n1628 = n1623 & n1624 ;
  assign n1629 = n1627 & n1628 ;
  assign n1630 = ~n1256 & ~n1629 ;
  assign n1632 = ~\data_o[121]_pad  & ~n1159 ;
  assign n1631 = ~\mix1_data_o_reg_reg[121]/NET0131  & n1159 ;
  assign n1633 = n1267 & ~n1631 ;
  assign n1634 = ~n1632 & n1633 ;
  assign n1635 = n1266 & n1634 ;
  assign n1636 = ~n1630 & ~n1635 ;
  assign n1637 = n973 & ~n1636 ;
  assign n1546 = \key_i[9]_pad  & ~n953 ;
  assign n1547 = \ks1_key_reg_reg[9]/NET0131  & n956 ;
  assign n1548 = ~n1546 & ~n1547 ;
  assign n1549 = ~n933 & ~n1548 ;
  assign n1551 = ~\key_i[9]_pad  & n951 ;
  assign n1550 = ~\ks1_key_reg_reg[9]/NET0131  & ~n951 ;
  assign n1552 = n933 & ~n1550 ;
  assign n1553 = ~n1551 & n1552 ;
  assign n1554 = ~n1549 & ~n1553 ;
  assign n1555 = n1274 & ~n1554 ;
  assign n1638 = \key_i[17]_pad  & ~n953 ;
  assign n1639 = \ks1_key_reg_reg[17]/NET0131  & n956 ;
  assign n1640 = ~n1638 & ~n1639 ;
  assign n1641 = ~n933 & ~n1640 ;
  assign n1643 = ~\key_i[17]_pad  & n951 ;
  assign n1642 = ~\ks1_key_reg_reg[17]/NET0131  & ~n951 ;
  assign n1644 = n933 & ~n1642 ;
  assign n1645 = ~n1643 & n1644 ;
  assign n1646 = ~n1641 & ~n1645 ;
  assign n1647 = n1286 & ~n1646 ;
  assign n1668 = ~n1555 & ~n1647 ;
  assign n1648 = \key_i[25]_pad  & ~n953 ;
  assign n1649 = \ks1_key_reg_reg[25]/NET0131  & n956 ;
  assign n1650 = ~n1648 & ~n1649 ;
  assign n1651 = ~n933 & ~n1650 ;
  assign n1653 = ~\key_i[25]_pad  & n951 ;
  assign n1652 = ~\ks1_key_reg_reg[25]/NET0131  & ~n951 ;
  assign n1654 = n933 & ~n1652 ;
  assign n1655 = ~n1653 & n1654 ;
  assign n1656 = ~n1651 & ~n1655 ;
  assign n1657 = n971 & ~n1656 ;
  assign n1658 = \key_i[1]_pad  & ~n953 ;
  assign n1659 = \ks1_key_reg_reg[1]/NET0131  & n956 ;
  assign n1660 = ~n1658 & ~n1659 ;
  assign n1661 = ~n933 & ~n1660 ;
  assign n1663 = ~\key_i[1]_pad  & n951 ;
  assign n1662 = ~\ks1_key_reg_reg[1]/NET0131  & ~n951 ;
  assign n1664 = n933 & ~n1662 ;
  assign n1665 = ~n1663 & n1664 ;
  assign n1666 = ~n1661 & ~n1665 ;
  assign n1667 = n1142 & ~n1666 ;
  assign n1669 = ~n1657 & ~n1667 ;
  assign n1670 = n1668 & n1669 ;
  assign n1671 = ~n1637 & n1670 ;
  assign n1673 = ~n1545 & ~n1671 ;
  assign n1672 = n1545 & n1671 ;
  assign n1674 = n974 & ~n1672 ;
  assign n1675 = ~n1673 & n1674 ;
  assign n1676 = ~n1311 & ~n1675 ;
  assign n1694 = ~\mix1_data_o_reg_reg[72]/NET0131  & n1159 ;
  assign n1693 = ~\data_o[72]_pad  & ~n1159 ;
  assign n1695 = n1232 & ~n1693 ;
  assign n1696 = ~n1694 & n1695 ;
  assign n1698 = ~\mix1_data_o_reg_reg[56]/NET0131  & n1159 ;
  assign n1697 = ~\data_o[56]_pad  & ~n1159 ;
  assign n1699 = n1184 & ~n1697 ;
  assign n1700 = ~n1698 & n1699 ;
  assign n1739 = ~n1696 & ~n1700 ;
  assign n1702 = ~\mix1_data_o_reg_reg[88]/NET0131  & n1159 ;
  assign n1701 = ~\data_o[88]_pad  & ~n1159 ;
  assign n1703 = n1227 & ~n1701 ;
  assign n1704 = ~n1702 & n1703 ;
  assign n1706 = ~\mix1_data_o_reg_reg[40]/NET0131  & n1159 ;
  assign n1705 = ~\data_o[40]_pad  & ~n1159 ;
  assign n1707 = n1195 & ~n1705 ;
  assign n1708 = ~n1706 & n1707 ;
  assign n1740 = ~n1704 & ~n1708 ;
  assign n1746 = n1739 & n1740 ;
  assign n1678 = ~\mix1_data_o_reg_reg[112]/NET0131  & n1159 ;
  assign n1677 = ~\data_o[112]_pad  & ~n1159 ;
  assign n1679 = n1189 & ~n1677 ;
  assign n1680 = ~n1678 & n1679 ;
  assign n1682 = ~\mix1_data_o_reg_reg[96]/NET0131  & n1159 ;
  assign n1681 = ~\data_o[96]_pad  & ~n1159 ;
  assign n1683 = n1166 & ~n1681 ;
  assign n1684 = ~n1682 & n1683 ;
  assign n1737 = ~n1680 & ~n1684 ;
  assign n1686 = ~\mix1_data_o_reg_reg[104]/NET0131  & n1159 ;
  assign n1685 = ~\data_o[104]_pad  & ~n1159 ;
  assign n1687 = n1237 & ~n1685 ;
  assign n1688 = ~n1686 & n1687 ;
  assign n1690 = ~\mix1_data_o_reg_reg[64]/NET0131  & n1159 ;
  assign n1689 = ~\data_o[64]_pad  & ~n1159 ;
  assign n1691 = n1206 & ~n1689 ;
  assign n1692 = ~n1690 & n1691 ;
  assign n1738 = ~n1688 & ~n1692 ;
  assign n1747 = n1737 & n1738 ;
  assign n1748 = n1746 & n1747 ;
  assign n1734 = ~\mix1_data_o_reg_reg[80]/NET0131  & n1159 ;
  assign n1733 = ~\data_o[80]_pad  & ~n1159 ;
  assign n1735 = n1222 & ~n1733 ;
  assign n1736 = ~n1734 & n1735 ;
  assign n1726 = ~\mix1_data_o_reg_reg[8]/NET0131  & n1159 ;
  assign n1725 = ~\data_o[8]_pad  & ~n1159 ;
  assign n1727 = n1155 & ~n1725 ;
  assign n1728 = ~n1726 & n1727 ;
  assign n1730 = ~\mix1_data_o_reg_reg[32]/NET0131  & n1159 ;
  assign n1729 = ~\data_o[32]_pad  & ~n1159 ;
  assign n1731 = n1211 & ~n1729 ;
  assign n1732 = ~n1730 & n1731 ;
  assign n1743 = ~n1728 & ~n1732 ;
  assign n1744 = ~n1736 & n1743 ;
  assign n1710 = ~\mix1_data_o_reg_reg[48]/NET0131  & n1159 ;
  assign n1709 = ~\data_o[48]_pad  & ~n1159 ;
  assign n1711 = n1216 & ~n1709 ;
  assign n1712 = ~n1710 & n1711 ;
  assign n1714 = ~\mix1_data_o_reg_reg[0]/NET0131  & n1159 ;
  assign n1713 = ~\data_o[0]_pad  & ~n1159 ;
  assign n1715 = n1201 & ~n1713 ;
  assign n1716 = ~n1714 & n1715 ;
  assign n1741 = ~n1712 & ~n1716 ;
  assign n1718 = ~\mix1_data_o_reg_reg[16]/NET0131  & n1159 ;
  assign n1717 = ~\data_o[16]_pad  & ~n1159 ;
  assign n1719 = n1178 & ~n1717 ;
  assign n1720 = ~n1718 & n1719 ;
  assign n1722 = ~\mix1_data_o_reg_reg[24]/NET0131  & n1159 ;
  assign n1721 = ~\data_o[24]_pad  & ~n1159 ;
  assign n1723 = n1172 & ~n1721 ;
  assign n1724 = ~n1722 & n1723 ;
  assign n1742 = ~n1720 & ~n1724 ;
  assign n1745 = n1741 & n1742 ;
  assign n1749 = n1744 & n1745 ;
  assign n1750 = n1748 & n1749 ;
  assign n1751 = ~n1256 & ~n1750 ;
  assign n1753 = ~\data_o[120]_pad  & ~n1159 ;
  assign n1752 = ~\mix1_data_o_reg_reg[120]/NET0131  & n1159 ;
  assign n1754 = n1267 & ~n1752 ;
  assign n1755 = ~n1753 & n1754 ;
  assign n1756 = n1266 & n1755 ;
  assign n1757 = ~n1751 & ~n1756 ;
  assign n1758 = n973 & ~n1757 ;
  assign n1759 = \key_i[16]_pad  & ~n1116 ;
  assign n1760 = \ks1_key_reg_reg[16]/NET0131  & n1116 ;
  assign n1761 = ~n1759 & ~n1760 ;
  assign n1762 = n1286 & ~n1761 ;
  assign n1763 = \key_i[8]_pad  & ~n953 ;
  assign n1764 = \ks1_key_reg_reg[8]/NET0131  & n956 ;
  assign n1765 = ~n1763 & ~n1764 ;
  assign n1766 = ~n933 & ~n1765 ;
  assign n1768 = ~\key_i[8]_pad  & n951 ;
  assign n1767 = ~\ks1_key_reg_reg[8]/NET0131  & ~n951 ;
  assign n1769 = n933 & ~n1767 ;
  assign n1770 = ~n1768 & n1769 ;
  assign n1771 = ~n1766 & ~n1770 ;
  assign n1772 = n1274 & ~n1771 ;
  assign n1793 = ~n1762 & ~n1772 ;
  assign n1773 = \key_i[24]_pad  & ~n953 ;
  assign n1774 = \ks1_key_reg_reg[24]/NET0131  & n956 ;
  assign n1775 = ~n1773 & ~n1774 ;
  assign n1776 = ~n933 & ~n1775 ;
  assign n1778 = ~\key_i[24]_pad  & n951 ;
  assign n1777 = ~\ks1_key_reg_reg[24]/NET0131  & ~n951 ;
  assign n1779 = n933 & ~n1777 ;
  assign n1780 = ~n1778 & n1779 ;
  assign n1781 = ~n1776 & ~n1780 ;
  assign n1782 = n971 & ~n1781 ;
  assign n1783 = \key_i[0]_pad  & ~n953 ;
  assign n1784 = \ks1_key_reg_reg[0]/NET0131  & n956 ;
  assign n1785 = ~n1783 & ~n1784 ;
  assign n1786 = ~n933 & ~n1785 ;
  assign n1788 = ~\key_i[0]_pad  & n951 ;
  assign n1787 = ~\ks1_key_reg_reg[0]/NET0131  & ~n951 ;
  assign n1789 = n933 & ~n1787 ;
  assign n1790 = ~n1788 & n1789 ;
  assign n1791 = ~n1786 & ~n1790 ;
  assign n1792 = n1142 & ~n1791 ;
  assign n1794 = ~n1782 & ~n1792 ;
  assign n1795 = n1793 & n1794 ;
  assign n1796 = ~n1758 & n1795 ;
  assign n1814 = ~\mix1_data_o_reg_reg[21]/NET0131  & n1159 ;
  assign n1813 = ~\data_o[21]_pad  & ~n1159 ;
  assign n1815 = n1178 & ~n1813 ;
  assign n1816 = ~n1814 & n1815 ;
  assign n1818 = ~\mix1_data_o_reg_reg[13]/NET0131  & n1159 ;
  assign n1817 = ~\data_o[13]_pad  & ~n1159 ;
  assign n1819 = n1155 & ~n1817 ;
  assign n1820 = ~n1818 & n1819 ;
  assign n1859 = ~n1816 & ~n1820 ;
  assign n1822 = ~\mix1_data_o_reg_reg[5]/NET0131  & n1159 ;
  assign n1821 = ~\data_o[5]_pad  & ~n1159 ;
  assign n1823 = n1201 & ~n1821 ;
  assign n1824 = ~n1822 & n1823 ;
  assign n1826 = ~\mix1_data_o_reg_reg[53]/NET0131  & n1159 ;
  assign n1825 = ~\data_o[53]_pad  & ~n1159 ;
  assign n1827 = n1216 & ~n1825 ;
  assign n1828 = ~n1826 & n1827 ;
  assign n1860 = ~n1824 & ~n1828 ;
  assign n1866 = n1859 & n1860 ;
  assign n1798 = ~\mix1_data_o_reg_reg[61]/NET0131  & n1159 ;
  assign n1797 = ~\data_o[61]_pad  & ~n1159 ;
  assign n1799 = n1184 & ~n1797 ;
  assign n1800 = ~n1798 & n1799 ;
  assign n1802 = ~\mix1_data_o_reg_reg[29]/NET0131  & n1159 ;
  assign n1801 = ~\data_o[29]_pad  & ~n1159 ;
  assign n1803 = n1172 & ~n1801 ;
  assign n1804 = ~n1802 & n1803 ;
  assign n1857 = ~n1800 & ~n1804 ;
  assign n1806 = ~\mix1_data_o_reg_reg[85]/NET0131  & n1159 ;
  assign n1805 = ~\data_o[85]_pad  & ~n1159 ;
  assign n1807 = n1222 & ~n1805 ;
  assign n1808 = ~n1806 & n1807 ;
  assign n1810 = ~\mix1_data_o_reg_reg[69]/NET0131  & n1159 ;
  assign n1809 = ~\data_o[69]_pad  & ~n1159 ;
  assign n1811 = n1206 & ~n1809 ;
  assign n1812 = ~n1810 & n1811 ;
  assign n1858 = ~n1808 & ~n1812 ;
  assign n1867 = n1857 & n1858 ;
  assign n1868 = n1866 & n1867 ;
  assign n1854 = ~\mix1_data_o_reg_reg[109]/NET0131  & n1159 ;
  assign n1853 = ~\data_o[109]_pad  & ~n1159 ;
  assign n1855 = n1237 & ~n1853 ;
  assign n1856 = ~n1854 & n1855 ;
  assign n1846 = ~\mix1_data_o_reg_reg[117]/NET0131  & n1159 ;
  assign n1845 = ~\data_o[117]_pad  & ~n1159 ;
  assign n1847 = n1189 & ~n1845 ;
  assign n1848 = ~n1846 & n1847 ;
  assign n1850 = ~\mix1_data_o_reg_reg[37]/NET0131  & n1159 ;
  assign n1849 = ~\data_o[37]_pad  & ~n1159 ;
  assign n1851 = n1211 & ~n1849 ;
  assign n1852 = ~n1850 & n1851 ;
  assign n1863 = ~n1848 & ~n1852 ;
  assign n1864 = ~n1856 & n1863 ;
  assign n1830 = ~\mix1_data_o_reg_reg[45]/NET0131  & n1159 ;
  assign n1829 = ~\data_o[45]_pad  & ~n1159 ;
  assign n1831 = n1195 & ~n1829 ;
  assign n1832 = ~n1830 & n1831 ;
  assign n1834 = ~\mix1_data_o_reg_reg[93]/NET0131  & n1159 ;
  assign n1833 = ~\data_o[93]_pad  & ~n1159 ;
  assign n1835 = n1227 & ~n1833 ;
  assign n1836 = ~n1834 & n1835 ;
  assign n1861 = ~n1832 & ~n1836 ;
  assign n1838 = ~\mix1_data_o_reg_reg[77]/NET0131  & n1159 ;
  assign n1837 = ~\data_o[77]_pad  & ~n1159 ;
  assign n1839 = n1232 & ~n1837 ;
  assign n1840 = ~n1838 & n1839 ;
  assign n1842 = ~\mix1_data_o_reg_reg[101]/NET0131  & n1159 ;
  assign n1841 = ~\data_o[101]_pad  & ~n1159 ;
  assign n1843 = n1166 & ~n1841 ;
  assign n1844 = ~n1842 & n1843 ;
  assign n1862 = ~n1840 & ~n1844 ;
  assign n1865 = n1861 & n1862 ;
  assign n1869 = n1864 & n1865 ;
  assign n1870 = n1868 & n1869 ;
  assign n1871 = ~n1256 & ~n1870 ;
  assign n1873 = ~\data_o[125]_pad  & ~n1159 ;
  assign n1872 = ~\mix1_data_o_reg_reg[125]/NET0131  & n1159 ;
  assign n1874 = n1267 & ~n1872 ;
  assign n1875 = ~n1873 & n1874 ;
  assign n1876 = n1266 & n1875 ;
  assign n1877 = ~n1871 & ~n1876 ;
  assign n1878 = n973 & ~n1877 ;
  assign n1879 = \key_i[5]_pad  & ~n1116 ;
  assign n1880 = \ks1_key_reg_reg[5]/NET0131  & n1116 ;
  assign n1881 = ~n1879 & ~n1880 ;
  assign n1882 = n1142 & ~n1881 ;
  assign n1883 = \key_i[21]_pad  & ~n953 ;
  assign n1884 = \ks1_key_reg_reg[21]/NET0131  & n956 ;
  assign n1885 = ~n1883 & ~n1884 ;
  assign n1886 = ~n933 & ~n1885 ;
  assign n1888 = ~\key_i[21]_pad  & n951 ;
  assign n1887 = ~\ks1_key_reg_reg[21]/NET0131  & ~n951 ;
  assign n1889 = n933 & ~n1887 ;
  assign n1890 = ~n1888 & n1889 ;
  assign n1891 = ~n1886 & ~n1890 ;
  assign n1892 = n1286 & ~n1891 ;
  assign n1913 = ~n1882 & ~n1892 ;
  assign n1893 = \key_i[29]_pad  & ~n953 ;
  assign n1894 = \ks1_key_reg_reg[29]/NET0131  & n956 ;
  assign n1895 = ~n1893 & ~n1894 ;
  assign n1896 = ~n933 & ~n1895 ;
  assign n1898 = ~\key_i[29]_pad  & n951 ;
  assign n1897 = ~\ks1_key_reg_reg[29]/NET0131  & ~n951 ;
  assign n1899 = n933 & ~n1897 ;
  assign n1900 = ~n1898 & n1899 ;
  assign n1901 = ~n1896 & ~n1900 ;
  assign n1902 = n971 & ~n1901 ;
  assign n1903 = \key_i[13]_pad  & ~n953 ;
  assign n1904 = \ks1_key_reg_reg[13]/NET0131  & n956 ;
  assign n1905 = ~n1903 & ~n1904 ;
  assign n1906 = ~n933 & ~n1905 ;
  assign n1908 = ~\key_i[13]_pad  & n951 ;
  assign n1907 = ~\ks1_key_reg_reg[13]/NET0131  & ~n951 ;
  assign n1909 = n933 & ~n1907 ;
  assign n1910 = ~n1908 & n1909 ;
  assign n1911 = ~n1906 & ~n1910 ;
  assign n1912 = n1274 & ~n1911 ;
  assign n1914 = ~n1902 & ~n1912 ;
  assign n1915 = n1913 & n1914 ;
  assign n1916 = ~n1878 & n1915 ;
  assign n1917 = n1796 & ~n1916 ;
  assign n1918 = ~n1796 & n1916 ;
  assign n1919 = ~n1917 & ~n1918 ;
  assign n1920 = n1542 & ~n1919 ;
  assign n1921 = ~n1542 & n1919 ;
  assign n1922 = ~n1920 & ~n1921 ;
  assign n1923 = n974 & ~n1922 ;
  assign n1924 = ~n974 & ~n1416 ;
  assign n1925 = ~n1923 & ~n1924 ;
  assign n1926 = n1676 & ~n1925 ;
  assign n1927 = ~n1676 & n1925 ;
  assign n1928 = ~n1926 & ~n1927 ;
  assign n1956 = ~\mix1_data_o_reg_reg[58]/NET0131  & n1159 ;
  assign n1955 = ~\data_o[58]_pad  & ~n1159 ;
  assign n1957 = n1184 & ~n1955 ;
  assign n1958 = ~n1956 & n1957 ;
  assign n1960 = ~\mix1_data_o_reg_reg[98]/NET0131  & n1159 ;
  assign n1959 = ~\data_o[98]_pad  & ~n1159 ;
  assign n1961 = n1166 & ~n1959 ;
  assign n1962 = ~n1960 & n1961 ;
  assign n2001 = ~n1958 & ~n1962 ;
  assign n1964 = ~\mix1_data_o_reg_reg[50]/NET0131  & n1159 ;
  assign n1963 = ~\data_o[50]_pad  & ~n1159 ;
  assign n1965 = n1216 & ~n1963 ;
  assign n1966 = ~n1964 & n1965 ;
  assign n1968 = ~\mix1_data_o_reg_reg[90]/NET0131  & n1159 ;
  assign n1967 = ~\data_o[90]_pad  & ~n1159 ;
  assign n1969 = n1227 & ~n1967 ;
  assign n1970 = ~n1968 & n1969 ;
  assign n2002 = ~n1966 & ~n1970 ;
  assign n2008 = n2001 & n2002 ;
  assign n1940 = ~\mix1_data_o_reg_reg[106]/NET0131  & n1159 ;
  assign n1939 = ~\data_o[106]_pad  & ~n1159 ;
  assign n1941 = n1237 & ~n1939 ;
  assign n1942 = ~n1940 & n1941 ;
  assign n1944 = ~\mix1_data_o_reg_reg[82]/NET0131  & n1159 ;
  assign n1943 = ~\data_o[82]_pad  & ~n1159 ;
  assign n1945 = n1222 & ~n1943 ;
  assign n1946 = ~n1944 & n1945 ;
  assign n1999 = ~n1942 & ~n1946 ;
  assign n1948 = ~\mix1_data_o_reg_reg[114]/NET0131  & n1159 ;
  assign n1947 = ~\data_o[114]_pad  & ~n1159 ;
  assign n1949 = n1189 & ~n1947 ;
  assign n1950 = ~n1948 & n1949 ;
  assign n1952 = ~\mix1_data_o_reg_reg[18]/NET0131  & n1159 ;
  assign n1951 = ~\data_o[18]_pad  & ~n1159 ;
  assign n1953 = n1178 & ~n1951 ;
  assign n1954 = ~n1952 & n1953 ;
  assign n2000 = ~n1950 & ~n1954 ;
  assign n2009 = n1999 & n2000 ;
  assign n2010 = n2008 & n2009 ;
  assign n1996 = ~\mix1_data_o_reg_reg[34]/NET0131  & n1159 ;
  assign n1995 = ~\data_o[34]_pad  & ~n1159 ;
  assign n1997 = n1211 & ~n1995 ;
  assign n1998 = ~n1996 & n1997 ;
  assign n1988 = ~\mix1_data_o_reg_reg[74]/NET0131  & n1159 ;
  assign n1987 = ~\data_o[74]_pad  & ~n1159 ;
  assign n1989 = n1232 & ~n1987 ;
  assign n1990 = ~n1988 & n1989 ;
  assign n1992 = ~\mix1_data_o_reg_reg[2]/NET0131  & n1159 ;
  assign n1991 = ~\data_o[2]_pad  & ~n1159 ;
  assign n1993 = n1201 & ~n1991 ;
  assign n1994 = ~n1992 & n1993 ;
  assign n2005 = ~n1990 & ~n1994 ;
  assign n2006 = ~n1998 & n2005 ;
  assign n1972 = ~\mix1_data_o_reg_reg[42]/NET0131  & n1159 ;
  assign n1971 = ~\data_o[42]_pad  & ~n1159 ;
  assign n1973 = n1195 & ~n1971 ;
  assign n1974 = ~n1972 & n1973 ;
  assign n1976 = ~\mix1_data_o_reg_reg[26]/NET0131  & n1159 ;
  assign n1975 = ~\data_o[26]_pad  & ~n1159 ;
  assign n1977 = n1172 & ~n1975 ;
  assign n1978 = ~n1976 & n1977 ;
  assign n2003 = ~n1974 & ~n1978 ;
  assign n1980 = ~\mix1_data_o_reg_reg[66]/NET0131  & n1159 ;
  assign n1979 = ~\data_o[66]_pad  & ~n1159 ;
  assign n1981 = n1206 & ~n1979 ;
  assign n1982 = ~n1980 & n1981 ;
  assign n1984 = ~\mix1_data_o_reg_reg[10]/NET0131  & n1159 ;
  assign n1983 = ~\data_o[10]_pad  & ~n1159 ;
  assign n1985 = n1155 & ~n1983 ;
  assign n1986 = ~n1984 & n1985 ;
  assign n2004 = ~n1982 & ~n1986 ;
  assign n2007 = n2003 & n2004 ;
  assign n2011 = n2006 & n2007 ;
  assign n2012 = n2010 & n2011 ;
  assign n2013 = ~n1256 & ~n2012 ;
  assign n2015 = ~\data_o[122]_pad  & ~n1159 ;
  assign n2014 = ~\mix1_data_o_reg_reg[122]/NET0131  & n1159 ;
  assign n2016 = n1267 & ~n2014 ;
  assign n2017 = ~n2015 & n2016 ;
  assign n2018 = n1266 & n2017 ;
  assign n2019 = ~n2013 & ~n2018 ;
  assign n2020 = n973 & ~n2019 ;
  assign n1929 = \key_i[26]_pad  & ~n953 ;
  assign n1930 = \ks1_key_reg_reg[26]/NET0131  & n956 ;
  assign n1931 = ~n1929 & ~n1930 ;
  assign n1932 = ~n933 & ~n1931 ;
  assign n1934 = ~\key_i[26]_pad  & n951 ;
  assign n1933 = ~\ks1_key_reg_reg[26]/NET0131  & ~n951 ;
  assign n1935 = n933 & ~n1933 ;
  assign n1936 = ~n1934 & n1935 ;
  assign n1937 = ~n1932 & ~n1936 ;
  assign n1938 = n971 & ~n1937 ;
  assign n2021 = \key_i[18]_pad  & ~n953 ;
  assign n2022 = \ks1_key_reg_reg[18]/NET0131  & n956 ;
  assign n2023 = ~n2021 & ~n2022 ;
  assign n2024 = ~n933 & ~n2023 ;
  assign n2026 = ~\key_i[18]_pad  & n951 ;
  assign n2025 = ~\ks1_key_reg_reg[18]/NET0131  & ~n951 ;
  assign n2027 = n933 & ~n2025 ;
  assign n2028 = ~n2026 & n2027 ;
  assign n2029 = ~n2024 & ~n2028 ;
  assign n2030 = n1286 & ~n2029 ;
  assign n2051 = ~n1938 & ~n2030 ;
  assign n2031 = \key_i[10]_pad  & ~n953 ;
  assign n2032 = \ks1_key_reg_reg[10]/NET0131  & n956 ;
  assign n2033 = ~n2031 & ~n2032 ;
  assign n2034 = ~n933 & ~n2033 ;
  assign n2036 = ~\key_i[10]_pad  & n951 ;
  assign n2035 = ~\ks1_key_reg_reg[10]/NET0131  & ~n951 ;
  assign n2037 = n933 & ~n2035 ;
  assign n2038 = ~n2036 & n2037 ;
  assign n2039 = ~n2034 & ~n2038 ;
  assign n2040 = n1274 & ~n2039 ;
  assign n2041 = \key_i[2]_pad  & ~n953 ;
  assign n2042 = \ks1_key_reg_reg[2]/NET0131  & n956 ;
  assign n2043 = ~n2041 & ~n2042 ;
  assign n2044 = ~n933 & ~n2043 ;
  assign n2046 = ~\key_i[2]_pad  & n951 ;
  assign n2045 = ~\ks1_key_reg_reg[2]/NET0131  & ~n951 ;
  assign n2047 = n933 & ~n2045 ;
  assign n2048 = ~n2046 & n2047 ;
  assign n2049 = ~n2044 & ~n2048 ;
  assign n2050 = n1142 & ~n2049 ;
  assign n2052 = ~n2040 & ~n2050 ;
  assign n2053 = n2051 & n2052 ;
  assign n2054 = ~n2020 & n2053 ;
  assign n2055 = ~n974 & ~n2054 ;
  assign n2056 = \key_i[23]_pad  & ~n953 ;
  assign n2057 = \ks1_key_reg_reg[23]/NET0131  & n956 ;
  assign n2058 = ~n2056 & ~n2057 ;
  assign n2059 = ~n933 & ~n2058 ;
  assign n2061 = ~\key_i[23]_pad  & n951 ;
  assign n2060 = ~\ks1_key_reg_reg[23]/NET0131  & ~n951 ;
  assign n2062 = n933 & ~n2060 ;
  assign n2063 = ~n2061 & n2062 ;
  assign n2064 = ~n2059 & ~n2063 ;
  assign n2065 = n1286 & ~n2064 ;
  assign n2066 = \key_i[7]_pad  & ~n953 ;
  assign n2067 = \ks1_key_reg_reg[7]/NET0131  & n956 ;
  assign n2068 = ~n2066 & ~n2067 ;
  assign n2069 = ~n933 & ~n2068 ;
  assign n2071 = ~\key_i[7]_pad  & n951 ;
  assign n2070 = ~\ks1_key_reg_reg[7]/NET0131  & ~n951 ;
  assign n2072 = n933 & ~n2070 ;
  assign n2073 = ~n2071 & n2072 ;
  assign n2074 = ~n2069 & ~n2073 ;
  assign n2075 = n1142 & ~n2074 ;
  assign n2096 = ~n2065 & ~n2075 ;
  assign n2076 = \key_i[15]_pad  & ~n953 ;
  assign n2077 = \ks1_key_reg_reg[15]/NET0131  & n956 ;
  assign n2078 = ~n2076 & ~n2077 ;
  assign n2079 = ~n933 & ~n2078 ;
  assign n2081 = ~\key_i[15]_pad  & n951 ;
  assign n2080 = ~\ks1_key_reg_reg[15]/NET0131  & ~n951 ;
  assign n2082 = n933 & ~n2080 ;
  assign n2083 = ~n2081 & n2082 ;
  assign n2084 = ~n2079 & ~n2083 ;
  assign n2085 = n1274 & ~n2084 ;
  assign n2086 = \key_i[31]_pad  & ~n953 ;
  assign n2087 = \ks1_key_reg_reg[31]/NET0131  & n956 ;
  assign n2088 = ~n2086 & ~n2087 ;
  assign n2089 = ~n933 & ~n2088 ;
  assign n2091 = ~\key_i[31]_pad  & n951 ;
  assign n2090 = ~\ks1_key_reg_reg[31]/NET0131  & ~n951 ;
  assign n2092 = n933 & ~n2090 ;
  assign n2093 = ~n2091 & n2092 ;
  assign n2094 = ~n2089 & ~n2093 ;
  assign n2095 = n971 & ~n2094 ;
  assign n2097 = ~n2085 & ~n2095 ;
  assign n2098 = n2096 & n2097 ;
  assign n2099 = ~n973 & ~n2098 ;
  assign n2117 = ~\mix1_data_o_reg_reg[87]/NET0131  & n1159 ;
  assign n2116 = ~\data_o[87]_pad  & ~n1159 ;
  assign n2118 = n1222 & ~n2116 ;
  assign n2119 = ~n2117 & n2118 ;
  assign n2121 = ~\mix1_data_o_reg_reg[63]/NET0131  & n1159 ;
  assign n2120 = ~\data_o[63]_pad  & ~n1159 ;
  assign n2122 = n1184 & ~n2120 ;
  assign n2123 = ~n2121 & n2122 ;
  assign n2162 = ~n2119 & ~n2123 ;
  assign n2125 = ~\mix1_data_o_reg_reg[55]/NET0131  & n1159 ;
  assign n2124 = ~\data_o[55]_pad  & ~n1159 ;
  assign n2126 = n1216 & ~n2124 ;
  assign n2127 = ~n2125 & n2126 ;
  assign n2129 = ~\mix1_data_o_reg_reg[95]/NET0131  & n1159 ;
  assign n2128 = ~\data_o[95]_pad  & ~n1159 ;
  assign n2130 = n1227 & ~n2128 ;
  assign n2131 = ~n2129 & n2130 ;
  assign n2163 = ~n2127 & ~n2131 ;
  assign n2169 = n2162 & n2163 ;
  assign n2101 = ~\mix1_data_o_reg_reg[15]/NET0131  & n1159 ;
  assign n2100 = ~\data_o[15]_pad  & ~n1159 ;
  assign n2102 = n1155 & ~n2100 ;
  assign n2103 = ~n2101 & n2102 ;
  assign n2105 = ~\mix1_data_o_reg_reg[39]/NET0131  & n1159 ;
  assign n2104 = ~\data_o[39]_pad  & ~n1159 ;
  assign n2106 = n1211 & ~n2104 ;
  assign n2107 = ~n2105 & n2106 ;
  assign n2160 = ~n2103 & ~n2107 ;
  assign n2109 = ~\mix1_data_o_reg_reg[31]/NET0131  & n1159 ;
  assign n2108 = ~\data_o[31]_pad  & ~n1159 ;
  assign n2110 = n1172 & ~n2108 ;
  assign n2111 = ~n2109 & n2110 ;
  assign n2113 = ~\mix1_data_o_reg_reg[23]/NET0131  & n1159 ;
  assign n2112 = ~\data_o[23]_pad  & ~n1159 ;
  assign n2114 = n1178 & ~n2112 ;
  assign n2115 = ~n2113 & n2114 ;
  assign n2161 = ~n2111 & ~n2115 ;
  assign n2170 = n2160 & n2161 ;
  assign n2171 = n2169 & n2170 ;
  assign n2157 = ~\mix1_data_o_reg_reg[119]/NET0131  & n1159 ;
  assign n2156 = ~\data_o[119]_pad  & ~n1159 ;
  assign n2158 = n1189 & ~n2156 ;
  assign n2159 = ~n2157 & n2158 ;
  assign n2149 = ~\mix1_data_o_reg_reg[79]/NET0131  & n1159 ;
  assign n2148 = ~\data_o[79]_pad  & ~n1159 ;
  assign n2150 = n1232 & ~n2148 ;
  assign n2151 = ~n2149 & n2150 ;
  assign n2153 = ~\mix1_data_o_reg_reg[7]/NET0131  & n1159 ;
  assign n2152 = ~\data_o[7]_pad  & ~n1159 ;
  assign n2154 = n1201 & ~n2152 ;
  assign n2155 = ~n2153 & n2154 ;
  assign n2166 = ~n2151 & ~n2155 ;
  assign n2167 = ~n2159 & n2166 ;
  assign n2133 = ~\mix1_data_o_reg_reg[47]/NET0131  & n1159 ;
  assign n2132 = ~\data_o[47]_pad  & ~n1159 ;
  assign n2134 = n1195 & ~n2132 ;
  assign n2135 = ~n2133 & n2134 ;
  assign n2137 = ~\mix1_data_o_reg_reg[103]/NET0131  & n1159 ;
  assign n2136 = ~\data_o[103]_pad  & ~n1159 ;
  assign n2138 = n1166 & ~n2136 ;
  assign n2139 = ~n2137 & n2138 ;
  assign n2164 = ~n2135 & ~n2139 ;
  assign n2141 = ~\mix1_data_o_reg_reg[71]/NET0131  & n1159 ;
  assign n2140 = ~\data_o[71]_pad  & ~n1159 ;
  assign n2142 = n1206 & ~n2140 ;
  assign n2143 = ~n2141 & n2142 ;
  assign n2145 = ~\mix1_data_o_reg_reg[111]/NET0131  & n1159 ;
  assign n2144 = ~\data_o[111]_pad  & ~n1159 ;
  assign n2146 = n1237 & ~n2144 ;
  assign n2147 = ~n2145 & n2146 ;
  assign n2165 = ~n2143 & ~n2147 ;
  assign n2168 = n2164 & n2165 ;
  assign n2172 = n2167 & n2168 ;
  assign n2173 = n2171 & n2172 ;
  assign n2174 = ~n1256 & ~n2173 ;
  assign n2176 = ~\data_o[127]_pad  & ~n1159 ;
  assign n2175 = ~\mix1_data_o_reg_reg[127]/NET0131  & n1159 ;
  assign n2177 = n1267 & ~n2175 ;
  assign n2178 = ~n2176 & n2177 ;
  assign n2179 = n1266 & n2178 ;
  assign n2180 = ~n2174 & ~n2179 ;
  assign n2181 = n973 & ~n2180 ;
  assign n2182 = ~n2099 & ~n2181 ;
  assign n2183 = ~n1310 & n1671 ;
  assign n2184 = n1310 & ~n1671 ;
  assign n2185 = ~n2183 & ~n2184 ;
  assign n2187 = n2182 & ~n2185 ;
  assign n2186 = ~n2182 & n2185 ;
  assign n2188 = n974 & ~n2186 ;
  assign n2189 = ~n2187 & n2188 ;
  assign n2190 = ~n2055 & ~n2189 ;
  assign n2191 = ~n1676 & ~n2190 ;
  assign n2192 = n1676 & n2190 ;
  assign n2193 = ~n2191 & ~n2192 ;
  assign n2194 = n2054 & ~n2182 ;
  assign n2195 = ~n2054 & n2182 ;
  assign n2196 = ~n2194 & ~n2195 ;
  assign n2197 = n1310 & ~n2196 ;
  assign n2198 = ~n1310 & n2196 ;
  assign n2199 = ~n2197 & ~n2198 ;
  assign n2200 = n974 & ~n2199 ;
  assign n2201 = ~n974 & ~n1916 ;
  assign n2202 = ~n2200 & ~n2201 ;
  assign n2203 = n1928 & ~n2202 ;
  assign n2204 = ~n1928 & n2202 ;
  assign n2205 = ~n2203 & ~n2204 ;
  assign n2206 = ~n2193 & n2205 ;
  assign n2207 = n2193 & ~n2205 ;
  assign n2208 = ~n2206 & ~n2207 ;
  assign n2209 = n1916 & ~n2196 ;
  assign n2210 = ~n1916 & n2196 ;
  assign n2211 = ~n2209 & ~n2210 ;
  assign n2212 = n974 & ~n2211 ;
  assign n2213 = ~n974 & n1796 ;
  assign n2214 = ~n2212 & ~n2213 ;
  assign n2215 = n2208 & ~n2214 ;
  assign n2216 = ~n2208 & n2214 ;
  assign n2217 = ~n2215 & ~n2216 ;
  assign n2218 = n1928 & ~n2217 ;
  assign n2219 = ~n974 & ~n1671 ;
  assign n2221 = ~n1545 & ~n1796 ;
  assign n2220 = n1545 & n1796 ;
  assign n2222 = n974 & ~n2220 ;
  assign n2223 = ~n2221 & n2222 ;
  assign n2224 = ~n2219 & ~n2223 ;
  assign n2225 = ~n974 & ~n2182 ;
  assign n2227 = ~n1416 & ~n2185 ;
  assign n2226 = n1416 & n2185 ;
  assign n2228 = n974 & ~n2226 ;
  assign n2229 = ~n2227 & n2228 ;
  assign n2230 = ~n2225 & ~n2229 ;
  assign n2231 = ~n2224 & ~n2230 ;
  assign n2232 = n2224 & n2230 ;
  assign n2233 = ~n2231 & ~n2232 ;
  assign n2234 = n2217 & ~n2233 ;
  assign n2235 = ~n2218 & ~n2234 ;
  assign n2236 = ~n2190 & ~n2224 ;
  assign n2237 = n2190 & n2224 ;
  assign n2238 = ~n2236 & ~n2237 ;
  assign n2239 = ~n2205 & ~n2238 ;
  assign n2240 = ~n2193 & ~n2233 ;
  assign n2241 = n2193 & n2233 ;
  assign n2242 = ~n2240 & ~n2241 ;
  assign n2243 = n2202 & ~n2230 ;
  assign n2244 = ~n2202 & n2230 ;
  assign n2245 = ~n2243 & ~n2244 ;
  assign n2246 = n1919 & ~n2054 ;
  assign n2247 = ~n1919 & n2054 ;
  assign n2248 = ~n2246 & ~n2247 ;
  assign n2249 = n974 & ~n2248 ;
  assign n2250 = ~n974 & ~n1542 ;
  assign n2251 = ~n2249 & ~n2250 ;
  assign n2252 = n2190 & ~n2251 ;
  assign n2253 = ~n2190 & n2251 ;
  assign n2254 = ~n2252 & ~n2253 ;
  assign n2255 = n2245 & n2254 ;
  assign n2256 = ~n2245 & ~n2254 ;
  assign n2257 = ~n2255 & ~n2256 ;
  assign n2258 = n2242 & n2257 ;
  assign n2259 = n2239 & ~n2258 ;
  assign n2260 = ~n2239 & n2258 ;
  assign n2261 = ~n2259 & ~n2260 ;
  assign n2262 = n2190 & ~n2243 ;
  assign n2263 = ~n2190 & ~n2244 ;
  assign n2264 = ~n2262 & ~n2263 ;
  assign n2265 = n2261 & ~n2264 ;
  assign n2266 = ~n2261 & n2264 ;
  assign n2267 = ~n2265 & ~n2266 ;
  assign n2268 = n2235 & n2267 ;
  assign n2269 = ~n2235 & ~n2267 ;
  assign n2270 = ~n2268 & ~n2269 ;
  assign n2271 = n2238 & n2257 ;
  assign n2272 = n2206 & ~n2271 ;
  assign n2273 = ~n2206 & n2271 ;
  assign n2274 = ~n2272 & ~n2273 ;
  assign n2275 = ~n1928 & ~n2233 ;
  assign n2276 = ~n2217 & ~n2245 ;
  assign n2277 = n2275 & ~n2276 ;
  assign n2278 = ~n2275 & n2276 ;
  assign n2279 = ~n2277 & ~n2278 ;
  assign n2280 = n2274 & n2279 ;
  assign n2281 = ~n2274 & ~n2279 ;
  assign n2282 = ~n2280 & ~n2281 ;
  assign n2283 = ~n2217 & n2257 ;
  assign n2284 = ~n2205 & n2233 ;
  assign n2285 = ~n2193 & ~n2245 ;
  assign n2286 = n2284 & ~n2285 ;
  assign n2287 = n2242 & ~n2245 ;
  assign n2288 = ~n2284 & n2287 ;
  assign n2289 = ~n2286 & ~n2288 ;
  assign n2290 = n2283 & ~n2289 ;
  assign n2291 = ~n2283 & n2289 ;
  assign n2292 = ~n2290 & ~n2291 ;
  assign n2293 = n1928 & n2233 ;
  assign n2294 = ~n2275 & ~n2293 ;
  assign n2295 = n2238 & ~n2294 ;
  assign n2296 = ~n1676 & n2295 ;
  assign n2297 = n1676 & ~n2295 ;
  assign n2298 = ~n2296 & ~n2297 ;
  assign n2299 = n2292 & n2298 ;
  assign n2300 = ~n2292 & ~n2298 ;
  assign n2301 = ~n2299 & ~n2300 ;
  assign n2302 = \sbox1_alph_reg[1]/NET0131  & n982 ;
  assign n2303 = \sbox1_alph_reg[3]/NET0131  & n999 ;
  assign n2304 = \sbox1_alph_reg[2]/NET0131  & ~n1007 ;
  assign n2305 = \sbox1_alph_reg[0]/NET0131  & ~n992 ;
  assign n2306 = n2304 & ~n2305 ;
  assign n2307 = ~n2304 & n2305 ;
  assign n2308 = ~n2306 & ~n2307 ;
  assign n2309 = n2303 & n2308 ;
  assign n2310 = ~n2303 & ~n2308 ;
  assign n2311 = ~n2309 & ~n2310 ;
  assign n2312 = n2302 & ~n2311 ;
  assign n2313 = ~n2302 & n2311 ;
  assign n2314 = ~n2312 & ~n2313 ;
  assign n2315 = n1017 & n2314 ;
  assign n2316 = ~n1017 & ~n2314 ;
  assign n2317 = ~n2315 & ~n2316 ;
  assign n2318 = ~n1017 & ~n1106 ;
  assign n2319 = n1017 & n1106 ;
  assign n2320 = ~n2318 & ~n2319 ;
  assign n2321 = \sbox1_ah_reg_reg[2]/NET0131  & ~n982 ;
  assign n2322 = n999 & ~n1026 ;
  assign n2323 = ~n2321 & n2322 ;
  assign n2324 = n2321 & ~n2322 ;
  assign n2325 = ~n2323 & ~n2324 ;
  assign n2326 = \sbox1_ah_reg_reg[1]/NET0131  & ~n992 ;
  assign n2327 = n2325 & ~n2326 ;
  assign n2328 = ~n2325 & n2326 ;
  assign n2329 = ~n2327 & ~n2328 ;
  assign n2330 = \sbox1_ah_reg_reg[3]/NET0131  & ~n1007 ;
  assign n2331 = \sbox1_ah_reg_reg[2]/NET0131  & n1007 ;
  assign n2332 = ~n2330 & ~n2331 ;
  assign n2333 = ~n1014 & n2332 ;
  assign n2334 = n1014 & ~n2332 ;
  assign n2335 = ~n2333 & ~n2334 ;
  assign n2336 = n2329 & n2335 ;
  assign n2337 = ~n2329 & ~n2335 ;
  assign n2338 = ~n2336 & ~n2337 ;
  assign n2339 = n2320 & n2338 ;
  assign n2340 = ~n2320 & ~n2338 ;
  assign n2341 = ~n2339 & ~n2340 ;
  assign n2343 = n1109 & n2341 ;
  assign n2342 = ~n1109 & ~n2341 ;
  assign n2344 = ~n974 & ~n2342 ;
  assign n2345 = ~n2343 & n2344 ;
  assign n2346 = n2317 & n2345 ;
  assign n2347 = ~n2317 & ~n2345 ;
  assign n2348 = ~n2346 & ~n2347 ;
  assign n2349 = ~\ks1_key_reg_reg[104]/NET0131  & n1116 ;
  assign n2350 = ~\key_i[104]_pad  & ~n1116 ;
  assign n2351 = ~n2349 & ~n2350 ;
  assign n2352 = n2348 & ~n2351 ;
  assign n2353 = ~n2348 & n2351 ;
  assign n2354 = ~n2352 & ~n2353 ;
  assign n2355 = ~\ks1_key_reg_reg[72]/P0002  & n1116 ;
  assign n2356 = ~\key_i[72]_pad  & ~n1116 ;
  assign n2357 = ~n2355 & ~n2356 ;
  assign n2358 = n2354 & ~n2357 ;
  assign n2359 = ~n2354 & n2357 ;
  assign n2360 = ~n2358 & ~n2359 ;
  assign n2361 = ~\ks1_key_reg_reg[40]/P0002  & n1116 ;
  assign n2362 = ~\key_i[40]_pad  & ~n1116 ;
  assign n2363 = ~n2361 & ~n2362 ;
  assign n2364 = n2360 & ~n2363 ;
  assign n2365 = ~n2360 & n2363 ;
  assign n2366 = ~n2364 & ~n2365 ;
  assign n2367 = n1771 & ~n2366 ;
  assign n2368 = ~n1771 & n2366 ;
  assign n2369 = ~n2367 & ~n2368 ;
  assign n2370 = n929 & ~n2369 ;
  assign n2371 = \ks1_key_reg_reg[8]/NET0131  & ~n929 ;
  assign n2372 = ~n2370 & ~n2371 ;
  assign n2373 = \ks1_key_reg_reg[10]/NET0131  & ~n929 ;
  assign n2374 = \key_i[74]_pad  & ~n1116 ;
  assign n2375 = \ks1_key_reg_reg[74]/NET0131  & n1116 ;
  assign n2376 = ~n2374 & ~n2375 ;
  assign n2377 = \key_i[106]_pad  & ~n953 ;
  assign n2378 = \ks1_key_reg_reg[106]/NET0131  & n956 ;
  assign n2379 = ~n2377 & ~n2378 ;
  assign n2380 = ~n933 & ~n2379 ;
  assign n2382 = ~\key_i[106]_pad  & n951 ;
  assign n2381 = ~\ks1_key_reg_reg[106]/NET0131  & ~n951 ;
  assign n2383 = n933 & ~n2381 ;
  assign n2384 = ~n2382 & n2383 ;
  assign n2385 = ~n2380 & ~n2384 ;
  assign n2386 = n1090 & n2317 ;
  assign n2387 = ~n1090 & ~n2317 ;
  assign n2388 = ~n2386 & ~n2387 ;
  assign n2389 = n1033 & n2338 ;
  assign n2390 = ~n1033 & ~n2338 ;
  assign n2391 = ~n2389 & ~n2390 ;
  assign n2392 = ~n2317 & ~n2391 ;
  assign n2393 = n2317 & n2391 ;
  assign n2394 = ~n2392 & ~n2393 ;
  assign n2395 = n974 & ~n2394 ;
  assign n2396 = ~n974 & n2341 ;
  assign n2397 = ~n2395 & ~n2396 ;
  assign n2398 = n2388 & ~n2397 ;
  assign n2399 = ~n2388 & n2397 ;
  assign n2400 = ~n2398 & ~n2399 ;
  assign n2401 = n2385 & n2400 ;
  assign n2402 = ~n2385 & ~n2400 ;
  assign n2403 = ~n2401 & ~n2402 ;
  assign n2404 = n2376 & n2403 ;
  assign n2405 = ~n2376 & ~n2403 ;
  assign n2406 = ~n2404 & ~n2405 ;
  assign n2407 = ~\ks1_key_reg_reg[42]/P0002  & n1116 ;
  assign n2408 = ~\key_i[42]_pad  & ~n1116 ;
  assign n2409 = ~n2407 & ~n2408 ;
  assign n2410 = n2406 & ~n2409 ;
  assign n2411 = ~n2406 & n2409 ;
  assign n2412 = ~n2410 & ~n2411 ;
  assign n2414 = ~n2039 & ~n2412 ;
  assign n2413 = n2039 & n2412 ;
  assign n2415 = n929 & ~n2413 ;
  assign n2416 = ~n2414 & n2415 ;
  assign n2417 = ~n2373 & ~n2416 ;
  assign n2424 = \sub1_state_reg[2]/NET0131  & ~n1171 ;
  assign n2425 = ~n1183 & ~n2424 ;
  assign n2426 = ~\sub1_state_reg[4]/NET0131  & n2425 ;
  assign n2427 = ~n1165 & ~n1171 ;
  assign n2428 = n2426 & ~n2427 ;
  assign n2429 = \sub1_state_reg[3]/NET0131  & ~n1183 ;
  assign n2430 = ~n1256 & ~n2429 ;
  assign n2431 = ~\sub1_state_reg[0]/NET0131  & n2430 ;
  assign n2432 = n2428 & n2431 ;
  assign n2434 = n1114 & n2432 ;
  assign n2433 = ~\sub1_data_reg_reg[102]/NET0131  & ~n2432 ;
  assign n2435 = ~n1256 & ~n2433 ;
  assign n2436 = ~n2434 & n2435 ;
  assign n2418 = \sub1_data_reg_reg[102]/NET0131  & n1267 ;
  assign n2419 = ~decrypt_i_pad & ~n1058 ;
  assign n2420 = decrypt_i_pad & ~\sub1_data_reg_reg[70]/NET0131  ;
  assign n2421 = \sub1_state_reg[4]/NET0131  & n1256 ;
  assign n2422 = ~n2420 & n2421 ;
  assign n2423 = ~n2419 & n2422 ;
  assign n2437 = ~n2418 & ~n2423 ;
  assign n2438 = ~n2436 & n2437 ;
  assign n2451 = n1072 & ~n2338 ;
  assign n2452 = ~n1072 & n2338 ;
  assign n2453 = ~n2451 & ~n2452 ;
  assign n2454 = n974 & ~n2453 ;
  assign n2440 = n1052 & n2338 ;
  assign n2441 = ~n1052 & ~n2338 ;
  assign n2442 = ~n2440 & ~n2441 ;
  assign n2443 = ~n1109 & ~n2442 ;
  assign n2444 = n1109 & n2442 ;
  assign n2445 = ~n2443 & ~n2444 ;
  assign n2455 = ~n974 & n2445 ;
  assign n2456 = ~n2454 & ~n2455 ;
  assign n2457 = n2432 & ~n2456 ;
  assign n2450 = ~\sub1_data_reg_reg[101]/NET0131  & ~n2432 ;
  assign n2458 = ~n1256 & ~n2450 ;
  assign n2459 = ~n2457 & n2458 ;
  assign n2439 = \sub1_data_reg_reg[101]/NET0131  & n1267 ;
  assign n2446 = ~decrypt_i_pad & n2445 ;
  assign n2447 = decrypt_i_pad & ~\sub1_data_reg_reg[69]/NET0131  ;
  assign n2448 = n2421 & ~n2447 ;
  assign n2449 = ~n2446 & n2448 ;
  assign n2460 = ~n2439 & ~n2449 ;
  assign n2461 = ~n2459 & n2460 ;
  assign n2467 = n2426 & n2427 ;
  assign n2468 = n2431 & n2467 ;
  assign n2470 = ~n2456 & n2468 ;
  assign n2469 = ~\sub1_data_reg_reg[117]/NET0131  & ~n2468 ;
  assign n2471 = ~n1256 & ~n2469 ;
  assign n2472 = ~n2470 & n2471 ;
  assign n2462 = \sub1_data_reg_reg[117]/NET0131  & n1267 ;
  assign n2463 = ~decrypt_i_pad & ~\sub1_data_reg_reg[85]/NET0131  ;
  assign n2464 = decrypt_i_pad & ~\sub1_data_reg_reg[21]/NET0131  ;
  assign n2465 = ~n2463 & ~n2464 ;
  assign n2466 = n2421 & n2465 ;
  assign n2473 = ~n2462 & ~n2466 ;
  assign n2474 = ~n2472 & n2473 ;
  assign n2481 = n1114 & n2468 ;
  assign n2480 = ~\sub1_data_reg_reg[118]/NET0131  & ~n2468 ;
  assign n2482 = ~n1256 & ~n2480 ;
  assign n2483 = ~n2481 & n2482 ;
  assign n2475 = \sub1_data_reg_reg[118]/NET0131  & n1267 ;
  assign n2476 = ~decrypt_i_pad & ~\sub1_data_reg_reg[86]/NET0131  ;
  assign n2477 = decrypt_i_pad & ~\sub1_data_reg_reg[22]/NET0131  ;
  assign n2478 = ~n2476 & ~n2477 ;
  assign n2479 = n2421 & n2478 ;
  assign n2484 = ~n2475 & ~n2479 ;
  assign n2485 = ~n2483 & n2484 ;
  assign n2491 = \sub1_state_reg[4]/NET0131  & ~n1256 ;
  assign n2492 = ~n1267 & ~n2425 ;
  assign n2493 = ~n2491 & n2492 ;
  assign n2494 = n2427 & n2493 ;
  assign n2495 = ~\sub1_state_reg[0]/NET0131  & ~n1267 ;
  assign n2496 = ~n2430 & n2495 ;
  assign n2497 = n2494 & n2496 ;
  assign n2499 = ~n2456 & n2497 ;
  assign n2498 = ~\sub1_data_reg_reg[21]/NET0131  & ~n2497 ;
  assign n2500 = ~n1256 & ~n2498 ;
  assign n2501 = ~n2499 & n2500 ;
  assign n2486 = \sub1_data_reg_reg[21]/NET0131  & n1267 ;
  assign n2487 = ~decrypt_i_pad & ~\sub1_data_reg_reg[117]/NET0131  ;
  assign n2488 = decrypt_i_pad & ~\sub1_data_reg_reg[53]/NET0131  ;
  assign n2489 = ~n2487 & ~n2488 ;
  assign n2490 = n2421 & n2489 ;
  assign n2502 = ~n2486 & ~n2490 ;
  assign n2503 = ~n2501 & n2502 ;
  assign n2510 = n1114 & n2497 ;
  assign n2509 = ~\sub1_data_reg_reg[22]/NET0131  & ~n2497 ;
  assign n2511 = ~n1256 & ~n2509 ;
  assign n2512 = ~n2510 & n2511 ;
  assign n2504 = \sub1_data_reg_reg[22]/NET0131  & n1267 ;
  assign n2505 = ~decrypt_i_pad & ~\sub1_data_reg_reg[118]/NET0131  ;
  assign n2506 = decrypt_i_pad & ~\sub1_data_reg_reg[54]/NET0131  ;
  assign n2507 = ~n2505 & ~n2506 ;
  assign n2508 = n2421 & n2507 ;
  assign n2513 = ~n2504 & ~n2508 ;
  assign n2514 = ~n2512 & n2513 ;
  assign n2515 = n2428 & n2496 ;
  assign n2516 = ~n2456 & n2515 ;
  assign n2517 = ~n1256 & ~n2516 ;
  assign n2519 = ~n1267 & ~n2517 ;
  assign n2520 = \sub1_data_reg_reg[37]/NET0131  & ~n2519 ;
  assign n2518 = n2515 & n2517 ;
  assign n2522 = decrypt_i_pad & ~n2456 ;
  assign n2521 = ~decrypt_i_pad & ~\sub1_data_reg_reg[69]/NET0131  ;
  assign n2523 = n2421 & ~n2521 ;
  assign n2524 = ~n2522 & n2523 ;
  assign n2525 = ~n2518 & ~n2524 ;
  assign n2526 = ~n2520 & n2525 ;
  assign n2533 = decrypt_i_pad & n1114 ;
  assign n2532 = ~decrypt_i_pad & ~\sub1_data_reg_reg[70]/NET0131  ;
  assign n2534 = n2421 & ~n2532 ;
  assign n2535 = ~n2533 & n2534 ;
  assign n2527 = \sub1_data_reg_reg[38]/NET0131  & n1267 ;
  assign n2529 = n1114 & n2515 ;
  assign n2528 = ~\sub1_data_reg_reg[38]/NET0131  & ~n2515 ;
  assign n2530 = ~n1256 & ~n2528 ;
  assign n2531 = ~n2529 & n2530 ;
  assign n2536 = ~n2527 & ~n2531 ;
  assign n2537 = ~n2535 & n2536 ;
  assign n2543 = n2467 & n2496 ;
  assign n2545 = ~n2456 & n2543 ;
  assign n2544 = ~\sub1_data_reg_reg[53]/NET0131  & ~n2543 ;
  assign n2546 = ~n1256 & ~n2544 ;
  assign n2547 = ~n2545 & n2546 ;
  assign n2538 = \sub1_data_reg_reg[53]/NET0131  & n1267 ;
  assign n2539 = ~decrypt_i_pad & ~\sub1_data_reg_reg[21]/NET0131  ;
  assign n2540 = decrypt_i_pad & ~\sub1_data_reg_reg[85]/NET0131  ;
  assign n2541 = ~n2539 & ~n2540 ;
  assign n2542 = n2421 & n2541 ;
  assign n2548 = ~n2538 & ~n2542 ;
  assign n2549 = ~n2547 & n2548 ;
  assign n2556 = n1114 & n2543 ;
  assign n2555 = ~\sub1_data_reg_reg[54]/NET0131  & ~n2543 ;
  assign n2557 = ~n1256 & ~n2555 ;
  assign n2558 = ~n2556 & n2557 ;
  assign n2550 = \sub1_data_reg_reg[54]/NET0131  & n1267 ;
  assign n2551 = ~decrypt_i_pad & ~\sub1_data_reg_reg[22]/NET0131  ;
  assign n2552 = decrypt_i_pad & ~\sub1_data_reg_reg[86]/NET0131  ;
  assign n2553 = ~n2551 & ~n2552 ;
  assign n2554 = n2421 & n2553 ;
  assign n2559 = ~n2550 & ~n2554 ;
  assign n2560 = ~n2558 & n2559 ;
  assign n2561 = ~n2427 & n2493 ;
  assign n2562 = n2496 & n2561 ;
  assign n2563 = \sub1_data_reg_reg[5]/NET0131  & ~n2562 ;
  assign n2564 = ~decrypt_i_pad & ~\sub1_data_reg_reg[37]/NET0131  ;
  assign n2565 = decrypt_i_pad & ~\sub1_data_reg_reg[101]/NET0131  ;
  assign n2566 = ~n2564 & ~n2565 ;
  assign n2567 = n2421 & n2566 ;
  assign n2568 = ~n2563 & ~n2567 ;
  assign n2569 = \sub1_data_reg_reg[6]/NET0131  & ~n2562 ;
  assign n2570 = ~decrypt_i_pad & ~\sub1_data_reg_reg[38]/NET0131  ;
  assign n2571 = decrypt_i_pad & ~\sub1_data_reg_reg[102]/NET0131  ;
  assign n2572 = ~n2570 & ~n2571 ;
  assign n2573 = n2421 & n2572 ;
  assign n2574 = ~n2569 & ~n2573 ;
  assign n2580 = n2431 & n2561 ;
  assign n2582 = ~n2456 & n2580 ;
  assign n2581 = ~\sub1_data_reg_reg[69]/NET0131  & ~n2580 ;
  assign n2583 = ~n1256 & ~n2581 ;
  assign n2584 = ~n2582 & n2583 ;
  assign n2575 = \sub1_data_reg_reg[69]/NET0131  & n1267 ;
  assign n2576 = ~decrypt_i_pad & ~\sub1_data_reg_reg[101]/NET0131  ;
  assign n2577 = decrypt_i_pad & ~\sub1_data_reg_reg[37]/NET0131  ;
  assign n2578 = ~n2576 & ~n2577 ;
  assign n2579 = n2421 & n2578 ;
  assign n2585 = ~n2575 & ~n2579 ;
  assign n2586 = ~n2584 & n2585 ;
  assign n2593 = n1114 & n2580 ;
  assign n2592 = ~\sub1_data_reg_reg[70]/NET0131  & ~n2580 ;
  assign n2594 = ~n1256 & ~n2592 ;
  assign n2595 = ~n2593 & n2594 ;
  assign n2587 = \sub1_data_reg_reg[70]/NET0131  & n1267 ;
  assign n2588 = ~decrypt_i_pad & ~\sub1_data_reg_reg[102]/NET0131  ;
  assign n2589 = decrypt_i_pad & ~\sub1_data_reg_reg[38]/NET0131  ;
  assign n2590 = ~n2588 & ~n2589 ;
  assign n2591 = n2421 & n2590 ;
  assign n2596 = ~n2587 & ~n2591 ;
  assign n2597 = ~n2595 & n2596 ;
  assign n2603 = n2431 & n2494 ;
  assign n2605 = ~n2456 & n2603 ;
  assign n2604 = ~\sub1_data_reg_reg[85]/NET0131  & ~n2603 ;
  assign n2606 = ~n1256 & ~n2604 ;
  assign n2607 = ~n2605 & n2606 ;
  assign n2598 = \sub1_data_reg_reg[85]/NET0131  & n1267 ;
  assign n2599 = ~decrypt_i_pad & ~\sub1_data_reg_reg[53]/NET0131  ;
  assign n2600 = decrypt_i_pad & ~\sub1_data_reg_reg[117]/NET0131  ;
  assign n2601 = ~n2599 & ~n2600 ;
  assign n2602 = n2421 & n2601 ;
  assign n2608 = ~n2598 & ~n2602 ;
  assign n2609 = ~n2607 & n2608 ;
  assign n2616 = n1114 & n2603 ;
  assign n2615 = ~\sub1_data_reg_reg[86]/NET0131  & ~n2603 ;
  assign n2617 = ~n1256 & ~n2615 ;
  assign n2618 = ~n2616 & n2617 ;
  assign n2610 = \sub1_data_reg_reg[86]/NET0131  & n1267 ;
  assign n2611 = ~decrypt_i_pad & ~\sub1_data_reg_reg[54]/NET0131  ;
  assign n2612 = decrypt_i_pad & ~\sub1_data_reg_reg[118]/NET0131  ;
  assign n2613 = ~n2611 & ~n2612 ;
  assign n2614 = n2421 & n2613 ;
  assign n2619 = ~n2610 & ~n2614 ;
  assign n2620 = ~n2618 & n2619 ;
  assign n2623 = \sub1_state_reg[0]/NET0131  & ~\sub1_state_reg[3]/NET0131  ;
  assign n2624 = n2428 & n2623 ;
  assign n2626 = ~n2456 & n2624 ;
  assign n2625 = ~\sub1_data_reg_reg[109]/NET0131  & ~n2624 ;
  assign n2627 = ~n1256 & ~n2625 ;
  assign n2628 = ~n2626 & n2627 ;
  assign n2621 = \sub1_data_reg_reg[45]/NET0131  & n2421 ;
  assign n2622 = \sub1_data_reg_reg[109]/NET0131  & n1267 ;
  assign n2629 = ~n2621 & ~n2622 ;
  assign n2630 = ~n2628 & n2629 ;
  assign n2634 = n1114 & n2624 ;
  assign n2633 = ~\sub1_data_reg_reg[110]/NET0131  & ~n2624 ;
  assign n2635 = ~n1256 & ~n2633 ;
  assign n2636 = ~n2634 & n2635 ;
  assign n2631 = \sub1_data_reg_reg[46]/NET0131  & n2421 ;
  assign n2632 = \sub1_data_reg_reg[110]/NET0131  & n1267 ;
  assign n2637 = ~n2631 & ~n2632 ;
  assign n2638 = ~n2636 & n2637 ;
  assign n2641 = \sub1_state_reg[0]/NET0131  & \sub1_state_reg[3]/NET0131  ;
  assign n2642 = n2561 & n2641 ;
  assign n2644 = ~n2456 & n2642 ;
  assign n2643 = ~\sub1_data_reg_reg[13]/NET0131  & ~n2642 ;
  assign n2645 = ~n1256 & ~n2643 ;
  assign n2646 = ~n2644 & n2645 ;
  assign n2639 = \sub1_data_reg_reg[77]/NET0131  & n2421 ;
  assign n2640 = \sub1_data_reg_reg[13]/NET0131  & n1267 ;
  assign n2647 = ~n2639 & ~n2640 ;
  assign n2648 = ~n2646 & n2647 ;
  assign n2652 = n1114 & n2642 ;
  assign n2651 = ~\sub1_data_reg_reg[14]/NET0131  & ~n2642 ;
  assign n2653 = ~n1256 & ~n2651 ;
  assign n2654 = ~n2652 & n2653 ;
  assign n2649 = \sub1_data_reg_reg[78]/NET0131  & n2421 ;
  assign n2650 = \sub1_data_reg_reg[14]/NET0131  & n1267 ;
  assign n2655 = ~n2649 & ~n2650 ;
  assign n2656 = ~n2654 & n2655 ;
  assign n2659 = n2428 & n2641 ;
  assign n2661 = ~n2456 & n2659 ;
  assign n2660 = ~\sub1_data_reg_reg[45]/NET0131  & ~n2659 ;
  assign n2662 = ~n1256 & ~n2660 ;
  assign n2663 = ~n2661 & n2662 ;
  assign n2657 = \sub1_data_reg_reg[109]/NET0131  & n2421 ;
  assign n2658 = \sub1_data_reg_reg[45]/NET0131  & n1267 ;
  assign n2664 = ~n2657 & ~n2658 ;
  assign n2665 = ~n2663 & n2664 ;
  assign n2669 = n1114 & n2659 ;
  assign n2668 = ~\sub1_data_reg_reg[46]/NET0131  & ~n2659 ;
  assign n2670 = ~n1256 & ~n2668 ;
  assign n2671 = ~n2669 & n2670 ;
  assign n2666 = \sub1_data_reg_reg[110]/NET0131  & n2421 ;
  assign n2667 = \sub1_data_reg_reg[46]/NET0131  & n1267 ;
  assign n2672 = ~n2666 & ~n2667 ;
  assign n2673 = ~n2671 & n2672 ;
  assign n2676 = n2561 & n2623 ;
  assign n2678 = ~n2456 & n2676 ;
  assign n2677 = ~\sub1_data_reg_reg[77]/NET0131  & ~n2676 ;
  assign n2679 = ~n1256 & ~n2677 ;
  assign n2680 = ~n2678 & n2679 ;
  assign n2674 = \sub1_data_reg_reg[13]/NET0131  & n2421 ;
  assign n2675 = \sub1_data_reg_reg[77]/NET0131  & n1267 ;
  assign n2681 = ~n2674 & ~n2675 ;
  assign n2682 = ~n2680 & n2681 ;
  assign n2686 = n1114 & n2676 ;
  assign n2685 = ~\sub1_data_reg_reg[78]/NET0131  & ~n2676 ;
  assign n2687 = ~n1256 & ~n2685 ;
  assign n2688 = ~n2686 & n2687 ;
  assign n2683 = \sub1_data_reg_reg[14]/NET0131  & n2421 ;
  assign n2684 = \sub1_data_reg_reg[78]/NET0131  & n1267 ;
  assign n2689 = ~n2683 & ~n2684 ;
  assign n2690 = ~n2688 & n2689 ;
  assign n2691 = ~decrypt_i_pad & \sub1_data_reg_reg[32]/NET0131  ;
  assign n2692 = decrypt_i_pad & \sub1_data_reg_reg[96]/NET0131  ;
  assign n2693 = ~n2691 & ~n2692 ;
  assign n2694 = n2421 & ~n2693 ;
  assign n2695 = \sub1_data_reg_reg[0]/NET0131  & ~n2421 ;
  assign n2696 = ~n2694 & ~n2695 ;
  assign n2697 = ~n1090 & ~n2442 ;
  assign n2698 = n1090 & n2442 ;
  assign n2699 = ~n2697 & ~n2698 ;
  assign n2701 = ~n1109 & ~n2699 ;
  assign n2700 = n1109 & n2699 ;
  assign n2702 = ~n974 & ~n2700 ;
  assign n2703 = ~n2701 & n2702 ;
  assign n2704 = ~n1113 & ~n2703 ;
  assign n2705 = ~n2341 & n2704 ;
  assign n2706 = n2341 & ~n2704 ;
  assign n2707 = ~n2705 & ~n2706 ;
  assign n2708 = n2432 & ~n2707 ;
  assign n2709 = ~n1256 & ~n2708 ;
  assign n2711 = ~n1267 & ~n2709 ;
  assign n2712 = \sub1_data_reg_reg[103]/NET0131  & ~n2711 ;
  assign n2710 = n2432 & n2709 ;
  assign n2713 = ~decrypt_i_pad & ~n2707 ;
  assign n2714 = decrypt_i_pad & ~\sub1_data_reg_reg[71]/NET0131  ;
  assign n2715 = n2421 & ~n2714 ;
  assign n2716 = ~n2713 & n2715 ;
  assign n2717 = ~n2710 & ~n2716 ;
  assign n2718 = ~n2712 & n2717 ;
  assign n2725 = ~n2348 & n2468 ;
  assign n2724 = ~\sub1_data_reg_reg[112]/NET0131  & ~n2468 ;
  assign n2726 = ~n1256 & ~n2724 ;
  assign n2727 = ~n2725 & n2726 ;
  assign n2719 = \sub1_data_reg_reg[112]/NET0131  & n1267 ;
  assign n2720 = ~decrypt_i_pad & ~\sub1_data_reg_reg[80]/NET0131  ;
  assign n2721 = decrypt_i_pad & ~\sub1_data_reg_reg[16]/NET0131  ;
  assign n2722 = ~n2720 & ~n2721 ;
  assign n2723 = n2421 & n2722 ;
  assign n2728 = ~n2719 & ~n2723 ;
  assign n2729 = ~n2727 & n2728 ;
  assign n2736 = n1075 & n2317 ;
  assign n2737 = ~n1075 & ~n2317 ;
  assign n2738 = ~n2736 & ~n2737 ;
  assign n2739 = n1052 & n2738 ;
  assign n2740 = ~n1052 & ~n2738 ;
  assign n2741 = ~n2739 & ~n2740 ;
  assign n2742 = ~n974 & ~n2741 ;
  assign n2743 = n974 & n2699 ;
  assign n2744 = ~n2742 & ~n2743 ;
  assign n2745 = n2468 & ~n2744 ;
  assign n2735 = ~\sub1_data_reg_reg[115]/NET0131  & ~n2468 ;
  assign n2746 = ~n1256 & ~n2735 ;
  assign n2747 = ~n2745 & n2746 ;
  assign n2730 = \sub1_data_reg_reg[115]/NET0131  & n1267 ;
  assign n2731 = ~decrypt_i_pad & ~\sub1_data_reg_reg[83]/NET0131  ;
  assign n2732 = decrypt_i_pad & ~\sub1_data_reg_reg[19]/NET0131  ;
  assign n2733 = ~n2731 & ~n2732 ;
  assign n2734 = n2421 & n2733 ;
  assign n2748 = ~n2730 & ~n2734 ;
  assign n2749 = ~n2747 & n2748 ;
  assign n2756 = ~n1106 & ~n2394 ;
  assign n2757 = n1106 & n2394 ;
  assign n2758 = ~n2756 & ~n2757 ;
  assign n2759 = n974 & ~n2317 ;
  assign n2760 = ~n974 & n2442 ;
  assign n2761 = ~n2759 & ~n2760 ;
  assign n2762 = n2758 & ~n2761 ;
  assign n2763 = ~n2758 & n2761 ;
  assign n2764 = ~n2762 & ~n2763 ;
  assign n2765 = n2468 & n2764 ;
  assign n2755 = ~\sub1_data_reg_reg[116]/NET0131  & ~n2468 ;
  assign n2766 = ~n1256 & ~n2755 ;
  assign n2767 = ~n2765 & n2766 ;
  assign n2750 = \sub1_data_reg_reg[116]/NET0131  & n1267 ;
  assign n2751 = ~decrypt_i_pad & ~\sub1_data_reg_reg[84]/NET0131  ;
  assign n2752 = decrypt_i_pad & ~\sub1_data_reg_reg[20]/NET0131  ;
  assign n2753 = ~n2751 & ~n2752 ;
  assign n2754 = n2421 & n2753 ;
  assign n2768 = ~n2750 & ~n2754 ;
  assign n2769 = ~n2767 & n2768 ;
  assign n2776 = n2468 & ~n2707 ;
  assign n2775 = ~\sub1_data_reg_reg[119]/NET0131  & ~n2468 ;
  assign n2777 = ~n1256 & ~n2775 ;
  assign n2778 = ~n2776 & n2777 ;
  assign n2770 = \sub1_data_reg_reg[119]/NET0131  & n1267 ;
  assign n2771 = ~decrypt_i_pad & ~\sub1_data_reg_reg[87]/NET0131  ;
  assign n2772 = decrypt_i_pad & ~\sub1_data_reg_reg[23]/NET0131  ;
  assign n2773 = ~n2771 & ~n2772 ;
  assign n2774 = n2421 & n2773 ;
  assign n2779 = ~n2770 & ~n2774 ;
  assign n2780 = ~n2778 & n2779 ;
  assign n2787 = ~n2348 & n2497 ;
  assign n2786 = ~\sub1_data_reg_reg[16]/NET0131  & ~n2497 ;
  assign n2788 = ~n1256 & ~n2786 ;
  assign n2789 = ~n2787 & n2788 ;
  assign n2781 = \sub1_data_reg_reg[16]/NET0131  & n1267 ;
  assign n2782 = ~decrypt_i_pad & ~\sub1_data_reg_reg[112]/NET0131  ;
  assign n2783 = decrypt_i_pad & ~\sub1_data_reg_reg[48]/NET0131  ;
  assign n2784 = ~n2782 & ~n2783 ;
  assign n2785 = n2421 & n2784 ;
  assign n2790 = ~n2781 & ~n2785 ;
  assign n2791 = ~n2789 & n2790 ;
  assign n2798 = n2497 & ~n2744 ;
  assign n2797 = ~\sub1_data_reg_reg[19]/NET0131  & ~n2497 ;
  assign n2799 = ~n1256 & ~n2797 ;
  assign n2800 = ~n2798 & n2799 ;
  assign n2792 = \sub1_data_reg_reg[19]/NET0131  & n1267 ;
  assign n2793 = ~decrypt_i_pad & ~\sub1_data_reg_reg[115]/NET0131  ;
  assign n2794 = decrypt_i_pad & ~\sub1_data_reg_reg[51]/NET0131  ;
  assign n2795 = ~n2793 & ~n2794 ;
  assign n2796 = n2421 & n2795 ;
  assign n2801 = ~n2792 & ~n2796 ;
  assign n2802 = ~n2800 & n2801 ;
  assign n2809 = n2497 & n2764 ;
  assign n2808 = ~\sub1_data_reg_reg[20]/NET0131  & ~n2497 ;
  assign n2810 = ~n1256 & ~n2808 ;
  assign n2811 = ~n2809 & n2810 ;
  assign n2803 = \sub1_data_reg_reg[20]/NET0131  & n1267 ;
  assign n2804 = ~decrypt_i_pad & ~\sub1_data_reg_reg[116]/NET0131  ;
  assign n2805 = decrypt_i_pad & ~\sub1_data_reg_reg[52]/NET0131  ;
  assign n2806 = ~n2804 & ~n2805 ;
  assign n2807 = n2421 & n2806 ;
  assign n2812 = ~n2803 & ~n2807 ;
  assign n2813 = ~n2811 & n2812 ;
  assign n2820 = n2497 & ~n2707 ;
  assign n2819 = ~\sub1_data_reg_reg[23]/NET0131  & ~n2497 ;
  assign n2821 = ~n1256 & ~n2819 ;
  assign n2822 = ~n2820 & n2821 ;
  assign n2814 = \sub1_data_reg_reg[23]/NET0131  & n1267 ;
  assign n2815 = ~decrypt_i_pad & ~\sub1_data_reg_reg[119]/NET0131  ;
  assign n2816 = decrypt_i_pad & ~\sub1_data_reg_reg[55]/NET0131  ;
  assign n2817 = ~n2815 & ~n2816 ;
  assign n2818 = n2421 & n2817 ;
  assign n2823 = ~n2814 & ~n2818 ;
  assign n2824 = ~n2822 & n2823 ;
  assign n2825 = n2515 & n2764 ;
  assign n2826 = ~n1256 & ~n2825 ;
  assign n2828 = ~n1267 & ~n2826 ;
  assign n2829 = \sub1_data_reg_reg[36]/NET0131  & ~n2828 ;
  assign n2827 = n2515 & n2826 ;
  assign n2831 = decrypt_i_pad & n2764 ;
  assign n2830 = ~decrypt_i_pad & ~\sub1_data_reg_reg[68]/NET0131  ;
  assign n2832 = n2421 & ~n2830 ;
  assign n2833 = ~n2831 & n2832 ;
  assign n2834 = ~n2827 & ~n2833 ;
  assign n2835 = ~n2829 & n2834 ;
  assign n2836 = \sub1_data_reg_reg[3]/NET0131  & ~n2562 ;
  assign n2837 = ~decrypt_i_pad & ~\sub1_data_reg_reg[35]/NET0131  ;
  assign n2838 = decrypt_i_pad & ~\sub1_data_reg_reg[99]/NET0131  ;
  assign n2839 = ~n2837 & ~n2838 ;
  assign n2840 = n2421 & n2839 ;
  assign n2841 = ~n2836 & ~n2840 ;
  assign n2848 = ~n2348 & n2543 ;
  assign n2847 = ~\sub1_data_reg_reg[48]/NET0131  & ~n2543 ;
  assign n2849 = ~n1256 & ~n2847 ;
  assign n2850 = ~n2848 & n2849 ;
  assign n2842 = \sub1_data_reg_reg[48]/NET0131  & n1267 ;
  assign n2843 = ~decrypt_i_pad & ~\sub1_data_reg_reg[16]/NET0131  ;
  assign n2844 = decrypt_i_pad & ~\sub1_data_reg_reg[80]/NET0131  ;
  assign n2845 = ~n2843 & ~n2844 ;
  assign n2846 = n2421 & n2845 ;
  assign n2851 = ~n2842 & ~n2846 ;
  assign n2852 = ~n2850 & n2851 ;
  assign n2853 = \sub1_data_reg_reg[4]/NET0131  & ~n2562 ;
  assign n2854 = ~decrypt_i_pad & ~\sub1_data_reg_reg[36]/NET0131  ;
  assign n2855 = decrypt_i_pad & ~\sub1_data_reg_reg[100]/NET0131  ;
  assign n2856 = ~n2854 & ~n2855 ;
  assign n2857 = n2421 & n2856 ;
  assign n2858 = ~n2853 & ~n2857 ;
  assign n2865 = n2543 & ~n2744 ;
  assign n2864 = ~\sub1_data_reg_reg[51]/NET0131  & ~n2543 ;
  assign n2866 = ~n1256 & ~n2864 ;
  assign n2867 = ~n2865 & n2866 ;
  assign n2859 = \sub1_data_reg_reg[51]/NET0131  & n1267 ;
  assign n2860 = ~decrypt_i_pad & ~\sub1_data_reg_reg[19]/NET0131  ;
  assign n2861 = decrypt_i_pad & ~\sub1_data_reg_reg[83]/NET0131  ;
  assign n2862 = ~n2860 & ~n2861 ;
  assign n2863 = n2421 & n2862 ;
  assign n2868 = ~n2859 & ~n2863 ;
  assign n2869 = ~n2867 & n2868 ;
  assign n2876 = n2543 & n2764 ;
  assign n2875 = ~\sub1_data_reg_reg[52]/NET0131  & ~n2543 ;
  assign n2877 = ~n1256 & ~n2875 ;
  assign n2878 = ~n2876 & n2877 ;
  assign n2870 = \sub1_data_reg_reg[52]/NET0131  & n1267 ;
  assign n2871 = ~decrypt_i_pad & ~\sub1_data_reg_reg[20]/NET0131  ;
  assign n2872 = decrypt_i_pad & ~\sub1_data_reg_reg[84]/NET0131  ;
  assign n2873 = ~n2871 & ~n2872 ;
  assign n2874 = n2421 & n2873 ;
  assign n2879 = ~n2870 & ~n2874 ;
  assign n2880 = ~n2878 & n2879 ;
  assign n2887 = n2543 & ~n2707 ;
  assign n2886 = ~\sub1_data_reg_reg[55]/NET0131  & ~n2543 ;
  assign n2888 = ~n1256 & ~n2886 ;
  assign n2889 = ~n2887 & n2888 ;
  assign n2881 = \sub1_data_reg_reg[55]/NET0131  & n1267 ;
  assign n2882 = ~decrypt_i_pad & ~\sub1_data_reg_reg[23]/NET0131  ;
  assign n2883 = decrypt_i_pad & ~\sub1_data_reg_reg[87]/NET0131  ;
  assign n2884 = ~n2882 & ~n2883 ;
  assign n2885 = n2421 & n2884 ;
  assign n2890 = ~n2881 & ~n2885 ;
  assign n2891 = ~n2889 & n2890 ;
  assign n2898 = ~n2348 & n2580 ;
  assign n2897 = ~\sub1_data_reg_reg[64]/NET0131  & ~n2580 ;
  assign n2899 = ~n1256 & ~n2897 ;
  assign n2900 = ~n2898 & n2899 ;
  assign n2892 = \sub1_data_reg_reg[64]/NET0131  & n1267 ;
  assign n2893 = ~decrypt_i_pad & ~\sub1_data_reg_reg[96]/NET0131  ;
  assign n2894 = decrypt_i_pad & ~\sub1_data_reg_reg[32]/NET0131  ;
  assign n2895 = ~n2893 & ~n2894 ;
  assign n2896 = n2421 & n2895 ;
  assign n2901 = ~n2892 & ~n2896 ;
  assign n2902 = ~n2900 & n2901 ;
  assign n2909 = n2580 & ~n2744 ;
  assign n2908 = ~\sub1_data_reg_reg[67]/NET0131  & ~n2580 ;
  assign n2910 = ~n1256 & ~n2908 ;
  assign n2911 = ~n2909 & n2910 ;
  assign n2903 = \sub1_data_reg_reg[67]/NET0131  & n1267 ;
  assign n2904 = ~decrypt_i_pad & ~\sub1_data_reg_reg[99]/NET0131  ;
  assign n2905 = decrypt_i_pad & ~\sub1_data_reg_reg[35]/NET0131  ;
  assign n2906 = ~n2904 & ~n2905 ;
  assign n2907 = n2421 & n2906 ;
  assign n2912 = ~n2903 & ~n2907 ;
  assign n2913 = ~n2911 & n2912 ;
  assign n2920 = n2580 & n2764 ;
  assign n2919 = ~\sub1_data_reg_reg[68]/NET0131  & ~n2580 ;
  assign n2921 = ~n1256 & ~n2919 ;
  assign n2922 = ~n2920 & n2921 ;
  assign n2914 = \sub1_data_reg_reg[68]/NET0131  & n1267 ;
  assign n2915 = ~decrypt_i_pad & ~\sub1_data_reg_reg[100]/NET0131  ;
  assign n2916 = decrypt_i_pad & ~\sub1_data_reg_reg[36]/NET0131  ;
  assign n2917 = ~n2915 & ~n2916 ;
  assign n2918 = n2421 & n2917 ;
  assign n2923 = ~n2914 & ~n2918 ;
  assign n2924 = ~n2922 & n2923 ;
  assign n2931 = n2580 & ~n2707 ;
  assign n2930 = ~\sub1_data_reg_reg[71]/NET0131  & ~n2580 ;
  assign n2932 = ~n1256 & ~n2930 ;
  assign n2933 = ~n2931 & n2932 ;
  assign n2925 = \sub1_data_reg_reg[71]/NET0131  & n1267 ;
  assign n2926 = ~decrypt_i_pad & ~\sub1_data_reg_reg[103]/NET0131  ;
  assign n2927 = decrypt_i_pad & ~\sub1_data_reg_reg[39]/NET0131  ;
  assign n2928 = ~n2926 & ~n2927 ;
  assign n2929 = n2421 & n2928 ;
  assign n2934 = ~n2925 & ~n2929 ;
  assign n2935 = ~n2933 & n2934 ;
  assign n2936 = \sub1_data_reg_reg[7]/NET0131  & ~n2562 ;
  assign n2937 = ~decrypt_i_pad & ~\sub1_data_reg_reg[39]/NET0131  ;
  assign n2938 = decrypt_i_pad & ~\sub1_data_reg_reg[103]/NET0131  ;
  assign n2939 = ~n2937 & ~n2938 ;
  assign n2940 = n2421 & n2939 ;
  assign n2941 = ~n2936 & ~n2940 ;
  assign n2948 = ~n2348 & n2603 ;
  assign n2947 = ~\sub1_data_reg_reg[80]/NET0131  & ~n2603 ;
  assign n2949 = ~n1256 & ~n2947 ;
  assign n2950 = ~n2948 & n2949 ;
  assign n2942 = \sub1_data_reg_reg[80]/NET0131  & n1267 ;
  assign n2943 = ~decrypt_i_pad & ~\sub1_data_reg_reg[48]/NET0131  ;
  assign n2944 = decrypt_i_pad & ~\sub1_data_reg_reg[112]/NET0131  ;
  assign n2945 = ~n2943 & ~n2944 ;
  assign n2946 = n2421 & n2945 ;
  assign n2951 = ~n2942 & ~n2946 ;
  assign n2952 = ~n2950 & n2951 ;
  assign n2959 = n2603 & ~n2744 ;
  assign n2958 = ~\sub1_data_reg_reg[83]/NET0131  & ~n2603 ;
  assign n2960 = ~n1256 & ~n2958 ;
  assign n2961 = ~n2959 & n2960 ;
  assign n2953 = \sub1_data_reg_reg[83]/NET0131  & n1267 ;
  assign n2954 = ~decrypt_i_pad & ~\sub1_data_reg_reg[51]/NET0131  ;
  assign n2955 = decrypt_i_pad & ~\sub1_data_reg_reg[115]/NET0131  ;
  assign n2956 = ~n2954 & ~n2955 ;
  assign n2957 = n2421 & n2956 ;
  assign n2962 = ~n2953 & ~n2957 ;
  assign n2963 = ~n2961 & n2962 ;
  assign n2970 = n2603 & n2764 ;
  assign n2969 = ~\sub1_data_reg_reg[84]/NET0131  & ~n2603 ;
  assign n2971 = ~n1256 & ~n2969 ;
  assign n2972 = ~n2970 & n2971 ;
  assign n2964 = \sub1_data_reg_reg[84]/NET0131  & n1267 ;
  assign n2965 = ~decrypt_i_pad & ~\sub1_data_reg_reg[52]/NET0131  ;
  assign n2966 = decrypt_i_pad & ~\sub1_data_reg_reg[116]/NET0131  ;
  assign n2967 = ~n2965 & ~n2966 ;
  assign n2968 = n2421 & n2967 ;
  assign n2973 = ~n2964 & ~n2968 ;
  assign n2974 = ~n2972 & n2973 ;
  assign n2981 = n2603 & ~n2707 ;
  assign n2980 = ~\sub1_data_reg_reg[87]/NET0131  & ~n2603 ;
  assign n2982 = ~n1256 & ~n2980 ;
  assign n2983 = ~n2981 & n2982 ;
  assign n2975 = \sub1_data_reg_reg[87]/NET0131  & n1267 ;
  assign n2976 = ~decrypt_i_pad & ~\sub1_data_reg_reg[55]/NET0131  ;
  assign n2977 = decrypt_i_pad & ~\sub1_data_reg_reg[119]/NET0131  ;
  assign n2978 = ~n2976 & ~n2977 ;
  assign n2979 = n2421 & n2978 ;
  assign n2984 = ~n2975 & ~n2979 ;
  assign n2985 = ~n2983 & n2984 ;
  assign n2992 = ~n2348 & n2432 ;
  assign n2991 = ~\sub1_data_reg_reg[96]/NET0131  & ~n2432 ;
  assign n2993 = ~n1256 & ~n2991 ;
  assign n2994 = ~n2992 & n2993 ;
  assign n2986 = \sub1_data_reg_reg[96]/NET0131  & n1267 ;
  assign n2987 = ~decrypt_i_pad & ~n2348 ;
  assign n2988 = decrypt_i_pad & ~\sub1_data_reg_reg[64]/NET0131  ;
  assign n2989 = n2421 & ~n2988 ;
  assign n2990 = ~n2987 & n2989 ;
  assign n2995 = ~n2986 & ~n2990 ;
  assign n2996 = ~n2994 & n2995 ;
  assign n3000 = ~n2348 & n2624 ;
  assign n2999 = ~\sub1_data_reg_reg[104]/NET0131  & ~n2624 ;
  assign n3001 = ~n1256 & ~n2999 ;
  assign n3002 = ~n3000 & n3001 ;
  assign n2997 = \sub1_data_reg_reg[40]/NET0131  & n2421 ;
  assign n2998 = \sub1_data_reg_reg[104]/NET0131  & n1267 ;
  assign n3003 = ~n2997 & ~n2998 ;
  assign n3004 = ~n3002 & n3003 ;
  assign n3008 = n2624 & ~n2744 ;
  assign n3007 = ~\sub1_data_reg_reg[107]/NET0131  & ~n2624 ;
  assign n3009 = ~n1256 & ~n3007 ;
  assign n3010 = ~n3008 & n3009 ;
  assign n3005 = \sub1_data_reg_reg[43]/NET0131  & n2421 ;
  assign n3006 = \sub1_data_reg_reg[107]/NET0131  & n1267 ;
  assign n3011 = ~n3005 & ~n3006 ;
  assign n3012 = ~n3010 & n3011 ;
  assign n3016 = n2624 & n2764 ;
  assign n3015 = ~\sub1_data_reg_reg[108]/NET0131  & ~n2624 ;
  assign n3017 = ~n1256 & ~n3015 ;
  assign n3018 = ~n3016 & n3017 ;
  assign n3013 = \sub1_data_reg_reg[44]/NET0131  & n2421 ;
  assign n3014 = \sub1_data_reg_reg[108]/NET0131  & n1267 ;
  assign n3019 = ~n3013 & ~n3014 ;
  assign n3020 = ~n3018 & n3019 ;
  assign n3024 = n2624 & ~n2707 ;
  assign n3023 = ~\sub1_data_reg_reg[111]/NET0131  & ~n2624 ;
  assign n3025 = ~n1256 & ~n3023 ;
  assign n3026 = ~n3024 & n3025 ;
  assign n3021 = \sub1_data_reg_reg[47]/NET0131  & n2421 ;
  assign n3022 = \sub1_data_reg_reg[111]/NET0131  & n1267 ;
  assign n3027 = ~n3021 & ~n3022 ;
  assign n3028 = ~n3026 & n3027 ;
  assign n3032 = n2642 & ~n2744 ;
  assign n3031 = ~\sub1_data_reg_reg[11]/NET0131  & ~n2642 ;
  assign n3033 = ~n1256 & ~n3031 ;
  assign n3034 = ~n3032 & n3033 ;
  assign n3029 = \sub1_data_reg_reg[75]/NET0131  & n2421 ;
  assign n3030 = \sub1_data_reg_reg[11]/NET0131  & n1267 ;
  assign n3035 = ~n3029 & ~n3030 ;
  assign n3036 = ~n3034 & n3035 ;
  assign n3037 = ~n1114 & n1274 ;
  assign n3038 = \ks1_col_reg[30]/NET0131  & ~n1274 ;
  assign n3039 = ~n3037 & ~n3038 ;
  assign n3040 = \ks1_col_reg[21]/NET0131  & ~n1142 ;
  assign n3041 = n1142 & n2456 ;
  assign n3042 = ~n3040 & ~n3041 ;
  assign n3046 = n2642 & n2764 ;
  assign n3045 = ~\sub1_data_reg_reg[12]/NET0131  & ~n2642 ;
  assign n3047 = ~n1256 & ~n3045 ;
  assign n3048 = ~n3046 & n3047 ;
  assign n3043 = \sub1_data_reg_reg[76]/NET0131  & n2421 ;
  assign n3044 = \sub1_data_reg_reg[12]/NET0131  & n1267 ;
  assign n3049 = ~n3043 & ~n3044 ;
  assign n3050 = ~n3048 & n3049 ;
  assign n3051 = ~n1114 & n1142 ;
  assign n3052 = \ks1_col_reg[22]/NET0131  & ~n1142 ;
  assign n3053 = ~n3051 & ~n3052 ;
  assign n3057 = n2642 & ~n2707 ;
  assign n3056 = ~\sub1_data_reg_reg[15]/NET0131  & ~n2642 ;
  assign n3058 = ~n1256 & ~n3056 ;
  assign n3059 = ~n3057 & n3058 ;
  assign n3054 = \sub1_data_reg_reg[79]/NET0131  & n2421 ;
  assign n3055 = \sub1_data_reg_reg[15]/NET0131  & n1267 ;
  assign n3060 = ~n3054 & ~n3055 ;
  assign n3061 = ~n3059 & n3060 ;
  assign n3062 = ~n1114 & n1286 ;
  assign n3063 = \ks1_col_reg[6]/NET0131  & ~n1286 ;
  assign n3064 = ~n3062 & ~n3063 ;
  assign n3065 = \ks1_col_reg[29]/NET0131  & ~n1274 ;
  assign n3066 = n1274 & n2456 ;
  assign n3067 = ~n3065 & ~n3066 ;
  assign n3068 = \ks1_col_reg[5]/NET0131  & ~n1286 ;
  assign n3069 = n1286 & n2456 ;
  assign n3070 = ~n3068 & ~n3069 ;
  assign n3074 = ~n2348 & n2659 ;
  assign n3073 = ~\sub1_data_reg_reg[40]/NET0131  & ~n2659 ;
  assign n3075 = ~n1256 & ~n3073 ;
  assign n3076 = ~n3074 & n3075 ;
  assign n3071 = \sub1_data_reg_reg[104]/NET0131  & n2421 ;
  assign n3072 = \sub1_data_reg_reg[40]/NET0131  & n1267 ;
  assign n3077 = ~n3071 & ~n3072 ;
  assign n3078 = ~n3076 & n3077 ;
  assign n3082 = n2659 & ~n2744 ;
  assign n3081 = ~\sub1_data_reg_reg[43]/NET0131  & ~n2659 ;
  assign n3083 = ~n1256 & ~n3081 ;
  assign n3084 = ~n3082 & n3083 ;
  assign n3079 = \sub1_data_reg_reg[107]/NET0131  & n2421 ;
  assign n3080 = \sub1_data_reg_reg[43]/NET0131  & n1267 ;
  assign n3085 = ~n3079 & ~n3080 ;
  assign n3086 = ~n3084 & n3085 ;
  assign n3090 = n2659 & n2764 ;
  assign n3089 = ~\sub1_data_reg_reg[44]/NET0131  & ~n2659 ;
  assign n3091 = ~n1256 & ~n3089 ;
  assign n3092 = ~n3090 & n3091 ;
  assign n3087 = \sub1_data_reg_reg[108]/NET0131  & n2421 ;
  assign n3088 = \sub1_data_reg_reg[44]/NET0131  & n1267 ;
  assign n3093 = ~n3087 & ~n3088 ;
  assign n3094 = ~n3092 & n3093 ;
  assign n3098 = n2659 & ~n2707 ;
  assign n3097 = ~\sub1_data_reg_reg[47]/NET0131  & ~n2659 ;
  assign n3099 = ~n1256 & ~n3097 ;
  assign n3100 = ~n3098 & n3099 ;
  assign n3095 = \sub1_data_reg_reg[111]/NET0131  & n2421 ;
  assign n3096 = \sub1_data_reg_reg[47]/NET0131  & n1267 ;
  assign n3101 = ~n3095 & ~n3096 ;
  assign n3102 = ~n3100 & n3101 ;
  assign n3106 = ~n2348 & n2676 ;
  assign n3105 = ~\sub1_data_reg_reg[72]/NET0131  & ~n2676 ;
  assign n3107 = ~n1256 & ~n3105 ;
  assign n3108 = ~n3106 & n3107 ;
  assign n3103 = \sub1_data_reg_reg[8]/NET0131  & n2421 ;
  assign n3104 = \sub1_data_reg_reg[72]/NET0131  & n1267 ;
  assign n3109 = ~n3103 & ~n3104 ;
  assign n3110 = ~n3108 & n3109 ;
  assign n3114 = n2676 & ~n2744 ;
  assign n3113 = ~\sub1_data_reg_reg[75]/NET0131  & ~n2676 ;
  assign n3115 = ~n1256 & ~n3113 ;
  assign n3116 = ~n3114 & n3115 ;
  assign n3111 = \sub1_data_reg_reg[11]/NET0131  & n2421 ;
  assign n3112 = \sub1_data_reg_reg[75]/NET0131  & n1267 ;
  assign n3117 = ~n3111 & ~n3112 ;
  assign n3118 = ~n3116 & n3117 ;
  assign n3122 = n2676 & n2764 ;
  assign n3121 = ~\sub1_data_reg_reg[76]/NET0131  & ~n2676 ;
  assign n3123 = ~n1256 & ~n3121 ;
  assign n3124 = ~n3122 & n3123 ;
  assign n3119 = \sub1_data_reg_reg[12]/NET0131  & n2421 ;
  assign n3120 = \sub1_data_reg_reg[76]/NET0131  & n1267 ;
  assign n3125 = ~n3119 & ~n3120 ;
  assign n3126 = ~n3124 & n3125 ;
  assign n3130 = n2676 & ~n2707 ;
  assign n3129 = ~\sub1_data_reg_reg[79]/NET0131  & ~n2676 ;
  assign n3131 = ~n1256 & ~n3129 ;
  assign n3132 = ~n3130 & n3131 ;
  assign n3127 = \sub1_data_reg_reg[15]/NET0131  & n2421 ;
  assign n3128 = \sub1_data_reg_reg[79]/NET0131  & n1267 ;
  assign n3133 = ~n3127 & ~n3128 ;
  assign n3134 = ~n3132 & n3133 ;
  assign n3138 = ~n2348 & n2642 ;
  assign n3137 = ~\sub1_data_reg_reg[8]/NET0131  & ~n2642 ;
  assign n3139 = ~n1256 & ~n3137 ;
  assign n3140 = ~n3138 & n3139 ;
  assign n3135 = \sub1_data_reg_reg[72]/NET0131  & n2421 ;
  assign n3136 = \sub1_data_reg_reg[8]/NET0131  & n1267 ;
  assign n3141 = ~n3135 & ~n3136 ;
  assign n3142 = ~n3140 & n3141 ;
  assign n3143 = ~n2348 & n2515 ;
  assign n3144 = ~n1256 & ~n3143 ;
  assign n3146 = ~n1267 & ~n3144 ;
  assign n3147 = \sub1_data_reg_reg[32]/NET0131  & ~n3146 ;
  assign n3145 = n2515 & n3144 ;
  assign n3149 = decrypt_i_pad & ~n2348 ;
  assign n3148 = ~decrypt_i_pad & ~\sub1_data_reg_reg[64]/NET0131  ;
  assign n3150 = n2421 & ~n3148 ;
  assign n3151 = ~n3149 & n3150 ;
  assign n3152 = ~n3145 & ~n3151 ;
  assign n3153 = ~n3147 & n3152 ;
  assign n3154 = n2515 & ~n2744 ;
  assign n3155 = ~n1256 & ~n3154 ;
  assign n3157 = ~n1267 & ~n3155 ;
  assign n3158 = \sub1_data_reg_reg[35]/NET0131  & ~n3157 ;
  assign n3156 = n2515 & n3155 ;
  assign n3160 = decrypt_i_pad & ~n2744 ;
  assign n3159 = ~decrypt_i_pad & ~\sub1_data_reg_reg[67]/NET0131  ;
  assign n3161 = n2421 & ~n3159 ;
  assign n3162 = ~n3160 & n3161 ;
  assign n3163 = ~n3156 & ~n3162 ;
  assign n3164 = ~n3158 & n3163 ;
  assign n3165 = n2515 & ~n2707 ;
  assign n3166 = ~n1256 & ~n3165 ;
  assign n3168 = ~n1267 & ~n3166 ;
  assign n3169 = \sub1_data_reg_reg[39]/NET0131  & ~n3168 ;
  assign n3167 = n2515 & n3166 ;
  assign n3171 = decrypt_i_pad & ~n2707 ;
  assign n3170 = ~decrypt_i_pad & ~\sub1_data_reg_reg[71]/NET0131  ;
  assign n3172 = n2421 & ~n3170 ;
  assign n3173 = ~n3171 & n3172 ;
  assign n3174 = ~n3167 & ~n3173 ;
  assign n3175 = ~n3169 & n3174 ;
  assign n3176 = n2432 & n2764 ;
  assign n3177 = ~n1256 & ~n3176 ;
  assign n3179 = ~n1267 & ~n3177 ;
  assign n3180 = \sub1_data_reg_reg[100]/NET0131  & ~n3179 ;
  assign n3178 = n2432 & n3177 ;
  assign n3181 = ~decrypt_i_pad & n2764 ;
  assign n3182 = decrypt_i_pad & ~\sub1_data_reg_reg[68]/NET0131  ;
  assign n3183 = n2421 & ~n3182 ;
  assign n3184 = ~n3181 & n3183 ;
  assign n3185 = ~n3178 & ~n3184 ;
  assign n3186 = ~n3180 & n3185 ;
  assign n3187 = n2432 & ~n2744 ;
  assign n3188 = ~n1256 & ~n3187 ;
  assign n3190 = ~n1267 & ~n3188 ;
  assign n3191 = \sub1_data_reg_reg[99]/NET0131  & ~n3190 ;
  assign n3189 = n2432 & n3188 ;
  assign n3192 = ~decrypt_i_pad & ~n2741 ;
  assign n3193 = decrypt_i_pad & ~\sub1_data_reg_reg[67]/NET0131  ;
  assign n3194 = n2421 & ~n3193 ;
  assign n3195 = ~n3192 & n3194 ;
  assign n3196 = ~n3189 & ~n3195 ;
  assign n3197 = ~n3191 & n3196 ;
  assign n3198 = n2467 & n2623 ;
  assign n3199 = \sub1_data_reg_reg[125]/NET0131  & ~n3198 ;
  assign n3200 = n2456 & n3198 ;
  assign n3201 = ~n3199 & ~n3200 ;
  assign n3202 = ~n1114 & n3198 ;
  assign n3203 = \sub1_data_reg_reg[126]/NET0131  & ~n3198 ;
  assign n3204 = ~n3202 & ~n3203 ;
  assign n3205 = n2494 & n2641 ;
  assign n3206 = \sub1_data_reg_reg[29]/NET0131  & ~n3205 ;
  assign n3207 = n2456 & n3205 ;
  assign n3208 = ~n3206 & ~n3207 ;
  assign n3209 = ~n1114 & n3205 ;
  assign n3210 = \sub1_data_reg_reg[30]/NET0131  & ~n3205 ;
  assign n3211 = ~n3209 & ~n3210 ;
  assign n3212 = n2467 & n2641 ;
  assign n3213 = \sub1_data_reg_reg[61]/NET0131  & ~n3212 ;
  assign n3214 = n2456 & n3212 ;
  assign n3215 = ~n3213 & ~n3214 ;
  assign n3216 = ~n1114 & n3212 ;
  assign n3217 = \sub1_data_reg_reg[62]/NET0131  & ~n3212 ;
  assign n3218 = ~n3216 & ~n3217 ;
  assign n3219 = n2494 & n2623 ;
  assign n3220 = \sub1_data_reg_reg[93]/NET0131  & ~n3219 ;
  assign n3221 = n2456 & n3219 ;
  assign n3222 = ~n3220 & ~n3221 ;
  assign n3223 = ~n1114 & n3219 ;
  assign n3224 = \sub1_data_reg_reg[94]/NET0131  & ~n3219 ;
  assign n3225 = ~n3223 & ~n3224 ;
  assign n3226 = \ks1_key_reg_reg[73]/NET0131  & ~n929 ;
  assign n3227 = \key_i[73]_pad  & ~n1116 ;
  assign n3228 = \ks1_key_reg_reg[73]/NET0131  & n1116 ;
  assign n3229 = ~n3227 & ~n3228 ;
  assign n3230 = n974 & ~n2391 ;
  assign n3231 = ~n2341 & n2738 ;
  assign n3232 = n2341 & ~n2738 ;
  assign n3233 = ~n3231 & ~n3232 ;
  assign n3234 = ~n974 & n3233 ;
  assign n3235 = ~n3230 & ~n3234 ;
  assign n3236 = ~\ks1_key_reg_reg[105]/NET0131  & n1116 ;
  assign n3237 = ~\key_i[105]_pad  & ~n1116 ;
  assign n3238 = ~n3236 & ~n3237 ;
  assign n3239 = n3235 & ~n3238 ;
  assign n3240 = ~n3235 & n3238 ;
  assign n3241 = ~n3239 & ~n3240 ;
  assign n3242 = n3229 & n3241 ;
  assign n3243 = ~n3229 & ~n3241 ;
  assign n3244 = ~n3242 & ~n3243 ;
  assign n3245 = n929 & ~n3244 ;
  assign n3246 = ~n3226 & ~n3245 ;
  assign n3247 = n929 & n2406 ;
  assign n3248 = \ks1_key_reg_reg[74]/NET0131  & ~n929 ;
  assign n3249 = ~n3247 & ~n3248 ;
  assign n3256 = n2468 & n3235 ;
  assign n3255 = ~\sub1_data_reg_reg[113]/NET0131  & ~n2468 ;
  assign n3257 = ~n1256 & ~n3255 ;
  assign n3258 = ~n3256 & n3257 ;
  assign n3250 = \sub1_data_reg_reg[113]/NET0131  & n1267 ;
  assign n3251 = ~decrypt_i_pad & ~\sub1_data_reg_reg[81]/NET0131  ;
  assign n3252 = decrypt_i_pad & ~\sub1_data_reg_reg[17]/NET0131  ;
  assign n3253 = ~n3251 & ~n3252 ;
  assign n3254 = n2421 & n3253 ;
  assign n3259 = ~n3250 & ~n3254 ;
  assign n3260 = ~n3258 & n3259 ;
  assign n3267 = ~n2400 & n2468 ;
  assign n3266 = ~\sub1_data_reg_reg[114]/NET0131  & ~n2468 ;
  assign n3268 = ~n1256 & ~n3266 ;
  assign n3269 = ~n3267 & n3268 ;
  assign n3261 = \sub1_data_reg_reg[114]/NET0131  & n1267 ;
  assign n3262 = ~decrypt_i_pad & ~\sub1_data_reg_reg[82]/NET0131  ;
  assign n3263 = decrypt_i_pad & ~\sub1_data_reg_reg[18]/NET0131  ;
  assign n3264 = ~n3262 & ~n3263 ;
  assign n3265 = n2421 & n3264 ;
  assign n3270 = ~n3261 & ~n3265 ;
  assign n3271 = ~n3269 & n3270 ;
  assign n3278 = n2497 & n3235 ;
  assign n3277 = ~\sub1_data_reg_reg[17]/NET0131  & ~n2497 ;
  assign n3279 = ~n1256 & ~n3277 ;
  assign n3280 = ~n3278 & n3279 ;
  assign n3272 = \sub1_data_reg_reg[17]/NET0131  & n1267 ;
  assign n3273 = ~decrypt_i_pad & ~\sub1_data_reg_reg[113]/NET0131  ;
  assign n3274 = decrypt_i_pad & ~\sub1_data_reg_reg[49]/NET0131  ;
  assign n3275 = ~n3273 & ~n3274 ;
  assign n3276 = n2421 & n3275 ;
  assign n3281 = ~n3272 & ~n3276 ;
  assign n3282 = ~n3280 & n3281 ;
  assign n3289 = ~n2400 & n2497 ;
  assign n3288 = ~\sub1_data_reg_reg[18]/NET0131  & ~n2497 ;
  assign n3290 = ~n1256 & ~n3288 ;
  assign n3291 = ~n3289 & n3290 ;
  assign n3283 = \sub1_data_reg_reg[18]/NET0131  & n1267 ;
  assign n3284 = ~decrypt_i_pad & ~\sub1_data_reg_reg[114]/NET0131  ;
  assign n3285 = decrypt_i_pad & ~\sub1_data_reg_reg[50]/NET0131  ;
  assign n3286 = ~n3284 & ~n3285 ;
  assign n3287 = n2421 & n3286 ;
  assign n3292 = ~n3283 & ~n3287 ;
  assign n3293 = ~n3291 & n3292 ;
  assign n3294 = ~decrypt_i_pad & \sub1_data_reg_reg[33]/NET0131  ;
  assign n3295 = decrypt_i_pad & \sub1_data_reg_reg[97]/NET0131  ;
  assign n3296 = ~n3294 & ~n3295 ;
  assign n3297 = n2421 & ~n3296 ;
  assign n3298 = \sub1_data_reg_reg[1]/NET0131  & ~n2421 ;
  assign n3299 = ~n3297 & ~n3298 ;
  assign n3300 = \sub1_data_reg_reg[2]/NET0131  & ~n2562 ;
  assign n3301 = ~decrypt_i_pad & ~\sub1_data_reg_reg[34]/NET0131  ;
  assign n3302 = decrypt_i_pad & ~\sub1_data_reg_reg[98]/NET0131  ;
  assign n3303 = ~n3301 & ~n3302 ;
  assign n3304 = n2421 & n3303 ;
  assign n3305 = ~n3300 & ~n3304 ;
  assign n3312 = n2543 & n3235 ;
  assign n3311 = ~\sub1_data_reg_reg[49]/NET0131  & ~n2543 ;
  assign n3313 = ~n1256 & ~n3311 ;
  assign n3314 = ~n3312 & n3313 ;
  assign n3306 = \sub1_data_reg_reg[49]/NET0131  & n1267 ;
  assign n3307 = ~decrypt_i_pad & ~\sub1_data_reg_reg[17]/NET0131  ;
  assign n3308 = decrypt_i_pad & ~\sub1_data_reg_reg[81]/NET0131  ;
  assign n3309 = ~n3307 & ~n3308 ;
  assign n3310 = n2421 & n3309 ;
  assign n3315 = ~n3306 & ~n3310 ;
  assign n3316 = ~n3314 & n3315 ;
  assign n3323 = ~n2400 & n2543 ;
  assign n3322 = ~\sub1_data_reg_reg[50]/NET0131  & ~n2543 ;
  assign n3324 = ~n1256 & ~n3322 ;
  assign n3325 = ~n3323 & n3324 ;
  assign n3317 = \sub1_data_reg_reg[50]/NET0131  & n1267 ;
  assign n3318 = ~decrypt_i_pad & ~\sub1_data_reg_reg[18]/NET0131  ;
  assign n3319 = decrypt_i_pad & ~\sub1_data_reg_reg[82]/NET0131  ;
  assign n3320 = ~n3318 & ~n3319 ;
  assign n3321 = n2421 & n3320 ;
  assign n3326 = ~n3317 & ~n3321 ;
  assign n3327 = ~n3325 & n3326 ;
  assign n3334 = n2580 & n3235 ;
  assign n3333 = ~\sub1_data_reg_reg[65]/NET0131  & ~n2580 ;
  assign n3335 = ~n1256 & ~n3333 ;
  assign n3336 = ~n3334 & n3335 ;
  assign n3328 = \sub1_data_reg_reg[65]/NET0131  & n1267 ;
  assign n3329 = ~decrypt_i_pad & ~\sub1_data_reg_reg[97]/NET0131  ;
  assign n3330 = decrypt_i_pad & ~\sub1_data_reg_reg[33]/NET0131  ;
  assign n3331 = ~n3329 & ~n3330 ;
  assign n3332 = n2421 & n3331 ;
  assign n3337 = ~n3328 & ~n3332 ;
  assign n3338 = ~n3336 & n3337 ;
  assign n3345 = ~n2400 & n2580 ;
  assign n3344 = ~\sub1_data_reg_reg[66]/NET0131  & ~n2580 ;
  assign n3346 = ~n1256 & ~n3344 ;
  assign n3347 = ~n3345 & n3346 ;
  assign n3339 = \sub1_data_reg_reg[66]/NET0131  & n1267 ;
  assign n3340 = ~decrypt_i_pad & ~\sub1_data_reg_reg[98]/NET0131  ;
  assign n3341 = decrypt_i_pad & ~\sub1_data_reg_reg[34]/NET0131  ;
  assign n3342 = ~n3340 & ~n3341 ;
  assign n3343 = n2421 & n3342 ;
  assign n3348 = ~n3339 & ~n3343 ;
  assign n3349 = ~n3347 & n3348 ;
  assign n3356 = n2603 & n3235 ;
  assign n3355 = ~\sub1_data_reg_reg[81]/NET0131  & ~n2603 ;
  assign n3357 = ~n1256 & ~n3355 ;
  assign n3358 = ~n3356 & n3357 ;
  assign n3350 = \sub1_data_reg_reg[81]/NET0131  & n1267 ;
  assign n3351 = ~decrypt_i_pad & ~\sub1_data_reg_reg[49]/NET0131  ;
  assign n3352 = decrypt_i_pad & ~\sub1_data_reg_reg[113]/NET0131  ;
  assign n3353 = ~n3351 & ~n3352 ;
  assign n3354 = n2421 & n3353 ;
  assign n3359 = ~n3350 & ~n3354 ;
  assign n3360 = ~n3358 & n3359 ;
  assign n3367 = ~n2400 & n2603 ;
  assign n3366 = ~\sub1_data_reg_reg[82]/NET0131  & ~n2603 ;
  assign n3368 = ~n1256 & ~n3366 ;
  assign n3369 = ~n3367 & n3368 ;
  assign n3361 = \sub1_data_reg_reg[82]/NET0131  & n1267 ;
  assign n3362 = ~decrypt_i_pad & ~\sub1_data_reg_reg[50]/NET0131  ;
  assign n3363 = decrypt_i_pad & ~\sub1_data_reg_reg[114]/NET0131  ;
  assign n3364 = ~n3362 & ~n3363 ;
  assign n3365 = n2421 & n3364 ;
  assign n3370 = ~n3361 & ~n3365 ;
  assign n3371 = ~n3369 & n3370 ;
  assign n3378 = n2432 & n3235 ;
  assign n3377 = ~\sub1_data_reg_reg[97]/NET0131  & ~n2432 ;
  assign n3379 = ~n1256 & ~n3377 ;
  assign n3380 = ~n3378 & n3379 ;
  assign n3372 = \sub1_data_reg_reg[97]/NET0131  & n1267 ;
  assign n3373 = ~decrypt_i_pad & ~n3233 ;
  assign n3374 = decrypt_i_pad & ~\sub1_data_reg_reg[65]/NET0131  ;
  assign n3375 = n2421 & ~n3374 ;
  assign n3376 = ~n3373 & n3375 ;
  assign n3381 = ~n3372 & ~n3376 ;
  assign n3382 = ~n3380 & n3381 ;
  assign n3383 = ~n2400 & n2432 ;
  assign n3384 = ~n1256 & ~n3383 ;
  assign n3386 = ~n1267 & ~n3384 ;
  assign n3387 = \sub1_data_reg_reg[98]/NET0131  & ~n3386 ;
  assign n3385 = n2432 & n3384 ;
  assign n3388 = ~decrypt_i_pad & ~n2400 ;
  assign n3389 = decrypt_i_pad & ~\sub1_data_reg_reg[66]/NET0131  ;
  assign n3390 = n2421 & ~n3389 ;
  assign n3391 = ~n3388 & n3390 ;
  assign n3392 = ~n3385 & ~n3391 ;
  assign n3393 = ~n3387 & n3392 ;
  assign n3397 = n2624 & n3235 ;
  assign n3396 = ~\sub1_data_reg_reg[105]/NET0131  & ~n2624 ;
  assign n3398 = ~n1256 & ~n3396 ;
  assign n3399 = ~n3397 & n3398 ;
  assign n3394 = \sub1_data_reg_reg[41]/NET0131  & n2421 ;
  assign n3395 = \sub1_data_reg_reg[105]/NET0131  & n1267 ;
  assign n3400 = ~n3394 & ~n3395 ;
  assign n3401 = ~n3399 & n3400 ;
  assign n3405 = ~n2400 & n2624 ;
  assign n3404 = ~\sub1_data_reg_reg[106]/NET0131  & ~n2624 ;
  assign n3406 = ~n1256 & ~n3404 ;
  assign n3407 = ~n3405 & n3406 ;
  assign n3402 = \sub1_data_reg_reg[42]/NET0131  & n2421 ;
  assign n3403 = \sub1_data_reg_reg[106]/NET0131  & n1267 ;
  assign n3408 = ~n3402 & ~n3403 ;
  assign n3409 = ~n3407 & n3408 ;
  assign n3410 = n1286 & ~n2348 ;
  assign n3411 = ~\ks1_col_reg[0]/NET0131  & ~n1286 ;
  assign n3412 = ~n3410 & ~n3411 ;
  assign n3413 = n1142 & ~n2744 ;
  assign n3414 = ~\ks1_col_reg[19]/NET0131  & ~n1142 ;
  assign n3415 = ~n3413 & ~n3414 ;
  assign n3416 = n1142 & ~n2348 ;
  assign n3417 = ~\ks1_col_reg[16]/NET0131  & ~n1142 ;
  assign n3418 = ~n3416 & ~n3417 ;
  assign n3419 = \ks1_col_reg[20]/NET0131  & ~n1142 ;
  assign n3420 = n1142 & ~n2764 ;
  assign n3421 = ~n3419 & ~n3420 ;
  assign n3425 = ~n2400 & n2642 ;
  assign n3424 = ~\sub1_data_reg_reg[10]/NET0131  & ~n2642 ;
  assign n3426 = ~n1256 & ~n3424 ;
  assign n3427 = ~n3425 & n3426 ;
  assign n3422 = \sub1_data_reg_reg[74]/NET0131  & n2421 ;
  assign n3423 = \sub1_data_reg_reg[10]/NET0131  & n1267 ;
  assign n3428 = ~n3422 & ~n3423 ;
  assign n3429 = ~n3427 & n3428 ;
  assign n3430 = n1142 & n2707 ;
  assign n3431 = \ks1_col_reg[23]/NET0131  & ~n1142 ;
  assign n3432 = ~n3430 & ~n3431 ;
  assign n3433 = n1274 & ~n2348 ;
  assign n3434 = ~\ks1_col_reg[24]/NET0131  & ~n1274 ;
  assign n3435 = ~n3433 & ~n3434 ;
  assign n3436 = n1274 & ~n2744 ;
  assign n3437 = ~\ks1_col_reg[27]/NET0131  & ~n1274 ;
  assign n3438 = ~n3436 & ~n3437 ;
  assign n3439 = \ks1_col_reg[28]/NET0131  & ~n1274 ;
  assign n3440 = n1274 & ~n2764 ;
  assign n3441 = ~n3439 & ~n3440 ;
  assign n3442 = n1274 & n2707 ;
  assign n3443 = \ks1_col_reg[31]/NET0131  & ~n1274 ;
  assign n3444 = ~n3442 & ~n3443 ;
  assign n3445 = n1286 & ~n2744 ;
  assign n3446 = ~\ks1_col_reg[3]/NET0131  & ~n1286 ;
  assign n3447 = ~n3445 & ~n3446 ;
  assign n3448 = \ks1_col_reg[4]/NET0131  & ~n1286 ;
  assign n3449 = n1286 & ~n2764 ;
  assign n3450 = ~n3448 & ~n3449 ;
  assign n3451 = n1286 & n2707 ;
  assign n3452 = \ks1_col_reg[7]/NET0131  & ~n1286 ;
  assign n3453 = ~n3451 & ~n3452 ;
  assign n3457 = n2659 & n3235 ;
  assign n3456 = ~\sub1_data_reg_reg[41]/NET0131  & ~n2659 ;
  assign n3458 = ~n1256 & ~n3456 ;
  assign n3459 = ~n3457 & n3458 ;
  assign n3454 = \sub1_data_reg_reg[105]/NET0131  & n2421 ;
  assign n3455 = \sub1_data_reg_reg[41]/NET0131  & n1267 ;
  assign n3460 = ~n3454 & ~n3455 ;
  assign n3461 = ~n3459 & n3460 ;
  assign n3465 = ~n2400 & n2659 ;
  assign n3464 = ~\sub1_data_reg_reg[42]/NET0131  & ~n2659 ;
  assign n3466 = ~n1256 & ~n3464 ;
  assign n3467 = ~n3465 & n3466 ;
  assign n3462 = \sub1_data_reg_reg[106]/NET0131  & n2421 ;
  assign n3463 = \sub1_data_reg_reg[42]/NET0131  & n1267 ;
  assign n3468 = ~n3462 & ~n3463 ;
  assign n3469 = ~n3467 & n3468 ;
  assign n3473 = n2676 & n3235 ;
  assign n3472 = ~\sub1_data_reg_reg[73]/NET0131  & ~n2676 ;
  assign n3474 = ~n1256 & ~n3472 ;
  assign n3475 = ~n3473 & n3474 ;
  assign n3470 = \sub1_data_reg_reg[9]/NET0131  & n2421 ;
  assign n3471 = \sub1_data_reg_reg[73]/NET0131  & n1267 ;
  assign n3476 = ~n3470 & ~n3471 ;
  assign n3477 = ~n3475 & n3476 ;
  assign n3481 = ~n2400 & n2676 ;
  assign n3480 = ~\sub1_data_reg_reg[74]/NET0131  & ~n2676 ;
  assign n3482 = ~n1256 & ~n3480 ;
  assign n3483 = ~n3481 & n3482 ;
  assign n3478 = \sub1_data_reg_reg[10]/NET0131  & n2421 ;
  assign n3479 = \sub1_data_reg_reg[74]/NET0131  & n1267 ;
  assign n3484 = ~n3478 & ~n3479 ;
  assign n3485 = ~n3483 & n3484 ;
  assign n3489 = n2642 & n3235 ;
  assign n3488 = ~\sub1_data_reg_reg[9]/NET0131  & ~n2642 ;
  assign n3490 = ~n1256 & ~n3488 ;
  assign n3491 = ~n3489 & n3490 ;
  assign n3486 = \sub1_data_reg_reg[73]/NET0131  & n2421 ;
  assign n3487 = \sub1_data_reg_reg[9]/NET0131  & n1267 ;
  assign n3492 = ~n3486 & ~n3487 ;
  assign n3493 = ~n3491 & n3492 ;
  assign n3494 = n2515 & n3235 ;
  assign n3495 = ~n1256 & ~n3494 ;
  assign n3497 = ~n1267 & ~n3495 ;
  assign n3498 = \sub1_data_reg_reg[33]/NET0131  & ~n3497 ;
  assign n3496 = n2515 & n3495 ;
  assign n3500 = decrypt_i_pad & n3235 ;
  assign n3499 = ~decrypt_i_pad & ~\sub1_data_reg_reg[65]/NET0131  ;
  assign n3501 = n2421 & ~n3499 ;
  assign n3502 = ~n3500 & n3501 ;
  assign n3503 = ~n3496 & ~n3502 ;
  assign n3504 = ~n3498 & n3503 ;
  assign n3505 = ~n2400 & n2515 ;
  assign n3506 = ~n1256 & ~n3505 ;
  assign n3508 = ~n1267 & ~n3506 ;
  assign n3509 = \sub1_data_reg_reg[34]/NET0131  & ~n3508 ;
  assign n3507 = n2515 & n3506 ;
  assign n3511 = decrypt_i_pad & ~n2400 ;
  assign n3510 = ~decrypt_i_pad & ~\sub1_data_reg_reg[66]/NET0131  ;
  assign n3512 = n2421 & ~n3510 ;
  assign n3513 = ~n3511 & n3512 ;
  assign n3514 = ~n3507 & ~n3513 ;
  assign n3515 = ~n3509 & n3514 ;
  assign n3516 = ~n2348 & n3198 ;
  assign n3517 = ~\sub1_data_reg_reg[120]/NET0131  & ~n3198 ;
  assign n3518 = ~n3516 & ~n3517 ;
  assign n3519 = ~n2348 & n3205 ;
  assign n3520 = ~\sub1_data_reg_reg[24]/NET0131  & ~n3205 ;
  assign n3521 = ~n3519 & ~n3520 ;
  assign n3522 = ~n2348 & n3212 ;
  assign n3523 = ~\sub1_data_reg_reg[56]/NET0131  & ~n3212 ;
  assign n3524 = ~n3522 & ~n3523 ;
  assign n3525 = ~n2348 & n3219 ;
  assign n3526 = ~\sub1_data_reg_reg[88]/NET0131  & ~n3219 ;
  assign n3527 = ~n3525 & ~n3526 ;
  assign n3528 = ~n2744 & n3198 ;
  assign n3529 = ~\sub1_data_reg_reg[123]/NET0131  & ~n3198 ;
  assign n3530 = ~n3528 & ~n3529 ;
  assign n3531 = \sub1_data_reg_reg[124]/NET0131  & ~n3198 ;
  assign n3532 = ~n2764 & n3198 ;
  assign n3533 = ~n3531 & ~n3532 ;
  assign n3534 = n2707 & n3198 ;
  assign n3535 = \sub1_data_reg_reg[127]/NET0131  & ~n3198 ;
  assign n3536 = ~n3534 & ~n3535 ;
  assign n3537 = ~n2744 & n3205 ;
  assign n3538 = ~\sub1_data_reg_reg[27]/NET0131  & ~n3205 ;
  assign n3539 = ~n3537 & ~n3538 ;
  assign n3540 = \sub1_data_reg_reg[28]/NET0131  & ~n3205 ;
  assign n3541 = ~n2764 & n3205 ;
  assign n3542 = ~n3540 & ~n3541 ;
  assign n3543 = n2707 & n3205 ;
  assign n3544 = \sub1_data_reg_reg[31]/NET0131  & ~n3205 ;
  assign n3545 = ~n3543 & ~n3544 ;
  assign n3546 = ~n2744 & n3212 ;
  assign n3547 = ~\sub1_data_reg_reg[59]/NET0131  & ~n3212 ;
  assign n3548 = ~n3546 & ~n3547 ;
  assign n3549 = \sub1_data_reg_reg[60]/NET0131  & ~n3212 ;
  assign n3550 = ~n2764 & n3212 ;
  assign n3551 = ~n3549 & ~n3550 ;
  assign n3552 = n2707 & n3212 ;
  assign n3553 = \sub1_data_reg_reg[63]/NET0131  & ~n3212 ;
  assign n3554 = ~n3552 & ~n3553 ;
  assign n3555 = ~n2744 & n3219 ;
  assign n3556 = ~\sub1_data_reg_reg[91]/NET0131  & ~n3219 ;
  assign n3557 = ~n3555 & ~n3556 ;
  assign n3558 = \sub1_data_reg_reg[92]/NET0131  & ~n3219 ;
  assign n3559 = ~n2764 & n3219 ;
  assign n3560 = ~n3558 & ~n3559 ;
  assign n3561 = n2707 & n3219 ;
  assign n3562 = \sub1_data_reg_reg[95]/NET0131  & ~n3219 ;
  assign n3563 = ~n3561 & ~n3562 ;
  assign n3564 = ~\ks1_key_reg_reg[111]/NET0131  & n1116 ;
  assign n3565 = ~\key_i[111]_pad  & ~n1116 ;
  assign n3566 = ~n3564 & ~n3565 ;
  assign n3567 = n2707 & ~n3566 ;
  assign n3568 = ~n2707 & n3566 ;
  assign n3569 = ~n3567 & ~n3568 ;
  assign n3570 = ~n2233 & n2257 ;
  assign n3571 = n2233 & ~n2257 ;
  assign n3572 = ~n3570 & ~n3571 ;
  assign n3573 = n1142 & n2400 ;
  assign n3574 = \ks1_col_reg[18]/NET0131  & ~n1142 ;
  assign n3575 = ~n3573 & ~n3574 ;
  assign n3576 = \ks1_col_reg[17]/NET0131  & ~n1142 ;
  assign n3577 = n1142 & ~n3235 ;
  assign n3578 = ~n3576 & ~n3577 ;
  assign n3579 = \ks1_col_reg[1]/NET0131  & ~n1286 ;
  assign n3580 = n1286 & ~n3235 ;
  assign n3581 = ~n3579 & ~n3580 ;
  assign n3582 = \ks1_col_reg[25]/NET0131  & ~n1274 ;
  assign n3583 = n1274 & ~n3235 ;
  assign n3584 = ~n3582 & ~n3583 ;
  assign n3585 = n1274 & n2400 ;
  assign n3586 = \ks1_col_reg[26]/NET0131  & ~n1274 ;
  assign n3587 = ~n3585 & ~n3586 ;
  assign n3588 = n1286 & n2400 ;
  assign n3589 = \ks1_col_reg[2]/NET0131  & ~n1286 ;
  assign n3590 = ~n3588 & ~n3589 ;
  assign n3591 = \sub1_data_reg_reg[121]/NET0131  & ~n3198 ;
  assign n3592 = n3198 & ~n3235 ;
  assign n3593 = ~n3591 & ~n3592 ;
  assign n3594 = \sub1_data_reg_reg[25]/NET0131  & ~n3205 ;
  assign n3595 = n3205 & ~n3235 ;
  assign n3596 = ~n3594 & ~n3595 ;
  assign n3597 = \sub1_data_reg_reg[57]/NET0131  & ~n3212 ;
  assign n3598 = n3212 & ~n3235 ;
  assign n3599 = ~n3597 & ~n3598 ;
  assign n3600 = \sub1_data_reg_reg[89]/NET0131  & ~n3219 ;
  assign n3601 = n3219 & ~n3235 ;
  assign n3602 = ~n3600 & ~n3601 ;
  assign n3603 = n2400 & n3198 ;
  assign n3604 = \sub1_data_reg_reg[122]/NET0131  & ~n3198 ;
  assign n3605 = ~n3603 & ~n3604 ;
  assign n3606 = n2400 & n3205 ;
  assign n3607 = \sub1_data_reg_reg[26]/NET0131  & ~n3205 ;
  assign n3608 = ~n3606 & ~n3607 ;
  assign n3609 = n2400 & n3212 ;
  assign n3610 = \sub1_data_reg_reg[58]/NET0131  & ~n3212 ;
  assign n3611 = ~n3609 & ~n3610 ;
  assign n3612 = n2400 & n3219 ;
  assign n3613 = \sub1_data_reg_reg[90]/NET0131  & ~n3219 ;
  assign n3614 = ~n3612 & ~n3613 ;
  assign n3615 = ~n2238 & n2294 ;
  assign n3616 = ~n2295 & ~n3615 ;
  assign n3617 = n2193 & n2245 ;
  assign n3618 = ~n2285 & ~n3617 ;
  assign n3622 = ~decrypt_i_pad & \round_reg[0]/NET0131  ;
  assign n3623 = ~\round_reg[1]/NET0131  & n3622 ;
  assign n3624 = n1156 & n3623 ;
  assign n3625 = ~n1260 & ~n3624 ;
  assign n3626 = \state_reg/NET0131  & ~n3625 ;
  assign n3619 = \addroundkey_ready_o_reg/NET0131  & n1159 ;
  assign n3620 = ~decrypt_i_pad & \sub1_ready_o_reg/NET0131  ;
  assign n3621 = ~n3619 & ~n3620 ;
  assign n3627 = ~\mix1_state_reg[0]/NET0131  & ~\mix1_state_reg[1]/NET0131  ;
  assign n3628 = ~n3621 & n3627 ;
  assign n3629 = ~n3626 & n3628 ;
  assign n3645 = ~\sub1_data_reg_reg[114]/NET0131  & ~n1159 ;
  assign n3646 = ~\data_o[114]_pad  & n1159 ;
  assign n3647 = ~n3645 & ~n3646 ;
  assign n3648 = n3629 & n3647 ;
  assign n3642 = ~\data_o[18]_pad  & n1159 ;
  assign n3640 = \mix1_state_reg[0]/NET0131  & \mix1_state_reg[1]/NET0131  ;
  assign n3641 = ~\sub1_data_reg_reg[18]/NET0131  & ~n1159 ;
  assign n3643 = n3640 & ~n3641 ;
  assign n3644 = ~n3642 & n3643 ;
  assign n3632 = ~\data_o[82]_pad  & n1159 ;
  assign n3630 = \mix1_state_reg[0]/NET0131  & ~\mix1_state_reg[1]/NET0131  ;
  assign n3631 = ~\sub1_data_reg_reg[82]/NET0131  & ~n1159 ;
  assign n3633 = n3630 & ~n3631 ;
  assign n3634 = ~n3632 & n3633 ;
  assign n3637 = ~\data_o[50]_pad  & n1159 ;
  assign n3635 = ~\mix1_state_reg[0]/NET0131  & \mix1_state_reg[1]/NET0131  ;
  assign n3636 = ~\sub1_data_reg_reg[50]/NET0131  & ~n1159 ;
  assign n3638 = n3635 & ~n3636 ;
  assign n3639 = ~n3637 & n3638 ;
  assign n3649 = ~n3634 & ~n3639 ;
  assign n3650 = ~n3644 & n3649 ;
  assign n3651 = ~n3648 & n3650 ;
  assign n3664 = ~\sub1_data_reg_reg[103]/NET0131  & ~n1159 ;
  assign n3665 = ~\data_o[103]_pad  & n1159 ;
  assign n3666 = ~n3664 & ~n3665 ;
  assign n3667 = n3629 & n3666 ;
  assign n3661 = ~\data_o[7]_pad  & n1159 ;
  assign n3660 = ~\sub1_data_reg_reg[7]/NET0131  & ~n1159 ;
  assign n3662 = n3640 & ~n3660 ;
  assign n3663 = ~n3661 & n3662 ;
  assign n3653 = ~\data_o[71]_pad  & n1159 ;
  assign n3652 = ~\sub1_data_reg_reg[71]/NET0131  & ~n1159 ;
  assign n3654 = n3630 & ~n3652 ;
  assign n3655 = ~n3653 & n3654 ;
  assign n3657 = ~\data_o[39]_pad  & n1159 ;
  assign n3656 = ~\sub1_data_reg_reg[39]/NET0131  & ~n1159 ;
  assign n3658 = n3635 & ~n3656 ;
  assign n3659 = ~n3657 & n3658 ;
  assign n3668 = ~n3655 & ~n3659 ;
  assign n3669 = ~n3663 & n3668 ;
  assign n3670 = ~n3667 & n3669 ;
  assign n3683 = ~\sub1_data_reg_reg[119]/NET0131  & ~n1159 ;
  assign n3684 = ~\data_o[119]_pad  & n1159 ;
  assign n3685 = ~n3683 & ~n3684 ;
  assign n3686 = n3629 & n3685 ;
  assign n3680 = ~\data_o[23]_pad  & n1159 ;
  assign n3679 = ~\sub1_data_reg_reg[23]/NET0131  & ~n1159 ;
  assign n3681 = n3640 & ~n3679 ;
  assign n3682 = ~n3680 & n3681 ;
  assign n3672 = ~\data_o[55]_pad  & n1159 ;
  assign n3671 = ~\sub1_data_reg_reg[55]/NET0131  & ~n1159 ;
  assign n3673 = n3635 & ~n3671 ;
  assign n3674 = ~n3672 & n3673 ;
  assign n3676 = ~\data_o[87]_pad  & n1159 ;
  assign n3675 = ~\sub1_data_reg_reg[87]/NET0131  & ~n1159 ;
  assign n3677 = n3630 & ~n3675 ;
  assign n3678 = ~n3676 & n3677 ;
  assign n3687 = ~n3674 & ~n3678 ;
  assign n3688 = ~n3682 & n3687 ;
  assign n3689 = ~n3686 & n3688 ;
  assign n3690 = n3670 & ~n3689 ;
  assign n3691 = ~n3670 & n3689 ;
  assign n3692 = ~n3690 & ~n3691 ;
  assign n3705 = ~\sub1_data_reg_reg[117]/NET0131  & ~n1159 ;
  assign n3706 = ~\data_o[117]_pad  & n1159 ;
  assign n3707 = ~n3705 & ~n3706 ;
  assign n3708 = n3629 & n3707 ;
  assign n3702 = ~\data_o[85]_pad  & n1159 ;
  assign n3701 = ~\sub1_data_reg_reg[85]/NET0131  & ~n1159 ;
  assign n3703 = n3630 & ~n3701 ;
  assign n3704 = ~n3702 & n3703 ;
  assign n3694 = ~\data_o[21]_pad  & n1159 ;
  assign n3693 = ~\sub1_data_reg_reg[21]/NET0131  & ~n1159 ;
  assign n3695 = n3640 & ~n3693 ;
  assign n3696 = ~n3694 & n3695 ;
  assign n3698 = ~\data_o[53]_pad  & n1159 ;
  assign n3697 = ~\sub1_data_reg_reg[53]/NET0131  & ~n1159 ;
  assign n3699 = n3635 & ~n3697 ;
  assign n3700 = ~n3698 & n3699 ;
  assign n3709 = ~n3696 & ~n3700 ;
  assign n3710 = ~n3704 & n3709 ;
  assign n3711 = ~n3708 & n3710 ;
  assign n3724 = ~\sub1_data_reg_reg[125]/NET0131  & ~n1159 ;
  assign n3725 = ~\data_o[125]_pad  & n1159 ;
  assign n3726 = ~n3724 & ~n3725 ;
  assign n3727 = n3629 & n3726 ;
  assign n3721 = ~\data_o[93]_pad  & n1159 ;
  assign n3720 = ~\sub1_data_reg_reg[93]/NET0131  & ~n1159 ;
  assign n3722 = n3630 & ~n3720 ;
  assign n3723 = ~n3721 & n3722 ;
  assign n3713 = ~\data_o[29]_pad  & n1159 ;
  assign n3712 = ~\sub1_data_reg_reg[29]/NET0131  & ~n1159 ;
  assign n3714 = n3640 & ~n3712 ;
  assign n3715 = ~n3713 & n3714 ;
  assign n3717 = ~\data_o[61]_pad  & n1159 ;
  assign n3716 = ~\sub1_data_reg_reg[61]/NET0131  & ~n1159 ;
  assign n3718 = n3635 & ~n3716 ;
  assign n3719 = ~n3717 & n3718 ;
  assign n3728 = ~n3715 & ~n3719 ;
  assign n3729 = ~n3723 & n3728 ;
  assign n3730 = ~n3727 & n3729 ;
  assign n3731 = n3711 & ~n3730 ;
  assign n3732 = ~n3711 & n3730 ;
  assign n3733 = ~n3731 & ~n3732 ;
  assign n3746 = ~\sub1_data_reg_reg[101]/NET0131  & ~n1159 ;
  assign n3747 = ~\data_o[101]_pad  & n1159 ;
  assign n3748 = ~n3746 & ~n3747 ;
  assign n3749 = n3629 & n3748 ;
  assign n3743 = ~\data_o[37]_pad  & n1159 ;
  assign n3742 = ~\sub1_data_reg_reg[37]/NET0131  & ~n1159 ;
  assign n3744 = n3635 & ~n3742 ;
  assign n3745 = ~n3743 & n3744 ;
  assign n3735 = ~\data_o[69]_pad  & n1159 ;
  assign n3734 = ~\sub1_data_reg_reg[69]/NET0131  & ~n1159 ;
  assign n3736 = n3630 & ~n3734 ;
  assign n3737 = ~n3735 & n3736 ;
  assign n3739 = ~\data_o[5]_pad  & n1159 ;
  assign n3738 = ~\sub1_data_reg_reg[5]/NET0131  & ~n1159 ;
  assign n3740 = n3640 & ~n3738 ;
  assign n3741 = ~n3739 & n3740 ;
  assign n3750 = ~n3737 & ~n3741 ;
  assign n3751 = ~n3745 & n3750 ;
  assign n3752 = ~n3749 & n3751 ;
  assign n3765 = ~\sub1_data_reg_reg[109]/NET0131  & ~n1159 ;
  assign n3766 = ~\data_o[109]_pad  & n1159 ;
  assign n3767 = ~n3765 & ~n3766 ;
  assign n3768 = n3629 & n3767 ;
  assign n3762 = ~\data_o[13]_pad  & n1159 ;
  assign n3761 = ~\sub1_data_reg_reg[13]/NET0131  & ~n1159 ;
  assign n3763 = n3640 & ~n3761 ;
  assign n3764 = ~n3762 & n3763 ;
  assign n3754 = ~\data_o[45]_pad  & n1159 ;
  assign n3753 = ~\sub1_data_reg_reg[45]/NET0131  & ~n1159 ;
  assign n3755 = n3635 & ~n3753 ;
  assign n3756 = ~n3754 & n3755 ;
  assign n3758 = ~\data_o[77]_pad  & n1159 ;
  assign n3757 = ~\sub1_data_reg_reg[77]/NET0131  & ~n1159 ;
  assign n3759 = n3630 & ~n3757 ;
  assign n3760 = ~n3758 & n3759 ;
  assign n3769 = ~n3756 & ~n3760 ;
  assign n3770 = ~n3764 & n3769 ;
  assign n3771 = ~n3768 & n3770 ;
  assign n3772 = n3752 & ~n3771 ;
  assign n3773 = ~n3752 & n3771 ;
  assign n3774 = ~n3772 & ~n3773 ;
  assign n3775 = n3733 & n3774 ;
  assign n3776 = ~n3733 & ~n3774 ;
  assign n3777 = ~n3775 & ~n3776 ;
  assign n3790 = ~\sub1_data_reg_reg[110]/NET0131  & ~n1159 ;
  assign n3791 = ~\data_o[110]_pad  & n1159 ;
  assign n3792 = ~n3790 & ~n3791 ;
  assign n3793 = n3629 & n3792 ;
  assign n3787 = ~\data_o[14]_pad  & n1159 ;
  assign n3786 = ~\sub1_data_reg_reg[14]/NET0131  & ~n1159 ;
  assign n3788 = n3640 & ~n3786 ;
  assign n3789 = ~n3787 & n3788 ;
  assign n3779 = ~\data_o[46]_pad  & n1159 ;
  assign n3778 = ~\sub1_data_reg_reg[46]/NET0131  & ~n1159 ;
  assign n3780 = n3635 & ~n3778 ;
  assign n3781 = ~n3779 & n3780 ;
  assign n3783 = ~\data_o[78]_pad  & n1159 ;
  assign n3782 = ~\sub1_data_reg_reg[78]/NET0131  & ~n1159 ;
  assign n3784 = n3630 & ~n3782 ;
  assign n3785 = ~n3783 & n3784 ;
  assign n3794 = ~n3781 & ~n3785 ;
  assign n3795 = ~n3789 & n3794 ;
  assign n3796 = ~n3793 & n3795 ;
  assign n3809 = ~\sub1_data_reg_reg[126]/NET0131  & ~n1159 ;
  assign n3810 = ~\data_o[126]_pad  & n1159 ;
  assign n3811 = ~n3809 & ~n3810 ;
  assign n3812 = n3629 & n3811 ;
  assign n3806 = ~\data_o[94]_pad  & n1159 ;
  assign n3805 = ~\sub1_data_reg_reg[94]/NET0131  & ~n1159 ;
  assign n3807 = n3630 & ~n3805 ;
  assign n3808 = ~n3806 & n3807 ;
  assign n3798 = ~\data_o[62]_pad  & n1159 ;
  assign n3797 = ~\sub1_data_reg_reg[62]/NET0131  & ~n1159 ;
  assign n3799 = n3635 & ~n3797 ;
  assign n3800 = ~n3798 & n3799 ;
  assign n3802 = ~\data_o[30]_pad  & n1159 ;
  assign n3801 = ~\sub1_data_reg_reg[30]/NET0131  & ~n1159 ;
  assign n3803 = n3640 & ~n3801 ;
  assign n3804 = ~n3802 & n3803 ;
  assign n3813 = ~n3800 & ~n3804 ;
  assign n3814 = ~n3808 & n3813 ;
  assign n3815 = ~n3812 & n3814 ;
  assign n3816 = n3796 & ~n3815 ;
  assign n3817 = ~n3796 & n3815 ;
  assign n3818 = ~n3816 & ~n3817 ;
  assign n3819 = n3777 & n3818 ;
  assign n3820 = ~n3777 & ~n3818 ;
  assign n3821 = ~n3819 & ~n3820 ;
  assign n3822 = ~n3692 & ~n3821 ;
  assign n3823 = n3692 & n3821 ;
  assign n3824 = ~n3822 & ~n3823 ;
  assign n3837 = ~\sub1_data_reg_reg[98]/NET0131  & ~n1159 ;
  assign n3838 = ~\data_o[98]_pad  & n1159 ;
  assign n3839 = ~n3837 & ~n3838 ;
  assign n3840 = n3629 & n3839 ;
  assign n3834 = ~\data_o[2]_pad  & n1159 ;
  assign n3833 = ~\sub1_data_reg_reg[2]/NET0131  & ~n1159 ;
  assign n3835 = n3640 & ~n3833 ;
  assign n3836 = ~n3834 & n3835 ;
  assign n3826 = ~\data_o[66]_pad  & n1159 ;
  assign n3825 = ~\sub1_data_reg_reg[66]/NET0131  & ~n1159 ;
  assign n3827 = n3630 & ~n3825 ;
  assign n3828 = ~n3826 & n3827 ;
  assign n3830 = ~\data_o[34]_pad  & n1159 ;
  assign n3829 = ~\sub1_data_reg_reg[34]/NET0131  & ~n1159 ;
  assign n3831 = n3635 & ~n3829 ;
  assign n3832 = ~n3830 & n3831 ;
  assign n3841 = ~n3828 & ~n3832 ;
  assign n3842 = ~n3836 & n3841 ;
  assign n3843 = ~n3840 & n3842 ;
  assign n3844 = n3824 & ~n3843 ;
  assign n3845 = ~n3824 & n3843 ;
  assign n3846 = ~n3844 & ~n3845 ;
  assign n3847 = n3651 & n3846 ;
  assign n3848 = ~n3651 & ~n3846 ;
  assign n3849 = ~n3847 & ~n3848 ;
  assign n3862 = ~\sub1_data_reg_reg[97]/NET0131  & ~n1159 ;
  assign n3863 = ~\data_o[97]_pad  & n1159 ;
  assign n3864 = ~n3862 & ~n3863 ;
  assign n3865 = n3629 & n3864 ;
  assign n3859 = ~\data_o[33]_pad  & n1159 ;
  assign n3858 = ~\sub1_data_reg_reg[33]/NET0131  & ~n1159 ;
  assign n3860 = n3635 & ~n3858 ;
  assign n3861 = ~n3859 & n3860 ;
  assign n3851 = ~\data_o[1]_pad  & n1159 ;
  assign n3850 = ~\sub1_data_reg_reg[1]/NET0131  & ~n1159 ;
  assign n3852 = n3640 & ~n3850 ;
  assign n3853 = ~n3851 & n3852 ;
  assign n3855 = ~\data_o[65]_pad  & n1159 ;
  assign n3854 = ~\sub1_data_reg_reg[65]/NET0131  & ~n1159 ;
  assign n3856 = n3630 & ~n3854 ;
  assign n3857 = ~n3855 & n3856 ;
  assign n3866 = ~n3853 & ~n3857 ;
  assign n3867 = ~n3861 & n3866 ;
  assign n3868 = ~n3865 & n3867 ;
  assign n3881 = ~\sub1_data_reg_reg[113]/NET0131  & ~n1159 ;
  assign n3882 = ~\data_o[113]_pad  & n1159 ;
  assign n3883 = ~n3881 & ~n3882 ;
  assign n3884 = n3629 & n3883 ;
  assign n3878 = ~\data_o[49]_pad  & n1159 ;
  assign n3877 = ~\sub1_data_reg_reg[49]/NET0131  & ~n1159 ;
  assign n3879 = n3635 & ~n3877 ;
  assign n3880 = ~n3878 & n3879 ;
  assign n3870 = ~\data_o[17]_pad  & n1159 ;
  assign n3869 = ~\sub1_data_reg_reg[17]/NET0131  & ~n1159 ;
  assign n3871 = n3640 & ~n3869 ;
  assign n3872 = ~n3870 & n3871 ;
  assign n3874 = ~\data_o[81]_pad  & n1159 ;
  assign n3873 = ~\sub1_data_reg_reg[81]/NET0131  & ~n1159 ;
  assign n3875 = n3630 & ~n3873 ;
  assign n3876 = ~n3874 & n3875 ;
  assign n3885 = ~n3872 & ~n3876 ;
  assign n3886 = ~n3880 & n3885 ;
  assign n3887 = ~n3884 & n3886 ;
  assign n3888 = n3868 & ~n3887 ;
  assign n3889 = ~n3868 & n3887 ;
  assign n3890 = ~n3888 & ~n3889 ;
  assign n3903 = ~\sub1_data_reg_reg[121]/NET0131  & ~n1159 ;
  assign n3904 = ~\data_o[121]_pad  & n1159 ;
  assign n3905 = ~n3903 & ~n3904 ;
  assign n3906 = n3629 & n3905 ;
  assign n3900 = ~\data_o[89]_pad  & n1159 ;
  assign n3899 = ~\sub1_data_reg_reg[89]/NET0131  & ~n1159 ;
  assign n3901 = n3630 & ~n3899 ;
  assign n3902 = ~n3900 & n3901 ;
  assign n3892 = ~\data_o[25]_pad  & n1159 ;
  assign n3891 = ~\sub1_data_reg_reg[25]/NET0131  & ~n1159 ;
  assign n3893 = n3640 & ~n3891 ;
  assign n3894 = ~n3892 & n3893 ;
  assign n3896 = ~\data_o[57]_pad  & n1159 ;
  assign n3895 = ~\sub1_data_reg_reg[57]/NET0131  & ~n1159 ;
  assign n3897 = n3635 & ~n3895 ;
  assign n3898 = ~n3896 & n3897 ;
  assign n3907 = ~n3894 & ~n3898 ;
  assign n3908 = ~n3902 & n3907 ;
  assign n3909 = ~n3906 & n3908 ;
  assign n3922 = ~\sub1_data_reg_reg[105]/NET0131  & ~n1159 ;
  assign n3923 = ~\data_o[105]_pad  & n1159 ;
  assign n3924 = ~n3922 & ~n3923 ;
  assign n3925 = n3629 & n3924 ;
  assign n3919 = ~\data_o[41]_pad  & n1159 ;
  assign n3918 = ~\sub1_data_reg_reg[41]/NET0131  & ~n1159 ;
  assign n3920 = n3635 & ~n3918 ;
  assign n3921 = ~n3919 & n3920 ;
  assign n3911 = ~\data_o[9]_pad  & n1159 ;
  assign n3910 = ~\sub1_data_reg_reg[9]/NET0131  & ~n1159 ;
  assign n3912 = n3640 & ~n3910 ;
  assign n3913 = ~n3911 & n3912 ;
  assign n3915 = ~\data_o[73]_pad  & n1159 ;
  assign n3914 = ~\sub1_data_reg_reg[73]/NET0131  & ~n1159 ;
  assign n3916 = n3630 & ~n3914 ;
  assign n3917 = ~n3915 & n3916 ;
  assign n3926 = ~n3913 & ~n3917 ;
  assign n3927 = ~n3921 & n3926 ;
  assign n3928 = ~n3925 & n3927 ;
  assign n3929 = n3909 & ~n3928 ;
  assign n3930 = ~n3909 & n3928 ;
  assign n3931 = ~n3929 & ~n3930 ;
  assign n3932 = n3890 & n3931 ;
  assign n3933 = ~n3890 & ~n3931 ;
  assign n3934 = ~n3932 & ~n3933 ;
  assign n3936 = n3849 & ~n3934 ;
  assign n3935 = ~n3849 & n3934 ;
  assign n3937 = decrypt_i_pad & ~n3935 ;
  assign n3938 = ~n3936 & n3937 ;
  assign n3951 = ~\sub1_data_reg_reg[116]/NET0131  & ~n1159 ;
  assign n3952 = ~\data_o[116]_pad  & n1159 ;
  assign n3953 = ~n3951 & ~n3952 ;
  assign n3954 = n3629 & n3953 ;
  assign n3948 = ~\data_o[52]_pad  & n1159 ;
  assign n3947 = ~\sub1_data_reg_reg[52]/NET0131  & ~n1159 ;
  assign n3949 = n3635 & ~n3947 ;
  assign n3950 = ~n3948 & n3949 ;
  assign n3940 = ~\data_o[84]_pad  & n1159 ;
  assign n3939 = ~\sub1_data_reg_reg[84]/NET0131  & ~n1159 ;
  assign n3941 = n3630 & ~n3939 ;
  assign n3942 = ~n3940 & n3941 ;
  assign n3944 = ~\data_o[20]_pad  & n1159 ;
  assign n3943 = ~\sub1_data_reg_reg[20]/NET0131  & ~n1159 ;
  assign n3945 = n3640 & ~n3943 ;
  assign n3946 = ~n3944 & n3945 ;
  assign n3955 = ~n3942 & ~n3946 ;
  assign n3956 = ~n3950 & n3955 ;
  assign n3957 = ~n3954 & n3956 ;
  assign n3970 = ~\sub1_data_reg_reg[124]/NET0131  & ~n1159 ;
  assign n3971 = ~\data_o[124]_pad  & n1159 ;
  assign n3972 = ~n3970 & ~n3971 ;
  assign n3973 = n3629 & n3972 ;
  assign n3967 = ~\data_o[60]_pad  & n1159 ;
  assign n3966 = ~\sub1_data_reg_reg[60]/NET0131  & ~n1159 ;
  assign n3968 = n3635 & ~n3966 ;
  assign n3969 = ~n3967 & n3968 ;
  assign n3959 = ~\data_o[28]_pad  & n1159 ;
  assign n3958 = ~\sub1_data_reg_reg[28]/NET0131  & ~n1159 ;
  assign n3960 = n3640 & ~n3958 ;
  assign n3961 = ~n3959 & n3960 ;
  assign n3963 = ~\data_o[92]_pad  & n1159 ;
  assign n3962 = ~\sub1_data_reg_reg[92]/NET0131  & ~n1159 ;
  assign n3964 = n3630 & ~n3962 ;
  assign n3965 = ~n3963 & n3964 ;
  assign n3974 = ~n3961 & ~n3965 ;
  assign n3975 = ~n3969 & n3974 ;
  assign n3976 = ~n3973 & n3975 ;
  assign n3989 = ~\sub1_data_reg_reg[108]/NET0131  & ~n1159 ;
  assign n3990 = ~\data_o[108]_pad  & n1159 ;
  assign n3991 = ~n3989 & ~n3990 ;
  assign n3992 = n3629 & n3991 ;
  assign n3986 = ~\data_o[44]_pad  & n1159 ;
  assign n3985 = ~\sub1_data_reg_reg[44]/NET0131  & ~n1159 ;
  assign n3987 = n3635 & ~n3985 ;
  assign n3988 = ~n3986 & n3987 ;
  assign n3978 = ~\data_o[12]_pad  & n1159 ;
  assign n3977 = ~\sub1_data_reg_reg[12]/NET0131  & ~n1159 ;
  assign n3979 = n3640 & ~n3977 ;
  assign n3980 = ~n3978 & n3979 ;
  assign n3982 = ~\data_o[76]_pad  & n1159 ;
  assign n3981 = ~\sub1_data_reg_reg[76]/NET0131  & ~n1159 ;
  assign n3983 = n3630 & ~n3981 ;
  assign n3984 = ~n3982 & n3983 ;
  assign n3993 = ~n3980 & ~n3984 ;
  assign n3994 = ~n3988 & n3993 ;
  assign n3995 = ~n3992 & n3994 ;
  assign n3996 = n3976 & ~n3995 ;
  assign n3997 = ~n3976 & n3995 ;
  assign n3998 = ~n3996 & ~n3997 ;
  assign n3999 = n3957 & n3998 ;
  assign n4000 = ~n3957 & ~n3998 ;
  assign n4001 = ~n3999 & ~n4000 ;
  assign n4014 = ~\sub1_data_reg_reg[123]/NET0131  & ~n1159 ;
  assign n4015 = ~\data_o[123]_pad  & n1159 ;
  assign n4016 = ~n4014 & ~n4015 ;
  assign n4017 = n3629 & n4016 ;
  assign n4011 = ~\data_o[27]_pad  & n1159 ;
  assign n4010 = ~\sub1_data_reg_reg[27]/NET0131  & ~n1159 ;
  assign n4012 = n3640 & ~n4010 ;
  assign n4013 = ~n4011 & n4012 ;
  assign n4003 = ~\data_o[91]_pad  & n1159 ;
  assign n4002 = ~\sub1_data_reg_reg[91]/NET0131  & ~n1159 ;
  assign n4004 = n3630 & ~n4002 ;
  assign n4005 = ~n4003 & n4004 ;
  assign n4007 = ~\data_o[59]_pad  & n1159 ;
  assign n4006 = ~\sub1_data_reg_reg[59]/NET0131  & ~n1159 ;
  assign n4008 = n3635 & ~n4006 ;
  assign n4009 = ~n4007 & n4008 ;
  assign n4018 = ~n4005 & ~n4009 ;
  assign n4019 = ~n4013 & n4018 ;
  assign n4020 = ~n4017 & n4019 ;
  assign n4033 = ~\sub1_data_reg_reg[99]/NET0131  & ~n1159 ;
  assign n4034 = ~\data_o[99]_pad  & n1159 ;
  assign n4035 = ~n4033 & ~n4034 ;
  assign n4036 = n3629 & n4035 ;
  assign n4030 = ~\data_o[3]_pad  & n1159 ;
  assign n4029 = ~\sub1_data_reg_reg[3]/NET0131  & ~n1159 ;
  assign n4031 = n3640 & ~n4029 ;
  assign n4032 = ~n4030 & n4031 ;
  assign n4022 = ~\data_o[35]_pad  & n1159 ;
  assign n4021 = ~\sub1_data_reg_reg[35]/NET0131  & ~n1159 ;
  assign n4023 = n3635 & ~n4021 ;
  assign n4024 = ~n4022 & n4023 ;
  assign n4026 = ~\data_o[67]_pad  & n1159 ;
  assign n4025 = ~\sub1_data_reg_reg[67]/NET0131  & ~n1159 ;
  assign n4027 = n3630 & ~n4025 ;
  assign n4028 = ~n4026 & n4027 ;
  assign n4037 = ~n4024 & ~n4028 ;
  assign n4038 = ~n4032 & n4037 ;
  assign n4039 = ~n4036 & n4038 ;
  assign n4040 = n4020 & ~n4039 ;
  assign n4041 = ~n4020 & n4039 ;
  assign n4042 = ~n4040 & ~n4041 ;
  assign n4055 = ~\sub1_data_reg_reg[127]/NET0131  & ~n1159 ;
  assign n4056 = ~\data_o[127]_pad  & n1159 ;
  assign n4057 = ~n4055 & ~n4056 ;
  assign n4058 = n3629 & n4057 ;
  assign n4052 = ~\data_o[63]_pad  & n1159 ;
  assign n4051 = ~\sub1_data_reg_reg[63]/NET0131  & ~n1159 ;
  assign n4053 = n3635 & ~n4051 ;
  assign n4054 = ~n4052 & n4053 ;
  assign n4044 = ~\data_o[95]_pad  & n1159 ;
  assign n4043 = ~\sub1_data_reg_reg[95]/NET0131  & ~n1159 ;
  assign n4045 = n3630 & ~n4043 ;
  assign n4046 = ~n4044 & n4045 ;
  assign n4048 = ~\data_o[31]_pad  & n1159 ;
  assign n4047 = ~\sub1_data_reg_reg[31]/NET0131  & ~n1159 ;
  assign n4049 = n3640 & ~n4047 ;
  assign n4050 = ~n4048 & n4049 ;
  assign n4059 = ~n4046 & ~n4050 ;
  assign n4060 = ~n4054 & n4059 ;
  assign n4061 = ~n4058 & n4060 ;
  assign n4062 = n3670 & ~n4061 ;
  assign n4063 = ~n3670 & n4061 ;
  assign n4064 = ~n4062 & ~n4063 ;
  assign n4065 = n4042 & n4064 ;
  assign n4066 = ~n4042 & ~n4064 ;
  assign n4067 = ~n4065 & ~n4066 ;
  assign n4068 = n4001 & ~n4067 ;
  assign n4069 = ~n4001 & n4067 ;
  assign n4070 = ~n4068 & ~n4069 ;
  assign n4071 = n3938 & n4070 ;
  assign n4072 = ~n3938 & ~n4070 ;
  assign n4073 = ~n4071 & ~n4072 ;
  assign n4074 = n3629 & ~n4073 ;
  assign n4075 = \mix1_data_reg_reg[100]/NET0131  & ~n3629 ;
  assign n4076 = ~n4074 & ~n4075 ;
  assign n4077 = n3771 & ~n3976 ;
  assign n4078 = ~n3771 & n3976 ;
  assign n4079 = ~n4077 & ~n4078 ;
  assign n4080 = n3733 & ~n4079 ;
  assign n4081 = ~n3733 & n4079 ;
  assign n4082 = ~n4080 & ~n4081 ;
  assign n4095 = ~\sub1_data_reg_reg[100]/NET0131  & ~n1159 ;
  assign n4096 = ~\data_o[100]_pad  & n1159 ;
  assign n4097 = ~n4095 & ~n4096 ;
  assign n4098 = n3629 & n4097 ;
  assign n4092 = ~\data_o[4]_pad  & n1159 ;
  assign n4091 = ~\sub1_data_reg_reg[4]/NET0131  & ~n1159 ;
  assign n4093 = n3640 & ~n4091 ;
  assign n4094 = ~n4092 & n4093 ;
  assign n4084 = ~\data_o[36]_pad  & n1159 ;
  assign n4083 = ~\sub1_data_reg_reg[36]/NET0131  & ~n1159 ;
  assign n4085 = n3635 & ~n4083 ;
  assign n4086 = ~n4084 & n4085 ;
  assign n4088 = ~\data_o[68]_pad  & n1159 ;
  assign n4087 = ~\sub1_data_reg_reg[68]/NET0131  & ~n1159 ;
  assign n4089 = n3630 & ~n4087 ;
  assign n4090 = ~n4088 & n4089 ;
  assign n4099 = ~n4086 & ~n4090 ;
  assign n4100 = ~n4094 & n4099 ;
  assign n4101 = ~n4098 & n4100 ;
  assign n4114 = ~\sub1_data_reg_reg[102]/NET0131  & ~n1159 ;
  assign n4115 = ~\data_o[102]_pad  & n1159 ;
  assign n4116 = ~n4114 & ~n4115 ;
  assign n4117 = n3629 & n4116 ;
  assign n4111 = ~\data_o[6]_pad  & n1159 ;
  assign n4110 = ~\sub1_data_reg_reg[6]/NET0131  & ~n1159 ;
  assign n4112 = n3640 & ~n4110 ;
  assign n4113 = ~n4111 & n4112 ;
  assign n4103 = ~\data_o[38]_pad  & n1159 ;
  assign n4102 = ~\sub1_data_reg_reg[38]/NET0131  & ~n1159 ;
  assign n4104 = n3635 & ~n4102 ;
  assign n4105 = ~n4103 & n4104 ;
  assign n4107 = ~\data_o[70]_pad  & n1159 ;
  assign n4106 = ~\sub1_data_reg_reg[70]/NET0131  & ~n1159 ;
  assign n4108 = n3630 & ~n4106 ;
  assign n4109 = ~n4107 & n4108 ;
  assign n4118 = ~n4105 & ~n4109 ;
  assign n4119 = ~n4113 & n4118 ;
  assign n4120 = ~n4117 & n4119 ;
  assign n4121 = n3815 & ~n4120 ;
  assign n4122 = ~n3815 & n4120 ;
  assign n4123 = ~n4121 & ~n4122 ;
  assign n4136 = ~\sub1_data_reg_reg[118]/NET0131  & ~n1159 ;
  assign n4137 = ~\data_o[118]_pad  & n1159 ;
  assign n4138 = ~n4136 & ~n4137 ;
  assign n4139 = n3629 & n4138 ;
  assign n4133 = ~\data_o[86]_pad  & n1159 ;
  assign n4132 = ~\sub1_data_reg_reg[86]/NET0131  & ~n1159 ;
  assign n4134 = n3630 & ~n4132 ;
  assign n4135 = ~n4133 & n4134 ;
  assign n4125 = ~\data_o[54]_pad  & n1159 ;
  assign n4124 = ~\sub1_data_reg_reg[54]/NET0131  & ~n1159 ;
  assign n4126 = n3635 & ~n4124 ;
  assign n4127 = ~n4125 & n4126 ;
  assign n4129 = ~\data_o[22]_pad  & n1159 ;
  assign n4128 = ~\sub1_data_reg_reg[22]/NET0131  & ~n1159 ;
  assign n4130 = n3640 & ~n4128 ;
  assign n4131 = ~n4129 & n4130 ;
  assign n4140 = ~n4127 & ~n4131 ;
  assign n4141 = ~n4135 & n4140 ;
  assign n4142 = ~n4139 & n4141 ;
  assign n4143 = ~n3796 & ~n4142 ;
  assign n4144 = n3796 & n4142 ;
  assign n4145 = ~n4143 & ~n4144 ;
  assign n4146 = n3692 & ~n4145 ;
  assign n4147 = ~n3692 & n4145 ;
  assign n4148 = ~n4146 & ~n4147 ;
  assign n4149 = n4123 & n4148 ;
  assign n4150 = ~n4123 & ~n4148 ;
  assign n4151 = ~n4149 & ~n4150 ;
  assign n4152 = n4039 & n4151 ;
  assign n4153 = ~n4039 & ~n4151 ;
  assign n4154 = ~n4152 & ~n4153 ;
  assign n4167 = ~\sub1_data_reg_reg[115]/NET0131  & ~n1159 ;
  assign n4168 = ~\data_o[115]_pad  & n1159 ;
  assign n4169 = ~n4167 & ~n4168 ;
  assign n4170 = n3629 & n4169 ;
  assign n4164 = ~\data_o[19]_pad  & n1159 ;
  assign n4163 = ~\sub1_data_reg_reg[19]/NET0131  & ~n1159 ;
  assign n4165 = n3640 & ~n4163 ;
  assign n4166 = ~n4164 & n4165 ;
  assign n4156 = ~\data_o[51]_pad  & n1159 ;
  assign n4155 = ~\sub1_data_reg_reg[51]/NET0131  & ~n1159 ;
  assign n4157 = n3635 & ~n4155 ;
  assign n4158 = ~n4156 & n4157 ;
  assign n4160 = ~\data_o[83]_pad  & n1159 ;
  assign n4159 = ~\sub1_data_reg_reg[83]/NET0131  & ~n1159 ;
  assign n4161 = n3630 & ~n4159 ;
  assign n4162 = ~n4160 & n4161 ;
  assign n4171 = ~n4158 & ~n4162 ;
  assign n4172 = ~n4166 & n4171 ;
  assign n4173 = ~n4170 & n4172 ;
  assign n4186 = ~\sub1_data_reg_reg[122]/NET0131  & ~n1159 ;
  assign n4187 = ~\data_o[122]_pad  & n1159 ;
  assign n4188 = ~n4186 & ~n4187 ;
  assign n4189 = n3629 & n4188 ;
  assign n4183 = ~\data_o[90]_pad  & n1159 ;
  assign n4182 = ~\sub1_data_reg_reg[90]/NET0131  & ~n1159 ;
  assign n4184 = n3630 & ~n4182 ;
  assign n4185 = ~n4183 & n4184 ;
  assign n4175 = ~\data_o[58]_pad  & n1159 ;
  assign n4174 = ~\sub1_data_reg_reg[58]/NET0131  & ~n1159 ;
  assign n4176 = n3635 & ~n4174 ;
  assign n4177 = ~n4175 & n4176 ;
  assign n4179 = ~\data_o[26]_pad  & n1159 ;
  assign n4178 = ~\sub1_data_reg_reg[26]/NET0131  & ~n1159 ;
  assign n4180 = n3640 & ~n4178 ;
  assign n4181 = ~n4179 & n4180 ;
  assign n4190 = ~n4177 & ~n4181 ;
  assign n4191 = ~n4185 & n4190 ;
  assign n4192 = ~n4189 & n4191 ;
  assign n4193 = n3843 & ~n4064 ;
  assign n4194 = ~n3843 & n4064 ;
  assign n4195 = ~n4193 & ~n4194 ;
  assign n4196 = n4192 & n4195 ;
  assign n4197 = ~n4192 & ~n4195 ;
  assign n4198 = ~n4196 & ~n4197 ;
  assign n4199 = n4173 & n4198 ;
  assign n4200 = ~n4173 & ~n4198 ;
  assign n4201 = ~n4199 & ~n4200 ;
  assign n4214 = ~\sub1_data_reg_reg[111]/NET0131  & ~n1159 ;
  assign n4215 = ~\data_o[111]_pad  & n1159 ;
  assign n4216 = ~n4214 & ~n4215 ;
  assign n4217 = n3629 & n4216 ;
  assign n4211 = ~\data_o[15]_pad  & n1159 ;
  assign n4210 = ~\sub1_data_reg_reg[15]/NET0131  & ~n1159 ;
  assign n4212 = n3640 & ~n4210 ;
  assign n4213 = ~n4211 & n4212 ;
  assign n4203 = ~\data_o[79]_pad  & n1159 ;
  assign n4202 = ~\sub1_data_reg_reg[79]/NET0131  & ~n1159 ;
  assign n4204 = n3630 & ~n4202 ;
  assign n4205 = ~n4203 & n4204 ;
  assign n4207 = ~\data_o[47]_pad  & n1159 ;
  assign n4206 = ~\sub1_data_reg_reg[47]/NET0131  & ~n1159 ;
  assign n4208 = n3635 & ~n4206 ;
  assign n4209 = ~n4207 & n4208 ;
  assign n4218 = ~n4205 & ~n4209 ;
  assign n4219 = ~n4213 & n4218 ;
  assign n4220 = ~n4217 & n4219 ;
  assign n4221 = n3689 & ~n4220 ;
  assign n4222 = ~n3689 & n4220 ;
  assign n4223 = ~n4221 & ~n4222 ;
  assign n4236 = ~\sub1_data_reg_reg[106]/NET0131  & ~n1159 ;
  assign n4237 = ~\data_o[106]_pad  & n1159 ;
  assign n4238 = ~n4236 & ~n4237 ;
  assign n4239 = n3629 & n4238 ;
  assign n4233 = ~\data_o[74]_pad  & n1159 ;
  assign n4232 = ~\sub1_data_reg_reg[74]/NET0131  & ~n1159 ;
  assign n4234 = n3630 & ~n4232 ;
  assign n4235 = ~n4233 & n4234 ;
  assign n4225 = ~\data_o[10]_pad  & n1159 ;
  assign n4224 = ~\sub1_data_reg_reg[10]/NET0131  & ~n1159 ;
  assign n4226 = n3640 & ~n4224 ;
  assign n4227 = ~n4225 & n4226 ;
  assign n4229 = ~\data_o[42]_pad  & n1159 ;
  assign n4228 = ~\sub1_data_reg_reg[42]/NET0131  & ~n1159 ;
  assign n4230 = n3635 & ~n4228 ;
  assign n4231 = ~n4229 & n4230 ;
  assign n4240 = ~n4227 & ~n4231 ;
  assign n4241 = ~n4235 & n4240 ;
  assign n4242 = ~n4239 & n4241 ;
  assign n4243 = ~n3651 & ~n4242 ;
  assign n4244 = n3651 & n4242 ;
  assign n4245 = ~n4243 & ~n4244 ;
  assign n4246 = n4223 & n4245 ;
  assign n4247 = ~n4223 & ~n4245 ;
  assign n4248 = ~n4246 & ~n4247 ;
  assign n4249 = n4201 & n4248 ;
  assign n4250 = ~n4201 & ~n4248 ;
  assign n4251 = ~n4249 & ~n4250 ;
  assign n4253 = n4154 & n4251 ;
  assign n4252 = ~n4154 & ~n4251 ;
  assign n4254 = decrypt_i_pad & ~n4252 ;
  assign n4255 = ~n4253 & n4254 ;
  assign n4256 = n4101 & ~n4255 ;
  assign n4257 = ~n4101 & n4255 ;
  assign n4258 = ~n4256 & ~n4257 ;
  assign n4259 = n4082 & n4258 ;
  assign n4260 = ~n4082 & ~n4258 ;
  assign n4261 = ~n4259 & ~n4260 ;
  assign n4262 = n3629 & ~n4261 ;
  assign n4263 = \mix1_data_reg_reg[101]/NET0131  & ~n3629 ;
  assign n4264 = ~n4262 & ~n4263 ;
  assign n4265 = \mix1_data_reg_reg[107]/NET0131  & ~n3629 ;
  assign n4266 = n3670 & ~n4220 ;
  assign n4267 = ~n3670 & n4220 ;
  assign n4268 = ~n4266 & ~n4267 ;
  assign n4269 = ~n3843 & ~n4242 ;
  assign n4270 = n3843 & n4242 ;
  assign n4271 = ~n4269 & ~n4270 ;
  assign n4272 = n4268 & n4271 ;
  assign n4273 = ~n4268 & ~n4271 ;
  assign n4274 = ~n4272 & ~n4273 ;
  assign n4287 = ~\sub1_data_reg_reg[104]/NET0131  & ~n1159 ;
  assign n4288 = ~\data_o[104]_pad  & n1159 ;
  assign n4289 = ~n4287 & ~n4288 ;
  assign n4290 = n3629 & n4289 ;
  assign n4284 = ~\data_o[72]_pad  & n1159 ;
  assign n4283 = ~\sub1_data_reg_reg[72]/NET0131  & ~n1159 ;
  assign n4285 = n3630 & ~n4283 ;
  assign n4286 = ~n4284 & n4285 ;
  assign n4276 = ~\data_o[8]_pad  & n1159 ;
  assign n4275 = ~\sub1_data_reg_reg[8]/NET0131  & ~n1159 ;
  assign n4277 = n3640 & ~n4275 ;
  assign n4278 = ~n4276 & n4277 ;
  assign n4280 = ~\data_o[40]_pad  & n1159 ;
  assign n4279 = ~\sub1_data_reg_reg[40]/NET0131  & ~n1159 ;
  assign n4281 = n3635 & ~n4279 ;
  assign n4282 = ~n4280 & n4281 ;
  assign n4291 = ~n4278 & ~n4282 ;
  assign n4292 = ~n4286 & n4291 ;
  assign n4293 = ~n4290 & n4292 ;
  assign n4306 = ~\sub1_data_reg_reg[96]/NET0131  & ~n1159 ;
  assign n4307 = ~\data_o[96]_pad  & n1159 ;
  assign n4308 = ~n4306 & ~n4307 ;
  assign n4309 = n3629 & n4308 ;
  assign n4303 = ~\data_o[0]_pad  & n1159 ;
  assign n4302 = ~\sub1_data_reg_reg[0]/NET0131  & ~n1159 ;
  assign n4304 = n3640 & ~n4302 ;
  assign n4305 = ~n4303 & n4304 ;
  assign n4295 = ~\data_o[32]_pad  & n1159 ;
  assign n4294 = ~\sub1_data_reg_reg[32]/NET0131  & ~n1159 ;
  assign n4296 = n3635 & ~n4294 ;
  assign n4297 = ~n4295 & n4296 ;
  assign n4299 = ~\data_o[64]_pad  & n1159 ;
  assign n4298 = ~\sub1_data_reg_reg[64]/NET0131  & ~n1159 ;
  assign n4300 = n3630 & ~n4298 ;
  assign n4301 = ~n4299 & n4300 ;
  assign n4310 = ~n4297 & ~n4301 ;
  assign n4311 = ~n4305 & n4310 ;
  assign n4312 = ~n4309 & n4311 ;
  assign n4313 = ~n4268 & ~n4312 ;
  assign n4314 = n4268 & n4312 ;
  assign n4315 = ~n4313 & ~n4314 ;
  assign n4316 = ~n4293 & ~n4315 ;
  assign n4317 = n4293 & n4315 ;
  assign n4318 = ~n4316 & ~n4317 ;
  assign n4319 = ~n3821 & ~n3909 ;
  assign n4320 = n3821 & n3909 ;
  assign n4321 = ~n4319 & ~n4320 ;
  assign n4322 = ~n3689 & ~n4061 ;
  assign n4323 = n3689 & n4061 ;
  assign n4324 = ~n4322 & ~n4323 ;
  assign n4337 = ~\sub1_data_reg_reg[112]/NET0131  & ~n1159 ;
  assign n4338 = ~\data_o[112]_pad  & n1159 ;
  assign n4339 = ~n4337 & ~n4338 ;
  assign n4340 = n3629 & n4339 ;
  assign n4334 = ~\data_o[16]_pad  & n1159 ;
  assign n4333 = ~\sub1_data_reg_reg[16]/NET0131  & ~n1159 ;
  assign n4335 = n3640 & ~n4333 ;
  assign n4336 = ~n4334 & n4335 ;
  assign n4326 = ~\data_o[80]_pad  & n1159 ;
  assign n4325 = ~\sub1_data_reg_reg[80]/NET0131  & ~n1159 ;
  assign n4327 = n3630 & ~n4325 ;
  assign n4328 = ~n4326 & n4327 ;
  assign n4330 = ~\data_o[48]_pad  & n1159 ;
  assign n4329 = ~\sub1_data_reg_reg[48]/NET0131  & ~n1159 ;
  assign n4331 = n3635 & ~n4329 ;
  assign n4332 = ~n4330 & n4331 ;
  assign n4341 = ~n4328 & ~n4332 ;
  assign n4342 = ~n4336 & n4341 ;
  assign n4343 = ~n4340 & n4342 ;
  assign n4356 = ~\sub1_data_reg_reg[120]/NET0131  & ~n1159 ;
  assign n4357 = ~\data_o[120]_pad  & n1159 ;
  assign n4358 = ~n4356 & ~n4357 ;
  assign n4359 = n3629 & n4358 ;
  assign n4353 = ~\data_o[56]_pad  & n1159 ;
  assign n4352 = ~\sub1_data_reg_reg[56]/NET0131  & ~n1159 ;
  assign n4354 = n3635 & ~n4352 ;
  assign n4355 = ~n4353 & n4354 ;
  assign n4345 = ~\data_o[24]_pad  & n1159 ;
  assign n4344 = ~\sub1_data_reg_reg[24]/NET0131  & ~n1159 ;
  assign n4346 = n3640 & ~n4344 ;
  assign n4347 = ~n4345 & n4346 ;
  assign n4349 = ~\data_o[88]_pad  & n1159 ;
  assign n4348 = ~\sub1_data_reg_reg[88]/NET0131  & ~n1159 ;
  assign n4350 = n3630 & ~n4348 ;
  assign n4351 = ~n4349 & n4350 ;
  assign n4360 = ~n4347 & ~n4351 ;
  assign n4361 = ~n4355 & n4360 ;
  assign n4362 = ~n4359 & n4361 ;
  assign n4363 = ~n4343 & ~n4362 ;
  assign n4364 = n4343 & n4362 ;
  assign n4365 = ~n4363 & ~n4364 ;
  assign n4366 = n3928 & ~n4365 ;
  assign n4367 = ~n3928 & n4365 ;
  assign n4368 = ~n4366 & ~n4367 ;
  assign n4369 = n4324 & n4368 ;
  assign n4370 = ~n4324 & ~n4368 ;
  assign n4371 = ~n4369 & ~n4370 ;
  assign n4372 = n4321 & n4371 ;
  assign n4373 = ~n4321 & ~n4371 ;
  assign n4374 = ~n4372 & ~n4373 ;
  assign n4376 = ~n4318 & n4374 ;
  assign n4375 = n4318 & ~n4374 ;
  assign n4377 = decrypt_i_pad & ~n4375 ;
  assign n4378 = ~n4376 & n4377 ;
  assign n4379 = n4173 & ~n4378 ;
  assign n4380 = ~n4173 & n4378 ;
  assign n4381 = ~n4379 & ~n4380 ;
  assign n4382 = n4042 & ~n4381 ;
  assign n4383 = ~n4042 & n4381 ;
  assign n4384 = ~n4382 & ~n4383 ;
  assign n4385 = n4274 & n4384 ;
  assign n4386 = ~n4274 & ~n4384 ;
  assign n4387 = ~n4385 & ~n4386 ;
  assign n4388 = n3629 & ~n4387 ;
  assign n4389 = ~n4265 & ~n4388 ;
  assign n4390 = ~n4192 & ~n4242 ;
  assign n4391 = n4192 & n4242 ;
  assign n4392 = ~n4390 & ~n4391 ;
  assign n4393 = ~n4145 & ~n4220 ;
  assign n4394 = n4145 & n4220 ;
  assign n4395 = ~n4393 & ~n4394 ;
  assign n4396 = ~n4061 & ~n4123 ;
  assign n4397 = n4061 & n4123 ;
  assign n4398 = ~n4396 & ~n4397 ;
  assign n4399 = n4395 & n4398 ;
  assign n4400 = ~n4395 & ~n4398 ;
  assign n4401 = ~n4399 & ~n4400 ;
  assign n4402 = n3821 & n4401 ;
  assign n4403 = ~n3821 & ~n4401 ;
  assign n4404 = ~n4402 & ~n4403 ;
  assign n4405 = n4392 & n4404 ;
  assign n4406 = ~n4392 & ~n4404 ;
  assign n4407 = ~n4405 & ~n4406 ;
  assign n4409 = n3934 & n4407 ;
  assign n4408 = ~n3934 & ~n4407 ;
  assign n4410 = decrypt_i_pad & ~n4408 ;
  assign n4411 = ~n4409 & n4410 ;
  assign n4412 = n4101 & ~n4411 ;
  assign n4413 = ~n4101 & n4411 ;
  assign n4414 = ~n4412 & ~n4413 ;
  assign n4415 = n4268 & ~n4414 ;
  assign n4416 = ~n4268 & n4414 ;
  assign n4417 = ~n4415 & ~n4416 ;
  assign n4430 = ~\sub1_data_reg_reg[107]/NET0131  & ~n1159 ;
  assign n4431 = ~\data_o[107]_pad  & n1159 ;
  assign n4432 = ~n4430 & ~n4431 ;
  assign n4433 = n3629 & n4432 ;
  assign n4427 = ~\data_o[75]_pad  & n1159 ;
  assign n4426 = ~\sub1_data_reg_reg[75]/NET0131  & ~n1159 ;
  assign n4428 = n3630 & ~n4426 ;
  assign n4429 = ~n4427 & n4428 ;
  assign n4419 = ~\data_o[11]_pad  & n1159 ;
  assign n4418 = ~\sub1_data_reg_reg[11]/NET0131  & ~n1159 ;
  assign n4420 = n3640 & ~n4418 ;
  assign n4421 = ~n4419 & n4420 ;
  assign n4423 = ~\data_o[43]_pad  & n1159 ;
  assign n4422 = ~\sub1_data_reg_reg[43]/NET0131  & ~n1159 ;
  assign n4424 = n3635 & ~n4422 ;
  assign n4425 = ~n4423 & n4424 ;
  assign n4434 = ~n4421 & ~n4425 ;
  assign n4435 = ~n4429 & n4434 ;
  assign n4436 = ~n4433 & n4435 ;
  assign n4437 = n4039 & ~n4436 ;
  assign n4438 = ~n4039 & n4436 ;
  assign n4439 = ~n4437 & ~n4438 ;
  assign n4440 = ~n3957 & n3976 ;
  assign n4441 = n3957 & ~n3976 ;
  assign n4442 = ~n4440 & ~n4441 ;
  assign n4443 = n4439 & ~n4442 ;
  assign n4444 = ~n4439 & n4442 ;
  assign n4445 = ~n4443 & ~n4444 ;
  assign n4446 = n4417 & n4445 ;
  assign n4447 = ~n4417 & ~n4445 ;
  assign n4448 = ~n4446 & ~n4447 ;
  assign n4449 = n3629 & ~n4448 ;
  assign n4450 = \mix1_data_reg_reg[108]/NET0131  & ~n3629 ;
  assign n4451 = ~n4449 & ~n4450 ;
  assign n4452 = n3711 & ~n3752 ;
  assign n4453 = ~n3711 & n3752 ;
  assign n4454 = ~n4452 & ~n4453 ;
  assign n4455 = ~n4101 & ~n4454 ;
  assign n4456 = n4101 & n4454 ;
  assign n4457 = ~n4455 & ~n4456 ;
  assign n4458 = n4401 & ~n4436 ;
  assign n4459 = ~n4401 & n4436 ;
  assign n4460 = ~n4458 & ~n4459 ;
  assign n4461 = n3651 & ~n4192 ;
  assign n4462 = ~n3651 & n4192 ;
  assign n4463 = ~n4461 & ~n4462 ;
  assign n4464 = n4324 & n4463 ;
  assign n4465 = ~n4324 & ~n4463 ;
  assign n4466 = ~n4464 & ~n4465 ;
  assign n4467 = n4274 & n4466 ;
  assign n4468 = ~n4274 & ~n4466 ;
  assign n4469 = ~n4467 & ~n4468 ;
  assign n4470 = n4020 & n4469 ;
  assign n4471 = ~n4020 & ~n4469 ;
  assign n4472 = ~n4470 & ~n4471 ;
  assign n4474 = ~n4460 & ~n4472 ;
  assign n4473 = n4460 & n4472 ;
  assign n4475 = decrypt_i_pad & ~n4473 ;
  assign n4476 = ~n4474 & n4475 ;
  assign n4477 = ~n4457 & ~n4476 ;
  assign n4478 = n4457 & n4476 ;
  assign n4479 = ~n4477 & ~n4478 ;
  assign n4480 = n3730 & ~n3995 ;
  assign n4481 = ~n3730 & n3995 ;
  assign n4482 = ~n4480 & ~n4481 ;
  assign n4483 = n4479 & n4482 ;
  assign n4484 = ~n4479 & ~n4482 ;
  assign n4485 = ~n4483 & ~n4484 ;
  assign n4486 = n3629 & ~n4485 ;
  assign n4487 = \mix1_data_reg_reg[109]/NET0131  & ~n3629 ;
  assign n4488 = ~n4486 & ~n4487 ;
  assign n4489 = ~n4120 & n4142 ;
  assign n4490 = n4120 & ~n4142 ;
  assign n4491 = ~n4489 & ~n4490 ;
  assign n4492 = n3777 & n4491 ;
  assign n4493 = ~n3777 & ~n4491 ;
  assign n4494 = ~n4492 & ~n4493 ;
  assign n4495 = n4064 & n4223 ;
  assign n4496 = ~n4064 & ~n4223 ;
  assign n4497 = ~n4495 & ~n4496 ;
  assign n4498 = n3890 & ~n4497 ;
  assign n4499 = ~n3890 & n4497 ;
  assign n4500 = ~n4498 & ~n4499 ;
  assign n4501 = n4494 & n4500 ;
  assign n4502 = ~n4494 & ~n4500 ;
  assign n4503 = ~n4501 & ~n4502 ;
  assign n4504 = n4293 & ~n4343 ;
  assign n4505 = ~n4293 & n4343 ;
  assign n4506 = ~n4504 & ~n4505 ;
  assign n4507 = n4312 & ~n4362 ;
  assign n4508 = ~n4312 & n4362 ;
  assign n4509 = ~n4507 & ~n4508 ;
  assign n4510 = n4506 & n4509 ;
  assign n4511 = ~n4506 & ~n4509 ;
  assign n4512 = ~n4510 & ~n4511 ;
  assign n4514 = n4503 & ~n4512 ;
  assign n4513 = ~n4503 & n4512 ;
  assign n4515 = decrypt_i_pad & ~n4513 ;
  assign n4516 = ~n4514 & n4515 ;
  assign n4517 = n4020 & ~n4436 ;
  assign n4518 = ~n4020 & n4436 ;
  assign n4519 = ~n4517 & ~n4518 ;
  assign n4520 = n4516 & n4519 ;
  assign n4521 = ~n4516 & ~n4519 ;
  assign n4522 = ~n4520 & ~n4521 ;
  assign n4523 = n4039 & n4248 ;
  assign n4524 = ~n4039 & ~n4248 ;
  assign n4525 = ~n4523 & ~n4524 ;
  assign n4526 = n4522 & n4525 ;
  assign n4527 = ~n4522 & ~n4525 ;
  assign n4528 = ~n4526 & ~n4527 ;
  assign n4529 = n3629 & ~n4528 ;
  assign n4530 = \mix1_data_reg_reg[115]/NET0131  & ~n3629 ;
  assign n4531 = ~n4529 & ~n4530 ;
  assign n4532 = ~n3998 & n4223 ;
  assign n4533 = n3998 & ~n4223 ;
  assign n4534 = ~n4532 & ~n4533 ;
  assign n4535 = ~n4101 & n4173 ;
  assign n4536 = n4101 & ~n4173 ;
  assign n4537 = ~n4535 & ~n4536 ;
  assign n4538 = n4436 & n4537 ;
  assign n4539 = ~n4436 & ~n4537 ;
  assign n4540 = ~n4538 & ~n4539 ;
  assign n4541 = n3938 & ~n4540 ;
  assign n4542 = ~n3938 & n4540 ;
  assign n4543 = ~n4541 & ~n4542 ;
  assign n4544 = n4534 & n4543 ;
  assign n4545 = ~n4534 & ~n4543 ;
  assign n4546 = ~n4544 & ~n4545 ;
  assign n4547 = n3629 & ~n4546 ;
  assign n4548 = ~\mix1_data_reg_reg[116]/NET0131  & ~n3629 ;
  assign n4549 = ~n4547 & ~n4548 ;
  assign n4550 = ~n3957 & ~n3995 ;
  assign n4551 = n3957 & n3995 ;
  assign n4552 = ~n4550 & ~n4551 ;
  assign n4553 = ~n4151 & ~n4173 ;
  assign n4554 = n4151 & n4173 ;
  assign n4555 = ~n4553 & ~n4554 ;
  assign n4556 = n4198 & n4525 ;
  assign n4557 = ~n4198 & ~n4525 ;
  assign n4558 = ~n4556 & ~n4557 ;
  assign n4560 = n4555 & n4558 ;
  assign n4559 = ~n4555 & ~n4558 ;
  assign n4561 = decrypt_i_pad & ~n4559 ;
  assign n4562 = ~n4560 & n4561 ;
  assign n4563 = ~n4552 & ~n4562 ;
  assign n4564 = n4552 & n4562 ;
  assign n4565 = ~n4563 & ~n4564 ;
  assign n4566 = n3730 & ~n4565 ;
  assign n4567 = ~n3730 & n4565 ;
  assign n4568 = ~n4566 & ~n4567 ;
  assign n4569 = n3774 & n4568 ;
  assign n4570 = ~n3774 & ~n4568 ;
  assign n4571 = ~n4569 & ~n4570 ;
  assign n4572 = n3629 & ~n4571 ;
  assign n4573 = \mix1_data_reg_reg[117]/NET0131  & ~n3629 ;
  assign n4574 = ~n4572 & ~n4573 ;
  assign n4575 = \mix1_data_reg_reg[123]/NET0131  & ~n3629 ;
  assign n4576 = n4381 & ~n4439 ;
  assign n4577 = ~n4381 & n4439 ;
  assign n4578 = ~n4576 & ~n4577 ;
  assign n4579 = n4466 & n4578 ;
  assign n4580 = ~n4466 & ~n4578 ;
  assign n4581 = ~n4579 & ~n4580 ;
  assign n4582 = n3629 & ~n4581 ;
  assign n4583 = ~n4575 & ~n4582 ;
  assign n4584 = n3957 & ~n4079 ;
  assign n4585 = ~n3957 & n4079 ;
  assign n4586 = ~n4584 & ~n4585 ;
  assign n4587 = ~n4020 & n4401 ;
  assign n4588 = n4020 & ~n4401 ;
  assign n4589 = ~n4587 & ~n4588 ;
  assign n4590 = n4436 & n4469 ;
  assign n4591 = ~n4436 & ~n4469 ;
  assign n4592 = ~n4590 & ~n4591 ;
  assign n4594 = n4589 & n4592 ;
  assign n4593 = ~n4589 & ~n4592 ;
  assign n4595 = decrypt_i_pad & ~n4593 ;
  assign n4596 = ~n4594 & n4595 ;
  assign n4597 = n4454 & ~n4596 ;
  assign n4598 = ~n4454 & n4596 ;
  assign n4599 = ~n4597 & ~n4598 ;
  assign n4600 = n4586 & n4599 ;
  assign n4601 = ~n4586 & ~n4599 ;
  assign n4602 = ~n4600 & ~n4601 ;
  assign n4603 = n3629 & ~n4602 ;
  assign n4604 = \mix1_data_reg_reg[125]/NET0131  & ~n3629 ;
  assign n4605 = ~n4603 & ~n4604 ;
  assign n4606 = n4020 & ~n4173 ;
  assign n4607 = ~n4020 & n4173 ;
  assign n4608 = ~n4606 & ~n4607 ;
  assign n4609 = ~n4324 & ~n4608 ;
  assign n4610 = n4324 & n4608 ;
  assign n4611 = ~n4609 & ~n4610 ;
  assign n4612 = n4552 & ~n4611 ;
  assign n4613 = ~n4552 & n4611 ;
  assign n4614 = ~n4612 & ~n4613 ;
  assign n4615 = n4414 & n4614 ;
  assign n4616 = ~n4414 & ~n4614 ;
  assign n4617 = ~n4615 & ~n4616 ;
  assign n4618 = n3629 & ~n4617 ;
  assign n4619 = ~\mix1_data_reg_reg[124]/NET0131  & ~n3629 ;
  assign n4620 = ~n4618 & ~n4619 ;
  assign n4621 = ~n4201 & ~n4522 ;
  assign n4622 = n4201 & n4522 ;
  assign n4623 = ~n4621 & ~n4622 ;
  assign n4624 = n3629 & n4623 ;
  assign n4625 = \mix1_data_reg_reg[99]/NET0131  & ~n3629 ;
  assign n4626 = ~n4624 & ~n4625 ;
  assign n4627 = ~n3730 & ~n3752 ;
  assign n4628 = n3730 & n3752 ;
  assign n4629 = ~n4627 & ~n4628 ;
  assign n4630 = n4142 & ~n4629 ;
  assign n4631 = ~n4142 & n4629 ;
  assign n4632 = ~n4630 & ~n4631 ;
  assign n4633 = n4067 & n4223 ;
  assign n4634 = ~n4067 & ~n4223 ;
  assign n4635 = ~n4633 & ~n4634 ;
  assign n4636 = n3957 & n4540 ;
  assign n4637 = ~n3957 & ~n4540 ;
  assign n4638 = ~n4636 & ~n4637 ;
  assign n4640 = n4635 & n4638 ;
  assign n4639 = ~n4635 & ~n4638 ;
  assign n4641 = decrypt_i_pad & ~n4639 ;
  assign n4642 = ~n4640 & n4641 ;
  assign n4643 = n3818 & ~n4642 ;
  assign n4644 = ~n3818 & n4642 ;
  assign n4645 = ~n4643 & ~n4644 ;
  assign n4646 = n4632 & n4645 ;
  assign n4647 = ~n4632 & ~n4645 ;
  assign n4648 = ~n4646 & ~n4647 ;
  assign n4649 = n3629 & ~n4648 ;
  assign n4650 = ~\mix1_data_reg_reg[102]/NET0131  & ~n3629 ;
  assign n4651 = ~n4649 & ~n4650 ;
  assign n4653 = ~n4001 & ~n4457 ;
  assign n4652 = n4001 & n4457 ;
  assign n4654 = decrypt_i_pad & ~n4652 ;
  assign n4655 = ~n4653 & n4654 ;
  assign n4656 = n4223 & ~n4398 ;
  assign n4657 = ~n4223 & n4398 ;
  assign n4658 = ~n4656 & ~n4657 ;
  assign n4659 = n4655 & n4658 ;
  assign n4660 = ~n4655 & ~n4658 ;
  assign n4661 = ~n4659 & ~n4660 ;
  assign n4662 = n3629 & n4661 ;
  assign n4663 = \mix1_data_reg_reg[103]/NET0131  & ~n3629 ;
  assign n4664 = ~n4662 & ~n4663 ;
  assign n4665 = decrypt_i_pad & n4404 ;
  assign n4666 = ~n3890 & n4665 ;
  assign n4667 = n3890 & ~n4665 ;
  assign n4668 = ~n4666 & ~n4667 ;
  assign n4669 = n3909 & ~n4668 ;
  assign n4670 = ~n3909 & n4668 ;
  assign n4671 = ~n4669 & ~n4670 ;
  assign n4672 = n4318 & n4671 ;
  assign n4673 = ~n4318 & ~n4671 ;
  assign n4674 = ~n4672 & ~n4673 ;
  assign n4675 = n3629 & ~n4674 ;
  assign n4676 = \mix1_data_reg_reg[105]/NET0131  & ~n3629 ;
  assign n4677 = ~n4675 & ~n4676 ;
  assign n4678 = ~n3843 & ~n3928 ;
  assign n4679 = n3843 & n3928 ;
  assign n4680 = ~n4678 & ~n4679 ;
  assign n4681 = n3868 & ~n4680 ;
  assign n4682 = ~n3868 & n4680 ;
  assign n4683 = ~n4681 & ~n4682 ;
  assign n4684 = ~n4223 & ~n4293 ;
  assign n4685 = n4223 & n4293 ;
  assign n4686 = ~n4684 & ~n4685 ;
  assign n4687 = ~n4064 & ~n4362 ;
  assign n4688 = n4064 & n4362 ;
  assign n4689 = ~n4687 & ~n4688 ;
  assign n4690 = ~n4686 & ~n4689 ;
  assign n4691 = n4686 & n4689 ;
  assign n4692 = ~n4690 & ~n4691 ;
  assign n4694 = n4401 & ~n4692 ;
  assign n4693 = ~n4401 & n4692 ;
  assign n4695 = decrypt_i_pad & ~n4693 ;
  assign n4696 = ~n4694 & n4695 ;
  assign n4697 = n4463 & ~n4696 ;
  assign n4698 = ~n4463 & n4696 ;
  assign n4699 = ~n4697 & ~n4698 ;
  assign n4700 = n4683 & n4699 ;
  assign n4701 = ~n4683 & ~n4699 ;
  assign n4702 = ~n4700 & ~n4701 ;
  assign n4703 = n3629 & ~n4702 ;
  assign n4704 = ~\mix1_data_reg_reg[106]/NET0131  & ~n3629 ;
  assign n4705 = ~n4703 & ~n4704 ;
  assign n4706 = ~n3815 & ~n4142 ;
  assign n4707 = n3815 & n4142 ;
  assign n4708 = ~n4706 & ~n4707 ;
  assign n4709 = n4439 & ~n4497 ;
  assign n4710 = ~n4439 & n4497 ;
  assign n4711 = ~n4709 & ~n4710 ;
  assign n4712 = n3998 & n4711 ;
  assign n4713 = ~n3998 & ~n4711 ;
  assign n4714 = ~n4712 & ~n4713 ;
  assign n4716 = n4608 & n4714 ;
  assign n4715 = ~n4608 & ~n4714 ;
  assign n4717 = decrypt_i_pad & ~n4715 ;
  assign n4718 = ~n4716 & n4717 ;
  assign n4719 = n4120 & ~n4718 ;
  assign n4720 = ~n4120 & n4718 ;
  assign n4721 = ~n4719 & ~n4720 ;
  assign n4722 = n3774 & ~n4721 ;
  assign n4723 = ~n3774 & n4721 ;
  assign n4724 = ~n4722 & ~n4723 ;
  assign n4725 = n4708 & n4724 ;
  assign n4726 = ~n4708 & ~n4724 ;
  assign n4727 = ~n4725 & ~n4726 ;
  assign n4728 = n3629 & n4727 ;
  assign n4729 = \mix1_data_reg_reg[110]/NET0131  & ~n3629 ;
  assign n4730 = ~n4728 & ~n4729 ;
  assign n4731 = n3771 & ~n4442 ;
  assign n4732 = ~n3771 & n4442 ;
  assign n4733 = ~n4731 & ~n4732 ;
  assign n4734 = n4482 & n4733 ;
  assign n4735 = ~n4482 & ~n4733 ;
  assign n4736 = ~n4734 & ~n4735 ;
  assign n4738 = ~n4101 & n4736 ;
  assign n4737 = n4101 & ~n4736 ;
  assign n4739 = decrypt_i_pad & ~n4737 ;
  assign n4740 = ~n4738 & n4739 ;
  assign n4741 = n3689 & ~n4740 ;
  assign n4742 = ~n3689 & n4740 ;
  assign n4743 = ~n4741 & ~n4742 ;
  assign n4744 = ~n4120 & ~n4743 ;
  assign n4745 = n4120 & n4743 ;
  assign n4746 = ~n4744 & ~n4745 ;
  assign n4747 = n3796 & ~n4746 ;
  assign n4748 = ~n3796 & n4746 ;
  assign n4749 = ~n4747 & ~n4748 ;
  assign n4750 = n4064 & n4749 ;
  assign n4751 = ~n4064 & ~n4749 ;
  assign n4752 = ~n4750 & ~n4751 ;
  assign n4753 = n3629 & ~n4752 ;
  assign n4754 = ~\mix1_data_reg_reg[111]/NET0131  & ~n3629 ;
  assign n4755 = ~n4753 & ~n4754 ;
  assign n4756 = decrypt_i_pad & n3824 ;
  assign n4757 = n3928 & ~n4756 ;
  assign n4758 = ~n3928 & n4756 ;
  assign n4759 = ~n4757 & ~n4758 ;
  assign n4760 = ~n3868 & n3909 ;
  assign n4761 = n3868 & ~n3909 ;
  assign n4762 = ~n4760 & ~n4761 ;
  assign n4763 = n4223 & ~n4762 ;
  assign n4764 = ~n4223 & n4762 ;
  assign n4765 = ~n4763 & ~n4764 ;
  assign n4766 = n4759 & ~n4765 ;
  assign n4767 = ~n4759 & n4765 ;
  assign n4768 = ~n4766 & ~n4767 ;
  assign n4769 = n4506 & n4768 ;
  assign n4770 = ~n4506 & ~n4768 ;
  assign n4771 = ~n4769 & ~n4770 ;
  assign n4772 = n3629 & ~n4771 ;
  assign n4773 = \mix1_data_reg_reg[113]/NET0131  & ~n3629 ;
  assign n4774 = ~n4772 & ~n4773 ;
  assign n4775 = \mix1_data_reg_reg[114]/NET0131  & ~n3629 ;
  assign n4776 = n3887 & ~n4680 ;
  assign n4777 = ~n3887 & n4680 ;
  assign n4778 = ~n4776 & ~n4777 ;
  assign n4779 = ~n4312 & n4343 ;
  assign n4780 = n4312 & ~n4343 ;
  assign n4781 = ~n4779 & ~n4780 ;
  assign n4782 = n4497 & n4781 ;
  assign n4783 = ~n4497 & ~n4781 ;
  assign n4784 = ~n4782 & ~n4783 ;
  assign n4786 = n4151 & n4784 ;
  assign n4785 = ~n4151 & ~n4784 ;
  assign n4787 = decrypt_i_pad & ~n4785 ;
  assign n4788 = ~n4786 & n4787 ;
  assign n4789 = n4392 & ~n4788 ;
  assign n4790 = ~n4392 & n4788 ;
  assign n4791 = ~n4789 & ~n4790 ;
  assign n4792 = n4778 & n4791 ;
  assign n4793 = ~n4778 & ~n4791 ;
  assign n4794 = ~n4792 & ~n4793 ;
  assign n4795 = n3629 & ~n4794 ;
  assign n4796 = ~n4775 & ~n4795 ;
  assign n4797 = ~n3771 & ~n3796 ;
  assign n4798 = n3771 & n3796 ;
  assign n4799 = ~n4797 & ~n4798 ;
  assign n4800 = n3711 & ~n4799 ;
  assign n4801 = ~n3711 & n4799 ;
  assign n4802 = ~n4800 & ~n4801 ;
  assign n4803 = n4123 & ~n4642 ;
  assign n4804 = ~n4123 & n4642 ;
  assign n4805 = ~n4803 & ~n4804 ;
  assign n4806 = n4802 & n4805 ;
  assign n4807 = ~n4802 & ~n4805 ;
  assign n4808 = ~n4806 & ~n4807 ;
  assign n4809 = n3629 & ~n4808 ;
  assign n4810 = ~\mix1_data_reg_reg[118]/NET0131  & ~n3629 ;
  assign n4811 = ~n4809 & ~n4810 ;
  assign n4812 = n4064 & ~n4395 ;
  assign n4813 = ~n4064 & n4395 ;
  assign n4814 = ~n4812 & ~n4813 ;
  assign n4815 = n4655 & n4814 ;
  assign n4816 = ~n4655 & ~n4814 ;
  assign n4817 = ~n4815 & ~n4816 ;
  assign n4818 = n3629 & ~n4817 ;
  assign n4819 = \mix1_data_reg_reg[119]/NET0131  & ~n3629 ;
  assign n4820 = ~n4818 & ~n4819 ;
  assign n4821 = n4371 & n4668 ;
  assign n4822 = ~n4371 & ~n4668 ;
  assign n4823 = ~n4821 & ~n4822 ;
  assign n4824 = n3629 & n4823 ;
  assign n4825 = \mix1_data_reg_reg[121]/NET0131  & ~n3629 ;
  assign n4826 = ~n4824 & ~n4825 ;
  assign n4827 = ~n3887 & n3909 ;
  assign n4828 = n3887 & ~n3909 ;
  assign n4829 = ~n4827 & ~n4828 ;
  assign n4830 = ~n4271 & n4696 ;
  assign n4831 = n4271 & ~n4696 ;
  assign n4832 = ~n4830 & ~n4831 ;
  assign n4833 = n3651 & ~n4832 ;
  assign n4834 = ~n3651 & n4832 ;
  assign n4835 = ~n4833 & ~n4834 ;
  assign n4836 = n4829 & n4835 ;
  assign n4837 = ~n4829 & ~n4835 ;
  assign n4838 = ~n4836 & ~n4837 ;
  assign n4839 = n3629 & n4838 ;
  assign n4840 = \mix1_data_reg_reg[122]/NET0131  & ~n3629 ;
  assign n4841 = ~n4839 & ~n4840 ;
  assign n4842 = n3733 & ~n4145 ;
  assign n4843 = ~n3733 & n4145 ;
  assign n4844 = ~n4842 & ~n4843 ;
  assign n4845 = n4721 & n4844 ;
  assign n4846 = ~n4721 & ~n4844 ;
  assign n4847 = ~n4845 & ~n4846 ;
  assign n4848 = n3629 & n4847 ;
  assign n4849 = \mix1_data_reg_reg[126]/NET0131  & ~n3629 ;
  assign n4850 = ~n4848 & ~n4849 ;
  assign n4851 = n4268 & ~n4743 ;
  assign n4852 = ~n4268 & n4743 ;
  assign n4853 = ~n4851 & ~n4852 ;
  assign n4854 = n4708 & n4853 ;
  assign n4855 = ~n4708 & ~n4853 ;
  assign n4856 = ~n4854 & ~n4855 ;
  assign n4857 = n3629 & n4856 ;
  assign n4858 = \mix1_data_reg_reg[127]/NET0131  & ~n3629 ;
  assign n4859 = ~n4857 & ~n4858 ;
  assign n4860 = n3635 & n4623 ;
  assign n4861 = \mix1_data_reg_reg[35]/NET0131  & ~n3635 ;
  assign n4862 = ~n4860 & ~n4861 ;
  assign n4863 = n3635 & ~n4073 ;
  assign n4864 = \mix1_data_reg_reg[36]/NET0131  & ~n3635 ;
  assign n4865 = ~n4863 & ~n4864 ;
  assign n4866 = n3635 & ~n4261 ;
  assign n4867 = \mix1_data_reg_reg[37]/NET0131  & ~n3635 ;
  assign n4868 = ~n4866 & ~n4867 ;
  assign n4869 = \mix1_data_reg_reg[43]/NET0131  & ~n3635 ;
  assign n4870 = n3635 & ~n4387 ;
  assign n4871 = ~n4869 & ~n4870 ;
  assign n4872 = n3635 & ~n4448 ;
  assign n4873 = \mix1_data_reg_reg[44]/NET0131  & ~n3635 ;
  assign n4874 = ~n4872 & ~n4873 ;
  assign n4875 = n3635 & ~n4485 ;
  assign n4876 = \mix1_data_reg_reg[45]/NET0131  & ~n3635 ;
  assign n4877 = ~n4875 & ~n4876 ;
  assign n4878 = n3635 & ~n4528 ;
  assign n4879 = \mix1_data_reg_reg[51]/NET0131  & ~n3635 ;
  assign n4880 = ~n4878 & ~n4879 ;
  assign n4881 = n3635 & ~n4571 ;
  assign n4882 = \mix1_data_reg_reg[53]/NET0131  & ~n3635 ;
  assign n4883 = ~n4881 & ~n4882 ;
  assign n4884 = n3635 & ~n4546 ;
  assign n4885 = ~\mix1_data_reg_reg[52]/NET0131  & ~n3635 ;
  assign n4886 = ~n4884 & ~n4885 ;
  assign n4887 = \mix1_data_reg_reg[59]/NET0131  & ~n3635 ;
  assign n4888 = n3635 & ~n4581 ;
  assign n4889 = ~n4887 & ~n4888 ;
  assign n4890 = n3635 & ~n4617 ;
  assign n4891 = ~\mix1_data_reg_reg[60]/NET0131  & ~n3635 ;
  assign n4892 = ~n4890 & ~n4891 ;
  assign n4893 = n3635 & ~n4602 ;
  assign n4894 = \mix1_data_reg_reg[61]/NET0131  & ~n3635 ;
  assign n4895 = ~n4893 & ~n4894 ;
  assign n4896 = n3630 & ~n4073 ;
  assign n4897 = \mix1_data_reg_reg[68]/NET0131  & ~n3630 ;
  assign n4898 = ~n4896 & ~n4897 ;
  assign n4899 = n3630 & ~n4261 ;
  assign n4900 = \mix1_data_reg_reg[69]/NET0131  & ~n3630 ;
  assign n4901 = ~n4899 & ~n4900 ;
  assign n4902 = n3630 & n4623 ;
  assign n4903 = \mix1_data_reg_reg[67]/NET0131  & ~n3630 ;
  assign n4904 = ~n4902 & ~n4903 ;
  assign n4905 = \mix1_data_reg_reg[75]/NET0131  & ~n3630 ;
  assign n4906 = n3630 & ~n4387 ;
  assign n4907 = ~n4905 & ~n4906 ;
  assign n4908 = n3630 & ~n4448 ;
  assign n4909 = \mix1_data_reg_reg[76]/NET0131  & ~n3630 ;
  assign n4910 = ~n4908 & ~n4909 ;
  assign n4911 = n3630 & ~n4485 ;
  assign n4912 = \mix1_data_reg_reg[77]/NET0131  & ~n3630 ;
  assign n4913 = ~n4911 & ~n4912 ;
  assign n4914 = n3630 & ~n4546 ;
  assign n4915 = ~\mix1_data_reg_reg[84]/NET0131  & ~n3630 ;
  assign n4916 = ~n4914 & ~n4915 ;
  assign n4917 = n3630 & ~n4571 ;
  assign n4918 = \mix1_data_reg_reg[85]/NET0131  & ~n3630 ;
  assign n4919 = ~n4917 & ~n4918 ;
  assign n4920 = n3630 & ~n4528 ;
  assign n4921 = \mix1_data_reg_reg[83]/NET0131  & ~n3630 ;
  assign n4922 = ~n4920 & ~n4921 ;
  assign n4923 = n3630 & ~n4617 ;
  assign n4924 = ~\mix1_data_reg_reg[92]/NET0131  & ~n3630 ;
  assign n4925 = ~n4923 & ~n4924 ;
  assign n4926 = \mix1_data_reg_reg[91]/NET0131  & ~n3630 ;
  assign n4927 = n3630 & ~n4581 ;
  assign n4928 = ~n4926 & ~n4927 ;
  assign n4929 = n3630 & ~n4602 ;
  assign n4930 = \mix1_data_reg_reg[93]/NET0131  & ~n3630 ;
  assign n4931 = ~n4929 & ~n4930 ;
  assign n4932 = ~n4245 & n4788 ;
  assign n4933 = n4245 & ~n4788 ;
  assign n4934 = ~n4932 & ~n4933 ;
  assign n4935 = n4192 & ~n4934 ;
  assign n4936 = ~n4192 & n4934 ;
  assign n4937 = ~n4935 & ~n4936 ;
  assign n4938 = n4762 & n4937 ;
  assign n4939 = ~n4762 & ~n4937 ;
  assign n4940 = ~n4938 & ~n4939 ;
  assign n4941 = n3629 & n4940 ;
  assign n4942 = \mix1_data_reg_reg[98]/NET0131  & ~n3629 ;
  assign n4943 = ~n4941 & ~n4942 ;
  assign n4944 = n4064 & ~n4829 ;
  assign n4945 = ~n4064 & n4829 ;
  assign n4946 = ~n4944 & ~n4945 ;
  assign n4947 = ~n4509 & n4759 ;
  assign n4948 = n4509 & ~n4759 ;
  assign n4949 = ~n4947 & ~n4948 ;
  assign n4950 = n4946 & n4949 ;
  assign n4951 = ~n4946 & ~n4949 ;
  assign n4952 = ~n4950 & ~n4951 ;
  assign n4953 = n3629 & ~n4952 ;
  assign n4954 = \mix1_data_reg_reg[97]/NET0131  & ~n3629 ;
  assign n4955 = ~n4953 & ~n4954 ;
  assign n4956 = \addroundkey_round_reg[3]/NET0131  & ~n949 ;
  assign n4957 = \addroundkey_round_reg[0]/NET0131  & \addroundkey_round_reg[1]/NET0131  ;
  assign n4958 = \addroundkey_round_reg[2]/NET0131  & n4957 ;
  assign n4959 = ~\addroundkey_round_reg[3]/NET0131  & ~n4958 ;
  assign n4960 = \addroundkey_round_reg[3]/NET0131  & n4958 ;
  assign n4961 = ~n4959 & ~n4960 ;
  assign n4962 = n949 & n4961 ;
  assign n4963 = ~n4956 & ~n4962 ;
  assign n4964 = ~\addroundkey_start_i_reg/NET0131  & ~n4963 ;
  assign n4965 = \addroundkey_round_reg[3]/NET0131  & n933 ;
  assign n4966 = ~n4964 & ~n4965 ;
  assign n4967 = \addroundkey_round_reg[1]/NET0131  & ~n949 ;
  assign n4968 = ~\addroundkey_round_reg[0]/NET0131  & ~\addroundkey_round_reg[1]/NET0131  ;
  assign n4969 = ~n4957 & ~n4968 ;
  assign n4970 = n949 & n4969 ;
  assign n4971 = ~n4967 & ~n4970 ;
  assign n4972 = ~\addroundkey_start_i_reg/NET0131  & ~n4971 ;
  assign n4973 = \addroundkey_round_reg[1]/NET0131  & n933 ;
  assign n4974 = ~n4972 & ~n4973 ;
  assign n4975 = \addroundkey_round_reg[0]/NET0131  & ~n968 ;
  assign n4976 = \addroundkey_round_reg[0]/NET0131  & ~n955 ;
  assign n4977 = ~n969 & ~n4976 ;
  assign n4978 = ~n4975 & ~n4977 ;
  assign n4979 = \addroundkey_round_reg[2]/NET0131  & ~n949 ;
  assign n4980 = ~\addroundkey_round_reg[2]/NET0131  & ~n4957 ;
  assign n4981 = ~n4958 & ~n4980 ;
  assign n4982 = n949 & n4981 ;
  assign n4983 = ~n4979 & ~n4982 ;
  assign n4984 = ~\addroundkey_start_i_reg/NET0131  & ~n4983 ;
  assign n4985 = \addroundkey_round_reg[2]/NET0131  & n933 ;
  assign n4986 = ~n4984 & ~n4985 ;
  assign n4993 = n4978 & n4986 ;
  assign n4994 = ~n4974 & n4993 ;
  assign n4995 = ~n4966 & n4994 ;
  assign n4987 = ~n4978 & n4986 ;
  assign n4988 = n4974 & n4987 ;
  assign n4989 = ~n4966 & n4988 ;
  assign n4990 = n4966 & ~n4986 ;
  assign n4991 = ~n4978 & n4990 ;
  assign n4992 = n4974 & n4991 ;
  assign n4996 = ~n4989 & ~n4992 ;
  assign n4997 = ~n4995 & n4996 ;
  assign n4998 = \ks1_col_reg[28]/NET0131  & ~n4997 ;
  assign n4999 = ~\ks1_col_reg[28]/NET0131  & n4997 ;
  assign n5000 = ~n4998 & ~n4999 ;
  assign n5001 = ~\ks1_key_reg_reg[124]/NET0131  & n1116 ;
  assign n5002 = ~\key_i[124]_pad  & ~n1116 ;
  assign n5003 = ~n5001 & ~n5002 ;
  assign n5004 = n5000 & ~n5003 ;
  assign n5005 = ~n5000 & n5003 ;
  assign n5006 = ~n5004 & ~n5005 ;
  assign n5007 = ~\ks1_key_reg_reg[92]/NET0131  & n1116 ;
  assign n5008 = ~\key_i[92]_pad  & ~n1116 ;
  assign n5009 = ~n5007 & ~n5008 ;
  assign n5010 = n5006 & ~n5009 ;
  assign n5011 = ~n5006 & n5009 ;
  assign n5012 = ~n5010 & ~n5011 ;
  assign n5013 = ~\ks1_key_reg_reg[60]/NET0131  & n1116 ;
  assign n5014 = ~\key_i[60]_pad  & ~n1116 ;
  assign n5015 = ~n5013 & ~n5014 ;
  assign n5016 = n5012 & ~n5015 ;
  assign n5017 = ~n5012 & n5015 ;
  assign n5018 = ~n5016 & ~n5017 ;
  assign n5019 = n929 & ~n5018 ;
  assign n5020 = \ks1_key_reg_reg[60]/NET0131  & ~n929 ;
  assign n5021 = ~n5019 & ~n5020 ;
  assign n5022 = n1305 & n5018 ;
  assign n5023 = ~n1305 & ~n5018 ;
  assign n5024 = ~n5022 & ~n5023 ;
  assign n5025 = \sub1_ready_o_reg/NET0131  & ~n3625 ;
  assign n5026 = n1261 & ~n5025 ;
  assign n5027 = ~decrypt_i_pad & \mix1_ready_o_reg/NET0131  ;
  assign n5028 = decrypt_i_pad & \sub1_ready_o_reg/NET0131  ;
  assign n5029 = ~decrypt_i_pad & ~n932 ;
  assign n5030 = ~\data_i[112]_pad  & ~n5029 ;
  assign n5031 = ~\mix1_data_o_reg_reg[112]/NET0131  & n5029 ;
  assign n5032 = ~n5030 & ~n5031 ;
  assign n5033 = ~n1159 & ~n5032 ;
  assign n5034 = ~\sub1_data_reg_reg[112]/NET0131  & n1159 ;
  assign n5035 = ~n5033 & ~n5034 ;
  assign n5036 = ~n5028 & ~n5035 ;
  assign n5037 = ~\sub1_data_reg_reg[112]/NET0131  & n5028 ;
  assign n5038 = ~n5036 & ~n5037 ;
  assign n5039 = ~n5027 & ~n5038 ;
  assign n5040 = ~\mix1_data_o_reg_reg[112]/NET0131  & n5027 ;
  assign n5041 = ~n5039 & ~n5040 ;
  assign n5042 = n5026 & ~n5041 ;
  assign n5043 = ~\sub1_data_reg_reg[112]/NET0131  & ~n5026 ;
  assign n5044 = ~n5042 & ~n5043 ;
  assign n5045 = \state_reg/NET0131  & ~n5044 ;
  assign n5046 = ~\state_reg/NET0131  & ~n5035 ;
  assign n5047 = ~n5045 & ~n5046 ;
  assign n5049 = \key_i[112]_pad  & n5047 ;
  assign n5048 = ~\key_i[112]_pad  & ~n5047 ;
  assign n5050 = n933 & ~n5048 ;
  assign n5051 = ~n5049 & n5050 ;
  assign n5052 = \ks1_ready_o_reg/NET0131  & ~n955 ;
  assign n5053 = n948 & n5052 ;
  assign n5055 = ~\ks1_key_reg_reg[112]/NET0131  & ~n5047 ;
  assign n5056 = \ks1_key_reg_reg[112]/NET0131  & n5047 ;
  assign n5057 = ~n5055 & ~n5056 ;
  assign n5058 = n5053 & ~n5057 ;
  assign n5054 = ~\data_o[112]_pad  & ~n5053 ;
  assign n5059 = ~n933 & ~n5054 ;
  assign n5060 = ~n5058 & n5059 ;
  assign n5061 = ~n5051 & ~n5060 ;
  assign n5062 = \data_i[61]_pad  & ~n5029 ;
  assign n5063 = \mix1_data_o_reg_reg[61]/NET0131  & n5029 ;
  assign n5064 = ~n5062 & ~n5063 ;
  assign n5065 = ~n1159 & ~n5064 ;
  assign n5066 = \sub1_data_reg_reg[61]/NET0131  & n1159 ;
  assign n5067 = ~n5065 & ~n5066 ;
  assign n5068 = ~n5028 & n5067 ;
  assign n5069 = ~\sub1_data_reg_reg[61]/NET0131  & n5028 ;
  assign n5070 = ~n5068 & ~n5069 ;
  assign n5071 = ~n5027 & ~n5070 ;
  assign n5072 = ~\mix1_data_o_reg_reg[61]/NET0131  & n5027 ;
  assign n5073 = ~n5071 & ~n5072 ;
  assign n5074 = n5026 & ~n5073 ;
  assign n5075 = ~\sub1_data_reg_reg[61]/NET0131  & ~n5026 ;
  assign n5076 = ~n5074 & ~n5075 ;
  assign n5077 = \state_reg/NET0131  & ~n5076 ;
  assign n5078 = ~\state_reg/NET0131  & n5067 ;
  assign n5079 = ~n5077 & ~n5078 ;
  assign n5081 = \key_i[61]_pad  & n5079 ;
  assign n5080 = ~\key_i[61]_pad  & ~n5079 ;
  assign n5082 = n933 & ~n5080 ;
  assign n5083 = ~n5081 & n5082 ;
  assign n5085 = ~\ks1_key_reg_reg[61]/NET0131  & ~n5079 ;
  assign n5086 = \ks1_key_reg_reg[61]/NET0131  & n5079 ;
  assign n5087 = ~n5085 & ~n5086 ;
  assign n5088 = n5053 & ~n5087 ;
  assign n5084 = ~\data_o[61]_pad  & ~n5053 ;
  assign n5089 = ~n933 & ~n5084 ;
  assign n5090 = ~n5088 & n5089 ;
  assign n5091 = ~n5083 & ~n5090 ;
  assign n5092 = ~\data_i[19]_pad  & ~n5029 ;
  assign n5093 = ~\mix1_data_o_reg_reg[19]/NET0131  & n5029 ;
  assign n5094 = ~n5092 & ~n5093 ;
  assign n5095 = ~n1159 & ~n5094 ;
  assign n5096 = ~\sub1_data_reg_reg[19]/NET0131  & n1159 ;
  assign n5097 = ~n5095 & ~n5096 ;
  assign n5098 = ~n5028 & ~n5097 ;
  assign n5099 = ~\sub1_data_reg_reg[19]/NET0131  & n5028 ;
  assign n5100 = ~n5098 & ~n5099 ;
  assign n5101 = ~n5027 & ~n5100 ;
  assign n5102 = ~\mix1_data_o_reg_reg[19]/NET0131  & n5027 ;
  assign n5103 = ~n5101 & ~n5102 ;
  assign n5104 = n5026 & ~n5103 ;
  assign n5105 = ~\sub1_data_reg_reg[19]/NET0131  & ~n5026 ;
  assign n5106 = ~n5104 & ~n5105 ;
  assign n5107 = \state_reg/NET0131  & ~n5106 ;
  assign n5108 = ~\state_reg/NET0131  & ~n5097 ;
  assign n5109 = ~n5107 & ~n5108 ;
  assign n5111 = \key_i[19]_pad  & n5109 ;
  assign n5110 = ~\key_i[19]_pad  & ~n5109 ;
  assign n5112 = n933 & ~n5110 ;
  assign n5113 = ~n5111 & n5112 ;
  assign n5115 = ~\ks1_key_reg_reg[19]/NET0131  & ~n5109 ;
  assign n5116 = \ks1_key_reg_reg[19]/NET0131  & n5109 ;
  assign n5117 = ~n5115 & ~n5116 ;
  assign n5118 = n5053 & ~n5117 ;
  assign n5114 = ~\data_o[19]_pad  & ~n5053 ;
  assign n5119 = ~n933 & ~n5114 ;
  assign n5120 = ~n5118 & n5119 ;
  assign n5121 = ~n5113 & ~n5120 ;
  assign n5122 = \data_i[62]_pad  & ~n5029 ;
  assign n5123 = \mix1_data_o_reg_reg[62]/NET0131  & n5029 ;
  assign n5124 = ~n5122 & ~n5123 ;
  assign n5125 = ~n1159 & ~n5124 ;
  assign n5126 = \sub1_data_reg_reg[62]/NET0131  & n1159 ;
  assign n5127 = ~n5125 & ~n5126 ;
  assign n5128 = ~n5028 & n5127 ;
  assign n5129 = ~\sub1_data_reg_reg[62]/NET0131  & n5028 ;
  assign n5130 = ~n5128 & ~n5129 ;
  assign n5131 = ~n5027 & ~n5130 ;
  assign n5132 = ~\mix1_data_o_reg_reg[62]/NET0131  & n5027 ;
  assign n5133 = ~n5131 & ~n5132 ;
  assign n5134 = n5026 & ~n5133 ;
  assign n5135 = ~\sub1_data_reg_reg[62]/NET0131  & ~n5026 ;
  assign n5136 = ~n5134 & ~n5135 ;
  assign n5137 = \state_reg/NET0131  & ~n5136 ;
  assign n5138 = ~\state_reg/NET0131  & n5127 ;
  assign n5139 = ~n5137 & ~n5138 ;
  assign n5141 = \key_i[62]_pad  & n5139 ;
  assign n5140 = ~\key_i[62]_pad  & ~n5139 ;
  assign n5142 = n933 & ~n5140 ;
  assign n5143 = ~n5141 & n5142 ;
  assign n5145 = ~\ks1_key_reg_reg[62]/NET0131  & ~n5139 ;
  assign n5146 = \ks1_key_reg_reg[62]/NET0131  & n5139 ;
  assign n5147 = ~n5145 & ~n5146 ;
  assign n5148 = n5053 & ~n5147 ;
  assign n5144 = ~\data_o[62]_pad  & ~n5053 ;
  assign n5149 = ~n933 & ~n5144 ;
  assign n5150 = ~n5148 & n5149 ;
  assign n5151 = ~n5143 & ~n5150 ;
  assign n5152 = \data_i[63]_pad  & ~n5029 ;
  assign n5153 = \mix1_data_o_reg_reg[63]/NET0131  & n5029 ;
  assign n5154 = ~n5152 & ~n5153 ;
  assign n5155 = ~n1159 & ~n5154 ;
  assign n5156 = \sub1_data_reg_reg[63]/NET0131  & n1159 ;
  assign n5157 = ~n5155 & ~n5156 ;
  assign n5158 = ~n5028 & n5157 ;
  assign n5159 = ~\sub1_data_reg_reg[63]/NET0131  & n5028 ;
  assign n5160 = ~n5158 & ~n5159 ;
  assign n5161 = ~n5027 & ~n5160 ;
  assign n5162 = ~\mix1_data_o_reg_reg[63]/NET0131  & n5027 ;
  assign n5163 = ~n5161 & ~n5162 ;
  assign n5164 = n5026 & ~n5163 ;
  assign n5165 = ~\sub1_data_reg_reg[63]/NET0131  & ~n5026 ;
  assign n5166 = ~n5164 & ~n5165 ;
  assign n5167 = \state_reg/NET0131  & ~n5166 ;
  assign n5168 = ~\state_reg/NET0131  & n5157 ;
  assign n5169 = ~n5167 & ~n5168 ;
  assign n5171 = \key_i[63]_pad  & n5169 ;
  assign n5170 = ~\key_i[63]_pad  & ~n5169 ;
  assign n5172 = n933 & ~n5170 ;
  assign n5173 = ~n5171 & n5172 ;
  assign n5175 = ~\ks1_key_reg_reg[63]/NET0131  & ~n5169 ;
  assign n5176 = \ks1_key_reg_reg[63]/NET0131  & n5169 ;
  assign n5177 = ~n5175 & ~n5176 ;
  assign n5178 = n5053 & ~n5177 ;
  assign n5174 = ~\data_o[63]_pad  & ~n5053 ;
  assign n5179 = ~n933 & ~n5174 ;
  assign n5180 = ~n5178 & n5179 ;
  assign n5181 = ~n5173 & ~n5180 ;
  assign n5182 = \data_i[1]_pad  & ~n5029 ;
  assign n5183 = \mix1_data_o_reg_reg[1]/NET0131  & n5029 ;
  assign n5184 = ~n5182 & ~n5183 ;
  assign n5185 = ~n1159 & ~n5184 ;
  assign n5186 = \sub1_data_reg_reg[1]/NET0131  & n1159 ;
  assign n5187 = ~n5185 & ~n5186 ;
  assign n5188 = ~n5028 & n5187 ;
  assign n5189 = ~\sub1_data_reg_reg[1]/NET0131  & n5028 ;
  assign n5190 = ~n5188 & ~n5189 ;
  assign n5191 = ~n5027 & ~n5190 ;
  assign n5192 = ~\mix1_data_o_reg_reg[1]/NET0131  & n5027 ;
  assign n5193 = ~n5191 & ~n5192 ;
  assign n5194 = n5026 & ~n5193 ;
  assign n5195 = ~\sub1_data_reg_reg[1]/NET0131  & ~n5026 ;
  assign n5196 = ~n5194 & ~n5195 ;
  assign n5197 = \state_reg/NET0131  & ~n5196 ;
  assign n5198 = ~\state_reg/NET0131  & n5187 ;
  assign n5199 = ~n5197 & ~n5198 ;
  assign n5201 = \key_i[1]_pad  & n5199 ;
  assign n5200 = ~\key_i[1]_pad  & ~n5199 ;
  assign n5202 = n933 & ~n5200 ;
  assign n5203 = ~n5201 & n5202 ;
  assign n5205 = ~\ks1_key_reg_reg[1]/NET0131  & ~n5199 ;
  assign n5206 = \ks1_key_reg_reg[1]/NET0131  & n5199 ;
  assign n5207 = ~n5205 & ~n5206 ;
  assign n5208 = n5053 & ~n5207 ;
  assign n5204 = ~\data_o[1]_pad  & ~n5053 ;
  assign n5209 = ~n933 & ~n5204 ;
  assign n5210 = ~n5208 & n5209 ;
  assign n5211 = ~n5203 & ~n5210 ;
  assign n5212 = ~\data_i[64]_pad  & ~n5029 ;
  assign n5213 = ~\mix1_data_o_reg_reg[64]/NET0131  & n5029 ;
  assign n5214 = ~n5212 & ~n5213 ;
  assign n5215 = ~n1159 & ~n5214 ;
  assign n5216 = ~\sub1_data_reg_reg[64]/NET0131  & n1159 ;
  assign n5217 = ~n5215 & ~n5216 ;
  assign n5218 = ~n5028 & ~n5217 ;
  assign n5219 = ~\sub1_data_reg_reg[64]/NET0131  & n5028 ;
  assign n5220 = ~n5218 & ~n5219 ;
  assign n5221 = ~n5027 & ~n5220 ;
  assign n5222 = ~\mix1_data_o_reg_reg[64]/NET0131  & n5027 ;
  assign n5223 = ~n5221 & ~n5222 ;
  assign n5224 = n5026 & ~n5223 ;
  assign n5225 = ~\sub1_data_reg_reg[64]/NET0131  & ~n5026 ;
  assign n5226 = ~n5224 & ~n5225 ;
  assign n5227 = \state_reg/NET0131  & ~n5226 ;
  assign n5228 = ~\state_reg/NET0131  & ~n5217 ;
  assign n5229 = ~n5227 & ~n5228 ;
  assign n5231 = \key_i[64]_pad  & n5229 ;
  assign n5230 = ~\key_i[64]_pad  & ~n5229 ;
  assign n5232 = n933 & ~n5230 ;
  assign n5233 = ~n5231 & n5232 ;
  assign n5235 = ~\ks1_key_reg_reg[64]/NET0131  & ~n5229 ;
  assign n5236 = \ks1_key_reg_reg[64]/NET0131  & n5229 ;
  assign n5237 = ~n5235 & ~n5236 ;
  assign n5238 = n5053 & ~n5237 ;
  assign n5234 = ~\data_o[64]_pad  & ~n5053 ;
  assign n5239 = ~n933 & ~n5234 ;
  assign n5240 = ~n5238 & n5239 ;
  assign n5241 = ~n5233 & ~n5240 ;
  assign n5242 = ~\data_i[101]_pad  & ~n5029 ;
  assign n5243 = ~\mix1_data_o_reg_reg[101]/NET0131  & n5029 ;
  assign n5244 = ~n5242 & ~n5243 ;
  assign n5245 = ~n1159 & ~n5244 ;
  assign n5246 = ~\sub1_data_reg_reg[101]/NET0131  & n1159 ;
  assign n5247 = ~n5245 & ~n5246 ;
  assign n5248 = ~n5028 & ~n5247 ;
  assign n5249 = ~\sub1_data_reg_reg[101]/NET0131  & n5028 ;
  assign n5250 = ~n5248 & ~n5249 ;
  assign n5251 = ~n5027 & ~n5250 ;
  assign n5252 = ~\mix1_data_o_reg_reg[101]/NET0131  & n5027 ;
  assign n5253 = ~n5251 & ~n5252 ;
  assign n5254 = n5026 & ~n5253 ;
  assign n5255 = ~\sub1_data_reg_reg[101]/NET0131  & ~n5026 ;
  assign n5256 = ~n5254 & ~n5255 ;
  assign n5257 = \state_reg/NET0131  & ~n5256 ;
  assign n5258 = ~\state_reg/NET0131  & ~n5247 ;
  assign n5259 = ~n5257 & ~n5258 ;
  assign n5261 = \key_i[101]_pad  & n5259 ;
  assign n5260 = ~\key_i[101]_pad  & ~n5259 ;
  assign n5262 = n933 & ~n5260 ;
  assign n5263 = ~n5261 & n5262 ;
  assign n5265 = ~\ks1_key_reg_reg[101]/NET0131  & ~n5259 ;
  assign n5266 = \ks1_key_reg_reg[101]/NET0131  & n5259 ;
  assign n5267 = ~n5265 & ~n5266 ;
  assign n5268 = n5053 & ~n5267 ;
  assign n5264 = ~\data_o[101]_pad  & ~n5053 ;
  assign n5269 = ~n933 & ~n5264 ;
  assign n5270 = ~n5268 & n5269 ;
  assign n5271 = ~n5263 & ~n5270 ;
  assign n5272 = ~\data_i[65]_pad  & ~n5029 ;
  assign n5273 = ~\mix1_data_o_reg_reg[65]/NET0131  & n5029 ;
  assign n5274 = ~n5272 & ~n5273 ;
  assign n5275 = ~n1159 & ~n5274 ;
  assign n5276 = ~\sub1_data_reg_reg[65]/NET0131  & n1159 ;
  assign n5277 = ~n5275 & ~n5276 ;
  assign n5278 = ~n5028 & ~n5277 ;
  assign n5279 = ~\sub1_data_reg_reg[65]/NET0131  & n5028 ;
  assign n5280 = ~n5278 & ~n5279 ;
  assign n5281 = ~n5027 & ~n5280 ;
  assign n5282 = ~\mix1_data_o_reg_reg[65]/NET0131  & n5027 ;
  assign n5283 = ~n5281 & ~n5282 ;
  assign n5284 = n5026 & ~n5283 ;
  assign n5285 = ~\sub1_data_reg_reg[65]/NET0131  & ~n5026 ;
  assign n5286 = ~n5284 & ~n5285 ;
  assign n5287 = \state_reg/NET0131  & ~n5286 ;
  assign n5288 = ~\state_reg/NET0131  & ~n5277 ;
  assign n5289 = ~n5287 & ~n5288 ;
  assign n5291 = \key_i[65]_pad  & n5289 ;
  assign n5290 = ~\key_i[65]_pad  & ~n5289 ;
  assign n5292 = n933 & ~n5290 ;
  assign n5293 = ~n5291 & n5292 ;
  assign n5295 = ~\ks1_key_reg_reg[65]/NET0131  & ~n5289 ;
  assign n5296 = \ks1_key_reg_reg[65]/NET0131  & n5289 ;
  assign n5297 = ~n5295 & ~n5296 ;
  assign n5298 = n5053 & ~n5297 ;
  assign n5294 = ~\data_o[65]_pad  & ~n5053 ;
  assign n5299 = ~n933 & ~n5294 ;
  assign n5300 = ~n5298 & n5299 ;
  assign n5301 = ~n5293 & ~n5300 ;
  assign n5302 = ~\data_i[66]_pad  & ~n5029 ;
  assign n5303 = ~\mix1_data_o_reg_reg[66]/NET0131  & n5029 ;
  assign n5304 = ~n5302 & ~n5303 ;
  assign n5305 = ~n1159 & ~n5304 ;
  assign n5306 = ~\sub1_data_reg_reg[66]/NET0131  & n1159 ;
  assign n5307 = ~n5305 & ~n5306 ;
  assign n5308 = ~n5028 & ~n5307 ;
  assign n5309 = ~\sub1_data_reg_reg[66]/NET0131  & n5028 ;
  assign n5310 = ~n5308 & ~n5309 ;
  assign n5311 = ~n5027 & ~n5310 ;
  assign n5312 = ~\mix1_data_o_reg_reg[66]/NET0131  & n5027 ;
  assign n5313 = ~n5311 & ~n5312 ;
  assign n5314 = n5026 & ~n5313 ;
  assign n5315 = ~\sub1_data_reg_reg[66]/NET0131  & ~n5026 ;
  assign n5316 = ~n5314 & ~n5315 ;
  assign n5317 = \state_reg/NET0131  & ~n5316 ;
  assign n5318 = ~\state_reg/NET0131  & ~n5307 ;
  assign n5319 = ~n5317 & ~n5318 ;
  assign n5321 = \key_i[66]_pad  & n5319 ;
  assign n5320 = ~\key_i[66]_pad  & ~n5319 ;
  assign n5322 = n933 & ~n5320 ;
  assign n5323 = ~n5321 & n5322 ;
  assign n5325 = ~\ks1_key_reg_reg[66]/NET0131  & ~n5319 ;
  assign n5326 = \ks1_key_reg_reg[66]/NET0131  & n5319 ;
  assign n5327 = ~n5325 & ~n5326 ;
  assign n5328 = n5053 & ~n5327 ;
  assign n5324 = ~\data_o[66]_pad  & ~n5053 ;
  assign n5329 = ~n933 & ~n5324 ;
  assign n5330 = ~n5328 & n5329 ;
  assign n5331 = ~n5323 & ~n5330 ;
  assign n5332 = ~\data_i[20]_pad  & ~n5029 ;
  assign n5333 = ~\mix1_data_o_reg_reg[20]/NET0131  & n5029 ;
  assign n5334 = ~n5332 & ~n5333 ;
  assign n5335 = ~n1159 & ~n5334 ;
  assign n5336 = ~\sub1_data_reg_reg[20]/NET0131  & n1159 ;
  assign n5337 = ~n5335 & ~n5336 ;
  assign n5338 = ~n5028 & ~n5337 ;
  assign n5339 = ~\sub1_data_reg_reg[20]/NET0131  & n5028 ;
  assign n5340 = ~n5338 & ~n5339 ;
  assign n5341 = ~n5027 & ~n5340 ;
  assign n5342 = ~\mix1_data_o_reg_reg[20]/NET0131  & n5027 ;
  assign n5343 = ~n5341 & ~n5342 ;
  assign n5344 = n5026 & ~n5343 ;
  assign n5345 = ~\sub1_data_reg_reg[20]/NET0131  & ~n5026 ;
  assign n5346 = ~n5344 & ~n5345 ;
  assign n5347 = \state_reg/NET0131  & ~n5346 ;
  assign n5348 = ~\state_reg/NET0131  & ~n5337 ;
  assign n5349 = ~n5347 & ~n5348 ;
  assign n5351 = \key_i[20]_pad  & n5349 ;
  assign n5350 = ~\key_i[20]_pad  & ~n5349 ;
  assign n5352 = n933 & ~n5350 ;
  assign n5353 = ~n5351 & n5352 ;
  assign n5355 = ~\ks1_key_reg_reg[20]/NET0131  & ~n5349 ;
  assign n5356 = \ks1_key_reg_reg[20]/NET0131  & n5349 ;
  assign n5357 = ~n5355 & ~n5356 ;
  assign n5358 = n5053 & ~n5357 ;
  assign n5354 = ~\data_o[20]_pad  & ~n5053 ;
  assign n5359 = ~n933 & ~n5354 ;
  assign n5360 = ~n5358 & n5359 ;
  assign n5361 = ~n5353 & ~n5360 ;
  assign n5362 = ~\data_i[67]_pad  & ~n5029 ;
  assign n5363 = ~\mix1_data_o_reg_reg[67]/NET0131  & n5029 ;
  assign n5364 = ~n5362 & ~n5363 ;
  assign n5365 = ~n1159 & ~n5364 ;
  assign n5366 = ~\sub1_data_reg_reg[67]/NET0131  & n1159 ;
  assign n5367 = ~n5365 & ~n5366 ;
  assign n5368 = ~n5028 & ~n5367 ;
  assign n5369 = ~\sub1_data_reg_reg[67]/NET0131  & n5028 ;
  assign n5370 = ~n5368 & ~n5369 ;
  assign n5371 = ~n5027 & ~n5370 ;
  assign n5372 = ~\mix1_data_o_reg_reg[67]/NET0131  & n5027 ;
  assign n5373 = ~n5371 & ~n5372 ;
  assign n5374 = n5026 & ~n5373 ;
  assign n5375 = ~\sub1_data_reg_reg[67]/NET0131  & ~n5026 ;
  assign n5376 = ~n5374 & ~n5375 ;
  assign n5377 = \state_reg/NET0131  & ~n5376 ;
  assign n5378 = ~\state_reg/NET0131  & ~n5367 ;
  assign n5379 = ~n5377 & ~n5378 ;
  assign n5381 = \key_i[67]_pad  & n5379 ;
  assign n5380 = ~\key_i[67]_pad  & ~n5379 ;
  assign n5382 = n933 & ~n5380 ;
  assign n5383 = ~n5381 & n5382 ;
  assign n5385 = ~\ks1_key_reg_reg[67]/NET0131  & ~n5379 ;
  assign n5386 = \ks1_key_reg_reg[67]/NET0131  & n5379 ;
  assign n5387 = ~n5385 & ~n5386 ;
  assign n5388 = n5053 & ~n5387 ;
  assign n5384 = ~\data_o[67]_pad  & ~n5053 ;
  assign n5389 = ~n933 & ~n5384 ;
  assign n5390 = ~n5388 & n5389 ;
  assign n5391 = ~n5383 & ~n5390 ;
  assign n5392 = ~\data_i[113]_pad  & ~n5029 ;
  assign n5393 = ~\mix1_data_o_reg_reg[113]/NET0131  & n5029 ;
  assign n5394 = ~n5392 & ~n5393 ;
  assign n5395 = ~n1159 & ~n5394 ;
  assign n5396 = ~\sub1_data_reg_reg[113]/NET0131  & n1159 ;
  assign n5397 = ~n5395 & ~n5396 ;
  assign n5398 = ~n5028 & ~n5397 ;
  assign n5399 = ~\sub1_data_reg_reg[113]/NET0131  & n5028 ;
  assign n5400 = ~n5398 & ~n5399 ;
  assign n5401 = ~n5027 & ~n5400 ;
  assign n5402 = ~\mix1_data_o_reg_reg[113]/NET0131  & n5027 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = n5026 & ~n5403 ;
  assign n5405 = ~\sub1_data_reg_reg[113]/NET0131  & ~n5026 ;
  assign n5406 = ~n5404 & ~n5405 ;
  assign n5407 = \state_reg/NET0131  & ~n5406 ;
  assign n5408 = ~\state_reg/NET0131  & ~n5397 ;
  assign n5409 = ~n5407 & ~n5408 ;
  assign n5411 = \key_i[113]_pad  & n5409 ;
  assign n5410 = ~\key_i[113]_pad  & ~n5409 ;
  assign n5412 = n933 & ~n5410 ;
  assign n5413 = ~n5411 & n5412 ;
  assign n5415 = ~\ks1_key_reg_reg[113]/NET0131  & ~n5409 ;
  assign n5416 = \ks1_key_reg_reg[113]/NET0131  & n5409 ;
  assign n5417 = ~n5415 & ~n5416 ;
  assign n5418 = n5053 & ~n5417 ;
  assign n5414 = ~\data_o[113]_pad  & ~n5053 ;
  assign n5419 = ~n933 & ~n5414 ;
  assign n5420 = ~n5418 & n5419 ;
  assign n5421 = ~n5413 & ~n5420 ;
  assign n5422 = ~\data_i[21]_pad  & ~n5029 ;
  assign n5423 = ~\mix1_data_o_reg_reg[21]/NET0131  & n5029 ;
  assign n5424 = ~n5422 & ~n5423 ;
  assign n5425 = ~n1159 & ~n5424 ;
  assign n5426 = ~\sub1_data_reg_reg[21]/NET0131  & n1159 ;
  assign n5427 = ~n5425 & ~n5426 ;
  assign n5428 = ~n5028 & ~n5427 ;
  assign n5429 = ~\sub1_data_reg_reg[21]/NET0131  & n5028 ;
  assign n5430 = ~n5428 & ~n5429 ;
  assign n5431 = ~n5027 & ~n5430 ;
  assign n5432 = ~\mix1_data_o_reg_reg[21]/NET0131  & n5027 ;
  assign n5433 = ~n5431 & ~n5432 ;
  assign n5434 = n5026 & ~n5433 ;
  assign n5435 = ~\sub1_data_reg_reg[21]/NET0131  & ~n5026 ;
  assign n5436 = ~n5434 & ~n5435 ;
  assign n5437 = \state_reg/NET0131  & ~n5436 ;
  assign n5438 = ~\state_reg/NET0131  & ~n5427 ;
  assign n5439 = ~n5437 & ~n5438 ;
  assign n5441 = \key_i[21]_pad  & n5439 ;
  assign n5440 = ~\key_i[21]_pad  & ~n5439 ;
  assign n5442 = n933 & ~n5440 ;
  assign n5443 = ~n5441 & n5442 ;
  assign n5445 = ~\ks1_key_reg_reg[21]/NET0131  & ~n5439 ;
  assign n5446 = \ks1_key_reg_reg[21]/NET0131  & n5439 ;
  assign n5447 = ~n5445 & ~n5446 ;
  assign n5448 = n5053 & ~n5447 ;
  assign n5444 = ~\data_o[21]_pad  & ~n5053 ;
  assign n5449 = ~n933 & ~n5444 ;
  assign n5450 = ~n5448 & n5449 ;
  assign n5451 = ~n5443 & ~n5450 ;
  assign n5452 = ~\data_i[68]_pad  & ~n5029 ;
  assign n5453 = ~\mix1_data_o_reg_reg[68]/NET0131  & n5029 ;
  assign n5454 = ~n5452 & ~n5453 ;
  assign n5455 = ~n1159 & ~n5454 ;
  assign n5456 = ~\sub1_data_reg_reg[68]/NET0131  & n1159 ;
  assign n5457 = ~n5455 & ~n5456 ;
  assign n5458 = ~n5028 & ~n5457 ;
  assign n5459 = ~\sub1_data_reg_reg[68]/NET0131  & n5028 ;
  assign n5460 = ~n5458 & ~n5459 ;
  assign n5461 = ~n5027 & ~n5460 ;
  assign n5462 = ~\mix1_data_o_reg_reg[68]/NET0131  & n5027 ;
  assign n5463 = ~n5461 & ~n5462 ;
  assign n5464 = n5026 & ~n5463 ;
  assign n5465 = ~\sub1_data_reg_reg[68]/NET0131  & ~n5026 ;
  assign n5466 = ~n5464 & ~n5465 ;
  assign n5467 = \state_reg/NET0131  & ~n5466 ;
  assign n5468 = ~\state_reg/NET0131  & ~n5457 ;
  assign n5469 = ~n5467 & ~n5468 ;
  assign n5471 = \key_i[68]_pad  & n5469 ;
  assign n5470 = ~\key_i[68]_pad  & ~n5469 ;
  assign n5472 = n933 & ~n5470 ;
  assign n5473 = ~n5471 & n5472 ;
  assign n5475 = ~\ks1_key_reg_reg[68]/NET0131  & ~n5469 ;
  assign n5476 = \ks1_key_reg_reg[68]/NET0131  & n5469 ;
  assign n5477 = ~n5475 & ~n5476 ;
  assign n5478 = n5053 & ~n5477 ;
  assign n5474 = ~\data_o[68]_pad  & ~n5053 ;
  assign n5479 = ~n933 & ~n5474 ;
  assign n5480 = ~n5478 & n5479 ;
  assign n5481 = ~n5473 & ~n5480 ;
  assign n5482 = ~\data_i[69]_pad  & ~n5029 ;
  assign n5483 = ~\mix1_data_o_reg_reg[69]/NET0131  & n5029 ;
  assign n5484 = ~n5482 & ~n5483 ;
  assign n5485 = ~n1159 & ~n5484 ;
  assign n5486 = ~\sub1_data_reg_reg[69]/NET0131  & n1159 ;
  assign n5487 = ~n5485 & ~n5486 ;
  assign n5488 = ~n5028 & ~n5487 ;
  assign n5489 = ~\sub1_data_reg_reg[69]/NET0131  & n5028 ;
  assign n5490 = ~n5488 & ~n5489 ;
  assign n5491 = ~n5027 & ~n5490 ;
  assign n5492 = ~\mix1_data_o_reg_reg[69]/NET0131  & n5027 ;
  assign n5493 = ~n5491 & ~n5492 ;
  assign n5494 = n5026 & ~n5493 ;
  assign n5495 = ~\sub1_data_reg_reg[69]/NET0131  & ~n5026 ;
  assign n5496 = ~n5494 & ~n5495 ;
  assign n5497 = \state_reg/NET0131  & ~n5496 ;
  assign n5498 = ~\state_reg/NET0131  & ~n5487 ;
  assign n5499 = ~n5497 & ~n5498 ;
  assign n5501 = \key_i[69]_pad  & n5499 ;
  assign n5500 = ~\key_i[69]_pad  & ~n5499 ;
  assign n5502 = n933 & ~n5500 ;
  assign n5503 = ~n5501 & n5502 ;
  assign n5505 = ~\ks1_key_reg_reg[69]/NET0131  & ~n5499 ;
  assign n5506 = \ks1_key_reg_reg[69]/NET0131  & n5499 ;
  assign n5507 = ~n5505 & ~n5506 ;
  assign n5508 = n5053 & ~n5507 ;
  assign n5504 = ~\data_o[69]_pad  & ~n5053 ;
  assign n5509 = ~n933 & ~n5504 ;
  assign n5510 = ~n5508 & n5509 ;
  assign n5511 = ~n5503 & ~n5510 ;
  assign n5512 = ~\data_i[102]_pad  & ~n5029 ;
  assign n5513 = ~\mix1_data_o_reg_reg[102]/NET0131  & n5029 ;
  assign n5514 = ~n5512 & ~n5513 ;
  assign n5515 = ~n1159 & ~n5514 ;
  assign n5516 = ~\sub1_data_reg_reg[102]/NET0131  & n1159 ;
  assign n5517 = ~n5515 & ~n5516 ;
  assign n5518 = ~n5028 & ~n5517 ;
  assign n5519 = ~\sub1_data_reg_reg[102]/NET0131  & n5028 ;
  assign n5520 = ~n5518 & ~n5519 ;
  assign n5521 = ~n5027 & ~n5520 ;
  assign n5522 = ~\mix1_data_o_reg_reg[102]/NET0131  & n5027 ;
  assign n5523 = ~n5521 & ~n5522 ;
  assign n5524 = n5026 & ~n5523 ;
  assign n5525 = ~\sub1_data_reg_reg[102]/NET0131  & ~n5026 ;
  assign n5526 = ~n5524 & ~n5525 ;
  assign n5527 = \state_reg/NET0131  & ~n5526 ;
  assign n5528 = ~\state_reg/NET0131  & ~n5517 ;
  assign n5529 = ~n5527 & ~n5528 ;
  assign n5531 = \key_i[102]_pad  & n5529 ;
  assign n5530 = ~\key_i[102]_pad  & ~n5529 ;
  assign n5532 = n933 & ~n5530 ;
  assign n5533 = ~n5531 & n5532 ;
  assign n5535 = ~\ks1_key_reg_reg[102]/NET0131  & ~n5529 ;
  assign n5536 = \ks1_key_reg_reg[102]/NET0131  & n5529 ;
  assign n5537 = ~n5535 & ~n5536 ;
  assign n5538 = n5053 & ~n5537 ;
  assign n5534 = ~\data_o[102]_pad  & ~n5053 ;
  assign n5539 = ~n933 & ~n5534 ;
  assign n5540 = ~n5538 & n5539 ;
  assign n5541 = ~n5533 & ~n5540 ;
  assign n5542 = ~\data_i[114]_pad  & ~n5029 ;
  assign n5543 = ~\mix1_data_o_reg_reg[114]/NET0131  & n5029 ;
  assign n5544 = ~n5542 & ~n5543 ;
  assign n5545 = ~n1159 & ~n5544 ;
  assign n5546 = ~\sub1_data_reg_reg[114]/NET0131  & n1159 ;
  assign n5547 = ~n5545 & ~n5546 ;
  assign n5548 = ~n5028 & ~n5547 ;
  assign n5549 = ~\sub1_data_reg_reg[114]/NET0131  & n5028 ;
  assign n5550 = ~n5548 & ~n5549 ;
  assign n5551 = ~n5027 & ~n5550 ;
  assign n5552 = ~\mix1_data_o_reg_reg[114]/NET0131  & n5027 ;
  assign n5553 = ~n5551 & ~n5552 ;
  assign n5554 = n5026 & ~n5553 ;
  assign n5555 = ~\sub1_data_reg_reg[114]/NET0131  & ~n5026 ;
  assign n5556 = ~n5554 & ~n5555 ;
  assign n5557 = \state_reg/NET0131  & ~n5556 ;
  assign n5558 = ~\state_reg/NET0131  & ~n5547 ;
  assign n5559 = ~n5557 & ~n5558 ;
  assign n5561 = \key_i[114]_pad  & n5559 ;
  assign n5560 = ~\key_i[114]_pad  & ~n5559 ;
  assign n5562 = n933 & ~n5560 ;
  assign n5563 = ~n5561 & n5562 ;
  assign n5565 = ~\ks1_key_reg_reg[114]/NET0131  & ~n5559 ;
  assign n5566 = \ks1_key_reg_reg[114]/NET0131  & n5559 ;
  assign n5567 = ~n5565 & ~n5566 ;
  assign n5568 = n5053 & ~n5567 ;
  assign n5564 = ~\data_o[114]_pad  & ~n5053 ;
  assign n5569 = ~n933 & ~n5564 ;
  assign n5570 = ~n5568 & n5569 ;
  assign n5571 = ~n5563 & ~n5570 ;
  assign n5572 = \data_i[6]_pad  & ~n5029 ;
  assign n5573 = \mix1_data_o_reg_reg[6]/NET0131  & n5029 ;
  assign n5574 = ~n5572 & ~n5573 ;
  assign n5575 = ~n1159 & ~n5574 ;
  assign n5576 = \sub1_data_reg_reg[6]/NET0131  & n1159 ;
  assign n5577 = ~n5575 & ~n5576 ;
  assign n5578 = ~n5028 & n5577 ;
  assign n5579 = ~\sub1_data_reg_reg[6]/NET0131  & n5028 ;
  assign n5580 = ~n5578 & ~n5579 ;
  assign n5581 = ~n5027 & ~n5580 ;
  assign n5582 = ~\mix1_data_o_reg_reg[6]/NET0131  & n5027 ;
  assign n5583 = ~n5581 & ~n5582 ;
  assign n5584 = n5026 & ~n5583 ;
  assign n5585 = ~\sub1_data_reg_reg[6]/NET0131  & ~n5026 ;
  assign n5586 = ~n5584 & ~n5585 ;
  assign n5587 = \state_reg/NET0131  & ~n5586 ;
  assign n5588 = ~\state_reg/NET0131  & n5577 ;
  assign n5589 = ~n5587 & ~n5588 ;
  assign n5591 = \key_i[6]_pad  & n5589 ;
  assign n5590 = ~\key_i[6]_pad  & ~n5589 ;
  assign n5592 = n933 & ~n5590 ;
  assign n5593 = ~n5591 & n5592 ;
  assign n5595 = ~\ks1_key_reg_reg[6]/NET0131  & ~n5589 ;
  assign n5596 = \ks1_key_reg_reg[6]/NET0131  & n5589 ;
  assign n5597 = ~n5595 & ~n5596 ;
  assign n5598 = n5053 & ~n5597 ;
  assign n5594 = ~\data_o[6]_pad  & ~n5053 ;
  assign n5599 = ~n933 & ~n5594 ;
  assign n5600 = ~n5598 & n5599 ;
  assign n5601 = ~n5593 & ~n5600 ;
  assign n5602 = ~\data_i[22]_pad  & ~n5029 ;
  assign n5603 = ~\mix1_data_o_reg_reg[22]/NET0131  & n5029 ;
  assign n5604 = ~n5602 & ~n5603 ;
  assign n5605 = ~n1159 & ~n5604 ;
  assign n5606 = ~\sub1_data_reg_reg[22]/NET0131  & n1159 ;
  assign n5607 = ~n5605 & ~n5606 ;
  assign n5608 = ~n5028 & ~n5607 ;
  assign n5609 = ~\sub1_data_reg_reg[22]/NET0131  & n5028 ;
  assign n5610 = ~n5608 & ~n5609 ;
  assign n5611 = ~n5027 & ~n5610 ;
  assign n5612 = ~\mix1_data_o_reg_reg[22]/NET0131  & n5027 ;
  assign n5613 = ~n5611 & ~n5612 ;
  assign n5614 = n5026 & ~n5613 ;
  assign n5615 = ~\sub1_data_reg_reg[22]/NET0131  & ~n5026 ;
  assign n5616 = ~n5614 & ~n5615 ;
  assign n5617 = \state_reg/NET0131  & ~n5616 ;
  assign n5618 = ~\state_reg/NET0131  & ~n5607 ;
  assign n5619 = ~n5617 & ~n5618 ;
  assign n5621 = \key_i[22]_pad  & n5619 ;
  assign n5620 = ~\key_i[22]_pad  & ~n5619 ;
  assign n5622 = n933 & ~n5620 ;
  assign n5623 = ~n5621 & n5622 ;
  assign n5625 = ~\ks1_key_reg_reg[22]/NET0131  & ~n5619 ;
  assign n5626 = \ks1_key_reg_reg[22]/NET0131  & n5619 ;
  assign n5627 = ~n5625 & ~n5626 ;
  assign n5628 = n5053 & ~n5627 ;
  assign n5624 = ~\data_o[22]_pad  & ~n5053 ;
  assign n5629 = ~n933 & ~n5624 ;
  assign n5630 = ~n5628 & n5629 ;
  assign n5631 = ~n5623 & ~n5630 ;
  assign n5632 = ~\data_i[70]_pad  & ~n5029 ;
  assign n5633 = ~\mix1_data_o_reg_reg[70]/NET0131  & n5029 ;
  assign n5634 = ~n5632 & ~n5633 ;
  assign n5635 = ~n1159 & ~n5634 ;
  assign n5636 = ~\sub1_data_reg_reg[70]/NET0131  & n1159 ;
  assign n5637 = ~n5635 & ~n5636 ;
  assign n5638 = ~n5028 & ~n5637 ;
  assign n5639 = ~\sub1_data_reg_reg[70]/NET0131  & n5028 ;
  assign n5640 = ~n5638 & ~n5639 ;
  assign n5641 = ~n5027 & ~n5640 ;
  assign n5642 = ~\mix1_data_o_reg_reg[70]/NET0131  & n5027 ;
  assign n5643 = ~n5641 & ~n5642 ;
  assign n5644 = n5026 & ~n5643 ;
  assign n5645 = ~\sub1_data_reg_reg[70]/NET0131  & ~n5026 ;
  assign n5646 = ~n5644 & ~n5645 ;
  assign n5647 = \state_reg/NET0131  & ~n5646 ;
  assign n5648 = ~\state_reg/NET0131  & ~n5637 ;
  assign n5649 = ~n5647 & ~n5648 ;
  assign n5651 = \key_i[70]_pad  & n5649 ;
  assign n5650 = ~\key_i[70]_pad  & ~n5649 ;
  assign n5652 = n933 & ~n5650 ;
  assign n5653 = ~n5651 & n5652 ;
  assign n5655 = ~\ks1_key_reg_reg[70]/NET0131  & ~n5649 ;
  assign n5656 = \ks1_key_reg_reg[70]/NET0131  & n5649 ;
  assign n5657 = ~n5655 & ~n5656 ;
  assign n5658 = n5053 & ~n5657 ;
  assign n5654 = ~\data_o[70]_pad  & ~n5053 ;
  assign n5659 = ~n933 & ~n5654 ;
  assign n5660 = ~n5658 & n5659 ;
  assign n5661 = ~n5653 & ~n5660 ;
  assign n5662 = ~\data_i[71]_pad  & ~n5029 ;
  assign n5663 = ~\mix1_data_o_reg_reg[71]/NET0131  & n5029 ;
  assign n5664 = ~n5662 & ~n5663 ;
  assign n5665 = ~n1159 & ~n5664 ;
  assign n5666 = ~\sub1_data_reg_reg[71]/NET0131  & n1159 ;
  assign n5667 = ~n5665 & ~n5666 ;
  assign n5668 = ~n5028 & ~n5667 ;
  assign n5669 = ~\sub1_data_reg_reg[71]/NET0131  & n5028 ;
  assign n5670 = ~n5668 & ~n5669 ;
  assign n5671 = ~n5027 & ~n5670 ;
  assign n5672 = ~\mix1_data_o_reg_reg[71]/NET0131  & n5027 ;
  assign n5673 = ~n5671 & ~n5672 ;
  assign n5674 = n5026 & ~n5673 ;
  assign n5675 = ~\sub1_data_reg_reg[71]/NET0131  & ~n5026 ;
  assign n5676 = ~n5674 & ~n5675 ;
  assign n5677 = \state_reg/NET0131  & ~n5676 ;
  assign n5678 = ~\state_reg/NET0131  & ~n5667 ;
  assign n5679 = ~n5677 & ~n5678 ;
  assign n5681 = \key_i[71]_pad  & n5679 ;
  assign n5680 = ~\key_i[71]_pad  & ~n5679 ;
  assign n5682 = n933 & ~n5680 ;
  assign n5683 = ~n5681 & n5682 ;
  assign n5685 = ~\ks1_key_reg_reg[71]/NET0131  & ~n5679 ;
  assign n5686 = \ks1_key_reg_reg[71]/NET0131  & n5679 ;
  assign n5687 = ~n5685 & ~n5686 ;
  assign n5688 = n5053 & ~n5687 ;
  assign n5684 = ~\data_o[71]_pad  & ~n5053 ;
  assign n5689 = ~n933 & ~n5684 ;
  assign n5690 = ~n5688 & n5689 ;
  assign n5691 = ~n5683 & ~n5690 ;
  assign n5692 = ~\data_i[23]_pad  & ~n5029 ;
  assign n5693 = ~\mix1_data_o_reg_reg[23]/NET0131  & n5029 ;
  assign n5694 = ~n5692 & ~n5693 ;
  assign n5695 = ~n1159 & ~n5694 ;
  assign n5696 = ~\sub1_data_reg_reg[23]/NET0131  & n1159 ;
  assign n5697 = ~n5695 & ~n5696 ;
  assign n5698 = ~n5028 & ~n5697 ;
  assign n5699 = ~\sub1_data_reg_reg[23]/NET0131  & n5028 ;
  assign n5700 = ~n5698 & ~n5699 ;
  assign n5701 = ~n5027 & ~n5700 ;
  assign n5702 = ~\mix1_data_o_reg_reg[23]/NET0131  & n5027 ;
  assign n5703 = ~n5701 & ~n5702 ;
  assign n5704 = n5026 & ~n5703 ;
  assign n5705 = ~\sub1_data_reg_reg[23]/NET0131  & ~n5026 ;
  assign n5706 = ~n5704 & ~n5705 ;
  assign n5707 = \state_reg/NET0131  & ~n5706 ;
  assign n5708 = ~\state_reg/NET0131  & ~n5697 ;
  assign n5709 = ~n5707 & ~n5708 ;
  assign n5711 = \key_i[23]_pad  & n5709 ;
  assign n5710 = ~\key_i[23]_pad  & ~n5709 ;
  assign n5712 = n933 & ~n5710 ;
  assign n5713 = ~n5711 & n5712 ;
  assign n5715 = ~\ks1_key_reg_reg[23]/NET0131  & ~n5709 ;
  assign n5716 = \ks1_key_reg_reg[23]/NET0131  & n5709 ;
  assign n5717 = ~n5715 & ~n5716 ;
  assign n5718 = n5053 & ~n5717 ;
  assign n5714 = ~\data_o[23]_pad  & ~n5053 ;
  assign n5719 = ~n933 & ~n5714 ;
  assign n5720 = ~n5718 & n5719 ;
  assign n5721 = ~n5713 & ~n5720 ;
  assign n5722 = ~\data_i[115]_pad  & ~n5029 ;
  assign n5723 = ~\mix1_data_o_reg_reg[115]/NET0131  & n5029 ;
  assign n5724 = ~n5722 & ~n5723 ;
  assign n5725 = ~n1159 & ~n5724 ;
  assign n5726 = ~\sub1_data_reg_reg[115]/NET0131  & n1159 ;
  assign n5727 = ~n5725 & ~n5726 ;
  assign n5728 = ~n5028 & ~n5727 ;
  assign n5729 = ~\sub1_data_reg_reg[115]/NET0131  & n5028 ;
  assign n5730 = ~n5728 & ~n5729 ;
  assign n5731 = ~n5027 & ~n5730 ;
  assign n5732 = ~\mix1_data_o_reg_reg[115]/NET0131  & n5027 ;
  assign n5733 = ~n5731 & ~n5732 ;
  assign n5734 = n5026 & ~n5733 ;
  assign n5735 = ~\sub1_data_reg_reg[115]/NET0131  & ~n5026 ;
  assign n5736 = ~n5734 & ~n5735 ;
  assign n5737 = \state_reg/NET0131  & ~n5736 ;
  assign n5738 = ~\state_reg/NET0131  & ~n5727 ;
  assign n5739 = ~n5737 & ~n5738 ;
  assign n5741 = \key_i[115]_pad  & n5739 ;
  assign n5740 = ~\key_i[115]_pad  & ~n5739 ;
  assign n5742 = n933 & ~n5740 ;
  assign n5743 = ~n5741 & n5742 ;
  assign n5745 = ~\ks1_key_reg_reg[115]/NET0131  & ~n5739 ;
  assign n5746 = \ks1_key_reg_reg[115]/NET0131  & n5739 ;
  assign n5747 = ~n5745 & ~n5746 ;
  assign n5748 = n5053 & ~n5747 ;
  assign n5744 = ~\data_o[115]_pad  & ~n5053 ;
  assign n5749 = ~n933 & ~n5744 ;
  assign n5750 = ~n5748 & n5749 ;
  assign n5751 = ~n5743 & ~n5750 ;
  assign n5752 = \data_i[72]_pad  & ~n5029 ;
  assign n5753 = \mix1_data_o_reg_reg[72]/NET0131  & n5029 ;
  assign n5754 = ~n5752 & ~n5753 ;
  assign n5755 = ~n1159 & ~n5754 ;
  assign n5756 = \sub1_data_reg_reg[72]/NET0131  & n1159 ;
  assign n5757 = ~n5755 & ~n5756 ;
  assign n5758 = ~n5028 & n5757 ;
  assign n5759 = ~\sub1_data_reg_reg[72]/NET0131  & n5028 ;
  assign n5760 = ~n5758 & ~n5759 ;
  assign n5761 = ~n5027 & ~n5760 ;
  assign n5762 = ~\mix1_data_o_reg_reg[72]/NET0131  & n5027 ;
  assign n5763 = ~n5761 & ~n5762 ;
  assign n5764 = n5026 & ~n5763 ;
  assign n5765 = ~\sub1_data_reg_reg[72]/NET0131  & ~n5026 ;
  assign n5766 = ~n5764 & ~n5765 ;
  assign n5767 = \state_reg/NET0131  & ~n5766 ;
  assign n5768 = ~\state_reg/NET0131  & n5757 ;
  assign n5769 = ~n5767 & ~n5768 ;
  assign n5771 = \key_i[72]_pad  & n5769 ;
  assign n5770 = ~\key_i[72]_pad  & ~n5769 ;
  assign n5772 = n933 & ~n5770 ;
  assign n5773 = ~n5771 & n5772 ;
  assign n5775 = ~\ks1_key_reg_reg[72]/P0002  & ~n5769 ;
  assign n5776 = \ks1_key_reg_reg[72]/P0002  & n5769 ;
  assign n5777 = ~n5775 & ~n5776 ;
  assign n5778 = n5053 & ~n5777 ;
  assign n5774 = ~\data_o[72]_pad  & ~n5053 ;
  assign n5779 = ~n933 & ~n5774 ;
  assign n5780 = ~n5778 & n5779 ;
  assign n5781 = ~n5773 & ~n5780 ;
  assign n5782 = \data_i[24]_pad  & ~n5029 ;
  assign n5783 = \mix1_data_o_reg_reg[24]/NET0131  & n5029 ;
  assign n5784 = ~n5782 & ~n5783 ;
  assign n5785 = ~n1159 & ~n5784 ;
  assign n5786 = \sub1_data_reg_reg[24]/NET0131  & n1159 ;
  assign n5787 = ~n5785 & ~n5786 ;
  assign n5788 = ~n5028 & n5787 ;
  assign n5789 = ~\sub1_data_reg_reg[24]/NET0131  & n5028 ;
  assign n5790 = ~n5788 & ~n5789 ;
  assign n5791 = ~n5027 & ~n5790 ;
  assign n5792 = ~\mix1_data_o_reg_reg[24]/NET0131  & n5027 ;
  assign n5793 = ~n5791 & ~n5792 ;
  assign n5794 = n5026 & ~n5793 ;
  assign n5795 = ~\sub1_data_reg_reg[24]/NET0131  & ~n5026 ;
  assign n5796 = ~n5794 & ~n5795 ;
  assign n5797 = \state_reg/NET0131  & ~n5796 ;
  assign n5798 = ~\state_reg/NET0131  & n5787 ;
  assign n5799 = ~n5797 & ~n5798 ;
  assign n5801 = \key_i[24]_pad  & n5799 ;
  assign n5800 = ~\key_i[24]_pad  & ~n5799 ;
  assign n5802 = n933 & ~n5800 ;
  assign n5803 = ~n5801 & n5802 ;
  assign n5805 = ~\ks1_key_reg_reg[24]/NET0131  & ~n5799 ;
  assign n5806 = \ks1_key_reg_reg[24]/NET0131  & n5799 ;
  assign n5807 = ~n5805 & ~n5806 ;
  assign n5808 = n5053 & ~n5807 ;
  assign n5804 = ~\data_o[24]_pad  & ~n5053 ;
  assign n5809 = ~n933 & ~n5804 ;
  assign n5810 = ~n5808 & n5809 ;
  assign n5811 = ~n5803 & ~n5810 ;
  assign n5812 = \data_i[73]_pad  & ~n5029 ;
  assign n5813 = \mix1_data_o_reg_reg[73]/NET0131  & n5029 ;
  assign n5814 = ~n5812 & ~n5813 ;
  assign n5815 = ~n1159 & ~n5814 ;
  assign n5816 = \sub1_data_reg_reg[73]/NET0131  & n1159 ;
  assign n5817 = ~n5815 & ~n5816 ;
  assign n5818 = ~n5028 & n5817 ;
  assign n5819 = ~\sub1_data_reg_reg[73]/NET0131  & n5028 ;
  assign n5820 = ~n5818 & ~n5819 ;
  assign n5821 = ~n5027 & ~n5820 ;
  assign n5822 = ~\mix1_data_o_reg_reg[73]/NET0131  & n5027 ;
  assign n5823 = ~n5821 & ~n5822 ;
  assign n5824 = n5026 & ~n5823 ;
  assign n5825 = ~\sub1_data_reg_reg[73]/NET0131  & ~n5026 ;
  assign n5826 = ~n5824 & ~n5825 ;
  assign n5827 = \state_reg/NET0131  & ~n5826 ;
  assign n5828 = ~\state_reg/NET0131  & n5817 ;
  assign n5829 = ~n5827 & ~n5828 ;
  assign n5831 = \key_i[73]_pad  & n5829 ;
  assign n5830 = ~\key_i[73]_pad  & ~n5829 ;
  assign n5832 = n933 & ~n5830 ;
  assign n5833 = ~n5831 & n5832 ;
  assign n5835 = ~\ks1_key_reg_reg[73]/NET0131  & ~n5829 ;
  assign n5836 = \ks1_key_reg_reg[73]/NET0131  & n5829 ;
  assign n5837 = ~n5835 & ~n5836 ;
  assign n5838 = n5053 & ~n5837 ;
  assign n5834 = ~\data_o[73]_pad  & ~n5053 ;
  assign n5839 = ~n933 & ~n5834 ;
  assign n5840 = ~n5838 & n5839 ;
  assign n5841 = ~n5833 & ~n5840 ;
  assign n5842 = \data_i[74]_pad  & ~n5029 ;
  assign n5843 = \mix1_data_o_reg_reg[74]/NET0131  & n5029 ;
  assign n5844 = ~n5842 & ~n5843 ;
  assign n5845 = ~n1159 & ~n5844 ;
  assign n5846 = \sub1_data_reg_reg[74]/NET0131  & n1159 ;
  assign n5847 = ~n5845 & ~n5846 ;
  assign n5848 = ~n5028 & n5847 ;
  assign n5849 = ~\sub1_data_reg_reg[74]/NET0131  & n5028 ;
  assign n5850 = ~n5848 & ~n5849 ;
  assign n5851 = ~n5027 & ~n5850 ;
  assign n5852 = ~\mix1_data_o_reg_reg[74]/NET0131  & n5027 ;
  assign n5853 = ~n5851 & ~n5852 ;
  assign n5854 = n5026 & ~n5853 ;
  assign n5855 = ~\sub1_data_reg_reg[74]/NET0131  & ~n5026 ;
  assign n5856 = ~n5854 & ~n5855 ;
  assign n5857 = \state_reg/NET0131  & ~n5856 ;
  assign n5858 = ~\state_reg/NET0131  & n5847 ;
  assign n5859 = ~n5857 & ~n5858 ;
  assign n5861 = \key_i[74]_pad  & n5859 ;
  assign n5860 = ~\key_i[74]_pad  & ~n5859 ;
  assign n5862 = n933 & ~n5860 ;
  assign n5863 = ~n5861 & n5862 ;
  assign n5865 = ~\ks1_key_reg_reg[74]/NET0131  & ~n5859 ;
  assign n5866 = \ks1_key_reg_reg[74]/NET0131  & n5859 ;
  assign n5867 = ~n5865 & ~n5866 ;
  assign n5868 = n5053 & ~n5867 ;
  assign n5864 = ~\data_o[74]_pad  & ~n5053 ;
  assign n5869 = ~n933 & ~n5864 ;
  assign n5870 = ~n5868 & n5869 ;
  assign n5871 = ~n5863 & ~n5870 ;
  assign n5872 = \data_i[25]_pad  & ~n5029 ;
  assign n5873 = \mix1_data_o_reg_reg[25]/NET0131  & n5029 ;
  assign n5874 = ~n5872 & ~n5873 ;
  assign n5875 = ~n1159 & ~n5874 ;
  assign n5876 = \sub1_data_reg_reg[25]/NET0131  & n1159 ;
  assign n5877 = ~n5875 & ~n5876 ;
  assign n5878 = ~n5028 & n5877 ;
  assign n5879 = ~\sub1_data_reg_reg[25]/NET0131  & n5028 ;
  assign n5880 = ~n5878 & ~n5879 ;
  assign n5881 = ~n5027 & ~n5880 ;
  assign n5882 = ~\mix1_data_o_reg_reg[25]/NET0131  & n5027 ;
  assign n5883 = ~n5881 & ~n5882 ;
  assign n5884 = n5026 & ~n5883 ;
  assign n5885 = ~\sub1_data_reg_reg[25]/NET0131  & ~n5026 ;
  assign n5886 = ~n5884 & ~n5885 ;
  assign n5887 = \state_reg/NET0131  & ~n5886 ;
  assign n5888 = ~\state_reg/NET0131  & n5877 ;
  assign n5889 = ~n5887 & ~n5888 ;
  assign n5891 = \key_i[25]_pad  & n5889 ;
  assign n5890 = ~\key_i[25]_pad  & ~n5889 ;
  assign n5892 = n933 & ~n5890 ;
  assign n5893 = ~n5891 & n5892 ;
  assign n5895 = ~\ks1_key_reg_reg[25]/NET0131  & ~n5889 ;
  assign n5896 = \ks1_key_reg_reg[25]/NET0131  & n5889 ;
  assign n5897 = ~n5895 & ~n5896 ;
  assign n5898 = n5053 & ~n5897 ;
  assign n5894 = ~\data_o[25]_pad  & ~n5053 ;
  assign n5899 = ~n933 & ~n5894 ;
  assign n5900 = ~n5898 & n5899 ;
  assign n5901 = ~n5893 & ~n5900 ;
  assign n5902 = \data_i[75]_pad  & ~n5029 ;
  assign n5903 = \mix1_data_o_reg_reg[75]/NET0131  & n5029 ;
  assign n5904 = ~n5902 & ~n5903 ;
  assign n5905 = ~n1159 & ~n5904 ;
  assign n5906 = \sub1_data_reg_reg[75]/NET0131  & n1159 ;
  assign n5907 = ~n5905 & ~n5906 ;
  assign n5908 = ~n5028 & n5907 ;
  assign n5909 = ~\sub1_data_reg_reg[75]/NET0131  & n5028 ;
  assign n5910 = ~n5908 & ~n5909 ;
  assign n5911 = ~n5027 & ~n5910 ;
  assign n5912 = ~\mix1_data_o_reg_reg[75]/NET0131  & n5027 ;
  assign n5913 = ~n5911 & ~n5912 ;
  assign n5914 = n5026 & ~n5913 ;
  assign n5915 = ~\sub1_data_reg_reg[75]/NET0131  & ~n5026 ;
  assign n5916 = ~n5914 & ~n5915 ;
  assign n5917 = \state_reg/NET0131  & ~n5916 ;
  assign n5918 = ~\state_reg/NET0131  & n5907 ;
  assign n5919 = ~n5917 & ~n5918 ;
  assign n5921 = \key_i[75]_pad  & n5919 ;
  assign n5920 = ~\key_i[75]_pad  & ~n5919 ;
  assign n5922 = n933 & ~n5920 ;
  assign n5923 = ~n5921 & n5922 ;
  assign n5925 = ~\ks1_key_reg_reg[75]/P0002  & ~n5919 ;
  assign n5926 = \ks1_key_reg_reg[75]/P0002  & n5919 ;
  assign n5927 = ~n5925 & ~n5926 ;
  assign n5928 = n5053 & ~n5927 ;
  assign n5924 = ~\data_o[75]_pad  & ~n5053 ;
  assign n5929 = ~n933 & ~n5924 ;
  assign n5930 = ~n5928 & n5929 ;
  assign n5931 = ~n5923 & ~n5930 ;
  assign n5932 = \data_i[76]_pad  & ~n5029 ;
  assign n5933 = \mix1_data_o_reg_reg[76]/NET0131  & n5029 ;
  assign n5934 = ~n5932 & ~n5933 ;
  assign n5935 = ~n1159 & ~n5934 ;
  assign n5936 = \sub1_data_reg_reg[76]/NET0131  & n1159 ;
  assign n5937 = ~n5935 & ~n5936 ;
  assign n5938 = ~n5028 & n5937 ;
  assign n5939 = ~\sub1_data_reg_reg[76]/NET0131  & n5028 ;
  assign n5940 = ~n5938 & ~n5939 ;
  assign n5941 = ~n5027 & ~n5940 ;
  assign n5942 = ~\mix1_data_o_reg_reg[76]/NET0131  & n5027 ;
  assign n5943 = ~n5941 & ~n5942 ;
  assign n5944 = n5026 & ~n5943 ;
  assign n5945 = ~\sub1_data_reg_reg[76]/NET0131  & ~n5026 ;
  assign n5946 = ~n5944 & ~n5945 ;
  assign n5947 = \state_reg/NET0131  & ~n5946 ;
  assign n5948 = ~\state_reg/NET0131  & n5937 ;
  assign n5949 = ~n5947 & ~n5948 ;
  assign n5951 = \key_i[76]_pad  & n5949 ;
  assign n5950 = ~\key_i[76]_pad  & ~n5949 ;
  assign n5952 = n933 & ~n5950 ;
  assign n5953 = ~n5951 & n5952 ;
  assign n5955 = ~\ks1_key_reg_reg[76]/P0002  & ~n5949 ;
  assign n5956 = \ks1_key_reg_reg[76]/P0002  & n5949 ;
  assign n5957 = ~n5955 & ~n5956 ;
  assign n5958 = n5053 & ~n5957 ;
  assign n5954 = ~\data_o[76]_pad  & ~n5053 ;
  assign n5959 = ~n933 & ~n5954 ;
  assign n5960 = ~n5958 & n5959 ;
  assign n5961 = ~n5953 & ~n5960 ;
  assign n5962 = \data_i[77]_pad  & ~n5029 ;
  assign n5963 = \mix1_data_o_reg_reg[77]/NET0131  & n5029 ;
  assign n5964 = ~n5962 & ~n5963 ;
  assign n5965 = ~n1159 & ~n5964 ;
  assign n5966 = \sub1_data_reg_reg[77]/NET0131  & n1159 ;
  assign n5967 = ~n5965 & ~n5966 ;
  assign n5968 = ~n5028 & n5967 ;
  assign n5969 = ~\sub1_data_reg_reg[77]/NET0131  & n5028 ;
  assign n5970 = ~n5968 & ~n5969 ;
  assign n5971 = ~n5027 & ~n5970 ;
  assign n5972 = ~\mix1_data_o_reg_reg[77]/NET0131  & n5027 ;
  assign n5973 = ~n5971 & ~n5972 ;
  assign n5974 = n5026 & ~n5973 ;
  assign n5975 = ~\sub1_data_reg_reg[77]/NET0131  & ~n5026 ;
  assign n5976 = ~n5974 & ~n5975 ;
  assign n5977 = \state_reg/NET0131  & ~n5976 ;
  assign n5978 = ~\state_reg/NET0131  & n5967 ;
  assign n5979 = ~n5977 & ~n5978 ;
  assign n5981 = \key_i[77]_pad  & n5979 ;
  assign n5980 = ~\key_i[77]_pad  & ~n5979 ;
  assign n5982 = n933 & ~n5980 ;
  assign n5983 = ~n5981 & n5982 ;
  assign n5985 = ~\ks1_key_reg_reg[77]/P0002  & ~n5979 ;
  assign n5986 = \ks1_key_reg_reg[77]/P0002  & n5979 ;
  assign n5987 = ~n5985 & ~n5986 ;
  assign n5988 = n5053 & ~n5987 ;
  assign n5984 = ~\data_o[77]_pad  & ~n5053 ;
  assign n5989 = ~n933 & ~n5984 ;
  assign n5990 = ~n5988 & n5989 ;
  assign n5991 = ~n5983 & ~n5990 ;
  assign n5992 = \data_i[26]_pad  & ~n5029 ;
  assign n5993 = \mix1_data_o_reg_reg[26]/NET0131  & n5029 ;
  assign n5994 = ~n5992 & ~n5993 ;
  assign n5995 = ~n1159 & ~n5994 ;
  assign n5996 = \sub1_data_reg_reg[26]/NET0131  & n1159 ;
  assign n5997 = ~n5995 & ~n5996 ;
  assign n5998 = ~n5028 & n5997 ;
  assign n5999 = ~\sub1_data_reg_reg[26]/NET0131  & n5028 ;
  assign n6000 = ~n5998 & ~n5999 ;
  assign n6001 = ~n5027 & ~n6000 ;
  assign n6002 = ~\mix1_data_o_reg_reg[26]/NET0131  & n5027 ;
  assign n6003 = ~n6001 & ~n6002 ;
  assign n6004 = n5026 & ~n6003 ;
  assign n6005 = ~\sub1_data_reg_reg[26]/NET0131  & ~n5026 ;
  assign n6006 = ~n6004 & ~n6005 ;
  assign n6007 = \state_reg/NET0131  & ~n6006 ;
  assign n6008 = ~\state_reg/NET0131  & n5997 ;
  assign n6009 = ~n6007 & ~n6008 ;
  assign n6011 = \key_i[26]_pad  & n6009 ;
  assign n6010 = ~\key_i[26]_pad  & ~n6009 ;
  assign n6012 = n933 & ~n6010 ;
  assign n6013 = ~n6011 & n6012 ;
  assign n6015 = ~\ks1_key_reg_reg[26]/NET0131  & ~n6009 ;
  assign n6016 = \ks1_key_reg_reg[26]/NET0131  & n6009 ;
  assign n6017 = ~n6015 & ~n6016 ;
  assign n6018 = n5053 & ~n6017 ;
  assign n6014 = ~\data_o[26]_pad  & ~n5053 ;
  assign n6019 = ~n933 & ~n6014 ;
  assign n6020 = ~n6018 & n6019 ;
  assign n6021 = ~n6013 & ~n6020 ;
  assign n6022 = ~\data_i[103]_pad  & ~n5029 ;
  assign n6023 = ~\mix1_data_o_reg_reg[103]/NET0131  & n5029 ;
  assign n6024 = ~n6022 & ~n6023 ;
  assign n6025 = ~n1159 & ~n6024 ;
  assign n6026 = ~\sub1_data_reg_reg[103]/NET0131  & n1159 ;
  assign n6027 = ~n6025 & ~n6026 ;
  assign n6028 = ~n5028 & ~n6027 ;
  assign n6029 = ~\sub1_data_reg_reg[103]/NET0131  & n5028 ;
  assign n6030 = ~n6028 & ~n6029 ;
  assign n6031 = ~n5027 & ~n6030 ;
  assign n6032 = ~\mix1_data_o_reg_reg[103]/NET0131  & n5027 ;
  assign n6033 = ~n6031 & ~n6032 ;
  assign n6034 = n5026 & ~n6033 ;
  assign n6035 = ~\sub1_data_reg_reg[103]/NET0131  & ~n5026 ;
  assign n6036 = ~n6034 & ~n6035 ;
  assign n6037 = \state_reg/NET0131  & ~n6036 ;
  assign n6038 = ~\state_reg/NET0131  & ~n6027 ;
  assign n6039 = ~n6037 & ~n6038 ;
  assign n6041 = \key_i[103]_pad  & n6039 ;
  assign n6040 = ~\key_i[103]_pad  & ~n6039 ;
  assign n6042 = n933 & ~n6040 ;
  assign n6043 = ~n6041 & n6042 ;
  assign n6045 = ~\ks1_key_reg_reg[103]/NET0131  & ~n6039 ;
  assign n6046 = \ks1_key_reg_reg[103]/NET0131  & n6039 ;
  assign n6047 = ~n6045 & ~n6046 ;
  assign n6048 = n5053 & ~n6047 ;
  assign n6044 = ~\data_o[103]_pad  & ~n5053 ;
  assign n6049 = ~n933 & ~n6044 ;
  assign n6050 = ~n6048 & n6049 ;
  assign n6051 = ~n6043 & ~n6050 ;
  assign n6052 = \data_i[78]_pad  & ~n5029 ;
  assign n6053 = \mix1_data_o_reg_reg[78]/NET0131  & n5029 ;
  assign n6054 = ~n6052 & ~n6053 ;
  assign n6055 = ~n1159 & ~n6054 ;
  assign n6056 = \sub1_data_reg_reg[78]/NET0131  & n1159 ;
  assign n6057 = ~n6055 & ~n6056 ;
  assign n6058 = ~n5028 & n6057 ;
  assign n6059 = ~\sub1_data_reg_reg[78]/NET0131  & n5028 ;
  assign n6060 = ~n6058 & ~n6059 ;
  assign n6061 = ~n5027 & ~n6060 ;
  assign n6062 = ~\mix1_data_o_reg_reg[78]/NET0131  & n5027 ;
  assign n6063 = ~n6061 & ~n6062 ;
  assign n6064 = n5026 & ~n6063 ;
  assign n6065 = ~\sub1_data_reg_reg[78]/NET0131  & ~n5026 ;
  assign n6066 = ~n6064 & ~n6065 ;
  assign n6067 = \state_reg/NET0131  & ~n6066 ;
  assign n6068 = ~\state_reg/NET0131  & n6057 ;
  assign n6069 = ~n6067 & ~n6068 ;
  assign n6071 = \key_i[78]_pad  & n6069 ;
  assign n6070 = ~\key_i[78]_pad  & ~n6069 ;
  assign n6072 = n933 & ~n6070 ;
  assign n6073 = ~n6071 & n6072 ;
  assign n6075 = ~\ks1_key_reg_reg[78]/P0002  & ~n6069 ;
  assign n6076 = \ks1_key_reg_reg[78]/P0002  & n6069 ;
  assign n6077 = ~n6075 & ~n6076 ;
  assign n6078 = n5053 & ~n6077 ;
  assign n6074 = ~\data_o[78]_pad  & ~n5053 ;
  assign n6079 = ~n933 & ~n6074 ;
  assign n6080 = ~n6078 & n6079 ;
  assign n6081 = ~n6073 & ~n6080 ;
  assign n6082 = ~\data_i[116]_pad  & ~n5029 ;
  assign n6083 = ~\mix1_data_o_reg_reg[116]/NET0131  & n5029 ;
  assign n6084 = ~n6082 & ~n6083 ;
  assign n6085 = ~n1159 & ~n6084 ;
  assign n6086 = ~\sub1_data_reg_reg[116]/NET0131  & n1159 ;
  assign n6087 = ~n6085 & ~n6086 ;
  assign n6088 = ~n5028 & ~n6087 ;
  assign n6089 = ~\sub1_data_reg_reg[116]/NET0131  & n5028 ;
  assign n6090 = ~n6088 & ~n6089 ;
  assign n6091 = ~n5027 & ~n6090 ;
  assign n6092 = ~\mix1_data_o_reg_reg[116]/NET0131  & n5027 ;
  assign n6093 = ~n6091 & ~n6092 ;
  assign n6094 = n5026 & ~n6093 ;
  assign n6095 = ~\sub1_data_reg_reg[116]/NET0131  & ~n5026 ;
  assign n6096 = ~n6094 & ~n6095 ;
  assign n6097 = \state_reg/NET0131  & ~n6096 ;
  assign n6098 = ~\state_reg/NET0131  & ~n6087 ;
  assign n6099 = ~n6097 & ~n6098 ;
  assign n6101 = \key_i[116]_pad  & n6099 ;
  assign n6100 = ~\key_i[116]_pad  & ~n6099 ;
  assign n6102 = n933 & ~n6100 ;
  assign n6103 = ~n6101 & n6102 ;
  assign n6105 = ~\ks1_key_reg_reg[116]/NET0131  & ~n6099 ;
  assign n6106 = \ks1_key_reg_reg[116]/NET0131  & n6099 ;
  assign n6107 = ~n6105 & ~n6106 ;
  assign n6108 = n5053 & ~n6107 ;
  assign n6104 = ~\data_o[116]_pad  & ~n5053 ;
  assign n6109 = ~n933 & ~n6104 ;
  assign n6110 = ~n6108 & n6109 ;
  assign n6111 = ~n6103 & ~n6110 ;
  assign n6112 = \data_i[79]_pad  & ~n5029 ;
  assign n6113 = \mix1_data_o_reg_reg[79]/NET0131  & n5029 ;
  assign n6114 = ~n6112 & ~n6113 ;
  assign n6115 = ~n1159 & ~n6114 ;
  assign n6116 = \sub1_data_reg_reg[79]/NET0131  & n1159 ;
  assign n6117 = ~n6115 & ~n6116 ;
  assign n6118 = ~n5028 & n6117 ;
  assign n6119 = ~\sub1_data_reg_reg[79]/NET0131  & n5028 ;
  assign n6120 = ~n6118 & ~n6119 ;
  assign n6121 = ~n5027 & ~n6120 ;
  assign n6122 = ~\mix1_data_o_reg_reg[79]/NET0131  & n5027 ;
  assign n6123 = ~n6121 & ~n6122 ;
  assign n6124 = n5026 & ~n6123 ;
  assign n6125 = ~\sub1_data_reg_reg[79]/NET0131  & ~n5026 ;
  assign n6126 = ~n6124 & ~n6125 ;
  assign n6127 = \state_reg/NET0131  & ~n6126 ;
  assign n6128 = ~\state_reg/NET0131  & n6117 ;
  assign n6129 = ~n6127 & ~n6128 ;
  assign n6131 = \key_i[79]_pad  & n6129 ;
  assign n6130 = ~\key_i[79]_pad  & ~n6129 ;
  assign n6132 = n933 & ~n6130 ;
  assign n6133 = ~n6131 & n6132 ;
  assign n6135 = ~\ks1_key_reg_reg[79]/P0002  & ~n6129 ;
  assign n6136 = \ks1_key_reg_reg[79]/P0002  & n6129 ;
  assign n6137 = ~n6135 & ~n6136 ;
  assign n6138 = n5053 & ~n6137 ;
  assign n6134 = ~\data_o[79]_pad  & ~n5053 ;
  assign n6139 = ~n933 & ~n6134 ;
  assign n6140 = ~n6138 & n6139 ;
  assign n6141 = ~n6133 & ~n6140 ;
  assign n6142 = \data_i[27]_pad  & ~n5029 ;
  assign n6143 = \mix1_data_o_reg_reg[27]/NET0131  & n5029 ;
  assign n6144 = ~n6142 & ~n6143 ;
  assign n6145 = ~n1159 & ~n6144 ;
  assign n6146 = \sub1_data_reg_reg[27]/NET0131  & n1159 ;
  assign n6147 = ~n6145 & ~n6146 ;
  assign n6148 = ~n5028 & n6147 ;
  assign n6149 = ~\sub1_data_reg_reg[27]/NET0131  & n5028 ;
  assign n6150 = ~n6148 & ~n6149 ;
  assign n6151 = ~n5027 & ~n6150 ;
  assign n6152 = ~\mix1_data_o_reg_reg[27]/NET0131  & n5027 ;
  assign n6153 = ~n6151 & ~n6152 ;
  assign n6154 = n5026 & ~n6153 ;
  assign n6155 = ~\sub1_data_reg_reg[27]/NET0131  & ~n5026 ;
  assign n6156 = ~n6154 & ~n6155 ;
  assign n6157 = \state_reg/NET0131  & ~n6156 ;
  assign n6158 = ~\state_reg/NET0131  & n6147 ;
  assign n6159 = ~n6157 & ~n6158 ;
  assign n6161 = \key_i[27]_pad  & n6159 ;
  assign n6160 = ~\key_i[27]_pad  & ~n6159 ;
  assign n6162 = n933 & ~n6160 ;
  assign n6163 = ~n6161 & n6162 ;
  assign n6165 = ~\ks1_key_reg_reg[27]/NET0131  & ~n6159 ;
  assign n6166 = \ks1_key_reg_reg[27]/NET0131  & n6159 ;
  assign n6167 = ~n6165 & ~n6166 ;
  assign n6168 = n5053 & ~n6167 ;
  assign n6164 = ~\data_o[27]_pad  & ~n5053 ;
  assign n6169 = ~n933 & ~n6164 ;
  assign n6170 = ~n6168 & n6169 ;
  assign n6171 = ~n6163 & ~n6170 ;
  assign n6172 = \data_i[7]_pad  & ~n5029 ;
  assign n6173 = \mix1_data_o_reg_reg[7]/NET0131  & n5029 ;
  assign n6174 = ~n6172 & ~n6173 ;
  assign n6175 = ~n1159 & ~n6174 ;
  assign n6176 = \sub1_data_reg_reg[7]/NET0131  & n1159 ;
  assign n6177 = ~n6175 & ~n6176 ;
  assign n6178 = ~n5028 & n6177 ;
  assign n6179 = ~\sub1_data_reg_reg[7]/NET0131  & n5028 ;
  assign n6180 = ~n6178 & ~n6179 ;
  assign n6181 = ~n5027 & ~n6180 ;
  assign n6182 = ~\mix1_data_o_reg_reg[7]/NET0131  & n5027 ;
  assign n6183 = ~n6181 & ~n6182 ;
  assign n6184 = n5026 & ~n6183 ;
  assign n6185 = ~\sub1_data_reg_reg[7]/NET0131  & ~n5026 ;
  assign n6186 = ~n6184 & ~n6185 ;
  assign n6187 = \state_reg/NET0131  & ~n6186 ;
  assign n6188 = ~\state_reg/NET0131  & n6177 ;
  assign n6189 = ~n6187 & ~n6188 ;
  assign n6191 = \key_i[7]_pad  & n6189 ;
  assign n6190 = ~\key_i[7]_pad  & ~n6189 ;
  assign n6192 = n933 & ~n6190 ;
  assign n6193 = ~n6191 & n6192 ;
  assign n6195 = ~\ks1_key_reg_reg[7]/NET0131  & ~n6189 ;
  assign n6196 = \ks1_key_reg_reg[7]/NET0131  & n6189 ;
  assign n6197 = ~n6195 & ~n6196 ;
  assign n6198 = n5053 & ~n6197 ;
  assign n6194 = ~\data_o[7]_pad  & ~n5053 ;
  assign n6199 = ~n933 & ~n6194 ;
  assign n6200 = ~n6198 & n6199 ;
  assign n6201 = ~n6193 & ~n6200 ;
  assign n6202 = ~\data_i[117]_pad  & ~n5029 ;
  assign n6203 = ~\mix1_data_o_reg_reg[117]/NET0131  & n5029 ;
  assign n6204 = ~n6202 & ~n6203 ;
  assign n6205 = ~n1159 & ~n6204 ;
  assign n6206 = ~\sub1_data_reg_reg[117]/NET0131  & n1159 ;
  assign n6207 = ~n6205 & ~n6206 ;
  assign n6208 = ~n5028 & ~n6207 ;
  assign n6209 = ~\sub1_data_reg_reg[117]/NET0131  & n5028 ;
  assign n6210 = ~n6208 & ~n6209 ;
  assign n6211 = ~n5027 & ~n6210 ;
  assign n6212 = ~\mix1_data_o_reg_reg[117]/NET0131  & n5027 ;
  assign n6213 = ~n6211 & ~n6212 ;
  assign n6214 = n5026 & ~n6213 ;
  assign n6215 = ~\sub1_data_reg_reg[117]/NET0131  & ~n5026 ;
  assign n6216 = ~n6214 & ~n6215 ;
  assign n6217 = \state_reg/NET0131  & ~n6216 ;
  assign n6218 = ~\state_reg/NET0131  & ~n6207 ;
  assign n6219 = ~n6217 & ~n6218 ;
  assign n6221 = \key_i[117]_pad  & n6219 ;
  assign n6220 = ~\key_i[117]_pad  & ~n6219 ;
  assign n6222 = n933 & ~n6220 ;
  assign n6223 = ~n6221 & n6222 ;
  assign n6225 = ~\ks1_key_reg_reg[117]/NET0131  & ~n6219 ;
  assign n6226 = \ks1_key_reg_reg[117]/NET0131  & n6219 ;
  assign n6227 = ~n6225 & ~n6226 ;
  assign n6228 = n5053 & ~n6227 ;
  assign n6224 = ~\data_o[117]_pad  & ~n5053 ;
  assign n6229 = ~n933 & ~n6224 ;
  assign n6230 = ~n6228 & n6229 ;
  assign n6231 = ~n6223 & ~n6230 ;
  assign n6232 = ~\data_i[80]_pad  & ~n5029 ;
  assign n6233 = ~\mix1_data_o_reg_reg[80]/NET0131  & n5029 ;
  assign n6234 = ~n6232 & ~n6233 ;
  assign n6235 = ~n1159 & ~n6234 ;
  assign n6236 = ~\sub1_data_reg_reg[80]/NET0131  & n1159 ;
  assign n6237 = ~n6235 & ~n6236 ;
  assign n6238 = ~n5028 & ~n6237 ;
  assign n6239 = ~\sub1_data_reg_reg[80]/NET0131  & n5028 ;
  assign n6240 = ~n6238 & ~n6239 ;
  assign n6241 = ~n5027 & ~n6240 ;
  assign n6242 = ~\mix1_data_o_reg_reg[80]/NET0131  & n5027 ;
  assign n6243 = ~n6241 & ~n6242 ;
  assign n6244 = n5026 & ~n6243 ;
  assign n6245 = ~\sub1_data_reg_reg[80]/NET0131  & ~n5026 ;
  assign n6246 = ~n6244 & ~n6245 ;
  assign n6247 = \state_reg/NET0131  & ~n6246 ;
  assign n6248 = ~\state_reg/NET0131  & ~n6237 ;
  assign n6249 = ~n6247 & ~n6248 ;
  assign n6251 = \key_i[80]_pad  & n6249 ;
  assign n6250 = ~\key_i[80]_pad  & ~n6249 ;
  assign n6252 = n933 & ~n6250 ;
  assign n6253 = ~n6251 & n6252 ;
  assign n6255 = ~\ks1_key_reg_reg[80]/NET0131  & ~n6249 ;
  assign n6256 = \ks1_key_reg_reg[80]/NET0131  & n6249 ;
  assign n6257 = ~n6255 & ~n6256 ;
  assign n6258 = n5053 & ~n6257 ;
  assign n6254 = ~\data_o[80]_pad  & ~n5053 ;
  assign n6259 = ~n933 & ~n6254 ;
  assign n6260 = ~n6258 & n6259 ;
  assign n6261 = ~n6253 & ~n6260 ;
  assign n6262 = \data_i[28]_pad  & ~n5029 ;
  assign n6263 = \mix1_data_o_reg_reg[28]/NET0131  & n5029 ;
  assign n6264 = ~n6262 & ~n6263 ;
  assign n6265 = ~n1159 & ~n6264 ;
  assign n6266 = \sub1_data_reg_reg[28]/NET0131  & n1159 ;
  assign n6267 = ~n6265 & ~n6266 ;
  assign n6268 = ~n5028 & n6267 ;
  assign n6269 = ~\sub1_data_reg_reg[28]/NET0131  & n5028 ;
  assign n6270 = ~n6268 & ~n6269 ;
  assign n6271 = ~n5027 & ~n6270 ;
  assign n6272 = ~\mix1_data_o_reg_reg[28]/NET0131  & n5027 ;
  assign n6273 = ~n6271 & ~n6272 ;
  assign n6274 = n5026 & ~n6273 ;
  assign n6275 = ~\sub1_data_reg_reg[28]/NET0131  & ~n5026 ;
  assign n6276 = ~n6274 & ~n6275 ;
  assign n6277 = \state_reg/NET0131  & ~n6276 ;
  assign n6278 = ~\state_reg/NET0131  & n6267 ;
  assign n6279 = ~n6277 & ~n6278 ;
  assign n6281 = \key_i[28]_pad  & n6279 ;
  assign n6280 = ~\key_i[28]_pad  & ~n6279 ;
  assign n6282 = n933 & ~n6280 ;
  assign n6283 = ~n6281 & n6282 ;
  assign n6285 = ~\ks1_key_reg_reg[28]/NET0131  & ~n6279 ;
  assign n6286 = \ks1_key_reg_reg[28]/NET0131  & n6279 ;
  assign n6287 = ~n6285 & ~n6286 ;
  assign n6288 = n5053 & ~n6287 ;
  assign n6284 = ~\data_o[28]_pad  & ~n5053 ;
  assign n6289 = ~n933 & ~n6284 ;
  assign n6290 = ~n6288 & n6289 ;
  assign n6291 = ~n6283 & ~n6290 ;
  assign n6292 = ~\data_i[81]_pad  & ~n5029 ;
  assign n6293 = ~\mix1_data_o_reg_reg[81]/NET0131  & n5029 ;
  assign n6294 = ~n6292 & ~n6293 ;
  assign n6295 = ~n1159 & ~n6294 ;
  assign n6296 = ~\sub1_data_reg_reg[81]/NET0131  & n1159 ;
  assign n6297 = ~n6295 & ~n6296 ;
  assign n6298 = ~n5028 & ~n6297 ;
  assign n6299 = ~\sub1_data_reg_reg[81]/NET0131  & n5028 ;
  assign n6300 = ~n6298 & ~n6299 ;
  assign n6301 = ~n5027 & ~n6300 ;
  assign n6302 = ~\mix1_data_o_reg_reg[81]/NET0131  & n5027 ;
  assign n6303 = ~n6301 & ~n6302 ;
  assign n6304 = n5026 & ~n6303 ;
  assign n6305 = ~\sub1_data_reg_reg[81]/NET0131  & ~n5026 ;
  assign n6306 = ~n6304 & ~n6305 ;
  assign n6307 = \state_reg/NET0131  & ~n6306 ;
  assign n6308 = ~\state_reg/NET0131  & ~n6297 ;
  assign n6309 = ~n6307 & ~n6308 ;
  assign n6311 = \key_i[81]_pad  & n6309 ;
  assign n6310 = ~\key_i[81]_pad  & ~n6309 ;
  assign n6312 = n933 & ~n6310 ;
  assign n6313 = ~n6311 & n6312 ;
  assign n6315 = ~\ks1_key_reg_reg[81]/NET0131  & ~n6309 ;
  assign n6316 = \ks1_key_reg_reg[81]/NET0131  & n6309 ;
  assign n6317 = ~n6315 & ~n6316 ;
  assign n6318 = n5053 & ~n6317 ;
  assign n6314 = ~\data_o[81]_pad  & ~n5053 ;
  assign n6319 = ~n933 & ~n6314 ;
  assign n6320 = ~n6318 & n6319 ;
  assign n6321 = ~n6313 & ~n6320 ;
  assign n6322 = ~\data_i[82]_pad  & ~n5029 ;
  assign n6323 = ~\mix1_data_o_reg_reg[82]/NET0131  & n5029 ;
  assign n6324 = ~n6322 & ~n6323 ;
  assign n6325 = ~n1159 & ~n6324 ;
  assign n6326 = ~\sub1_data_reg_reg[82]/NET0131  & n1159 ;
  assign n6327 = ~n6325 & ~n6326 ;
  assign n6328 = ~n5028 & ~n6327 ;
  assign n6329 = ~\sub1_data_reg_reg[82]/NET0131  & n5028 ;
  assign n6330 = ~n6328 & ~n6329 ;
  assign n6331 = ~n5027 & ~n6330 ;
  assign n6332 = ~\mix1_data_o_reg_reg[82]/NET0131  & n5027 ;
  assign n6333 = ~n6331 & ~n6332 ;
  assign n6334 = n5026 & ~n6333 ;
  assign n6335 = ~\sub1_data_reg_reg[82]/NET0131  & ~n5026 ;
  assign n6336 = ~n6334 & ~n6335 ;
  assign n6337 = \state_reg/NET0131  & ~n6336 ;
  assign n6338 = ~\state_reg/NET0131  & ~n6327 ;
  assign n6339 = ~n6337 & ~n6338 ;
  assign n6341 = \key_i[82]_pad  & n6339 ;
  assign n6340 = ~\key_i[82]_pad  & ~n6339 ;
  assign n6342 = n933 & ~n6340 ;
  assign n6343 = ~n6341 & n6342 ;
  assign n6345 = ~\ks1_key_reg_reg[82]/NET0131  & ~n6339 ;
  assign n6346 = \ks1_key_reg_reg[82]/NET0131  & n6339 ;
  assign n6347 = ~n6345 & ~n6346 ;
  assign n6348 = n5053 & ~n6347 ;
  assign n6344 = ~\data_o[82]_pad  & ~n5053 ;
  assign n6349 = ~n933 & ~n6344 ;
  assign n6350 = ~n6348 & n6349 ;
  assign n6351 = ~n6343 & ~n6350 ;
  assign n6352 = \data_i[29]_pad  & ~n5029 ;
  assign n6353 = \mix1_data_o_reg_reg[29]/NET0131  & n5029 ;
  assign n6354 = ~n6352 & ~n6353 ;
  assign n6355 = ~n1159 & ~n6354 ;
  assign n6356 = \sub1_data_reg_reg[29]/NET0131  & n1159 ;
  assign n6357 = ~n6355 & ~n6356 ;
  assign n6358 = ~n5028 & n6357 ;
  assign n6359 = ~\sub1_data_reg_reg[29]/NET0131  & n5028 ;
  assign n6360 = ~n6358 & ~n6359 ;
  assign n6361 = ~n5027 & ~n6360 ;
  assign n6362 = ~\mix1_data_o_reg_reg[29]/NET0131  & n5027 ;
  assign n6363 = ~n6361 & ~n6362 ;
  assign n6364 = n5026 & ~n6363 ;
  assign n6365 = ~\sub1_data_reg_reg[29]/NET0131  & ~n5026 ;
  assign n6366 = ~n6364 & ~n6365 ;
  assign n6367 = \state_reg/NET0131  & ~n6366 ;
  assign n6368 = ~\state_reg/NET0131  & n6357 ;
  assign n6369 = ~n6367 & ~n6368 ;
  assign n6371 = \key_i[29]_pad  & n6369 ;
  assign n6370 = ~\key_i[29]_pad  & ~n6369 ;
  assign n6372 = n933 & ~n6370 ;
  assign n6373 = ~n6371 & n6372 ;
  assign n6375 = ~\ks1_key_reg_reg[29]/NET0131  & ~n6369 ;
  assign n6376 = \ks1_key_reg_reg[29]/NET0131  & n6369 ;
  assign n6377 = ~n6375 & ~n6376 ;
  assign n6378 = n5053 & ~n6377 ;
  assign n6374 = ~\data_o[29]_pad  & ~n5053 ;
  assign n6379 = ~n933 & ~n6374 ;
  assign n6380 = ~n6378 & n6379 ;
  assign n6381 = ~n6373 & ~n6380 ;
  assign n6382 = ~\data_i[83]_pad  & ~n5029 ;
  assign n6383 = ~\mix1_data_o_reg_reg[83]/NET0131  & n5029 ;
  assign n6384 = ~n6382 & ~n6383 ;
  assign n6385 = ~n1159 & ~n6384 ;
  assign n6386 = ~\sub1_data_reg_reg[83]/NET0131  & n1159 ;
  assign n6387 = ~n6385 & ~n6386 ;
  assign n6388 = ~n5028 & ~n6387 ;
  assign n6389 = ~\sub1_data_reg_reg[83]/NET0131  & n5028 ;
  assign n6390 = ~n6388 & ~n6389 ;
  assign n6391 = ~n5027 & ~n6390 ;
  assign n6392 = ~\mix1_data_o_reg_reg[83]/NET0131  & n5027 ;
  assign n6393 = ~n6391 & ~n6392 ;
  assign n6394 = n5026 & ~n6393 ;
  assign n6395 = ~\sub1_data_reg_reg[83]/NET0131  & ~n5026 ;
  assign n6396 = ~n6394 & ~n6395 ;
  assign n6397 = \state_reg/NET0131  & ~n6396 ;
  assign n6398 = ~\state_reg/NET0131  & ~n6387 ;
  assign n6399 = ~n6397 & ~n6398 ;
  assign n6401 = \key_i[83]_pad  & n6399 ;
  assign n6400 = ~\key_i[83]_pad  & ~n6399 ;
  assign n6402 = n933 & ~n6400 ;
  assign n6403 = ~n6401 & n6402 ;
  assign n6405 = ~\ks1_key_reg_reg[83]/NET0131  & ~n6399 ;
  assign n6406 = \ks1_key_reg_reg[83]/NET0131  & n6399 ;
  assign n6407 = ~n6405 & ~n6406 ;
  assign n6408 = n5053 & ~n6407 ;
  assign n6404 = ~\data_o[83]_pad  & ~n5053 ;
  assign n6409 = ~n933 & ~n6404 ;
  assign n6410 = ~n6408 & n6409 ;
  assign n6411 = ~n6403 & ~n6410 ;
  assign n6412 = ~\data_i[84]_pad  & ~n5029 ;
  assign n6413 = ~\mix1_data_o_reg_reg[84]/NET0131  & n5029 ;
  assign n6414 = ~n6412 & ~n6413 ;
  assign n6415 = ~n1159 & ~n6414 ;
  assign n6416 = ~\sub1_data_reg_reg[84]/NET0131  & n1159 ;
  assign n6417 = ~n6415 & ~n6416 ;
  assign n6418 = ~n5028 & ~n6417 ;
  assign n6419 = ~\sub1_data_reg_reg[84]/NET0131  & n5028 ;
  assign n6420 = ~n6418 & ~n6419 ;
  assign n6421 = ~n5027 & ~n6420 ;
  assign n6422 = ~\mix1_data_o_reg_reg[84]/NET0131  & n5027 ;
  assign n6423 = ~n6421 & ~n6422 ;
  assign n6424 = n5026 & ~n6423 ;
  assign n6425 = ~\sub1_data_reg_reg[84]/NET0131  & ~n5026 ;
  assign n6426 = ~n6424 & ~n6425 ;
  assign n6427 = \state_reg/NET0131  & ~n6426 ;
  assign n6428 = ~\state_reg/NET0131  & ~n6417 ;
  assign n6429 = ~n6427 & ~n6428 ;
  assign n6431 = \key_i[84]_pad  & n6429 ;
  assign n6430 = ~\key_i[84]_pad  & ~n6429 ;
  assign n6432 = n933 & ~n6430 ;
  assign n6433 = ~n6431 & n6432 ;
  assign n6435 = ~\ks1_key_reg_reg[84]/NET0131  & ~n6429 ;
  assign n6436 = \ks1_key_reg_reg[84]/NET0131  & n6429 ;
  assign n6437 = ~n6435 & ~n6436 ;
  assign n6438 = n5053 & ~n6437 ;
  assign n6434 = ~\data_o[84]_pad  & ~n5053 ;
  assign n6439 = ~n933 & ~n6434 ;
  assign n6440 = ~n6438 & n6439 ;
  assign n6441 = ~n6433 & ~n6440 ;
  assign n6442 = ~\data_i[118]_pad  & ~n5029 ;
  assign n6443 = ~\mix1_data_o_reg_reg[118]/NET0131  & n5029 ;
  assign n6444 = ~n6442 & ~n6443 ;
  assign n6445 = ~n1159 & ~n6444 ;
  assign n6446 = ~\sub1_data_reg_reg[118]/NET0131  & n1159 ;
  assign n6447 = ~n6445 & ~n6446 ;
  assign n6448 = ~n5028 & ~n6447 ;
  assign n6449 = ~\sub1_data_reg_reg[118]/NET0131  & n5028 ;
  assign n6450 = ~n6448 & ~n6449 ;
  assign n6451 = ~n5027 & ~n6450 ;
  assign n6452 = ~\mix1_data_o_reg_reg[118]/NET0131  & n5027 ;
  assign n6453 = ~n6451 & ~n6452 ;
  assign n6454 = n5026 & ~n6453 ;
  assign n6455 = ~\sub1_data_reg_reg[118]/NET0131  & ~n5026 ;
  assign n6456 = ~n6454 & ~n6455 ;
  assign n6457 = \state_reg/NET0131  & ~n6456 ;
  assign n6458 = ~\state_reg/NET0131  & ~n6447 ;
  assign n6459 = ~n6457 & ~n6458 ;
  assign n6461 = \key_i[118]_pad  & n6459 ;
  assign n6460 = ~\key_i[118]_pad  & ~n6459 ;
  assign n6462 = n933 & ~n6460 ;
  assign n6463 = ~n6461 & n6462 ;
  assign n6465 = ~\ks1_key_reg_reg[118]/NET0131  & ~n6459 ;
  assign n6466 = \ks1_key_reg_reg[118]/NET0131  & n6459 ;
  assign n6467 = ~n6465 & ~n6466 ;
  assign n6468 = n5053 & ~n6467 ;
  assign n6464 = ~\data_o[118]_pad  & ~n5053 ;
  assign n6469 = ~n933 & ~n6464 ;
  assign n6470 = ~n6468 & n6469 ;
  assign n6471 = ~n6463 & ~n6470 ;
  assign n6472 = \data_i[2]_pad  & ~n5029 ;
  assign n6473 = \mix1_data_o_reg_reg[2]/NET0131  & n5029 ;
  assign n6474 = ~n6472 & ~n6473 ;
  assign n6475 = ~n1159 & ~n6474 ;
  assign n6476 = \sub1_data_reg_reg[2]/NET0131  & n1159 ;
  assign n6477 = ~n6475 & ~n6476 ;
  assign n6478 = ~n5028 & n6477 ;
  assign n6479 = ~\sub1_data_reg_reg[2]/NET0131  & n5028 ;
  assign n6480 = ~n6478 & ~n6479 ;
  assign n6481 = ~n5027 & ~n6480 ;
  assign n6482 = ~\mix1_data_o_reg_reg[2]/NET0131  & n5027 ;
  assign n6483 = ~n6481 & ~n6482 ;
  assign n6484 = n5026 & ~n6483 ;
  assign n6485 = ~\sub1_data_reg_reg[2]/NET0131  & ~n5026 ;
  assign n6486 = ~n6484 & ~n6485 ;
  assign n6487 = \state_reg/NET0131  & ~n6486 ;
  assign n6488 = ~\state_reg/NET0131  & n6477 ;
  assign n6489 = ~n6487 & ~n6488 ;
  assign n6491 = \key_i[2]_pad  & n6489 ;
  assign n6490 = ~\key_i[2]_pad  & ~n6489 ;
  assign n6492 = n933 & ~n6490 ;
  assign n6493 = ~n6491 & n6492 ;
  assign n6495 = ~\ks1_key_reg_reg[2]/NET0131  & ~n6489 ;
  assign n6496 = \ks1_key_reg_reg[2]/NET0131  & n6489 ;
  assign n6497 = ~n6495 & ~n6496 ;
  assign n6498 = n5053 & ~n6497 ;
  assign n6494 = ~\data_o[2]_pad  & ~n5053 ;
  assign n6499 = ~n933 & ~n6494 ;
  assign n6500 = ~n6498 & n6499 ;
  assign n6501 = ~n6493 & ~n6500 ;
  assign n6502 = ~\data_i[85]_pad  & ~n5029 ;
  assign n6503 = ~\mix1_data_o_reg_reg[85]/NET0131  & n5029 ;
  assign n6504 = ~n6502 & ~n6503 ;
  assign n6505 = ~n1159 & ~n6504 ;
  assign n6506 = ~\sub1_data_reg_reg[85]/NET0131  & n1159 ;
  assign n6507 = ~n6505 & ~n6506 ;
  assign n6508 = ~n5028 & ~n6507 ;
  assign n6509 = ~\sub1_data_reg_reg[85]/NET0131  & n5028 ;
  assign n6510 = ~n6508 & ~n6509 ;
  assign n6511 = ~n5027 & ~n6510 ;
  assign n6512 = ~\mix1_data_o_reg_reg[85]/NET0131  & n5027 ;
  assign n6513 = ~n6511 & ~n6512 ;
  assign n6514 = n5026 & ~n6513 ;
  assign n6515 = ~\sub1_data_reg_reg[85]/NET0131  & ~n5026 ;
  assign n6516 = ~n6514 & ~n6515 ;
  assign n6517 = \state_reg/NET0131  & ~n6516 ;
  assign n6518 = ~\state_reg/NET0131  & ~n6507 ;
  assign n6519 = ~n6517 & ~n6518 ;
  assign n6521 = \key_i[85]_pad  & n6519 ;
  assign n6520 = ~\key_i[85]_pad  & ~n6519 ;
  assign n6522 = n933 & ~n6520 ;
  assign n6523 = ~n6521 & n6522 ;
  assign n6525 = ~\ks1_key_reg_reg[85]/NET0131  & ~n6519 ;
  assign n6526 = \ks1_key_reg_reg[85]/NET0131  & n6519 ;
  assign n6527 = ~n6525 & ~n6526 ;
  assign n6528 = n5053 & ~n6527 ;
  assign n6524 = ~\data_o[85]_pad  & ~n5053 ;
  assign n6529 = ~n933 & ~n6524 ;
  assign n6530 = ~n6528 & n6529 ;
  assign n6531 = ~n6523 & ~n6530 ;
  assign n6532 = \data_i[30]_pad  & ~n5029 ;
  assign n6533 = \mix1_data_o_reg_reg[30]/NET0131  & n5029 ;
  assign n6534 = ~n6532 & ~n6533 ;
  assign n6535 = ~n1159 & ~n6534 ;
  assign n6536 = \sub1_data_reg_reg[30]/NET0131  & n1159 ;
  assign n6537 = ~n6535 & ~n6536 ;
  assign n6538 = ~n5028 & n6537 ;
  assign n6539 = ~\sub1_data_reg_reg[30]/NET0131  & n5028 ;
  assign n6540 = ~n6538 & ~n6539 ;
  assign n6541 = ~n5027 & ~n6540 ;
  assign n6542 = ~\mix1_data_o_reg_reg[30]/NET0131  & n5027 ;
  assign n6543 = ~n6541 & ~n6542 ;
  assign n6544 = n5026 & ~n6543 ;
  assign n6545 = ~\sub1_data_reg_reg[30]/NET0131  & ~n5026 ;
  assign n6546 = ~n6544 & ~n6545 ;
  assign n6547 = \state_reg/NET0131  & ~n6546 ;
  assign n6548 = ~\state_reg/NET0131  & n6537 ;
  assign n6549 = ~n6547 & ~n6548 ;
  assign n6551 = \key_i[30]_pad  & n6549 ;
  assign n6550 = ~\key_i[30]_pad  & ~n6549 ;
  assign n6552 = n933 & ~n6550 ;
  assign n6553 = ~n6551 & n6552 ;
  assign n6555 = ~\ks1_key_reg_reg[30]/NET0131  & ~n6549 ;
  assign n6556 = \ks1_key_reg_reg[30]/NET0131  & n6549 ;
  assign n6557 = ~n6555 & ~n6556 ;
  assign n6558 = n5053 & ~n6557 ;
  assign n6554 = ~\data_o[30]_pad  & ~n5053 ;
  assign n6559 = ~n933 & ~n6554 ;
  assign n6560 = ~n6558 & n6559 ;
  assign n6561 = ~n6553 & ~n6560 ;
  assign n6562 = ~\data_i[86]_pad  & ~n5029 ;
  assign n6563 = ~\mix1_data_o_reg_reg[86]/NET0131  & n5029 ;
  assign n6564 = ~n6562 & ~n6563 ;
  assign n6565 = ~n1159 & ~n6564 ;
  assign n6566 = ~\sub1_data_reg_reg[86]/NET0131  & n1159 ;
  assign n6567 = ~n6565 & ~n6566 ;
  assign n6568 = ~n5028 & ~n6567 ;
  assign n6569 = ~\sub1_data_reg_reg[86]/NET0131  & n5028 ;
  assign n6570 = ~n6568 & ~n6569 ;
  assign n6571 = ~n5027 & ~n6570 ;
  assign n6572 = ~\mix1_data_o_reg_reg[86]/NET0131  & n5027 ;
  assign n6573 = ~n6571 & ~n6572 ;
  assign n6574 = n5026 & ~n6573 ;
  assign n6575 = ~\sub1_data_reg_reg[86]/NET0131  & ~n5026 ;
  assign n6576 = ~n6574 & ~n6575 ;
  assign n6577 = \state_reg/NET0131  & ~n6576 ;
  assign n6578 = ~\state_reg/NET0131  & ~n6567 ;
  assign n6579 = ~n6577 & ~n6578 ;
  assign n6581 = \key_i[86]_pad  & n6579 ;
  assign n6580 = ~\key_i[86]_pad  & ~n6579 ;
  assign n6582 = n933 & ~n6580 ;
  assign n6583 = ~n6581 & n6582 ;
  assign n6585 = ~\ks1_key_reg_reg[86]/NET0131  & ~n6579 ;
  assign n6586 = \ks1_key_reg_reg[86]/NET0131  & n6579 ;
  assign n6587 = ~n6585 & ~n6586 ;
  assign n6588 = n5053 & ~n6587 ;
  assign n6584 = ~\data_o[86]_pad  & ~n5053 ;
  assign n6589 = ~n933 & ~n6584 ;
  assign n6590 = ~n6588 & n6589 ;
  assign n6591 = ~n6583 & ~n6590 ;
  assign n6592 = ~\data_i[87]_pad  & ~n5029 ;
  assign n6593 = ~\mix1_data_o_reg_reg[87]/NET0131  & n5029 ;
  assign n6594 = ~n6592 & ~n6593 ;
  assign n6595 = ~n1159 & ~n6594 ;
  assign n6596 = ~\sub1_data_reg_reg[87]/NET0131  & n1159 ;
  assign n6597 = ~n6595 & ~n6596 ;
  assign n6598 = ~n5028 & ~n6597 ;
  assign n6599 = ~\sub1_data_reg_reg[87]/NET0131  & n5028 ;
  assign n6600 = ~n6598 & ~n6599 ;
  assign n6601 = ~n5027 & ~n6600 ;
  assign n6602 = ~\mix1_data_o_reg_reg[87]/NET0131  & n5027 ;
  assign n6603 = ~n6601 & ~n6602 ;
  assign n6604 = n5026 & ~n6603 ;
  assign n6605 = ~\sub1_data_reg_reg[87]/NET0131  & ~n5026 ;
  assign n6606 = ~n6604 & ~n6605 ;
  assign n6607 = \state_reg/NET0131  & ~n6606 ;
  assign n6608 = ~\state_reg/NET0131  & ~n6597 ;
  assign n6609 = ~n6607 & ~n6608 ;
  assign n6611 = \key_i[87]_pad  & n6609 ;
  assign n6610 = ~\key_i[87]_pad  & ~n6609 ;
  assign n6612 = n933 & ~n6610 ;
  assign n6613 = ~n6611 & n6612 ;
  assign n6615 = ~\ks1_key_reg_reg[87]/NET0131  & ~n6609 ;
  assign n6616 = \ks1_key_reg_reg[87]/NET0131  & n6609 ;
  assign n6617 = ~n6615 & ~n6616 ;
  assign n6618 = n5053 & ~n6617 ;
  assign n6614 = ~\data_o[87]_pad  & ~n5053 ;
  assign n6619 = ~n933 & ~n6614 ;
  assign n6620 = ~n6618 & n6619 ;
  assign n6621 = ~n6613 & ~n6620 ;
  assign n6622 = \data_i[31]_pad  & ~n5029 ;
  assign n6623 = \mix1_data_o_reg_reg[31]/NET0131  & n5029 ;
  assign n6624 = ~n6622 & ~n6623 ;
  assign n6625 = ~n1159 & ~n6624 ;
  assign n6626 = \sub1_data_reg_reg[31]/NET0131  & n1159 ;
  assign n6627 = ~n6625 & ~n6626 ;
  assign n6628 = ~n5028 & n6627 ;
  assign n6629 = ~\sub1_data_reg_reg[31]/NET0131  & n5028 ;
  assign n6630 = ~n6628 & ~n6629 ;
  assign n6631 = ~n5027 & ~n6630 ;
  assign n6632 = ~\mix1_data_o_reg_reg[31]/NET0131  & n5027 ;
  assign n6633 = ~n6631 & ~n6632 ;
  assign n6634 = n5026 & ~n6633 ;
  assign n6635 = ~\sub1_data_reg_reg[31]/NET0131  & ~n5026 ;
  assign n6636 = ~n6634 & ~n6635 ;
  assign n6637 = \state_reg/NET0131  & ~n6636 ;
  assign n6638 = ~\state_reg/NET0131  & n6627 ;
  assign n6639 = ~n6637 & ~n6638 ;
  assign n6641 = \key_i[31]_pad  & n6639 ;
  assign n6640 = ~\key_i[31]_pad  & ~n6639 ;
  assign n6642 = n933 & ~n6640 ;
  assign n6643 = ~n6641 & n6642 ;
  assign n6645 = ~\ks1_key_reg_reg[31]/NET0131  & ~n6639 ;
  assign n6646 = \ks1_key_reg_reg[31]/NET0131  & n6639 ;
  assign n6647 = ~n6645 & ~n6646 ;
  assign n6648 = n5053 & ~n6647 ;
  assign n6644 = ~\data_o[31]_pad  & ~n5053 ;
  assign n6649 = ~n933 & ~n6644 ;
  assign n6650 = ~n6648 & n6649 ;
  assign n6651 = ~n6643 & ~n6650 ;
  assign n6652 = \data_i[88]_pad  & ~n5029 ;
  assign n6653 = \mix1_data_o_reg_reg[88]/NET0131  & n5029 ;
  assign n6654 = ~n6652 & ~n6653 ;
  assign n6655 = ~n1159 & ~n6654 ;
  assign n6656 = \sub1_data_reg_reg[88]/NET0131  & n1159 ;
  assign n6657 = ~n6655 & ~n6656 ;
  assign n6658 = ~n5028 & n6657 ;
  assign n6659 = ~\sub1_data_reg_reg[88]/NET0131  & n5028 ;
  assign n6660 = ~n6658 & ~n6659 ;
  assign n6661 = ~n5027 & ~n6660 ;
  assign n6662 = ~\mix1_data_o_reg_reg[88]/NET0131  & n5027 ;
  assign n6663 = ~n6661 & ~n6662 ;
  assign n6664 = n5026 & ~n6663 ;
  assign n6665 = ~\sub1_data_reg_reg[88]/NET0131  & ~n5026 ;
  assign n6666 = ~n6664 & ~n6665 ;
  assign n6667 = \state_reg/NET0131  & ~n6666 ;
  assign n6668 = ~\state_reg/NET0131  & n6657 ;
  assign n6669 = ~n6667 & ~n6668 ;
  assign n6671 = \key_i[88]_pad  & n6669 ;
  assign n6670 = ~\key_i[88]_pad  & ~n6669 ;
  assign n6672 = n933 & ~n6670 ;
  assign n6673 = ~n6671 & n6672 ;
  assign n6675 = ~\ks1_key_reg_reg[88]/NET0131  & ~n6669 ;
  assign n6676 = \ks1_key_reg_reg[88]/NET0131  & n6669 ;
  assign n6677 = ~n6675 & ~n6676 ;
  assign n6678 = n5053 & ~n6677 ;
  assign n6674 = ~\data_o[88]_pad  & ~n5053 ;
  assign n6679 = ~n933 & ~n6674 ;
  assign n6680 = ~n6678 & n6679 ;
  assign n6681 = ~n6673 & ~n6680 ;
  assign n6682 = ~\data_i[119]_pad  & ~n5029 ;
  assign n6683 = ~\mix1_data_o_reg_reg[119]/NET0131  & n5029 ;
  assign n6684 = ~n6682 & ~n6683 ;
  assign n6685 = ~n1159 & ~n6684 ;
  assign n6686 = ~\sub1_data_reg_reg[119]/NET0131  & n1159 ;
  assign n6687 = ~n6685 & ~n6686 ;
  assign n6688 = ~n5028 & ~n6687 ;
  assign n6689 = ~\sub1_data_reg_reg[119]/NET0131  & n5028 ;
  assign n6690 = ~n6688 & ~n6689 ;
  assign n6691 = ~n5027 & ~n6690 ;
  assign n6692 = ~\mix1_data_o_reg_reg[119]/NET0131  & n5027 ;
  assign n6693 = ~n6691 & ~n6692 ;
  assign n6694 = n5026 & ~n6693 ;
  assign n6695 = ~\sub1_data_reg_reg[119]/NET0131  & ~n5026 ;
  assign n6696 = ~n6694 & ~n6695 ;
  assign n6697 = \state_reg/NET0131  & ~n6696 ;
  assign n6698 = ~\state_reg/NET0131  & ~n6687 ;
  assign n6699 = ~n6697 & ~n6698 ;
  assign n6701 = \key_i[119]_pad  & n6699 ;
  assign n6700 = ~\key_i[119]_pad  & ~n6699 ;
  assign n6702 = n933 & ~n6700 ;
  assign n6703 = ~n6701 & n6702 ;
  assign n6705 = ~\ks1_key_reg_reg[119]/NET0131  & ~n6699 ;
  assign n6706 = \ks1_key_reg_reg[119]/NET0131  & n6699 ;
  assign n6707 = ~n6705 & ~n6706 ;
  assign n6708 = n5053 & ~n6707 ;
  assign n6704 = ~\data_o[119]_pad  & ~n5053 ;
  assign n6709 = ~n933 & ~n6704 ;
  assign n6710 = ~n6708 & n6709 ;
  assign n6711 = ~n6703 & ~n6710 ;
  assign n6712 = \data_i[89]_pad  & ~n5029 ;
  assign n6713 = \mix1_data_o_reg_reg[89]/NET0131  & n5029 ;
  assign n6714 = ~n6712 & ~n6713 ;
  assign n6715 = ~n1159 & ~n6714 ;
  assign n6716 = \sub1_data_reg_reg[89]/NET0131  & n1159 ;
  assign n6717 = ~n6715 & ~n6716 ;
  assign n6718 = ~n5028 & n6717 ;
  assign n6719 = ~\sub1_data_reg_reg[89]/NET0131  & n5028 ;
  assign n6720 = ~n6718 & ~n6719 ;
  assign n6721 = ~n5027 & ~n6720 ;
  assign n6722 = ~\mix1_data_o_reg_reg[89]/NET0131  & n5027 ;
  assign n6723 = ~n6721 & ~n6722 ;
  assign n6724 = n5026 & ~n6723 ;
  assign n6725 = ~\sub1_data_reg_reg[89]/NET0131  & ~n5026 ;
  assign n6726 = ~n6724 & ~n6725 ;
  assign n6727 = \state_reg/NET0131  & ~n6726 ;
  assign n6728 = ~\state_reg/NET0131  & n6717 ;
  assign n6729 = ~n6727 & ~n6728 ;
  assign n6731 = \key_i[89]_pad  & n6729 ;
  assign n6730 = ~\key_i[89]_pad  & ~n6729 ;
  assign n6732 = n933 & ~n6730 ;
  assign n6733 = ~n6731 & n6732 ;
  assign n6735 = ~\ks1_key_reg_reg[89]/NET0131  & ~n6729 ;
  assign n6736 = \ks1_key_reg_reg[89]/NET0131  & n6729 ;
  assign n6737 = ~n6735 & ~n6736 ;
  assign n6738 = n5053 & ~n6737 ;
  assign n6734 = ~\data_o[89]_pad  & ~n5053 ;
  assign n6739 = ~n933 & ~n6734 ;
  assign n6740 = ~n6738 & n6739 ;
  assign n6741 = ~n6733 & ~n6740 ;
  assign n6742 = \data_i[8]_pad  & ~n5029 ;
  assign n6743 = \mix1_data_o_reg_reg[8]/NET0131  & n5029 ;
  assign n6744 = ~n6742 & ~n6743 ;
  assign n6745 = ~n1159 & ~n6744 ;
  assign n6746 = \sub1_data_reg_reg[8]/NET0131  & n1159 ;
  assign n6747 = ~n6745 & ~n6746 ;
  assign n6748 = ~n5028 & n6747 ;
  assign n6749 = ~\sub1_data_reg_reg[8]/NET0131  & n5028 ;
  assign n6750 = ~n6748 & ~n6749 ;
  assign n6751 = ~n5027 & ~n6750 ;
  assign n6752 = ~\mix1_data_o_reg_reg[8]/NET0131  & n5027 ;
  assign n6753 = ~n6751 & ~n6752 ;
  assign n6754 = n5026 & ~n6753 ;
  assign n6755 = ~\sub1_data_reg_reg[8]/NET0131  & ~n5026 ;
  assign n6756 = ~n6754 & ~n6755 ;
  assign n6757 = \state_reg/NET0131  & ~n6756 ;
  assign n6758 = ~\state_reg/NET0131  & n6747 ;
  assign n6759 = ~n6757 & ~n6758 ;
  assign n6761 = \key_i[8]_pad  & n6759 ;
  assign n6760 = ~\key_i[8]_pad  & ~n6759 ;
  assign n6762 = n933 & ~n6760 ;
  assign n6763 = ~n6761 & n6762 ;
  assign n6765 = ~\ks1_key_reg_reg[8]/NET0131  & ~n6759 ;
  assign n6766 = \ks1_key_reg_reg[8]/NET0131  & n6759 ;
  assign n6767 = ~n6765 & ~n6766 ;
  assign n6768 = n5053 & ~n6767 ;
  assign n6764 = ~\data_o[8]_pad  & ~n5053 ;
  assign n6769 = ~n933 & ~n6764 ;
  assign n6770 = ~n6768 & n6769 ;
  assign n6771 = ~n6763 & ~n6770 ;
  assign n6772 = ~\data_i[32]_pad  & ~n5029 ;
  assign n6773 = ~\mix1_data_o_reg_reg[32]/NET0131  & n5029 ;
  assign n6774 = ~n6772 & ~n6773 ;
  assign n6775 = ~n1159 & ~n6774 ;
  assign n6776 = ~\sub1_data_reg_reg[32]/NET0131  & n1159 ;
  assign n6777 = ~n6775 & ~n6776 ;
  assign n6778 = ~n5028 & ~n6777 ;
  assign n6779 = ~\sub1_data_reg_reg[32]/NET0131  & n5028 ;
  assign n6780 = ~n6778 & ~n6779 ;
  assign n6781 = ~n5027 & ~n6780 ;
  assign n6782 = ~\mix1_data_o_reg_reg[32]/NET0131  & n5027 ;
  assign n6783 = ~n6781 & ~n6782 ;
  assign n6784 = n5026 & ~n6783 ;
  assign n6785 = ~\sub1_data_reg_reg[32]/NET0131  & ~n5026 ;
  assign n6786 = ~n6784 & ~n6785 ;
  assign n6787 = \state_reg/NET0131  & ~n6786 ;
  assign n6788 = ~\state_reg/NET0131  & ~n6777 ;
  assign n6789 = ~n6787 & ~n6788 ;
  assign n6791 = \key_i[32]_pad  & n6789 ;
  assign n6790 = ~\key_i[32]_pad  & ~n6789 ;
  assign n6792 = n933 & ~n6790 ;
  assign n6793 = ~n6791 & n6792 ;
  assign n6795 = ~\ks1_key_reg_reg[32]/NET0131  & ~n6789 ;
  assign n6796 = \ks1_key_reg_reg[32]/NET0131  & n6789 ;
  assign n6797 = ~n6795 & ~n6796 ;
  assign n6798 = n5053 & ~n6797 ;
  assign n6794 = ~\data_o[32]_pad  & ~n5053 ;
  assign n6799 = ~n933 & ~n6794 ;
  assign n6800 = ~n6798 & n6799 ;
  assign n6801 = ~n6793 & ~n6800 ;
  assign n6802 = \data_i[104]_pad  & ~n5029 ;
  assign n6803 = \mix1_data_o_reg_reg[104]/NET0131  & n5029 ;
  assign n6804 = ~n6802 & ~n6803 ;
  assign n6805 = ~n1159 & ~n6804 ;
  assign n6806 = \sub1_data_reg_reg[104]/NET0131  & n1159 ;
  assign n6807 = ~n6805 & ~n6806 ;
  assign n6808 = ~n5028 & n6807 ;
  assign n6809 = ~\sub1_data_reg_reg[104]/NET0131  & n5028 ;
  assign n6810 = ~n6808 & ~n6809 ;
  assign n6811 = ~n5027 & ~n6810 ;
  assign n6812 = ~\mix1_data_o_reg_reg[104]/NET0131  & n5027 ;
  assign n6813 = ~n6811 & ~n6812 ;
  assign n6814 = n5026 & ~n6813 ;
  assign n6815 = ~\sub1_data_reg_reg[104]/NET0131  & ~n5026 ;
  assign n6816 = ~n6814 & ~n6815 ;
  assign n6817 = \state_reg/NET0131  & ~n6816 ;
  assign n6818 = ~\state_reg/NET0131  & n6807 ;
  assign n6819 = ~n6817 & ~n6818 ;
  assign n6821 = \key_i[104]_pad  & n6819 ;
  assign n6820 = ~\key_i[104]_pad  & ~n6819 ;
  assign n6822 = n933 & ~n6820 ;
  assign n6823 = ~n6821 & n6822 ;
  assign n6825 = ~\ks1_key_reg_reg[104]/NET0131  & ~n6819 ;
  assign n6826 = \ks1_key_reg_reg[104]/NET0131  & n6819 ;
  assign n6827 = ~n6825 & ~n6826 ;
  assign n6828 = n5053 & ~n6827 ;
  assign n6824 = ~\data_o[104]_pad  & ~n5053 ;
  assign n6829 = ~n933 & ~n6824 ;
  assign n6830 = ~n6828 & n6829 ;
  assign n6831 = ~n6823 & ~n6830 ;
  assign n6832 = \data_i[90]_pad  & ~n5029 ;
  assign n6833 = \mix1_data_o_reg_reg[90]/NET0131  & n5029 ;
  assign n6834 = ~n6832 & ~n6833 ;
  assign n6835 = ~n1159 & ~n6834 ;
  assign n6836 = \sub1_data_reg_reg[90]/NET0131  & n1159 ;
  assign n6837 = ~n6835 & ~n6836 ;
  assign n6838 = ~n5028 & n6837 ;
  assign n6839 = ~\sub1_data_reg_reg[90]/NET0131  & n5028 ;
  assign n6840 = ~n6838 & ~n6839 ;
  assign n6841 = ~n5027 & ~n6840 ;
  assign n6842 = ~\mix1_data_o_reg_reg[90]/NET0131  & n5027 ;
  assign n6843 = ~n6841 & ~n6842 ;
  assign n6844 = n5026 & ~n6843 ;
  assign n6845 = ~\sub1_data_reg_reg[90]/NET0131  & ~n5026 ;
  assign n6846 = ~n6844 & ~n6845 ;
  assign n6847 = \state_reg/NET0131  & ~n6846 ;
  assign n6848 = ~\state_reg/NET0131  & n6837 ;
  assign n6849 = ~n6847 & ~n6848 ;
  assign n6851 = \key_i[90]_pad  & n6849 ;
  assign n6850 = ~\key_i[90]_pad  & ~n6849 ;
  assign n6852 = n933 & ~n6850 ;
  assign n6853 = ~n6851 & n6852 ;
  assign n6855 = ~\ks1_key_reg_reg[90]/NET0131  & ~n6849 ;
  assign n6856 = \ks1_key_reg_reg[90]/NET0131  & n6849 ;
  assign n6857 = ~n6855 & ~n6856 ;
  assign n6858 = n5053 & ~n6857 ;
  assign n6854 = ~\data_o[90]_pad  & ~n5053 ;
  assign n6859 = ~n933 & ~n6854 ;
  assign n6860 = ~n6858 & n6859 ;
  assign n6861 = ~n6853 & ~n6860 ;
  assign n6862 = \data_i[105]_pad  & ~n5029 ;
  assign n6863 = \mix1_data_o_reg_reg[105]/NET0131  & n5029 ;
  assign n6864 = ~n6862 & ~n6863 ;
  assign n6865 = ~n1159 & ~n6864 ;
  assign n6866 = \sub1_data_reg_reg[105]/NET0131  & n1159 ;
  assign n6867 = ~n6865 & ~n6866 ;
  assign n6868 = ~n5028 & n6867 ;
  assign n6869 = ~\sub1_data_reg_reg[105]/NET0131  & n5028 ;
  assign n6870 = ~n6868 & ~n6869 ;
  assign n6871 = ~n5027 & ~n6870 ;
  assign n6872 = ~\mix1_data_o_reg_reg[105]/NET0131  & n5027 ;
  assign n6873 = ~n6871 & ~n6872 ;
  assign n6874 = n5026 & ~n6873 ;
  assign n6875 = ~\sub1_data_reg_reg[105]/NET0131  & ~n5026 ;
  assign n6876 = ~n6874 & ~n6875 ;
  assign n6877 = \state_reg/NET0131  & ~n6876 ;
  assign n6878 = ~\state_reg/NET0131  & n6867 ;
  assign n6879 = ~n6877 & ~n6878 ;
  assign n6881 = \key_i[105]_pad  & n6879 ;
  assign n6880 = ~\key_i[105]_pad  & ~n6879 ;
  assign n6882 = n933 & ~n6880 ;
  assign n6883 = ~n6881 & n6882 ;
  assign n6885 = ~\ks1_key_reg_reg[105]/NET0131  & ~n6879 ;
  assign n6886 = \ks1_key_reg_reg[105]/NET0131  & n6879 ;
  assign n6887 = ~n6885 & ~n6886 ;
  assign n6888 = n5053 & ~n6887 ;
  assign n6884 = ~\data_o[105]_pad  & ~n5053 ;
  assign n6889 = ~n933 & ~n6884 ;
  assign n6890 = ~n6888 & n6889 ;
  assign n6891 = ~n6883 & ~n6890 ;
  assign n6892 = \data_i[91]_pad  & ~n5029 ;
  assign n6893 = \mix1_data_o_reg_reg[91]/NET0131  & n5029 ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6895 = ~n1159 & ~n6894 ;
  assign n6896 = \sub1_data_reg_reg[91]/NET0131  & n1159 ;
  assign n6897 = ~n6895 & ~n6896 ;
  assign n6898 = ~n5028 & n6897 ;
  assign n6899 = ~\sub1_data_reg_reg[91]/NET0131  & n5028 ;
  assign n6900 = ~n6898 & ~n6899 ;
  assign n6901 = ~n5027 & ~n6900 ;
  assign n6902 = ~\mix1_data_o_reg_reg[91]/NET0131  & n5027 ;
  assign n6903 = ~n6901 & ~n6902 ;
  assign n6904 = n5026 & ~n6903 ;
  assign n6905 = ~\sub1_data_reg_reg[91]/NET0131  & ~n5026 ;
  assign n6906 = ~n6904 & ~n6905 ;
  assign n6907 = \state_reg/NET0131  & ~n6906 ;
  assign n6908 = ~\state_reg/NET0131  & n6897 ;
  assign n6909 = ~n6907 & ~n6908 ;
  assign n6911 = \key_i[91]_pad  & n6909 ;
  assign n6910 = ~\key_i[91]_pad  & ~n6909 ;
  assign n6912 = n933 & ~n6910 ;
  assign n6913 = ~n6911 & n6912 ;
  assign n6915 = ~\ks1_key_reg_reg[91]/NET0131  & ~n6909 ;
  assign n6916 = \ks1_key_reg_reg[91]/NET0131  & n6909 ;
  assign n6917 = ~n6915 & ~n6916 ;
  assign n6918 = n5053 & ~n6917 ;
  assign n6914 = ~\data_o[91]_pad  & ~n5053 ;
  assign n6919 = ~n933 & ~n6914 ;
  assign n6920 = ~n6918 & n6919 ;
  assign n6921 = ~n6913 & ~n6920 ;
  assign n6922 = ~\data_i[33]_pad  & ~n5029 ;
  assign n6923 = ~\mix1_data_o_reg_reg[33]/NET0131  & n5029 ;
  assign n6924 = ~n6922 & ~n6923 ;
  assign n6925 = ~n1159 & ~n6924 ;
  assign n6926 = ~\sub1_data_reg_reg[33]/NET0131  & n1159 ;
  assign n6927 = ~n6925 & ~n6926 ;
  assign n6928 = ~n5028 & ~n6927 ;
  assign n6929 = ~\sub1_data_reg_reg[33]/NET0131  & n5028 ;
  assign n6930 = ~n6928 & ~n6929 ;
  assign n6931 = ~n5027 & ~n6930 ;
  assign n6932 = ~\mix1_data_o_reg_reg[33]/NET0131  & n5027 ;
  assign n6933 = ~n6931 & ~n6932 ;
  assign n6934 = n5026 & ~n6933 ;
  assign n6935 = ~\sub1_data_reg_reg[33]/NET0131  & ~n5026 ;
  assign n6936 = ~n6934 & ~n6935 ;
  assign n6937 = \state_reg/NET0131  & ~n6936 ;
  assign n6938 = ~\state_reg/NET0131  & ~n6927 ;
  assign n6939 = ~n6937 & ~n6938 ;
  assign n6941 = \key_i[33]_pad  & n6939 ;
  assign n6940 = ~\key_i[33]_pad  & ~n6939 ;
  assign n6942 = n933 & ~n6940 ;
  assign n6943 = ~n6941 & n6942 ;
  assign n6945 = ~\ks1_key_reg_reg[33]/NET0131  & ~n6939 ;
  assign n6946 = \ks1_key_reg_reg[33]/NET0131  & n6939 ;
  assign n6947 = ~n6945 & ~n6946 ;
  assign n6948 = n5053 & ~n6947 ;
  assign n6944 = ~\data_o[33]_pad  & ~n5053 ;
  assign n6949 = ~n933 & ~n6944 ;
  assign n6950 = ~n6948 & n6949 ;
  assign n6951 = ~n6943 & ~n6950 ;
  assign n6952 = \data_i[11]_pad  & ~n5029 ;
  assign n6953 = \mix1_data_o_reg_reg[11]/NET0131  & n5029 ;
  assign n6954 = ~n6952 & ~n6953 ;
  assign n6955 = ~n1159 & ~n6954 ;
  assign n6956 = \sub1_data_reg_reg[11]/NET0131  & n1159 ;
  assign n6957 = ~n6955 & ~n6956 ;
  assign n6958 = ~n5028 & n6957 ;
  assign n6959 = ~\sub1_data_reg_reg[11]/NET0131  & n5028 ;
  assign n6960 = ~n6958 & ~n6959 ;
  assign n6961 = ~n5027 & ~n6960 ;
  assign n6962 = ~\mix1_data_o_reg_reg[11]/NET0131  & n5027 ;
  assign n6963 = ~n6961 & ~n6962 ;
  assign n6964 = n5026 & ~n6963 ;
  assign n6965 = ~\sub1_data_reg_reg[11]/NET0131  & ~n5026 ;
  assign n6966 = ~n6964 & ~n6965 ;
  assign n6967 = \state_reg/NET0131  & ~n6966 ;
  assign n6968 = ~\state_reg/NET0131  & n6957 ;
  assign n6969 = ~n6967 & ~n6968 ;
  assign n6971 = \key_i[11]_pad  & n6969 ;
  assign n6970 = ~\key_i[11]_pad  & ~n6969 ;
  assign n6972 = n933 & ~n6970 ;
  assign n6973 = ~n6971 & n6972 ;
  assign n6975 = ~\ks1_key_reg_reg[11]/NET0131  & ~n6969 ;
  assign n6976 = \ks1_key_reg_reg[11]/NET0131  & n6969 ;
  assign n6977 = ~n6975 & ~n6976 ;
  assign n6978 = n5053 & ~n6977 ;
  assign n6974 = ~\data_o[11]_pad  & ~n5053 ;
  assign n6979 = ~n933 & ~n6974 ;
  assign n6980 = ~n6978 & n6979 ;
  assign n6981 = ~n6973 & ~n6980 ;
  assign n6982 = \data_i[92]_pad  & ~n5029 ;
  assign n6983 = \mix1_data_o_reg_reg[92]/NET0131  & n5029 ;
  assign n6984 = ~n6982 & ~n6983 ;
  assign n6985 = ~n1159 & ~n6984 ;
  assign n6986 = \sub1_data_reg_reg[92]/NET0131  & n1159 ;
  assign n6987 = ~n6985 & ~n6986 ;
  assign n6988 = ~n5028 & n6987 ;
  assign n6989 = ~\sub1_data_reg_reg[92]/NET0131  & n5028 ;
  assign n6990 = ~n6988 & ~n6989 ;
  assign n6991 = ~n5027 & ~n6990 ;
  assign n6992 = ~\mix1_data_o_reg_reg[92]/NET0131  & n5027 ;
  assign n6993 = ~n6991 & ~n6992 ;
  assign n6994 = n5026 & ~n6993 ;
  assign n6995 = ~\sub1_data_reg_reg[92]/NET0131  & ~n5026 ;
  assign n6996 = ~n6994 & ~n6995 ;
  assign n6997 = \state_reg/NET0131  & ~n6996 ;
  assign n6998 = ~\state_reg/NET0131  & n6987 ;
  assign n6999 = ~n6997 & ~n6998 ;
  assign n7001 = \key_i[92]_pad  & n6999 ;
  assign n7000 = ~\key_i[92]_pad  & ~n6999 ;
  assign n7002 = n933 & ~n7000 ;
  assign n7003 = ~n7001 & n7002 ;
  assign n7005 = ~\ks1_key_reg_reg[92]/NET0131  & ~n6999 ;
  assign n7006 = \ks1_key_reg_reg[92]/NET0131  & n6999 ;
  assign n7007 = ~n7005 & ~n7006 ;
  assign n7008 = n5053 & ~n7007 ;
  assign n7004 = ~\data_o[92]_pad  & ~n5053 ;
  assign n7009 = ~n933 & ~n7004 ;
  assign n7010 = ~n7008 & n7009 ;
  assign n7011 = ~n7003 & ~n7010 ;
  assign n7012 = \data_i[93]_pad  & ~n5029 ;
  assign n7013 = \mix1_data_o_reg_reg[93]/NET0131  & n5029 ;
  assign n7014 = ~n7012 & ~n7013 ;
  assign n7015 = ~n1159 & ~n7014 ;
  assign n7016 = \sub1_data_reg_reg[93]/NET0131  & n1159 ;
  assign n7017 = ~n7015 & ~n7016 ;
  assign n7018 = ~n5028 & n7017 ;
  assign n7019 = ~\sub1_data_reg_reg[93]/NET0131  & n5028 ;
  assign n7020 = ~n7018 & ~n7019 ;
  assign n7021 = ~n5027 & ~n7020 ;
  assign n7022 = ~\mix1_data_o_reg_reg[93]/NET0131  & n5027 ;
  assign n7023 = ~n7021 & ~n7022 ;
  assign n7024 = n5026 & ~n7023 ;
  assign n7025 = ~\sub1_data_reg_reg[93]/NET0131  & ~n5026 ;
  assign n7026 = ~n7024 & ~n7025 ;
  assign n7027 = \state_reg/NET0131  & ~n7026 ;
  assign n7028 = ~\state_reg/NET0131  & n7017 ;
  assign n7029 = ~n7027 & ~n7028 ;
  assign n7031 = \key_i[93]_pad  & n7029 ;
  assign n7030 = ~\key_i[93]_pad  & ~n7029 ;
  assign n7032 = n933 & ~n7030 ;
  assign n7033 = ~n7031 & n7032 ;
  assign n7035 = ~\ks1_key_reg_reg[93]/NET0131  & ~n7029 ;
  assign n7036 = \ks1_key_reg_reg[93]/NET0131  & n7029 ;
  assign n7037 = ~n7035 & ~n7036 ;
  assign n7038 = n5053 & ~n7037 ;
  assign n7034 = ~\data_o[93]_pad  & ~n5053 ;
  assign n7039 = ~n933 & ~n7034 ;
  assign n7040 = ~n7038 & n7039 ;
  assign n7041 = ~n7033 & ~n7040 ;
  assign n7042 = ~\data_i[34]_pad  & ~n5029 ;
  assign n7043 = ~\mix1_data_o_reg_reg[34]/NET0131  & n5029 ;
  assign n7044 = ~n7042 & ~n7043 ;
  assign n7045 = ~n1159 & ~n7044 ;
  assign n7046 = ~\sub1_data_reg_reg[34]/NET0131  & n1159 ;
  assign n7047 = ~n7045 & ~n7046 ;
  assign n7048 = ~n5028 & ~n7047 ;
  assign n7049 = ~\sub1_data_reg_reg[34]/NET0131  & n5028 ;
  assign n7050 = ~n7048 & ~n7049 ;
  assign n7051 = ~n5027 & ~n7050 ;
  assign n7052 = ~\mix1_data_o_reg_reg[34]/NET0131  & n5027 ;
  assign n7053 = ~n7051 & ~n7052 ;
  assign n7054 = n5026 & ~n7053 ;
  assign n7055 = ~\sub1_data_reg_reg[34]/NET0131  & ~n5026 ;
  assign n7056 = ~n7054 & ~n7055 ;
  assign n7057 = \state_reg/NET0131  & ~n7056 ;
  assign n7058 = ~\state_reg/NET0131  & ~n7047 ;
  assign n7059 = ~n7057 & ~n7058 ;
  assign n7061 = \key_i[34]_pad  & n7059 ;
  assign n7060 = ~\key_i[34]_pad  & ~n7059 ;
  assign n7062 = n933 & ~n7060 ;
  assign n7063 = ~n7061 & n7062 ;
  assign n7065 = ~\ks1_key_reg_reg[34]/NET0131  & ~n7059 ;
  assign n7066 = \ks1_key_reg_reg[34]/NET0131  & n7059 ;
  assign n7067 = ~n7065 & ~n7066 ;
  assign n7068 = n5053 & ~n7067 ;
  assign n7064 = ~\data_o[34]_pad  & ~n5053 ;
  assign n7069 = ~n933 & ~n7064 ;
  assign n7070 = ~n7068 & n7069 ;
  assign n7071 = ~n7063 & ~n7070 ;
  assign n7072 = \data_i[94]_pad  & ~n5029 ;
  assign n7073 = \mix1_data_o_reg_reg[94]/NET0131  & n5029 ;
  assign n7074 = ~n7072 & ~n7073 ;
  assign n7075 = ~n1159 & ~n7074 ;
  assign n7076 = \sub1_data_reg_reg[94]/NET0131  & n1159 ;
  assign n7077 = ~n7075 & ~n7076 ;
  assign n7078 = ~n5028 & n7077 ;
  assign n7079 = ~\sub1_data_reg_reg[94]/NET0131  & n5028 ;
  assign n7080 = ~n7078 & ~n7079 ;
  assign n7081 = ~n5027 & ~n7080 ;
  assign n7082 = ~\mix1_data_o_reg_reg[94]/NET0131  & n5027 ;
  assign n7083 = ~n7081 & ~n7082 ;
  assign n7084 = n5026 & ~n7083 ;
  assign n7085 = ~\sub1_data_reg_reg[94]/NET0131  & ~n5026 ;
  assign n7086 = ~n7084 & ~n7085 ;
  assign n7087 = \state_reg/NET0131  & ~n7086 ;
  assign n7088 = ~\state_reg/NET0131  & n7077 ;
  assign n7089 = ~n7087 & ~n7088 ;
  assign n7091 = \key_i[94]_pad  & n7089 ;
  assign n7090 = ~\key_i[94]_pad  & ~n7089 ;
  assign n7092 = n933 & ~n7090 ;
  assign n7093 = ~n7091 & n7092 ;
  assign n7095 = ~\ks1_key_reg_reg[94]/NET0131  & ~n7089 ;
  assign n7096 = \ks1_key_reg_reg[94]/NET0131  & n7089 ;
  assign n7097 = ~n7095 & ~n7096 ;
  assign n7098 = n5053 & ~n7097 ;
  assign n7094 = ~\data_o[94]_pad  & ~n5053 ;
  assign n7099 = ~n933 & ~n7094 ;
  assign n7100 = ~n7098 & n7099 ;
  assign n7101 = ~n7093 & ~n7100 ;
  assign n7102 = \data_i[95]_pad  & ~n5029 ;
  assign n7103 = \mix1_data_o_reg_reg[95]/NET0131  & n5029 ;
  assign n7104 = ~n7102 & ~n7103 ;
  assign n7105 = ~n1159 & ~n7104 ;
  assign n7106 = \sub1_data_reg_reg[95]/NET0131  & n1159 ;
  assign n7107 = ~n7105 & ~n7106 ;
  assign n7108 = ~n5028 & n7107 ;
  assign n7109 = ~\sub1_data_reg_reg[95]/NET0131  & n5028 ;
  assign n7110 = ~n7108 & ~n7109 ;
  assign n7111 = ~n5027 & ~n7110 ;
  assign n7112 = ~\mix1_data_o_reg_reg[95]/NET0131  & n5027 ;
  assign n7113 = ~n7111 & ~n7112 ;
  assign n7114 = n5026 & ~n7113 ;
  assign n7115 = ~\sub1_data_reg_reg[95]/NET0131  & ~n5026 ;
  assign n7116 = ~n7114 & ~n7115 ;
  assign n7117 = \state_reg/NET0131  & ~n7116 ;
  assign n7118 = ~\state_reg/NET0131  & n7107 ;
  assign n7119 = ~n7117 & ~n7118 ;
  assign n7121 = \key_i[95]_pad  & n7119 ;
  assign n7120 = ~\key_i[95]_pad  & ~n7119 ;
  assign n7122 = n933 & ~n7120 ;
  assign n7123 = ~n7121 & n7122 ;
  assign n7125 = ~\ks1_key_reg_reg[95]/NET0131  & ~n7119 ;
  assign n7126 = \ks1_key_reg_reg[95]/NET0131  & n7119 ;
  assign n7127 = ~n7125 & ~n7126 ;
  assign n7128 = n5053 & ~n7127 ;
  assign n7124 = ~\data_o[95]_pad  & ~n5053 ;
  assign n7129 = ~n933 & ~n7124 ;
  assign n7130 = ~n7128 & n7129 ;
  assign n7131 = ~n7123 & ~n7130 ;
  assign n7132 = ~\data_i[35]_pad  & ~n5029 ;
  assign n7133 = ~\mix1_data_o_reg_reg[35]/NET0131  & n5029 ;
  assign n7134 = ~n7132 & ~n7133 ;
  assign n7135 = ~n1159 & ~n7134 ;
  assign n7136 = ~\sub1_data_reg_reg[35]/NET0131  & n1159 ;
  assign n7137 = ~n7135 & ~n7136 ;
  assign n7138 = ~n5028 & ~n7137 ;
  assign n7139 = ~\sub1_data_reg_reg[35]/NET0131  & n5028 ;
  assign n7140 = ~n7138 & ~n7139 ;
  assign n7141 = ~n5027 & ~n7140 ;
  assign n7142 = ~\mix1_data_o_reg_reg[35]/NET0131  & n5027 ;
  assign n7143 = ~n7141 & ~n7142 ;
  assign n7144 = n5026 & ~n7143 ;
  assign n7145 = ~\sub1_data_reg_reg[35]/NET0131  & ~n5026 ;
  assign n7146 = ~n7144 & ~n7145 ;
  assign n7147 = \state_reg/NET0131  & ~n7146 ;
  assign n7148 = ~\state_reg/NET0131  & ~n7137 ;
  assign n7149 = ~n7147 & ~n7148 ;
  assign n7151 = \key_i[35]_pad  & n7149 ;
  assign n7150 = ~\key_i[35]_pad  & ~n7149 ;
  assign n7152 = n933 & ~n7150 ;
  assign n7153 = ~n7151 & n7152 ;
  assign n7155 = ~\ks1_key_reg_reg[35]/NET0131  & ~n7149 ;
  assign n7156 = \ks1_key_reg_reg[35]/NET0131  & n7149 ;
  assign n7157 = ~n7155 & ~n7156 ;
  assign n7158 = n5053 & ~n7157 ;
  assign n7154 = ~\data_o[35]_pad  & ~n5053 ;
  assign n7159 = ~n933 & ~n7154 ;
  assign n7160 = ~n7158 & n7159 ;
  assign n7161 = ~n7153 & ~n7160 ;
  assign n7162 = ~n1159 & ~n5029 ;
  assign n7163 = \data_i[96]_pad  & n7162 ;
  assign n7164 = \mix1_data_o_reg_reg[96]/NET0131  & n5029 ;
  assign n7165 = \sub1_data_reg_reg[96]/NET0131  & n1159 ;
  assign n7166 = ~n7164 & ~n7165 ;
  assign n7167 = ~n7163 & n7166 ;
  assign n7168 = ~n5028 & ~n7167 ;
  assign n7169 = \sub1_ready_o_reg/NET0131  & n2692 ;
  assign n7170 = ~n5027 & ~n7169 ;
  assign n7171 = ~n7168 & n7170 ;
  assign n7172 = ~\mix1_data_o_reg_reg[96]/NET0131  & n5027 ;
  assign n7173 = ~n7171 & ~n7172 ;
  assign n7174 = n5026 & ~n7173 ;
  assign n7175 = ~\sub1_data_reg_reg[96]/NET0131  & ~n5026 ;
  assign n7176 = ~n7174 & ~n7175 ;
  assign n7177 = \state_reg/NET0131  & ~n7176 ;
  assign n7178 = ~\state_reg/NET0131  & n7167 ;
  assign n7179 = ~n7177 & ~n7178 ;
  assign n7181 = \key_i[96]_pad  & n7179 ;
  assign n7180 = ~\key_i[96]_pad  & ~n7179 ;
  assign n7182 = n933 & ~n7180 ;
  assign n7183 = ~n7181 & n7182 ;
  assign n7185 = ~\ks1_key_reg_reg[96]/NET0131  & ~n7179 ;
  assign n7186 = \ks1_key_reg_reg[96]/NET0131  & n7179 ;
  assign n7187 = ~n7185 & ~n7186 ;
  assign n7188 = n5053 & ~n7187 ;
  assign n7184 = ~\data_o[96]_pad  & ~n5053 ;
  assign n7189 = ~n933 & ~n7184 ;
  assign n7190 = ~n7188 & n7189 ;
  assign n7191 = ~n7183 & ~n7190 ;
  assign n7192 = \data_i[120]_pad  & ~n5029 ;
  assign n7193 = \mix1_data_o_reg_reg[120]/NET0131  & n5029 ;
  assign n7194 = ~n7192 & ~n7193 ;
  assign n7195 = ~n1159 & ~n7194 ;
  assign n7196 = \sub1_data_reg_reg[120]/NET0131  & n1159 ;
  assign n7197 = ~n7195 & ~n7196 ;
  assign n7198 = ~n5028 & n7197 ;
  assign n7199 = ~\sub1_data_reg_reg[120]/NET0131  & n5028 ;
  assign n7200 = ~n7198 & ~n7199 ;
  assign n7201 = ~n5027 & ~n7200 ;
  assign n7202 = ~\mix1_data_o_reg_reg[120]/NET0131  & n5027 ;
  assign n7203 = ~n7201 & ~n7202 ;
  assign n7204 = n5026 & ~n7203 ;
  assign n7205 = ~\sub1_data_reg_reg[120]/NET0131  & ~n5026 ;
  assign n7206 = ~n7204 & ~n7205 ;
  assign n7207 = \state_reg/NET0131  & ~n7206 ;
  assign n7208 = ~\state_reg/NET0131  & n7197 ;
  assign n7209 = ~n7207 & ~n7208 ;
  assign n7211 = \key_i[120]_pad  & n7209 ;
  assign n7210 = ~\key_i[120]_pad  & ~n7209 ;
  assign n7212 = n933 & ~n7210 ;
  assign n7213 = ~n7211 & n7212 ;
  assign n7215 = ~\ks1_key_reg_reg[120]/NET0131  & ~n7209 ;
  assign n7216 = \ks1_key_reg_reg[120]/NET0131  & n7209 ;
  assign n7217 = ~n7215 & ~n7216 ;
  assign n7218 = n5053 & ~n7217 ;
  assign n7214 = ~\data_o[120]_pad  & ~n5053 ;
  assign n7219 = ~n933 & ~n7214 ;
  assign n7220 = ~n7218 & n7219 ;
  assign n7221 = ~n7213 & ~n7220 ;
  assign n7222 = ~\data_i[36]_pad  & ~n5029 ;
  assign n7223 = ~\mix1_data_o_reg_reg[36]/NET0131  & n5029 ;
  assign n7224 = ~n7222 & ~n7223 ;
  assign n7225 = ~n1159 & ~n7224 ;
  assign n7226 = ~\sub1_data_reg_reg[36]/NET0131  & n1159 ;
  assign n7227 = ~n7225 & ~n7226 ;
  assign n7228 = ~n5028 & ~n7227 ;
  assign n7229 = ~\sub1_data_reg_reg[36]/NET0131  & n5028 ;
  assign n7230 = ~n7228 & ~n7229 ;
  assign n7231 = ~n5027 & ~n7230 ;
  assign n7232 = ~\mix1_data_o_reg_reg[36]/NET0131  & n5027 ;
  assign n7233 = ~n7231 & ~n7232 ;
  assign n7234 = n5026 & ~n7233 ;
  assign n7235 = ~\sub1_data_reg_reg[36]/NET0131  & ~n5026 ;
  assign n7236 = ~n7234 & ~n7235 ;
  assign n7237 = \state_reg/NET0131  & ~n7236 ;
  assign n7238 = ~\state_reg/NET0131  & ~n7227 ;
  assign n7239 = ~n7237 & ~n7238 ;
  assign n7241 = \key_i[36]_pad  & n7239 ;
  assign n7240 = ~\key_i[36]_pad  & ~n7239 ;
  assign n7242 = n933 & ~n7240 ;
  assign n7243 = ~n7241 & n7242 ;
  assign n7245 = ~\ks1_key_reg_reg[36]/NET0131  & ~n7239 ;
  assign n7246 = \ks1_key_reg_reg[36]/NET0131  & n7239 ;
  assign n7247 = ~n7245 & ~n7246 ;
  assign n7248 = n5053 & ~n7247 ;
  assign n7244 = ~\data_o[36]_pad  & ~n5053 ;
  assign n7249 = ~n933 & ~n7244 ;
  assign n7250 = ~n7248 & n7249 ;
  assign n7251 = ~n7243 & ~n7250 ;
  assign n7252 = \data_i[97]_pad  & n7162 ;
  assign n7253 = \mix1_data_o_reg_reg[97]/NET0131  & n5029 ;
  assign n7254 = \sub1_data_reg_reg[97]/NET0131  & n1159 ;
  assign n7255 = ~n7253 & ~n7254 ;
  assign n7256 = ~n7252 & n7255 ;
  assign n7257 = ~n5028 & ~n7256 ;
  assign n7258 = \sub1_ready_o_reg/NET0131  & n3295 ;
  assign n7259 = ~n5027 & ~n7258 ;
  assign n7260 = ~n7257 & n7259 ;
  assign n7261 = ~\mix1_data_o_reg_reg[97]/NET0131  & n5027 ;
  assign n7262 = ~n7260 & ~n7261 ;
  assign n7263 = n5026 & ~n7262 ;
  assign n7264 = ~\sub1_data_reg_reg[97]/NET0131  & ~n5026 ;
  assign n7265 = ~n7263 & ~n7264 ;
  assign n7266 = \state_reg/NET0131  & ~n7265 ;
  assign n7267 = ~\state_reg/NET0131  & n7256 ;
  assign n7268 = ~n7266 & ~n7267 ;
  assign n7270 = \key_i[97]_pad  & n7268 ;
  assign n7269 = ~\key_i[97]_pad  & ~n7268 ;
  assign n7271 = n933 & ~n7269 ;
  assign n7272 = ~n7270 & n7271 ;
  assign n7274 = ~\ks1_key_reg_reg[97]/NET0131  & ~n7268 ;
  assign n7275 = \ks1_key_reg_reg[97]/NET0131  & n7268 ;
  assign n7276 = ~n7274 & ~n7275 ;
  assign n7277 = n5053 & ~n7276 ;
  assign n7273 = ~\data_o[97]_pad  & ~n5053 ;
  assign n7278 = ~n933 & ~n7273 ;
  assign n7279 = ~n7277 & n7278 ;
  assign n7280 = ~n7272 & ~n7279 ;
  assign n7281 = ~\data_i[98]_pad  & ~n5029 ;
  assign n7282 = ~\mix1_data_o_reg_reg[98]/NET0131  & n5029 ;
  assign n7283 = ~n7281 & ~n7282 ;
  assign n7284 = ~n1159 & ~n7283 ;
  assign n7285 = ~\sub1_data_reg_reg[98]/NET0131  & n1159 ;
  assign n7286 = ~n7284 & ~n7285 ;
  assign n7287 = ~n5028 & ~n7286 ;
  assign n7288 = ~\sub1_data_reg_reg[98]/NET0131  & n5028 ;
  assign n7289 = ~n7287 & ~n7288 ;
  assign n7290 = ~n5027 & ~n7289 ;
  assign n7291 = ~\mix1_data_o_reg_reg[98]/NET0131  & n5027 ;
  assign n7292 = ~n7290 & ~n7291 ;
  assign n7293 = n5026 & ~n7292 ;
  assign n7294 = ~\sub1_data_reg_reg[98]/NET0131  & ~n5026 ;
  assign n7295 = ~n7293 & ~n7294 ;
  assign n7296 = \state_reg/NET0131  & ~n7295 ;
  assign n7297 = ~\state_reg/NET0131  & ~n7286 ;
  assign n7298 = ~n7296 & ~n7297 ;
  assign n7300 = \key_i[98]_pad  & n7298 ;
  assign n7299 = ~\key_i[98]_pad  & ~n7298 ;
  assign n7301 = n933 & ~n7299 ;
  assign n7302 = ~n7300 & n7301 ;
  assign n7304 = ~\ks1_key_reg_reg[98]/NET0131  & ~n7298 ;
  assign n7305 = \ks1_key_reg_reg[98]/NET0131  & n7298 ;
  assign n7306 = ~n7304 & ~n7305 ;
  assign n7307 = n5053 & ~n7306 ;
  assign n7303 = ~\data_o[98]_pad  & ~n5053 ;
  assign n7308 = ~n933 & ~n7303 ;
  assign n7309 = ~n7307 & n7308 ;
  assign n7310 = ~n7302 & ~n7309 ;
  assign n7311 = ~\data_i[37]_pad  & ~n5029 ;
  assign n7312 = ~\mix1_data_o_reg_reg[37]/NET0131  & n5029 ;
  assign n7313 = ~n7311 & ~n7312 ;
  assign n7314 = ~n1159 & ~n7313 ;
  assign n7315 = ~\sub1_data_reg_reg[37]/NET0131  & n1159 ;
  assign n7316 = ~n7314 & ~n7315 ;
  assign n7317 = ~n5028 & ~n7316 ;
  assign n7318 = ~\sub1_data_reg_reg[37]/NET0131  & n5028 ;
  assign n7319 = ~n7317 & ~n7318 ;
  assign n7320 = ~n5027 & ~n7319 ;
  assign n7321 = ~\mix1_data_o_reg_reg[37]/NET0131  & n5027 ;
  assign n7322 = ~n7320 & ~n7321 ;
  assign n7323 = n5026 & ~n7322 ;
  assign n7324 = ~\sub1_data_reg_reg[37]/NET0131  & ~n5026 ;
  assign n7325 = ~n7323 & ~n7324 ;
  assign n7326 = \state_reg/NET0131  & ~n7325 ;
  assign n7327 = ~\state_reg/NET0131  & ~n7316 ;
  assign n7328 = ~n7326 & ~n7327 ;
  assign n7330 = \key_i[37]_pad  & n7328 ;
  assign n7329 = ~\key_i[37]_pad  & ~n7328 ;
  assign n7331 = n933 & ~n7329 ;
  assign n7332 = ~n7330 & n7331 ;
  assign n7334 = ~\ks1_key_reg_reg[37]/NET0131  & ~n7328 ;
  assign n7335 = \ks1_key_reg_reg[37]/NET0131  & n7328 ;
  assign n7336 = ~n7334 & ~n7335 ;
  assign n7337 = n5053 & ~n7336 ;
  assign n7333 = ~\data_o[37]_pad  & ~n5053 ;
  assign n7338 = ~n933 & ~n7333 ;
  assign n7339 = ~n7337 & n7338 ;
  assign n7340 = ~n7332 & ~n7339 ;
  assign n7341 = ~\data_i[99]_pad  & ~n5029 ;
  assign n7342 = ~\mix1_data_o_reg_reg[99]/NET0131  & n5029 ;
  assign n7343 = ~n7341 & ~n7342 ;
  assign n7344 = ~n1159 & ~n7343 ;
  assign n7345 = ~\sub1_data_reg_reg[99]/NET0131  & n1159 ;
  assign n7346 = ~n7344 & ~n7345 ;
  assign n7347 = ~n5028 & ~n7346 ;
  assign n7348 = ~\sub1_data_reg_reg[99]/NET0131  & n5028 ;
  assign n7349 = ~n7347 & ~n7348 ;
  assign n7350 = ~n5027 & ~n7349 ;
  assign n7351 = ~\mix1_data_o_reg_reg[99]/NET0131  & n5027 ;
  assign n7352 = ~n7350 & ~n7351 ;
  assign n7353 = n5026 & ~n7352 ;
  assign n7354 = ~\sub1_data_reg_reg[99]/NET0131  & ~n5026 ;
  assign n7355 = ~n7353 & ~n7354 ;
  assign n7356 = \state_reg/NET0131  & ~n7355 ;
  assign n7357 = ~\state_reg/NET0131  & ~n7346 ;
  assign n7358 = ~n7356 & ~n7357 ;
  assign n7360 = \key_i[99]_pad  & n7358 ;
  assign n7359 = ~\key_i[99]_pad  & ~n7358 ;
  assign n7361 = n933 & ~n7359 ;
  assign n7362 = ~n7360 & n7361 ;
  assign n7364 = ~\ks1_key_reg_reg[99]/NET0131  & ~n7358 ;
  assign n7365 = \ks1_key_reg_reg[99]/NET0131  & n7358 ;
  assign n7366 = ~n7364 & ~n7365 ;
  assign n7367 = n5053 & ~n7366 ;
  assign n7363 = ~\data_o[99]_pad  & ~n5053 ;
  assign n7368 = ~n933 & ~n7363 ;
  assign n7369 = ~n7367 & n7368 ;
  assign n7370 = ~n7362 & ~n7369 ;
  assign n7371 = \data_i[121]_pad  & ~n5029 ;
  assign n7372 = \mix1_data_o_reg_reg[121]/NET0131  & n5029 ;
  assign n7373 = ~n7371 & ~n7372 ;
  assign n7374 = ~n1159 & ~n7373 ;
  assign n7375 = \sub1_data_reg_reg[121]/NET0131  & n1159 ;
  assign n7376 = ~n7374 & ~n7375 ;
  assign n7377 = ~n5028 & n7376 ;
  assign n7378 = ~\sub1_data_reg_reg[121]/NET0131  & n5028 ;
  assign n7379 = ~n7377 & ~n7378 ;
  assign n7380 = ~n5027 & ~n7379 ;
  assign n7381 = ~\mix1_data_o_reg_reg[121]/NET0131  & n5027 ;
  assign n7382 = ~n7380 & ~n7381 ;
  assign n7383 = n5026 & ~n7382 ;
  assign n7384 = ~\sub1_data_reg_reg[121]/NET0131  & ~n5026 ;
  assign n7385 = ~n7383 & ~n7384 ;
  assign n7386 = \state_reg/NET0131  & ~n7385 ;
  assign n7387 = ~\state_reg/NET0131  & n7376 ;
  assign n7388 = ~n7386 & ~n7387 ;
  assign n7390 = \key_i[121]_pad  & n7388 ;
  assign n7389 = ~\key_i[121]_pad  & ~n7388 ;
  assign n7391 = n933 & ~n7389 ;
  assign n7392 = ~n7390 & n7391 ;
  assign n7394 = ~\ks1_key_reg_reg[121]/NET0131  & ~n7388 ;
  assign n7395 = \ks1_key_reg_reg[121]/NET0131  & n7388 ;
  assign n7396 = ~n7394 & ~n7395 ;
  assign n7397 = n5053 & ~n7396 ;
  assign n7393 = ~\data_o[121]_pad  & ~n5053 ;
  assign n7398 = ~n933 & ~n7393 ;
  assign n7399 = ~n7397 & n7398 ;
  assign n7400 = ~n7392 & ~n7399 ;
  assign n7401 = \data_i[9]_pad  & ~n5029 ;
  assign n7402 = \mix1_data_o_reg_reg[9]/NET0131  & n5029 ;
  assign n7403 = ~n7401 & ~n7402 ;
  assign n7404 = ~n1159 & ~n7403 ;
  assign n7405 = \sub1_data_reg_reg[9]/NET0131  & n1159 ;
  assign n7406 = ~n7404 & ~n7405 ;
  assign n7407 = ~n5028 & n7406 ;
  assign n7408 = ~\sub1_data_reg_reg[9]/NET0131  & n5028 ;
  assign n7409 = ~n7407 & ~n7408 ;
  assign n7410 = ~n5027 & ~n7409 ;
  assign n7411 = ~\mix1_data_o_reg_reg[9]/NET0131  & n5027 ;
  assign n7412 = ~n7410 & ~n7411 ;
  assign n7413 = n5026 & ~n7412 ;
  assign n7414 = ~\sub1_data_reg_reg[9]/NET0131  & ~n5026 ;
  assign n7415 = ~n7413 & ~n7414 ;
  assign n7416 = \state_reg/NET0131  & ~n7415 ;
  assign n7417 = ~\state_reg/NET0131  & n7406 ;
  assign n7418 = ~n7416 & ~n7417 ;
  assign n7420 = \key_i[9]_pad  & n7418 ;
  assign n7419 = ~\key_i[9]_pad  & ~n7418 ;
  assign n7421 = n933 & ~n7419 ;
  assign n7422 = ~n7420 & n7421 ;
  assign n7424 = ~\ks1_key_reg_reg[9]/NET0131  & ~n7418 ;
  assign n7425 = \ks1_key_reg_reg[9]/NET0131  & n7418 ;
  assign n7426 = ~n7424 & ~n7425 ;
  assign n7427 = n5053 & ~n7426 ;
  assign n7423 = ~\data_o[9]_pad  & ~n5053 ;
  assign n7428 = ~n933 & ~n7423 ;
  assign n7429 = ~n7427 & n7428 ;
  assign n7430 = ~n7422 & ~n7429 ;
  assign n7431 = ~\data_i[38]_pad  & ~n5029 ;
  assign n7432 = ~\mix1_data_o_reg_reg[38]/NET0131  & n5029 ;
  assign n7433 = ~n7431 & ~n7432 ;
  assign n7434 = ~n1159 & ~n7433 ;
  assign n7435 = ~\sub1_data_reg_reg[38]/NET0131  & n1159 ;
  assign n7436 = ~n7434 & ~n7435 ;
  assign n7437 = ~n5028 & ~n7436 ;
  assign n7438 = ~\sub1_data_reg_reg[38]/NET0131  & n5028 ;
  assign n7439 = ~n7437 & ~n7438 ;
  assign n7440 = ~n5027 & ~n7439 ;
  assign n7441 = ~\mix1_data_o_reg_reg[38]/NET0131  & n5027 ;
  assign n7442 = ~n7440 & ~n7441 ;
  assign n7443 = n5026 & ~n7442 ;
  assign n7444 = ~\sub1_data_reg_reg[38]/NET0131  & ~n5026 ;
  assign n7445 = ~n7443 & ~n7444 ;
  assign n7446 = \state_reg/NET0131  & ~n7445 ;
  assign n7447 = ~\state_reg/NET0131  & ~n7436 ;
  assign n7448 = ~n7446 & ~n7447 ;
  assign n7450 = \key_i[38]_pad  & n7448 ;
  assign n7449 = ~\key_i[38]_pad  & ~n7448 ;
  assign n7451 = n933 & ~n7449 ;
  assign n7452 = ~n7450 & n7451 ;
  assign n7454 = ~\ks1_key_reg_reg[38]/NET0131  & ~n7448 ;
  assign n7455 = \ks1_key_reg_reg[38]/NET0131  & n7448 ;
  assign n7456 = ~n7454 & ~n7455 ;
  assign n7457 = n5053 & ~n7456 ;
  assign n7453 = ~\data_o[38]_pad  & ~n5053 ;
  assign n7458 = ~n933 & ~n7453 ;
  assign n7459 = ~n7457 & n7458 ;
  assign n7460 = ~n7452 & ~n7459 ;
  assign n7461 = \data_i[106]_pad  & ~n5029 ;
  assign n7462 = \mix1_data_o_reg_reg[106]/NET0131  & n5029 ;
  assign n7463 = ~n7461 & ~n7462 ;
  assign n7464 = ~n1159 & ~n7463 ;
  assign n7465 = \sub1_data_reg_reg[106]/NET0131  & n1159 ;
  assign n7466 = ~n7464 & ~n7465 ;
  assign n7467 = ~n5028 & n7466 ;
  assign n7468 = ~\sub1_data_reg_reg[106]/NET0131  & n5028 ;
  assign n7469 = ~n7467 & ~n7468 ;
  assign n7470 = ~n5027 & ~n7469 ;
  assign n7471 = ~\mix1_data_o_reg_reg[106]/NET0131  & n5027 ;
  assign n7472 = ~n7470 & ~n7471 ;
  assign n7473 = n5026 & ~n7472 ;
  assign n7474 = ~\sub1_data_reg_reg[106]/NET0131  & ~n5026 ;
  assign n7475 = ~n7473 & ~n7474 ;
  assign n7476 = \state_reg/NET0131  & ~n7475 ;
  assign n7477 = ~\state_reg/NET0131  & n7466 ;
  assign n7478 = ~n7476 & ~n7477 ;
  assign n7480 = \key_i[106]_pad  & n7478 ;
  assign n7479 = ~\key_i[106]_pad  & ~n7478 ;
  assign n7481 = n933 & ~n7479 ;
  assign n7482 = ~n7480 & n7481 ;
  assign n7484 = ~\ks1_key_reg_reg[106]/NET0131  & ~n7478 ;
  assign n7485 = \ks1_key_reg_reg[106]/NET0131  & n7478 ;
  assign n7486 = ~n7484 & ~n7485 ;
  assign n7487 = n5053 & ~n7486 ;
  assign n7483 = ~\data_o[106]_pad  & ~n5053 ;
  assign n7488 = ~n933 & ~n7483 ;
  assign n7489 = ~n7487 & n7488 ;
  assign n7490 = ~n7482 & ~n7489 ;
  assign n7491 = \data_i[122]_pad  & ~n5029 ;
  assign n7492 = \mix1_data_o_reg_reg[122]/NET0131  & n5029 ;
  assign n7493 = ~n7491 & ~n7492 ;
  assign n7494 = ~n1159 & ~n7493 ;
  assign n7495 = \sub1_data_reg_reg[122]/NET0131  & n1159 ;
  assign n7496 = ~n7494 & ~n7495 ;
  assign n7497 = ~n5028 & n7496 ;
  assign n7498 = ~\sub1_data_reg_reg[122]/NET0131  & n5028 ;
  assign n7499 = ~n7497 & ~n7498 ;
  assign n7500 = ~n5027 & ~n7499 ;
  assign n7501 = ~\mix1_data_o_reg_reg[122]/NET0131  & n5027 ;
  assign n7502 = ~n7500 & ~n7501 ;
  assign n7503 = n5026 & ~n7502 ;
  assign n7504 = ~\sub1_data_reg_reg[122]/NET0131  & ~n5026 ;
  assign n7505 = ~n7503 & ~n7504 ;
  assign n7506 = \state_reg/NET0131  & ~n7505 ;
  assign n7507 = ~\state_reg/NET0131  & n7496 ;
  assign n7508 = ~n7506 & ~n7507 ;
  assign n7510 = \key_i[122]_pad  & n7508 ;
  assign n7509 = ~\key_i[122]_pad  & ~n7508 ;
  assign n7511 = n933 & ~n7509 ;
  assign n7512 = ~n7510 & n7511 ;
  assign n7514 = ~\ks1_key_reg_reg[122]/NET0131  & ~n7508 ;
  assign n7515 = \ks1_key_reg_reg[122]/NET0131  & n7508 ;
  assign n7516 = ~n7514 & ~n7515 ;
  assign n7517 = n5053 & ~n7516 ;
  assign n7513 = ~\data_o[122]_pad  & ~n5053 ;
  assign n7518 = ~n933 & ~n7513 ;
  assign n7519 = ~n7517 & n7518 ;
  assign n7520 = ~n7512 & ~n7519 ;
  assign n7521 = ~\data_i[39]_pad  & ~n5029 ;
  assign n7522 = ~\mix1_data_o_reg_reg[39]/NET0131  & n5029 ;
  assign n7523 = ~n7521 & ~n7522 ;
  assign n7524 = ~n1159 & ~n7523 ;
  assign n7525 = ~\sub1_data_reg_reg[39]/NET0131  & n1159 ;
  assign n7526 = ~n7524 & ~n7525 ;
  assign n7527 = ~n5028 & ~n7526 ;
  assign n7528 = ~\sub1_data_reg_reg[39]/NET0131  & n5028 ;
  assign n7529 = ~n7527 & ~n7528 ;
  assign n7530 = ~n5027 & ~n7529 ;
  assign n7531 = ~\mix1_data_o_reg_reg[39]/NET0131  & n5027 ;
  assign n7532 = ~n7530 & ~n7531 ;
  assign n7533 = n5026 & ~n7532 ;
  assign n7534 = ~\sub1_data_reg_reg[39]/NET0131  & ~n5026 ;
  assign n7535 = ~n7533 & ~n7534 ;
  assign n7536 = \state_reg/NET0131  & ~n7535 ;
  assign n7537 = ~\state_reg/NET0131  & ~n7526 ;
  assign n7538 = ~n7536 & ~n7537 ;
  assign n7540 = \key_i[39]_pad  & n7538 ;
  assign n7539 = ~\key_i[39]_pad  & ~n7538 ;
  assign n7541 = n933 & ~n7539 ;
  assign n7542 = ~n7540 & n7541 ;
  assign n7544 = ~\ks1_key_reg_reg[39]/NET0131  & ~n7538 ;
  assign n7545 = \ks1_key_reg_reg[39]/NET0131  & n7538 ;
  assign n7546 = ~n7544 & ~n7545 ;
  assign n7547 = n5053 & ~n7546 ;
  assign n7543 = ~\data_o[39]_pad  & ~n5053 ;
  assign n7548 = ~n933 & ~n7543 ;
  assign n7549 = ~n7547 & n7548 ;
  assign n7550 = ~n7542 & ~n7549 ;
  assign n7551 = \data_i[3]_pad  & ~n5029 ;
  assign n7552 = \mix1_data_o_reg_reg[3]/NET0131  & n5029 ;
  assign n7553 = ~n7551 & ~n7552 ;
  assign n7554 = ~n1159 & ~n7553 ;
  assign n7555 = \sub1_data_reg_reg[3]/NET0131  & n1159 ;
  assign n7556 = ~n7554 & ~n7555 ;
  assign n7557 = ~n5028 & n7556 ;
  assign n7558 = ~\sub1_data_reg_reg[3]/NET0131  & n5028 ;
  assign n7559 = ~n7557 & ~n7558 ;
  assign n7560 = ~n5027 & ~n7559 ;
  assign n7561 = ~\mix1_data_o_reg_reg[3]/NET0131  & n5027 ;
  assign n7562 = ~n7560 & ~n7561 ;
  assign n7563 = n5026 & ~n7562 ;
  assign n7564 = ~\sub1_data_reg_reg[3]/NET0131  & ~n5026 ;
  assign n7565 = ~n7563 & ~n7564 ;
  assign n7566 = \state_reg/NET0131  & ~n7565 ;
  assign n7567 = ~\state_reg/NET0131  & n7556 ;
  assign n7568 = ~n7566 & ~n7567 ;
  assign n7570 = \key_i[3]_pad  & n7568 ;
  assign n7569 = ~\key_i[3]_pad  & ~n7568 ;
  assign n7571 = n933 & ~n7569 ;
  assign n7572 = ~n7570 & n7571 ;
  assign n7574 = ~\ks1_key_reg_reg[3]/NET0131  & ~n7568 ;
  assign n7575 = \ks1_key_reg_reg[3]/NET0131  & n7568 ;
  assign n7576 = ~n7574 & ~n7575 ;
  assign n7577 = n5053 & ~n7576 ;
  assign n7573 = ~\data_o[3]_pad  & ~n5053 ;
  assign n7578 = ~n933 & ~n7573 ;
  assign n7579 = ~n7577 & n7578 ;
  assign n7580 = ~n7572 & ~n7579 ;
  assign n7581 = \data_i[0]_pad  & ~n5029 ;
  assign n7582 = \mix1_data_o_reg_reg[0]/NET0131  & n5029 ;
  assign n7583 = ~n7581 & ~n7582 ;
  assign n7584 = ~n1159 & ~n7583 ;
  assign n7585 = \sub1_data_reg_reg[0]/NET0131  & n1159 ;
  assign n7586 = ~n7584 & ~n7585 ;
  assign n7587 = ~n5028 & n7586 ;
  assign n7588 = ~\sub1_data_reg_reg[0]/NET0131  & n5028 ;
  assign n7589 = ~n7587 & ~n7588 ;
  assign n7590 = ~n5027 & ~n7589 ;
  assign n7591 = ~\mix1_data_o_reg_reg[0]/NET0131  & n5027 ;
  assign n7592 = ~n7590 & ~n7591 ;
  assign n7593 = n5026 & ~n7592 ;
  assign n7594 = ~\sub1_data_reg_reg[0]/NET0131  & ~n5026 ;
  assign n7595 = ~n7593 & ~n7594 ;
  assign n7596 = \state_reg/NET0131  & ~n7595 ;
  assign n7597 = ~\state_reg/NET0131  & n7586 ;
  assign n7598 = ~n7596 & ~n7597 ;
  assign n7600 = \key_i[0]_pad  & n7598 ;
  assign n7599 = ~\key_i[0]_pad  & ~n7598 ;
  assign n7601 = n933 & ~n7599 ;
  assign n7602 = ~n7600 & n7601 ;
  assign n7604 = ~\ks1_key_reg_reg[0]/NET0131  & ~n7598 ;
  assign n7605 = \ks1_key_reg_reg[0]/NET0131  & n7598 ;
  assign n7606 = ~n7604 & ~n7605 ;
  assign n7607 = n5053 & ~n7606 ;
  assign n7603 = ~\data_o[0]_pad  & ~n5053 ;
  assign n7608 = ~n933 & ~n7603 ;
  assign n7609 = ~n7607 & n7608 ;
  assign n7610 = ~n7602 & ~n7609 ;
  assign n7611 = \data_i[40]_pad  & ~n5029 ;
  assign n7612 = \mix1_data_o_reg_reg[40]/NET0131  & n5029 ;
  assign n7613 = ~n7611 & ~n7612 ;
  assign n7614 = ~n1159 & ~n7613 ;
  assign n7615 = \sub1_data_reg_reg[40]/NET0131  & n1159 ;
  assign n7616 = ~n7614 & ~n7615 ;
  assign n7617 = ~n5028 & n7616 ;
  assign n7618 = ~\sub1_data_reg_reg[40]/NET0131  & n5028 ;
  assign n7619 = ~n7617 & ~n7618 ;
  assign n7620 = ~n5027 & ~n7619 ;
  assign n7621 = ~\mix1_data_o_reg_reg[40]/NET0131  & n5027 ;
  assign n7622 = ~n7620 & ~n7621 ;
  assign n7623 = n5026 & ~n7622 ;
  assign n7624 = ~\sub1_data_reg_reg[40]/NET0131  & ~n5026 ;
  assign n7625 = ~n7623 & ~n7624 ;
  assign n7626 = \state_reg/NET0131  & ~n7625 ;
  assign n7627 = ~\state_reg/NET0131  & n7616 ;
  assign n7628 = ~n7626 & ~n7627 ;
  assign n7630 = \key_i[40]_pad  & n7628 ;
  assign n7629 = ~\key_i[40]_pad  & ~n7628 ;
  assign n7631 = n933 & ~n7629 ;
  assign n7632 = ~n7630 & n7631 ;
  assign n7634 = ~\ks1_key_reg_reg[40]/P0002  & ~n7628 ;
  assign n7635 = \ks1_key_reg_reg[40]/P0002  & n7628 ;
  assign n7636 = ~n7634 & ~n7635 ;
  assign n7637 = n5053 & ~n7636 ;
  assign n7633 = ~\data_o[40]_pad  & ~n5053 ;
  assign n7638 = ~n933 & ~n7633 ;
  assign n7639 = ~n7637 & n7638 ;
  assign n7640 = ~n7632 & ~n7639 ;
  assign n7641 = \data_i[123]_pad  & ~n5029 ;
  assign n7642 = \mix1_data_o_reg_reg[123]/NET0131  & n5029 ;
  assign n7643 = ~n7641 & ~n7642 ;
  assign n7644 = ~n1159 & ~n7643 ;
  assign n7645 = \sub1_data_reg_reg[123]/NET0131  & n1159 ;
  assign n7646 = ~n7644 & ~n7645 ;
  assign n7647 = ~n5028 & n7646 ;
  assign n7648 = ~\sub1_data_reg_reg[123]/NET0131  & n5028 ;
  assign n7649 = ~n7647 & ~n7648 ;
  assign n7650 = ~n5027 & ~n7649 ;
  assign n7651 = ~\mix1_data_o_reg_reg[123]/NET0131  & n5027 ;
  assign n7652 = ~n7650 & ~n7651 ;
  assign n7653 = n5026 & ~n7652 ;
  assign n7654 = ~\sub1_data_reg_reg[123]/NET0131  & ~n5026 ;
  assign n7655 = ~n7653 & ~n7654 ;
  assign n7656 = \state_reg/NET0131  & ~n7655 ;
  assign n7657 = ~\state_reg/NET0131  & n7646 ;
  assign n7658 = ~n7656 & ~n7657 ;
  assign n7660 = \key_i[123]_pad  & n7658 ;
  assign n7659 = ~\key_i[123]_pad  & ~n7658 ;
  assign n7661 = n933 & ~n7659 ;
  assign n7662 = ~n7660 & n7661 ;
  assign n7664 = ~\ks1_key_reg_reg[123]/NET0131  & ~n7658 ;
  assign n7665 = \ks1_key_reg_reg[123]/NET0131  & n7658 ;
  assign n7666 = ~n7664 & ~n7665 ;
  assign n7667 = n5053 & ~n7666 ;
  assign n7663 = ~\data_o[123]_pad  & ~n5053 ;
  assign n7668 = ~n933 & ~n7663 ;
  assign n7669 = ~n7667 & n7668 ;
  assign n7670 = ~n7662 & ~n7669 ;
  assign n7671 = \data_i[41]_pad  & ~n5029 ;
  assign n7672 = \mix1_data_o_reg_reg[41]/NET0131  & n5029 ;
  assign n7673 = ~n7671 & ~n7672 ;
  assign n7674 = ~n1159 & ~n7673 ;
  assign n7675 = \sub1_data_reg_reg[41]/NET0131  & n1159 ;
  assign n7676 = ~n7674 & ~n7675 ;
  assign n7677 = ~n5028 & n7676 ;
  assign n7678 = ~\sub1_data_reg_reg[41]/NET0131  & n5028 ;
  assign n7679 = ~n7677 & ~n7678 ;
  assign n7680 = ~n5027 & ~n7679 ;
  assign n7681 = ~\mix1_data_o_reg_reg[41]/NET0131  & n5027 ;
  assign n7682 = ~n7680 & ~n7681 ;
  assign n7683 = n5026 & ~n7682 ;
  assign n7684 = ~\sub1_data_reg_reg[41]/NET0131  & ~n5026 ;
  assign n7685 = ~n7683 & ~n7684 ;
  assign n7686 = \state_reg/NET0131  & ~n7685 ;
  assign n7687 = ~\state_reg/NET0131  & n7676 ;
  assign n7688 = ~n7686 & ~n7687 ;
  assign n7690 = \key_i[41]_pad  & n7688 ;
  assign n7689 = ~\key_i[41]_pad  & ~n7688 ;
  assign n7691 = n933 & ~n7689 ;
  assign n7692 = ~n7690 & n7691 ;
  assign n7694 = ~\ks1_key_reg_reg[41]/P0002  & ~n7688 ;
  assign n7695 = \ks1_key_reg_reg[41]/P0002  & n7688 ;
  assign n7696 = ~n7694 & ~n7695 ;
  assign n7697 = n5053 & ~n7696 ;
  assign n7693 = ~\data_o[41]_pad  & ~n5053 ;
  assign n7698 = ~n933 & ~n7693 ;
  assign n7699 = ~n7697 & n7698 ;
  assign n7700 = ~n7692 & ~n7699 ;
  assign n7701 = \data_i[47]_pad  & ~n5029 ;
  assign n7702 = \mix1_data_o_reg_reg[47]/NET0131  & n5029 ;
  assign n7703 = ~n7701 & ~n7702 ;
  assign n7704 = ~n1159 & ~n7703 ;
  assign n7705 = \sub1_data_reg_reg[47]/NET0131  & n1159 ;
  assign n7706 = ~n7704 & ~n7705 ;
  assign n7707 = ~n5028 & n7706 ;
  assign n7708 = ~\sub1_data_reg_reg[47]/NET0131  & n5028 ;
  assign n7709 = ~n7707 & ~n7708 ;
  assign n7710 = ~n5027 & ~n7709 ;
  assign n7711 = ~\mix1_data_o_reg_reg[47]/NET0131  & n5027 ;
  assign n7712 = ~n7710 & ~n7711 ;
  assign n7713 = n5026 & ~n7712 ;
  assign n7714 = ~\sub1_data_reg_reg[47]/NET0131  & ~n5026 ;
  assign n7715 = ~n7713 & ~n7714 ;
  assign n7716 = \state_reg/NET0131  & ~n7715 ;
  assign n7717 = ~\state_reg/NET0131  & n7706 ;
  assign n7718 = ~n7716 & ~n7717 ;
  assign n7720 = \key_i[47]_pad  & n7718 ;
  assign n7719 = ~\key_i[47]_pad  & ~n7718 ;
  assign n7721 = n933 & ~n7719 ;
  assign n7722 = ~n7720 & n7721 ;
  assign n7724 = ~\ks1_key_reg_reg[47]/P0002  & ~n7718 ;
  assign n7725 = \ks1_key_reg_reg[47]/P0002  & n7718 ;
  assign n7726 = ~n7724 & ~n7725 ;
  assign n7727 = n5053 & ~n7726 ;
  assign n7723 = ~\data_o[47]_pad  & ~n5053 ;
  assign n7728 = ~n933 & ~n7723 ;
  assign n7729 = ~n7727 & n7728 ;
  assign n7730 = ~n7722 & ~n7729 ;
  assign n7731 = \data_i[42]_pad  & ~n5029 ;
  assign n7732 = \mix1_data_o_reg_reg[42]/NET0131  & n5029 ;
  assign n7733 = ~n7731 & ~n7732 ;
  assign n7734 = ~n1159 & ~n7733 ;
  assign n7735 = \sub1_data_reg_reg[42]/NET0131  & n1159 ;
  assign n7736 = ~n7734 & ~n7735 ;
  assign n7737 = ~n5028 & n7736 ;
  assign n7738 = ~\sub1_data_reg_reg[42]/NET0131  & n5028 ;
  assign n7739 = ~n7737 & ~n7738 ;
  assign n7740 = ~n5027 & ~n7739 ;
  assign n7741 = ~\mix1_data_o_reg_reg[42]/NET0131  & n5027 ;
  assign n7742 = ~n7740 & ~n7741 ;
  assign n7743 = n5026 & ~n7742 ;
  assign n7744 = ~\sub1_data_reg_reg[42]/NET0131  & ~n5026 ;
  assign n7745 = ~n7743 & ~n7744 ;
  assign n7746 = \state_reg/NET0131  & ~n7745 ;
  assign n7747 = ~\state_reg/NET0131  & n7736 ;
  assign n7748 = ~n7746 & ~n7747 ;
  assign n7750 = \key_i[42]_pad  & n7748 ;
  assign n7749 = ~\key_i[42]_pad  & ~n7748 ;
  assign n7751 = n933 & ~n7749 ;
  assign n7752 = ~n7750 & n7751 ;
  assign n7754 = ~\ks1_key_reg_reg[42]/P0002  & ~n7748 ;
  assign n7755 = \ks1_key_reg_reg[42]/P0002  & n7748 ;
  assign n7756 = ~n7754 & ~n7755 ;
  assign n7757 = n5053 & ~n7756 ;
  assign n7753 = ~\data_o[42]_pad  & ~n5053 ;
  assign n7758 = ~n933 & ~n7753 ;
  assign n7759 = ~n7757 & n7758 ;
  assign n7760 = ~n7752 & ~n7759 ;
  assign n7761 = \data_i[124]_pad  & ~n5029 ;
  assign n7762 = \mix1_data_o_reg_reg[124]/NET0131  & n5029 ;
  assign n7763 = ~n7761 & ~n7762 ;
  assign n7764 = ~n1159 & ~n7763 ;
  assign n7765 = \sub1_data_reg_reg[124]/NET0131  & n1159 ;
  assign n7766 = ~n7764 & ~n7765 ;
  assign n7767 = ~n5028 & n7766 ;
  assign n7768 = ~\sub1_data_reg_reg[124]/NET0131  & n5028 ;
  assign n7769 = ~n7767 & ~n7768 ;
  assign n7770 = ~n5027 & ~n7769 ;
  assign n7771 = ~\mix1_data_o_reg_reg[124]/NET0131  & n5027 ;
  assign n7772 = ~n7770 & ~n7771 ;
  assign n7773 = n5026 & ~n7772 ;
  assign n7774 = ~\sub1_data_reg_reg[124]/NET0131  & ~n5026 ;
  assign n7775 = ~n7773 & ~n7774 ;
  assign n7776 = \state_reg/NET0131  & ~n7775 ;
  assign n7777 = ~\state_reg/NET0131  & n7766 ;
  assign n7778 = ~n7776 & ~n7777 ;
  assign n7780 = \key_i[124]_pad  & n7778 ;
  assign n7779 = ~\key_i[124]_pad  & ~n7778 ;
  assign n7781 = n933 & ~n7779 ;
  assign n7782 = ~n7780 & n7781 ;
  assign n7784 = ~\ks1_key_reg_reg[124]/NET0131  & ~n7778 ;
  assign n7785 = \ks1_key_reg_reg[124]/NET0131  & n7778 ;
  assign n7786 = ~n7784 & ~n7785 ;
  assign n7787 = n5053 & ~n7786 ;
  assign n7783 = ~\data_o[124]_pad  & ~n5053 ;
  assign n7788 = ~n933 & ~n7783 ;
  assign n7789 = ~n7787 & n7788 ;
  assign n7790 = ~n7782 & ~n7789 ;
  assign n7791 = \data_i[43]_pad  & ~n5029 ;
  assign n7792 = \mix1_data_o_reg_reg[43]/NET0131  & n5029 ;
  assign n7793 = ~n7791 & ~n7792 ;
  assign n7794 = ~n1159 & ~n7793 ;
  assign n7795 = \sub1_data_reg_reg[43]/NET0131  & n1159 ;
  assign n7796 = ~n7794 & ~n7795 ;
  assign n7797 = ~n5028 & n7796 ;
  assign n7798 = ~\sub1_data_reg_reg[43]/NET0131  & n5028 ;
  assign n7799 = ~n7797 & ~n7798 ;
  assign n7800 = ~n5027 & ~n7799 ;
  assign n7801 = ~\mix1_data_o_reg_reg[43]/NET0131  & n5027 ;
  assign n7802 = ~n7800 & ~n7801 ;
  assign n7803 = n5026 & ~n7802 ;
  assign n7804 = ~\sub1_data_reg_reg[43]/NET0131  & ~n5026 ;
  assign n7805 = ~n7803 & ~n7804 ;
  assign n7806 = \state_reg/NET0131  & ~n7805 ;
  assign n7807 = ~\state_reg/NET0131  & n7796 ;
  assign n7808 = ~n7806 & ~n7807 ;
  assign n7810 = \key_i[43]_pad  & n7808 ;
  assign n7809 = ~\key_i[43]_pad  & ~n7808 ;
  assign n7811 = n933 & ~n7809 ;
  assign n7812 = ~n7810 & n7811 ;
  assign n7814 = ~\ks1_key_reg_reg[43]/P0002  & ~n7808 ;
  assign n7815 = \ks1_key_reg_reg[43]/P0002  & n7808 ;
  assign n7816 = ~n7814 & ~n7815 ;
  assign n7817 = n5053 & ~n7816 ;
  assign n7813 = ~\data_o[43]_pad  & ~n5053 ;
  assign n7818 = ~n933 & ~n7813 ;
  assign n7819 = ~n7817 & n7818 ;
  assign n7820 = ~n7812 & ~n7819 ;
  assign n7821 = \data_i[107]_pad  & ~n5029 ;
  assign n7822 = \mix1_data_o_reg_reg[107]/NET0131  & n5029 ;
  assign n7823 = ~n7821 & ~n7822 ;
  assign n7824 = ~n1159 & ~n7823 ;
  assign n7825 = \sub1_data_reg_reg[107]/NET0131  & n1159 ;
  assign n7826 = ~n7824 & ~n7825 ;
  assign n7827 = ~n5028 & n7826 ;
  assign n7828 = ~\sub1_data_reg_reg[107]/NET0131  & n5028 ;
  assign n7829 = ~n7827 & ~n7828 ;
  assign n7830 = ~n5027 & ~n7829 ;
  assign n7831 = ~\mix1_data_o_reg_reg[107]/NET0131  & n5027 ;
  assign n7832 = ~n7830 & ~n7831 ;
  assign n7833 = n5026 & ~n7832 ;
  assign n7834 = ~\sub1_data_reg_reg[107]/NET0131  & ~n5026 ;
  assign n7835 = ~n7833 & ~n7834 ;
  assign n7836 = \state_reg/NET0131  & ~n7835 ;
  assign n7837 = ~\state_reg/NET0131  & n7826 ;
  assign n7838 = ~n7836 & ~n7837 ;
  assign n7840 = \key_i[107]_pad  & n7838 ;
  assign n7839 = ~\key_i[107]_pad  & ~n7838 ;
  assign n7841 = n933 & ~n7839 ;
  assign n7842 = ~n7840 & n7841 ;
  assign n7844 = ~\ks1_key_reg_reg[107]/NET0131  & ~n7838 ;
  assign n7845 = \ks1_key_reg_reg[107]/NET0131  & n7838 ;
  assign n7846 = ~n7844 & ~n7845 ;
  assign n7847 = n5053 & ~n7846 ;
  assign n7843 = ~\data_o[107]_pad  & ~n5053 ;
  assign n7848 = ~n933 & ~n7843 ;
  assign n7849 = ~n7847 & n7848 ;
  assign n7850 = ~n7842 & ~n7849 ;
  assign n7851 = \data_i[125]_pad  & ~n5029 ;
  assign n7852 = \mix1_data_o_reg_reg[125]/NET0131  & n5029 ;
  assign n7853 = ~n7851 & ~n7852 ;
  assign n7854 = ~n1159 & ~n7853 ;
  assign n7855 = \sub1_data_reg_reg[125]/NET0131  & n1159 ;
  assign n7856 = ~n7854 & ~n7855 ;
  assign n7857 = ~n5028 & n7856 ;
  assign n7858 = ~\sub1_data_reg_reg[125]/NET0131  & n5028 ;
  assign n7859 = ~n7857 & ~n7858 ;
  assign n7860 = ~n5027 & ~n7859 ;
  assign n7861 = ~\mix1_data_o_reg_reg[125]/NET0131  & n5027 ;
  assign n7862 = ~n7860 & ~n7861 ;
  assign n7863 = n5026 & ~n7862 ;
  assign n7864 = ~\sub1_data_reg_reg[125]/NET0131  & ~n5026 ;
  assign n7865 = ~n7863 & ~n7864 ;
  assign n7866 = \state_reg/NET0131  & ~n7865 ;
  assign n7867 = ~\state_reg/NET0131  & n7856 ;
  assign n7868 = ~n7866 & ~n7867 ;
  assign n7870 = \key_i[125]_pad  & n7868 ;
  assign n7869 = ~\key_i[125]_pad  & ~n7868 ;
  assign n7871 = n933 & ~n7869 ;
  assign n7872 = ~n7870 & n7871 ;
  assign n7874 = ~\ks1_key_reg_reg[125]/NET0131  & ~n7868 ;
  assign n7875 = \ks1_key_reg_reg[125]/NET0131  & n7868 ;
  assign n7876 = ~n7874 & ~n7875 ;
  assign n7877 = n5053 & ~n7876 ;
  assign n7873 = ~\data_o[125]_pad  & ~n5053 ;
  assign n7878 = ~n933 & ~n7873 ;
  assign n7879 = ~n7877 & n7878 ;
  assign n7880 = ~n7872 & ~n7879 ;
  assign n7881 = \data_i[44]_pad  & ~n5029 ;
  assign n7882 = \mix1_data_o_reg_reg[44]/NET0131  & n5029 ;
  assign n7883 = ~n7881 & ~n7882 ;
  assign n7884 = ~n1159 & ~n7883 ;
  assign n7885 = \sub1_data_reg_reg[44]/NET0131  & n1159 ;
  assign n7886 = ~n7884 & ~n7885 ;
  assign n7887 = ~n5028 & n7886 ;
  assign n7888 = ~\sub1_data_reg_reg[44]/NET0131  & n5028 ;
  assign n7889 = ~n7887 & ~n7888 ;
  assign n7890 = ~n5027 & ~n7889 ;
  assign n7891 = ~\mix1_data_o_reg_reg[44]/NET0131  & n5027 ;
  assign n7892 = ~n7890 & ~n7891 ;
  assign n7893 = n5026 & ~n7892 ;
  assign n7894 = ~\sub1_data_reg_reg[44]/NET0131  & ~n5026 ;
  assign n7895 = ~n7893 & ~n7894 ;
  assign n7896 = \state_reg/NET0131  & ~n7895 ;
  assign n7897 = ~\state_reg/NET0131  & n7886 ;
  assign n7898 = ~n7896 & ~n7897 ;
  assign n7900 = \key_i[44]_pad  & n7898 ;
  assign n7899 = ~\key_i[44]_pad  & ~n7898 ;
  assign n7901 = n933 & ~n7899 ;
  assign n7902 = ~n7900 & n7901 ;
  assign n7904 = ~\ks1_key_reg_reg[44]/P0002  & ~n7898 ;
  assign n7905 = \ks1_key_reg_reg[44]/P0002  & n7898 ;
  assign n7906 = ~n7904 & ~n7905 ;
  assign n7907 = n5053 & ~n7906 ;
  assign n7903 = ~\data_o[44]_pad  & ~n5053 ;
  assign n7908 = ~n933 & ~n7903 ;
  assign n7909 = ~n7907 & n7908 ;
  assign n7910 = ~n7902 & ~n7909 ;
  assign n7911 = \data_i[108]_pad  & ~n5029 ;
  assign n7912 = \mix1_data_o_reg_reg[108]/NET0131  & n5029 ;
  assign n7913 = ~n7911 & ~n7912 ;
  assign n7914 = ~n1159 & ~n7913 ;
  assign n7915 = \sub1_data_reg_reg[108]/NET0131  & n1159 ;
  assign n7916 = ~n7914 & ~n7915 ;
  assign n7917 = ~n5028 & n7916 ;
  assign n7918 = ~\sub1_data_reg_reg[108]/NET0131  & n5028 ;
  assign n7919 = ~n7917 & ~n7918 ;
  assign n7920 = ~n5027 & ~n7919 ;
  assign n7921 = ~\mix1_data_o_reg_reg[108]/NET0131  & n5027 ;
  assign n7922 = ~n7920 & ~n7921 ;
  assign n7923 = n5026 & ~n7922 ;
  assign n7924 = ~\sub1_data_reg_reg[108]/NET0131  & ~n5026 ;
  assign n7925 = ~n7923 & ~n7924 ;
  assign n7926 = \state_reg/NET0131  & ~n7925 ;
  assign n7927 = ~\state_reg/NET0131  & n7916 ;
  assign n7928 = ~n7926 & ~n7927 ;
  assign n7930 = \key_i[108]_pad  & n7928 ;
  assign n7929 = ~\key_i[108]_pad  & ~n7928 ;
  assign n7931 = n933 & ~n7929 ;
  assign n7932 = ~n7930 & n7931 ;
  assign n7934 = ~\ks1_key_reg_reg[108]/NET0131  & ~n7928 ;
  assign n7935 = \ks1_key_reg_reg[108]/NET0131  & n7928 ;
  assign n7936 = ~n7934 & ~n7935 ;
  assign n7937 = n5053 & ~n7936 ;
  assign n7933 = ~\data_o[108]_pad  & ~n5053 ;
  assign n7938 = ~n933 & ~n7933 ;
  assign n7939 = ~n7937 & n7938 ;
  assign n7940 = ~n7932 & ~n7939 ;
  assign n7941 = \data_i[45]_pad  & ~n5029 ;
  assign n7942 = \mix1_data_o_reg_reg[45]/NET0131  & n5029 ;
  assign n7943 = ~n7941 & ~n7942 ;
  assign n7944 = ~n1159 & ~n7943 ;
  assign n7945 = \sub1_data_reg_reg[45]/NET0131  & n1159 ;
  assign n7946 = ~n7944 & ~n7945 ;
  assign n7947 = ~n5028 & n7946 ;
  assign n7948 = ~\sub1_data_reg_reg[45]/NET0131  & n5028 ;
  assign n7949 = ~n7947 & ~n7948 ;
  assign n7950 = ~n5027 & ~n7949 ;
  assign n7951 = ~\mix1_data_o_reg_reg[45]/NET0131  & n5027 ;
  assign n7952 = ~n7950 & ~n7951 ;
  assign n7953 = n5026 & ~n7952 ;
  assign n7954 = ~\sub1_data_reg_reg[45]/NET0131  & ~n5026 ;
  assign n7955 = ~n7953 & ~n7954 ;
  assign n7956 = \state_reg/NET0131  & ~n7955 ;
  assign n7957 = ~\state_reg/NET0131  & n7946 ;
  assign n7958 = ~n7956 & ~n7957 ;
  assign n7960 = \key_i[45]_pad  & n7958 ;
  assign n7959 = ~\key_i[45]_pad  & ~n7958 ;
  assign n7961 = n933 & ~n7959 ;
  assign n7962 = ~n7960 & n7961 ;
  assign n7964 = ~\ks1_key_reg_reg[45]/P0002  & ~n7958 ;
  assign n7965 = \ks1_key_reg_reg[45]/P0002  & n7958 ;
  assign n7966 = ~n7964 & ~n7965 ;
  assign n7967 = n5053 & ~n7966 ;
  assign n7963 = ~\data_o[45]_pad  & ~n5053 ;
  assign n7968 = ~n933 & ~n7963 ;
  assign n7969 = ~n7967 & n7968 ;
  assign n7970 = ~n7962 & ~n7969 ;
  assign n7971 = \data_i[46]_pad  & ~n5029 ;
  assign n7972 = \mix1_data_o_reg_reg[46]/NET0131  & n5029 ;
  assign n7973 = ~n7971 & ~n7972 ;
  assign n7974 = ~n1159 & ~n7973 ;
  assign n7975 = \sub1_data_reg_reg[46]/NET0131  & n1159 ;
  assign n7976 = ~n7974 & ~n7975 ;
  assign n7977 = ~n5028 & n7976 ;
  assign n7978 = ~\sub1_data_reg_reg[46]/NET0131  & n5028 ;
  assign n7979 = ~n7977 & ~n7978 ;
  assign n7980 = ~n5027 & ~n7979 ;
  assign n7981 = ~\mix1_data_o_reg_reg[46]/NET0131  & n5027 ;
  assign n7982 = ~n7980 & ~n7981 ;
  assign n7983 = n5026 & ~n7982 ;
  assign n7984 = ~\sub1_data_reg_reg[46]/NET0131  & ~n5026 ;
  assign n7985 = ~n7983 & ~n7984 ;
  assign n7986 = \state_reg/NET0131  & ~n7985 ;
  assign n7987 = ~\state_reg/NET0131  & n7976 ;
  assign n7988 = ~n7986 & ~n7987 ;
  assign n7990 = \key_i[46]_pad  & n7988 ;
  assign n7989 = ~\key_i[46]_pad  & ~n7988 ;
  assign n7991 = n933 & ~n7989 ;
  assign n7992 = ~n7990 & n7991 ;
  assign n7994 = ~\ks1_key_reg_reg[46]/P0002  & ~n7988 ;
  assign n7995 = \ks1_key_reg_reg[46]/P0002  & n7988 ;
  assign n7996 = ~n7994 & ~n7995 ;
  assign n7997 = n5053 & ~n7996 ;
  assign n7993 = ~\data_o[46]_pad  & ~n5053 ;
  assign n7998 = ~n933 & ~n7993 ;
  assign n7999 = ~n7997 & n7998 ;
  assign n8000 = ~n7992 & ~n7999 ;
  assign n8001 = \data_i[126]_pad  & ~n5029 ;
  assign n8002 = \mix1_data_o_reg_reg[126]/NET0131  & n5029 ;
  assign n8003 = ~n8001 & ~n8002 ;
  assign n8004 = ~n1159 & ~n8003 ;
  assign n8005 = \sub1_data_reg_reg[126]/NET0131  & n1159 ;
  assign n8006 = ~n8004 & ~n8005 ;
  assign n8007 = ~n5028 & n8006 ;
  assign n8008 = ~\sub1_data_reg_reg[126]/NET0131  & n5028 ;
  assign n8009 = ~n8007 & ~n8008 ;
  assign n8010 = ~n5027 & ~n8009 ;
  assign n8011 = ~\mix1_data_o_reg_reg[126]/NET0131  & n5027 ;
  assign n8012 = ~n8010 & ~n8011 ;
  assign n8013 = n5026 & ~n8012 ;
  assign n8014 = ~\sub1_data_reg_reg[126]/NET0131  & ~n5026 ;
  assign n8015 = ~n8013 & ~n8014 ;
  assign n8016 = \state_reg/NET0131  & ~n8015 ;
  assign n8017 = ~\state_reg/NET0131  & n8006 ;
  assign n8018 = ~n8016 & ~n8017 ;
  assign n8020 = \key_i[126]_pad  & n8018 ;
  assign n8019 = ~\key_i[126]_pad  & ~n8018 ;
  assign n8021 = n933 & ~n8019 ;
  assign n8022 = ~n8020 & n8021 ;
  assign n8024 = ~\ks1_key_reg_reg[126]/NET0131  & ~n8018 ;
  assign n8025 = \ks1_key_reg_reg[126]/NET0131  & n8018 ;
  assign n8026 = ~n8024 & ~n8025 ;
  assign n8027 = n5053 & ~n8026 ;
  assign n8023 = ~\data_o[126]_pad  & ~n5053 ;
  assign n8028 = ~n933 & ~n8023 ;
  assign n8029 = ~n8027 & n8028 ;
  assign n8030 = ~n8022 & ~n8029 ;
  assign n8031 = ~\data_i[48]_pad  & ~n5029 ;
  assign n8032 = ~\mix1_data_o_reg_reg[48]/NET0131  & n5029 ;
  assign n8033 = ~n8031 & ~n8032 ;
  assign n8034 = ~n1159 & ~n8033 ;
  assign n8035 = ~\sub1_data_reg_reg[48]/NET0131  & n1159 ;
  assign n8036 = ~n8034 & ~n8035 ;
  assign n8037 = ~n5028 & ~n8036 ;
  assign n8038 = ~\sub1_data_reg_reg[48]/NET0131  & n5028 ;
  assign n8039 = ~n8037 & ~n8038 ;
  assign n8040 = ~n5027 & ~n8039 ;
  assign n8041 = ~\mix1_data_o_reg_reg[48]/NET0131  & n5027 ;
  assign n8042 = ~n8040 & ~n8041 ;
  assign n8043 = n5026 & ~n8042 ;
  assign n8044 = ~\sub1_data_reg_reg[48]/NET0131  & ~n5026 ;
  assign n8045 = ~n8043 & ~n8044 ;
  assign n8046 = \state_reg/NET0131  & ~n8045 ;
  assign n8047 = ~\state_reg/NET0131  & ~n8036 ;
  assign n8048 = ~n8046 & ~n8047 ;
  assign n8050 = \key_i[48]_pad  & n8048 ;
  assign n8049 = ~\key_i[48]_pad  & ~n8048 ;
  assign n8051 = n933 & ~n8049 ;
  assign n8052 = ~n8050 & n8051 ;
  assign n8054 = ~\ks1_key_reg_reg[48]/NET0131  & ~n8048 ;
  assign n8055 = \ks1_key_reg_reg[48]/NET0131  & n8048 ;
  assign n8056 = ~n8054 & ~n8055 ;
  assign n8057 = n5053 & ~n8056 ;
  assign n8053 = ~\data_o[48]_pad  & ~n5053 ;
  assign n8058 = ~n933 & ~n8053 ;
  assign n8059 = ~n8057 & n8058 ;
  assign n8060 = ~n8052 & ~n8059 ;
  assign n8061 = \data_i[127]_pad  & ~n5029 ;
  assign n8062 = \mix1_data_o_reg_reg[127]/NET0131  & n5029 ;
  assign n8063 = ~n8061 & ~n8062 ;
  assign n8064 = ~n1159 & ~n8063 ;
  assign n8065 = \sub1_data_reg_reg[127]/NET0131  & n1159 ;
  assign n8066 = ~n8064 & ~n8065 ;
  assign n8067 = ~n5028 & n8066 ;
  assign n8068 = ~\sub1_data_reg_reg[127]/NET0131  & n5028 ;
  assign n8069 = ~n8067 & ~n8068 ;
  assign n8070 = ~n5027 & ~n8069 ;
  assign n8071 = ~\mix1_data_o_reg_reg[127]/NET0131  & n5027 ;
  assign n8072 = ~n8070 & ~n8071 ;
  assign n8073 = n5026 & ~n8072 ;
  assign n8074 = ~\sub1_data_reg_reg[127]/NET0131  & ~n5026 ;
  assign n8075 = ~n8073 & ~n8074 ;
  assign n8076 = \state_reg/NET0131  & ~n8075 ;
  assign n8077 = ~\state_reg/NET0131  & n8066 ;
  assign n8078 = ~n8076 & ~n8077 ;
  assign n8080 = \key_i[127]_pad  & n8078 ;
  assign n8079 = ~\key_i[127]_pad  & ~n8078 ;
  assign n8081 = n933 & ~n8079 ;
  assign n8082 = ~n8080 & n8081 ;
  assign n8084 = ~\ks1_key_reg_reg[127]/NET0131  & ~n8078 ;
  assign n8085 = \ks1_key_reg_reg[127]/NET0131  & n8078 ;
  assign n8086 = ~n8084 & ~n8085 ;
  assign n8087 = n5053 & ~n8086 ;
  assign n8083 = ~\data_o[127]_pad  & ~n5053 ;
  assign n8088 = ~n933 & ~n8083 ;
  assign n8089 = ~n8087 & n8088 ;
  assign n8090 = ~n8082 & ~n8089 ;
  assign n8091 = ~\data_i[49]_pad  & ~n5029 ;
  assign n8092 = ~\mix1_data_o_reg_reg[49]/NET0131  & n5029 ;
  assign n8093 = ~n8091 & ~n8092 ;
  assign n8094 = ~n1159 & ~n8093 ;
  assign n8095 = ~\sub1_data_reg_reg[49]/NET0131  & n1159 ;
  assign n8096 = ~n8094 & ~n8095 ;
  assign n8097 = ~n5028 & ~n8096 ;
  assign n8098 = ~\sub1_data_reg_reg[49]/NET0131  & n5028 ;
  assign n8099 = ~n8097 & ~n8098 ;
  assign n8100 = ~n5027 & ~n8099 ;
  assign n8101 = ~\mix1_data_o_reg_reg[49]/NET0131  & n5027 ;
  assign n8102 = ~n8100 & ~n8101 ;
  assign n8103 = n5026 & ~n8102 ;
  assign n8104 = ~\sub1_data_reg_reg[49]/NET0131  & ~n5026 ;
  assign n8105 = ~n8103 & ~n8104 ;
  assign n8106 = \state_reg/NET0131  & ~n8105 ;
  assign n8107 = ~\state_reg/NET0131  & ~n8096 ;
  assign n8108 = ~n8106 & ~n8107 ;
  assign n8110 = \key_i[49]_pad  & n8108 ;
  assign n8109 = ~\key_i[49]_pad  & ~n8108 ;
  assign n8111 = n933 & ~n8109 ;
  assign n8112 = ~n8110 & n8111 ;
  assign n8114 = ~\ks1_key_reg_reg[49]/NET0131  & ~n8108 ;
  assign n8115 = \ks1_key_reg_reg[49]/NET0131  & n8108 ;
  assign n8116 = ~n8114 & ~n8115 ;
  assign n8117 = n5053 & ~n8116 ;
  assign n8113 = ~\data_o[49]_pad  & ~n5053 ;
  assign n8118 = ~n933 & ~n8113 ;
  assign n8119 = ~n8117 & n8118 ;
  assign n8120 = ~n8112 & ~n8119 ;
  assign n8121 = \data_i[109]_pad  & ~n5029 ;
  assign n8122 = \mix1_data_o_reg_reg[109]/NET0131  & n5029 ;
  assign n8123 = ~n8121 & ~n8122 ;
  assign n8124 = ~n1159 & ~n8123 ;
  assign n8125 = \sub1_data_reg_reg[109]/NET0131  & n1159 ;
  assign n8126 = ~n8124 & ~n8125 ;
  assign n8127 = ~n5028 & n8126 ;
  assign n8128 = ~\sub1_data_reg_reg[109]/NET0131  & n5028 ;
  assign n8129 = ~n8127 & ~n8128 ;
  assign n8130 = ~n5027 & ~n8129 ;
  assign n8131 = ~\mix1_data_o_reg_reg[109]/NET0131  & n5027 ;
  assign n8132 = ~n8130 & ~n8131 ;
  assign n8133 = n5026 & ~n8132 ;
  assign n8134 = ~\sub1_data_reg_reg[109]/NET0131  & ~n5026 ;
  assign n8135 = ~n8133 & ~n8134 ;
  assign n8136 = \state_reg/NET0131  & ~n8135 ;
  assign n8137 = ~\state_reg/NET0131  & n8126 ;
  assign n8138 = ~n8136 & ~n8137 ;
  assign n8140 = \key_i[109]_pad  & n8138 ;
  assign n8139 = ~\key_i[109]_pad  & ~n8138 ;
  assign n8141 = n933 & ~n8139 ;
  assign n8142 = ~n8140 & n8141 ;
  assign n8144 = ~\ks1_key_reg_reg[109]/P0002  & ~n8138 ;
  assign n8145 = \ks1_key_reg_reg[109]/P0002  & n8138 ;
  assign n8146 = ~n8144 & ~n8145 ;
  assign n8147 = n5053 & ~n8146 ;
  assign n8143 = ~\data_o[109]_pad  & ~n5053 ;
  assign n8148 = ~n933 & ~n8143 ;
  assign n8149 = ~n8147 & n8148 ;
  assign n8150 = ~n8142 & ~n8149 ;
  assign n8151 = \data_i[4]_pad  & ~n5029 ;
  assign n8152 = \mix1_data_o_reg_reg[4]/NET0131  & n5029 ;
  assign n8153 = ~n8151 & ~n8152 ;
  assign n8154 = ~n1159 & ~n8153 ;
  assign n8155 = \sub1_data_reg_reg[4]/NET0131  & n1159 ;
  assign n8156 = ~n8154 & ~n8155 ;
  assign n8157 = ~n5028 & n8156 ;
  assign n8158 = ~\sub1_data_reg_reg[4]/NET0131  & n5028 ;
  assign n8159 = ~n8157 & ~n8158 ;
  assign n8160 = ~n5027 & ~n8159 ;
  assign n8161 = ~\mix1_data_o_reg_reg[4]/NET0131  & n5027 ;
  assign n8162 = ~n8160 & ~n8161 ;
  assign n8163 = n5026 & ~n8162 ;
  assign n8164 = ~\sub1_data_reg_reg[4]/NET0131  & ~n5026 ;
  assign n8165 = ~n8163 & ~n8164 ;
  assign n8166 = \state_reg/NET0131  & ~n8165 ;
  assign n8167 = ~\state_reg/NET0131  & n8156 ;
  assign n8168 = ~n8166 & ~n8167 ;
  assign n8170 = \key_i[4]_pad  & n8168 ;
  assign n8169 = ~\key_i[4]_pad  & ~n8168 ;
  assign n8171 = n933 & ~n8169 ;
  assign n8172 = ~n8170 & n8171 ;
  assign n8174 = ~\ks1_key_reg_reg[4]/NET0131  & ~n8168 ;
  assign n8175 = \ks1_key_reg_reg[4]/NET0131  & n8168 ;
  assign n8176 = ~n8174 & ~n8175 ;
  assign n8177 = n5053 & ~n8176 ;
  assign n8173 = ~\data_o[4]_pad  & ~n5053 ;
  assign n8178 = ~n933 & ~n8173 ;
  assign n8179 = ~n8177 & n8178 ;
  assign n8180 = ~n8172 & ~n8179 ;
  assign n8181 = \data_i[12]_pad  & ~n5029 ;
  assign n8182 = \mix1_data_o_reg_reg[12]/NET0131  & n5029 ;
  assign n8183 = ~n8181 & ~n8182 ;
  assign n8184 = ~n1159 & ~n8183 ;
  assign n8185 = \sub1_data_reg_reg[12]/NET0131  & n1159 ;
  assign n8186 = ~n8184 & ~n8185 ;
  assign n8187 = ~n5028 & n8186 ;
  assign n8188 = ~\sub1_data_reg_reg[12]/NET0131  & n5028 ;
  assign n8189 = ~n8187 & ~n8188 ;
  assign n8190 = ~n5027 & ~n8189 ;
  assign n8191 = ~\mix1_data_o_reg_reg[12]/NET0131  & n5027 ;
  assign n8192 = ~n8190 & ~n8191 ;
  assign n8193 = n5026 & ~n8192 ;
  assign n8194 = ~\sub1_data_reg_reg[12]/NET0131  & ~n5026 ;
  assign n8195 = ~n8193 & ~n8194 ;
  assign n8196 = \state_reg/NET0131  & ~n8195 ;
  assign n8197 = ~\state_reg/NET0131  & n8186 ;
  assign n8198 = ~n8196 & ~n8197 ;
  assign n8200 = \key_i[12]_pad  & n8198 ;
  assign n8199 = ~\key_i[12]_pad  & ~n8198 ;
  assign n8201 = n933 & ~n8199 ;
  assign n8202 = ~n8200 & n8201 ;
  assign n8204 = ~\ks1_key_reg_reg[12]/NET0131  & ~n8198 ;
  assign n8205 = \ks1_key_reg_reg[12]/NET0131  & n8198 ;
  assign n8206 = ~n8204 & ~n8205 ;
  assign n8207 = n5053 & ~n8206 ;
  assign n8203 = ~\data_o[12]_pad  & ~n5053 ;
  assign n8208 = ~n933 & ~n8203 ;
  assign n8209 = ~n8207 & n8208 ;
  assign n8210 = ~n8202 & ~n8209 ;
  assign n8211 = ~\data_i[50]_pad  & ~n5029 ;
  assign n8212 = ~\mix1_data_o_reg_reg[50]/NET0131  & n5029 ;
  assign n8213 = ~n8211 & ~n8212 ;
  assign n8214 = ~n1159 & ~n8213 ;
  assign n8215 = ~\sub1_data_reg_reg[50]/NET0131  & n1159 ;
  assign n8216 = ~n8214 & ~n8215 ;
  assign n8217 = ~n5028 & ~n8216 ;
  assign n8218 = ~\sub1_data_reg_reg[50]/NET0131  & n5028 ;
  assign n8219 = ~n8217 & ~n8218 ;
  assign n8220 = ~n5027 & ~n8219 ;
  assign n8221 = ~\mix1_data_o_reg_reg[50]/NET0131  & n5027 ;
  assign n8222 = ~n8220 & ~n8221 ;
  assign n8223 = n5026 & ~n8222 ;
  assign n8224 = ~\sub1_data_reg_reg[50]/NET0131  & ~n5026 ;
  assign n8225 = ~n8223 & ~n8224 ;
  assign n8226 = \state_reg/NET0131  & ~n8225 ;
  assign n8227 = ~\state_reg/NET0131  & ~n8216 ;
  assign n8228 = ~n8226 & ~n8227 ;
  assign n8230 = \key_i[50]_pad  & n8228 ;
  assign n8229 = ~\key_i[50]_pad  & ~n8228 ;
  assign n8231 = n933 & ~n8229 ;
  assign n8232 = ~n8230 & n8231 ;
  assign n8234 = ~\ks1_key_reg_reg[50]/NET0131  & ~n8228 ;
  assign n8235 = \ks1_key_reg_reg[50]/NET0131  & n8228 ;
  assign n8236 = ~n8234 & ~n8235 ;
  assign n8237 = n5053 & ~n8236 ;
  assign n8233 = ~\data_o[50]_pad  & ~n5053 ;
  assign n8238 = ~n933 & ~n8233 ;
  assign n8239 = ~n8237 & n8238 ;
  assign n8240 = ~n8232 & ~n8239 ;
  assign n8241 = \data_i[10]_pad  & ~n5029 ;
  assign n8242 = \mix1_data_o_reg_reg[10]/NET0131  & n5029 ;
  assign n8243 = ~n8241 & ~n8242 ;
  assign n8244 = ~n1159 & ~n8243 ;
  assign n8245 = \sub1_data_reg_reg[10]/NET0131  & n1159 ;
  assign n8246 = ~n8244 & ~n8245 ;
  assign n8247 = ~n5028 & n8246 ;
  assign n8248 = ~\sub1_data_reg_reg[10]/NET0131  & n5028 ;
  assign n8249 = ~n8247 & ~n8248 ;
  assign n8250 = ~n5027 & ~n8249 ;
  assign n8251 = ~\mix1_data_o_reg_reg[10]/NET0131  & n5027 ;
  assign n8252 = ~n8250 & ~n8251 ;
  assign n8253 = n5026 & ~n8252 ;
  assign n8254 = ~\sub1_data_reg_reg[10]/NET0131  & ~n5026 ;
  assign n8255 = ~n8253 & ~n8254 ;
  assign n8256 = \state_reg/NET0131  & ~n8255 ;
  assign n8257 = ~\state_reg/NET0131  & n8246 ;
  assign n8258 = ~n8256 & ~n8257 ;
  assign n8260 = \key_i[10]_pad  & n8258 ;
  assign n8259 = ~\key_i[10]_pad  & ~n8258 ;
  assign n8261 = n933 & ~n8259 ;
  assign n8262 = ~n8260 & n8261 ;
  assign n8264 = ~\ks1_key_reg_reg[10]/NET0131  & ~n8258 ;
  assign n8265 = \ks1_key_reg_reg[10]/NET0131  & n8258 ;
  assign n8266 = ~n8264 & ~n8265 ;
  assign n8267 = n5053 & ~n8266 ;
  assign n8263 = ~\data_o[10]_pad  & ~n5053 ;
  assign n8268 = ~n933 & ~n8263 ;
  assign n8269 = ~n8267 & n8268 ;
  assign n8270 = ~n8262 & ~n8269 ;
  assign n8271 = \data_i[13]_pad  & ~n5029 ;
  assign n8272 = \mix1_data_o_reg_reg[13]/NET0131  & n5029 ;
  assign n8273 = ~n8271 & ~n8272 ;
  assign n8274 = ~n1159 & ~n8273 ;
  assign n8275 = \sub1_data_reg_reg[13]/NET0131  & n1159 ;
  assign n8276 = ~n8274 & ~n8275 ;
  assign n8277 = ~n5028 & n8276 ;
  assign n8278 = ~\sub1_data_reg_reg[13]/NET0131  & n5028 ;
  assign n8279 = ~n8277 & ~n8278 ;
  assign n8280 = ~n5027 & ~n8279 ;
  assign n8281 = ~\mix1_data_o_reg_reg[13]/NET0131  & n5027 ;
  assign n8282 = ~n8280 & ~n8281 ;
  assign n8283 = n5026 & ~n8282 ;
  assign n8284 = ~\sub1_data_reg_reg[13]/NET0131  & ~n5026 ;
  assign n8285 = ~n8283 & ~n8284 ;
  assign n8286 = \state_reg/NET0131  & ~n8285 ;
  assign n8287 = ~\state_reg/NET0131  & n8276 ;
  assign n8288 = ~n8286 & ~n8287 ;
  assign n8290 = \key_i[13]_pad  & n8288 ;
  assign n8289 = ~\key_i[13]_pad  & ~n8288 ;
  assign n8291 = n933 & ~n8289 ;
  assign n8292 = ~n8290 & n8291 ;
  assign n8294 = ~\ks1_key_reg_reg[13]/NET0131  & ~n8288 ;
  assign n8295 = \ks1_key_reg_reg[13]/NET0131  & n8288 ;
  assign n8296 = ~n8294 & ~n8295 ;
  assign n8297 = n5053 & ~n8296 ;
  assign n8293 = ~\data_o[13]_pad  & ~n5053 ;
  assign n8298 = ~n933 & ~n8293 ;
  assign n8299 = ~n8297 & n8298 ;
  assign n8300 = ~n8292 & ~n8299 ;
  assign n8301 = ~\data_i[51]_pad  & ~n5029 ;
  assign n8302 = ~\mix1_data_o_reg_reg[51]/NET0131  & n5029 ;
  assign n8303 = ~n8301 & ~n8302 ;
  assign n8304 = ~n1159 & ~n8303 ;
  assign n8305 = ~\sub1_data_reg_reg[51]/NET0131  & n1159 ;
  assign n8306 = ~n8304 & ~n8305 ;
  assign n8307 = ~n5028 & ~n8306 ;
  assign n8308 = ~\sub1_data_reg_reg[51]/NET0131  & n5028 ;
  assign n8309 = ~n8307 & ~n8308 ;
  assign n8310 = ~n5027 & ~n8309 ;
  assign n8311 = ~\mix1_data_o_reg_reg[51]/NET0131  & n5027 ;
  assign n8312 = ~n8310 & ~n8311 ;
  assign n8313 = n5026 & ~n8312 ;
  assign n8314 = ~\sub1_data_reg_reg[51]/NET0131  & ~n5026 ;
  assign n8315 = ~n8313 & ~n8314 ;
  assign n8316 = \state_reg/NET0131  & ~n8315 ;
  assign n8317 = ~\state_reg/NET0131  & ~n8306 ;
  assign n8318 = ~n8316 & ~n8317 ;
  assign n8320 = \key_i[51]_pad  & n8318 ;
  assign n8319 = ~\key_i[51]_pad  & ~n8318 ;
  assign n8321 = n933 & ~n8319 ;
  assign n8322 = ~n8320 & n8321 ;
  assign n8324 = ~\ks1_key_reg_reg[51]/NET0131  & ~n8318 ;
  assign n8325 = \ks1_key_reg_reg[51]/NET0131  & n8318 ;
  assign n8326 = ~n8324 & ~n8325 ;
  assign n8327 = n5053 & ~n8326 ;
  assign n8323 = ~\data_o[51]_pad  & ~n5053 ;
  assign n8328 = ~n933 & ~n8323 ;
  assign n8329 = ~n8327 & n8328 ;
  assign n8330 = ~n8322 & ~n8329 ;
  assign n8331 = ~\data_i[52]_pad  & ~n5029 ;
  assign n8332 = ~\mix1_data_o_reg_reg[52]/NET0131  & n5029 ;
  assign n8333 = ~n8331 & ~n8332 ;
  assign n8334 = ~n1159 & ~n8333 ;
  assign n8335 = ~\sub1_data_reg_reg[52]/NET0131  & n1159 ;
  assign n8336 = ~n8334 & ~n8335 ;
  assign n8337 = ~n5028 & ~n8336 ;
  assign n8338 = ~\sub1_data_reg_reg[52]/NET0131  & n5028 ;
  assign n8339 = ~n8337 & ~n8338 ;
  assign n8340 = ~n5027 & ~n8339 ;
  assign n8341 = ~\mix1_data_o_reg_reg[52]/NET0131  & n5027 ;
  assign n8342 = ~n8340 & ~n8341 ;
  assign n8343 = n5026 & ~n8342 ;
  assign n8344 = ~\sub1_data_reg_reg[52]/NET0131  & ~n5026 ;
  assign n8345 = ~n8343 & ~n8344 ;
  assign n8346 = \state_reg/NET0131  & ~n8345 ;
  assign n8347 = ~\state_reg/NET0131  & ~n8336 ;
  assign n8348 = ~n8346 & ~n8347 ;
  assign n8350 = \key_i[52]_pad  & n8348 ;
  assign n8349 = ~\key_i[52]_pad  & ~n8348 ;
  assign n8351 = n933 & ~n8349 ;
  assign n8352 = ~n8350 & n8351 ;
  assign n8354 = ~\ks1_key_reg_reg[52]/NET0131  & ~n8348 ;
  assign n8355 = \ks1_key_reg_reg[52]/NET0131  & n8348 ;
  assign n8356 = ~n8354 & ~n8355 ;
  assign n8357 = n5053 & ~n8356 ;
  assign n8353 = ~\data_o[52]_pad  & ~n5053 ;
  assign n8358 = ~n933 & ~n8353 ;
  assign n8359 = ~n8357 & n8358 ;
  assign n8360 = ~n8352 & ~n8359 ;
  assign n8361 = ~\data_i[53]_pad  & ~n5029 ;
  assign n8362 = ~\mix1_data_o_reg_reg[53]/NET0131  & n5029 ;
  assign n8363 = ~n8361 & ~n8362 ;
  assign n8364 = ~n1159 & ~n8363 ;
  assign n8365 = ~\sub1_data_reg_reg[53]/NET0131  & n1159 ;
  assign n8366 = ~n8364 & ~n8365 ;
  assign n8367 = ~n5028 & ~n8366 ;
  assign n8368 = ~\sub1_data_reg_reg[53]/NET0131  & n5028 ;
  assign n8369 = ~n8367 & ~n8368 ;
  assign n8370 = ~n5027 & ~n8369 ;
  assign n8371 = ~\mix1_data_o_reg_reg[53]/NET0131  & n5027 ;
  assign n8372 = ~n8370 & ~n8371 ;
  assign n8373 = n5026 & ~n8372 ;
  assign n8374 = ~\sub1_data_reg_reg[53]/NET0131  & ~n5026 ;
  assign n8375 = ~n8373 & ~n8374 ;
  assign n8376 = \state_reg/NET0131  & ~n8375 ;
  assign n8377 = ~\state_reg/NET0131  & ~n8366 ;
  assign n8378 = ~n8376 & ~n8377 ;
  assign n8380 = \key_i[53]_pad  & n8378 ;
  assign n8379 = ~\key_i[53]_pad  & ~n8378 ;
  assign n8381 = n933 & ~n8379 ;
  assign n8382 = ~n8380 & n8381 ;
  assign n8384 = ~\ks1_key_reg_reg[53]/NET0131  & ~n8378 ;
  assign n8385 = \ks1_key_reg_reg[53]/NET0131  & n8378 ;
  assign n8386 = ~n8384 & ~n8385 ;
  assign n8387 = n5053 & ~n8386 ;
  assign n8383 = ~\data_o[53]_pad  & ~n5053 ;
  assign n8388 = ~n933 & ~n8383 ;
  assign n8389 = ~n8387 & n8388 ;
  assign n8390 = ~n8382 & ~n8389 ;
  assign n8391 = \data_i[14]_pad  & ~n5029 ;
  assign n8392 = \mix1_data_o_reg_reg[14]/NET0131  & n5029 ;
  assign n8393 = ~n8391 & ~n8392 ;
  assign n8394 = ~n1159 & ~n8393 ;
  assign n8395 = \sub1_data_reg_reg[14]/NET0131  & n1159 ;
  assign n8396 = ~n8394 & ~n8395 ;
  assign n8397 = ~n5028 & n8396 ;
  assign n8398 = ~\sub1_data_reg_reg[14]/NET0131  & n5028 ;
  assign n8399 = ~n8397 & ~n8398 ;
  assign n8400 = ~n5027 & ~n8399 ;
  assign n8401 = ~\mix1_data_o_reg_reg[14]/NET0131  & n5027 ;
  assign n8402 = ~n8400 & ~n8401 ;
  assign n8403 = n5026 & ~n8402 ;
  assign n8404 = ~\sub1_data_reg_reg[14]/NET0131  & ~n5026 ;
  assign n8405 = ~n8403 & ~n8404 ;
  assign n8406 = \state_reg/NET0131  & ~n8405 ;
  assign n8407 = ~\state_reg/NET0131  & n8396 ;
  assign n8408 = ~n8406 & ~n8407 ;
  assign n8410 = \key_i[14]_pad  & n8408 ;
  assign n8409 = ~\key_i[14]_pad  & ~n8408 ;
  assign n8411 = n933 & ~n8409 ;
  assign n8412 = ~n8410 & n8411 ;
  assign n8414 = ~\ks1_key_reg_reg[14]/NET0131  & ~n8408 ;
  assign n8415 = \ks1_key_reg_reg[14]/NET0131  & n8408 ;
  assign n8416 = ~n8414 & ~n8415 ;
  assign n8417 = n5053 & ~n8416 ;
  assign n8413 = ~\data_o[14]_pad  & ~n5053 ;
  assign n8418 = ~n933 & ~n8413 ;
  assign n8419 = ~n8417 & n8418 ;
  assign n8420 = ~n8412 & ~n8419 ;
  assign n8421 = ~\data_i[100]_pad  & ~n5029 ;
  assign n8422 = ~\mix1_data_o_reg_reg[100]/NET0131  & n5029 ;
  assign n8423 = ~n8421 & ~n8422 ;
  assign n8424 = ~n1159 & ~n8423 ;
  assign n8425 = ~\sub1_data_reg_reg[100]/NET0131  & n1159 ;
  assign n8426 = ~n8424 & ~n8425 ;
  assign n8427 = ~n5028 & ~n8426 ;
  assign n8428 = ~\sub1_data_reg_reg[100]/NET0131  & n5028 ;
  assign n8429 = ~n8427 & ~n8428 ;
  assign n8430 = ~n5027 & ~n8429 ;
  assign n8431 = ~\mix1_data_o_reg_reg[100]/NET0131  & n5027 ;
  assign n8432 = ~n8430 & ~n8431 ;
  assign n8433 = n5026 & ~n8432 ;
  assign n8434 = ~\sub1_data_reg_reg[100]/NET0131  & ~n5026 ;
  assign n8435 = ~n8433 & ~n8434 ;
  assign n8436 = \state_reg/NET0131  & ~n8435 ;
  assign n8437 = ~\state_reg/NET0131  & ~n8426 ;
  assign n8438 = ~n8436 & ~n8437 ;
  assign n8440 = \key_i[100]_pad  & n8438 ;
  assign n8439 = ~\key_i[100]_pad  & ~n8438 ;
  assign n8441 = n933 & ~n8439 ;
  assign n8442 = ~n8440 & n8441 ;
  assign n8444 = ~\ks1_key_reg_reg[100]/NET0131  & ~n8438 ;
  assign n8445 = \ks1_key_reg_reg[100]/NET0131  & n8438 ;
  assign n8446 = ~n8444 & ~n8445 ;
  assign n8447 = n5053 & ~n8446 ;
  assign n8443 = ~\data_o[100]_pad  & ~n5053 ;
  assign n8448 = ~n933 & ~n8443 ;
  assign n8449 = ~n8447 & n8448 ;
  assign n8450 = ~n8442 & ~n8449 ;
  assign n8451 = ~\data_i[54]_pad  & ~n5029 ;
  assign n8452 = ~\mix1_data_o_reg_reg[54]/NET0131  & n5029 ;
  assign n8453 = ~n8451 & ~n8452 ;
  assign n8454 = ~n1159 & ~n8453 ;
  assign n8455 = ~\sub1_data_reg_reg[54]/NET0131  & n1159 ;
  assign n8456 = ~n8454 & ~n8455 ;
  assign n8457 = ~n5028 & ~n8456 ;
  assign n8458 = ~\sub1_data_reg_reg[54]/NET0131  & n5028 ;
  assign n8459 = ~n8457 & ~n8458 ;
  assign n8460 = ~n5027 & ~n8459 ;
  assign n8461 = ~\mix1_data_o_reg_reg[54]/NET0131  & n5027 ;
  assign n8462 = ~n8460 & ~n8461 ;
  assign n8463 = n5026 & ~n8462 ;
  assign n8464 = ~\sub1_data_reg_reg[54]/NET0131  & ~n5026 ;
  assign n8465 = ~n8463 & ~n8464 ;
  assign n8466 = \state_reg/NET0131  & ~n8465 ;
  assign n8467 = ~\state_reg/NET0131  & ~n8456 ;
  assign n8468 = ~n8466 & ~n8467 ;
  assign n8470 = \key_i[54]_pad  & n8468 ;
  assign n8469 = ~\key_i[54]_pad  & ~n8468 ;
  assign n8471 = n933 & ~n8469 ;
  assign n8472 = ~n8470 & n8471 ;
  assign n8474 = ~\ks1_key_reg_reg[54]/NET0131  & ~n8468 ;
  assign n8475 = \ks1_key_reg_reg[54]/NET0131  & n8468 ;
  assign n8476 = ~n8474 & ~n8475 ;
  assign n8477 = n5053 & ~n8476 ;
  assign n8473 = ~\data_o[54]_pad  & ~n5053 ;
  assign n8478 = ~n933 & ~n8473 ;
  assign n8479 = ~n8477 & n8478 ;
  assign n8480 = ~n8472 & ~n8479 ;
  assign n8481 = ~\data_i[55]_pad  & ~n5029 ;
  assign n8482 = ~\mix1_data_o_reg_reg[55]/NET0131  & n5029 ;
  assign n8483 = ~n8481 & ~n8482 ;
  assign n8484 = ~n1159 & ~n8483 ;
  assign n8485 = ~\sub1_data_reg_reg[55]/NET0131  & n1159 ;
  assign n8486 = ~n8484 & ~n8485 ;
  assign n8487 = ~n5028 & ~n8486 ;
  assign n8488 = ~\sub1_data_reg_reg[55]/NET0131  & n5028 ;
  assign n8489 = ~n8487 & ~n8488 ;
  assign n8490 = ~n5027 & ~n8489 ;
  assign n8491 = ~\mix1_data_o_reg_reg[55]/NET0131  & n5027 ;
  assign n8492 = ~n8490 & ~n8491 ;
  assign n8493 = n5026 & ~n8492 ;
  assign n8494 = ~\sub1_data_reg_reg[55]/NET0131  & ~n5026 ;
  assign n8495 = ~n8493 & ~n8494 ;
  assign n8496 = \state_reg/NET0131  & ~n8495 ;
  assign n8497 = ~\state_reg/NET0131  & ~n8486 ;
  assign n8498 = ~n8496 & ~n8497 ;
  assign n8500 = \key_i[55]_pad  & n8498 ;
  assign n8499 = ~\key_i[55]_pad  & ~n8498 ;
  assign n8501 = n933 & ~n8499 ;
  assign n8502 = ~n8500 & n8501 ;
  assign n8504 = ~\ks1_key_reg_reg[55]/NET0131  & ~n8498 ;
  assign n8505 = \ks1_key_reg_reg[55]/NET0131  & n8498 ;
  assign n8506 = ~n8504 & ~n8505 ;
  assign n8507 = n5053 & ~n8506 ;
  assign n8503 = ~\data_o[55]_pad  & ~n5053 ;
  assign n8508 = ~n933 & ~n8503 ;
  assign n8509 = ~n8507 & n8508 ;
  assign n8510 = ~n8502 & ~n8509 ;
  assign n8511 = \data_i[15]_pad  & ~n5029 ;
  assign n8512 = \mix1_data_o_reg_reg[15]/NET0131  & n5029 ;
  assign n8513 = ~n8511 & ~n8512 ;
  assign n8514 = ~n1159 & ~n8513 ;
  assign n8515 = \sub1_data_reg_reg[15]/NET0131  & n1159 ;
  assign n8516 = ~n8514 & ~n8515 ;
  assign n8517 = ~n5028 & n8516 ;
  assign n8518 = ~\sub1_data_reg_reg[15]/NET0131  & n5028 ;
  assign n8519 = ~n8517 & ~n8518 ;
  assign n8520 = ~n5027 & ~n8519 ;
  assign n8521 = ~\mix1_data_o_reg_reg[15]/NET0131  & n5027 ;
  assign n8522 = ~n8520 & ~n8521 ;
  assign n8523 = n5026 & ~n8522 ;
  assign n8524 = ~\sub1_data_reg_reg[15]/NET0131  & ~n5026 ;
  assign n8525 = ~n8523 & ~n8524 ;
  assign n8526 = \state_reg/NET0131  & ~n8525 ;
  assign n8527 = ~\state_reg/NET0131  & n8516 ;
  assign n8528 = ~n8526 & ~n8527 ;
  assign n8530 = \key_i[15]_pad  & n8528 ;
  assign n8529 = ~\key_i[15]_pad  & ~n8528 ;
  assign n8531 = n933 & ~n8529 ;
  assign n8532 = ~n8530 & n8531 ;
  assign n8534 = ~\ks1_key_reg_reg[15]/NET0131  & ~n8528 ;
  assign n8535 = \ks1_key_reg_reg[15]/NET0131  & n8528 ;
  assign n8536 = ~n8534 & ~n8535 ;
  assign n8537 = n5053 & ~n8536 ;
  assign n8533 = ~\data_o[15]_pad  & ~n5053 ;
  assign n8538 = ~n933 & ~n8533 ;
  assign n8539 = ~n8537 & n8538 ;
  assign n8540 = ~n8532 & ~n8539 ;
  assign n8541 = \data_i[110]_pad  & ~n5029 ;
  assign n8542 = \mix1_data_o_reg_reg[110]/NET0131  & n5029 ;
  assign n8543 = ~n8541 & ~n8542 ;
  assign n8544 = ~n1159 & ~n8543 ;
  assign n8545 = \sub1_data_reg_reg[110]/NET0131  & n1159 ;
  assign n8546 = ~n8544 & ~n8545 ;
  assign n8547 = ~n5028 & n8546 ;
  assign n8548 = ~\sub1_data_reg_reg[110]/NET0131  & n5028 ;
  assign n8549 = ~n8547 & ~n8548 ;
  assign n8550 = ~n5027 & ~n8549 ;
  assign n8551 = ~\mix1_data_o_reg_reg[110]/NET0131  & n5027 ;
  assign n8552 = ~n8550 & ~n8551 ;
  assign n8553 = n5026 & ~n8552 ;
  assign n8554 = ~\sub1_data_reg_reg[110]/NET0131  & ~n5026 ;
  assign n8555 = ~n8553 & ~n8554 ;
  assign n8556 = \state_reg/NET0131  & ~n8555 ;
  assign n8557 = ~\state_reg/NET0131  & n8546 ;
  assign n8558 = ~n8556 & ~n8557 ;
  assign n8560 = \key_i[110]_pad  & n8558 ;
  assign n8559 = ~\key_i[110]_pad  & ~n8558 ;
  assign n8561 = n933 & ~n8559 ;
  assign n8562 = ~n8560 & n8561 ;
  assign n8564 = ~\ks1_key_reg_reg[110]/P0002  & ~n8558 ;
  assign n8565 = \ks1_key_reg_reg[110]/P0002  & n8558 ;
  assign n8566 = ~n8564 & ~n8565 ;
  assign n8567 = n5053 & ~n8566 ;
  assign n8563 = ~\data_o[110]_pad  & ~n5053 ;
  assign n8568 = ~n933 & ~n8563 ;
  assign n8569 = ~n8567 & n8568 ;
  assign n8570 = ~n8562 & ~n8569 ;
  assign n8571 = \data_i[56]_pad  & ~n5029 ;
  assign n8572 = \mix1_data_o_reg_reg[56]/NET0131  & n5029 ;
  assign n8573 = ~n8571 & ~n8572 ;
  assign n8574 = ~n1159 & ~n8573 ;
  assign n8575 = \sub1_data_reg_reg[56]/NET0131  & n1159 ;
  assign n8576 = ~n8574 & ~n8575 ;
  assign n8577 = ~n5028 & n8576 ;
  assign n8578 = ~\sub1_data_reg_reg[56]/NET0131  & n5028 ;
  assign n8579 = ~n8577 & ~n8578 ;
  assign n8580 = ~n5027 & ~n8579 ;
  assign n8581 = ~\mix1_data_o_reg_reg[56]/NET0131  & n5027 ;
  assign n8582 = ~n8580 & ~n8581 ;
  assign n8583 = n5026 & ~n8582 ;
  assign n8584 = ~\sub1_data_reg_reg[56]/NET0131  & ~n5026 ;
  assign n8585 = ~n8583 & ~n8584 ;
  assign n8586 = \state_reg/NET0131  & ~n8585 ;
  assign n8587 = ~\state_reg/NET0131  & n8576 ;
  assign n8588 = ~n8586 & ~n8587 ;
  assign n8590 = \key_i[56]_pad  & n8588 ;
  assign n8589 = ~\key_i[56]_pad  & ~n8588 ;
  assign n8591 = n933 & ~n8589 ;
  assign n8592 = ~n8590 & n8591 ;
  assign n8594 = ~\ks1_key_reg_reg[56]/NET0131  & ~n8588 ;
  assign n8595 = \ks1_key_reg_reg[56]/NET0131  & n8588 ;
  assign n8596 = ~n8594 & ~n8595 ;
  assign n8597 = n5053 & ~n8596 ;
  assign n8593 = ~\data_o[56]_pad  & ~n5053 ;
  assign n8598 = ~n933 & ~n8593 ;
  assign n8599 = ~n8597 & n8598 ;
  assign n8600 = ~n8592 & ~n8599 ;
  assign n8601 = \data_i[57]_pad  & ~n5029 ;
  assign n8602 = \mix1_data_o_reg_reg[57]/NET0131  & n5029 ;
  assign n8603 = ~n8601 & ~n8602 ;
  assign n8604 = ~n1159 & ~n8603 ;
  assign n8605 = \sub1_data_reg_reg[57]/NET0131  & n1159 ;
  assign n8606 = ~n8604 & ~n8605 ;
  assign n8607 = ~n5028 & n8606 ;
  assign n8608 = ~\sub1_data_reg_reg[57]/NET0131  & n5028 ;
  assign n8609 = ~n8607 & ~n8608 ;
  assign n8610 = ~n5027 & ~n8609 ;
  assign n8611 = ~\mix1_data_o_reg_reg[57]/NET0131  & n5027 ;
  assign n8612 = ~n8610 & ~n8611 ;
  assign n8613 = n5026 & ~n8612 ;
  assign n8614 = ~\sub1_data_reg_reg[57]/NET0131  & ~n5026 ;
  assign n8615 = ~n8613 & ~n8614 ;
  assign n8616 = \state_reg/NET0131  & ~n8615 ;
  assign n8617 = ~\state_reg/NET0131  & n8606 ;
  assign n8618 = ~n8616 & ~n8617 ;
  assign n8620 = \key_i[57]_pad  & n8618 ;
  assign n8619 = ~\key_i[57]_pad  & ~n8618 ;
  assign n8621 = n933 & ~n8619 ;
  assign n8622 = ~n8620 & n8621 ;
  assign n8624 = ~\ks1_key_reg_reg[57]/NET0131  & ~n8618 ;
  assign n8625 = \ks1_key_reg_reg[57]/NET0131  & n8618 ;
  assign n8626 = ~n8624 & ~n8625 ;
  assign n8627 = n5053 & ~n8626 ;
  assign n8623 = ~\data_o[57]_pad  & ~n5053 ;
  assign n8628 = ~n933 & ~n8623 ;
  assign n8629 = ~n8627 & n8628 ;
  assign n8630 = ~n8622 & ~n8629 ;
  assign n8631 = ~\data_i[16]_pad  & ~n5029 ;
  assign n8632 = ~\mix1_data_o_reg_reg[16]/NET0131  & n5029 ;
  assign n8633 = ~n8631 & ~n8632 ;
  assign n8634 = ~n1159 & ~n8633 ;
  assign n8635 = ~\sub1_data_reg_reg[16]/NET0131  & n1159 ;
  assign n8636 = ~n8634 & ~n8635 ;
  assign n8637 = ~n5028 & ~n8636 ;
  assign n8638 = ~\sub1_data_reg_reg[16]/NET0131  & n5028 ;
  assign n8639 = ~n8637 & ~n8638 ;
  assign n8640 = ~n5027 & ~n8639 ;
  assign n8641 = ~\mix1_data_o_reg_reg[16]/NET0131  & n5027 ;
  assign n8642 = ~n8640 & ~n8641 ;
  assign n8643 = n5026 & ~n8642 ;
  assign n8644 = ~\sub1_data_reg_reg[16]/NET0131  & ~n5026 ;
  assign n8645 = ~n8643 & ~n8644 ;
  assign n8646 = \state_reg/NET0131  & ~n8645 ;
  assign n8647 = ~\state_reg/NET0131  & ~n8636 ;
  assign n8648 = ~n8646 & ~n8647 ;
  assign n8650 = \key_i[16]_pad  & n8648 ;
  assign n8649 = ~\key_i[16]_pad  & ~n8648 ;
  assign n8651 = n933 & ~n8649 ;
  assign n8652 = ~n8650 & n8651 ;
  assign n8654 = ~\ks1_key_reg_reg[16]/NET0131  & ~n8648 ;
  assign n8655 = \ks1_key_reg_reg[16]/NET0131  & n8648 ;
  assign n8656 = ~n8654 & ~n8655 ;
  assign n8657 = n5053 & ~n8656 ;
  assign n8653 = ~\data_o[16]_pad  & ~n5053 ;
  assign n8658 = ~n933 & ~n8653 ;
  assign n8659 = ~n8657 & n8658 ;
  assign n8660 = ~n8652 & ~n8659 ;
  assign n8661 = \data_i[58]_pad  & ~n5029 ;
  assign n8662 = \mix1_data_o_reg_reg[58]/NET0131  & n5029 ;
  assign n8663 = ~n8661 & ~n8662 ;
  assign n8664 = ~n1159 & ~n8663 ;
  assign n8665 = \sub1_data_reg_reg[58]/NET0131  & n1159 ;
  assign n8666 = ~n8664 & ~n8665 ;
  assign n8667 = ~n5028 & n8666 ;
  assign n8668 = ~\sub1_data_reg_reg[58]/NET0131  & n5028 ;
  assign n8669 = ~n8667 & ~n8668 ;
  assign n8670 = ~n5027 & ~n8669 ;
  assign n8671 = ~\mix1_data_o_reg_reg[58]/NET0131  & n5027 ;
  assign n8672 = ~n8670 & ~n8671 ;
  assign n8673 = n5026 & ~n8672 ;
  assign n8674 = ~\sub1_data_reg_reg[58]/NET0131  & ~n5026 ;
  assign n8675 = ~n8673 & ~n8674 ;
  assign n8676 = \state_reg/NET0131  & ~n8675 ;
  assign n8677 = ~\state_reg/NET0131  & n8666 ;
  assign n8678 = ~n8676 & ~n8677 ;
  assign n8680 = \key_i[58]_pad  & n8678 ;
  assign n8679 = ~\key_i[58]_pad  & ~n8678 ;
  assign n8681 = n933 & ~n8679 ;
  assign n8682 = ~n8680 & n8681 ;
  assign n8684 = ~\ks1_key_reg_reg[58]/NET0131  & ~n8678 ;
  assign n8685 = \ks1_key_reg_reg[58]/NET0131  & n8678 ;
  assign n8686 = ~n8684 & ~n8685 ;
  assign n8687 = n5053 & ~n8686 ;
  assign n8683 = ~\data_o[58]_pad  & ~n5053 ;
  assign n8688 = ~n933 & ~n8683 ;
  assign n8689 = ~n8687 & n8688 ;
  assign n8690 = ~n8682 & ~n8689 ;
  assign n8691 = \data_i[59]_pad  & ~n5029 ;
  assign n8692 = \mix1_data_o_reg_reg[59]/NET0131  & n5029 ;
  assign n8693 = ~n8691 & ~n8692 ;
  assign n8694 = ~n1159 & ~n8693 ;
  assign n8695 = \sub1_data_reg_reg[59]/NET0131  & n1159 ;
  assign n8696 = ~n8694 & ~n8695 ;
  assign n8697 = ~n5028 & n8696 ;
  assign n8698 = ~\sub1_data_reg_reg[59]/NET0131  & n5028 ;
  assign n8699 = ~n8697 & ~n8698 ;
  assign n8700 = ~n5027 & ~n8699 ;
  assign n8701 = ~\mix1_data_o_reg_reg[59]/NET0131  & n5027 ;
  assign n8702 = ~n8700 & ~n8701 ;
  assign n8703 = n5026 & ~n8702 ;
  assign n8704 = ~\sub1_data_reg_reg[59]/NET0131  & ~n5026 ;
  assign n8705 = ~n8703 & ~n8704 ;
  assign n8706 = \state_reg/NET0131  & ~n8705 ;
  assign n8707 = ~\state_reg/NET0131  & n8696 ;
  assign n8708 = ~n8706 & ~n8707 ;
  assign n8710 = \key_i[59]_pad  & n8708 ;
  assign n8709 = ~\key_i[59]_pad  & ~n8708 ;
  assign n8711 = n933 & ~n8709 ;
  assign n8712 = ~n8710 & n8711 ;
  assign n8714 = ~\ks1_key_reg_reg[59]/NET0131  & ~n8708 ;
  assign n8715 = \ks1_key_reg_reg[59]/NET0131  & n8708 ;
  assign n8716 = ~n8714 & ~n8715 ;
  assign n8717 = n5053 & ~n8716 ;
  assign n8713 = ~\data_o[59]_pad  & ~n5053 ;
  assign n8718 = ~n933 & ~n8713 ;
  assign n8719 = ~n8717 & n8718 ;
  assign n8720 = ~n8712 & ~n8719 ;
  assign n8721 = \data_i[111]_pad  & ~n5029 ;
  assign n8722 = \mix1_data_o_reg_reg[111]/NET0131  & n5029 ;
  assign n8723 = ~n8721 & ~n8722 ;
  assign n8724 = ~n1159 & ~n8723 ;
  assign n8725 = \sub1_data_reg_reg[111]/NET0131  & n1159 ;
  assign n8726 = ~n8724 & ~n8725 ;
  assign n8727 = ~n5028 & n8726 ;
  assign n8728 = ~\sub1_data_reg_reg[111]/NET0131  & n5028 ;
  assign n8729 = ~n8727 & ~n8728 ;
  assign n8730 = ~n5027 & ~n8729 ;
  assign n8731 = ~\mix1_data_o_reg_reg[111]/NET0131  & n5027 ;
  assign n8732 = ~n8730 & ~n8731 ;
  assign n8733 = n5026 & ~n8732 ;
  assign n8734 = ~\sub1_data_reg_reg[111]/NET0131  & ~n5026 ;
  assign n8735 = ~n8733 & ~n8734 ;
  assign n8736 = \state_reg/NET0131  & ~n8735 ;
  assign n8737 = ~\state_reg/NET0131  & n8726 ;
  assign n8738 = ~n8736 & ~n8737 ;
  assign n8740 = \key_i[111]_pad  & n8738 ;
  assign n8739 = ~\key_i[111]_pad  & ~n8738 ;
  assign n8741 = n933 & ~n8739 ;
  assign n8742 = ~n8740 & n8741 ;
  assign n8744 = ~\ks1_key_reg_reg[111]/NET0131  & ~n8738 ;
  assign n8745 = \ks1_key_reg_reg[111]/NET0131  & n8738 ;
  assign n8746 = ~n8744 & ~n8745 ;
  assign n8747 = n5053 & ~n8746 ;
  assign n8743 = ~\data_o[111]_pad  & ~n5053 ;
  assign n8748 = ~n933 & ~n8743 ;
  assign n8749 = ~n8747 & n8748 ;
  assign n8750 = ~n8742 & ~n8749 ;
  assign n8751 = ~\data_i[17]_pad  & ~n5029 ;
  assign n8752 = ~\mix1_data_o_reg_reg[17]/NET0131  & n5029 ;
  assign n8753 = ~n8751 & ~n8752 ;
  assign n8754 = ~n1159 & ~n8753 ;
  assign n8755 = ~\sub1_data_reg_reg[17]/NET0131  & n1159 ;
  assign n8756 = ~n8754 & ~n8755 ;
  assign n8757 = ~n5028 & ~n8756 ;
  assign n8758 = ~\sub1_data_reg_reg[17]/NET0131  & n5028 ;
  assign n8759 = ~n8757 & ~n8758 ;
  assign n8760 = ~n5027 & ~n8759 ;
  assign n8761 = ~\mix1_data_o_reg_reg[17]/NET0131  & n5027 ;
  assign n8762 = ~n8760 & ~n8761 ;
  assign n8763 = n5026 & ~n8762 ;
  assign n8764 = ~\sub1_data_reg_reg[17]/NET0131  & ~n5026 ;
  assign n8765 = ~n8763 & ~n8764 ;
  assign n8766 = \state_reg/NET0131  & ~n8765 ;
  assign n8767 = ~\state_reg/NET0131  & ~n8756 ;
  assign n8768 = ~n8766 & ~n8767 ;
  assign n8770 = \key_i[17]_pad  & n8768 ;
  assign n8769 = ~\key_i[17]_pad  & ~n8768 ;
  assign n8771 = n933 & ~n8769 ;
  assign n8772 = ~n8770 & n8771 ;
  assign n8774 = ~\ks1_key_reg_reg[17]/NET0131  & ~n8768 ;
  assign n8775 = \ks1_key_reg_reg[17]/NET0131  & n8768 ;
  assign n8776 = ~n8774 & ~n8775 ;
  assign n8777 = n5053 & ~n8776 ;
  assign n8773 = ~\data_o[17]_pad  & ~n5053 ;
  assign n8778 = ~n933 & ~n8773 ;
  assign n8779 = ~n8777 & n8778 ;
  assign n8780 = ~n8772 & ~n8779 ;
  assign n8781 = \data_i[5]_pad  & ~n5029 ;
  assign n8782 = \mix1_data_o_reg_reg[5]/NET0131  & n5029 ;
  assign n8783 = ~n8781 & ~n8782 ;
  assign n8784 = ~n1159 & ~n8783 ;
  assign n8785 = \sub1_data_reg_reg[5]/NET0131  & n1159 ;
  assign n8786 = ~n8784 & ~n8785 ;
  assign n8787 = ~n5028 & n8786 ;
  assign n8788 = ~\sub1_data_reg_reg[5]/NET0131  & n5028 ;
  assign n8789 = ~n8787 & ~n8788 ;
  assign n8790 = ~n5027 & ~n8789 ;
  assign n8791 = ~\mix1_data_o_reg_reg[5]/NET0131  & n5027 ;
  assign n8792 = ~n8790 & ~n8791 ;
  assign n8793 = n5026 & ~n8792 ;
  assign n8794 = ~\sub1_data_reg_reg[5]/NET0131  & ~n5026 ;
  assign n8795 = ~n8793 & ~n8794 ;
  assign n8796 = \state_reg/NET0131  & ~n8795 ;
  assign n8797 = ~\state_reg/NET0131  & n8786 ;
  assign n8798 = ~n8796 & ~n8797 ;
  assign n8800 = \key_i[5]_pad  & n8798 ;
  assign n8799 = ~\key_i[5]_pad  & ~n8798 ;
  assign n8801 = n933 & ~n8799 ;
  assign n8802 = ~n8800 & n8801 ;
  assign n8804 = ~\ks1_key_reg_reg[5]/NET0131  & ~n8798 ;
  assign n8805 = \ks1_key_reg_reg[5]/NET0131  & n8798 ;
  assign n8806 = ~n8804 & ~n8805 ;
  assign n8807 = n5053 & ~n8806 ;
  assign n8803 = ~\data_o[5]_pad  & ~n5053 ;
  assign n8808 = ~n933 & ~n8803 ;
  assign n8809 = ~n8807 & n8808 ;
  assign n8810 = ~n8802 & ~n8809 ;
  assign n8811 = \data_i[60]_pad  & ~n5029 ;
  assign n8812 = \mix1_data_o_reg_reg[60]/NET0131  & n5029 ;
  assign n8813 = ~n8811 & ~n8812 ;
  assign n8814 = ~n1159 & ~n8813 ;
  assign n8815 = \sub1_data_reg_reg[60]/NET0131  & n1159 ;
  assign n8816 = ~n8814 & ~n8815 ;
  assign n8817 = ~n5028 & n8816 ;
  assign n8818 = ~\sub1_data_reg_reg[60]/NET0131  & n5028 ;
  assign n8819 = ~n8817 & ~n8818 ;
  assign n8820 = ~n5027 & ~n8819 ;
  assign n8821 = ~\mix1_data_o_reg_reg[60]/NET0131  & n5027 ;
  assign n8822 = ~n8820 & ~n8821 ;
  assign n8823 = n5026 & ~n8822 ;
  assign n8824 = ~\sub1_data_reg_reg[60]/NET0131  & ~n5026 ;
  assign n8825 = ~n8823 & ~n8824 ;
  assign n8826 = \state_reg/NET0131  & ~n8825 ;
  assign n8827 = ~\state_reg/NET0131  & n8816 ;
  assign n8828 = ~n8826 & ~n8827 ;
  assign n8830 = \key_i[60]_pad  & n8828 ;
  assign n8829 = ~\key_i[60]_pad  & ~n8828 ;
  assign n8831 = n933 & ~n8829 ;
  assign n8832 = ~n8830 & n8831 ;
  assign n8834 = ~\ks1_key_reg_reg[60]/NET0131  & ~n8828 ;
  assign n8835 = \ks1_key_reg_reg[60]/NET0131  & n8828 ;
  assign n8836 = ~n8834 & ~n8835 ;
  assign n8837 = n5053 & ~n8836 ;
  assign n8833 = ~\data_o[60]_pad  & ~n5053 ;
  assign n8838 = ~n933 & ~n8833 ;
  assign n8839 = ~n8837 & n8838 ;
  assign n8840 = ~n8832 & ~n8839 ;
  assign n8841 = ~\data_i[18]_pad  & ~n5029 ;
  assign n8842 = ~\mix1_data_o_reg_reg[18]/NET0131  & n5029 ;
  assign n8843 = ~n8841 & ~n8842 ;
  assign n8844 = ~n1159 & ~n8843 ;
  assign n8845 = ~\sub1_data_reg_reg[18]/NET0131  & n1159 ;
  assign n8846 = ~n8844 & ~n8845 ;
  assign n8847 = ~n5028 & ~n8846 ;
  assign n8848 = ~\sub1_data_reg_reg[18]/NET0131  & n5028 ;
  assign n8849 = ~n8847 & ~n8848 ;
  assign n8850 = ~n5027 & ~n8849 ;
  assign n8851 = ~\mix1_data_o_reg_reg[18]/NET0131  & n5027 ;
  assign n8852 = ~n8850 & ~n8851 ;
  assign n8853 = n5026 & ~n8852 ;
  assign n8854 = ~\sub1_data_reg_reg[18]/NET0131  & ~n5026 ;
  assign n8855 = ~n8853 & ~n8854 ;
  assign n8856 = \state_reg/NET0131  & ~n8855 ;
  assign n8857 = ~\state_reg/NET0131  & ~n8846 ;
  assign n8858 = ~n8856 & ~n8857 ;
  assign n8860 = \key_i[18]_pad  & n8858 ;
  assign n8859 = ~\key_i[18]_pad  & ~n8858 ;
  assign n8861 = n933 & ~n8859 ;
  assign n8862 = ~n8860 & n8861 ;
  assign n8864 = ~\ks1_key_reg_reg[18]/NET0131  & ~n8858 ;
  assign n8865 = \ks1_key_reg_reg[18]/NET0131  & n8858 ;
  assign n8866 = ~n8864 & ~n8865 ;
  assign n8867 = n5053 & ~n8866 ;
  assign n8863 = ~\data_o[18]_pad  & ~n5053 ;
  assign n8868 = ~n933 & ~n8863 ;
  assign n8869 = ~n8867 & n8868 ;
  assign n8870 = ~n8862 & ~n8869 ;
  assign n8871 = \mix1_data_o_reg_reg[11]/NET0131  & ~n3640 ;
  assign n8872 = n3640 & ~n4387 ;
  assign n8873 = ~n8871 & ~n8872 ;
  assign n8874 = n3640 & ~n4448 ;
  assign n8875 = \mix1_data_o_reg_reg[12]/NET0131  & ~n3640 ;
  assign n8876 = ~n8874 & ~n8875 ;
  assign n8877 = n3640 & ~n4485 ;
  assign n8878 = \mix1_data_o_reg_reg[13]/NET0131  & ~n3640 ;
  assign n8879 = ~n8877 & ~n8878 ;
  assign n8880 = n3640 & ~n4528 ;
  assign n8881 = \mix1_data_o_reg_reg[19]/NET0131  & ~n3640 ;
  assign n8882 = ~n8880 & ~n8881 ;
  assign n8883 = n3640 & ~n4546 ;
  assign n8884 = ~\mix1_data_o_reg_reg[20]/NET0131  & ~n3640 ;
  assign n8885 = ~n8883 & ~n8884 ;
  assign n8886 = n3640 & ~n4571 ;
  assign n8887 = \mix1_data_o_reg_reg[21]/NET0131  & ~n3640 ;
  assign n8888 = ~n8886 & ~n8887 ;
  assign n8889 = \mix1_data_o_reg_reg[27]/NET0131  & ~n3640 ;
  assign n8890 = n3640 & ~n4581 ;
  assign n8891 = ~n8889 & ~n8890 ;
  assign n8892 = n3640 & ~n4617 ;
  assign n8893 = ~\mix1_data_o_reg_reg[28]/NET0131  & ~n3640 ;
  assign n8894 = ~n8892 & ~n8893 ;
  assign n8895 = n3640 & ~n4602 ;
  assign n8896 = \mix1_data_o_reg_reg[29]/NET0131  & ~n3640 ;
  assign n8897 = ~n8895 & ~n8896 ;
  assign n8898 = n3640 & n4623 ;
  assign n8899 = \mix1_data_o_reg_reg[3]/NET0131  & ~n3640 ;
  assign n8900 = ~n8898 & ~n8899 ;
  assign n8901 = n3640 & ~n4073 ;
  assign n8902 = \mix1_data_o_reg_reg[4]/NET0131  & ~n3640 ;
  assign n8903 = ~n8901 & ~n8902 ;
  assign n8904 = n3640 & ~n4261 ;
  assign n8905 = \mix1_data_o_reg_reg[5]/NET0131  & ~n3640 ;
  assign n8906 = ~n8904 & ~n8905 ;
  assign n8907 = ~n4989 & ~n4994 ;
  assign n8908 = \ks1_col_reg[25]/NET0131  & ~n8907 ;
  assign n8909 = ~\ks1_col_reg[25]/NET0131  & n8907 ;
  assign n8910 = ~n8908 & ~n8909 ;
  assign n8911 = ~\ks1_key_reg_reg[121]/NET0131  & n1116 ;
  assign n8912 = ~\key_i[121]_pad  & ~n1116 ;
  assign n8913 = ~n8911 & ~n8912 ;
  assign n8914 = n8910 & ~n8913 ;
  assign n8915 = ~n8910 & n8913 ;
  assign n8916 = ~n8914 & ~n8915 ;
  assign n8917 = ~\ks1_key_reg_reg[89]/NET0131  & n1116 ;
  assign n8918 = ~\key_i[89]_pad  & ~n1116 ;
  assign n8919 = ~n8917 & ~n8918 ;
  assign n8920 = n8916 & ~n8919 ;
  assign n8921 = ~n8916 & n8919 ;
  assign n8922 = ~n8920 & ~n8921 ;
  assign n8923 = ~\ks1_key_reg_reg[57]/NET0131  & n1116 ;
  assign n8924 = ~\key_i[57]_pad  & ~n1116 ;
  assign n8925 = ~n8923 & ~n8924 ;
  assign n8926 = n8922 & ~n8925 ;
  assign n8927 = ~n8922 & n8925 ;
  assign n8928 = ~n8926 & ~n8927 ;
  assign n8929 = n1656 & n8928 ;
  assign n8930 = ~n1656 & ~n8928 ;
  assign n8931 = ~n8929 & ~n8930 ;
  assign n8932 = n4966 & ~n4974 ;
  assign n8933 = n4987 & n8932 ;
  assign n8934 = ~n4995 & ~n8933 ;
  assign n8935 = \ks1_col_reg[26]/NET0131  & ~n8934 ;
  assign n8936 = ~\ks1_col_reg[26]/NET0131  & n8934 ;
  assign n8937 = ~n8935 & ~n8936 ;
  assign n8938 = ~\ks1_key_reg_reg[122]/NET0131  & n1116 ;
  assign n8939 = ~\key_i[122]_pad  & ~n1116 ;
  assign n8940 = ~n8938 & ~n8939 ;
  assign n8941 = n8937 & ~n8940 ;
  assign n8942 = ~n8937 & n8940 ;
  assign n8943 = ~n8941 & ~n8942 ;
  assign n8944 = ~\ks1_key_reg_reg[90]/NET0131  & n1116 ;
  assign n8945 = ~\key_i[90]_pad  & ~n1116 ;
  assign n8946 = ~n8944 & ~n8945 ;
  assign n8947 = n8943 & ~n8946 ;
  assign n8948 = ~n8943 & n8946 ;
  assign n8949 = ~n8947 & ~n8948 ;
  assign n8950 = ~\ks1_key_reg_reg[58]/NET0131  & n1116 ;
  assign n8951 = ~\key_i[58]_pad  & ~n1116 ;
  assign n8952 = ~n8950 & ~n8951 ;
  assign n8953 = n8949 & ~n8952 ;
  assign n8954 = ~n8949 & n8952 ;
  assign n8955 = ~n8953 & ~n8954 ;
  assign n8956 = n1937 & n8955 ;
  assign n8957 = ~n1937 & ~n8955 ;
  assign n8958 = ~n8956 & ~n8957 ;
  assign n8959 = n4978 & n4990 ;
  assign n8960 = n4974 & n8959 ;
  assign n8961 = ~n4989 & ~n8960 ;
  assign n8962 = \ks1_col_reg[27]/NET0131  & ~n8961 ;
  assign n8963 = ~\ks1_col_reg[27]/NET0131  & n8961 ;
  assign n8964 = ~n8962 & ~n8963 ;
  assign n8965 = ~\ks1_key_reg_reg[123]/NET0131  & n1116 ;
  assign n8966 = ~\key_i[123]_pad  & ~n1116 ;
  assign n8967 = ~n8965 & ~n8966 ;
  assign n8968 = n8964 & ~n8967 ;
  assign n8969 = ~n8964 & n8967 ;
  assign n8970 = ~n8968 & ~n8969 ;
  assign n8971 = ~\ks1_key_reg_reg[91]/NET0131  & n1116 ;
  assign n8972 = ~\key_i[91]_pad  & ~n1116 ;
  assign n8973 = ~n8971 & ~n8972 ;
  assign n8974 = n8970 & ~n8973 ;
  assign n8975 = ~n8970 & n8973 ;
  assign n8976 = ~n8974 & ~n8975 ;
  assign n8977 = ~\ks1_key_reg_reg[59]/NET0131  & n1116 ;
  assign n8978 = ~\key_i[59]_pad  & ~n1116 ;
  assign n8979 = ~n8977 & ~n8978 ;
  assign n8980 = n8976 & ~n8979 ;
  assign n8981 = ~n8976 & n8979 ;
  assign n8982 = ~n8980 & ~n8981 ;
  assign n8983 = n1537 & n8982 ;
  assign n8984 = ~n1537 & ~n8982 ;
  assign n8985 = ~n8983 & ~n8984 ;
  assign n8986 = ~n4974 & n8959 ;
  assign n8987 = ~n4995 & ~n8986 ;
  assign n8988 = \ks1_col_reg[29]/NET0131  & ~n8987 ;
  assign n8989 = ~\ks1_col_reg[29]/NET0131  & n8987 ;
  assign n8990 = ~n8988 & ~n8989 ;
  assign n8991 = ~\ks1_key_reg_reg[125]/NET0131  & n1116 ;
  assign n8992 = ~\key_i[125]_pad  & ~n1116 ;
  assign n8993 = ~n8991 & ~n8992 ;
  assign n8994 = n8990 & ~n8993 ;
  assign n8995 = ~n8990 & n8993 ;
  assign n8996 = ~n8994 & ~n8995 ;
  assign n8997 = ~\ks1_key_reg_reg[93]/NET0131  & n1116 ;
  assign n8998 = ~\key_i[93]_pad  & ~n1116 ;
  assign n8999 = ~n8997 & ~n8998 ;
  assign n9000 = n8996 & ~n8999 ;
  assign n9001 = ~n8996 & n8999 ;
  assign n9002 = ~n9000 & ~n9001 ;
  assign n9003 = ~\ks1_key_reg_reg[61]/NET0131  & n1116 ;
  assign n9004 = ~\key_i[61]_pad  & ~n1116 ;
  assign n9005 = ~n9003 & ~n9004 ;
  assign n9006 = n9002 & ~n9005 ;
  assign n9007 = ~n9002 & n9005 ;
  assign n9008 = ~n9006 & ~n9007 ;
  assign n9009 = n1901 & n9008 ;
  assign n9010 = ~n1901 & ~n9008 ;
  assign n9011 = ~n9009 & ~n9010 ;
  assign n9012 = \key_i[94]_pad  & ~n953 ;
  assign n9013 = \ks1_key_reg_reg[94]/NET0131  & n956 ;
  assign n9014 = ~n9012 & ~n9013 ;
  assign n9015 = ~n933 & ~n9014 ;
  assign n9017 = ~\key_i[94]_pad  & n951 ;
  assign n9016 = ~\ks1_key_reg_reg[94]/NET0131  & ~n951 ;
  assign n9018 = n933 & ~n9016 ;
  assign n9019 = ~n9017 & n9018 ;
  assign n9020 = ~n9015 & ~n9019 ;
  assign n9021 = ~n4974 & n4991 ;
  assign n9022 = \ks1_col_reg[30]/NET0131  & ~n9021 ;
  assign n9023 = ~\ks1_col_reg[30]/NET0131  & n9021 ;
  assign n9024 = ~n9022 & ~n9023 ;
  assign n9025 = ~\ks1_key_reg_reg[126]/NET0131  & n1116 ;
  assign n9026 = ~\key_i[126]_pad  & ~n1116 ;
  assign n9027 = ~n9025 & ~n9026 ;
  assign n9028 = n9024 & ~n9027 ;
  assign n9029 = ~n9024 & n9027 ;
  assign n9030 = ~n9028 & ~n9029 ;
  assign n9031 = n9020 & n9030 ;
  assign n9032 = ~n9020 & ~n9030 ;
  assign n9033 = ~n9031 & ~n9032 ;
  assign n9034 = ~\ks1_key_reg_reg[62]/NET0131  & n1116 ;
  assign n9035 = ~\key_i[62]_pad  & ~n1116 ;
  assign n9036 = ~n9034 & ~n9035 ;
  assign n9037 = n9033 & ~n9036 ;
  assign n9038 = ~n9033 & n9036 ;
  assign n9039 = ~n9037 & ~n9038 ;
  assign n9040 = n1402 & n9039 ;
  assign n9041 = ~n1402 & ~n9039 ;
  assign n9042 = ~n9040 & ~n9041 ;
  assign n9043 = \key_i[95]_pad  & ~n953 ;
  assign n9044 = \ks1_key_reg_reg[95]/NET0131  & n956 ;
  assign n9045 = ~n9043 & ~n9044 ;
  assign n9046 = ~n933 & ~n9045 ;
  assign n9048 = ~\key_i[95]_pad  & n951 ;
  assign n9047 = ~\ks1_key_reg_reg[95]/NET0131  & ~n951 ;
  assign n9049 = n933 & ~n9047 ;
  assign n9050 = ~n9048 & n9049 ;
  assign n9051 = ~n9046 & ~n9050 ;
  assign n9052 = ~n4966 & n4974 ;
  assign n9053 = n4993 & n9052 ;
  assign n9054 = \ks1_col_reg[31]/NET0131  & ~n9053 ;
  assign n9055 = ~\ks1_col_reg[31]/NET0131  & n9053 ;
  assign n9056 = ~n9054 & ~n9055 ;
  assign n9057 = ~\ks1_key_reg_reg[127]/NET0131  & n1116 ;
  assign n9058 = ~\key_i[127]_pad  & ~n1116 ;
  assign n9059 = ~n9057 & ~n9058 ;
  assign n9060 = n9056 & ~n9059 ;
  assign n9061 = ~n9056 & n9059 ;
  assign n9062 = ~n9060 & ~n9061 ;
  assign n9063 = n9051 & n9062 ;
  assign n9064 = ~n9051 & ~n9062 ;
  assign n9065 = ~n9063 & ~n9064 ;
  assign n9066 = ~\ks1_key_reg_reg[63]/NET0131  & n1116 ;
  assign n9067 = ~\key_i[63]_pad  & ~n1116 ;
  assign n9068 = ~n9066 & ~n9067 ;
  assign n9069 = n9065 & ~n9068 ;
  assign n9070 = ~n9065 & n9068 ;
  assign n9071 = ~n9069 & ~n9070 ;
  assign n9072 = n2094 & n9071 ;
  assign n9073 = ~n2094 & ~n9071 ;
  assign n9074 = ~n9072 & ~n9073 ;
  assign n9075 = \key_i[88]_pad  & ~n953 ;
  assign n9076 = \ks1_key_reg_reg[88]/NET0131  & n956 ;
  assign n9077 = ~n9075 & ~n9076 ;
  assign n9078 = ~n933 & ~n9077 ;
  assign n9080 = ~\key_i[88]_pad  & n951 ;
  assign n9079 = ~\ks1_key_reg_reg[88]/NET0131  & ~n951 ;
  assign n9081 = n933 & ~n9079 ;
  assign n9082 = ~n9080 & n9081 ;
  assign n9083 = ~n9078 & ~n9082 ;
  assign n9084 = \ks1_col_reg[24]/NET0131  & ~n4988 ;
  assign n9085 = ~\ks1_col_reg[24]/NET0131  & n4988 ;
  assign n9086 = ~n9084 & ~n9085 ;
  assign n9087 = ~\ks1_key_reg_reg[120]/NET0131  & n1116 ;
  assign n9088 = ~\key_i[120]_pad  & ~n1116 ;
  assign n9089 = ~n9087 & ~n9088 ;
  assign n9090 = n9086 & ~n9089 ;
  assign n9091 = ~n9086 & n9089 ;
  assign n9092 = ~n9090 & ~n9091 ;
  assign n9093 = n9083 & n9092 ;
  assign n9094 = ~n9083 & ~n9092 ;
  assign n9095 = ~n9093 & ~n9094 ;
  assign n9096 = ~\ks1_key_reg_reg[56]/NET0131  & n1116 ;
  assign n9097 = ~\key_i[56]_pad  & ~n1116 ;
  assign n9098 = ~n9096 & ~n9097 ;
  assign n9099 = n9095 & ~n9098 ;
  assign n9100 = ~n9095 & n9098 ;
  assign n9101 = ~n9099 & ~n9100 ;
  assign n9102 = n1781 & n9101 ;
  assign n9103 = ~n1781 & ~n9101 ;
  assign n9104 = ~n9102 & ~n9103 ;
  assign n9105 = decrypt_i_pad & ~n3821 ;
  assign n9106 = n4365 & ~n9105 ;
  assign n9107 = ~n4365 & n9105 ;
  assign n9108 = ~n9106 & ~n9107 ;
  assign n9109 = n4315 & n9108 ;
  assign n9110 = ~n4315 & ~n9108 ;
  assign n9111 = ~n9109 & ~n9110 ;
  assign n9112 = n3629 & ~n9111 ;
  assign n9113 = \mix1_data_reg_reg[104]/NET0131  & ~n3629 ;
  assign n9114 = ~n9112 & ~n9113 ;
  assign n9115 = decrypt_i_pad & ~n4494 ;
  assign n9116 = n4686 & ~n9115 ;
  assign n9117 = ~n4686 & n9115 ;
  assign n9118 = ~n9116 & ~n9117 ;
  assign n9119 = n4509 & n9118 ;
  assign n9120 = ~n4509 & ~n9118 ;
  assign n9121 = ~n9119 & ~n9120 ;
  assign n9122 = n3629 & n9121 ;
  assign n9123 = \mix1_data_reg_reg[112]/NET0131  & ~n3629 ;
  assign n9124 = ~n9122 & ~n9123 ;
  assign n9125 = ~n4324 & n9105 ;
  assign n9126 = n4324 & ~n9105 ;
  assign n9127 = ~n9125 & ~n9126 ;
  assign n9128 = n4312 & ~n9127 ;
  assign n9129 = ~n4312 & n9127 ;
  assign n9130 = ~n9128 & ~n9129 ;
  assign n9131 = n4506 & n9130 ;
  assign n9132 = ~n4506 & ~n9130 ;
  assign n9133 = ~n9131 & ~n9132 ;
  assign n9134 = n3629 & n9133 ;
  assign n9135 = \mix1_data_reg_reg[120]/NET0131  & ~n3629 ;
  assign n9136 = ~n9134 & ~n9135 ;
  assign n9137 = n3635 & ~n4952 ;
  assign n9138 = \mix1_data_reg_reg[33]/NET0131  & ~n3635 ;
  assign n9139 = ~n9137 & ~n9138 ;
  assign n9140 = n3635 & n4940 ;
  assign n9141 = \mix1_data_reg_reg[34]/NET0131  & ~n3635 ;
  assign n9142 = ~n9140 & ~n9141 ;
  assign n9143 = n3635 & ~n4648 ;
  assign n9144 = ~\mix1_data_reg_reg[38]/NET0131  & ~n3635 ;
  assign n9145 = ~n9143 & ~n9144 ;
  assign n9146 = n3635 & n4661 ;
  assign n9147 = \mix1_data_reg_reg[39]/NET0131  & ~n3635 ;
  assign n9148 = ~n9146 & ~n9147 ;
  assign n9149 = n3635 & ~n4674 ;
  assign n9150 = \mix1_data_reg_reg[41]/NET0131  & ~n3635 ;
  assign n9151 = ~n9149 & ~n9150 ;
  assign n9152 = n3635 & ~n4702 ;
  assign n9153 = ~\mix1_data_reg_reg[42]/NET0131  & ~n3635 ;
  assign n9154 = ~n9152 & ~n9153 ;
  assign n9155 = n3635 & n4727 ;
  assign n9156 = \mix1_data_reg_reg[46]/NET0131  & ~n3635 ;
  assign n9157 = ~n9155 & ~n9156 ;
  assign n9158 = n3635 & ~n4752 ;
  assign n9159 = ~\mix1_data_reg_reg[47]/NET0131  & ~n3635 ;
  assign n9160 = ~n9158 & ~n9159 ;
  assign n9161 = n3635 & ~n4771 ;
  assign n9162 = \mix1_data_reg_reg[49]/NET0131  & ~n3635 ;
  assign n9163 = ~n9161 & ~n9162 ;
  assign n9164 = \mix1_data_reg_reg[50]/NET0131  & ~n3635 ;
  assign n9165 = n3635 & ~n4794 ;
  assign n9166 = ~n9164 & ~n9165 ;
  assign n9167 = n3635 & ~n4808 ;
  assign n9168 = ~\mix1_data_reg_reg[54]/NET0131  & ~n3635 ;
  assign n9169 = ~n9167 & ~n9168 ;
  assign n9170 = n3635 & ~n4817 ;
  assign n9171 = \mix1_data_reg_reg[55]/NET0131  & ~n3635 ;
  assign n9172 = ~n9170 & ~n9171 ;
  assign n9173 = n3635 & n4823 ;
  assign n9174 = \mix1_data_reg_reg[57]/NET0131  & ~n3635 ;
  assign n9175 = ~n9173 & ~n9174 ;
  assign n9176 = n3635 & n4838 ;
  assign n9177 = \mix1_data_reg_reg[58]/NET0131  & ~n3635 ;
  assign n9178 = ~n9176 & ~n9177 ;
  assign n9179 = n3635 & n4847 ;
  assign n9180 = \mix1_data_reg_reg[62]/NET0131  & ~n3635 ;
  assign n9181 = ~n9179 & ~n9180 ;
  assign n9182 = n3635 & n4856 ;
  assign n9183 = \mix1_data_reg_reg[63]/NET0131  & ~n3635 ;
  assign n9184 = ~n9182 & ~n9183 ;
  assign n9185 = n3630 & ~n4952 ;
  assign n9186 = \mix1_data_reg_reg[65]/NET0131  & ~n3630 ;
  assign n9187 = ~n9185 & ~n9186 ;
  assign n9188 = n3630 & n4940 ;
  assign n9189 = \mix1_data_reg_reg[66]/NET0131  & ~n3630 ;
  assign n9190 = ~n9188 & ~n9189 ;
  assign n9191 = n3630 & ~n4648 ;
  assign n9192 = ~\mix1_data_reg_reg[70]/NET0131  & ~n3630 ;
  assign n9193 = ~n9191 & ~n9192 ;
  assign n9194 = n3630 & n4661 ;
  assign n9195 = \mix1_data_reg_reg[71]/NET0131  & ~n3630 ;
  assign n9196 = ~n9194 & ~n9195 ;
  assign n9197 = n3630 & ~n4674 ;
  assign n9198 = \mix1_data_reg_reg[73]/NET0131  & ~n3630 ;
  assign n9199 = ~n9197 & ~n9198 ;
  assign n9200 = n3630 & ~n4702 ;
  assign n9201 = ~\mix1_data_reg_reg[74]/NET0131  & ~n3630 ;
  assign n9202 = ~n9200 & ~n9201 ;
  assign n9203 = n3630 & n4727 ;
  assign n9204 = \mix1_data_reg_reg[78]/NET0131  & ~n3630 ;
  assign n9205 = ~n9203 & ~n9204 ;
  assign n9206 = n3630 & ~n4752 ;
  assign n9207 = ~\mix1_data_reg_reg[79]/NET0131  & ~n3630 ;
  assign n9208 = ~n9206 & ~n9207 ;
  assign n9209 = n3630 & ~n4771 ;
  assign n9210 = \mix1_data_reg_reg[81]/NET0131  & ~n3630 ;
  assign n9211 = ~n9209 & ~n9210 ;
  assign n9212 = \mix1_data_reg_reg[82]/NET0131  & ~n3630 ;
  assign n9213 = n3630 & ~n4794 ;
  assign n9214 = ~n9212 & ~n9213 ;
  assign n9215 = n3630 & ~n4808 ;
  assign n9216 = ~\mix1_data_reg_reg[86]/NET0131  & ~n3630 ;
  assign n9217 = ~n9215 & ~n9216 ;
  assign n9218 = n3630 & ~n4817 ;
  assign n9219 = \mix1_data_reg_reg[87]/NET0131  & ~n3630 ;
  assign n9220 = ~n9218 & ~n9219 ;
  assign n9221 = n3630 & n4823 ;
  assign n9222 = \mix1_data_reg_reg[89]/NET0131  & ~n3630 ;
  assign n9223 = ~n9221 & ~n9222 ;
  assign n9224 = n3630 & n4838 ;
  assign n9225 = \mix1_data_reg_reg[90]/NET0131  & ~n3630 ;
  assign n9226 = ~n9224 & ~n9225 ;
  assign n9227 = n3630 & n4847 ;
  assign n9228 = \mix1_data_reg_reg[94]/NET0131  & ~n3630 ;
  assign n9229 = ~n9227 & ~n9228 ;
  assign n9230 = n3630 & n4856 ;
  assign n9231 = \mix1_data_reg_reg[95]/NET0131  & ~n3630 ;
  assign n9232 = ~n9230 & ~n9231 ;
  assign n9233 = ~n4506 & n4689 ;
  assign n9234 = n4506 & ~n4689 ;
  assign n9235 = ~n9233 & ~n9234 ;
  assign n9236 = n9115 & n9235 ;
  assign n9237 = ~n9115 & ~n9235 ;
  assign n9238 = ~n9236 & ~n9237 ;
  assign n9239 = n3629 & ~n9238 ;
  assign n9240 = ~\mix1_data_reg_reg[96]/NET0131  & ~n3629 ;
  assign n9241 = ~n9239 & ~n9240 ;
  assign n9242 = n3640 & ~n4702 ;
  assign n9243 = ~\mix1_data_o_reg_reg[10]/NET0131  & ~n3640 ;
  assign n9244 = ~n9242 & ~n9243 ;
  assign n9245 = n3640 & n4727 ;
  assign n9246 = \mix1_data_o_reg_reg[14]/NET0131  & ~n3640 ;
  assign n9247 = ~n9245 & ~n9246 ;
  assign n9248 = n3640 & ~n4752 ;
  assign n9249 = ~\mix1_data_o_reg_reg[15]/NET0131  & ~n3640 ;
  assign n9250 = ~n9248 & ~n9249 ;
  assign n9251 = n3640 & ~n4771 ;
  assign n9252 = \mix1_data_o_reg_reg[17]/NET0131  & ~n3640 ;
  assign n9253 = ~n9251 & ~n9252 ;
  assign n9254 = \mix1_data_o_reg_reg[18]/NET0131  & ~n3640 ;
  assign n9255 = n3640 & ~n4794 ;
  assign n9256 = ~n9254 & ~n9255 ;
  assign n9257 = n3640 & ~n4952 ;
  assign n9258 = \mix1_data_o_reg_reg[1]/NET0131  & ~n3640 ;
  assign n9259 = ~n9257 & ~n9258 ;
  assign n9260 = n3640 & ~n4808 ;
  assign n9261 = ~\mix1_data_o_reg_reg[22]/NET0131  & ~n3640 ;
  assign n9262 = ~n9260 & ~n9261 ;
  assign n9263 = n3640 & ~n4817 ;
  assign n9264 = \mix1_data_o_reg_reg[23]/NET0131  & ~n3640 ;
  assign n9265 = ~n9263 & ~n9264 ;
  assign n9266 = n3640 & n4823 ;
  assign n9267 = \mix1_data_o_reg_reg[25]/NET0131  & ~n3640 ;
  assign n9268 = ~n9266 & ~n9267 ;
  assign n9269 = n3640 & n4838 ;
  assign n9270 = \mix1_data_o_reg_reg[26]/NET0131  & ~n3640 ;
  assign n9271 = ~n9269 & ~n9270 ;
  assign n9272 = n3640 & n4940 ;
  assign n9273 = \mix1_data_o_reg_reg[2]/NET0131  & ~n3640 ;
  assign n9274 = ~n9272 & ~n9273 ;
  assign n9275 = n3640 & n4847 ;
  assign n9276 = \mix1_data_o_reg_reg[30]/NET0131  & ~n3640 ;
  assign n9277 = ~n9275 & ~n9276 ;
  assign n9278 = n3640 & n4856 ;
  assign n9279 = \mix1_data_o_reg_reg[31]/NET0131  & ~n3640 ;
  assign n9280 = ~n9278 & ~n9279 ;
  assign n9281 = n3640 & ~n4648 ;
  assign n9282 = ~\mix1_data_o_reg_reg[6]/NET0131  & ~n3640 ;
  assign n9283 = ~n9281 & ~n9282 ;
  assign n9284 = n3640 & n4661 ;
  assign n9285 = \mix1_data_o_reg_reg[7]/NET0131  & ~n3640 ;
  assign n9286 = ~n9284 & ~n9285 ;
  assign n9287 = n3640 & ~n4674 ;
  assign n9288 = \mix1_data_o_reg_reg[9]/NET0131  & ~n3640 ;
  assign n9289 = ~n9287 & ~n9288 ;
  assign n9290 = n929 & n8949 ;
  assign n9291 = \ks1_key_reg_reg[90]/NET0131  & ~n929 ;
  assign n9292 = ~n9290 & ~n9291 ;
  assign n9293 = n929 & ~n9002 ;
  assign n9294 = ~\ks1_key_reg_reg[93]/NET0131  & ~n929 ;
  assign n9295 = ~n9293 & ~n9294 ;
  assign n9296 = n3635 & ~n9238 ;
  assign n9297 = ~\mix1_data_reg_reg[32]/NET0131  & ~n3635 ;
  assign n9298 = ~n9296 & ~n9297 ;
  assign n9299 = n3635 & ~n9111 ;
  assign n9300 = \mix1_data_reg_reg[40]/NET0131  & ~n3635 ;
  assign n9301 = ~n9299 & ~n9300 ;
  assign n9302 = n3635 & n9121 ;
  assign n9303 = \mix1_data_reg_reg[48]/NET0131  & ~n3635 ;
  assign n9304 = ~n9302 & ~n9303 ;
  assign n9305 = n3635 & n9133 ;
  assign n9306 = \mix1_data_reg_reg[56]/NET0131  & ~n3635 ;
  assign n9307 = ~n9305 & ~n9306 ;
  assign n9308 = n3630 & ~n9238 ;
  assign n9309 = ~\mix1_data_reg_reg[64]/NET0131  & ~n3630 ;
  assign n9310 = ~n9308 & ~n9309 ;
  assign n9311 = n3630 & ~n9111 ;
  assign n9312 = \mix1_data_reg_reg[72]/NET0131  & ~n3630 ;
  assign n9313 = ~n9311 & ~n9312 ;
  assign n9314 = n3630 & n9121 ;
  assign n9315 = \mix1_data_reg_reg[80]/NET0131  & ~n3630 ;
  assign n9316 = ~n9314 & ~n9315 ;
  assign n9317 = n3630 & n9133 ;
  assign n9318 = \mix1_data_reg_reg[88]/NET0131  & ~n3630 ;
  assign n9319 = ~n9317 & ~n9318 ;
  assign n9320 = \key_i[64]_pad  & ~n953 ;
  assign n9321 = \ks1_key_reg_reg[64]/NET0131  & n956 ;
  assign n9322 = ~n9320 & ~n9321 ;
  assign n9323 = ~n933 & ~n9322 ;
  assign n9325 = ~\key_i[64]_pad  & n951 ;
  assign n9324 = ~\ks1_key_reg_reg[64]/NET0131  & ~n951 ;
  assign n9326 = n933 & ~n9324 ;
  assign n9327 = ~n9325 & n9326 ;
  assign n9328 = ~n9323 & ~n9327 ;
  assign n9329 = ~\ks1_key_reg_reg[96]/NET0131  & n1116 ;
  assign n9330 = ~\key_i[96]_pad  & ~n1116 ;
  assign n9331 = ~n9329 & ~n9330 ;
  assign n9332 = \ks1_col_reg[0]/NET0131  & ~n9331 ;
  assign n9333 = ~\ks1_col_reg[0]/NET0131  & n9331 ;
  assign n9334 = ~n9332 & ~n9333 ;
  assign n9335 = n9328 & n9334 ;
  assign n9336 = ~n9328 & ~n9334 ;
  assign n9337 = ~n9335 & ~n9336 ;
  assign n9338 = ~\ks1_key_reg_reg[32]/NET0131  & n1116 ;
  assign n9339 = ~\key_i[32]_pad  & ~n1116 ;
  assign n9340 = ~n9338 & ~n9339 ;
  assign n9341 = n9337 & ~n9340 ;
  assign n9342 = ~n9337 & n9340 ;
  assign n9343 = ~n9341 & ~n9342 ;
  assign n9344 = n929 & ~n9343 ;
  assign n9345 = \ks1_key_reg_reg[32]/NET0131  & ~n929 ;
  assign n9346 = ~n9344 & ~n9345 ;
  assign n9347 = \key_i[65]_pad  & ~n953 ;
  assign n9348 = \ks1_key_reg_reg[65]/NET0131  & n956 ;
  assign n9349 = ~n9347 & ~n9348 ;
  assign n9350 = ~n933 & ~n9349 ;
  assign n9352 = ~\key_i[65]_pad  & n951 ;
  assign n9351 = ~\ks1_key_reg_reg[65]/NET0131  & ~n951 ;
  assign n9353 = n933 & ~n9351 ;
  assign n9354 = ~n9352 & n9353 ;
  assign n9355 = ~n9350 & ~n9354 ;
  assign n9356 = ~\ks1_key_reg_reg[97]/NET0131  & n1116 ;
  assign n9357 = ~\key_i[97]_pad  & ~n1116 ;
  assign n9358 = ~n9356 & ~n9357 ;
  assign n9359 = \ks1_col_reg[1]/NET0131  & ~n9358 ;
  assign n9360 = ~\ks1_col_reg[1]/NET0131  & n9358 ;
  assign n9361 = ~n9359 & ~n9360 ;
  assign n9362 = n9355 & n9361 ;
  assign n9363 = ~n9355 & ~n9361 ;
  assign n9364 = ~n9362 & ~n9363 ;
  assign n9365 = ~\ks1_key_reg_reg[33]/NET0131  & n1116 ;
  assign n9366 = ~\key_i[33]_pad  & ~n1116 ;
  assign n9367 = ~n9365 & ~n9366 ;
  assign n9368 = n9364 & ~n9367 ;
  assign n9369 = ~n9364 & n9367 ;
  assign n9370 = ~n9368 & ~n9369 ;
  assign n9371 = n929 & ~n9370 ;
  assign n9372 = \ks1_key_reg_reg[33]/NET0131  & ~n929 ;
  assign n9373 = ~n9371 & ~n9372 ;
  assign n9374 = \key_i[66]_pad  & ~n953 ;
  assign n9375 = \ks1_key_reg_reg[66]/NET0131  & n956 ;
  assign n9376 = ~n9374 & ~n9375 ;
  assign n9377 = ~n933 & ~n9376 ;
  assign n9379 = ~\key_i[66]_pad  & n951 ;
  assign n9378 = ~\ks1_key_reg_reg[66]/NET0131  & ~n951 ;
  assign n9380 = n933 & ~n9378 ;
  assign n9381 = ~n9379 & n9380 ;
  assign n9382 = ~n9377 & ~n9381 ;
  assign n9383 = ~\ks1_key_reg_reg[98]/NET0131  & n1116 ;
  assign n9384 = ~\key_i[98]_pad  & ~n1116 ;
  assign n9385 = ~n9383 & ~n9384 ;
  assign n9386 = \ks1_col_reg[2]/NET0131  & ~n9385 ;
  assign n9387 = ~\ks1_col_reg[2]/NET0131  & n9385 ;
  assign n9388 = ~n9386 & ~n9387 ;
  assign n9389 = n9382 & n9388 ;
  assign n9390 = ~n9382 & ~n9388 ;
  assign n9391 = ~n9389 & ~n9390 ;
  assign n9392 = ~\ks1_key_reg_reg[34]/NET0131  & n1116 ;
  assign n9393 = ~\key_i[34]_pad  & ~n1116 ;
  assign n9394 = ~n9392 & ~n9393 ;
  assign n9395 = n9391 & ~n9394 ;
  assign n9396 = ~n9391 & n9394 ;
  assign n9397 = ~n9395 & ~n9396 ;
  assign n9398 = n929 & ~n9397 ;
  assign n9399 = \ks1_key_reg_reg[34]/NET0131  & ~n929 ;
  assign n9400 = ~n9398 & ~n9399 ;
  assign n9401 = ~\ks1_key_reg_reg[99]/NET0131  & n1116 ;
  assign n9402 = ~\key_i[99]_pad  & ~n1116 ;
  assign n9403 = ~n9401 & ~n9402 ;
  assign n9404 = \ks1_col_reg[3]/NET0131  & ~n9403 ;
  assign n9405 = ~\ks1_col_reg[3]/NET0131  & n9403 ;
  assign n9406 = ~n9404 & ~n9405 ;
  assign n9407 = ~\ks1_key_reg_reg[67]/NET0131  & n1116 ;
  assign n9408 = ~\key_i[67]_pad  & ~n1116 ;
  assign n9409 = ~n9407 & ~n9408 ;
  assign n9410 = n9406 & ~n9409 ;
  assign n9411 = ~n9406 & n9409 ;
  assign n9412 = ~n9410 & ~n9411 ;
  assign n9413 = ~\ks1_key_reg_reg[35]/NET0131  & n1116 ;
  assign n9414 = ~\key_i[35]_pad  & ~n1116 ;
  assign n9415 = ~n9413 & ~n9414 ;
  assign n9416 = n9412 & ~n9415 ;
  assign n9417 = ~n9412 & n9415 ;
  assign n9418 = ~n9416 & ~n9417 ;
  assign n9419 = n929 & ~n9418 ;
  assign n9420 = \ks1_key_reg_reg[35]/NET0131  & ~n929 ;
  assign n9421 = ~n9419 & ~n9420 ;
  assign n9422 = ~\ks1_key_reg_reg[100]/NET0131  & n1116 ;
  assign n9423 = ~\key_i[100]_pad  & ~n1116 ;
  assign n9424 = ~n9422 & ~n9423 ;
  assign n9425 = \ks1_col_reg[4]/NET0131  & ~n9424 ;
  assign n9426 = ~\ks1_col_reg[4]/NET0131  & n9424 ;
  assign n9427 = ~n9425 & ~n9426 ;
  assign n9428 = ~\ks1_key_reg_reg[68]/NET0131  & n1116 ;
  assign n9429 = ~\key_i[68]_pad  & ~n1116 ;
  assign n9430 = ~n9428 & ~n9429 ;
  assign n9431 = n9427 & ~n9430 ;
  assign n9432 = ~n9427 & n9430 ;
  assign n9433 = ~n9431 & ~n9432 ;
  assign n9434 = ~\ks1_key_reg_reg[36]/NET0131  & n1116 ;
  assign n9435 = ~\key_i[36]_pad  & ~n1116 ;
  assign n9436 = ~n9434 & ~n9435 ;
  assign n9437 = n9433 & ~n9436 ;
  assign n9438 = ~n9433 & n9436 ;
  assign n9439 = ~n9437 & ~n9438 ;
  assign n9440 = n929 & ~n9439 ;
  assign n9441 = \ks1_key_reg_reg[36]/NET0131  & ~n929 ;
  assign n9442 = ~n9440 & ~n9441 ;
  assign n9443 = ~\ks1_key_reg_reg[101]/NET0131  & n1116 ;
  assign n9444 = ~\key_i[101]_pad  & ~n1116 ;
  assign n9445 = ~n9443 & ~n9444 ;
  assign n9446 = \ks1_col_reg[5]/NET0131  & ~n9445 ;
  assign n9447 = ~\ks1_col_reg[5]/NET0131  & n9445 ;
  assign n9448 = ~n9446 & ~n9447 ;
  assign n9449 = ~\ks1_key_reg_reg[69]/NET0131  & n1116 ;
  assign n9450 = ~\key_i[69]_pad  & ~n1116 ;
  assign n9451 = ~n9449 & ~n9450 ;
  assign n9452 = n9448 & ~n9451 ;
  assign n9453 = ~n9448 & n9451 ;
  assign n9454 = ~n9452 & ~n9453 ;
  assign n9455 = ~\ks1_key_reg_reg[37]/NET0131  & n1116 ;
  assign n9456 = ~\key_i[37]_pad  & ~n1116 ;
  assign n9457 = ~n9455 & ~n9456 ;
  assign n9458 = n9454 & ~n9457 ;
  assign n9459 = ~n9454 & n9457 ;
  assign n9460 = ~n9458 & ~n9459 ;
  assign n9461 = n929 & ~n9460 ;
  assign n9462 = \ks1_key_reg_reg[37]/NET0131  & ~n929 ;
  assign n9463 = ~n9461 & ~n9462 ;
  assign n9464 = ~\ks1_key_reg_reg[102]/NET0131  & n1116 ;
  assign n9465 = ~\key_i[102]_pad  & ~n1116 ;
  assign n9466 = ~n9464 & ~n9465 ;
  assign n9467 = \ks1_col_reg[6]/NET0131  & ~n9466 ;
  assign n9468 = ~\ks1_col_reg[6]/NET0131  & n9466 ;
  assign n9469 = ~n9467 & ~n9468 ;
  assign n9470 = ~\ks1_key_reg_reg[70]/NET0131  & n1116 ;
  assign n9471 = ~\key_i[70]_pad  & ~n1116 ;
  assign n9472 = ~n9470 & ~n9471 ;
  assign n9473 = n9469 & ~n9472 ;
  assign n9474 = ~n9469 & n9472 ;
  assign n9475 = ~n9473 & ~n9474 ;
  assign n9476 = ~\ks1_key_reg_reg[38]/NET0131  & n1116 ;
  assign n9477 = ~\key_i[38]_pad  & ~n1116 ;
  assign n9478 = ~n9476 & ~n9477 ;
  assign n9479 = n9475 & ~n9478 ;
  assign n9480 = ~n9475 & n9478 ;
  assign n9481 = ~n9479 & ~n9480 ;
  assign n9482 = n929 & ~n9481 ;
  assign n9483 = \ks1_key_reg_reg[38]/NET0131  & ~n929 ;
  assign n9484 = ~n9482 & ~n9483 ;
  assign n9485 = ~\ks1_key_reg_reg[103]/NET0131  & n1116 ;
  assign n9486 = ~\key_i[103]_pad  & ~n1116 ;
  assign n9487 = ~n9485 & ~n9486 ;
  assign n9488 = \ks1_col_reg[7]/NET0131  & ~n9487 ;
  assign n9489 = ~\ks1_col_reg[7]/NET0131  & n9487 ;
  assign n9490 = ~n9488 & ~n9489 ;
  assign n9491 = ~\ks1_key_reg_reg[71]/NET0131  & n1116 ;
  assign n9492 = ~\key_i[71]_pad  & ~n1116 ;
  assign n9493 = ~n9491 & ~n9492 ;
  assign n9494 = n9490 & ~n9493 ;
  assign n9495 = ~n9490 & n9493 ;
  assign n9496 = ~n9494 & ~n9495 ;
  assign n9497 = ~\ks1_key_reg_reg[39]/NET0131  & n1116 ;
  assign n9498 = ~\key_i[39]_pad  & ~n1116 ;
  assign n9499 = ~n9497 & ~n9498 ;
  assign n9500 = n9496 & ~n9499 ;
  assign n9501 = ~n9496 & n9499 ;
  assign n9502 = ~n9500 & ~n9501 ;
  assign n9503 = n929 & ~n9502 ;
  assign n9504 = \ks1_key_reg_reg[39]/NET0131  & ~n929 ;
  assign n9505 = ~n9503 & ~n9504 ;
  assign n9506 = \key_i[80]_pad  & ~n953 ;
  assign n9507 = \ks1_key_reg_reg[80]/NET0131  & n956 ;
  assign n9508 = ~n9506 & ~n9507 ;
  assign n9509 = ~n933 & ~n9508 ;
  assign n9511 = ~\key_i[80]_pad  & n951 ;
  assign n9510 = ~\ks1_key_reg_reg[80]/NET0131  & ~n951 ;
  assign n9512 = n933 & ~n9510 ;
  assign n9513 = ~n9511 & n9512 ;
  assign n9514 = ~n9509 & ~n9513 ;
  assign n9515 = ~\ks1_key_reg_reg[112]/NET0131  & n1116 ;
  assign n9516 = ~\key_i[112]_pad  & ~n1116 ;
  assign n9517 = ~n9515 & ~n9516 ;
  assign n9518 = \ks1_col_reg[16]/NET0131  & ~n9517 ;
  assign n9519 = ~\ks1_col_reg[16]/NET0131  & n9517 ;
  assign n9520 = ~n9518 & ~n9519 ;
  assign n9521 = n9514 & n9520 ;
  assign n9522 = ~n9514 & ~n9520 ;
  assign n9523 = ~n9521 & ~n9522 ;
  assign n9524 = ~\ks1_key_reg_reg[48]/NET0131  & n1116 ;
  assign n9525 = ~\key_i[48]_pad  & ~n1116 ;
  assign n9526 = ~n9524 & ~n9525 ;
  assign n9527 = n9523 & ~n9526 ;
  assign n9528 = ~n9523 & n9526 ;
  assign n9529 = ~n9527 & ~n9528 ;
  assign n9530 = n929 & ~n9529 ;
  assign n9531 = \ks1_key_reg_reg[48]/NET0131  & ~n929 ;
  assign n9532 = ~n9530 & ~n9531 ;
  assign n9533 = \key_i[81]_pad  & ~n953 ;
  assign n9534 = \ks1_key_reg_reg[81]/NET0131  & n956 ;
  assign n9535 = ~n9533 & ~n9534 ;
  assign n9536 = ~n933 & ~n9535 ;
  assign n9538 = ~\key_i[81]_pad  & n951 ;
  assign n9537 = ~\ks1_key_reg_reg[81]/NET0131  & ~n951 ;
  assign n9539 = n933 & ~n9537 ;
  assign n9540 = ~n9538 & n9539 ;
  assign n9541 = ~n9536 & ~n9540 ;
  assign n9542 = ~\ks1_key_reg_reg[113]/NET0131  & n1116 ;
  assign n9543 = ~\key_i[113]_pad  & ~n1116 ;
  assign n9544 = ~n9542 & ~n9543 ;
  assign n9545 = \ks1_col_reg[17]/NET0131  & ~n9544 ;
  assign n9546 = ~\ks1_col_reg[17]/NET0131  & n9544 ;
  assign n9547 = ~n9545 & ~n9546 ;
  assign n9548 = n9541 & n9547 ;
  assign n9549 = ~n9541 & ~n9547 ;
  assign n9550 = ~n9548 & ~n9549 ;
  assign n9551 = ~\ks1_key_reg_reg[49]/NET0131  & n1116 ;
  assign n9552 = ~\key_i[49]_pad  & ~n1116 ;
  assign n9553 = ~n9551 & ~n9552 ;
  assign n9554 = n9550 & ~n9553 ;
  assign n9555 = ~n9550 & n9553 ;
  assign n9556 = ~n9554 & ~n9555 ;
  assign n9557 = n929 & ~n9556 ;
  assign n9558 = \ks1_key_reg_reg[49]/NET0131  & ~n929 ;
  assign n9559 = ~n9557 & ~n9558 ;
  assign n9560 = \key_i[82]_pad  & ~n953 ;
  assign n9561 = \ks1_key_reg_reg[82]/NET0131  & n956 ;
  assign n9562 = ~n9560 & ~n9561 ;
  assign n9563 = ~n933 & ~n9562 ;
  assign n9565 = ~\key_i[82]_pad  & n951 ;
  assign n9564 = ~\ks1_key_reg_reg[82]/NET0131  & ~n951 ;
  assign n9566 = n933 & ~n9564 ;
  assign n9567 = ~n9565 & n9566 ;
  assign n9568 = ~n9563 & ~n9567 ;
  assign n9569 = ~\ks1_key_reg_reg[114]/NET0131  & n1116 ;
  assign n9570 = ~\key_i[114]_pad  & ~n1116 ;
  assign n9571 = ~n9569 & ~n9570 ;
  assign n9572 = \ks1_col_reg[18]/NET0131  & ~n9571 ;
  assign n9573 = ~\ks1_col_reg[18]/NET0131  & n9571 ;
  assign n9574 = ~n9572 & ~n9573 ;
  assign n9575 = n9568 & n9574 ;
  assign n9576 = ~n9568 & ~n9574 ;
  assign n9577 = ~n9575 & ~n9576 ;
  assign n9578 = ~\ks1_key_reg_reg[50]/NET0131  & n1116 ;
  assign n9579 = ~\key_i[50]_pad  & ~n1116 ;
  assign n9580 = ~n9578 & ~n9579 ;
  assign n9581 = n9577 & ~n9580 ;
  assign n9582 = ~n9577 & n9580 ;
  assign n9583 = ~n9581 & ~n9582 ;
  assign n9584 = n929 & ~n9583 ;
  assign n9585 = \ks1_key_reg_reg[50]/NET0131  & ~n929 ;
  assign n9586 = ~n9584 & ~n9585 ;
  assign n9587 = \key_i[83]_pad  & ~n953 ;
  assign n9588 = \ks1_key_reg_reg[83]/NET0131  & n956 ;
  assign n9589 = ~n9587 & ~n9588 ;
  assign n9590 = ~n933 & ~n9589 ;
  assign n9592 = ~\key_i[83]_pad  & n951 ;
  assign n9591 = ~\ks1_key_reg_reg[83]/NET0131  & ~n951 ;
  assign n9593 = n933 & ~n9591 ;
  assign n9594 = ~n9592 & n9593 ;
  assign n9595 = ~n9590 & ~n9594 ;
  assign n9596 = ~\ks1_key_reg_reg[115]/NET0131  & n1116 ;
  assign n9597 = ~\key_i[115]_pad  & ~n1116 ;
  assign n9598 = ~n9596 & ~n9597 ;
  assign n9599 = \ks1_col_reg[19]/NET0131  & ~n9598 ;
  assign n9600 = ~\ks1_col_reg[19]/NET0131  & n9598 ;
  assign n9601 = ~n9599 & ~n9600 ;
  assign n9602 = n9595 & n9601 ;
  assign n9603 = ~n9595 & ~n9601 ;
  assign n9604 = ~n9602 & ~n9603 ;
  assign n9605 = ~\ks1_key_reg_reg[51]/NET0131  & n1116 ;
  assign n9606 = ~\key_i[51]_pad  & ~n1116 ;
  assign n9607 = ~n9605 & ~n9606 ;
  assign n9608 = n9604 & ~n9607 ;
  assign n9609 = ~n9604 & n9607 ;
  assign n9610 = ~n9608 & ~n9609 ;
  assign n9611 = n929 & ~n9610 ;
  assign n9612 = \ks1_key_reg_reg[51]/NET0131  & ~n929 ;
  assign n9613 = ~n9611 & ~n9612 ;
  assign n9614 = \key_i[84]_pad  & ~n953 ;
  assign n9615 = \ks1_key_reg_reg[84]/NET0131  & n956 ;
  assign n9616 = ~n9614 & ~n9615 ;
  assign n9617 = ~n933 & ~n9616 ;
  assign n9619 = ~\key_i[84]_pad  & n951 ;
  assign n9618 = ~\ks1_key_reg_reg[84]/NET0131  & ~n951 ;
  assign n9620 = n933 & ~n9618 ;
  assign n9621 = ~n9619 & n9620 ;
  assign n9622 = ~n9617 & ~n9621 ;
  assign n9623 = ~\ks1_key_reg_reg[116]/NET0131  & n1116 ;
  assign n9624 = ~\key_i[116]_pad  & ~n1116 ;
  assign n9625 = ~n9623 & ~n9624 ;
  assign n9626 = \ks1_col_reg[20]/NET0131  & ~n9625 ;
  assign n9627 = ~\ks1_col_reg[20]/NET0131  & n9625 ;
  assign n9628 = ~n9626 & ~n9627 ;
  assign n9629 = n9622 & n9628 ;
  assign n9630 = ~n9622 & ~n9628 ;
  assign n9631 = ~n9629 & ~n9630 ;
  assign n9632 = ~\ks1_key_reg_reg[52]/NET0131  & n1116 ;
  assign n9633 = ~\key_i[52]_pad  & ~n1116 ;
  assign n9634 = ~n9632 & ~n9633 ;
  assign n9635 = n9631 & ~n9634 ;
  assign n9636 = ~n9631 & n9634 ;
  assign n9637 = ~n9635 & ~n9636 ;
  assign n9638 = n929 & ~n9637 ;
  assign n9639 = \ks1_key_reg_reg[52]/NET0131  & ~n929 ;
  assign n9640 = ~n9638 & ~n9639 ;
  assign n9641 = \key_i[85]_pad  & ~n953 ;
  assign n9642 = \ks1_key_reg_reg[85]/NET0131  & n956 ;
  assign n9643 = ~n9641 & ~n9642 ;
  assign n9644 = ~n933 & ~n9643 ;
  assign n9646 = ~\key_i[85]_pad  & n951 ;
  assign n9645 = ~\ks1_key_reg_reg[85]/NET0131  & ~n951 ;
  assign n9647 = n933 & ~n9645 ;
  assign n9648 = ~n9646 & n9647 ;
  assign n9649 = ~n9644 & ~n9648 ;
  assign n9650 = ~\ks1_key_reg_reg[117]/NET0131  & n1116 ;
  assign n9651 = ~\key_i[117]_pad  & ~n1116 ;
  assign n9652 = ~n9650 & ~n9651 ;
  assign n9653 = \ks1_col_reg[21]/NET0131  & ~n9652 ;
  assign n9654 = ~\ks1_col_reg[21]/NET0131  & n9652 ;
  assign n9655 = ~n9653 & ~n9654 ;
  assign n9656 = n9649 & n9655 ;
  assign n9657 = ~n9649 & ~n9655 ;
  assign n9658 = ~n9656 & ~n9657 ;
  assign n9659 = ~\ks1_key_reg_reg[53]/NET0131  & n1116 ;
  assign n9660 = ~\key_i[53]_pad  & ~n1116 ;
  assign n9661 = ~n9659 & ~n9660 ;
  assign n9662 = n9658 & ~n9661 ;
  assign n9663 = ~n9658 & n9661 ;
  assign n9664 = ~n9662 & ~n9663 ;
  assign n9665 = n929 & ~n9664 ;
  assign n9666 = \ks1_key_reg_reg[53]/NET0131  & ~n929 ;
  assign n9667 = ~n9665 & ~n9666 ;
  assign n9668 = \key_i[86]_pad  & ~n953 ;
  assign n9669 = \ks1_key_reg_reg[86]/NET0131  & n956 ;
  assign n9670 = ~n9668 & ~n9669 ;
  assign n9671 = ~n933 & ~n9670 ;
  assign n9673 = ~\key_i[86]_pad  & n951 ;
  assign n9672 = ~\ks1_key_reg_reg[86]/NET0131  & ~n951 ;
  assign n9674 = n933 & ~n9672 ;
  assign n9675 = ~n9673 & n9674 ;
  assign n9676 = ~n9671 & ~n9675 ;
  assign n9677 = ~\ks1_key_reg_reg[118]/NET0131  & n1116 ;
  assign n9678 = ~\key_i[118]_pad  & ~n1116 ;
  assign n9679 = ~n9677 & ~n9678 ;
  assign n9680 = \ks1_col_reg[22]/NET0131  & ~n9679 ;
  assign n9681 = ~\ks1_col_reg[22]/NET0131  & n9679 ;
  assign n9682 = ~n9680 & ~n9681 ;
  assign n9683 = n9676 & n9682 ;
  assign n9684 = ~n9676 & ~n9682 ;
  assign n9685 = ~n9683 & ~n9684 ;
  assign n9686 = ~\ks1_key_reg_reg[54]/NET0131  & n1116 ;
  assign n9687 = ~\key_i[54]_pad  & ~n1116 ;
  assign n9688 = ~n9686 & ~n9687 ;
  assign n9689 = n9685 & ~n9688 ;
  assign n9690 = ~n9685 & n9688 ;
  assign n9691 = ~n9689 & ~n9690 ;
  assign n9692 = n929 & ~n9691 ;
  assign n9693 = \ks1_key_reg_reg[54]/NET0131  & ~n929 ;
  assign n9694 = ~n9692 & ~n9693 ;
  assign n9695 = \key_i[87]_pad  & ~n953 ;
  assign n9696 = \ks1_key_reg_reg[87]/NET0131  & n956 ;
  assign n9697 = ~n9695 & ~n9696 ;
  assign n9698 = ~n933 & ~n9697 ;
  assign n9700 = ~\key_i[87]_pad  & n951 ;
  assign n9699 = ~\ks1_key_reg_reg[87]/NET0131  & ~n951 ;
  assign n9701 = n933 & ~n9699 ;
  assign n9702 = ~n9700 & n9701 ;
  assign n9703 = ~n9698 & ~n9702 ;
  assign n9704 = ~\ks1_key_reg_reg[119]/NET0131  & n1116 ;
  assign n9705 = ~\key_i[119]_pad  & ~n1116 ;
  assign n9706 = ~n9704 & ~n9705 ;
  assign n9707 = \ks1_col_reg[23]/NET0131  & ~n9706 ;
  assign n9708 = ~\ks1_col_reg[23]/NET0131  & n9706 ;
  assign n9709 = ~n9707 & ~n9708 ;
  assign n9710 = n9703 & n9709 ;
  assign n9711 = ~n9703 & ~n9709 ;
  assign n9712 = ~n9710 & ~n9711 ;
  assign n9713 = ~\ks1_key_reg_reg[55]/NET0131  & n1116 ;
  assign n9714 = ~\key_i[55]_pad  & ~n1116 ;
  assign n9715 = ~n9713 & ~n9714 ;
  assign n9716 = n9712 & ~n9715 ;
  assign n9717 = ~n9712 & n9715 ;
  assign n9718 = ~n9716 & ~n9717 ;
  assign n9719 = n929 & ~n9718 ;
  assign n9720 = \ks1_key_reg_reg[55]/NET0131  & ~n929 ;
  assign n9721 = ~n9719 & ~n9720 ;
  assign n9722 = n1507 & n9418 ;
  assign n9723 = ~n1507 & ~n9418 ;
  assign n9724 = ~n9722 & ~n9723 ;
  assign n9725 = n1151 & n9439 ;
  assign n9726 = ~n1151 & ~n9439 ;
  assign n9727 = ~n9725 & ~n9726 ;
  assign n9728 = n1881 & n9460 ;
  assign n9729 = ~n1881 & ~n9460 ;
  assign n9730 = ~n9728 & ~n9729 ;
  assign n9731 = n1406 & n9481 ;
  assign n9732 = ~n1406 & ~n9481 ;
  assign n9733 = ~n9731 & ~n9732 ;
  assign n9734 = n2074 & n9502 ;
  assign n9735 = ~n2074 & ~n9502 ;
  assign n9736 = ~n9734 & ~n9735 ;
  assign n9737 = n1791 & n9343 ;
  assign n9738 = ~n1791 & ~n9343 ;
  assign n9739 = ~n9737 & ~n9738 ;
  assign n9740 = n1761 & n9529 ;
  assign n9741 = ~n1761 & ~n9529 ;
  assign n9742 = ~n9740 & ~n9741 ;
  assign n9743 = n1646 & n9556 ;
  assign n9744 = ~n1646 & ~n9556 ;
  assign n9745 = ~n9743 & ~n9744 ;
  assign n9746 = n2029 & n9583 ;
  assign n9747 = ~n2029 & ~n9583 ;
  assign n9748 = ~n9746 & ~n9747 ;
  assign n9749 = n1517 & n9610 ;
  assign n9750 = ~n1517 & ~n9610 ;
  assign n9751 = ~n9749 & ~n9750 ;
  assign n9752 = n1666 & n9370 ;
  assign n9753 = ~n1666 & ~n9370 ;
  assign n9754 = ~n9752 & ~n9753 ;
  assign n9755 = n1295 & n9637 ;
  assign n9756 = ~n1295 & ~n9637 ;
  assign n9757 = ~n9755 & ~n9756 ;
  assign n9758 = n1891 & n9664 ;
  assign n9759 = ~n1891 & ~n9664 ;
  assign n9760 = ~n9758 & ~n9759 ;
  assign n9761 = n1410 & n9691 ;
  assign n9762 = ~n1410 & ~n9691 ;
  assign n9763 = ~n9761 & ~n9762 ;
  assign n9764 = n2064 & n9718 ;
  assign n9765 = ~n2064 & ~n9718 ;
  assign n9766 = ~n9764 & ~n9765 ;
  assign n9767 = n2049 & n9397 ;
  assign n9768 = ~n2049 & ~n9397 ;
  assign n9769 = ~n9767 & ~n9768 ;
  assign n9770 = n3640 & ~n9238 ;
  assign n9771 = ~\mix1_data_o_reg_reg[0]/NET0131  & ~n3640 ;
  assign n9772 = ~n9770 & ~n9771 ;
  assign n9773 = n3640 & n9121 ;
  assign n9774 = \mix1_data_o_reg_reg[16]/NET0131  & ~n3640 ;
  assign n9775 = ~n9773 & ~n9774 ;
  assign n9776 = n3640 & n9133 ;
  assign n9777 = \mix1_data_o_reg_reg[24]/NET0131  & ~n3640 ;
  assign n9778 = ~n9776 & ~n9777 ;
  assign n9779 = n3640 & ~n9111 ;
  assign n9780 = \mix1_data_o_reg_reg[8]/NET0131  & ~n3640 ;
  assign n9781 = ~n9779 & ~n9780 ;
  assign n9782 = ~n971 & ~n1274 ;
  assign n9783 = \addroundkey_round_reg[0]/NET0131  & ~n967 ;
  assign n9784 = ~n4977 & ~n9783 ;
  assign n9785 = \addroundkey_round_reg[3]/NET0131  & ~\ks1_ready_o_reg/NET0131  ;
  assign n9786 = ~n4962 & ~n9785 ;
  assign n9787 = ~\addroundkey_start_i_reg/NET0131  & ~n9786 ;
  assign n9788 = ~n4965 & ~n9787 ;
  assign n9789 = \addroundkey_round_reg[1]/NET0131  & ~\ks1_ready_o_reg/NET0131  ;
  assign n9790 = ~n4970 & ~n9789 ;
  assign n9791 = ~\addroundkey_start_i_reg/NET0131  & ~n9790 ;
  assign n9792 = ~n4973 & ~n9791 ;
  assign n9793 = \addroundkey_round_reg[2]/NET0131  & ~\ks1_ready_o_reg/NET0131  ;
  assign n9794 = ~n4982 & ~n9793 ;
  assign n9795 = ~\addroundkey_start_i_reg/NET0131  & ~n9794 ;
  assign n9796 = ~n4985 & ~n9795 ;
  assign n9797 = ~n933 & ~n5053 ;
  assign n9802 = ~n5025 & ~n5027 ;
  assign n9811 = \round_reg[0]/NET0131  & \round_reg[1]/NET0131  ;
  assign n9812 = \round_reg[2]/NET0131  & n9811 ;
  assign n9813 = \round_reg[3]/NET0131  & ~n9812 ;
  assign n9814 = ~\round_reg[3]/NET0131  & n9812 ;
  assign n9815 = ~n9813 & ~n9814 ;
  assign n9816 = ~n9802 & n9815 ;
  assign n9803 = n930 & n5028 ;
  assign n9804 = ~\round_reg[2]/NET0131  & n9803 ;
  assign n9805 = \round_reg[3]/NET0131  & ~n9804 ;
  assign n9806 = \sub1_ready_o_reg/NET0131  & n1260 ;
  assign n9807 = ~n9805 & ~n9806 ;
  assign n9808 = n9802 & n9807 ;
  assign n9809 = \addroundkey_ready_o_reg/NET0131  & ~n1261 ;
  assign n9810 = \state_reg/NET0131  & ~n9809 ;
  assign n9817 = ~n9808 & n9810 ;
  assign n9818 = ~n9816 & n9817 ;
  assign n9798 = ~load_i_pad & ~\state_reg/NET0131  ;
  assign n9799 = \round_reg[3]/NET0131  & n9798 ;
  assign n9800 = load_i_pad & ~\state_reg/NET0131  ;
  assign n9801 = decrypt_i_pad & n9800 ;
  assign n9819 = ~n9799 & ~n9801 ;
  assign n9820 = ~n9818 & n9819 ;
  assign n9822 = ~n930 & ~n9811 ;
  assign n9823 = ~\round_reg[0]/NET0131  & ~n5028 ;
  assign n9824 = n9802 & ~n9823 ;
  assign n9826 = ~n9822 & ~n9824 ;
  assign n9825 = n9822 & n9824 ;
  assign n9827 = n9810 & ~n9825 ;
  assign n9828 = ~n9826 & n9827 ;
  assign n9821 = \round_reg[1]/NET0131  & n9798 ;
  assign n9829 = ~n9801 & ~n9821 ;
  assign n9830 = ~n9828 & n9829 ;
  assign n9831 = ~n3629 & ~n3635 ;
  assign n9832 = ~n3630 & ~n3635 ;
  assign n9833 = \first_round_reg_reg/NET0131  & ~\state_reg/NET0131  ;
  assign n9834 = ~\first_round_reg_reg/NET0131  & ~n5027 ;
  assign n9835 = ~n5028 & n9834 ;
  assign n9836 = n3625 & ~n9835 ;
  assign n9837 = ~n5025 & ~n9836 ;
  assign n9838 = n9810 & ~n9837 ;
  assign n9839 = ~n9833 & ~n9838 ;
  assign n9840 = ~\sub1_state_reg[0]/NET0131  & ~n1256 ;
  assign n9841 = ~\sub1_state_reg[0]/NET0131  & ~n1266 ;
  assign n9842 = n1267 & ~n9841 ;
  assign n9843 = ~n9840 & ~n9842 ;
  assign n9844 = \round_reg[2]/NET0131  & n9798 ;
  assign n9845 = \round_reg[2]/NET0131  & ~n9803 ;
  assign n9846 = ~n5027 & ~n9804 ;
  assign n9847 = ~n9845 & n9846 ;
  assign n9848 = ~\round_reg[2]/NET0131  & ~n9811 ;
  assign n9849 = ~n9812 & ~n9848 ;
  assign n9850 = n5027 & ~n9849 ;
  assign n9851 = n3625 & ~n9850 ;
  assign n9852 = ~n9847 & n9851 ;
  assign n9853 = n9810 & n9852 ;
  assign n9854 = ~n9844 & ~n9853 ;
  assign n9855 = ~n1201 & ~n2491 ;
  assign n9856 = \sub1_state_reg[4]/NET0131  & n1201 ;
  assign n9857 = ~n9855 & ~n9856 ;
  assign n9858 = ~\sub1_state_reg[2]/NET0131  & ~n1165 ;
  assign n9859 = ~n1200 & ~n9858 ;
  assign n9860 = ~n5028 & n9802 ;
  assign n9861 = n9810 & ~n9860 ;
  assign n9862 = ~\round_reg[0]/NET0131  & ~n9861 ;
  assign n9863 = n9810 & n9860 ;
  assign n9864 = \round_reg[0]/NET0131  & ~n9798 ;
  assign n9865 = ~n9863 & n9864 ;
  assign n9866 = ~n9862 & ~n9865 ;
  assign n9867 = ~n9800 & ~n9810 ;
  assign n9868 = \addroundkey_ready_o_reg/NET0131  & n1262 ;
  assign n9869 = \sub1_state_reg[3]/NET0131  & ~n1200 ;
  assign n9870 = ~n1206 & ~n9869 ;
  assign n9871 = \mix1_data_o_reg_reg[89]/NET0131  & ~n3640 ;
  assign n9872 = \mix1_data_reg_reg[89]/NET0131  & n3640 ;
  assign n9873 = ~n9871 & ~n9872 ;
  assign n9874 = \mix1_data_o_reg_reg[99]/NET0131  & ~n3640 ;
  assign n9875 = \mix1_data_reg_reg[99]/NET0131  & n3640 ;
  assign n9876 = ~n9874 & ~n9875 ;
  assign n9877 = \mix1_data_o_reg_reg[37]/NET0131  & ~n3640 ;
  assign n9878 = \mix1_data_reg_reg[37]/NET0131  & n3640 ;
  assign n9879 = ~n9877 & ~n9878 ;
  assign n9880 = \mix1_data_o_reg_reg[110]/NET0131  & ~n3640 ;
  assign n9881 = \mix1_data_reg_reg[110]/NET0131  & n3640 ;
  assign n9882 = ~n9880 & ~n9881 ;
  assign n9883 = \mix1_data_o_reg_reg[40]/NET0131  & ~n3640 ;
  assign n9884 = \mix1_data_reg_reg[40]/NET0131  & n3640 ;
  assign n9885 = ~n9883 & ~n9884 ;
  assign n9886 = \mix1_data_o_reg_reg[34]/NET0131  & ~n3640 ;
  assign n9887 = \mix1_data_reg_reg[34]/NET0131  & n3640 ;
  assign n9888 = ~n9886 & ~n9887 ;
  assign n9889 = \mix1_data_o_reg_reg[48]/NET0131  & ~n3640 ;
  assign n9890 = \mix1_data_reg_reg[48]/NET0131  & n3640 ;
  assign n9891 = ~n9889 & ~n9890 ;
  assign n9892 = \mix1_data_o_reg_reg[105]/NET0131  & ~n3640 ;
  assign n9893 = \mix1_data_reg_reg[105]/NET0131  & n3640 ;
  assign n9894 = ~n9892 & ~n9893 ;
  assign n9895 = \mix1_data_o_reg_reg[43]/NET0131  & ~n3640 ;
  assign n9896 = \mix1_data_reg_reg[43]/NET0131  & n3640 ;
  assign n9897 = ~n9895 & ~n9896 ;
  assign n9898 = \mix1_data_o_reg_reg[95]/NET0131  & ~n3640 ;
  assign n9899 = \mix1_data_reg_reg[95]/NET0131  & n3640 ;
  assign n9900 = ~n9898 & ~n9899 ;
  assign n9901 = \mix1_data_o_reg_reg[93]/NET0131  & ~n3640 ;
  assign n9902 = \mix1_data_reg_reg[93]/NET0131  & n3640 ;
  assign n9903 = ~n9901 & ~n9902 ;
  assign n9904 = \mix1_data_o_reg_reg[97]/NET0131  & ~n3640 ;
  assign n9905 = \mix1_data_reg_reg[97]/NET0131  & n3640 ;
  assign n9906 = ~n9904 & ~n9905 ;
  assign n9907 = \mix1_data_o_reg_reg[35]/NET0131  & ~n3640 ;
  assign n9908 = \mix1_data_reg_reg[35]/NET0131  & n3640 ;
  assign n9909 = ~n9907 & ~n9908 ;
  assign n9910 = \mix1_data_o_reg_reg[106]/NET0131  & ~n3640 ;
  assign n9911 = \mix1_data_reg_reg[106]/NET0131  & n3640 ;
  assign n9912 = ~n9910 & ~n9911 ;
  assign n9913 = \mix1_data_o_reg_reg[107]/NET0131  & ~n3640 ;
  assign n9914 = \mix1_data_reg_reg[107]/NET0131  & n3640 ;
  assign n9915 = ~n9913 & ~n9914 ;
  assign n9916 = \mix1_data_o_reg_reg[108]/NET0131  & ~n3640 ;
  assign n9917 = \mix1_data_reg_reg[108]/NET0131  & n3640 ;
  assign n9918 = ~n9916 & ~n9917 ;
  assign n9919 = \mix1_data_o_reg_reg[91]/NET0131  & ~n3640 ;
  assign n9920 = \mix1_data_reg_reg[91]/NET0131  & n3640 ;
  assign n9921 = ~n9919 & ~n9920 ;
  assign n9922 = \mix1_data_o_reg_reg[111]/NET0131  & ~n3640 ;
  assign n9923 = \mix1_data_reg_reg[111]/NET0131  & n3640 ;
  assign n9924 = ~n9922 & ~n9923 ;
  assign n9925 = \mix1_data_o_reg_reg[33]/NET0131  & ~n3640 ;
  assign n9926 = \mix1_data_reg_reg[33]/NET0131  & n3640 ;
  assign n9927 = ~n9925 & ~n9926 ;
  assign n9928 = \mix1_data_o_reg_reg[114]/NET0131  & ~n3640 ;
  assign n9929 = \mix1_data_reg_reg[114]/NET0131  & n3640 ;
  assign n9930 = ~n9928 & ~n9929 ;
  assign n9931 = \mix1_data_o_reg_reg[115]/NET0131  & ~n3640 ;
  assign n9932 = \mix1_data_reg_reg[115]/NET0131  & n3640 ;
  assign n9933 = ~n9931 & ~n9932 ;
  assign n9934 = \mix1_data_o_reg_reg[116]/NET0131  & ~n3640 ;
  assign n9935 = \mix1_data_reg_reg[116]/NET0131  & n3640 ;
  assign n9936 = ~n9934 & ~n9935 ;
  assign n9937 = \mix1_data_o_reg_reg[118]/NET0131  & ~n3640 ;
  assign n9938 = \mix1_data_reg_reg[118]/NET0131  & n3640 ;
  assign n9939 = ~n9937 & ~n9938 ;
  assign n9940 = \mix1_data_o_reg_reg[120]/NET0131  & ~n3640 ;
  assign n9941 = \mix1_data_reg_reg[120]/NET0131  & n3640 ;
  assign n9942 = ~n9940 & ~n9941 ;
  assign n9943 = \mix1_data_o_reg_reg[112]/NET0131  & ~n3640 ;
  assign n9944 = \mix1_data_reg_reg[112]/NET0131  & n3640 ;
  assign n9945 = ~n9943 & ~n9944 ;
  assign n9946 = \mix1_data_o_reg_reg[124]/NET0131  & ~n3640 ;
  assign n9947 = \mix1_data_reg_reg[124]/NET0131  & n3640 ;
  assign n9948 = ~n9946 & ~n9947 ;
  assign n9949 = \mix1_data_o_reg_reg[83]/NET0131  & ~n3640 ;
  assign n9950 = \mix1_data_reg_reg[83]/NET0131  & n3640 ;
  assign n9951 = ~n9949 & ~n9950 ;
  assign n9952 = \mix1_data_o_reg_reg[81]/NET0131  & ~n3640 ;
  assign n9953 = \mix1_data_reg_reg[81]/NET0131  & n3640 ;
  assign n9954 = ~n9952 & ~n9953 ;
  assign n9955 = \mix1_data_o_reg_reg[42]/NET0131  & ~n3640 ;
  assign n9956 = \mix1_data_reg_reg[42]/NET0131  & n3640 ;
  assign n9957 = ~n9955 & ~n9956 ;
  assign n9958 = \mix1_data_o_reg_reg[32]/NET0131  & ~n3640 ;
  assign n9959 = \mix1_data_reg_reg[32]/NET0131  & n3640 ;
  assign n9960 = ~n9958 & ~n9959 ;
  assign n9961 = \mix1_data_o_reg_reg[113]/NET0131  & ~n3640 ;
  assign n9962 = \mix1_data_reg_reg[113]/NET0131  & n3640 ;
  assign n9963 = ~n9961 & ~n9962 ;
  assign n9964 = \mix1_data_o_reg_reg[38]/NET0131  & ~n3640 ;
  assign n9965 = \mix1_data_reg_reg[38]/NET0131  & n3640 ;
  assign n9966 = ~n9964 & ~n9965 ;
  assign n9967 = \mix1_data_o_reg_reg[41]/NET0131  & ~n3640 ;
  assign n9968 = \mix1_data_reg_reg[41]/NET0131  & n3640 ;
  assign n9969 = ~n9967 & ~n9968 ;
  assign n9970 = \mix1_data_o_reg_reg[45]/NET0131  & ~n3640 ;
  assign n9971 = \mix1_data_reg_reg[45]/NET0131  & n3640 ;
  assign n9972 = ~n9970 & ~n9971 ;
  assign n9973 = \mix1_data_o_reg_reg[49]/NET0131  & ~n3640 ;
  assign n9974 = \mix1_data_reg_reg[49]/NET0131  & n3640 ;
  assign n9975 = ~n9973 & ~n9974 ;
  assign n9976 = \mix1_data_o_reg_reg[52]/NET0131  & ~n3640 ;
  assign n9977 = \mix1_data_reg_reg[52]/NET0131  & n3640 ;
  assign n9978 = ~n9976 & ~n9977 ;
  assign n9979 = \mix1_data_o_reg_reg[56]/NET0131  & ~n3640 ;
  assign n9980 = \mix1_data_reg_reg[56]/NET0131  & n3640 ;
  assign n9981 = ~n9979 & ~n9980 ;
  assign n9982 = \mix1_data_o_reg_reg[61]/NET0131  & ~n3640 ;
  assign n9983 = \mix1_data_reg_reg[61]/NET0131  & n3640 ;
  assign n9984 = ~n9982 & ~n9983 ;
  assign n9985 = \mix1_data_o_reg_reg[62]/NET0131  & ~n3640 ;
  assign n9986 = \mix1_data_reg_reg[62]/NET0131  & n3640 ;
  assign n9987 = ~n9985 & ~n9986 ;
  assign n9988 = \mix1_data_o_reg_reg[64]/NET0131  & ~n3640 ;
  assign n9989 = \mix1_data_reg_reg[64]/NET0131  & n3640 ;
  assign n9990 = ~n9988 & ~n9989 ;
  assign n9991 = \mix1_data_o_reg_reg[125]/NET0131  & ~n3640 ;
  assign n9992 = \mix1_data_reg_reg[125]/NET0131  & n3640 ;
  assign n9993 = ~n9991 & ~n9992 ;
  assign n9994 = \mix1_data_o_reg_reg[71]/NET0131  & ~n3640 ;
  assign n9995 = \mix1_data_reg_reg[71]/NET0131  & n3640 ;
  assign n9996 = ~n9994 & ~n9995 ;
  assign n9997 = \mix1_data_o_reg_reg[75]/NET0131  & ~n3640 ;
  assign n9998 = \mix1_data_reg_reg[75]/NET0131  & n3640 ;
  assign n9999 = ~n9997 & ~n9998 ;
  assign n10000 = \mix1_data_o_reg_reg[77]/NET0131  & ~n3640 ;
  assign n10001 = \mix1_data_reg_reg[77]/NET0131  & n3640 ;
  assign n10002 = ~n10000 & ~n10001 ;
  assign n10003 = \mix1_data_o_reg_reg[80]/NET0131  & ~n3640 ;
  assign n10004 = \mix1_data_reg_reg[80]/NET0131  & n3640 ;
  assign n10005 = ~n10003 & ~n10004 ;
  assign n10006 = \mix1_data_o_reg_reg[98]/NET0131  & ~n3640 ;
  assign n10007 = \mix1_data_reg_reg[98]/NET0131  & n3640 ;
  assign n10008 = ~n10006 & ~n10007 ;
  assign n10009 = \mix1_data_o_reg_reg[84]/NET0131  & ~n3640 ;
  assign n10010 = \mix1_data_reg_reg[84]/NET0131  & n3640 ;
  assign n10011 = ~n10009 & ~n10010 ;
  assign n10012 = \mix1_data_o_reg_reg[90]/NET0131  & ~n3640 ;
  assign n10013 = \mix1_data_reg_reg[90]/NET0131  & n3640 ;
  assign n10014 = ~n10012 & ~n10013 ;
  assign n10015 = \mix1_data_o_reg_reg[92]/NET0131  & ~n3640 ;
  assign n10016 = \mix1_data_reg_reg[92]/NET0131  & n3640 ;
  assign n10017 = ~n10015 & ~n10016 ;
  assign n10018 = \mix1_data_o_reg_reg[94]/NET0131  & ~n3640 ;
  assign n10019 = \mix1_data_reg_reg[94]/NET0131  & n3640 ;
  assign n10020 = ~n10018 & ~n10019 ;
  assign n10021 = \mix1_data_o_reg_reg[76]/NET0131  & ~n3640 ;
  assign n10022 = \mix1_data_reg_reg[76]/NET0131  & n3640 ;
  assign n10023 = ~n10021 & ~n10022 ;
  assign n10024 = \mix1_data_o_reg_reg[127]/NET0131  & ~n3640 ;
  assign n10025 = \mix1_data_reg_reg[127]/NET0131  & n3640 ;
  assign n10026 = ~n10024 & ~n10025 ;
  assign n10027 = \mix1_data_o_reg_reg[109]/NET0131  & ~n3640 ;
  assign n10028 = \mix1_data_reg_reg[109]/NET0131  & n3640 ;
  assign n10029 = ~n10027 & ~n10028 ;
  assign n10030 = \mix1_data_o_reg_reg[78]/NET0131  & ~n3640 ;
  assign n10031 = \mix1_data_reg_reg[78]/NET0131  & n3640 ;
  assign n10032 = ~n10030 & ~n10031 ;
  assign n10033 = \mix1_data_o_reg_reg[72]/NET0131  & ~n3640 ;
  assign n10034 = \mix1_data_reg_reg[72]/NET0131  & n3640 ;
  assign n10035 = ~n10033 & ~n10034 ;
  assign n10036 = \mix1_data_o_reg_reg[50]/NET0131  & ~n3640 ;
  assign n10037 = \mix1_data_reg_reg[50]/NET0131  & n3640 ;
  assign n10038 = ~n10036 & ~n10037 ;
  assign n10039 = \mix1_data_o_reg_reg[87]/NET0131  & ~n3640 ;
  assign n10040 = \mix1_data_reg_reg[87]/NET0131  & n3640 ;
  assign n10041 = ~n10039 & ~n10040 ;
  assign n10042 = \mix1_data_o_reg_reg[123]/NET0131  & ~n3640 ;
  assign n10043 = \mix1_data_reg_reg[123]/NET0131  & n3640 ;
  assign n10044 = ~n10042 & ~n10043 ;
  assign n10045 = \mix1_data_o_reg_reg[70]/NET0131  & ~n3640 ;
  assign n10046 = \mix1_data_reg_reg[70]/NET0131  & n3640 ;
  assign n10047 = ~n10045 & ~n10046 ;
  assign n10048 = \mix1_data_o_reg_reg[39]/NET0131  & ~n3640 ;
  assign n10049 = \mix1_data_reg_reg[39]/NET0131  & n3640 ;
  assign n10050 = ~n10048 & ~n10049 ;
  assign n10051 = \mix1_data_o_reg_reg[122]/NET0131  & ~n3640 ;
  assign n10052 = \mix1_data_reg_reg[122]/NET0131  & n3640 ;
  assign n10053 = ~n10051 & ~n10052 ;
  assign n10054 = \mix1_data_o_reg_reg[121]/NET0131  & ~n3640 ;
  assign n10055 = \mix1_data_reg_reg[121]/NET0131  & n3640 ;
  assign n10056 = ~n10054 & ~n10055 ;
  assign n10057 = \mix1_data_o_reg_reg[79]/NET0131  & ~n3640 ;
  assign n10058 = \mix1_data_reg_reg[79]/NET0131  & n3640 ;
  assign n10059 = ~n10057 & ~n10058 ;
  assign n10060 = \mix1_data_o_reg_reg[88]/NET0131  & ~n3640 ;
  assign n10061 = \mix1_data_reg_reg[88]/NET0131  & n3640 ;
  assign n10062 = ~n10060 & ~n10061 ;
  assign n10063 = \mix1_data_o_reg_reg[85]/NET0131  & ~n3640 ;
  assign n10064 = \mix1_data_reg_reg[85]/NET0131  & n3640 ;
  assign n10065 = ~n10063 & ~n10064 ;
  assign n10066 = \mix1_data_o_reg_reg[103]/NET0131  & ~n3640 ;
  assign n10067 = \mix1_data_reg_reg[103]/NET0131  & n3640 ;
  assign n10068 = ~n10066 & ~n10067 ;
  assign n10069 = \mix1_data_o_reg_reg[69]/NET0131  & ~n3640 ;
  assign n10070 = \mix1_data_reg_reg[69]/NET0131  & n3640 ;
  assign n10071 = ~n10069 & ~n10070 ;
  assign n10072 = \mix1_data_o_reg_reg[73]/NET0131  & ~n3640 ;
  assign n10073 = \mix1_data_reg_reg[73]/NET0131  & n3640 ;
  assign n10074 = ~n10072 & ~n10073 ;
  assign n10075 = \mix1_data_o_reg_reg[104]/NET0131  & ~n3640 ;
  assign n10076 = \mix1_data_reg_reg[104]/NET0131  & n3640 ;
  assign n10077 = ~n10075 & ~n10076 ;
  assign n10078 = \mix1_data_o_reg_reg[68]/NET0131  & ~n3640 ;
  assign n10079 = \mix1_data_reg_reg[68]/NET0131  & n3640 ;
  assign n10080 = ~n10078 & ~n10079 ;
  assign n10081 = \mix1_data_o_reg_reg[82]/NET0131  & ~n3640 ;
  assign n10082 = \mix1_data_reg_reg[82]/NET0131  & n3640 ;
  assign n10083 = ~n10081 & ~n10082 ;
  assign n10084 = \mix1_data_o_reg_reg[65]/NET0131  & ~n3640 ;
  assign n10085 = \mix1_data_reg_reg[65]/NET0131  & n3640 ;
  assign n10086 = ~n10084 & ~n10085 ;
  assign n10087 = \mix1_data_o_reg_reg[66]/NET0131  & ~n3640 ;
  assign n10088 = \mix1_data_reg_reg[66]/NET0131  & n3640 ;
  assign n10089 = ~n10087 & ~n10088 ;
  assign n10090 = \mix1_data_o_reg_reg[58]/NET0131  & ~n3640 ;
  assign n10091 = \mix1_data_reg_reg[58]/NET0131  & n3640 ;
  assign n10092 = ~n10090 & ~n10091 ;
  assign n10093 = \mix1_data_o_reg_reg[63]/NET0131  & ~n3640 ;
  assign n10094 = \mix1_data_reg_reg[63]/NET0131  & n3640 ;
  assign n10095 = ~n10093 & ~n10094 ;
  assign n10096 = \mix1_data_o_reg_reg[36]/NET0131  & ~n3640 ;
  assign n10097 = \mix1_data_reg_reg[36]/NET0131  & n3640 ;
  assign n10098 = ~n10096 & ~n10097 ;
  assign n10099 = \mix1_data_o_reg_reg[47]/NET0131  & ~n3640 ;
  assign n10100 = \mix1_data_reg_reg[47]/NET0131  & n3640 ;
  assign n10101 = ~n10099 & ~n10100 ;
  assign n10102 = \mix1_data_o_reg_reg[60]/NET0131  & ~n3640 ;
  assign n10103 = \mix1_data_reg_reg[60]/NET0131  & n3640 ;
  assign n10104 = ~n10102 & ~n10103 ;
  assign n10105 = \mix1_data_o_reg_reg[86]/NET0131  & ~n3640 ;
  assign n10106 = \mix1_data_reg_reg[86]/NET0131  & n3640 ;
  assign n10107 = ~n10105 & ~n10106 ;
  assign n10108 = \mix1_data_o_reg_reg[46]/NET0131  & ~n3640 ;
  assign n10109 = \mix1_data_reg_reg[46]/NET0131  & n3640 ;
  assign n10110 = ~n10108 & ~n10109 ;
  assign n10111 = \mix1_data_o_reg_reg[101]/NET0131  & ~n3640 ;
  assign n10112 = \mix1_data_reg_reg[101]/NET0131  & n3640 ;
  assign n10113 = ~n10111 & ~n10112 ;
  assign n10114 = \mix1_data_o_reg_reg[44]/NET0131  & ~n3640 ;
  assign n10115 = \mix1_data_reg_reg[44]/NET0131  & n3640 ;
  assign n10116 = ~n10114 & ~n10115 ;
  assign n10117 = \mix1_data_o_reg_reg[119]/NET0131  & ~n3640 ;
  assign n10118 = \mix1_data_reg_reg[119]/NET0131  & n3640 ;
  assign n10119 = ~n10117 & ~n10118 ;
  assign n10120 = \mix1_data_o_reg_reg[53]/NET0131  & ~n3640 ;
  assign n10121 = \mix1_data_reg_reg[53]/NET0131  & n3640 ;
  assign n10122 = ~n10120 & ~n10121 ;
  assign n10123 = \mix1_data_o_reg_reg[100]/NET0131  & ~n3640 ;
  assign n10124 = \mix1_data_reg_reg[100]/NET0131  & n3640 ;
  assign n10125 = ~n10123 & ~n10124 ;
  assign n10126 = \mix1_data_o_reg_reg[74]/NET0131  & ~n3640 ;
  assign n10127 = \mix1_data_reg_reg[74]/NET0131  & n3640 ;
  assign n10128 = ~n10126 & ~n10127 ;
  assign n10129 = \mix1_data_o_reg_reg[117]/NET0131  & ~n3640 ;
  assign n10130 = \mix1_data_reg_reg[117]/NET0131  & n3640 ;
  assign n10131 = ~n10129 & ~n10130 ;
  assign n10132 = \mix1_data_o_reg_reg[67]/NET0131  & ~n3640 ;
  assign n10133 = \mix1_data_reg_reg[67]/NET0131  & n3640 ;
  assign n10134 = ~n10132 & ~n10133 ;
  assign n10135 = \mix1_data_o_reg_reg[54]/NET0131  & ~n3640 ;
  assign n10136 = \mix1_data_reg_reg[54]/NET0131  & n3640 ;
  assign n10137 = ~n10135 & ~n10136 ;
  assign n10138 = \mix1_data_o_reg_reg[59]/NET0131  & ~n3640 ;
  assign n10139 = \mix1_data_reg_reg[59]/NET0131  & n3640 ;
  assign n10140 = ~n10138 & ~n10139 ;
  assign n10141 = \mix1_data_o_reg_reg[51]/NET0131  & ~n3640 ;
  assign n10142 = \mix1_data_reg_reg[51]/NET0131  & n3640 ;
  assign n10143 = ~n10141 & ~n10142 ;
  assign n10144 = \mix1_data_o_reg_reg[96]/NET0131  & ~n3640 ;
  assign n10145 = \mix1_data_reg_reg[96]/NET0131  & n3640 ;
  assign n10146 = ~n10144 & ~n10145 ;
  assign n10147 = \mix1_data_o_reg_reg[126]/NET0131  & ~n3640 ;
  assign n10148 = \mix1_data_reg_reg[126]/NET0131  & n3640 ;
  assign n10149 = ~n10147 & ~n10148 ;
  assign n10150 = \mix1_data_o_reg_reg[57]/NET0131  & ~n3640 ;
  assign n10151 = \mix1_data_reg_reg[57]/NET0131  & n3640 ;
  assign n10152 = ~n10150 & ~n10151 ;
  assign n10153 = \mix1_data_o_reg_reg[102]/NET0131  & ~n3640 ;
  assign n10154 = \mix1_data_reg_reg[102]/NET0131  & n3640 ;
  assign n10155 = ~n10153 & ~n10154 ;
  assign n10156 = \mix1_data_o_reg_reg[55]/NET0131  & ~n3640 ;
  assign n10157 = \mix1_data_reg_reg[55]/NET0131  & n3640 ;
  assign n10158 = ~n10156 & ~n10157 ;
  assign n10159 = ~n1274 & ~n1286 ;
  assign n10160 = \key_i[41]_pad  & ~n1116 ;
  assign n10161 = \ks1_key_reg_reg[41]/P0002  & n1116 ;
  assign n10162 = ~n10160 & ~n10161 ;
  assign n10163 = n3244 & n10162 ;
  assign n10164 = ~n3244 & ~n10162 ;
  assign n10165 = ~n10163 & ~n10164 ;
  assign n10166 = ~n1554 & ~n10165 ;
  assign n10167 = n1554 & n10165 ;
  assign n10168 = ~n10166 & ~n10167 ;
  assign n10169 = n929 & ~n10168 ;
  assign n10170 = \ks1_key_reg_reg[9]/NET0131  & ~n929 ;
  assign n10171 = ~n10169 & ~n10170 ;
  assign n10172 = ~\ks1_key_reg_reg[108]/NET0131  & n1116 ;
  assign n10173 = ~\key_i[108]_pad  & ~n1116 ;
  assign n10174 = ~n10172 & ~n10173 ;
  assign n10175 = n2764 & ~n10174 ;
  assign n10176 = ~n2764 & n10174 ;
  assign n10177 = ~n10175 & ~n10176 ;
  assign n10178 = ~\ks1_key_reg_reg[107]/NET0131  & n1116 ;
  assign n10179 = ~\key_i[107]_pad  & ~n1116 ;
  assign n10180 = ~n10178 & ~n10179 ;
  assign n10181 = n2744 & ~n10180 ;
  assign n10182 = ~n2744 & n10180 ;
  assign n10183 = ~n10181 & ~n10182 ;
  assign n10184 = \key_i[44]_pad  & ~n1116 ;
  assign n10185 = \ks1_key_reg_reg[44]/P0002  & n1116 ;
  assign n10186 = ~n10184 & ~n10185 ;
  assign n10187 = \key_i[76]_pad  & ~n1116 ;
  assign n10188 = \ks1_key_reg_reg[76]/P0002  & n1116 ;
  assign n10189 = ~n10187 & ~n10188 ;
  assign n10190 = n10177 & n10189 ;
  assign n10191 = ~n10177 & ~n10189 ;
  assign n10192 = ~n10190 & ~n10191 ;
  assign n10193 = n10186 & n10192 ;
  assign n10194 = ~n10186 & ~n10192 ;
  assign n10195 = ~n10193 & ~n10194 ;
  assign n10196 = ~n1283 & ~n10195 ;
  assign n10197 = n1283 & n10195 ;
  assign n10198 = ~n10196 & ~n10197 ;
  assign n10199 = n929 & ~n10198 ;
  assign n10200 = \ks1_key_reg_reg[12]/NET0131  & ~n929 ;
  assign n10201 = ~n10199 & ~n10200 ;
  assign n10202 = ~\ks1_key_reg_reg[75]/P0002  & n1116 ;
  assign n10203 = ~\key_i[75]_pad  & ~n1116 ;
  assign n10204 = ~n10202 & ~n10203 ;
  assign n10205 = n10183 & ~n10204 ;
  assign n10206 = ~n10183 & n10204 ;
  assign n10207 = ~n10205 & ~n10206 ;
  assign n10208 = ~\ks1_key_reg_reg[43]/P0002  & n1116 ;
  assign n10209 = ~\key_i[43]_pad  & ~n1116 ;
  assign n10210 = ~n10208 & ~n10209 ;
  assign n10211 = n10207 & ~n10210 ;
  assign n10212 = ~n10207 & n10210 ;
  assign n10213 = ~n10211 & ~n10212 ;
  assign n10214 = n1527 & ~n10213 ;
  assign n10215 = ~n1527 & n10213 ;
  assign n10216 = ~n10214 & ~n10215 ;
  assign n10217 = n929 & ~n10216 ;
  assign n10218 = \ks1_key_reg_reg[11]/NET0131  & ~n929 ;
  assign n10219 = ~n10217 & ~n10218 ;
  assign n10220 = ~\ks1_key_reg_reg[109]/P0002  & n1116 ;
  assign n10221 = ~\key_i[109]_pad  & ~n1116 ;
  assign n10222 = ~n10220 & ~n10221 ;
  assign n10223 = n2456 & ~n10222 ;
  assign n10224 = ~n2456 & n10222 ;
  assign n10225 = ~n10223 & ~n10224 ;
  assign n10226 = ~\ks1_key_reg_reg[77]/P0002  & n1116 ;
  assign n10227 = ~\key_i[77]_pad  & ~n1116 ;
  assign n10228 = ~n10226 & ~n10227 ;
  assign n10229 = n10225 & ~n10228 ;
  assign n10230 = ~n10225 & n10228 ;
  assign n10231 = ~n10229 & ~n10230 ;
  assign n10232 = ~\ks1_key_reg_reg[45]/P0002  & n1116 ;
  assign n10233 = ~\key_i[45]_pad  & ~n1116 ;
  assign n10234 = ~n10232 & ~n10233 ;
  assign n10235 = n10231 & ~n10234 ;
  assign n10236 = ~n10231 & n10234 ;
  assign n10237 = ~n10235 & ~n10236 ;
  assign n10238 = n1911 & ~n10237 ;
  assign n10239 = ~n1911 & n10237 ;
  assign n10240 = ~n10238 & ~n10239 ;
  assign n10241 = n929 & ~n10240 ;
  assign n10242 = \ks1_key_reg_reg[13]/NET0131  & ~n929 ;
  assign n10243 = ~n10241 & ~n10242 ;
  assign n10244 = ~\ks1_key_reg_reg[79]/P0002  & n1116 ;
  assign n10245 = ~\key_i[79]_pad  & ~n1116 ;
  assign n10246 = ~n10244 & ~n10245 ;
  assign n10247 = n3569 & ~n10246 ;
  assign n10248 = ~n3569 & n10246 ;
  assign n10249 = ~n10247 & ~n10248 ;
  assign n10250 = ~n2202 & n2214 ;
  assign n10251 = n1928 & ~n2214 ;
  assign n10252 = ~n10250 & ~n10251 ;
  assign n10253 = n2193 & ~n2294 ;
  assign n10254 = n2238 & ~n2245 ;
  assign n10255 = n3570 & ~n10254 ;
  assign n10256 = ~n3570 & n10254 ;
  assign n10257 = ~n10255 & ~n10256 ;
  assign n10258 = n10253 & ~n10257 ;
  assign n10259 = ~n10253 & n10257 ;
  assign n10260 = ~n10258 & ~n10259 ;
  assign n10261 = n10252 & n10260 ;
  assign n10262 = ~n10252 & ~n10260 ;
  assign n10263 = ~n10261 & ~n10262 ;
  assign n10264 = ~\ks1_key_reg_reg[47]/P0002  & n1116 ;
  assign n10265 = ~\key_i[47]_pad  & ~n1116 ;
  assign n10266 = ~n10264 & ~n10265 ;
  assign n10267 = n10249 & ~n10266 ;
  assign n10268 = ~n10249 & n10266 ;
  assign n10269 = ~n10267 & ~n10268 ;
  assign n10270 = n2084 & ~n10269 ;
  assign n10271 = ~n2084 & n10269 ;
  assign n10272 = ~n10270 & ~n10271 ;
  assign n10273 = n929 & ~n10272 ;
  assign n10274 = \ks1_key_reg_reg[15]/NET0131  & ~n929 ;
  assign n10275 = ~n10273 & ~n10274 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g27929/_0_  = n1140 ;
  assign \g27942/_3_  = n2270 ;
  assign \g27943/_3_  = ~n2282 ;
  assign \g27944/_3_  = n2301 ;
  assign \g27945/_0_  = ~n2372 ;
  assign \g27995/_0_  = ~n2417 ;
  assign \g27998/_0_  = n1134 ;
  assign \g28019/_0_  = ~n2438 ;
  assign \g28020/_0_  = ~n2461 ;
  assign \g28021/_0_  = ~n2474 ;
  assign \g28022/_0_  = ~n2485 ;
  assign \g28023/_0_  = ~n2503 ;
  assign \g28024/_0_  = ~n2514 ;
  assign \g28025/_0_  = ~n2526 ;
  assign \g28026/_0_  = ~n2537 ;
  assign \g28027/_0_  = ~n2549 ;
  assign \g28028/_0_  = ~n2560 ;
  assign \g28029/_0_  = ~n2568 ;
  assign \g28030/_0_  = ~n2574 ;
  assign \g28031/_0_  = ~n2586 ;
  assign \g28032/_0_  = ~n2597 ;
  assign \g28033/_0_  = ~n2609 ;
  assign \g28034/_0_  = ~n2620 ;
  assign \g28044/_0_  = ~n2630 ;
  assign \g28045/_0_  = ~n2638 ;
  assign \g28046/_0_  = ~n2648 ;
  assign \g28047/_0_  = ~n2656 ;
  assign \g28048/_0_  = ~n2665 ;
  assign \g28049/_0_  = ~n2673 ;
  assign \g28050/_0_  = ~n2682 ;
  assign \g28051/_0_  = ~n2690 ;
  assign \g28151/_0_  = ~n1128 ;
  assign \g28177/_0_  = ~n2696 ;
  assign \g28178/_0_  = ~n2718 ;
  assign \g28179/_0_  = ~n2729 ;
  assign \g28180/_0_  = ~n2749 ;
  assign \g28181/_0_  = ~n2769 ;
  assign \g28182/_0_  = ~n2780 ;
  assign \g28183/_0_  = ~n2791 ;
  assign \g28184/_0_  = ~n2802 ;
  assign \g28185/_0_  = ~n2813 ;
  assign \g28186/_0_  = ~n2824 ;
  assign \g28187/_0_  = ~n2835 ;
  assign \g28188/_0_  = ~n2841 ;
  assign \g28189/_0_  = ~n2852 ;
  assign \g28190/_0_  = ~n2858 ;
  assign \g28191/_0_  = ~n2869 ;
  assign \g28192/_0_  = ~n2880 ;
  assign \g28193/_0_  = ~n2891 ;
  assign \g28194/_0_  = ~n2902 ;
  assign \g28195/_0_  = ~n2913 ;
  assign \g28196/_0_  = ~n2924 ;
  assign \g28197/_0_  = ~n2935 ;
  assign \g28198/_0_  = ~n2941 ;
  assign \g28199/_0_  = ~n2952 ;
  assign \g28200/_0_  = ~n2963 ;
  assign \g28201/_0_  = ~n2974 ;
  assign \g28202/_0_  = ~n2985 ;
  assign \g28203/_0_  = ~n2996 ;
  assign \g28253/_0_  = ~n3004 ;
  assign \g28254/_0_  = ~n3012 ;
  assign \g28255/_0_  = ~n3020 ;
  assign \g28256/_0_  = ~n3028 ;
  assign \g28257/_0_  = ~n3036 ;
  assign \g28258/_0_  = ~n3039 ;
  assign \g28259/_0_  = ~n3042 ;
  assign \g28260/_0_  = ~n3050 ;
  assign \g28261/_0_  = ~n3053 ;
  assign \g28262/_0_  = ~n3061 ;
  assign \g28263/_0_  = ~n3064 ;
  assign \g28264/_0_  = ~n3067 ;
  assign \g28265/_0_  = ~n3070 ;
  assign \g28266/_0_  = ~n3078 ;
  assign \g28267/_0_  = ~n3086 ;
  assign \g28268/_0_  = ~n3094 ;
  assign \g28269/_0_  = ~n3102 ;
  assign \g28270/_0_  = ~n3110 ;
  assign \g28271/_0_  = ~n3118 ;
  assign \g28272/_0_  = ~n3126 ;
  assign \g28273/_0_  = ~n3134 ;
  assign \g28274/_0_  = ~n3142 ;
  assign \g28275/_0_  = ~n3153 ;
  assign \g28276/_0_  = ~n3164 ;
  assign \g28277/_0_  = ~n3175 ;
  assign \g28278/_0_  = ~n3186 ;
  assign \g28279/_0_  = ~n3197 ;
  assign \g28384/_2_  = ~n3201 ;
  assign \g28385/_2_  = ~n3204 ;
  assign \g28388/_2_  = ~n3208 ;
  assign \g28389/_2_  = ~n3211 ;
  assign \g28394/_2_  = ~n3215 ;
  assign \g28395/_2_  = ~n3218 ;
  assign \g28401/_2_  = ~n3222 ;
  assign \g28402/_2_  = ~n3225 ;
  assign \g28403/_0_  = ~n3246 ;
  assign \g28404/_0_  = ~n3249 ;
  assign \g28408/_0_  = ~n2412 ;
  assign \g28410/_0_  = n2360 ;
  assign \g28440/_0_  = ~n3260 ;
  assign \g28441/_0_  = ~n3271 ;
  assign \g28442/_0_  = ~n3282 ;
  assign \g28443/_0_  = ~n3293 ;
  assign \g28444/_0_  = ~n3299 ;
  assign \g28445/_0_  = ~n3305 ;
  assign \g28446/_0_  = ~n3316 ;
  assign \g28447/_0_  = ~n3327 ;
  assign \g28448/_0_  = ~n3338 ;
  assign \g28449/_0_  = ~n3349 ;
  assign \g28450/_0_  = ~n3360 ;
  assign \g28451/_0_  = ~n3371 ;
  assign \g28452/_0_  = ~n3382 ;
  assign \g28453/_0_  = ~n3393 ;
  assign \g28538/_0_  = ~n3401 ;
  assign \g28539/_0_  = ~n3409 ;
  assign \g28540/_0_  = n3412 ;
  assign \g28541/_0_  = n3415 ;
  assign \g28542/_0_  = n3418 ;
  assign \g28543/_0_  = ~n3421 ;
  assign \g28544/_0_  = ~n3429 ;
  assign \g28545/_0_  = ~n3432 ;
  assign \g28546/_0_  = n3435 ;
  assign \g28547/_0_  = n3438 ;
  assign \g28548/_0_  = ~n3441 ;
  assign \g28549/_0_  = ~n3444 ;
  assign \g28550/_0_  = n3447 ;
  assign \g28551/_0_  = ~n3450 ;
  assign \g28552/_0_  = ~n3453 ;
  assign \g28557/_0_  = ~n3461 ;
  assign \g28558/_0_  = ~n3469 ;
  assign \g28563/_0_  = ~n3477 ;
  assign \g28564/_0_  = ~n3485 ;
  assign \g28565/_0_  = ~n3493 ;
  assign \g28566/_0_  = ~n3504 ;
  assign \g28567/_0_  = ~n3515 ;
  assign \g28625/_2_  = n3518 ;
  assign \g28626/_2_  = n3521 ;
  assign \g28633/_2_  = n3524 ;
  assign \g28639/_2_  = n3527 ;
  assign \g28655/_2_  = n3530 ;
  assign \g28656/_2_  = ~n3533 ;
  assign \g28657/_2_  = ~n3536 ;
  assign \g28660/_2_  = n3539 ;
  assign \g28661/_2_  = ~n3542 ;
  assign \g28662/_2_  = ~n3545 ;
  assign \g28666/_2_  = n3548 ;
  assign \g28667/_2_  = ~n3551 ;
  assign \g28668/_2_  = ~n3554 ;
  assign \g28678/_2_  = n3557 ;
  assign \g28679/_2_  = ~n3560 ;
  assign \g28680/_2_  = ~n3563 ;
  assign \g28690/_0_  = ~n3569 ;
  assign \g28710/_0_  = ~n2354 ;
  assign \g28716/_0_  = ~n3572 ;
  assign \g28795/_0_  = ~n3575 ;
  assign \g28796/_0_  = ~n3578 ;
  assign \g28798/_0_  = ~n3581 ;
  assign \g28799/_0_  = ~n3584 ;
  assign \g28800/_0_  = ~n3587 ;
  assign \g28801/_0_  = ~n3590 ;
  assign \g28804/_0_  = n2214 ;
  assign \g28825/_2_  = ~n3593 ;
  assign \g28826/_2_  = ~n3596 ;
  assign \g28830/_2_  = ~n3599 ;
  assign \g28834/_2_  = ~n3602 ;
  assign \g28842/_2_  = ~n3605 ;
  assign \g28843/_2_  = ~n3608 ;
  assign \g28845/_2_  = ~n3611 ;
  assign \g28848/_2_  = ~n3614 ;
  assign \g28890/_0_  = n3241 ;
  assign \g28936/_0_  = n3616 ;
  assign \g28982/_0_  = ~n3618 ;
  assign \g29050/_0_  = ~n4076 ;
  assign \g29051/_0_  = ~n4264 ;
  assign \g29052/_0_  = ~n4389 ;
  assign \g29053/_0_  = ~n4451 ;
  assign \g29054/_0_  = ~n4488 ;
  assign \g29055/_0_  = ~n4531 ;
  assign \g29056/_0_  = n4549 ;
  assign \g29057/_0_  = ~n4574 ;
  assign \g29058/_0_  = ~n4583 ;
  assign \g29059/_0_  = ~n4605 ;
  assign \g29060/_0_  = n4620 ;
  assign \g29061/_0_  = ~n4626 ;
  assign \g29328/_0_  = n4651 ;
  assign \g29329/_0_  = ~n4664 ;
  assign \g29330/_0_  = ~n4677 ;
  assign \g29331/_0_  = n4705 ;
  assign \g29332/_0_  = ~n4730 ;
  assign \g29333/_0_  = n4755 ;
  assign \g29334/_0_  = ~n4774 ;
  assign \g29335/_0_  = ~n4796 ;
  assign \g29336/_0_  = n4811 ;
  assign \g29337/_0_  = ~n4820 ;
  assign \g29338/_0_  = ~n4826 ;
  assign \g29339/_0_  = ~n4841 ;
  assign \g29340/_0_  = ~n4850 ;
  assign \g29341/_0_  = ~n4859 ;
  assign \g29342/_0_  = ~n4862 ;
  assign \g29343/_0_  = ~n4865 ;
  assign \g29344/_0_  = ~n4868 ;
  assign \g29345/_0_  = ~n4871 ;
  assign \g29346/_0_  = ~n4874 ;
  assign \g29347/_0_  = ~n4877 ;
  assign \g29348/_0_  = ~n4880 ;
  assign \g29349/_0_  = ~n4883 ;
  assign \g29350/_0_  = n4886 ;
  assign \g29351/_0_  = ~n4889 ;
  assign \g29352/_0_  = n4892 ;
  assign \g29353/_0_  = ~n4895 ;
  assign \g29354/_0_  = ~n4898 ;
  assign \g29355/_0_  = ~n4901 ;
  assign \g29356/_0_  = ~n4904 ;
  assign \g29357/_0_  = ~n4907 ;
  assign \g29358/_0_  = ~n4910 ;
  assign \g29359/_0_  = ~n4913 ;
  assign \g29360/_0_  = n4916 ;
  assign \g29361/_0_  = ~n4919 ;
  assign \g29362/_0_  = ~n4922 ;
  assign \g29363/_0_  = n4925 ;
  assign \g29364/_0_  = ~n4928 ;
  assign \g29365/_0_  = ~n4931 ;
  assign \g29366/_0_  = ~n4943 ;
  assign \g29367/_0_  = ~n4955 ;
  assign \g29395/_0_  = ~n5021 ;
  assign \g29396/_0_  = n5024 ;
  assign \g29453/_0_  = ~n5061 ;
  assign \g29454/_0_  = ~n5091 ;
  assign \g29455/_0_  = ~n5121 ;
  assign \g29456/_0_  = ~n5151 ;
  assign \g29457/_0_  = ~n5181 ;
  assign \g29458/_0_  = ~n5211 ;
  assign \g29459/_0_  = ~n5241 ;
  assign \g29460/_0_  = ~n5271 ;
  assign \g29461/_0_  = ~n5301 ;
  assign \g29462/_0_  = ~n5331 ;
  assign \g29463/_0_  = ~n5361 ;
  assign \g29464/_0_  = ~n5391 ;
  assign \g29465/_0_  = ~n5421 ;
  assign \g29466/_0_  = ~n5451 ;
  assign \g29467/_0_  = ~n5481 ;
  assign \g29468/_0_  = ~n5511 ;
  assign \g29469/_0_  = ~n5541 ;
  assign \g29470/_0_  = ~n5571 ;
  assign \g29471/_0_  = ~n5601 ;
  assign \g29472/_0_  = ~n5631 ;
  assign \g29473/_0_  = ~n5661 ;
  assign \g29474/_0_  = ~n5691 ;
  assign \g29475/_0_  = ~n5721 ;
  assign \g29476/_0_  = ~n5751 ;
  assign \g29477/_0_  = ~n5781 ;
  assign \g29478/_0_  = ~n5811 ;
  assign \g29479/_0_  = ~n5841 ;
  assign \g29480/_0_  = ~n5871 ;
  assign \g29481/_0_  = ~n5901 ;
  assign \g29482/_0_  = ~n5931 ;
  assign \g29483/_0_  = ~n5961 ;
  assign \g29484/_0_  = ~n5991 ;
  assign \g29485/_0_  = ~n6021 ;
  assign \g29486/_0_  = ~n6051 ;
  assign \g29487/_0_  = ~n6081 ;
  assign \g29488/_0_  = ~n6111 ;
  assign \g29489/_0_  = ~n6141 ;
  assign \g29490/_0_  = ~n6171 ;
  assign \g29491/_0_  = ~n6201 ;
  assign \g29492/_0_  = ~n6231 ;
  assign \g29493/_0_  = ~n6261 ;
  assign \g29494/_0_  = ~n6291 ;
  assign \g29495/_0_  = ~n6321 ;
  assign \g29496/_0_  = ~n6351 ;
  assign \g29497/_0_  = ~n6381 ;
  assign \g29498/_0_  = ~n6411 ;
  assign \g29499/_0_  = ~n6441 ;
  assign \g29500/_0_  = ~n6471 ;
  assign \g29501/_0_  = ~n6501 ;
  assign \g29502/_0_  = ~n6531 ;
  assign \g29503/_0_  = ~n6561 ;
  assign \g29504/_0_  = ~n6591 ;
  assign \g29505/_0_  = ~n6621 ;
  assign \g29506/_0_  = ~n6651 ;
  assign \g29507/_0_  = ~n6681 ;
  assign \g29508/_0_  = ~n6711 ;
  assign \g29509/_0_  = ~n6741 ;
  assign \g29510/_0_  = ~n6771 ;
  assign \g29511/_0_  = ~n6801 ;
  assign \g29512/_0_  = ~n6831 ;
  assign \g29513/_0_  = ~n6861 ;
  assign \g29514/_0_  = ~n6891 ;
  assign \g29515/_0_  = ~n6921 ;
  assign \g29516/_0_  = ~n6951 ;
  assign \g29517/_0_  = ~n6981 ;
  assign \g29518/_0_  = ~n7011 ;
  assign \g29519/_0_  = ~n7041 ;
  assign \g29520/_0_  = ~n7071 ;
  assign \g29521/_0_  = ~n7101 ;
  assign \g29522/_0_  = ~n7131 ;
  assign \g29523/_0_  = ~n7161 ;
  assign \g29524/_0_  = ~n7191 ;
  assign \g29525/_0_  = ~n7221 ;
  assign \g29526/_0_  = ~n7251 ;
  assign \g29527/_0_  = ~n7280 ;
  assign \g29528/_0_  = ~n7310 ;
  assign \g29529/_0_  = ~n7340 ;
  assign \g29530/_0_  = ~n7370 ;
  assign \g29531/_0_  = ~n7400 ;
  assign \g29532/_0_  = ~n7430 ;
  assign \g29533/_0_  = ~n7460 ;
  assign \g29534/_0_  = ~n7490 ;
  assign \g29535/_0_  = ~n7520 ;
  assign \g29536/_0_  = ~n7550 ;
  assign \g29537/_0_  = ~n7580 ;
  assign \g29538/_0_  = ~n7610 ;
  assign \g29539/_0_  = ~n7640 ;
  assign \g29540/_0_  = ~n7670 ;
  assign \g29541/_0_  = ~n7700 ;
  assign \g29542/_0_  = ~n7730 ;
  assign \g29543/_0_  = ~n7760 ;
  assign \g29544/_0_  = ~n7790 ;
  assign \g29545/_0_  = ~n7820 ;
  assign \g29546/_0_  = ~n7850 ;
  assign \g29547/_0_  = ~n7880 ;
  assign \g29548/_0_  = ~n7910 ;
  assign \g29549/_0_  = ~n7940 ;
  assign \g29550/_0_  = ~n7970 ;
  assign \g29551/_0_  = ~n8000 ;
  assign \g29552/_0_  = ~n8030 ;
  assign \g29553/_0_  = ~n8060 ;
  assign \g29554/_0_  = ~n8090 ;
  assign \g29555/_0_  = ~n8120 ;
  assign \g29556/_0_  = ~n8150 ;
  assign \g29557/_0_  = ~n8180 ;
  assign \g29558/_0_  = ~n8210 ;
  assign \g29559/_0_  = ~n8240 ;
  assign \g29560/_0_  = ~n8270 ;
  assign \g29561/_0_  = ~n8300 ;
  assign \g29562/_0_  = ~n8330 ;
  assign \g29563/_0_  = ~n8360 ;
  assign \g29564/_0_  = ~n8390 ;
  assign \g29565/_0_  = ~n8420 ;
  assign \g29566/_0_  = ~n8450 ;
  assign \g29567/_0_  = ~n8480 ;
  assign \g29568/_0_  = ~n8510 ;
  assign \g29569/_0_  = ~n8540 ;
  assign \g29570/_0_  = ~n8570 ;
  assign \g29571/_0_  = ~n8600 ;
  assign \g29572/_0_  = ~n8630 ;
  assign \g29573/_0_  = ~n8660 ;
  assign \g29574/_0_  = ~n8690 ;
  assign \g29575/_0_  = ~n8720 ;
  assign \g29576/_0_  = ~n8750 ;
  assign \g29577/_0_  = ~n8780 ;
  assign \g29578/_0_  = ~n8810 ;
  assign \g29579/_0_  = ~n8840 ;
  assign \g29580/_0_  = ~n8870 ;
  assign \g29582/_0_  = ~n8873 ;
  assign \g29583/_0_  = ~n8876 ;
  assign \g29584/_0_  = ~n8879 ;
  assign \g29585/_0_  = ~n8882 ;
  assign \g29586/_0_  = n8885 ;
  assign \g29587/_0_  = ~n8888 ;
  assign \g29588/_0_  = ~n8891 ;
  assign \g29589/_0_  = n8894 ;
  assign \g29590/_0_  = ~n8897 ;
  assign \g29591/_0_  = ~n8900 ;
  assign \g29592/_0_  = ~n8903 ;
  assign \g29593/_0_  = ~n8906 ;
  assign \g29634/_0_  = n8931 ;
  assign \g29635/_0_  = n8958 ;
  assign \g29636/_0_  = n8985 ;
  assign \g29637/_0_  = n9011 ;
  assign \g29645/_0_  = ~n9042 ;
  assign \g29646/_0_  = ~n9074 ;
  assign \g29647/_0_  = ~n9104 ;
  assign \g29824/_0_  = ~n9114 ;
  assign \g29828/_0_  = ~n9124 ;
  assign \g29832/_0_  = ~n9136 ;
  assign \g29836/_0_  = ~n9139 ;
  assign \g29837/_0_  = ~n9142 ;
  assign \g29838/_0_  = n9145 ;
  assign \g29839/_0_  = ~n9148 ;
  assign \g29840/_0_  = ~n9151 ;
  assign \g29841/_0_  = n9154 ;
  assign \g29842/_0_  = ~n9157 ;
  assign \g29843/_0_  = n9160 ;
  assign \g29844/_0_  = ~n9163 ;
  assign \g29845/_0_  = ~n9166 ;
  assign \g29846/_0_  = n9169 ;
  assign \g29847/_0_  = ~n9172 ;
  assign \g29848/_0_  = ~n9175 ;
  assign \g29849/_0_  = ~n9178 ;
  assign \g29850/_0_  = ~n9181 ;
  assign \g29851/_0_  = ~n9184 ;
  assign \g29852/_0_  = ~n9187 ;
  assign \g29853/_0_  = ~n9190 ;
  assign \g29854/_0_  = n9193 ;
  assign \g29855/_0_  = ~n9196 ;
  assign \g29856/_0_  = ~n9199 ;
  assign \g29857/_0_  = n9202 ;
  assign \g29858/_0_  = ~n9205 ;
  assign \g29859/_0_  = n9208 ;
  assign \g29860/_0_  = ~n9211 ;
  assign \g29861/_0_  = ~n9214 ;
  assign \g29862/_0_  = n9217 ;
  assign \g29863/_0_  = ~n9220 ;
  assign \g29864/_0_  = ~n9223 ;
  assign \g29865/_0_  = ~n9226 ;
  assign \g29866/_0_  = ~n9229 ;
  assign \g29867/_0_  = ~n9232 ;
  assign \g29868/_0_  = n9241 ;
  assign \g30081/_0_  = n9244 ;
  assign \g30082/_0_  = ~n9247 ;
  assign \g30083/_0_  = n9250 ;
  assign \g30084/_0_  = ~n9253 ;
  assign \g30085/_0_  = ~n9256 ;
  assign \g30086/_0_  = ~n9259 ;
  assign \g30087/_0_  = n9262 ;
  assign \g30088/_0_  = ~n9265 ;
  assign \g30089/_0_  = ~n9268 ;
  assign \g30090/_0_  = ~n9271 ;
  assign \g30091/_0_  = ~n9274 ;
  assign \g30092/_0_  = ~n9277 ;
  assign \g30093/_0_  = ~n9280 ;
  assign \g30094/_0_  = n9283 ;
  assign \g30095/_0_  = ~n9286 ;
  assign \g30096/_0_  = ~n9289 ;
  assign \g30135/_0_  = ~n9292 ;
  assign \g30137/_0_  = n9295 ;
  assign \g30164/_0_  = n9039 ;
  assign \g30165/_0_  = n9071 ;
  assign \g30166/_0_  = n9101 ;
  assign \g30167/_0_  = ~n8928 ;
  assign \g30168/_0_  = ~n8955 ;
  assign \g30169/_0_  = ~n8982 ;
  assign \g30170/_0_  = ~n9008 ;
  assign \g30231/_0_  = n9298 ;
  assign \g30232/_0_  = ~n9301 ;
  assign \g30233/_0_  = ~n9304 ;
  assign \g30234/_0_  = ~n9307 ;
  assign \g30235/_0_  = n9310 ;
  assign \g30236/_0_  = ~n9313 ;
  assign \g30237/_0_  = ~n9316 ;
  assign \g30238/_0_  = ~n9319 ;
  assign \g30286/_0_  = ~n9346 ;
  assign \g30287/_0_  = ~n9373 ;
  assign \g30288/_0_  = ~n9400 ;
  assign \g30289/_0_  = ~n9421 ;
  assign \g30290/_0_  = ~n9442 ;
  assign \g30291/_0_  = ~n9463 ;
  assign \g30292/_0_  = ~n9484 ;
  assign \g30293/_0_  = ~n9505 ;
  assign \g30294/_0_  = ~n9532 ;
  assign \g30295/_0_  = ~n9559 ;
  assign \g30296/_0_  = ~n9586 ;
  assign \g30297/_0_  = ~n9613 ;
  assign \g30298/_0_  = ~n9640 ;
  assign \g30299/_0_  = ~n9667 ;
  assign \g30300/_0_  = ~n9694 ;
  assign \g30301/_0_  = ~n9721 ;
  assign \g30303/_0_  = n9724 ;
  assign \g30304/_0_  = n9727 ;
  assign \g30305/_0_  = n9730 ;
  assign \g30306/_0_  = n9733 ;
  assign \g30307/_0_  = n9736 ;
  assign \g30308/_0_  = n9739 ;
  assign \g30309/_0_  = n9742 ;
  assign \g30310/_0_  = n9745 ;
  assign \g30311/_0_  = n9748 ;
  assign \g30312/_0_  = n9751 ;
  assign \g30313/_0_  = n9754 ;
  assign \g30314/_0_  = n9757 ;
  assign \g30315/_0_  = n9760 ;
  assign \g30316/_0_  = n9763 ;
  assign \g30317/_0_  = n9766 ;
  assign \g30318/_0_  = n5012 ;
  assign \g30319/_0_  = n9769 ;
  assign \g30481/_0_  = n9772 ;
  assign \g30482/_0_  = ~n9775 ;
  assign \g30483/_0_  = ~n9778 ;
  assign \g30484/_0_  = ~n9781 ;
  assign \g30493/_0_  = n8922 ;
  assign \g30495/_0_  = n8976 ;
  assign \g30536/_0_  = ~n9033 ;
  assign \g30537/_0_  = ~n9065 ;
  assign \g30538/_0_  = ~n9095 ;
  assign \g30735/_0_  = ~n5006 ;
  assign \g30927/_0_  = n9092 ;
  assign \g30928/_0_  = n9030 ;
  assign \g30929/_0_  = n9062 ;
  assign \g30971/_0_  = ~n8996 ;
  assign \g30972/_0_  = ~n8916 ;
  assign \g30973/_0_  = ~n8943 ;
  assign \g30974/_0_  = ~n8970 ;
  assign \g31129/_0_  = n9412 ;
  assign \g31130/_0_  = n9433 ;
  assign \g31131/_0_  = n9454 ;
  assign \g31132/_0_  = n9475 ;
  assign \g31133/_0_  = n9496 ;
  assign \g31134/_0_  = n9337 ;
  assign \g31135/_0_  = n9523 ;
  assign \g31136/_0_  = n9550 ;
  assign \g31137/_0_  = n9577 ;
  assign \g31138/_0_  = n9604 ;
  assign \g31139/_0_  = n9364 ;
  assign \g31140/_0_  = n9631 ;
  assign \g31141/_0_  = n9658 ;
  assign \g31142/_0_  = n9685 ;
  assign \g31143/_0_  = n9712 ;
  assign \g31144/_0_  = n9391 ;
  assign \g31352/_0_  = ~n9406 ;
  assign \g31353/_0_  = ~n9547 ;
  assign \g31354/_0_  = ~n9334 ;
  assign \g31355/_0_  = ~n9655 ;
  assign \g31356/_0_  = ~n9427 ;
  assign \g31357/_0_  = ~n9448 ;
  assign \g31358/_0_  = ~n9469 ;
  assign \g31359/_0_  = ~n9490 ;
  assign \g31360/_0_  = ~n9520 ;
  assign \g31361/_0_  = ~n9574 ;
  assign \g31362/_0_  = ~n9628 ;
  assign \g31363/_0_  = ~n9682 ;
  assign \g31364/_0_  = ~n9709 ;
  assign \g31365/_0_  = ~n9601 ;
  assign \g31366/_0_  = ~n9361 ;
  assign \g31367/_0_  = ~n9388 ;
  assign \g31706/_0_  = ~n9782 ;
  assign \g32001/_0_  = ~n9784 ;
  assign \g32008/_0_  = ~n9788 ;
  assign \g32009/_0_  = ~n9792 ;
  assign \g32010/_0_  = ~n9796 ;
  assign \g32011/_0_  = ~n9797 ;
  assign \g32118/_0_  = ~n9820 ;
  assign \g33261/_0_  = ~n9830 ;
  assign \g33262/_0_  = ~n9831 ;
  assign \g33263/_0_  = ~n9832 ;
  assign \g33264/_0_  = ~n9839 ;
  assign \g33265/_0_  = ~n9843 ;
  assign \g33266/_0_  = ~n9854 ;
  assign \g33450/_0_  = n9857 ;
  assign \g33451/_0_  = n9859 ;
  assign \g33453/_0_  = n9866 ;
  assign \g33485/_0_  = ~n9867 ;
  assign \g33679/_2_  = n9868 ;
  assign \g34838/_2_  = ~n9870 ;
  assign \g34971/_0_  = ~n9873 ;
  assign \g34972/_0_  = ~n9876 ;
  assign \g34973/_0_  = ~n9879 ;
  assign \g34974/_0_  = ~n9882 ;
  assign \g34975/_0_  = ~n9885 ;
  assign \g34976/_0_  = ~n9888 ;
  assign \g34977/_0_  = ~n9891 ;
  assign \g34978/_0_  = ~n9894 ;
  assign \g34979/_0_  = ~n9897 ;
  assign \g34980/_0_  = ~n9900 ;
  assign \g34981/_0_  = ~n9903 ;
  assign \g34982/_0_  = ~n9906 ;
  assign \g34983/_0_  = ~n9909 ;
  assign \g34984/_0_  = ~n9912 ;
  assign \g34985/_0_  = ~n9915 ;
  assign \g34986/_0_  = ~n9918 ;
  assign \g34987/_0_  = ~n9921 ;
  assign \g34988/_0_  = ~n9924 ;
  assign \g34989/_0_  = ~n9927 ;
  assign \g34990/_0_  = ~n9930 ;
  assign \g34991/_0_  = ~n9933 ;
  assign \g34992/_0_  = ~n9936 ;
  assign \g34993/_0_  = ~n9939 ;
  assign \g34994/_0_  = ~n9942 ;
  assign \g34995/_0_  = ~n9945 ;
  assign \g34996/_0_  = ~n9948 ;
  assign \g34997/_0_  = ~n9951 ;
  assign \g34998/_0_  = ~n9954 ;
  assign \g34999/_0_  = ~n9957 ;
  assign \g35000/_0_  = ~n9960 ;
  assign \g35001/_0_  = ~n9963 ;
  assign \g35002/_0_  = ~n9966 ;
  assign \g35003/_0_  = ~n9969 ;
  assign \g35004/_0_  = ~n9972 ;
  assign \g35005/_0_  = ~n9975 ;
  assign \g35006/_0_  = ~n9978 ;
  assign \g35007/_0_  = ~n9981 ;
  assign \g35008/_0_  = ~n9984 ;
  assign \g35009/_0_  = ~n9987 ;
  assign \g35010/_0_  = ~n9990 ;
  assign \g35011/_0_  = ~n9993 ;
  assign \g35012/_0_  = ~n9996 ;
  assign \g35013/_0_  = ~n9999 ;
  assign \g35014/_0_  = ~n10002 ;
  assign \g35015/_0_  = ~n10005 ;
  assign \g35016/_0_  = ~n10008 ;
  assign \g35017/_0_  = ~n10011 ;
  assign \g35018/_0_  = ~n10014 ;
  assign \g35019/_0_  = ~n10017 ;
  assign \g35020/_0_  = ~n10020 ;
  assign \g35021/_0_  = ~n10023 ;
  assign \g35022/_0_  = ~n10026 ;
  assign \g35023/_0_  = ~n10029 ;
  assign \g35024/_0_  = ~n10032 ;
  assign \g35025/_0_  = ~n10035 ;
  assign \g35026/_0_  = ~n10038 ;
  assign \g35027/_0_  = ~n10041 ;
  assign \g35028/_0_  = ~n10044 ;
  assign \g35029/_0_  = ~n10047 ;
  assign \g35030/_0_  = ~n10050 ;
  assign \g35031/_0_  = ~n10053 ;
  assign \g35032/_0_  = ~n10056 ;
  assign \g35033/_0_  = ~n10059 ;
  assign \g35034/_0_  = ~n10062 ;
  assign \g35035/_0_  = ~n10065 ;
  assign \g35036/_0_  = ~n10068 ;
  assign \g35037/_0_  = ~n10071 ;
  assign \g35038/_0_  = ~n10074 ;
  assign \g35039/_0_  = ~n10077 ;
  assign \g35040/_0_  = ~n10080 ;
  assign \g35041/_0_  = ~n10083 ;
  assign \g35042/_0_  = ~n10086 ;
  assign \g35043/_0_  = ~n10089 ;
  assign \g35044/_0_  = ~n10092 ;
  assign \g35045/_0_  = ~n10095 ;
  assign \g35046/_0_  = ~n10098 ;
  assign \g35047/_0_  = ~n10101 ;
  assign \g35048/_0_  = ~n10104 ;
  assign \g35049/_0_  = ~n10107 ;
  assign \g35050/_0_  = ~n10110 ;
  assign \g35051/_0_  = ~n10113 ;
  assign \g35052/_0_  = ~n10116 ;
  assign \g35053/_0_  = ~n10119 ;
  assign \g35054/_0_  = ~n10122 ;
  assign \g35055/_0_  = ~n10125 ;
  assign \g35056/_0_  = ~n10128 ;
  assign \g35057/_0_  = ~n10131 ;
  assign \g35058/_0_  = ~n10134 ;
  assign \g35059/_0_  = ~n10137 ;
  assign \g35060/_0_  = ~n10140 ;
  assign \g35061/_0_  = ~n10143 ;
  assign \g35062/_0_  = ~n10146 ;
  assign \g35063/_0_  = ~n10149 ;
  assign \g35064/_0_  = ~n10152 ;
  assign \g35065/_0_  = ~n10155 ;
  assign \g35066/_0_  = ~n10158 ;
  assign \g35538/_0_  = ~n10159 ;
  assign \g35956/_0_  = n2421 ;
  assign \g36298/_1_  = n9800 ;
  assign \g36324/_0_  = n929 ;
  assign \g36375/_0_  = n2427 ;
  assign \g38269/_0_  = ~n10171 ;
  assign \g38473/_0_  = n10177 ;
  assign \g38501/_0_  = ~n10183 ;
  assign \g38569/_0_  = ~n10201 ;
  assign \g38629/_0_  = ~n10219 ;
  assign \g38721_dup/_3_  = ~n10225 ;
  assign \g38735/_0_  = ~n10243 ;
  assign \g38753/_0_  = n1142 ;
  assign \g38849/_3_  = ~n2205 ;
  assign \g39071/_0_  = ~n10237 ;
  assign \g39073/_0_  = n10231 ;
  assign \g39077/_0_  = n10195 ;
  assign \g39080/_0_  = ~n10192 ;
  assign \g39135/_0_  = ~n10213 ;
  assign \g39138/_0_  = n10207 ;
  assign \g39182/_0_  = n10249 ;
  assign \g39197/_3_  = n10165 ;
  assign \g39207/_3_  = n1122 ;
  assign \g39241/_0_  = n10263 ;
  assign \g39272/_0_  = ~n10275 ;
  assign \g39307/_0_  = n2257 ;
  assign \g39308/_0_  = ~n2245 ;
  assign \g39361/_0_  = ~n2294 ;
  assign \g39494/_0_  = n3640 ;
  assign \g39558/_0_  = ~n2403 ;
  assign \g39575/_0_  = ~n10269 ;
  assign \g39583/_0_  = ~n2366 ;
endmodule
