module top (\CM_rd0[0]_pad , \CM_rd0[10]_pad , \CM_rd0[11]_pad , \CM_rd0[12]_pad , \CM_rd0[13]_pad , \CM_rd0[14]_pad , \CM_rd0[15]_pad , \CM_rd0[16]_pad , \CM_rd0[17]_pad , \CM_rd0[18]_pad , \CM_rd0[19]_pad , \CM_rd0[1]_pad , \CM_rd0[20]_pad , \CM_rd0[21]_pad , \CM_rd0[22]_pad , \CM_rd0[23]_pad , \CM_rd0[2]_pad , \CM_rd0[3]_pad , \CM_rd0[4]_pad , \CM_rd0[5]_pad , \CM_rd0[6]_pad , \CM_rd0[7]_pad , \CM_rd0[8]_pad , \CM_rd0[9]_pad , \CM_rd1[0]_pad , \CM_rd1[10]_pad , \CM_rd1[11]_pad , \CM_rd1[12]_pad , \CM_rd1[13]_pad , \CM_rd1[14]_pad , \CM_rd1[15]_pad , \CM_rd1[16]_pad , \CM_rd1[17]_pad , \CM_rd1[18]_pad , \CM_rd1[19]_pad , \CM_rd1[1]_pad , \CM_rd1[20]_pad , \CM_rd1[21]_pad , \CM_rd1[22]_pad , \CM_rd1[23]_pad , \CM_rd1[2]_pad , \CM_rd1[3]_pad , \CM_rd1[4]_pad , \CM_rd1[5]_pad , \CM_rd1[6]_pad , \CM_rd1[7]_pad , \CM_rd1[8]_pad , \CM_rd1[9]_pad , \CM_rd2[0]_pad , \CM_rd2[10]_pad , \CM_rd2[11]_pad , \CM_rd2[12]_pad , \CM_rd2[13]_pad , \CM_rd2[14]_pad , \CM_rd2[15]_pad , \CM_rd2[16]_pad , \CM_rd2[17]_pad , \CM_rd2[18]_pad , \CM_rd2[19]_pad , \CM_rd2[1]_pad , \CM_rd2[20]_pad , \CM_rd2[21]_pad , \CM_rd2[22]_pad , \CM_rd2[23]_pad , \CM_rd2[2]_pad , \CM_rd2[3]_pad , \CM_rd2[4]_pad , \CM_rd2[5]_pad , \CM_rd2[6]_pad , \CM_rd2[7]_pad , \CM_rd2[8]_pad , \CM_rd2[9]_pad , \CM_rd3[0]_pad , \CM_rd3[10]_pad , \CM_rd3[11]_pad , \CM_rd3[12]_pad , \CM_rd3[13]_pad , \CM_rd3[14]_pad , \CM_rd3[15]_pad , \CM_rd3[16]_pad , \CM_rd3[17]_pad , \CM_rd3[18]_pad , \CM_rd3[19]_pad , \CM_rd3[1]_pad , \CM_rd3[20]_pad , \CM_rd3[21]_pad , \CM_rd3[22]_pad , \CM_rd3[23]_pad , \CM_rd3[2]_pad , \CM_rd3[3]_pad , \CM_rd3[4]_pad , \CM_rd3[5]_pad , \CM_rd3[6]_pad , \CM_rd3[7]_pad , \CM_rd3[8]_pad , \CM_rd3[9]_pad , \CM_rd4[0]_pad , \CM_rd4[10]_pad , \CM_rd4[11]_pad , \CM_rd4[12]_pad , \CM_rd4[13]_pad , \CM_rd4[14]_pad , \CM_rd4[15]_pad , \CM_rd4[16]_pad , \CM_rd4[17]_pad , \CM_rd4[18]_pad , \CM_rd4[19]_pad , \CM_rd4[1]_pad , \CM_rd4[20]_pad , \CM_rd4[21]_pad , \CM_rd4[22]_pad , \CM_rd4[23]_pad , \CM_rd4[2]_pad , \CM_rd4[3]_pad , \CM_rd4[4]_pad , \CM_rd4[5]_pad , \CM_rd4[6]_pad , \CM_rd4[7]_pad , \CM_rd4[8]_pad , \CM_rd4[9]_pad , \CM_rd5[0]_pad , \CM_rd5[10]_pad , \CM_rd5[11]_pad , \CM_rd5[12]_pad , \CM_rd5[13]_pad , \CM_rd5[14]_pad , \CM_rd5[15]_pad , \CM_rd5[16]_pad , \CM_rd5[17]_pad , \CM_rd5[18]_pad , \CM_rd5[19]_pad , \CM_rd5[1]_pad , \CM_rd5[20]_pad , \CM_rd5[21]_pad , \CM_rd5[22]_pad , \CM_rd5[23]_pad , \CM_rd5[2]_pad , \CM_rd5[3]_pad , \CM_rd5[4]_pad , \CM_rd5[5]_pad , \CM_rd5[6]_pad , \CM_rd5[7]_pad , \CM_rd5[8]_pad , \CM_rd5[9]_pad , \CM_rd6[0]_pad , \CM_rd6[10]_pad , \CM_rd6[11]_pad , \CM_rd6[12]_pad , \CM_rd6[13]_pad , \CM_rd6[14]_pad , \CM_rd6[15]_pad , \CM_rd6[16]_pad , \CM_rd6[17]_pad , \CM_rd6[18]_pad , \CM_rd6[19]_pad , \CM_rd6[1]_pad , \CM_rd6[20]_pad , \CM_rd6[21]_pad , \CM_rd6[22]_pad , \CM_rd6[23]_pad , \CM_rd6[2]_pad , \CM_rd6[3]_pad , \CM_rd6[4]_pad , \CM_rd6[5]_pad , \CM_rd6[6]_pad , \CM_rd6[7]_pad , \CM_rd6[8]_pad , \CM_rd6[9]_pad , \CM_rd7[0]_pad , \CM_rd7[10]_pad , \CM_rd7[11]_pad , \CM_rd7[12]_pad , \CM_rd7[13]_pad , \CM_rd7[14]_pad , \CM_rd7[15]_pad , \CM_rd7[16]_pad , \CM_rd7[17]_pad , \CM_rd7[18]_pad , \CM_rd7[19]_pad , \CM_rd7[1]_pad , \CM_rd7[20]_pad , \CM_rd7[21]_pad , \CM_rd7[22]_pad , \CM_rd7[23]_pad , \CM_rd7[2]_pad , \CM_rd7[3]_pad , \CM_rd7[4]_pad , \CM_rd7[5]_pad , \CM_rd7[6]_pad , \CM_rd7[7]_pad , \CM_rd7[8]_pad , \CM_rd7[9]_pad , \CM_rdm[0]_pad , \CM_rdm[10]_pad , \CM_rdm[11]_pad , \CM_rdm[12]_pad , \CM_rdm[13]_pad , \CM_rdm[14]_pad , \CM_rdm[15]_pad , \CM_rdm[16]_pad , \CM_rdm[17]_pad , \CM_rdm[18]_pad , \CM_rdm[19]_pad , \CM_rdm[1]_pad , \CM_rdm[20]_pad , \CM_rdm[21]_pad , \CM_rdm[22]_pad , \CM_rdm[23]_pad , \CM_rdm[2]_pad , \CM_rdm[3]_pad , \CM_rdm[4]_pad , \CM_rdm[5]_pad , \CM_rdm[6]_pad , \CM_rdm[7]_pad , \CM_rdm[8]_pad , \CM_rdm[9]_pad , \DM_rd0[0]_pad , \DM_rd0[10]_pad , \DM_rd0[11]_pad , \DM_rd0[12]_pad , \DM_rd0[13]_pad , \DM_rd0[14]_pad , \DM_rd0[15]_pad , \DM_rd0[1]_pad , \DM_rd0[2]_pad , \DM_rd0[3]_pad , \DM_rd0[4]_pad , \DM_rd0[5]_pad , \DM_rd0[6]_pad , \DM_rd0[7]_pad , \DM_rd0[8]_pad , \DM_rd0[9]_pad , \DM_rd1[0]_pad , \DM_rd1[10]_pad , \DM_rd1[11]_pad , \DM_rd1[12]_pad , \DM_rd1[13]_pad , \DM_rd1[14]_pad , \DM_rd1[15]_pad , \DM_rd1[1]_pad , \DM_rd1[2]_pad , \DM_rd1[3]_pad , \DM_rd1[4]_pad , \DM_rd1[5]_pad , \DM_rd1[6]_pad , \DM_rd1[7]_pad , \DM_rd1[8]_pad , \DM_rd1[9]_pad , \DM_rd2[0]_pad , \DM_rd2[10]_pad , \DM_rd2[11]_pad , \DM_rd2[12]_pad , \DM_rd2[13]_pad , \DM_rd2[14]_pad , \DM_rd2[15]_pad , \DM_rd2[1]_pad , \DM_rd2[2]_pad , \DM_rd2[3]_pad , \DM_rd2[4]_pad , \DM_rd2[5]_pad , \DM_rd2[6]_pad , \DM_rd2[7]_pad , \DM_rd2[8]_pad , \DM_rd2[9]_pad , \DM_rd3[0]_pad , \DM_rd3[10]_pad , \DM_rd3[11]_pad , \DM_rd3[12]_pad , \DM_rd3[13]_pad , \DM_rd3[14]_pad , \DM_rd3[15]_pad , \DM_rd3[1]_pad , \DM_rd3[2]_pad , \DM_rd3[3]_pad , \DM_rd3[4]_pad , \DM_rd3[5]_pad , \DM_rd3[6]_pad , \DM_rd3[7]_pad , \DM_rd3[8]_pad , \DM_rd3[9]_pad , \DM_rd4[0]_pad , \DM_rd4[10]_pad , \DM_rd4[11]_pad , \DM_rd4[12]_pad , \DM_rd4[13]_pad , \DM_rd4[14]_pad , \DM_rd4[15]_pad , \DM_rd4[1]_pad , \DM_rd4[2]_pad , \DM_rd4[3]_pad , \DM_rd4[4]_pad , \DM_rd4[5]_pad , \DM_rd4[6]_pad , \DM_rd4[7]_pad , \DM_rd4[8]_pad , \DM_rd4[9]_pad , \DM_rd5[0]_pad , \DM_rd5[10]_pad , \DM_rd5[11]_pad , \DM_rd5[12]_pad , \DM_rd5[13]_pad , \DM_rd5[14]_pad , \DM_rd5[15]_pad , \DM_rd5[1]_pad , \DM_rd5[2]_pad , \DM_rd5[3]_pad , \DM_rd5[4]_pad , \DM_rd5[5]_pad , \DM_rd5[6]_pad , \DM_rd5[7]_pad , \DM_rd5[8]_pad , \DM_rd5[9]_pad , \DM_rd6[0]_pad , \DM_rd6[10]_pad , \DM_rd6[11]_pad , \DM_rd6[12]_pad , \DM_rd6[13]_pad , \DM_rd6[14]_pad , \DM_rd6[15]_pad , \DM_rd6[1]_pad , \DM_rd6[2]_pad , \DM_rd6[3]_pad , \DM_rd6[4]_pad , \DM_rd6[5]_pad , \DM_rd6[6]_pad , \DM_rd6[7]_pad , \DM_rd6[8]_pad , \DM_rd6[9]_pad , \DM_rd7[0]_pad , \DM_rd7[10]_pad , \DM_rd7[11]_pad , \DM_rd7[12]_pad , \DM_rd7[13]_pad , \DM_rd7[14]_pad , \DM_rd7[15]_pad , \DM_rd7[1]_pad , \DM_rd7[2]_pad , \DM_rd7[3]_pad , \DM_rd7[4]_pad , \DM_rd7[5]_pad , \DM_rd7[6]_pad , \DM_rd7[7]_pad , \DM_rd7[8]_pad , \DM_rd7[9]_pad , \DM_rdm[0]_pad , \DM_rdm[10]_pad , \DM_rdm[11]_pad , \DM_rdm[12]_pad , \DM_rdm[13]_pad , \DM_rdm[14]_pad , \DM_rdm[15]_pad , \DM_rdm[1]_pad , \DM_rdm[2]_pad , \DM_rdm[3]_pad , \DM_rdm[4]_pad , \DM_rdm[5]_pad , \DM_rdm[6]_pad , \DM_rdm[7]_pad , \DM_rdm[8]_pad , \DM_rdm[9]_pad , IACKn_pad, \IRFS0_pad , \IRFS1_pad , \ISCLK0_pad , \ISCLK1_pad , \ITFS0_pad , \ITFS1_pad , \PIO_oe[0]_pad , \PIO_oe[10]_pad , \PIO_oe[11]_pad , \PIO_oe[1]_pad , \PIO_oe[2]_pad , \PIO_oe[3]_pad , \PIO_oe[4]_pad , \PIO_oe[5]_pad , \PIO_oe[6]_pad , \PIO_oe[7]_pad , \PIO_oe[8]_pad , \PIO_oe[9]_pad , \PIO_out[0]_pad , \PIO_out[10]_pad , \PIO_out[11]_pad , \PIO_out[1]_pad , \PIO_out[2]_pad , \PIO_out[3]_pad , \PIO_out[4]_pad , \PIO_out[5]_pad , \PIO_out[6]_pad , \PIO_out[7]_pad , \PIO_out[8]_pad , \PIO_out[9]_pad , PM_bdry_sel_pad, \PM_rd0[0]_pad , \PM_rd0[10]_pad , \PM_rd0[11]_pad , \PM_rd0[12]_pad , \PM_rd0[13]_pad , \PM_rd0[14]_pad , \PM_rd0[15]_pad , \PM_rd0[1]_pad , \PM_rd0[2]_pad , \PM_rd0[3]_pad , \PM_rd0[4]_pad , \PM_rd0[5]_pad , \PM_rd0[6]_pad , \PM_rd0[7]_pad , \PM_rd0[8]_pad , \PM_rd0[9]_pad , \PM_rd1[0]_pad , \PM_rd1[10]_pad , \PM_rd1[11]_pad , \PM_rd1[12]_pad , \PM_rd1[13]_pad , \PM_rd1[14]_pad , \PM_rd1[15]_pad , \PM_rd1[1]_pad , \PM_rd1[2]_pad , \PM_rd1[3]_pad , \PM_rd1[4]_pad , \PM_rd1[5]_pad , \PM_rd1[6]_pad , \PM_rd1[7]_pad , \PM_rd1[8]_pad , \PM_rd1[9]_pad , \PM_rd2[0]_pad , \PM_rd2[10]_pad , \PM_rd2[11]_pad , \PM_rd2[12]_pad , \PM_rd2[13]_pad , \PM_rd2[14]_pad , \PM_rd2[15]_pad , \PM_rd2[1]_pad , \PM_rd2[2]_pad , \PM_rd2[3]_pad , \PM_rd2[4]_pad , \PM_rd2[5]_pad , \PM_rd2[6]_pad , \PM_rd2[7]_pad , \PM_rd2[8]_pad , \PM_rd2[9]_pad , \PM_rd3[0]_pad , \PM_rd3[10]_pad , \PM_rd3[11]_pad , \PM_rd3[12]_pad , \PM_rd3[13]_pad , \PM_rd3[14]_pad , \PM_rd3[15]_pad , \PM_rd3[1]_pad , \PM_rd3[2]_pad , \PM_rd3[3]_pad , \PM_rd3[4]_pad , \PM_rd3[5]_pad , \PM_rd3[6]_pad , \PM_rd3[7]_pad , \PM_rd3[8]_pad , \PM_rd3[9]_pad , \PM_rd4[0]_pad , \PM_rd4[10]_pad , \PM_rd4[11]_pad , \PM_rd4[12]_pad , \PM_rd4[13]_pad , \PM_rd4[14]_pad , \PM_rd4[15]_pad , \PM_rd4[1]_pad , \PM_rd4[2]_pad , \PM_rd4[3]_pad , \PM_rd4[4]_pad , \PM_rd4[5]_pad , \PM_rd4[6]_pad , \PM_rd4[7]_pad , \PM_rd4[8]_pad , \PM_rd4[9]_pad , \PM_rd5[0]_pad , \PM_rd5[10]_pad , \PM_rd5[11]_pad , \PM_rd5[12]_pad , \PM_rd5[13]_pad , \PM_rd5[14]_pad , \PM_rd5[15]_pad , \PM_rd5[1]_pad , \PM_rd5[2]_pad , \PM_rd5[3]_pad , \PM_rd5[4]_pad , \PM_rd5[5]_pad , \PM_rd5[6]_pad , \PM_rd5[7]_pad , \PM_rd5[8]_pad , \PM_rd5[9]_pad , \PM_rd6[0]_pad , \PM_rd6[10]_pad , \PM_rd6[11]_pad , \PM_rd6[12]_pad , \PM_rd6[13]_pad , \PM_rd6[14]_pad , \PM_rd6[15]_pad , \PM_rd6[1]_pad , \PM_rd6[2]_pad , \PM_rd6[3]_pad , \PM_rd6[4]_pad , \PM_rd6[5]_pad , \PM_rd6[6]_pad , \PM_rd6[7]_pad , \PM_rd6[8]_pad , \PM_rd6[9]_pad , \PM_rd7[0]_pad , \PM_rd7[10]_pad , \PM_rd7[11]_pad , \PM_rd7[12]_pad , \PM_rd7[13]_pad , \PM_rd7[14]_pad , \PM_rd7[15]_pad , \PM_rd7[1]_pad , \PM_rd7[2]_pad , \PM_rd7[3]_pad , \PM_rd7[4]_pad , \PM_rd7[5]_pad , \PM_rd7[6]_pad , \PM_rd7[7]_pad , \PM_rd7[8]_pad , \PM_rd7[9]_pad , PWDACK_pad, T_BMODE_pad, T_BRn_pad, T_CLKI_OSC_pad, T_CLKI_PLL_pad, \T_ED[0]_pad , \T_ED[10]_pad , \T_ED[11]_pad , \T_ED[12]_pad , \T_ED[13]_pad , \T_ED[14]_pad , \T_ED[15]_pad , \T_ED[1]_pad , \T_ED[2]_pad , \T_ED[3]_pad , \T_ED[4]_pad , \T_ED[5]_pad , \T_ED[6]_pad , \T_ED[7]_pad , \T_ED[8]_pad , \T_ED[9]_pad , T_ICE_RSTn_pad, T_ID_pad, T_IMS_pad, T_IRDn_pad, \T_IRQ0n_pad , \T_IRQ1n_pad , \T_IRQ2n_pad , \T_IRQE0n_pad , \T_IRQE1n_pad , \T_IRQL1n_pad , T_ISn_pad, T_IWRn_pad, T_MMAP_pad, \T_PIOin[0]_pad , \T_PIOin[10]_pad , \T_PIOin[11]_pad , \T_PIOin[1]_pad , \T_PIOin[2]_pad , \T_PIOin[3]_pad , \T_PIOin[4]_pad , \T_PIOin[5]_pad , \T_PIOin[6]_pad , \T_PIOin[7]_pad , \T_PIOin[8]_pad , \T_PIOin[9]_pad , T_PWDn_pad, \T_RD0_pad , \T_RD1_pad , \T_RFS0_pad , \T_RFS1_pad , T_RSTn_pad, \T_SCLK0_pad , \T_SCLK1_pad , T_Sel_PLL_pad, \T_TFS0_pad , \T_TFS1_pad , \T_TMODE[0]_pad , \T_TMODE[1]_pad , \auctl_BSack_reg/NET0131 , \auctl_DSack_reg/NET0131 , \auctl_R0Sack_reg/NET0131 , \auctl_R1Sack_reg/NET0131 , \auctl_RST_reg/P0001 , \auctl_STEAL_reg/NET0131 , \auctl_T0Sack_reg/NET0131 , \auctl_T1Sack_reg/NET0131 , \bdma_BCTL_reg[0]/NET0131 , \bdma_BCTL_reg[10]/NET0131 , \bdma_BCTL_reg[11]/NET0131 , \bdma_BCTL_reg[12]/NET0131 , \bdma_BCTL_reg[13]/NET0131 , \bdma_BCTL_reg[14]/NET0131 , \bdma_BCTL_reg[15]/NET0131 , \bdma_BCTL_reg[1]/NET0131 , \bdma_BCTL_reg[2]/NET0131 , \bdma_BCTL_reg[3]/NET0131 , \bdma_BCTL_reg[4]/NET0131 , \bdma_BCTL_reg[5]/NET0131 , \bdma_BCTL_reg[6]/NET0131 , \bdma_BCTL_reg[7]/NET0131 , \bdma_BCTL_reg[8]/NET0131 , \bdma_BCTL_reg[9]/NET0131 , \bdma_BDMA_boot_reg/NET0131_reg_syn_10 , \bdma_BDMA_boot_reg/NET0131_reg_syn_2 , \bdma_BDMA_boot_reg/NET0131_reg_syn_8 , \bdma_BDMAmode_reg/NET0131 , \bdma_BEAD_reg[0]/NET0131 , \bdma_BEAD_reg[10]/NET0131 , \bdma_BEAD_reg[11]/NET0131 , \bdma_BEAD_reg[12]/NET0131 , \bdma_BEAD_reg[13]/NET0131 , \bdma_BEAD_reg[1]/NET0131 , \bdma_BEAD_reg[2]/NET0131 , \bdma_BEAD_reg[3]/NET0131 , \bdma_BEAD_reg[4]/NET0131 , \bdma_BEAD_reg[5]/NET0131 , \bdma_BEAD_reg[6]/NET0131 , \bdma_BEAD_reg[7]/NET0131 , \bdma_BEAD_reg[8]/NET0131 , \bdma_BEAD_reg[9]/NET0131 , \bdma_BIAD_reg[0]/NET0131 , \bdma_BIAD_reg[10]/NET0131 , \bdma_BIAD_reg[11]/NET0131 , \bdma_BIAD_reg[12]/NET0131 , \bdma_BIAD_reg[13]/NET0131 , \bdma_BIAD_reg[1]/NET0131 , \bdma_BIAD_reg[2]/NET0131 , \bdma_BIAD_reg[3]/NET0131 , \bdma_BIAD_reg[4]/NET0131 , \bdma_BIAD_reg[5]/NET0131 , \bdma_BIAD_reg[6]/NET0131 , \bdma_BIAD_reg[7]/NET0131 , \bdma_BIAD_reg[8]/NET0131 , \bdma_BIAD_reg[9]/NET0131 , \bdma_BM_cyc_reg/P0001 , \bdma_BMcyc_del_reg/P0001 , \bdma_BOVL_reg[0]/NET0131 , \bdma_BOVL_reg[10]/NET0131 , \bdma_BOVL_reg[11]/NET0131 , \bdma_BOVL_reg[1]/NET0131 , \bdma_BOVL_reg[2]/NET0131 , \bdma_BOVL_reg[3]/NET0131 , \bdma_BOVL_reg[4]/NET0131 , \bdma_BOVL_reg[5]/NET0131 , \bdma_BOVL_reg[6]/NET0131 , \bdma_BOVL_reg[7]/NET0131 , \bdma_BOVL_reg[8]/NET0131 , \bdma_BOVL_reg[9]/NET0131 , \bdma_BRST_s2_reg/NET0131 , \bdma_BRdataBUF_reg[0]/P0001 , \bdma_BRdataBUF_reg[10]/P0001 , \bdma_BRdataBUF_reg[11]/P0001 , \bdma_BRdataBUF_reg[12]/P0001 , \bdma_BRdataBUF_reg[13]/P0001 , \bdma_BRdataBUF_reg[14]/P0001 , \bdma_BRdataBUF_reg[15]/P0001 , \bdma_BRdataBUF_reg[16]/P0001 , \bdma_BRdataBUF_reg[17]/P0001 , \bdma_BRdataBUF_reg[18]/P0001 , \bdma_BRdataBUF_reg[19]/P0001 , \bdma_BRdataBUF_reg[1]/P0001 , \bdma_BRdataBUF_reg[20]/P0001 , \bdma_BRdataBUF_reg[21]/P0001 , \bdma_BRdataBUF_reg[22]/P0001 , \bdma_BRdataBUF_reg[23]/P0001 , \bdma_BRdataBUF_reg[2]/P0001 , \bdma_BRdataBUF_reg[3]/P0001 , \bdma_BRdataBUF_reg[4]/P0001 , \bdma_BRdataBUF_reg[5]/P0001 , \bdma_BRdataBUF_reg[6]/P0001 , \bdma_BRdataBUF_reg[7]/P0001 , \bdma_BRdataBUF_reg[8]/P0001 , \bdma_BRdataBUF_reg[9]/P0001 , \bdma_BSreq_reg/NET0131 , \bdma_BWCOUNT_reg[0]/NET0131 , \bdma_BWCOUNT_reg[10]/NET0131 , \bdma_BWCOUNT_reg[11]/NET0131 , \bdma_BWCOUNT_reg[12]/NET0131 , \bdma_BWCOUNT_reg[13]/NET0131 , \bdma_BWCOUNT_reg[1]/NET0131 , \bdma_BWCOUNT_reg[2]/NET0131 , \bdma_BWCOUNT_reg[3]/NET0131 , \bdma_BWCOUNT_reg[4]/NET0131 , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2 , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8 , \bdma_BWCOUNT_reg[6]/NET0131 , \bdma_BWCOUNT_reg[7]/NET0131 , \bdma_BWCOUNT_reg[8]/NET0131 , \bdma_BWCOUNT_reg[9]/NET0131 , \bdma_BWRn_reg/NET0131 , \bdma_BWcnt_reg[0]/NET0131 , \bdma_BWcnt_reg[1]/NET0131 , \bdma_BWcnt_reg[2]/NET0131 , \bdma_BWcnt_reg[3]/NET0131 , \bdma_BWcnt_reg[4]/NET0131 , \bdma_BWdataBUF_h_reg[0]/P0001 , \bdma_BWdataBUF_h_reg[10]/P0001 , \bdma_BWdataBUF_h_reg[11]/P0001 , \bdma_BWdataBUF_h_reg[12]/P0001 , \bdma_BWdataBUF_h_reg[13]/P0001 , \bdma_BWdataBUF_h_reg[14]/P0001 , \bdma_BWdataBUF_h_reg[15]/P0001 , \bdma_BWdataBUF_h_reg[16]/P0001 , \bdma_BWdataBUF_h_reg[17]/P0001 , \bdma_BWdataBUF_h_reg[18]/P0001 , \bdma_BWdataBUF_h_reg[19]/P0001 , \bdma_BWdataBUF_h_reg[1]/P0001 , \bdma_BWdataBUF_h_reg[20]/P0001 , \bdma_BWdataBUF_h_reg[21]/P0001 , \bdma_BWdataBUF_h_reg[22]/P0001 , \bdma_BWdataBUF_h_reg[23]/P0001 , \bdma_BWdataBUF_h_reg[2]/P0001 , \bdma_BWdataBUF_h_reg[3]/P0001 , \bdma_BWdataBUF_h_reg[4]/P0001 , \bdma_BWdataBUF_h_reg[5]/P0001 , \bdma_BWdataBUF_h_reg[6]/P0001 , \bdma_BWdataBUF_h_reg[7]/P0001 , \bdma_BWdataBUF_h_reg[8]/P0001 , \bdma_BWdataBUF_h_reg[9]/P0001 , \bdma_BWdataBUF_reg[0]/P0001 , \bdma_BWdataBUF_reg[1]/P0001 , \bdma_BWdataBUF_reg[2]/P0001 , \bdma_BWdataBUF_reg[3]/P0001 , \bdma_BWdataBUF_reg[4]/P0001 , \bdma_BWdataBUF_reg[5]/P0001 , \bdma_BWdataBUF_reg[6]/P0001 , \bdma_BWdataBUF_reg[7]/P0001 , \bdma_CMcnt_reg[0]/NET0131 , \bdma_CMcnt_reg[1]/NET0131 , \bdma_DM_2nd_reg/NET0131 , \bdma_RST_pin_reg/P0001 , \bdma_WRlat_reg/P0001 , \clkc_Awake_reg/NET0131 , \clkc_CLKOUT_reg/NET0131 , \clkc_CTR_cnt_reg[0]/NET0131 , \clkc_CTR_cnt_reg[1]/NET0131 , \clkc_Cnt128_reg/NET0131 , \clkc_Cnt4096_reg/NET0131 , \clkc_Cnt4096_s1_reg/NET0131 , \clkc_Cnt4096_s2_reg/NET0131 , \clkc_DSPoff_reg/NET0131 , \clkc_OSCoff_reg/NET0131 , \clkc_OSCoff_set_reg/P0001 , \clkc_OUTcnt_reg[0]/NET0131 , \clkc_OUTcnt_reg[1]/NET0131 , \clkc_OUTcnt_reg[2]/NET0131 , \clkc_OUTcnt_reg[3]/NET0131 , \clkc_OUTcnt_reg[4]/NET0131 , \clkc_OUTcnt_reg[5]/NET0131 , \clkc_OUTcnt_reg[6]/NET0131 , \clkc_RSTtext_reg/P0001 , \clkc_SIDLE_s1_reg/NET0131 , \clkc_SIDLE_s2_reg/NET0131 , \clkc_SLEEP_reg/NET0131 , \clkc_STBY_reg/NET0131 , \clkc_STDcnt_reg[0]/NET0131 , \clkc_STDcnt_reg[10]/NET0131 , \clkc_STDcnt_reg[1]/NET0131 , \clkc_STDcnt_reg[2]/NET0131 , \clkc_STDcnt_reg[3]/NET0131 , \clkc_STDcnt_reg[4]/NET0131 , \clkc_STDcnt_reg[5]/NET0131 , \clkc_STDcnt_reg[6]/NET0131 , \clkc_STDcnt_reg[7]/NET0131 , \clkc_STDcnt_reg[8]/NET0131 , \clkc_STDcnt_reg[9]/NET0131 , \clkc_SlowDn_reg/NET0131 , \clkc_SlowDn_s1_reg/P0001 , \clkc_SlowDn_s2_reg/P0001 , \clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131 , \clkc_ckr_reg_DO_reg[0]/NET0131 , \clkc_ckr_reg_DO_reg[10]/NET0131 , \clkc_ckr_reg_DO_reg[11]/NET0131 , \clkc_ckr_reg_DO_reg[12]/NET0131 , \clkc_ckr_reg_DO_reg[13]/NET0131 , \clkc_ckr_reg_DO_reg[14]/NET0131 , \clkc_ckr_reg_DO_reg[15]/NET0131 , \clkc_ckr_reg_DO_reg[1]/NET0131 , \clkc_ckr_reg_DO_reg[2]/NET0131 , \clkc_ckr_reg_DO_reg[3]/NET0131 , \clkc_ckr_reg_DO_reg[4]/NET0131 , \clkc_ckr_reg_DO_reg[5]/NET0131 , \clkc_ckr_reg_DO_reg[6]/NET0131 , \clkc_ckr_reg_DO_reg[7]/NET0131 , \clkc_ckr_reg_DO_reg[8]/NET0131 , \clkc_ckr_reg_DO_reg[9]/NET0131 , \clkc_oscntr_reg_DO_reg[0]/NET0131 , \clkc_oscntr_reg_DO_reg[10]/NET0131 , \clkc_oscntr_reg_DO_reg[11]/NET0131 , \clkc_oscntr_reg_DO_reg[1]/NET0131 , \clkc_oscntr_reg_DO_reg[2]/NET0131 , \clkc_oscntr_reg_DO_reg[3]/NET0131 , \clkc_oscntr_reg_DO_reg[4]/NET0131 , \clkc_oscntr_reg_DO_reg[5]/NET0131 , \clkc_oscntr_reg_DO_reg[6]/NET0131 , \clkc_oscntr_reg_DO_reg[7]/NET0131 , \clkc_oscntr_reg_DO_reg[8]/NET0131 , \clkc_oscntr_reg_DO_reg[9]/NET0131 , \core_c_dec_ALUop_E_reg/P0001 , \core_c_dec_BR_Ed_reg/P0001 , \core_c_dec_Call_Ed_reg/P0001 , \core_c_dec_DIVQ_E_reg/P0001 , \core_c_dec_DIVS_E_reg/P0001 , \core_c_dec_DU_Eg_reg/P0001 , \core_c_dec_Double_E_reg/P0001 , \core_c_dec_Dummy_E_reg/NET0131 , \core_c_dec_EXIT_E_reg/P0001 , \core_c_dec_IDLE_Eg_reg/P0001 , \core_c_dec_IRE_reg[0]/NET0131 , \core_c_dec_IRE_reg[10]/NET0131 , \core_c_dec_IRE_reg[11]/NET0131 , \core_c_dec_IRE_reg[12]/NET0131 , \core_c_dec_IRE_reg[13]/NET0131 , \core_c_dec_IRE_reg[14]/NET0131 , \core_c_dec_IRE_reg[15]/NET0131 , \core_c_dec_IRE_reg[16]/NET0131 , \core_c_dec_IRE_reg[17]/NET0131 , \core_c_dec_IRE_reg[18]/NET0131 , \core_c_dec_IRE_reg[19]/NET0131 , \core_c_dec_IRE_reg[1]/NET0131 , \core_c_dec_IRE_reg[2]/NET0131 , \core_c_dec_IRE_reg[3]/NET0131 , \core_c_dec_IRE_reg[4]/NET0131 , \core_c_dec_IRE_reg[5]/NET0131 , \core_c_dec_IRE_reg[6]/NET0131 , \core_c_dec_IRE_reg[7]/NET0131 , \core_c_dec_IRE_reg[8]/NET0131 , \core_c_dec_IRE_reg[9]/NET0131 , \core_c_dec_IR_reg[0]/NET0131 , \core_c_dec_IR_reg[10]/NET0131 , \core_c_dec_IR_reg[11]/NET0131 , \core_c_dec_IR_reg[12]/NET0131 , \core_c_dec_IR_reg[13]/NET0131 , \core_c_dec_IR_reg[14]/NET0131 , \core_c_dec_IR_reg[15]/NET0131 , \core_c_dec_IR_reg[16]/NET0131 , \core_c_dec_IR_reg[17]/NET0131 , \core_c_dec_IR_reg[18]/NET0131 , \core_c_dec_IR_reg[19]/NET0131 , \core_c_dec_IR_reg[1]/NET0131 , \core_c_dec_IR_reg[20]/NET0131 , \core_c_dec_IR_reg[21]/NET0131 , \core_c_dec_IR_reg[22]/NET0131 , \core_c_dec_IR_reg[23]/NET0131 , \core_c_dec_IR_reg[2]/NET0131 , \core_c_dec_IR_reg[3]/NET0131 , \core_c_dec_IR_reg[4]/NET0131 , \core_c_dec_IR_reg[5]/NET0131 , \core_c_dec_IR_reg[6]/NET0131 , \core_c_dec_IR_reg[7]/NET0131 , \core_c_dec_IR_reg[8]/NET0131 , \core_c_dec_IR_reg[9]/NET0131 , \core_c_dec_Long_Cg_reg/P0001 , \core_c_dec_Long_Eg_reg/P0001 , \core_c_dec_MACdep_Eg_reg/P0001 , \core_c_dec_MACop_E_reg/P0001 , \core_c_dec_MFALU_Ei_reg/NET0131 , \core_c_dec_MFAR_E_reg/P0001 , \core_c_dec_MFASTAT_E_reg/P0001 , \core_c_dec_MFAX0_E_reg/P0001 , \core_c_dec_MFAX1_E_reg/P0001 , \core_c_dec_MFAY0_E_reg/P0001 , \core_c_dec_MFAY1_E_reg/P0001 , \core_c_dec_MFCNTR_E_reg/P0001 , \core_c_dec_MFDAG1_Ei_reg/NET0131 , \core_c_dec_MFDAG2_Ei_reg/NET0131 , \core_c_dec_MFDMOVL_E_reg/P0001 , \core_c_dec_MFICNTL_E_reg/P0001 , \core_c_dec_MFIDR_E_reg/P0001 , \core_c_dec_MFIMASK_E_reg/P0001 , \core_c_dec_MFIreg_E_reg[0]/P0001 , \core_c_dec_MFIreg_E_reg[1]/P0001 , \core_c_dec_MFIreg_E_reg[2]/P0001 , \core_c_dec_MFIreg_E_reg[3]/P0001 , \core_c_dec_MFIreg_E_reg[4]/P0001 , \core_c_dec_MFIreg_E_reg[5]/P0001 , \core_c_dec_MFIreg_E_reg[6]/P0001 , \core_c_dec_MFIreg_E_reg[7]/P0001 , \core_c_dec_MFLreg_E_reg[0]/P0001 , \core_c_dec_MFLreg_E_reg[1]/P0001 , \core_c_dec_MFLreg_E_reg[2]/P0001 , \core_c_dec_MFLreg_E_reg[3]/P0001 , \core_c_dec_MFLreg_E_reg[4]/P0001 , \core_c_dec_MFLreg_E_reg[5]/P0001 , \core_c_dec_MFLreg_E_reg[6]/P0001 , \core_c_dec_MFLreg_E_reg[7]/P0001 , \core_c_dec_MFMAC_Ei_reg/NET0131 , \core_c_dec_MFMR0_E_reg/P0001 , \core_c_dec_MFMR1_E_reg/P0001 , \core_c_dec_MFMR2_E_reg/P0001 , \core_c_dec_MFMSTAT_E_reg/P0001 , \core_c_dec_MFMX0_E_reg/P0001 , \core_c_dec_MFMX1_E_reg/P0001 , \core_c_dec_MFMY0_E_reg/P0001 , \core_c_dec_MFMY1_E_reg/P0001 , \core_c_dec_MFMreg_E_reg[0]/P0001 , \core_c_dec_MFMreg_E_reg[1]/P0001 , \core_c_dec_MFMreg_E_reg[2]/P0001 , \core_c_dec_MFMreg_E_reg[3]/P0001 , \core_c_dec_MFMreg_E_reg[4]/P0001 , \core_c_dec_MFMreg_E_reg[5]/P0001 , \core_c_dec_MFMreg_E_reg[6]/P0001 , \core_c_dec_MFMreg_E_reg[7]/P0001 , \core_c_dec_MFPMOVL_E_reg/P0001 , \core_c_dec_MFPSQ_Ei_reg/NET0131 , \core_c_dec_MFRX0_E_reg/P0001 , \core_c_dec_MFRX1_E_reg/P0001 , \core_c_dec_MFSB_E_reg/P0001 , \core_c_dec_MFSE_E_reg/P0001 , \core_c_dec_MFSHT_Ei_reg/NET0131 , \core_c_dec_MFSI_E_reg/P0001 , \core_c_dec_MFSPT_Ei_reg/NET0131 , \core_c_dec_MFSR0_E_reg/P0001 , \core_c_dec_MFSR1_E_reg/P0001 , \core_c_dec_MFSSTAT_E_reg/P0001 , \core_c_dec_MFTX0_E_reg/P0001 , \core_c_dec_MFTX1_E_reg/P0001 , \core_c_dec_MFtoppcs_Eg_reg/P0001 , \core_c_dec_MTAR_E_reg/P0001 , \core_c_dec_MTASTAT_E_reg/P0001 , \core_c_dec_MTAX0_E_reg/P0001 , \core_c_dec_MTAX1_E_reg/P0001 , \core_c_dec_MTAY0_E_reg/P0001 , \core_c_dec_MTAY1_E_reg/P0001 , \core_c_dec_MTCNTR_Eg_reg/P0001 , \core_c_dec_MTDMOVL_E_reg/P0001 , \core_c_dec_MTICNTL_Eg_reg/P0001 , \core_c_dec_MTIDR_E_reg/P0001 , \core_c_dec_MTIFC_Eg_reg/P0001 , \core_c_dec_MTIMASK_Eg_reg/P0001 , \core_c_dec_MTIreg_E_reg[0]/P0001 , \core_c_dec_MTIreg_E_reg[1]/P0001 , \core_c_dec_MTIreg_E_reg[2]/P0001 , \core_c_dec_MTIreg_E_reg[3]/P0001 , \core_c_dec_MTIreg_E_reg[4]/P0001 , \core_c_dec_MTIreg_E_reg[5]/P0001 , \core_c_dec_MTIreg_E_reg[6]/P0001 , \core_c_dec_MTIreg_E_reg[7]/P0001 , \core_c_dec_MTLreg_E_reg[0]/P0001 , \core_c_dec_MTLreg_E_reg[1]/P0001 , \core_c_dec_MTLreg_E_reg[2]/P0001 , \core_c_dec_MTLreg_E_reg[3]/P0001 , \core_c_dec_MTLreg_E_reg[4]/P0001 , \core_c_dec_MTLreg_E_reg[5]/P0001 , \core_c_dec_MTLreg_E_reg[6]/P0001 , \core_c_dec_MTLreg_E_reg[7]/P0001 , \core_c_dec_MTMR0_E_reg/P0001 , \core_c_dec_MTMR1_E_reg/P0001 , \core_c_dec_MTMR2_E_reg/P0001 , \core_c_dec_MTMSTAT_Eg_reg/P0001 , \core_c_dec_MTMX0_E_reg/P0001 , \core_c_dec_MTMX1_E_reg/P0001 , \core_c_dec_MTMY0_E_reg/P0001 , \core_c_dec_MTMY1_E_reg/P0001 , \core_c_dec_MTMreg_E_reg[0]/P0001 , \core_c_dec_MTMreg_E_reg[1]/P0001 , \core_c_dec_MTMreg_E_reg[2]/P0001 , \core_c_dec_MTMreg_E_reg[3]/P0001 , \core_c_dec_MTMreg_E_reg[4]/P0001 , \core_c_dec_MTMreg_E_reg[5]/P0001 , \core_c_dec_MTMreg_E_reg[6]/P0001 , \core_c_dec_MTMreg_E_reg[7]/P0001 , \core_c_dec_MTOWRCNTR_Eg_reg/P0001 , \core_c_dec_MTPMOVL_E_reg/P0001 , \core_c_dec_MTRX0_E_reg/P0001 , \core_c_dec_MTRX1_E_reg/P0001 , \core_c_dec_MTSB_E_reg/P0001 , \core_c_dec_MTSE_E_reg/P0001 , \core_c_dec_MTSI_E_reg/P0001 , \core_c_dec_MTSR0_E_reg/P0001 , \core_c_dec_MTSR1_E_reg/P0001 , \core_c_dec_MTTX0_E_reg/P0001 , \core_c_dec_MTTX1_E_reg/P0001 , \core_c_dec_MTtoppcs_Eg_reg/P0001 , \core_c_dec_Modctl_Eg_reg/P0001 , \core_c_dec_MpopLP_Eg_reg/P0001 , \core_c_dec_NOP_E_reg/P0001 , \core_c_dec_Nrti_Ed_reg/P0001 , \core_c_dec_Nseq_Ed_reg/P0001 , \core_c_dec_PPclr_reg/P0001 , \core_c_dec_Post1_E_reg/P0001 , \core_c_dec_Post2_E_reg/P0001 , \core_c_dec_Prderr_Cg_reg/NET0131 , \core_c_dec_RET_Ed_reg/P0001 , \core_c_dec_RTI_Ed_reg/P0001 , \core_c_dec_SHTop_E_reg/P0001 , \core_c_dec_Stkctl_Eg_reg/P0001 , \core_c_dec_Usecond_E_reg/P0001 , \core_c_dec_accCM_E_reg/NET0131 , \core_c_dec_accPM_E_reg/P0001 , \core_c_dec_cdAM_E_reg/P0001 , \core_c_dec_imSHT_E_reg/P0001 , \core_c_dec_imm14_E_reg/P0001 , \core_c_dec_imm16_E_reg/P0001 , \core_c_dec_pMFALU_Ei_reg/NET0131 , \core_c_dec_pMFMAC_Ei_reg/NET0131 , \core_c_dec_pMFSHT_Ei_reg/NET0131 , \core_c_dec_rdCM_E_reg/NET0131 , \core_c_dec_satMR_E_reg/P0001 , \core_c_dec_updAF_E_reg/P0001 , \core_c_dec_updAR_E_reg/P0001 , \core_c_dec_updMF_E_reg/P0001 , \core_c_dec_updMR_E_reg/P0001 , \core_c_dec_updSR_E_reg/P0001 , \core_c_psq_CE_reg/NET0131 , \core_c_psq_CNTR_reg_DO_reg[0]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[10]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[11]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[12]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[13]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[1]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[2]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[3]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[4]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[5]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[6]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[7]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[8]/NET0131 , \core_c_psq_CNTR_reg_DO_reg[9]/NET0131 , \core_c_psq_CNTRval_reg/NET0131 , \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 , \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 , \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 , \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 , \core_c_psq_DRA_reg[0]/P0001 , \core_c_psq_DRA_reg[10]/P0001 , \core_c_psq_DRA_reg[11]/P0001 , \core_c_psq_DRA_reg[12]/P0001 , \core_c_psq_DRA_reg[13]/P0001 , \core_c_psq_DRA_reg[1]/P0001 , \core_c_psq_DRA_reg[2]/P0001 , \core_c_psq_DRA_reg[3]/P0001 , \core_c_psq_DRA_reg[4]/P0001 , \core_c_psq_DRA_reg[5]/P0001 , \core_c_psq_DRA_reg[6]/P0001 , \core_c_psq_DRA_reg[7]/P0001 , \core_c_psq_DRA_reg[8]/P0001 , \core_c_psq_DRA_reg[9]/P0001 , \core_c_psq_ECYC_reg/P0001 , \core_c_psq_EXA_reg[0]/P0001 , \core_c_psq_EXA_reg[10]/P0001 , \core_c_psq_EXA_reg[11]/P0001 , \core_c_psq_EXA_reg[12]/P0001 , \core_c_psq_EXA_reg[13]/P0001 , \core_c_psq_EXA_reg[1]/P0001 , \core_c_psq_EXA_reg[2]/P0001 , \core_c_psq_EXA_reg[3]/P0001 , \core_c_psq_EXA_reg[4]/P0001 , \core_c_psq_EXA_reg[5]/P0001 , \core_c_psq_EXA_reg[6]/P0001 , \core_c_psq_EXA_reg[7]/P0001 , \core_c_psq_EXA_reg[8]/P0001 , \core_c_psq_EXA_reg[9]/P0001 , \core_c_psq_Eqend_D_reg/P0001 , \core_c_psq_Eqend_Ed_reg/P0001 , \core_c_psq_ICNTL_reg_DO_reg[0]/NET0131 , \core_c_psq_ICNTL_reg_DO_reg[1]/NET0131 , \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 , \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 , \core_c_psq_IFA_reg[0]/P0001 , \core_c_psq_IFA_reg[10]/P0001 , \core_c_psq_IFA_reg[11]/P0001 , \core_c_psq_IFA_reg[12]/P0001 , \core_c_psq_IFA_reg[13]/P0001 , \core_c_psq_IFA_reg[1]/P0001 , \core_c_psq_IFA_reg[2]/P0001 , \core_c_psq_IFA_reg[3]/P0001 , \core_c_psq_IFA_reg[4]/P0001 , \core_c_psq_IFA_reg[5]/P0001 , \core_c_psq_IFA_reg[6]/P0001 , \core_c_psq_IFA_reg[7]/P0001 , \core_c_psq_IFA_reg[8]/P0001 , \core_c_psq_IFA_reg[9]/P0001 , \core_c_psq_IFC_reg[0]/NET0131 , \core_c_psq_IFC_reg[10]/NET0131 , \core_c_psq_IFC_reg[11]/NET0131 , \core_c_psq_IFC_reg[12]/NET0131 , \core_c_psq_IFC_reg[13]/NET0131 , \core_c_psq_IFC_reg[14]/NET0131 , \core_c_psq_IFC_reg[15]/NET0131 , \core_c_psq_IFC_reg[1]/NET0131 , \core_c_psq_IFC_reg[2]/NET0131 , \core_c_psq_IFC_reg[3]/NET0131 , \core_c_psq_IFC_reg[4]/NET0131 , \core_c_psq_IFC_reg[5]/NET0131 , \core_c_psq_IFC_reg[6]/NET0131 , \core_c_psq_IFC_reg[7]/NET0131 , \core_c_psq_IFC_reg[8]/NET0131 , \core_c_psq_IFC_reg[9]/NET0131 , \core_c_psq_IMASK_reg[0]/NET0131 , \core_c_psq_IMASK_reg[1]/NET0131 , \core_c_psq_IMASK_reg[2]/NET0131 , \core_c_psq_IMASK_reg[3]/NET0131 , \core_c_psq_IMASK_reg[4]/NET0131 , \core_c_psq_IMASK_reg[5]/NET0131 , \core_c_psq_IMASK_reg[6]/NET0131 , \core_c_psq_IMASK_reg[7]/NET0131 , \core_c_psq_IMASK_reg[8]/NET0131 , \core_c_psq_IMASK_reg[9]/NET0131 , \core_c_psq_INT_en_reg/NET0131 , \core_c_psq_Iact_E_reg[0]/NET0131 , \core_c_psq_Iact_E_reg[10]/NET0131 , \core_c_psq_Iact_E_reg[1]/NET0131 , \core_c_psq_Iact_E_reg[2]/NET0131 , \core_c_psq_Iact_E_reg[3]/NET0131 , \core_c_psq_Iact_E_reg[4]/NET0131 , \core_c_psq_Iact_E_reg[5]/NET0131 , \core_c_psq_Iact_E_reg[6]/NET0131 , \core_c_psq_Iact_E_reg[7]/NET0131 , \core_c_psq_Iact_E_reg[8]/NET0131 , \core_c_psq_Iact_E_reg[9]/NET0131 , \core_c_psq_Iflag_reg[0]/NET0131 , \core_c_psq_Iflag_reg[10]/NET0131 , \core_c_psq_Iflag_reg[11]/NET0131 , \core_c_psq_Iflag_reg[12]/NET0131 , \core_c_psq_Iflag_reg[1]/NET0131 , \core_c_psq_Iflag_reg[2]/NET0131 , \core_c_psq_Iflag_reg[3]/NET0131 , \core_c_psq_Iflag_reg[4]/NET0131 , \core_c_psq_Iflag_reg[5]/NET0131 , \core_c_psq_Iflag_reg[6]/NET0131 , \core_c_psq_Iflag_reg[7]/NET0131 , \core_c_psq_Iflag_reg[8]/NET0131 , \core_c_psq_Iflag_reg[9]/NET0131 , \core_c_psq_MGNT_reg/NET0131 , \core_c_psq_MREQ_reg/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[0]/P0002 , \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 , \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 , \core_c_psq_PCS2or3_reg/NET0131 , \core_c_psq_PCS_reg[0]/NET0131 , \core_c_psq_PCS_reg[10]/NET0131 , \core_c_psq_PCS_reg[11]/NET0131 , \core_c_psq_PCS_reg[12]/NET0131 , \core_c_psq_PCS_reg[13]/NET0131 , \core_c_psq_PCS_reg[14]/NET0131 , \core_c_psq_PCS_reg[15]/NET0131 , \core_c_psq_PCS_reg[1]/NET0131 , \core_c_psq_PCS_reg[2]/NET0131 , \core_c_psq_PCS_reg[3]/NET0131 , \core_c_psq_PCS_reg[4]/NET0131 , \core_c_psq_PCS_reg[5]/NET0131 , \core_c_psq_PCS_reg[6]/NET0131 , \core_c_psq_PCS_reg[7]/NET0131 , \core_c_psq_PCS_reg[8]/NET0131 , \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 , \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 , \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 , \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 , \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 , \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 , \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 , \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 , \core_c_psq_SRST_reg/P0001 , \core_c_psq_SSTAT_reg[0]/NET0131 , \core_c_psq_SSTAT_reg[1]/NET0131 , \core_c_psq_SSTAT_reg[2]/NET0131 , \core_c_psq_SSTAT_reg[3]/NET0131 , \core_c_psq_SSTAT_reg[4]/NET0131 , \core_c_psq_SSTAT_reg[5]/NET0131 , \core_c_psq_SSTAT_reg[6]/NET0131 , \core_c_psq_SSTAT_reg[7]/NET0131 , \core_c_psq_TRAP_Eg_reg/NET0131 , \core_c_psq_TRAP_R_L_reg/NET0131 , \core_c_psq_T_IRQ0_s1_reg/P0001 , \core_c_psq_T_IRQ0p_reg/P0001 , \core_c_psq_T_IRQ1_s1_reg/P0001 , \core_c_psq_T_IRQ1p_reg/P0001 , \core_c_psq_T_IRQ2_s1_reg/P0001 , \core_c_psq_T_IRQ2p_reg/P0001 , \core_c_psq_T_IRQE0_reg/P0001 , \core_c_psq_T_IRQE0_s1_reg/P0001 , \core_c_psq_T_IRQE1_reg/P0001 , \core_c_psq_T_IRQE1_s1_reg/P0001 , \core_c_psq_T_IRQL0p_reg/P0001 , \core_c_psq_T_IRQL1p_reg/P0001 , \core_c_psq_T_PWRDN_reg/P0001 , \core_c_psq_T_PWRDN_s1_reg/P0001 , \core_c_psq_Taddr_Eb_reg[0]/P0001 , \core_c_psq_Taddr_Eb_reg[10]/P0001 , \core_c_psq_Taddr_Eb_reg[11]/P0001 , \core_c_psq_Taddr_Eb_reg[12]/P0001 , \core_c_psq_Taddr_Eb_reg[13]/P0001 , \core_c_psq_Taddr_Eb_reg[1]/P0001 , \core_c_psq_Taddr_Eb_reg[2]/P0001 , \core_c_psq_Taddr_Eb_reg[3]/P0001 , \core_c_psq_Taddr_Eb_reg[4]/P0001 , \core_c_psq_Taddr_Eb_reg[5]/P0001 , \core_c_psq_Taddr_Eb_reg[6]/P0001 , \core_c_psq_Taddr_Eb_reg[7]/P0001 , \core_c_psq_Taddr_Eb_reg[8]/P0001 , \core_c_psq_Taddr_Eb_reg[9]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001 , \core_c_psq_cntstk_ptr_reg[0]/NET0131 , \core_c_psq_cntstk_ptr_reg[1]/NET0131 , \core_c_psq_cntstk_ptr_reg[2]/NET0131 , \core_c_psq_irq0_de_IN_syn_reg/P0001 , \core_c_psq_irq0_de_OUT_reg/P0001 , \core_c_psq_irq1_de_IN_syn_reg/P0001 , \core_c_psq_irq1_de_OUT_reg/P0001 , \core_c_psq_irq2_de_IN_syn_reg/P0001 , \core_c_psq_irq2_de_OUT_reg/P0001 , \core_c_psq_irql0_de_IN_syn_reg/P0001 , \core_c_psq_irql0_de_OUT_reg/P0001 , \core_c_psq_irql1_de_IN_syn_reg/P0001 , \core_c_psq_irql1_de_OUT_reg/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001 , \core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001 , \core_c_psq_lpstk_ptr_reg[0]/NET0131 , \core_c_psq_lpstk_ptr_reg[1]/NET0131 , \core_c_psq_lpstk_ptr_reg[2]/NET0131 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001 , \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001 , \core_c_psq_pcstk_ptr_reg[0]/NET0131 , \core_c_psq_pcstk_ptr_reg[1]/NET0131 , \core_c_psq_pcstk_ptr_reg[2]/NET0131 , \core_c_psq_pcstk_ptr_reg[3]/NET0131 , \core_c_psq_pcstk_ptr_reg[4]/NET0131 , \core_c_psq_ststk_ptr_reg[0]/NET0131 , \core_c_psq_ststk_ptr_reg[1]/NET0131 , \core_c_psq_ststk_ptr_reg[2]/NET0131 , \core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001 , \core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001 , \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 , \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_I_reg[0]/NET0131 , \core_dag_ilm1reg_I_reg[10]/NET0131 , \core_dag_ilm1reg_I_reg[11]/NET0131 , \core_dag_ilm1reg_I_reg[12]/NET0131 , \core_dag_ilm1reg_I_reg[13]/NET0131 , \core_dag_ilm1reg_I_reg[1]/NET0131 , \core_dag_ilm1reg_I_reg[2]/NET0131 , \core_dag_ilm1reg_I_reg[3]/NET0131 , \core_dag_ilm1reg_I_reg[4]/NET0131 , \core_dag_ilm1reg_I_reg[5]/NET0131 , \core_dag_ilm1reg_I_reg[6]/NET0131 , \core_dag_ilm1reg_I_reg[7]/NET0131 , \core_dag_ilm1reg_I_reg[8]/NET0131 , \core_dag_ilm1reg_I_reg[9]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_L_reg[0]/NET0131 , \core_dag_ilm1reg_L_reg[10]/NET0131 , \core_dag_ilm1reg_L_reg[11]/NET0131 , \core_dag_ilm1reg_L_reg[12]/NET0131 , \core_dag_ilm1reg_L_reg[13]/NET0131 , \core_dag_ilm1reg_L_reg[1]/NET0131 , \core_dag_ilm1reg_L_reg[2]/NET0131 , \core_dag_ilm1reg_L_reg[3]/NET0131 , \core_dag_ilm1reg_L_reg[4]/NET0131 , \core_dag_ilm1reg_L_reg[5]/NET0131 , \core_dag_ilm1reg_L_reg[6]/NET0131 , \core_dag_ilm1reg_L_reg[7]/NET0131 , \core_dag_ilm1reg_L_reg[8]/NET0131 , \core_dag_ilm1reg_L_reg[9]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131 , \core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131 , \core_dag_ilm1reg_M_reg[0]/NET0131 , \core_dag_ilm1reg_M_reg[10]/NET0131 , \core_dag_ilm1reg_M_reg[11]/NET0131 , \core_dag_ilm1reg_M_reg[12]/NET0131 , \core_dag_ilm1reg_M_reg[13]/NET0131 , \core_dag_ilm1reg_M_reg[1]/NET0131 , \core_dag_ilm1reg_M_reg[2]/NET0131 , \core_dag_ilm1reg_M_reg[3]/NET0131 , \core_dag_ilm1reg_M_reg[4]/NET0131 , \core_dag_ilm1reg_M_reg[5]/NET0131 , \core_dag_ilm1reg_M_reg[6]/NET0131 , \core_dag_ilm1reg_M_reg[7]/NET0131 , \core_dag_ilm1reg_M_reg[8]/NET0131 , \core_dag_ilm1reg_M_reg[9]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131 , \core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131 , \core_dag_ilm1reg_STEALI_E_reg[0]/P0001 , \core_dag_ilm1reg_STEALI_E_reg[1]/P0001 , \core_dag_ilm1reg_STEALI_E_reg[2]/P0001 , \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_IL_E_reg[0]/P0001 , \core_dag_ilm2reg_IL_E_reg[1]/P0001 , \core_dag_ilm2reg_I_reg[0]/NET0131 , \core_dag_ilm2reg_I_reg[10]/NET0131 , \core_dag_ilm2reg_I_reg[11]/NET0131 , \core_dag_ilm2reg_I_reg[12]/NET0131 , \core_dag_ilm2reg_I_reg[13]/NET0131 , \core_dag_ilm2reg_I_reg[1]/NET0131 , \core_dag_ilm2reg_I_reg[2]/NET0131 , \core_dag_ilm2reg_I_reg[3]/NET0131 , \core_dag_ilm2reg_I_reg[4]/NET0131 , \core_dag_ilm2reg_I_reg[5]/NET0131 , \core_dag_ilm2reg_I_reg[6]/NET0131 , \core_dag_ilm2reg_I_reg[7]/NET0131 , \core_dag_ilm2reg_I_reg[8]/NET0131 , \core_dag_ilm2reg_I_reg[9]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_L_reg[0]/NET0131 , \core_dag_ilm2reg_L_reg[10]/NET0131 , \core_dag_ilm2reg_L_reg[11]/NET0131 , \core_dag_ilm2reg_L_reg[12]/NET0131 , \core_dag_ilm2reg_L_reg[13]/NET0131 , \core_dag_ilm2reg_L_reg[1]/NET0131 , \core_dag_ilm2reg_L_reg[2]/NET0131 , \core_dag_ilm2reg_L_reg[3]/NET0131 , \core_dag_ilm2reg_L_reg[4]/NET0131 , \core_dag_ilm2reg_L_reg[5]/NET0131 , \core_dag_ilm2reg_L_reg[6]/NET0131 , \core_dag_ilm2reg_L_reg[7]/NET0131 , \core_dag_ilm2reg_L_reg[8]/NET0131 , \core_dag_ilm2reg_L_reg[9]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131 , \core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131 , \core_dag_ilm2reg_M_E_reg[0]/NET0131 , \core_dag_ilm2reg_M_E_reg[1]/NET0131 , \core_dag_ilm2reg_M_reg[0]/NET0131 , \core_dag_ilm2reg_M_reg[10]/NET0131 , \core_dag_ilm2reg_M_reg[11]/NET0131 , \core_dag_ilm2reg_M_reg[12]/NET0131 , \core_dag_ilm2reg_M_reg[13]/NET0131 , \core_dag_ilm2reg_M_reg[1]/NET0131 , \core_dag_ilm2reg_M_reg[2]/NET0131 , \core_dag_ilm2reg_M_reg[3]/NET0131 , \core_dag_ilm2reg_M_reg[4]/NET0131 , \core_dag_ilm2reg_M_reg[5]/NET0131 , \core_dag_ilm2reg_M_reg[6]/NET0131 , \core_dag_ilm2reg_M_reg[7]/NET0131 , \core_dag_ilm2reg_M_reg[8]/NET0131 , \core_dag_ilm2reg_M_reg[9]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 , \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 , \core_dag_modulo1_R0wrap_reg/P0001 , \core_dag_modulo1_R1wrap_reg/P0001 , \core_dag_modulo1_T0wrap_reg/P0001 , \core_dag_modulo1_T1wrap_reg/P0001 , \core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 , \core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 , \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 , \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 , \core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001 , \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001 , \core_eu_ec_cun_AC_reg/P0001 , \core_eu_ec_cun_AN_reg/P0001 , \core_eu_ec_cun_AQ_reg/P0001 , \core_eu_ec_cun_AS_reg/P0001 , \core_eu_ec_cun_AV_reg/P0001 , \core_eu_ec_cun_AZ_reg/P0001 , \core_eu_ec_cun_COND_E_reg[0]/P0001 , \core_eu_ec_cun_COND_E_reg[1]/P0001 , \core_eu_ec_cun_COND_E_reg[2]/P0001 , \core_eu_ec_cun_COND_E_reg[3]/P0001 , \core_eu_ec_cun_MV_reg/P0000_reg_syn_2 , \core_eu_ec_cun_MVi_pre_C_reg/P0001 , \core_eu_ec_cun_SS_reg/P0001 , \core_eu_ec_cun_TERM_E_reg[0]/P0001 , \core_eu_ec_cun_TERM_E_reg[1]/P0001 , \core_eu_ec_cun_TERM_E_reg[2]/P0001 , \core_eu_ec_cun_TERM_E_reg[3]/P0001 , \core_eu_ec_cun_condOK_CE_reg/P0001 , \core_eu_ec_cun_mven_FFout_reg/NET0131 , \core_eu_ec_cun_termOK_CE_reg/P0001 , \core_eu_ec_cun_updateMV_C_reg/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 , \core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_Sq_E_reg/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 , \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 , \core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 , \core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2 , \core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2 , \core_eu_es_sht_es_reg_SBr_reg[0]/P0001 , \core_eu_es_sht_es_reg_SBr_reg[1]/P0001 , \core_eu_es_sht_es_reg_SBr_reg[2]/P0001 , \core_eu_es_sht_es_reg_SBr_reg[3]/P0001 , \core_eu_es_sht_es_reg_SBr_reg[4]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[0]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[1]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[2]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[3]/P0001 , \core_eu_es_sht_es_reg_SBs_reg[4]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 , \core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 , \emc_DMDoe_reg/NET0131 , \emc_DMDreg_reg[0]/P0001 , \emc_DMDreg_reg[10]/P0001 , \emc_DMDreg_reg[11]/P0001 , \emc_DMDreg_reg[12]/P0001 , \emc_DMDreg_reg[13]/P0001 , \emc_DMDreg_reg[14]/P0001 , \emc_DMDreg_reg[15]/P0001 , \emc_DMDreg_reg[1]/P0001 , \emc_DMDreg_reg[2]/P0001 , \emc_DMDreg_reg[3]/P0001 , \emc_DMDreg_reg[4]/P0001 , \emc_DMDreg_reg[5]/P0001 , \emc_DMDreg_reg[6]/P0001 , \emc_DMDreg_reg[7]/P0001 , \emc_DMDreg_reg[8]/P0001 , \emc_DMDreg_reg[9]/P0001 , \emc_DMcst_reg/NET0131 , \emc_ECMA_reg[0]/P0001 , \emc_ECMA_reg[10]/P0001 , \emc_ECMA_reg[11]/P0001 , \emc_ECMA_reg[12]/P0001 , \emc_ECMA_reg[1]/P0001 , \emc_ECMA_reg[2]/P0001 , \emc_ECMA_reg[3]/P0001 , \emc_ECMA_reg[4]/P0001 , \emc_ECMA_reg[5]/P0001 , \emc_ECMA_reg[6]/P0001 , \emc_ECMA_reg[7]/P0001 , \emc_ECMA_reg[8]/P0001 , \emc_ECMA_reg[9]/P0001 , \emc_ECMDreg_reg[0]/P0001 , \emc_ECMDreg_reg[10]/P0001 , \emc_ECMDreg_reg[11]/P0001 , \emc_ECMDreg_reg[12]/P0001 , \emc_ECMDreg_reg[13]/P0001 , \emc_ECMDreg_reg[14]/P0001 , \emc_ECMDreg_reg[15]/P0001 , \emc_ECMDreg_reg[16]/P0001 , \emc_ECMDreg_reg[17]/P0001 , \emc_ECMDreg_reg[18]/P0001 , \emc_ECMDreg_reg[19]/P0001 , \emc_ECMDreg_reg[1]/P0001 , \emc_ECMDreg_reg[20]/P0001 , \emc_ECMDreg_reg[21]/P0001 , \emc_ECMDreg_reg[22]/P0001 , \emc_ECMDreg_reg[23]/P0001 , \emc_ECMDreg_reg[2]/P0001 , \emc_ECMDreg_reg[3]/P0001 , \emc_ECMDreg_reg[4]/P0001 , \emc_ECMDreg_reg[5]/P0001 , \emc_ECMDreg_reg[6]/P0001 , \emc_ECMDreg_reg[7]/P0001 , \emc_ECMDreg_reg[8]/P0001 , \emc_ECMDreg_reg[9]/P0001 , \emc_ECMcs_reg/NET0131 , \emc_ECS_reg[0]/NET0131 , \emc_ECS_reg[1]/NET0131 , \emc_ECS_reg[2]/NET0131 , \emc_ECS_reg[3]/NET0131 , \emc_ED_oei_reg/P0001 , \emc_EXTC_Eg_syn_reg/P0001 , \emc_IOcst_reg/NET0131 , \emc_PMDoe_reg/NET0131 , \emc_PMDreg_reg[0]/P0001 , \emc_PMDreg_reg[10]/P0001 , \emc_PMDreg_reg[11]/P0001 , \emc_PMDreg_reg[12]/P0001 , \emc_PMDreg_reg[13]/P0001 , \emc_PMDreg_reg[14]/P0001 , \emc_PMDreg_reg[15]/P0001 , \emc_PMDreg_reg[1]/P0001 , \emc_PMDreg_reg[2]/P0001 , \emc_PMDreg_reg[3]/P0001 , \emc_PMDreg_reg[4]/P0001 , \emc_PMDreg_reg[5]/P0001 , \emc_PMDreg_reg[6]/P0001 , \emc_PMDreg_reg[7]/P0001 , \emc_PMDreg_reg[8]/P0001 , \emc_PMDreg_reg[9]/P0001 , \emc_PMcst_reg/NET0131 , \emc_RWcnt_reg[0]/P0001 , \emc_RWcnt_reg[1]/P0001 , \emc_RWcnt_reg[2]/P0001 , \emc_RWcnt_reg[3]/P0001 , \emc_RWcnt_reg[4]/P0001 , \emc_RWcnt_reg[5]/P0001 , \emc_WRn_h_reg/P0001 , \emc_WSCRext_reg_DO_reg[0]/NET0131 , \emc_WSCRext_reg_DO_reg[1]/NET0131 , \emc_WSCRext_reg_DO_reg[2]/NET0131 , \emc_WSCRext_reg_DO_reg[3]/NET0131 , \emc_WSCRext_reg_DO_reg[4]/NET0131 , \emc_WSCRext_reg_DO_reg[5]/NET0131 , \emc_WSCRext_reg_DO_reg[6]/NET0131 , \emc_WSCRext_reg_DO_reg[7]/NET0131 , \emc_WSCRreg_DO_reg[0]/NET0131 , \emc_WSCRreg_DO_reg[10]/NET0131 , \emc_WSCRreg_DO_reg[11]/NET0131 , \emc_WSCRreg_DO_reg[12]/NET0131 , \emc_WSCRreg_DO_reg[13]/NET0131 , \emc_WSCRreg_DO_reg[14]/NET0131 , \emc_WSCRreg_DO_reg[1]/NET0131 , \emc_WSCRreg_DO_reg[2]/NET0131 , \emc_WSCRreg_DO_reg[3]/NET0131 , \emc_WSCRreg_DO_reg[4]/NET0131 , \emc_WSCRreg_DO_reg[5]/NET0131 , \emc_WSCRreg_DO_reg[6]/NET0131 , \emc_WSCRreg_DO_reg[7]/NET0131 , \emc_WSCRreg_DO_reg[8]/NET0131 , \emc_WSCRreg_DO_reg[9]/NET0131 , \emc_eRDY_reg/NET0131 , \emc_selDMDi_reg/P0001 , \emc_selPMDi_reg/P0001 , \idma_CM_oe_reg/P0001 , \idma_CMo_oe0_reg/P0001 , \idma_CMo_oe1_reg/P0001 , \idma_CMo_oe2_reg/P0001 , \idma_CMo_oe3_reg/P0001 , \idma_CMo_oe4_reg/P0001 , \idma_CMo_oe5_reg/P0001 , \idma_CMo_oe6_reg/P0001 , \idma_CMo_oe7_reg/P0001 , \idma_DCTL_reg[0]/NET0131 , \idma_DCTL_reg[10]/NET0131 , \idma_DCTL_reg[11]/NET0131 , \idma_DCTL_reg[12]/NET0131 , \idma_DCTL_reg[13]/NET0131 , \idma_DCTL_reg[14]/NET0131 , \idma_DCTL_reg[1]/NET0131 , \idma_DCTL_reg[2]/NET0131 , \idma_DCTL_reg[3]/NET0131 , \idma_DCTL_reg[4]/NET0131 , \idma_DCTL_reg[5]/NET0131 , \idma_DCTL_reg[6]/NET0131 , \idma_DCTL_reg[7]/NET0131 , \idma_DCTL_reg[8]/NET0131 , \idma_DCTL_reg[9]/NET0131 , \idma_DOVL_reg[0]/NET0131 , \idma_DOVL_reg[10]/NET0131 , \idma_DOVL_reg[11]/NET0131 , \idma_DOVL_reg[1]/NET0131 , \idma_DOVL_reg[2]/NET0131 , \idma_DOVL_reg[3]/NET0131 , \idma_DOVL_reg[4]/NET0131 , \idma_DOVL_reg[5]/NET0131 , \idma_DOVL_reg[6]/NET0131 , \idma_DOVL_reg[7]/NET0131 , \idma_DOVL_reg[8]/NET0131 , \idma_DOVL_reg[9]/NET0131 , \idma_DSreq_reg/NET0131 , \idma_DTMP_H_reg[0]/P0001 , \idma_DTMP_H_reg[10]/P0001 , \idma_DTMP_H_reg[11]/P0001 , \idma_DTMP_H_reg[12]/P0001 , \idma_DTMP_H_reg[13]/P0001 , \idma_DTMP_H_reg[14]/P0001 , \idma_DTMP_H_reg[15]/P0001 , \idma_DTMP_H_reg[1]/P0001 , \idma_DTMP_H_reg[2]/P0001 , \idma_DTMP_H_reg[3]/P0001 , \idma_DTMP_H_reg[4]/P0001 , \idma_DTMP_H_reg[5]/P0001 , \idma_DTMP_H_reg[6]/P0001 , \idma_DTMP_H_reg[7]/P0001 , \idma_DTMP_H_reg[8]/P0001 , \idma_DTMP_H_reg[9]/P0001 , \idma_DTMP_L_reg[0]/P0001 , \idma_DTMP_L_reg[1]/P0001 , \idma_DTMP_L_reg[2]/P0001 , \idma_DTMP_L_reg[3]/P0001 , \idma_DTMP_L_reg[4]/P0001 , \idma_DTMP_L_reg[5]/P0001 , \idma_DTMP_L_reg[6]/P0001 , \idma_DTMP_L_reg[7]/P0001 , \idma_IADi_reg[0]/P0001 , \idma_IADi_reg[10]/P0001 , \idma_IADi_reg[11]/P0001 , \idma_IADi_reg[12]/P0001 , \idma_IADi_reg[13]/P0001 , \idma_IADi_reg[14]/P0001 , \idma_IADi_reg[15]/P0001 , \idma_IADi_reg[1]/P0001 , \idma_IADi_reg[2]/P0001 , \idma_IADi_reg[3]/P0001 , \idma_IADi_reg[4]/P0001 , \idma_IADi_reg[5]/P0001 , \idma_IADi_reg[6]/P0001 , \idma_IADi_reg[7]/P0001 , \idma_IADi_reg[8]/P0001 , \idma_IADi_reg[9]/P0001 , \idma_IAL_reg/P0001 , \idma_IDMA_boot_reg/NET0131_reg_syn_10 , \idma_IDMA_boot_reg/NET0131_reg_syn_2 , \idma_IDMA_boot_reg/NET0131_reg_syn_8 , \idma_IRDn_reg/P0001 , \idma_ISn_reg/P0001 , \idma_IWRn_reg/P0001 , \idma_PCrd_1st_reg/NET0131 , \idma_PM_1st_reg/NET0131 , \idma_RDCMD_d1_reg/P0001 , \idma_RDCMD_reg/P0001 , \idma_RDcnt_reg[0]/NET0131 , \idma_RDcnt_reg[1]/NET0131 , \idma_RDcnt_reg[2]/NET0131 , \idma_RDcyc_reg/NET0131 , \idma_WRCMD_d1_reg/P0001 , \idma_WRCMD_reg/P0001 , \idma_WRcnt_reg[0]/NET0131 , \idma_WRcnt_reg[1]/NET0131 , \idma_WRcnt_reg[2]/NET0131 , \idma_WRcyc_reg/NET0131 , \idma_WRtrue_reg/NET0131 , \memc_DM_oe_reg/P0001 , \memc_DMo_oe0_reg/P0001 , \memc_DMo_oe1_reg/P0001 , \memc_DMo_oe2_reg/P0001 , \memc_DMo_oe3_reg/P0001 , \memc_DMo_oe4_reg/P0001 , \memc_DMo_oe5_reg/P0001 , \memc_DMo_oe6_reg/P0001 , \memc_DMo_oe7_reg/P0001 , \memc_Dread_E_reg/NET0131 , \memc_Dwrite_C_reg/NET0131 , \memc_Dwrite_E_reg/NET0131 , \memc_EXTC_E_reg/NET0131 , \memc_EXTC_Eg_reg/NET0131_reg_syn_10 , \memc_EXTC_Eg_reg/NET0131_reg_syn_2 , \memc_EXTC_Eg_reg/NET0131_reg_syn_8 , \memc_IOcmd_E_reg/NET0131 , \memc_LDaST_Eg_reg/NET0131 , \memc_MMR_web_reg/NET0131 , \memc_PMo_oe0_reg/P0001 , \memc_PMo_oe1_reg/P0001 , \memc_PMo_oe2_reg/P0001 , \memc_PMo_oe3_reg/P0001 , \memc_PMo_oe4_reg/P0001 , \memc_PMo_oe5_reg/P0001 , \memc_PMo_oe6_reg/P0001 , \memc_PMo_oe7_reg/P0001 , \memc_Pread_E_reg/NET0131 , \memc_Pwrite_C_reg/NET0131 , \memc_Pwrite_E_reg/NET0131 , \memc_STI_Cg_reg/NET0131 , \memc_accDM_E_reg/NET0131 , \memc_accPM_E_reg/NET0131 , \memc_ldSREG_E_reg/NET0131 , \memc_selMIO_E_reg/P0001 , \memc_usysr_DO_reg[0]/NET0131 , \memc_usysr_DO_reg[10]/NET0131 , \memc_usysr_DO_reg[11]/NET0131 , \memc_usysr_DO_reg[12]/NET0131 , \memc_usysr_DO_reg[13]/NET0131 , \memc_usysr_DO_reg[14]/NET0131 , \memc_usysr_DO_reg[15]/NET0131 , \memc_usysr_DO_reg[1]/NET0131 , \memc_usysr_DO_reg[2]/NET0131 , \memc_usysr_DO_reg[3]/NET0131 , \memc_usysr_DO_reg[4]/NET0131 , \memc_usysr_DO_reg[5]/NET0131 , \memc_usysr_DO_reg[6]/NET0131 , \memc_usysr_DO_reg[7]/NET0131 , \memc_usysr_DO_reg[8]/NET0131 , \memc_usysr_DO_reg[9]/NET0131 , \pio_PINT_reg[0]/NET0131 , \pio_PINT_reg[10]/NET0131 , \pio_PINT_reg[11]/NET0131 , \pio_PINT_reg[1]/NET0131 , \pio_PINT_reg[2]/NET0131 , \pio_PINT_reg[3]/NET0131 , \pio_PINT_reg[4]/NET0131 , \pio_PINT_reg[5]/NET0131 , \pio_PINT_reg[6]/NET0131 , \pio_PINT_reg[7]/NET0131 , \pio_PINT_reg[8]/NET0131 , \pio_PINT_reg[9]/NET0131 , \pio_PIO_IN_P_reg[0]/P0001 , \pio_PIO_IN_P_reg[10]/P0001 , \pio_PIO_IN_P_reg[11]/P0001 , \pio_PIO_IN_P_reg[1]/P0001 , \pio_PIO_IN_P_reg[2]/P0001 , \pio_PIO_IN_P_reg[3]/P0001 , \pio_PIO_IN_P_reg[4]/P0001 , \pio_PIO_IN_P_reg[5]/P0001 , \pio_PIO_IN_P_reg[6]/P0001 , \pio_PIO_IN_P_reg[7]/P0001 , \pio_PIO_IN_P_reg[8]/P0001 , \pio_PIO_IN_P_reg[9]/P0001 , \pio_PIO_RES_OUT_reg[0]/P0001 , \pio_PIO_RES_OUT_reg[10]/P0001 , \pio_PIO_RES_OUT_reg[11]/P0001 , \pio_PIO_RES_OUT_reg[1]/P0001 , \pio_PIO_RES_OUT_reg[2]/P0001 , \pio_PIO_RES_OUT_reg[3]/P0001 , \pio_PIO_RES_OUT_reg[4]/P0001 , \pio_PIO_RES_OUT_reg[5]/P0001 , \pio_PIO_RES_OUT_reg[6]/P0001 , \pio_PIO_RES_OUT_reg[7]/P0001 , \pio_PIO_RES_OUT_reg[8]/P0001 , \pio_PIO_RES_OUT_reg[9]/P0001 , \pio_PIO_RES_reg[0]/NET0131 , \pio_PIO_RES_reg[10]/NET0131 , \pio_PIO_RES_reg[11]/NET0131 , \pio_PIO_RES_reg[1]/NET0131 , \pio_PIO_RES_reg[2]/NET0131 , \pio_PIO_RES_reg[3]/NET0131 , \pio_PIO_RES_reg[4]/NET0131 , \pio_PIO_RES_reg[5]/NET0131 , \pio_PIO_RES_reg[6]/NET0131 , \pio_PIO_RES_reg[7]/NET0131 , \pio_PIO_RES_reg[8]/NET0131 , \pio_PIO_RES_reg[9]/NET0131 , \pio_pmask_reg_DO_reg[0]/NET0131 , \pio_pmask_reg_DO_reg[10]/NET0131 , \pio_pmask_reg_DO_reg[11]/NET0131 , \pio_pmask_reg_DO_reg[1]/NET0131 , \pio_pmask_reg_DO_reg[2]/NET0131 , \pio_pmask_reg_DO_reg[3]/NET0131 , \pio_pmask_reg_DO_reg[4]/NET0131 , \pio_pmask_reg_DO_reg[5]/NET0131 , \pio_pmask_reg_DO_reg[6]/NET0131 , \pio_pmask_reg_DO_reg[7]/NET0131 , \pio_pmask_reg_DO_reg[8]/NET0131 , \pio_pmask_reg_DO_reg[9]/NET0131 , \regout_STD_C_reg[0]/P0001 , \regout_STD_C_reg[10]/P0001 , \regout_STD_C_reg[11]/P0001 , \regout_STD_C_reg[12]/P0001 , \regout_STD_C_reg[13]/P0001 , \regout_STD_C_reg[14]/P0001 , \regout_STD_C_reg[15]/P0001 , \regout_STD_C_reg[1]/P0001 , \regout_STD_C_reg[2]/P0001 , \regout_STD_C_reg[3]/P0001 , \regout_STD_C_reg[4]/P0001 , \regout_STD_C_reg[5]/P0001 , \regout_STD_C_reg[6]/P0001 , \regout_STD_C_reg[7]/P0001 , \regout_STD_C_reg[8]/P0001 , \regout_STD_C_reg[9]/P0001 , \sice_CLR_I_reg/NET0131 , \sice_CLR_M_reg/NET0131 , \sice_CMRW_reg/NET0131 , \sice_DBR1_reg[0]/P0001 , \sice_DBR1_reg[10]/P0001 , \sice_DBR1_reg[11]/P0001 , \sice_DBR1_reg[12]/P0001 , \sice_DBR1_reg[13]/P0001 , \sice_DBR1_reg[14]/P0001 , \sice_DBR1_reg[15]/P0001 , \sice_DBR1_reg[16]/P0001 , \sice_DBR1_reg[17]/P0001 , \sice_DBR1_reg[18]/P0001 , \sice_DBR1_reg[1]/P0001 , \sice_DBR1_reg[2]/P0001 , \sice_DBR1_reg[3]/P0001 , \sice_DBR1_reg[4]/P0001 , \sice_DBR1_reg[5]/P0001 , \sice_DBR1_reg[6]/P0001 , \sice_DBR1_reg[7]/P0001 , \sice_DBR1_reg[8]/P0001 , \sice_DBR1_reg[9]/P0001 , \sice_DBR2_reg[0]/P0001 , \sice_DBR2_reg[10]/P0001 , \sice_DBR2_reg[11]/P0001 , \sice_DBR2_reg[12]/P0001 , \sice_DBR2_reg[13]/P0001 , \sice_DBR2_reg[14]/P0001 , \sice_DBR2_reg[15]/P0001 , \sice_DBR2_reg[16]/P0001 , \sice_DBR2_reg[17]/P0001 , \sice_DBR2_reg[18]/P0001 , \sice_DBR2_reg[1]/P0001 , \sice_DBR2_reg[2]/P0001 , \sice_DBR2_reg[3]/P0001 , \sice_DBR2_reg[4]/P0001 , \sice_DBR2_reg[5]/P0001 , \sice_DBR2_reg[6]/P0001 , \sice_DBR2_reg[7]/P0001 , \sice_DBR2_reg[8]/P0001 , \sice_DBR2_reg[9]/P0001 , \sice_DMR1_reg[0]/NET0131 , \sice_DMR1_reg[10]/NET0131 , \sice_DMR1_reg[11]/NET0131 , \sice_DMR1_reg[12]/NET0131 , \sice_DMR1_reg[13]/NET0131 , \sice_DMR1_reg[14]/NET0131 , \sice_DMR1_reg[15]/NET0131 , \sice_DMR1_reg[16]/NET0131 , \sice_DMR1_reg[17]/NET0131 , \sice_DMR1_reg[1]/NET0131 , \sice_DMR1_reg[2]/NET0131 , \sice_DMR1_reg[3]/NET0131 , \sice_DMR1_reg[4]/NET0131 , \sice_DMR1_reg[5]/NET0131 , \sice_DMR1_reg[6]/NET0131 , \sice_DMR1_reg[7]/NET0131 , \sice_DMR1_reg[8]/NET0131 , \sice_DMR1_reg[9]/NET0131 , \sice_DMR2_reg[0]/NET0131 , \sice_DMR2_reg[10]/NET0131 , \sice_DMR2_reg[11]/NET0131 , \sice_DMR2_reg[12]/NET0131 , \sice_DMR2_reg[13]/NET0131 , \sice_DMR2_reg[14]/NET0131 , \sice_DMR2_reg[15]/NET0131 , \sice_DMR2_reg[16]/NET0131 , \sice_DMR2_reg[17]/NET0131 , \sice_DMR2_reg[1]/NET0131 , \sice_DMR2_reg[2]/NET0131 , \sice_DMR2_reg[3]/NET0131 , \sice_DMR2_reg[4]/NET0131 , \sice_DMR2_reg[5]/NET0131 , \sice_DMR2_reg[6]/NET0131 , \sice_DMR2_reg[7]/NET0131 , \sice_DMR2_reg[8]/NET0131 , \sice_DMR2_reg[9]/NET0131 , \sice_GOICE_1_reg/NET0131 , \sice_GOICE_2_reg/NET0131 , \sice_GOICE_s1_reg/NET0131 , \sice_GOICE_syn_reg/P0001 , \sice_GO_NX_reg/NET0131 , \sice_GO_NXi_reg/NET0131 , \sice_HALT_E_reg/P0001 , \sice_IAR_reg[0]/NET0131 , \sice_IAR_reg[1]/NET0131 , \sice_IAR_reg[2]/NET0131 , \sice_IAR_reg[3]/NET0131 , \sice_IBR1_reg[0]/P0001 , \sice_IBR1_reg[10]/P0001 , \sice_IBR1_reg[11]/P0001 , \sice_IBR1_reg[12]/P0001 , \sice_IBR1_reg[13]/P0001 , \sice_IBR1_reg[14]/P0001 , \sice_IBR1_reg[15]/P0001 , \sice_IBR1_reg[16]/P0001 , \sice_IBR1_reg[17]/P0001 , \sice_IBR1_reg[1]/P0001 , \sice_IBR1_reg[2]/P0001 , \sice_IBR1_reg[3]/P0001 , \sice_IBR1_reg[4]/P0001 , \sice_IBR1_reg[5]/P0001 , \sice_IBR1_reg[6]/P0001 , \sice_IBR1_reg[7]/P0001 , \sice_IBR1_reg[8]/P0001 , \sice_IBR1_reg[9]/P0001 , \sice_IBR2_reg[0]/P0001 , \sice_IBR2_reg[10]/P0001 , \sice_IBR2_reg[11]/P0001 , \sice_IBR2_reg[12]/P0001 , \sice_IBR2_reg[13]/P0001 , \sice_IBR2_reg[14]/P0001 , \sice_IBR2_reg[15]/P0001 , \sice_IBR2_reg[16]/P0001 , \sice_IBR2_reg[17]/P0001 , \sice_IBR2_reg[1]/P0001 , \sice_IBR2_reg[2]/P0001 , \sice_IBR2_reg[3]/P0001 , \sice_IBR2_reg[4]/P0001 , \sice_IBR2_reg[5]/P0001 , \sice_IBR2_reg[6]/P0001 , \sice_IBR2_reg[7]/P0001 , \sice_IBR2_reg[8]/P0001 , \sice_IBR2_reg[9]/P0001 , \sice_ICS_reg[0]/NET0131 , \sice_ICS_reg[1]/NET0131 , \sice_ICS_reg[2]/NET0131 , \sice_ICYC_clr_reg/NET0131 , \sice_ICYC_en_reg/NET0131 , \sice_ICYC_en_syn_reg/P0001 , \sice_ICYC_reg[0]/NET0131 , \sice_ICYC_reg[10]/NET0131 , \sice_ICYC_reg[11]/NET0131 , \sice_ICYC_reg[12]/NET0131 , \sice_ICYC_reg[13]/NET0131 , \sice_ICYC_reg[14]/NET0131 , \sice_ICYC_reg[15]/NET0131 , \sice_ICYC_reg[16]/NET0131 , \sice_ICYC_reg[17]/NET0131 , \sice_ICYC_reg[18]/NET0131 , \sice_ICYC_reg[19]/NET0131 , \sice_ICYC_reg[1]/NET0131 , \sice_ICYC_reg[20]/NET0131 , \sice_ICYC_reg[21]/NET0131 , \sice_ICYC_reg[22]/NET0131 , \sice_ICYC_reg[23]/NET0131 , \sice_ICYC_reg[2]/NET0131 , \sice_ICYC_reg[3]/NET0131 , \sice_ICYC_reg[4]/NET0131 , \sice_ICYC_reg[5]/NET0131 , \sice_ICYC_reg[6]/NET0131 , \sice_ICYC_reg[7]/NET0131 , \sice_ICYC_reg[8]/NET0131 , \sice_ICYC_reg[9]/NET0131 , \sice_IDONE_reg/NET0131 , \sice_IIRC_reg[0]/NET0131 , \sice_IIRC_reg[10]/NET0131 , \sice_IIRC_reg[11]/NET0131 , \sice_IIRC_reg[12]/NET0131 , \sice_IIRC_reg[13]/NET0131 , \sice_IIRC_reg[14]/NET0131 , \sice_IIRC_reg[15]/NET0131 , \sice_IIRC_reg[16]/NET0131 , \sice_IIRC_reg[17]/NET0131 , \sice_IIRC_reg[18]/NET0131 , \sice_IIRC_reg[19]/NET0131 , \sice_IIRC_reg[1]/NET0131 , \sice_IIRC_reg[20]/NET0131 , \sice_IIRC_reg[21]/NET0131 , \sice_IIRC_reg[22]/NET0131 , \sice_IIRC_reg[23]/NET0131 , \sice_IIRC_reg[2]/NET0131 , \sice_IIRC_reg[3]/NET0131 , \sice_IIRC_reg[4]/NET0131 , \sice_IIRC_reg[5]/NET0131 , \sice_IIRC_reg[6]/NET0131 , \sice_IIRC_reg[7]/NET0131 , \sice_IIRC_reg[8]/NET0131 , \sice_IIRC_reg[9]/NET0131 , \sice_IMR1_reg[0]/NET0131 , \sice_IMR1_reg[10]/NET0131 , \sice_IMR1_reg[11]/NET0131 , \sice_IMR1_reg[12]/NET0131 , \sice_IMR1_reg[13]/NET0131 , \sice_IMR1_reg[14]/NET0131 , \sice_IMR1_reg[15]/NET0131 , \sice_IMR1_reg[16]/NET0131 , \sice_IMR1_reg[17]/NET0131 , \sice_IMR1_reg[1]/NET0131 , \sice_IMR1_reg[2]/NET0131 , \sice_IMR1_reg[3]/NET0131 , \sice_IMR1_reg[4]/NET0131 , \sice_IMR1_reg[5]/NET0131 , \sice_IMR1_reg[6]/NET0131 , \sice_IMR1_reg[7]/NET0131 , \sice_IMR1_reg[8]/NET0131 , \sice_IMR1_reg[9]/NET0131 , \sice_IMR2_reg[0]/NET0131 , \sice_IMR2_reg[10]/NET0131 , \sice_IMR2_reg[11]/NET0131 , \sice_IMR2_reg[12]/NET0131 , \sice_IMR2_reg[13]/NET0131 , \sice_IMR2_reg[14]/NET0131 , \sice_IMR2_reg[15]/NET0131 , \sice_IMR2_reg[16]/NET0131 , \sice_IMR2_reg[17]/NET0131 , \sice_IMR2_reg[1]/NET0131 , \sice_IMR2_reg[2]/NET0131 , \sice_IMR2_reg[3]/NET0131 , \sice_IMR2_reg[4]/NET0131 , \sice_IMR2_reg[5]/NET0131 , \sice_IMR2_reg[6]/NET0131 , \sice_IMR2_reg[7]/NET0131 , \sice_IMR2_reg[8]/NET0131 , \sice_IMR2_reg[9]/NET0131 , \sice_IRR_reg[0]/P0001 , \sice_IRR_reg[10]/P0001 , \sice_IRR_reg[11]/P0001 , \sice_IRR_reg[12]/P0001 , \sice_IRR_reg[13]/P0001 , \sice_IRR_reg[1]/P0001 , \sice_IRR_reg[2]/P0001 , \sice_IRR_reg[3]/P0001 , \sice_IRR_reg[4]/P0001 , \sice_IRR_reg[5]/P0001 , \sice_IRR_reg[6]/P0001 , \sice_IRR_reg[7]/P0001 , \sice_IRR_reg[8]/P0001 , \sice_IRR_reg[9]/P0001 , \sice_IRST_reg/NET0131 , \sice_IRST_syn_reg/P0001 , \sice_ITR_reg[0]/NET0131 , \sice_ITR_reg[1]/NET0131 , \sice_ITR_reg[2]/NET0131 , \sice_OE_reg/P0001 , \sice_RCS_reg[0]/NET0131 , \sice_RCS_reg[1]/NET0131 , \sice_RST_req_reg/NET0131 , \sice_SPC_reg[0]/P0001 , \sice_SPC_reg[10]/P0001 , \sice_SPC_reg[11]/P0001 , \sice_SPC_reg[12]/P0001 , \sice_SPC_reg[13]/P0001 , \sice_SPC_reg[14]/P0001 , \sice_SPC_reg[15]/P0001 , \sice_SPC_reg[16]/P0001 , \sice_SPC_reg[17]/P0001 , \sice_SPC_reg[18]/P0001 , \sice_SPC_reg[19]/P0001 , \sice_SPC_reg[1]/P0001 , \sice_SPC_reg[20]/P0001 , \sice_SPC_reg[21]/P0001 , \sice_SPC_reg[22]/P0001 , \sice_SPC_reg[23]/P0001 , \sice_SPC_reg[2]/P0001 , \sice_SPC_reg[3]/P0001 , \sice_SPC_reg[4]/P0001 , \sice_SPC_reg[5]/P0001 , \sice_SPC_reg[6]/P0001 , \sice_SPC_reg[7]/P0001 , \sice_SPC_reg[8]/P0001 , \sice_SPC_reg[9]/P0001 , \sice_UpdDR_sd1_reg/P0001 , \sice_UpdDR_sd2_reg/P0001 , \sice_idr0_reg_DO_reg[0]/P0001 , \sice_idr0_reg_DO_reg[10]/P0001 , \sice_idr0_reg_DO_reg[11]/P0001 , \sice_idr0_reg_DO_reg[1]/P0001 , \sice_idr0_reg_DO_reg[2]/P0001 , \sice_idr0_reg_DO_reg[3]/P0001 , \sice_idr0_reg_DO_reg[4]/P0001 , \sice_idr0_reg_DO_reg[5]/P0001 , \sice_idr0_reg_DO_reg[6]/P0001 , \sice_idr0_reg_DO_reg[7]/P0001 , \sice_idr0_reg_DO_reg[8]/P0001 , \sice_idr0_reg_DO_reg[9]/P0001 , \sice_idr1_reg_DO_reg[0]/P0001 , \sice_idr1_reg_DO_reg[10]/P0001 , \sice_idr1_reg_DO_reg[11]/P0001 , \sice_idr1_reg_DO_reg[1]/P0001 , \sice_idr1_reg_DO_reg[2]/P0001 , \sice_idr1_reg_DO_reg[3]/P0001 , \sice_idr1_reg_DO_reg[4]/P0001 , \sice_idr1_reg_DO_reg[5]/P0001 , \sice_idr1_reg_DO_reg[6]/P0001 , \sice_idr1_reg_DO_reg[7]/P0001 , \sice_idr1_reg_DO_reg[8]/P0001 , \sice_idr1_reg_DO_reg[9]/P0001 , \sport0_cfg_FSi_cnt_reg[0]/NET0131 , \sport0_cfg_FSi_cnt_reg[10]/NET0131 , \sport0_cfg_FSi_cnt_reg[11]/NET0131 , \sport0_cfg_FSi_cnt_reg[12]/NET0131 , \sport0_cfg_FSi_cnt_reg[13]/NET0131 , \sport0_cfg_FSi_cnt_reg[14]/NET0131 , \sport0_cfg_FSi_cnt_reg[15]/NET0131 , \sport0_cfg_FSi_cnt_reg[1]/NET0131 , \sport0_cfg_FSi_cnt_reg[2]/NET0131 , \sport0_cfg_FSi_cnt_reg[3]/NET0131 , \sport0_cfg_FSi_cnt_reg[4]/NET0131 , \sport0_cfg_FSi_cnt_reg[5]/NET0131 , \sport0_cfg_FSi_cnt_reg[6]/NET0131 , \sport0_cfg_FSi_cnt_reg[7]/NET0131 , \sport0_cfg_FSi_cnt_reg[8]/NET0131 , \sport0_cfg_FSi_cnt_reg[9]/NET0131 , \sport0_cfg_FSi_reg/NET0131 , \sport0_cfg_RFSg_d1_reg/NET0131 , \sport0_cfg_RFSg_d2_reg/NET0131 , \sport0_cfg_RFSg_d3_reg/NET0131 , \sport0_cfg_RFSgi_d_reg/NET0131 , \sport0_cfg_SCLKi_cnt_reg[0]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[10]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[11]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[12]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[13]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[14]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[15]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[1]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[2]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[3]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[4]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[5]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[6]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[7]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[8]/NET0131 , \sport0_cfg_SCLKi_cnt_reg[9]/NET0131 , \sport0_cfg_SCLKi_h_reg/NET0131 , \sport0_cfg_SP_ENg_D1_reg/P0001 , \sport0_cfg_SP_ENg_reg/NET0131 , \sport0_cfg_TFSg_d1_reg/NET0131 , \sport0_cfg_TFSg_d2_reg/NET0131 , \sport0_cfg_TFSg_d3_reg/NET0131 , \sport0_cfg_TFSgi_d_reg/NET0131 , \sport0_regs_AUTO_a_reg[12]/NET0131 , \sport0_regs_AUTO_a_reg[13]/NET0131 , \sport0_regs_AUTO_a_reg[14]/NET0131 , \sport0_regs_AUTO_a_reg[15]/NET0131 , \sport0_regs_AUTOreg_DO_reg[0]/NET0131 , \sport0_regs_AUTOreg_DO_reg[10]/NET0131 , \sport0_regs_AUTOreg_DO_reg[11]/NET0131 , \sport0_regs_AUTOreg_DO_reg[1]/NET0131 , \sport0_regs_AUTOreg_DO_reg[2]/NET0131 , \sport0_regs_AUTOreg_DO_reg[3]/NET0131 , \sport0_regs_AUTOreg_DO_reg[4]/NET0131 , \sport0_regs_AUTOreg_DO_reg[5]/NET0131 , \sport0_regs_AUTOreg_DO_reg[6]/NET0131 , \sport0_regs_AUTOreg_DO_reg[7]/NET0131 , \sport0_regs_AUTOreg_DO_reg[8]/NET0131 , \sport0_regs_AUTOreg_DO_reg[9]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[0]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[10]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[11]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[12]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[13]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[14]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[15]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[1]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[2]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[3]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[4]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[5]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[6]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[7]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[8]/NET0131 , \sport0_regs_FSDIVreg_DO_reg[9]/NET0131 , \sport0_regs_MWORDreg_DO_reg[0]/NET0131 , \sport0_regs_MWORDreg_DO_reg[10]/NET0131 , \sport0_regs_MWORDreg_DO_reg[1]/NET0131 , \sport0_regs_MWORDreg_DO_reg[2]/NET0131 , \sport0_regs_MWORDreg_DO_reg[3]/NET0131 , \sport0_regs_MWORDreg_DO_reg[4]/NET0131 , \sport0_regs_MWORDreg_DO_reg[5]/NET0131 , \sport0_regs_MWORDreg_DO_reg[6]/NET0131 , \sport0_regs_MWORDreg_DO_reg[7]/NET0131 , \sport0_regs_MWORDreg_DO_reg[8]/NET0131 , \sport0_regs_MWORDreg_DO_reg[9]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 , \sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 , \sport0_regs_SCTLreg_DO_reg[0]/NET0131 , \sport0_regs_SCTLreg_DO_reg[10]/NET0131 , \sport0_regs_SCTLreg_DO_reg[11]/NET0131 , \sport0_regs_SCTLreg_DO_reg[12]/NET0131 , \sport0_regs_SCTLreg_DO_reg[13]/NET0131 , \sport0_regs_SCTLreg_DO_reg[15]/NET0131 , \sport0_regs_SCTLreg_DO_reg[1]/NET0131 , \sport0_regs_SCTLreg_DO_reg[2]/NET0131 , \sport0_regs_SCTLreg_DO_reg[3]/NET0131 , \sport0_regs_SCTLreg_DO_reg[4]/NET0131 , \sport0_regs_SCTLreg_DO_reg[5]/NET0131 , \sport0_regs_SCTLreg_DO_reg[6]/NET0131 , \sport0_regs_SCTLreg_DO_reg[7]/NET0131 , \sport0_rxctl_Bcnt_reg[0]/NET0131 , \sport0_rxctl_Bcnt_reg[1]/NET0131 , \sport0_rxctl_Bcnt_reg[2]/NET0131 , \sport0_rxctl_Bcnt_reg[3]/NET0131 , \sport0_rxctl_Bcnt_reg[4]/NET0131 , \sport0_rxctl_ISRa_reg/P0001 , \sport0_rxctl_LMcnt_reg[0]/NET0131 , \sport0_rxctl_LMcnt_reg[1]/NET0131 , \sport0_rxctl_LMcnt_reg[2]/NET0131 , \sport0_rxctl_LMcnt_reg[3]/NET0131 , \sport0_rxctl_LMcnt_reg[4]/NET0131 , \sport0_rxctl_RCS_reg[0]/NET0131 , \sport0_rxctl_RCS_reg[1]/NET0131 , \sport0_rxctl_RCS_reg[2]/NET0131 , \sport0_rxctl_RSreq_reg/NET0131 , \sport0_rxctl_RXSHT_reg[0]/P0001 , \sport0_rxctl_RXSHT_reg[10]/P0001 , \sport0_rxctl_RXSHT_reg[11]/P0001 , \sport0_rxctl_RXSHT_reg[12]/P0001 , \sport0_rxctl_RXSHT_reg[13]/P0001 , \sport0_rxctl_RXSHT_reg[14]/P0001 , \sport0_rxctl_RXSHT_reg[15]/P0001 , \sport0_rxctl_RXSHT_reg[1]/P0001 , \sport0_rxctl_RXSHT_reg[2]/P0001 , \sport0_rxctl_RXSHT_reg[3]/P0001 , \sport0_rxctl_RXSHT_reg[4]/P0001 , \sport0_rxctl_RXSHT_reg[5]/P0001 , \sport0_rxctl_RXSHT_reg[6]/P0001 , \sport0_rxctl_RXSHT_reg[7]/P0001 , \sport0_rxctl_RXSHT_reg[8]/P0001 , \sport0_rxctl_RXSHT_reg[9]/P0001 , \sport0_rxctl_RX_reg[0]/P0001 , \sport0_rxctl_RX_reg[10]/P0001 , \sport0_rxctl_RX_reg[11]/P0001 , \sport0_rxctl_RX_reg[12]/P0001 , \sport0_rxctl_RX_reg[13]/P0001 , \sport0_rxctl_RX_reg[14]/P0001 , \sport0_rxctl_RX_reg[15]/P0001 , \sport0_rxctl_RX_reg[1]/P0001 , \sport0_rxctl_RX_reg[2]/P0001 , \sport0_rxctl_RX_reg[3]/P0001 , \sport0_rxctl_RX_reg[4]/P0001 , \sport0_rxctl_RX_reg[5]/P0001 , \sport0_rxctl_RX_reg[6]/P0001 , \sport0_rxctl_RX_reg[7]/P0001 , \sport0_rxctl_RX_reg[8]/P0001 , \sport0_rxctl_RX_reg[9]/P0001 , \sport0_rxctl_SLOT1_EXT_reg[2]/NET0131 , \sport0_rxctl_SLOT1_EXT_reg[3]/NET0131 , \sport0_rxctl_TAG_SLOT_reg/P0001 , \sport0_rxctl_Wcnt_reg[0]/NET0131 , \sport0_rxctl_Wcnt_reg[1]/NET0131 , \sport0_rxctl_Wcnt_reg[2]/NET0131 , \sport0_rxctl_Wcnt_reg[3]/NET0131 , \sport0_rxctl_Wcnt_reg[4]/NET0131 , \sport0_rxctl_Wcnt_reg[5]/NET0131 , \sport0_rxctl_Wcnt_reg[6]/NET0131 , \sport0_rxctl_Wcnt_reg[7]/NET0131 , \sport0_rxctl_a_sync1_reg/P0001 , \sport0_rxctl_a_sync2_reg/P0001 , \sport0_rxctl_ldRX_cmp_reg/P0001 , \sport0_rxctl_sht2nd_reg/P0001 , \sport0_txctl_Bcnt_reg[0]/NET0131 , \sport0_txctl_Bcnt_reg[1]/NET0131 , \sport0_txctl_Bcnt_reg[2]/NET0131 , \sport0_txctl_Bcnt_reg[3]/NET0131 , \sport0_txctl_Bcnt_reg[4]/NET0131 , \sport0_txctl_SP_EN_D1_reg/P0001 , \sport0_txctl_TCS_reg[0]/NET0131 , \sport0_txctl_TCS_reg[1]/NET0131 , \sport0_txctl_TCS_reg[2]/NET0131 , \sport0_txctl_TSreq_reg/NET0131 , \sport0_txctl_TSreqi_reg/NET0131 , \sport0_txctl_TXSHT_reg[0]/P0001 , \sport0_txctl_TXSHT_reg[10]/P0001 , \sport0_txctl_TXSHT_reg[11]/P0001 , \sport0_txctl_TXSHT_reg[12]/P0001 , \sport0_txctl_TXSHT_reg[13]/P0001 , \sport0_txctl_TXSHT_reg[14]/P0001 , \sport0_txctl_TXSHT_reg[15]/P0001 , \sport0_txctl_TXSHT_reg[1]/P0001 , \sport0_txctl_TXSHT_reg[2]/P0001 , \sport0_txctl_TXSHT_reg[3]/P0001 , \sport0_txctl_TXSHT_reg[4]/P0001 , \sport0_txctl_TXSHT_reg[5]/P0001 , \sport0_txctl_TXSHT_reg[6]/P0001 , \sport0_txctl_TXSHT_reg[7]/P0001 , \sport0_txctl_TXSHT_reg[8]/P0001 , \sport0_txctl_TXSHT_reg[9]/P0001 , \sport0_txctl_TX_reg[0]/P0001 , \sport0_txctl_TX_reg[10]/P0001 , \sport0_txctl_TX_reg[11]/P0001 , \sport0_txctl_TX_reg[12]/P0001 , \sport0_txctl_TX_reg[13]/P0001 , \sport0_txctl_TX_reg[14]/P0001 , \sport0_txctl_TX_reg[15]/P0001 , \sport0_txctl_TX_reg[1]/P0001 , \sport0_txctl_TX_reg[2]/P0001 , \sport0_txctl_TX_reg[3]/P0001 , \sport0_txctl_TX_reg[4]/P0001 , \sport0_txctl_TX_reg[5]/P0001 , \sport0_txctl_TX_reg[6]/P0001 , \sport0_txctl_TX_reg[7]/P0001 , \sport0_txctl_TX_reg[8]/P0001 , \sport0_txctl_TX_reg[9]/P0001 , \sport0_txctl_Wcnt_reg[0]/NET0131 , \sport0_txctl_Wcnt_reg[1]/NET0131 , \sport0_txctl_Wcnt_reg[2]/NET0131 , \sport0_txctl_Wcnt_reg[3]/NET0131 , \sport0_txctl_Wcnt_reg[4]/NET0131 , \sport0_txctl_Wcnt_reg[5]/NET0131 , \sport0_txctl_Wcnt_reg[6]/NET0131 , \sport0_txctl_Wcnt_reg[7]/NET0131 , \sport0_txctl_b_sync1_reg/P0001 , \sport0_txctl_c_sync1_reg/P0001 , \sport0_txctl_c_sync2_reg/P0001 , \sport0_txctl_ldTX_cmp_reg/P0001 , \sport1_cfg_FSi_cnt_reg[0]/NET0131 , \sport1_cfg_FSi_cnt_reg[10]/NET0131 , \sport1_cfg_FSi_cnt_reg[11]/NET0131 , \sport1_cfg_FSi_cnt_reg[12]/NET0131 , \sport1_cfg_FSi_cnt_reg[13]/NET0131 , \sport1_cfg_FSi_cnt_reg[14]/NET0131 , \sport1_cfg_FSi_cnt_reg[15]/NET0131 , \sport1_cfg_FSi_cnt_reg[1]/NET0131 , \sport1_cfg_FSi_cnt_reg[2]/NET0131 , \sport1_cfg_FSi_cnt_reg[3]/NET0131 , \sport1_cfg_FSi_cnt_reg[4]/NET0131 , \sport1_cfg_FSi_cnt_reg[5]/NET0131 , \sport1_cfg_FSi_cnt_reg[6]/NET0131 , \sport1_cfg_FSi_cnt_reg[7]/NET0131 , \sport1_cfg_FSi_cnt_reg[8]/NET0131 , \sport1_cfg_FSi_cnt_reg[9]/NET0131 , \sport1_cfg_FSi_reg/NET0131 , \sport1_cfg_RFSg_d1_reg/NET0131 , \sport1_cfg_RFSg_d2_reg/NET0131 , \sport1_cfg_RFSg_d3_reg/NET0131 , \sport1_cfg_RFSgi_d_reg/NET0131 , \sport1_cfg_SCLKi_cnt_reg[0]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[10]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[11]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[12]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[13]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[14]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[15]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[1]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[2]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[3]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[4]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[5]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[6]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[7]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[8]/NET0131 , \sport1_cfg_SCLKi_cnt_reg[9]/NET0131 , \sport1_cfg_SCLKi_h_reg/NET0131 , \sport1_cfg_SP_ENg_D1_reg/P0001 , \sport1_cfg_SP_ENg_reg/NET0131 , \sport1_cfg_TFSg_d1_reg/NET0131 , \sport1_cfg_TFSg_d2_reg/NET0131 , \sport1_cfg_TFSg_d3_reg/NET0131 , \sport1_cfg_TFSgi_d_reg/NET0131 , \sport1_regs_AUTOreg_DO_reg[0]/NET0131 , \sport1_regs_AUTOreg_DO_reg[10]/NET0131 , \sport1_regs_AUTOreg_DO_reg[11]/NET0131 , \sport1_regs_AUTOreg_DO_reg[1]/NET0131 , \sport1_regs_AUTOreg_DO_reg[2]/NET0131 , \sport1_regs_AUTOreg_DO_reg[3]/NET0131 , \sport1_regs_AUTOreg_DO_reg[4]/NET0131 , \sport1_regs_AUTOreg_DO_reg[5]/NET0131 , \sport1_regs_AUTOreg_DO_reg[6]/NET0131 , \sport1_regs_AUTOreg_DO_reg[7]/NET0131 , \sport1_regs_AUTOreg_DO_reg[8]/NET0131 , \sport1_regs_AUTOreg_DO_reg[9]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[0]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[10]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[11]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[12]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[13]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[14]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[15]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[1]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[2]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[3]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[4]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[5]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[6]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[7]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[8]/NET0131 , \sport1_regs_FSDIVreg_DO_reg[9]/NET0131 , \sport1_regs_MWORDreg_DO_reg[0]/NET0131 , \sport1_regs_MWORDreg_DO_reg[10]/NET0131 , \sport1_regs_MWORDreg_DO_reg[1]/NET0131 , \sport1_regs_MWORDreg_DO_reg[2]/NET0131 , \sport1_regs_MWORDreg_DO_reg[3]/NET0131 , \sport1_regs_MWORDreg_DO_reg[4]/NET0131 , \sport1_regs_MWORDreg_DO_reg[5]/NET0131 , \sport1_regs_MWORDreg_DO_reg[6]/NET0131 , \sport1_regs_MWORDreg_DO_reg[7]/NET0131 , \sport1_regs_MWORDreg_DO_reg[8]/NET0131 , \sport1_regs_MWORDreg_DO_reg[9]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 , \sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 , \sport1_regs_SCTLreg_DO_reg[0]/NET0131 , \sport1_regs_SCTLreg_DO_reg[10]/NET0131 , \sport1_regs_SCTLreg_DO_reg[11]/NET0131 , \sport1_regs_SCTLreg_DO_reg[12]/NET0131 , \sport1_regs_SCTLreg_DO_reg[13]/NET0131 , \sport1_regs_SCTLreg_DO_reg[15]/NET0131 , \sport1_regs_SCTLreg_DO_reg[1]/NET0131 , \sport1_regs_SCTLreg_DO_reg[2]/NET0131 , \sport1_regs_SCTLreg_DO_reg[3]/NET0131 , \sport1_regs_SCTLreg_DO_reg[4]/NET0131 , \sport1_regs_SCTLreg_DO_reg[5]/NET0131 , \sport1_regs_SCTLreg_DO_reg[6]/NET0131 , \sport1_regs_SCTLreg_DO_reg[7]/NET0131 , \sport1_rxctl_Bcnt_reg[0]/NET0131 , \sport1_rxctl_Bcnt_reg[1]/NET0131 , \sport1_rxctl_Bcnt_reg[2]/NET0131 , \sport1_rxctl_Bcnt_reg[3]/NET0131 , \sport1_rxctl_Bcnt_reg[4]/NET0131 , \sport1_rxctl_ISRa_reg/P0001 , \sport1_rxctl_LMcnt_reg[0]/NET0131 , \sport1_rxctl_LMcnt_reg[1]/NET0131 , \sport1_rxctl_LMcnt_reg[2]/NET0131 , \sport1_rxctl_LMcnt_reg[3]/NET0131 , \sport1_rxctl_LMcnt_reg[4]/NET0131 , \sport1_rxctl_RCS_reg[0]/NET0131 , \sport1_rxctl_RCS_reg[1]/NET0131 , \sport1_rxctl_RCS_reg[2]/NET0131 , \sport1_rxctl_RSreq_reg/NET0131 , \sport1_rxctl_RXSHT_reg[0]/P0001 , \sport1_rxctl_RXSHT_reg[10]/P0001 , \sport1_rxctl_RXSHT_reg[11]/P0001 , \sport1_rxctl_RXSHT_reg[12]/P0001 , \sport1_rxctl_RXSHT_reg[13]/P0001 , \sport1_rxctl_RXSHT_reg[14]/P0001 , \sport1_rxctl_RXSHT_reg[15]/P0001 , \sport1_rxctl_RXSHT_reg[1]/P0001 , \sport1_rxctl_RXSHT_reg[2]/P0001 , \sport1_rxctl_RXSHT_reg[3]/P0001 , \sport1_rxctl_RXSHT_reg[4]/P0001 , \sport1_rxctl_RXSHT_reg[5]/P0001 , \sport1_rxctl_RXSHT_reg[6]/P0001 , \sport1_rxctl_RXSHT_reg[7]/P0001 , \sport1_rxctl_RXSHT_reg[8]/P0001 , \sport1_rxctl_RXSHT_reg[9]/P0001 , \sport1_rxctl_RX_reg[0]/P0001 , \sport1_rxctl_RX_reg[10]/P0001 , \sport1_rxctl_RX_reg[11]/P0001 , \sport1_rxctl_RX_reg[12]/P0001 , \sport1_rxctl_RX_reg[13]/P0001 , \sport1_rxctl_RX_reg[14]/P0001 , \sport1_rxctl_RX_reg[15]/P0001 , \sport1_rxctl_RX_reg[1]/P0001 , \sport1_rxctl_RX_reg[2]/P0001 , \sport1_rxctl_RX_reg[3]/P0001 , \sport1_rxctl_RX_reg[4]/P0001 , \sport1_rxctl_RX_reg[5]/P0001 , \sport1_rxctl_RX_reg[6]/P0001 , \sport1_rxctl_RX_reg[7]/P0001 , \sport1_rxctl_RX_reg[8]/P0001 , \sport1_rxctl_RX_reg[9]/P0001 , \sport1_rxctl_SLOT1_EXT_reg[2]/NET0131 , \sport1_rxctl_SLOT1_EXT_reg[3]/NET0131 , \sport1_rxctl_TAG_SLOT_reg/P0001 , \sport1_rxctl_Wcnt_reg[0]/NET0131 , \sport1_rxctl_Wcnt_reg[1]/NET0131 , \sport1_rxctl_Wcnt_reg[2]/NET0131 , \sport1_rxctl_Wcnt_reg[3]/NET0131 , \sport1_rxctl_Wcnt_reg[4]/NET0131 , \sport1_rxctl_Wcnt_reg[5]/NET0131 , \sport1_rxctl_Wcnt_reg[6]/NET0131 , \sport1_rxctl_Wcnt_reg[7]/NET0131 , \sport1_rxctl_a_sync1_reg/P0001 , \sport1_rxctl_a_sync2_reg/P0001 , \sport1_rxctl_sht2nd_reg/P0001 , \sport1_txctl_Bcnt_reg[0]/NET0131 , \sport1_txctl_Bcnt_reg[1]/NET0131 , \sport1_txctl_Bcnt_reg[2]/NET0131 , \sport1_txctl_Bcnt_reg[3]/NET0131 , \sport1_txctl_Bcnt_reg[4]/NET0131 , \sport1_txctl_SP_EN_D1_reg/P0001 , \sport1_txctl_TCS_reg[0]/NET0131 , \sport1_txctl_TCS_reg[1]/NET0131 , \sport1_txctl_TCS_reg[2]/NET0131 , \sport1_txctl_TSreq_reg/NET0131 , \sport1_txctl_TSreqi_reg/NET0131 , \sport1_txctl_TXSHT_reg[0]/P0001 , \sport1_txctl_TXSHT_reg[10]/P0001 , \sport1_txctl_TXSHT_reg[11]/P0001 , \sport1_txctl_TXSHT_reg[12]/P0001 , \sport1_txctl_TXSHT_reg[13]/P0001 , \sport1_txctl_TXSHT_reg[14]/P0001 , \sport1_txctl_TXSHT_reg[15]/P0001 , \sport1_txctl_TXSHT_reg[1]/P0001 , \sport1_txctl_TXSHT_reg[2]/P0001 , \sport1_txctl_TXSHT_reg[3]/P0001 , \sport1_txctl_TXSHT_reg[4]/P0001 , \sport1_txctl_TXSHT_reg[5]/P0001 , \sport1_txctl_TXSHT_reg[6]/P0001 , \sport1_txctl_TXSHT_reg[7]/P0001 , \sport1_txctl_TXSHT_reg[8]/P0001 , \sport1_txctl_TXSHT_reg[9]/P0001 , \sport1_txctl_TX_reg[0]/P0001 , \sport1_txctl_TX_reg[10]/P0001 , \sport1_txctl_TX_reg[11]/P0001 , \sport1_txctl_TX_reg[12]/P0001 , \sport1_txctl_TX_reg[13]/P0001 , \sport1_txctl_TX_reg[14]/P0001 , \sport1_txctl_TX_reg[15]/P0001 , \sport1_txctl_TX_reg[1]/P0001 , \sport1_txctl_TX_reg[2]/P0001 , \sport1_txctl_TX_reg[3]/P0001 , \sport1_txctl_TX_reg[4]/P0001 , \sport1_txctl_TX_reg[5]/P0001 , \sport1_txctl_TX_reg[6]/P0001 , \sport1_txctl_TX_reg[7]/P0001 , \sport1_txctl_TX_reg[8]/P0001 , \sport1_txctl_TX_reg[9]/P0001 , \sport1_txctl_Wcnt_reg[0]/NET0131 , \sport1_txctl_Wcnt_reg[1]/NET0131 , \sport1_txctl_Wcnt_reg[2]/NET0131 , \sport1_txctl_Wcnt_reg[3]/NET0131 , \sport1_txctl_Wcnt_reg[4]/NET0131 , \sport1_txctl_Wcnt_reg[5]/NET0131 , \sport1_txctl_Wcnt_reg[6]/NET0131 , \sport1_txctl_Wcnt_reg[7]/NET0131 , \sport1_txctl_c_sync1_reg/P0001 , \sport1_txctl_c_sync2_reg/P0001 , \tm_MSTAT5_syn_reg/NET0131 , \tm_TCR_TMP_reg[0]/NET0131 , \tm_TCR_TMP_reg[10]/NET0131 , \tm_TCR_TMP_reg[11]/NET0131 , \tm_TCR_TMP_reg[12]/NET0131 , \tm_TCR_TMP_reg[13]/NET0131 , \tm_TCR_TMP_reg[14]/NET0131 , \tm_TCR_TMP_reg[15]/NET0131 , \tm_TCR_TMP_reg[1]/NET0131 , \tm_TCR_TMP_reg[2]/NET0131 , \tm_TCR_TMP_reg[3]/NET0131 , \tm_TCR_TMP_reg[4]/NET0131 , \tm_TCR_TMP_reg[5]/NET0131 , \tm_TCR_TMP_reg[6]/NET0131 , \tm_TCR_TMP_reg[7]/NET0131 , \tm_TCR_TMP_reg[8]/NET0131 , \tm_TCR_TMP_reg[9]/NET0131 , \tm_TINT_GEN1_reg/NET0131 , \tm_TINT_GEN2_reg/NET0131 , \tm_TSR_TMP_reg[0]/NET0131 , \tm_TSR_TMP_reg[1]/NET0131 , \tm_TSR_TMP_reg[2]/NET0131 , \tm_TSR_TMP_reg[3]/NET0131 , \tm_TSR_TMP_reg[4]/NET0131 , \tm_TSR_TMP_reg[5]/NET0131 , \tm_TSR_TMP_reg[6]/NET0131 , \tm_TSR_TMP_reg[7]/NET0131 , \tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131 , \tm_WR_TCR_TMP_GEN1_reg/P0001 , \tm_WR_TCR_TMP_GEN2_reg/P0001 , \tm_WR_TCR_p_reg/P0001 , \tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131 , \tm_WR_TSR_TMP_GEN1_reg/P0001 , \tm_WR_TSR_TMP_GEN2_reg/P0001 , \tm_WR_TSR_p_reg/P0001 , \tm_tcr_reg_DO_reg[0]/NET0131 , \tm_tcr_reg_DO_reg[10]/NET0131 , \tm_tcr_reg_DO_reg[11]/NET0131 , \tm_tcr_reg_DO_reg[12]/NET0131 , \tm_tcr_reg_DO_reg[13]/NET0131 , \tm_tcr_reg_DO_reg[14]/NET0131 , \tm_tcr_reg_DO_reg[15]/NET0131 , \tm_tcr_reg_DO_reg[1]/NET0131 , \tm_tcr_reg_DO_reg[2]/NET0131 , \tm_tcr_reg_DO_reg[3]/NET0131 , \tm_tcr_reg_DO_reg[4]/NET0131 , \tm_tcr_reg_DO_reg[5]/NET0131 , \tm_tcr_reg_DO_reg[6]/NET0131 , \tm_tcr_reg_DO_reg[7]/NET0131 , \tm_tcr_reg_DO_reg[8]/NET0131 , \tm_tcr_reg_DO_reg[9]/NET0131 , \tm_tpr_reg_DO_reg[0]/NET0131 , \tm_tpr_reg_DO_reg[10]/NET0131 , \tm_tpr_reg_DO_reg[11]/NET0131 , \tm_tpr_reg_DO_reg[12]/NET0131 , \tm_tpr_reg_DO_reg[13]/NET0131 , \tm_tpr_reg_DO_reg[14]/NET0131 , \tm_tpr_reg_DO_reg[15]/NET0131 , \tm_tpr_reg_DO_reg[1]/NET0131 , \tm_tpr_reg_DO_reg[2]/NET0131 , \tm_tpr_reg_DO_reg[3]/NET0131 , \tm_tpr_reg_DO_reg[4]/NET0131 , \tm_tpr_reg_DO_reg[5]/NET0131 , \tm_tpr_reg_DO_reg[6]/NET0131 , \tm_tpr_reg_DO_reg[7]/NET0131 , \tm_tpr_reg_DO_reg[8]/NET0131 , \tm_tpr_reg_DO_reg[9]/NET0131 , \tm_tsr_reg_DO_reg[0]/NET0131 , \tm_tsr_reg_DO_reg[1]/NET0131 , \tm_tsr_reg_DO_reg[2]/NET0131 , \tm_tsr_reg_DO_reg[3]/NET0131 , \tm_tsr_reg_DO_reg[4]/NET0131 , \tm_tsr_reg_DO_reg[5]/NET0131 , \tm_tsr_reg_DO_reg[6]/NET0131 , \tm_tsr_reg_DO_reg[7]/NET0131 , \tm_tsr_reg_DO_reg[8]/NET0131 , CLKO_pad, \CMAinx[0]_pad , \CMAinx[10]_pad , \CMAinx[11]_pad , \CMAinx[1]_pad , \CMAinx[2]_pad , \CMAinx[3]_pad , \CMAinx[4]_pad , \CMAinx[5]_pad , \CMAinx[6]_pad , \CMAinx[7]_pad , \CMAinx[8]_pad , \CMAinx[9]_pad , CMSn_pad, CM_cs_pad, \CM_wd[0]_pad , \CM_wd[10]_pad , \CM_wd[11]_pad , \CM_wd[12]_pad , \CM_wd[13]_pad , \CM_wd[14]_pad , \CM_wd[15]_pad , \CM_wd[16]_pad , \CM_wd[17]_pad , \CM_wd[18]_pad , \CM_wd[19]_pad , \CM_wd[1]_pad , \CM_wd[20]_pad , \CM_wd[21]_pad , \CM_wd[22]_pad , \CM_wd[23]_pad , \CM_wd[2]_pad , \CM_wd[3]_pad , \CM_wd[4]_pad , \CM_wd[5]_pad , \CM_wd[6]_pad , \CM_wd[7]_pad , \CM_wd[8]_pad , \CM_wd[9]_pad , CM_web_pad, \CMo_cs0_pad , \CMo_cs1_pad , \CMo_cs2_pad , \CMo_cs3_pad , \CMo_cs4_pad , \CMo_cs5_pad , \CMo_cs6_pad , \CMo_cs7_pad , \DMAinx[0]_pad , \DMAinx[10]_pad , \DMAinx[11]_pad , \DMAinx[12]_pad , \DMAinx[13]_pad , \DMAinx[1]_pad , \DMAinx[2]_pad , \DMAinx[3]_pad , \DMAinx[4]_pad , \DMAinx[5]_pad , \DMAinx[6]_pad , \DMAinx[7]_pad , \DMAinx[8]_pad , \DMAinx[9]_pad , DMSn_pad, DM_cs_pad, \DM_wd[0]_pad , \DM_wd[10]_pad , \DM_wd[11]_pad , \DM_wd[12]_pad , \DM_wd[13]_pad , \DM_wd[14]_pad , \DM_wd[15]_pad , \DM_wd[1]_pad , \DM_wd[2]_pad , \DM_wd[3]_pad , \DM_wd[4]_pad , \DM_wd[5]_pad , \DM_wd[6]_pad , \DM_wd[7]_pad , \DM_wd[8]_pad , \DM_wd[9]_pad , \DMo_cs0_pad , \DMo_cs1_pad , \DMo_cs2_pad , \DMo_cs3_pad , \DMo_cs4_pad , \DMo_cs5_pad , \DMo_cs6_pad , \DMo_cs7_pad , \DSPCLK_cm1_pad , \EA_do[0]_pad , \EA_do[10]_pad , \EA_do[12]_pad , \EA_do[13]_pad , \EA_do[14]_pad , \EA_do[1]_pad , \EA_do[2]_pad , \EA_do[3]_pad , \EA_do[4]_pad , \EA_do[5]_pad , \EA_do[6]_pad , \EA_do[7]_pad , \EA_do[8]_pad , \EA_do[9]_pad , EA_oe_pad, \ED_do[0]_pad , \ED_do[10]_pad , \ED_do[11]_pad , \ED_do[12]_pad , \ED_do[13]_pad , \ED_do[14]_pad , \ED_do[15]_pad , \ED_do[1]_pad , \ED_do[2]_pad , \ED_do[3]_pad , \ED_do[4]_pad , \ED_do[5]_pad , \ED_do[6]_pad , \ED_do[7]_pad , \ED_do[8]_pad , \ED_do[9]_pad , \ED_oe_14_8_pad , \ED_oe_7_0_pad , \IAD_do[0]_pad , \IAD_do[10]_pad , \IAD_do[11]_pad , \IAD_do[12]_pad , \IAD_do[13]_pad , \IAD_do[14]_pad , \IAD_do[15]_pad , \IAD_do[1]_pad , \IAD_do[2]_pad , \IAD_do[3]_pad , \IAD_do[4]_pad , \IAD_do[5]_pad , \IAD_do[6]_pad , \IAD_do[7]_pad , \IAD_do[8]_pad , \IAD_do[9]_pad , IAD_oe_pad, IDoe_pad, IOSn_pad, \PMAinx[0]_pad , \PMAinx[10]_pad , \PMAinx[11]_pad , \PMAinx[1]_pad , \PMAinx[2]_pad , \PMAinx[3]_pad , \PMAinx[4]_pad , \PMAinx[5]_pad , \PMAinx[6]_pad , \PMAinx[7]_pad , \PMAinx[8]_pad , \PMAinx[9]_pad , \PM_wd[0]_pad , \PM_wd[10]_pad , \PM_wd[11]_pad , \PM_wd[12]_pad , \PM_wd[13]_pad , \PM_wd[14]_pad , \PM_wd[15]_pad , \PM_wd[1]_pad , \PM_wd[2]_pad , \PM_wd[3]_pad , \PM_wd[4]_pad , \PM_wd[5]_pad , \PM_wd[6]_pad , \PM_wd[7]_pad , \PM_wd[8]_pad , \PM_wd[9]_pad , \PMo_cs0_pad , \PMo_cs1_pad , \PMo_cs2_pad , \PMo_cs3_pad , \PMo_cs4_pad , \PMo_cs5_pad , \PMo_cs6_pad , \PMo_cs7_pad , \PMo_oe0_pad , \RFS0_pad , \RFS1_pad , \SCLK0_pad , \SCLK1_pad , \TD0_pad , \TD1_pad , \TFS0_pad , \TFS1_pad , \T_ISn_syn_2 , WRn_pad, XTALoffn_pad, \_al_n0 , \bdma_BDMA_boot_reg/NET0131_reg_syn_3 , \bdma_BDMA_boot_reg/n0 , \bdma_BM_cyc_reg/P0000 , \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3 , \core_c_psq_MGNT_reg/P0001 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3 , \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3 , \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3 , \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3 , \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3 , \emc_DMDreg_reg[8]/P0001_reg_syn_3 , \emc_DMDreg_reg[9]/P0001_reg_syn_3 , \emc_ECMcs_reg/P0001 , \emc_PMDreg_reg[8]/P0001_reg_syn_3 , \emc_PMDreg_reg[9]/P0001_reg_syn_3 , \g10/_0_ , \g1000/_0_ , \g10000/_0_ , \g10001/_0_ , \g10002/_0_ , \g10003/_0_ , \g10004/_0_ , \g10005/_0_ , \g10007/_0_ , \g10008/_0_ , \g10009/_0_ , \g1001/_3_ , \g10010/_0_ , \g10011/_0_ , \g10012/_0_ , \g10013/_0_ , \g10014/_0_ , \g10015/_0_ , \g10016/_0_ , \g10017/_0_ , \g10018/_0_ , \g10019/_0_ , \g1002/_3_ , \g10020/_0_ , \g10021/_0_ , \g10022/_0_ , \g10023/_0_ , \g10024/_0_ , \g10025/_0_ , \g10026/_0_ , \g10027/_0_ , \g10028/_0_ , \g10029/_0_ , \g1003/_0_ , \g10030/_0_ , \g10031/_0_ , \g10032/_0_ , \g10033/_0_ , \g10034/_0_ , \g10035/_0_ , \g10036/_0_ , \g10037/_0_ , \g10038/_0_ , \g10039/_0_ , \g10040/_0_ , \g10041/_0_ , \g10042/_0_ , \g10043/_0_ , \g10044/_0_ , \g10045/_0_ , \g10046/_0_ , \g10047/_0_ , \g10048/_0_ , \g10049/_0_ , \g10050/_0_ , \g10051/_0_ , \g10052/_0_ , \g10053/_0_ , \g10054/_0_ , \g10055/_0_ , \g10056/_0_ , \g10057/_0_ , \g10058/_0_ , \g10059/_0_ , \g10060/_0_ , \g10061/_0_ , \g10062/_0_ , \g10063/_0_ , \g10064/_0_ , \g10065/_0_ , \g10066/_0_ , \g10067/_0_ , \g10068/_0_ , \g10069/_0_ , \g10070/_0_ , \g10071/_0_ , \g10072/_0_ , \g10073/_0_ , \g10074/_0_ , \g10075/_0_ , \g10076/_0_ , \g10077/_0_ , \g10078/_0_ , \g10080/_0_ , \g10081/_0_ , \g10083/_0_ , \g10089/_0_ , \g1009/_0_ , \g10090/_0_ , \g10091/_0_ , \g10092/_0_ , \g10093/_0_ , \g10094/_0_ , \g1010/_0_ , \g10108/_3_ , \g1011/_0_ , \g10110/_0_ , \g10111/_0_ , \g10113/_3_ , \g10115/_3_ , \g1013/_0_ , \g1014/_0_ , \g10152/_0_ , \g10153/_0_ , \g10154/_0_ , \g10155/_0_ , \g10156/_0_ , \g10157/_0_ , \g10158/_0_ , \g10159/_0_ , \g1016/_0_ , \g10160/_0_ , \g10161/_0_ , \g10162/_0_ , \g10163/_0_ , \g10164/_0_ , \g10165/_0_ , \g1017/_0_ , \g10170/_3_ , \g1018/_0_ , \g10190/_3_ , \g10194/_3_ , \g10198/_0_ , \g10199/_0_ , \g102/_0_ , \g103/_0_ , \g104/_0_ , \g105/_0_ , \g10598/_0_ , \g106/_0_ , \g10667/_0_ , \g10683/_0_ , \g10685/_0_ , \g107/_0_ , \g10721/_0_ , \g10758/_0_ , \g10765/_0_ , \g10778/_0_ , \g10791/_0_ , \g108/_0_ , \g10887/_0_ , \g1089/_0_ , \g109/_0_ , \g1090/_0_ , \g1091/_0_ , \g1092/_0_ , \g10923/_0_ , \g1093/_0_ , \g10930/_0_ , \g10931/_0_ , \g10936/_0_ , \g1097/_0_ , \g11/_0_ , \g110/_0_ , \g1101/_0_ , \g11013/_0_ , \g1102/_0_ , \g1103/_0_ , \g11032/_0_ , \g1104/_0_ , \g1105/_0_ , \g1107/_0_ , \g11074/_0_ , \g11077/_0_ , \g1108/_0_ , \g1109/_0_ , \g11112/_0_ , \g11115/_0_ , \g11116/_0_ , \g11119/_0_ , \g11120/_0_ , \g1113/_0_ , \g1115/_0_ , \g1116/_0_ , \g1117/_0_ , \g11267/_0_ , \g11281/_0_ , \g11287/_0_ , \g11300/_0_ , \g11323/_0_ , \g11325/_2__syn_2 , \g11345/_2_ , \g11470/_0_ , \g11471/_0_ , \g11472/_0_ , \g11473/_0_ , \g11474/_0_ , \g11476/_0_ , \g11477/_0_ , \g11496/_0_ , \g11497/_0_ , \g11498/_0_ , \g11499/_0_ , \g11500/_0_ , \g11501/_0_ , \g11502/_0_ , \g11503/_0_ , \g11504/_0_ , \g11505/_0_ , \g11506/_0_ , \g11507/_0_ , \g11509/_0_ , \g11510/_0_ , \g11515/_0_ , \g11516/_0_ , \g11520/_0_ , \g11521/_0_ , \g11576/_0_ , \g11577/_0_ , \g11578/_0_ , \g11579/_0_ , \g11580/_0_ , \g11581/_0_ , \g11582/_0_ , \g11583/_0_ , \g11584/_0_ , \g11585/_0_ , \g11586/_0_ , \g11587/_0_ , \g11588/_0_ , \g11589/_0_ , \g11591/_0_ , \g11593/_0_ , \g11595/_0_ , \g11596/_0_ , \g11597/_0_ , \g11605/_0_ , \g11606/_0_ , \g11607/_0_ , \g11608/_0_ , \g11609/_0_ , \g11610/_0_ , \g11611/_0_ , \g11612/_0_ , \g11613/_0_ , \g11615/_0_ , \g11616/_0_ , \g11617/_0_ , \g11651/_3_ , \g11704/_0_ , \g11705/_0_ , \g11709/_0_ , \g11722/_0_ , \g11723/_0_ , \g119/_0_ , \g1192/_0_ , \g11994/_0_ , \g120/_0_ , \g1200/_0_ , \g12003/_0_ , \g1201/_0_ , \g12019/_0_ , \g1203/_3_ , \g1204/_3_ , \g1207/_0_ , \g1208/_0_ , \g12092/_0_ , \g1210/_0_ , \g1211/_0_ , \g1212/_0_ , \g1213/_0_ , \g12145/_0_ , \g12155/_0_ , \g12186/_0_ , \g12187/_0_ , \g12192/_0_ , \g12201/_0_ , \g12202/_0_ , \g12203/_0_ , \g12204/_0_ , \g12207/_0_ , \g12229/_3_ , \g12267/_0_ , \g12276/_0_ , \g12278/_0_ , \g12279/_0_ , \g12280/_0_ , \g12302/_0_ , \g12316/_0_ , \g12317/_0_ , \g12319/_0_ , \g12328/_3_ , \g1233/_0_ , \g12348/_0_ , \g12351/_0_ , \g12352/_0_ , \g12353/_0_ , \g12354/_0_ , \g12355/_0_ , \g1237/_0_ , \g124/_0_ , \g12444/_0_ , \g125/_0_ , \g12637/_0_ , \g12639/_0_ , \g12658/_0_ , \g12659/_0_ , \g12660/_0_ , \g12663/_0_ , \g12664/_0_ , \g12665/_0_ , \g12672/_3_ , \g12673/_3_ , \g12674/_3_ , \g12675/_3_ , \g12676/_3_ , \g12677/_3_ , \g12678/_0_ , \g12679/_3_ , \g12697/_3_ , \g12701/_3_ , \g12711/_2_ , \g12713/_2_ , \g12715/_2_ , \g12717/_2_ , \g12718/_2__syn_2 , \g1272/_0_ , \g12728/_1__syn_2 , \g12730/_3_ , \g12741/_1__syn_2 , \g12746/_0__syn_2 , \g12748/_0_ , \g12749/_0_ , \g12759/_1__syn_2 , \g12760/_0_ , \g12762/_0_ , \g12763/_0_ , \g12764/_0_ , \g12765/_0_ , \g12766/_0_ , \g12767/_0_ , \g12768/_0_ , \g12769/_0_ , \g12770/_0_ , \g12771/_0_ , \g12772/_0_ , \g12773/_0_ , \g12774/_0_ , \g12775/_0_ , \g12776/_0_ , \g12777/_0_ , \g12778/_0_ , \g12779/_0_ , \g1278/_0_ , \g12780/_0_ , \g12781/_0_ , \g12782/_0_ , \g12783/_0_ , \g12784/_0_ , \g12785/_0_ , \g12786/_0_ , \g12787/_0_ , \g12788/_0_ , \g12789/_0_ , \g12790/_0_ , \g12791/_0_ , \g12792/_0_ , \g12793/_0_ , \g12794/_0_ , \g12795/_0_ , \g12796/_0_ , \g12797/_0_ , \g12798/_0_ , \g12799/_0_ , \g12800/_0_ , \g12801/_0_ , \g12802/_0_ , \g12803/_0_ , \g12804/_0_ , \g12805/_0_ , \g12806/_0_ , \g12807/_0_ , \g12808/_0_ , \g12809/_0_ , \g1281/_0_ , \g12810/_0_ , \g12811/_0_ , \g12812/_0_ , \g12813/_0_ , \g12814/_0_ , \g12815/_0_ , \g12816/_0_ , \g12817/_0_ , \g12818/_0_ , \g12819/_0_ , \g1282/_0_ , \g12820/_0_ , \g12821/_0_ , \g12822/_0_ , \g12823/_0_ , \g12824/_0_ , \g12825/_0_ , \g12826/_0_ , \g12827/_0_ , \g12828/_0_ , \g12829/_0_ , \g12830/_0_ , \g12831/_0_ , \g12832/_0_ , \g12833/_0_ , \g12835/_0_ , \g12836/_0_ , \g12838/_0_ , \g12848/_0_ , \g12849/_0_ , \g1285/_0_ , \g12850/_0_ , \g12857/_0_ , \g12858/_0_ , \g12859/_0_ , \g12861/_0_ , \g12862/_0_ , \g12868/_0_ , \g12869/_0_ , \g1287/_0_ , \g12870/_0_ , \g12871/_0_ , \g12872/_0_ , \g12873/_0_ , \g12874/_0_ , \g12875/_0_ , \g12876/_0_ , \g12877/_0_ , \g12878/_0_ , \g12879/_0_ , \g12880/_0_ , \g12881/_0_ , \g12882/_0_ , \g12883/_0_ , \g12884/_0_ , \g12885/_0_ , \g12886/_0_ , \g12887/_0_ , \g12888/_0_ , \g12889/_0_ , \g1289/_0_ , \g12890/_0_ , \g12891/_0_ , \g12894/_0_ , \g12898/_0_ , \g12899/_0_ , \g12900/_0_ , \g12901/_0_ , \g12902/_0_ , \g12903/_0_ , \g12906/_0_ , \g12907/_0_ , \g12908/_0_ , \g12912/_0_ , \g12913/_0_ , \g12914/_0_ , \g12915/_0_ , \g12916/_0_ , \g12917/_0_ , \g12918/_0_ , \g12919/_0_ , \g12920/_0_ , \g12921/_0_ , \g12922/_0_ , \g12923/_0_ , \g12924/_0_ , \g12925/_0_ , \g12926/_0_ , \g12932/_0_ , \g12933/_0_ , \g12936/_0_ , \g12955/_0_ , \g13015/_0_ , \g13016/_0_ , \g13017/_0_ , \g13018/_0_ , \g13019/_0_ , \g13020/_0_ , \g13021/_0_ , \g13024/_0_ , \g13025/_0_ , \g13027/_0_ , \g13028/_0_ , \g13030/_0_ , \g13031/_0_ , \g13033/_0_ , \g13047/_0_ , \g13060/_0_ , \g13062/_0_ , \g13063/_0_ , \g13064/_0_ , \g13067/_0_ , \g13068/_0_ , \g13069/_0_ , \g13070/_0_ , \g13072/_0_ , \g13094/_0_ , \g13104/_0_ , \g13110/_0_ , \g13114/_0_ , \g13115/_0_ , \g13116/_0_ , \g13117/_0_ , \g13118/_0_ , \g13119/_0_ , \g13120/_0_ , \g13121/_0_ , \g13124/_0_ , \g13125/_0_ , \g13127/_0_ , \g13128/_0_ , \g13129/_0_ , \g13130/_0_ , \g13131/_0_ , \g13132/_0_ , \g13133/_0_ , \g13134/_0_ , \g13138/_0_ , \g13139/_0_ , \g13140/_0_ , \g13141/_0_ , \g13142/_0_ , \g13143/_0_ , \g13144/_0_ , \g13146/_0_ , \g13150/_0_ , \g13152/_0_ , \g13154/_0_ , \g13155/_0_ , \g13156/_0_ , \g13157/_0_ , \g13158/_0_ , \g1320/_3_ , \g13266/_0_ , \g13269/_0_ , \g13274/_0_ , \g13277/_0_ , \g13280/_0_ , \g13283/_0_ , \g13294/_0_ , \g13330/_0_ , \g13333/_0_ , \g13334/_0_ , \g13335/_0_ , \g13336/_0_ , \g13337/_0_ , \g13338/_0_ , \g13345/_0_ , \g13346/_0_ , \g13347/_0_ , \g13348/_0_ , \g13349/_0_ , \g13350/_0_ , \g13351/_0_ , \g13352/_0_ , \g13486/_0_ , \g13488/_0_ , \g13508/_0_ , \g13509/_0_ , \g13510/_0_ , \g13511/_0_ , \g13512/_0_ , \g13513/_0_ , \g13514/_0_ , \g13515/_0_ , \g13516/_0_ , \g13517/_0_ , \g13518/_0_ , \g13519/_0_ , \g13520/_0_ , \g13521/_0_ , \g13540/_0_ , \g13541/_0_ , \g13542/_0_ , \g13543/_0_ , \g13544/_0_ , \g13545/_0_ , \g13546/_0_ , \g13547/_0_ , \g13548/_0_ , \g13549/_0_ , \g13550/_0_ , \g13551/_0_ , \g13552/_0_ , \g13553/_0_ , \g13554/_0_ , \g13555/_0_ , \g13556/_0_ , \g13557/_0_ , \g13558/_0_ , \g13559/_0_ , \g13560/_0_ , \g13561/_0_ , \g13562/_0_ , \g13563/_0_ , \g13564/_0_ , \g13565/_0_ , \g13566/_0_ , \g13567/_0_ , \g13568/_0_ , \g13569/_0_ , \g13570/_0_ , \g13571/_0_ , \g13572/_0_ , \g137/_3_ , \g1387/_3_ , \g1388/_3_ , \g1389/_0_ , \g139/_0_ , \g1390/_0_ , \g1393/_0_ , \g140/_0_ , \g141/_0_ , \g14173/_0_ , \g14176/_0_ , \g142/_3_ , \g14273/_1__syn_2 , \g14274/_0_ , \g14280/_0_ , \g14281/_0_ , \g143/_3_ , \g14354/_3__syn_2 , \g14370/_0_ , \g14385/_0_ , \g14386/_0_ , \g144/_3_ , \g14407/_0_ , \g14412/_0_ , \g14435/_0_ , \g14439/_0_ , \g145/_0_ , \g14522/_0_ , \g14528/_0_ , \g14533/_0_ , \g14581/_1_ , \g14582/_0_ , \g146/_3_ , \g14671/_0_ , \g14672/_0_ , \g147/_0_ , \g1473/_0_ , \g148/_0_ , \g14826/_0_ , \g149/_0_ , \g14908/_0_ , \g14911/_0_ , \g14936/_2_ , \g1494/_0_ , \g1495/_0_ , \g14950/_2_ , \g14953/_2_ , \g15003/_0_ , \g15004/_0_ , \g15006/_0_ , \g15007/_0_ , \g15008/_0_ , \g15009/_0_ , \g15010/_0_ , \g15011/_0_ , \g15012/_0_ , \g15013/_0_ , \g15014/_0_ , \g15015/_0_ , \g15016/_0_ , \g15017/_0_ , \g15018/_0_ , \g15019/_0_ , \g15035/_0_ , \g15036/_0_ , \g15038/_0_ , \g15039/_0_ , \g15040/_0_ , \g15041/_0_ , \g15042/_0_ , \g15043/_0_ , \g15044/_0_ , \g15045/_0_ , \g15046/_0_ , \g15056/_00_ , \g151/_0_ , \g15193/_0_ , \g152/_0_ , \g15256/_0_ , \g153/_0_ , \g15393/_0_ , \g15394/_0_ , \g15395/_0_ , \g15396/_0_ , \g15397/_0_ , \g15398/_0_ , \g15399/_0_ , \g154/_0_ , \g15400/_0_ , \g15401/_0_ , \g15402/_0_ , \g15403/_0_ , \g15404/_0_ , \g15405/_0_ , \g15406/_0_ , \g15407/_0_ , \g15408/_0_ , \g15473/_0_ , \g15650/_0_ , \g15651/_0_ , \g15652/_0_ , \g15653/_0_ , \g15662/_0_ , \g15663/_0_ , \g15664/_0_ , \g15665/_0_ , \g15666/_0_ , \g15667/_0_ , \g15668/_0_ , \g15669/_0_ , \g15670/_0_ , \g15671/_0_ , \g15672/_0_ , \g15673/_0_ , \g15674/_0_ , \g15675/_0_ , \g1569/_0_ , \g1570/_0_ , \g1575/_0_ , \g1576/_0_ , \g15922/_1_ , \g15970/_0_ , \g16059/_0_ , \g1606/_3_ , \g16124/_0_ , \g16144/_0_ , \g16202/_0_ , \g16214/_0_ , \g16247/_0_ , \g16257/_0_ , \g16274/_1_ , \g16324/_0_ , \g16343/_1__syn_2 , \g16381/_0_ , \g16383/_0_ , \g16386/_0_ , \g16414/_1__syn_2 , \g16416/_0__syn_2 , \g16448/_0_ , \g16460/_1_ , \g16625/_3_ , \g16662/_0_ , \g16668/_1__syn_2 , \g16692/_0_ , \g16721/_0_ , \g16723/_0_ , \g16725/_0_ , \g16726/_0_ , \g16727/_0_ , \g16728/_0_ , \g16729/_0_ , \g16730/_0_ , \g16731/_0_ , \g16732/_0_ , \g16733/_0_ , \g16734/_0_ , \g16735/_0_ , \g16736/_0_ , \g16737/_0_ , \g16738/_0_ , \g16739/_0_ , \g16740/_0_ , \g16741/_0_ , \g16742/_0_ , \g16743/_0_ , \g16747/_0_ , \g16748/_0_ , \g16749/_0_ , \g16750/_0_ , \g16753/_0_ , \g16754/_0_ , \g16755/_0_ , \g16756/_0_ , \g16757/_0_ , \g16758/_0_ , \g16761/_0_ , \g16765/_0_ , \g16766/_0_ , \g16767/_0_ , \g16768/_0_ , \g16769/_0_ , \g16772/_0_ , \g16785/_0_ , \g16786/_0_ , \g16787/_0_ , \g16788/_0_ , \g16789/_0_ , \g16790/_0_ , \g16791/_0_ , \g16804/_0_ , \g16805/_0_ , \g16806/_0_ , \g16807/_0_ , \g16808/_0_ , \g16809/_0_ , \g16810/_0_ , \g16811/_0_ , \g16812/_0_ , \g16813/_0_ , \g16814/_0_ , \g16815/_0_ , \g16816/_0_ , \g16817/_0_ , \g16819/_0_ , \g16822/_0_ , \g16823/_0_ , \g16824/_0_ , \g16825/_0_ , \g16828/_0_ , \g16829/_0_ , \g16830/_0_ , \g16831/_0_ , \g16832/_0_ , \g16833/_0_ , \g16834/_0_ , \g16835/_0_ , \g16836/_0_ , \g16837/_0_ , \g16840/_0_ , \g16841/_0_ , \g16842/_0_ , \g16843/_0_ , \g16846/_0_ , \g16847/_0_ , \g16848/_0_ , \g16849/_0_ , \g16850/_0_ , \g16851/_0_ , \g16852/_0_ , \g16853/_0_ , \g16854/_0_ , \g16855/_0_ , \g16856/_0_ , \g16857/_0_ , \g16859/_0_ , \g16862/_0_ , \g16865/_0_ , \g16866/_0_ , \g16867/_0_ , \g16868/_0_ , \g16869/_0_ , \g16870/_0_ , \g16871/_0_ , \g16872/_0_ , \g16873/_0_ , \g16874/_0_ , \g16875/_0_ , \g16876/_0_ , \g16877/_0_ , \g16878/_0_ , \g16879/_0_ , \g16880/_0_ , \g16881/_0_ , \g16882/_0_ , \g16884/_0_ , \g16887/_0_ , \g16891/_0_ , \g16892/_0_ , \g16893/_0_ , \g16894/_0_ , \g16895/_0_ , \g16897/_0_ , \g16898/_0_ , \g16899/_0_ , \g16900/_0_ , \g16901/_0_ , \g16902/_0_ , \g16903/_0_ , \g16904/_0_ , \g16905/_0_ , \g16906/_0_ , \g16907/_0_ , \g16908/_0_ , \g16909/_0_ , \g16910/_0_ , \g16912/_0_ , \g16914/_0_ , \g16915/_0_ , \g16950/_0_ , \g16951/_0_ , \g16952/_0_ , \g16953/_0_ , \g16954/_0_ , \g16955/_0_ , \g16956/_0_ , \g16957/_0_ , \g16958/_0_ , \g16959/_0_ , \g16960/_0_ , \g16961/_0_ , \g16962/_0_ , \g16963/_0_ , \g16964/_0_ , \g16965/_0_ , \g16966/_0_ , \g16967/_0_ , \g16968/_0_ , \g16970/_0_ , \g17102/_3_ , \g17106/_0_ , \g17107/_0_ , \g17109/_0_ , \g17110/_0_ , \g17111/_0_ , \g17112/_0_ , \g17115/_0_ , \g17116/_0_ , \g17119/_0_ , \g17120/_0_ , \g17122/_0_ , \g17123/_0_ , \g17124/_0_ , \g17125/_0_ , \g17126/_0_ , \g17127/_0_ , \g17128/_0_ , \g17130/_0_ , \g17131/_0_ , \g17132/_0_ , \g17133/_0_ , \g17134/_0_ , \g17135/_0_ , \g17136/_0_ , \g17137/_0_ , \g17138/_0_ , \g17140/_0_ , \g17141/_0_ , \g17142/_0_ , \g17143/_0_ , \g17144/_0_ , \g17145/_0_ , \g17146/_0_ , \g17147/_0_ , \g17148/_0_ , \g17149/_0_ , \g17150/_0_ , \g17151/_0_ , \g17152/_0_ , \g17153/_0_ , \g17154/_0_ , \g17155/_0_ , \g17157/_0_ , \g17159/_0_ , \g17160/_0_ , \g17161/_0_ , \g17162/_0_ , \g17163/_0_ , \g17164/_0_ , \g17165/_0_ , \g17166/_0_ , \g17168/_0_ , \g17171/_0_ , \g17173/_0_ , \g17177/_0_ , \g17178/_0_ , \g17179/_0_ , \g17180/_0_ , \g17182/_0_ , \g17183/_0_ , \g17184/_0_ , \g17185/_0_ , \g17186/_0_ , \g17188/_0_ , \g17189/_0_ , \g17190/_0_ , \g17191/_0_ , \g17193/_0_ , \g17194/_0_ , \g17195/_0_ , \g17196/_0_ , \g17197/_0_ , \g17198/_0_ , \g17199/_0_ , \g17200/_0_ , \g17201/_0_ , \g17202/_0_ , \g17203/_0_ , \g17204/_0_ , \g17205/_0_ , \g17206/_0_ , \g17207/_0_ , \g17208/_0_ , \g17209/_0_ , \g17210/_0_ , \g17211/_0_ , \g17212/_0_ , \g17213/_0_ , \g17214/_0_ , \g17215/_0_ , \g17216/_0_ , \g17217/_0_ , \g17218/_0_ , \g17219/_0_ , \g17223/_0_ , \g17224/_0_ , \g17225/_0_ , \g17226/_0_ , \g17227/_0_ , \g17228/_0_ , \g17229/_0_ , \g17231/_0_ , \g17232/_0_ , \g17233/_0_ , \g17234/_0_ , \g17237/_0_ , \g17239/_0_ , \g17240/_0_ , \g17243/_0_ , \g17246/_0_ , \g17247/_0_ , \g17248/_0_ , \g17249/_0_ , \g17250/_0_ , \g17251/_0_ , \g17252/_0_ , \g17253/_0_ , \g17254/_0_ , \g17258/_0_ , \g17261/_0_ , \g17262/_0_ , \g17269/_0_ , \g17271/_0_ , \g17274/_0_ , \g17275/_0_ , \g17276/_0_ , \g17277/_0_ , \g17278/_0_ , \g17279/_0_ , \g17280/_0_ , \g17281/_0_ , \g17282/_0_ , \g17283/_0_ , \g17285/_0_ , \g17290/_0_ , \g17292/_0_ , \g17293/_0_ , \g17296/_0_ , \g17297/_0_ , \g17298/_0_ , \g173/_0_ , \g17303/_0_ , \g17304/_0_ , \g17305/_0_ , \g17306/_0_ , \g17307/_0_ , \g17308/_0_ , \g17309/_0_ , \g17310/_0_ , \g17311/_0_ , \g17312/_0_ , \g17314/_0_ , \g17315/_0_ , \g17316/_0_ , \g17317/_0_ , \g17318/_0_ , \g17319/_0_ , \g17320/_0_ , \g17321/_0_ , \g17322/_0_ , \g17323/_0_ , \g17324/_0_ , \g17325/_0_ , \g17326/_0_ , \g17327/_0_ , \g17328/_0_ , \g17329/_0_ , \g17330/_0_ , \g17331/_0_ , \g17332/_0_ , \g17333/_0_ , \g17335/_0_ , \g17336/_0_ , \g17337/_0_ , \g17338/_0_ , \g17339/_0_ , \g17340/_0_ , \g17342/_0_ , \g17343/_0_ , \g17347/_0_ , \g17350/_0_ , \g17354/_0_ , \g17356/_0_ , \g17357/_0_ , \g17358/_0_ , \g17359/_0_ , \g17360/_0_ , \g17415/_0_ , \g17441/_0_ , \g17442/_0_ , \g17451/_0_ , \g17457/_0_ , \g17458/_0_ , \g17459/_0_ , \g17460/_0_ , \g17461/_0_ , \g17462/_0_ , \g17463/_0_ , \g17464/_0_ , \g17465/_0_ , \g17466/_0_ , \g17467/_0_ , \g17468/_0_ , \g17469/_0_ , \g17470/_0_ , \g17471/_0_ , \g17472/_0_ , \g175/_3_ , \g1750/_0_ , \g176/_3_ , \g17619/_0_ , \g17620/_0_ , \g1763/_3_ , \g1764/_3_ , \g1768/_0_ , \g1769/_0_ , \g177/_3_ , \g17737/_0_ , \g17747/_0_ , \g178/_3_ , \g17814/_1_ , \g17815/_0_ , \g17821/_1_ , \g17821/_1__syn_2 , \g17872/_0_ , \g179/_3_ , \g17902/_0_ , \g180/_3_ , \g18020/_1_ , \g18057/_0_ , \g18096/_0_ , \g18099/_0_ , \g18107/_0_ , \g18133/_0_ , \g18140/_1_ , \g18153/_0_ , \g182/_0_ , \g18218/_0_ , \g18244/_0_ , \g18262/_0_ , \g18267/_0_ , \g18387/_1__syn_2 , \g184/_0_ , \g18478/_1_ , \g18585/_3_ , \g18608/_0_ , \g18609/_0_ , \g18613/_0_ , \g18618/_0_ , \g18647/_0_ , \g18687/_2_ , \g18707/_0_ , \g18748/_0_ , \g18753/_0_ , \g18758/_0_ , \g18759/_0_ , \g18760/_0_ , \g18761/_0_ , \g18762/_0_ , \g18763/_0_ , \g18764/_0_ , \g18765/_0_ , \g18766/_0_ , \g18767/_0_ , \g18768/_0_ , \g18770/_0_ , \g18771/_0_ , \g18788/_0_ , \g18796/_0_ , \g18800/_0_ , \g18801/_0_ , \g18802/_0_ , \g18803/_0_ , \g18804/_0_ , \g18805/_0_ , \g18807/_0_ , \g18840/_0_ , \g18843/_0_ , \g18844/_0_ , \g18846/_0_ , \g18847/_0_ , \g18848/_0_ , \g18849/_0_ , \g18850/_0_ , \g18851/_0_ , \g18852/_0_ , \g18853/_0_ , \g18854/_0_ , \g18855/_0_ , \g18856/_0_ , \g18858/_0_ , \g18860/_0_ , \g18861/_0_ , \g18863/_0_ , \g18864/_0_ , \g18866/_0_ , \g18867/_0_ , \g18868/_0_ , \g18869/_0_ , \g18870/_0_ , \g18871/_0_ , \g18872/_0_ , \g18873/_0_ , \g18874/_0_ , \g18875/_0_ , \g18876/_0_ , \g18877/_0_ , \g18878/_0_ , \g18879/_0_ , \g18880/_0_ , \g18881/_0_ , \g18882/_0_ , \g18883/_0_ , \g18888/_0_ , \g18892/_0_ , \g18895/_0_ , \g18896/_0_ , \g18897/_0_ , \g18905/_0_ , \g18908/_0_ , \g18909/_0_ , \g18912/_0_ , \g18918/_0_ , \g18919/_0_ , \g18920/_0_ , \g18921/_0_ , \g18922/_0_ , \g18924/_0_ , \g18925/_0_ , \g18927/_0_ , \g18930/_0_ , \g18966/_0_ , \g18968/_0_ , \g18970/_0_ , \g18974/_0_ , \g18975/_0_ , \g18977/_0_ , \g18981/_0_ , \g18983/_0_ , \g18985/_0_ , \g18987/_0_ , \g18989/_0_ , \g18991/_0_ , \g18992/_0_ , \g18993/_0_ , \g18994/_0_ , \g18995/_0_ , \g18996/_0_ , \g18997/_0_ , \g18998/_0_ , \g18999/_0_ , \g19001/_0_ , \g19003/_0_ , \g19005/_0_ , \g19006/_0_ , \g19014/_0_ , \g19016/_0_ , \g19018/_0_ , \g19020/_0_ , \g19022/_0_ , \g19056/_3_ , \g19058/_3_ , \g19060/_3_ , \g19062/_3_ , \g1910/_0_ , \g19186/_0_ , \g19188/_0_ , \g19235/_0_ , \g19239/_0_ , \g19244/_0_ , \g19253/_0_ , \g19254/_0_ , \g19259/_0_ , \g19261/_0_ , \g19267/_0_ , \g19277/_0_ , \g19278/_0_ , \g19280/_0_ , \g19281/_0_ , \g19282/_0_ , \g19283/_0_ , \g19284/_0_ , \g19285/_0_ , \g19286/_0_ , \g19287/_0_ , \g19288/_0_ , \g19289/_0_ , \g19290/_0_ , \g19291/_0_ , \g19292/_0_ , \g19293/_0_ , \g19294/_0_ , \g19295/_0_ , \g19296/_0_ , \g19297/_0_ , \g19298/_0_ , \g19299/_0_ , \g19300/_0_ , \g19301/_0_ , \g19302/_0_ , \g19303/_0_ , \g19304/_0_ , \g19305/_0_ , \g19306/_0_ , \g19307/_0_ , \g19308/_0_ , \g19315/_0_ , \g19316/_0_ , \g19317/_0_ , \g19318/_0_ , \g19319/_0_ , \g19320/_0_ , \g19321/_0_ , \g19322/_0_ , \g19323/_0_ , \g19325/_3_ , \g19326/_3_ , \g19333/_3_ , \g19341/_3_ , \g19347/_3_ , \g19377/_3_ , \g19381/_3_ , \g19393/_0_ , \g19401/_0_ , \g19402/_0_ , \g195/_2_ , \g19513/_0_ , \g19514/_0_ , \g19515/_0_ , \g19516/_0_ , \g1952/_3_ , \g19529/_0_ , \g19530/_0_ , \g19531/_0_ , \g19532/_0_ , \g19533/_0_ , \g19534/_0_ , \g19535/_0_ , \g19536/_0_ , \g19537/_0_ , \g19539/_0_ , \g19546/_0_ , \g19552/_0_ , \g19553/_0_ , \g19562/_0_ , \g19563/_0_ , \g19564/_0_ , \g19572/_0_ , \g19575/_0_ , \g19615/_0_ , \g19686/_0_ , \g19688/_0_ , \g197/_0_ , \g19729/_0_ , \g19774/_0_ , \g19777/_0_ , \g19791/_0_ , \g19818/_0_ , \g19819/_0_ , \g19828/_0_ , \g19852/_1_ , \g19860/_0_ , \g19861/_0_ , \g19864/_0_ , \g19886/_0_ , \g19887/_0_ , \g199/_0_ , \g19908/_0_ , \g19918/_0_ , \g19927/_0_ , \g19933/_0_ , \g200/_0_ , \g20019/_0_ , \g20046/_0_ , \g20068/_1_ , \g20080/_1_ , \g201/_0_ , \g20137/_0_ , \g20139/_0_ , \g20141/_0_ , \g20152/_1_ , \g20154/_00_ , \g202/_0_ , \g20206/_0_ , \g20211/_2_ , \g20217/_2_ , \g20239/_0_ , \g20265/_2_ , \g20266/_0_ , \g20272/_2_ , \g20278/_2_ , \g20283/_0_ , \g20285/_2_ , \g20288/_2__syn_2 , \g20293/_0_ , \g20295/_2_ , \g203/_0_ , \g20302/_2_ , \g20303/_2_ , \g20304/_2_ , \g20311/_2_ , \g20326/_0_ , \g20330/_0_ , \g2034/_0_ , \g20345/_0_ , \g20346/_0_ , \g2035/_0_ , \g20363/_0_ , \g20364/_0_ , \g204/_0_ , \g2047/_0_ , \g20483/_0_ , \g20493/_00_ , \g205/_0_ , \g20569/_0_ , \g20570/_0_ , \g20571/_0_ , \g206/_0_ , \g20613/_0_ , \g20615/_0_ , \g20657/_1__syn_2 , \g20660/_0_ , \g20685/_0_ , \g207/_0_ , \g20713/_1_ , \g20747/_1_ , \g20784/_0_ , \g20820/_1_ , \g20859/_0_ , \g20873/_2_ , \g20886/_0_ , \g20887/_0_ , \g20891/_2__syn_2 , \g20907/_2_ , \g20936/_2__syn_2 , \g20937/_1_ , \g20955/_0_ , \g20959/_2__syn_2 , \g20967/_0_ , \g20971/_2__syn_2 , \g20974/_1__syn_2 , \g21015/_1_ , \g21051/_2_ , \g21079/_1_ , \g21081/_1_ , \g21087/_2__syn_2 , \g21114/_1_ , \g21116/_1_ , \g21120/_2__syn_2 , \g21147/_0_ , \g21179/_1_ , \g21185/_1_ , \g21223/_0_ , \g21242/_0_ , \g21253/_0_ , \g21257/_0_ , \g21323/_1_ , \g21324/_1_ , \g21366/_0_ , \g21385/_2_ , \g21464/_0_ , \g21475/_3_ , \g21481/_0_ , \g21482/_0_ , \g21494/_3_ , \g21500/_3_ , \g21507/_3_ , \g21511/_3_ , \g21537/_1_ , \g21568/_0_ , \g21591/_0_ , \g21604/_0_ , \g21605/_3_ , \g21606/_0_ , \g21607/_0_ , \g21608/_0_ , \g21609/_0_ , \g21610/_0_ , \g21611/_0_ , \g21612/_0_ , \g21613/_0_ , \g21614/_0_ , \g21615/_0_ , \g21616/_0_ , \g21617/_0_ , \g21618/_0_ , \g21621/_0_ , \g21640/_0_ , \g21678/_0_ , \g21679/_0_ , \g21686/_0_ , \g21692/_3_ , \g21696/_0_ , \g21698/_0_ , \g21702/_3_ , \g21707/_0_ , \g21709/_0_ , \g21728/_0_ , \g21729/_0_ , \g21731/_0_ , \g21732/_0_ , \g21733/_0_ , \g21736/_0_ , \g21744/_3_ , \g21753/_0_ , \g21754/_0_ , \g21755/_0_ , \g21756/_0_ , \g21757/_0_ , \g21759/_0_ , \g21761/_0_ , \g21763/_0_ , \g21764/_0_ , \g21766/_0_ , \g2180/_0_ , \g21853/_3_ , \g21861/_3_ , \g21863/_3_ , \g21869/_3_ , \g2187/_0_ , \g21875/_3_ , \g21877/_3_ , \g21879/_3_ , \g2188/_0_ , \g21900/_0_ , \g22080/_0_ , \g22082/_0_ , \g22135/_0_ , \g22145/_1_ , \g22225/_0_ , \g223/_0_ , \g22354/_0_ , \g224/_0_ , \g22412/_0_ , \g22415/_1__syn_2 , \g225/_0_ , \g2257/_0_ , \g226/_3_ , \g22624/_0_ , \g227/_3_ , \g22702/_0_ , \g22919/_1__syn_2 , \g22933/_0_ , \g22954/_0_ , \g22989/_1_ , \g23529/_0_ , \g23539/_0_ , \g2362/_2_ , \g23766/_0_ , \g24/_3_ , \g24018/_0_ , \g2416/_0_ , \g2420/_0_ , \g24213/_0_ , \g24301/_0_ , \g2479/_0_ , \g248/_3_ , \g2480/_0_ , \g2481/_0_ , \g2482/_0_ , \g2483/_0_ , \g2484/_0_ , \g2485/_0_ , \g2486/_0_ , \g2487/_0_ , \g2488/_0_ , \g249/_3_ , \g2490/_0_ , \g2491/_0_ , \g2492/_0_ , \g2493/_0_ , \g2494/_0_ , \g2495/_0_ , \g2496/_0_ , \g2497/_0_ , \g2507/_0_ , \g2508/_0_ , \g2509/_0_ , \g2510/_0_ , \g2511/_0_ , \g2512/_0_ , \g2513/_0_ , \g2514/_0_ , \g2515/_0_ , \g2516/_0_ , \g25237/_0_ , \g2558/_0_ , \g2562/_0_ , \g2563/_0_ , \g2564/_0_ , \g2565/_0_ , \g2566/_0_ , \g2567/_0_ , \g2699/_0_ , \g27/_2_ , \g271/_0_ , \g272/_3_ , \g273/_3_ , \g274/_3_ , \g275/_3_ , \g276/_3_ , \g277/_3_ , \g2787/_3_ , \g2788/_3_ , \g279/_0_ , \g2795/_0_ , \g2796/_0_ , \g280/_0_ , \g2842/_3_ , \g29/_1_ , \g2927/_0_ , \g2978/_0_ , \g2979/_0_ , \g2980/_0_ , \g2981/_0_ , \g2982/_0_ , \g2983/_0_ , \g2984/_0_ , \g2985/_0_ , \g3021/_3_ , \g3022/_3_ , \g3023/_3_ , \g3024/_3_ , \g3025/_3_ , \g3026/_3_ , \g3027/_3_ , \g3028/_3_ , \g3029/_3_ , \g3030/_3_ , \g3031/_3_ , \g3032/_3_ , \g3033/_3_ , \g3034/_3_ , \g3035/_3_ , \g3036/_3_ , \g3037/_3_ , \g3038/_3_ , \g3039/_3_ , \g3040/_3_ , \g3041/_3_ , \g3042/_3_ , \g3049/_0_ , \g3050/_0_ , \g3051/_0_ , \g3052/_0_ , \g3053/_0_ , \g3054/_0_ , \g3058/_0_ , \g3059/_0_ , \g3088/_0_ , \g3089/_0_ , \g3090/_0_ , \g3091/_0_ , \g3092/_0_ , \g3093/_0_ , \g3094/_0_ , \g3095/_0_ , \g314/_0_ , \g3147/_3_ , \g3148/_3_ , \g3189/_0_ , \g3190/_0_ , \g3191/_0_ , \g3192/_0_ , \g3193/_0_ , \g3194/_0_ , \g3195/_0_ , \g3196/_0_ , \g3197/_0_ , \g3198/_0_ , \g3199/_0_ , \g32/_0_ , \g320/_3_ , \g3200/_0_ , \g3201/_0_ , \g3202/_0_ , \g3203/_0_ , \g3204/_0_ , \g321/_3_ , \g325/_3_ , \g3271/_2_ , \g33/_0_ , \g3363/_0_ , \g3413/_0_ , \g3414/_0_ , \g352/_0_ , \g355/_0_ , \g356/_3_ , \g357/_3_ , \g35_dup/_1_ , \g36/_3_ , \g365/_3_ , \g366/_3_ , \g367/_3_ , \g368/_3_ , \g3687/_0_ , \g369/_3_ , \g37/_3_ , \g370/_3_ , \g372/_3_ , \g374/_3_ , \g3740/_0_ , \g375/_3_ , \g376/_3_ , \g3878/_0_ , \g3879/_0_ , \g388/_3_ , \g3880/_0_ , \g3881/_0_ , \g3882/_0_ , \g389/_3_ , \g3894/_0_ , \g3895/_0_ , \g3896/_0_ , \g3897/_0_ , \g3898/_0_ , \g392/_3_ , \g393/_3_ , \g394/_3_ , \g395/_3_ , \g396/_3_ , \g397/_3_ , \g398/_3_ , \g399/_3_ , \g401/_3_ , \g402/_3_ , \g404/_3_ , \g4048/_0_ , \g405/_3_ , \g4050/_0_ , \g406/_3_ , \g407/_3_ , \g410/_3_ , \g411/_3_ , \g412/_3_ , \g413/_3_ , \g415/_3_ , \g416/_3_ , \g42/_0_ , \g4216/_3_ , \g4217/_3_ , \g4218/_3_ , \g4219/_3_ , \g4296/_0_ , \g4297/_0_ , \g4298/_0_ , \g4299/_0_ , \g43/_0_ , \g4300/_0_ , \g4301/_0_ , \g4302/_0_ , \g4303/_0_ , \g4304/_0_ , \g4305/_0_ , \g4306/_0_ , \g4307/_0_ , \g4308/_0_ , \g4309/_0_ , \g4310/_0_ , \g4311/_0_ , \g4312/_0_ , \g4313/_0_ , \g4314/_0_ , \g4315/_0_ , \g4316/_0_ , \g4317/_0_ , \g4318/_0_ , \g4319/_0_ , \g4320/_0_ , \g4321/_0_ , \g4322/_0_ , \g4323/_0_ , \g436/_0_ , \g44/_0_ , \g448/_3_ , \g45/_0_ , \g4587/_0_ , \g4588/_0_ , \g46/_0_ , \g4601/_0_ , \g4602/_0_ , \g4613/_3_ , \g4614/_3_ , \g4615/_3_ , \g463/_0_ , \g465/_0_ , \g4653/_0_ , \g4654/_0_ , \g4655/_0_ , \g4656/_0_ , \g4659/_0_ , \g466/_0_ , \g468/_3_ , \g469/_3_ , \g4697/_0_ , \g47/_3_ , \g470/_0_ , \g471/_0_ , \g4755/_0_ , \g476/_0_ , \g48/_3_ , \g480/_00_ , \g4839/_0_ , \g4840/_0_ , \g485/_3_ , \g4854/_0_ , \g4855/_0_ , \g4859/_0_ , \g486/_3_ , \g4860/_0_ , \g4880/_0_ , \g4881/_0_ , \g4882/_0_ , \g4883/_0_ , \g4884/_0_ , \g4885/_0_ , \g4886/_0_ , \g4887/_0_ , \g4888/_0_ , \g49/_0_ , \g494/_0_ , \g499/_1_ , \g50/_0_ , \g5002/_0_ , \g5003/_0_ , \g5009/_0_ , \g5010/_0_ , \g5011/_0_ , \g5014/_0_ , \g51/_0_ , \g5105/_0_ , \g5129/_2_ , \g5132/_0_ , \g5135/_0_ , \g5168/_0_ , \g5169/_0_ , \g5173/_0_ , \g5224/_0_ , \g5225/_0_ , \g5226/_0_ , \g5227/_0_ , \g5334/_0_ , \g5335/_0_ , \g5336/_0_ , \g5337/_0_ , \g5338/_0_ , \g5339/_0_ , \g5340/_0_ , \g5341/_0_ , \g5342/_0_ , \g5343/_0_ , \g5344/_0_ , \g5345/_0_ , \g5346/_0_ , \g5347/_0_ , \g5348/_0_ , \g5349/_0_ , \g5395/_0_ , \g54/_0_ , \g5434/_0_ , \g5447/_0_ , \g5450/_0_ , \g5451/_0_ , \g5452/_0_ , \g5453/_0_ , \g5454/_0_ , \g5461/_0_ , \g5483/_0_ , \g5484/_0_ , \g5492/_0_ , \g5493/_0_ , \g5496/_3_ , \g5497/_3_ , \g55/_0_ , \g5500/_0_ , \g5502/_0_ , \g5503/_0_ , \g5506/_0_ , \g5511/_0_ , \g5518/_0_ , \g5519/_0_ , \g5520/_0_ , \g5522/_0_ , \g5523/_0_ , \g5524/_0_ , \g5525/_0_ , \g5532/_0_ , \g5533/_0_ , \g5534/_0_ , \g5535/_0_ , \g5536/_0_ , \g5537/_0_ , \g5538/_0_ , \g5546/_0_ , \g5555/_00_ , \g5593/_0_ , \g5614/_2_ , \g567/_0_ , \g5677/_0_ , \g5678/_0_ , \g5682/_0_ , \g5683/_0_ , \g5684/_0_ , \g5686/_0_ , \g5687/_0_ , \g5689/_0_ , \g5690/_0_ , \g5691/_0_ , \g5692/_0_ , \g5698/_0_ , \g5699/_0_ , \g5700/_0_ , \g5701/_0_ , \g5702/_0_ , \g5703/_0_ , \g5704/_0_ , \g5709/_0_ , \g5711/_0_ , \g5714/_0_ , \g572/_0_ , \g5723/_0_ , \g5724/_0_ , \g5725/_0_ , \g573/_0_ , \g5739/_0_ , \g5740/_0_ , \g575/_0_ , \g5756/_0_ , \g5757/_0_ , \g5758/_0_ , \g5759/_0_ , \g576/_0_ , \g5760/_0_ , \g5761/_0_ , \g5762/_0_ , \g5763/_0_ , \g577/_0_ , \g5772/_0_ , \g5773/_0_ , \g5774/_0_ , \g5775/_0_ , \g5776/_0_ , \g5777/_0_ , \g578/_0_ , \g5781/_0_ , \g5783/_0_ , \g5784/_0_ , \g5785/_0_ , \g5786/_0_ , \g5787/_0_ , \g5788/_0_ , \g5789/_0_ , \g579/_0_ , \g5790/_0_ , \g5791/_0_ , \g5792/_0_ , \g5794/_0_ , \g5795/_0_ , \g5796/_0_ , \g580/_0_ , \g5801/_0_ , \g5802/_0_ , \g5803/_0_ , \g5804/_0_ , \g5805/_0_ , \g581/_0_ , \g5814/_0_ , \g582/_0_ , \g583/_0_ , \g5849/_3_ , \g585/_0_ , \g586/_0_ , \g587/_0_ , \g588/_0_ , \g589/_0_ , \g590/_0_ , \g591/_0_ , \g592/_0_ , \g593/_0_ , \g594/_0_ , \g595/_0_ , \g596/_0_ , \g597/_0_ , \g5971/_0_ , \g5972/_0_ , \g5976/_0_ , \g598/_0_ , \g5989/_0_ , \g599/_0_ , \g600/_0_ , \g601/_0_ , \g602/_0_ , \g603/_0_ , \g604/_0_ , \g605/_0_ , \g6092/_0_ , \g6093/_2_ , \g6094/_0_ , \g6114/_0_ , \g614/_3_ , \g6148/_0_ , \g6149/_0_ , \g6171/_0_ , \g6172/_0_ , \g6173/_0_ , \g6174/_0_ , \g6175/_0_ , \g6176/_0_ , \g6177/_0_ , \g6178/_0_ , \g6179/_0_ , \g6180/_0_ , \g6181/_0_ , \g6182/_0_ , \g6183/_0_ , \g6184/_0_ , \g6185/_0_ , \g6186/_0_ , \g6187/_0_ , \g6193/_0_ , \g6196/_0_ , \g6197/_0_ , \g6198/_3_ , \g6200/_2_ , \g6202/_2_ , \g6203/_3_ , \g6204/_3_ , \g6209/_0_ , \g6211/_0_ , \g6215/_0_ , \g6217/_0_ , \g6219/_0_ , \g6220/_0_ , \g6222/_0_ , \g6224/_0_ , \g6228/_0_ , \g6238/_0_ , \g6239/_0_ , \g6240/_0_ , \g6242/_0_ , \g6243/_0_ , \g6244/_0_ , \g6245/_0_ , \g6246/_0_ , \g6248/_0_ , \g6249/_0_ , \g6259/_0_ , \g6260/_0_ , \g6261/_0_ , \g6262/_0_ , \g6263/_0_ , \g6264/_0_ , \g6265/_0_ , \g6266/_0_ , \g6267/_0_ , \g6268/_0_ , \g6269/_0_ , \g6270/_0_ , \g6271/_0_ , \g6272/_0_ , \g6277/_0_ , \g6318/_0_ , \g6326/_0_ , \g6329/_0_ , \g6330/_0_ , \g6331/_0_ , \g6332/_0_ , \g6333/_0_ , \g6334/_0_ , \g6335/_0_ , \g6336/_0_ , \g6337/_0_ , \g6338/_0_ , \g6339/_0_ , \g6340/_0_ , \g6341/_0_ , \g6342/_0_ , \g6343/_0_ , \g6344/_0_ , \g6345/_0_ , \g6346/_0_ , \g6347/_0_ , \g6348/_0_ , \g6349/_0_ , \g6350/_0_ , \g6351/_0_ , \g6352/_0_ , \g6353/_0_ , \g6354/_0_ , \g6355/_0_ , \g6361/_0_ , \g637/_0_ , \g638/_0_ , \g639/_3_ , \g64/_3_ , \g640/_3_ , \g6419/_0_ , \g6442/_0_ , \g6442/_1_ , \g6489/_0_ , \g6490/_0_ , \g65/_3_ , \g6513/_0_ , \g6515/_0_ , \g6571/_0_ , \g6588/_0_ , \g6589/_0_ , \g6638/_0_ , \g6639/_0_ , \g6653/_0_ , \g6654/_3_ , \g6655/_0_ , \g6656/_0_ , \g6657/_0_ , \g6687/_0_ , \g6688/_0_ , \g6689/_0_ , \g6690/_0_ , \g6691/_0_ , \g6692/_0_ , \g6693/_0_ , \g6694/_0_ , \g6701/_0_ , \g6706/_0_ , \g6711/_0_ , \g6727/_0_ , \g6728/_0_ , \g6736/_0_ , \g6739/_0_ , \g6742/_0_ , \g6746/_0_ , \g6752/_0_ , \g6771/_0_ , \g684/_0_ , \g685/_0_ , \g686/_0_ , \g687/_0_ , \g688/_0_ , \g689/_0_ , \g690/_0_ , \g691/_0_ , \g692/_0_ , \g693/_0_ , \g696/_3_ , \g697/_3_ , \g699/_0_ , \g7/_0_ , \g700/_0_ , \g7005/_0_ , \g7056/_0_ , \g7057/_0_ , \g7058/_0_ , \g7060/_0_ , \g7075/_0_ , \g7086/_0_ , \g7087/_0_ , \g7089/_0_ , \g7108/_0_ , \g7109/_0_ , \g7112/_0_ , \g7172/_2_ , \g7210/_2_ , \g7211/_0_ , \g7212/_0_ , \g7213/_0_ , \g7214/_0_ , \g7215/_0_ , \g7216/_0_ , \g7217/_3_ , \g7218/_0_ , \g7219/_0_ , \g7220/_0_ , \g7222/_0_ , \g7227/_2_ , \g723/_3_ , \g7234/_0_ , \g7237/_3_ , \g7238/_3_ , \g7239/_3_ , \g724/_3_ , \g7240/_3_ , \g7241/_3_ , \g7242/_3_ , \g7243/_3_ , \g7244/_0_ , \g7245/_0_ , \g7246/_0_ , \g7247/_0_ , \g7248/_0_ , \g7249/_0_ , \g7250/_0_ , \g7251/_0_ , \g7253/_0_ , \g7254/_0_ , \g7255/_0_ , \g7256/_0_ , \g7257/_0_ , \g7258/_0_ , \g7261/_0_ , \g7264/_0_ , \g7265/_0_ , \g7266/_0_ , \g7267/_0_ , \g7268/_0_ , \g7269/_0_ , \g7278/_0_ , \g7279/_0_ , \g7280/_0_ , \g7281/_0_ , \g7282/_0_ , \g7283/_0_ , \g7284/_0_ , \g7285/_0_ , \g7286/_3_ , \g7288/_3_ , \g7291/_0_ , \g7296/_3_ , \g73/_0_ , \g7302/_3_ , \g7306/_3_ , \g7310/_3_ , \g7311/_3_ , \g7312/_3_ , \g7313/_3_ , \g7314/_3_ , \g7315/_3_ , \g7316/_3_ , \g7317/_3_ , \g7323/_3_ , \g7324/_3_ , \g7325/_3_ , \g7327/_0_ , \g7362/_0_ , \g74/_0_ , \g75/_0_ , \g7512/_0_ , \g7513/_0_ , \g7514/_0_ , \g7515/_0_ , \g7516/_0_ , \g7518/_0_ , \g7528/_0_ , \g7529/_0_ , \g7548/_0_ , \g7549/_0_ , \g7550/_0_ , \g7575/_0_ , \g7576/_0_ , \g7577/_0_ , \g7578/_0_ , \g7579/_0_ , \g7580/_0_ , \g7581/_0_ , \g7582/_0_ , \g7583/_0_ , \g7584/_0_ , \g7585/_0_ , \g7586/_0_ , \g7587/_0_ , \g7588/_0_ , \g7589/_0_ , \g7590/_0_ , \g7591/_0_ , \g7592/_0_ , \g7593/_0_ , \g7594/_0_ , \g7595/_0_ , \g7596/_0_ , \g7597/_0_ , \g7598/_0_ , \g7599/_0_ , \g76/_0_ , \g7600/_0_ , \g7601/_0_ , \g7602/_0_ , \g7603/_0_ , \g7604/_0_ , \g7614/_0_ , \g7618/_0_ , \g762/_0_ , \g7634/_0_ , \g766/_0_ , \g767/_0_ , \g768/_0_ , \g769/_0_ , \g77/_0_ , \g770/_3_ , \g771/_3_ , \g7715/_0_ , \g774/_0_ , \g7746/_0_ , \g7753/_0_ , \g7754/_0_ , \g7755/_0_ , \g7756/_0_ , \g7757/_0_ , \g7758/_0_ , \g7759/_0_ , \g7760/_0_ , \g7761/_0_ , \g7762/_0_ , \g7763/_0_ , \g7764/_0_ , \g7765/_0_ , \g7766/_0_ , \g7778/_0_ , \g7779/_0_ , \g7780/_0_ , \g7781/_0_ , \g7782/_0_ , \g7784/_0_ , \g78/_0_ , \g7800/_0_ , \g7823/_3_ , \g7837/_0_ , \g7841/_0_ , \g7842/_0_ , \g7843/_0_ , \g7844/_0_ , \g7845/_0_ , \g7846/_0_ , \g7847/_0_ , \g7849/_0_ , \g7850/_0_ , \g7852/_0_ , \g7854/_0_ , \g7855/_0_ , \g7857/_0_ , \g7858/_0_ , \g7859/_0_ , \g7860/_0_ , \g7861/_0_ , \g7862/_0_ , \g7863/_0_ , \g7864/_0_ , \g7865/_0_ , \g7866/_0_ , \g7867/_0_ , \g7868/_0_ , \g7869/_0_ , \g7870/_0_ , \g7871/_0_ , \g79211/_3_ , \g79258/_3_ , \g79299/_3_ , \g79316/_2_ , \g79342/_3_ , \g79401/_3_ , \g79452/_3_ , \g79457/_3_ , \g7951/_0_ , \g79541/_3_ , \g7958/_0_ , \g79598/_3_ , \g79654/_3_ , \g79675/_3_ , \g7971/_0_ , \g7972/_0_ , \g7973/_3_ , \g79753/_3_ , \g7976/_3_ , \g79855/_3_ , \g79858/_3_ , \g79997/_3_ , \g8/_0_ , \g80008/_3_ , \g80011/_0_ , \g80104/_0_ , \g80172/_1_ , \g80195/_3_ , \g80238/_3_ , \g80290/_2_ , \g80294/_0_ , \g80302/_0_ , \g80327/_0_ , \g80360/_3_ , \g80373/_0_ , \g80401/_0_ , \g80410/_0_ , \g80475/_0_ , \g80476/_0_ , \g80516/_3_ , \g80536/_0_ , \g80537/_0_ , \g80572/_0_ , \g80573/_0_ , \g80609/_2_ , \g80610/_2_ , \g80676/_0_ , \g80798/_0_ , \g80807/_0_ , \g80890/_2_ , \g80904/_0_ , \g81719/_2_ , \g81746/_0_ , \g81775/_0_ , \g81872/_0_ , \g81961/_0_ , \g81968/_0_ , \g82096/_0_ , \g82123/_0_ , \g82147/_0_ , \g82147/_1_ , \g82335/_0_ , \g82338/_2_ , \g82368/_0_ , \g82460/_2_ , \g82469/_0_ , \g82481/_0_ , \g82625/_1_ , \g82711/_0_ , \g82772/_0_ , \g82946/_0_ , \g82947/_0_ , \g82956/_0_ , \g83003/_0_ , \g83006/_1_ , \g83415/_0_ , \g83498/_0_ , \g837/_0_ , \g838/_0_ , \g83863/_0_ , \g839/_0_ , \g84049/_3_ , \g84050/_3_ , \g84077/_2_ , \g842/_0_ , \g84245/_0_ , \g843/_0_ , \g844/_0_ , \g84448/_0_ , \g84478/_3_ , \g845/_0_ , \g846/_0_ , \g847/_0_ , \g848/_0_ , \g8487/_0_ , \g8488/_0_ , \g8489/_0_ , \g849/_0_ , \g8490/_0_ , \g84904/_0_ , \g8491/_0_ , \g8492/_0_ , \g8493/_0_ , \g8494/_0_ , \g8496/_0_ , \g8517/_0_ , \g8534/_0_ , \g8538/_0_ , \g8540/_0_ , \g8576/_2_ , \g8597/_0_ , \g8598/_0_ , \g8599/_0_ , \g8600/_0_ , \g8601/_0_ , \g8602/_0_ , \g8603/_0_ , \g8605/_0_ , \g8606/_0_ , \g8607/_0_ , \g8608/_0_ , \g8609/_0_ , \g8610/_0_ , \g8611/_0_ , \g8612/_0_ , \g8613/_0_ , \g8614/_0_ , \g8615/_0_ , \g8617/_0_ , \g8643/_0_ , \g8644/_0_ , \g8645/_0_ , \g8646/_0_ , \g8647/_0_ , \g8648/_0_ , \g8650/_0_ , \g8651/_0_ , \g8652/_0_ , \g8653/_0_ , \g8654/_0_ , \g8655/_0_ , \g8656/_0_ , \g8657/_0_ , \g8658/_0_ , \g8659/_0_ , \g8660/_0_ , \g8665/_00_ , \g8666/_00_ , \g8667/_00_ , \g8668/_00_ , \g8669/_00_ , \g86715/_0_ , \g86745/_3_ , \g8691/_0_ , \g8700/_0_ , \g8701/_0_ , \g8702/_0_ , \g8703/_0_ , \g8704/_0_ , \g8705/_0_ , \g87063/_0_ , \g87114/_0_ , \g8712/_0_ , \g8713/_0_ , \g8714/_0_ , \g87171/_1_ , \g87252/_1_ , \g87298/_0_ , \g8730/_0_ , \g8741/_0_ , \g8747/_0_ , \g87480/_0_ , \g87484/_2_ , \g87488/_1__syn_2 , \g8761/_0_ , \g8762/_0_ , \g8763/_0_ , \g8764/_0_ , \g8765/_0_ , \g8775/_0_ , \g8776/_0_ , \g8777/_0_ , \g8778/_0_ , \g8784/_0_ , \g8804/_0_ , \g8807/_0_ , \g8808/_0_ , \g8809/_0_ , \g8810/_0_ , \g8811/_0_ , \g8812/_0_ , \g8813/_0_ , \g8814/_0_ , \g8815/_0_ , \g8816/_0_ , \g8817/_0_ , \g8818/_0_ , \g8819/_0_ , \g8820/_0_ , \g8821/_0_ , \g8822/_0_ , \g8823/_0_ , \g8824/_0_ , \g8825/_0_ , \g8826/_0_ , \g8827/_0_ , \g8828/_0_ , \g8829/_0_ , \g8830/_0_ , \g8831/_0_ , \g8832/_0_ , \g8833/_0_ , \g8834/_0_ , \g8835/_0_ , \g8836/_0_ , \g8837/_0_ , \g8838/_0_ , \g8839/_0_ , \g8840/_0_ , \g8842/_0_ , \g8843/_0_ , \g8846/_0_ , \g8848/_0_ , \g8857/_0_ , \g8895/_0_ , \g8902/_3_ , \g8903/_3_ , \g8904/_3_ , \g8905/_3_ , \g8906/_3_ , \g8909/_0_ , \g8910/_0_ , \g8911/_0_ , \g8924/_3_ , \g8926/_3_ , \g8927/_3_ , \g8943/_0_ , \g8944/_0_ , \g8958/_3_ , \g8960/_00_ , \g8961/_3_ , \g8965/_0_ , \g8966/_0_ , \g8967/_0_ , \g8968/_0_ , \g9/_0_ , \g9123/_0_ , \g9125/_0_ , \g9126/_0_ , \g913/_0_ , \g915/_0_ , \g916/_0_ , \g917/_0_ , \g918/_0_ , \g919/_0_ , \g920/_3_ , \g921/_3_ , \g925/_0_ , \g926/_0_ , \g927/_0_ , \g928/_0_ , \g929/_0_ , \g930/_0_ , \g9336/_0_ , \g9337/_0_ , \g939/_3_ , \g9396/_0_ , \g9397/_0_ , \g9399/_0_ , \g9400/_0_ , \g9401/_0_ , \g9402/_0_ , \g9403/_0_ , \g9404/_0_ , \g9415/_0_ , \g9418/_0_ , \g9419/_0_ , \g9420/_0_ , \g9446/_0_ , \g9465/_0_ , \g9493/_0_ , \g9536/_0_ , \g9537/_0_ , \g9538/_0_ , \g9539/_0_ , \g9540/_0_ , \g9541/_0_ , \g9542/_0_ , \g955/_2_ , \g9561/_0_ , \g9562/_0_ , \g9563/_0_ , \g9564/_0_ , \g9565/_0_ , \g9566/_0_ , \g9567/_0_ , \g9568/_0_ , \g9569/_0_ , \g9570/_0_ , \g9571/_0_ , \g9572/_0_ , \g9573/_0_ , \g9574/_0_ , \g9575/_0_ , \g9576/_0_ , \g9577/_0_ , \g9578/_0_ , \g9579/_0_ , \g9580/_0_ , \g9581/_0_ , \g9582/_0_ , \g9583/_0_ , \g9584/_0_ , \g9585/_0_ , \g9586/_0_ , \g9587/_0_ , \g9588/_0_ , \g9589/_0_ , \g9590/_0_ , \g9591/_0_ , \g9592/_0_ , \g9593/_0_ , \g9594/_0_ , \g9595/_0_ , \g9596/_0_ , \g9597/_0_ , \g9598/_0_ , \g9599/_0_ , \g9600/_0_ , \g9601/_0_ , \g9602/_0_ , \g9603/_0_ , \g9604/_0_ , \g9605/_0_ , \g9606/_0_ , \g9607/_0_ , \g9608/_0_ , \g9609/_0_ , \g9610/_0_ , \g9611/_0_ , \g9612/_0_ , \g9613/_0_ , \g9614/_0_ , \g9615/_0_ , \g9616/_0_ , \g9617/_0_ , \g9618/_0_ , \g9619/_0_ , \g9620/_0_ , \g9621/_0_ , \g9622/_0_ , \g9623/_0_ , \g9624/_0_ , \g9625/_0_ , \g9626/_0_ , \g9627/_0_ , \g9628/_0_ , \g9629/_0_ , \g9630/_0_ , \g9631/_0_ , \g9632/_0_ , \g9633/_0_ , \g9634/_0_ , \g9635/_0_ , \g9636/_0_ , \g9637/_0_ , \g9638/_0_ , \g9639/_0_ , \g9640/_0_ , \g9641/_0_ , \g9642/_0_ , \g9643/_0_ , \g9644/_0_ , \g9645/_0_ , \g9646/_0_ , \g9647/_0_ , \g9648/_0_ , \g9649/_0_ , \g9650/_0_ , \g9651/_0_ , \g9652/_0_ , \g9653/_0_ , \g9654/_0_ , \g9655/_0_ , \g9656/_0_ , \g9657/_0_ , \g9658/_0_ , \g9659/_0_ , \g9660/_0_ , \g9661/_0_ , \g9662/_0_ , \g9663/_0_ , \g9664/_0_ , \g9665/_0_ , \g9666/_0_ , \g9667/_0_ , \g9668/_0_ , \g9669/_0_ , \g9670/_0_ , \g9671/_0_ , \g9672/_0_ , \g9673/_0_ , \g9674/_0_ , \g9675/_0_ , \g9676/_0_ , \g9677/_0_ , \g9678/_0_ , \g9681/_0_ , \g9683/_0_ , \g9689/_0_ , \g9692/_0_ , \g9694/_0_ , \g9695/_0_ , \g9701/_0_ , \g9702/_0_ , \g9703/_0_ , \g9704/_0_ , \g9709/_0_ , \g9710/_0_ , \g9711/_0_ , \g9712/_0_ , \g9720/_0_ , \g9721/_0_ , \g9722/_0_ , \g9726/_0_ , \g9733/_0_ , \g9734/_0_ , \g9735/_0_ , \g9736/_0_ , \g9737/_0_ , \g9738/_0_ , \g9739/_0_ , \g9740/_0_ , \g9741/_0_ , \g9742/_0_ , \g9743/_0_ , \g9744/_0_ , \g9745/_0_ , \g9746/_0_ , \g9747/_0_ , \g9748/_0_ , \g9749/_0_ , \g9750/_0_ , \g9751/_0_ , \g9752/_0_ , \g9753/_0_ , \g9754/_0_ , \g9755/_0_ , \g9756/_0_ , \g9757/_0_ , \g9758/_0_ , \g9759/_0_ , \g9760/_0_ , \g9761/_0_ , \g9762/_0_ , \g9763/_0_ , \g9764/_0_ , \g9765/_0_ , \g9766/_0_ , \g9767/_0_ , \g9768/_0_ , \g9769/_0_ , \g9770/_0_ , \g9771/_0_ , \g9772/_0_ , \g9773/_0_ , \g9774/_0_ , \g9775/_0_ , \g9776/_0_ , \g9777/_0_ , \g9778/_0_ , \g9779/_0_ , \g9780/_0_ , \g9781/_0_ , \g9782/_0_ , \g9783/_0_ , \g9784/_0_ , \g9785/_0_ , \g9786/_0_ , \g9787/_0_ , \g9788/_0_ , \g9789/_0_ , \g9790/_0_ , \g9791/_0_ , \g9792/_0_ , \g9793/_0_ , \g9794/_0_ , \g9795/_0_ , \g9796/_0_ , \g9797/_0_ , \g9798/_0_ , \g9799/_0_ , \g9800/_0_ , \g9801/_0_ , \g9802/_0_ , \g9803/_0_ , \g9804/_0_ , \g9805/_0_ , \g9806/_0_ , \g9807/_0_ , \g9808/_0_ , \g9809/_0_ , \g9810/_0_ , \g9811/_0_ , \g9812/_0_ , \g9813/_0_ , \g9814/_0_ , \g9815/_0_ , \g9816/_0_ , \g9817/_0_ , \g9818/_0_ , \g9819/_0_ , \g9820/_0_ , \g9821/_0_ , \g9822/_0_ , \g9823/_0_ , \g9824/_0_ , \g9825/_0_ , \g9826/_0_ , \g9827/_0_ , \g9828/_0_ , \g9829/_0_ , \g9830/_0_ , \g9831/_0_ , \g9832/_0_ , \g9833/_0_ , \g9835/_0_ , \g9836/_0_ , \g9837/_0_ , \g9838/_0_ , \g9839/_0_ , \g9840/_0_ , \g9841/_0_ , \g9842/_0_ , \g9844/_0_ , \g9845/_0_ , \g9846/_0_ , \g9848/_0_ , \g9849/_0_ , \g9850/_0_ , \g9851/_0_ , \g9853/_0_ , \g9854/_0_ , \g9855/_0_ , \g9856/_0_ , \g9857/_0_ , \g9858/_0_ , \g9859/_0_ , \g9860/_0_ , \g9862/_0_ , \g9863/_0_ , \g9864/_0_ , \g9865/_0_ , \g9867/_0_ , \g9868/_0_ , \g9876/_0_ , \g9877/_0_ , \g9878/_0_ , \g9879/_0_ , \g9880/_0_ , \g9881/_0_ , \g9898/_0_ , \g9900/_0_ , \g9901/_0_ , \g9902/_0_ , \g9903/_0_ , \g9904/_0_ , \g9905/_0_ , \g9906/_0_ , \g9907/_0_ , \g9908/_0_ , \g9909/_0_ , \g9910/_0_ , \g9911/_0_ , \g9912/_0_ , \g9913/_0_ , \g9914/_0_ , \g9915/_0_ , \g9916/_0_ , \g9917/_0_ , \g9918/_0_ , \g9919/_0_ , \g992/_0_ , \g9920/_0_ , \g9921/_0_ , \g9922/_0_ , \g9923/_0_ , \g9924/_0_ , \g9925/_0_ , \g9926/_0_ , \g9927/_0_ , \g9928/_0_ , \g9929/_0_ , \g9930/_0_ , \g9931/_0_ , \g9932/_0_ , \g9933/_0_ , \g9934/_0_ , \g9935/_0_ , \g9936/_0_ , \g9937/_0_ , \g9938/_0_ , \g9939/_0_ , \g9940/_0_ , \g9941/_0_ , \g9942/_0_ , \g9943/_0_ , \g9944/_0_ , \g9945/_0_ , \g9946/_0_ , \g9947/_0_ , \g9948/_0_ , \g9949/_0_ , \g9950/_0_ , \g9951/_0_ , \g9952/_0_ , \g9953/_0_ , \g9954/_0_ , \g9955/_0_ , \g9956/_0_ , \g9957/_0_ , \g9958/_0_ , \g9959/_0_ , \g9960/_0_ , \g9961/_0_ , \g9962/_0_ , \g9963/_0_ , \g9964/_0_ , \g9965/_0_ , \g9966/_0_ , \g9967/_0_ , \g9968/_0_ , \g9969/_0_ , \g9970/_0_ , \g9971/_0_ , \g9972/_0_ , \g9973/_0_ , \g9974/_0_ , \g9975/_0_ , \g9976/_0_ , \g9977/_0_ , \g9978/_0_ , \g9979/_0_ , \g9980/_0_ , \g9981/_0_ , \g9982/_0_ , \g9983/_0_ , \g9984/_0_ , \g9985/_0_ , \g9987/_0_ , \g9988/_0_ , \g9989/_0_ , \g999/_0_ , \g9990/_0_ , \g9991/_0_ , \g9992/_0_ , \g9993/_0_ , \g9994/_0_ , \g9995/_0_ , \g9996/_0_ , \g9997/_0_ , \g9998/_0_ , \g9999/_0_ , \idma_IDMA_boot_reg/NET0131_reg_syn_3 , \memc_EXTC_Eg_reg/NET0131 , \memc_EXTC_Eg_reg/NET0131_reg_syn_3 , \memc_EXTC_Eg_reg/n0 , \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3 , \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3 , \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3 , \sice_GO_NXi_reg/NET0131_reg_syn_3 , \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3 , \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3 , \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3 , \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3 );
	input \CM_rd0[0]_pad  ;
	input \CM_rd0[10]_pad  ;
	input \CM_rd0[11]_pad  ;
	input \CM_rd0[12]_pad  ;
	input \CM_rd0[13]_pad  ;
	input \CM_rd0[14]_pad  ;
	input \CM_rd0[15]_pad  ;
	input \CM_rd0[16]_pad  ;
	input \CM_rd0[17]_pad  ;
	input \CM_rd0[18]_pad  ;
	input \CM_rd0[19]_pad  ;
	input \CM_rd0[1]_pad  ;
	input \CM_rd0[20]_pad  ;
	input \CM_rd0[21]_pad  ;
	input \CM_rd0[22]_pad  ;
	input \CM_rd0[23]_pad  ;
	input \CM_rd0[2]_pad  ;
	input \CM_rd0[3]_pad  ;
	input \CM_rd0[4]_pad  ;
	input \CM_rd0[5]_pad  ;
	input \CM_rd0[6]_pad  ;
	input \CM_rd0[7]_pad  ;
	input \CM_rd0[8]_pad  ;
	input \CM_rd0[9]_pad  ;
	input \CM_rd1[0]_pad  ;
	input \CM_rd1[10]_pad  ;
	input \CM_rd1[11]_pad  ;
	input \CM_rd1[12]_pad  ;
	input \CM_rd1[13]_pad  ;
	input \CM_rd1[14]_pad  ;
	input \CM_rd1[15]_pad  ;
	input \CM_rd1[16]_pad  ;
	input \CM_rd1[17]_pad  ;
	input \CM_rd1[18]_pad  ;
	input \CM_rd1[19]_pad  ;
	input \CM_rd1[1]_pad  ;
	input \CM_rd1[20]_pad  ;
	input \CM_rd1[21]_pad  ;
	input \CM_rd1[22]_pad  ;
	input \CM_rd1[23]_pad  ;
	input \CM_rd1[2]_pad  ;
	input \CM_rd1[3]_pad  ;
	input \CM_rd1[4]_pad  ;
	input \CM_rd1[5]_pad  ;
	input \CM_rd1[6]_pad  ;
	input \CM_rd1[7]_pad  ;
	input \CM_rd1[8]_pad  ;
	input \CM_rd1[9]_pad  ;
	input \CM_rd2[0]_pad  ;
	input \CM_rd2[10]_pad  ;
	input \CM_rd2[11]_pad  ;
	input \CM_rd2[12]_pad  ;
	input \CM_rd2[13]_pad  ;
	input \CM_rd2[14]_pad  ;
	input \CM_rd2[15]_pad  ;
	input \CM_rd2[16]_pad  ;
	input \CM_rd2[17]_pad  ;
	input \CM_rd2[18]_pad  ;
	input \CM_rd2[19]_pad  ;
	input \CM_rd2[1]_pad  ;
	input \CM_rd2[20]_pad  ;
	input \CM_rd2[21]_pad  ;
	input \CM_rd2[22]_pad  ;
	input \CM_rd2[23]_pad  ;
	input \CM_rd2[2]_pad  ;
	input \CM_rd2[3]_pad  ;
	input \CM_rd2[4]_pad  ;
	input \CM_rd2[5]_pad  ;
	input \CM_rd2[6]_pad  ;
	input \CM_rd2[7]_pad  ;
	input \CM_rd2[8]_pad  ;
	input \CM_rd2[9]_pad  ;
	input \CM_rd3[0]_pad  ;
	input \CM_rd3[10]_pad  ;
	input \CM_rd3[11]_pad  ;
	input \CM_rd3[12]_pad  ;
	input \CM_rd3[13]_pad  ;
	input \CM_rd3[14]_pad  ;
	input \CM_rd3[15]_pad  ;
	input \CM_rd3[16]_pad  ;
	input \CM_rd3[17]_pad  ;
	input \CM_rd3[18]_pad  ;
	input \CM_rd3[19]_pad  ;
	input \CM_rd3[1]_pad  ;
	input \CM_rd3[20]_pad  ;
	input \CM_rd3[21]_pad  ;
	input \CM_rd3[22]_pad  ;
	input \CM_rd3[23]_pad  ;
	input \CM_rd3[2]_pad  ;
	input \CM_rd3[3]_pad  ;
	input \CM_rd3[4]_pad  ;
	input \CM_rd3[5]_pad  ;
	input \CM_rd3[6]_pad  ;
	input \CM_rd3[7]_pad  ;
	input \CM_rd3[8]_pad  ;
	input \CM_rd3[9]_pad  ;
	input \CM_rd4[0]_pad  ;
	input \CM_rd4[10]_pad  ;
	input \CM_rd4[11]_pad  ;
	input \CM_rd4[12]_pad  ;
	input \CM_rd4[13]_pad  ;
	input \CM_rd4[14]_pad  ;
	input \CM_rd4[15]_pad  ;
	input \CM_rd4[16]_pad  ;
	input \CM_rd4[17]_pad  ;
	input \CM_rd4[18]_pad  ;
	input \CM_rd4[19]_pad  ;
	input \CM_rd4[1]_pad  ;
	input \CM_rd4[20]_pad  ;
	input \CM_rd4[21]_pad  ;
	input \CM_rd4[22]_pad  ;
	input \CM_rd4[23]_pad  ;
	input \CM_rd4[2]_pad  ;
	input \CM_rd4[3]_pad  ;
	input \CM_rd4[4]_pad  ;
	input \CM_rd4[5]_pad  ;
	input \CM_rd4[6]_pad  ;
	input \CM_rd4[7]_pad  ;
	input \CM_rd4[8]_pad  ;
	input \CM_rd4[9]_pad  ;
	input \CM_rd5[0]_pad  ;
	input \CM_rd5[10]_pad  ;
	input \CM_rd5[11]_pad  ;
	input \CM_rd5[12]_pad  ;
	input \CM_rd5[13]_pad  ;
	input \CM_rd5[14]_pad  ;
	input \CM_rd5[15]_pad  ;
	input \CM_rd5[16]_pad  ;
	input \CM_rd5[17]_pad  ;
	input \CM_rd5[18]_pad  ;
	input \CM_rd5[19]_pad  ;
	input \CM_rd5[1]_pad  ;
	input \CM_rd5[20]_pad  ;
	input \CM_rd5[21]_pad  ;
	input \CM_rd5[22]_pad  ;
	input \CM_rd5[23]_pad  ;
	input \CM_rd5[2]_pad  ;
	input \CM_rd5[3]_pad  ;
	input \CM_rd5[4]_pad  ;
	input \CM_rd5[5]_pad  ;
	input \CM_rd5[6]_pad  ;
	input \CM_rd5[7]_pad  ;
	input \CM_rd5[8]_pad  ;
	input \CM_rd5[9]_pad  ;
	input \CM_rd6[0]_pad  ;
	input \CM_rd6[10]_pad  ;
	input \CM_rd6[11]_pad  ;
	input \CM_rd6[12]_pad  ;
	input \CM_rd6[13]_pad  ;
	input \CM_rd6[14]_pad  ;
	input \CM_rd6[15]_pad  ;
	input \CM_rd6[16]_pad  ;
	input \CM_rd6[17]_pad  ;
	input \CM_rd6[18]_pad  ;
	input \CM_rd6[19]_pad  ;
	input \CM_rd6[1]_pad  ;
	input \CM_rd6[20]_pad  ;
	input \CM_rd6[21]_pad  ;
	input \CM_rd6[22]_pad  ;
	input \CM_rd6[23]_pad  ;
	input \CM_rd6[2]_pad  ;
	input \CM_rd6[3]_pad  ;
	input \CM_rd6[4]_pad  ;
	input \CM_rd6[5]_pad  ;
	input \CM_rd6[6]_pad  ;
	input \CM_rd6[7]_pad  ;
	input \CM_rd6[8]_pad  ;
	input \CM_rd6[9]_pad  ;
	input \CM_rd7[0]_pad  ;
	input \CM_rd7[10]_pad  ;
	input \CM_rd7[11]_pad  ;
	input \CM_rd7[12]_pad  ;
	input \CM_rd7[13]_pad  ;
	input \CM_rd7[14]_pad  ;
	input \CM_rd7[15]_pad  ;
	input \CM_rd7[16]_pad  ;
	input \CM_rd7[17]_pad  ;
	input \CM_rd7[18]_pad  ;
	input \CM_rd7[19]_pad  ;
	input \CM_rd7[1]_pad  ;
	input \CM_rd7[20]_pad  ;
	input \CM_rd7[21]_pad  ;
	input \CM_rd7[22]_pad  ;
	input \CM_rd7[23]_pad  ;
	input \CM_rd7[2]_pad  ;
	input \CM_rd7[3]_pad  ;
	input \CM_rd7[4]_pad  ;
	input \CM_rd7[5]_pad  ;
	input \CM_rd7[6]_pad  ;
	input \CM_rd7[7]_pad  ;
	input \CM_rd7[8]_pad  ;
	input \CM_rd7[9]_pad  ;
	input \CM_rdm[0]_pad  ;
	input \CM_rdm[10]_pad  ;
	input \CM_rdm[11]_pad  ;
	input \CM_rdm[12]_pad  ;
	input \CM_rdm[13]_pad  ;
	input \CM_rdm[14]_pad  ;
	input \CM_rdm[15]_pad  ;
	input \CM_rdm[16]_pad  ;
	input \CM_rdm[17]_pad  ;
	input \CM_rdm[18]_pad  ;
	input \CM_rdm[19]_pad  ;
	input \CM_rdm[1]_pad  ;
	input \CM_rdm[20]_pad  ;
	input \CM_rdm[21]_pad  ;
	input \CM_rdm[22]_pad  ;
	input \CM_rdm[23]_pad  ;
	input \CM_rdm[2]_pad  ;
	input \CM_rdm[3]_pad  ;
	input \CM_rdm[4]_pad  ;
	input \CM_rdm[5]_pad  ;
	input \CM_rdm[6]_pad  ;
	input \CM_rdm[7]_pad  ;
	input \CM_rdm[8]_pad  ;
	input \CM_rdm[9]_pad  ;
	input \DM_rd0[0]_pad  ;
	input \DM_rd0[10]_pad  ;
	input \DM_rd0[11]_pad  ;
	input \DM_rd0[12]_pad  ;
	input \DM_rd0[13]_pad  ;
	input \DM_rd0[14]_pad  ;
	input \DM_rd0[15]_pad  ;
	input \DM_rd0[1]_pad  ;
	input \DM_rd0[2]_pad  ;
	input \DM_rd0[3]_pad  ;
	input \DM_rd0[4]_pad  ;
	input \DM_rd0[5]_pad  ;
	input \DM_rd0[6]_pad  ;
	input \DM_rd0[7]_pad  ;
	input \DM_rd0[8]_pad  ;
	input \DM_rd0[9]_pad  ;
	input \DM_rd1[0]_pad  ;
	input \DM_rd1[10]_pad  ;
	input \DM_rd1[11]_pad  ;
	input \DM_rd1[12]_pad  ;
	input \DM_rd1[13]_pad  ;
	input \DM_rd1[14]_pad  ;
	input \DM_rd1[15]_pad  ;
	input \DM_rd1[1]_pad  ;
	input \DM_rd1[2]_pad  ;
	input \DM_rd1[3]_pad  ;
	input \DM_rd1[4]_pad  ;
	input \DM_rd1[5]_pad  ;
	input \DM_rd1[6]_pad  ;
	input \DM_rd1[7]_pad  ;
	input \DM_rd1[8]_pad  ;
	input \DM_rd1[9]_pad  ;
	input \DM_rd2[0]_pad  ;
	input \DM_rd2[10]_pad  ;
	input \DM_rd2[11]_pad  ;
	input \DM_rd2[12]_pad  ;
	input \DM_rd2[13]_pad  ;
	input \DM_rd2[14]_pad  ;
	input \DM_rd2[15]_pad  ;
	input \DM_rd2[1]_pad  ;
	input \DM_rd2[2]_pad  ;
	input \DM_rd2[3]_pad  ;
	input \DM_rd2[4]_pad  ;
	input \DM_rd2[5]_pad  ;
	input \DM_rd2[6]_pad  ;
	input \DM_rd2[7]_pad  ;
	input \DM_rd2[8]_pad  ;
	input \DM_rd2[9]_pad  ;
	input \DM_rd3[0]_pad  ;
	input \DM_rd3[10]_pad  ;
	input \DM_rd3[11]_pad  ;
	input \DM_rd3[12]_pad  ;
	input \DM_rd3[13]_pad  ;
	input \DM_rd3[14]_pad  ;
	input \DM_rd3[15]_pad  ;
	input \DM_rd3[1]_pad  ;
	input \DM_rd3[2]_pad  ;
	input \DM_rd3[3]_pad  ;
	input \DM_rd3[4]_pad  ;
	input \DM_rd3[5]_pad  ;
	input \DM_rd3[6]_pad  ;
	input \DM_rd3[7]_pad  ;
	input \DM_rd3[8]_pad  ;
	input \DM_rd3[9]_pad  ;
	input \DM_rd4[0]_pad  ;
	input \DM_rd4[10]_pad  ;
	input \DM_rd4[11]_pad  ;
	input \DM_rd4[12]_pad  ;
	input \DM_rd4[13]_pad  ;
	input \DM_rd4[14]_pad  ;
	input \DM_rd4[15]_pad  ;
	input \DM_rd4[1]_pad  ;
	input \DM_rd4[2]_pad  ;
	input \DM_rd4[3]_pad  ;
	input \DM_rd4[4]_pad  ;
	input \DM_rd4[5]_pad  ;
	input \DM_rd4[6]_pad  ;
	input \DM_rd4[7]_pad  ;
	input \DM_rd4[8]_pad  ;
	input \DM_rd4[9]_pad  ;
	input \DM_rd5[0]_pad  ;
	input \DM_rd5[10]_pad  ;
	input \DM_rd5[11]_pad  ;
	input \DM_rd5[12]_pad  ;
	input \DM_rd5[13]_pad  ;
	input \DM_rd5[14]_pad  ;
	input \DM_rd5[15]_pad  ;
	input \DM_rd5[1]_pad  ;
	input \DM_rd5[2]_pad  ;
	input \DM_rd5[3]_pad  ;
	input \DM_rd5[4]_pad  ;
	input \DM_rd5[5]_pad  ;
	input \DM_rd5[6]_pad  ;
	input \DM_rd5[7]_pad  ;
	input \DM_rd5[8]_pad  ;
	input \DM_rd5[9]_pad  ;
	input \DM_rd6[0]_pad  ;
	input \DM_rd6[10]_pad  ;
	input \DM_rd6[11]_pad  ;
	input \DM_rd6[12]_pad  ;
	input \DM_rd6[13]_pad  ;
	input \DM_rd6[14]_pad  ;
	input \DM_rd6[15]_pad  ;
	input \DM_rd6[1]_pad  ;
	input \DM_rd6[2]_pad  ;
	input \DM_rd6[3]_pad  ;
	input \DM_rd6[4]_pad  ;
	input \DM_rd6[5]_pad  ;
	input \DM_rd6[6]_pad  ;
	input \DM_rd6[7]_pad  ;
	input \DM_rd6[8]_pad  ;
	input \DM_rd6[9]_pad  ;
	input \DM_rd7[0]_pad  ;
	input \DM_rd7[10]_pad  ;
	input \DM_rd7[11]_pad  ;
	input \DM_rd7[12]_pad  ;
	input \DM_rd7[13]_pad  ;
	input \DM_rd7[14]_pad  ;
	input \DM_rd7[15]_pad  ;
	input \DM_rd7[1]_pad  ;
	input \DM_rd7[2]_pad  ;
	input \DM_rd7[3]_pad  ;
	input \DM_rd7[4]_pad  ;
	input \DM_rd7[5]_pad  ;
	input \DM_rd7[6]_pad  ;
	input \DM_rd7[7]_pad  ;
	input \DM_rd7[8]_pad  ;
	input \DM_rd7[9]_pad  ;
	input \DM_rdm[0]_pad  ;
	input \DM_rdm[10]_pad  ;
	input \DM_rdm[11]_pad  ;
	input \DM_rdm[12]_pad  ;
	input \DM_rdm[13]_pad  ;
	input \DM_rdm[14]_pad  ;
	input \DM_rdm[15]_pad  ;
	input \DM_rdm[1]_pad  ;
	input \DM_rdm[2]_pad  ;
	input \DM_rdm[3]_pad  ;
	input \DM_rdm[4]_pad  ;
	input \DM_rdm[5]_pad  ;
	input \DM_rdm[6]_pad  ;
	input \DM_rdm[7]_pad  ;
	input \DM_rdm[8]_pad  ;
	input \DM_rdm[9]_pad  ;
	input IACKn_pad ;
	input \IRFS0_pad  ;
	input \IRFS1_pad  ;
	input \ISCLK0_pad  ;
	input \ISCLK1_pad  ;
	input \ITFS0_pad  ;
	input \ITFS1_pad  ;
	input \PIO_oe[0]_pad  ;
	input \PIO_oe[10]_pad  ;
	input \PIO_oe[11]_pad  ;
	input \PIO_oe[1]_pad  ;
	input \PIO_oe[2]_pad  ;
	input \PIO_oe[3]_pad  ;
	input \PIO_oe[4]_pad  ;
	input \PIO_oe[5]_pad  ;
	input \PIO_oe[6]_pad  ;
	input \PIO_oe[7]_pad  ;
	input \PIO_oe[8]_pad  ;
	input \PIO_oe[9]_pad  ;
	input \PIO_out[0]_pad  ;
	input \PIO_out[10]_pad  ;
	input \PIO_out[11]_pad  ;
	input \PIO_out[1]_pad  ;
	input \PIO_out[2]_pad  ;
	input \PIO_out[3]_pad  ;
	input \PIO_out[4]_pad  ;
	input \PIO_out[5]_pad  ;
	input \PIO_out[6]_pad  ;
	input \PIO_out[7]_pad  ;
	input \PIO_out[8]_pad  ;
	input \PIO_out[9]_pad  ;
	input PM_bdry_sel_pad ;
	input \PM_rd0[0]_pad  ;
	input \PM_rd0[10]_pad  ;
	input \PM_rd0[11]_pad  ;
	input \PM_rd0[12]_pad  ;
	input \PM_rd0[13]_pad  ;
	input \PM_rd0[14]_pad  ;
	input \PM_rd0[15]_pad  ;
	input \PM_rd0[1]_pad  ;
	input \PM_rd0[2]_pad  ;
	input \PM_rd0[3]_pad  ;
	input \PM_rd0[4]_pad  ;
	input \PM_rd0[5]_pad  ;
	input \PM_rd0[6]_pad  ;
	input \PM_rd0[7]_pad  ;
	input \PM_rd0[8]_pad  ;
	input \PM_rd0[9]_pad  ;
	input \PM_rd1[0]_pad  ;
	input \PM_rd1[10]_pad  ;
	input \PM_rd1[11]_pad  ;
	input \PM_rd1[12]_pad  ;
	input \PM_rd1[13]_pad  ;
	input \PM_rd1[14]_pad  ;
	input \PM_rd1[15]_pad  ;
	input \PM_rd1[1]_pad  ;
	input \PM_rd1[2]_pad  ;
	input \PM_rd1[3]_pad  ;
	input \PM_rd1[4]_pad  ;
	input \PM_rd1[5]_pad  ;
	input \PM_rd1[6]_pad  ;
	input \PM_rd1[7]_pad  ;
	input \PM_rd1[8]_pad  ;
	input \PM_rd1[9]_pad  ;
	input \PM_rd2[0]_pad  ;
	input \PM_rd2[10]_pad  ;
	input \PM_rd2[11]_pad  ;
	input \PM_rd2[12]_pad  ;
	input \PM_rd2[13]_pad  ;
	input \PM_rd2[14]_pad  ;
	input \PM_rd2[15]_pad  ;
	input \PM_rd2[1]_pad  ;
	input \PM_rd2[2]_pad  ;
	input \PM_rd2[3]_pad  ;
	input \PM_rd2[4]_pad  ;
	input \PM_rd2[5]_pad  ;
	input \PM_rd2[6]_pad  ;
	input \PM_rd2[7]_pad  ;
	input \PM_rd2[8]_pad  ;
	input \PM_rd2[9]_pad  ;
	input \PM_rd3[0]_pad  ;
	input \PM_rd3[10]_pad  ;
	input \PM_rd3[11]_pad  ;
	input \PM_rd3[12]_pad  ;
	input \PM_rd3[13]_pad  ;
	input \PM_rd3[14]_pad  ;
	input \PM_rd3[15]_pad  ;
	input \PM_rd3[1]_pad  ;
	input \PM_rd3[2]_pad  ;
	input \PM_rd3[3]_pad  ;
	input \PM_rd3[4]_pad  ;
	input \PM_rd3[5]_pad  ;
	input \PM_rd3[6]_pad  ;
	input \PM_rd3[7]_pad  ;
	input \PM_rd3[8]_pad  ;
	input \PM_rd3[9]_pad  ;
	input \PM_rd4[0]_pad  ;
	input \PM_rd4[10]_pad  ;
	input \PM_rd4[11]_pad  ;
	input \PM_rd4[12]_pad  ;
	input \PM_rd4[13]_pad  ;
	input \PM_rd4[14]_pad  ;
	input \PM_rd4[15]_pad  ;
	input \PM_rd4[1]_pad  ;
	input \PM_rd4[2]_pad  ;
	input \PM_rd4[3]_pad  ;
	input \PM_rd4[4]_pad  ;
	input \PM_rd4[5]_pad  ;
	input \PM_rd4[6]_pad  ;
	input \PM_rd4[7]_pad  ;
	input \PM_rd4[8]_pad  ;
	input \PM_rd4[9]_pad  ;
	input \PM_rd5[0]_pad  ;
	input \PM_rd5[10]_pad  ;
	input \PM_rd5[11]_pad  ;
	input \PM_rd5[12]_pad  ;
	input \PM_rd5[13]_pad  ;
	input \PM_rd5[14]_pad  ;
	input \PM_rd5[15]_pad  ;
	input \PM_rd5[1]_pad  ;
	input \PM_rd5[2]_pad  ;
	input \PM_rd5[3]_pad  ;
	input \PM_rd5[4]_pad  ;
	input \PM_rd5[5]_pad  ;
	input \PM_rd5[6]_pad  ;
	input \PM_rd5[7]_pad  ;
	input \PM_rd5[8]_pad  ;
	input \PM_rd5[9]_pad  ;
	input \PM_rd6[0]_pad  ;
	input \PM_rd6[10]_pad  ;
	input \PM_rd6[11]_pad  ;
	input \PM_rd6[12]_pad  ;
	input \PM_rd6[13]_pad  ;
	input \PM_rd6[14]_pad  ;
	input \PM_rd6[15]_pad  ;
	input \PM_rd6[1]_pad  ;
	input \PM_rd6[2]_pad  ;
	input \PM_rd6[3]_pad  ;
	input \PM_rd6[4]_pad  ;
	input \PM_rd6[5]_pad  ;
	input \PM_rd6[6]_pad  ;
	input \PM_rd6[7]_pad  ;
	input \PM_rd6[8]_pad  ;
	input \PM_rd6[9]_pad  ;
	input \PM_rd7[0]_pad  ;
	input \PM_rd7[10]_pad  ;
	input \PM_rd7[11]_pad  ;
	input \PM_rd7[12]_pad  ;
	input \PM_rd7[13]_pad  ;
	input \PM_rd7[14]_pad  ;
	input \PM_rd7[15]_pad  ;
	input \PM_rd7[1]_pad  ;
	input \PM_rd7[2]_pad  ;
	input \PM_rd7[3]_pad  ;
	input \PM_rd7[4]_pad  ;
	input \PM_rd7[5]_pad  ;
	input \PM_rd7[6]_pad  ;
	input \PM_rd7[7]_pad  ;
	input \PM_rd7[8]_pad  ;
	input \PM_rd7[9]_pad  ;
	input PWDACK_pad ;
	input T_BMODE_pad ;
	input T_BRn_pad ;
	input T_CLKI_OSC_pad ;
	input T_CLKI_PLL_pad ;
	input \T_ED[0]_pad  ;
	input \T_ED[10]_pad  ;
	input \T_ED[11]_pad  ;
	input \T_ED[12]_pad  ;
	input \T_ED[13]_pad  ;
	input \T_ED[14]_pad  ;
	input \T_ED[15]_pad  ;
	input \T_ED[1]_pad  ;
	input \T_ED[2]_pad  ;
	input \T_ED[3]_pad  ;
	input \T_ED[4]_pad  ;
	input \T_ED[5]_pad  ;
	input \T_ED[6]_pad  ;
	input \T_ED[7]_pad  ;
	input \T_ED[8]_pad  ;
	input \T_ED[9]_pad  ;
	input T_ICE_RSTn_pad ;
	input T_ID_pad ;
	input T_IMS_pad ;
	input T_IRDn_pad ;
	input \T_IRQ0n_pad  ;
	input \T_IRQ1n_pad  ;
	input \T_IRQ2n_pad  ;
	input \T_IRQE0n_pad  ;
	input \T_IRQE1n_pad  ;
	input \T_IRQL1n_pad  ;
	input T_ISn_pad ;
	input T_IWRn_pad ;
	input T_MMAP_pad ;
	input \T_PIOin[0]_pad  ;
	input \T_PIOin[10]_pad  ;
	input \T_PIOin[11]_pad  ;
	input \T_PIOin[1]_pad  ;
	input \T_PIOin[2]_pad  ;
	input \T_PIOin[3]_pad  ;
	input \T_PIOin[4]_pad  ;
	input \T_PIOin[5]_pad  ;
	input \T_PIOin[6]_pad  ;
	input \T_PIOin[7]_pad  ;
	input \T_PIOin[8]_pad  ;
	input \T_PIOin[9]_pad  ;
	input T_PWDn_pad ;
	input \T_RD0_pad  ;
	input \T_RD1_pad  ;
	input \T_RFS0_pad  ;
	input \T_RFS1_pad  ;
	input T_RSTn_pad ;
	input \T_SCLK0_pad  ;
	input \T_SCLK1_pad  ;
	input T_Sel_PLL_pad ;
	input \T_TFS0_pad  ;
	input \T_TFS1_pad  ;
	input \T_TMODE[0]_pad  ;
	input \T_TMODE[1]_pad  ;
	input \auctl_BSack_reg/NET0131  ;
	input \auctl_DSack_reg/NET0131  ;
	input \auctl_R0Sack_reg/NET0131  ;
	input \auctl_R1Sack_reg/NET0131  ;
	input \auctl_RST_reg/P0001  ;
	input \auctl_STEAL_reg/NET0131  ;
	input \auctl_T0Sack_reg/NET0131  ;
	input \auctl_T1Sack_reg/NET0131  ;
	input \bdma_BCTL_reg[0]/NET0131  ;
	input \bdma_BCTL_reg[10]/NET0131  ;
	input \bdma_BCTL_reg[11]/NET0131  ;
	input \bdma_BCTL_reg[12]/NET0131  ;
	input \bdma_BCTL_reg[13]/NET0131  ;
	input \bdma_BCTL_reg[14]/NET0131  ;
	input \bdma_BCTL_reg[15]/NET0131  ;
	input \bdma_BCTL_reg[1]/NET0131  ;
	input \bdma_BCTL_reg[2]/NET0131  ;
	input \bdma_BCTL_reg[3]/NET0131  ;
	input \bdma_BCTL_reg[4]/NET0131  ;
	input \bdma_BCTL_reg[5]/NET0131  ;
	input \bdma_BCTL_reg[6]/NET0131  ;
	input \bdma_BCTL_reg[7]/NET0131  ;
	input \bdma_BCTL_reg[8]/NET0131  ;
	input \bdma_BCTL_reg[9]/NET0131  ;
	input \bdma_BDMA_boot_reg/NET0131_reg_syn_10  ;
	input \bdma_BDMA_boot_reg/NET0131_reg_syn_2  ;
	input \bdma_BDMA_boot_reg/NET0131_reg_syn_8  ;
	input \bdma_BDMAmode_reg/NET0131  ;
	input \bdma_BEAD_reg[0]/NET0131  ;
	input \bdma_BEAD_reg[10]/NET0131  ;
	input \bdma_BEAD_reg[11]/NET0131  ;
	input \bdma_BEAD_reg[12]/NET0131  ;
	input \bdma_BEAD_reg[13]/NET0131  ;
	input \bdma_BEAD_reg[1]/NET0131  ;
	input \bdma_BEAD_reg[2]/NET0131  ;
	input \bdma_BEAD_reg[3]/NET0131  ;
	input \bdma_BEAD_reg[4]/NET0131  ;
	input \bdma_BEAD_reg[5]/NET0131  ;
	input \bdma_BEAD_reg[6]/NET0131  ;
	input \bdma_BEAD_reg[7]/NET0131  ;
	input \bdma_BEAD_reg[8]/NET0131  ;
	input \bdma_BEAD_reg[9]/NET0131  ;
	input \bdma_BIAD_reg[0]/NET0131  ;
	input \bdma_BIAD_reg[10]/NET0131  ;
	input \bdma_BIAD_reg[11]/NET0131  ;
	input \bdma_BIAD_reg[12]/NET0131  ;
	input \bdma_BIAD_reg[13]/NET0131  ;
	input \bdma_BIAD_reg[1]/NET0131  ;
	input \bdma_BIAD_reg[2]/NET0131  ;
	input \bdma_BIAD_reg[3]/NET0131  ;
	input \bdma_BIAD_reg[4]/NET0131  ;
	input \bdma_BIAD_reg[5]/NET0131  ;
	input \bdma_BIAD_reg[6]/NET0131  ;
	input \bdma_BIAD_reg[7]/NET0131  ;
	input \bdma_BIAD_reg[8]/NET0131  ;
	input \bdma_BIAD_reg[9]/NET0131  ;
	input \bdma_BM_cyc_reg/P0001  ;
	input \bdma_BMcyc_del_reg/P0001  ;
	input \bdma_BOVL_reg[0]/NET0131  ;
	input \bdma_BOVL_reg[10]/NET0131  ;
	input \bdma_BOVL_reg[11]/NET0131  ;
	input \bdma_BOVL_reg[1]/NET0131  ;
	input \bdma_BOVL_reg[2]/NET0131  ;
	input \bdma_BOVL_reg[3]/NET0131  ;
	input \bdma_BOVL_reg[4]/NET0131  ;
	input \bdma_BOVL_reg[5]/NET0131  ;
	input \bdma_BOVL_reg[6]/NET0131  ;
	input \bdma_BOVL_reg[7]/NET0131  ;
	input \bdma_BOVL_reg[8]/NET0131  ;
	input \bdma_BOVL_reg[9]/NET0131  ;
	input \bdma_BRST_s2_reg/NET0131  ;
	input \bdma_BRdataBUF_reg[0]/P0001  ;
	input \bdma_BRdataBUF_reg[10]/P0001  ;
	input \bdma_BRdataBUF_reg[11]/P0001  ;
	input \bdma_BRdataBUF_reg[12]/P0001  ;
	input \bdma_BRdataBUF_reg[13]/P0001  ;
	input \bdma_BRdataBUF_reg[14]/P0001  ;
	input \bdma_BRdataBUF_reg[15]/P0001  ;
	input \bdma_BRdataBUF_reg[16]/P0001  ;
	input \bdma_BRdataBUF_reg[17]/P0001  ;
	input \bdma_BRdataBUF_reg[18]/P0001  ;
	input \bdma_BRdataBUF_reg[19]/P0001  ;
	input \bdma_BRdataBUF_reg[1]/P0001  ;
	input \bdma_BRdataBUF_reg[20]/P0001  ;
	input \bdma_BRdataBUF_reg[21]/P0001  ;
	input \bdma_BRdataBUF_reg[22]/P0001  ;
	input \bdma_BRdataBUF_reg[23]/P0001  ;
	input \bdma_BRdataBUF_reg[2]/P0001  ;
	input \bdma_BRdataBUF_reg[3]/P0001  ;
	input \bdma_BRdataBUF_reg[4]/P0001  ;
	input \bdma_BRdataBUF_reg[5]/P0001  ;
	input \bdma_BRdataBUF_reg[6]/P0001  ;
	input \bdma_BRdataBUF_reg[7]/P0001  ;
	input \bdma_BRdataBUF_reg[8]/P0001  ;
	input \bdma_BRdataBUF_reg[9]/P0001  ;
	input \bdma_BSreq_reg/NET0131  ;
	input \bdma_BWCOUNT_reg[0]/NET0131  ;
	input \bdma_BWCOUNT_reg[10]/NET0131  ;
	input \bdma_BWCOUNT_reg[11]/NET0131  ;
	input \bdma_BWCOUNT_reg[12]/NET0131  ;
	input \bdma_BWCOUNT_reg[13]/NET0131  ;
	input \bdma_BWCOUNT_reg[1]/NET0131  ;
	input \bdma_BWCOUNT_reg[2]/NET0131  ;
	input \bdma_BWCOUNT_reg[3]/NET0131  ;
	input \bdma_BWCOUNT_reg[4]/NET0131  ;
	input \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2  ;
	input \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8  ;
	input \bdma_BWCOUNT_reg[6]/NET0131  ;
	input \bdma_BWCOUNT_reg[7]/NET0131  ;
	input \bdma_BWCOUNT_reg[8]/NET0131  ;
	input \bdma_BWCOUNT_reg[9]/NET0131  ;
	input \bdma_BWRn_reg/NET0131  ;
	input \bdma_BWcnt_reg[0]/NET0131  ;
	input \bdma_BWcnt_reg[1]/NET0131  ;
	input \bdma_BWcnt_reg[2]/NET0131  ;
	input \bdma_BWcnt_reg[3]/NET0131  ;
	input \bdma_BWcnt_reg[4]/NET0131  ;
	input \bdma_BWdataBUF_h_reg[0]/P0001  ;
	input \bdma_BWdataBUF_h_reg[10]/P0001  ;
	input \bdma_BWdataBUF_h_reg[11]/P0001  ;
	input \bdma_BWdataBUF_h_reg[12]/P0001  ;
	input \bdma_BWdataBUF_h_reg[13]/P0001  ;
	input \bdma_BWdataBUF_h_reg[14]/P0001  ;
	input \bdma_BWdataBUF_h_reg[15]/P0001  ;
	input \bdma_BWdataBUF_h_reg[16]/P0001  ;
	input \bdma_BWdataBUF_h_reg[17]/P0001  ;
	input \bdma_BWdataBUF_h_reg[18]/P0001  ;
	input \bdma_BWdataBUF_h_reg[19]/P0001  ;
	input \bdma_BWdataBUF_h_reg[1]/P0001  ;
	input \bdma_BWdataBUF_h_reg[20]/P0001  ;
	input \bdma_BWdataBUF_h_reg[21]/P0001  ;
	input \bdma_BWdataBUF_h_reg[22]/P0001  ;
	input \bdma_BWdataBUF_h_reg[23]/P0001  ;
	input \bdma_BWdataBUF_h_reg[2]/P0001  ;
	input \bdma_BWdataBUF_h_reg[3]/P0001  ;
	input \bdma_BWdataBUF_h_reg[4]/P0001  ;
	input \bdma_BWdataBUF_h_reg[5]/P0001  ;
	input \bdma_BWdataBUF_h_reg[6]/P0001  ;
	input \bdma_BWdataBUF_h_reg[7]/P0001  ;
	input \bdma_BWdataBUF_h_reg[8]/P0001  ;
	input \bdma_BWdataBUF_h_reg[9]/P0001  ;
	input \bdma_BWdataBUF_reg[0]/P0001  ;
	input \bdma_BWdataBUF_reg[1]/P0001  ;
	input \bdma_BWdataBUF_reg[2]/P0001  ;
	input \bdma_BWdataBUF_reg[3]/P0001  ;
	input \bdma_BWdataBUF_reg[4]/P0001  ;
	input \bdma_BWdataBUF_reg[5]/P0001  ;
	input \bdma_BWdataBUF_reg[6]/P0001  ;
	input \bdma_BWdataBUF_reg[7]/P0001  ;
	input \bdma_CMcnt_reg[0]/NET0131  ;
	input \bdma_CMcnt_reg[1]/NET0131  ;
	input \bdma_DM_2nd_reg/NET0131  ;
	input \bdma_RST_pin_reg/P0001  ;
	input \bdma_WRlat_reg/P0001  ;
	input \clkc_Awake_reg/NET0131  ;
	input \clkc_CLKOUT_reg/NET0131  ;
	input \clkc_CTR_cnt_reg[0]/NET0131  ;
	input \clkc_CTR_cnt_reg[1]/NET0131  ;
	input \clkc_Cnt128_reg/NET0131  ;
	input \clkc_Cnt4096_reg/NET0131  ;
	input \clkc_Cnt4096_s1_reg/NET0131  ;
	input \clkc_Cnt4096_s2_reg/NET0131  ;
	input \clkc_DSPoff_reg/NET0131  ;
	input \clkc_OSCoff_reg/NET0131  ;
	input \clkc_OSCoff_set_reg/P0001  ;
	input \clkc_OUTcnt_reg[0]/NET0131  ;
	input \clkc_OUTcnt_reg[1]/NET0131  ;
	input \clkc_OUTcnt_reg[2]/NET0131  ;
	input \clkc_OUTcnt_reg[3]/NET0131  ;
	input \clkc_OUTcnt_reg[4]/NET0131  ;
	input \clkc_OUTcnt_reg[5]/NET0131  ;
	input \clkc_OUTcnt_reg[6]/NET0131  ;
	input \clkc_RSTtext_reg/P0001  ;
	input \clkc_SIDLE_s1_reg/NET0131  ;
	input \clkc_SIDLE_s2_reg/NET0131  ;
	input \clkc_SLEEP_reg/NET0131  ;
	input \clkc_STBY_reg/NET0131  ;
	input \clkc_STDcnt_reg[0]/NET0131  ;
	input \clkc_STDcnt_reg[10]/NET0131  ;
	input \clkc_STDcnt_reg[1]/NET0131  ;
	input \clkc_STDcnt_reg[2]/NET0131  ;
	input \clkc_STDcnt_reg[3]/NET0131  ;
	input \clkc_STDcnt_reg[4]/NET0131  ;
	input \clkc_STDcnt_reg[5]/NET0131  ;
	input \clkc_STDcnt_reg[6]/NET0131  ;
	input \clkc_STDcnt_reg[7]/NET0131  ;
	input \clkc_STDcnt_reg[8]/NET0131  ;
	input \clkc_STDcnt_reg[9]/NET0131  ;
	input \clkc_SlowDn_reg/NET0131  ;
	input \clkc_SlowDn_s1_reg/P0001  ;
	input \clkc_SlowDn_s2_reg/P0001  ;
	input \clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131  ;
	input \clkc_ckr_reg_DO_reg[0]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[10]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[11]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[12]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[13]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[14]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[15]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[1]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[2]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[3]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[4]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[5]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[6]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[7]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[8]/NET0131  ;
	input \clkc_ckr_reg_DO_reg[9]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[0]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[10]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[11]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[1]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[2]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[3]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[4]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[5]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[6]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[7]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[8]/NET0131  ;
	input \clkc_oscntr_reg_DO_reg[9]/NET0131  ;
	input \core_c_dec_ALUop_E_reg/P0001  ;
	input \core_c_dec_BR_Ed_reg/P0001  ;
	input \core_c_dec_Call_Ed_reg/P0001  ;
	input \core_c_dec_DIVQ_E_reg/P0001  ;
	input \core_c_dec_DIVS_E_reg/P0001  ;
	input \core_c_dec_DU_Eg_reg/P0001  ;
	input \core_c_dec_Double_E_reg/P0001  ;
	input \core_c_dec_Dummy_E_reg/NET0131  ;
	input \core_c_dec_EXIT_E_reg/P0001  ;
	input \core_c_dec_IDLE_Eg_reg/P0001  ;
	input \core_c_dec_IRE_reg[0]/NET0131  ;
	input \core_c_dec_IRE_reg[10]/NET0131  ;
	input \core_c_dec_IRE_reg[11]/NET0131  ;
	input \core_c_dec_IRE_reg[12]/NET0131  ;
	input \core_c_dec_IRE_reg[13]/NET0131  ;
	input \core_c_dec_IRE_reg[14]/NET0131  ;
	input \core_c_dec_IRE_reg[15]/NET0131  ;
	input \core_c_dec_IRE_reg[16]/NET0131  ;
	input \core_c_dec_IRE_reg[17]/NET0131  ;
	input \core_c_dec_IRE_reg[18]/NET0131  ;
	input \core_c_dec_IRE_reg[19]/NET0131  ;
	input \core_c_dec_IRE_reg[1]/NET0131  ;
	input \core_c_dec_IRE_reg[2]/NET0131  ;
	input \core_c_dec_IRE_reg[3]/NET0131  ;
	input \core_c_dec_IRE_reg[4]/NET0131  ;
	input \core_c_dec_IRE_reg[5]/NET0131  ;
	input \core_c_dec_IRE_reg[6]/NET0131  ;
	input \core_c_dec_IRE_reg[7]/NET0131  ;
	input \core_c_dec_IRE_reg[8]/NET0131  ;
	input \core_c_dec_IRE_reg[9]/NET0131  ;
	input \core_c_dec_IR_reg[0]/NET0131  ;
	input \core_c_dec_IR_reg[10]/NET0131  ;
	input \core_c_dec_IR_reg[11]/NET0131  ;
	input \core_c_dec_IR_reg[12]/NET0131  ;
	input \core_c_dec_IR_reg[13]/NET0131  ;
	input \core_c_dec_IR_reg[14]/NET0131  ;
	input \core_c_dec_IR_reg[15]/NET0131  ;
	input \core_c_dec_IR_reg[16]/NET0131  ;
	input \core_c_dec_IR_reg[17]/NET0131  ;
	input \core_c_dec_IR_reg[18]/NET0131  ;
	input \core_c_dec_IR_reg[19]/NET0131  ;
	input \core_c_dec_IR_reg[1]/NET0131  ;
	input \core_c_dec_IR_reg[20]/NET0131  ;
	input \core_c_dec_IR_reg[21]/NET0131  ;
	input \core_c_dec_IR_reg[22]/NET0131  ;
	input \core_c_dec_IR_reg[23]/NET0131  ;
	input \core_c_dec_IR_reg[2]/NET0131  ;
	input \core_c_dec_IR_reg[3]/NET0131  ;
	input \core_c_dec_IR_reg[4]/NET0131  ;
	input \core_c_dec_IR_reg[5]/NET0131  ;
	input \core_c_dec_IR_reg[6]/NET0131  ;
	input \core_c_dec_IR_reg[7]/NET0131  ;
	input \core_c_dec_IR_reg[8]/NET0131  ;
	input \core_c_dec_IR_reg[9]/NET0131  ;
	input \core_c_dec_Long_Cg_reg/P0001  ;
	input \core_c_dec_Long_Eg_reg/P0001  ;
	input \core_c_dec_MACdep_Eg_reg/P0001  ;
	input \core_c_dec_MACop_E_reg/P0001  ;
	input \core_c_dec_MFALU_Ei_reg/NET0131  ;
	input \core_c_dec_MFAR_E_reg/P0001  ;
	input \core_c_dec_MFASTAT_E_reg/P0001  ;
	input \core_c_dec_MFAX0_E_reg/P0001  ;
	input \core_c_dec_MFAX1_E_reg/P0001  ;
	input \core_c_dec_MFAY0_E_reg/P0001  ;
	input \core_c_dec_MFAY1_E_reg/P0001  ;
	input \core_c_dec_MFCNTR_E_reg/P0001  ;
	input \core_c_dec_MFDAG1_Ei_reg/NET0131  ;
	input \core_c_dec_MFDAG2_Ei_reg/NET0131  ;
	input \core_c_dec_MFDMOVL_E_reg/P0001  ;
	input \core_c_dec_MFICNTL_E_reg/P0001  ;
	input \core_c_dec_MFIDR_E_reg/P0001  ;
	input \core_c_dec_MFIMASK_E_reg/P0001  ;
	input \core_c_dec_MFIreg_E_reg[0]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[1]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[2]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[3]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[4]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[5]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[6]/P0001  ;
	input \core_c_dec_MFIreg_E_reg[7]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[0]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[1]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[2]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[3]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[4]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[5]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[6]/P0001  ;
	input \core_c_dec_MFLreg_E_reg[7]/P0001  ;
	input \core_c_dec_MFMAC_Ei_reg/NET0131  ;
	input \core_c_dec_MFMR0_E_reg/P0001  ;
	input \core_c_dec_MFMR1_E_reg/P0001  ;
	input \core_c_dec_MFMR2_E_reg/P0001  ;
	input \core_c_dec_MFMSTAT_E_reg/P0001  ;
	input \core_c_dec_MFMX0_E_reg/P0001  ;
	input \core_c_dec_MFMX1_E_reg/P0001  ;
	input \core_c_dec_MFMY0_E_reg/P0001  ;
	input \core_c_dec_MFMY1_E_reg/P0001  ;
	input \core_c_dec_MFMreg_E_reg[0]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[1]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[2]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[3]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[4]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[5]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[6]/P0001  ;
	input \core_c_dec_MFMreg_E_reg[7]/P0001  ;
	input \core_c_dec_MFPMOVL_E_reg/P0001  ;
	input \core_c_dec_MFPSQ_Ei_reg/NET0131  ;
	input \core_c_dec_MFRX0_E_reg/P0001  ;
	input \core_c_dec_MFRX1_E_reg/P0001  ;
	input \core_c_dec_MFSB_E_reg/P0001  ;
	input \core_c_dec_MFSE_E_reg/P0001  ;
	input \core_c_dec_MFSHT_Ei_reg/NET0131  ;
	input \core_c_dec_MFSI_E_reg/P0001  ;
	input \core_c_dec_MFSPT_Ei_reg/NET0131  ;
	input \core_c_dec_MFSR0_E_reg/P0001  ;
	input \core_c_dec_MFSR1_E_reg/P0001  ;
	input \core_c_dec_MFSSTAT_E_reg/P0001  ;
	input \core_c_dec_MFTX0_E_reg/P0001  ;
	input \core_c_dec_MFTX1_E_reg/P0001  ;
	input \core_c_dec_MFtoppcs_Eg_reg/P0001  ;
	input \core_c_dec_MTAR_E_reg/P0001  ;
	input \core_c_dec_MTASTAT_E_reg/P0001  ;
	input \core_c_dec_MTAX0_E_reg/P0001  ;
	input \core_c_dec_MTAX1_E_reg/P0001  ;
	input \core_c_dec_MTAY0_E_reg/P0001  ;
	input \core_c_dec_MTAY1_E_reg/P0001  ;
	input \core_c_dec_MTCNTR_Eg_reg/P0001  ;
	input \core_c_dec_MTDMOVL_E_reg/P0001  ;
	input \core_c_dec_MTICNTL_Eg_reg/P0001  ;
	input \core_c_dec_MTIDR_E_reg/P0001  ;
	input \core_c_dec_MTIFC_Eg_reg/P0001  ;
	input \core_c_dec_MTIMASK_Eg_reg/P0001  ;
	input \core_c_dec_MTIreg_E_reg[0]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[1]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[2]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[3]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[4]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[5]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[6]/P0001  ;
	input \core_c_dec_MTIreg_E_reg[7]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[0]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[1]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[2]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[3]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[4]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[5]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[6]/P0001  ;
	input \core_c_dec_MTLreg_E_reg[7]/P0001  ;
	input \core_c_dec_MTMR0_E_reg/P0001  ;
	input \core_c_dec_MTMR1_E_reg/P0001  ;
	input \core_c_dec_MTMR2_E_reg/P0001  ;
	input \core_c_dec_MTMSTAT_Eg_reg/P0001  ;
	input \core_c_dec_MTMX0_E_reg/P0001  ;
	input \core_c_dec_MTMX1_E_reg/P0001  ;
	input \core_c_dec_MTMY0_E_reg/P0001  ;
	input \core_c_dec_MTMY1_E_reg/P0001  ;
	input \core_c_dec_MTMreg_E_reg[0]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[1]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[2]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[3]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[4]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[5]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[6]/P0001  ;
	input \core_c_dec_MTMreg_E_reg[7]/P0001  ;
	input \core_c_dec_MTOWRCNTR_Eg_reg/P0001  ;
	input \core_c_dec_MTPMOVL_E_reg/P0001  ;
	input \core_c_dec_MTRX0_E_reg/P0001  ;
	input \core_c_dec_MTRX1_E_reg/P0001  ;
	input \core_c_dec_MTSB_E_reg/P0001  ;
	input \core_c_dec_MTSE_E_reg/P0001  ;
	input \core_c_dec_MTSI_E_reg/P0001  ;
	input \core_c_dec_MTSR0_E_reg/P0001  ;
	input \core_c_dec_MTSR1_E_reg/P0001  ;
	input \core_c_dec_MTTX0_E_reg/P0001  ;
	input \core_c_dec_MTTX1_E_reg/P0001  ;
	input \core_c_dec_MTtoppcs_Eg_reg/P0001  ;
	input \core_c_dec_Modctl_Eg_reg/P0001  ;
	input \core_c_dec_MpopLP_Eg_reg/P0001  ;
	input \core_c_dec_NOP_E_reg/P0001  ;
	input \core_c_dec_Nrti_Ed_reg/P0001  ;
	input \core_c_dec_Nseq_Ed_reg/P0001  ;
	input \core_c_dec_PPclr_reg/P0001  ;
	input \core_c_dec_Post1_E_reg/P0001  ;
	input \core_c_dec_Post2_E_reg/P0001  ;
	input \core_c_dec_Prderr_Cg_reg/NET0131  ;
	input \core_c_dec_RET_Ed_reg/P0001  ;
	input \core_c_dec_RTI_Ed_reg/P0001  ;
	input \core_c_dec_SHTop_E_reg/P0001  ;
	input \core_c_dec_Stkctl_Eg_reg/P0001  ;
	input \core_c_dec_Usecond_E_reg/P0001  ;
	input \core_c_dec_accCM_E_reg/NET0131  ;
	input \core_c_dec_accPM_E_reg/P0001  ;
	input \core_c_dec_cdAM_E_reg/P0001  ;
	input \core_c_dec_imSHT_E_reg/P0001  ;
	input \core_c_dec_imm14_E_reg/P0001  ;
	input \core_c_dec_imm16_E_reg/P0001  ;
	input \core_c_dec_pMFALU_Ei_reg/NET0131  ;
	input \core_c_dec_pMFMAC_Ei_reg/NET0131  ;
	input \core_c_dec_pMFSHT_Ei_reg/NET0131  ;
	input \core_c_dec_rdCM_E_reg/NET0131  ;
	input \core_c_dec_satMR_E_reg/P0001  ;
	input \core_c_dec_updAF_E_reg/P0001  ;
	input \core_c_dec_updAR_E_reg/P0001  ;
	input \core_c_dec_updMF_E_reg/P0001  ;
	input \core_c_dec_updMR_E_reg/P0001  ;
	input \core_c_dec_updSR_E_reg/P0001  ;
	input \core_c_psq_CE_reg/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[0]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[10]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[11]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[12]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[13]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[1]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[2]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[3]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[4]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[5]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[6]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[7]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[8]/NET0131  ;
	input \core_c_psq_CNTR_reg_DO_reg[9]/NET0131  ;
	input \core_c_psq_CNTRval_reg/NET0131  ;
	input \core_c_psq_DMOVL_reg_DO_reg[0]/NET0131  ;
	input \core_c_psq_DMOVL_reg_DO_reg[1]/NET0131  ;
	input \core_c_psq_DMOVL_reg_DO_reg[2]/NET0131  ;
	input \core_c_psq_DMOVL_reg_DO_reg[3]/NET0131  ;
	input \core_c_psq_DRA_reg[0]/P0001  ;
	input \core_c_psq_DRA_reg[10]/P0001  ;
	input \core_c_psq_DRA_reg[11]/P0001  ;
	input \core_c_psq_DRA_reg[12]/P0001  ;
	input \core_c_psq_DRA_reg[13]/P0001  ;
	input \core_c_psq_DRA_reg[1]/P0001  ;
	input \core_c_psq_DRA_reg[2]/P0001  ;
	input \core_c_psq_DRA_reg[3]/P0001  ;
	input \core_c_psq_DRA_reg[4]/P0001  ;
	input \core_c_psq_DRA_reg[5]/P0001  ;
	input \core_c_psq_DRA_reg[6]/P0001  ;
	input \core_c_psq_DRA_reg[7]/P0001  ;
	input \core_c_psq_DRA_reg[8]/P0001  ;
	input \core_c_psq_DRA_reg[9]/P0001  ;
	input \core_c_psq_ECYC_reg/P0001  ;
	input \core_c_psq_EXA_reg[0]/P0001  ;
	input \core_c_psq_EXA_reg[10]/P0001  ;
	input \core_c_psq_EXA_reg[11]/P0001  ;
	input \core_c_psq_EXA_reg[12]/P0001  ;
	input \core_c_psq_EXA_reg[13]/P0001  ;
	input \core_c_psq_EXA_reg[1]/P0001  ;
	input \core_c_psq_EXA_reg[2]/P0001  ;
	input \core_c_psq_EXA_reg[3]/P0001  ;
	input \core_c_psq_EXA_reg[4]/P0001  ;
	input \core_c_psq_EXA_reg[5]/P0001  ;
	input \core_c_psq_EXA_reg[6]/P0001  ;
	input \core_c_psq_EXA_reg[7]/P0001  ;
	input \core_c_psq_EXA_reg[8]/P0001  ;
	input \core_c_psq_EXA_reg[9]/P0001  ;
	input \core_c_psq_Eqend_D_reg/P0001  ;
	input \core_c_psq_Eqend_Ed_reg/P0001  ;
	input \core_c_psq_ICNTL_reg_DO_reg[0]/NET0131  ;
	input \core_c_psq_ICNTL_reg_DO_reg[1]/NET0131  ;
	input \core_c_psq_ICNTL_reg_DO_reg[2]/NET0131  ;
	input \core_c_psq_ICNTL_reg_DO_reg[4]/NET0131  ;
	input \core_c_psq_IFA_reg[0]/P0001  ;
	input \core_c_psq_IFA_reg[10]/P0001  ;
	input \core_c_psq_IFA_reg[11]/P0001  ;
	input \core_c_psq_IFA_reg[12]/P0001  ;
	input \core_c_psq_IFA_reg[13]/P0001  ;
	input \core_c_psq_IFA_reg[1]/P0001  ;
	input \core_c_psq_IFA_reg[2]/P0001  ;
	input \core_c_psq_IFA_reg[3]/P0001  ;
	input \core_c_psq_IFA_reg[4]/P0001  ;
	input \core_c_psq_IFA_reg[5]/P0001  ;
	input \core_c_psq_IFA_reg[6]/P0001  ;
	input \core_c_psq_IFA_reg[7]/P0001  ;
	input \core_c_psq_IFA_reg[8]/P0001  ;
	input \core_c_psq_IFA_reg[9]/P0001  ;
	input \core_c_psq_IFC_reg[0]/NET0131  ;
	input \core_c_psq_IFC_reg[10]/NET0131  ;
	input \core_c_psq_IFC_reg[11]/NET0131  ;
	input \core_c_psq_IFC_reg[12]/NET0131  ;
	input \core_c_psq_IFC_reg[13]/NET0131  ;
	input \core_c_psq_IFC_reg[14]/NET0131  ;
	input \core_c_psq_IFC_reg[15]/NET0131  ;
	input \core_c_psq_IFC_reg[1]/NET0131  ;
	input \core_c_psq_IFC_reg[2]/NET0131  ;
	input \core_c_psq_IFC_reg[3]/NET0131  ;
	input \core_c_psq_IFC_reg[4]/NET0131  ;
	input \core_c_psq_IFC_reg[5]/NET0131  ;
	input \core_c_psq_IFC_reg[6]/NET0131  ;
	input \core_c_psq_IFC_reg[7]/NET0131  ;
	input \core_c_psq_IFC_reg[8]/NET0131  ;
	input \core_c_psq_IFC_reg[9]/NET0131  ;
	input \core_c_psq_IMASK_reg[0]/NET0131  ;
	input \core_c_psq_IMASK_reg[1]/NET0131  ;
	input \core_c_psq_IMASK_reg[2]/NET0131  ;
	input \core_c_psq_IMASK_reg[3]/NET0131  ;
	input \core_c_psq_IMASK_reg[4]/NET0131  ;
	input \core_c_psq_IMASK_reg[5]/NET0131  ;
	input \core_c_psq_IMASK_reg[6]/NET0131  ;
	input \core_c_psq_IMASK_reg[7]/NET0131  ;
	input \core_c_psq_IMASK_reg[8]/NET0131  ;
	input \core_c_psq_IMASK_reg[9]/NET0131  ;
	input \core_c_psq_INT_en_reg/NET0131  ;
	input \core_c_psq_Iact_E_reg[0]/NET0131  ;
	input \core_c_psq_Iact_E_reg[10]/NET0131  ;
	input \core_c_psq_Iact_E_reg[1]/NET0131  ;
	input \core_c_psq_Iact_E_reg[2]/NET0131  ;
	input \core_c_psq_Iact_E_reg[3]/NET0131  ;
	input \core_c_psq_Iact_E_reg[4]/NET0131  ;
	input \core_c_psq_Iact_E_reg[5]/NET0131  ;
	input \core_c_psq_Iact_E_reg[6]/NET0131  ;
	input \core_c_psq_Iact_E_reg[7]/NET0131  ;
	input \core_c_psq_Iact_E_reg[8]/NET0131  ;
	input \core_c_psq_Iact_E_reg[9]/NET0131  ;
	input \core_c_psq_Iflag_reg[0]/NET0131  ;
	input \core_c_psq_Iflag_reg[10]/NET0131  ;
	input \core_c_psq_Iflag_reg[11]/NET0131  ;
	input \core_c_psq_Iflag_reg[12]/NET0131  ;
	input \core_c_psq_Iflag_reg[1]/NET0131  ;
	input \core_c_psq_Iflag_reg[2]/NET0131  ;
	input \core_c_psq_Iflag_reg[3]/NET0131  ;
	input \core_c_psq_Iflag_reg[4]/NET0131  ;
	input \core_c_psq_Iflag_reg[5]/NET0131  ;
	input \core_c_psq_Iflag_reg[6]/NET0131  ;
	input \core_c_psq_Iflag_reg[7]/NET0131  ;
	input \core_c_psq_Iflag_reg[8]/NET0131  ;
	input \core_c_psq_Iflag_reg[9]/NET0131  ;
	input \core_c_psq_MGNT_reg/NET0131  ;
	input \core_c_psq_MREQ_reg/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[0]/P0002  ;
	input \core_c_psq_MSTAT_reg_DO_reg[1]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[2]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[3]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[4]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[5]/NET0131  ;
	input \core_c_psq_MSTAT_reg_DO_reg[6]/NET0131  ;
	input \core_c_psq_PCS2or3_reg/NET0131  ;
	input \core_c_psq_PCS_reg[0]/NET0131  ;
	input \core_c_psq_PCS_reg[10]/NET0131  ;
	input \core_c_psq_PCS_reg[11]/NET0131  ;
	input \core_c_psq_PCS_reg[12]/NET0131  ;
	input \core_c_psq_PCS_reg[13]/NET0131  ;
	input \core_c_psq_PCS_reg[14]/NET0131  ;
	input \core_c_psq_PCS_reg[15]/NET0131  ;
	input \core_c_psq_PCS_reg[1]/NET0131  ;
	input \core_c_psq_PCS_reg[2]/NET0131  ;
	input \core_c_psq_PCS_reg[3]/NET0131  ;
	input \core_c_psq_PCS_reg[4]/NET0131  ;
	input \core_c_psq_PCS_reg[5]/NET0131  ;
	input \core_c_psq_PCS_reg[6]/NET0131  ;
	input \core_c_psq_PCS_reg[7]/NET0131  ;
	input \core_c_psq_PCS_reg[8]/NET0131  ;
	input \core_c_psq_PMOVL_regh_DO_reg[0]/NET0131  ;
	input \core_c_psq_PMOVL_regh_DO_reg[1]/NET0131  ;
	input \core_c_psq_PMOVL_regh_DO_reg[2]/NET0131  ;
	input \core_c_psq_PMOVL_regh_DO_reg[3]/NET0131  ;
	input \core_c_psq_PMOVL_regl_DO_reg[0]/NET0131  ;
	input \core_c_psq_PMOVL_regl_DO_reg[1]/NET0131  ;
	input \core_c_psq_PMOVL_regl_DO_reg[2]/NET0131  ;
	input \core_c_psq_PMOVL_regl_DO_reg[3]/NET0131  ;
	input \core_c_psq_SRST_reg/P0001  ;
	input \core_c_psq_SSTAT_reg[0]/NET0131  ;
	input \core_c_psq_SSTAT_reg[1]/NET0131  ;
	input \core_c_psq_SSTAT_reg[2]/NET0131  ;
	input \core_c_psq_SSTAT_reg[3]/NET0131  ;
	input \core_c_psq_SSTAT_reg[4]/NET0131  ;
	input \core_c_psq_SSTAT_reg[5]/NET0131  ;
	input \core_c_psq_SSTAT_reg[6]/NET0131  ;
	input \core_c_psq_SSTAT_reg[7]/NET0131  ;
	input \core_c_psq_TRAP_Eg_reg/NET0131  ;
	input \core_c_psq_TRAP_R_L_reg/NET0131  ;
	input \core_c_psq_T_IRQ0_s1_reg/P0001  ;
	input \core_c_psq_T_IRQ0p_reg/P0001  ;
	input \core_c_psq_T_IRQ1_s1_reg/P0001  ;
	input \core_c_psq_T_IRQ1p_reg/P0001  ;
	input \core_c_psq_T_IRQ2_s1_reg/P0001  ;
	input \core_c_psq_T_IRQ2p_reg/P0001  ;
	input \core_c_psq_T_IRQE0_reg/P0001  ;
	input \core_c_psq_T_IRQE0_s1_reg/P0001  ;
	input \core_c_psq_T_IRQE1_reg/P0001  ;
	input \core_c_psq_T_IRQE1_s1_reg/P0001  ;
	input \core_c_psq_T_IRQL0p_reg/P0001  ;
	input \core_c_psq_T_IRQL1p_reg/P0001  ;
	input \core_c_psq_T_PWRDN_reg/P0001  ;
	input \core_c_psq_T_PWRDN_s1_reg/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[0]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[10]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[11]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[12]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[13]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[1]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[2]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[3]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[4]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[5]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[6]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[7]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[8]/P0001  ;
	input \core_c_psq_Taddr_Eb_reg[9]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001  ;
	input \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001  ;
	input \core_c_psq_cntstk_ptr_reg[0]/NET0131  ;
	input \core_c_psq_cntstk_ptr_reg[1]/NET0131  ;
	input \core_c_psq_cntstk_ptr_reg[2]/NET0131  ;
	input \core_c_psq_irq0_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irq0_de_OUT_reg/P0001  ;
	input \core_c_psq_irq1_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irq1_de_OUT_reg/P0001  ;
	input \core_c_psq_irq2_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irq2_de_OUT_reg/P0001  ;
	input \core_c_psq_irql0_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irql0_de_OUT_reg/P0001  ;
	input \core_c_psq_irql1_de_IN_syn_reg/P0001  ;
	input \core_c_psq_irql1_de_OUT_reg/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001  ;
	input \core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001  ;
	input \core_c_psq_lpstk_ptr_reg[0]/NET0131  ;
	input \core_c_psq_lpstk_ptr_reg[1]/NET0131  ;
	input \core_c_psq_lpstk_ptr_reg[2]/NET0131  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001  ;
	input \core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001  ;
	input \core_c_psq_pcstk_ptr_reg[0]/NET0131  ;
	input \core_c_psq_pcstk_ptr_reg[1]/NET0131  ;
	input \core_c_psq_pcstk_ptr_reg[2]/NET0131  ;
	input \core_c_psq_pcstk_ptr_reg[3]/NET0131  ;
	input \core_c_psq_pcstk_ptr_reg[4]/NET0131  ;
	input \core_c_psq_ststk_ptr_reg[0]/NET0131  ;
	input \core_c_psq_ststk_ptr_reg[1]/NET0131  ;
	input \core_c_psq_ststk_ptr_reg[2]/NET0131  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001  ;
	input \core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_I_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_L_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_M_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131  ;
	input \core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131  ;
	input \core_dag_ilm1reg_STEALI_E_reg[0]/P0001  ;
	input \core_dag_ilm1reg_STEALI_E_reg[1]/P0001  ;
	input \core_dag_ilm1reg_STEALI_E_reg[2]/P0001  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_IL_E_reg[0]/P0001  ;
	input \core_dag_ilm2reg_IL_E_reg[1]/P0001  ;
	input \core_dag_ilm2reg_I_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_I_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_L_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_M_E_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M_E_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_M_reg[9]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131  ;
	input \core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131  ;
	input \core_dag_modulo1_R0wrap_reg/P0001  ;
	input \core_dag_modulo1_R1wrap_reg/P0001  ;
	input \core_dag_modulo1_T0wrap_reg/P0001  ;
	input \core_dag_modulo1_T1wrap_reg/P0001  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001  ;
	input \core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001  ;
	input \core_eu_ec_cun_AC_reg/P0001  ;
	input \core_eu_ec_cun_AN_reg/P0001  ;
	input \core_eu_ec_cun_AQ_reg/P0001  ;
	input \core_eu_ec_cun_AS_reg/P0001  ;
	input \core_eu_ec_cun_AV_reg/P0001  ;
	input \core_eu_ec_cun_AZ_reg/P0001  ;
	input \core_eu_ec_cun_COND_E_reg[0]/P0001  ;
	input \core_eu_ec_cun_COND_E_reg[1]/P0001  ;
	input \core_eu_ec_cun_COND_E_reg[2]/P0001  ;
	input \core_eu_ec_cun_COND_E_reg[3]/P0001  ;
	input \core_eu_ec_cun_MV_reg/P0000_reg_syn_2  ;
	input \core_eu_ec_cun_MVi_pre_C_reg/P0001  ;
	input \core_eu_ec_cun_SS_reg/P0001  ;
	input \core_eu_ec_cun_TERM_E_reg[0]/P0001  ;
	input \core_eu_ec_cun_TERM_E_reg[1]/P0001  ;
	input \core_eu_ec_cun_TERM_E_reg[2]/P0001  ;
	input \core_eu_ec_cun_TERM_E_reg[3]/P0001  ;
	input \core_eu_ec_cun_condOK_CE_reg/P0001  ;
	input \core_eu_ec_cun_mven_FFout_reg/NET0131  ;
	input \core_eu_ec_cun_termOK_CE_reg/P0001  ;
	input \core_eu_ec_cun_updateMV_C_reg/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_Sq_E_reg/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001  ;
	input \core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001  ;
	input \core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2  ;
	input \core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2  ;
	input \core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2  ;
	input \core_eu_es_sht_es_reg_SBr_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_SBr_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_SBr_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_SBr_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_SBr_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_SBs_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001  ;
	input \core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001  ;
	input \emc_DMDoe_reg/NET0131  ;
	input \emc_DMDreg_reg[0]/P0001  ;
	input \emc_DMDreg_reg[10]/P0001  ;
	input \emc_DMDreg_reg[11]/P0001  ;
	input \emc_DMDreg_reg[12]/P0001  ;
	input \emc_DMDreg_reg[13]/P0001  ;
	input \emc_DMDreg_reg[14]/P0001  ;
	input \emc_DMDreg_reg[15]/P0001  ;
	input \emc_DMDreg_reg[1]/P0001  ;
	input \emc_DMDreg_reg[2]/P0001  ;
	input \emc_DMDreg_reg[3]/P0001  ;
	input \emc_DMDreg_reg[4]/P0001  ;
	input \emc_DMDreg_reg[5]/P0001  ;
	input \emc_DMDreg_reg[6]/P0001  ;
	input \emc_DMDreg_reg[7]/P0001  ;
	input \emc_DMDreg_reg[8]/P0001  ;
	input \emc_DMDreg_reg[9]/P0001  ;
	input \emc_DMcst_reg/NET0131  ;
	input \emc_ECMA_reg[0]/P0001  ;
	input \emc_ECMA_reg[10]/P0001  ;
	input \emc_ECMA_reg[11]/P0001  ;
	input \emc_ECMA_reg[12]/P0001  ;
	input \emc_ECMA_reg[1]/P0001  ;
	input \emc_ECMA_reg[2]/P0001  ;
	input \emc_ECMA_reg[3]/P0001  ;
	input \emc_ECMA_reg[4]/P0001  ;
	input \emc_ECMA_reg[5]/P0001  ;
	input \emc_ECMA_reg[6]/P0001  ;
	input \emc_ECMA_reg[7]/P0001  ;
	input \emc_ECMA_reg[8]/P0001  ;
	input \emc_ECMA_reg[9]/P0001  ;
	input \emc_ECMDreg_reg[0]/P0001  ;
	input \emc_ECMDreg_reg[10]/P0001  ;
	input \emc_ECMDreg_reg[11]/P0001  ;
	input \emc_ECMDreg_reg[12]/P0001  ;
	input \emc_ECMDreg_reg[13]/P0001  ;
	input \emc_ECMDreg_reg[14]/P0001  ;
	input \emc_ECMDreg_reg[15]/P0001  ;
	input \emc_ECMDreg_reg[16]/P0001  ;
	input \emc_ECMDreg_reg[17]/P0001  ;
	input \emc_ECMDreg_reg[18]/P0001  ;
	input \emc_ECMDreg_reg[19]/P0001  ;
	input \emc_ECMDreg_reg[1]/P0001  ;
	input \emc_ECMDreg_reg[20]/P0001  ;
	input \emc_ECMDreg_reg[21]/P0001  ;
	input \emc_ECMDreg_reg[22]/P0001  ;
	input \emc_ECMDreg_reg[23]/P0001  ;
	input \emc_ECMDreg_reg[2]/P0001  ;
	input \emc_ECMDreg_reg[3]/P0001  ;
	input \emc_ECMDreg_reg[4]/P0001  ;
	input \emc_ECMDreg_reg[5]/P0001  ;
	input \emc_ECMDreg_reg[6]/P0001  ;
	input \emc_ECMDreg_reg[7]/P0001  ;
	input \emc_ECMDreg_reg[8]/P0001  ;
	input \emc_ECMDreg_reg[9]/P0001  ;
	input \emc_ECMcs_reg/NET0131  ;
	input \emc_ECS_reg[0]/NET0131  ;
	input \emc_ECS_reg[1]/NET0131  ;
	input \emc_ECS_reg[2]/NET0131  ;
	input \emc_ECS_reg[3]/NET0131  ;
	input \emc_ED_oei_reg/P0001  ;
	input \emc_EXTC_Eg_syn_reg/P0001  ;
	input \emc_IOcst_reg/NET0131  ;
	input \emc_PMDoe_reg/NET0131  ;
	input \emc_PMDreg_reg[0]/P0001  ;
	input \emc_PMDreg_reg[10]/P0001  ;
	input \emc_PMDreg_reg[11]/P0001  ;
	input \emc_PMDreg_reg[12]/P0001  ;
	input \emc_PMDreg_reg[13]/P0001  ;
	input \emc_PMDreg_reg[14]/P0001  ;
	input \emc_PMDreg_reg[15]/P0001  ;
	input \emc_PMDreg_reg[1]/P0001  ;
	input \emc_PMDreg_reg[2]/P0001  ;
	input \emc_PMDreg_reg[3]/P0001  ;
	input \emc_PMDreg_reg[4]/P0001  ;
	input \emc_PMDreg_reg[5]/P0001  ;
	input \emc_PMDreg_reg[6]/P0001  ;
	input \emc_PMDreg_reg[7]/P0001  ;
	input \emc_PMDreg_reg[8]/P0001  ;
	input \emc_PMDreg_reg[9]/P0001  ;
	input \emc_PMcst_reg/NET0131  ;
	input \emc_RWcnt_reg[0]/P0001  ;
	input \emc_RWcnt_reg[1]/P0001  ;
	input \emc_RWcnt_reg[2]/P0001  ;
	input \emc_RWcnt_reg[3]/P0001  ;
	input \emc_RWcnt_reg[4]/P0001  ;
	input \emc_RWcnt_reg[5]/P0001  ;
	input \emc_WRn_h_reg/P0001  ;
	input \emc_WSCRext_reg_DO_reg[0]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[1]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[2]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[3]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[4]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[5]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[6]/NET0131  ;
	input \emc_WSCRext_reg_DO_reg[7]/NET0131  ;
	input \emc_WSCRreg_DO_reg[0]/NET0131  ;
	input \emc_WSCRreg_DO_reg[10]/NET0131  ;
	input \emc_WSCRreg_DO_reg[11]/NET0131  ;
	input \emc_WSCRreg_DO_reg[12]/NET0131  ;
	input \emc_WSCRreg_DO_reg[13]/NET0131  ;
	input \emc_WSCRreg_DO_reg[14]/NET0131  ;
	input \emc_WSCRreg_DO_reg[1]/NET0131  ;
	input \emc_WSCRreg_DO_reg[2]/NET0131  ;
	input \emc_WSCRreg_DO_reg[3]/NET0131  ;
	input \emc_WSCRreg_DO_reg[4]/NET0131  ;
	input \emc_WSCRreg_DO_reg[5]/NET0131  ;
	input \emc_WSCRreg_DO_reg[6]/NET0131  ;
	input \emc_WSCRreg_DO_reg[7]/NET0131  ;
	input \emc_WSCRreg_DO_reg[8]/NET0131  ;
	input \emc_WSCRreg_DO_reg[9]/NET0131  ;
	input \emc_eRDY_reg/NET0131  ;
	input \emc_selDMDi_reg/P0001  ;
	input \emc_selPMDi_reg/P0001  ;
	input \idma_CM_oe_reg/P0001  ;
	input \idma_CMo_oe0_reg/P0001  ;
	input \idma_CMo_oe1_reg/P0001  ;
	input \idma_CMo_oe2_reg/P0001  ;
	input \idma_CMo_oe3_reg/P0001  ;
	input \idma_CMo_oe4_reg/P0001  ;
	input \idma_CMo_oe5_reg/P0001  ;
	input \idma_CMo_oe6_reg/P0001  ;
	input \idma_CMo_oe7_reg/P0001  ;
	input \idma_DCTL_reg[0]/NET0131  ;
	input \idma_DCTL_reg[10]/NET0131  ;
	input \idma_DCTL_reg[11]/NET0131  ;
	input \idma_DCTL_reg[12]/NET0131  ;
	input \idma_DCTL_reg[13]/NET0131  ;
	input \idma_DCTL_reg[14]/NET0131  ;
	input \idma_DCTL_reg[1]/NET0131  ;
	input \idma_DCTL_reg[2]/NET0131  ;
	input \idma_DCTL_reg[3]/NET0131  ;
	input \idma_DCTL_reg[4]/NET0131  ;
	input \idma_DCTL_reg[5]/NET0131  ;
	input \idma_DCTL_reg[6]/NET0131  ;
	input \idma_DCTL_reg[7]/NET0131  ;
	input \idma_DCTL_reg[8]/NET0131  ;
	input \idma_DCTL_reg[9]/NET0131  ;
	input \idma_DOVL_reg[0]/NET0131  ;
	input \idma_DOVL_reg[10]/NET0131  ;
	input \idma_DOVL_reg[11]/NET0131  ;
	input \idma_DOVL_reg[1]/NET0131  ;
	input \idma_DOVL_reg[2]/NET0131  ;
	input \idma_DOVL_reg[3]/NET0131  ;
	input \idma_DOVL_reg[4]/NET0131  ;
	input \idma_DOVL_reg[5]/NET0131  ;
	input \idma_DOVL_reg[6]/NET0131  ;
	input \idma_DOVL_reg[7]/NET0131  ;
	input \idma_DOVL_reg[8]/NET0131  ;
	input \idma_DOVL_reg[9]/NET0131  ;
	input \idma_DSreq_reg/NET0131  ;
	input \idma_DTMP_H_reg[0]/P0001  ;
	input \idma_DTMP_H_reg[10]/P0001  ;
	input \idma_DTMP_H_reg[11]/P0001  ;
	input \idma_DTMP_H_reg[12]/P0001  ;
	input \idma_DTMP_H_reg[13]/P0001  ;
	input \idma_DTMP_H_reg[14]/P0001  ;
	input \idma_DTMP_H_reg[15]/P0001  ;
	input \idma_DTMP_H_reg[1]/P0001  ;
	input \idma_DTMP_H_reg[2]/P0001  ;
	input \idma_DTMP_H_reg[3]/P0001  ;
	input \idma_DTMP_H_reg[4]/P0001  ;
	input \idma_DTMP_H_reg[5]/P0001  ;
	input \idma_DTMP_H_reg[6]/P0001  ;
	input \idma_DTMP_H_reg[7]/P0001  ;
	input \idma_DTMP_H_reg[8]/P0001  ;
	input \idma_DTMP_H_reg[9]/P0001  ;
	input \idma_DTMP_L_reg[0]/P0001  ;
	input \idma_DTMP_L_reg[1]/P0001  ;
	input \idma_DTMP_L_reg[2]/P0001  ;
	input \idma_DTMP_L_reg[3]/P0001  ;
	input \idma_DTMP_L_reg[4]/P0001  ;
	input \idma_DTMP_L_reg[5]/P0001  ;
	input \idma_DTMP_L_reg[6]/P0001  ;
	input \idma_DTMP_L_reg[7]/P0001  ;
	input \idma_IADi_reg[0]/P0001  ;
	input \idma_IADi_reg[10]/P0001  ;
	input \idma_IADi_reg[11]/P0001  ;
	input \idma_IADi_reg[12]/P0001  ;
	input \idma_IADi_reg[13]/P0001  ;
	input \idma_IADi_reg[14]/P0001  ;
	input \idma_IADi_reg[15]/P0001  ;
	input \idma_IADi_reg[1]/P0001  ;
	input \idma_IADi_reg[2]/P0001  ;
	input \idma_IADi_reg[3]/P0001  ;
	input \idma_IADi_reg[4]/P0001  ;
	input \idma_IADi_reg[5]/P0001  ;
	input \idma_IADi_reg[6]/P0001  ;
	input \idma_IADi_reg[7]/P0001  ;
	input \idma_IADi_reg[8]/P0001  ;
	input \idma_IADi_reg[9]/P0001  ;
	input \idma_IAL_reg/P0001  ;
	input \idma_IDMA_boot_reg/NET0131_reg_syn_10  ;
	input \idma_IDMA_boot_reg/NET0131_reg_syn_2  ;
	input \idma_IDMA_boot_reg/NET0131_reg_syn_8  ;
	input \idma_IRDn_reg/P0001  ;
	input \idma_ISn_reg/P0001  ;
	input \idma_IWRn_reg/P0001  ;
	input \idma_PCrd_1st_reg/NET0131  ;
	input \idma_PM_1st_reg/NET0131  ;
	input \idma_RDCMD_d1_reg/P0001  ;
	input \idma_RDCMD_reg/P0001  ;
	input \idma_RDcnt_reg[0]/NET0131  ;
	input \idma_RDcnt_reg[1]/NET0131  ;
	input \idma_RDcnt_reg[2]/NET0131  ;
	input \idma_RDcyc_reg/NET0131  ;
	input \idma_WRCMD_d1_reg/P0001  ;
	input \idma_WRCMD_reg/P0001  ;
	input \idma_WRcnt_reg[0]/NET0131  ;
	input \idma_WRcnt_reg[1]/NET0131  ;
	input \idma_WRcnt_reg[2]/NET0131  ;
	input \idma_WRcyc_reg/NET0131  ;
	input \idma_WRtrue_reg/NET0131  ;
	input \memc_DM_oe_reg/P0001  ;
	input \memc_DMo_oe0_reg/P0001  ;
	input \memc_DMo_oe1_reg/P0001  ;
	input \memc_DMo_oe2_reg/P0001  ;
	input \memc_DMo_oe3_reg/P0001  ;
	input \memc_DMo_oe4_reg/P0001  ;
	input \memc_DMo_oe5_reg/P0001  ;
	input \memc_DMo_oe6_reg/P0001  ;
	input \memc_DMo_oe7_reg/P0001  ;
	input \memc_Dread_E_reg/NET0131  ;
	input \memc_Dwrite_C_reg/NET0131  ;
	input \memc_Dwrite_E_reg/NET0131  ;
	input \memc_EXTC_E_reg/NET0131  ;
	input \memc_EXTC_Eg_reg/NET0131_reg_syn_10  ;
	input \memc_EXTC_Eg_reg/NET0131_reg_syn_2  ;
	input \memc_EXTC_Eg_reg/NET0131_reg_syn_8  ;
	input \memc_IOcmd_E_reg/NET0131  ;
	input \memc_LDaST_Eg_reg/NET0131  ;
	input \memc_MMR_web_reg/NET0131  ;
	input \memc_PMo_oe0_reg/P0001  ;
	input \memc_PMo_oe1_reg/P0001  ;
	input \memc_PMo_oe2_reg/P0001  ;
	input \memc_PMo_oe3_reg/P0001  ;
	input \memc_PMo_oe4_reg/P0001  ;
	input \memc_PMo_oe5_reg/P0001  ;
	input \memc_PMo_oe6_reg/P0001  ;
	input \memc_PMo_oe7_reg/P0001  ;
	input \memc_Pread_E_reg/NET0131  ;
	input \memc_Pwrite_C_reg/NET0131  ;
	input \memc_Pwrite_E_reg/NET0131  ;
	input \memc_STI_Cg_reg/NET0131  ;
	input \memc_accDM_E_reg/NET0131  ;
	input \memc_accPM_E_reg/NET0131  ;
	input \memc_ldSREG_E_reg/NET0131  ;
	input \memc_selMIO_E_reg/P0001  ;
	input \memc_usysr_DO_reg[0]/NET0131  ;
	input \memc_usysr_DO_reg[10]/NET0131  ;
	input \memc_usysr_DO_reg[11]/NET0131  ;
	input \memc_usysr_DO_reg[12]/NET0131  ;
	input \memc_usysr_DO_reg[13]/NET0131  ;
	input \memc_usysr_DO_reg[14]/NET0131  ;
	input \memc_usysr_DO_reg[15]/NET0131  ;
	input \memc_usysr_DO_reg[1]/NET0131  ;
	input \memc_usysr_DO_reg[2]/NET0131  ;
	input \memc_usysr_DO_reg[3]/NET0131  ;
	input \memc_usysr_DO_reg[4]/NET0131  ;
	input \memc_usysr_DO_reg[5]/NET0131  ;
	input \memc_usysr_DO_reg[6]/NET0131  ;
	input \memc_usysr_DO_reg[7]/NET0131  ;
	input \memc_usysr_DO_reg[8]/NET0131  ;
	input \memc_usysr_DO_reg[9]/NET0131  ;
	input \pio_PINT_reg[0]/NET0131  ;
	input \pio_PINT_reg[10]/NET0131  ;
	input \pio_PINT_reg[11]/NET0131  ;
	input \pio_PINT_reg[1]/NET0131  ;
	input \pio_PINT_reg[2]/NET0131  ;
	input \pio_PINT_reg[3]/NET0131  ;
	input \pio_PINT_reg[4]/NET0131  ;
	input \pio_PINT_reg[5]/NET0131  ;
	input \pio_PINT_reg[6]/NET0131  ;
	input \pio_PINT_reg[7]/NET0131  ;
	input \pio_PINT_reg[8]/NET0131  ;
	input \pio_PINT_reg[9]/NET0131  ;
	input \pio_PIO_IN_P_reg[0]/P0001  ;
	input \pio_PIO_IN_P_reg[10]/P0001  ;
	input \pio_PIO_IN_P_reg[11]/P0001  ;
	input \pio_PIO_IN_P_reg[1]/P0001  ;
	input \pio_PIO_IN_P_reg[2]/P0001  ;
	input \pio_PIO_IN_P_reg[3]/P0001  ;
	input \pio_PIO_IN_P_reg[4]/P0001  ;
	input \pio_PIO_IN_P_reg[5]/P0001  ;
	input \pio_PIO_IN_P_reg[6]/P0001  ;
	input \pio_PIO_IN_P_reg[7]/P0001  ;
	input \pio_PIO_IN_P_reg[8]/P0001  ;
	input \pio_PIO_IN_P_reg[9]/P0001  ;
	input \pio_PIO_RES_OUT_reg[0]/P0001  ;
	input \pio_PIO_RES_OUT_reg[10]/P0001  ;
	input \pio_PIO_RES_OUT_reg[11]/P0001  ;
	input \pio_PIO_RES_OUT_reg[1]/P0001  ;
	input \pio_PIO_RES_OUT_reg[2]/P0001  ;
	input \pio_PIO_RES_OUT_reg[3]/P0001  ;
	input \pio_PIO_RES_OUT_reg[4]/P0001  ;
	input \pio_PIO_RES_OUT_reg[5]/P0001  ;
	input \pio_PIO_RES_OUT_reg[6]/P0001  ;
	input \pio_PIO_RES_OUT_reg[7]/P0001  ;
	input \pio_PIO_RES_OUT_reg[8]/P0001  ;
	input \pio_PIO_RES_OUT_reg[9]/P0001  ;
	input \pio_PIO_RES_reg[0]/NET0131  ;
	input \pio_PIO_RES_reg[10]/NET0131  ;
	input \pio_PIO_RES_reg[11]/NET0131  ;
	input \pio_PIO_RES_reg[1]/NET0131  ;
	input \pio_PIO_RES_reg[2]/NET0131  ;
	input \pio_PIO_RES_reg[3]/NET0131  ;
	input \pio_PIO_RES_reg[4]/NET0131  ;
	input \pio_PIO_RES_reg[5]/NET0131  ;
	input \pio_PIO_RES_reg[6]/NET0131  ;
	input \pio_PIO_RES_reg[7]/NET0131  ;
	input \pio_PIO_RES_reg[8]/NET0131  ;
	input \pio_PIO_RES_reg[9]/NET0131  ;
	input \pio_pmask_reg_DO_reg[0]/NET0131  ;
	input \pio_pmask_reg_DO_reg[10]/NET0131  ;
	input \pio_pmask_reg_DO_reg[11]/NET0131  ;
	input \pio_pmask_reg_DO_reg[1]/NET0131  ;
	input \pio_pmask_reg_DO_reg[2]/NET0131  ;
	input \pio_pmask_reg_DO_reg[3]/NET0131  ;
	input \pio_pmask_reg_DO_reg[4]/NET0131  ;
	input \pio_pmask_reg_DO_reg[5]/NET0131  ;
	input \pio_pmask_reg_DO_reg[6]/NET0131  ;
	input \pio_pmask_reg_DO_reg[7]/NET0131  ;
	input \pio_pmask_reg_DO_reg[8]/NET0131  ;
	input \pio_pmask_reg_DO_reg[9]/NET0131  ;
	input \regout_STD_C_reg[0]/P0001  ;
	input \regout_STD_C_reg[10]/P0001  ;
	input \regout_STD_C_reg[11]/P0001  ;
	input \regout_STD_C_reg[12]/P0001  ;
	input \regout_STD_C_reg[13]/P0001  ;
	input \regout_STD_C_reg[14]/P0001  ;
	input \regout_STD_C_reg[15]/P0001  ;
	input \regout_STD_C_reg[1]/P0001  ;
	input \regout_STD_C_reg[2]/P0001  ;
	input \regout_STD_C_reg[3]/P0001  ;
	input \regout_STD_C_reg[4]/P0001  ;
	input \regout_STD_C_reg[5]/P0001  ;
	input \regout_STD_C_reg[6]/P0001  ;
	input \regout_STD_C_reg[7]/P0001  ;
	input \regout_STD_C_reg[8]/P0001  ;
	input \regout_STD_C_reg[9]/P0001  ;
	input \sice_CLR_I_reg/NET0131  ;
	input \sice_CLR_M_reg/NET0131  ;
	input \sice_CMRW_reg/NET0131  ;
	input \sice_DBR1_reg[0]/P0001  ;
	input \sice_DBR1_reg[10]/P0001  ;
	input \sice_DBR1_reg[11]/P0001  ;
	input \sice_DBR1_reg[12]/P0001  ;
	input \sice_DBR1_reg[13]/P0001  ;
	input \sice_DBR1_reg[14]/P0001  ;
	input \sice_DBR1_reg[15]/P0001  ;
	input \sice_DBR1_reg[16]/P0001  ;
	input \sice_DBR1_reg[17]/P0001  ;
	input \sice_DBR1_reg[18]/P0001  ;
	input \sice_DBR1_reg[1]/P0001  ;
	input \sice_DBR1_reg[2]/P0001  ;
	input \sice_DBR1_reg[3]/P0001  ;
	input \sice_DBR1_reg[4]/P0001  ;
	input \sice_DBR1_reg[5]/P0001  ;
	input \sice_DBR1_reg[6]/P0001  ;
	input \sice_DBR1_reg[7]/P0001  ;
	input \sice_DBR1_reg[8]/P0001  ;
	input \sice_DBR1_reg[9]/P0001  ;
	input \sice_DBR2_reg[0]/P0001  ;
	input \sice_DBR2_reg[10]/P0001  ;
	input \sice_DBR2_reg[11]/P0001  ;
	input \sice_DBR2_reg[12]/P0001  ;
	input \sice_DBR2_reg[13]/P0001  ;
	input \sice_DBR2_reg[14]/P0001  ;
	input \sice_DBR2_reg[15]/P0001  ;
	input \sice_DBR2_reg[16]/P0001  ;
	input \sice_DBR2_reg[17]/P0001  ;
	input \sice_DBR2_reg[18]/P0001  ;
	input \sice_DBR2_reg[1]/P0001  ;
	input \sice_DBR2_reg[2]/P0001  ;
	input \sice_DBR2_reg[3]/P0001  ;
	input \sice_DBR2_reg[4]/P0001  ;
	input \sice_DBR2_reg[5]/P0001  ;
	input \sice_DBR2_reg[6]/P0001  ;
	input \sice_DBR2_reg[7]/P0001  ;
	input \sice_DBR2_reg[8]/P0001  ;
	input \sice_DBR2_reg[9]/P0001  ;
	input \sice_DMR1_reg[0]/NET0131  ;
	input \sice_DMR1_reg[10]/NET0131  ;
	input \sice_DMR1_reg[11]/NET0131  ;
	input \sice_DMR1_reg[12]/NET0131  ;
	input \sice_DMR1_reg[13]/NET0131  ;
	input \sice_DMR1_reg[14]/NET0131  ;
	input \sice_DMR1_reg[15]/NET0131  ;
	input \sice_DMR1_reg[16]/NET0131  ;
	input \sice_DMR1_reg[17]/NET0131  ;
	input \sice_DMR1_reg[1]/NET0131  ;
	input \sice_DMR1_reg[2]/NET0131  ;
	input \sice_DMR1_reg[3]/NET0131  ;
	input \sice_DMR1_reg[4]/NET0131  ;
	input \sice_DMR1_reg[5]/NET0131  ;
	input \sice_DMR1_reg[6]/NET0131  ;
	input \sice_DMR1_reg[7]/NET0131  ;
	input \sice_DMR1_reg[8]/NET0131  ;
	input \sice_DMR1_reg[9]/NET0131  ;
	input \sice_DMR2_reg[0]/NET0131  ;
	input \sice_DMR2_reg[10]/NET0131  ;
	input \sice_DMR2_reg[11]/NET0131  ;
	input \sice_DMR2_reg[12]/NET0131  ;
	input \sice_DMR2_reg[13]/NET0131  ;
	input \sice_DMR2_reg[14]/NET0131  ;
	input \sice_DMR2_reg[15]/NET0131  ;
	input \sice_DMR2_reg[16]/NET0131  ;
	input \sice_DMR2_reg[17]/NET0131  ;
	input \sice_DMR2_reg[1]/NET0131  ;
	input \sice_DMR2_reg[2]/NET0131  ;
	input \sice_DMR2_reg[3]/NET0131  ;
	input \sice_DMR2_reg[4]/NET0131  ;
	input \sice_DMR2_reg[5]/NET0131  ;
	input \sice_DMR2_reg[6]/NET0131  ;
	input \sice_DMR2_reg[7]/NET0131  ;
	input \sice_DMR2_reg[8]/NET0131  ;
	input \sice_DMR2_reg[9]/NET0131  ;
	input \sice_GOICE_1_reg/NET0131  ;
	input \sice_GOICE_2_reg/NET0131  ;
	input \sice_GOICE_s1_reg/NET0131  ;
	input \sice_GOICE_syn_reg/P0001  ;
	input \sice_GO_NX_reg/NET0131  ;
	input \sice_GO_NXi_reg/NET0131  ;
	input \sice_HALT_E_reg/P0001  ;
	input \sice_IAR_reg[0]/NET0131  ;
	input \sice_IAR_reg[1]/NET0131  ;
	input \sice_IAR_reg[2]/NET0131  ;
	input \sice_IAR_reg[3]/NET0131  ;
	input \sice_IBR1_reg[0]/P0001  ;
	input \sice_IBR1_reg[10]/P0001  ;
	input \sice_IBR1_reg[11]/P0001  ;
	input \sice_IBR1_reg[12]/P0001  ;
	input \sice_IBR1_reg[13]/P0001  ;
	input \sice_IBR1_reg[14]/P0001  ;
	input \sice_IBR1_reg[15]/P0001  ;
	input \sice_IBR1_reg[16]/P0001  ;
	input \sice_IBR1_reg[17]/P0001  ;
	input \sice_IBR1_reg[1]/P0001  ;
	input \sice_IBR1_reg[2]/P0001  ;
	input \sice_IBR1_reg[3]/P0001  ;
	input \sice_IBR1_reg[4]/P0001  ;
	input \sice_IBR1_reg[5]/P0001  ;
	input \sice_IBR1_reg[6]/P0001  ;
	input \sice_IBR1_reg[7]/P0001  ;
	input \sice_IBR1_reg[8]/P0001  ;
	input \sice_IBR1_reg[9]/P0001  ;
	input \sice_IBR2_reg[0]/P0001  ;
	input \sice_IBR2_reg[10]/P0001  ;
	input \sice_IBR2_reg[11]/P0001  ;
	input \sice_IBR2_reg[12]/P0001  ;
	input \sice_IBR2_reg[13]/P0001  ;
	input \sice_IBR2_reg[14]/P0001  ;
	input \sice_IBR2_reg[15]/P0001  ;
	input \sice_IBR2_reg[16]/P0001  ;
	input \sice_IBR2_reg[17]/P0001  ;
	input \sice_IBR2_reg[1]/P0001  ;
	input \sice_IBR2_reg[2]/P0001  ;
	input \sice_IBR2_reg[3]/P0001  ;
	input \sice_IBR2_reg[4]/P0001  ;
	input \sice_IBR2_reg[5]/P0001  ;
	input \sice_IBR2_reg[6]/P0001  ;
	input \sice_IBR2_reg[7]/P0001  ;
	input \sice_IBR2_reg[8]/P0001  ;
	input \sice_IBR2_reg[9]/P0001  ;
	input \sice_ICS_reg[0]/NET0131  ;
	input \sice_ICS_reg[1]/NET0131  ;
	input \sice_ICS_reg[2]/NET0131  ;
	input \sice_ICYC_clr_reg/NET0131  ;
	input \sice_ICYC_en_reg/NET0131  ;
	input \sice_ICYC_en_syn_reg/P0001  ;
	input \sice_ICYC_reg[0]/NET0131  ;
	input \sice_ICYC_reg[10]/NET0131  ;
	input \sice_ICYC_reg[11]/NET0131  ;
	input \sice_ICYC_reg[12]/NET0131  ;
	input \sice_ICYC_reg[13]/NET0131  ;
	input \sice_ICYC_reg[14]/NET0131  ;
	input \sice_ICYC_reg[15]/NET0131  ;
	input \sice_ICYC_reg[16]/NET0131  ;
	input \sice_ICYC_reg[17]/NET0131  ;
	input \sice_ICYC_reg[18]/NET0131  ;
	input \sice_ICYC_reg[19]/NET0131  ;
	input \sice_ICYC_reg[1]/NET0131  ;
	input \sice_ICYC_reg[20]/NET0131  ;
	input \sice_ICYC_reg[21]/NET0131  ;
	input \sice_ICYC_reg[22]/NET0131  ;
	input \sice_ICYC_reg[23]/NET0131  ;
	input \sice_ICYC_reg[2]/NET0131  ;
	input \sice_ICYC_reg[3]/NET0131  ;
	input \sice_ICYC_reg[4]/NET0131  ;
	input \sice_ICYC_reg[5]/NET0131  ;
	input \sice_ICYC_reg[6]/NET0131  ;
	input \sice_ICYC_reg[7]/NET0131  ;
	input \sice_ICYC_reg[8]/NET0131  ;
	input \sice_ICYC_reg[9]/NET0131  ;
	input \sice_IDONE_reg/NET0131  ;
	input \sice_IIRC_reg[0]/NET0131  ;
	input \sice_IIRC_reg[10]/NET0131  ;
	input \sice_IIRC_reg[11]/NET0131  ;
	input \sice_IIRC_reg[12]/NET0131  ;
	input \sice_IIRC_reg[13]/NET0131  ;
	input \sice_IIRC_reg[14]/NET0131  ;
	input \sice_IIRC_reg[15]/NET0131  ;
	input \sice_IIRC_reg[16]/NET0131  ;
	input \sice_IIRC_reg[17]/NET0131  ;
	input \sice_IIRC_reg[18]/NET0131  ;
	input \sice_IIRC_reg[19]/NET0131  ;
	input \sice_IIRC_reg[1]/NET0131  ;
	input \sice_IIRC_reg[20]/NET0131  ;
	input \sice_IIRC_reg[21]/NET0131  ;
	input \sice_IIRC_reg[22]/NET0131  ;
	input \sice_IIRC_reg[23]/NET0131  ;
	input \sice_IIRC_reg[2]/NET0131  ;
	input \sice_IIRC_reg[3]/NET0131  ;
	input \sice_IIRC_reg[4]/NET0131  ;
	input \sice_IIRC_reg[5]/NET0131  ;
	input \sice_IIRC_reg[6]/NET0131  ;
	input \sice_IIRC_reg[7]/NET0131  ;
	input \sice_IIRC_reg[8]/NET0131  ;
	input \sice_IIRC_reg[9]/NET0131  ;
	input \sice_IMR1_reg[0]/NET0131  ;
	input \sice_IMR1_reg[10]/NET0131  ;
	input \sice_IMR1_reg[11]/NET0131  ;
	input \sice_IMR1_reg[12]/NET0131  ;
	input \sice_IMR1_reg[13]/NET0131  ;
	input \sice_IMR1_reg[14]/NET0131  ;
	input \sice_IMR1_reg[15]/NET0131  ;
	input \sice_IMR1_reg[16]/NET0131  ;
	input \sice_IMR1_reg[17]/NET0131  ;
	input \sice_IMR1_reg[1]/NET0131  ;
	input \sice_IMR1_reg[2]/NET0131  ;
	input \sice_IMR1_reg[3]/NET0131  ;
	input \sice_IMR1_reg[4]/NET0131  ;
	input \sice_IMR1_reg[5]/NET0131  ;
	input \sice_IMR1_reg[6]/NET0131  ;
	input \sice_IMR1_reg[7]/NET0131  ;
	input \sice_IMR1_reg[8]/NET0131  ;
	input \sice_IMR1_reg[9]/NET0131  ;
	input \sice_IMR2_reg[0]/NET0131  ;
	input \sice_IMR2_reg[10]/NET0131  ;
	input \sice_IMR2_reg[11]/NET0131  ;
	input \sice_IMR2_reg[12]/NET0131  ;
	input \sice_IMR2_reg[13]/NET0131  ;
	input \sice_IMR2_reg[14]/NET0131  ;
	input \sice_IMR2_reg[15]/NET0131  ;
	input \sice_IMR2_reg[16]/NET0131  ;
	input \sice_IMR2_reg[17]/NET0131  ;
	input \sice_IMR2_reg[1]/NET0131  ;
	input \sice_IMR2_reg[2]/NET0131  ;
	input \sice_IMR2_reg[3]/NET0131  ;
	input \sice_IMR2_reg[4]/NET0131  ;
	input \sice_IMR2_reg[5]/NET0131  ;
	input \sice_IMR2_reg[6]/NET0131  ;
	input \sice_IMR2_reg[7]/NET0131  ;
	input \sice_IMR2_reg[8]/NET0131  ;
	input \sice_IMR2_reg[9]/NET0131  ;
	input \sice_IRR_reg[0]/P0001  ;
	input \sice_IRR_reg[10]/P0001  ;
	input \sice_IRR_reg[11]/P0001  ;
	input \sice_IRR_reg[12]/P0001  ;
	input \sice_IRR_reg[13]/P0001  ;
	input \sice_IRR_reg[1]/P0001  ;
	input \sice_IRR_reg[2]/P0001  ;
	input \sice_IRR_reg[3]/P0001  ;
	input \sice_IRR_reg[4]/P0001  ;
	input \sice_IRR_reg[5]/P0001  ;
	input \sice_IRR_reg[6]/P0001  ;
	input \sice_IRR_reg[7]/P0001  ;
	input \sice_IRR_reg[8]/P0001  ;
	input \sice_IRR_reg[9]/P0001  ;
	input \sice_IRST_reg/NET0131  ;
	input \sice_IRST_syn_reg/P0001  ;
	input \sice_ITR_reg[0]/NET0131  ;
	input \sice_ITR_reg[1]/NET0131  ;
	input \sice_ITR_reg[2]/NET0131  ;
	input \sice_OE_reg/P0001  ;
	input \sice_RCS_reg[0]/NET0131  ;
	input \sice_RCS_reg[1]/NET0131  ;
	input \sice_RST_req_reg/NET0131  ;
	input \sice_SPC_reg[0]/P0001  ;
	input \sice_SPC_reg[10]/P0001  ;
	input \sice_SPC_reg[11]/P0001  ;
	input \sice_SPC_reg[12]/P0001  ;
	input \sice_SPC_reg[13]/P0001  ;
	input \sice_SPC_reg[14]/P0001  ;
	input \sice_SPC_reg[15]/P0001  ;
	input \sice_SPC_reg[16]/P0001  ;
	input \sice_SPC_reg[17]/P0001  ;
	input \sice_SPC_reg[18]/P0001  ;
	input \sice_SPC_reg[19]/P0001  ;
	input \sice_SPC_reg[1]/P0001  ;
	input \sice_SPC_reg[20]/P0001  ;
	input \sice_SPC_reg[21]/P0001  ;
	input \sice_SPC_reg[22]/P0001  ;
	input \sice_SPC_reg[23]/P0001  ;
	input \sice_SPC_reg[2]/P0001  ;
	input \sice_SPC_reg[3]/P0001  ;
	input \sice_SPC_reg[4]/P0001  ;
	input \sice_SPC_reg[5]/P0001  ;
	input \sice_SPC_reg[6]/P0001  ;
	input \sice_SPC_reg[7]/P0001  ;
	input \sice_SPC_reg[8]/P0001  ;
	input \sice_SPC_reg[9]/P0001  ;
	input \sice_UpdDR_sd1_reg/P0001  ;
	input \sice_UpdDR_sd2_reg/P0001  ;
	input \sice_idr0_reg_DO_reg[0]/P0001  ;
	input \sice_idr0_reg_DO_reg[10]/P0001  ;
	input \sice_idr0_reg_DO_reg[11]/P0001  ;
	input \sice_idr0_reg_DO_reg[1]/P0001  ;
	input \sice_idr0_reg_DO_reg[2]/P0001  ;
	input \sice_idr0_reg_DO_reg[3]/P0001  ;
	input \sice_idr0_reg_DO_reg[4]/P0001  ;
	input \sice_idr0_reg_DO_reg[5]/P0001  ;
	input \sice_idr0_reg_DO_reg[6]/P0001  ;
	input \sice_idr0_reg_DO_reg[7]/P0001  ;
	input \sice_idr0_reg_DO_reg[8]/P0001  ;
	input \sice_idr0_reg_DO_reg[9]/P0001  ;
	input \sice_idr1_reg_DO_reg[0]/P0001  ;
	input \sice_idr1_reg_DO_reg[10]/P0001  ;
	input \sice_idr1_reg_DO_reg[11]/P0001  ;
	input \sice_idr1_reg_DO_reg[1]/P0001  ;
	input \sice_idr1_reg_DO_reg[2]/P0001  ;
	input \sice_idr1_reg_DO_reg[3]/P0001  ;
	input \sice_idr1_reg_DO_reg[4]/P0001  ;
	input \sice_idr1_reg_DO_reg[5]/P0001  ;
	input \sice_idr1_reg_DO_reg[6]/P0001  ;
	input \sice_idr1_reg_DO_reg[7]/P0001  ;
	input \sice_idr1_reg_DO_reg[8]/P0001  ;
	input \sice_idr1_reg_DO_reg[9]/P0001  ;
	input \sport0_cfg_FSi_cnt_reg[0]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[10]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[11]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[12]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[13]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[14]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[15]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[1]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[2]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[3]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[4]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[5]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[6]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[7]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[8]/NET0131  ;
	input \sport0_cfg_FSi_cnt_reg[9]/NET0131  ;
	input \sport0_cfg_FSi_reg/NET0131  ;
	input \sport0_cfg_RFSg_d1_reg/NET0131  ;
	input \sport0_cfg_RFSg_d2_reg/NET0131  ;
	input \sport0_cfg_RFSg_d3_reg/NET0131  ;
	input \sport0_cfg_RFSgi_d_reg/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[0]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[10]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[11]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[12]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[13]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[14]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[15]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[1]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[2]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[3]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[4]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[5]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[6]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[7]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[8]/NET0131  ;
	input \sport0_cfg_SCLKi_cnt_reg[9]/NET0131  ;
	input \sport0_cfg_SCLKi_h_reg/NET0131  ;
	input \sport0_cfg_SP_ENg_D1_reg/P0001  ;
	input \sport0_cfg_SP_ENg_reg/NET0131  ;
	input \sport0_cfg_TFSg_d1_reg/NET0131  ;
	input \sport0_cfg_TFSg_d2_reg/NET0131  ;
	input \sport0_cfg_TFSg_d3_reg/NET0131  ;
	input \sport0_cfg_TFSgi_d_reg/NET0131  ;
	input \sport0_regs_AUTO_a_reg[12]/NET0131  ;
	input \sport0_regs_AUTO_a_reg[13]/NET0131  ;
	input \sport0_regs_AUTO_a_reg[14]/NET0131  ;
	input \sport0_regs_AUTO_a_reg[15]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[11]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[7]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[8]/NET0131  ;
	input \sport0_regs_AUTOreg_DO_reg[9]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[11]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[12]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[13]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[14]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[15]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[7]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[8]/NET0131  ;
	input \sport0_regs_FSDIVreg_DO_reg[9]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[7]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[8]/NET0131  ;
	input \sport0_regs_MWORDreg_DO_reg[9]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
	input \sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[0]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[10]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[11]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[12]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[13]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[15]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[1]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[2]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[3]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[4]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[5]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[6]/NET0131  ;
	input \sport0_regs_SCTLreg_DO_reg[7]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[0]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[1]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[2]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[3]/NET0131  ;
	input \sport0_rxctl_Bcnt_reg[4]/NET0131  ;
	input \sport0_rxctl_ISRa_reg/P0001  ;
	input \sport0_rxctl_LMcnt_reg[0]/NET0131  ;
	input \sport0_rxctl_LMcnt_reg[1]/NET0131  ;
	input \sport0_rxctl_LMcnt_reg[2]/NET0131  ;
	input \sport0_rxctl_LMcnt_reg[3]/NET0131  ;
	input \sport0_rxctl_LMcnt_reg[4]/NET0131  ;
	input \sport0_rxctl_RCS_reg[0]/NET0131  ;
	input \sport0_rxctl_RCS_reg[1]/NET0131  ;
	input \sport0_rxctl_RCS_reg[2]/NET0131  ;
	input \sport0_rxctl_RSreq_reg/NET0131  ;
	input \sport0_rxctl_RXSHT_reg[0]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[10]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[11]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[12]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[13]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[14]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[15]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[1]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[2]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[3]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[4]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[5]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[6]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[7]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[8]/P0001  ;
	input \sport0_rxctl_RXSHT_reg[9]/P0001  ;
	input \sport0_rxctl_RX_reg[0]/P0001  ;
	input \sport0_rxctl_RX_reg[10]/P0001  ;
	input \sport0_rxctl_RX_reg[11]/P0001  ;
	input \sport0_rxctl_RX_reg[12]/P0001  ;
	input \sport0_rxctl_RX_reg[13]/P0001  ;
	input \sport0_rxctl_RX_reg[14]/P0001  ;
	input \sport0_rxctl_RX_reg[15]/P0001  ;
	input \sport0_rxctl_RX_reg[1]/P0001  ;
	input \sport0_rxctl_RX_reg[2]/P0001  ;
	input \sport0_rxctl_RX_reg[3]/P0001  ;
	input \sport0_rxctl_RX_reg[4]/P0001  ;
	input \sport0_rxctl_RX_reg[5]/P0001  ;
	input \sport0_rxctl_RX_reg[6]/P0001  ;
	input \sport0_rxctl_RX_reg[7]/P0001  ;
	input \sport0_rxctl_RX_reg[8]/P0001  ;
	input \sport0_rxctl_RX_reg[9]/P0001  ;
	input \sport0_rxctl_SLOT1_EXT_reg[2]/NET0131  ;
	input \sport0_rxctl_SLOT1_EXT_reg[3]/NET0131  ;
	input \sport0_rxctl_TAG_SLOT_reg/P0001  ;
	input \sport0_rxctl_Wcnt_reg[0]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[1]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[2]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[3]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[4]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[5]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[6]/NET0131  ;
	input \sport0_rxctl_Wcnt_reg[7]/NET0131  ;
	input \sport0_rxctl_a_sync1_reg/P0001  ;
	input \sport0_rxctl_a_sync2_reg/P0001  ;
	input \sport0_rxctl_ldRX_cmp_reg/P0001  ;
	input \sport0_rxctl_sht2nd_reg/P0001  ;
	input \sport0_txctl_Bcnt_reg[0]/NET0131  ;
	input \sport0_txctl_Bcnt_reg[1]/NET0131  ;
	input \sport0_txctl_Bcnt_reg[2]/NET0131  ;
	input \sport0_txctl_Bcnt_reg[3]/NET0131  ;
	input \sport0_txctl_Bcnt_reg[4]/NET0131  ;
	input \sport0_txctl_SP_EN_D1_reg/P0001  ;
	input \sport0_txctl_TCS_reg[0]/NET0131  ;
	input \sport0_txctl_TCS_reg[1]/NET0131  ;
	input \sport0_txctl_TCS_reg[2]/NET0131  ;
	input \sport0_txctl_TSreq_reg/NET0131  ;
	input \sport0_txctl_TSreqi_reg/NET0131  ;
	input \sport0_txctl_TXSHT_reg[0]/P0001  ;
	input \sport0_txctl_TXSHT_reg[10]/P0001  ;
	input \sport0_txctl_TXSHT_reg[11]/P0001  ;
	input \sport0_txctl_TXSHT_reg[12]/P0001  ;
	input \sport0_txctl_TXSHT_reg[13]/P0001  ;
	input \sport0_txctl_TXSHT_reg[14]/P0001  ;
	input \sport0_txctl_TXSHT_reg[15]/P0001  ;
	input \sport0_txctl_TXSHT_reg[1]/P0001  ;
	input \sport0_txctl_TXSHT_reg[2]/P0001  ;
	input \sport0_txctl_TXSHT_reg[3]/P0001  ;
	input \sport0_txctl_TXSHT_reg[4]/P0001  ;
	input \sport0_txctl_TXSHT_reg[5]/P0001  ;
	input \sport0_txctl_TXSHT_reg[6]/P0001  ;
	input \sport0_txctl_TXSHT_reg[7]/P0001  ;
	input \sport0_txctl_TXSHT_reg[8]/P0001  ;
	input \sport0_txctl_TXSHT_reg[9]/P0001  ;
	input \sport0_txctl_TX_reg[0]/P0001  ;
	input \sport0_txctl_TX_reg[10]/P0001  ;
	input \sport0_txctl_TX_reg[11]/P0001  ;
	input \sport0_txctl_TX_reg[12]/P0001  ;
	input \sport0_txctl_TX_reg[13]/P0001  ;
	input \sport0_txctl_TX_reg[14]/P0001  ;
	input \sport0_txctl_TX_reg[15]/P0001  ;
	input \sport0_txctl_TX_reg[1]/P0001  ;
	input \sport0_txctl_TX_reg[2]/P0001  ;
	input \sport0_txctl_TX_reg[3]/P0001  ;
	input \sport0_txctl_TX_reg[4]/P0001  ;
	input \sport0_txctl_TX_reg[5]/P0001  ;
	input \sport0_txctl_TX_reg[6]/P0001  ;
	input \sport0_txctl_TX_reg[7]/P0001  ;
	input \sport0_txctl_TX_reg[8]/P0001  ;
	input \sport0_txctl_TX_reg[9]/P0001  ;
	input \sport0_txctl_Wcnt_reg[0]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[1]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[2]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[3]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[4]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[5]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[6]/NET0131  ;
	input \sport0_txctl_Wcnt_reg[7]/NET0131  ;
	input \sport0_txctl_b_sync1_reg/P0001  ;
	input \sport0_txctl_c_sync1_reg/P0001  ;
	input \sport0_txctl_c_sync2_reg/P0001  ;
	input \sport0_txctl_ldTX_cmp_reg/P0001  ;
	input \sport1_cfg_FSi_cnt_reg[0]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[10]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[11]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[12]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[13]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[14]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[15]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[1]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[2]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[3]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[4]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[5]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[6]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[7]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[8]/NET0131  ;
	input \sport1_cfg_FSi_cnt_reg[9]/NET0131  ;
	input \sport1_cfg_FSi_reg/NET0131  ;
	input \sport1_cfg_RFSg_d1_reg/NET0131  ;
	input \sport1_cfg_RFSg_d2_reg/NET0131  ;
	input \sport1_cfg_RFSg_d3_reg/NET0131  ;
	input \sport1_cfg_RFSgi_d_reg/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[0]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[10]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[11]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[12]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[13]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[14]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[15]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[1]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[2]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[3]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[4]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[5]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[6]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[7]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[8]/NET0131  ;
	input \sport1_cfg_SCLKi_cnt_reg[9]/NET0131  ;
	input \sport1_cfg_SCLKi_h_reg/NET0131  ;
	input \sport1_cfg_SP_ENg_D1_reg/P0001  ;
	input \sport1_cfg_SP_ENg_reg/NET0131  ;
	input \sport1_cfg_TFSg_d1_reg/NET0131  ;
	input \sport1_cfg_TFSg_d2_reg/NET0131  ;
	input \sport1_cfg_TFSg_d3_reg/NET0131  ;
	input \sport1_cfg_TFSgi_d_reg/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[11]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[7]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[8]/NET0131  ;
	input \sport1_regs_AUTOreg_DO_reg[9]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[11]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[12]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[13]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[14]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[15]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[7]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[8]/NET0131  ;
	input \sport1_regs_FSDIVreg_DO_reg[9]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[7]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[8]/NET0131  ;
	input \sport1_regs_MWORDreg_DO_reg[9]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131  ;
	input \sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[0]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[10]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[11]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[12]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[13]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[15]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[1]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[2]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[3]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[4]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[5]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[6]/NET0131  ;
	input \sport1_regs_SCTLreg_DO_reg[7]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[0]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[1]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[2]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[3]/NET0131  ;
	input \sport1_rxctl_Bcnt_reg[4]/NET0131  ;
	input \sport1_rxctl_ISRa_reg/P0001  ;
	input \sport1_rxctl_LMcnt_reg[0]/NET0131  ;
	input \sport1_rxctl_LMcnt_reg[1]/NET0131  ;
	input \sport1_rxctl_LMcnt_reg[2]/NET0131  ;
	input \sport1_rxctl_LMcnt_reg[3]/NET0131  ;
	input \sport1_rxctl_LMcnt_reg[4]/NET0131  ;
	input \sport1_rxctl_RCS_reg[0]/NET0131  ;
	input \sport1_rxctl_RCS_reg[1]/NET0131  ;
	input \sport1_rxctl_RCS_reg[2]/NET0131  ;
	input \sport1_rxctl_RSreq_reg/NET0131  ;
	input \sport1_rxctl_RXSHT_reg[0]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[10]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[11]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[12]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[13]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[14]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[15]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[1]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[2]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[3]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[4]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[5]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[6]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[7]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[8]/P0001  ;
	input \sport1_rxctl_RXSHT_reg[9]/P0001  ;
	input \sport1_rxctl_RX_reg[0]/P0001  ;
	input \sport1_rxctl_RX_reg[10]/P0001  ;
	input \sport1_rxctl_RX_reg[11]/P0001  ;
	input \sport1_rxctl_RX_reg[12]/P0001  ;
	input \sport1_rxctl_RX_reg[13]/P0001  ;
	input \sport1_rxctl_RX_reg[14]/P0001  ;
	input \sport1_rxctl_RX_reg[15]/P0001  ;
	input \sport1_rxctl_RX_reg[1]/P0001  ;
	input \sport1_rxctl_RX_reg[2]/P0001  ;
	input \sport1_rxctl_RX_reg[3]/P0001  ;
	input \sport1_rxctl_RX_reg[4]/P0001  ;
	input \sport1_rxctl_RX_reg[5]/P0001  ;
	input \sport1_rxctl_RX_reg[6]/P0001  ;
	input \sport1_rxctl_RX_reg[7]/P0001  ;
	input \sport1_rxctl_RX_reg[8]/P0001  ;
	input \sport1_rxctl_RX_reg[9]/P0001  ;
	input \sport1_rxctl_SLOT1_EXT_reg[2]/NET0131  ;
	input \sport1_rxctl_SLOT1_EXT_reg[3]/NET0131  ;
	input \sport1_rxctl_TAG_SLOT_reg/P0001  ;
	input \sport1_rxctl_Wcnt_reg[0]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[1]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[2]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[3]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[4]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[5]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[6]/NET0131  ;
	input \sport1_rxctl_Wcnt_reg[7]/NET0131  ;
	input \sport1_rxctl_a_sync1_reg/P0001  ;
	input \sport1_rxctl_a_sync2_reg/P0001  ;
	input \sport1_rxctl_sht2nd_reg/P0001  ;
	input \sport1_txctl_Bcnt_reg[0]/NET0131  ;
	input \sport1_txctl_Bcnt_reg[1]/NET0131  ;
	input \sport1_txctl_Bcnt_reg[2]/NET0131  ;
	input \sport1_txctl_Bcnt_reg[3]/NET0131  ;
	input \sport1_txctl_Bcnt_reg[4]/NET0131  ;
	input \sport1_txctl_SP_EN_D1_reg/P0001  ;
	input \sport1_txctl_TCS_reg[0]/NET0131  ;
	input \sport1_txctl_TCS_reg[1]/NET0131  ;
	input \sport1_txctl_TCS_reg[2]/NET0131  ;
	input \sport1_txctl_TSreq_reg/NET0131  ;
	input \sport1_txctl_TSreqi_reg/NET0131  ;
	input \sport1_txctl_TXSHT_reg[0]/P0001  ;
	input \sport1_txctl_TXSHT_reg[10]/P0001  ;
	input \sport1_txctl_TXSHT_reg[11]/P0001  ;
	input \sport1_txctl_TXSHT_reg[12]/P0001  ;
	input \sport1_txctl_TXSHT_reg[13]/P0001  ;
	input \sport1_txctl_TXSHT_reg[14]/P0001  ;
	input \sport1_txctl_TXSHT_reg[15]/P0001  ;
	input \sport1_txctl_TXSHT_reg[1]/P0001  ;
	input \sport1_txctl_TXSHT_reg[2]/P0001  ;
	input \sport1_txctl_TXSHT_reg[3]/P0001  ;
	input \sport1_txctl_TXSHT_reg[4]/P0001  ;
	input \sport1_txctl_TXSHT_reg[5]/P0001  ;
	input \sport1_txctl_TXSHT_reg[6]/P0001  ;
	input \sport1_txctl_TXSHT_reg[7]/P0001  ;
	input \sport1_txctl_TXSHT_reg[8]/P0001  ;
	input \sport1_txctl_TXSHT_reg[9]/P0001  ;
	input \sport1_txctl_TX_reg[0]/P0001  ;
	input \sport1_txctl_TX_reg[10]/P0001  ;
	input \sport1_txctl_TX_reg[11]/P0001  ;
	input \sport1_txctl_TX_reg[12]/P0001  ;
	input \sport1_txctl_TX_reg[13]/P0001  ;
	input \sport1_txctl_TX_reg[14]/P0001  ;
	input \sport1_txctl_TX_reg[15]/P0001  ;
	input \sport1_txctl_TX_reg[1]/P0001  ;
	input \sport1_txctl_TX_reg[2]/P0001  ;
	input \sport1_txctl_TX_reg[3]/P0001  ;
	input \sport1_txctl_TX_reg[4]/P0001  ;
	input \sport1_txctl_TX_reg[5]/P0001  ;
	input \sport1_txctl_TX_reg[6]/P0001  ;
	input \sport1_txctl_TX_reg[7]/P0001  ;
	input \sport1_txctl_TX_reg[8]/P0001  ;
	input \sport1_txctl_TX_reg[9]/P0001  ;
	input \sport1_txctl_Wcnt_reg[0]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[1]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[2]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[3]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[4]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[5]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[6]/NET0131  ;
	input \sport1_txctl_Wcnt_reg[7]/NET0131  ;
	input \sport1_txctl_c_sync1_reg/P0001  ;
	input \sport1_txctl_c_sync2_reg/P0001  ;
	input \tm_MSTAT5_syn_reg/NET0131  ;
	input \tm_TCR_TMP_reg[0]/NET0131  ;
	input \tm_TCR_TMP_reg[10]/NET0131  ;
	input \tm_TCR_TMP_reg[11]/NET0131  ;
	input \tm_TCR_TMP_reg[12]/NET0131  ;
	input \tm_TCR_TMP_reg[13]/NET0131  ;
	input \tm_TCR_TMP_reg[14]/NET0131  ;
	input \tm_TCR_TMP_reg[15]/NET0131  ;
	input \tm_TCR_TMP_reg[1]/NET0131  ;
	input \tm_TCR_TMP_reg[2]/NET0131  ;
	input \tm_TCR_TMP_reg[3]/NET0131  ;
	input \tm_TCR_TMP_reg[4]/NET0131  ;
	input \tm_TCR_TMP_reg[5]/NET0131  ;
	input \tm_TCR_TMP_reg[6]/NET0131  ;
	input \tm_TCR_TMP_reg[7]/NET0131  ;
	input \tm_TCR_TMP_reg[8]/NET0131  ;
	input \tm_TCR_TMP_reg[9]/NET0131  ;
	input \tm_TINT_GEN1_reg/NET0131  ;
	input \tm_TINT_GEN2_reg/NET0131  ;
	input \tm_TSR_TMP_reg[0]/NET0131  ;
	input \tm_TSR_TMP_reg[1]/NET0131  ;
	input \tm_TSR_TMP_reg[2]/NET0131  ;
	input \tm_TSR_TMP_reg[3]/NET0131  ;
	input \tm_TSR_TMP_reg[4]/NET0131  ;
	input \tm_TSR_TMP_reg[5]/NET0131  ;
	input \tm_TSR_TMP_reg[6]/NET0131  ;
	input \tm_TSR_TMP_reg[7]/NET0131  ;
	input \tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131  ;
	input \tm_WR_TCR_TMP_GEN1_reg/P0001  ;
	input \tm_WR_TCR_TMP_GEN2_reg/P0001  ;
	input \tm_WR_TCR_p_reg/P0001  ;
	input \tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131  ;
	input \tm_WR_TSR_TMP_GEN1_reg/P0001  ;
	input \tm_WR_TSR_TMP_GEN2_reg/P0001  ;
	input \tm_WR_TSR_p_reg/P0001  ;
	input \tm_tcr_reg_DO_reg[0]/NET0131  ;
	input \tm_tcr_reg_DO_reg[10]/NET0131  ;
	input \tm_tcr_reg_DO_reg[11]/NET0131  ;
	input \tm_tcr_reg_DO_reg[12]/NET0131  ;
	input \tm_tcr_reg_DO_reg[13]/NET0131  ;
	input \tm_tcr_reg_DO_reg[14]/NET0131  ;
	input \tm_tcr_reg_DO_reg[15]/NET0131  ;
	input \tm_tcr_reg_DO_reg[1]/NET0131  ;
	input \tm_tcr_reg_DO_reg[2]/NET0131  ;
	input \tm_tcr_reg_DO_reg[3]/NET0131  ;
	input \tm_tcr_reg_DO_reg[4]/NET0131  ;
	input \tm_tcr_reg_DO_reg[5]/NET0131  ;
	input \tm_tcr_reg_DO_reg[6]/NET0131  ;
	input \tm_tcr_reg_DO_reg[7]/NET0131  ;
	input \tm_tcr_reg_DO_reg[8]/NET0131  ;
	input \tm_tcr_reg_DO_reg[9]/NET0131  ;
	input \tm_tpr_reg_DO_reg[0]/NET0131  ;
	input \tm_tpr_reg_DO_reg[10]/NET0131  ;
	input \tm_tpr_reg_DO_reg[11]/NET0131  ;
	input \tm_tpr_reg_DO_reg[12]/NET0131  ;
	input \tm_tpr_reg_DO_reg[13]/NET0131  ;
	input \tm_tpr_reg_DO_reg[14]/NET0131  ;
	input \tm_tpr_reg_DO_reg[15]/NET0131  ;
	input \tm_tpr_reg_DO_reg[1]/NET0131  ;
	input \tm_tpr_reg_DO_reg[2]/NET0131  ;
	input \tm_tpr_reg_DO_reg[3]/NET0131  ;
	input \tm_tpr_reg_DO_reg[4]/NET0131  ;
	input \tm_tpr_reg_DO_reg[5]/NET0131  ;
	input \tm_tpr_reg_DO_reg[6]/NET0131  ;
	input \tm_tpr_reg_DO_reg[7]/NET0131  ;
	input \tm_tpr_reg_DO_reg[8]/NET0131  ;
	input \tm_tpr_reg_DO_reg[9]/NET0131  ;
	input \tm_tsr_reg_DO_reg[0]/NET0131  ;
	input \tm_tsr_reg_DO_reg[1]/NET0131  ;
	input \tm_tsr_reg_DO_reg[2]/NET0131  ;
	input \tm_tsr_reg_DO_reg[3]/NET0131  ;
	input \tm_tsr_reg_DO_reg[4]/NET0131  ;
	input \tm_tsr_reg_DO_reg[5]/NET0131  ;
	input \tm_tsr_reg_DO_reg[6]/NET0131  ;
	input \tm_tsr_reg_DO_reg[7]/NET0131  ;
	input \tm_tsr_reg_DO_reg[8]/NET0131  ;
	output CLKO_pad ;
	output \CMAinx[0]_pad  ;
	output \CMAinx[10]_pad  ;
	output \CMAinx[11]_pad  ;
	output \CMAinx[1]_pad  ;
	output \CMAinx[2]_pad  ;
	output \CMAinx[3]_pad  ;
	output \CMAinx[4]_pad  ;
	output \CMAinx[5]_pad  ;
	output \CMAinx[6]_pad  ;
	output \CMAinx[7]_pad  ;
	output \CMAinx[8]_pad  ;
	output \CMAinx[9]_pad  ;
	output CMSn_pad ;
	output CM_cs_pad ;
	output \CM_wd[0]_pad  ;
	output \CM_wd[10]_pad  ;
	output \CM_wd[11]_pad  ;
	output \CM_wd[12]_pad  ;
	output \CM_wd[13]_pad  ;
	output \CM_wd[14]_pad  ;
	output \CM_wd[15]_pad  ;
	output \CM_wd[16]_pad  ;
	output \CM_wd[17]_pad  ;
	output \CM_wd[18]_pad  ;
	output \CM_wd[19]_pad  ;
	output \CM_wd[1]_pad  ;
	output \CM_wd[20]_pad  ;
	output \CM_wd[21]_pad  ;
	output \CM_wd[22]_pad  ;
	output \CM_wd[23]_pad  ;
	output \CM_wd[2]_pad  ;
	output \CM_wd[3]_pad  ;
	output \CM_wd[4]_pad  ;
	output \CM_wd[5]_pad  ;
	output \CM_wd[6]_pad  ;
	output \CM_wd[7]_pad  ;
	output \CM_wd[8]_pad  ;
	output \CM_wd[9]_pad  ;
	output CM_web_pad ;
	output \CMo_cs0_pad  ;
	output \CMo_cs1_pad  ;
	output \CMo_cs2_pad  ;
	output \CMo_cs3_pad  ;
	output \CMo_cs4_pad  ;
	output \CMo_cs5_pad  ;
	output \CMo_cs6_pad  ;
	output \CMo_cs7_pad  ;
	output \DMAinx[0]_pad  ;
	output \DMAinx[10]_pad  ;
	output \DMAinx[11]_pad  ;
	output \DMAinx[12]_pad  ;
	output \DMAinx[13]_pad  ;
	output \DMAinx[1]_pad  ;
	output \DMAinx[2]_pad  ;
	output \DMAinx[3]_pad  ;
	output \DMAinx[4]_pad  ;
	output \DMAinx[5]_pad  ;
	output \DMAinx[6]_pad  ;
	output \DMAinx[7]_pad  ;
	output \DMAinx[8]_pad  ;
	output \DMAinx[9]_pad  ;
	output DMSn_pad ;
	output DM_cs_pad ;
	output \DM_wd[0]_pad  ;
	output \DM_wd[10]_pad  ;
	output \DM_wd[11]_pad  ;
	output \DM_wd[12]_pad  ;
	output \DM_wd[13]_pad  ;
	output \DM_wd[14]_pad  ;
	output \DM_wd[15]_pad  ;
	output \DM_wd[1]_pad  ;
	output \DM_wd[2]_pad  ;
	output \DM_wd[3]_pad  ;
	output \DM_wd[4]_pad  ;
	output \DM_wd[5]_pad  ;
	output \DM_wd[6]_pad  ;
	output \DM_wd[7]_pad  ;
	output \DM_wd[8]_pad  ;
	output \DM_wd[9]_pad  ;
	output \DMo_cs0_pad  ;
	output \DMo_cs1_pad  ;
	output \DMo_cs2_pad  ;
	output \DMo_cs3_pad  ;
	output \DMo_cs4_pad  ;
	output \DMo_cs5_pad  ;
	output \DMo_cs6_pad  ;
	output \DMo_cs7_pad  ;
	output \DSPCLK_cm1_pad  ;
	output \EA_do[0]_pad  ;
	output \EA_do[10]_pad  ;
	output \EA_do[12]_pad  ;
	output \EA_do[13]_pad  ;
	output \EA_do[14]_pad  ;
	output \EA_do[1]_pad  ;
	output \EA_do[2]_pad  ;
	output \EA_do[3]_pad  ;
	output \EA_do[4]_pad  ;
	output \EA_do[5]_pad  ;
	output \EA_do[6]_pad  ;
	output \EA_do[7]_pad  ;
	output \EA_do[8]_pad  ;
	output \EA_do[9]_pad  ;
	output EA_oe_pad ;
	output \ED_do[0]_pad  ;
	output \ED_do[10]_pad  ;
	output \ED_do[11]_pad  ;
	output \ED_do[12]_pad  ;
	output \ED_do[13]_pad  ;
	output \ED_do[14]_pad  ;
	output \ED_do[15]_pad  ;
	output \ED_do[1]_pad  ;
	output \ED_do[2]_pad  ;
	output \ED_do[3]_pad  ;
	output \ED_do[4]_pad  ;
	output \ED_do[5]_pad  ;
	output \ED_do[6]_pad  ;
	output \ED_do[7]_pad  ;
	output \ED_do[8]_pad  ;
	output \ED_do[9]_pad  ;
	output \ED_oe_14_8_pad  ;
	output \ED_oe_7_0_pad  ;
	output \IAD_do[0]_pad  ;
	output \IAD_do[10]_pad  ;
	output \IAD_do[11]_pad  ;
	output \IAD_do[12]_pad  ;
	output \IAD_do[13]_pad  ;
	output \IAD_do[14]_pad  ;
	output \IAD_do[15]_pad  ;
	output \IAD_do[1]_pad  ;
	output \IAD_do[2]_pad  ;
	output \IAD_do[3]_pad  ;
	output \IAD_do[4]_pad  ;
	output \IAD_do[5]_pad  ;
	output \IAD_do[6]_pad  ;
	output \IAD_do[7]_pad  ;
	output \IAD_do[8]_pad  ;
	output \IAD_do[9]_pad  ;
	output IAD_oe_pad ;
	output IDoe_pad ;
	output IOSn_pad ;
	output \PMAinx[0]_pad  ;
	output \PMAinx[10]_pad  ;
	output \PMAinx[11]_pad  ;
	output \PMAinx[1]_pad  ;
	output \PMAinx[2]_pad  ;
	output \PMAinx[3]_pad  ;
	output \PMAinx[4]_pad  ;
	output \PMAinx[5]_pad  ;
	output \PMAinx[6]_pad  ;
	output \PMAinx[7]_pad  ;
	output \PMAinx[8]_pad  ;
	output \PMAinx[9]_pad  ;
	output \PM_wd[0]_pad  ;
	output \PM_wd[10]_pad  ;
	output \PM_wd[11]_pad  ;
	output \PM_wd[12]_pad  ;
	output \PM_wd[13]_pad  ;
	output \PM_wd[14]_pad  ;
	output \PM_wd[15]_pad  ;
	output \PM_wd[1]_pad  ;
	output \PM_wd[2]_pad  ;
	output \PM_wd[3]_pad  ;
	output \PM_wd[4]_pad  ;
	output \PM_wd[5]_pad  ;
	output \PM_wd[6]_pad  ;
	output \PM_wd[7]_pad  ;
	output \PM_wd[8]_pad  ;
	output \PM_wd[9]_pad  ;
	output \PMo_cs0_pad  ;
	output \PMo_cs1_pad  ;
	output \PMo_cs2_pad  ;
	output \PMo_cs3_pad  ;
	output \PMo_cs4_pad  ;
	output \PMo_cs5_pad  ;
	output \PMo_cs6_pad  ;
	output \PMo_cs7_pad  ;
	output \PMo_oe0_pad  ;
	output \RFS0_pad  ;
	output \RFS1_pad  ;
	output \SCLK0_pad  ;
	output \SCLK1_pad  ;
	output \TD0_pad  ;
	output \TD1_pad  ;
	output \TFS0_pad  ;
	output \TFS1_pad  ;
	output \T_ISn_syn_2  ;
	output WRn_pad ;
	output XTALoffn_pad ;
	output \_al_n0  ;
	output \bdma_BDMA_boot_reg/NET0131_reg_syn_3  ;
	output \bdma_BDMA_boot_reg/n0  ;
	output \bdma_BM_cyc_reg/P0000  ;
	output \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3  ;
	output \core_c_psq_MGNT_reg/P0001  ;
	output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3  ;
	output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3  ;
	output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3  ;
	output \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3  ;
	output \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3  ;
	output \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3  ;
	output \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3  ;
	output \emc_DMDreg_reg[8]/P0001_reg_syn_3  ;
	output \emc_DMDreg_reg[9]/P0001_reg_syn_3  ;
	output \emc_ECMcs_reg/P0001  ;
	output \emc_PMDreg_reg[8]/P0001_reg_syn_3  ;
	output \emc_PMDreg_reg[9]/P0001_reg_syn_3  ;
	output \g10/_0_  ;
	output \g1000/_0_  ;
	output \g10000/_0_  ;
	output \g10001/_0_  ;
	output \g10002/_0_  ;
	output \g10003/_0_  ;
	output \g10004/_0_  ;
	output \g10005/_0_  ;
	output \g10007/_0_  ;
	output \g10008/_0_  ;
	output \g10009/_0_  ;
	output \g1001/_3_  ;
	output \g10010/_0_  ;
	output \g10011/_0_  ;
	output \g10012/_0_  ;
	output \g10013/_0_  ;
	output \g10014/_0_  ;
	output \g10015/_0_  ;
	output \g10016/_0_  ;
	output \g10017/_0_  ;
	output \g10018/_0_  ;
	output \g10019/_0_  ;
	output \g1002/_3_  ;
	output \g10020/_0_  ;
	output \g10021/_0_  ;
	output \g10022/_0_  ;
	output \g10023/_0_  ;
	output \g10024/_0_  ;
	output \g10025/_0_  ;
	output \g10026/_0_  ;
	output \g10027/_0_  ;
	output \g10028/_0_  ;
	output \g10029/_0_  ;
	output \g1003/_0_  ;
	output \g10030/_0_  ;
	output \g10031/_0_  ;
	output \g10032/_0_  ;
	output \g10033/_0_  ;
	output \g10034/_0_  ;
	output \g10035/_0_  ;
	output \g10036/_0_  ;
	output \g10037/_0_  ;
	output \g10038/_0_  ;
	output \g10039/_0_  ;
	output \g10040/_0_  ;
	output \g10041/_0_  ;
	output \g10042/_0_  ;
	output \g10043/_0_  ;
	output \g10044/_0_  ;
	output \g10045/_0_  ;
	output \g10046/_0_  ;
	output \g10047/_0_  ;
	output \g10048/_0_  ;
	output \g10049/_0_  ;
	output \g10050/_0_  ;
	output \g10051/_0_  ;
	output \g10052/_0_  ;
	output \g10053/_0_  ;
	output \g10054/_0_  ;
	output \g10055/_0_  ;
	output \g10056/_0_  ;
	output \g10057/_0_  ;
	output \g10058/_0_  ;
	output \g10059/_0_  ;
	output \g10060/_0_  ;
	output \g10061/_0_  ;
	output \g10062/_0_  ;
	output \g10063/_0_  ;
	output \g10064/_0_  ;
	output \g10065/_0_  ;
	output \g10066/_0_  ;
	output \g10067/_0_  ;
	output \g10068/_0_  ;
	output \g10069/_0_  ;
	output \g10070/_0_  ;
	output \g10071/_0_  ;
	output \g10072/_0_  ;
	output \g10073/_0_  ;
	output \g10074/_0_  ;
	output \g10075/_0_  ;
	output \g10076/_0_  ;
	output \g10077/_0_  ;
	output \g10078/_0_  ;
	output \g10080/_0_  ;
	output \g10081/_0_  ;
	output \g10083/_0_  ;
	output \g10089/_0_  ;
	output \g1009/_0_  ;
	output \g10090/_0_  ;
	output \g10091/_0_  ;
	output \g10092/_0_  ;
	output \g10093/_0_  ;
	output \g10094/_0_  ;
	output \g1010/_0_  ;
	output \g10108/_3_  ;
	output \g1011/_0_  ;
	output \g10110/_0_  ;
	output \g10111/_0_  ;
	output \g10113/_3_  ;
	output \g10115/_3_  ;
	output \g1013/_0_  ;
	output \g1014/_0_  ;
	output \g10152/_0_  ;
	output \g10153/_0_  ;
	output \g10154/_0_  ;
	output \g10155/_0_  ;
	output \g10156/_0_  ;
	output \g10157/_0_  ;
	output \g10158/_0_  ;
	output \g10159/_0_  ;
	output \g1016/_0_  ;
	output \g10160/_0_  ;
	output \g10161/_0_  ;
	output \g10162/_0_  ;
	output \g10163/_0_  ;
	output \g10164/_0_  ;
	output \g10165/_0_  ;
	output \g1017/_0_  ;
	output \g10170/_3_  ;
	output \g1018/_0_  ;
	output \g10190/_3_  ;
	output \g10194/_3_  ;
	output \g10198/_0_  ;
	output \g10199/_0_  ;
	output \g102/_0_  ;
	output \g103/_0_  ;
	output \g104/_0_  ;
	output \g105/_0_  ;
	output \g10598/_0_  ;
	output \g106/_0_  ;
	output \g10667/_0_  ;
	output \g10683/_0_  ;
	output \g10685/_0_  ;
	output \g107/_0_  ;
	output \g10721/_0_  ;
	output \g10758/_0_  ;
	output \g10765/_0_  ;
	output \g10778/_0_  ;
	output \g10791/_0_  ;
	output \g108/_0_  ;
	output \g10887/_0_  ;
	output \g1089/_0_  ;
	output \g109/_0_  ;
	output \g1090/_0_  ;
	output \g1091/_0_  ;
	output \g1092/_0_  ;
	output \g10923/_0_  ;
	output \g1093/_0_  ;
	output \g10930/_0_  ;
	output \g10931/_0_  ;
	output \g10936/_0_  ;
	output \g1097/_0_  ;
	output \g11/_0_  ;
	output \g110/_0_  ;
	output \g1101/_0_  ;
	output \g11013/_0_  ;
	output \g1102/_0_  ;
	output \g1103/_0_  ;
	output \g11032/_0_  ;
	output \g1104/_0_  ;
	output \g1105/_0_  ;
	output \g1107/_0_  ;
	output \g11074/_0_  ;
	output \g11077/_0_  ;
	output \g1108/_0_  ;
	output \g1109/_0_  ;
	output \g11112/_0_  ;
	output \g11115/_0_  ;
	output \g11116/_0_  ;
	output \g11119/_0_  ;
	output \g11120/_0_  ;
	output \g1113/_0_  ;
	output \g1115/_0_  ;
	output \g1116/_0_  ;
	output \g1117/_0_  ;
	output \g11267/_0_  ;
	output \g11281/_0_  ;
	output \g11287/_0_  ;
	output \g11300/_0_  ;
	output \g11323/_0_  ;
	output \g11325/_2__syn_2  ;
	output \g11345/_2_  ;
	output \g11470/_0_  ;
	output \g11471/_0_  ;
	output \g11472/_0_  ;
	output \g11473/_0_  ;
	output \g11474/_0_  ;
	output \g11476/_0_  ;
	output \g11477/_0_  ;
	output \g11496/_0_  ;
	output \g11497/_0_  ;
	output \g11498/_0_  ;
	output \g11499/_0_  ;
	output \g11500/_0_  ;
	output \g11501/_0_  ;
	output \g11502/_0_  ;
	output \g11503/_0_  ;
	output \g11504/_0_  ;
	output \g11505/_0_  ;
	output \g11506/_0_  ;
	output \g11507/_0_  ;
	output \g11509/_0_  ;
	output \g11510/_0_  ;
	output \g11515/_0_  ;
	output \g11516/_0_  ;
	output \g11520/_0_  ;
	output \g11521/_0_  ;
	output \g11576/_0_  ;
	output \g11577/_0_  ;
	output \g11578/_0_  ;
	output \g11579/_0_  ;
	output \g11580/_0_  ;
	output \g11581/_0_  ;
	output \g11582/_0_  ;
	output \g11583/_0_  ;
	output \g11584/_0_  ;
	output \g11585/_0_  ;
	output \g11586/_0_  ;
	output \g11587/_0_  ;
	output \g11588/_0_  ;
	output \g11589/_0_  ;
	output \g11591/_0_  ;
	output \g11593/_0_  ;
	output \g11595/_0_  ;
	output \g11596/_0_  ;
	output \g11597/_0_  ;
	output \g11605/_0_  ;
	output \g11606/_0_  ;
	output \g11607/_0_  ;
	output \g11608/_0_  ;
	output \g11609/_0_  ;
	output \g11610/_0_  ;
	output \g11611/_0_  ;
	output \g11612/_0_  ;
	output \g11613/_0_  ;
	output \g11615/_0_  ;
	output \g11616/_0_  ;
	output \g11617/_0_  ;
	output \g11651/_3_  ;
	output \g11704/_0_  ;
	output \g11705/_0_  ;
	output \g11709/_0_  ;
	output \g11722/_0_  ;
	output \g11723/_0_  ;
	output \g119/_0_  ;
	output \g1192/_0_  ;
	output \g11994/_0_  ;
	output \g120/_0_  ;
	output \g1200/_0_  ;
	output \g12003/_0_  ;
	output \g1201/_0_  ;
	output \g12019/_0_  ;
	output \g1203/_3_  ;
	output \g1204/_3_  ;
	output \g1207/_0_  ;
	output \g1208/_0_  ;
	output \g12092/_0_  ;
	output \g1210/_0_  ;
	output \g1211/_0_  ;
	output \g1212/_0_  ;
	output \g1213/_0_  ;
	output \g12145/_0_  ;
	output \g12155/_0_  ;
	output \g12186/_0_  ;
	output \g12187/_0_  ;
	output \g12192/_0_  ;
	output \g12201/_0_  ;
	output \g12202/_0_  ;
	output \g12203/_0_  ;
	output \g12204/_0_  ;
	output \g12207/_0_  ;
	output \g12229/_3_  ;
	output \g12267/_0_  ;
	output \g12276/_0_  ;
	output \g12278/_0_  ;
	output \g12279/_0_  ;
	output \g12280/_0_  ;
	output \g12302/_0_  ;
	output \g12316/_0_  ;
	output \g12317/_0_  ;
	output \g12319/_0_  ;
	output \g12328/_3_  ;
	output \g1233/_0_  ;
	output \g12348/_0_  ;
	output \g12351/_0_  ;
	output \g12352/_0_  ;
	output \g12353/_0_  ;
	output \g12354/_0_  ;
	output \g12355/_0_  ;
	output \g1237/_0_  ;
	output \g124/_0_  ;
	output \g12444/_0_  ;
	output \g125/_0_  ;
	output \g12637/_0_  ;
	output \g12639/_0_  ;
	output \g12658/_0_  ;
	output \g12659/_0_  ;
	output \g12660/_0_  ;
	output \g12663/_0_  ;
	output \g12664/_0_  ;
	output \g12665/_0_  ;
	output \g12672/_3_  ;
	output \g12673/_3_  ;
	output \g12674/_3_  ;
	output \g12675/_3_  ;
	output \g12676/_3_  ;
	output \g12677/_3_  ;
	output \g12678/_0_  ;
	output \g12679/_3_  ;
	output \g12697/_3_  ;
	output \g12701/_3_  ;
	output \g12711/_2_  ;
	output \g12713/_2_  ;
	output \g12715/_2_  ;
	output \g12717/_2_  ;
	output \g12718/_2__syn_2  ;
	output \g1272/_0_  ;
	output \g12728/_1__syn_2  ;
	output \g12730/_3_  ;
	output \g12741/_1__syn_2  ;
	output \g12746/_0__syn_2  ;
	output \g12748/_0_  ;
	output \g12749/_0_  ;
	output \g12759/_1__syn_2  ;
	output \g12760/_0_  ;
	output \g12762/_0_  ;
	output \g12763/_0_  ;
	output \g12764/_0_  ;
	output \g12765/_0_  ;
	output \g12766/_0_  ;
	output \g12767/_0_  ;
	output \g12768/_0_  ;
	output \g12769/_0_  ;
	output \g12770/_0_  ;
	output \g12771/_0_  ;
	output \g12772/_0_  ;
	output \g12773/_0_  ;
	output \g12774/_0_  ;
	output \g12775/_0_  ;
	output \g12776/_0_  ;
	output \g12777/_0_  ;
	output \g12778/_0_  ;
	output \g12779/_0_  ;
	output \g1278/_0_  ;
	output \g12780/_0_  ;
	output \g12781/_0_  ;
	output \g12782/_0_  ;
	output \g12783/_0_  ;
	output \g12784/_0_  ;
	output \g12785/_0_  ;
	output \g12786/_0_  ;
	output \g12787/_0_  ;
	output \g12788/_0_  ;
	output \g12789/_0_  ;
	output \g12790/_0_  ;
	output \g12791/_0_  ;
	output \g12792/_0_  ;
	output \g12793/_0_  ;
	output \g12794/_0_  ;
	output \g12795/_0_  ;
	output \g12796/_0_  ;
	output \g12797/_0_  ;
	output \g12798/_0_  ;
	output \g12799/_0_  ;
	output \g12800/_0_  ;
	output \g12801/_0_  ;
	output \g12802/_0_  ;
	output \g12803/_0_  ;
	output \g12804/_0_  ;
	output \g12805/_0_  ;
	output \g12806/_0_  ;
	output \g12807/_0_  ;
	output \g12808/_0_  ;
	output \g12809/_0_  ;
	output \g1281/_0_  ;
	output \g12810/_0_  ;
	output \g12811/_0_  ;
	output \g12812/_0_  ;
	output \g12813/_0_  ;
	output \g12814/_0_  ;
	output \g12815/_0_  ;
	output \g12816/_0_  ;
	output \g12817/_0_  ;
	output \g12818/_0_  ;
	output \g12819/_0_  ;
	output \g1282/_0_  ;
	output \g12820/_0_  ;
	output \g12821/_0_  ;
	output \g12822/_0_  ;
	output \g12823/_0_  ;
	output \g12824/_0_  ;
	output \g12825/_0_  ;
	output \g12826/_0_  ;
	output \g12827/_0_  ;
	output \g12828/_0_  ;
	output \g12829/_0_  ;
	output \g12830/_0_  ;
	output \g12831/_0_  ;
	output \g12832/_0_  ;
	output \g12833/_0_  ;
	output \g12835/_0_  ;
	output \g12836/_0_  ;
	output \g12838/_0_  ;
	output \g12848/_0_  ;
	output \g12849/_0_  ;
	output \g1285/_0_  ;
	output \g12850/_0_  ;
	output \g12857/_0_  ;
	output \g12858/_0_  ;
	output \g12859/_0_  ;
	output \g12861/_0_  ;
	output \g12862/_0_  ;
	output \g12868/_0_  ;
	output \g12869/_0_  ;
	output \g1287/_0_  ;
	output \g12870/_0_  ;
	output \g12871/_0_  ;
	output \g12872/_0_  ;
	output \g12873/_0_  ;
	output \g12874/_0_  ;
	output \g12875/_0_  ;
	output \g12876/_0_  ;
	output \g12877/_0_  ;
	output \g12878/_0_  ;
	output \g12879/_0_  ;
	output \g12880/_0_  ;
	output \g12881/_0_  ;
	output \g12882/_0_  ;
	output \g12883/_0_  ;
	output \g12884/_0_  ;
	output \g12885/_0_  ;
	output \g12886/_0_  ;
	output \g12887/_0_  ;
	output \g12888/_0_  ;
	output \g12889/_0_  ;
	output \g1289/_0_  ;
	output \g12890/_0_  ;
	output \g12891/_0_  ;
	output \g12894/_0_  ;
	output \g12898/_0_  ;
	output \g12899/_0_  ;
	output \g12900/_0_  ;
	output \g12901/_0_  ;
	output \g12902/_0_  ;
	output \g12903/_0_  ;
	output \g12906/_0_  ;
	output \g12907/_0_  ;
	output \g12908/_0_  ;
	output \g12912/_0_  ;
	output \g12913/_0_  ;
	output \g12914/_0_  ;
	output \g12915/_0_  ;
	output \g12916/_0_  ;
	output \g12917/_0_  ;
	output \g12918/_0_  ;
	output \g12919/_0_  ;
	output \g12920/_0_  ;
	output \g12921/_0_  ;
	output \g12922/_0_  ;
	output \g12923/_0_  ;
	output \g12924/_0_  ;
	output \g12925/_0_  ;
	output \g12926/_0_  ;
	output \g12932/_0_  ;
	output \g12933/_0_  ;
	output \g12936/_0_  ;
	output \g12955/_0_  ;
	output \g13015/_0_  ;
	output \g13016/_0_  ;
	output \g13017/_0_  ;
	output \g13018/_0_  ;
	output \g13019/_0_  ;
	output \g13020/_0_  ;
	output \g13021/_0_  ;
	output \g13024/_0_  ;
	output \g13025/_0_  ;
	output \g13027/_0_  ;
	output \g13028/_0_  ;
	output \g13030/_0_  ;
	output \g13031/_0_  ;
	output \g13033/_0_  ;
	output \g13047/_0_  ;
	output \g13060/_0_  ;
	output \g13062/_0_  ;
	output \g13063/_0_  ;
	output \g13064/_0_  ;
	output \g13067/_0_  ;
	output \g13068/_0_  ;
	output \g13069/_0_  ;
	output \g13070/_0_  ;
	output \g13072/_0_  ;
	output \g13094/_0_  ;
	output \g13104/_0_  ;
	output \g13110/_0_  ;
	output \g13114/_0_  ;
	output \g13115/_0_  ;
	output \g13116/_0_  ;
	output \g13117/_0_  ;
	output \g13118/_0_  ;
	output \g13119/_0_  ;
	output \g13120/_0_  ;
	output \g13121/_0_  ;
	output \g13124/_0_  ;
	output \g13125/_0_  ;
	output \g13127/_0_  ;
	output \g13128/_0_  ;
	output \g13129/_0_  ;
	output \g13130/_0_  ;
	output \g13131/_0_  ;
	output \g13132/_0_  ;
	output \g13133/_0_  ;
	output \g13134/_0_  ;
	output \g13138/_0_  ;
	output \g13139/_0_  ;
	output \g13140/_0_  ;
	output \g13141/_0_  ;
	output \g13142/_0_  ;
	output \g13143/_0_  ;
	output \g13144/_0_  ;
	output \g13146/_0_  ;
	output \g13150/_0_  ;
	output \g13152/_0_  ;
	output \g13154/_0_  ;
	output \g13155/_0_  ;
	output \g13156/_0_  ;
	output \g13157/_0_  ;
	output \g13158/_0_  ;
	output \g1320/_3_  ;
	output \g13266/_0_  ;
	output \g13269/_0_  ;
	output \g13274/_0_  ;
	output \g13277/_0_  ;
	output \g13280/_0_  ;
	output \g13283/_0_  ;
	output \g13294/_0_  ;
	output \g13330/_0_  ;
	output \g13333/_0_  ;
	output \g13334/_0_  ;
	output \g13335/_0_  ;
	output \g13336/_0_  ;
	output \g13337/_0_  ;
	output \g13338/_0_  ;
	output \g13345/_0_  ;
	output \g13346/_0_  ;
	output \g13347/_0_  ;
	output \g13348/_0_  ;
	output \g13349/_0_  ;
	output \g13350/_0_  ;
	output \g13351/_0_  ;
	output \g13352/_0_  ;
	output \g13486/_0_  ;
	output \g13488/_0_  ;
	output \g13508/_0_  ;
	output \g13509/_0_  ;
	output \g13510/_0_  ;
	output \g13511/_0_  ;
	output \g13512/_0_  ;
	output \g13513/_0_  ;
	output \g13514/_0_  ;
	output \g13515/_0_  ;
	output \g13516/_0_  ;
	output \g13517/_0_  ;
	output \g13518/_0_  ;
	output \g13519/_0_  ;
	output \g13520/_0_  ;
	output \g13521/_0_  ;
	output \g13540/_0_  ;
	output \g13541/_0_  ;
	output \g13542/_0_  ;
	output \g13543/_0_  ;
	output \g13544/_0_  ;
	output \g13545/_0_  ;
	output \g13546/_0_  ;
	output \g13547/_0_  ;
	output \g13548/_0_  ;
	output \g13549/_0_  ;
	output \g13550/_0_  ;
	output \g13551/_0_  ;
	output \g13552/_0_  ;
	output \g13553/_0_  ;
	output \g13554/_0_  ;
	output \g13555/_0_  ;
	output \g13556/_0_  ;
	output \g13557/_0_  ;
	output \g13558/_0_  ;
	output \g13559/_0_  ;
	output \g13560/_0_  ;
	output \g13561/_0_  ;
	output \g13562/_0_  ;
	output \g13563/_0_  ;
	output \g13564/_0_  ;
	output \g13565/_0_  ;
	output \g13566/_0_  ;
	output \g13567/_0_  ;
	output \g13568/_0_  ;
	output \g13569/_0_  ;
	output \g13570/_0_  ;
	output \g13571/_0_  ;
	output \g13572/_0_  ;
	output \g137/_3_  ;
	output \g1387/_3_  ;
	output \g1388/_3_  ;
	output \g1389/_0_  ;
	output \g139/_0_  ;
	output \g1390/_0_  ;
	output \g1393/_0_  ;
	output \g140/_0_  ;
	output \g141/_0_  ;
	output \g14173/_0_  ;
	output \g14176/_0_  ;
	output \g142/_3_  ;
	output \g14273/_1__syn_2  ;
	output \g14274/_0_  ;
	output \g14280/_0_  ;
	output \g14281/_0_  ;
	output \g143/_3_  ;
	output \g14354/_3__syn_2  ;
	output \g14370/_0_  ;
	output \g14385/_0_  ;
	output \g14386/_0_  ;
	output \g144/_3_  ;
	output \g14407/_0_  ;
	output \g14412/_0_  ;
	output \g14435/_0_  ;
	output \g14439/_0_  ;
	output \g145/_0_  ;
	output \g14522/_0_  ;
	output \g14528/_0_  ;
	output \g14533/_0_  ;
	output \g14581/_1_  ;
	output \g14582/_0_  ;
	output \g146/_3_  ;
	output \g14671/_0_  ;
	output \g14672/_0_  ;
	output \g147/_0_  ;
	output \g1473/_0_  ;
	output \g148/_0_  ;
	output \g14826/_0_  ;
	output \g149/_0_  ;
	output \g14908/_0_  ;
	output \g14911/_0_  ;
	output \g14936/_2_  ;
	output \g1494/_0_  ;
	output \g1495/_0_  ;
	output \g14950/_2_  ;
	output \g14953/_2_  ;
	output \g15003/_0_  ;
	output \g15004/_0_  ;
	output \g15006/_0_  ;
	output \g15007/_0_  ;
	output \g15008/_0_  ;
	output \g15009/_0_  ;
	output \g15010/_0_  ;
	output \g15011/_0_  ;
	output \g15012/_0_  ;
	output \g15013/_0_  ;
	output \g15014/_0_  ;
	output \g15015/_0_  ;
	output \g15016/_0_  ;
	output \g15017/_0_  ;
	output \g15018/_0_  ;
	output \g15019/_0_  ;
	output \g15035/_0_  ;
	output \g15036/_0_  ;
	output \g15038/_0_  ;
	output \g15039/_0_  ;
	output \g15040/_0_  ;
	output \g15041/_0_  ;
	output \g15042/_0_  ;
	output \g15043/_0_  ;
	output \g15044/_0_  ;
	output \g15045/_0_  ;
	output \g15046/_0_  ;
	output \g15056/_00_  ;
	output \g151/_0_  ;
	output \g15193/_0_  ;
	output \g152/_0_  ;
	output \g15256/_0_  ;
	output \g153/_0_  ;
	output \g15393/_0_  ;
	output \g15394/_0_  ;
	output \g15395/_0_  ;
	output \g15396/_0_  ;
	output \g15397/_0_  ;
	output \g15398/_0_  ;
	output \g15399/_0_  ;
	output \g154/_0_  ;
	output \g15400/_0_  ;
	output \g15401/_0_  ;
	output \g15402/_0_  ;
	output \g15403/_0_  ;
	output \g15404/_0_  ;
	output \g15405/_0_  ;
	output \g15406/_0_  ;
	output \g15407/_0_  ;
	output \g15408/_0_  ;
	output \g15473/_0_  ;
	output \g15650/_0_  ;
	output \g15651/_0_  ;
	output \g15652/_0_  ;
	output \g15653/_0_  ;
	output \g15662/_0_  ;
	output \g15663/_0_  ;
	output \g15664/_0_  ;
	output \g15665/_0_  ;
	output \g15666/_0_  ;
	output \g15667/_0_  ;
	output \g15668/_0_  ;
	output \g15669/_0_  ;
	output \g15670/_0_  ;
	output \g15671/_0_  ;
	output \g15672/_0_  ;
	output \g15673/_0_  ;
	output \g15674/_0_  ;
	output \g15675/_0_  ;
	output \g1569/_0_  ;
	output \g1570/_0_  ;
	output \g1575/_0_  ;
	output \g1576/_0_  ;
	output \g15922/_1_  ;
	output \g15970/_0_  ;
	output \g16059/_0_  ;
	output \g1606/_3_  ;
	output \g16124/_0_  ;
	output \g16144/_0_  ;
	output \g16202/_0_  ;
	output \g16214/_0_  ;
	output \g16247/_0_  ;
	output \g16257/_0_  ;
	output \g16274/_1_  ;
	output \g16324/_0_  ;
	output \g16343/_1__syn_2  ;
	output \g16381/_0_  ;
	output \g16383/_0_  ;
	output \g16386/_0_  ;
	output \g16414/_1__syn_2  ;
	output \g16416/_0__syn_2  ;
	output \g16448/_0_  ;
	output \g16460/_1_  ;
	output \g16625/_3_  ;
	output \g16662/_0_  ;
	output \g16668/_1__syn_2  ;
	output \g16692/_0_  ;
	output \g16721/_0_  ;
	output \g16723/_0_  ;
	output \g16725/_0_  ;
	output \g16726/_0_  ;
	output \g16727/_0_  ;
	output \g16728/_0_  ;
	output \g16729/_0_  ;
	output \g16730/_0_  ;
	output \g16731/_0_  ;
	output \g16732/_0_  ;
	output \g16733/_0_  ;
	output \g16734/_0_  ;
	output \g16735/_0_  ;
	output \g16736/_0_  ;
	output \g16737/_0_  ;
	output \g16738/_0_  ;
	output \g16739/_0_  ;
	output \g16740/_0_  ;
	output \g16741/_0_  ;
	output \g16742/_0_  ;
	output \g16743/_0_  ;
	output \g16747/_0_  ;
	output \g16748/_0_  ;
	output \g16749/_0_  ;
	output \g16750/_0_  ;
	output \g16753/_0_  ;
	output \g16754/_0_  ;
	output \g16755/_0_  ;
	output \g16756/_0_  ;
	output \g16757/_0_  ;
	output \g16758/_0_  ;
	output \g16761/_0_  ;
	output \g16765/_0_  ;
	output \g16766/_0_  ;
	output \g16767/_0_  ;
	output \g16768/_0_  ;
	output \g16769/_0_  ;
	output \g16772/_0_  ;
	output \g16785/_0_  ;
	output \g16786/_0_  ;
	output \g16787/_0_  ;
	output \g16788/_0_  ;
	output \g16789/_0_  ;
	output \g16790/_0_  ;
	output \g16791/_0_  ;
	output \g16804/_0_  ;
	output \g16805/_0_  ;
	output \g16806/_0_  ;
	output \g16807/_0_  ;
	output \g16808/_0_  ;
	output \g16809/_0_  ;
	output \g16810/_0_  ;
	output \g16811/_0_  ;
	output \g16812/_0_  ;
	output \g16813/_0_  ;
	output \g16814/_0_  ;
	output \g16815/_0_  ;
	output \g16816/_0_  ;
	output \g16817/_0_  ;
	output \g16819/_0_  ;
	output \g16822/_0_  ;
	output \g16823/_0_  ;
	output \g16824/_0_  ;
	output \g16825/_0_  ;
	output \g16828/_0_  ;
	output \g16829/_0_  ;
	output \g16830/_0_  ;
	output \g16831/_0_  ;
	output \g16832/_0_  ;
	output \g16833/_0_  ;
	output \g16834/_0_  ;
	output \g16835/_0_  ;
	output \g16836/_0_  ;
	output \g16837/_0_  ;
	output \g16840/_0_  ;
	output \g16841/_0_  ;
	output \g16842/_0_  ;
	output \g16843/_0_  ;
	output \g16846/_0_  ;
	output \g16847/_0_  ;
	output \g16848/_0_  ;
	output \g16849/_0_  ;
	output \g16850/_0_  ;
	output \g16851/_0_  ;
	output \g16852/_0_  ;
	output \g16853/_0_  ;
	output \g16854/_0_  ;
	output \g16855/_0_  ;
	output \g16856/_0_  ;
	output \g16857/_0_  ;
	output \g16859/_0_  ;
	output \g16862/_0_  ;
	output \g16865/_0_  ;
	output \g16866/_0_  ;
	output \g16867/_0_  ;
	output \g16868/_0_  ;
	output \g16869/_0_  ;
	output \g16870/_0_  ;
	output \g16871/_0_  ;
	output \g16872/_0_  ;
	output \g16873/_0_  ;
	output \g16874/_0_  ;
	output \g16875/_0_  ;
	output \g16876/_0_  ;
	output \g16877/_0_  ;
	output \g16878/_0_  ;
	output \g16879/_0_  ;
	output \g16880/_0_  ;
	output \g16881/_0_  ;
	output \g16882/_0_  ;
	output \g16884/_0_  ;
	output \g16887/_0_  ;
	output \g16891/_0_  ;
	output \g16892/_0_  ;
	output \g16893/_0_  ;
	output \g16894/_0_  ;
	output \g16895/_0_  ;
	output \g16897/_0_  ;
	output \g16898/_0_  ;
	output \g16899/_0_  ;
	output \g16900/_0_  ;
	output \g16901/_0_  ;
	output \g16902/_0_  ;
	output \g16903/_0_  ;
	output \g16904/_0_  ;
	output \g16905/_0_  ;
	output \g16906/_0_  ;
	output \g16907/_0_  ;
	output \g16908/_0_  ;
	output \g16909/_0_  ;
	output \g16910/_0_  ;
	output \g16912/_0_  ;
	output \g16914/_0_  ;
	output \g16915/_0_  ;
	output \g16950/_0_  ;
	output \g16951/_0_  ;
	output \g16952/_0_  ;
	output \g16953/_0_  ;
	output \g16954/_0_  ;
	output \g16955/_0_  ;
	output \g16956/_0_  ;
	output \g16957/_0_  ;
	output \g16958/_0_  ;
	output \g16959/_0_  ;
	output \g16960/_0_  ;
	output \g16961/_0_  ;
	output \g16962/_0_  ;
	output \g16963/_0_  ;
	output \g16964/_0_  ;
	output \g16965/_0_  ;
	output \g16966/_0_  ;
	output \g16967/_0_  ;
	output \g16968/_0_  ;
	output \g16970/_0_  ;
	output \g17102/_3_  ;
	output \g17106/_0_  ;
	output \g17107/_0_  ;
	output \g17109/_0_  ;
	output \g17110/_0_  ;
	output \g17111/_0_  ;
	output \g17112/_0_  ;
	output \g17115/_0_  ;
	output \g17116/_0_  ;
	output \g17119/_0_  ;
	output \g17120/_0_  ;
	output \g17122/_0_  ;
	output \g17123/_0_  ;
	output \g17124/_0_  ;
	output \g17125/_0_  ;
	output \g17126/_0_  ;
	output \g17127/_0_  ;
	output \g17128/_0_  ;
	output \g17130/_0_  ;
	output \g17131/_0_  ;
	output \g17132/_0_  ;
	output \g17133/_0_  ;
	output \g17134/_0_  ;
	output \g17135/_0_  ;
	output \g17136/_0_  ;
	output \g17137/_0_  ;
	output \g17138/_0_  ;
	output \g17140/_0_  ;
	output \g17141/_0_  ;
	output \g17142/_0_  ;
	output \g17143/_0_  ;
	output \g17144/_0_  ;
	output \g17145/_0_  ;
	output \g17146/_0_  ;
	output \g17147/_0_  ;
	output \g17148/_0_  ;
	output \g17149/_0_  ;
	output \g17150/_0_  ;
	output \g17151/_0_  ;
	output \g17152/_0_  ;
	output \g17153/_0_  ;
	output \g17154/_0_  ;
	output \g17155/_0_  ;
	output \g17157/_0_  ;
	output \g17159/_0_  ;
	output \g17160/_0_  ;
	output \g17161/_0_  ;
	output \g17162/_0_  ;
	output \g17163/_0_  ;
	output \g17164/_0_  ;
	output \g17165/_0_  ;
	output \g17166/_0_  ;
	output \g17168/_0_  ;
	output \g17171/_0_  ;
	output \g17173/_0_  ;
	output \g17177/_0_  ;
	output \g17178/_0_  ;
	output \g17179/_0_  ;
	output \g17180/_0_  ;
	output \g17182/_0_  ;
	output \g17183/_0_  ;
	output \g17184/_0_  ;
	output \g17185/_0_  ;
	output \g17186/_0_  ;
	output \g17188/_0_  ;
	output \g17189/_0_  ;
	output \g17190/_0_  ;
	output \g17191/_0_  ;
	output \g17193/_0_  ;
	output \g17194/_0_  ;
	output \g17195/_0_  ;
	output \g17196/_0_  ;
	output \g17197/_0_  ;
	output \g17198/_0_  ;
	output \g17199/_0_  ;
	output \g17200/_0_  ;
	output \g17201/_0_  ;
	output \g17202/_0_  ;
	output \g17203/_0_  ;
	output \g17204/_0_  ;
	output \g17205/_0_  ;
	output \g17206/_0_  ;
	output \g17207/_0_  ;
	output \g17208/_0_  ;
	output \g17209/_0_  ;
	output \g17210/_0_  ;
	output \g17211/_0_  ;
	output \g17212/_0_  ;
	output \g17213/_0_  ;
	output \g17214/_0_  ;
	output \g17215/_0_  ;
	output \g17216/_0_  ;
	output \g17217/_0_  ;
	output \g17218/_0_  ;
	output \g17219/_0_  ;
	output \g17223/_0_  ;
	output \g17224/_0_  ;
	output \g17225/_0_  ;
	output \g17226/_0_  ;
	output \g17227/_0_  ;
	output \g17228/_0_  ;
	output \g17229/_0_  ;
	output \g17231/_0_  ;
	output \g17232/_0_  ;
	output \g17233/_0_  ;
	output \g17234/_0_  ;
	output \g17237/_0_  ;
	output \g17239/_0_  ;
	output \g17240/_0_  ;
	output \g17243/_0_  ;
	output \g17246/_0_  ;
	output \g17247/_0_  ;
	output \g17248/_0_  ;
	output \g17249/_0_  ;
	output \g17250/_0_  ;
	output \g17251/_0_  ;
	output \g17252/_0_  ;
	output \g17253/_0_  ;
	output \g17254/_0_  ;
	output \g17258/_0_  ;
	output \g17261/_0_  ;
	output \g17262/_0_  ;
	output \g17269/_0_  ;
	output \g17271/_0_  ;
	output \g17274/_0_  ;
	output \g17275/_0_  ;
	output \g17276/_0_  ;
	output \g17277/_0_  ;
	output \g17278/_0_  ;
	output \g17279/_0_  ;
	output \g17280/_0_  ;
	output \g17281/_0_  ;
	output \g17282/_0_  ;
	output \g17283/_0_  ;
	output \g17285/_0_  ;
	output \g17290/_0_  ;
	output \g17292/_0_  ;
	output \g17293/_0_  ;
	output \g17296/_0_  ;
	output \g17297/_0_  ;
	output \g17298/_0_  ;
	output \g173/_0_  ;
	output \g17303/_0_  ;
	output \g17304/_0_  ;
	output \g17305/_0_  ;
	output \g17306/_0_  ;
	output \g17307/_0_  ;
	output \g17308/_0_  ;
	output \g17309/_0_  ;
	output \g17310/_0_  ;
	output \g17311/_0_  ;
	output \g17312/_0_  ;
	output \g17314/_0_  ;
	output \g17315/_0_  ;
	output \g17316/_0_  ;
	output \g17317/_0_  ;
	output \g17318/_0_  ;
	output \g17319/_0_  ;
	output \g17320/_0_  ;
	output \g17321/_0_  ;
	output \g17322/_0_  ;
	output \g17323/_0_  ;
	output \g17324/_0_  ;
	output \g17325/_0_  ;
	output \g17326/_0_  ;
	output \g17327/_0_  ;
	output \g17328/_0_  ;
	output \g17329/_0_  ;
	output \g17330/_0_  ;
	output \g17331/_0_  ;
	output \g17332/_0_  ;
	output \g17333/_0_  ;
	output \g17335/_0_  ;
	output \g17336/_0_  ;
	output \g17337/_0_  ;
	output \g17338/_0_  ;
	output \g17339/_0_  ;
	output \g17340/_0_  ;
	output \g17342/_0_  ;
	output \g17343/_0_  ;
	output \g17347/_0_  ;
	output \g17350/_0_  ;
	output \g17354/_0_  ;
	output \g17356/_0_  ;
	output \g17357/_0_  ;
	output \g17358/_0_  ;
	output \g17359/_0_  ;
	output \g17360/_0_  ;
	output \g17415/_0_  ;
	output \g17441/_0_  ;
	output \g17442/_0_  ;
	output \g17451/_0_  ;
	output \g17457/_0_  ;
	output \g17458/_0_  ;
	output \g17459/_0_  ;
	output \g17460/_0_  ;
	output \g17461/_0_  ;
	output \g17462/_0_  ;
	output \g17463/_0_  ;
	output \g17464/_0_  ;
	output \g17465/_0_  ;
	output \g17466/_0_  ;
	output \g17467/_0_  ;
	output \g17468/_0_  ;
	output \g17469/_0_  ;
	output \g17470/_0_  ;
	output \g17471/_0_  ;
	output \g17472/_0_  ;
	output \g175/_3_  ;
	output \g1750/_0_  ;
	output \g176/_3_  ;
	output \g17619/_0_  ;
	output \g17620/_0_  ;
	output \g1763/_3_  ;
	output \g1764/_3_  ;
	output \g1768/_0_  ;
	output \g1769/_0_  ;
	output \g177/_3_  ;
	output \g17737/_0_  ;
	output \g17747/_0_  ;
	output \g178/_3_  ;
	output \g17814/_1_  ;
	output \g17815/_0_  ;
	output \g17821/_1_  ;
	output \g17821/_1__syn_2  ;
	output \g17872/_0_  ;
	output \g179/_3_  ;
	output \g17902/_0_  ;
	output \g180/_3_  ;
	output \g18020/_1_  ;
	output \g18057/_0_  ;
	output \g18096/_0_  ;
	output \g18099/_0_  ;
	output \g18107/_0_  ;
	output \g18133/_0_  ;
	output \g18140/_1_  ;
	output \g18153/_0_  ;
	output \g182/_0_  ;
	output \g18218/_0_  ;
	output \g18244/_0_  ;
	output \g18262/_0_  ;
	output \g18267/_0_  ;
	output \g18387/_1__syn_2  ;
	output \g184/_0_  ;
	output \g18478/_1_  ;
	output \g18585/_3_  ;
	output \g18608/_0_  ;
	output \g18609/_0_  ;
	output \g18613/_0_  ;
	output \g18618/_0_  ;
	output \g18647/_0_  ;
	output \g18687/_2_  ;
	output \g18707/_0_  ;
	output \g18748/_0_  ;
	output \g18753/_0_  ;
	output \g18758/_0_  ;
	output \g18759/_0_  ;
	output \g18760/_0_  ;
	output \g18761/_0_  ;
	output \g18762/_0_  ;
	output \g18763/_0_  ;
	output \g18764/_0_  ;
	output \g18765/_0_  ;
	output \g18766/_0_  ;
	output \g18767/_0_  ;
	output \g18768/_0_  ;
	output \g18770/_0_  ;
	output \g18771/_0_  ;
	output \g18788/_0_  ;
	output \g18796/_0_  ;
	output \g18800/_0_  ;
	output \g18801/_0_  ;
	output \g18802/_0_  ;
	output \g18803/_0_  ;
	output \g18804/_0_  ;
	output \g18805/_0_  ;
	output \g18807/_0_  ;
	output \g18840/_0_  ;
	output \g18843/_0_  ;
	output \g18844/_0_  ;
	output \g18846/_0_  ;
	output \g18847/_0_  ;
	output \g18848/_0_  ;
	output \g18849/_0_  ;
	output \g18850/_0_  ;
	output \g18851/_0_  ;
	output \g18852/_0_  ;
	output \g18853/_0_  ;
	output \g18854/_0_  ;
	output \g18855/_0_  ;
	output \g18856/_0_  ;
	output \g18858/_0_  ;
	output \g18860/_0_  ;
	output \g18861/_0_  ;
	output \g18863/_0_  ;
	output \g18864/_0_  ;
	output \g18866/_0_  ;
	output \g18867/_0_  ;
	output \g18868/_0_  ;
	output \g18869/_0_  ;
	output \g18870/_0_  ;
	output \g18871/_0_  ;
	output \g18872/_0_  ;
	output \g18873/_0_  ;
	output \g18874/_0_  ;
	output \g18875/_0_  ;
	output \g18876/_0_  ;
	output \g18877/_0_  ;
	output \g18878/_0_  ;
	output \g18879/_0_  ;
	output \g18880/_0_  ;
	output \g18881/_0_  ;
	output \g18882/_0_  ;
	output \g18883/_0_  ;
	output \g18888/_0_  ;
	output \g18892/_0_  ;
	output \g18895/_0_  ;
	output \g18896/_0_  ;
	output \g18897/_0_  ;
	output \g18905/_0_  ;
	output \g18908/_0_  ;
	output \g18909/_0_  ;
	output \g18912/_0_  ;
	output \g18918/_0_  ;
	output \g18919/_0_  ;
	output \g18920/_0_  ;
	output \g18921/_0_  ;
	output \g18922/_0_  ;
	output \g18924/_0_  ;
	output \g18925/_0_  ;
	output \g18927/_0_  ;
	output \g18930/_0_  ;
	output \g18966/_0_  ;
	output \g18968/_0_  ;
	output \g18970/_0_  ;
	output \g18974/_0_  ;
	output \g18975/_0_  ;
	output \g18977/_0_  ;
	output \g18981/_0_  ;
	output \g18983/_0_  ;
	output \g18985/_0_  ;
	output \g18987/_0_  ;
	output \g18989/_0_  ;
	output \g18991/_0_  ;
	output \g18992/_0_  ;
	output \g18993/_0_  ;
	output \g18994/_0_  ;
	output \g18995/_0_  ;
	output \g18996/_0_  ;
	output \g18997/_0_  ;
	output \g18998/_0_  ;
	output \g18999/_0_  ;
	output \g19001/_0_  ;
	output \g19003/_0_  ;
	output \g19005/_0_  ;
	output \g19006/_0_  ;
	output \g19014/_0_  ;
	output \g19016/_0_  ;
	output \g19018/_0_  ;
	output \g19020/_0_  ;
	output \g19022/_0_  ;
	output \g19056/_3_  ;
	output \g19058/_3_  ;
	output \g19060/_3_  ;
	output \g19062/_3_  ;
	output \g1910/_0_  ;
	output \g19186/_0_  ;
	output \g19188/_0_  ;
	output \g19235/_0_  ;
	output \g19239/_0_  ;
	output \g19244/_0_  ;
	output \g19253/_0_  ;
	output \g19254/_0_  ;
	output \g19259/_0_  ;
	output \g19261/_0_  ;
	output \g19267/_0_  ;
	output \g19277/_0_  ;
	output \g19278/_0_  ;
	output \g19280/_0_  ;
	output \g19281/_0_  ;
	output \g19282/_0_  ;
	output \g19283/_0_  ;
	output \g19284/_0_  ;
	output \g19285/_0_  ;
	output \g19286/_0_  ;
	output \g19287/_0_  ;
	output \g19288/_0_  ;
	output \g19289/_0_  ;
	output \g19290/_0_  ;
	output \g19291/_0_  ;
	output \g19292/_0_  ;
	output \g19293/_0_  ;
	output \g19294/_0_  ;
	output \g19295/_0_  ;
	output \g19296/_0_  ;
	output \g19297/_0_  ;
	output \g19298/_0_  ;
	output \g19299/_0_  ;
	output \g19300/_0_  ;
	output \g19301/_0_  ;
	output \g19302/_0_  ;
	output \g19303/_0_  ;
	output \g19304/_0_  ;
	output \g19305/_0_  ;
	output \g19306/_0_  ;
	output \g19307/_0_  ;
	output \g19308/_0_  ;
	output \g19315/_0_  ;
	output \g19316/_0_  ;
	output \g19317/_0_  ;
	output \g19318/_0_  ;
	output \g19319/_0_  ;
	output \g19320/_0_  ;
	output \g19321/_0_  ;
	output \g19322/_0_  ;
	output \g19323/_0_  ;
	output \g19325/_3_  ;
	output \g19326/_3_  ;
	output \g19333/_3_  ;
	output \g19341/_3_  ;
	output \g19347/_3_  ;
	output \g19377/_3_  ;
	output \g19381/_3_  ;
	output \g19393/_0_  ;
	output \g19401/_0_  ;
	output \g19402/_0_  ;
	output \g195/_2_  ;
	output \g19513/_0_  ;
	output \g19514/_0_  ;
	output \g19515/_0_  ;
	output \g19516/_0_  ;
	output \g1952/_3_  ;
	output \g19529/_0_  ;
	output \g19530/_0_  ;
	output \g19531/_0_  ;
	output \g19532/_0_  ;
	output \g19533/_0_  ;
	output \g19534/_0_  ;
	output \g19535/_0_  ;
	output \g19536/_0_  ;
	output \g19537/_0_  ;
	output \g19539/_0_  ;
	output \g19546/_0_  ;
	output \g19552/_0_  ;
	output \g19553/_0_  ;
	output \g19562/_0_  ;
	output \g19563/_0_  ;
	output \g19564/_0_  ;
	output \g19572/_0_  ;
	output \g19575/_0_  ;
	output \g19615/_0_  ;
	output \g19686/_0_  ;
	output \g19688/_0_  ;
	output \g197/_0_  ;
	output \g19729/_0_  ;
	output \g19774/_0_  ;
	output \g19777/_0_  ;
	output \g19791/_0_  ;
	output \g19818/_0_  ;
	output \g19819/_0_  ;
	output \g19828/_0_  ;
	output \g19852/_1_  ;
	output \g19860/_0_  ;
	output \g19861/_0_  ;
	output \g19864/_0_  ;
	output \g19886/_0_  ;
	output \g19887/_0_  ;
	output \g199/_0_  ;
	output \g19908/_0_  ;
	output \g19918/_0_  ;
	output \g19927/_0_  ;
	output \g19933/_0_  ;
	output \g200/_0_  ;
	output \g20019/_0_  ;
	output \g20046/_0_  ;
	output \g20068/_1_  ;
	output \g20080/_1_  ;
	output \g201/_0_  ;
	output \g20137/_0_  ;
	output \g20139/_0_  ;
	output \g20141/_0_  ;
	output \g20152/_1_  ;
	output \g20154/_00_  ;
	output \g202/_0_  ;
	output \g20206/_0_  ;
	output \g20211/_2_  ;
	output \g20217/_2_  ;
	output \g20239/_0_  ;
	output \g20265/_2_  ;
	output \g20266/_0_  ;
	output \g20272/_2_  ;
	output \g20278/_2_  ;
	output \g20283/_0_  ;
	output \g20285/_2_  ;
	output \g20288/_2__syn_2  ;
	output \g20293/_0_  ;
	output \g20295/_2_  ;
	output \g203/_0_  ;
	output \g20302/_2_  ;
	output \g20303/_2_  ;
	output \g20304/_2_  ;
	output \g20311/_2_  ;
	output \g20326/_0_  ;
	output \g20330/_0_  ;
	output \g2034/_0_  ;
	output \g20345/_0_  ;
	output \g20346/_0_  ;
	output \g2035/_0_  ;
	output \g20363/_0_  ;
	output \g20364/_0_  ;
	output \g204/_0_  ;
	output \g2047/_0_  ;
	output \g20483/_0_  ;
	output \g20493/_00_  ;
	output \g205/_0_  ;
	output \g20569/_0_  ;
	output \g20570/_0_  ;
	output \g20571/_0_  ;
	output \g206/_0_  ;
	output \g20613/_0_  ;
	output \g20615/_0_  ;
	output \g20657/_1__syn_2  ;
	output \g20660/_0_  ;
	output \g20685/_0_  ;
	output \g207/_0_  ;
	output \g20713/_1_  ;
	output \g20747/_1_  ;
	output \g20784/_0_  ;
	output \g20820/_1_  ;
	output \g20859/_0_  ;
	output \g20873/_2_  ;
	output \g20886/_0_  ;
	output \g20887/_0_  ;
	output \g20891/_2__syn_2  ;
	output \g20907/_2_  ;
	output \g20936/_2__syn_2  ;
	output \g20937/_1_  ;
	output \g20955/_0_  ;
	output \g20959/_2__syn_2  ;
	output \g20967/_0_  ;
	output \g20971/_2__syn_2  ;
	output \g20974/_1__syn_2  ;
	output \g21015/_1_  ;
	output \g21051/_2_  ;
	output \g21079/_1_  ;
	output \g21081/_1_  ;
	output \g21087/_2__syn_2  ;
	output \g21114/_1_  ;
	output \g21116/_1_  ;
	output \g21120/_2__syn_2  ;
	output \g21147/_0_  ;
	output \g21179/_1_  ;
	output \g21185/_1_  ;
	output \g21223/_0_  ;
	output \g21242/_0_  ;
	output \g21253/_0_  ;
	output \g21257/_0_  ;
	output \g21323/_1_  ;
	output \g21324/_1_  ;
	output \g21366/_0_  ;
	output \g21385/_2_  ;
	output \g21464/_0_  ;
	output \g21475/_3_  ;
	output \g21481/_0_  ;
	output \g21482/_0_  ;
	output \g21494/_3_  ;
	output \g21500/_3_  ;
	output \g21507/_3_  ;
	output \g21511/_3_  ;
	output \g21537/_1_  ;
	output \g21568/_0_  ;
	output \g21591/_0_  ;
	output \g21604/_0_  ;
	output \g21605/_3_  ;
	output \g21606/_0_  ;
	output \g21607/_0_  ;
	output \g21608/_0_  ;
	output \g21609/_0_  ;
	output \g21610/_0_  ;
	output \g21611/_0_  ;
	output \g21612/_0_  ;
	output \g21613/_0_  ;
	output \g21614/_0_  ;
	output \g21615/_0_  ;
	output \g21616/_0_  ;
	output \g21617/_0_  ;
	output \g21618/_0_  ;
	output \g21621/_0_  ;
	output \g21640/_0_  ;
	output \g21678/_0_  ;
	output \g21679/_0_  ;
	output \g21686/_0_  ;
	output \g21692/_3_  ;
	output \g21696/_0_  ;
	output \g21698/_0_  ;
	output \g21702/_3_  ;
	output \g21707/_0_  ;
	output \g21709/_0_  ;
	output \g21728/_0_  ;
	output \g21729/_0_  ;
	output \g21731/_0_  ;
	output \g21732/_0_  ;
	output \g21733/_0_  ;
	output \g21736/_0_  ;
	output \g21744/_3_  ;
	output \g21753/_0_  ;
	output \g21754/_0_  ;
	output \g21755/_0_  ;
	output \g21756/_0_  ;
	output \g21757/_0_  ;
	output \g21759/_0_  ;
	output \g21761/_0_  ;
	output \g21763/_0_  ;
	output \g21764/_0_  ;
	output \g21766/_0_  ;
	output \g2180/_0_  ;
	output \g21853/_3_  ;
	output \g21861/_3_  ;
	output \g21863/_3_  ;
	output \g21869/_3_  ;
	output \g2187/_0_  ;
	output \g21875/_3_  ;
	output \g21877/_3_  ;
	output \g21879/_3_  ;
	output \g2188/_0_  ;
	output \g21900/_0_  ;
	output \g22080/_0_  ;
	output \g22082/_0_  ;
	output \g22135/_0_  ;
	output \g22145/_1_  ;
	output \g22225/_0_  ;
	output \g223/_0_  ;
	output \g22354/_0_  ;
	output \g224/_0_  ;
	output \g22412/_0_  ;
	output \g22415/_1__syn_2  ;
	output \g225/_0_  ;
	output \g2257/_0_  ;
	output \g226/_3_  ;
	output \g22624/_0_  ;
	output \g227/_3_  ;
	output \g22702/_0_  ;
	output \g22919/_1__syn_2  ;
	output \g22933/_0_  ;
	output \g22954/_0_  ;
	output \g22989/_1_  ;
	output \g23529/_0_  ;
	output \g23539/_0_  ;
	output \g2362/_2_  ;
	output \g23766/_0_  ;
	output \g24/_3_  ;
	output \g24018/_0_  ;
	output \g2416/_0_  ;
	output \g2420/_0_  ;
	output \g24213/_0_  ;
	output \g24301/_0_  ;
	output \g2479/_0_  ;
	output \g248/_3_  ;
	output \g2480/_0_  ;
	output \g2481/_0_  ;
	output \g2482/_0_  ;
	output \g2483/_0_  ;
	output \g2484/_0_  ;
	output \g2485/_0_  ;
	output \g2486/_0_  ;
	output \g2487/_0_  ;
	output \g2488/_0_  ;
	output \g249/_3_  ;
	output \g2490/_0_  ;
	output \g2491/_0_  ;
	output \g2492/_0_  ;
	output \g2493/_0_  ;
	output \g2494/_0_  ;
	output \g2495/_0_  ;
	output \g2496/_0_  ;
	output \g2497/_0_  ;
	output \g2507/_0_  ;
	output \g2508/_0_  ;
	output \g2509/_0_  ;
	output \g2510/_0_  ;
	output \g2511/_0_  ;
	output \g2512/_0_  ;
	output \g2513/_0_  ;
	output \g2514/_0_  ;
	output \g2515/_0_  ;
	output \g2516/_0_  ;
	output \g25237/_0_  ;
	output \g2558/_0_  ;
	output \g2562/_0_  ;
	output \g2563/_0_  ;
	output \g2564/_0_  ;
	output \g2565/_0_  ;
	output \g2566/_0_  ;
	output \g2567/_0_  ;
	output \g2699/_0_  ;
	output \g27/_2_  ;
	output \g271/_0_  ;
	output \g272/_3_  ;
	output \g273/_3_  ;
	output \g274/_3_  ;
	output \g275/_3_  ;
	output \g276/_3_  ;
	output \g277/_3_  ;
	output \g2787/_3_  ;
	output \g2788/_3_  ;
	output \g279/_0_  ;
	output \g2795/_0_  ;
	output \g2796/_0_  ;
	output \g280/_0_  ;
	output \g2842/_3_  ;
	output \g29/_1_  ;
	output \g2927/_0_  ;
	output \g2978/_0_  ;
	output \g2979/_0_  ;
	output \g2980/_0_  ;
	output \g2981/_0_  ;
	output \g2982/_0_  ;
	output \g2983/_0_  ;
	output \g2984/_0_  ;
	output \g2985/_0_  ;
	output \g3021/_3_  ;
	output \g3022/_3_  ;
	output \g3023/_3_  ;
	output \g3024/_3_  ;
	output \g3025/_3_  ;
	output \g3026/_3_  ;
	output \g3027/_3_  ;
	output \g3028/_3_  ;
	output \g3029/_3_  ;
	output \g3030/_3_  ;
	output \g3031/_3_  ;
	output \g3032/_3_  ;
	output \g3033/_3_  ;
	output \g3034/_3_  ;
	output \g3035/_3_  ;
	output \g3036/_3_  ;
	output \g3037/_3_  ;
	output \g3038/_3_  ;
	output \g3039/_3_  ;
	output \g3040/_3_  ;
	output \g3041/_3_  ;
	output \g3042/_3_  ;
	output \g3049/_0_  ;
	output \g3050/_0_  ;
	output \g3051/_0_  ;
	output \g3052/_0_  ;
	output \g3053/_0_  ;
	output \g3054/_0_  ;
	output \g3058/_0_  ;
	output \g3059/_0_  ;
	output \g3088/_0_  ;
	output \g3089/_0_  ;
	output \g3090/_0_  ;
	output \g3091/_0_  ;
	output \g3092/_0_  ;
	output \g3093/_0_  ;
	output \g3094/_0_  ;
	output \g3095/_0_  ;
	output \g314/_0_  ;
	output \g3147/_3_  ;
	output \g3148/_3_  ;
	output \g3189/_0_  ;
	output \g3190/_0_  ;
	output \g3191/_0_  ;
	output \g3192/_0_  ;
	output \g3193/_0_  ;
	output \g3194/_0_  ;
	output \g3195/_0_  ;
	output \g3196/_0_  ;
	output \g3197/_0_  ;
	output \g3198/_0_  ;
	output \g3199/_0_  ;
	output \g32/_0_  ;
	output \g320/_3_  ;
	output \g3200/_0_  ;
	output \g3201/_0_  ;
	output \g3202/_0_  ;
	output \g3203/_0_  ;
	output \g3204/_0_  ;
	output \g321/_3_  ;
	output \g325/_3_  ;
	output \g3271/_2_  ;
	output \g33/_0_  ;
	output \g3363/_0_  ;
	output \g3413/_0_  ;
	output \g3414/_0_  ;
	output \g352/_0_  ;
	output \g355/_0_  ;
	output \g356/_3_  ;
	output \g357/_3_  ;
	output \g35_dup/_1_  ;
	output \g36/_3_  ;
	output \g365/_3_  ;
	output \g366/_3_  ;
	output \g367/_3_  ;
	output \g368/_3_  ;
	output \g3687/_0_  ;
	output \g369/_3_  ;
	output \g37/_3_  ;
	output \g370/_3_  ;
	output \g372/_3_  ;
	output \g374/_3_  ;
	output \g3740/_0_  ;
	output \g375/_3_  ;
	output \g376/_3_  ;
	output \g3878/_0_  ;
	output \g3879/_0_  ;
	output \g388/_3_  ;
	output \g3880/_0_  ;
	output \g3881/_0_  ;
	output \g3882/_0_  ;
	output \g389/_3_  ;
	output \g3894/_0_  ;
	output \g3895/_0_  ;
	output \g3896/_0_  ;
	output \g3897/_0_  ;
	output \g3898/_0_  ;
	output \g392/_3_  ;
	output \g393/_3_  ;
	output \g394/_3_  ;
	output \g395/_3_  ;
	output \g396/_3_  ;
	output \g397/_3_  ;
	output \g398/_3_  ;
	output \g399/_3_  ;
	output \g401/_3_  ;
	output \g402/_3_  ;
	output \g404/_3_  ;
	output \g4048/_0_  ;
	output \g405/_3_  ;
	output \g4050/_0_  ;
	output \g406/_3_  ;
	output \g407/_3_  ;
	output \g410/_3_  ;
	output \g411/_3_  ;
	output \g412/_3_  ;
	output \g413/_3_  ;
	output \g415/_3_  ;
	output \g416/_3_  ;
	output \g42/_0_  ;
	output \g4216/_3_  ;
	output \g4217/_3_  ;
	output \g4218/_3_  ;
	output \g4219/_3_  ;
	output \g4296/_0_  ;
	output \g4297/_0_  ;
	output \g4298/_0_  ;
	output \g4299/_0_  ;
	output \g43/_0_  ;
	output \g4300/_0_  ;
	output \g4301/_0_  ;
	output \g4302/_0_  ;
	output \g4303/_0_  ;
	output \g4304/_0_  ;
	output \g4305/_0_  ;
	output \g4306/_0_  ;
	output \g4307/_0_  ;
	output \g4308/_0_  ;
	output \g4309/_0_  ;
	output \g4310/_0_  ;
	output \g4311/_0_  ;
	output \g4312/_0_  ;
	output \g4313/_0_  ;
	output \g4314/_0_  ;
	output \g4315/_0_  ;
	output \g4316/_0_  ;
	output \g4317/_0_  ;
	output \g4318/_0_  ;
	output \g4319/_0_  ;
	output \g4320/_0_  ;
	output \g4321/_0_  ;
	output \g4322/_0_  ;
	output \g4323/_0_  ;
	output \g436/_0_  ;
	output \g44/_0_  ;
	output \g448/_3_  ;
	output \g45/_0_  ;
	output \g4587/_0_  ;
	output \g4588/_0_  ;
	output \g46/_0_  ;
	output \g4601/_0_  ;
	output \g4602/_0_  ;
	output \g4613/_3_  ;
	output \g4614/_3_  ;
	output \g4615/_3_  ;
	output \g463/_0_  ;
	output \g465/_0_  ;
	output \g4653/_0_  ;
	output \g4654/_0_  ;
	output \g4655/_0_  ;
	output \g4656/_0_  ;
	output \g4659/_0_  ;
	output \g466/_0_  ;
	output \g468/_3_  ;
	output \g469/_3_  ;
	output \g4697/_0_  ;
	output \g47/_3_  ;
	output \g470/_0_  ;
	output \g471/_0_  ;
	output \g4755/_0_  ;
	output \g476/_0_  ;
	output \g48/_3_  ;
	output \g480/_00_  ;
	output \g4839/_0_  ;
	output \g4840/_0_  ;
	output \g485/_3_  ;
	output \g4854/_0_  ;
	output \g4855/_0_  ;
	output \g4859/_0_  ;
	output \g486/_3_  ;
	output \g4860/_0_  ;
	output \g4880/_0_  ;
	output \g4881/_0_  ;
	output \g4882/_0_  ;
	output \g4883/_0_  ;
	output \g4884/_0_  ;
	output \g4885/_0_  ;
	output \g4886/_0_  ;
	output \g4887/_0_  ;
	output \g4888/_0_  ;
	output \g49/_0_  ;
	output \g494/_0_  ;
	output \g499/_1_  ;
	output \g50/_0_  ;
	output \g5002/_0_  ;
	output \g5003/_0_  ;
	output \g5009/_0_  ;
	output \g5010/_0_  ;
	output \g5011/_0_  ;
	output \g5014/_0_  ;
	output \g51/_0_  ;
	output \g5105/_0_  ;
	output \g5129/_2_  ;
	output \g5132/_0_  ;
	output \g5135/_0_  ;
	output \g5168/_0_  ;
	output \g5169/_0_  ;
	output \g5173/_0_  ;
	output \g5224/_0_  ;
	output \g5225/_0_  ;
	output \g5226/_0_  ;
	output \g5227/_0_  ;
	output \g5334/_0_  ;
	output \g5335/_0_  ;
	output \g5336/_0_  ;
	output \g5337/_0_  ;
	output \g5338/_0_  ;
	output \g5339/_0_  ;
	output \g5340/_0_  ;
	output \g5341/_0_  ;
	output \g5342/_0_  ;
	output \g5343/_0_  ;
	output \g5344/_0_  ;
	output \g5345/_0_  ;
	output \g5346/_0_  ;
	output \g5347/_0_  ;
	output \g5348/_0_  ;
	output \g5349/_0_  ;
	output \g5395/_0_  ;
	output \g54/_0_  ;
	output \g5434/_0_  ;
	output \g5447/_0_  ;
	output \g5450/_0_  ;
	output \g5451/_0_  ;
	output \g5452/_0_  ;
	output \g5453/_0_  ;
	output \g5454/_0_  ;
	output \g5461/_0_  ;
	output \g5483/_0_  ;
	output \g5484/_0_  ;
	output \g5492/_0_  ;
	output \g5493/_0_  ;
	output \g5496/_3_  ;
	output \g5497/_3_  ;
	output \g55/_0_  ;
	output \g5500/_0_  ;
	output \g5502/_0_  ;
	output \g5503/_0_  ;
	output \g5506/_0_  ;
	output \g5511/_0_  ;
	output \g5518/_0_  ;
	output \g5519/_0_  ;
	output \g5520/_0_  ;
	output \g5522/_0_  ;
	output \g5523/_0_  ;
	output \g5524/_0_  ;
	output \g5525/_0_  ;
	output \g5532/_0_  ;
	output \g5533/_0_  ;
	output \g5534/_0_  ;
	output \g5535/_0_  ;
	output \g5536/_0_  ;
	output \g5537/_0_  ;
	output \g5538/_0_  ;
	output \g5546/_0_  ;
	output \g5555/_00_  ;
	output \g5593/_0_  ;
	output \g5614/_2_  ;
	output \g567/_0_  ;
	output \g5677/_0_  ;
	output \g5678/_0_  ;
	output \g5682/_0_  ;
	output \g5683/_0_  ;
	output \g5684/_0_  ;
	output \g5686/_0_  ;
	output \g5687/_0_  ;
	output \g5689/_0_  ;
	output \g5690/_0_  ;
	output \g5691/_0_  ;
	output \g5692/_0_  ;
	output \g5698/_0_  ;
	output \g5699/_0_  ;
	output \g5700/_0_  ;
	output \g5701/_0_  ;
	output \g5702/_0_  ;
	output \g5703/_0_  ;
	output \g5704/_0_  ;
	output \g5709/_0_  ;
	output \g5711/_0_  ;
	output \g5714/_0_  ;
	output \g572/_0_  ;
	output \g5723/_0_  ;
	output \g5724/_0_  ;
	output \g5725/_0_  ;
	output \g573/_0_  ;
	output \g5739/_0_  ;
	output \g5740/_0_  ;
	output \g575/_0_  ;
	output \g5756/_0_  ;
	output \g5757/_0_  ;
	output \g5758/_0_  ;
	output \g5759/_0_  ;
	output \g576/_0_  ;
	output \g5760/_0_  ;
	output \g5761/_0_  ;
	output \g5762/_0_  ;
	output \g5763/_0_  ;
	output \g577/_0_  ;
	output \g5772/_0_  ;
	output \g5773/_0_  ;
	output \g5774/_0_  ;
	output \g5775/_0_  ;
	output \g5776/_0_  ;
	output \g5777/_0_  ;
	output \g578/_0_  ;
	output \g5781/_0_  ;
	output \g5783/_0_  ;
	output \g5784/_0_  ;
	output \g5785/_0_  ;
	output \g5786/_0_  ;
	output \g5787/_0_  ;
	output \g5788/_0_  ;
	output \g5789/_0_  ;
	output \g579/_0_  ;
	output \g5790/_0_  ;
	output \g5791/_0_  ;
	output \g5792/_0_  ;
	output \g5794/_0_  ;
	output \g5795/_0_  ;
	output \g5796/_0_  ;
	output \g580/_0_  ;
	output \g5801/_0_  ;
	output \g5802/_0_  ;
	output \g5803/_0_  ;
	output \g5804/_0_  ;
	output \g5805/_0_  ;
	output \g581/_0_  ;
	output \g5814/_0_  ;
	output \g582/_0_  ;
	output \g583/_0_  ;
	output \g5849/_3_  ;
	output \g585/_0_  ;
	output \g586/_0_  ;
	output \g587/_0_  ;
	output \g588/_0_  ;
	output \g589/_0_  ;
	output \g590/_0_  ;
	output \g591/_0_  ;
	output \g592/_0_  ;
	output \g593/_0_  ;
	output \g594/_0_  ;
	output \g595/_0_  ;
	output \g596/_0_  ;
	output \g597/_0_  ;
	output \g5971/_0_  ;
	output \g5972/_0_  ;
	output \g5976/_0_  ;
	output \g598/_0_  ;
	output \g5989/_0_  ;
	output \g599/_0_  ;
	output \g600/_0_  ;
	output \g601/_0_  ;
	output \g602/_0_  ;
	output \g603/_0_  ;
	output \g604/_0_  ;
	output \g605/_0_  ;
	output \g6092/_0_  ;
	output \g6093/_2_  ;
	output \g6094/_0_  ;
	output \g6114/_0_  ;
	output \g614/_3_  ;
	output \g6148/_0_  ;
	output \g6149/_0_  ;
	output \g6171/_0_  ;
	output \g6172/_0_  ;
	output \g6173/_0_  ;
	output \g6174/_0_  ;
	output \g6175/_0_  ;
	output \g6176/_0_  ;
	output \g6177/_0_  ;
	output \g6178/_0_  ;
	output \g6179/_0_  ;
	output \g6180/_0_  ;
	output \g6181/_0_  ;
	output \g6182/_0_  ;
	output \g6183/_0_  ;
	output \g6184/_0_  ;
	output \g6185/_0_  ;
	output \g6186/_0_  ;
	output \g6187/_0_  ;
	output \g6193/_0_  ;
	output \g6196/_0_  ;
	output \g6197/_0_  ;
	output \g6198/_3_  ;
	output \g6200/_2_  ;
	output \g6202/_2_  ;
	output \g6203/_3_  ;
	output \g6204/_3_  ;
	output \g6209/_0_  ;
	output \g6211/_0_  ;
	output \g6215/_0_  ;
	output \g6217/_0_  ;
	output \g6219/_0_  ;
	output \g6220/_0_  ;
	output \g6222/_0_  ;
	output \g6224/_0_  ;
	output \g6228/_0_  ;
	output \g6238/_0_  ;
	output \g6239/_0_  ;
	output \g6240/_0_  ;
	output \g6242/_0_  ;
	output \g6243/_0_  ;
	output \g6244/_0_  ;
	output \g6245/_0_  ;
	output \g6246/_0_  ;
	output \g6248/_0_  ;
	output \g6249/_0_  ;
	output \g6259/_0_  ;
	output \g6260/_0_  ;
	output \g6261/_0_  ;
	output \g6262/_0_  ;
	output \g6263/_0_  ;
	output \g6264/_0_  ;
	output \g6265/_0_  ;
	output \g6266/_0_  ;
	output \g6267/_0_  ;
	output \g6268/_0_  ;
	output \g6269/_0_  ;
	output \g6270/_0_  ;
	output \g6271/_0_  ;
	output \g6272/_0_  ;
	output \g6277/_0_  ;
	output \g6318/_0_  ;
	output \g6326/_0_  ;
	output \g6329/_0_  ;
	output \g6330/_0_  ;
	output \g6331/_0_  ;
	output \g6332/_0_  ;
	output \g6333/_0_  ;
	output \g6334/_0_  ;
	output \g6335/_0_  ;
	output \g6336/_0_  ;
	output \g6337/_0_  ;
	output \g6338/_0_  ;
	output \g6339/_0_  ;
	output \g6340/_0_  ;
	output \g6341/_0_  ;
	output \g6342/_0_  ;
	output \g6343/_0_  ;
	output \g6344/_0_  ;
	output \g6345/_0_  ;
	output \g6346/_0_  ;
	output \g6347/_0_  ;
	output \g6348/_0_  ;
	output \g6349/_0_  ;
	output \g6350/_0_  ;
	output \g6351/_0_  ;
	output \g6352/_0_  ;
	output \g6353/_0_  ;
	output \g6354/_0_  ;
	output \g6355/_0_  ;
	output \g6361/_0_  ;
	output \g637/_0_  ;
	output \g638/_0_  ;
	output \g639/_3_  ;
	output \g64/_3_  ;
	output \g640/_3_  ;
	output \g6419/_0_  ;
	output \g6442/_0_  ;
	output \g6442/_1_  ;
	output \g6489/_0_  ;
	output \g6490/_0_  ;
	output \g65/_3_  ;
	output \g6513/_0_  ;
	output \g6515/_0_  ;
	output \g6571/_0_  ;
	output \g6588/_0_  ;
	output \g6589/_0_  ;
	output \g6638/_0_  ;
	output \g6639/_0_  ;
	output \g6653/_0_  ;
	output \g6654/_3_  ;
	output \g6655/_0_  ;
	output \g6656/_0_  ;
	output \g6657/_0_  ;
	output \g6687/_0_  ;
	output \g6688/_0_  ;
	output \g6689/_0_  ;
	output \g6690/_0_  ;
	output \g6691/_0_  ;
	output \g6692/_0_  ;
	output \g6693/_0_  ;
	output \g6694/_0_  ;
	output \g6701/_0_  ;
	output \g6706/_0_  ;
	output \g6711/_0_  ;
	output \g6727/_0_  ;
	output \g6728/_0_  ;
	output \g6736/_0_  ;
	output \g6739/_0_  ;
	output \g6742/_0_  ;
	output \g6746/_0_  ;
	output \g6752/_0_  ;
	output \g6771/_0_  ;
	output \g684/_0_  ;
	output \g685/_0_  ;
	output \g686/_0_  ;
	output \g687/_0_  ;
	output \g688/_0_  ;
	output \g689/_0_  ;
	output \g690/_0_  ;
	output \g691/_0_  ;
	output \g692/_0_  ;
	output \g693/_0_  ;
	output \g696/_3_  ;
	output \g697/_3_  ;
	output \g699/_0_  ;
	output \g7/_0_  ;
	output \g700/_0_  ;
	output \g7005/_0_  ;
	output \g7056/_0_  ;
	output \g7057/_0_  ;
	output \g7058/_0_  ;
	output \g7060/_0_  ;
	output \g7075/_0_  ;
	output \g7086/_0_  ;
	output \g7087/_0_  ;
	output \g7089/_0_  ;
	output \g7108/_0_  ;
	output \g7109/_0_  ;
	output \g7112/_0_  ;
	output \g7172/_2_  ;
	output \g7210/_2_  ;
	output \g7211/_0_  ;
	output \g7212/_0_  ;
	output \g7213/_0_  ;
	output \g7214/_0_  ;
	output \g7215/_0_  ;
	output \g7216/_0_  ;
	output \g7217/_3_  ;
	output \g7218/_0_  ;
	output \g7219/_0_  ;
	output \g7220/_0_  ;
	output \g7222/_0_  ;
	output \g7227/_2_  ;
	output \g723/_3_  ;
	output \g7234/_0_  ;
	output \g7237/_3_  ;
	output \g7238/_3_  ;
	output \g7239/_3_  ;
	output \g724/_3_  ;
	output \g7240/_3_  ;
	output \g7241/_3_  ;
	output \g7242/_3_  ;
	output \g7243/_3_  ;
	output \g7244/_0_  ;
	output \g7245/_0_  ;
	output \g7246/_0_  ;
	output \g7247/_0_  ;
	output \g7248/_0_  ;
	output \g7249/_0_  ;
	output \g7250/_0_  ;
	output \g7251/_0_  ;
	output \g7253/_0_  ;
	output \g7254/_0_  ;
	output \g7255/_0_  ;
	output \g7256/_0_  ;
	output \g7257/_0_  ;
	output \g7258/_0_  ;
	output \g7261/_0_  ;
	output \g7264/_0_  ;
	output \g7265/_0_  ;
	output \g7266/_0_  ;
	output \g7267/_0_  ;
	output \g7268/_0_  ;
	output \g7269/_0_  ;
	output \g7278/_0_  ;
	output \g7279/_0_  ;
	output \g7280/_0_  ;
	output \g7281/_0_  ;
	output \g7282/_0_  ;
	output \g7283/_0_  ;
	output \g7284/_0_  ;
	output \g7285/_0_  ;
	output \g7286/_3_  ;
	output \g7288/_3_  ;
	output \g7291/_0_  ;
	output \g7296/_3_  ;
	output \g73/_0_  ;
	output \g7302/_3_  ;
	output \g7306/_3_  ;
	output \g7310/_3_  ;
	output \g7311/_3_  ;
	output \g7312/_3_  ;
	output \g7313/_3_  ;
	output \g7314/_3_  ;
	output \g7315/_3_  ;
	output \g7316/_3_  ;
	output \g7317/_3_  ;
	output \g7323/_3_  ;
	output \g7324/_3_  ;
	output \g7325/_3_  ;
	output \g7327/_0_  ;
	output \g7362/_0_  ;
	output \g74/_0_  ;
	output \g75/_0_  ;
	output \g7512/_0_  ;
	output \g7513/_0_  ;
	output \g7514/_0_  ;
	output \g7515/_0_  ;
	output \g7516/_0_  ;
	output \g7518/_0_  ;
	output \g7528/_0_  ;
	output \g7529/_0_  ;
	output \g7548/_0_  ;
	output \g7549/_0_  ;
	output \g7550/_0_  ;
	output \g7575/_0_  ;
	output \g7576/_0_  ;
	output \g7577/_0_  ;
	output \g7578/_0_  ;
	output \g7579/_0_  ;
	output \g7580/_0_  ;
	output \g7581/_0_  ;
	output \g7582/_0_  ;
	output \g7583/_0_  ;
	output \g7584/_0_  ;
	output \g7585/_0_  ;
	output \g7586/_0_  ;
	output \g7587/_0_  ;
	output \g7588/_0_  ;
	output \g7589/_0_  ;
	output \g7590/_0_  ;
	output \g7591/_0_  ;
	output \g7592/_0_  ;
	output \g7593/_0_  ;
	output \g7594/_0_  ;
	output \g7595/_0_  ;
	output \g7596/_0_  ;
	output \g7597/_0_  ;
	output \g7598/_0_  ;
	output \g7599/_0_  ;
	output \g76/_0_  ;
	output \g7600/_0_  ;
	output \g7601/_0_  ;
	output \g7602/_0_  ;
	output \g7603/_0_  ;
	output \g7604/_0_  ;
	output \g7614/_0_  ;
	output \g7618/_0_  ;
	output \g762/_0_  ;
	output \g7634/_0_  ;
	output \g766/_0_  ;
	output \g767/_0_  ;
	output \g768/_0_  ;
	output \g769/_0_  ;
	output \g77/_0_  ;
	output \g770/_3_  ;
	output \g771/_3_  ;
	output \g7715/_0_  ;
	output \g774/_0_  ;
	output \g7746/_0_  ;
	output \g7753/_0_  ;
	output \g7754/_0_  ;
	output \g7755/_0_  ;
	output \g7756/_0_  ;
	output \g7757/_0_  ;
	output \g7758/_0_  ;
	output \g7759/_0_  ;
	output \g7760/_0_  ;
	output \g7761/_0_  ;
	output \g7762/_0_  ;
	output \g7763/_0_  ;
	output \g7764/_0_  ;
	output \g7765/_0_  ;
	output \g7766/_0_  ;
	output \g7778/_0_  ;
	output \g7779/_0_  ;
	output \g7780/_0_  ;
	output \g7781/_0_  ;
	output \g7782/_0_  ;
	output \g7784/_0_  ;
	output \g78/_0_  ;
	output \g7800/_0_  ;
	output \g7823/_3_  ;
	output \g7837/_0_  ;
	output \g7841/_0_  ;
	output \g7842/_0_  ;
	output \g7843/_0_  ;
	output \g7844/_0_  ;
	output \g7845/_0_  ;
	output \g7846/_0_  ;
	output \g7847/_0_  ;
	output \g7849/_0_  ;
	output \g7850/_0_  ;
	output \g7852/_0_  ;
	output \g7854/_0_  ;
	output \g7855/_0_  ;
	output \g7857/_0_  ;
	output \g7858/_0_  ;
	output \g7859/_0_  ;
	output \g7860/_0_  ;
	output \g7861/_0_  ;
	output \g7862/_0_  ;
	output \g7863/_0_  ;
	output \g7864/_0_  ;
	output \g7865/_0_  ;
	output \g7866/_0_  ;
	output \g7867/_0_  ;
	output \g7868/_0_  ;
	output \g7869/_0_  ;
	output \g7870/_0_  ;
	output \g7871/_0_  ;
	output \g79211/_3_  ;
	output \g79258/_3_  ;
	output \g79299/_3_  ;
	output \g79316/_2_  ;
	output \g79342/_3_  ;
	output \g79401/_3_  ;
	output \g79452/_3_  ;
	output \g79457/_3_  ;
	output \g7951/_0_  ;
	output \g79541/_3_  ;
	output \g7958/_0_  ;
	output \g79598/_3_  ;
	output \g79654/_3_  ;
	output \g79675/_3_  ;
	output \g7971/_0_  ;
	output \g7972/_0_  ;
	output \g7973/_3_  ;
	output \g79753/_3_  ;
	output \g7976/_3_  ;
	output \g79855/_3_  ;
	output \g79858/_3_  ;
	output \g79997/_3_  ;
	output \g8/_0_  ;
	output \g80008/_3_  ;
	output \g80011/_0_  ;
	output \g80104/_0_  ;
	output \g80172/_1_  ;
	output \g80195/_3_  ;
	output \g80238/_3_  ;
	output \g80290/_2_  ;
	output \g80294/_0_  ;
	output \g80302/_0_  ;
	output \g80327/_0_  ;
	output \g80360/_3_  ;
	output \g80373/_0_  ;
	output \g80401/_0_  ;
	output \g80410/_0_  ;
	output \g80475/_0_  ;
	output \g80476/_0_  ;
	output \g80516/_3_  ;
	output \g80536/_0_  ;
	output \g80537/_0_  ;
	output \g80572/_0_  ;
	output \g80573/_0_  ;
	output \g80609/_2_  ;
	output \g80610/_2_  ;
	output \g80676/_0_  ;
	output \g80798/_0_  ;
	output \g80807/_0_  ;
	output \g80890/_2_  ;
	output \g80904/_0_  ;
	output \g81719/_2_  ;
	output \g81746/_0_  ;
	output \g81775/_0_  ;
	output \g81872/_0_  ;
	output \g81961/_0_  ;
	output \g81968/_0_  ;
	output \g82096/_0_  ;
	output \g82123/_0_  ;
	output \g82147/_0_  ;
	output \g82147/_1_  ;
	output \g82335/_0_  ;
	output \g82338/_2_  ;
	output \g82368/_0_  ;
	output \g82460/_2_  ;
	output \g82469/_0_  ;
	output \g82481/_0_  ;
	output \g82625/_1_  ;
	output \g82711/_0_  ;
	output \g82772/_0_  ;
	output \g82946/_0_  ;
	output \g82947/_0_  ;
	output \g82956/_0_  ;
	output \g83003/_0_  ;
	output \g83006/_1_  ;
	output \g83415/_0_  ;
	output \g83498/_0_  ;
	output \g837/_0_  ;
	output \g838/_0_  ;
	output \g83863/_0_  ;
	output \g839/_0_  ;
	output \g84049/_3_  ;
	output \g84050/_3_  ;
	output \g84077/_2_  ;
	output \g842/_0_  ;
	output \g84245/_0_  ;
	output \g843/_0_  ;
	output \g844/_0_  ;
	output \g84448/_0_  ;
	output \g84478/_3_  ;
	output \g845/_0_  ;
	output \g846/_0_  ;
	output \g847/_0_  ;
	output \g848/_0_  ;
	output \g8487/_0_  ;
	output \g8488/_0_  ;
	output \g8489/_0_  ;
	output \g849/_0_  ;
	output \g8490/_0_  ;
	output \g84904/_0_  ;
	output \g8491/_0_  ;
	output \g8492/_0_  ;
	output \g8493/_0_  ;
	output \g8494/_0_  ;
	output \g8496/_0_  ;
	output \g8517/_0_  ;
	output \g8534/_0_  ;
	output \g8538/_0_  ;
	output \g8540/_0_  ;
	output \g8576/_2_  ;
	output \g8597/_0_  ;
	output \g8598/_0_  ;
	output \g8599/_0_  ;
	output \g8600/_0_  ;
	output \g8601/_0_  ;
	output \g8602/_0_  ;
	output \g8603/_0_  ;
	output \g8605/_0_  ;
	output \g8606/_0_  ;
	output \g8607/_0_  ;
	output \g8608/_0_  ;
	output \g8609/_0_  ;
	output \g8610/_0_  ;
	output \g8611/_0_  ;
	output \g8612/_0_  ;
	output \g8613/_0_  ;
	output \g8614/_0_  ;
	output \g8615/_0_  ;
	output \g8617/_0_  ;
	output \g8643/_0_  ;
	output \g8644/_0_  ;
	output \g8645/_0_  ;
	output \g8646/_0_  ;
	output \g8647/_0_  ;
	output \g8648/_0_  ;
	output \g8650/_0_  ;
	output \g8651/_0_  ;
	output \g8652/_0_  ;
	output \g8653/_0_  ;
	output \g8654/_0_  ;
	output \g8655/_0_  ;
	output \g8656/_0_  ;
	output \g8657/_0_  ;
	output \g8658/_0_  ;
	output \g8659/_0_  ;
	output \g8660/_0_  ;
	output \g8665/_00_  ;
	output \g8666/_00_  ;
	output \g8667/_00_  ;
	output \g8668/_00_  ;
	output \g8669/_00_  ;
	output \g86715/_0_  ;
	output \g86745/_3_  ;
	output \g8691/_0_  ;
	output \g8700/_0_  ;
	output \g8701/_0_  ;
	output \g8702/_0_  ;
	output \g8703/_0_  ;
	output \g8704/_0_  ;
	output \g8705/_0_  ;
	output \g87063/_0_  ;
	output \g87114/_0_  ;
	output \g8712/_0_  ;
	output \g8713/_0_  ;
	output \g8714/_0_  ;
	output \g87171/_1_  ;
	output \g87252/_1_  ;
	output \g87298/_0_  ;
	output \g8730/_0_  ;
	output \g8741/_0_  ;
	output \g8747/_0_  ;
	output \g87480/_0_  ;
	output \g87484/_2_  ;
	output \g87488/_1__syn_2  ;
	output \g8761/_0_  ;
	output \g8762/_0_  ;
	output \g8763/_0_  ;
	output \g8764/_0_  ;
	output \g8765/_0_  ;
	output \g8775/_0_  ;
	output \g8776/_0_  ;
	output \g8777/_0_  ;
	output \g8778/_0_  ;
	output \g8784/_0_  ;
	output \g8804/_0_  ;
	output \g8807/_0_  ;
	output \g8808/_0_  ;
	output \g8809/_0_  ;
	output \g8810/_0_  ;
	output \g8811/_0_  ;
	output \g8812/_0_  ;
	output \g8813/_0_  ;
	output \g8814/_0_  ;
	output \g8815/_0_  ;
	output \g8816/_0_  ;
	output \g8817/_0_  ;
	output \g8818/_0_  ;
	output \g8819/_0_  ;
	output \g8820/_0_  ;
	output \g8821/_0_  ;
	output \g8822/_0_  ;
	output \g8823/_0_  ;
	output \g8824/_0_  ;
	output \g8825/_0_  ;
	output \g8826/_0_  ;
	output \g8827/_0_  ;
	output \g8828/_0_  ;
	output \g8829/_0_  ;
	output \g8830/_0_  ;
	output \g8831/_0_  ;
	output \g8832/_0_  ;
	output \g8833/_0_  ;
	output \g8834/_0_  ;
	output \g8835/_0_  ;
	output \g8836/_0_  ;
	output \g8837/_0_  ;
	output \g8838/_0_  ;
	output \g8839/_0_  ;
	output \g8840/_0_  ;
	output \g8842/_0_  ;
	output \g8843/_0_  ;
	output \g8846/_0_  ;
	output \g8848/_0_  ;
	output \g8857/_0_  ;
	output \g8895/_0_  ;
	output \g8902/_3_  ;
	output \g8903/_3_  ;
	output \g8904/_3_  ;
	output \g8905/_3_  ;
	output \g8906/_3_  ;
	output \g8909/_0_  ;
	output \g8910/_0_  ;
	output \g8911/_0_  ;
	output \g8924/_3_  ;
	output \g8926/_3_  ;
	output \g8927/_3_  ;
	output \g8943/_0_  ;
	output \g8944/_0_  ;
	output \g8958/_3_  ;
	output \g8960/_00_  ;
	output \g8961/_3_  ;
	output \g8965/_0_  ;
	output \g8966/_0_  ;
	output \g8967/_0_  ;
	output \g8968/_0_  ;
	output \g9/_0_  ;
	output \g9123/_0_  ;
	output \g9125/_0_  ;
	output \g9126/_0_  ;
	output \g913/_0_  ;
	output \g915/_0_  ;
	output \g916/_0_  ;
	output \g917/_0_  ;
	output \g918/_0_  ;
	output \g919/_0_  ;
	output \g920/_3_  ;
	output \g921/_3_  ;
	output \g925/_0_  ;
	output \g926/_0_  ;
	output \g927/_0_  ;
	output \g928/_0_  ;
	output \g929/_0_  ;
	output \g930/_0_  ;
	output \g9336/_0_  ;
	output \g9337/_0_  ;
	output \g939/_3_  ;
	output \g9396/_0_  ;
	output \g9397/_0_  ;
	output \g9399/_0_  ;
	output \g9400/_0_  ;
	output \g9401/_0_  ;
	output \g9402/_0_  ;
	output \g9403/_0_  ;
	output \g9404/_0_  ;
	output \g9415/_0_  ;
	output \g9418/_0_  ;
	output \g9419/_0_  ;
	output \g9420/_0_  ;
	output \g9446/_0_  ;
	output \g9465/_0_  ;
	output \g9493/_0_  ;
	output \g9536/_0_  ;
	output \g9537/_0_  ;
	output \g9538/_0_  ;
	output \g9539/_0_  ;
	output \g9540/_0_  ;
	output \g9541/_0_  ;
	output \g9542/_0_  ;
	output \g955/_2_  ;
	output \g9561/_0_  ;
	output \g9562/_0_  ;
	output \g9563/_0_  ;
	output \g9564/_0_  ;
	output \g9565/_0_  ;
	output \g9566/_0_  ;
	output \g9567/_0_  ;
	output \g9568/_0_  ;
	output \g9569/_0_  ;
	output \g9570/_0_  ;
	output \g9571/_0_  ;
	output \g9572/_0_  ;
	output \g9573/_0_  ;
	output \g9574/_0_  ;
	output \g9575/_0_  ;
	output \g9576/_0_  ;
	output \g9577/_0_  ;
	output \g9578/_0_  ;
	output \g9579/_0_  ;
	output \g9580/_0_  ;
	output \g9581/_0_  ;
	output \g9582/_0_  ;
	output \g9583/_0_  ;
	output \g9584/_0_  ;
	output \g9585/_0_  ;
	output \g9586/_0_  ;
	output \g9587/_0_  ;
	output \g9588/_0_  ;
	output \g9589/_0_  ;
	output \g9590/_0_  ;
	output \g9591/_0_  ;
	output \g9592/_0_  ;
	output \g9593/_0_  ;
	output \g9594/_0_  ;
	output \g9595/_0_  ;
	output \g9596/_0_  ;
	output \g9597/_0_  ;
	output \g9598/_0_  ;
	output \g9599/_0_  ;
	output \g9600/_0_  ;
	output \g9601/_0_  ;
	output \g9602/_0_  ;
	output \g9603/_0_  ;
	output \g9604/_0_  ;
	output \g9605/_0_  ;
	output \g9606/_0_  ;
	output \g9607/_0_  ;
	output \g9608/_0_  ;
	output \g9609/_0_  ;
	output \g9610/_0_  ;
	output \g9611/_0_  ;
	output \g9612/_0_  ;
	output \g9613/_0_  ;
	output \g9614/_0_  ;
	output \g9615/_0_  ;
	output \g9616/_0_  ;
	output \g9617/_0_  ;
	output \g9618/_0_  ;
	output \g9619/_0_  ;
	output \g9620/_0_  ;
	output \g9621/_0_  ;
	output \g9622/_0_  ;
	output \g9623/_0_  ;
	output \g9624/_0_  ;
	output \g9625/_0_  ;
	output \g9626/_0_  ;
	output \g9627/_0_  ;
	output \g9628/_0_  ;
	output \g9629/_0_  ;
	output \g9630/_0_  ;
	output \g9631/_0_  ;
	output \g9632/_0_  ;
	output \g9633/_0_  ;
	output \g9634/_0_  ;
	output \g9635/_0_  ;
	output \g9636/_0_  ;
	output \g9637/_0_  ;
	output \g9638/_0_  ;
	output \g9639/_0_  ;
	output \g9640/_0_  ;
	output \g9641/_0_  ;
	output \g9642/_0_  ;
	output \g9643/_0_  ;
	output \g9644/_0_  ;
	output \g9645/_0_  ;
	output \g9646/_0_  ;
	output \g9647/_0_  ;
	output \g9648/_0_  ;
	output \g9649/_0_  ;
	output \g9650/_0_  ;
	output \g9651/_0_  ;
	output \g9652/_0_  ;
	output \g9653/_0_  ;
	output \g9654/_0_  ;
	output \g9655/_0_  ;
	output \g9656/_0_  ;
	output \g9657/_0_  ;
	output \g9658/_0_  ;
	output \g9659/_0_  ;
	output \g9660/_0_  ;
	output \g9661/_0_  ;
	output \g9662/_0_  ;
	output \g9663/_0_  ;
	output \g9664/_0_  ;
	output \g9665/_0_  ;
	output \g9666/_0_  ;
	output \g9667/_0_  ;
	output \g9668/_0_  ;
	output \g9669/_0_  ;
	output \g9670/_0_  ;
	output \g9671/_0_  ;
	output \g9672/_0_  ;
	output \g9673/_0_  ;
	output \g9674/_0_  ;
	output \g9675/_0_  ;
	output \g9676/_0_  ;
	output \g9677/_0_  ;
	output \g9678/_0_  ;
	output \g9681/_0_  ;
	output \g9683/_0_  ;
	output \g9689/_0_  ;
	output \g9692/_0_  ;
	output \g9694/_0_  ;
	output \g9695/_0_  ;
	output \g9701/_0_  ;
	output \g9702/_0_  ;
	output \g9703/_0_  ;
	output \g9704/_0_  ;
	output \g9709/_0_  ;
	output \g9710/_0_  ;
	output \g9711/_0_  ;
	output \g9712/_0_  ;
	output \g9720/_0_  ;
	output \g9721/_0_  ;
	output \g9722/_0_  ;
	output \g9726/_0_  ;
	output \g9733/_0_  ;
	output \g9734/_0_  ;
	output \g9735/_0_  ;
	output \g9736/_0_  ;
	output \g9737/_0_  ;
	output \g9738/_0_  ;
	output \g9739/_0_  ;
	output \g9740/_0_  ;
	output \g9741/_0_  ;
	output \g9742/_0_  ;
	output \g9743/_0_  ;
	output \g9744/_0_  ;
	output \g9745/_0_  ;
	output \g9746/_0_  ;
	output \g9747/_0_  ;
	output \g9748/_0_  ;
	output \g9749/_0_  ;
	output \g9750/_0_  ;
	output \g9751/_0_  ;
	output \g9752/_0_  ;
	output \g9753/_0_  ;
	output \g9754/_0_  ;
	output \g9755/_0_  ;
	output \g9756/_0_  ;
	output \g9757/_0_  ;
	output \g9758/_0_  ;
	output \g9759/_0_  ;
	output \g9760/_0_  ;
	output \g9761/_0_  ;
	output \g9762/_0_  ;
	output \g9763/_0_  ;
	output \g9764/_0_  ;
	output \g9765/_0_  ;
	output \g9766/_0_  ;
	output \g9767/_0_  ;
	output \g9768/_0_  ;
	output \g9769/_0_  ;
	output \g9770/_0_  ;
	output \g9771/_0_  ;
	output \g9772/_0_  ;
	output \g9773/_0_  ;
	output \g9774/_0_  ;
	output \g9775/_0_  ;
	output \g9776/_0_  ;
	output \g9777/_0_  ;
	output \g9778/_0_  ;
	output \g9779/_0_  ;
	output \g9780/_0_  ;
	output \g9781/_0_  ;
	output \g9782/_0_  ;
	output \g9783/_0_  ;
	output \g9784/_0_  ;
	output \g9785/_0_  ;
	output \g9786/_0_  ;
	output \g9787/_0_  ;
	output \g9788/_0_  ;
	output \g9789/_0_  ;
	output \g9790/_0_  ;
	output \g9791/_0_  ;
	output \g9792/_0_  ;
	output \g9793/_0_  ;
	output \g9794/_0_  ;
	output \g9795/_0_  ;
	output \g9796/_0_  ;
	output \g9797/_0_  ;
	output \g9798/_0_  ;
	output \g9799/_0_  ;
	output \g9800/_0_  ;
	output \g9801/_0_  ;
	output \g9802/_0_  ;
	output \g9803/_0_  ;
	output \g9804/_0_  ;
	output \g9805/_0_  ;
	output \g9806/_0_  ;
	output \g9807/_0_  ;
	output \g9808/_0_  ;
	output \g9809/_0_  ;
	output \g9810/_0_  ;
	output \g9811/_0_  ;
	output \g9812/_0_  ;
	output \g9813/_0_  ;
	output \g9814/_0_  ;
	output \g9815/_0_  ;
	output \g9816/_0_  ;
	output \g9817/_0_  ;
	output \g9818/_0_  ;
	output \g9819/_0_  ;
	output \g9820/_0_  ;
	output \g9821/_0_  ;
	output \g9822/_0_  ;
	output \g9823/_0_  ;
	output \g9824/_0_  ;
	output \g9825/_0_  ;
	output \g9826/_0_  ;
	output \g9827/_0_  ;
	output \g9828/_0_  ;
	output \g9829/_0_  ;
	output \g9830/_0_  ;
	output \g9831/_0_  ;
	output \g9832/_0_  ;
	output \g9833/_0_  ;
	output \g9835/_0_  ;
	output \g9836/_0_  ;
	output \g9837/_0_  ;
	output \g9838/_0_  ;
	output \g9839/_0_  ;
	output \g9840/_0_  ;
	output \g9841/_0_  ;
	output \g9842/_0_  ;
	output \g9844/_0_  ;
	output \g9845/_0_  ;
	output \g9846/_0_  ;
	output \g9848/_0_  ;
	output \g9849/_0_  ;
	output \g9850/_0_  ;
	output \g9851/_0_  ;
	output \g9853/_0_  ;
	output \g9854/_0_  ;
	output \g9855/_0_  ;
	output \g9856/_0_  ;
	output \g9857/_0_  ;
	output \g9858/_0_  ;
	output \g9859/_0_  ;
	output \g9860/_0_  ;
	output \g9862/_0_  ;
	output \g9863/_0_  ;
	output \g9864/_0_  ;
	output \g9865/_0_  ;
	output \g9867/_0_  ;
	output \g9868/_0_  ;
	output \g9876/_0_  ;
	output \g9877/_0_  ;
	output \g9878/_0_  ;
	output \g9879/_0_  ;
	output \g9880/_0_  ;
	output \g9881/_0_  ;
	output \g9898/_0_  ;
	output \g9900/_0_  ;
	output \g9901/_0_  ;
	output \g9902/_0_  ;
	output \g9903/_0_  ;
	output \g9904/_0_  ;
	output \g9905/_0_  ;
	output \g9906/_0_  ;
	output \g9907/_0_  ;
	output \g9908/_0_  ;
	output \g9909/_0_  ;
	output \g9910/_0_  ;
	output \g9911/_0_  ;
	output \g9912/_0_  ;
	output \g9913/_0_  ;
	output \g9914/_0_  ;
	output \g9915/_0_  ;
	output \g9916/_0_  ;
	output \g9917/_0_  ;
	output \g9918/_0_  ;
	output \g9919/_0_  ;
	output \g992/_0_  ;
	output \g9920/_0_  ;
	output \g9921/_0_  ;
	output \g9922/_0_  ;
	output \g9923/_0_  ;
	output \g9924/_0_  ;
	output \g9925/_0_  ;
	output \g9926/_0_  ;
	output \g9927/_0_  ;
	output \g9928/_0_  ;
	output \g9929/_0_  ;
	output \g9930/_0_  ;
	output \g9931/_0_  ;
	output \g9932/_0_  ;
	output \g9933/_0_  ;
	output \g9934/_0_  ;
	output \g9935/_0_  ;
	output \g9936/_0_  ;
	output \g9937/_0_  ;
	output \g9938/_0_  ;
	output \g9939/_0_  ;
	output \g9940/_0_  ;
	output \g9941/_0_  ;
	output \g9942/_0_  ;
	output \g9943/_0_  ;
	output \g9944/_0_  ;
	output \g9945/_0_  ;
	output \g9946/_0_  ;
	output \g9947/_0_  ;
	output \g9948/_0_  ;
	output \g9949/_0_  ;
	output \g9950/_0_  ;
	output \g9951/_0_  ;
	output \g9952/_0_  ;
	output \g9953/_0_  ;
	output \g9954/_0_  ;
	output \g9955/_0_  ;
	output \g9956/_0_  ;
	output \g9957/_0_  ;
	output \g9958/_0_  ;
	output \g9959/_0_  ;
	output \g9960/_0_  ;
	output \g9961/_0_  ;
	output \g9962/_0_  ;
	output \g9963/_0_  ;
	output \g9964/_0_  ;
	output \g9965/_0_  ;
	output \g9966/_0_  ;
	output \g9967/_0_  ;
	output \g9968/_0_  ;
	output \g9969/_0_  ;
	output \g9970/_0_  ;
	output \g9971/_0_  ;
	output \g9972/_0_  ;
	output \g9973/_0_  ;
	output \g9974/_0_  ;
	output \g9975/_0_  ;
	output \g9976/_0_  ;
	output \g9977/_0_  ;
	output \g9978/_0_  ;
	output \g9979/_0_  ;
	output \g9980/_0_  ;
	output \g9981/_0_  ;
	output \g9982/_0_  ;
	output \g9983/_0_  ;
	output \g9984/_0_  ;
	output \g9985/_0_  ;
	output \g9987/_0_  ;
	output \g9988/_0_  ;
	output \g9989/_0_  ;
	output \g999/_0_  ;
	output \g9990/_0_  ;
	output \g9991/_0_  ;
	output \g9992/_0_  ;
	output \g9993/_0_  ;
	output \g9994/_0_  ;
	output \g9995/_0_  ;
	output \g9996/_0_  ;
	output \g9997/_0_  ;
	output \g9998/_0_  ;
	output \g9999/_0_  ;
	output \idma_IDMA_boot_reg/NET0131_reg_syn_3  ;
	output \memc_EXTC_Eg_reg/NET0131  ;
	output \memc_EXTC_Eg_reg/NET0131_reg_syn_3  ;
	output \memc_EXTC_Eg_reg/n0  ;
	output \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3  ;
	output \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3  ;
	output \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3  ;
	output \sice_GO_NXi_reg/NET0131_reg_syn_3  ;
	output \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  ;
	output \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  ;
	output \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  ;
	output \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  ;
	wire _w38588_ ;
	wire _w38587_ ;
	wire _w38586_ ;
	wire _w38585_ ;
	wire _w38584_ ;
	wire _w38583_ ;
	wire _w38582_ ;
	wire _w38581_ ;
	wire _w38580_ ;
	wire _w38579_ ;
	wire _w38578_ ;
	wire _w38577_ ;
	wire _w38576_ ;
	wire _w38575_ ;
	wire _w38574_ ;
	wire _w38573_ ;
	wire _w38572_ ;
	wire _w38571_ ;
	wire _w38570_ ;
	wire _w38569_ ;
	wire _w38568_ ;
	wire _w38567_ ;
	wire _w38566_ ;
	wire _w38565_ ;
	wire _w38564_ ;
	wire _w38563_ ;
	wire _w38562_ ;
	wire _w38561_ ;
	wire _w38560_ ;
	wire _w38559_ ;
	wire _w38558_ ;
	wire _w38557_ ;
	wire _w38556_ ;
	wire _w38555_ ;
	wire _w38554_ ;
	wire _w38553_ ;
	wire _w38552_ ;
	wire _w38551_ ;
	wire _w38550_ ;
	wire _w38549_ ;
	wire _w38548_ ;
	wire _w38547_ ;
	wire _w38546_ ;
	wire _w38545_ ;
	wire _w38544_ ;
	wire _w38543_ ;
	wire _w38542_ ;
	wire _w38541_ ;
	wire _w38540_ ;
	wire _w38539_ ;
	wire _w38538_ ;
	wire _w38537_ ;
	wire _w38536_ ;
	wire _w38535_ ;
	wire _w38534_ ;
	wire _w38533_ ;
	wire _w38532_ ;
	wire _w38531_ ;
	wire _w38530_ ;
	wire _w38529_ ;
	wire _w38528_ ;
	wire _w38527_ ;
	wire _w38526_ ;
	wire _w38525_ ;
	wire _w38524_ ;
	wire _w38523_ ;
	wire _w38522_ ;
	wire _w38521_ ;
	wire _w38520_ ;
	wire _w38519_ ;
	wire _w38518_ ;
	wire _w38517_ ;
	wire _w38516_ ;
	wire _w38515_ ;
	wire _w38514_ ;
	wire _w38513_ ;
	wire _w38512_ ;
	wire _w38511_ ;
	wire _w38510_ ;
	wire _w38509_ ;
	wire _w38508_ ;
	wire _w38507_ ;
	wire _w38506_ ;
	wire _w38505_ ;
	wire _w38504_ ;
	wire _w38503_ ;
	wire _w38502_ ;
	wire _w38501_ ;
	wire _w38500_ ;
	wire _w38499_ ;
	wire _w38498_ ;
	wire _w38497_ ;
	wire _w38496_ ;
	wire _w38495_ ;
	wire _w38494_ ;
	wire _w38493_ ;
	wire _w38492_ ;
	wire _w38491_ ;
	wire _w38490_ ;
	wire _w38489_ ;
	wire _w38488_ ;
	wire _w38487_ ;
	wire _w38486_ ;
	wire _w38485_ ;
	wire _w38484_ ;
	wire _w38483_ ;
	wire _w38482_ ;
	wire _w38481_ ;
	wire _w38480_ ;
	wire _w38479_ ;
	wire _w38478_ ;
	wire _w38477_ ;
	wire _w38476_ ;
	wire _w38475_ ;
	wire _w38474_ ;
	wire _w38473_ ;
	wire _w38472_ ;
	wire _w38471_ ;
	wire _w38470_ ;
	wire _w38469_ ;
	wire _w38468_ ;
	wire _w38467_ ;
	wire _w38466_ ;
	wire _w38465_ ;
	wire _w38464_ ;
	wire _w38463_ ;
	wire _w38462_ ;
	wire _w38461_ ;
	wire _w38460_ ;
	wire _w38459_ ;
	wire _w38458_ ;
	wire _w38457_ ;
	wire _w38456_ ;
	wire _w38455_ ;
	wire _w38454_ ;
	wire _w38453_ ;
	wire _w38452_ ;
	wire _w38451_ ;
	wire _w38450_ ;
	wire _w38449_ ;
	wire _w38448_ ;
	wire _w38447_ ;
	wire _w38446_ ;
	wire _w38445_ ;
	wire _w38444_ ;
	wire _w38443_ ;
	wire _w38442_ ;
	wire _w38441_ ;
	wire _w38440_ ;
	wire _w38439_ ;
	wire _w38438_ ;
	wire _w38437_ ;
	wire _w38436_ ;
	wire _w38435_ ;
	wire _w38434_ ;
	wire _w38433_ ;
	wire _w38432_ ;
	wire _w38431_ ;
	wire _w38430_ ;
	wire _w38429_ ;
	wire _w38428_ ;
	wire _w38427_ ;
	wire _w38426_ ;
	wire _w38425_ ;
	wire _w38424_ ;
	wire _w38423_ ;
	wire _w38422_ ;
	wire _w38421_ ;
	wire _w38420_ ;
	wire _w38419_ ;
	wire _w38418_ ;
	wire _w38417_ ;
	wire _w38416_ ;
	wire _w38415_ ;
	wire _w38414_ ;
	wire _w38413_ ;
	wire _w38412_ ;
	wire _w38411_ ;
	wire _w38410_ ;
	wire _w38409_ ;
	wire _w38408_ ;
	wire _w38407_ ;
	wire _w38406_ ;
	wire _w38405_ ;
	wire _w38404_ ;
	wire _w38403_ ;
	wire _w38402_ ;
	wire _w38401_ ;
	wire _w38400_ ;
	wire _w38399_ ;
	wire _w38398_ ;
	wire _w38397_ ;
	wire _w38396_ ;
	wire _w38395_ ;
	wire _w38394_ ;
	wire _w38393_ ;
	wire _w38392_ ;
	wire _w38391_ ;
	wire _w38390_ ;
	wire _w38389_ ;
	wire _w38388_ ;
	wire _w38387_ ;
	wire _w38386_ ;
	wire _w38385_ ;
	wire _w38384_ ;
	wire _w38383_ ;
	wire _w38382_ ;
	wire _w38381_ ;
	wire _w38380_ ;
	wire _w38379_ ;
	wire _w38378_ ;
	wire _w38377_ ;
	wire _w38376_ ;
	wire _w38375_ ;
	wire _w38374_ ;
	wire _w38373_ ;
	wire _w38372_ ;
	wire _w38371_ ;
	wire _w38370_ ;
	wire _w38369_ ;
	wire _w38368_ ;
	wire _w38367_ ;
	wire _w38366_ ;
	wire _w38365_ ;
	wire _w38364_ ;
	wire _w38363_ ;
	wire _w38362_ ;
	wire _w38361_ ;
	wire _w38360_ ;
	wire _w38359_ ;
	wire _w38358_ ;
	wire _w38357_ ;
	wire _w38356_ ;
	wire _w38355_ ;
	wire _w38354_ ;
	wire _w38353_ ;
	wire _w38352_ ;
	wire _w38351_ ;
	wire _w38350_ ;
	wire _w38349_ ;
	wire _w38348_ ;
	wire _w38347_ ;
	wire _w38346_ ;
	wire _w38345_ ;
	wire _w38344_ ;
	wire _w38343_ ;
	wire _w38342_ ;
	wire _w38341_ ;
	wire _w38340_ ;
	wire _w38339_ ;
	wire _w38338_ ;
	wire _w38337_ ;
	wire _w38336_ ;
	wire _w38335_ ;
	wire _w38334_ ;
	wire _w38333_ ;
	wire _w38332_ ;
	wire _w38331_ ;
	wire _w38330_ ;
	wire _w38329_ ;
	wire _w38328_ ;
	wire _w38327_ ;
	wire _w38326_ ;
	wire _w38325_ ;
	wire _w38324_ ;
	wire _w38323_ ;
	wire _w38322_ ;
	wire _w38321_ ;
	wire _w38320_ ;
	wire _w38319_ ;
	wire _w38318_ ;
	wire _w38317_ ;
	wire _w38316_ ;
	wire _w38315_ ;
	wire _w38314_ ;
	wire _w38313_ ;
	wire _w38312_ ;
	wire _w38311_ ;
	wire _w38310_ ;
	wire _w38309_ ;
	wire _w38308_ ;
	wire _w38307_ ;
	wire _w38306_ ;
	wire _w38305_ ;
	wire _w38304_ ;
	wire _w38303_ ;
	wire _w38302_ ;
	wire _w38301_ ;
	wire _w38300_ ;
	wire _w38299_ ;
	wire _w38298_ ;
	wire _w38297_ ;
	wire _w38296_ ;
	wire _w38295_ ;
	wire _w38294_ ;
	wire _w38293_ ;
	wire _w38292_ ;
	wire _w38291_ ;
	wire _w38290_ ;
	wire _w38289_ ;
	wire _w38288_ ;
	wire _w38287_ ;
	wire _w38286_ ;
	wire _w38285_ ;
	wire _w38284_ ;
	wire _w38283_ ;
	wire _w38282_ ;
	wire _w38281_ ;
	wire _w38280_ ;
	wire _w38279_ ;
	wire _w38278_ ;
	wire _w38277_ ;
	wire _w38276_ ;
	wire _w38275_ ;
	wire _w38274_ ;
	wire _w38273_ ;
	wire _w38272_ ;
	wire _w38271_ ;
	wire _w38270_ ;
	wire _w38269_ ;
	wire _w38268_ ;
	wire _w38267_ ;
	wire _w38266_ ;
	wire _w38265_ ;
	wire _w38264_ ;
	wire _w38263_ ;
	wire _w38262_ ;
	wire _w38261_ ;
	wire _w38260_ ;
	wire _w38259_ ;
	wire _w38258_ ;
	wire _w38257_ ;
	wire _w38256_ ;
	wire _w38255_ ;
	wire _w38254_ ;
	wire _w38253_ ;
	wire _w38252_ ;
	wire _w38251_ ;
	wire _w38250_ ;
	wire _w38249_ ;
	wire _w38248_ ;
	wire _w38247_ ;
	wire _w38246_ ;
	wire _w38245_ ;
	wire _w38244_ ;
	wire _w38243_ ;
	wire _w38242_ ;
	wire _w38241_ ;
	wire _w38240_ ;
	wire _w38239_ ;
	wire _w38238_ ;
	wire _w38237_ ;
	wire _w38236_ ;
	wire _w38235_ ;
	wire _w38234_ ;
	wire _w38233_ ;
	wire _w38232_ ;
	wire _w38231_ ;
	wire _w38230_ ;
	wire _w38229_ ;
	wire _w38228_ ;
	wire _w38227_ ;
	wire _w38226_ ;
	wire _w38225_ ;
	wire _w38224_ ;
	wire _w38223_ ;
	wire _w38222_ ;
	wire _w38221_ ;
	wire _w38220_ ;
	wire _w38219_ ;
	wire _w38218_ ;
	wire _w38217_ ;
	wire _w38216_ ;
	wire _w38215_ ;
	wire _w38214_ ;
	wire _w38213_ ;
	wire _w38212_ ;
	wire _w38211_ ;
	wire _w38210_ ;
	wire _w38209_ ;
	wire _w38208_ ;
	wire _w38207_ ;
	wire _w38206_ ;
	wire _w38205_ ;
	wire _w38204_ ;
	wire _w38203_ ;
	wire _w38202_ ;
	wire _w38201_ ;
	wire _w38200_ ;
	wire _w38199_ ;
	wire _w38198_ ;
	wire _w38197_ ;
	wire _w38196_ ;
	wire _w38195_ ;
	wire _w38194_ ;
	wire _w38193_ ;
	wire _w38192_ ;
	wire _w38191_ ;
	wire _w38190_ ;
	wire _w38189_ ;
	wire _w38188_ ;
	wire _w38187_ ;
	wire _w38186_ ;
	wire _w38185_ ;
	wire _w38184_ ;
	wire _w38183_ ;
	wire _w38182_ ;
	wire _w38181_ ;
	wire _w38180_ ;
	wire _w38179_ ;
	wire _w38178_ ;
	wire _w38177_ ;
	wire _w38176_ ;
	wire _w38175_ ;
	wire _w38174_ ;
	wire _w38173_ ;
	wire _w38172_ ;
	wire _w38171_ ;
	wire _w38170_ ;
	wire _w38169_ ;
	wire _w38168_ ;
	wire _w38167_ ;
	wire _w38166_ ;
	wire _w38165_ ;
	wire _w38164_ ;
	wire _w38163_ ;
	wire _w38162_ ;
	wire _w38161_ ;
	wire _w38160_ ;
	wire _w38159_ ;
	wire _w38158_ ;
	wire _w38157_ ;
	wire _w38156_ ;
	wire _w38155_ ;
	wire _w38154_ ;
	wire _w38153_ ;
	wire _w38152_ ;
	wire _w38151_ ;
	wire _w38150_ ;
	wire _w38149_ ;
	wire _w38148_ ;
	wire _w38147_ ;
	wire _w38146_ ;
	wire _w38145_ ;
	wire _w38144_ ;
	wire _w38143_ ;
	wire _w38142_ ;
	wire _w38141_ ;
	wire _w38140_ ;
	wire _w38139_ ;
	wire _w38138_ ;
	wire _w38137_ ;
	wire _w38136_ ;
	wire _w38135_ ;
	wire _w38134_ ;
	wire _w38133_ ;
	wire _w38132_ ;
	wire _w38131_ ;
	wire _w38130_ ;
	wire _w38129_ ;
	wire _w38128_ ;
	wire _w38127_ ;
	wire _w38126_ ;
	wire _w38125_ ;
	wire _w38124_ ;
	wire _w38123_ ;
	wire _w38122_ ;
	wire _w38121_ ;
	wire _w38120_ ;
	wire _w38119_ ;
	wire _w38118_ ;
	wire _w38117_ ;
	wire _w38116_ ;
	wire _w38115_ ;
	wire _w38114_ ;
	wire _w38113_ ;
	wire _w38112_ ;
	wire _w38111_ ;
	wire _w38110_ ;
	wire _w38109_ ;
	wire _w38108_ ;
	wire _w38107_ ;
	wire _w38106_ ;
	wire _w38105_ ;
	wire _w38104_ ;
	wire _w38103_ ;
	wire _w38102_ ;
	wire _w38101_ ;
	wire _w38100_ ;
	wire _w38099_ ;
	wire _w38098_ ;
	wire _w38097_ ;
	wire _w38096_ ;
	wire _w38095_ ;
	wire _w38094_ ;
	wire _w38093_ ;
	wire _w38092_ ;
	wire _w38091_ ;
	wire _w38090_ ;
	wire _w38089_ ;
	wire _w38088_ ;
	wire _w38087_ ;
	wire _w38086_ ;
	wire _w38085_ ;
	wire _w38084_ ;
	wire _w38083_ ;
	wire _w38082_ ;
	wire _w38081_ ;
	wire _w38080_ ;
	wire _w38079_ ;
	wire _w38078_ ;
	wire _w38077_ ;
	wire _w38076_ ;
	wire _w38075_ ;
	wire _w38074_ ;
	wire _w38073_ ;
	wire _w38072_ ;
	wire _w38071_ ;
	wire _w38070_ ;
	wire _w38069_ ;
	wire _w38068_ ;
	wire _w38067_ ;
	wire _w38066_ ;
	wire _w38065_ ;
	wire _w38064_ ;
	wire _w38063_ ;
	wire _w38062_ ;
	wire _w38061_ ;
	wire _w38060_ ;
	wire _w38059_ ;
	wire _w38058_ ;
	wire _w38057_ ;
	wire _w38056_ ;
	wire _w38055_ ;
	wire _w38054_ ;
	wire _w38053_ ;
	wire _w38052_ ;
	wire _w38051_ ;
	wire _w38050_ ;
	wire _w38049_ ;
	wire _w38048_ ;
	wire _w38047_ ;
	wire _w38046_ ;
	wire _w38045_ ;
	wire _w38044_ ;
	wire _w38043_ ;
	wire _w38042_ ;
	wire _w38041_ ;
	wire _w38040_ ;
	wire _w38039_ ;
	wire _w38038_ ;
	wire _w38037_ ;
	wire _w38036_ ;
	wire _w38035_ ;
	wire _w38034_ ;
	wire _w38033_ ;
	wire _w38032_ ;
	wire _w38031_ ;
	wire _w38030_ ;
	wire _w38029_ ;
	wire _w38028_ ;
	wire _w38027_ ;
	wire _w38026_ ;
	wire _w38025_ ;
	wire _w38024_ ;
	wire _w38023_ ;
	wire _w38022_ ;
	wire _w38021_ ;
	wire _w38020_ ;
	wire _w38019_ ;
	wire _w38018_ ;
	wire _w38017_ ;
	wire _w38016_ ;
	wire _w38015_ ;
	wire _w38014_ ;
	wire _w38013_ ;
	wire _w38012_ ;
	wire _w38011_ ;
	wire _w38010_ ;
	wire _w38009_ ;
	wire _w38008_ ;
	wire _w38007_ ;
	wire _w38006_ ;
	wire _w38005_ ;
	wire _w38004_ ;
	wire _w38003_ ;
	wire _w38002_ ;
	wire _w38001_ ;
	wire _w38000_ ;
	wire _w37999_ ;
	wire _w37998_ ;
	wire _w37997_ ;
	wire _w37996_ ;
	wire _w37995_ ;
	wire _w37994_ ;
	wire _w37993_ ;
	wire _w37992_ ;
	wire _w37991_ ;
	wire _w37990_ ;
	wire _w37989_ ;
	wire _w37988_ ;
	wire _w37987_ ;
	wire _w37986_ ;
	wire _w37985_ ;
	wire _w37984_ ;
	wire _w37983_ ;
	wire _w37982_ ;
	wire _w37981_ ;
	wire _w37980_ ;
	wire _w37979_ ;
	wire _w37978_ ;
	wire _w37977_ ;
	wire _w37976_ ;
	wire _w37975_ ;
	wire _w37974_ ;
	wire _w37973_ ;
	wire _w37972_ ;
	wire _w37971_ ;
	wire _w37970_ ;
	wire _w37969_ ;
	wire _w37968_ ;
	wire _w37967_ ;
	wire _w37966_ ;
	wire _w37965_ ;
	wire _w37964_ ;
	wire _w37963_ ;
	wire _w37962_ ;
	wire _w37961_ ;
	wire _w37960_ ;
	wire _w37959_ ;
	wire _w37958_ ;
	wire _w37957_ ;
	wire _w37956_ ;
	wire _w37955_ ;
	wire _w37954_ ;
	wire _w37953_ ;
	wire _w37952_ ;
	wire _w37951_ ;
	wire _w37950_ ;
	wire _w37949_ ;
	wire _w37948_ ;
	wire _w37947_ ;
	wire _w37946_ ;
	wire _w37945_ ;
	wire _w37944_ ;
	wire _w37943_ ;
	wire _w37942_ ;
	wire _w37941_ ;
	wire _w37940_ ;
	wire _w37939_ ;
	wire _w37938_ ;
	wire _w37937_ ;
	wire _w37936_ ;
	wire _w37935_ ;
	wire _w37934_ ;
	wire _w37933_ ;
	wire _w37932_ ;
	wire _w37931_ ;
	wire _w37930_ ;
	wire _w37929_ ;
	wire _w37928_ ;
	wire _w37927_ ;
	wire _w37926_ ;
	wire _w37925_ ;
	wire _w37924_ ;
	wire _w37923_ ;
	wire _w37922_ ;
	wire _w37921_ ;
	wire _w37920_ ;
	wire _w37919_ ;
	wire _w37918_ ;
	wire _w37917_ ;
	wire _w37916_ ;
	wire _w37915_ ;
	wire _w37914_ ;
	wire _w37913_ ;
	wire _w37912_ ;
	wire _w37911_ ;
	wire _w37910_ ;
	wire _w37909_ ;
	wire _w37908_ ;
	wire _w37907_ ;
	wire _w37906_ ;
	wire _w37905_ ;
	wire _w37904_ ;
	wire _w37903_ ;
	wire _w37902_ ;
	wire _w37901_ ;
	wire _w37900_ ;
	wire _w37899_ ;
	wire _w37898_ ;
	wire _w37897_ ;
	wire _w37896_ ;
	wire _w37895_ ;
	wire _w37894_ ;
	wire _w37893_ ;
	wire _w37892_ ;
	wire _w37891_ ;
	wire _w37890_ ;
	wire _w37889_ ;
	wire _w37888_ ;
	wire _w37887_ ;
	wire _w37886_ ;
	wire _w37885_ ;
	wire _w37884_ ;
	wire _w37883_ ;
	wire _w37882_ ;
	wire _w37881_ ;
	wire _w37880_ ;
	wire _w37879_ ;
	wire _w37878_ ;
	wire _w37877_ ;
	wire _w37876_ ;
	wire _w37875_ ;
	wire _w37874_ ;
	wire _w37873_ ;
	wire _w37872_ ;
	wire _w37871_ ;
	wire _w37870_ ;
	wire _w37869_ ;
	wire _w37868_ ;
	wire _w37867_ ;
	wire _w37866_ ;
	wire _w37865_ ;
	wire _w37864_ ;
	wire _w37863_ ;
	wire _w37862_ ;
	wire _w37861_ ;
	wire _w37860_ ;
	wire _w37859_ ;
	wire _w37858_ ;
	wire _w37857_ ;
	wire _w37856_ ;
	wire _w37855_ ;
	wire _w37854_ ;
	wire _w37853_ ;
	wire _w37852_ ;
	wire _w37851_ ;
	wire _w37850_ ;
	wire _w37849_ ;
	wire _w37848_ ;
	wire _w37847_ ;
	wire _w37846_ ;
	wire _w37845_ ;
	wire _w37844_ ;
	wire _w37843_ ;
	wire _w37842_ ;
	wire _w37841_ ;
	wire _w37840_ ;
	wire _w37839_ ;
	wire _w37838_ ;
	wire _w37837_ ;
	wire _w37836_ ;
	wire _w37835_ ;
	wire _w37834_ ;
	wire _w37833_ ;
	wire _w37832_ ;
	wire _w37831_ ;
	wire _w37830_ ;
	wire _w37829_ ;
	wire _w37828_ ;
	wire _w37827_ ;
	wire _w37826_ ;
	wire _w37825_ ;
	wire _w37824_ ;
	wire _w37823_ ;
	wire _w37822_ ;
	wire _w37821_ ;
	wire _w37820_ ;
	wire _w37819_ ;
	wire _w37818_ ;
	wire _w37817_ ;
	wire _w37816_ ;
	wire _w37815_ ;
	wire _w37814_ ;
	wire _w37813_ ;
	wire _w37812_ ;
	wire _w37811_ ;
	wire _w37810_ ;
	wire _w37809_ ;
	wire _w37808_ ;
	wire _w37807_ ;
	wire _w37806_ ;
	wire _w37805_ ;
	wire _w37804_ ;
	wire _w37803_ ;
	wire _w37802_ ;
	wire _w37801_ ;
	wire _w37800_ ;
	wire _w37799_ ;
	wire _w37798_ ;
	wire _w37797_ ;
	wire _w37796_ ;
	wire _w37795_ ;
	wire _w37794_ ;
	wire _w37793_ ;
	wire _w37792_ ;
	wire _w37791_ ;
	wire _w37790_ ;
	wire _w37789_ ;
	wire _w37788_ ;
	wire _w37787_ ;
	wire _w37786_ ;
	wire _w37785_ ;
	wire _w37784_ ;
	wire _w37783_ ;
	wire _w37782_ ;
	wire _w37781_ ;
	wire _w37780_ ;
	wire _w37779_ ;
	wire _w37778_ ;
	wire _w37777_ ;
	wire _w37776_ ;
	wire _w37775_ ;
	wire _w37774_ ;
	wire _w37773_ ;
	wire _w37772_ ;
	wire _w37771_ ;
	wire _w37770_ ;
	wire _w37769_ ;
	wire _w37768_ ;
	wire _w37767_ ;
	wire _w37766_ ;
	wire _w37765_ ;
	wire _w37764_ ;
	wire _w37763_ ;
	wire _w37762_ ;
	wire _w37761_ ;
	wire _w37760_ ;
	wire _w37759_ ;
	wire _w37758_ ;
	wire _w37757_ ;
	wire _w37756_ ;
	wire _w37755_ ;
	wire _w37754_ ;
	wire _w37753_ ;
	wire _w37752_ ;
	wire _w37751_ ;
	wire _w37750_ ;
	wire _w37749_ ;
	wire _w37748_ ;
	wire _w37747_ ;
	wire _w37746_ ;
	wire _w37745_ ;
	wire _w37744_ ;
	wire _w37743_ ;
	wire _w37742_ ;
	wire _w37741_ ;
	wire _w37740_ ;
	wire _w37739_ ;
	wire _w37738_ ;
	wire _w37737_ ;
	wire _w37736_ ;
	wire _w37735_ ;
	wire _w37734_ ;
	wire _w37733_ ;
	wire _w37732_ ;
	wire _w37731_ ;
	wire _w37730_ ;
	wire _w37729_ ;
	wire _w37728_ ;
	wire _w37727_ ;
	wire _w37726_ ;
	wire _w37725_ ;
	wire _w37724_ ;
	wire _w37723_ ;
	wire _w37722_ ;
	wire _w37721_ ;
	wire _w37720_ ;
	wire _w37719_ ;
	wire _w37718_ ;
	wire _w37717_ ;
	wire _w37716_ ;
	wire _w37715_ ;
	wire _w37714_ ;
	wire _w37713_ ;
	wire _w37712_ ;
	wire _w37711_ ;
	wire _w37710_ ;
	wire _w37709_ ;
	wire _w37708_ ;
	wire _w37707_ ;
	wire _w37706_ ;
	wire _w37705_ ;
	wire _w37704_ ;
	wire _w37703_ ;
	wire _w37702_ ;
	wire _w37701_ ;
	wire _w37700_ ;
	wire _w37699_ ;
	wire _w37698_ ;
	wire _w37697_ ;
	wire _w37696_ ;
	wire _w37695_ ;
	wire _w37694_ ;
	wire _w37693_ ;
	wire _w37692_ ;
	wire _w37691_ ;
	wire _w37690_ ;
	wire _w37689_ ;
	wire _w37688_ ;
	wire _w37687_ ;
	wire _w37686_ ;
	wire _w37685_ ;
	wire _w37684_ ;
	wire _w37683_ ;
	wire _w37682_ ;
	wire _w37681_ ;
	wire _w37680_ ;
	wire _w37679_ ;
	wire _w37678_ ;
	wire _w37677_ ;
	wire _w37676_ ;
	wire _w37675_ ;
	wire _w37674_ ;
	wire _w37673_ ;
	wire _w37672_ ;
	wire _w37671_ ;
	wire _w37670_ ;
	wire _w37669_ ;
	wire _w37668_ ;
	wire _w37667_ ;
	wire _w37666_ ;
	wire _w37665_ ;
	wire _w37664_ ;
	wire _w37663_ ;
	wire _w37662_ ;
	wire _w37661_ ;
	wire _w37660_ ;
	wire _w37659_ ;
	wire _w37658_ ;
	wire _w37657_ ;
	wire _w37656_ ;
	wire _w37655_ ;
	wire _w37654_ ;
	wire _w37653_ ;
	wire _w37652_ ;
	wire _w37651_ ;
	wire _w37650_ ;
	wire _w37649_ ;
	wire _w37648_ ;
	wire _w37647_ ;
	wire _w37646_ ;
	wire _w37645_ ;
	wire _w37644_ ;
	wire _w37643_ ;
	wire _w37642_ ;
	wire _w37641_ ;
	wire _w37640_ ;
	wire _w37639_ ;
	wire _w37638_ ;
	wire _w37637_ ;
	wire _w37636_ ;
	wire _w37635_ ;
	wire _w37634_ ;
	wire _w37633_ ;
	wire _w37632_ ;
	wire _w37631_ ;
	wire _w37630_ ;
	wire _w37629_ ;
	wire _w37628_ ;
	wire _w37627_ ;
	wire _w37626_ ;
	wire _w37625_ ;
	wire _w37624_ ;
	wire _w37623_ ;
	wire _w37622_ ;
	wire _w37621_ ;
	wire _w37620_ ;
	wire _w37619_ ;
	wire _w37618_ ;
	wire _w37617_ ;
	wire _w37616_ ;
	wire _w37615_ ;
	wire _w37614_ ;
	wire _w37613_ ;
	wire _w37612_ ;
	wire _w37611_ ;
	wire _w37610_ ;
	wire _w37609_ ;
	wire _w37608_ ;
	wire _w37607_ ;
	wire _w37606_ ;
	wire _w37605_ ;
	wire _w37604_ ;
	wire _w37603_ ;
	wire _w37602_ ;
	wire _w37601_ ;
	wire _w37600_ ;
	wire _w37599_ ;
	wire _w37598_ ;
	wire _w37597_ ;
	wire _w37596_ ;
	wire _w37595_ ;
	wire _w37594_ ;
	wire _w37593_ ;
	wire _w37592_ ;
	wire _w37591_ ;
	wire _w37590_ ;
	wire _w37589_ ;
	wire _w37588_ ;
	wire _w37587_ ;
	wire _w37586_ ;
	wire _w37585_ ;
	wire _w37584_ ;
	wire _w37583_ ;
	wire _w37582_ ;
	wire _w37581_ ;
	wire _w37580_ ;
	wire _w37579_ ;
	wire _w37578_ ;
	wire _w37577_ ;
	wire _w37576_ ;
	wire _w37575_ ;
	wire _w37574_ ;
	wire _w37573_ ;
	wire _w37572_ ;
	wire _w37571_ ;
	wire _w37570_ ;
	wire _w37569_ ;
	wire _w37568_ ;
	wire _w37567_ ;
	wire _w37566_ ;
	wire _w37565_ ;
	wire _w37564_ ;
	wire _w37563_ ;
	wire _w37562_ ;
	wire _w37561_ ;
	wire _w37560_ ;
	wire _w37559_ ;
	wire _w37558_ ;
	wire _w37557_ ;
	wire _w37556_ ;
	wire _w37555_ ;
	wire _w37554_ ;
	wire _w37553_ ;
	wire _w37552_ ;
	wire _w37551_ ;
	wire _w37550_ ;
	wire _w37549_ ;
	wire _w37548_ ;
	wire _w37547_ ;
	wire _w37546_ ;
	wire _w37545_ ;
	wire _w37544_ ;
	wire _w37543_ ;
	wire _w37542_ ;
	wire _w37541_ ;
	wire _w37540_ ;
	wire _w37539_ ;
	wire _w37538_ ;
	wire _w37537_ ;
	wire _w37536_ ;
	wire _w37535_ ;
	wire _w37534_ ;
	wire _w37533_ ;
	wire _w37532_ ;
	wire _w37531_ ;
	wire _w37530_ ;
	wire _w37529_ ;
	wire _w37528_ ;
	wire _w37527_ ;
	wire _w37526_ ;
	wire _w37525_ ;
	wire _w37524_ ;
	wire _w37523_ ;
	wire _w37522_ ;
	wire _w37521_ ;
	wire _w37520_ ;
	wire _w37519_ ;
	wire _w37518_ ;
	wire _w37517_ ;
	wire _w37516_ ;
	wire _w37515_ ;
	wire _w37514_ ;
	wire _w37513_ ;
	wire _w37512_ ;
	wire _w37511_ ;
	wire _w37510_ ;
	wire _w37509_ ;
	wire _w37508_ ;
	wire _w37507_ ;
	wire _w37506_ ;
	wire _w37505_ ;
	wire _w37504_ ;
	wire _w37503_ ;
	wire _w37502_ ;
	wire _w37501_ ;
	wire _w37500_ ;
	wire _w37499_ ;
	wire _w37498_ ;
	wire _w37497_ ;
	wire _w37496_ ;
	wire _w37495_ ;
	wire _w37494_ ;
	wire _w37493_ ;
	wire _w37492_ ;
	wire _w37491_ ;
	wire _w37490_ ;
	wire _w37489_ ;
	wire _w37488_ ;
	wire _w37487_ ;
	wire _w37486_ ;
	wire _w37485_ ;
	wire _w37484_ ;
	wire _w37483_ ;
	wire _w37482_ ;
	wire _w37481_ ;
	wire _w37480_ ;
	wire _w37479_ ;
	wire _w37478_ ;
	wire _w37477_ ;
	wire _w37476_ ;
	wire _w37475_ ;
	wire _w37474_ ;
	wire _w37473_ ;
	wire _w37472_ ;
	wire _w37471_ ;
	wire _w37470_ ;
	wire _w37469_ ;
	wire _w37468_ ;
	wire _w37467_ ;
	wire _w37466_ ;
	wire _w37465_ ;
	wire _w37464_ ;
	wire _w37463_ ;
	wire _w37462_ ;
	wire _w37461_ ;
	wire _w37460_ ;
	wire _w37459_ ;
	wire _w37458_ ;
	wire _w37457_ ;
	wire _w37456_ ;
	wire _w37455_ ;
	wire _w37454_ ;
	wire _w37453_ ;
	wire _w37452_ ;
	wire _w37451_ ;
	wire _w37450_ ;
	wire _w37449_ ;
	wire _w37448_ ;
	wire _w37447_ ;
	wire _w37446_ ;
	wire _w37445_ ;
	wire _w37444_ ;
	wire _w37443_ ;
	wire _w37442_ ;
	wire _w37441_ ;
	wire _w37440_ ;
	wire _w37439_ ;
	wire _w37438_ ;
	wire _w37437_ ;
	wire _w37436_ ;
	wire _w37435_ ;
	wire _w37434_ ;
	wire _w37433_ ;
	wire _w37432_ ;
	wire _w37431_ ;
	wire _w37430_ ;
	wire _w37429_ ;
	wire _w37428_ ;
	wire _w37427_ ;
	wire _w37426_ ;
	wire _w37425_ ;
	wire _w37424_ ;
	wire _w37423_ ;
	wire _w37422_ ;
	wire _w37421_ ;
	wire _w37420_ ;
	wire _w37419_ ;
	wire _w37418_ ;
	wire _w37417_ ;
	wire _w37416_ ;
	wire _w37415_ ;
	wire _w37414_ ;
	wire _w37413_ ;
	wire _w37412_ ;
	wire _w37411_ ;
	wire _w37410_ ;
	wire _w37409_ ;
	wire _w37408_ ;
	wire _w37407_ ;
	wire _w37406_ ;
	wire _w37405_ ;
	wire _w37404_ ;
	wire _w37403_ ;
	wire _w37402_ ;
	wire _w37401_ ;
	wire _w37400_ ;
	wire _w37399_ ;
	wire _w37398_ ;
	wire _w37397_ ;
	wire _w37396_ ;
	wire _w37395_ ;
	wire _w37394_ ;
	wire _w37393_ ;
	wire _w37392_ ;
	wire _w37391_ ;
	wire _w37390_ ;
	wire _w37389_ ;
	wire _w37388_ ;
	wire _w37387_ ;
	wire _w37386_ ;
	wire _w37385_ ;
	wire _w37384_ ;
	wire _w37383_ ;
	wire _w37382_ ;
	wire _w37381_ ;
	wire _w37380_ ;
	wire _w37379_ ;
	wire _w37378_ ;
	wire _w37377_ ;
	wire _w37376_ ;
	wire _w37375_ ;
	wire _w37374_ ;
	wire _w37373_ ;
	wire _w37372_ ;
	wire _w37371_ ;
	wire _w37370_ ;
	wire _w37369_ ;
	wire _w37368_ ;
	wire _w37367_ ;
	wire _w37366_ ;
	wire _w37365_ ;
	wire _w37364_ ;
	wire _w37363_ ;
	wire _w37362_ ;
	wire _w37361_ ;
	wire _w37360_ ;
	wire _w37359_ ;
	wire _w37358_ ;
	wire _w37357_ ;
	wire _w37356_ ;
	wire _w37355_ ;
	wire _w37354_ ;
	wire _w37353_ ;
	wire _w37352_ ;
	wire _w37351_ ;
	wire _w37350_ ;
	wire _w37349_ ;
	wire _w37348_ ;
	wire _w37347_ ;
	wire _w37346_ ;
	wire _w37345_ ;
	wire _w37344_ ;
	wire _w37343_ ;
	wire _w37342_ ;
	wire _w37341_ ;
	wire _w37340_ ;
	wire _w37339_ ;
	wire _w37338_ ;
	wire _w37337_ ;
	wire _w37336_ ;
	wire _w37335_ ;
	wire _w37334_ ;
	wire _w37333_ ;
	wire _w37332_ ;
	wire _w37331_ ;
	wire _w37330_ ;
	wire _w37329_ ;
	wire _w37328_ ;
	wire _w37327_ ;
	wire _w37326_ ;
	wire _w37325_ ;
	wire _w37324_ ;
	wire _w37323_ ;
	wire _w37322_ ;
	wire _w37321_ ;
	wire _w37320_ ;
	wire _w37319_ ;
	wire _w37318_ ;
	wire _w37317_ ;
	wire _w37316_ ;
	wire _w37315_ ;
	wire _w37314_ ;
	wire _w37313_ ;
	wire _w37312_ ;
	wire _w37311_ ;
	wire _w37310_ ;
	wire _w37309_ ;
	wire _w37308_ ;
	wire _w37307_ ;
	wire _w37306_ ;
	wire _w37305_ ;
	wire _w37304_ ;
	wire _w37303_ ;
	wire _w37302_ ;
	wire _w37301_ ;
	wire _w37300_ ;
	wire _w37299_ ;
	wire _w37298_ ;
	wire _w37297_ ;
	wire _w37296_ ;
	wire _w37295_ ;
	wire _w37294_ ;
	wire _w37293_ ;
	wire _w37292_ ;
	wire _w37291_ ;
	wire _w37290_ ;
	wire _w37289_ ;
	wire _w37288_ ;
	wire _w37287_ ;
	wire _w37286_ ;
	wire _w37285_ ;
	wire _w37284_ ;
	wire _w37283_ ;
	wire _w37282_ ;
	wire _w37281_ ;
	wire _w37280_ ;
	wire _w37279_ ;
	wire _w37278_ ;
	wire _w37277_ ;
	wire _w37276_ ;
	wire _w37275_ ;
	wire _w37274_ ;
	wire _w37273_ ;
	wire _w37272_ ;
	wire _w37271_ ;
	wire _w37270_ ;
	wire _w37269_ ;
	wire _w37268_ ;
	wire _w37267_ ;
	wire _w37266_ ;
	wire _w37265_ ;
	wire _w37264_ ;
	wire _w37263_ ;
	wire _w37262_ ;
	wire _w37261_ ;
	wire _w37260_ ;
	wire _w37259_ ;
	wire _w37258_ ;
	wire _w37257_ ;
	wire _w37256_ ;
	wire _w37255_ ;
	wire _w37254_ ;
	wire _w37253_ ;
	wire _w37252_ ;
	wire _w37251_ ;
	wire _w37250_ ;
	wire _w37249_ ;
	wire _w37248_ ;
	wire _w37247_ ;
	wire _w37246_ ;
	wire _w37245_ ;
	wire _w37244_ ;
	wire _w37243_ ;
	wire _w37242_ ;
	wire _w37241_ ;
	wire _w37240_ ;
	wire _w37239_ ;
	wire _w37238_ ;
	wire _w37237_ ;
	wire _w37236_ ;
	wire _w37235_ ;
	wire _w37234_ ;
	wire _w37233_ ;
	wire _w37232_ ;
	wire _w37231_ ;
	wire _w37230_ ;
	wire _w37229_ ;
	wire _w37228_ ;
	wire _w37227_ ;
	wire _w37226_ ;
	wire _w37225_ ;
	wire _w37224_ ;
	wire _w37223_ ;
	wire _w37222_ ;
	wire _w37221_ ;
	wire _w37220_ ;
	wire _w37219_ ;
	wire _w37218_ ;
	wire _w37217_ ;
	wire _w37216_ ;
	wire _w37215_ ;
	wire _w37214_ ;
	wire _w37213_ ;
	wire _w37212_ ;
	wire _w37211_ ;
	wire _w37210_ ;
	wire _w37209_ ;
	wire _w37208_ ;
	wire _w37207_ ;
	wire _w37206_ ;
	wire _w37205_ ;
	wire _w37204_ ;
	wire _w37203_ ;
	wire _w37202_ ;
	wire _w37201_ ;
	wire _w37200_ ;
	wire _w37199_ ;
	wire _w37198_ ;
	wire _w37197_ ;
	wire _w37196_ ;
	wire _w37195_ ;
	wire _w37194_ ;
	wire _w37193_ ;
	wire _w37192_ ;
	wire _w37191_ ;
	wire _w37190_ ;
	wire _w37189_ ;
	wire _w37188_ ;
	wire _w37187_ ;
	wire _w37186_ ;
	wire _w37185_ ;
	wire _w37184_ ;
	wire _w37183_ ;
	wire _w37182_ ;
	wire _w37181_ ;
	wire _w37180_ ;
	wire _w37179_ ;
	wire _w37178_ ;
	wire _w37177_ ;
	wire _w37176_ ;
	wire _w37175_ ;
	wire _w37174_ ;
	wire _w37173_ ;
	wire _w37172_ ;
	wire _w37171_ ;
	wire _w37170_ ;
	wire _w37169_ ;
	wire _w37168_ ;
	wire _w37167_ ;
	wire _w37166_ ;
	wire _w37165_ ;
	wire _w37164_ ;
	wire _w37163_ ;
	wire _w37162_ ;
	wire _w37161_ ;
	wire _w37160_ ;
	wire _w37159_ ;
	wire _w37158_ ;
	wire _w37157_ ;
	wire _w37156_ ;
	wire _w37155_ ;
	wire _w37154_ ;
	wire _w37153_ ;
	wire _w37152_ ;
	wire _w37151_ ;
	wire _w37150_ ;
	wire _w37149_ ;
	wire _w37148_ ;
	wire _w37147_ ;
	wire _w37146_ ;
	wire _w37145_ ;
	wire _w37144_ ;
	wire _w37143_ ;
	wire _w37142_ ;
	wire _w37141_ ;
	wire _w37140_ ;
	wire _w37139_ ;
	wire _w37138_ ;
	wire _w37137_ ;
	wire _w37136_ ;
	wire _w37135_ ;
	wire _w37134_ ;
	wire _w37133_ ;
	wire _w37132_ ;
	wire _w37131_ ;
	wire _w37130_ ;
	wire _w37129_ ;
	wire _w37128_ ;
	wire _w37127_ ;
	wire _w37126_ ;
	wire _w37125_ ;
	wire _w37124_ ;
	wire _w37123_ ;
	wire _w37122_ ;
	wire _w37121_ ;
	wire _w37120_ ;
	wire _w37119_ ;
	wire _w37118_ ;
	wire _w37117_ ;
	wire _w37116_ ;
	wire _w37115_ ;
	wire _w37114_ ;
	wire _w37113_ ;
	wire _w37112_ ;
	wire _w37111_ ;
	wire _w37110_ ;
	wire _w37109_ ;
	wire _w37108_ ;
	wire _w37107_ ;
	wire _w37106_ ;
	wire _w37105_ ;
	wire _w37104_ ;
	wire _w37103_ ;
	wire _w37102_ ;
	wire _w37101_ ;
	wire _w37100_ ;
	wire _w37099_ ;
	wire _w37098_ ;
	wire _w37097_ ;
	wire _w37096_ ;
	wire _w37095_ ;
	wire _w37094_ ;
	wire _w37093_ ;
	wire _w37092_ ;
	wire _w37091_ ;
	wire _w37090_ ;
	wire _w37089_ ;
	wire _w37088_ ;
	wire _w37087_ ;
	wire _w37086_ ;
	wire _w37085_ ;
	wire _w37084_ ;
	wire _w37083_ ;
	wire _w37082_ ;
	wire _w37081_ ;
	wire _w37080_ ;
	wire _w37079_ ;
	wire _w37078_ ;
	wire _w37077_ ;
	wire _w37076_ ;
	wire _w37075_ ;
	wire _w37074_ ;
	wire _w37073_ ;
	wire _w37072_ ;
	wire _w37071_ ;
	wire _w37070_ ;
	wire _w37069_ ;
	wire _w37068_ ;
	wire _w37067_ ;
	wire _w37066_ ;
	wire _w37065_ ;
	wire _w37064_ ;
	wire _w37063_ ;
	wire _w37062_ ;
	wire _w37061_ ;
	wire _w37060_ ;
	wire _w37059_ ;
	wire _w37058_ ;
	wire _w37057_ ;
	wire _w37056_ ;
	wire _w37055_ ;
	wire _w37054_ ;
	wire _w37053_ ;
	wire _w37052_ ;
	wire _w37051_ ;
	wire _w37050_ ;
	wire _w37049_ ;
	wire _w37048_ ;
	wire _w37047_ ;
	wire _w37046_ ;
	wire _w37045_ ;
	wire _w37044_ ;
	wire _w37043_ ;
	wire _w37042_ ;
	wire _w37041_ ;
	wire _w37040_ ;
	wire _w37039_ ;
	wire _w37038_ ;
	wire _w37037_ ;
	wire _w37036_ ;
	wire _w37035_ ;
	wire _w37034_ ;
	wire _w37033_ ;
	wire _w37032_ ;
	wire _w37031_ ;
	wire _w37030_ ;
	wire _w37029_ ;
	wire _w37028_ ;
	wire _w37027_ ;
	wire _w37026_ ;
	wire _w37025_ ;
	wire _w37024_ ;
	wire _w37023_ ;
	wire _w37022_ ;
	wire _w37021_ ;
	wire _w37020_ ;
	wire _w37019_ ;
	wire _w37018_ ;
	wire _w37017_ ;
	wire _w37016_ ;
	wire _w37015_ ;
	wire _w37014_ ;
	wire _w37013_ ;
	wire _w37012_ ;
	wire _w37011_ ;
	wire _w37010_ ;
	wire _w37009_ ;
	wire _w37008_ ;
	wire _w37007_ ;
	wire _w37006_ ;
	wire _w37005_ ;
	wire _w37004_ ;
	wire _w37003_ ;
	wire _w37002_ ;
	wire _w37001_ ;
	wire _w37000_ ;
	wire _w36999_ ;
	wire _w36998_ ;
	wire _w36997_ ;
	wire _w36996_ ;
	wire _w36995_ ;
	wire _w36994_ ;
	wire _w36993_ ;
	wire _w36992_ ;
	wire _w36991_ ;
	wire _w36990_ ;
	wire _w36989_ ;
	wire _w36988_ ;
	wire _w36987_ ;
	wire _w36986_ ;
	wire _w36985_ ;
	wire _w36984_ ;
	wire _w36983_ ;
	wire _w36982_ ;
	wire _w36981_ ;
	wire _w36980_ ;
	wire _w36979_ ;
	wire _w36978_ ;
	wire _w36977_ ;
	wire _w36976_ ;
	wire _w36975_ ;
	wire _w36974_ ;
	wire _w36973_ ;
	wire _w36972_ ;
	wire _w36971_ ;
	wire _w36970_ ;
	wire _w36969_ ;
	wire _w36968_ ;
	wire _w36967_ ;
	wire _w36966_ ;
	wire _w36965_ ;
	wire _w36964_ ;
	wire _w36963_ ;
	wire _w36962_ ;
	wire _w36961_ ;
	wire _w36960_ ;
	wire _w36959_ ;
	wire _w36958_ ;
	wire _w36957_ ;
	wire _w36956_ ;
	wire _w36955_ ;
	wire _w36954_ ;
	wire _w36953_ ;
	wire _w36952_ ;
	wire _w36951_ ;
	wire _w36950_ ;
	wire _w36949_ ;
	wire _w36948_ ;
	wire _w36947_ ;
	wire _w36946_ ;
	wire _w36945_ ;
	wire _w36944_ ;
	wire _w36943_ ;
	wire _w36942_ ;
	wire _w36941_ ;
	wire _w36940_ ;
	wire _w36939_ ;
	wire _w36938_ ;
	wire _w36937_ ;
	wire _w36936_ ;
	wire _w36935_ ;
	wire _w36934_ ;
	wire _w36933_ ;
	wire _w36932_ ;
	wire _w36931_ ;
	wire _w36930_ ;
	wire _w36929_ ;
	wire _w36928_ ;
	wire _w36927_ ;
	wire _w36926_ ;
	wire _w36925_ ;
	wire _w36924_ ;
	wire _w36923_ ;
	wire _w36922_ ;
	wire _w36921_ ;
	wire _w36920_ ;
	wire _w36919_ ;
	wire _w36918_ ;
	wire _w36917_ ;
	wire _w36916_ ;
	wire _w36915_ ;
	wire _w36914_ ;
	wire _w36913_ ;
	wire _w36912_ ;
	wire _w36911_ ;
	wire _w36910_ ;
	wire _w36909_ ;
	wire _w36908_ ;
	wire _w36907_ ;
	wire _w36906_ ;
	wire _w36905_ ;
	wire _w36904_ ;
	wire _w36903_ ;
	wire _w36902_ ;
	wire _w36901_ ;
	wire _w36900_ ;
	wire _w36899_ ;
	wire _w36898_ ;
	wire _w36897_ ;
	wire _w36896_ ;
	wire _w36895_ ;
	wire _w36894_ ;
	wire _w36893_ ;
	wire _w36892_ ;
	wire _w36891_ ;
	wire _w36890_ ;
	wire _w36889_ ;
	wire _w36888_ ;
	wire _w36887_ ;
	wire _w36886_ ;
	wire _w36885_ ;
	wire _w36884_ ;
	wire _w36883_ ;
	wire _w36882_ ;
	wire _w36881_ ;
	wire _w36880_ ;
	wire _w36879_ ;
	wire _w36878_ ;
	wire _w36877_ ;
	wire _w36876_ ;
	wire _w36875_ ;
	wire _w36874_ ;
	wire _w36873_ ;
	wire _w36872_ ;
	wire _w36871_ ;
	wire _w36870_ ;
	wire _w36869_ ;
	wire _w36868_ ;
	wire _w36867_ ;
	wire _w36866_ ;
	wire _w36865_ ;
	wire _w36864_ ;
	wire _w36863_ ;
	wire _w36862_ ;
	wire _w36861_ ;
	wire _w36860_ ;
	wire _w36859_ ;
	wire _w36858_ ;
	wire _w36857_ ;
	wire _w36856_ ;
	wire _w36855_ ;
	wire _w36854_ ;
	wire _w36853_ ;
	wire _w36852_ ;
	wire _w36851_ ;
	wire _w36850_ ;
	wire _w36849_ ;
	wire _w36848_ ;
	wire _w36847_ ;
	wire _w36846_ ;
	wire _w36845_ ;
	wire _w36844_ ;
	wire _w36843_ ;
	wire _w36842_ ;
	wire _w36841_ ;
	wire _w36840_ ;
	wire _w36839_ ;
	wire _w36838_ ;
	wire _w36837_ ;
	wire _w36836_ ;
	wire _w36835_ ;
	wire _w36834_ ;
	wire _w36833_ ;
	wire _w36832_ ;
	wire _w36831_ ;
	wire _w36830_ ;
	wire _w36829_ ;
	wire _w36828_ ;
	wire _w36827_ ;
	wire _w36826_ ;
	wire _w36825_ ;
	wire _w36824_ ;
	wire _w36823_ ;
	wire _w36822_ ;
	wire _w36821_ ;
	wire _w36820_ ;
	wire _w36819_ ;
	wire _w36818_ ;
	wire _w36817_ ;
	wire _w36816_ ;
	wire _w36815_ ;
	wire _w36814_ ;
	wire _w36813_ ;
	wire _w36812_ ;
	wire _w36811_ ;
	wire _w36810_ ;
	wire _w36809_ ;
	wire _w36808_ ;
	wire _w36807_ ;
	wire _w36806_ ;
	wire _w36805_ ;
	wire _w36804_ ;
	wire _w36803_ ;
	wire _w36802_ ;
	wire _w36801_ ;
	wire _w36800_ ;
	wire _w36799_ ;
	wire _w36798_ ;
	wire _w36797_ ;
	wire _w36796_ ;
	wire _w36795_ ;
	wire _w36794_ ;
	wire _w36793_ ;
	wire _w36792_ ;
	wire _w36791_ ;
	wire _w36790_ ;
	wire _w36789_ ;
	wire _w36788_ ;
	wire _w36787_ ;
	wire _w36786_ ;
	wire _w36785_ ;
	wire _w36784_ ;
	wire _w36783_ ;
	wire _w36782_ ;
	wire _w36781_ ;
	wire _w36780_ ;
	wire _w36779_ ;
	wire _w36778_ ;
	wire _w36777_ ;
	wire _w36776_ ;
	wire _w36775_ ;
	wire _w36774_ ;
	wire _w36773_ ;
	wire _w36772_ ;
	wire _w36771_ ;
	wire _w36770_ ;
	wire _w36769_ ;
	wire _w36768_ ;
	wire _w36767_ ;
	wire _w36766_ ;
	wire _w36765_ ;
	wire _w36764_ ;
	wire _w36763_ ;
	wire _w36762_ ;
	wire _w36761_ ;
	wire _w36760_ ;
	wire _w36759_ ;
	wire _w36758_ ;
	wire _w36757_ ;
	wire _w36756_ ;
	wire _w36755_ ;
	wire _w36754_ ;
	wire _w36753_ ;
	wire _w36752_ ;
	wire _w36751_ ;
	wire _w36750_ ;
	wire _w36749_ ;
	wire _w36748_ ;
	wire _w36747_ ;
	wire _w36746_ ;
	wire _w36745_ ;
	wire _w36744_ ;
	wire _w36743_ ;
	wire _w36742_ ;
	wire _w36741_ ;
	wire _w36740_ ;
	wire _w36739_ ;
	wire _w36738_ ;
	wire _w36737_ ;
	wire _w36736_ ;
	wire _w36735_ ;
	wire _w36734_ ;
	wire _w36733_ ;
	wire _w36732_ ;
	wire _w36731_ ;
	wire _w36730_ ;
	wire _w36729_ ;
	wire _w36728_ ;
	wire _w36727_ ;
	wire _w36726_ ;
	wire _w36725_ ;
	wire _w36724_ ;
	wire _w36723_ ;
	wire _w36722_ ;
	wire _w36721_ ;
	wire _w36720_ ;
	wire _w36719_ ;
	wire _w36718_ ;
	wire _w36717_ ;
	wire _w36716_ ;
	wire _w36715_ ;
	wire _w36714_ ;
	wire _w36713_ ;
	wire _w36712_ ;
	wire _w36711_ ;
	wire _w36710_ ;
	wire _w36709_ ;
	wire _w36708_ ;
	wire _w36707_ ;
	wire _w36706_ ;
	wire _w36705_ ;
	wire _w36704_ ;
	wire _w36703_ ;
	wire _w36702_ ;
	wire _w36701_ ;
	wire _w36700_ ;
	wire _w36699_ ;
	wire _w36698_ ;
	wire _w36697_ ;
	wire _w36696_ ;
	wire _w36695_ ;
	wire _w36694_ ;
	wire _w36693_ ;
	wire _w36692_ ;
	wire _w36691_ ;
	wire _w36690_ ;
	wire _w36689_ ;
	wire _w36688_ ;
	wire _w36687_ ;
	wire _w36686_ ;
	wire _w36685_ ;
	wire _w36684_ ;
	wire _w36683_ ;
	wire _w36682_ ;
	wire _w36681_ ;
	wire _w36680_ ;
	wire _w36679_ ;
	wire _w36678_ ;
	wire _w36677_ ;
	wire _w36676_ ;
	wire _w36675_ ;
	wire _w36674_ ;
	wire _w36673_ ;
	wire _w36672_ ;
	wire _w36671_ ;
	wire _w36670_ ;
	wire _w36669_ ;
	wire _w36668_ ;
	wire _w36667_ ;
	wire _w36666_ ;
	wire _w36665_ ;
	wire _w36664_ ;
	wire _w36663_ ;
	wire _w36662_ ;
	wire _w36661_ ;
	wire _w36660_ ;
	wire _w36659_ ;
	wire _w36658_ ;
	wire _w36657_ ;
	wire _w36656_ ;
	wire _w36655_ ;
	wire _w36654_ ;
	wire _w36653_ ;
	wire _w36652_ ;
	wire _w36651_ ;
	wire _w36650_ ;
	wire _w36649_ ;
	wire _w36648_ ;
	wire _w36647_ ;
	wire _w36646_ ;
	wire _w36645_ ;
	wire _w36644_ ;
	wire _w36643_ ;
	wire _w36642_ ;
	wire _w36641_ ;
	wire _w36640_ ;
	wire _w36639_ ;
	wire _w36638_ ;
	wire _w36637_ ;
	wire _w36636_ ;
	wire _w36635_ ;
	wire _w36634_ ;
	wire _w36633_ ;
	wire _w36632_ ;
	wire _w36631_ ;
	wire _w36630_ ;
	wire _w36629_ ;
	wire _w36628_ ;
	wire _w36627_ ;
	wire _w36626_ ;
	wire _w36625_ ;
	wire _w36624_ ;
	wire _w36623_ ;
	wire _w36622_ ;
	wire _w36621_ ;
	wire _w36620_ ;
	wire _w36619_ ;
	wire _w36618_ ;
	wire _w36617_ ;
	wire _w36616_ ;
	wire _w36615_ ;
	wire _w36614_ ;
	wire _w36613_ ;
	wire _w36612_ ;
	wire _w36611_ ;
	wire _w36610_ ;
	wire _w36609_ ;
	wire _w36608_ ;
	wire _w36607_ ;
	wire _w36606_ ;
	wire _w36605_ ;
	wire _w36604_ ;
	wire _w36603_ ;
	wire _w36602_ ;
	wire _w36601_ ;
	wire _w36600_ ;
	wire _w36599_ ;
	wire _w36598_ ;
	wire _w36597_ ;
	wire _w36596_ ;
	wire _w36595_ ;
	wire _w36594_ ;
	wire _w36593_ ;
	wire _w36592_ ;
	wire _w36591_ ;
	wire _w36590_ ;
	wire _w36589_ ;
	wire _w36588_ ;
	wire _w36587_ ;
	wire _w36586_ ;
	wire _w36585_ ;
	wire _w36584_ ;
	wire _w36583_ ;
	wire _w36582_ ;
	wire _w36581_ ;
	wire _w36580_ ;
	wire _w36579_ ;
	wire _w36578_ ;
	wire _w36577_ ;
	wire _w36576_ ;
	wire _w36575_ ;
	wire _w36574_ ;
	wire _w36573_ ;
	wire _w36572_ ;
	wire _w36571_ ;
	wire _w36570_ ;
	wire _w36569_ ;
	wire _w36568_ ;
	wire _w36567_ ;
	wire _w36566_ ;
	wire _w36565_ ;
	wire _w36564_ ;
	wire _w36563_ ;
	wire _w36562_ ;
	wire _w36561_ ;
	wire _w36560_ ;
	wire _w36559_ ;
	wire _w36558_ ;
	wire _w36557_ ;
	wire _w36556_ ;
	wire _w36555_ ;
	wire _w36554_ ;
	wire _w36553_ ;
	wire _w36552_ ;
	wire _w36551_ ;
	wire _w36550_ ;
	wire _w36549_ ;
	wire _w36548_ ;
	wire _w36547_ ;
	wire _w36546_ ;
	wire _w36545_ ;
	wire _w36544_ ;
	wire _w36543_ ;
	wire _w36542_ ;
	wire _w36541_ ;
	wire _w36540_ ;
	wire _w36539_ ;
	wire _w36538_ ;
	wire _w36537_ ;
	wire _w36536_ ;
	wire _w36535_ ;
	wire _w36534_ ;
	wire _w36533_ ;
	wire _w36532_ ;
	wire _w36531_ ;
	wire _w36530_ ;
	wire _w36529_ ;
	wire _w36528_ ;
	wire _w36527_ ;
	wire _w36526_ ;
	wire _w36525_ ;
	wire _w36524_ ;
	wire _w36523_ ;
	wire _w36522_ ;
	wire _w36521_ ;
	wire _w36520_ ;
	wire _w36519_ ;
	wire _w36518_ ;
	wire _w36517_ ;
	wire _w36516_ ;
	wire _w36515_ ;
	wire _w36514_ ;
	wire _w36513_ ;
	wire _w36512_ ;
	wire _w36511_ ;
	wire _w36510_ ;
	wire _w36509_ ;
	wire _w36508_ ;
	wire _w36507_ ;
	wire _w36506_ ;
	wire _w36505_ ;
	wire _w36504_ ;
	wire _w36503_ ;
	wire _w36502_ ;
	wire _w36501_ ;
	wire _w36500_ ;
	wire _w36499_ ;
	wire _w36498_ ;
	wire _w36497_ ;
	wire _w36496_ ;
	wire _w36495_ ;
	wire _w36494_ ;
	wire _w36493_ ;
	wire _w36492_ ;
	wire _w36491_ ;
	wire _w36490_ ;
	wire _w36489_ ;
	wire _w36488_ ;
	wire _w36487_ ;
	wire _w36486_ ;
	wire _w36485_ ;
	wire _w36484_ ;
	wire _w36483_ ;
	wire _w36482_ ;
	wire _w36481_ ;
	wire _w36480_ ;
	wire _w36479_ ;
	wire _w36478_ ;
	wire _w36477_ ;
	wire _w36476_ ;
	wire _w36475_ ;
	wire _w36474_ ;
	wire _w36473_ ;
	wire _w36472_ ;
	wire _w36471_ ;
	wire _w36470_ ;
	wire _w36469_ ;
	wire _w36468_ ;
	wire _w36467_ ;
	wire _w36466_ ;
	wire _w36465_ ;
	wire _w36464_ ;
	wire _w36463_ ;
	wire _w36462_ ;
	wire _w36461_ ;
	wire _w36460_ ;
	wire _w36459_ ;
	wire _w36458_ ;
	wire _w36457_ ;
	wire _w36456_ ;
	wire _w36455_ ;
	wire _w36454_ ;
	wire _w36453_ ;
	wire _w36452_ ;
	wire _w36451_ ;
	wire _w36450_ ;
	wire _w36449_ ;
	wire _w36448_ ;
	wire _w36447_ ;
	wire _w36446_ ;
	wire _w36445_ ;
	wire _w36444_ ;
	wire _w36443_ ;
	wire _w36442_ ;
	wire _w36441_ ;
	wire _w36440_ ;
	wire _w36439_ ;
	wire _w36438_ ;
	wire _w36437_ ;
	wire _w36436_ ;
	wire _w36435_ ;
	wire _w36434_ ;
	wire _w36433_ ;
	wire _w36432_ ;
	wire _w36431_ ;
	wire _w36430_ ;
	wire _w36429_ ;
	wire _w36428_ ;
	wire _w36427_ ;
	wire _w36426_ ;
	wire _w36425_ ;
	wire _w36424_ ;
	wire _w36423_ ;
	wire _w36422_ ;
	wire _w36421_ ;
	wire _w36420_ ;
	wire _w36419_ ;
	wire _w36418_ ;
	wire _w36417_ ;
	wire _w36416_ ;
	wire _w36415_ ;
	wire _w36414_ ;
	wire _w36413_ ;
	wire _w36412_ ;
	wire _w36411_ ;
	wire _w36410_ ;
	wire _w36409_ ;
	wire _w36408_ ;
	wire _w36407_ ;
	wire _w36406_ ;
	wire _w36405_ ;
	wire _w36404_ ;
	wire _w36403_ ;
	wire _w36402_ ;
	wire _w36401_ ;
	wire _w36400_ ;
	wire _w36399_ ;
	wire _w36398_ ;
	wire _w36397_ ;
	wire _w36396_ ;
	wire _w36395_ ;
	wire _w36394_ ;
	wire _w36393_ ;
	wire _w36392_ ;
	wire _w36391_ ;
	wire _w36390_ ;
	wire _w36389_ ;
	wire _w36388_ ;
	wire _w36387_ ;
	wire _w36386_ ;
	wire _w36385_ ;
	wire _w36384_ ;
	wire _w36383_ ;
	wire _w36382_ ;
	wire _w36381_ ;
	wire _w36380_ ;
	wire _w36379_ ;
	wire _w36378_ ;
	wire _w36377_ ;
	wire _w36376_ ;
	wire _w36375_ ;
	wire _w36374_ ;
	wire _w36373_ ;
	wire _w36372_ ;
	wire _w36371_ ;
	wire _w36370_ ;
	wire _w36369_ ;
	wire _w36368_ ;
	wire _w36367_ ;
	wire _w36366_ ;
	wire _w36365_ ;
	wire _w36364_ ;
	wire _w36363_ ;
	wire _w36362_ ;
	wire _w36361_ ;
	wire _w36360_ ;
	wire _w36359_ ;
	wire _w36358_ ;
	wire _w36357_ ;
	wire _w36356_ ;
	wire _w36355_ ;
	wire _w36354_ ;
	wire _w36353_ ;
	wire _w36352_ ;
	wire _w36351_ ;
	wire _w36350_ ;
	wire _w36349_ ;
	wire _w36348_ ;
	wire _w36347_ ;
	wire _w36346_ ;
	wire _w36345_ ;
	wire _w36344_ ;
	wire _w36343_ ;
	wire _w36342_ ;
	wire _w36341_ ;
	wire _w36340_ ;
	wire _w36339_ ;
	wire _w36338_ ;
	wire _w36337_ ;
	wire _w36336_ ;
	wire _w36335_ ;
	wire _w36334_ ;
	wire _w36333_ ;
	wire _w36332_ ;
	wire _w36331_ ;
	wire _w36330_ ;
	wire _w36329_ ;
	wire _w36328_ ;
	wire _w36327_ ;
	wire _w36326_ ;
	wire _w36325_ ;
	wire _w36324_ ;
	wire _w36323_ ;
	wire _w36322_ ;
	wire _w36321_ ;
	wire _w36320_ ;
	wire _w36319_ ;
	wire _w36318_ ;
	wire _w36317_ ;
	wire _w36316_ ;
	wire _w36315_ ;
	wire _w36314_ ;
	wire _w36313_ ;
	wire _w36312_ ;
	wire _w36311_ ;
	wire _w36310_ ;
	wire _w36309_ ;
	wire _w36308_ ;
	wire _w36307_ ;
	wire _w36306_ ;
	wire _w36305_ ;
	wire _w36304_ ;
	wire _w36303_ ;
	wire _w36302_ ;
	wire _w36301_ ;
	wire _w36300_ ;
	wire _w36299_ ;
	wire _w36298_ ;
	wire _w36297_ ;
	wire _w36296_ ;
	wire _w36295_ ;
	wire _w36294_ ;
	wire _w36293_ ;
	wire _w36292_ ;
	wire _w36291_ ;
	wire _w36290_ ;
	wire _w36289_ ;
	wire _w36288_ ;
	wire _w36287_ ;
	wire _w36286_ ;
	wire _w36285_ ;
	wire _w36284_ ;
	wire _w36283_ ;
	wire _w36282_ ;
	wire _w36281_ ;
	wire _w36280_ ;
	wire _w36279_ ;
	wire _w36278_ ;
	wire _w36277_ ;
	wire _w36276_ ;
	wire _w36275_ ;
	wire _w36274_ ;
	wire _w36273_ ;
	wire _w36272_ ;
	wire _w36271_ ;
	wire _w36270_ ;
	wire _w36269_ ;
	wire _w36268_ ;
	wire _w36267_ ;
	wire _w36266_ ;
	wire _w36265_ ;
	wire _w36264_ ;
	wire _w36263_ ;
	wire _w36262_ ;
	wire _w36261_ ;
	wire _w36260_ ;
	wire _w36259_ ;
	wire _w36258_ ;
	wire _w36257_ ;
	wire _w36256_ ;
	wire _w36255_ ;
	wire _w36254_ ;
	wire _w36253_ ;
	wire _w36252_ ;
	wire _w36251_ ;
	wire _w36250_ ;
	wire _w36249_ ;
	wire _w36248_ ;
	wire _w36247_ ;
	wire _w36246_ ;
	wire _w36245_ ;
	wire _w36244_ ;
	wire _w36243_ ;
	wire _w36242_ ;
	wire _w36241_ ;
	wire _w36240_ ;
	wire _w36239_ ;
	wire _w36238_ ;
	wire _w36237_ ;
	wire _w36236_ ;
	wire _w36235_ ;
	wire _w36234_ ;
	wire _w36233_ ;
	wire _w36232_ ;
	wire _w36231_ ;
	wire _w36230_ ;
	wire _w36229_ ;
	wire _w36228_ ;
	wire _w36227_ ;
	wire _w36226_ ;
	wire _w36225_ ;
	wire _w36224_ ;
	wire _w36223_ ;
	wire _w36222_ ;
	wire _w36221_ ;
	wire _w36220_ ;
	wire _w36219_ ;
	wire _w36218_ ;
	wire _w36217_ ;
	wire _w36216_ ;
	wire _w36215_ ;
	wire _w36214_ ;
	wire _w36213_ ;
	wire _w36212_ ;
	wire _w36211_ ;
	wire _w36210_ ;
	wire _w36209_ ;
	wire _w36208_ ;
	wire _w36207_ ;
	wire _w36206_ ;
	wire _w36205_ ;
	wire _w36204_ ;
	wire _w36203_ ;
	wire _w36202_ ;
	wire _w36201_ ;
	wire _w36200_ ;
	wire _w36199_ ;
	wire _w36198_ ;
	wire _w36197_ ;
	wire _w36196_ ;
	wire _w36195_ ;
	wire _w36194_ ;
	wire _w36193_ ;
	wire _w36192_ ;
	wire _w36191_ ;
	wire _w36190_ ;
	wire _w36189_ ;
	wire _w36188_ ;
	wire _w36187_ ;
	wire _w36186_ ;
	wire _w36185_ ;
	wire _w36184_ ;
	wire _w36183_ ;
	wire _w36182_ ;
	wire _w36181_ ;
	wire _w36180_ ;
	wire _w36179_ ;
	wire _w36178_ ;
	wire _w36177_ ;
	wire _w36176_ ;
	wire _w36175_ ;
	wire _w36174_ ;
	wire _w36173_ ;
	wire _w36172_ ;
	wire _w36171_ ;
	wire _w36170_ ;
	wire _w36169_ ;
	wire _w36168_ ;
	wire _w36167_ ;
	wire _w36166_ ;
	wire _w36165_ ;
	wire _w36164_ ;
	wire _w36163_ ;
	wire _w36162_ ;
	wire _w36161_ ;
	wire _w36160_ ;
	wire _w36159_ ;
	wire _w36158_ ;
	wire _w36157_ ;
	wire _w36156_ ;
	wire _w36155_ ;
	wire _w36154_ ;
	wire _w36153_ ;
	wire _w36152_ ;
	wire _w36151_ ;
	wire _w36150_ ;
	wire _w36149_ ;
	wire _w36148_ ;
	wire _w36147_ ;
	wire _w36146_ ;
	wire _w36145_ ;
	wire _w36144_ ;
	wire _w36143_ ;
	wire _w36142_ ;
	wire _w36141_ ;
	wire _w36140_ ;
	wire _w36139_ ;
	wire _w36138_ ;
	wire _w36137_ ;
	wire _w36136_ ;
	wire _w36135_ ;
	wire _w36134_ ;
	wire _w36133_ ;
	wire _w36132_ ;
	wire _w36131_ ;
	wire _w36130_ ;
	wire _w36129_ ;
	wire _w36128_ ;
	wire _w36127_ ;
	wire _w36126_ ;
	wire _w36125_ ;
	wire _w36124_ ;
	wire _w36123_ ;
	wire _w36122_ ;
	wire _w36121_ ;
	wire _w36120_ ;
	wire _w36119_ ;
	wire _w36118_ ;
	wire _w36117_ ;
	wire _w36116_ ;
	wire _w36115_ ;
	wire _w36114_ ;
	wire _w36113_ ;
	wire _w36112_ ;
	wire _w36111_ ;
	wire _w36110_ ;
	wire _w36109_ ;
	wire _w36108_ ;
	wire _w36107_ ;
	wire _w36106_ ;
	wire _w36105_ ;
	wire _w36104_ ;
	wire _w36103_ ;
	wire _w36102_ ;
	wire _w36101_ ;
	wire _w36100_ ;
	wire _w36099_ ;
	wire _w36098_ ;
	wire _w36097_ ;
	wire _w36096_ ;
	wire _w36095_ ;
	wire _w36094_ ;
	wire _w36093_ ;
	wire _w36092_ ;
	wire _w36091_ ;
	wire _w36090_ ;
	wire _w36089_ ;
	wire _w36088_ ;
	wire _w36087_ ;
	wire _w36086_ ;
	wire _w36085_ ;
	wire _w36084_ ;
	wire _w36083_ ;
	wire _w36082_ ;
	wire _w36081_ ;
	wire _w36080_ ;
	wire _w36079_ ;
	wire _w36078_ ;
	wire _w36077_ ;
	wire _w36076_ ;
	wire _w36075_ ;
	wire _w36074_ ;
	wire _w36073_ ;
	wire _w36072_ ;
	wire _w36071_ ;
	wire _w36070_ ;
	wire _w36069_ ;
	wire _w36068_ ;
	wire _w36067_ ;
	wire _w36066_ ;
	wire _w36065_ ;
	wire _w36064_ ;
	wire _w36063_ ;
	wire _w36062_ ;
	wire _w36061_ ;
	wire _w36060_ ;
	wire _w36059_ ;
	wire _w36058_ ;
	wire _w36057_ ;
	wire _w36056_ ;
	wire _w36055_ ;
	wire _w36054_ ;
	wire _w36053_ ;
	wire _w36052_ ;
	wire _w36051_ ;
	wire _w36050_ ;
	wire _w36049_ ;
	wire _w36048_ ;
	wire _w36047_ ;
	wire _w36046_ ;
	wire _w36045_ ;
	wire _w36044_ ;
	wire _w36043_ ;
	wire _w36042_ ;
	wire _w36041_ ;
	wire _w36040_ ;
	wire _w36039_ ;
	wire _w36038_ ;
	wire _w36037_ ;
	wire _w36036_ ;
	wire _w36035_ ;
	wire _w36034_ ;
	wire _w36033_ ;
	wire _w36032_ ;
	wire _w36031_ ;
	wire _w36030_ ;
	wire _w36029_ ;
	wire _w36028_ ;
	wire _w36027_ ;
	wire _w36026_ ;
	wire _w36025_ ;
	wire _w36024_ ;
	wire _w36023_ ;
	wire _w36022_ ;
	wire _w36021_ ;
	wire _w36020_ ;
	wire _w36019_ ;
	wire _w36018_ ;
	wire _w36017_ ;
	wire _w36016_ ;
	wire _w36015_ ;
	wire _w36014_ ;
	wire _w36013_ ;
	wire _w36012_ ;
	wire _w36011_ ;
	wire _w36010_ ;
	wire _w36009_ ;
	wire _w36008_ ;
	wire _w36007_ ;
	wire _w36006_ ;
	wire _w36005_ ;
	wire _w36004_ ;
	wire _w36003_ ;
	wire _w36002_ ;
	wire _w36001_ ;
	wire _w36000_ ;
	wire _w35999_ ;
	wire _w35998_ ;
	wire _w35997_ ;
	wire _w35996_ ;
	wire _w35995_ ;
	wire _w35994_ ;
	wire _w35993_ ;
	wire _w35992_ ;
	wire _w35991_ ;
	wire _w35990_ ;
	wire _w35989_ ;
	wire _w35988_ ;
	wire _w35987_ ;
	wire _w35986_ ;
	wire _w35985_ ;
	wire _w35984_ ;
	wire _w35983_ ;
	wire _w35982_ ;
	wire _w35981_ ;
	wire _w35980_ ;
	wire _w35979_ ;
	wire _w35978_ ;
	wire _w35977_ ;
	wire _w35976_ ;
	wire _w35975_ ;
	wire _w35974_ ;
	wire _w35973_ ;
	wire _w35972_ ;
	wire _w35971_ ;
	wire _w35970_ ;
	wire _w35969_ ;
	wire _w35968_ ;
	wire _w35967_ ;
	wire _w35966_ ;
	wire _w35965_ ;
	wire _w35964_ ;
	wire _w35963_ ;
	wire _w35962_ ;
	wire _w35961_ ;
	wire _w35960_ ;
	wire _w35959_ ;
	wire _w35958_ ;
	wire _w35957_ ;
	wire _w35956_ ;
	wire _w35955_ ;
	wire _w35954_ ;
	wire _w35953_ ;
	wire _w35952_ ;
	wire _w35951_ ;
	wire _w35950_ ;
	wire _w35949_ ;
	wire _w35948_ ;
	wire _w35947_ ;
	wire _w35946_ ;
	wire _w35945_ ;
	wire _w35944_ ;
	wire _w35943_ ;
	wire _w35942_ ;
	wire _w35941_ ;
	wire _w35940_ ;
	wire _w35939_ ;
	wire _w35938_ ;
	wire _w35937_ ;
	wire _w35936_ ;
	wire _w35935_ ;
	wire _w35934_ ;
	wire _w35933_ ;
	wire _w35932_ ;
	wire _w35931_ ;
	wire _w35930_ ;
	wire _w35929_ ;
	wire _w35928_ ;
	wire _w35927_ ;
	wire _w35926_ ;
	wire _w35925_ ;
	wire _w35924_ ;
	wire _w35923_ ;
	wire _w35922_ ;
	wire _w35921_ ;
	wire _w35920_ ;
	wire _w35919_ ;
	wire _w35918_ ;
	wire _w35917_ ;
	wire _w35916_ ;
	wire _w35915_ ;
	wire _w35914_ ;
	wire _w35913_ ;
	wire _w35912_ ;
	wire _w35911_ ;
	wire _w35910_ ;
	wire _w35909_ ;
	wire _w35908_ ;
	wire _w35907_ ;
	wire _w35906_ ;
	wire _w35905_ ;
	wire _w35904_ ;
	wire _w35903_ ;
	wire _w35902_ ;
	wire _w35901_ ;
	wire _w35900_ ;
	wire _w35899_ ;
	wire _w35898_ ;
	wire _w35897_ ;
	wire _w35896_ ;
	wire _w35895_ ;
	wire _w35894_ ;
	wire _w35893_ ;
	wire _w35892_ ;
	wire _w35891_ ;
	wire _w35890_ ;
	wire _w35889_ ;
	wire _w35888_ ;
	wire _w35887_ ;
	wire _w35886_ ;
	wire _w35885_ ;
	wire _w35884_ ;
	wire _w35883_ ;
	wire _w35882_ ;
	wire _w35881_ ;
	wire _w35880_ ;
	wire _w35879_ ;
	wire _w35878_ ;
	wire _w35877_ ;
	wire _w35876_ ;
	wire _w35875_ ;
	wire _w35874_ ;
	wire _w35873_ ;
	wire _w35872_ ;
	wire _w35871_ ;
	wire _w35870_ ;
	wire _w35869_ ;
	wire _w35868_ ;
	wire _w35867_ ;
	wire _w35866_ ;
	wire _w35865_ ;
	wire _w35864_ ;
	wire _w35863_ ;
	wire _w35862_ ;
	wire _w35861_ ;
	wire _w35860_ ;
	wire _w35859_ ;
	wire _w35858_ ;
	wire _w35857_ ;
	wire _w35856_ ;
	wire _w35855_ ;
	wire _w35854_ ;
	wire _w35853_ ;
	wire _w35852_ ;
	wire _w35851_ ;
	wire _w35850_ ;
	wire _w35849_ ;
	wire _w35848_ ;
	wire _w35847_ ;
	wire _w35846_ ;
	wire _w35845_ ;
	wire _w35844_ ;
	wire _w35843_ ;
	wire _w35842_ ;
	wire _w35841_ ;
	wire _w35840_ ;
	wire _w35839_ ;
	wire _w35838_ ;
	wire _w35837_ ;
	wire _w35836_ ;
	wire _w35835_ ;
	wire _w35834_ ;
	wire _w35833_ ;
	wire _w35832_ ;
	wire _w35831_ ;
	wire _w35830_ ;
	wire _w35829_ ;
	wire _w35828_ ;
	wire _w35827_ ;
	wire _w35826_ ;
	wire _w35825_ ;
	wire _w35824_ ;
	wire _w35823_ ;
	wire _w35822_ ;
	wire _w35821_ ;
	wire _w35820_ ;
	wire _w35819_ ;
	wire _w35818_ ;
	wire _w35817_ ;
	wire _w35816_ ;
	wire _w35815_ ;
	wire _w35814_ ;
	wire _w35813_ ;
	wire _w35812_ ;
	wire _w35811_ ;
	wire _w35810_ ;
	wire _w35809_ ;
	wire _w35808_ ;
	wire _w35807_ ;
	wire _w35806_ ;
	wire _w35805_ ;
	wire _w35804_ ;
	wire _w35803_ ;
	wire _w35802_ ;
	wire _w35801_ ;
	wire _w35800_ ;
	wire _w35799_ ;
	wire _w35798_ ;
	wire _w35797_ ;
	wire _w35796_ ;
	wire _w35795_ ;
	wire _w35794_ ;
	wire _w35793_ ;
	wire _w35792_ ;
	wire _w35791_ ;
	wire _w35790_ ;
	wire _w35789_ ;
	wire _w35788_ ;
	wire _w35787_ ;
	wire _w35786_ ;
	wire _w35785_ ;
	wire _w35784_ ;
	wire _w35783_ ;
	wire _w35782_ ;
	wire _w35781_ ;
	wire _w35780_ ;
	wire _w35779_ ;
	wire _w35778_ ;
	wire _w35777_ ;
	wire _w35776_ ;
	wire _w35775_ ;
	wire _w35774_ ;
	wire _w35773_ ;
	wire _w35772_ ;
	wire _w35771_ ;
	wire _w35770_ ;
	wire _w35769_ ;
	wire _w35768_ ;
	wire _w35767_ ;
	wire _w35766_ ;
	wire _w35765_ ;
	wire _w35764_ ;
	wire _w35763_ ;
	wire _w35762_ ;
	wire _w35761_ ;
	wire _w35760_ ;
	wire _w35759_ ;
	wire _w35758_ ;
	wire _w35757_ ;
	wire _w35756_ ;
	wire _w35755_ ;
	wire _w35754_ ;
	wire _w35753_ ;
	wire _w35752_ ;
	wire _w35751_ ;
	wire _w35750_ ;
	wire _w35749_ ;
	wire _w35748_ ;
	wire _w35747_ ;
	wire _w35746_ ;
	wire _w35745_ ;
	wire _w35744_ ;
	wire _w35743_ ;
	wire _w35742_ ;
	wire _w35741_ ;
	wire _w35740_ ;
	wire _w35739_ ;
	wire _w35738_ ;
	wire _w35737_ ;
	wire _w35736_ ;
	wire _w35735_ ;
	wire _w35734_ ;
	wire _w35733_ ;
	wire _w35732_ ;
	wire _w35731_ ;
	wire _w35730_ ;
	wire _w35729_ ;
	wire _w35728_ ;
	wire _w35727_ ;
	wire _w35726_ ;
	wire _w35725_ ;
	wire _w35724_ ;
	wire _w35723_ ;
	wire _w35722_ ;
	wire _w35721_ ;
	wire _w35720_ ;
	wire _w35719_ ;
	wire _w35718_ ;
	wire _w35717_ ;
	wire _w35716_ ;
	wire _w35715_ ;
	wire _w35714_ ;
	wire _w35713_ ;
	wire _w35712_ ;
	wire _w35711_ ;
	wire _w35710_ ;
	wire _w35709_ ;
	wire _w35708_ ;
	wire _w35707_ ;
	wire _w35706_ ;
	wire _w35705_ ;
	wire _w35704_ ;
	wire _w35703_ ;
	wire _w35702_ ;
	wire _w35701_ ;
	wire _w35700_ ;
	wire _w35699_ ;
	wire _w35698_ ;
	wire _w35697_ ;
	wire _w35696_ ;
	wire _w35695_ ;
	wire _w35694_ ;
	wire _w35693_ ;
	wire _w35692_ ;
	wire _w35691_ ;
	wire _w35690_ ;
	wire _w35689_ ;
	wire _w35688_ ;
	wire _w35687_ ;
	wire _w35686_ ;
	wire _w35685_ ;
	wire _w35684_ ;
	wire _w35683_ ;
	wire _w35682_ ;
	wire _w35681_ ;
	wire _w35680_ ;
	wire _w35679_ ;
	wire _w35678_ ;
	wire _w35677_ ;
	wire _w35676_ ;
	wire _w35675_ ;
	wire _w35674_ ;
	wire _w35673_ ;
	wire _w35672_ ;
	wire _w35671_ ;
	wire _w35670_ ;
	wire _w35669_ ;
	wire _w35668_ ;
	wire _w35667_ ;
	wire _w35666_ ;
	wire _w35665_ ;
	wire _w35664_ ;
	wire _w35663_ ;
	wire _w35662_ ;
	wire _w35661_ ;
	wire _w35660_ ;
	wire _w35659_ ;
	wire _w35658_ ;
	wire _w35657_ ;
	wire _w35656_ ;
	wire _w35655_ ;
	wire _w35654_ ;
	wire _w35653_ ;
	wire _w35652_ ;
	wire _w35651_ ;
	wire _w35650_ ;
	wire _w35649_ ;
	wire _w35648_ ;
	wire _w35647_ ;
	wire _w35646_ ;
	wire _w35645_ ;
	wire _w35644_ ;
	wire _w35643_ ;
	wire _w35642_ ;
	wire _w35641_ ;
	wire _w35640_ ;
	wire _w35639_ ;
	wire _w35638_ ;
	wire _w35637_ ;
	wire _w35636_ ;
	wire _w35635_ ;
	wire _w35634_ ;
	wire _w35633_ ;
	wire _w35632_ ;
	wire _w35631_ ;
	wire _w35630_ ;
	wire _w35629_ ;
	wire _w35628_ ;
	wire _w35627_ ;
	wire _w35626_ ;
	wire _w35625_ ;
	wire _w35624_ ;
	wire _w35623_ ;
	wire _w35622_ ;
	wire _w35621_ ;
	wire _w35620_ ;
	wire _w35619_ ;
	wire _w35618_ ;
	wire _w35617_ ;
	wire _w35616_ ;
	wire _w35615_ ;
	wire _w35614_ ;
	wire _w35613_ ;
	wire _w35612_ ;
	wire _w35611_ ;
	wire _w35610_ ;
	wire _w35609_ ;
	wire _w35608_ ;
	wire _w35607_ ;
	wire _w35606_ ;
	wire _w35605_ ;
	wire _w35604_ ;
	wire _w35603_ ;
	wire _w35602_ ;
	wire _w35601_ ;
	wire _w35600_ ;
	wire _w35599_ ;
	wire _w35598_ ;
	wire _w35597_ ;
	wire _w35596_ ;
	wire _w35595_ ;
	wire _w35594_ ;
	wire _w35593_ ;
	wire _w35592_ ;
	wire _w35591_ ;
	wire _w35590_ ;
	wire _w35589_ ;
	wire _w35588_ ;
	wire _w35587_ ;
	wire _w35586_ ;
	wire _w35585_ ;
	wire _w35584_ ;
	wire _w35583_ ;
	wire _w35582_ ;
	wire _w35581_ ;
	wire _w35580_ ;
	wire _w35579_ ;
	wire _w35578_ ;
	wire _w35577_ ;
	wire _w35576_ ;
	wire _w35575_ ;
	wire _w35574_ ;
	wire _w35573_ ;
	wire _w35572_ ;
	wire _w35571_ ;
	wire _w35570_ ;
	wire _w35569_ ;
	wire _w35568_ ;
	wire _w35567_ ;
	wire _w35566_ ;
	wire _w35565_ ;
	wire _w35564_ ;
	wire _w35563_ ;
	wire _w35562_ ;
	wire _w35561_ ;
	wire _w35560_ ;
	wire _w35559_ ;
	wire _w35558_ ;
	wire _w35557_ ;
	wire _w35556_ ;
	wire _w35555_ ;
	wire _w35554_ ;
	wire _w35553_ ;
	wire _w35552_ ;
	wire _w35551_ ;
	wire _w35550_ ;
	wire _w35549_ ;
	wire _w35548_ ;
	wire _w35547_ ;
	wire _w35546_ ;
	wire _w35545_ ;
	wire _w35544_ ;
	wire _w35543_ ;
	wire _w35542_ ;
	wire _w35541_ ;
	wire _w35540_ ;
	wire _w35539_ ;
	wire _w35538_ ;
	wire _w35537_ ;
	wire _w35536_ ;
	wire _w35535_ ;
	wire _w35534_ ;
	wire _w35533_ ;
	wire _w35532_ ;
	wire _w35531_ ;
	wire _w35530_ ;
	wire _w35529_ ;
	wire _w35528_ ;
	wire _w35527_ ;
	wire _w35526_ ;
	wire _w35525_ ;
	wire _w35524_ ;
	wire _w35523_ ;
	wire _w35522_ ;
	wire _w35521_ ;
	wire _w35520_ ;
	wire _w35519_ ;
	wire _w35518_ ;
	wire _w35517_ ;
	wire _w35516_ ;
	wire _w35515_ ;
	wire _w35514_ ;
	wire _w35513_ ;
	wire _w35512_ ;
	wire _w35511_ ;
	wire _w35510_ ;
	wire _w35509_ ;
	wire _w35508_ ;
	wire _w35507_ ;
	wire _w35506_ ;
	wire _w35505_ ;
	wire _w35504_ ;
	wire _w35503_ ;
	wire _w35502_ ;
	wire _w35501_ ;
	wire _w35500_ ;
	wire _w35499_ ;
	wire _w35498_ ;
	wire _w35497_ ;
	wire _w35496_ ;
	wire _w35495_ ;
	wire _w35494_ ;
	wire _w35493_ ;
	wire _w35492_ ;
	wire _w35491_ ;
	wire _w35490_ ;
	wire _w35489_ ;
	wire _w35488_ ;
	wire _w35487_ ;
	wire _w35486_ ;
	wire _w35485_ ;
	wire _w35484_ ;
	wire _w35483_ ;
	wire _w35482_ ;
	wire _w35481_ ;
	wire _w35480_ ;
	wire _w35479_ ;
	wire _w35478_ ;
	wire _w35477_ ;
	wire _w35476_ ;
	wire _w35475_ ;
	wire _w35474_ ;
	wire _w35473_ ;
	wire _w35472_ ;
	wire _w35471_ ;
	wire _w35470_ ;
	wire _w35469_ ;
	wire _w35468_ ;
	wire _w35467_ ;
	wire _w35466_ ;
	wire _w35465_ ;
	wire _w35464_ ;
	wire _w35463_ ;
	wire _w35462_ ;
	wire _w35461_ ;
	wire _w35460_ ;
	wire _w35459_ ;
	wire _w35458_ ;
	wire _w35457_ ;
	wire _w35456_ ;
	wire _w35455_ ;
	wire _w35454_ ;
	wire _w35453_ ;
	wire _w35452_ ;
	wire _w35451_ ;
	wire _w35450_ ;
	wire _w35449_ ;
	wire _w35448_ ;
	wire _w35447_ ;
	wire _w35446_ ;
	wire _w35445_ ;
	wire _w35444_ ;
	wire _w35443_ ;
	wire _w35442_ ;
	wire _w35441_ ;
	wire _w35440_ ;
	wire _w35439_ ;
	wire _w35438_ ;
	wire _w35437_ ;
	wire _w35436_ ;
	wire _w35435_ ;
	wire _w35434_ ;
	wire _w35433_ ;
	wire _w35432_ ;
	wire _w35431_ ;
	wire _w35430_ ;
	wire _w35429_ ;
	wire _w35428_ ;
	wire _w35427_ ;
	wire _w35426_ ;
	wire _w35425_ ;
	wire _w35424_ ;
	wire _w35423_ ;
	wire _w35422_ ;
	wire _w35421_ ;
	wire _w35420_ ;
	wire _w35419_ ;
	wire _w35418_ ;
	wire _w35417_ ;
	wire _w35416_ ;
	wire _w35415_ ;
	wire _w35414_ ;
	wire _w35413_ ;
	wire _w35412_ ;
	wire _w35411_ ;
	wire _w35410_ ;
	wire _w35409_ ;
	wire _w35408_ ;
	wire _w35407_ ;
	wire _w35406_ ;
	wire _w35405_ ;
	wire _w35404_ ;
	wire _w35403_ ;
	wire _w35402_ ;
	wire _w35401_ ;
	wire _w35400_ ;
	wire _w35399_ ;
	wire _w35398_ ;
	wire _w35397_ ;
	wire _w35396_ ;
	wire _w35395_ ;
	wire _w35394_ ;
	wire _w35393_ ;
	wire _w35392_ ;
	wire _w35391_ ;
	wire _w35390_ ;
	wire _w35389_ ;
	wire _w35388_ ;
	wire _w35387_ ;
	wire _w35386_ ;
	wire _w35385_ ;
	wire _w35384_ ;
	wire _w35383_ ;
	wire _w35382_ ;
	wire _w35381_ ;
	wire _w35380_ ;
	wire _w35379_ ;
	wire _w35378_ ;
	wire _w35377_ ;
	wire _w35376_ ;
	wire _w35375_ ;
	wire _w35374_ ;
	wire _w35373_ ;
	wire _w35372_ ;
	wire _w35371_ ;
	wire _w35370_ ;
	wire _w35369_ ;
	wire _w35368_ ;
	wire _w35367_ ;
	wire _w35366_ ;
	wire _w35365_ ;
	wire _w35364_ ;
	wire _w35363_ ;
	wire _w35362_ ;
	wire _w35361_ ;
	wire _w35360_ ;
	wire _w35359_ ;
	wire _w35358_ ;
	wire _w35357_ ;
	wire _w35356_ ;
	wire _w35355_ ;
	wire _w35354_ ;
	wire _w35353_ ;
	wire _w35352_ ;
	wire _w35351_ ;
	wire _w35350_ ;
	wire _w35349_ ;
	wire _w35348_ ;
	wire _w35347_ ;
	wire _w35346_ ;
	wire _w35345_ ;
	wire _w35344_ ;
	wire _w35343_ ;
	wire _w35342_ ;
	wire _w35341_ ;
	wire _w35340_ ;
	wire _w35339_ ;
	wire _w35338_ ;
	wire _w35337_ ;
	wire _w35336_ ;
	wire _w35335_ ;
	wire _w35334_ ;
	wire _w35333_ ;
	wire _w35332_ ;
	wire _w35331_ ;
	wire _w35330_ ;
	wire _w35329_ ;
	wire _w35328_ ;
	wire _w35327_ ;
	wire _w35326_ ;
	wire _w35325_ ;
	wire _w35324_ ;
	wire _w35323_ ;
	wire _w35322_ ;
	wire _w35321_ ;
	wire _w35320_ ;
	wire _w35319_ ;
	wire _w35318_ ;
	wire _w35317_ ;
	wire _w35316_ ;
	wire _w35315_ ;
	wire _w35314_ ;
	wire _w35313_ ;
	wire _w35312_ ;
	wire _w35311_ ;
	wire _w35310_ ;
	wire _w35309_ ;
	wire _w35308_ ;
	wire _w35307_ ;
	wire _w35306_ ;
	wire _w35305_ ;
	wire _w35304_ ;
	wire _w35303_ ;
	wire _w35302_ ;
	wire _w35301_ ;
	wire _w35300_ ;
	wire _w35299_ ;
	wire _w35298_ ;
	wire _w35297_ ;
	wire _w35296_ ;
	wire _w35295_ ;
	wire _w35294_ ;
	wire _w35293_ ;
	wire _w35292_ ;
	wire _w35291_ ;
	wire _w35290_ ;
	wire _w35289_ ;
	wire _w35288_ ;
	wire _w35287_ ;
	wire _w35286_ ;
	wire _w35285_ ;
	wire _w35284_ ;
	wire _w35283_ ;
	wire _w35282_ ;
	wire _w35281_ ;
	wire _w35280_ ;
	wire _w35279_ ;
	wire _w35278_ ;
	wire _w35277_ ;
	wire _w35276_ ;
	wire _w35275_ ;
	wire _w35274_ ;
	wire _w35273_ ;
	wire _w35272_ ;
	wire _w35271_ ;
	wire _w35270_ ;
	wire _w35269_ ;
	wire _w35268_ ;
	wire _w35267_ ;
	wire _w35266_ ;
	wire _w35265_ ;
	wire _w35264_ ;
	wire _w35263_ ;
	wire _w35262_ ;
	wire _w35261_ ;
	wire _w35260_ ;
	wire _w35259_ ;
	wire _w35258_ ;
	wire _w35257_ ;
	wire _w35256_ ;
	wire _w35255_ ;
	wire _w35254_ ;
	wire _w35253_ ;
	wire _w35252_ ;
	wire _w35251_ ;
	wire _w35250_ ;
	wire _w35249_ ;
	wire _w35248_ ;
	wire _w35247_ ;
	wire _w35246_ ;
	wire _w35245_ ;
	wire _w35244_ ;
	wire _w35243_ ;
	wire _w35242_ ;
	wire _w35241_ ;
	wire _w35240_ ;
	wire _w35239_ ;
	wire _w35238_ ;
	wire _w35237_ ;
	wire _w35236_ ;
	wire _w35235_ ;
	wire _w35234_ ;
	wire _w35233_ ;
	wire _w35232_ ;
	wire _w35231_ ;
	wire _w35230_ ;
	wire _w35229_ ;
	wire _w35228_ ;
	wire _w35227_ ;
	wire _w35226_ ;
	wire _w35225_ ;
	wire _w35224_ ;
	wire _w35223_ ;
	wire _w35222_ ;
	wire _w35221_ ;
	wire _w35220_ ;
	wire _w35219_ ;
	wire _w35218_ ;
	wire _w35217_ ;
	wire _w35216_ ;
	wire _w35215_ ;
	wire _w35214_ ;
	wire _w35213_ ;
	wire _w35212_ ;
	wire _w35211_ ;
	wire _w35210_ ;
	wire _w35209_ ;
	wire _w35208_ ;
	wire _w35207_ ;
	wire _w35206_ ;
	wire _w35205_ ;
	wire _w35204_ ;
	wire _w35203_ ;
	wire _w35202_ ;
	wire _w35201_ ;
	wire _w35200_ ;
	wire _w35199_ ;
	wire _w35198_ ;
	wire _w35197_ ;
	wire _w35196_ ;
	wire _w35195_ ;
	wire _w35194_ ;
	wire _w35193_ ;
	wire _w35192_ ;
	wire _w35191_ ;
	wire _w35190_ ;
	wire _w35189_ ;
	wire _w35188_ ;
	wire _w35187_ ;
	wire _w35186_ ;
	wire _w35185_ ;
	wire _w35184_ ;
	wire _w35183_ ;
	wire _w35182_ ;
	wire _w35181_ ;
	wire _w35180_ ;
	wire _w35179_ ;
	wire _w35178_ ;
	wire _w35177_ ;
	wire _w35176_ ;
	wire _w35175_ ;
	wire _w35174_ ;
	wire _w35173_ ;
	wire _w35172_ ;
	wire _w35171_ ;
	wire _w35170_ ;
	wire _w35169_ ;
	wire _w35168_ ;
	wire _w35167_ ;
	wire _w35166_ ;
	wire _w35165_ ;
	wire _w35164_ ;
	wire _w35163_ ;
	wire _w35162_ ;
	wire _w35161_ ;
	wire _w35160_ ;
	wire _w35159_ ;
	wire _w35158_ ;
	wire _w35157_ ;
	wire _w35156_ ;
	wire _w35155_ ;
	wire _w35154_ ;
	wire _w35153_ ;
	wire _w35152_ ;
	wire _w35151_ ;
	wire _w35150_ ;
	wire _w35149_ ;
	wire _w35148_ ;
	wire _w35147_ ;
	wire _w35146_ ;
	wire _w35145_ ;
	wire _w35144_ ;
	wire _w35143_ ;
	wire _w35142_ ;
	wire _w35141_ ;
	wire _w35140_ ;
	wire _w35139_ ;
	wire _w35138_ ;
	wire _w35137_ ;
	wire _w35136_ ;
	wire _w35135_ ;
	wire _w35134_ ;
	wire _w35133_ ;
	wire _w35132_ ;
	wire _w35131_ ;
	wire _w35130_ ;
	wire _w35129_ ;
	wire _w35128_ ;
	wire _w35127_ ;
	wire _w35126_ ;
	wire _w35125_ ;
	wire _w35124_ ;
	wire _w35123_ ;
	wire _w35122_ ;
	wire _w35121_ ;
	wire _w35120_ ;
	wire _w35119_ ;
	wire _w35118_ ;
	wire _w35117_ ;
	wire _w35116_ ;
	wire _w35115_ ;
	wire _w35114_ ;
	wire _w35113_ ;
	wire _w35112_ ;
	wire _w35111_ ;
	wire _w35110_ ;
	wire _w35109_ ;
	wire _w35108_ ;
	wire _w35107_ ;
	wire _w35106_ ;
	wire _w35105_ ;
	wire _w35104_ ;
	wire _w35103_ ;
	wire _w35102_ ;
	wire _w35101_ ;
	wire _w35100_ ;
	wire _w35099_ ;
	wire _w35098_ ;
	wire _w35097_ ;
	wire _w35096_ ;
	wire _w35095_ ;
	wire _w35094_ ;
	wire _w35093_ ;
	wire _w35092_ ;
	wire _w35091_ ;
	wire _w35090_ ;
	wire _w35089_ ;
	wire _w35088_ ;
	wire _w35087_ ;
	wire _w35086_ ;
	wire _w35085_ ;
	wire _w35084_ ;
	wire _w35083_ ;
	wire _w35082_ ;
	wire _w35081_ ;
	wire _w35080_ ;
	wire _w35079_ ;
	wire _w35078_ ;
	wire _w35077_ ;
	wire _w35076_ ;
	wire _w35075_ ;
	wire _w35074_ ;
	wire _w35073_ ;
	wire _w35072_ ;
	wire _w35071_ ;
	wire _w35070_ ;
	wire _w35069_ ;
	wire _w35068_ ;
	wire _w35067_ ;
	wire _w35066_ ;
	wire _w35065_ ;
	wire _w35064_ ;
	wire _w35063_ ;
	wire _w35062_ ;
	wire _w35061_ ;
	wire _w35060_ ;
	wire _w35059_ ;
	wire _w35058_ ;
	wire _w35057_ ;
	wire _w35056_ ;
	wire _w35055_ ;
	wire _w35054_ ;
	wire _w35053_ ;
	wire _w35052_ ;
	wire _w35051_ ;
	wire _w35050_ ;
	wire _w35049_ ;
	wire _w35048_ ;
	wire _w35047_ ;
	wire _w35046_ ;
	wire _w35045_ ;
	wire _w35044_ ;
	wire _w35043_ ;
	wire _w35042_ ;
	wire _w35041_ ;
	wire _w35040_ ;
	wire _w35039_ ;
	wire _w35038_ ;
	wire _w35037_ ;
	wire _w35036_ ;
	wire _w35035_ ;
	wire _w35034_ ;
	wire _w35033_ ;
	wire _w35032_ ;
	wire _w35031_ ;
	wire _w35030_ ;
	wire _w35029_ ;
	wire _w35028_ ;
	wire _w35027_ ;
	wire _w35026_ ;
	wire _w35025_ ;
	wire _w35024_ ;
	wire _w35023_ ;
	wire _w35022_ ;
	wire _w35021_ ;
	wire _w35020_ ;
	wire _w35019_ ;
	wire _w35018_ ;
	wire _w35017_ ;
	wire _w35016_ ;
	wire _w35015_ ;
	wire _w35014_ ;
	wire _w35013_ ;
	wire _w35012_ ;
	wire _w35011_ ;
	wire _w35010_ ;
	wire _w35009_ ;
	wire _w35008_ ;
	wire _w35007_ ;
	wire _w35006_ ;
	wire _w35005_ ;
	wire _w35004_ ;
	wire _w35003_ ;
	wire _w35002_ ;
	wire _w35001_ ;
	wire _w35000_ ;
	wire _w34999_ ;
	wire _w34998_ ;
	wire _w34997_ ;
	wire _w34996_ ;
	wire _w34995_ ;
	wire _w34994_ ;
	wire _w34993_ ;
	wire _w34992_ ;
	wire _w34991_ ;
	wire _w34990_ ;
	wire _w34989_ ;
	wire _w34988_ ;
	wire _w34987_ ;
	wire _w34986_ ;
	wire _w34985_ ;
	wire _w34984_ ;
	wire _w34983_ ;
	wire _w34982_ ;
	wire _w34981_ ;
	wire _w34980_ ;
	wire _w34979_ ;
	wire _w34978_ ;
	wire _w34977_ ;
	wire _w34976_ ;
	wire _w34975_ ;
	wire _w34974_ ;
	wire _w34973_ ;
	wire _w34972_ ;
	wire _w34971_ ;
	wire _w34970_ ;
	wire _w34969_ ;
	wire _w34968_ ;
	wire _w34967_ ;
	wire _w34966_ ;
	wire _w34965_ ;
	wire _w34964_ ;
	wire _w34963_ ;
	wire _w34962_ ;
	wire _w34961_ ;
	wire _w34960_ ;
	wire _w34959_ ;
	wire _w34958_ ;
	wire _w34957_ ;
	wire _w34956_ ;
	wire _w34955_ ;
	wire _w34954_ ;
	wire _w34953_ ;
	wire _w34952_ ;
	wire _w34951_ ;
	wire _w34950_ ;
	wire _w34949_ ;
	wire _w34948_ ;
	wire _w34947_ ;
	wire _w34946_ ;
	wire _w34945_ ;
	wire _w34944_ ;
	wire _w34943_ ;
	wire _w34942_ ;
	wire _w34941_ ;
	wire _w34940_ ;
	wire _w34939_ ;
	wire _w34938_ ;
	wire _w34937_ ;
	wire _w34936_ ;
	wire _w34935_ ;
	wire _w34934_ ;
	wire _w34933_ ;
	wire _w34932_ ;
	wire _w34931_ ;
	wire _w34930_ ;
	wire _w34929_ ;
	wire _w34928_ ;
	wire _w34927_ ;
	wire _w34926_ ;
	wire _w34925_ ;
	wire _w34924_ ;
	wire _w34923_ ;
	wire _w34922_ ;
	wire _w34921_ ;
	wire _w34920_ ;
	wire _w34919_ ;
	wire _w34918_ ;
	wire _w34917_ ;
	wire _w34916_ ;
	wire _w34915_ ;
	wire _w34914_ ;
	wire _w34913_ ;
	wire _w34912_ ;
	wire _w34911_ ;
	wire _w34910_ ;
	wire _w34909_ ;
	wire _w34908_ ;
	wire _w34907_ ;
	wire _w34906_ ;
	wire _w34905_ ;
	wire _w34904_ ;
	wire _w34903_ ;
	wire _w34902_ ;
	wire _w34901_ ;
	wire _w34900_ ;
	wire _w34899_ ;
	wire _w34898_ ;
	wire _w34897_ ;
	wire _w34896_ ;
	wire _w34895_ ;
	wire _w34894_ ;
	wire _w34893_ ;
	wire _w34892_ ;
	wire _w34891_ ;
	wire _w34890_ ;
	wire _w34889_ ;
	wire _w34888_ ;
	wire _w34887_ ;
	wire _w34886_ ;
	wire _w34885_ ;
	wire _w34884_ ;
	wire _w34883_ ;
	wire _w34882_ ;
	wire _w34881_ ;
	wire _w34880_ ;
	wire _w34879_ ;
	wire _w34878_ ;
	wire _w34877_ ;
	wire _w34876_ ;
	wire _w34875_ ;
	wire _w34874_ ;
	wire _w34873_ ;
	wire _w34872_ ;
	wire _w34871_ ;
	wire _w34870_ ;
	wire _w34869_ ;
	wire _w34868_ ;
	wire _w34867_ ;
	wire _w34866_ ;
	wire _w34865_ ;
	wire _w34864_ ;
	wire _w34863_ ;
	wire _w34862_ ;
	wire _w34861_ ;
	wire _w34860_ ;
	wire _w34859_ ;
	wire _w34858_ ;
	wire _w34857_ ;
	wire _w34856_ ;
	wire _w34855_ ;
	wire _w34854_ ;
	wire _w34853_ ;
	wire _w34852_ ;
	wire _w34851_ ;
	wire _w34850_ ;
	wire _w34849_ ;
	wire _w34848_ ;
	wire _w34847_ ;
	wire _w34846_ ;
	wire _w34845_ ;
	wire _w34844_ ;
	wire _w34843_ ;
	wire _w34842_ ;
	wire _w34841_ ;
	wire _w34840_ ;
	wire _w34839_ ;
	wire _w34838_ ;
	wire _w34837_ ;
	wire _w34836_ ;
	wire _w34835_ ;
	wire _w34834_ ;
	wire _w34833_ ;
	wire _w34832_ ;
	wire _w34831_ ;
	wire _w34830_ ;
	wire _w34829_ ;
	wire _w34828_ ;
	wire _w34827_ ;
	wire _w34826_ ;
	wire _w34825_ ;
	wire _w34824_ ;
	wire _w34823_ ;
	wire _w34822_ ;
	wire _w34821_ ;
	wire _w34820_ ;
	wire _w34819_ ;
	wire _w34818_ ;
	wire _w34817_ ;
	wire _w34816_ ;
	wire _w34815_ ;
	wire _w34814_ ;
	wire _w34813_ ;
	wire _w34812_ ;
	wire _w34811_ ;
	wire _w34810_ ;
	wire _w34809_ ;
	wire _w34808_ ;
	wire _w34807_ ;
	wire _w34806_ ;
	wire _w34805_ ;
	wire _w34804_ ;
	wire _w34803_ ;
	wire _w34802_ ;
	wire _w34801_ ;
	wire _w34800_ ;
	wire _w34799_ ;
	wire _w34798_ ;
	wire _w34797_ ;
	wire _w34796_ ;
	wire _w34795_ ;
	wire _w34794_ ;
	wire _w34793_ ;
	wire _w34792_ ;
	wire _w34791_ ;
	wire _w34790_ ;
	wire _w34789_ ;
	wire _w34788_ ;
	wire _w34787_ ;
	wire _w34786_ ;
	wire _w34785_ ;
	wire _w34784_ ;
	wire _w34783_ ;
	wire _w34782_ ;
	wire _w34781_ ;
	wire _w34780_ ;
	wire _w34779_ ;
	wire _w34778_ ;
	wire _w34777_ ;
	wire _w34776_ ;
	wire _w34775_ ;
	wire _w34774_ ;
	wire _w34773_ ;
	wire _w34772_ ;
	wire _w34771_ ;
	wire _w34770_ ;
	wire _w34769_ ;
	wire _w34768_ ;
	wire _w34767_ ;
	wire _w34766_ ;
	wire _w34765_ ;
	wire _w34764_ ;
	wire _w34763_ ;
	wire _w34762_ ;
	wire _w34761_ ;
	wire _w34760_ ;
	wire _w34759_ ;
	wire _w34758_ ;
	wire _w34757_ ;
	wire _w34756_ ;
	wire _w34755_ ;
	wire _w34754_ ;
	wire _w34753_ ;
	wire _w34752_ ;
	wire _w34751_ ;
	wire _w34750_ ;
	wire _w34749_ ;
	wire _w34748_ ;
	wire _w34747_ ;
	wire _w34746_ ;
	wire _w34745_ ;
	wire _w34744_ ;
	wire _w34743_ ;
	wire _w34742_ ;
	wire _w34741_ ;
	wire _w34740_ ;
	wire _w34739_ ;
	wire _w34738_ ;
	wire _w34737_ ;
	wire _w34736_ ;
	wire _w34735_ ;
	wire _w34734_ ;
	wire _w34733_ ;
	wire _w34732_ ;
	wire _w34731_ ;
	wire _w34730_ ;
	wire _w34729_ ;
	wire _w34728_ ;
	wire _w34727_ ;
	wire _w34726_ ;
	wire _w34725_ ;
	wire _w34724_ ;
	wire _w34723_ ;
	wire _w34722_ ;
	wire _w34721_ ;
	wire _w34720_ ;
	wire _w34719_ ;
	wire _w34718_ ;
	wire _w34717_ ;
	wire _w34716_ ;
	wire _w34715_ ;
	wire _w34714_ ;
	wire _w34713_ ;
	wire _w34712_ ;
	wire _w34711_ ;
	wire _w34710_ ;
	wire _w34709_ ;
	wire _w34708_ ;
	wire _w34707_ ;
	wire _w34706_ ;
	wire _w34705_ ;
	wire _w34704_ ;
	wire _w34703_ ;
	wire _w34702_ ;
	wire _w34701_ ;
	wire _w34700_ ;
	wire _w34699_ ;
	wire _w34698_ ;
	wire _w34697_ ;
	wire _w34696_ ;
	wire _w34695_ ;
	wire _w34694_ ;
	wire _w34693_ ;
	wire _w34692_ ;
	wire _w34691_ ;
	wire _w34690_ ;
	wire _w34689_ ;
	wire _w34688_ ;
	wire _w34687_ ;
	wire _w34686_ ;
	wire _w34685_ ;
	wire _w34684_ ;
	wire _w34683_ ;
	wire _w34682_ ;
	wire _w34681_ ;
	wire _w34680_ ;
	wire _w34679_ ;
	wire _w34678_ ;
	wire _w34677_ ;
	wire _w34676_ ;
	wire _w34675_ ;
	wire _w34674_ ;
	wire _w34673_ ;
	wire _w34672_ ;
	wire _w34671_ ;
	wire _w34670_ ;
	wire _w34669_ ;
	wire _w34668_ ;
	wire _w34667_ ;
	wire _w34666_ ;
	wire _w34665_ ;
	wire _w34664_ ;
	wire _w34663_ ;
	wire _w34662_ ;
	wire _w34661_ ;
	wire _w34660_ ;
	wire _w34659_ ;
	wire _w34658_ ;
	wire _w34657_ ;
	wire _w34656_ ;
	wire _w34655_ ;
	wire _w34654_ ;
	wire _w34653_ ;
	wire _w34652_ ;
	wire _w34651_ ;
	wire _w34650_ ;
	wire _w34649_ ;
	wire _w34648_ ;
	wire _w34647_ ;
	wire _w34646_ ;
	wire _w34645_ ;
	wire _w34644_ ;
	wire _w34643_ ;
	wire _w34642_ ;
	wire _w34641_ ;
	wire _w34640_ ;
	wire _w34639_ ;
	wire _w34638_ ;
	wire _w34637_ ;
	wire _w34636_ ;
	wire _w34635_ ;
	wire _w34634_ ;
	wire _w34633_ ;
	wire _w34632_ ;
	wire _w34631_ ;
	wire _w34630_ ;
	wire _w34629_ ;
	wire _w34628_ ;
	wire _w34627_ ;
	wire _w34626_ ;
	wire _w34625_ ;
	wire _w34624_ ;
	wire _w34623_ ;
	wire _w34622_ ;
	wire _w34621_ ;
	wire _w34620_ ;
	wire _w34619_ ;
	wire _w34618_ ;
	wire _w34617_ ;
	wire _w34616_ ;
	wire _w34615_ ;
	wire _w34614_ ;
	wire _w34613_ ;
	wire _w34612_ ;
	wire _w34611_ ;
	wire _w34610_ ;
	wire _w34609_ ;
	wire _w34608_ ;
	wire _w34607_ ;
	wire _w34606_ ;
	wire _w34605_ ;
	wire _w34604_ ;
	wire _w34603_ ;
	wire _w34602_ ;
	wire _w34601_ ;
	wire _w34600_ ;
	wire _w34599_ ;
	wire _w34598_ ;
	wire _w34597_ ;
	wire _w34596_ ;
	wire _w34595_ ;
	wire _w34594_ ;
	wire _w34593_ ;
	wire _w34592_ ;
	wire _w34591_ ;
	wire _w34590_ ;
	wire _w34589_ ;
	wire _w34588_ ;
	wire _w34587_ ;
	wire _w34586_ ;
	wire _w34585_ ;
	wire _w34584_ ;
	wire _w34583_ ;
	wire _w34582_ ;
	wire _w34581_ ;
	wire _w34580_ ;
	wire _w34579_ ;
	wire _w34578_ ;
	wire _w34577_ ;
	wire _w34576_ ;
	wire _w34575_ ;
	wire _w34574_ ;
	wire _w34573_ ;
	wire _w34572_ ;
	wire _w34571_ ;
	wire _w34570_ ;
	wire _w34569_ ;
	wire _w34568_ ;
	wire _w34567_ ;
	wire _w34566_ ;
	wire _w34565_ ;
	wire _w34564_ ;
	wire _w34563_ ;
	wire _w34562_ ;
	wire _w34561_ ;
	wire _w34560_ ;
	wire _w34559_ ;
	wire _w34558_ ;
	wire _w34557_ ;
	wire _w34556_ ;
	wire _w34555_ ;
	wire _w34554_ ;
	wire _w34553_ ;
	wire _w34552_ ;
	wire _w34551_ ;
	wire _w34550_ ;
	wire _w34549_ ;
	wire _w34548_ ;
	wire _w34547_ ;
	wire _w34546_ ;
	wire _w34545_ ;
	wire _w34544_ ;
	wire _w34543_ ;
	wire _w34542_ ;
	wire _w34541_ ;
	wire _w34540_ ;
	wire _w34539_ ;
	wire _w34538_ ;
	wire _w34537_ ;
	wire _w34536_ ;
	wire _w34535_ ;
	wire _w34534_ ;
	wire _w34533_ ;
	wire _w34532_ ;
	wire _w34531_ ;
	wire _w34530_ ;
	wire _w34529_ ;
	wire _w34528_ ;
	wire _w34527_ ;
	wire _w34526_ ;
	wire _w34525_ ;
	wire _w34524_ ;
	wire _w34523_ ;
	wire _w34522_ ;
	wire _w34521_ ;
	wire _w34520_ ;
	wire _w34519_ ;
	wire _w34518_ ;
	wire _w34517_ ;
	wire _w34516_ ;
	wire _w34515_ ;
	wire _w34514_ ;
	wire _w34513_ ;
	wire _w34512_ ;
	wire _w34511_ ;
	wire _w34510_ ;
	wire _w34509_ ;
	wire _w34508_ ;
	wire _w34507_ ;
	wire _w34506_ ;
	wire _w34505_ ;
	wire _w34504_ ;
	wire _w34503_ ;
	wire _w34502_ ;
	wire _w34501_ ;
	wire _w34500_ ;
	wire _w34499_ ;
	wire _w34498_ ;
	wire _w34497_ ;
	wire _w34496_ ;
	wire _w34495_ ;
	wire _w34494_ ;
	wire _w34493_ ;
	wire _w34492_ ;
	wire _w34491_ ;
	wire _w34490_ ;
	wire _w34489_ ;
	wire _w34488_ ;
	wire _w34487_ ;
	wire _w34486_ ;
	wire _w34485_ ;
	wire _w34484_ ;
	wire _w34483_ ;
	wire _w34482_ ;
	wire _w34481_ ;
	wire _w34480_ ;
	wire _w34479_ ;
	wire _w34478_ ;
	wire _w34477_ ;
	wire _w34476_ ;
	wire _w34475_ ;
	wire _w34474_ ;
	wire _w34473_ ;
	wire _w34472_ ;
	wire _w34471_ ;
	wire _w34470_ ;
	wire _w34469_ ;
	wire _w34468_ ;
	wire _w34467_ ;
	wire _w34466_ ;
	wire _w34465_ ;
	wire _w34464_ ;
	wire _w34463_ ;
	wire _w34462_ ;
	wire _w34461_ ;
	wire _w34460_ ;
	wire _w34459_ ;
	wire _w34458_ ;
	wire _w34457_ ;
	wire _w34456_ ;
	wire _w34455_ ;
	wire _w34454_ ;
	wire _w34453_ ;
	wire _w34452_ ;
	wire _w34451_ ;
	wire _w34450_ ;
	wire _w34449_ ;
	wire _w34448_ ;
	wire _w34447_ ;
	wire _w34446_ ;
	wire _w34445_ ;
	wire _w34444_ ;
	wire _w34443_ ;
	wire _w34442_ ;
	wire _w34441_ ;
	wire _w34440_ ;
	wire _w34439_ ;
	wire _w34438_ ;
	wire _w34437_ ;
	wire _w34436_ ;
	wire _w34435_ ;
	wire _w34434_ ;
	wire _w34433_ ;
	wire _w34432_ ;
	wire _w34431_ ;
	wire _w34430_ ;
	wire _w34429_ ;
	wire _w34428_ ;
	wire _w34427_ ;
	wire _w34426_ ;
	wire _w34425_ ;
	wire _w34424_ ;
	wire _w34423_ ;
	wire _w34422_ ;
	wire _w34421_ ;
	wire _w34420_ ;
	wire _w34419_ ;
	wire _w34418_ ;
	wire _w34417_ ;
	wire _w34416_ ;
	wire _w34415_ ;
	wire _w34414_ ;
	wire _w34413_ ;
	wire _w34412_ ;
	wire _w34411_ ;
	wire _w34410_ ;
	wire _w34409_ ;
	wire _w34408_ ;
	wire _w34407_ ;
	wire _w34406_ ;
	wire _w34405_ ;
	wire _w34404_ ;
	wire _w34403_ ;
	wire _w34402_ ;
	wire _w34401_ ;
	wire _w34400_ ;
	wire _w34399_ ;
	wire _w34398_ ;
	wire _w34397_ ;
	wire _w34396_ ;
	wire _w34395_ ;
	wire _w34394_ ;
	wire _w34393_ ;
	wire _w34392_ ;
	wire _w34391_ ;
	wire _w34390_ ;
	wire _w34389_ ;
	wire _w34388_ ;
	wire _w34387_ ;
	wire _w34386_ ;
	wire _w34385_ ;
	wire _w34384_ ;
	wire _w34383_ ;
	wire _w34382_ ;
	wire _w34381_ ;
	wire _w34380_ ;
	wire _w34379_ ;
	wire _w34378_ ;
	wire _w34377_ ;
	wire _w34376_ ;
	wire _w34375_ ;
	wire _w34374_ ;
	wire _w34373_ ;
	wire _w34372_ ;
	wire _w34371_ ;
	wire _w34370_ ;
	wire _w34369_ ;
	wire _w34368_ ;
	wire _w34367_ ;
	wire _w34366_ ;
	wire _w34365_ ;
	wire _w34364_ ;
	wire _w34363_ ;
	wire _w34362_ ;
	wire _w34361_ ;
	wire _w34360_ ;
	wire _w34359_ ;
	wire _w34358_ ;
	wire _w34357_ ;
	wire _w34356_ ;
	wire _w34355_ ;
	wire _w34354_ ;
	wire _w34353_ ;
	wire _w34352_ ;
	wire _w34351_ ;
	wire _w34350_ ;
	wire _w34349_ ;
	wire _w34348_ ;
	wire _w34347_ ;
	wire _w34346_ ;
	wire _w34345_ ;
	wire _w34344_ ;
	wire _w34343_ ;
	wire _w34342_ ;
	wire _w34341_ ;
	wire _w34340_ ;
	wire _w34339_ ;
	wire _w34338_ ;
	wire _w34337_ ;
	wire _w34336_ ;
	wire _w34335_ ;
	wire _w34334_ ;
	wire _w34333_ ;
	wire _w34332_ ;
	wire _w34331_ ;
	wire _w34330_ ;
	wire _w34329_ ;
	wire _w34328_ ;
	wire _w34327_ ;
	wire _w34326_ ;
	wire _w34325_ ;
	wire _w34324_ ;
	wire _w34323_ ;
	wire _w34322_ ;
	wire _w34321_ ;
	wire _w34320_ ;
	wire _w34319_ ;
	wire _w34318_ ;
	wire _w34317_ ;
	wire _w34316_ ;
	wire _w34315_ ;
	wire _w34314_ ;
	wire _w34313_ ;
	wire _w34312_ ;
	wire _w34311_ ;
	wire _w34310_ ;
	wire _w34309_ ;
	wire _w34308_ ;
	wire _w34307_ ;
	wire _w34306_ ;
	wire _w34305_ ;
	wire _w34304_ ;
	wire _w34303_ ;
	wire _w34302_ ;
	wire _w34301_ ;
	wire _w34300_ ;
	wire _w34299_ ;
	wire _w34298_ ;
	wire _w34297_ ;
	wire _w34296_ ;
	wire _w34295_ ;
	wire _w34294_ ;
	wire _w34293_ ;
	wire _w34292_ ;
	wire _w34291_ ;
	wire _w34290_ ;
	wire _w34289_ ;
	wire _w34288_ ;
	wire _w34287_ ;
	wire _w34286_ ;
	wire _w34285_ ;
	wire _w34284_ ;
	wire _w34283_ ;
	wire _w34282_ ;
	wire _w34281_ ;
	wire _w34280_ ;
	wire _w34279_ ;
	wire _w34278_ ;
	wire _w34277_ ;
	wire _w34276_ ;
	wire _w34275_ ;
	wire _w34274_ ;
	wire _w34273_ ;
	wire _w34272_ ;
	wire _w34271_ ;
	wire _w34270_ ;
	wire _w34269_ ;
	wire _w34268_ ;
	wire _w34267_ ;
	wire _w34266_ ;
	wire _w34265_ ;
	wire _w34264_ ;
	wire _w34263_ ;
	wire _w34262_ ;
	wire _w34261_ ;
	wire _w34260_ ;
	wire _w34259_ ;
	wire _w34258_ ;
	wire _w34257_ ;
	wire _w34256_ ;
	wire _w34255_ ;
	wire _w34254_ ;
	wire _w34253_ ;
	wire _w34252_ ;
	wire _w34251_ ;
	wire _w34250_ ;
	wire _w34249_ ;
	wire _w34248_ ;
	wire _w34247_ ;
	wire _w34246_ ;
	wire _w34245_ ;
	wire _w34244_ ;
	wire _w34243_ ;
	wire _w34242_ ;
	wire _w34241_ ;
	wire _w34240_ ;
	wire _w34239_ ;
	wire _w34238_ ;
	wire _w34237_ ;
	wire _w34236_ ;
	wire _w34235_ ;
	wire _w34234_ ;
	wire _w34233_ ;
	wire _w34232_ ;
	wire _w34231_ ;
	wire _w34230_ ;
	wire _w34229_ ;
	wire _w34228_ ;
	wire _w34227_ ;
	wire _w34226_ ;
	wire _w34225_ ;
	wire _w34224_ ;
	wire _w34223_ ;
	wire _w34222_ ;
	wire _w34221_ ;
	wire _w34220_ ;
	wire _w34219_ ;
	wire _w34218_ ;
	wire _w34217_ ;
	wire _w34216_ ;
	wire _w34215_ ;
	wire _w34214_ ;
	wire _w34213_ ;
	wire _w34212_ ;
	wire _w34211_ ;
	wire _w34210_ ;
	wire _w34209_ ;
	wire _w34208_ ;
	wire _w34207_ ;
	wire _w34206_ ;
	wire _w34205_ ;
	wire _w34204_ ;
	wire _w34203_ ;
	wire _w34202_ ;
	wire _w34201_ ;
	wire _w34200_ ;
	wire _w34199_ ;
	wire _w34198_ ;
	wire _w34197_ ;
	wire _w34196_ ;
	wire _w34195_ ;
	wire _w34194_ ;
	wire _w34193_ ;
	wire _w34192_ ;
	wire _w34191_ ;
	wire _w34190_ ;
	wire _w34189_ ;
	wire _w34188_ ;
	wire _w34187_ ;
	wire _w34186_ ;
	wire _w34185_ ;
	wire _w34184_ ;
	wire _w34183_ ;
	wire _w34182_ ;
	wire _w34181_ ;
	wire _w34180_ ;
	wire _w34179_ ;
	wire _w34178_ ;
	wire _w34177_ ;
	wire _w34176_ ;
	wire _w34175_ ;
	wire _w34174_ ;
	wire _w34173_ ;
	wire _w34172_ ;
	wire _w34171_ ;
	wire _w34170_ ;
	wire _w34169_ ;
	wire _w34168_ ;
	wire _w34167_ ;
	wire _w34166_ ;
	wire _w34165_ ;
	wire _w34164_ ;
	wire _w34163_ ;
	wire _w34162_ ;
	wire _w34161_ ;
	wire _w34160_ ;
	wire _w34159_ ;
	wire _w34158_ ;
	wire _w34157_ ;
	wire _w34156_ ;
	wire _w34155_ ;
	wire _w34154_ ;
	wire _w34153_ ;
	wire _w34152_ ;
	wire _w34151_ ;
	wire _w34150_ ;
	wire _w34149_ ;
	wire _w34148_ ;
	wire _w34147_ ;
	wire _w34146_ ;
	wire _w34145_ ;
	wire _w34144_ ;
	wire _w34143_ ;
	wire _w34142_ ;
	wire _w34141_ ;
	wire _w34140_ ;
	wire _w34139_ ;
	wire _w34138_ ;
	wire _w34137_ ;
	wire _w34136_ ;
	wire _w34135_ ;
	wire _w34134_ ;
	wire _w34133_ ;
	wire _w34132_ ;
	wire _w34131_ ;
	wire _w34130_ ;
	wire _w34129_ ;
	wire _w34128_ ;
	wire _w34127_ ;
	wire _w34126_ ;
	wire _w34125_ ;
	wire _w34124_ ;
	wire _w34123_ ;
	wire _w34122_ ;
	wire _w34121_ ;
	wire _w34120_ ;
	wire _w34119_ ;
	wire _w34118_ ;
	wire _w34117_ ;
	wire _w34116_ ;
	wire _w34115_ ;
	wire _w34114_ ;
	wire _w34113_ ;
	wire _w34112_ ;
	wire _w34111_ ;
	wire _w34110_ ;
	wire _w34109_ ;
	wire _w34108_ ;
	wire _w34107_ ;
	wire _w34106_ ;
	wire _w34105_ ;
	wire _w34104_ ;
	wire _w34103_ ;
	wire _w34102_ ;
	wire _w34101_ ;
	wire _w34100_ ;
	wire _w34099_ ;
	wire _w34098_ ;
	wire _w34097_ ;
	wire _w34096_ ;
	wire _w34095_ ;
	wire _w34094_ ;
	wire _w34093_ ;
	wire _w34092_ ;
	wire _w34091_ ;
	wire _w34090_ ;
	wire _w34089_ ;
	wire _w34088_ ;
	wire _w34087_ ;
	wire _w34086_ ;
	wire _w34085_ ;
	wire _w34084_ ;
	wire _w34083_ ;
	wire _w34082_ ;
	wire _w34081_ ;
	wire _w34080_ ;
	wire _w34079_ ;
	wire _w34078_ ;
	wire _w34077_ ;
	wire _w34076_ ;
	wire _w34075_ ;
	wire _w34074_ ;
	wire _w34073_ ;
	wire _w34072_ ;
	wire _w34071_ ;
	wire _w34070_ ;
	wire _w34069_ ;
	wire _w34068_ ;
	wire _w34067_ ;
	wire _w34066_ ;
	wire _w34065_ ;
	wire _w34064_ ;
	wire _w34063_ ;
	wire _w34062_ ;
	wire _w34061_ ;
	wire _w34060_ ;
	wire _w34059_ ;
	wire _w34058_ ;
	wire _w34057_ ;
	wire _w34056_ ;
	wire _w34055_ ;
	wire _w34054_ ;
	wire _w34053_ ;
	wire _w34052_ ;
	wire _w34051_ ;
	wire _w34050_ ;
	wire _w34049_ ;
	wire _w34048_ ;
	wire _w34047_ ;
	wire _w34046_ ;
	wire _w34045_ ;
	wire _w34044_ ;
	wire _w34043_ ;
	wire _w34042_ ;
	wire _w34041_ ;
	wire _w34040_ ;
	wire _w34039_ ;
	wire _w34038_ ;
	wire _w34037_ ;
	wire _w34036_ ;
	wire _w34035_ ;
	wire _w34034_ ;
	wire _w34033_ ;
	wire _w34032_ ;
	wire _w34031_ ;
	wire _w34030_ ;
	wire _w34029_ ;
	wire _w34028_ ;
	wire _w34027_ ;
	wire _w34026_ ;
	wire _w34025_ ;
	wire _w34024_ ;
	wire _w34023_ ;
	wire _w34022_ ;
	wire _w34021_ ;
	wire _w34020_ ;
	wire _w34019_ ;
	wire _w34018_ ;
	wire _w34017_ ;
	wire _w34016_ ;
	wire _w34015_ ;
	wire _w34014_ ;
	wire _w34013_ ;
	wire _w34012_ ;
	wire _w34011_ ;
	wire _w34010_ ;
	wire _w34009_ ;
	wire _w34008_ ;
	wire _w34007_ ;
	wire _w34006_ ;
	wire _w34005_ ;
	wire _w34004_ ;
	wire _w34003_ ;
	wire _w34002_ ;
	wire _w34001_ ;
	wire _w34000_ ;
	wire _w33999_ ;
	wire _w33998_ ;
	wire _w33997_ ;
	wire _w33996_ ;
	wire _w33995_ ;
	wire _w33994_ ;
	wire _w33993_ ;
	wire _w33992_ ;
	wire _w33991_ ;
	wire _w33990_ ;
	wire _w33989_ ;
	wire _w33988_ ;
	wire _w33987_ ;
	wire _w33986_ ;
	wire _w33985_ ;
	wire _w33984_ ;
	wire _w33983_ ;
	wire _w33982_ ;
	wire _w33981_ ;
	wire _w33980_ ;
	wire _w33979_ ;
	wire _w33978_ ;
	wire _w33977_ ;
	wire _w33976_ ;
	wire _w33975_ ;
	wire _w33974_ ;
	wire _w33973_ ;
	wire _w33972_ ;
	wire _w33971_ ;
	wire _w33970_ ;
	wire _w33969_ ;
	wire _w33968_ ;
	wire _w33967_ ;
	wire _w33966_ ;
	wire _w33965_ ;
	wire _w33964_ ;
	wire _w33963_ ;
	wire _w33962_ ;
	wire _w33961_ ;
	wire _w33960_ ;
	wire _w33959_ ;
	wire _w33958_ ;
	wire _w33957_ ;
	wire _w33956_ ;
	wire _w33955_ ;
	wire _w33954_ ;
	wire _w33953_ ;
	wire _w33952_ ;
	wire _w33951_ ;
	wire _w33950_ ;
	wire _w33949_ ;
	wire _w33948_ ;
	wire _w33947_ ;
	wire _w33946_ ;
	wire _w33945_ ;
	wire _w33944_ ;
	wire _w33943_ ;
	wire _w33942_ ;
	wire _w33941_ ;
	wire _w33940_ ;
	wire _w33939_ ;
	wire _w33938_ ;
	wire _w33937_ ;
	wire _w33936_ ;
	wire _w33935_ ;
	wire _w33934_ ;
	wire _w33933_ ;
	wire _w33932_ ;
	wire _w33931_ ;
	wire _w33930_ ;
	wire _w33929_ ;
	wire _w33928_ ;
	wire _w33927_ ;
	wire _w33926_ ;
	wire _w33925_ ;
	wire _w33924_ ;
	wire _w33923_ ;
	wire _w33922_ ;
	wire _w33921_ ;
	wire _w33920_ ;
	wire _w33919_ ;
	wire _w33918_ ;
	wire _w33917_ ;
	wire _w33916_ ;
	wire _w33915_ ;
	wire _w33914_ ;
	wire _w33913_ ;
	wire _w33912_ ;
	wire _w33911_ ;
	wire _w33910_ ;
	wire _w33909_ ;
	wire _w33908_ ;
	wire _w33907_ ;
	wire _w33906_ ;
	wire _w33905_ ;
	wire _w33904_ ;
	wire _w33903_ ;
	wire _w33902_ ;
	wire _w33901_ ;
	wire _w33900_ ;
	wire _w33899_ ;
	wire _w33898_ ;
	wire _w33897_ ;
	wire _w33896_ ;
	wire _w33895_ ;
	wire _w33894_ ;
	wire _w33893_ ;
	wire _w33892_ ;
	wire _w33891_ ;
	wire _w33890_ ;
	wire _w33889_ ;
	wire _w33888_ ;
	wire _w33887_ ;
	wire _w33886_ ;
	wire _w33885_ ;
	wire _w33884_ ;
	wire _w33883_ ;
	wire _w33882_ ;
	wire _w33881_ ;
	wire _w33880_ ;
	wire _w33879_ ;
	wire _w33878_ ;
	wire _w33877_ ;
	wire _w33876_ ;
	wire _w33875_ ;
	wire _w33874_ ;
	wire _w33873_ ;
	wire _w33872_ ;
	wire _w33871_ ;
	wire _w33870_ ;
	wire _w33869_ ;
	wire _w33868_ ;
	wire _w33867_ ;
	wire _w33866_ ;
	wire _w33865_ ;
	wire _w33864_ ;
	wire _w33863_ ;
	wire _w33862_ ;
	wire _w33861_ ;
	wire _w33860_ ;
	wire _w33859_ ;
	wire _w33858_ ;
	wire _w33857_ ;
	wire _w33856_ ;
	wire _w33855_ ;
	wire _w33854_ ;
	wire _w33853_ ;
	wire _w33852_ ;
	wire _w33851_ ;
	wire _w33850_ ;
	wire _w33849_ ;
	wire _w33848_ ;
	wire _w33847_ ;
	wire _w33846_ ;
	wire _w33845_ ;
	wire _w33844_ ;
	wire _w33843_ ;
	wire _w33842_ ;
	wire _w33841_ ;
	wire _w33840_ ;
	wire _w33839_ ;
	wire _w33838_ ;
	wire _w33837_ ;
	wire _w33836_ ;
	wire _w33835_ ;
	wire _w33834_ ;
	wire _w33833_ ;
	wire _w33832_ ;
	wire _w33831_ ;
	wire _w33830_ ;
	wire _w33829_ ;
	wire _w33828_ ;
	wire _w33827_ ;
	wire _w33826_ ;
	wire _w33825_ ;
	wire _w33824_ ;
	wire _w33823_ ;
	wire _w33822_ ;
	wire _w33821_ ;
	wire _w33820_ ;
	wire _w33819_ ;
	wire _w33818_ ;
	wire _w33817_ ;
	wire _w33816_ ;
	wire _w33815_ ;
	wire _w33814_ ;
	wire _w33813_ ;
	wire _w33812_ ;
	wire _w33811_ ;
	wire _w33810_ ;
	wire _w33809_ ;
	wire _w33808_ ;
	wire _w33807_ ;
	wire _w33806_ ;
	wire _w33805_ ;
	wire _w33804_ ;
	wire _w33803_ ;
	wire _w33802_ ;
	wire _w33801_ ;
	wire _w33800_ ;
	wire _w33799_ ;
	wire _w33798_ ;
	wire _w33797_ ;
	wire _w33796_ ;
	wire _w33795_ ;
	wire _w33794_ ;
	wire _w33793_ ;
	wire _w33792_ ;
	wire _w33791_ ;
	wire _w33790_ ;
	wire _w33789_ ;
	wire _w33788_ ;
	wire _w33787_ ;
	wire _w33786_ ;
	wire _w33785_ ;
	wire _w33784_ ;
	wire _w33783_ ;
	wire _w33782_ ;
	wire _w33781_ ;
	wire _w33780_ ;
	wire _w33779_ ;
	wire _w33778_ ;
	wire _w33777_ ;
	wire _w33776_ ;
	wire _w33775_ ;
	wire _w33774_ ;
	wire _w33773_ ;
	wire _w33772_ ;
	wire _w33771_ ;
	wire _w33770_ ;
	wire _w33769_ ;
	wire _w33768_ ;
	wire _w33767_ ;
	wire _w33766_ ;
	wire _w33765_ ;
	wire _w33764_ ;
	wire _w33763_ ;
	wire _w33762_ ;
	wire _w33761_ ;
	wire _w33760_ ;
	wire _w33759_ ;
	wire _w33758_ ;
	wire _w33757_ ;
	wire _w33756_ ;
	wire _w33755_ ;
	wire _w33754_ ;
	wire _w33753_ ;
	wire _w33752_ ;
	wire _w33751_ ;
	wire _w33750_ ;
	wire _w33749_ ;
	wire _w33748_ ;
	wire _w33747_ ;
	wire _w33746_ ;
	wire _w33745_ ;
	wire _w33744_ ;
	wire _w33743_ ;
	wire _w33742_ ;
	wire _w33741_ ;
	wire _w33740_ ;
	wire _w33739_ ;
	wire _w33738_ ;
	wire _w33737_ ;
	wire _w33736_ ;
	wire _w33735_ ;
	wire _w33734_ ;
	wire _w33733_ ;
	wire _w33732_ ;
	wire _w33731_ ;
	wire _w33730_ ;
	wire _w33729_ ;
	wire _w33728_ ;
	wire _w33727_ ;
	wire _w33726_ ;
	wire _w33725_ ;
	wire _w33724_ ;
	wire _w33723_ ;
	wire _w33722_ ;
	wire _w33721_ ;
	wire _w33720_ ;
	wire _w33719_ ;
	wire _w33718_ ;
	wire _w33717_ ;
	wire _w33716_ ;
	wire _w33715_ ;
	wire _w33714_ ;
	wire _w33713_ ;
	wire _w33712_ ;
	wire _w33711_ ;
	wire _w33710_ ;
	wire _w33709_ ;
	wire _w33708_ ;
	wire _w33707_ ;
	wire _w33706_ ;
	wire _w33705_ ;
	wire _w33704_ ;
	wire _w33703_ ;
	wire _w33702_ ;
	wire _w33701_ ;
	wire _w33700_ ;
	wire _w33699_ ;
	wire _w33698_ ;
	wire _w33697_ ;
	wire _w33696_ ;
	wire _w33695_ ;
	wire _w33694_ ;
	wire _w33693_ ;
	wire _w33692_ ;
	wire _w33691_ ;
	wire _w33690_ ;
	wire _w33689_ ;
	wire _w33688_ ;
	wire _w33687_ ;
	wire _w33686_ ;
	wire _w33685_ ;
	wire _w33684_ ;
	wire _w33683_ ;
	wire _w33682_ ;
	wire _w33681_ ;
	wire _w33680_ ;
	wire _w33679_ ;
	wire _w33678_ ;
	wire _w33677_ ;
	wire _w33676_ ;
	wire _w33675_ ;
	wire _w33674_ ;
	wire _w33673_ ;
	wire _w33672_ ;
	wire _w33671_ ;
	wire _w33670_ ;
	wire _w33669_ ;
	wire _w33668_ ;
	wire _w33667_ ;
	wire _w33666_ ;
	wire _w33665_ ;
	wire _w33664_ ;
	wire _w33663_ ;
	wire _w33662_ ;
	wire _w33661_ ;
	wire _w33660_ ;
	wire _w33659_ ;
	wire _w33658_ ;
	wire _w33657_ ;
	wire _w33656_ ;
	wire _w33655_ ;
	wire _w33654_ ;
	wire _w33653_ ;
	wire _w33652_ ;
	wire _w33651_ ;
	wire _w33650_ ;
	wire _w33649_ ;
	wire _w33648_ ;
	wire _w33647_ ;
	wire _w33646_ ;
	wire _w33645_ ;
	wire _w33644_ ;
	wire _w33643_ ;
	wire _w33642_ ;
	wire _w33641_ ;
	wire _w33640_ ;
	wire _w33639_ ;
	wire _w33638_ ;
	wire _w33637_ ;
	wire _w33636_ ;
	wire _w33635_ ;
	wire _w33634_ ;
	wire _w33633_ ;
	wire _w33632_ ;
	wire _w33631_ ;
	wire _w33630_ ;
	wire _w33629_ ;
	wire _w33628_ ;
	wire _w33627_ ;
	wire _w33626_ ;
	wire _w33625_ ;
	wire _w33624_ ;
	wire _w33623_ ;
	wire _w33622_ ;
	wire _w33621_ ;
	wire _w33620_ ;
	wire _w33619_ ;
	wire _w33618_ ;
	wire _w33617_ ;
	wire _w33616_ ;
	wire _w33615_ ;
	wire _w33614_ ;
	wire _w33613_ ;
	wire _w33612_ ;
	wire _w33611_ ;
	wire _w33610_ ;
	wire _w33609_ ;
	wire _w33608_ ;
	wire _w33607_ ;
	wire _w33606_ ;
	wire _w33605_ ;
	wire _w33604_ ;
	wire _w33603_ ;
	wire _w33602_ ;
	wire _w33601_ ;
	wire _w33600_ ;
	wire _w33599_ ;
	wire _w33598_ ;
	wire _w33597_ ;
	wire _w33596_ ;
	wire _w33595_ ;
	wire _w33594_ ;
	wire _w33593_ ;
	wire _w33592_ ;
	wire _w33591_ ;
	wire _w33590_ ;
	wire _w33589_ ;
	wire _w33588_ ;
	wire _w33587_ ;
	wire _w33586_ ;
	wire _w33585_ ;
	wire _w33584_ ;
	wire _w33583_ ;
	wire _w33582_ ;
	wire _w33581_ ;
	wire _w33580_ ;
	wire _w33579_ ;
	wire _w33578_ ;
	wire _w33577_ ;
	wire _w33576_ ;
	wire _w33575_ ;
	wire _w33574_ ;
	wire _w33573_ ;
	wire _w33572_ ;
	wire _w33571_ ;
	wire _w33570_ ;
	wire _w33569_ ;
	wire _w33568_ ;
	wire _w33567_ ;
	wire _w33566_ ;
	wire _w33565_ ;
	wire _w33564_ ;
	wire _w33563_ ;
	wire _w33562_ ;
	wire _w33561_ ;
	wire _w33560_ ;
	wire _w33559_ ;
	wire _w33558_ ;
	wire _w33557_ ;
	wire _w33556_ ;
	wire _w33555_ ;
	wire _w33554_ ;
	wire _w33553_ ;
	wire _w33552_ ;
	wire _w33551_ ;
	wire _w33550_ ;
	wire _w33549_ ;
	wire _w33548_ ;
	wire _w33547_ ;
	wire _w33546_ ;
	wire _w33545_ ;
	wire _w33544_ ;
	wire _w33543_ ;
	wire _w33542_ ;
	wire _w33541_ ;
	wire _w33540_ ;
	wire _w33539_ ;
	wire _w33538_ ;
	wire _w33537_ ;
	wire _w33536_ ;
	wire _w33535_ ;
	wire _w33534_ ;
	wire _w33533_ ;
	wire _w33532_ ;
	wire _w33531_ ;
	wire _w33530_ ;
	wire _w33529_ ;
	wire _w33528_ ;
	wire _w33527_ ;
	wire _w33526_ ;
	wire _w33525_ ;
	wire _w33524_ ;
	wire _w33523_ ;
	wire _w33522_ ;
	wire _w33521_ ;
	wire _w33520_ ;
	wire _w33519_ ;
	wire _w33518_ ;
	wire _w33517_ ;
	wire _w33516_ ;
	wire _w33515_ ;
	wire _w33514_ ;
	wire _w33513_ ;
	wire _w33512_ ;
	wire _w33511_ ;
	wire _w33510_ ;
	wire _w33509_ ;
	wire _w33508_ ;
	wire _w33507_ ;
	wire _w33506_ ;
	wire _w33505_ ;
	wire _w33504_ ;
	wire _w33503_ ;
	wire _w33502_ ;
	wire _w33501_ ;
	wire _w33500_ ;
	wire _w33499_ ;
	wire _w33498_ ;
	wire _w33497_ ;
	wire _w33496_ ;
	wire _w33495_ ;
	wire _w33494_ ;
	wire _w33493_ ;
	wire _w33492_ ;
	wire _w33491_ ;
	wire _w33490_ ;
	wire _w33489_ ;
	wire _w33488_ ;
	wire _w33487_ ;
	wire _w33486_ ;
	wire _w33485_ ;
	wire _w33484_ ;
	wire _w33483_ ;
	wire _w33482_ ;
	wire _w33481_ ;
	wire _w33480_ ;
	wire _w33479_ ;
	wire _w33478_ ;
	wire _w33477_ ;
	wire _w33476_ ;
	wire _w33475_ ;
	wire _w33474_ ;
	wire _w33473_ ;
	wire _w33472_ ;
	wire _w33471_ ;
	wire _w33470_ ;
	wire _w33469_ ;
	wire _w33468_ ;
	wire _w33467_ ;
	wire _w33466_ ;
	wire _w33465_ ;
	wire _w33464_ ;
	wire _w33463_ ;
	wire _w33462_ ;
	wire _w33461_ ;
	wire _w33460_ ;
	wire _w33459_ ;
	wire _w33458_ ;
	wire _w33457_ ;
	wire _w33456_ ;
	wire _w33455_ ;
	wire _w33454_ ;
	wire _w33453_ ;
	wire _w33452_ ;
	wire _w33451_ ;
	wire _w33450_ ;
	wire _w33449_ ;
	wire _w33448_ ;
	wire _w33447_ ;
	wire _w33446_ ;
	wire _w33445_ ;
	wire _w33444_ ;
	wire _w33443_ ;
	wire _w33442_ ;
	wire _w33441_ ;
	wire _w33440_ ;
	wire _w33439_ ;
	wire _w33438_ ;
	wire _w33437_ ;
	wire _w33436_ ;
	wire _w33435_ ;
	wire _w33434_ ;
	wire _w33433_ ;
	wire _w33432_ ;
	wire _w33431_ ;
	wire _w33430_ ;
	wire _w33429_ ;
	wire _w33428_ ;
	wire _w33427_ ;
	wire _w33426_ ;
	wire _w33425_ ;
	wire _w33424_ ;
	wire _w33423_ ;
	wire _w33422_ ;
	wire _w33421_ ;
	wire _w33420_ ;
	wire _w33419_ ;
	wire _w33418_ ;
	wire _w33417_ ;
	wire _w33416_ ;
	wire _w33415_ ;
	wire _w33414_ ;
	wire _w33413_ ;
	wire _w33412_ ;
	wire _w33411_ ;
	wire _w33410_ ;
	wire _w33409_ ;
	wire _w33408_ ;
	wire _w33407_ ;
	wire _w33406_ ;
	wire _w33405_ ;
	wire _w33404_ ;
	wire _w33403_ ;
	wire _w33402_ ;
	wire _w33401_ ;
	wire _w33400_ ;
	wire _w33399_ ;
	wire _w33398_ ;
	wire _w33397_ ;
	wire _w33396_ ;
	wire _w33395_ ;
	wire _w33394_ ;
	wire _w33393_ ;
	wire _w33392_ ;
	wire _w33391_ ;
	wire _w33390_ ;
	wire _w33389_ ;
	wire _w33388_ ;
	wire _w33387_ ;
	wire _w33386_ ;
	wire _w33385_ ;
	wire _w33384_ ;
	wire _w33383_ ;
	wire _w33382_ ;
	wire _w33381_ ;
	wire _w33380_ ;
	wire _w33379_ ;
	wire _w33378_ ;
	wire _w33377_ ;
	wire _w33376_ ;
	wire _w33375_ ;
	wire _w33374_ ;
	wire _w33373_ ;
	wire _w33372_ ;
	wire _w33371_ ;
	wire _w33370_ ;
	wire _w33369_ ;
	wire _w33368_ ;
	wire _w33367_ ;
	wire _w33366_ ;
	wire _w33365_ ;
	wire _w33364_ ;
	wire _w33363_ ;
	wire _w33362_ ;
	wire _w33361_ ;
	wire _w33360_ ;
	wire _w33359_ ;
	wire _w33358_ ;
	wire _w33357_ ;
	wire _w33356_ ;
	wire _w33355_ ;
	wire _w33354_ ;
	wire _w33353_ ;
	wire _w33352_ ;
	wire _w33351_ ;
	wire _w33350_ ;
	wire _w33349_ ;
	wire _w33348_ ;
	wire _w33347_ ;
	wire _w33346_ ;
	wire _w33345_ ;
	wire _w33344_ ;
	wire _w33343_ ;
	wire _w33342_ ;
	wire _w33341_ ;
	wire _w33340_ ;
	wire _w33339_ ;
	wire _w33338_ ;
	wire _w33337_ ;
	wire _w33336_ ;
	wire _w33335_ ;
	wire _w33334_ ;
	wire _w33333_ ;
	wire _w33332_ ;
	wire _w33331_ ;
	wire _w33330_ ;
	wire _w33329_ ;
	wire _w33328_ ;
	wire _w33327_ ;
	wire _w33326_ ;
	wire _w33325_ ;
	wire _w33324_ ;
	wire _w33323_ ;
	wire _w33322_ ;
	wire _w33321_ ;
	wire _w33320_ ;
	wire _w33319_ ;
	wire _w33318_ ;
	wire _w33317_ ;
	wire _w33316_ ;
	wire _w33315_ ;
	wire _w33314_ ;
	wire _w33313_ ;
	wire _w33312_ ;
	wire _w33311_ ;
	wire _w33310_ ;
	wire _w33309_ ;
	wire _w33308_ ;
	wire _w33307_ ;
	wire _w33306_ ;
	wire _w33305_ ;
	wire _w33304_ ;
	wire _w33303_ ;
	wire _w33302_ ;
	wire _w33301_ ;
	wire _w33300_ ;
	wire _w33299_ ;
	wire _w33298_ ;
	wire _w33297_ ;
	wire _w33296_ ;
	wire _w33295_ ;
	wire _w33294_ ;
	wire _w33293_ ;
	wire _w33292_ ;
	wire _w33291_ ;
	wire _w33290_ ;
	wire _w33289_ ;
	wire _w33288_ ;
	wire _w33287_ ;
	wire _w33286_ ;
	wire _w33285_ ;
	wire _w33284_ ;
	wire _w33283_ ;
	wire _w33282_ ;
	wire _w33281_ ;
	wire _w33280_ ;
	wire _w33279_ ;
	wire _w33278_ ;
	wire _w33277_ ;
	wire _w33276_ ;
	wire _w33275_ ;
	wire _w33274_ ;
	wire _w33273_ ;
	wire _w33272_ ;
	wire _w33271_ ;
	wire _w33270_ ;
	wire _w33269_ ;
	wire _w33268_ ;
	wire _w33267_ ;
	wire _w33266_ ;
	wire _w33265_ ;
	wire _w33264_ ;
	wire _w33263_ ;
	wire _w33262_ ;
	wire _w33261_ ;
	wire _w33260_ ;
	wire _w33259_ ;
	wire _w33258_ ;
	wire _w33257_ ;
	wire _w33256_ ;
	wire _w33255_ ;
	wire _w33254_ ;
	wire _w33253_ ;
	wire _w33252_ ;
	wire _w33251_ ;
	wire _w33250_ ;
	wire _w33249_ ;
	wire _w33248_ ;
	wire _w33247_ ;
	wire _w33246_ ;
	wire _w33245_ ;
	wire _w33244_ ;
	wire _w33243_ ;
	wire _w33242_ ;
	wire _w33241_ ;
	wire _w33240_ ;
	wire _w33239_ ;
	wire _w33238_ ;
	wire _w33237_ ;
	wire _w33236_ ;
	wire _w33235_ ;
	wire _w33234_ ;
	wire _w33233_ ;
	wire _w33232_ ;
	wire _w33231_ ;
	wire _w33230_ ;
	wire _w33229_ ;
	wire _w33228_ ;
	wire _w33227_ ;
	wire _w33226_ ;
	wire _w33225_ ;
	wire _w33224_ ;
	wire _w33223_ ;
	wire _w33222_ ;
	wire _w33221_ ;
	wire _w33220_ ;
	wire _w33219_ ;
	wire _w33218_ ;
	wire _w33217_ ;
	wire _w33216_ ;
	wire _w33215_ ;
	wire _w33214_ ;
	wire _w33213_ ;
	wire _w33212_ ;
	wire _w33211_ ;
	wire _w33210_ ;
	wire _w33209_ ;
	wire _w33208_ ;
	wire _w33207_ ;
	wire _w33206_ ;
	wire _w33205_ ;
	wire _w33204_ ;
	wire _w33203_ ;
	wire _w33202_ ;
	wire _w33201_ ;
	wire _w33200_ ;
	wire _w33199_ ;
	wire _w33198_ ;
	wire _w33197_ ;
	wire _w33196_ ;
	wire _w33195_ ;
	wire _w33194_ ;
	wire _w33193_ ;
	wire _w33192_ ;
	wire _w33191_ ;
	wire _w33190_ ;
	wire _w33189_ ;
	wire _w33188_ ;
	wire _w33187_ ;
	wire _w33186_ ;
	wire _w33185_ ;
	wire _w33184_ ;
	wire _w33183_ ;
	wire _w33182_ ;
	wire _w33181_ ;
	wire _w33180_ ;
	wire _w33179_ ;
	wire _w33178_ ;
	wire _w33177_ ;
	wire _w33176_ ;
	wire _w33175_ ;
	wire _w33174_ ;
	wire _w33173_ ;
	wire _w33172_ ;
	wire _w33171_ ;
	wire _w33170_ ;
	wire _w33169_ ;
	wire _w33168_ ;
	wire _w33167_ ;
	wire _w33166_ ;
	wire _w33165_ ;
	wire _w33164_ ;
	wire _w33163_ ;
	wire _w33162_ ;
	wire _w33161_ ;
	wire _w33160_ ;
	wire _w33159_ ;
	wire _w33158_ ;
	wire _w33157_ ;
	wire _w33156_ ;
	wire _w33155_ ;
	wire _w33154_ ;
	wire _w33153_ ;
	wire _w33152_ ;
	wire _w33151_ ;
	wire _w33150_ ;
	wire _w33149_ ;
	wire _w33148_ ;
	wire _w33147_ ;
	wire _w33146_ ;
	wire _w33145_ ;
	wire _w33144_ ;
	wire _w33143_ ;
	wire _w33142_ ;
	wire _w33141_ ;
	wire _w33140_ ;
	wire _w33139_ ;
	wire _w33138_ ;
	wire _w33137_ ;
	wire _w33136_ ;
	wire _w33135_ ;
	wire _w33134_ ;
	wire _w33133_ ;
	wire _w33132_ ;
	wire _w33131_ ;
	wire _w33130_ ;
	wire _w33129_ ;
	wire _w33128_ ;
	wire _w33127_ ;
	wire _w33126_ ;
	wire _w33125_ ;
	wire _w33124_ ;
	wire _w33123_ ;
	wire _w33122_ ;
	wire _w33121_ ;
	wire _w33120_ ;
	wire _w33119_ ;
	wire _w33118_ ;
	wire _w33117_ ;
	wire _w33116_ ;
	wire _w33115_ ;
	wire _w33114_ ;
	wire _w33113_ ;
	wire _w33112_ ;
	wire _w33111_ ;
	wire _w33110_ ;
	wire _w33109_ ;
	wire _w33108_ ;
	wire _w33107_ ;
	wire _w33106_ ;
	wire _w33105_ ;
	wire _w33104_ ;
	wire _w33103_ ;
	wire _w33102_ ;
	wire _w33101_ ;
	wire _w33100_ ;
	wire _w33099_ ;
	wire _w33098_ ;
	wire _w33097_ ;
	wire _w33096_ ;
	wire _w33095_ ;
	wire _w33094_ ;
	wire _w33093_ ;
	wire _w33092_ ;
	wire _w33091_ ;
	wire _w33090_ ;
	wire _w33089_ ;
	wire _w33088_ ;
	wire _w33087_ ;
	wire _w33086_ ;
	wire _w33085_ ;
	wire _w33084_ ;
	wire _w33083_ ;
	wire _w33082_ ;
	wire _w33081_ ;
	wire _w33080_ ;
	wire _w33079_ ;
	wire _w33078_ ;
	wire _w33077_ ;
	wire _w33076_ ;
	wire _w33075_ ;
	wire _w33074_ ;
	wire _w33073_ ;
	wire _w33072_ ;
	wire _w33071_ ;
	wire _w33070_ ;
	wire _w33069_ ;
	wire _w33068_ ;
	wire _w33067_ ;
	wire _w33066_ ;
	wire _w33065_ ;
	wire _w33064_ ;
	wire _w33063_ ;
	wire _w33062_ ;
	wire _w33061_ ;
	wire _w33060_ ;
	wire _w33059_ ;
	wire _w33058_ ;
	wire _w33057_ ;
	wire _w33056_ ;
	wire _w33055_ ;
	wire _w33054_ ;
	wire _w33053_ ;
	wire _w33052_ ;
	wire _w33051_ ;
	wire _w33050_ ;
	wire _w33049_ ;
	wire _w33048_ ;
	wire _w33047_ ;
	wire _w33046_ ;
	wire _w33045_ ;
	wire _w33044_ ;
	wire _w33043_ ;
	wire _w33042_ ;
	wire _w33041_ ;
	wire _w33040_ ;
	wire _w33039_ ;
	wire _w33038_ ;
	wire _w33037_ ;
	wire _w33036_ ;
	wire _w33035_ ;
	wire _w33034_ ;
	wire _w33033_ ;
	wire _w33032_ ;
	wire _w33031_ ;
	wire _w33030_ ;
	wire _w33029_ ;
	wire _w33028_ ;
	wire _w33027_ ;
	wire _w33026_ ;
	wire _w33025_ ;
	wire _w33024_ ;
	wire _w33023_ ;
	wire _w33022_ ;
	wire _w33021_ ;
	wire _w33020_ ;
	wire _w33019_ ;
	wire _w33018_ ;
	wire _w33017_ ;
	wire _w33016_ ;
	wire _w33015_ ;
	wire _w33014_ ;
	wire _w33013_ ;
	wire _w33012_ ;
	wire _w33011_ ;
	wire _w33010_ ;
	wire _w33009_ ;
	wire _w33008_ ;
	wire _w33007_ ;
	wire _w33006_ ;
	wire _w33005_ ;
	wire _w33004_ ;
	wire _w33003_ ;
	wire _w33002_ ;
	wire _w33001_ ;
	wire _w33000_ ;
	wire _w32999_ ;
	wire _w32998_ ;
	wire _w32997_ ;
	wire _w32996_ ;
	wire _w32995_ ;
	wire _w32994_ ;
	wire _w32993_ ;
	wire _w32992_ ;
	wire _w32991_ ;
	wire _w32990_ ;
	wire _w32989_ ;
	wire _w32988_ ;
	wire _w32987_ ;
	wire _w32986_ ;
	wire _w32985_ ;
	wire _w32984_ ;
	wire _w32983_ ;
	wire _w32982_ ;
	wire _w32981_ ;
	wire _w32980_ ;
	wire _w32979_ ;
	wire _w32978_ ;
	wire _w32977_ ;
	wire _w32976_ ;
	wire _w32975_ ;
	wire _w32974_ ;
	wire _w32973_ ;
	wire _w32972_ ;
	wire _w32971_ ;
	wire _w32970_ ;
	wire _w32969_ ;
	wire _w32968_ ;
	wire _w32967_ ;
	wire _w32966_ ;
	wire _w32965_ ;
	wire _w32964_ ;
	wire _w32963_ ;
	wire _w32962_ ;
	wire _w32961_ ;
	wire _w32960_ ;
	wire _w32959_ ;
	wire _w32958_ ;
	wire _w32957_ ;
	wire _w32956_ ;
	wire _w32955_ ;
	wire _w32954_ ;
	wire _w32953_ ;
	wire _w32952_ ;
	wire _w32951_ ;
	wire _w32950_ ;
	wire _w32949_ ;
	wire _w32948_ ;
	wire _w32947_ ;
	wire _w32946_ ;
	wire _w32945_ ;
	wire _w32944_ ;
	wire _w32943_ ;
	wire _w32942_ ;
	wire _w32941_ ;
	wire _w32940_ ;
	wire _w32939_ ;
	wire _w32938_ ;
	wire _w32937_ ;
	wire _w32936_ ;
	wire _w32935_ ;
	wire _w32934_ ;
	wire _w32933_ ;
	wire _w32932_ ;
	wire _w32931_ ;
	wire _w32930_ ;
	wire _w32929_ ;
	wire _w32928_ ;
	wire _w32927_ ;
	wire _w32926_ ;
	wire _w32925_ ;
	wire _w32924_ ;
	wire _w32923_ ;
	wire _w32922_ ;
	wire _w32921_ ;
	wire _w32920_ ;
	wire _w32919_ ;
	wire _w32918_ ;
	wire _w32917_ ;
	wire _w32916_ ;
	wire _w32915_ ;
	wire _w32914_ ;
	wire _w32913_ ;
	wire _w32912_ ;
	wire _w32911_ ;
	wire _w32910_ ;
	wire _w32909_ ;
	wire _w32908_ ;
	wire _w32907_ ;
	wire _w32906_ ;
	wire _w32905_ ;
	wire _w32904_ ;
	wire _w32903_ ;
	wire _w32902_ ;
	wire _w32901_ ;
	wire _w32900_ ;
	wire _w32899_ ;
	wire _w32898_ ;
	wire _w32897_ ;
	wire _w32896_ ;
	wire _w32895_ ;
	wire _w32894_ ;
	wire _w32893_ ;
	wire _w32892_ ;
	wire _w32891_ ;
	wire _w32890_ ;
	wire _w32889_ ;
	wire _w32888_ ;
	wire _w32887_ ;
	wire _w32886_ ;
	wire _w32885_ ;
	wire _w32884_ ;
	wire _w32883_ ;
	wire _w32882_ ;
	wire _w32881_ ;
	wire _w32880_ ;
	wire _w32879_ ;
	wire _w32878_ ;
	wire _w32877_ ;
	wire _w32876_ ;
	wire _w32875_ ;
	wire _w32874_ ;
	wire _w32873_ ;
	wire _w32872_ ;
	wire _w32871_ ;
	wire _w32870_ ;
	wire _w32869_ ;
	wire _w32868_ ;
	wire _w32867_ ;
	wire _w32866_ ;
	wire _w32865_ ;
	wire _w32864_ ;
	wire _w32863_ ;
	wire _w32862_ ;
	wire _w32861_ ;
	wire _w32860_ ;
	wire _w32859_ ;
	wire _w32858_ ;
	wire _w32857_ ;
	wire _w32856_ ;
	wire _w32855_ ;
	wire _w32854_ ;
	wire _w32853_ ;
	wire _w32852_ ;
	wire _w32851_ ;
	wire _w32850_ ;
	wire _w32849_ ;
	wire _w32848_ ;
	wire _w32847_ ;
	wire _w32846_ ;
	wire _w32845_ ;
	wire _w32844_ ;
	wire _w32843_ ;
	wire _w32842_ ;
	wire _w32841_ ;
	wire _w32840_ ;
	wire _w32839_ ;
	wire _w32838_ ;
	wire _w32837_ ;
	wire _w32836_ ;
	wire _w32835_ ;
	wire _w32834_ ;
	wire _w32833_ ;
	wire _w32832_ ;
	wire _w32831_ ;
	wire _w32830_ ;
	wire _w32829_ ;
	wire _w32828_ ;
	wire _w32827_ ;
	wire _w32826_ ;
	wire _w32825_ ;
	wire _w32824_ ;
	wire _w32823_ ;
	wire _w32822_ ;
	wire _w32821_ ;
	wire _w32820_ ;
	wire _w32819_ ;
	wire _w32818_ ;
	wire _w32817_ ;
	wire _w32816_ ;
	wire _w32815_ ;
	wire _w32814_ ;
	wire _w32813_ ;
	wire _w32812_ ;
	wire _w32811_ ;
	wire _w32810_ ;
	wire _w32809_ ;
	wire _w32808_ ;
	wire _w32807_ ;
	wire _w32806_ ;
	wire _w32805_ ;
	wire _w32804_ ;
	wire _w32803_ ;
	wire _w32802_ ;
	wire _w32801_ ;
	wire _w32800_ ;
	wire _w32799_ ;
	wire _w32798_ ;
	wire _w32797_ ;
	wire _w32796_ ;
	wire _w32795_ ;
	wire _w32794_ ;
	wire _w32793_ ;
	wire _w32792_ ;
	wire _w32791_ ;
	wire _w32790_ ;
	wire _w32789_ ;
	wire _w32788_ ;
	wire _w32787_ ;
	wire _w32786_ ;
	wire _w32785_ ;
	wire _w32784_ ;
	wire _w32783_ ;
	wire _w32782_ ;
	wire _w32781_ ;
	wire _w32780_ ;
	wire _w32779_ ;
	wire _w32778_ ;
	wire _w32777_ ;
	wire _w32776_ ;
	wire _w32775_ ;
	wire _w32774_ ;
	wire _w32773_ ;
	wire _w32772_ ;
	wire _w32771_ ;
	wire _w32770_ ;
	wire _w32769_ ;
	wire _w32768_ ;
	wire _w32767_ ;
	wire _w32766_ ;
	wire _w32765_ ;
	wire _w32764_ ;
	wire _w32763_ ;
	wire _w32762_ ;
	wire _w32761_ ;
	wire _w32760_ ;
	wire _w32759_ ;
	wire _w32758_ ;
	wire _w32757_ ;
	wire _w32756_ ;
	wire _w32755_ ;
	wire _w32754_ ;
	wire _w32753_ ;
	wire _w32752_ ;
	wire _w32751_ ;
	wire _w32750_ ;
	wire _w32749_ ;
	wire _w32748_ ;
	wire _w32747_ ;
	wire _w32746_ ;
	wire _w32745_ ;
	wire _w32744_ ;
	wire _w32743_ ;
	wire _w32742_ ;
	wire _w32741_ ;
	wire _w32740_ ;
	wire _w32739_ ;
	wire _w32738_ ;
	wire _w32737_ ;
	wire _w32736_ ;
	wire _w32735_ ;
	wire _w32734_ ;
	wire _w32733_ ;
	wire _w32732_ ;
	wire _w32731_ ;
	wire _w32730_ ;
	wire _w32729_ ;
	wire _w32728_ ;
	wire _w32727_ ;
	wire _w32726_ ;
	wire _w32725_ ;
	wire _w32724_ ;
	wire _w32723_ ;
	wire _w32722_ ;
	wire _w32721_ ;
	wire _w32720_ ;
	wire _w32719_ ;
	wire _w32718_ ;
	wire _w32717_ ;
	wire _w32716_ ;
	wire _w32715_ ;
	wire _w32714_ ;
	wire _w32713_ ;
	wire _w32712_ ;
	wire _w32711_ ;
	wire _w32710_ ;
	wire _w32709_ ;
	wire _w32708_ ;
	wire _w32707_ ;
	wire _w32706_ ;
	wire _w32705_ ;
	wire _w32704_ ;
	wire _w32703_ ;
	wire _w32702_ ;
	wire _w32701_ ;
	wire _w32700_ ;
	wire _w32699_ ;
	wire _w32698_ ;
	wire _w32697_ ;
	wire _w32696_ ;
	wire _w32695_ ;
	wire _w32694_ ;
	wire _w32693_ ;
	wire _w32692_ ;
	wire _w32691_ ;
	wire _w32690_ ;
	wire _w32689_ ;
	wire _w32688_ ;
	wire _w32687_ ;
	wire _w32686_ ;
	wire _w32685_ ;
	wire _w32684_ ;
	wire _w32683_ ;
	wire _w32682_ ;
	wire _w32681_ ;
	wire _w32680_ ;
	wire _w32679_ ;
	wire _w32678_ ;
	wire _w32677_ ;
	wire _w32676_ ;
	wire _w32675_ ;
	wire _w32674_ ;
	wire _w32673_ ;
	wire _w32672_ ;
	wire _w32671_ ;
	wire _w32670_ ;
	wire _w32669_ ;
	wire _w32668_ ;
	wire _w32667_ ;
	wire _w32666_ ;
	wire _w32665_ ;
	wire _w32664_ ;
	wire _w32663_ ;
	wire _w32662_ ;
	wire _w32661_ ;
	wire _w32660_ ;
	wire _w32659_ ;
	wire _w32658_ ;
	wire _w32657_ ;
	wire _w32656_ ;
	wire _w32655_ ;
	wire _w32654_ ;
	wire _w32653_ ;
	wire _w32652_ ;
	wire _w32651_ ;
	wire _w32650_ ;
	wire _w32649_ ;
	wire _w32648_ ;
	wire _w32647_ ;
	wire _w32646_ ;
	wire _w32645_ ;
	wire _w32644_ ;
	wire _w32643_ ;
	wire _w32642_ ;
	wire _w32641_ ;
	wire _w32640_ ;
	wire _w32639_ ;
	wire _w32638_ ;
	wire _w32637_ ;
	wire _w32636_ ;
	wire _w32635_ ;
	wire _w32634_ ;
	wire _w32633_ ;
	wire _w32632_ ;
	wire _w32631_ ;
	wire _w32630_ ;
	wire _w32629_ ;
	wire _w32628_ ;
	wire _w32627_ ;
	wire _w32626_ ;
	wire _w32625_ ;
	wire _w32624_ ;
	wire _w32623_ ;
	wire _w32622_ ;
	wire _w32621_ ;
	wire _w32620_ ;
	wire _w32619_ ;
	wire _w32618_ ;
	wire _w32617_ ;
	wire _w32616_ ;
	wire _w32615_ ;
	wire _w32614_ ;
	wire _w32613_ ;
	wire _w32612_ ;
	wire _w32611_ ;
	wire _w32610_ ;
	wire _w32609_ ;
	wire _w32608_ ;
	wire _w32607_ ;
	wire _w32606_ ;
	wire _w32605_ ;
	wire _w32604_ ;
	wire _w32603_ ;
	wire _w32602_ ;
	wire _w32601_ ;
	wire _w32600_ ;
	wire _w32599_ ;
	wire _w32598_ ;
	wire _w32597_ ;
	wire _w32596_ ;
	wire _w32595_ ;
	wire _w32594_ ;
	wire _w32593_ ;
	wire _w32592_ ;
	wire _w32591_ ;
	wire _w32590_ ;
	wire _w32589_ ;
	wire _w32588_ ;
	wire _w32587_ ;
	wire _w32586_ ;
	wire _w32585_ ;
	wire _w32584_ ;
	wire _w32583_ ;
	wire _w32582_ ;
	wire _w32581_ ;
	wire _w32580_ ;
	wire _w32579_ ;
	wire _w32578_ ;
	wire _w32577_ ;
	wire _w32576_ ;
	wire _w32575_ ;
	wire _w32574_ ;
	wire _w32573_ ;
	wire _w32572_ ;
	wire _w32571_ ;
	wire _w32570_ ;
	wire _w32569_ ;
	wire _w32568_ ;
	wire _w32567_ ;
	wire _w32566_ ;
	wire _w32565_ ;
	wire _w32564_ ;
	wire _w32563_ ;
	wire _w32562_ ;
	wire _w32561_ ;
	wire _w32560_ ;
	wire _w32559_ ;
	wire _w32558_ ;
	wire _w32557_ ;
	wire _w32556_ ;
	wire _w32555_ ;
	wire _w32554_ ;
	wire _w32553_ ;
	wire _w32552_ ;
	wire _w32551_ ;
	wire _w32550_ ;
	wire _w32549_ ;
	wire _w32548_ ;
	wire _w32547_ ;
	wire _w32546_ ;
	wire _w32545_ ;
	wire _w32544_ ;
	wire _w32543_ ;
	wire _w32542_ ;
	wire _w32541_ ;
	wire _w32540_ ;
	wire _w32539_ ;
	wire _w32538_ ;
	wire _w32537_ ;
	wire _w32536_ ;
	wire _w32535_ ;
	wire _w32534_ ;
	wire _w32533_ ;
	wire _w32532_ ;
	wire _w32531_ ;
	wire _w32530_ ;
	wire _w32529_ ;
	wire _w32528_ ;
	wire _w32527_ ;
	wire _w32526_ ;
	wire _w32525_ ;
	wire _w32524_ ;
	wire _w32523_ ;
	wire _w32522_ ;
	wire _w32521_ ;
	wire _w32520_ ;
	wire _w32519_ ;
	wire _w32518_ ;
	wire _w32517_ ;
	wire _w32516_ ;
	wire _w32515_ ;
	wire _w32514_ ;
	wire _w32513_ ;
	wire _w32512_ ;
	wire _w32511_ ;
	wire _w32510_ ;
	wire _w32509_ ;
	wire _w32508_ ;
	wire _w32507_ ;
	wire _w32506_ ;
	wire _w32505_ ;
	wire _w32504_ ;
	wire _w32503_ ;
	wire _w32502_ ;
	wire _w32501_ ;
	wire _w32500_ ;
	wire _w32499_ ;
	wire _w32498_ ;
	wire _w32497_ ;
	wire _w32496_ ;
	wire _w32495_ ;
	wire _w32494_ ;
	wire _w32493_ ;
	wire _w32492_ ;
	wire _w32491_ ;
	wire _w32490_ ;
	wire _w32489_ ;
	wire _w32488_ ;
	wire _w32487_ ;
	wire _w32486_ ;
	wire _w32485_ ;
	wire _w32484_ ;
	wire _w32483_ ;
	wire _w32482_ ;
	wire _w32481_ ;
	wire _w32480_ ;
	wire _w32479_ ;
	wire _w32478_ ;
	wire _w32477_ ;
	wire _w32476_ ;
	wire _w32475_ ;
	wire _w32474_ ;
	wire _w32473_ ;
	wire _w32472_ ;
	wire _w32471_ ;
	wire _w32470_ ;
	wire _w32469_ ;
	wire _w32468_ ;
	wire _w32467_ ;
	wire _w32466_ ;
	wire _w32465_ ;
	wire _w32464_ ;
	wire _w32463_ ;
	wire _w32462_ ;
	wire _w32461_ ;
	wire _w32460_ ;
	wire _w32459_ ;
	wire _w32458_ ;
	wire _w32457_ ;
	wire _w32456_ ;
	wire _w32455_ ;
	wire _w32454_ ;
	wire _w32453_ ;
	wire _w32452_ ;
	wire _w32451_ ;
	wire _w32450_ ;
	wire _w32449_ ;
	wire _w32448_ ;
	wire _w32447_ ;
	wire _w32446_ ;
	wire _w32445_ ;
	wire _w32444_ ;
	wire _w32443_ ;
	wire _w32442_ ;
	wire _w32441_ ;
	wire _w32440_ ;
	wire _w32439_ ;
	wire _w32438_ ;
	wire _w32437_ ;
	wire _w32436_ ;
	wire _w32435_ ;
	wire _w32434_ ;
	wire _w32433_ ;
	wire _w32432_ ;
	wire _w32431_ ;
	wire _w32430_ ;
	wire _w32429_ ;
	wire _w32428_ ;
	wire _w32427_ ;
	wire _w32426_ ;
	wire _w32425_ ;
	wire _w32424_ ;
	wire _w32423_ ;
	wire _w32422_ ;
	wire _w32421_ ;
	wire _w32420_ ;
	wire _w32419_ ;
	wire _w32418_ ;
	wire _w32417_ ;
	wire _w32416_ ;
	wire _w32415_ ;
	wire _w32414_ ;
	wire _w32413_ ;
	wire _w32412_ ;
	wire _w32411_ ;
	wire _w32410_ ;
	wire _w32409_ ;
	wire _w32408_ ;
	wire _w32407_ ;
	wire _w32406_ ;
	wire _w32405_ ;
	wire _w32404_ ;
	wire _w32403_ ;
	wire _w32402_ ;
	wire _w32401_ ;
	wire _w32400_ ;
	wire _w32399_ ;
	wire _w32398_ ;
	wire _w32397_ ;
	wire _w32396_ ;
	wire _w32395_ ;
	wire _w32394_ ;
	wire _w32393_ ;
	wire _w32392_ ;
	wire _w32391_ ;
	wire _w32390_ ;
	wire _w32389_ ;
	wire _w32388_ ;
	wire _w32387_ ;
	wire _w32386_ ;
	wire _w32385_ ;
	wire _w32384_ ;
	wire _w32383_ ;
	wire _w32382_ ;
	wire _w32381_ ;
	wire _w32380_ ;
	wire _w32379_ ;
	wire _w32378_ ;
	wire _w32377_ ;
	wire _w32376_ ;
	wire _w32375_ ;
	wire _w32374_ ;
	wire _w32373_ ;
	wire _w32372_ ;
	wire _w32371_ ;
	wire _w32370_ ;
	wire _w32369_ ;
	wire _w32368_ ;
	wire _w32367_ ;
	wire _w32366_ ;
	wire _w32365_ ;
	wire _w32364_ ;
	wire _w32363_ ;
	wire _w32362_ ;
	wire _w32361_ ;
	wire _w32360_ ;
	wire _w32359_ ;
	wire _w32358_ ;
	wire _w32357_ ;
	wire _w32356_ ;
	wire _w32355_ ;
	wire _w32354_ ;
	wire _w32353_ ;
	wire _w32352_ ;
	wire _w32351_ ;
	wire _w32350_ ;
	wire _w32349_ ;
	wire _w32348_ ;
	wire _w32347_ ;
	wire _w32346_ ;
	wire _w32345_ ;
	wire _w32344_ ;
	wire _w32343_ ;
	wire _w32342_ ;
	wire _w32341_ ;
	wire _w32340_ ;
	wire _w32339_ ;
	wire _w32338_ ;
	wire _w32337_ ;
	wire _w32336_ ;
	wire _w32335_ ;
	wire _w32334_ ;
	wire _w32333_ ;
	wire _w32332_ ;
	wire _w32331_ ;
	wire _w32330_ ;
	wire _w32329_ ;
	wire _w32328_ ;
	wire _w32327_ ;
	wire _w32326_ ;
	wire _w32325_ ;
	wire _w32324_ ;
	wire _w32323_ ;
	wire _w32322_ ;
	wire _w32321_ ;
	wire _w32320_ ;
	wire _w32319_ ;
	wire _w32318_ ;
	wire _w32317_ ;
	wire _w32316_ ;
	wire _w32315_ ;
	wire _w32314_ ;
	wire _w32313_ ;
	wire _w32312_ ;
	wire _w32311_ ;
	wire _w32310_ ;
	wire _w32309_ ;
	wire _w32308_ ;
	wire _w32307_ ;
	wire _w32306_ ;
	wire _w32305_ ;
	wire _w32304_ ;
	wire _w32303_ ;
	wire _w32302_ ;
	wire _w32301_ ;
	wire _w32300_ ;
	wire _w32299_ ;
	wire _w32298_ ;
	wire _w32297_ ;
	wire _w32296_ ;
	wire _w32295_ ;
	wire _w32294_ ;
	wire _w32293_ ;
	wire _w32292_ ;
	wire _w32291_ ;
	wire _w32290_ ;
	wire _w32289_ ;
	wire _w32288_ ;
	wire _w32287_ ;
	wire _w32286_ ;
	wire _w32285_ ;
	wire _w32284_ ;
	wire _w32283_ ;
	wire _w32282_ ;
	wire _w32281_ ;
	wire _w32280_ ;
	wire _w32279_ ;
	wire _w32278_ ;
	wire _w32277_ ;
	wire _w32276_ ;
	wire _w32275_ ;
	wire _w32274_ ;
	wire _w32273_ ;
	wire _w32272_ ;
	wire _w32271_ ;
	wire _w32270_ ;
	wire _w32269_ ;
	wire _w32268_ ;
	wire _w32267_ ;
	wire _w32266_ ;
	wire _w32265_ ;
	wire _w32264_ ;
	wire _w32263_ ;
	wire _w32262_ ;
	wire _w32261_ ;
	wire _w32260_ ;
	wire _w32259_ ;
	wire _w32258_ ;
	wire _w32257_ ;
	wire _w32256_ ;
	wire _w32255_ ;
	wire _w32254_ ;
	wire _w32253_ ;
	wire _w32252_ ;
	wire _w32251_ ;
	wire _w32250_ ;
	wire _w32249_ ;
	wire _w32248_ ;
	wire _w32247_ ;
	wire _w32246_ ;
	wire _w32245_ ;
	wire _w32244_ ;
	wire _w32243_ ;
	wire _w32242_ ;
	wire _w32241_ ;
	wire _w32240_ ;
	wire _w32239_ ;
	wire _w32238_ ;
	wire _w32237_ ;
	wire _w32236_ ;
	wire _w32235_ ;
	wire _w32234_ ;
	wire _w32233_ ;
	wire _w32232_ ;
	wire _w32231_ ;
	wire _w32230_ ;
	wire _w32229_ ;
	wire _w32228_ ;
	wire _w32227_ ;
	wire _w32226_ ;
	wire _w32225_ ;
	wire _w32224_ ;
	wire _w32223_ ;
	wire _w32222_ ;
	wire _w32221_ ;
	wire _w32220_ ;
	wire _w32219_ ;
	wire _w32218_ ;
	wire _w32217_ ;
	wire _w32216_ ;
	wire _w32215_ ;
	wire _w32214_ ;
	wire _w32213_ ;
	wire _w32212_ ;
	wire _w32211_ ;
	wire _w32210_ ;
	wire _w32209_ ;
	wire _w32208_ ;
	wire _w32207_ ;
	wire _w32206_ ;
	wire _w32205_ ;
	wire _w32204_ ;
	wire _w32203_ ;
	wire _w32202_ ;
	wire _w32201_ ;
	wire _w32200_ ;
	wire _w32199_ ;
	wire _w32198_ ;
	wire _w32197_ ;
	wire _w32196_ ;
	wire _w32195_ ;
	wire _w32194_ ;
	wire _w32193_ ;
	wire _w32192_ ;
	wire _w32191_ ;
	wire _w32190_ ;
	wire _w32189_ ;
	wire _w32188_ ;
	wire _w32187_ ;
	wire _w32186_ ;
	wire _w32185_ ;
	wire _w32184_ ;
	wire _w32183_ ;
	wire _w32182_ ;
	wire _w32181_ ;
	wire _w32180_ ;
	wire _w32179_ ;
	wire _w32178_ ;
	wire _w32177_ ;
	wire _w32176_ ;
	wire _w32175_ ;
	wire _w32174_ ;
	wire _w32173_ ;
	wire _w32172_ ;
	wire _w32171_ ;
	wire _w32170_ ;
	wire _w32169_ ;
	wire _w32168_ ;
	wire _w32167_ ;
	wire _w32166_ ;
	wire _w32165_ ;
	wire _w32164_ ;
	wire _w32163_ ;
	wire _w32162_ ;
	wire _w32161_ ;
	wire _w32160_ ;
	wire _w32159_ ;
	wire _w32158_ ;
	wire _w32157_ ;
	wire _w32156_ ;
	wire _w32155_ ;
	wire _w32154_ ;
	wire _w32153_ ;
	wire _w32152_ ;
	wire _w32151_ ;
	wire _w32150_ ;
	wire _w32149_ ;
	wire _w32148_ ;
	wire _w32147_ ;
	wire _w32146_ ;
	wire _w32145_ ;
	wire _w32144_ ;
	wire _w32143_ ;
	wire _w32142_ ;
	wire _w32141_ ;
	wire _w32140_ ;
	wire _w32139_ ;
	wire _w32138_ ;
	wire _w32137_ ;
	wire _w32136_ ;
	wire _w32135_ ;
	wire _w32134_ ;
	wire _w32133_ ;
	wire _w32132_ ;
	wire _w32131_ ;
	wire _w32130_ ;
	wire _w32129_ ;
	wire _w32128_ ;
	wire _w32127_ ;
	wire _w32126_ ;
	wire _w32125_ ;
	wire _w32124_ ;
	wire _w32123_ ;
	wire _w32122_ ;
	wire _w32121_ ;
	wire _w32120_ ;
	wire _w32119_ ;
	wire _w32118_ ;
	wire _w32117_ ;
	wire _w32116_ ;
	wire _w32115_ ;
	wire _w32114_ ;
	wire _w32113_ ;
	wire _w32112_ ;
	wire _w32111_ ;
	wire _w32110_ ;
	wire _w32109_ ;
	wire _w32108_ ;
	wire _w32107_ ;
	wire _w32106_ ;
	wire _w32105_ ;
	wire _w32104_ ;
	wire _w32103_ ;
	wire _w32102_ ;
	wire _w32101_ ;
	wire _w32100_ ;
	wire _w32099_ ;
	wire _w32098_ ;
	wire _w32097_ ;
	wire _w32096_ ;
	wire _w32095_ ;
	wire _w32094_ ;
	wire _w32093_ ;
	wire _w32092_ ;
	wire _w32091_ ;
	wire _w32090_ ;
	wire _w32089_ ;
	wire _w32088_ ;
	wire _w32087_ ;
	wire _w32086_ ;
	wire _w32085_ ;
	wire _w32084_ ;
	wire _w32083_ ;
	wire _w32082_ ;
	wire _w32081_ ;
	wire _w32080_ ;
	wire _w32079_ ;
	wire _w32078_ ;
	wire _w32077_ ;
	wire _w32076_ ;
	wire _w32075_ ;
	wire _w32074_ ;
	wire _w32073_ ;
	wire _w32072_ ;
	wire _w32071_ ;
	wire _w32070_ ;
	wire _w32069_ ;
	wire _w32068_ ;
	wire _w32067_ ;
	wire _w32066_ ;
	wire _w32065_ ;
	wire _w32064_ ;
	wire _w32063_ ;
	wire _w32062_ ;
	wire _w32061_ ;
	wire _w32060_ ;
	wire _w32059_ ;
	wire _w32058_ ;
	wire _w32057_ ;
	wire _w32056_ ;
	wire _w32055_ ;
	wire _w32054_ ;
	wire _w32053_ ;
	wire _w32052_ ;
	wire _w32051_ ;
	wire _w32050_ ;
	wire _w32049_ ;
	wire _w32048_ ;
	wire _w32047_ ;
	wire _w32046_ ;
	wire _w32045_ ;
	wire _w32044_ ;
	wire _w32043_ ;
	wire _w32042_ ;
	wire _w32041_ ;
	wire _w32040_ ;
	wire _w32039_ ;
	wire _w32038_ ;
	wire _w32037_ ;
	wire _w32036_ ;
	wire _w32035_ ;
	wire _w32034_ ;
	wire _w32033_ ;
	wire _w32032_ ;
	wire _w32031_ ;
	wire _w32030_ ;
	wire _w32029_ ;
	wire _w32028_ ;
	wire _w32027_ ;
	wire _w32026_ ;
	wire _w32025_ ;
	wire _w32024_ ;
	wire _w32023_ ;
	wire _w32022_ ;
	wire _w32021_ ;
	wire _w32020_ ;
	wire _w32019_ ;
	wire _w32018_ ;
	wire _w32017_ ;
	wire _w32016_ ;
	wire _w32015_ ;
	wire _w32014_ ;
	wire _w32013_ ;
	wire _w32012_ ;
	wire _w32011_ ;
	wire _w32010_ ;
	wire _w32009_ ;
	wire _w32008_ ;
	wire _w32007_ ;
	wire _w32006_ ;
	wire _w32005_ ;
	wire _w32004_ ;
	wire _w32003_ ;
	wire _w32002_ ;
	wire _w32001_ ;
	wire _w32000_ ;
	wire _w31999_ ;
	wire _w31998_ ;
	wire _w31997_ ;
	wire _w31996_ ;
	wire _w31995_ ;
	wire _w31994_ ;
	wire _w31993_ ;
	wire _w31992_ ;
	wire _w31991_ ;
	wire _w31990_ ;
	wire _w31989_ ;
	wire _w31988_ ;
	wire _w31987_ ;
	wire _w31986_ ;
	wire _w31985_ ;
	wire _w31984_ ;
	wire _w31983_ ;
	wire _w31982_ ;
	wire _w31981_ ;
	wire _w31980_ ;
	wire _w31979_ ;
	wire _w31978_ ;
	wire _w31977_ ;
	wire _w31976_ ;
	wire _w31975_ ;
	wire _w31974_ ;
	wire _w31973_ ;
	wire _w31972_ ;
	wire _w31971_ ;
	wire _w31970_ ;
	wire _w31969_ ;
	wire _w31968_ ;
	wire _w31967_ ;
	wire _w31966_ ;
	wire _w31965_ ;
	wire _w31964_ ;
	wire _w31963_ ;
	wire _w31962_ ;
	wire _w31961_ ;
	wire _w31960_ ;
	wire _w31959_ ;
	wire _w31958_ ;
	wire _w31957_ ;
	wire _w31956_ ;
	wire _w31955_ ;
	wire _w31954_ ;
	wire _w31953_ ;
	wire _w31952_ ;
	wire _w31951_ ;
	wire _w31950_ ;
	wire _w31949_ ;
	wire _w31948_ ;
	wire _w31947_ ;
	wire _w31946_ ;
	wire _w31945_ ;
	wire _w31944_ ;
	wire _w31943_ ;
	wire _w31942_ ;
	wire _w31941_ ;
	wire _w31940_ ;
	wire _w31939_ ;
	wire _w31938_ ;
	wire _w31937_ ;
	wire _w31936_ ;
	wire _w31935_ ;
	wire _w31934_ ;
	wire _w31933_ ;
	wire _w31932_ ;
	wire _w31931_ ;
	wire _w31930_ ;
	wire _w31929_ ;
	wire _w31928_ ;
	wire _w31927_ ;
	wire _w31926_ ;
	wire _w31925_ ;
	wire _w31924_ ;
	wire _w31923_ ;
	wire _w31922_ ;
	wire _w31921_ ;
	wire _w31920_ ;
	wire _w31919_ ;
	wire _w31918_ ;
	wire _w31917_ ;
	wire _w31916_ ;
	wire _w31915_ ;
	wire _w31914_ ;
	wire _w31913_ ;
	wire _w31912_ ;
	wire _w31911_ ;
	wire _w31910_ ;
	wire _w31909_ ;
	wire _w31908_ ;
	wire _w31907_ ;
	wire _w31906_ ;
	wire _w31905_ ;
	wire _w31904_ ;
	wire _w31903_ ;
	wire _w31902_ ;
	wire _w31901_ ;
	wire _w31900_ ;
	wire _w31899_ ;
	wire _w31898_ ;
	wire _w31897_ ;
	wire _w31896_ ;
	wire _w31895_ ;
	wire _w31894_ ;
	wire _w31893_ ;
	wire _w31892_ ;
	wire _w31891_ ;
	wire _w31890_ ;
	wire _w31889_ ;
	wire _w31888_ ;
	wire _w31887_ ;
	wire _w31886_ ;
	wire _w31885_ ;
	wire _w31884_ ;
	wire _w31883_ ;
	wire _w31882_ ;
	wire _w31881_ ;
	wire _w31880_ ;
	wire _w31879_ ;
	wire _w31878_ ;
	wire _w31877_ ;
	wire _w31876_ ;
	wire _w31875_ ;
	wire _w31874_ ;
	wire _w31873_ ;
	wire _w31872_ ;
	wire _w31871_ ;
	wire _w31870_ ;
	wire _w31869_ ;
	wire _w31868_ ;
	wire _w31867_ ;
	wire _w31866_ ;
	wire _w31865_ ;
	wire _w31864_ ;
	wire _w31863_ ;
	wire _w31862_ ;
	wire _w31861_ ;
	wire _w31860_ ;
	wire _w31859_ ;
	wire _w31858_ ;
	wire _w31857_ ;
	wire _w31856_ ;
	wire _w31855_ ;
	wire _w31854_ ;
	wire _w31853_ ;
	wire _w31852_ ;
	wire _w31851_ ;
	wire _w31850_ ;
	wire _w31849_ ;
	wire _w31848_ ;
	wire _w31847_ ;
	wire _w31846_ ;
	wire _w31845_ ;
	wire _w31844_ ;
	wire _w31843_ ;
	wire _w31842_ ;
	wire _w31841_ ;
	wire _w31840_ ;
	wire _w31839_ ;
	wire _w31838_ ;
	wire _w31837_ ;
	wire _w31836_ ;
	wire _w31835_ ;
	wire _w31834_ ;
	wire _w31833_ ;
	wire _w31832_ ;
	wire _w31831_ ;
	wire _w31830_ ;
	wire _w31829_ ;
	wire _w31828_ ;
	wire _w31827_ ;
	wire _w31826_ ;
	wire _w31825_ ;
	wire _w31824_ ;
	wire _w31823_ ;
	wire _w31822_ ;
	wire _w31821_ ;
	wire _w31820_ ;
	wire _w31819_ ;
	wire _w31818_ ;
	wire _w31817_ ;
	wire _w31816_ ;
	wire _w31815_ ;
	wire _w31814_ ;
	wire _w31813_ ;
	wire _w31812_ ;
	wire _w31811_ ;
	wire _w31810_ ;
	wire _w31809_ ;
	wire _w31808_ ;
	wire _w31807_ ;
	wire _w31806_ ;
	wire _w31805_ ;
	wire _w31804_ ;
	wire _w31803_ ;
	wire _w31802_ ;
	wire _w31801_ ;
	wire _w31800_ ;
	wire _w31799_ ;
	wire _w31798_ ;
	wire _w31797_ ;
	wire _w31796_ ;
	wire _w31795_ ;
	wire _w31794_ ;
	wire _w31793_ ;
	wire _w31792_ ;
	wire _w31791_ ;
	wire _w31790_ ;
	wire _w31789_ ;
	wire _w31788_ ;
	wire _w31787_ ;
	wire _w31786_ ;
	wire _w31785_ ;
	wire _w31784_ ;
	wire _w31783_ ;
	wire _w31782_ ;
	wire _w31781_ ;
	wire _w31780_ ;
	wire _w31779_ ;
	wire _w31778_ ;
	wire _w31777_ ;
	wire _w31776_ ;
	wire _w31775_ ;
	wire _w31774_ ;
	wire _w31773_ ;
	wire _w31772_ ;
	wire _w31771_ ;
	wire _w31770_ ;
	wire _w31769_ ;
	wire _w31768_ ;
	wire _w31767_ ;
	wire _w31766_ ;
	wire _w31765_ ;
	wire _w31764_ ;
	wire _w31763_ ;
	wire _w31762_ ;
	wire _w31761_ ;
	wire _w31760_ ;
	wire _w31759_ ;
	wire _w31758_ ;
	wire _w31757_ ;
	wire _w31756_ ;
	wire _w31755_ ;
	wire _w31754_ ;
	wire _w31753_ ;
	wire _w31752_ ;
	wire _w31751_ ;
	wire _w31750_ ;
	wire _w31749_ ;
	wire _w31748_ ;
	wire _w31747_ ;
	wire _w31746_ ;
	wire _w31745_ ;
	wire _w31744_ ;
	wire _w31743_ ;
	wire _w31742_ ;
	wire _w31741_ ;
	wire _w31740_ ;
	wire _w31739_ ;
	wire _w31738_ ;
	wire _w31737_ ;
	wire _w31736_ ;
	wire _w31735_ ;
	wire _w31734_ ;
	wire _w31733_ ;
	wire _w31732_ ;
	wire _w31731_ ;
	wire _w31730_ ;
	wire _w31729_ ;
	wire _w31728_ ;
	wire _w31727_ ;
	wire _w31726_ ;
	wire _w31725_ ;
	wire _w31724_ ;
	wire _w31723_ ;
	wire _w31722_ ;
	wire _w31721_ ;
	wire _w31720_ ;
	wire _w31719_ ;
	wire _w31718_ ;
	wire _w31717_ ;
	wire _w31716_ ;
	wire _w31715_ ;
	wire _w31714_ ;
	wire _w31713_ ;
	wire _w31712_ ;
	wire _w31711_ ;
	wire _w31710_ ;
	wire _w31709_ ;
	wire _w31708_ ;
	wire _w31707_ ;
	wire _w31706_ ;
	wire _w31705_ ;
	wire _w31704_ ;
	wire _w31703_ ;
	wire _w31702_ ;
	wire _w31701_ ;
	wire _w31700_ ;
	wire _w31699_ ;
	wire _w31698_ ;
	wire _w31697_ ;
	wire _w31696_ ;
	wire _w31695_ ;
	wire _w31694_ ;
	wire _w31693_ ;
	wire _w31692_ ;
	wire _w31691_ ;
	wire _w31690_ ;
	wire _w31689_ ;
	wire _w31688_ ;
	wire _w31687_ ;
	wire _w31686_ ;
	wire _w31685_ ;
	wire _w31684_ ;
	wire _w31683_ ;
	wire _w31682_ ;
	wire _w31681_ ;
	wire _w31680_ ;
	wire _w31679_ ;
	wire _w31678_ ;
	wire _w31677_ ;
	wire _w31676_ ;
	wire _w31675_ ;
	wire _w31674_ ;
	wire _w31673_ ;
	wire _w31672_ ;
	wire _w31671_ ;
	wire _w31670_ ;
	wire _w31669_ ;
	wire _w31668_ ;
	wire _w31667_ ;
	wire _w31666_ ;
	wire _w31665_ ;
	wire _w31664_ ;
	wire _w31663_ ;
	wire _w31662_ ;
	wire _w31661_ ;
	wire _w31660_ ;
	wire _w31659_ ;
	wire _w31658_ ;
	wire _w31657_ ;
	wire _w31656_ ;
	wire _w31655_ ;
	wire _w31654_ ;
	wire _w31653_ ;
	wire _w31652_ ;
	wire _w31651_ ;
	wire _w31650_ ;
	wire _w31649_ ;
	wire _w31648_ ;
	wire _w31647_ ;
	wire _w31646_ ;
	wire _w31645_ ;
	wire _w31644_ ;
	wire _w31643_ ;
	wire _w31642_ ;
	wire _w31641_ ;
	wire _w31640_ ;
	wire _w31639_ ;
	wire _w31638_ ;
	wire _w31637_ ;
	wire _w31636_ ;
	wire _w31635_ ;
	wire _w31634_ ;
	wire _w31633_ ;
	wire _w31632_ ;
	wire _w31631_ ;
	wire _w31630_ ;
	wire _w31629_ ;
	wire _w31628_ ;
	wire _w31627_ ;
	wire _w31626_ ;
	wire _w31625_ ;
	wire _w31624_ ;
	wire _w31623_ ;
	wire _w31622_ ;
	wire _w31621_ ;
	wire _w31620_ ;
	wire _w31619_ ;
	wire _w31618_ ;
	wire _w31617_ ;
	wire _w31616_ ;
	wire _w31615_ ;
	wire _w31614_ ;
	wire _w31613_ ;
	wire _w31612_ ;
	wire _w31611_ ;
	wire _w31610_ ;
	wire _w31609_ ;
	wire _w31608_ ;
	wire _w31607_ ;
	wire _w31606_ ;
	wire _w31605_ ;
	wire _w31604_ ;
	wire _w31603_ ;
	wire _w31602_ ;
	wire _w31601_ ;
	wire _w31600_ ;
	wire _w31599_ ;
	wire _w31598_ ;
	wire _w31597_ ;
	wire _w31596_ ;
	wire _w31595_ ;
	wire _w31594_ ;
	wire _w31593_ ;
	wire _w31592_ ;
	wire _w31591_ ;
	wire _w31590_ ;
	wire _w31589_ ;
	wire _w31588_ ;
	wire _w31587_ ;
	wire _w31586_ ;
	wire _w31585_ ;
	wire _w31584_ ;
	wire _w31583_ ;
	wire _w31582_ ;
	wire _w31581_ ;
	wire _w31580_ ;
	wire _w31579_ ;
	wire _w31578_ ;
	wire _w31577_ ;
	wire _w31576_ ;
	wire _w31575_ ;
	wire _w31574_ ;
	wire _w31573_ ;
	wire _w31572_ ;
	wire _w31571_ ;
	wire _w31570_ ;
	wire _w31569_ ;
	wire _w31568_ ;
	wire _w31567_ ;
	wire _w31566_ ;
	wire _w31565_ ;
	wire _w31564_ ;
	wire _w31563_ ;
	wire _w31562_ ;
	wire _w31561_ ;
	wire _w31560_ ;
	wire _w31559_ ;
	wire _w31558_ ;
	wire _w31557_ ;
	wire _w31556_ ;
	wire _w31555_ ;
	wire _w31554_ ;
	wire _w31553_ ;
	wire _w31552_ ;
	wire _w31551_ ;
	wire _w31550_ ;
	wire _w31549_ ;
	wire _w31548_ ;
	wire _w31547_ ;
	wire _w31546_ ;
	wire _w31545_ ;
	wire _w31544_ ;
	wire _w31543_ ;
	wire _w31542_ ;
	wire _w31541_ ;
	wire _w31540_ ;
	wire _w31539_ ;
	wire _w31538_ ;
	wire _w31537_ ;
	wire _w31536_ ;
	wire _w31535_ ;
	wire _w31534_ ;
	wire _w31533_ ;
	wire _w31532_ ;
	wire _w31531_ ;
	wire _w31530_ ;
	wire _w31529_ ;
	wire _w31528_ ;
	wire _w31527_ ;
	wire _w31526_ ;
	wire _w31525_ ;
	wire _w31524_ ;
	wire _w31523_ ;
	wire _w31522_ ;
	wire _w31521_ ;
	wire _w31520_ ;
	wire _w31519_ ;
	wire _w31518_ ;
	wire _w31517_ ;
	wire _w31516_ ;
	wire _w31515_ ;
	wire _w31514_ ;
	wire _w31513_ ;
	wire _w31512_ ;
	wire _w31511_ ;
	wire _w31510_ ;
	wire _w31509_ ;
	wire _w31508_ ;
	wire _w31507_ ;
	wire _w31506_ ;
	wire _w31505_ ;
	wire _w31504_ ;
	wire _w31503_ ;
	wire _w31502_ ;
	wire _w31501_ ;
	wire _w31500_ ;
	wire _w31499_ ;
	wire _w31498_ ;
	wire _w31497_ ;
	wire _w31496_ ;
	wire _w31495_ ;
	wire _w31494_ ;
	wire _w31493_ ;
	wire _w31492_ ;
	wire _w31491_ ;
	wire _w31490_ ;
	wire _w31489_ ;
	wire _w31488_ ;
	wire _w31487_ ;
	wire _w31486_ ;
	wire _w31485_ ;
	wire _w31484_ ;
	wire _w31483_ ;
	wire _w31482_ ;
	wire _w31481_ ;
	wire _w31480_ ;
	wire _w31479_ ;
	wire _w31478_ ;
	wire _w31477_ ;
	wire _w31476_ ;
	wire _w31475_ ;
	wire _w31474_ ;
	wire _w31473_ ;
	wire _w31472_ ;
	wire _w31471_ ;
	wire _w31470_ ;
	wire _w31469_ ;
	wire _w31468_ ;
	wire _w31467_ ;
	wire _w31466_ ;
	wire _w31465_ ;
	wire _w31464_ ;
	wire _w31463_ ;
	wire _w31462_ ;
	wire _w31461_ ;
	wire _w31460_ ;
	wire _w31459_ ;
	wire _w31458_ ;
	wire _w31457_ ;
	wire _w31456_ ;
	wire _w31455_ ;
	wire _w31454_ ;
	wire _w31453_ ;
	wire _w31452_ ;
	wire _w31451_ ;
	wire _w31450_ ;
	wire _w31449_ ;
	wire _w31448_ ;
	wire _w31447_ ;
	wire _w31446_ ;
	wire _w31445_ ;
	wire _w31444_ ;
	wire _w31443_ ;
	wire _w31442_ ;
	wire _w31441_ ;
	wire _w31440_ ;
	wire _w31439_ ;
	wire _w31438_ ;
	wire _w31437_ ;
	wire _w31436_ ;
	wire _w31435_ ;
	wire _w31434_ ;
	wire _w31433_ ;
	wire _w31432_ ;
	wire _w31431_ ;
	wire _w31430_ ;
	wire _w31429_ ;
	wire _w31428_ ;
	wire _w31427_ ;
	wire _w31426_ ;
	wire _w31425_ ;
	wire _w31424_ ;
	wire _w31423_ ;
	wire _w31422_ ;
	wire _w31421_ ;
	wire _w31420_ ;
	wire _w31419_ ;
	wire _w31418_ ;
	wire _w31417_ ;
	wire _w31416_ ;
	wire _w31415_ ;
	wire _w31414_ ;
	wire _w31413_ ;
	wire _w31412_ ;
	wire _w31411_ ;
	wire _w31410_ ;
	wire _w31409_ ;
	wire _w31408_ ;
	wire _w31407_ ;
	wire _w31406_ ;
	wire _w31405_ ;
	wire _w31404_ ;
	wire _w31403_ ;
	wire _w31402_ ;
	wire _w31401_ ;
	wire _w31400_ ;
	wire _w31399_ ;
	wire _w31398_ ;
	wire _w31397_ ;
	wire _w31396_ ;
	wire _w31395_ ;
	wire _w31394_ ;
	wire _w31393_ ;
	wire _w31392_ ;
	wire _w31391_ ;
	wire _w31390_ ;
	wire _w31389_ ;
	wire _w31388_ ;
	wire _w31387_ ;
	wire _w31386_ ;
	wire _w31385_ ;
	wire _w31384_ ;
	wire _w31383_ ;
	wire _w31382_ ;
	wire _w31381_ ;
	wire _w31380_ ;
	wire _w31379_ ;
	wire _w31378_ ;
	wire _w31377_ ;
	wire _w31376_ ;
	wire _w31375_ ;
	wire _w31374_ ;
	wire _w31373_ ;
	wire _w31372_ ;
	wire _w31371_ ;
	wire _w31370_ ;
	wire _w31369_ ;
	wire _w31368_ ;
	wire _w31367_ ;
	wire _w31366_ ;
	wire _w31365_ ;
	wire _w31364_ ;
	wire _w31363_ ;
	wire _w31362_ ;
	wire _w31361_ ;
	wire _w31360_ ;
	wire _w31359_ ;
	wire _w31358_ ;
	wire _w31357_ ;
	wire _w31356_ ;
	wire _w31355_ ;
	wire _w31354_ ;
	wire _w31353_ ;
	wire _w31352_ ;
	wire _w31351_ ;
	wire _w31350_ ;
	wire _w31349_ ;
	wire _w31348_ ;
	wire _w31347_ ;
	wire _w31346_ ;
	wire _w31345_ ;
	wire _w31344_ ;
	wire _w31343_ ;
	wire _w31342_ ;
	wire _w31341_ ;
	wire _w31340_ ;
	wire _w31339_ ;
	wire _w31338_ ;
	wire _w31337_ ;
	wire _w31336_ ;
	wire _w31335_ ;
	wire _w31334_ ;
	wire _w31333_ ;
	wire _w31332_ ;
	wire _w31331_ ;
	wire _w31330_ ;
	wire _w31329_ ;
	wire _w31328_ ;
	wire _w31327_ ;
	wire _w31326_ ;
	wire _w31325_ ;
	wire _w31324_ ;
	wire _w31323_ ;
	wire _w31322_ ;
	wire _w31321_ ;
	wire _w31320_ ;
	wire _w31319_ ;
	wire _w31318_ ;
	wire _w31317_ ;
	wire _w31316_ ;
	wire _w31315_ ;
	wire _w31314_ ;
	wire _w31313_ ;
	wire _w31312_ ;
	wire _w31311_ ;
	wire _w31310_ ;
	wire _w31309_ ;
	wire _w31308_ ;
	wire _w31307_ ;
	wire _w31306_ ;
	wire _w31305_ ;
	wire _w31304_ ;
	wire _w31303_ ;
	wire _w31302_ ;
	wire _w31301_ ;
	wire _w31300_ ;
	wire _w31299_ ;
	wire _w31298_ ;
	wire _w31297_ ;
	wire _w31296_ ;
	wire _w31295_ ;
	wire _w31294_ ;
	wire _w31293_ ;
	wire _w31292_ ;
	wire _w31291_ ;
	wire _w31290_ ;
	wire _w31289_ ;
	wire _w31288_ ;
	wire _w31287_ ;
	wire _w31286_ ;
	wire _w31285_ ;
	wire _w31284_ ;
	wire _w31283_ ;
	wire _w31282_ ;
	wire _w31281_ ;
	wire _w31280_ ;
	wire _w31279_ ;
	wire _w31278_ ;
	wire _w31277_ ;
	wire _w31276_ ;
	wire _w31275_ ;
	wire _w31274_ ;
	wire _w31273_ ;
	wire _w31272_ ;
	wire _w31271_ ;
	wire _w31270_ ;
	wire _w31269_ ;
	wire _w31268_ ;
	wire _w31267_ ;
	wire _w31266_ ;
	wire _w31265_ ;
	wire _w31264_ ;
	wire _w31263_ ;
	wire _w31262_ ;
	wire _w31261_ ;
	wire _w31260_ ;
	wire _w31259_ ;
	wire _w31258_ ;
	wire _w31257_ ;
	wire _w31256_ ;
	wire _w31255_ ;
	wire _w31254_ ;
	wire _w31253_ ;
	wire _w31252_ ;
	wire _w31251_ ;
	wire _w31250_ ;
	wire _w31249_ ;
	wire _w31248_ ;
	wire _w31247_ ;
	wire _w31246_ ;
	wire _w31245_ ;
	wire _w31244_ ;
	wire _w31243_ ;
	wire _w31242_ ;
	wire _w31241_ ;
	wire _w31240_ ;
	wire _w31239_ ;
	wire _w31238_ ;
	wire _w31237_ ;
	wire _w31236_ ;
	wire _w31235_ ;
	wire _w31234_ ;
	wire _w31233_ ;
	wire _w31232_ ;
	wire _w31231_ ;
	wire _w31230_ ;
	wire _w31229_ ;
	wire _w31228_ ;
	wire _w31227_ ;
	wire _w31226_ ;
	wire _w31225_ ;
	wire _w31224_ ;
	wire _w31223_ ;
	wire _w31222_ ;
	wire _w31221_ ;
	wire _w31220_ ;
	wire _w31219_ ;
	wire _w31218_ ;
	wire _w31217_ ;
	wire _w31216_ ;
	wire _w31215_ ;
	wire _w31214_ ;
	wire _w31213_ ;
	wire _w31212_ ;
	wire _w31211_ ;
	wire _w31210_ ;
	wire _w31209_ ;
	wire _w31208_ ;
	wire _w31207_ ;
	wire _w31206_ ;
	wire _w31205_ ;
	wire _w31204_ ;
	wire _w31203_ ;
	wire _w31202_ ;
	wire _w31201_ ;
	wire _w31200_ ;
	wire _w31199_ ;
	wire _w31198_ ;
	wire _w31197_ ;
	wire _w31196_ ;
	wire _w31195_ ;
	wire _w31194_ ;
	wire _w31193_ ;
	wire _w31192_ ;
	wire _w31191_ ;
	wire _w31190_ ;
	wire _w31189_ ;
	wire _w31188_ ;
	wire _w31187_ ;
	wire _w31186_ ;
	wire _w31185_ ;
	wire _w31184_ ;
	wire _w31183_ ;
	wire _w31182_ ;
	wire _w31181_ ;
	wire _w31180_ ;
	wire _w31179_ ;
	wire _w31178_ ;
	wire _w31177_ ;
	wire _w31176_ ;
	wire _w31175_ ;
	wire _w31174_ ;
	wire _w31173_ ;
	wire _w31172_ ;
	wire _w31171_ ;
	wire _w31170_ ;
	wire _w31169_ ;
	wire _w31168_ ;
	wire _w31167_ ;
	wire _w31166_ ;
	wire _w31165_ ;
	wire _w31164_ ;
	wire _w31163_ ;
	wire _w31162_ ;
	wire _w31161_ ;
	wire _w31160_ ;
	wire _w31159_ ;
	wire _w31158_ ;
	wire _w31157_ ;
	wire _w31156_ ;
	wire _w31155_ ;
	wire _w31154_ ;
	wire _w31153_ ;
	wire _w31152_ ;
	wire _w31151_ ;
	wire _w31150_ ;
	wire _w31149_ ;
	wire _w31148_ ;
	wire _w31147_ ;
	wire _w31146_ ;
	wire _w31145_ ;
	wire _w31144_ ;
	wire _w31143_ ;
	wire _w31142_ ;
	wire _w31141_ ;
	wire _w31140_ ;
	wire _w31139_ ;
	wire _w31138_ ;
	wire _w31137_ ;
	wire _w31136_ ;
	wire _w31135_ ;
	wire _w31134_ ;
	wire _w31133_ ;
	wire _w31132_ ;
	wire _w31131_ ;
	wire _w31130_ ;
	wire _w31129_ ;
	wire _w31128_ ;
	wire _w31127_ ;
	wire _w31126_ ;
	wire _w31125_ ;
	wire _w31124_ ;
	wire _w31123_ ;
	wire _w31122_ ;
	wire _w31121_ ;
	wire _w31120_ ;
	wire _w31119_ ;
	wire _w31118_ ;
	wire _w31117_ ;
	wire _w31116_ ;
	wire _w31115_ ;
	wire _w31114_ ;
	wire _w31113_ ;
	wire _w31112_ ;
	wire _w31111_ ;
	wire _w31110_ ;
	wire _w31109_ ;
	wire _w31108_ ;
	wire _w31107_ ;
	wire _w31106_ ;
	wire _w31105_ ;
	wire _w31104_ ;
	wire _w31103_ ;
	wire _w31102_ ;
	wire _w31101_ ;
	wire _w31100_ ;
	wire _w31099_ ;
	wire _w31098_ ;
	wire _w31097_ ;
	wire _w31096_ ;
	wire _w31095_ ;
	wire _w31094_ ;
	wire _w31093_ ;
	wire _w31092_ ;
	wire _w31091_ ;
	wire _w31090_ ;
	wire _w31089_ ;
	wire _w31088_ ;
	wire _w31087_ ;
	wire _w31086_ ;
	wire _w31085_ ;
	wire _w31084_ ;
	wire _w31083_ ;
	wire _w31082_ ;
	wire _w31081_ ;
	wire _w31080_ ;
	wire _w31079_ ;
	wire _w31078_ ;
	wire _w31077_ ;
	wire _w31076_ ;
	wire _w31075_ ;
	wire _w31074_ ;
	wire _w31073_ ;
	wire _w31072_ ;
	wire _w31071_ ;
	wire _w31070_ ;
	wire _w31069_ ;
	wire _w31068_ ;
	wire _w31067_ ;
	wire _w31066_ ;
	wire _w31065_ ;
	wire _w31064_ ;
	wire _w31063_ ;
	wire _w31062_ ;
	wire _w31061_ ;
	wire _w31060_ ;
	wire _w31059_ ;
	wire _w31058_ ;
	wire _w31057_ ;
	wire _w31056_ ;
	wire _w31055_ ;
	wire _w31054_ ;
	wire _w31053_ ;
	wire _w31052_ ;
	wire _w31051_ ;
	wire _w31050_ ;
	wire _w31049_ ;
	wire _w31048_ ;
	wire _w31047_ ;
	wire _w31046_ ;
	wire _w31045_ ;
	wire _w31044_ ;
	wire _w31043_ ;
	wire _w31042_ ;
	wire _w31041_ ;
	wire _w31040_ ;
	wire _w31039_ ;
	wire _w31038_ ;
	wire _w31037_ ;
	wire _w31036_ ;
	wire _w31035_ ;
	wire _w31034_ ;
	wire _w31033_ ;
	wire _w31032_ ;
	wire _w31031_ ;
	wire _w31030_ ;
	wire _w31029_ ;
	wire _w31028_ ;
	wire _w31027_ ;
	wire _w31026_ ;
	wire _w31025_ ;
	wire _w31024_ ;
	wire _w31023_ ;
	wire _w31022_ ;
	wire _w31021_ ;
	wire _w31020_ ;
	wire _w31019_ ;
	wire _w31018_ ;
	wire _w31017_ ;
	wire _w31016_ ;
	wire _w31015_ ;
	wire _w31014_ ;
	wire _w31013_ ;
	wire _w31012_ ;
	wire _w31011_ ;
	wire _w31010_ ;
	wire _w31009_ ;
	wire _w31008_ ;
	wire _w31007_ ;
	wire _w31006_ ;
	wire _w31005_ ;
	wire _w31004_ ;
	wire _w31003_ ;
	wire _w31002_ ;
	wire _w31001_ ;
	wire _w31000_ ;
	wire _w30999_ ;
	wire _w30998_ ;
	wire _w30997_ ;
	wire _w30996_ ;
	wire _w30995_ ;
	wire _w30994_ ;
	wire _w30993_ ;
	wire _w30992_ ;
	wire _w30991_ ;
	wire _w30990_ ;
	wire _w30989_ ;
	wire _w30988_ ;
	wire _w30987_ ;
	wire _w30986_ ;
	wire _w30985_ ;
	wire _w30984_ ;
	wire _w30983_ ;
	wire _w30982_ ;
	wire _w30981_ ;
	wire _w30980_ ;
	wire _w30979_ ;
	wire _w30978_ ;
	wire _w30977_ ;
	wire _w30976_ ;
	wire _w30975_ ;
	wire _w30974_ ;
	wire _w30973_ ;
	wire _w30972_ ;
	wire _w30971_ ;
	wire _w30970_ ;
	wire _w30969_ ;
	wire _w30968_ ;
	wire _w30967_ ;
	wire _w30966_ ;
	wire _w30965_ ;
	wire _w30964_ ;
	wire _w30963_ ;
	wire _w30962_ ;
	wire _w30961_ ;
	wire _w30960_ ;
	wire _w30959_ ;
	wire _w30958_ ;
	wire _w30957_ ;
	wire _w30956_ ;
	wire _w30955_ ;
	wire _w30954_ ;
	wire _w30953_ ;
	wire _w30952_ ;
	wire _w30951_ ;
	wire _w30950_ ;
	wire _w30949_ ;
	wire _w30948_ ;
	wire _w30947_ ;
	wire _w30946_ ;
	wire _w30945_ ;
	wire _w30944_ ;
	wire _w30943_ ;
	wire _w30942_ ;
	wire _w30941_ ;
	wire _w30940_ ;
	wire _w30939_ ;
	wire _w30938_ ;
	wire _w30937_ ;
	wire _w30936_ ;
	wire _w30935_ ;
	wire _w30934_ ;
	wire _w30933_ ;
	wire _w30932_ ;
	wire _w30931_ ;
	wire _w30930_ ;
	wire _w30929_ ;
	wire _w30928_ ;
	wire _w30927_ ;
	wire _w30926_ ;
	wire _w30925_ ;
	wire _w30924_ ;
	wire _w30923_ ;
	wire _w30922_ ;
	wire _w30921_ ;
	wire _w30920_ ;
	wire _w30919_ ;
	wire _w30918_ ;
	wire _w30917_ ;
	wire _w30916_ ;
	wire _w30915_ ;
	wire _w30914_ ;
	wire _w30913_ ;
	wire _w30912_ ;
	wire _w30911_ ;
	wire _w30910_ ;
	wire _w30909_ ;
	wire _w30908_ ;
	wire _w30907_ ;
	wire _w30906_ ;
	wire _w30905_ ;
	wire _w30904_ ;
	wire _w30903_ ;
	wire _w30902_ ;
	wire _w30901_ ;
	wire _w30900_ ;
	wire _w30899_ ;
	wire _w30898_ ;
	wire _w30897_ ;
	wire _w30896_ ;
	wire _w30895_ ;
	wire _w30894_ ;
	wire _w30893_ ;
	wire _w30892_ ;
	wire _w30891_ ;
	wire _w30890_ ;
	wire _w30889_ ;
	wire _w30888_ ;
	wire _w30887_ ;
	wire _w30886_ ;
	wire _w30885_ ;
	wire _w30884_ ;
	wire _w30883_ ;
	wire _w30882_ ;
	wire _w30881_ ;
	wire _w30880_ ;
	wire _w30879_ ;
	wire _w30878_ ;
	wire _w30877_ ;
	wire _w30876_ ;
	wire _w30875_ ;
	wire _w30874_ ;
	wire _w30873_ ;
	wire _w30872_ ;
	wire _w30871_ ;
	wire _w30870_ ;
	wire _w30869_ ;
	wire _w30868_ ;
	wire _w30867_ ;
	wire _w30866_ ;
	wire _w30865_ ;
	wire _w30864_ ;
	wire _w30863_ ;
	wire _w30862_ ;
	wire _w30861_ ;
	wire _w30860_ ;
	wire _w30859_ ;
	wire _w30858_ ;
	wire _w30857_ ;
	wire _w30856_ ;
	wire _w30855_ ;
	wire _w30854_ ;
	wire _w30853_ ;
	wire _w30852_ ;
	wire _w30851_ ;
	wire _w30850_ ;
	wire _w30849_ ;
	wire _w30848_ ;
	wire _w30847_ ;
	wire _w30846_ ;
	wire _w30845_ ;
	wire _w30844_ ;
	wire _w30843_ ;
	wire _w30842_ ;
	wire _w30841_ ;
	wire _w30840_ ;
	wire _w30839_ ;
	wire _w30838_ ;
	wire _w30837_ ;
	wire _w30836_ ;
	wire _w30835_ ;
	wire _w30834_ ;
	wire _w30833_ ;
	wire _w30832_ ;
	wire _w30831_ ;
	wire _w30830_ ;
	wire _w30829_ ;
	wire _w30828_ ;
	wire _w30827_ ;
	wire _w30826_ ;
	wire _w30825_ ;
	wire _w30824_ ;
	wire _w30823_ ;
	wire _w30822_ ;
	wire _w30821_ ;
	wire _w30820_ ;
	wire _w30819_ ;
	wire _w30818_ ;
	wire _w30817_ ;
	wire _w30816_ ;
	wire _w30815_ ;
	wire _w30814_ ;
	wire _w30813_ ;
	wire _w30812_ ;
	wire _w30811_ ;
	wire _w30810_ ;
	wire _w30809_ ;
	wire _w30808_ ;
	wire _w30807_ ;
	wire _w30806_ ;
	wire _w30805_ ;
	wire _w30804_ ;
	wire _w30803_ ;
	wire _w30802_ ;
	wire _w30801_ ;
	wire _w30800_ ;
	wire _w30799_ ;
	wire _w30798_ ;
	wire _w30797_ ;
	wire _w30796_ ;
	wire _w30795_ ;
	wire _w30794_ ;
	wire _w30793_ ;
	wire _w30792_ ;
	wire _w30791_ ;
	wire _w30790_ ;
	wire _w30789_ ;
	wire _w30788_ ;
	wire _w30787_ ;
	wire _w30786_ ;
	wire _w30785_ ;
	wire _w30784_ ;
	wire _w30783_ ;
	wire _w30782_ ;
	wire _w30781_ ;
	wire _w30780_ ;
	wire _w30779_ ;
	wire _w30778_ ;
	wire _w30777_ ;
	wire _w30776_ ;
	wire _w30775_ ;
	wire _w30774_ ;
	wire _w30773_ ;
	wire _w30772_ ;
	wire _w30771_ ;
	wire _w30770_ ;
	wire _w30769_ ;
	wire _w30768_ ;
	wire _w30767_ ;
	wire _w30766_ ;
	wire _w30765_ ;
	wire _w30764_ ;
	wire _w30763_ ;
	wire _w30762_ ;
	wire _w30761_ ;
	wire _w30760_ ;
	wire _w30759_ ;
	wire _w30758_ ;
	wire _w30757_ ;
	wire _w30756_ ;
	wire _w30755_ ;
	wire _w30754_ ;
	wire _w30753_ ;
	wire _w30752_ ;
	wire _w30751_ ;
	wire _w30750_ ;
	wire _w30749_ ;
	wire _w30748_ ;
	wire _w30747_ ;
	wire _w30746_ ;
	wire _w30745_ ;
	wire _w30744_ ;
	wire _w30743_ ;
	wire _w30742_ ;
	wire _w30741_ ;
	wire _w30740_ ;
	wire _w30739_ ;
	wire _w30738_ ;
	wire _w30737_ ;
	wire _w30736_ ;
	wire _w30735_ ;
	wire _w30734_ ;
	wire _w30733_ ;
	wire _w30732_ ;
	wire _w30731_ ;
	wire _w30730_ ;
	wire _w30729_ ;
	wire _w30728_ ;
	wire _w30727_ ;
	wire _w30726_ ;
	wire _w30725_ ;
	wire _w30724_ ;
	wire _w30723_ ;
	wire _w30722_ ;
	wire _w30721_ ;
	wire _w30720_ ;
	wire _w30719_ ;
	wire _w30718_ ;
	wire _w30717_ ;
	wire _w30716_ ;
	wire _w30715_ ;
	wire _w30714_ ;
	wire _w30713_ ;
	wire _w30712_ ;
	wire _w30711_ ;
	wire _w30710_ ;
	wire _w30709_ ;
	wire _w30708_ ;
	wire _w30707_ ;
	wire _w30706_ ;
	wire _w30705_ ;
	wire _w30704_ ;
	wire _w30703_ ;
	wire _w30702_ ;
	wire _w30701_ ;
	wire _w30700_ ;
	wire _w30699_ ;
	wire _w30698_ ;
	wire _w30697_ ;
	wire _w30696_ ;
	wire _w30695_ ;
	wire _w30694_ ;
	wire _w30693_ ;
	wire _w30692_ ;
	wire _w30691_ ;
	wire _w30690_ ;
	wire _w30689_ ;
	wire _w30688_ ;
	wire _w30687_ ;
	wire _w30686_ ;
	wire _w30685_ ;
	wire _w30684_ ;
	wire _w30683_ ;
	wire _w30682_ ;
	wire _w30681_ ;
	wire _w30680_ ;
	wire _w30679_ ;
	wire _w30678_ ;
	wire _w30677_ ;
	wire _w30676_ ;
	wire _w30675_ ;
	wire _w30674_ ;
	wire _w30673_ ;
	wire _w30672_ ;
	wire _w30671_ ;
	wire _w30670_ ;
	wire _w30669_ ;
	wire _w30668_ ;
	wire _w30667_ ;
	wire _w30666_ ;
	wire _w30665_ ;
	wire _w30664_ ;
	wire _w30663_ ;
	wire _w30662_ ;
	wire _w30661_ ;
	wire _w30660_ ;
	wire _w30659_ ;
	wire _w30658_ ;
	wire _w30657_ ;
	wire _w30656_ ;
	wire _w30655_ ;
	wire _w30654_ ;
	wire _w30653_ ;
	wire _w30652_ ;
	wire _w30651_ ;
	wire _w30650_ ;
	wire _w30649_ ;
	wire _w30648_ ;
	wire _w30647_ ;
	wire _w30646_ ;
	wire _w30645_ ;
	wire _w30644_ ;
	wire _w30643_ ;
	wire _w30642_ ;
	wire _w30641_ ;
	wire _w30640_ ;
	wire _w30639_ ;
	wire _w30638_ ;
	wire _w30637_ ;
	wire _w30636_ ;
	wire _w30635_ ;
	wire _w30634_ ;
	wire _w30633_ ;
	wire _w30632_ ;
	wire _w30631_ ;
	wire _w30630_ ;
	wire _w30629_ ;
	wire _w30628_ ;
	wire _w30627_ ;
	wire _w30626_ ;
	wire _w30625_ ;
	wire _w30624_ ;
	wire _w30623_ ;
	wire _w30622_ ;
	wire _w30621_ ;
	wire _w30620_ ;
	wire _w30619_ ;
	wire _w30618_ ;
	wire _w30617_ ;
	wire _w30616_ ;
	wire _w30615_ ;
	wire _w30614_ ;
	wire _w30613_ ;
	wire _w30612_ ;
	wire _w30611_ ;
	wire _w30610_ ;
	wire _w30609_ ;
	wire _w30608_ ;
	wire _w30607_ ;
	wire _w30606_ ;
	wire _w30605_ ;
	wire _w30604_ ;
	wire _w30603_ ;
	wire _w30602_ ;
	wire _w30601_ ;
	wire _w30600_ ;
	wire _w30599_ ;
	wire _w30598_ ;
	wire _w30597_ ;
	wire _w30596_ ;
	wire _w30595_ ;
	wire _w30594_ ;
	wire _w30593_ ;
	wire _w30592_ ;
	wire _w30591_ ;
	wire _w30590_ ;
	wire _w30589_ ;
	wire _w30588_ ;
	wire _w30587_ ;
	wire _w30586_ ;
	wire _w30585_ ;
	wire _w30584_ ;
	wire _w30583_ ;
	wire _w30582_ ;
	wire _w30581_ ;
	wire _w30580_ ;
	wire _w30579_ ;
	wire _w30578_ ;
	wire _w30577_ ;
	wire _w30576_ ;
	wire _w30575_ ;
	wire _w30574_ ;
	wire _w30573_ ;
	wire _w30572_ ;
	wire _w30571_ ;
	wire _w30570_ ;
	wire _w30569_ ;
	wire _w30568_ ;
	wire _w30567_ ;
	wire _w30566_ ;
	wire _w30565_ ;
	wire _w30564_ ;
	wire _w30563_ ;
	wire _w30562_ ;
	wire _w30561_ ;
	wire _w30560_ ;
	wire _w30559_ ;
	wire _w30558_ ;
	wire _w30557_ ;
	wire _w30556_ ;
	wire _w30555_ ;
	wire _w30554_ ;
	wire _w30553_ ;
	wire _w30552_ ;
	wire _w30551_ ;
	wire _w30550_ ;
	wire _w30549_ ;
	wire _w30548_ ;
	wire _w30547_ ;
	wire _w30546_ ;
	wire _w30545_ ;
	wire _w30544_ ;
	wire _w30543_ ;
	wire _w30542_ ;
	wire _w30541_ ;
	wire _w30540_ ;
	wire _w30539_ ;
	wire _w30538_ ;
	wire _w30537_ ;
	wire _w30536_ ;
	wire _w30535_ ;
	wire _w30534_ ;
	wire _w30533_ ;
	wire _w30532_ ;
	wire _w30531_ ;
	wire _w30530_ ;
	wire _w30529_ ;
	wire _w30528_ ;
	wire _w30527_ ;
	wire _w30526_ ;
	wire _w30525_ ;
	wire _w30524_ ;
	wire _w30523_ ;
	wire _w30522_ ;
	wire _w30521_ ;
	wire _w30520_ ;
	wire _w30519_ ;
	wire _w30518_ ;
	wire _w30517_ ;
	wire _w30516_ ;
	wire _w30515_ ;
	wire _w30514_ ;
	wire _w30513_ ;
	wire _w30512_ ;
	wire _w30511_ ;
	wire _w30510_ ;
	wire _w30509_ ;
	wire _w30508_ ;
	wire _w30507_ ;
	wire _w30506_ ;
	wire _w30505_ ;
	wire _w30504_ ;
	wire _w30503_ ;
	wire _w30502_ ;
	wire _w30501_ ;
	wire _w30500_ ;
	wire _w30499_ ;
	wire _w30498_ ;
	wire _w30497_ ;
	wire _w30496_ ;
	wire _w30495_ ;
	wire _w30494_ ;
	wire _w30493_ ;
	wire _w30492_ ;
	wire _w30491_ ;
	wire _w30490_ ;
	wire _w30489_ ;
	wire _w30488_ ;
	wire _w30487_ ;
	wire _w30486_ ;
	wire _w30485_ ;
	wire _w30484_ ;
	wire _w30483_ ;
	wire _w30482_ ;
	wire _w30481_ ;
	wire _w30480_ ;
	wire _w30479_ ;
	wire _w30478_ ;
	wire _w30477_ ;
	wire _w30476_ ;
	wire _w30475_ ;
	wire _w30474_ ;
	wire _w30473_ ;
	wire _w30472_ ;
	wire _w30471_ ;
	wire _w30470_ ;
	wire _w30469_ ;
	wire _w30468_ ;
	wire _w30467_ ;
	wire _w30466_ ;
	wire _w30465_ ;
	wire _w30464_ ;
	wire _w30463_ ;
	wire _w30462_ ;
	wire _w30461_ ;
	wire _w30460_ ;
	wire _w30459_ ;
	wire _w30458_ ;
	wire _w30457_ ;
	wire _w30456_ ;
	wire _w30455_ ;
	wire _w30454_ ;
	wire _w30453_ ;
	wire _w30452_ ;
	wire _w30451_ ;
	wire _w30450_ ;
	wire _w30449_ ;
	wire _w30448_ ;
	wire _w30447_ ;
	wire _w30446_ ;
	wire _w30445_ ;
	wire _w30444_ ;
	wire _w30443_ ;
	wire _w30442_ ;
	wire _w30441_ ;
	wire _w30440_ ;
	wire _w30439_ ;
	wire _w30438_ ;
	wire _w30437_ ;
	wire _w30436_ ;
	wire _w30435_ ;
	wire _w30434_ ;
	wire _w30433_ ;
	wire _w30432_ ;
	wire _w30431_ ;
	wire _w30430_ ;
	wire _w30429_ ;
	wire _w30428_ ;
	wire _w30427_ ;
	wire _w30426_ ;
	wire _w30425_ ;
	wire _w30424_ ;
	wire _w30423_ ;
	wire _w30422_ ;
	wire _w30421_ ;
	wire _w30420_ ;
	wire _w30419_ ;
	wire _w30418_ ;
	wire _w30417_ ;
	wire _w30416_ ;
	wire _w30415_ ;
	wire _w30414_ ;
	wire _w30413_ ;
	wire _w30412_ ;
	wire _w30411_ ;
	wire _w30410_ ;
	wire _w30409_ ;
	wire _w30408_ ;
	wire _w30407_ ;
	wire _w30406_ ;
	wire _w30405_ ;
	wire _w30404_ ;
	wire _w30403_ ;
	wire _w30402_ ;
	wire _w30401_ ;
	wire _w30400_ ;
	wire _w30399_ ;
	wire _w30398_ ;
	wire _w30397_ ;
	wire _w30396_ ;
	wire _w30395_ ;
	wire _w30394_ ;
	wire _w30393_ ;
	wire _w30392_ ;
	wire _w30391_ ;
	wire _w30390_ ;
	wire _w30389_ ;
	wire _w30388_ ;
	wire _w30387_ ;
	wire _w30386_ ;
	wire _w30385_ ;
	wire _w30384_ ;
	wire _w30383_ ;
	wire _w30382_ ;
	wire _w30381_ ;
	wire _w30380_ ;
	wire _w30379_ ;
	wire _w30378_ ;
	wire _w30377_ ;
	wire _w30376_ ;
	wire _w30375_ ;
	wire _w30374_ ;
	wire _w30373_ ;
	wire _w30372_ ;
	wire _w30371_ ;
	wire _w30370_ ;
	wire _w30369_ ;
	wire _w30368_ ;
	wire _w30367_ ;
	wire _w30366_ ;
	wire _w30365_ ;
	wire _w30364_ ;
	wire _w30363_ ;
	wire _w30362_ ;
	wire _w30361_ ;
	wire _w30360_ ;
	wire _w30359_ ;
	wire _w30358_ ;
	wire _w30357_ ;
	wire _w30356_ ;
	wire _w30355_ ;
	wire _w30354_ ;
	wire _w30353_ ;
	wire _w30352_ ;
	wire _w30351_ ;
	wire _w30350_ ;
	wire _w30349_ ;
	wire _w30348_ ;
	wire _w30347_ ;
	wire _w30346_ ;
	wire _w30345_ ;
	wire _w30344_ ;
	wire _w30343_ ;
	wire _w30342_ ;
	wire _w30341_ ;
	wire _w30340_ ;
	wire _w30339_ ;
	wire _w30338_ ;
	wire _w30337_ ;
	wire _w30336_ ;
	wire _w30335_ ;
	wire _w30334_ ;
	wire _w30333_ ;
	wire _w30332_ ;
	wire _w30331_ ;
	wire _w30330_ ;
	wire _w30329_ ;
	wire _w30328_ ;
	wire _w30327_ ;
	wire _w30326_ ;
	wire _w30325_ ;
	wire _w30324_ ;
	wire _w30323_ ;
	wire _w30322_ ;
	wire _w30321_ ;
	wire _w30320_ ;
	wire _w30319_ ;
	wire _w30318_ ;
	wire _w30317_ ;
	wire _w30316_ ;
	wire _w30315_ ;
	wire _w30314_ ;
	wire _w30313_ ;
	wire _w30312_ ;
	wire _w30311_ ;
	wire _w30310_ ;
	wire _w30309_ ;
	wire _w30308_ ;
	wire _w30307_ ;
	wire _w30306_ ;
	wire _w30305_ ;
	wire _w30304_ ;
	wire _w30303_ ;
	wire _w30302_ ;
	wire _w30301_ ;
	wire _w30300_ ;
	wire _w30299_ ;
	wire _w30298_ ;
	wire _w30297_ ;
	wire _w30296_ ;
	wire _w30295_ ;
	wire _w30294_ ;
	wire _w30293_ ;
	wire _w30292_ ;
	wire _w30291_ ;
	wire _w30290_ ;
	wire _w30289_ ;
	wire _w30288_ ;
	wire _w30287_ ;
	wire _w30286_ ;
	wire _w30285_ ;
	wire _w30284_ ;
	wire _w30283_ ;
	wire _w30282_ ;
	wire _w30281_ ;
	wire _w30280_ ;
	wire _w30279_ ;
	wire _w30278_ ;
	wire _w30277_ ;
	wire _w30276_ ;
	wire _w30275_ ;
	wire _w30274_ ;
	wire _w30273_ ;
	wire _w30272_ ;
	wire _w30271_ ;
	wire _w30270_ ;
	wire _w30269_ ;
	wire _w30268_ ;
	wire _w30267_ ;
	wire _w30266_ ;
	wire _w30265_ ;
	wire _w30264_ ;
	wire _w30263_ ;
	wire _w30262_ ;
	wire _w30261_ ;
	wire _w30260_ ;
	wire _w30259_ ;
	wire _w30258_ ;
	wire _w30257_ ;
	wire _w30256_ ;
	wire _w30255_ ;
	wire _w30254_ ;
	wire _w30253_ ;
	wire _w30252_ ;
	wire _w30251_ ;
	wire _w30250_ ;
	wire _w30249_ ;
	wire _w30248_ ;
	wire _w30247_ ;
	wire _w30246_ ;
	wire _w30245_ ;
	wire _w30244_ ;
	wire _w30243_ ;
	wire _w30242_ ;
	wire _w30241_ ;
	wire _w30240_ ;
	wire _w30239_ ;
	wire _w30238_ ;
	wire _w30237_ ;
	wire _w30236_ ;
	wire _w30235_ ;
	wire _w30234_ ;
	wire _w30233_ ;
	wire _w30232_ ;
	wire _w30231_ ;
	wire _w30230_ ;
	wire _w30229_ ;
	wire _w30228_ ;
	wire _w30227_ ;
	wire _w30226_ ;
	wire _w30225_ ;
	wire _w30224_ ;
	wire _w30223_ ;
	wire _w30222_ ;
	wire _w30221_ ;
	wire _w30220_ ;
	wire _w30219_ ;
	wire _w30218_ ;
	wire _w30217_ ;
	wire _w30216_ ;
	wire _w30215_ ;
	wire _w30214_ ;
	wire _w30213_ ;
	wire _w30212_ ;
	wire _w30211_ ;
	wire _w30210_ ;
	wire _w30209_ ;
	wire _w30208_ ;
	wire _w30207_ ;
	wire _w30206_ ;
	wire _w30205_ ;
	wire _w30204_ ;
	wire _w30203_ ;
	wire _w30202_ ;
	wire _w30201_ ;
	wire _w30200_ ;
	wire _w30199_ ;
	wire _w30198_ ;
	wire _w30197_ ;
	wire _w30196_ ;
	wire _w30195_ ;
	wire _w30194_ ;
	wire _w30193_ ;
	wire _w30192_ ;
	wire _w30191_ ;
	wire _w30190_ ;
	wire _w30189_ ;
	wire _w30188_ ;
	wire _w30187_ ;
	wire _w30186_ ;
	wire _w30185_ ;
	wire _w30184_ ;
	wire _w30183_ ;
	wire _w30182_ ;
	wire _w30181_ ;
	wire _w30180_ ;
	wire _w30179_ ;
	wire _w30178_ ;
	wire _w30177_ ;
	wire _w30176_ ;
	wire _w30175_ ;
	wire _w30174_ ;
	wire _w30173_ ;
	wire _w30172_ ;
	wire _w30171_ ;
	wire _w30170_ ;
	wire _w30169_ ;
	wire _w30168_ ;
	wire _w30167_ ;
	wire _w30166_ ;
	wire _w30165_ ;
	wire _w30164_ ;
	wire _w30163_ ;
	wire _w30162_ ;
	wire _w30161_ ;
	wire _w30160_ ;
	wire _w30159_ ;
	wire _w30158_ ;
	wire _w30157_ ;
	wire _w30156_ ;
	wire _w30155_ ;
	wire _w30154_ ;
	wire _w30153_ ;
	wire _w30152_ ;
	wire _w30151_ ;
	wire _w30150_ ;
	wire _w30149_ ;
	wire _w30148_ ;
	wire _w30147_ ;
	wire _w30146_ ;
	wire _w30145_ ;
	wire _w30144_ ;
	wire _w30143_ ;
	wire _w30142_ ;
	wire _w30141_ ;
	wire _w30140_ ;
	wire _w30139_ ;
	wire _w30138_ ;
	wire _w30137_ ;
	wire _w30136_ ;
	wire _w30135_ ;
	wire _w30134_ ;
	wire _w30133_ ;
	wire _w30132_ ;
	wire _w30131_ ;
	wire _w30130_ ;
	wire _w30129_ ;
	wire _w30128_ ;
	wire _w30127_ ;
	wire _w30126_ ;
	wire _w30125_ ;
	wire _w30124_ ;
	wire _w30123_ ;
	wire _w30122_ ;
	wire _w30121_ ;
	wire _w30120_ ;
	wire _w30119_ ;
	wire _w30118_ ;
	wire _w30117_ ;
	wire _w30116_ ;
	wire _w30115_ ;
	wire _w30114_ ;
	wire _w30113_ ;
	wire _w30112_ ;
	wire _w30111_ ;
	wire _w30110_ ;
	wire _w30109_ ;
	wire _w30108_ ;
	wire _w30107_ ;
	wire _w30106_ ;
	wire _w30105_ ;
	wire _w30104_ ;
	wire _w30103_ ;
	wire _w30102_ ;
	wire _w30101_ ;
	wire _w30100_ ;
	wire _w30099_ ;
	wire _w30098_ ;
	wire _w30097_ ;
	wire _w30096_ ;
	wire _w30095_ ;
	wire _w30094_ ;
	wire _w30093_ ;
	wire _w30092_ ;
	wire _w30091_ ;
	wire _w30090_ ;
	wire _w30089_ ;
	wire _w30088_ ;
	wire _w30087_ ;
	wire _w30086_ ;
	wire _w30085_ ;
	wire _w30084_ ;
	wire _w30083_ ;
	wire _w30082_ ;
	wire _w30081_ ;
	wire _w30080_ ;
	wire _w30079_ ;
	wire _w30078_ ;
	wire _w30077_ ;
	wire _w30076_ ;
	wire _w30075_ ;
	wire _w30074_ ;
	wire _w30073_ ;
	wire _w30072_ ;
	wire _w30071_ ;
	wire _w30070_ ;
	wire _w30069_ ;
	wire _w30068_ ;
	wire _w30067_ ;
	wire _w30066_ ;
	wire _w30065_ ;
	wire _w30064_ ;
	wire _w30063_ ;
	wire _w30062_ ;
	wire _w30061_ ;
	wire _w30060_ ;
	wire _w30059_ ;
	wire _w30058_ ;
	wire _w30057_ ;
	wire _w30056_ ;
	wire _w30055_ ;
	wire _w30054_ ;
	wire _w30053_ ;
	wire _w30052_ ;
	wire _w30051_ ;
	wire _w30050_ ;
	wire _w30049_ ;
	wire _w30048_ ;
	wire _w30047_ ;
	wire _w30046_ ;
	wire _w30045_ ;
	wire _w30044_ ;
	wire _w30043_ ;
	wire _w30042_ ;
	wire _w30041_ ;
	wire _w30040_ ;
	wire _w30039_ ;
	wire _w30038_ ;
	wire _w30037_ ;
	wire _w30036_ ;
	wire _w30035_ ;
	wire _w30034_ ;
	wire _w30033_ ;
	wire _w30032_ ;
	wire _w30031_ ;
	wire _w30030_ ;
	wire _w30029_ ;
	wire _w30028_ ;
	wire _w30027_ ;
	wire _w30026_ ;
	wire _w30025_ ;
	wire _w30024_ ;
	wire _w30023_ ;
	wire _w30022_ ;
	wire _w30021_ ;
	wire _w30020_ ;
	wire _w30019_ ;
	wire _w30018_ ;
	wire _w30017_ ;
	wire _w30016_ ;
	wire _w30015_ ;
	wire _w30014_ ;
	wire _w30013_ ;
	wire _w30012_ ;
	wire _w30011_ ;
	wire _w30010_ ;
	wire _w30009_ ;
	wire _w30008_ ;
	wire _w30007_ ;
	wire _w30006_ ;
	wire _w30005_ ;
	wire _w30004_ ;
	wire _w30003_ ;
	wire _w30002_ ;
	wire _w30001_ ;
	wire _w30000_ ;
	wire _w29999_ ;
	wire _w29998_ ;
	wire _w29997_ ;
	wire _w29996_ ;
	wire _w29995_ ;
	wire _w29994_ ;
	wire _w29993_ ;
	wire _w29992_ ;
	wire _w29991_ ;
	wire _w29990_ ;
	wire _w29989_ ;
	wire _w29988_ ;
	wire _w29987_ ;
	wire _w29986_ ;
	wire _w29985_ ;
	wire _w29984_ ;
	wire _w29983_ ;
	wire _w29982_ ;
	wire _w29981_ ;
	wire _w29980_ ;
	wire _w29979_ ;
	wire _w29978_ ;
	wire _w29977_ ;
	wire _w29976_ ;
	wire _w29975_ ;
	wire _w29974_ ;
	wire _w29973_ ;
	wire _w29972_ ;
	wire _w29971_ ;
	wire _w29970_ ;
	wire _w29969_ ;
	wire _w29968_ ;
	wire _w29967_ ;
	wire _w29966_ ;
	wire _w29965_ ;
	wire _w29964_ ;
	wire _w29963_ ;
	wire _w29962_ ;
	wire _w29961_ ;
	wire _w29960_ ;
	wire _w29959_ ;
	wire _w29958_ ;
	wire _w29957_ ;
	wire _w29956_ ;
	wire _w29955_ ;
	wire _w29954_ ;
	wire _w29953_ ;
	wire _w29952_ ;
	wire _w29951_ ;
	wire _w29950_ ;
	wire _w29949_ ;
	wire _w29948_ ;
	wire _w29947_ ;
	wire _w29946_ ;
	wire _w29945_ ;
	wire _w29944_ ;
	wire _w29943_ ;
	wire _w29942_ ;
	wire _w29941_ ;
	wire _w29940_ ;
	wire _w29939_ ;
	wire _w29938_ ;
	wire _w29937_ ;
	wire _w29936_ ;
	wire _w29935_ ;
	wire _w29934_ ;
	wire _w29933_ ;
	wire _w29932_ ;
	wire _w29931_ ;
	wire _w29930_ ;
	wire _w29929_ ;
	wire _w29928_ ;
	wire _w29927_ ;
	wire _w29926_ ;
	wire _w29925_ ;
	wire _w29924_ ;
	wire _w29923_ ;
	wire _w29922_ ;
	wire _w29921_ ;
	wire _w29920_ ;
	wire _w29919_ ;
	wire _w29918_ ;
	wire _w29917_ ;
	wire _w29916_ ;
	wire _w29915_ ;
	wire _w29914_ ;
	wire _w29913_ ;
	wire _w29912_ ;
	wire _w29911_ ;
	wire _w29910_ ;
	wire _w29909_ ;
	wire _w29908_ ;
	wire _w29907_ ;
	wire _w29906_ ;
	wire _w29905_ ;
	wire _w29904_ ;
	wire _w29903_ ;
	wire _w29902_ ;
	wire _w29901_ ;
	wire _w29900_ ;
	wire _w29899_ ;
	wire _w29898_ ;
	wire _w29897_ ;
	wire _w29896_ ;
	wire _w29895_ ;
	wire _w29894_ ;
	wire _w29893_ ;
	wire _w29892_ ;
	wire _w29891_ ;
	wire _w29890_ ;
	wire _w29889_ ;
	wire _w29888_ ;
	wire _w29887_ ;
	wire _w29886_ ;
	wire _w29885_ ;
	wire _w29884_ ;
	wire _w29883_ ;
	wire _w29882_ ;
	wire _w29881_ ;
	wire _w29880_ ;
	wire _w29879_ ;
	wire _w29878_ ;
	wire _w29877_ ;
	wire _w29876_ ;
	wire _w29875_ ;
	wire _w29874_ ;
	wire _w29873_ ;
	wire _w29872_ ;
	wire _w29871_ ;
	wire _w29870_ ;
	wire _w29869_ ;
	wire _w29868_ ;
	wire _w29867_ ;
	wire _w29866_ ;
	wire _w29865_ ;
	wire _w29864_ ;
	wire _w29863_ ;
	wire _w29862_ ;
	wire _w29861_ ;
	wire _w29860_ ;
	wire _w29859_ ;
	wire _w29858_ ;
	wire _w29857_ ;
	wire _w29856_ ;
	wire _w29855_ ;
	wire _w29854_ ;
	wire _w29853_ ;
	wire _w29852_ ;
	wire _w29851_ ;
	wire _w29850_ ;
	wire _w29849_ ;
	wire _w29848_ ;
	wire _w29847_ ;
	wire _w29846_ ;
	wire _w29845_ ;
	wire _w29844_ ;
	wire _w29843_ ;
	wire _w29842_ ;
	wire _w29841_ ;
	wire _w29840_ ;
	wire _w29839_ ;
	wire _w29838_ ;
	wire _w29837_ ;
	wire _w29836_ ;
	wire _w29835_ ;
	wire _w29834_ ;
	wire _w29833_ ;
	wire _w29832_ ;
	wire _w29831_ ;
	wire _w29830_ ;
	wire _w29829_ ;
	wire _w29828_ ;
	wire _w29827_ ;
	wire _w29826_ ;
	wire _w29825_ ;
	wire _w29824_ ;
	wire _w29823_ ;
	wire _w29822_ ;
	wire _w29821_ ;
	wire _w29820_ ;
	wire _w29819_ ;
	wire _w29818_ ;
	wire _w29817_ ;
	wire _w29816_ ;
	wire _w29815_ ;
	wire _w29814_ ;
	wire _w29813_ ;
	wire _w29812_ ;
	wire _w29811_ ;
	wire _w29810_ ;
	wire _w29809_ ;
	wire _w29808_ ;
	wire _w29807_ ;
	wire _w29806_ ;
	wire _w29805_ ;
	wire _w29804_ ;
	wire _w29803_ ;
	wire _w29802_ ;
	wire _w29801_ ;
	wire _w29800_ ;
	wire _w29799_ ;
	wire _w29798_ ;
	wire _w29797_ ;
	wire _w29796_ ;
	wire _w29795_ ;
	wire _w29794_ ;
	wire _w29793_ ;
	wire _w29792_ ;
	wire _w29791_ ;
	wire _w29790_ ;
	wire _w29789_ ;
	wire _w29788_ ;
	wire _w29787_ ;
	wire _w29786_ ;
	wire _w29785_ ;
	wire _w29784_ ;
	wire _w29783_ ;
	wire _w29782_ ;
	wire _w29781_ ;
	wire _w29780_ ;
	wire _w29779_ ;
	wire _w29778_ ;
	wire _w29777_ ;
	wire _w29776_ ;
	wire _w29775_ ;
	wire _w29774_ ;
	wire _w29773_ ;
	wire _w29772_ ;
	wire _w29771_ ;
	wire _w29770_ ;
	wire _w29769_ ;
	wire _w29768_ ;
	wire _w29767_ ;
	wire _w29766_ ;
	wire _w29765_ ;
	wire _w29764_ ;
	wire _w29763_ ;
	wire _w29762_ ;
	wire _w29761_ ;
	wire _w29760_ ;
	wire _w29759_ ;
	wire _w29758_ ;
	wire _w29757_ ;
	wire _w29756_ ;
	wire _w29755_ ;
	wire _w29754_ ;
	wire _w29753_ ;
	wire _w29752_ ;
	wire _w29751_ ;
	wire _w29750_ ;
	wire _w29749_ ;
	wire _w29748_ ;
	wire _w29747_ ;
	wire _w29746_ ;
	wire _w29745_ ;
	wire _w29744_ ;
	wire _w29743_ ;
	wire _w29742_ ;
	wire _w29741_ ;
	wire _w29740_ ;
	wire _w29739_ ;
	wire _w29738_ ;
	wire _w29737_ ;
	wire _w29736_ ;
	wire _w29735_ ;
	wire _w29734_ ;
	wire _w29733_ ;
	wire _w29732_ ;
	wire _w29731_ ;
	wire _w29730_ ;
	wire _w29729_ ;
	wire _w29728_ ;
	wire _w29727_ ;
	wire _w29726_ ;
	wire _w29725_ ;
	wire _w29724_ ;
	wire _w29723_ ;
	wire _w29722_ ;
	wire _w29721_ ;
	wire _w29720_ ;
	wire _w29719_ ;
	wire _w29718_ ;
	wire _w29717_ ;
	wire _w29716_ ;
	wire _w29715_ ;
	wire _w29714_ ;
	wire _w29713_ ;
	wire _w29712_ ;
	wire _w29711_ ;
	wire _w29710_ ;
	wire _w29709_ ;
	wire _w29708_ ;
	wire _w29707_ ;
	wire _w29706_ ;
	wire _w29705_ ;
	wire _w29704_ ;
	wire _w29703_ ;
	wire _w29702_ ;
	wire _w29701_ ;
	wire _w29700_ ;
	wire _w29699_ ;
	wire _w29698_ ;
	wire _w29697_ ;
	wire _w29696_ ;
	wire _w29695_ ;
	wire _w29694_ ;
	wire _w29693_ ;
	wire _w29692_ ;
	wire _w29691_ ;
	wire _w29690_ ;
	wire _w29689_ ;
	wire _w29688_ ;
	wire _w29687_ ;
	wire _w29686_ ;
	wire _w29685_ ;
	wire _w29684_ ;
	wire _w29683_ ;
	wire _w29682_ ;
	wire _w29681_ ;
	wire _w29680_ ;
	wire _w29679_ ;
	wire _w29678_ ;
	wire _w29677_ ;
	wire _w29676_ ;
	wire _w29675_ ;
	wire _w29674_ ;
	wire _w29673_ ;
	wire _w29672_ ;
	wire _w29671_ ;
	wire _w29670_ ;
	wire _w29669_ ;
	wire _w29668_ ;
	wire _w29667_ ;
	wire _w29666_ ;
	wire _w29665_ ;
	wire _w29664_ ;
	wire _w29663_ ;
	wire _w29662_ ;
	wire _w29661_ ;
	wire _w29660_ ;
	wire _w29659_ ;
	wire _w29658_ ;
	wire _w29657_ ;
	wire _w29656_ ;
	wire _w29655_ ;
	wire _w29654_ ;
	wire _w29653_ ;
	wire _w29652_ ;
	wire _w29651_ ;
	wire _w29650_ ;
	wire _w29649_ ;
	wire _w29648_ ;
	wire _w29647_ ;
	wire _w29646_ ;
	wire _w29645_ ;
	wire _w29644_ ;
	wire _w29643_ ;
	wire _w29642_ ;
	wire _w29641_ ;
	wire _w29640_ ;
	wire _w29639_ ;
	wire _w29638_ ;
	wire _w29637_ ;
	wire _w29636_ ;
	wire _w29635_ ;
	wire _w29634_ ;
	wire _w29633_ ;
	wire _w29632_ ;
	wire _w29631_ ;
	wire _w29630_ ;
	wire _w29629_ ;
	wire _w29628_ ;
	wire _w29627_ ;
	wire _w29626_ ;
	wire _w29625_ ;
	wire _w29624_ ;
	wire _w29623_ ;
	wire _w29622_ ;
	wire _w29621_ ;
	wire _w29620_ ;
	wire _w29619_ ;
	wire _w29618_ ;
	wire _w29617_ ;
	wire _w29616_ ;
	wire _w29615_ ;
	wire _w29614_ ;
	wire _w29613_ ;
	wire _w29612_ ;
	wire _w29611_ ;
	wire _w29610_ ;
	wire _w29609_ ;
	wire _w29608_ ;
	wire _w29607_ ;
	wire _w29606_ ;
	wire _w29605_ ;
	wire _w29604_ ;
	wire _w29603_ ;
	wire _w29602_ ;
	wire _w29601_ ;
	wire _w29600_ ;
	wire _w29599_ ;
	wire _w29598_ ;
	wire _w29597_ ;
	wire _w29596_ ;
	wire _w29595_ ;
	wire _w29594_ ;
	wire _w29593_ ;
	wire _w29592_ ;
	wire _w29591_ ;
	wire _w29590_ ;
	wire _w29589_ ;
	wire _w29588_ ;
	wire _w29587_ ;
	wire _w29586_ ;
	wire _w29585_ ;
	wire _w29584_ ;
	wire _w29583_ ;
	wire _w29582_ ;
	wire _w29581_ ;
	wire _w29580_ ;
	wire _w29579_ ;
	wire _w29578_ ;
	wire _w29577_ ;
	wire _w29576_ ;
	wire _w29575_ ;
	wire _w29574_ ;
	wire _w29573_ ;
	wire _w29572_ ;
	wire _w29571_ ;
	wire _w29570_ ;
	wire _w29569_ ;
	wire _w29568_ ;
	wire _w29567_ ;
	wire _w29566_ ;
	wire _w29565_ ;
	wire _w29564_ ;
	wire _w29563_ ;
	wire _w29562_ ;
	wire _w29561_ ;
	wire _w29560_ ;
	wire _w29559_ ;
	wire _w29558_ ;
	wire _w29557_ ;
	wire _w29556_ ;
	wire _w29555_ ;
	wire _w29554_ ;
	wire _w29553_ ;
	wire _w29552_ ;
	wire _w29551_ ;
	wire _w29550_ ;
	wire _w29549_ ;
	wire _w29548_ ;
	wire _w29547_ ;
	wire _w29546_ ;
	wire _w29545_ ;
	wire _w29544_ ;
	wire _w29543_ ;
	wire _w29542_ ;
	wire _w29541_ ;
	wire _w29540_ ;
	wire _w29539_ ;
	wire _w29538_ ;
	wire _w29537_ ;
	wire _w29536_ ;
	wire _w29535_ ;
	wire _w29534_ ;
	wire _w29533_ ;
	wire _w29532_ ;
	wire _w29531_ ;
	wire _w29530_ ;
	wire _w29529_ ;
	wire _w29528_ ;
	wire _w29527_ ;
	wire _w29526_ ;
	wire _w29525_ ;
	wire _w29524_ ;
	wire _w29523_ ;
	wire _w29522_ ;
	wire _w29521_ ;
	wire _w29520_ ;
	wire _w29519_ ;
	wire _w29518_ ;
	wire _w29517_ ;
	wire _w29516_ ;
	wire _w29515_ ;
	wire _w29514_ ;
	wire _w29513_ ;
	wire _w29512_ ;
	wire _w29511_ ;
	wire _w29510_ ;
	wire _w29509_ ;
	wire _w29508_ ;
	wire _w29507_ ;
	wire _w29506_ ;
	wire _w29505_ ;
	wire _w29504_ ;
	wire _w29503_ ;
	wire _w29502_ ;
	wire _w29501_ ;
	wire _w29500_ ;
	wire _w29499_ ;
	wire _w29498_ ;
	wire _w29497_ ;
	wire _w29496_ ;
	wire _w29495_ ;
	wire _w29494_ ;
	wire _w29493_ ;
	wire _w29492_ ;
	wire _w29491_ ;
	wire _w29490_ ;
	wire _w29489_ ;
	wire _w29488_ ;
	wire _w29487_ ;
	wire _w29486_ ;
	wire _w29485_ ;
	wire _w29484_ ;
	wire _w29483_ ;
	wire _w29482_ ;
	wire _w29481_ ;
	wire _w29480_ ;
	wire _w29479_ ;
	wire _w29478_ ;
	wire _w29477_ ;
	wire _w29476_ ;
	wire _w29475_ ;
	wire _w29474_ ;
	wire _w29473_ ;
	wire _w29472_ ;
	wire _w29471_ ;
	wire _w29470_ ;
	wire _w29469_ ;
	wire _w29468_ ;
	wire _w29467_ ;
	wire _w29466_ ;
	wire _w29465_ ;
	wire _w29464_ ;
	wire _w29463_ ;
	wire _w29462_ ;
	wire _w29461_ ;
	wire _w29460_ ;
	wire _w29459_ ;
	wire _w29458_ ;
	wire _w29457_ ;
	wire _w29456_ ;
	wire _w29455_ ;
	wire _w29454_ ;
	wire _w29453_ ;
	wire _w29452_ ;
	wire _w29451_ ;
	wire _w29450_ ;
	wire _w29449_ ;
	wire _w29448_ ;
	wire _w29447_ ;
	wire _w29446_ ;
	wire _w29445_ ;
	wire _w29444_ ;
	wire _w29443_ ;
	wire _w29442_ ;
	wire _w29441_ ;
	wire _w29440_ ;
	wire _w29439_ ;
	wire _w29438_ ;
	wire _w29437_ ;
	wire _w29436_ ;
	wire _w29435_ ;
	wire _w29434_ ;
	wire _w29433_ ;
	wire _w29432_ ;
	wire _w29431_ ;
	wire _w29430_ ;
	wire _w29429_ ;
	wire _w29428_ ;
	wire _w29427_ ;
	wire _w29426_ ;
	wire _w29425_ ;
	wire _w29424_ ;
	wire _w29423_ ;
	wire _w29422_ ;
	wire _w29421_ ;
	wire _w29420_ ;
	wire _w29419_ ;
	wire _w29418_ ;
	wire _w29417_ ;
	wire _w29416_ ;
	wire _w29415_ ;
	wire _w29414_ ;
	wire _w29413_ ;
	wire _w29412_ ;
	wire _w29411_ ;
	wire _w29410_ ;
	wire _w29409_ ;
	wire _w29408_ ;
	wire _w29407_ ;
	wire _w29406_ ;
	wire _w29405_ ;
	wire _w29404_ ;
	wire _w29403_ ;
	wire _w29402_ ;
	wire _w29401_ ;
	wire _w29400_ ;
	wire _w29399_ ;
	wire _w29398_ ;
	wire _w29397_ ;
	wire _w29396_ ;
	wire _w29395_ ;
	wire _w29394_ ;
	wire _w29393_ ;
	wire _w29392_ ;
	wire _w29391_ ;
	wire _w29390_ ;
	wire _w29389_ ;
	wire _w29388_ ;
	wire _w29387_ ;
	wire _w29386_ ;
	wire _w29385_ ;
	wire _w29384_ ;
	wire _w29383_ ;
	wire _w29382_ ;
	wire _w29381_ ;
	wire _w29380_ ;
	wire _w29379_ ;
	wire _w29378_ ;
	wire _w29377_ ;
	wire _w29376_ ;
	wire _w29375_ ;
	wire _w29374_ ;
	wire _w29373_ ;
	wire _w29372_ ;
	wire _w29371_ ;
	wire _w29370_ ;
	wire _w29369_ ;
	wire _w29368_ ;
	wire _w29367_ ;
	wire _w29366_ ;
	wire _w29365_ ;
	wire _w29364_ ;
	wire _w29363_ ;
	wire _w29362_ ;
	wire _w29361_ ;
	wire _w29360_ ;
	wire _w29359_ ;
	wire _w29358_ ;
	wire _w29357_ ;
	wire _w29356_ ;
	wire _w29355_ ;
	wire _w29354_ ;
	wire _w29353_ ;
	wire _w29352_ ;
	wire _w29351_ ;
	wire _w29350_ ;
	wire _w29349_ ;
	wire _w29348_ ;
	wire _w29347_ ;
	wire _w29346_ ;
	wire _w29345_ ;
	wire _w29344_ ;
	wire _w29343_ ;
	wire _w29342_ ;
	wire _w29341_ ;
	wire _w29340_ ;
	wire _w29339_ ;
	wire _w29338_ ;
	wire _w29337_ ;
	wire _w29336_ ;
	wire _w29335_ ;
	wire _w29334_ ;
	wire _w29333_ ;
	wire _w29332_ ;
	wire _w29331_ ;
	wire _w29330_ ;
	wire _w29329_ ;
	wire _w29328_ ;
	wire _w29327_ ;
	wire _w29326_ ;
	wire _w29325_ ;
	wire _w29324_ ;
	wire _w29323_ ;
	wire _w29322_ ;
	wire _w29321_ ;
	wire _w29320_ ;
	wire _w29319_ ;
	wire _w29318_ ;
	wire _w29317_ ;
	wire _w29316_ ;
	wire _w29315_ ;
	wire _w29314_ ;
	wire _w29313_ ;
	wire _w29312_ ;
	wire _w29311_ ;
	wire _w29310_ ;
	wire _w29309_ ;
	wire _w29308_ ;
	wire _w29307_ ;
	wire _w29306_ ;
	wire _w29305_ ;
	wire _w29304_ ;
	wire _w29303_ ;
	wire _w29302_ ;
	wire _w29301_ ;
	wire _w29300_ ;
	wire _w29299_ ;
	wire _w29298_ ;
	wire _w29297_ ;
	wire _w29296_ ;
	wire _w29295_ ;
	wire _w29294_ ;
	wire _w29293_ ;
	wire _w29292_ ;
	wire _w29291_ ;
	wire _w29290_ ;
	wire _w29289_ ;
	wire _w29288_ ;
	wire _w29287_ ;
	wire _w29286_ ;
	wire _w29285_ ;
	wire _w29284_ ;
	wire _w29283_ ;
	wire _w29282_ ;
	wire _w29281_ ;
	wire _w29280_ ;
	wire _w29279_ ;
	wire _w29278_ ;
	wire _w29277_ ;
	wire _w29276_ ;
	wire _w29275_ ;
	wire _w29274_ ;
	wire _w29273_ ;
	wire _w29272_ ;
	wire _w29271_ ;
	wire _w29270_ ;
	wire _w29269_ ;
	wire _w29268_ ;
	wire _w29267_ ;
	wire _w29266_ ;
	wire _w29265_ ;
	wire _w29264_ ;
	wire _w29263_ ;
	wire _w29262_ ;
	wire _w29261_ ;
	wire _w29260_ ;
	wire _w29259_ ;
	wire _w29258_ ;
	wire _w29257_ ;
	wire _w29256_ ;
	wire _w29255_ ;
	wire _w29254_ ;
	wire _w29253_ ;
	wire _w29252_ ;
	wire _w29251_ ;
	wire _w29250_ ;
	wire _w29249_ ;
	wire _w29248_ ;
	wire _w29247_ ;
	wire _w29246_ ;
	wire _w29245_ ;
	wire _w29244_ ;
	wire _w29243_ ;
	wire _w29242_ ;
	wire _w29241_ ;
	wire _w29240_ ;
	wire _w29239_ ;
	wire _w29238_ ;
	wire _w29237_ ;
	wire _w29236_ ;
	wire _w29235_ ;
	wire _w29234_ ;
	wire _w29233_ ;
	wire _w29232_ ;
	wire _w29231_ ;
	wire _w29230_ ;
	wire _w29229_ ;
	wire _w29228_ ;
	wire _w29227_ ;
	wire _w29226_ ;
	wire _w29225_ ;
	wire _w29224_ ;
	wire _w29223_ ;
	wire _w29222_ ;
	wire _w29221_ ;
	wire _w29220_ ;
	wire _w29219_ ;
	wire _w29218_ ;
	wire _w29217_ ;
	wire _w29216_ ;
	wire _w29215_ ;
	wire _w29214_ ;
	wire _w29213_ ;
	wire _w29212_ ;
	wire _w29211_ ;
	wire _w29210_ ;
	wire _w29209_ ;
	wire _w29208_ ;
	wire _w29207_ ;
	wire _w29206_ ;
	wire _w29205_ ;
	wire _w29204_ ;
	wire _w29203_ ;
	wire _w29202_ ;
	wire _w29201_ ;
	wire _w29200_ ;
	wire _w29199_ ;
	wire _w29198_ ;
	wire _w29197_ ;
	wire _w29196_ ;
	wire _w29195_ ;
	wire _w29194_ ;
	wire _w29193_ ;
	wire _w29192_ ;
	wire _w29191_ ;
	wire _w29190_ ;
	wire _w29189_ ;
	wire _w29188_ ;
	wire _w29187_ ;
	wire _w29186_ ;
	wire _w29185_ ;
	wire _w29184_ ;
	wire _w29183_ ;
	wire _w29182_ ;
	wire _w29181_ ;
	wire _w29180_ ;
	wire _w29179_ ;
	wire _w29178_ ;
	wire _w29177_ ;
	wire _w29176_ ;
	wire _w29175_ ;
	wire _w29174_ ;
	wire _w29173_ ;
	wire _w29172_ ;
	wire _w29171_ ;
	wire _w29170_ ;
	wire _w29169_ ;
	wire _w29168_ ;
	wire _w29167_ ;
	wire _w29166_ ;
	wire _w29165_ ;
	wire _w29164_ ;
	wire _w29163_ ;
	wire _w29162_ ;
	wire _w29161_ ;
	wire _w29160_ ;
	wire _w29159_ ;
	wire _w29158_ ;
	wire _w29157_ ;
	wire _w29156_ ;
	wire _w29155_ ;
	wire _w29154_ ;
	wire _w29153_ ;
	wire _w29152_ ;
	wire _w29151_ ;
	wire _w29150_ ;
	wire _w29149_ ;
	wire _w29148_ ;
	wire _w29147_ ;
	wire _w29146_ ;
	wire _w29145_ ;
	wire _w29144_ ;
	wire _w29143_ ;
	wire _w29142_ ;
	wire _w29141_ ;
	wire _w29140_ ;
	wire _w29139_ ;
	wire _w29138_ ;
	wire _w29137_ ;
	wire _w29136_ ;
	wire _w29135_ ;
	wire _w29134_ ;
	wire _w29133_ ;
	wire _w29132_ ;
	wire _w29131_ ;
	wire _w29130_ ;
	wire _w29129_ ;
	wire _w29128_ ;
	wire _w29127_ ;
	wire _w29126_ ;
	wire _w29125_ ;
	wire _w29124_ ;
	wire _w29123_ ;
	wire _w29122_ ;
	wire _w29121_ ;
	wire _w29120_ ;
	wire _w29119_ ;
	wire _w29118_ ;
	wire _w29117_ ;
	wire _w29116_ ;
	wire _w29115_ ;
	wire _w29114_ ;
	wire _w29113_ ;
	wire _w29112_ ;
	wire _w29111_ ;
	wire _w29110_ ;
	wire _w29109_ ;
	wire _w29108_ ;
	wire _w29107_ ;
	wire _w29106_ ;
	wire _w29105_ ;
	wire _w29104_ ;
	wire _w29103_ ;
	wire _w29102_ ;
	wire _w29101_ ;
	wire _w29100_ ;
	wire _w29099_ ;
	wire _w29098_ ;
	wire _w29097_ ;
	wire _w29096_ ;
	wire _w29095_ ;
	wire _w29094_ ;
	wire _w29093_ ;
	wire _w29092_ ;
	wire _w29091_ ;
	wire _w29090_ ;
	wire _w29089_ ;
	wire _w29088_ ;
	wire _w29087_ ;
	wire _w29086_ ;
	wire _w29085_ ;
	wire _w29084_ ;
	wire _w29083_ ;
	wire _w29082_ ;
	wire _w29081_ ;
	wire _w29080_ ;
	wire _w29079_ ;
	wire _w29078_ ;
	wire _w29077_ ;
	wire _w29076_ ;
	wire _w29075_ ;
	wire _w29074_ ;
	wire _w29073_ ;
	wire _w29072_ ;
	wire _w29071_ ;
	wire _w29070_ ;
	wire _w29069_ ;
	wire _w29068_ ;
	wire _w29067_ ;
	wire _w29066_ ;
	wire _w29065_ ;
	wire _w29064_ ;
	wire _w29063_ ;
	wire _w29062_ ;
	wire _w29061_ ;
	wire _w29060_ ;
	wire _w29059_ ;
	wire _w29058_ ;
	wire _w29057_ ;
	wire _w29056_ ;
	wire _w29055_ ;
	wire _w29054_ ;
	wire _w29053_ ;
	wire _w29052_ ;
	wire _w29051_ ;
	wire _w29050_ ;
	wire _w29049_ ;
	wire _w29048_ ;
	wire _w29047_ ;
	wire _w29046_ ;
	wire _w29045_ ;
	wire _w29044_ ;
	wire _w29043_ ;
	wire _w29042_ ;
	wire _w29041_ ;
	wire _w29040_ ;
	wire _w29039_ ;
	wire _w29038_ ;
	wire _w29037_ ;
	wire _w29036_ ;
	wire _w29035_ ;
	wire _w29034_ ;
	wire _w29033_ ;
	wire _w29032_ ;
	wire _w29031_ ;
	wire _w29030_ ;
	wire _w29029_ ;
	wire _w29028_ ;
	wire _w29027_ ;
	wire _w29026_ ;
	wire _w29025_ ;
	wire _w29024_ ;
	wire _w29023_ ;
	wire _w29022_ ;
	wire _w29021_ ;
	wire _w29020_ ;
	wire _w29019_ ;
	wire _w29018_ ;
	wire _w29017_ ;
	wire _w29016_ ;
	wire _w29015_ ;
	wire _w29014_ ;
	wire _w29013_ ;
	wire _w29012_ ;
	wire _w29011_ ;
	wire _w29010_ ;
	wire _w29009_ ;
	wire _w29008_ ;
	wire _w29007_ ;
	wire _w29006_ ;
	wire _w29005_ ;
	wire _w29004_ ;
	wire _w29003_ ;
	wire _w29002_ ;
	wire _w29001_ ;
	wire _w29000_ ;
	wire _w28999_ ;
	wire _w28998_ ;
	wire _w28997_ ;
	wire _w28996_ ;
	wire _w28995_ ;
	wire _w28994_ ;
	wire _w28993_ ;
	wire _w28992_ ;
	wire _w28991_ ;
	wire _w28990_ ;
	wire _w28989_ ;
	wire _w28988_ ;
	wire _w28987_ ;
	wire _w28986_ ;
	wire _w28985_ ;
	wire _w28984_ ;
	wire _w28983_ ;
	wire _w28982_ ;
	wire _w28981_ ;
	wire _w28980_ ;
	wire _w28979_ ;
	wire _w28978_ ;
	wire _w28977_ ;
	wire _w28976_ ;
	wire _w28975_ ;
	wire _w28974_ ;
	wire _w28973_ ;
	wire _w28972_ ;
	wire _w28971_ ;
	wire _w28970_ ;
	wire _w28969_ ;
	wire _w28968_ ;
	wire _w28967_ ;
	wire _w28966_ ;
	wire _w28965_ ;
	wire _w28964_ ;
	wire _w28963_ ;
	wire _w28962_ ;
	wire _w28961_ ;
	wire _w28960_ ;
	wire _w28959_ ;
	wire _w28958_ ;
	wire _w28957_ ;
	wire _w28956_ ;
	wire _w28955_ ;
	wire _w28954_ ;
	wire _w28953_ ;
	wire _w28952_ ;
	wire _w28951_ ;
	wire _w28950_ ;
	wire _w28949_ ;
	wire _w28948_ ;
	wire _w28947_ ;
	wire _w28946_ ;
	wire _w28945_ ;
	wire _w28944_ ;
	wire _w28943_ ;
	wire _w28942_ ;
	wire _w28941_ ;
	wire _w28940_ ;
	wire _w28939_ ;
	wire _w28938_ ;
	wire _w28937_ ;
	wire _w28936_ ;
	wire _w28935_ ;
	wire _w28934_ ;
	wire _w28933_ ;
	wire _w28932_ ;
	wire _w28931_ ;
	wire _w28930_ ;
	wire _w28929_ ;
	wire _w28928_ ;
	wire _w28927_ ;
	wire _w28926_ ;
	wire _w28925_ ;
	wire _w28924_ ;
	wire _w28923_ ;
	wire _w28922_ ;
	wire _w28921_ ;
	wire _w28920_ ;
	wire _w28919_ ;
	wire _w28918_ ;
	wire _w28917_ ;
	wire _w28916_ ;
	wire _w28915_ ;
	wire _w28914_ ;
	wire _w28913_ ;
	wire _w28912_ ;
	wire _w28911_ ;
	wire _w28910_ ;
	wire _w28909_ ;
	wire _w28908_ ;
	wire _w28907_ ;
	wire _w28906_ ;
	wire _w28905_ ;
	wire _w28904_ ;
	wire _w28903_ ;
	wire _w28902_ ;
	wire _w28901_ ;
	wire _w28900_ ;
	wire _w28899_ ;
	wire _w28898_ ;
	wire _w28897_ ;
	wire _w28896_ ;
	wire _w28895_ ;
	wire _w28894_ ;
	wire _w28893_ ;
	wire _w28892_ ;
	wire _w28891_ ;
	wire _w28890_ ;
	wire _w28889_ ;
	wire _w28888_ ;
	wire _w28887_ ;
	wire _w28886_ ;
	wire _w28885_ ;
	wire _w28884_ ;
	wire _w28883_ ;
	wire _w28882_ ;
	wire _w28881_ ;
	wire _w28880_ ;
	wire _w28879_ ;
	wire _w28878_ ;
	wire _w28877_ ;
	wire _w28876_ ;
	wire _w28875_ ;
	wire _w28874_ ;
	wire _w28873_ ;
	wire _w28872_ ;
	wire _w28871_ ;
	wire _w28870_ ;
	wire _w28869_ ;
	wire _w28868_ ;
	wire _w28867_ ;
	wire _w28866_ ;
	wire _w28865_ ;
	wire _w28864_ ;
	wire _w28863_ ;
	wire _w28862_ ;
	wire _w28861_ ;
	wire _w28860_ ;
	wire _w28859_ ;
	wire _w28858_ ;
	wire _w28857_ ;
	wire _w28856_ ;
	wire _w28855_ ;
	wire _w28854_ ;
	wire _w28853_ ;
	wire _w28852_ ;
	wire _w28851_ ;
	wire _w28850_ ;
	wire _w28849_ ;
	wire _w28848_ ;
	wire _w28847_ ;
	wire _w28846_ ;
	wire _w28845_ ;
	wire _w28844_ ;
	wire _w28843_ ;
	wire _w28842_ ;
	wire _w28841_ ;
	wire _w28840_ ;
	wire _w28839_ ;
	wire _w28838_ ;
	wire _w28837_ ;
	wire _w28836_ ;
	wire _w28835_ ;
	wire _w28834_ ;
	wire _w28833_ ;
	wire _w28832_ ;
	wire _w28831_ ;
	wire _w28830_ ;
	wire _w28829_ ;
	wire _w28828_ ;
	wire _w28827_ ;
	wire _w28826_ ;
	wire _w28825_ ;
	wire _w28824_ ;
	wire _w28823_ ;
	wire _w28822_ ;
	wire _w28821_ ;
	wire _w28820_ ;
	wire _w28819_ ;
	wire _w28818_ ;
	wire _w28817_ ;
	wire _w28816_ ;
	wire _w28815_ ;
	wire _w28814_ ;
	wire _w28813_ ;
	wire _w28812_ ;
	wire _w28811_ ;
	wire _w28810_ ;
	wire _w28809_ ;
	wire _w28808_ ;
	wire _w28807_ ;
	wire _w28806_ ;
	wire _w28805_ ;
	wire _w28804_ ;
	wire _w28803_ ;
	wire _w28802_ ;
	wire _w28801_ ;
	wire _w28800_ ;
	wire _w28799_ ;
	wire _w28798_ ;
	wire _w28797_ ;
	wire _w28796_ ;
	wire _w28795_ ;
	wire _w28794_ ;
	wire _w28793_ ;
	wire _w28792_ ;
	wire _w28791_ ;
	wire _w28790_ ;
	wire _w28789_ ;
	wire _w28788_ ;
	wire _w28787_ ;
	wire _w28786_ ;
	wire _w28785_ ;
	wire _w28784_ ;
	wire _w28783_ ;
	wire _w28782_ ;
	wire _w28781_ ;
	wire _w28780_ ;
	wire _w28779_ ;
	wire _w28778_ ;
	wire _w28777_ ;
	wire _w28776_ ;
	wire _w28775_ ;
	wire _w28774_ ;
	wire _w28773_ ;
	wire _w28772_ ;
	wire _w28771_ ;
	wire _w28770_ ;
	wire _w28769_ ;
	wire _w28768_ ;
	wire _w28767_ ;
	wire _w28766_ ;
	wire _w28765_ ;
	wire _w28764_ ;
	wire _w28763_ ;
	wire _w28762_ ;
	wire _w28761_ ;
	wire _w28760_ ;
	wire _w28759_ ;
	wire _w28758_ ;
	wire _w28757_ ;
	wire _w28756_ ;
	wire _w28755_ ;
	wire _w28754_ ;
	wire _w28753_ ;
	wire _w28752_ ;
	wire _w28751_ ;
	wire _w28750_ ;
	wire _w28749_ ;
	wire _w28748_ ;
	wire _w28747_ ;
	wire _w28746_ ;
	wire _w28745_ ;
	wire _w28744_ ;
	wire _w28743_ ;
	wire _w28742_ ;
	wire _w28741_ ;
	wire _w28740_ ;
	wire _w28739_ ;
	wire _w28738_ ;
	wire _w28737_ ;
	wire _w28736_ ;
	wire _w28735_ ;
	wire _w28734_ ;
	wire _w28733_ ;
	wire _w28732_ ;
	wire _w28731_ ;
	wire _w28730_ ;
	wire _w28729_ ;
	wire _w28728_ ;
	wire _w28727_ ;
	wire _w28726_ ;
	wire _w28725_ ;
	wire _w28724_ ;
	wire _w28723_ ;
	wire _w28722_ ;
	wire _w28721_ ;
	wire _w28720_ ;
	wire _w28719_ ;
	wire _w28718_ ;
	wire _w28717_ ;
	wire _w28716_ ;
	wire _w28715_ ;
	wire _w28714_ ;
	wire _w28713_ ;
	wire _w28712_ ;
	wire _w28711_ ;
	wire _w28710_ ;
	wire _w28709_ ;
	wire _w28708_ ;
	wire _w28707_ ;
	wire _w28706_ ;
	wire _w28705_ ;
	wire _w28704_ ;
	wire _w28703_ ;
	wire _w28702_ ;
	wire _w28701_ ;
	wire _w28700_ ;
	wire _w28699_ ;
	wire _w28698_ ;
	wire _w28697_ ;
	wire _w28696_ ;
	wire _w28695_ ;
	wire _w28694_ ;
	wire _w28693_ ;
	wire _w28692_ ;
	wire _w28691_ ;
	wire _w28690_ ;
	wire _w28689_ ;
	wire _w28688_ ;
	wire _w28687_ ;
	wire _w28686_ ;
	wire _w28685_ ;
	wire _w28684_ ;
	wire _w28683_ ;
	wire _w28682_ ;
	wire _w28681_ ;
	wire _w28680_ ;
	wire _w28679_ ;
	wire _w28678_ ;
	wire _w28677_ ;
	wire _w28676_ ;
	wire _w28675_ ;
	wire _w28674_ ;
	wire _w28673_ ;
	wire _w28672_ ;
	wire _w28671_ ;
	wire _w28670_ ;
	wire _w28669_ ;
	wire _w28668_ ;
	wire _w28667_ ;
	wire _w28666_ ;
	wire _w28665_ ;
	wire _w28664_ ;
	wire _w28663_ ;
	wire _w28662_ ;
	wire _w28661_ ;
	wire _w28660_ ;
	wire _w28659_ ;
	wire _w28658_ ;
	wire _w28657_ ;
	wire _w28656_ ;
	wire _w28655_ ;
	wire _w28654_ ;
	wire _w28653_ ;
	wire _w28652_ ;
	wire _w28651_ ;
	wire _w28650_ ;
	wire _w28649_ ;
	wire _w28648_ ;
	wire _w28647_ ;
	wire _w28646_ ;
	wire _w28645_ ;
	wire _w28644_ ;
	wire _w28643_ ;
	wire _w28642_ ;
	wire _w28641_ ;
	wire _w28640_ ;
	wire _w28639_ ;
	wire _w28638_ ;
	wire _w28637_ ;
	wire _w28636_ ;
	wire _w28635_ ;
	wire _w28634_ ;
	wire _w28633_ ;
	wire _w28632_ ;
	wire _w28631_ ;
	wire _w28630_ ;
	wire _w28629_ ;
	wire _w28628_ ;
	wire _w28627_ ;
	wire _w28626_ ;
	wire _w28625_ ;
	wire _w28624_ ;
	wire _w28623_ ;
	wire _w28622_ ;
	wire _w28621_ ;
	wire _w28620_ ;
	wire _w28619_ ;
	wire _w28618_ ;
	wire _w28617_ ;
	wire _w28616_ ;
	wire _w28615_ ;
	wire _w28614_ ;
	wire _w28613_ ;
	wire _w28612_ ;
	wire _w28611_ ;
	wire _w28610_ ;
	wire _w28609_ ;
	wire _w28608_ ;
	wire _w28607_ ;
	wire _w28606_ ;
	wire _w28605_ ;
	wire _w28604_ ;
	wire _w28603_ ;
	wire _w28602_ ;
	wire _w28601_ ;
	wire _w28600_ ;
	wire _w28599_ ;
	wire _w28598_ ;
	wire _w28597_ ;
	wire _w28596_ ;
	wire _w28595_ ;
	wire _w28594_ ;
	wire _w28593_ ;
	wire _w28592_ ;
	wire _w28591_ ;
	wire _w28590_ ;
	wire _w28589_ ;
	wire _w28588_ ;
	wire _w28587_ ;
	wire _w28586_ ;
	wire _w28585_ ;
	wire _w28584_ ;
	wire _w28583_ ;
	wire _w28582_ ;
	wire _w28581_ ;
	wire _w28580_ ;
	wire _w28579_ ;
	wire _w28578_ ;
	wire _w28577_ ;
	wire _w28576_ ;
	wire _w28575_ ;
	wire _w28574_ ;
	wire _w28573_ ;
	wire _w28572_ ;
	wire _w28571_ ;
	wire _w28570_ ;
	wire _w28569_ ;
	wire _w28568_ ;
	wire _w28567_ ;
	wire _w28566_ ;
	wire _w28565_ ;
	wire _w28564_ ;
	wire _w28563_ ;
	wire _w28562_ ;
	wire _w28561_ ;
	wire _w28560_ ;
	wire _w28559_ ;
	wire _w28558_ ;
	wire _w28557_ ;
	wire _w28556_ ;
	wire _w28555_ ;
	wire _w28554_ ;
	wire _w28553_ ;
	wire _w28552_ ;
	wire _w28551_ ;
	wire _w28550_ ;
	wire _w28549_ ;
	wire _w28548_ ;
	wire _w28547_ ;
	wire _w28546_ ;
	wire _w28545_ ;
	wire _w28544_ ;
	wire _w28543_ ;
	wire _w28542_ ;
	wire _w28541_ ;
	wire _w28540_ ;
	wire _w28539_ ;
	wire _w28538_ ;
	wire _w28537_ ;
	wire _w28536_ ;
	wire _w28535_ ;
	wire _w28534_ ;
	wire _w28533_ ;
	wire _w28532_ ;
	wire _w28531_ ;
	wire _w28530_ ;
	wire _w28529_ ;
	wire _w28528_ ;
	wire _w28527_ ;
	wire _w28526_ ;
	wire _w28525_ ;
	wire _w28524_ ;
	wire _w28523_ ;
	wire _w28522_ ;
	wire _w28521_ ;
	wire _w28520_ ;
	wire _w28519_ ;
	wire _w28518_ ;
	wire _w28517_ ;
	wire _w28516_ ;
	wire _w28515_ ;
	wire _w28514_ ;
	wire _w28513_ ;
	wire _w28512_ ;
	wire _w28511_ ;
	wire _w28510_ ;
	wire _w28509_ ;
	wire _w28508_ ;
	wire _w28507_ ;
	wire _w28506_ ;
	wire _w28505_ ;
	wire _w28504_ ;
	wire _w28503_ ;
	wire _w28502_ ;
	wire _w28501_ ;
	wire _w28500_ ;
	wire _w28499_ ;
	wire _w28498_ ;
	wire _w28497_ ;
	wire _w28496_ ;
	wire _w28495_ ;
	wire _w28494_ ;
	wire _w28493_ ;
	wire _w28492_ ;
	wire _w28491_ ;
	wire _w28490_ ;
	wire _w28489_ ;
	wire _w28488_ ;
	wire _w28487_ ;
	wire _w28486_ ;
	wire _w28485_ ;
	wire _w28484_ ;
	wire _w28483_ ;
	wire _w28482_ ;
	wire _w28481_ ;
	wire _w28480_ ;
	wire _w28479_ ;
	wire _w28478_ ;
	wire _w28477_ ;
	wire _w28476_ ;
	wire _w28475_ ;
	wire _w28474_ ;
	wire _w28473_ ;
	wire _w28472_ ;
	wire _w28471_ ;
	wire _w28470_ ;
	wire _w28469_ ;
	wire _w28468_ ;
	wire _w28467_ ;
	wire _w28466_ ;
	wire _w28465_ ;
	wire _w28464_ ;
	wire _w28463_ ;
	wire _w28462_ ;
	wire _w28461_ ;
	wire _w28460_ ;
	wire _w28459_ ;
	wire _w28458_ ;
	wire _w28457_ ;
	wire _w28456_ ;
	wire _w28455_ ;
	wire _w28454_ ;
	wire _w28453_ ;
	wire _w28452_ ;
	wire _w28451_ ;
	wire _w28450_ ;
	wire _w28449_ ;
	wire _w28448_ ;
	wire _w28447_ ;
	wire _w28446_ ;
	wire _w28445_ ;
	wire _w28444_ ;
	wire _w28443_ ;
	wire _w28442_ ;
	wire _w28441_ ;
	wire _w28440_ ;
	wire _w28439_ ;
	wire _w28438_ ;
	wire _w28437_ ;
	wire _w28436_ ;
	wire _w28435_ ;
	wire _w28434_ ;
	wire _w28433_ ;
	wire _w28432_ ;
	wire _w28431_ ;
	wire _w28430_ ;
	wire _w28429_ ;
	wire _w28428_ ;
	wire _w28427_ ;
	wire _w28426_ ;
	wire _w28425_ ;
	wire _w28424_ ;
	wire _w28423_ ;
	wire _w28422_ ;
	wire _w28421_ ;
	wire _w28420_ ;
	wire _w28419_ ;
	wire _w28418_ ;
	wire _w28417_ ;
	wire _w28416_ ;
	wire _w28415_ ;
	wire _w28414_ ;
	wire _w28413_ ;
	wire _w28412_ ;
	wire _w28411_ ;
	wire _w28410_ ;
	wire _w28409_ ;
	wire _w28408_ ;
	wire _w28407_ ;
	wire _w28406_ ;
	wire _w28405_ ;
	wire _w28404_ ;
	wire _w28403_ ;
	wire _w28402_ ;
	wire _w28401_ ;
	wire _w28400_ ;
	wire _w28399_ ;
	wire _w28398_ ;
	wire _w28397_ ;
	wire _w28396_ ;
	wire _w28395_ ;
	wire _w28394_ ;
	wire _w28393_ ;
	wire _w28392_ ;
	wire _w28391_ ;
	wire _w28390_ ;
	wire _w28389_ ;
	wire _w28388_ ;
	wire _w28387_ ;
	wire _w28386_ ;
	wire _w28385_ ;
	wire _w28384_ ;
	wire _w28383_ ;
	wire _w28382_ ;
	wire _w28381_ ;
	wire _w28380_ ;
	wire _w28379_ ;
	wire _w28378_ ;
	wire _w28377_ ;
	wire _w28376_ ;
	wire _w28375_ ;
	wire _w28374_ ;
	wire _w28373_ ;
	wire _w28372_ ;
	wire _w28371_ ;
	wire _w28370_ ;
	wire _w28369_ ;
	wire _w28368_ ;
	wire _w28367_ ;
	wire _w28366_ ;
	wire _w28365_ ;
	wire _w28364_ ;
	wire _w28363_ ;
	wire _w28362_ ;
	wire _w28361_ ;
	wire _w28360_ ;
	wire _w28359_ ;
	wire _w28358_ ;
	wire _w28357_ ;
	wire _w28356_ ;
	wire _w28355_ ;
	wire _w28354_ ;
	wire _w28353_ ;
	wire _w28352_ ;
	wire _w28351_ ;
	wire _w28350_ ;
	wire _w28349_ ;
	wire _w28348_ ;
	wire _w28347_ ;
	wire _w28346_ ;
	wire _w28345_ ;
	wire _w28344_ ;
	wire _w28343_ ;
	wire _w28342_ ;
	wire _w28341_ ;
	wire _w28340_ ;
	wire _w28339_ ;
	wire _w28338_ ;
	wire _w28337_ ;
	wire _w28336_ ;
	wire _w28335_ ;
	wire _w28334_ ;
	wire _w28333_ ;
	wire _w28332_ ;
	wire _w28331_ ;
	wire _w28330_ ;
	wire _w28329_ ;
	wire _w28328_ ;
	wire _w28327_ ;
	wire _w28326_ ;
	wire _w28325_ ;
	wire _w28324_ ;
	wire _w28323_ ;
	wire _w28322_ ;
	wire _w28321_ ;
	wire _w28320_ ;
	wire _w28319_ ;
	wire _w28318_ ;
	wire _w28317_ ;
	wire _w28316_ ;
	wire _w28315_ ;
	wire _w28314_ ;
	wire _w28313_ ;
	wire _w28312_ ;
	wire _w28311_ ;
	wire _w28310_ ;
	wire _w28309_ ;
	wire _w28308_ ;
	wire _w28307_ ;
	wire _w28306_ ;
	wire _w28305_ ;
	wire _w28304_ ;
	wire _w28303_ ;
	wire _w28302_ ;
	wire _w28301_ ;
	wire _w28300_ ;
	wire _w28299_ ;
	wire _w28298_ ;
	wire _w28297_ ;
	wire _w28296_ ;
	wire _w28295_ ;
	wire _w28294_ ;
	wire _w28293_ ;
	wire _w28292_ ;
	wire _w28291_ ;
	wire _w28290_ ;
	wire _w28289_ ;
	wire _w28288_ ;
	wire _w28287_ ;
	wire _w28286_ ;
	wire _w28285_ ;
	wire _w28284_ ;
	wire _w28283_ ;
	wire _w28282_ ;
	wire _w28281_ ;
	wire _w28280_ ;
	wire _w28279_ ;
	wire _w28278_ ;
	wire _w28277_ ;
	wire _w28276_ ;
	wire _w28275_ ;
	wire _w28274_ ;
	wire _w28273_ ;
	wire _w28272_ ;
	wire _w28271_ ;
	wire _w28270_ ;
	wire _w28269_ ;
	wire _w28268_ ;
	wire _w28267_ ;
	wire _w28266_ ;
	wire _w28265_ ;
	wire _w28264_ ;
	wire _w28263_ ;
	wire _w28262_ ;
	wire _w28261_ ;
	wire _w28260_ ;
	wire _w28259_ ;
	wire _w28258_ ;
	wire _w28257_ ;
	wire _w28256_ ;
	wire _w28255_ ;
	wire _w28254_ ;
	wire _w28253_ ;
	wire _w28252_ ;
	wire _w28251_ ;
	wire _w28250_ ;
	wire _w28249_ ;
	wire _w28248_ ;
	wire _w28247_ ;
	wire _w28246_ ;
	wire _w28245_ ;
	wire _w28244_ ;
	wire _w28243_ ;
	wire _w28242_ ;
	wire _w28241_ ;
	wire _w28240_ ;
	wire _w28239_ ;
	wire _w28238_ ;
	wire _w28237_ ;
	wire _w28236_ ;
	wire _w28235_ ;
	wire _w28234_ ;
	wire _w28233_ ;
	wire _w28232_ ;
	wire _w28231_ ;
	wire _w28230_ ;
	wire _w28229_ ;
	wire _w28228_ ;
	wire _w28227_ ;
	wire _w28226_ ;
	wire _w28225_ ;
	wire _w28224_ ;
	wire _w28223_ ;
	wire _w28222_ ;
	wire _w28221_ ;
	wire _w28220_ ;
	wire _w28219_ ;
	wire _w28218_ ;
	wire _w28217_ ;
	wire _w28216_ ;
	wire _w28215_ ;
	wire _w28214_ ;
	wire _w28213_ ;
	wire _w28212_ ;
	wire _w28211_ ;
	wire _w28210_ ;
	wire _w28209_ ;
	wire _w28208_ ;
	wire _w28207_ ;
	wire _w28206_ ;
	wire _w28205_ ;
	wire _w28204_ ;
	wire _w28203_ ;
	wire _w28202_ ;
	wire _w28201_ ;
	wire _w28200_ ;
	wire _w28199_ ;
	wire _w28198_ ;
	wire _w28197_ ;
	wire _w28196_ ;
	wire _w28195_ ;
	wire _w28194_ ;
	wire _w28193_ ;
	wire _w28192_ ;
	wire _w28191_ ;
	wire _w28190_ ;
	wire _w28189_ ;
	wire _w28188_ ;
	wire _w28187_ ;
	wire _w28186_ ;
	wire _w28185_ ;
	wire _w28184_ ;
	wire _w28183_ ;
	wire _w28182_ ;
	wire _w28181_ ;
	wire _w28180_ ;
	wire _w28179_ ;
	wire _w28178_ ;
	wire _w28177_ ;
	wire _w28176_ ;
	wire _w28175_ ;
	wire _w28174_ ;
	wire _w28173_ ;
	wire _w28172_ ;
	wire _w28171_ ;
	wire _w28170_ ;
	wire _w28169_ ;
	wire _w28168_ ;
	wire _w28167_ ;
	wire _w28166_ ;
	wire _w28165_ ;
	wire _w28164_ ;
	wire _w28163_ ;
	wire _w28162_ ;
	wire _w28161_ ;
	wire _w28160_ ;
	wire _w28159_ ;
	wire _w28158_ ;
	wire _w28157_ ;
	wire _w28156_ ;
	wire _w28155_ ;
	wire _w28154_ ;
	wire _w28153_ ;
	wire _w28152_ ;
	wire _w28151_ ;
	wire _w28150_ ;
	wire _w28149_ ;
	wire _w28148_ ;
	wire _w28147_ ;
	wire _w28146_ ;
	wire _w28145_ ;
	wire _w28144_ ;
	wire _w28143_ ;
	wire _w28142_ ;
	wire _w28141_ ;
	wire _w28140_ ;
	wire _w28139_ ;
	wire _w28138_ ;
	wire _w28137_ ;
	wire _w28136_ ;
	wire _w28135_ ;
	wire _w28134_ ;
	wire _w28133_ ;
	wire _w28132_ ;
	wire _w28131_ ;
	wire _w28130_ ;
	wire _w28129_ ;
	wire _w28128_ ;
	wire _w28127_ ;
	wire _w28126_ ;
	wire _w28125_ ;
	wire _w28124_ ;
	wire _w28123_ ;
	wire _w28122_ ;
	wire _w28121_ ;
	wire _w28120_ ;
	wire _w28119_ ;
	wire _w28118_ ;
	wire _w28117_ ;
	wire _w28116_ ;
	wire _w28115_ ;
	wire _w28114_ ;
	wire _w28113_ ;
	wire _w28112_ ;
	wire _w28111_ ;
	wire _w28110_ ;
	wire _w28109_ ;
	wire _w28108_ ;
	wire _w28107_ ;
	wire _w28106_ ;
	wire _w28105_ ;
	wire _w28104_ ;
	wire _w28103_ ;
	wire _w28102_ ;
	wire _w28101_ ;
	wire _w28100_ ;
	wire _w28099_ ;
	wire _w28098_ ;
	wire _w28097_ ;
	wire _w28096_ ;
	wire _w28095_ ;
	wire _w28094_ ;
	wire _w28093_ ;
	wire _w28092_ ;
	wire _w28091_ ;
	wire _w28090_ ;
	wire _w28089_ ;
	wire _w28088_ ;
	wire _w28087_ ;
	wire _w28086_ ;
	wire _w28085_ ;
	wire _w28084_ ;
	wire _w28083_ ;
	wire _w28082_ ;
	wire _w28081_ ;
	wire _w28080_ ;
	wire _w28079_ ;
	wire _w28078_ ;
	wire _w28077_ ;
	wire _w28076_ ;
	wire _w28075_ ;
	wire _w28074_ ;
	wire _w28073_ ;
	wire _w28072_ ;
	wire _w28071_ ;
	wire _w28070_ ;
	wire _w28069_ ;
	wire _w28068_ ;
	wire _w28067_ ;
	wire _w28066_ ;
	wire _w28065_ ;
	wire _w28064_ ;
	wire _w28063_ ;
	wire _w28062_ ;
	wire _w28061_ ;
	wire _w28060_ ;
	wire _w28059_ ;
	wire _w28058_ ;
	wire _w28057_ ;
	wire _w28056_ ;
	wire _w28055_ ;
	wire _w28054_ ;
	wire _w28053_ ;
	wire _w28052_ ;
	wire _w28051_ ;
	wire _w28050_ ;
	wire _w28049_ ;
	wire _w28048_ ;
	wire _w28047_ ;
	wire _w28046_ ;
	wire _w28045_ ;
	wire _w28044_ ;
	wire _w28043_ ;
	wire _w28042_ ;
	wire _w28041_ ;
	wire _w28040_ ;
	wire _w28039_ ;
	wire _w28038_ ;
	wire _w28037_ ;
	wire _w28036_ ;
	wire _w28035_ ;
	wire _w28034_ ;
	wire _w28033_ ;
	wire _w28032_ ;
	wire _w28031_ ;
	wire _w28030_ ;
	wire _w28029_ ;
	wire _w28028_ ;
	wire _w28027_ ;
	wire _w28026_ ;
	wire _w28025_ ;
	wire _w28024_ ;
	wire _w28023_ ;
	wire _w28022_ ;
	wire _w28021_ ;
	wire _w28020_ ;
	wire _w28019_ ;
	wire _w28018_ ;
	wire _w28017_ ;
	wire _w28016_ ;
	wire _w28015_ ;
	wire _w28014_ ;
	wire _w28013_ ;
	wire _w28012_ ;
	wire _w28011_ ;
	wire _w28010_ ;
	wire _w28009_ ;
	wire _w28008_ ;
	wire _w28007_ ;
	wire _w28006_ ;
	wire _w28005_ ;
	wire _w28004_ ;
	wire _w28003_ ;
	wire _w28002_ ;
	wire _w28001_ ;
	wire _w28000_ ;
	wire _w27999_ ;
	wire _w27998_ ;
	wire _w27997_ ;
	wire _w27996_ ;
	wire _w27995_ ;
	wire _w27994_ ;
	wire _w27993_ ;
	wire _w27992_ ;
	wire _w27991_ ;
	wire _w27990_ ;
	wire _w27989_ ;
	wire _w27988_ ;
	wire _w27987_ ;
	wire _w27986_ ;
	wire _w27985_ ;
	wire _w27984_ ;
	wire _w27983_ ;
	wire _w27982_ ;
	wire _w27981_ ;
	wire _w27980_ ;
	wire _w27979_ ;
	wire _w27978_ ;
	wire _w27977_ ;
	wire _w27976_ ;
	wire _w27975_ ;
	wire _w27974_ ;
	wire _w27973_ ;
	wire _w27972_ ;
	wire _w27971_ ;
	wire _w27970_ ;
	wire _w27969_ ;
	wire _w27968_ ;
	wire _w27967_ ;
	wire _w27966_ ;
	wire _w27965_ ;
	wire _w27964_ ;
	wire _w27963_ ;
	wire _w27962_ ;
	wire _w27961_ ;
	wire _w27960_ ;
	wire _w27959_ ;
	wire _w27958_ ;
	wire _w27957_ ;
	wire _w27956_ ;
	wire _w27955_ ;
	wire _w27954_ ;
	wire _w27953_ ;
	wire _w27952_ ;
	wire _w27951_ ;
	wire _w27950_ ;
	wire _w27949_ ;
	wire _w27948_ ;
	wire _w27947_ ;
	wire _w27946_ ;
	wire _w27945_ ;
	wire _w27944_ ;
	wire _w27943_ ;
	wire _w27942_ ;
	wire _w27941_ ;
	wire _w27940_ ;
	wire _w27939_ ;
	wire _w27938_ ;
	wire _w27937_ ;
	wire _w27936_ ;
	wire _w27935_ ;
	wire _w27934_ ;
	wire _w27933_ ;
	wire _w27932_ ;
	wire _w27931_ ;
	wire _w27930_ ;
	wire _w27929_ ;
	wire _w27928_ ;
	wire _w27927_ ;
	wire _w27926_ ;
	wire _w27925_ ;
	wire _w27924_ ;
	wire _w27923_ ;
	wire _w27922_ ;
	wire _w27921_ ;
	wire _w27920_ ;
	wire _w27919_ ;
	wire _w27918_ ;
	wire _w27917_ ;
	wire _w27916_ ;
	wire _w27915_ ;
	wire _w27914_ ;
	wire _w27913_ ;
	wire _w27912_ ;
	wire _w27911_ ;
	wire _w27910_ ;
	wire _w27909_ ;
	wire _w27908_ ;
	wire _w27907_ ;
	wire _w27906_ ;
	wire _w27905_ ;
	wire _w27904_ ;
	wire _w27903_ ;
	wire _w27902_ ;
	wire _w27901_ ;
	wire _w27900_ ;
	wire _w27899_ ;
	wire _w27898_ ;
	wire _w27897_ ;
	wire _w27896_ ;
	wire _w27895_ ;
	wire _w27894_ ;
	wire _w27893_ ;
	wire _w27892_ ;
	wire _w27891_ ;
	wire _w27890_ ;
	wire _w27889_ ;
	wire _w27888_ ;
	wire _w27887_ ;
	wire _w27886_ ;
	wire _w27885_ ;
	wire _w27884_ ;
	wire _w27883_ ;
	wire _w27882_ ;
	wire _w27881_ ;
	wire _w27880_ ;
	wire _w27879_ ;
	wire _w27878_ ;
	wire _w27877_ ;
	wire _w27876_ ;
	wire _w27875_ ;
	wire _w27874_ ;
	wire _w27873_ ;
	wire _w27872_ ;
	wire _w27871_ ;
	wire _w27870_ ;
	wire _w27869_ ;
	wire _w27868_ ;
	wire _w27867_ ;
	wire _w27866_ ;
	wire _w27865_ ;
	wire _w27864_ ;
	wire _w27863_ ;
	wire _w27862_ ;
	wire _w27861_ ;
	wire _w27860_ ;
	wire _w27859_ ;
	wire _w27858_ ;
	wire _w27857_ ;
	wire _w27856_ ;
	wire _w27855_ ;
	wire _w27854_ ;
	wire _w27853_ ;
	wire _w27852_ ;
	wire _w27851_ ;
	wire _w27850_ ;
	wire _w27849_ ;
	wire _w27848_ ;
	wire _w27847_ ;
	wire _w27846_ ;
	wire _w27845_ ;
	wire _w27844_ ;
	wire _w27843_ ;
	wire _w27842_ ;
	wire _w27841_ ;
	wire _w27840_ ;
	wire _w27839_ ;
	wire _w27838_ ;
	wire _w27837_ ;
	wire _w27836_ ;
	wire _w27835_ ;
	wire _w27834_ ;
	wire _w27833_ ;
	wire _w27832_ ;
	wire _w27831_ ;
	wire _w27830_ ;
	wire _w27829_ ;
	wire _w27828_ ;
	wire _w27827_ ;
	wire _w27826_ ;
	wire _w27825_ ;
	wire _w27824_ ;
	wire _w27823_ ;
	wire _w27822_ ;
	wire _w27821_ ;
	wire _w27820_ ;
	wire _w27819_ ;
	wire _w27818_ ;
	wire _w27817_ ;
	wire _w27816_ ;
	wire _w27815_ ;
	wire _w27814_ ;
	wire _w27813_ ;
	wire _w27812_ ;
	wire _w27811_ ;
	wire _w27810_ ;
	wire _w27809_ ;
	wire _w27808_ ;
	wire _w27807_ ;
	wire _w27806_ ;
	wire _w27805_ ;
	wire _w27804_ ;
	wire _w27803_ ;
	wire _w27802_ ;
	wire _w27801_ ;
	wire _w27800_ ;
	wire _w27799_ ;
	wire _w27798_ ;
	wire _w27797_ ;
	wire _w27796_ ;
	wire _w27795_ ;
	wire _w27794_ ;
	wire _w27793_ ;
	wire _w27792_ ;
	wire _w27791_ ;
	wire _w27790_ ;
	wire _w27789_ ;
	wire _w27788_ ;
	wire _w27787_ ;
	wire _w27786_ ;
	wire _w27785_ ;
	wire _w27784_ ;
	wire _w27783_ ;
	wire _w27782_ ;
	wire _w27781_ ;
	wire _w27780_ ;
	wire _w27779_ ;
	wire _w27778_ ;
	wire _w27777_ ;
	wire _w27776_ ;
	wire _w27775_ ;
	wire _w27774_ ;
	wire _w27773_ ;
	wire _w27772_ ;
	wire _w27771_ ;
	wire _w27770_ ;
	wire _w27769_ ;
	wire _w27768_ ;
	wire _w27767_ ;
	wire _w27766_ ;
	wire _w27765_ ;
	wire _w27764_ ;
	wire _w27763_ ;
	wire _w27762_ ;
	wire _w27761_ ;
	wire _w27760_ ;
	wire _w27759_ ;
	wire _w27758_ ;
	wire _w27757_ ;
	wire _w27756_ ;
	wire _w27755_ ;
	wire _w27754_ ;
	wire _w27753_ ;
	wire _w27752_ ;
	wire _w27751_ ;
	wire _w27750_ ;
	wire _w27749_ ;
	wire _w27748_ ;
	wire _w27747_ ;
	wire _w27746_ ;
	wire _w27745_ ;
	wire _w27744_ ;
	wire _w27743_ ;
	wire _w27742_ ;
	wire _w27741_ ;
	wire _w27740_ ;
	wire _w27739_ ;
	wire _w27738_ ;
	wire _w27737_ ;
	wire _w27736_ ;
	wire _w27735_ ;
	wire _w27734_ ;
	wire _w27733_ ;
	wire _w27732_ ;
	wire _w27731_ ;
	wire _w27730_ ;
	wire _w27729_ ;
	wire _w27728_ ;
	wire _w27727_ ;
	wire _w27726_ ;
	wire _w27725_ ;
	wire _w27724_ ;
	wire _w27723_ ;
	wire _w27722_ ;
	wire _w27721_ ;
	wire _w27720_ ;
	wire _w27719_ ;
	wire _w27718_ ;
	wire _w27717_ ;
	wire _w27716_ ;
	wire _w27715_ ;
	wire _w27714_ ;
	wire _w27713_ ;
	wire _w27712_ ;
	wire _w27711_ ;
	wire _w27710_ ;
	wire _w27709_ ;
	wire _w27708_ ;
	wire _w27707_ ;
	wire _w27706_ ;
	wire _w27705_ ;
	wire _w27704_ ;
	wire _w27703_ ;
	wire _w27702_ ;
	wire _w27701_ ;
	wire _w27700_ ;
	wire _w27699_ ;
	wire _w27698_ ;
	wire _w27697_ ;
	wire _w27696_ ;
	wire _w27695_ ;
	wire _w27694_ ;
	wire _w27693_ ;
	wire _w27692_ ;
	wire _w27691_ ;
	wire _w27690_ ;
	wire _w27689_ ;
	wire _w27688_ ;
	wire _w27687_ ;
	wire _w27686_ ;
	wire _w27685_ ;
	wire _w27684_ ;
	wire _w27683_ ;
	wire _w27682_ ;
	wire _w27681_ ;
	wire _w27680_ ;
	wire _w27679_ ;
	wire _w27678_ ;
	wire _w27677_ ;
	wire _w27676_ ;
	wire _w27675_ ;
	wire _w27674_ ;
	wire _w27673_ ;
	wire _w27672_ ;
	wire _w27671_ ;
	wire _w27670_ ;
	wire _w27669_ ;
	wire _w27668_ ;
	wire _w27667_ ;
	wire _w27666_ ;
	wire _w27665_ ;
	wire _w27664_ ;
	wire _w27663_ ;
	wire _w27662_ ;
	wire _w27661_ ;
	wire _w27660_ ;
	wire _w27659_ ;
	wire _w27658_ ;
	wire _w27657_ ;
	wire _w27656_ ;
	wire _w27655_ ;
	wire _w27654_ ;
	wire _w27653_ ;
	wire _w27652_ ;
	wire _w27651_ ;
	wire _w27650_ ;
	wire _w27649_ ;
	wire _w27648_ ;
	wire _w27647_ ;
	wire _w27646_ ;
	wire _w27645_ ;
	wire _w27644_ ;
	wire _w27643_ ;
	wire _w27642_ ;
	wire _w27641_ ;
	wire _w27640_ ;
	wire _w27639_ ;
	wire _w27638_ ;
	wire _w27637_ ;
	wire _w27636_ ;
	wire _w27635_ ;
	wire _w27634_ ;
	wire _w27633_ ;
	wire _w27632_ ;
	wire _w27631_ ;
	wire _w27630_ ;
	wire _w27629_ ;
	wire _w27628_ ;
	wire _w27627_ ;
	wire _w27626_ ;
	wire _w27625_ ;
	wire _w27624_ ;
	wire _w27623_ ;
	wire _w27622_ ;
	wire _w27621_ ;
	wire _w27620_ ;
	wire _w27619_ ;
	wire _w27618_ ;
	wire _w27617_ ;
	wire _w27616_ ;
	wire _w27615_ ;
	wire _w27614_ ;
	wire _w27613_ ;
	wire _w27612_ ;
	wire _w27611_ ;
	wire _w27610_ ;
	wire _w27609_ ;
	wire _w27608_ ;
	wire _w27607_ ;
	wire _w27606_ ;
	wire _w27605_ ;
	wire _w27604_ ;
	wire _w27603_ ;
	wire _w27602_ ;
	wire _w27601_ ;
	wire _w27600_ ;
	wire _w27599_ ;
	wire _w27598_ ;
	wire _w27597_ ;
	wire _w27596_ ;
	wire _w27595_ ;
	wire _w27594_ ;
	wire _w27593_ ;
	wire _w27592_ ;
	wire _w27591_ ;
	wire _w27590_ ;
	wire _w27589_ ;
	wire _w27588_ ;
	wire _w27587_ ;
	wire _w27586_ ;
	wire _w27585_ ;
	wire _w27584_ ;
	wire _w27583_ ;
	wire _w27582_ ;
	wire _w27581_ ;
	wire _w27580_ ;
	wire _w27579_ ;
	wire _w27578_ ;
	wire _w27577_ ;
	wire _w27576_ ;
	wire _w27575_ ;
	wire _w27574_ ;
	wire _w27573_ ;
	wire _w27572_ ;
	wire _w27571_ ;
	wire _w27570_ ;
	wire _w27569_ ;
	wire _w27568_ ;
	wire _w27567_ ;
	wire _w27566_ ;
	wire _w27565_ ;
	wire _w27564_ ;
	wire _w27563_ ;
	wire _w27562_ ;
	wire _w27561_ ;
	wire _w27560_ ;
	wire _w27559_ ;
	wire _w27558_ ;
	wire _w27557_ ;
	wire _w27556_ ;
	wire _w27555_ ;
	wire _w27554_ ;
	wire _w27553_ ;
	wire _w27552_ ;
	wire _w27551_ ;
	wire _w27550_ ;
	wire _w27549_ ;
	wire _w27548_ ;
	wire _w27547_ ;
	wire _w27546_ ;
	wire _w27545_ ;
	wire _w27544_ ;
	wire _w27543_ ;
	wire _w27542_ ;
	wire _w27541_ ;
	wire _w27540_ ;
	wire _w27539_ ;
	wire _w27538_ ;
	wire _w27537_ ;
	wire _w27536_ ;
	wire _w27535_ ;
	wire _w27534_ ;
	wire _w27533_ ;
	wire _w27532_ ;
	wire _w27531_ ;
	wire _w27530_ ;
	wire _w27529_ ;
	wire _w27528_ ;
	wire _w27527_ ;
	wire _w27526_ ;
	wire _w27525_ ;
	wire _w27524_ ;
	wire _w27523_ ;
	wire _w27522_ ;
	wire _w27521_ ;
	wire _w27520_ ;
	wire _w27519_ ;
	wire _w27518_ ;
	wire _w27517_ ;
	wire _w27516_ ;
	wire _w27515_ ;
	wire _w27514_ ;
	wire _w27513_ ;
	wire _w27512_ ;
	wire _w27511_ ;
	wire _w27510_ ;
	wire _w27509_ ;
	wire _w27508_ ;
	wire _w27507_ ;
	wire _w27506_ ;
	wire _w27505_ ;
	wire _w27504_ ;
	wire _w27503_ ;
	wire _w27502_ ;
	wire _w27501_ ;
	wire _w27500_ ;
	wire _w27499_ ;
	wire _w27498_ ;
	wire _w27497_ ;
	wire _w27496_ ;
	wire _w27495_ ;
	wire _w27494_ ;
	wire _w27493_ ;
	wire _w27492_ ;
	wire _w27491_ ;
	wire _w27490_ ;
	wire _w27489_ ;
	wire _w27488_ ;
	wire _w27487_ ;
	wire _w27486_ ;
	wire _w27485_ ;
	wire _w27484_ ;
	wire _w27483_ ;
	wire _w27482_ ;
	wire _w27481_ ;
	wire _w27480_ ;
	wire _w27479_ ;
	wire _w27478_ ;
	wire _w27477_ ;
	wire _w27476_ ;
	wire _w27475_ ;
	wire _w27474_ ;
	wire _w27473_ ;
	wire _w27472_ ;
	wire _w27471_ ;
	wire _w27470_ ;
	wire _w27469_ ;
	wire _w27468_ ;
	wire _w27467_ ;
	wire _w27466_ ;
	wire _w27465_ ;
	wire _w27464_ ;
	wire _w27463_ ;
	wire _w27462_ ;
	wire _w27461_ ;
	wire _w27460_ ;
	wire _w27459_ ;
	wire _w27458_ ;
	wire _w27457_ ;
	wire _w27456_ ;
	wire _w27455_ ;
	wire _w27454_ ;
	wire _w27453_ ;
	wire _w27452_ ;
	wire _w27451_ ;
	wire _w27450_ ;
	wire _w27449_ ;
	wire _w27448_ ;
	wire _w27447_ ;
	wire _w27446_ ;
	wire _w27445_ ;
	wire _w27444_ ;
	wire _w27443_ ;
	wire _w27442_ ;
	wire _w27441_ ;
	wire _w27440_ ;
	wire _w27439_ ;
	wire _w27438_ ;
	wire _w27437_ ;
	wire _w27436_ ;
	wire _w27435_ ;
	wire _w27434_ ;
	wire _w27433_ ;
	wire _w27432_ ;
	wire _w27431_ ;
	wire _w27430_ ;
	wire _w27429_ ;
	wire _w27428_ ;
	wire _w27427_ ;
	wire _w27426_ ;
	wire _w27425_ ;
	wire _w27424_ ;
	wire _w27423_ ;
	wire _w27422_ ;
	wire _w27421_ ;
	wire _w27420_ ;
	wire _w27419_ ;
	wire _w27418_ ;
	wire _w27417_ ;
	wire _w27416_ ;
	wire _w27415_ ;
	wire _w27414_ ;
	wire _w27413_ ;
	wire _w27412_ ;
	wire _w27411_ ;
	wire _w27410_ ;
	wire _w27409_ ;
	wire _w27408_ ;
	wire _w27407_ ;
	wire _w27406_ ;
	wire _w27405_ ;
	wire _w27404_ ;
	wire _w27403_ ;
	wire _w27402_ ;
	wire _w27401_ ;
	wire _w27400_ ;
	wire _w27399_ ;
	wire _w27398_ ;
	wire _w27397_ ;
	wire _w27396_ ;
	wire _w27395_ ;
	wire _w27394_ ;
	wire _w27393_ ;
	wire _w27392_ ;
	wire _w27391_ ;
	wire _w27390_ ;
	wire _w27389_ ;
	wire _w27388_ ;
	wire _w27387_ ;
	wire _w27386_ ;
	wire _w27385_ ;
	wire _w27384_ ;
	wire _w27383_ ;
	wire _w27382_ ;
	wire _w27381_ ;
	wire _w27380_ ;
	wire _w27379_ ;
	wire _w27378_ ;
	wire _w27377_ ;
	wire _w27376_ ;
	wire _w27375_ ;
	wire _w27374_ ;
	wire _w27373_ ;
	wire _w27372_ ;
	wire _w27371_ ;
	wire _w27370_ ;
	wire _w27369_ ;
	wire _w27368_ ;
	wire _w27367_ ;
	wire _w27366_ ;
	wire _w27365_ ;
	wire _w27364_ ;
	wire _w27363_ ;
	wire _w27362_ ;
	wire _w27361_ ;
	wire _w27360_ ;
	wire _w27359_ ;
	wire _w27358_ ;
	wire _w27357_ ;
	wire _w27356_ ;
	wire _w27355_ ;
	wire _w27354_ ;
	wire _w27353_ ;
	wire _w27352_ ;
	wire _w27351_ ;
	wire _w27350_ ;
	wire _w27349_ ;
	wire _w27348_ ;
	wire _w27347_ ;
	wire _w27346_ ;
	wire _w27345_ ;
	wire _w27344_ ;
	wire _w27343_ ;
	wire _w27342_ ;
	wire _w27341_ ;
	wire _w27340_ ;
	wire _w27339_ ;
	wire _w27338_ ;
	wire _w27337_ ;
	wire _w27336_ ;
	wire _w27335_ ;
	wire _w27334_ ;
	wire _w27333_ ;
	wire _w27332_ ;
	wire _w27331_ ;
	wire _w27330_ ;
	wire _w27329_ ;
	wire _w27328_ ;
	wire _w27327_ ;
	wire _w27326_ ;
	wire _w27325_ ;
	wire _w27324_ ;
	wire _w27323_ ;
	wire _w27322_ ;
	wire _w27321_ ;
	wire _w27320_ ;
	wire _w27319_ ;
	wire _w27318_ ;
	wire _w27317_ ;
	wire _w27316_ ;
	wire _w27315_ ;
	wire _w27314_ ;
	wire _w27313_ ;
	wire _w27312_ ;
	wire _w27311_ ;
	wire _w27310_ ;
	wire _w27309_ ;
	wire _w27308_ ;
	wire _w27307_ ;
	wire _w27306_ ;
	wire _w27305_ ;
	wire _w27304_ ;
	wire _w27303_ ;
	wire _w27302_ ;
	wire _w27301_ ;
	wire _w27300_ ;
	wire _w27299_ ;
	wire _w27298_ ;
	wire _w27297_ ;
	wire _w27296_ ;
	wire _w27295_ ;
	wire _w27294_ ;
	wire _w27293_ ;
	wire _w27292_ ;
	wire _w27291_ ;
	wire _w27290_ ;
	wire _w27289_ ;
	wire _w27288_ ;
	wire _w27287_ ;
	wire _w27286_ ;
	wire _w27285_ ;
	wire _w27284_ ;
	wire _w27283_ ;
	wire _w27282_ ;
	wire _w27281_ ;
	wire _w27280_ ;
	wire _w27279_ ;
	wire _w27278_ ;
	wire _w27277_ ;
	wire _w27276_ ;
	wire _w27275_ ;
	wire _w27274_ ;
	wire _w27273_ ;
	wire _w27272_ ;
	wire _w27271_ ;
	wire _w27270_ ;
	wire _w27269_ ;
	wire _w27268_ ;
	wire _w27267_ ;
	wire _w27266_ ;
	wire _w27265_ ;
	wire _w27264_ ;
	wire _w27263_ ;
	wire _w27262_ ;
	wire _w27261_ ;
	wire _w27260_ ;
	wire _w27259_ ;
	wire _w27258_ ;
	wire _w27257_ ;
	wire _w27256_ ;
	wire _w27255_ ;
	wire _w27254_ ;
	wire _w27253_ ;
	wire _w27252_ ;
	wire _w27251_ ;
	wire _w27250_ ;
	wire _w27249_ ;
	wire _w27248_ ;
	wire _w27247_ ;
	wire _w27246_ ;
	wire _w27245_ ;
	wire _w27244_ ;
	wire _w27243_ ;
	wire _w27242_ ;
	wire _w27241_ ;
	wire _w27240_ ;
	wire _w27239_ ;
	wire _w27238_ ;
	wire _w27237_ ;
	wire _w27236_ ;
	wire _w27235_ ;
	wire _w27234_ ;
	wire _w27233_ ;
	wire _w27232_ ;
	wire _w27231_ ;
	wire _w27230_ ;
	wire _w27229_ ;
	wire _w27228_ ;
	wire _w27227_ ;
	wire _w27226_ ;
	wire _w27225_ ;
	wire _w27224_ ;
	wire _w27223_ ;
	wire _w27222_ ;
	wire _w27221_ ;
	wire _w27220_ ;
	wire _w27219_ ;
	wire _w27218_ ;
	wire _w27217_ ;
	wire _w27216_ ;
	wire _w27215_ ;
	wire _w27214_ ;
	wire _w27213_ ;
	wire _w27212_ ;
	wire _w27211_ ;
	wire _w27210_ ;
	wire _w27209_ ;
	wire _w27208_ ;
	wire _w27207_ ;
	wire _w27206_ ;
	wire _w27205_ ;
	wire _w27204_ ;
	wire _w27203_ ;
	wire _w27202_ ;
	wire _w27201_ ;
	wire _w27200_ ;
	wire _w27199_ ;
	wire _w27198_ ;
	wire _w27197_ ;
	wire _w27196_ ;
	wire _w27195_ ;
	wire _w27194_ ;
	wire _w27193_ ;
	wire _w27192_ ;
	wire _w27191_ ;
	wire _w27190_ ;
	wire _w27189_ ;
	wire _w27188_ ;
	wire _w27187_ ;
	wire _w27186_ ;
	wire _w27185_ ;
	wire _w27184_ ;
	wire _w27183_ ;
	wire _w27182_ ;
	wire _w27181_ ;
	wire _w27180_ ;
	wire _w27179_ ;
	wire _w27178_ ;
	wire _w27177_ ;
	wire _w27176_ ;
	wire _w27175_ ;
	wire _w27174_ ;
	wire _w27173_ ;
	wire _w27172_ ;
	wire _w27171_ ;
	wire _w27170_ ;
	wire _w27169_ ;
	wire _w27168_ ;
	wire _w27167_ ;
	wire _w27166_ ;
	wire _w27165_ ;
	wire _w27164_ ;
	wire _w27163_ ;
	wire _w27162_ ;
	wire _w27161_ ;
	wire _w27160_ ;
	wire _w27159_ ;
	wire _w27158_ ;
	wire _w27157_ ;
	wire _w27156_ ;
	wire _w27155_ ;
	wire _w27154_ ;
	wire _w27153_ ;
	wire _w27152_ ;
	wire _w27151_ ;
	wire _w27150_ ;
	wire _w27149_ ;
	wire _w27148_ ;
	wire _w27147_ ;
	wire _w27146_ ;
	wire _w27145_ ;
	wire _w27144_ ;
	wire _w27143_ ;
	wire _w27142_ ;
	wire _w27141_ ;
	wire _w27140_ ;
	wire _w27139_ ;
	wire _w27138_ ;
	wire _w27137_ ;
	wire _w27136_ ;
	wire _w27135_ ;
	wire _w27134_ ;
	wire _w27133_ ;
	wire _w27132_ ;
	wire _w27131_ ;
	wire _w27130_ ;
	wire _w27129_ ;
	wire _w27128_ ;
	wire _w27127_ ;
	wire _w27126_ ;
	wire _w27125_ ;
	wire _w27124_ ;
	wire _w27123_ ;
	wire _w27122_ ;
	wire _w27121_ ;
	wire _w27120_ ;
	wire _w27119_ ;
	wire _w27118_ ;
	wire _w27117_ ;
	wire _w27116_ ;
	wire _w27115_ ;
	wire _w27114_ ;
	wire _w27113_ ;
	wire _w27112_ ;
	wire _w27111_ ;
	wire _w27110_ ;
	wire _w27109_ ;
	wire _w27108_ ;
	wire _w27107_ ;
	wire _w27106_ ;
	wire _w27105_ ;
	wire _w27104_ ;
	wire _w27103_ ;
	wire _w27102_ ;
	wire _w27101_ ;
	wire _w27100_ ;
	wire _w27099_ ;
	wire _w27098_ ;
	wire _w27097_ ;
	wire _w27096_ ;
	wire _w27095_ ;
	wire _w27094_ ;
	wire _w27093_ ;
	wire _w27092_ ;
	wire _w27091_ ;
	wire _w27090_ ;
	wire _w27089_ ;
	wire _w27088_ ;
	wire _w27087_ ;
	wire _w27086_ ;
	wire _w27085_ ;
	wire _w27084_ ;
	wire _w27083_ ;
	wire _w27082_ ;
	wire _w27081_ ;
	wire _w27080_ ;
	wire _w27079_ ;
	wire _w27078_ ;
	wire _w27077_ ;
	wire _w27076_ ;
	wire _w27075_ ;
	wire _w27074_ ;
	wire _w27073_ ;
	wire _w27072_ ;
	wire _w27071_ ;
	wire _w27070_ ;
	wire _w27069_ ;
	wire _w27068_ ;
	wire _w27067_ ;
	wire _w27066_ ;
	wire _w27065_ ;
	wire _w27064_ ;
	wire _w27063_ ;
	wire _w27062_ ;
	wire _w27061_ ;
	wire _w27060_ ;
	wire _w27059_ ;
	wire _w27058_ ;
	wire _w27057_ ;
	wire _w27056_ ;
	wire _w27055_ ;
	wire _w27054_ ;
	wire _w27053_ ;
	wire _w27052_ ;
	wire _w27051_ ;
	wire _w27050_ ;
	wire _w27049_ ;
	wire _w27048_ ;
	wire _w27047_ ;
	wire _w27046_ ;
	wire _w27045_ ;
	wire _w27044_ ;
	wire _w27043_ ;
	wire _w27042_ ;
	wire _w27041_ ;
	wire _w27040_ ;
	wire _w27039_ ;
	wire _w27038_ ;
	wire _w27037_ ;
	wire _w27036_ ;
	wire _w27035_ ;
	wire _w27034_ ;
	wire _w27033_ ;
	wire _w27032_ ;
	wire _w27031_ ;
	wire _w27030_ ;
	wire _w27029_ ;
	wire _w27028_ ;
	wire _w27027_ ;
	wire _w27026_ ;
	wire _w27025_ ;
	wire _w27024_ ;
	wire _w27023_ ;
	wire _w27022_ ;
	wire _w27021_ ;
	wire _w27020_ ;
	wire _w27019_ ;
	wire _w27018_ ;
	wire _w27017_ ;
	wire _w27016_ ;
	wire _w27015_ ;
	wire _w27014_ ;
	wire _w27013_ ;
	wire _w27012_ ;
	wire _w27011_ ;
	wire _w27010_ ;
	wire _w27009_ ;
	wire _w27008_ ;
	wire _w27007_ ;
	wire _w27006_ ;
	wire _w27005_ ;
	wire _w27004_ ;
	wire _w27003_ ;
	wire _w27002_ ;
	wire _w27001_ ;
	wire _w27000_ ;
	wire _w26999_ ;
	wire _w26998_ ;
	wire _w26997_ ;
	wire _w26996_ ;
	wire _w26995_ ;
	wire _w26994_ ;
	wire _w26993_ ;
	wire _w26992_ ;
	wire _w26991_ ;
	wire _w26990_ ;
	wire _w26989_ ;
	wire _w26988_ ;
	wire _w26987_ ;
	wire _w26986_ ;
	wire _w26985_ ;
	wire _w26984_ ;
	wire _w26983_ ;
	wire _w26982_ ;
	wire _w26981_ ;
	wire _w26980_ ;
	wire _w26979_ ;
	wire _w26978_ ;
	wire _w26977_ ;
	wire _w26976_ ;
	wire _w26975_ ;
	wire _w26974_ ;
	wire _w26973_ ;
	wire _w26972_ ;
	wire _w26971_ ;
	wire _w26970_ ;
	wire _w26969_ ;
	wire _w26968_ ;
	wire _w26967_ ;
	wire _w26966_ ;
	wire _w26965_ ;
	wire _w26964_ ;
	wire _w26963_ ;
	wire _w26962_ ;
	wire _w26961_ ;
	wire _w26960_ ;
	wire _w26959_ ;
	wire _w26958_ ;
	wire _w26957_ ;
	wire _w26956_ ;
	wire _w26955_ ;
	wire _w26954_ ;
	wire _w26953_ ;
	wire _w26952_ ;
	wire _w26951_ ;
	wire _w26950_ ;
	wire _w26949_ ;
	wire _w26948_ ;
	wire _w26947_ ;
	wire _w26946_ ;
	wire _w26945_ ;
	wire _w26944_ ;
	wire _w26943_ ;
	wire _w26942_ ;
	wire _w26941_ ;
	wire _w26940_ ;
	wire _w26939_ ;
	wire _w26938_ ;
	wire _w26937_ ;
	wire _w26936_ ;
	wire _w26935_ ;
	wire _w26934_ ;
	wire _w26933_ ;
	wire _w26932_ ;
	wire _w26931_ ;
	wire _w26930_ ;
	wire _w26929_ ;
	wire _w26928_ ;
	wire _w26927_ ;
	wire _w26926_ ;
	wire _w26925_ ;
	wire _w26924_ ;
	wire _w26923_ ;
	wire _w26922_ ;
	wire _w26921_ ;
	wire _w26920_ ;
	wire _w26919_ ;
	wire _w26918_ ;
	wire _w26917_ ;
	wire _w26916_ ;
	wire _w26915_ ;
	wire _w26914_ ;
	wire _w26913_ ;
	wire _w26912_ ;
	wire _w26911_ ;
	wire _w26910_ ;
	wire _w26909_ ;
	wire _w26908_ ;
	wire _w26907_ ;
	wire _w26906_ ;
	wire _w26905_ ;
	wire _w26904_ ;
	wire _w26903_ ;
	wire _w26902_ ;
	wire _w26901_ ;
	wire _w26900_ ;
	wire _w26899_ ;
	wire _w26898_ ;
	wire _w26897_ ;
	wire _w26896_ ;
	wire _w26895_ ;
	wire _w26894_ ;
	wire _w26893_ ;
	wire _w26892_ ;
	wire _w26891_ ;
	wire _w26890_ ;
	wire _w26889_ ;
	wire _w26888_ ;
	wire _w26887_ ;
	wire _w26886_ ;
	wire _w26885_ ;
	wire _w26884_ ;
	wire _w26883_ ;
	wire _w26882_ ;
	wire _w26881_ ;
	wire _w26880_ ;
	wire _w26879_ ;
	wire _w26878_ ;
	wire _w26877_ ;
	wire _w26876_ ;
	wire _w26875_ ;
	wire _w26874_ ;
	wire _w26873_ ;
	wire _w26872_ ;
	wire _w26871_ ;
	wire _w26870_ ;
	wire _w26869_ ;
	wire _w26868_ ;
	wire _w26867_ ;
	wire _w26866_ ;
	wire _w26865_ ;
	wire _w26864_ ;
	wire _w26863_ ;
	wire _w26862_ ;
	wire _w26861_ ;
	wire _w26860_ ;
	wire _w26859_ ;
	wire _w26858_ ;
	wire _w26857_ ;
	wire _w26856_ ;
	wire _w26855_ ;
	wire _w26854_ ;
	wire _w26853_ ;
	wire _w26852_ ;
	wire _w26851_ ;
	wire _w26850_ ;
	wire _w26849_ ;
	wire _w26848_ ;
	wire _w26847_ ;
	wire _w26846_ ;
	wire _w26845_ ;
	wire _w26844_ ;
	wire _w26843_ ;
	wire _w26842_ ;
	wire _w26841_ ;
	wire _w26840_ ;
	wire _w26839_ ;
	wire _w26838_ ;
	wire _w26837_ ;
	wire _w26836_ ;
	wire _w26835_ ;
	wire _w26834_ ;
	wire _w26833_ ;
	wire _w26832_ ;
	wire _w26831_ ;
	wire _w26830_ ;
	wire _w26829_ ;
	wire _w26828_ ;
	wire _w26827_ ;
	wire _w26826_ ;
	wire _w26825_ ;
	wire _w26824_ ;
	wire _w26823_ ;
	wire _w26822_ ;
	wire _w26821_ ;
	wire _w26820_ ;
	wire _w26819_ ;
	wire _w26818_ ;
	wire _w26817_ ;
	wire _w26816_ ;
	wire _w26815_ ;
	wire _w26814_ ;
	wire _w26813_ ;
	wire _w26812_ ;
	wire _w26811_ ;
	wire _w26810_ ;
	wire _w26809_ ;
	wire _w26808_ ;
	wire _w26807_ ;
	wire _w26806_ ;
	wire _w26805_ ;
	wire _w26804_ ;
	wire _w26803_ ;
	wire _w26802_ ;
	wire _w26801_ ;
	wire _w26800_ ;
	wire _w26799_ ;
	wire _w26798_ ;
	wire _w26797_ ;
	wire _w26796_ ;
	wire _w26795_ ;
	wire _w26794_ ;
	wire _w26793_ ;
	wire _w26792_ ;
	wire _w26791_ ;
	wire _w26790_ ;
	wire _w26789_ ;
	wire _w26788_ ;
	wire _w26787_ ;
	wire _w26786_ ;
	wire _w26785_ ;
	wire _w26784_ ;
	wire _w26783_ ;
	wire _w26782_ ;
	wire _w26781_ ;
	wire _w26780_ ;
	wire _w26779_ ;
	wire _w26778_ ;
	wire _w26777_ ;
	wire _w26776_ ;
	wire _w26775_ ;
	wire _w26774_ ;
	wire _w26773_ ;
	wire _w26772_ ;
	wire _w26771_ ;
	wire _w26770_ ;
	wire _w26769_ ;
	wire _w26768_ ;
	wire _w26767_ ;
	wire _w26766_ ;
	wire _w26765_ ;
	wire _w26764_ ;
	wire _w26763_ ;
	wire _w26762_ ;
	wire _w26761_ ;
	wire _w26760_ ;
	wire _w26759_ ;
	wire _w26758_ ;
	wire _w26757_ ;
	wire _w26756_ ;
	wire _w26755_ ;
	wire _w26754_ ;
	wire _w26753_ ;
	wire _w26752_ ;
	wire _w26751_ ;
	wire _w26750_ ;
	wire _w26749_ ;
	wire _w26748_ ;
	wire _w26747_ ;
	wire _w26746_ ;
	wire _w26745_ ;
	wire _w26744_ ;
	wire _w26743_ ;
	wire _w26742_ ;
	wire _w26741_ ;
	wire _w26740_ ;
	wire _w26739_ ;
	wire _w26738_ ;
	wire _w26737_ ;
	wire _w26736_ ;
	wire _w26735_ ;
	wire _w26734_ ;
	wire _w26733_ ;
	wire _w26732_ ;
	wire _w26731_ ;
	wire _w26730_ ;
	wire _w26729_ ;
	wire _w26728_ ;
	wire _w26727_ ;
	wire _w26726_ ;
	wire _w26725_ ;
	wire _w26724_ ;
	wire _w26723_ ;
	wire _w26722_ ;
	wire _w26721_ ;
	wire _w26720_ ;
	wire _w26719_ ;
	wire _w26718_ ;
	wire _w26717_ ;
	wire _w26716_ ;
	wire _w26715_ ;
	wire _w26714_ ;
	wire _w26713_ ;
	wire _w26712_ ;
	wire _w26711_ ;
	wire _w26710_ ;
	wire _w26709_ ;
	wire _w26708_ ;
	wire _w26707_ ;
	wire _w26706_ ;
	wire _w26705_ ;
	wire _w26704_ ;
	wire _w26703_ ;
	wire _w26702_ ;
	wire _w26701_ ;
	wire _w26700_ ;
	wire _w26699_ ;
	wire _w26698_ ;
	wire _w26697_ ;
	wire _w26696_ ;
	wire _w26695_ ;
	wire _w26694_ ;
	wire _w26693_ ;
	wire _w26692_ ;
	wire _w26691_ ;
	wire _w26690_ ;
	wire _w26689_ ;
	wire _w26688_ ;
	wire _w26687_ ;
	wire _w26686_ ;
	wire _w26685_ ;
	wire _w26684_ ;
	wire _w26683_ ;
	wire _w26682_ ;
	wire _w26681_ ;
	wire _w26680_ ;
	wire _w26679_ ;
	wire _w26678_ ;
	wire _w26677_ ;
	wire _w26676_ ;
	wire _w26675_ ;
	wire _w26674_ ;
	wire _w26673_ ;
	wire _w26672_ ;
	wire _w26671_ ;
	wire _w26670_ ;
	wire _w26669_ ;
	wire _w26668_ ;
	wire _w26667_ ;
	wire _w26666_ ;
	wire _w26665_ ;
	wire _w26664_ ;
	wire _w26663_ ;
	wire _w26662_ ;
	wire _w26661_ ;
	wire _w26660_ ;
	wire _w26659_ ;
	wire _w26658_ ;
	wire _w26657_ ;
	wire _w26656_ ;
	wire _w26655_ ;
	wire _w26654_ ;
	wire _w26653_ ;
	wire _w26652_ ;
	wire _w26651_ ;
	wire _w26650_ ;
	wire _w26649_ ;
	wire _w26648_ ;
	wire _w26647_ ;
	wire _w26646_ ;
	wire _w26645_ ;
	wire _w26644_ ;
	wire _w26643_ ;
	wire _w26642_ ;
	wire _w26641_ ;
	wire _w26640_ ;
	wire _w26639_ ;
	wire _w26638_ ;
	wire _w26637_ ;
	wire _w26636_ ;
	wire _w26635_ ;
	wire _w26634_ ;
	wire _w26633_ ;
	wire _w26632_ ;
	wire _w26631_ ;
	wire _w26630_ ;
	wire _w26629_ ;
	wire _w26628_ ;
	wire _w26627_ ;
	wire _w26626_ ;
	wire _w26625_ ;
	wire _w26624_ ;
	wire _w26623_ ;
	wire _w26622_ ;
	wire _w26621_ ;
	wire _w26620_ ;
	wire _w26619_ ;
	wire _w26618_ ;
	wire _w26617_ ;
	wire _w26616_ ;
	wire _w26615_ ;
	wire _w26614_ ;
	wire _w26613_ ;
	wire _w26612_ ;
	wire _w26611_ ;
	wire _w26610_ ;
	wire _w26609_ ;
	wire _w26608_ ;
	wire _w26607_ ;
	wire _w26606_ ;
	wire _w26605_ ;
	wire _w26604_ ;
	wire _w26603_ ;
	wire _w26602_ ;
	wire _w26601_ ;
	wire _w26600_ ;
	wire _w26599_ ;
	wire _w26598_ ;
	wire _w26597_ ;
	wire _w26596_ ;
	wire _w26595_ ;
	wire _w26594_ ;
	wire _w26593_ ;
	wire _w26592_ ;
	wire _w26591_ ;
	wire _w26590_ ;
	wire _w26589_ ;
	wire _w26588_ ;
	wire _w26587_ ;
	wire _w26586_ ;
	wire _w26585_ ;
	wire _w26584_ ;
	wire _w26583_ ;
	wire _w26582_ ;
	wire _w26581_ ;
	wire _w26580_ ;
	wire _w26579_ ;
	wire _w26578_ ;
	wire _w26577_ ;
	wire _w26576_ ;
	wire _w26575_ ;
	wire _w26574_ ;
	wire _w26573_ ;
	wire _w26572_ ;
	wire _w26571_ ;
	wire _w26570_ ;
	wire _w26569_ ;
	wire _w26568_ ;
	wire _w26567_ ;
	wire _w26566_ ;
	wire _w26565_ ;
	wire _w26564_ ;
	wire _w26563_ ;
	wire _w26562_ ;
	wire _w26561_ ;
	wire _w26560_ ;
	wire _w26559_ ;
	wire _w26558_ ;
	wire _w26557_ ;
	wire _w26556_ ;
	wire _w26555_ ;
	wire _w26554_ ;
	wire _w26553_ ;
	wire _w26552_ ;
	wire _w26551_ ;
	wire _w26550_ ;
	wire _w26549_ ;
	wire _w26548_ ;
	wire _w26547_ ;
	wire _w26546_ ;
	wire _w26545_ ;
	wire _w26544_ ;
	wire _w26543_ ;
	wire _w26542_ ;
	wire _w26541_ ;
	wire _w26540_ ;
	wire _w26539_ ;
	wire _w26538_ ;
	wire _w26537_ ;
	wire _w26536_ ;
	wire _w26535_ ;
	wire _w26534_ ;
	wire _w26533_ ;
	wire _w26532_ ;
	wire _w26531_ ;
	wire _w26530_ ;
	wire _w26529_ ;
	wire _w26528_ ;
	wire _w26527_ ;
	wire _w26526_ ;
	wire _w26525_ ;
	wire _w26524_ ;
	wire _w26523_ ;
	wire _w26522_ ;
	wire _w26521_ ;
	wire _w26520_ ;
	wire _w26519_ ;
	wire _w26518_ ;
	wire _w26517_ ;
	wire _w26516_ ;
	wire _w26515_ ;
	wire _w26514_ ;
	wire _w26513_ ;
	wire _w26512_ ;
	wire _w26511_ ;
	wire _w26510_ ;
	wire _w26509_ ;
	wire _w26508_ ;
	wire _w26507_ ;
	wire _w26506_ ;
	wire _w26505_ ;
	wire _w26504_ ;
	wire _w26503_ ;
	wire _w26502_ ;
	wire _w26501_ ;
	wire _w26500_ ;
	wire _w26499_ ;
	wire _w26498_ ;
	wire _w26497_ ;
	wire _w26496_ ;
	wire _w26495_ ;
	wire _w26494_ ;
	wire _w26493_ ;
	wire _w26492_ ;
	wire _w26491_ ;
	wire _w26490_ ;
	wire _w26489_ ;
	wire _w26488_ ;
	wire _w26487_ ;
	wire _w26486_ ;
	wire _w26485_ ;
	wire _w26484_ ;
	wire _w26483_ ;
	wire _w26482_ ;
	wire _w26481_ ;
	wire _w26480_ ;
	wire _w26479_ ;
	wire _w26478_ ;
	wire _w26477_ ;
	wire _w26476_ ;
	wire _w26475_ ;
	wire _w26474_ ;
	wire _w26473_ ;
	wire _w26472_ ;
	wire _w26471_ ;
	wire _w26470_ ;
	wire _w26469_ ;
	wire _w26468_ ;
	wire _w26467_ ;
	wire _w26466_ ;
	wire _w26465_ ;
	wire _w26464_ ;
	wire _w26463_ ;
	wire _w26462_ ;
	wire _w26461_ ;
	wire _w26460_ ;
	wire _w26459_ ;
	wire _w26458_ ;
	wire _w26457_ ;
	wire _w26456_ ;
	wire _w26455_ ;
	wire _w26454_ ;
	wire _w26453_ ;
	wire _w26452_ ;
	wire _w26451_ ;
	wire _w26450_ ;
	wire _w26449_ ;
	wire _w26448_ ;
	wire _w26447_ ;
	wire _w26446_ ;
	wire _w26445_ ;
	wire _w26444_ ;
	wire _w26443_ ;
	wire _w26442_ ;
	wire _w26441_ ;
	wire _w26440_ ;
	wire _w26439_ ;
	wire _w26438_ ;
	wire _w26437_ ;
	wire _w26436_ ;
	wire _w26435_ ;
	wire _w26434_ ;
	wire _w26433_ ;
	wire _w26432_ ;
	wire _w26431_ ;
	wire _w26430_ ;
	wire _w26429_ ;
	wire _w26428_ ;
	wire _w26427_ ;
	wire _w26426_ ;
	wire _w26425_ ;
	wire _w26424_ ;
	wire _w26423_ ;
	wire _w26422_ ;
	wire _w26421_ ;
	wire _w26420_ ;
	wire _w26419_ ;
	wire _w26418_ ;
	wire _w26417_ ;
	wire _w26416_ ;
	wire _w26415_ ;
	wire _w26414_ ;
	wire _w26413_ ;
	wire _w26412_ ;
	wire _w26411_ ;
	wire _w26410_ ;
	wire _w26409_ ;
	wire _w26408_ ;
	wire _w26407_ ;
	wire _w26406_ ;
	wire _w26405_ ;
	wire _w26404_ ;
	wire _w26403_ ;
	wire _w26402_ ;
	wire _w26401_ ;
	wire _w26400_ ;
	wire _w26399_ ;
	wire _w26398_ ;
	wire _w26397_ ;
	wire _w26396_ ;
	wire _w26395_ ;
	wire _w26394_ ;
	wire _w26393_ ;
	wire _w26392_ ;
	wire _w26391_ ;
	wire _w26390_ ;
	wire _w26389_ ;
	wire _w26388_ ;
	wire _w26387_ ;
	wire _w26386_ ;
	wire _w26385_ ;
	wire _w26384_ ;
	wire _w26383_ ;
	wire _w26382_ ;
	wire _w26381_ ;
	wire _w26380_ ;
	wire _w26379_ ;
	wire _w26378_ ;
	wire _w26377_ ;
	wire _w26376_ ;
	wire _w26375_ ;
	wire _w26374_ ;
	wire _w26373_ ;
	wire _w26372_ ;
	wire _w26371_ ;
	wire _w26370_ ;
	wire _w26369_ ;
	wire _w26368_ ;
	wire _w26367_ ;
	wire _w26366_ ;
	wire _w26365_ ;
	wire _w26364_ ;
	wire _w26363_ ;
	wire _w26362_ ;
	wire _w26361_ ;
	wire _w26360_ ;
	wire _w26359_ ;
	wire _w26358_ ;
	wire _w26357_ ;
	wire _w26356_ ;
	wire _w26355_ ;
	wire _w26354_ ;
	wire _w26353_ ;
	wire _w26352_ ;
	wire _w26351_ ;
	wire _w26350_ ;
	wire _w26349_ ;
	wire _w26348_ ;
	wire _w26347_ ;
	wire _w26346_ ;
	wire _w26345_ ;
	wire _w26344_ ;
	wire _w26343_ ;
	wire _w26342_ ;
	wire _w26341_ ;
	wire _w26340_ ;
	wire _w26339_ ;
	wire _w26338_ ;
	wire _w26337_ ;
	wire _w26336_ ;
	wire _w26335_ ;
	wire _w26334_ ;
	wire _w26333_ ;
	wire _w26332_ ;
	wire _w26331_ ;
	wire _w26330_ ;
	wire _w26329_ ;
	wire _w26328_ ;
	wire _w26327_ ;
	wire _w26326_ ;
	wire _w26325_ ;
	wire _w26324_ ;
	wire _w26323_ ;
	wire _w26322_ ;
	wire _w26321_ ;
	wire _w26320_ ;
	wire _w26319_ ;
	wire _w26318_ ;
	wire _w26317_ ;
	wire _w26316_ ;
	wire _w26315_ ;
	wire _w26314_ ;
	wire _w26313_ ;
	wire _w26312_ ;
	wire _w26311_ ;
	wire _w26310_ ;
	wire _w26309_ ;
	wire _w26308_ ;
	wire _w26307_ ;
	wire _w26306_ ;
	wire _w26305_ ;
	wire _w26304_ ;
	wire _w26303_ ;
	wire _w26302_ ;
	wire _w26301_ ;
	wire _w26300_ ;
	wire _w26299_ ;
	wire _w26298_ ;
	wire _w26297_ ;
	wire _w26296_ ;
	wire _w26295_ ;
	wire _w26294_ ;
	wire _w26293_ ;
	wire _w26292_ ;
	wire _w26291_ ;
	wire _w26290_ ;
	wire _w26289_ ;
	wire _w26288_ ;
	wire _w26287_ ;
	wire _w26286_ ;
	wire _w26285_ ;
	wire _w26284_ ;
	wire _w26283_ ;
	wire _w26282_ ;
	wire _w26281_ ;
	wire _w26280_ ;
	wire _w26279_ ;
	wire _w26278_ ;
	wire _w26277_ ;
	wire _w26276_ ;
	wire _w26275_ ;
	wire _w26274_ ;
	wire _w26273_ ;
	wire _w26272_ ;
	wire _w26271_ ;
	wire _w26270_ ;
	wire _w26269_ ;
	wire _w26268_ ;
	wire _w26267_ ;
	wire _w26266_ ;
	wire _w26265_ ;
	wire _w26264_ ;
	wire _w26263_ ;
	wire _w26262_ ;
	wire _w26261_ ;
	wire _w26260_ ;
	wire _w26259_ ;
	wire _w26258_ ;
	wire _w26257_ ;
	wire _w26256_ ;
	wire _w26255_ ;
	wire _w26254_ ;
	wire _w26253_ ;
	wire _w26252_ ;
	wire _w26251_ ;
	wire _w26250_ ;
	wire _w26249_ ;
	wire _w26248_ ;
	wire _w26247_ ;
	wire _w26246_ ;
	wire _w26245_ ;
	wire _w26244_ ;
	wire _w26243_ ;
	wire _w26242_ ;
	wire _w26241_ ;
	wire _w26240_ ;
	wire _w26239_ ;
	wire _w26238_ ;
	wire _w26237_ ;
	wire _w26236_ ;
	wire _w26235_ ;
	wire _w26234_ ;
	wire _w26233_ ;
	wire _w26232_ ;
	wire _w26231_ ;
	wire _w26230_ ;
	wire _w26229_ ;
	wire _w26228_ ;
	wire _w26227_ ;
	wire _w26226_ ;
	wire _w26225_ ;
	wire _w26224_ ;
	wire _w26223_ ;
	wire _w26222_ ;
	wire _w26221_ ;
	wire _w26220_ ;
	wire _w26219_ ;
	wire _w26218_ ;
	wire _w26217_ ;
	wire _w26216_ ;
	wire _w26215_ ;
	wire _w26214_ ;
	wire _w26213_ ;
	wire _w26212_ ;
	wire _w26211_ ;
	wire _w26210_ ;
	wire _w26209_ ;
	wire _w26208_ ;
	wire _w26207_ ;
	wire _w26206_ ;
	wire _w26205_ ;
	wire _w26204_ ;
	wire _w26203_ ;
	wire _w26202_ ;
	wire _w26201_ ;
	wire _w26200_ ;
	wire _w26199_ ;
	wire _w26198_ ;
	wire _w26197_ ;
	wire _w26196_ ;
	wire _w26195_ ;
	wire _w26194_ ;
	wire _w26193_ ;
	wire _w26192_ ;
	wire _w26191_ ;
	wire _w26190_ ;
	wire _w26189_ ;
	wire _w26188_ ;
	wire _w26187_ ;
	wire _w26186_ ;
	wire _w26185_ ;
	wire _w26184_ ;
	wire _w26183_ ;
	wire _w26182_ ;
	wire _w26181_ ;
	wire _w26180_ ;
	wire _w26179_ ;
	wire _w26178_ ;
	wire _w26177_ ;
	wire _w26176_ ;
	wire _w26175_ ;
	wire _w26174_ ;
	wire _w26173_ ;
	wire _w26172_ ;
	wire _w26171_ ;
	wire _w26170_ ;
	wire _w26169_ ;
	wire _w26168_ ;
	wire _w26167_ ;
	wire _w26166_ ;
	wire _w26165_ ;
	wire _w26164_ ;
	wire _w26163_ ;
	wire _w26162_ ;
	wire _w26161_ ;
	wire _w26160_ ;
	wire _w26159_ ;
	wire _w26158_ ;
	wire _w26157_ ;
	wire _w26156_ ;
	wire _w26155_ ;
	wire _w26154_ ;
	wire _w26153_ ;
	wire _w26152_ ;
	wire _w26151_ ;
	wire _w26150_ ;
	wire _w26149_ ;
	wire _w26148_ ;
	wire _w26147_ ;
	wire _w26146_ ;
	wire _w26145_ ;
	wire _w26144_ ;
	wire _w26143_ ;
	wire _w26142_ ;
	wire _w26141_ ;
	wire _w26140_ ;
	wire _w26139_ ;
	wire _w26138_ ;
	wire _w26137_ ;
	wire _w26136_ ;
	wire _w26135_ ;
	wire _w26134_ ;
	wire _w26133_ ;
	wire _w26132_ ;
	wire _w26131_ ;
	wire _w26130_ ;
	wire _w26129_ ;
	wire _w26128_ ;
	wire _w26127_ ;
	wire _w26126_ ;
	wire _w26125_ ;
	wire _w26124_ ;
	wire _w26123_ ;
	wire _w26122_ ;
	wire _w26121_ ;
	wire _w26120_ ;
	wire _w26119_ ;
	wire _w26118_ ;
	wire _w26117_ ;
	wire _w26116_ ;
	wire _w26115_ ;
	wire _w26114_ ;
	wire _w26113_ ;
	wire _w26112_ ;
	wire _w26111_ ;
	wire _w26110_ ;
	wire _w26109_ ;
	wire _w26108_ ;
	wire _w26107_ ;
	wire _w26106_ ;
	wire _w26105_ ;
	wire _w26104_ ;
	wire _w26103_ ;
	wire _w26102_ ;
	wire _w26101_ ;
	wire _w26100_ ;
	wire _w26099_ ;
	wire _w26098_ ;
	wire _w26097_ ;
	wire _w26096_ ;
	wire _w26095_ ;
	wire _w26094_ ;
	wire _w26093_ ;
	wire _w26092_ ;
	wire _w26091_ ;
	wire _w26090_ ;
	wire _w26089_ ;
	wire _w26088_ ;
	wire _w26087_ ;
	wire _w26086_ ;
	wire _w26085_ ;
	wire _w26084_ ;
	wire _w26083_ ;
	wire _w26082_ ;
	wire _w26081_ ;
	wire _w26080_ ;
	wire _w26079_ ;
	wire _w26078_ ;
	wire _w26077_ ;
	wire _w26076_ ;
	wire _w26075_ ;
	wire _w26074_ ;
	wire _w26073_ ;
	wire _w26072_ ;
	wire _w26071_ ;
	wire _w26070_ ;
	wire _w26069_ ;
	wire _w26068_ ;
	wire _w26067_ ;
	wire _w26066_ ;
	wire _w26065_ ;
	wire _w26064_ ;
	wire _w26063_ ;
	wire _w26062_ ;
	wire _w26061_ ;
	wire _w26060_ ;
	wire _w26059_ ;
	wire _w26058_ ;
	wire _w26057_ ;
	wire _w26056_ ;
	wire _w26055_ ;
	wire _w26054_ ;
	wire _w26053_ ;
	wire _w26052_ ;
	wire _w26051_ ;
	wire _w26050_ ;
	wire _w26049_ ;
	wire _w26048_ ;
	wire _w26047_ ;
	wire _w26046_ ;
	wire _w26045_ ;
	wire _w26044_ ;
	wire _w26043_ ;
	wire _w26042_ ;
	wire _w26041_ ;
	wire _w26040_ ;
	wire _w26039_ ;
	wire _w26038_ ;
	wire _w26037_ ;
	wire _w26036_ ;
	wire _w26035_ ;
	wire _w26034_ ;
	wire _w26033_ ;
	wire _w26032_ ;
	wire _w26031_ ;
	wire _w26030_ ;
	wire _w26029_ ;
	wire _w26028_ ;
	wire _w26027_ ;
	wire _w26026_ ;
	wire _w26025_ ;
	wire _w26024_ ;
	wire _w26023_ ;
	wire _w26022_ ;
	wire _w26021_ ;
	wire _w26020_ ;
	wire _w26019_ ;
	wire _w26018_ ;
	wire _w26017_ ;
	wire _w26016_ ;
	wire _w26015_ ;
	wire _w26014_ ;
	wire _w26013_ ;
	wire _w26012_ ;
	wire _w26011_ ;
	wire _w26010_ ;
	wire _w26009_ ;
	wire _w26008_ ;
	wire _w26007_ ;
	wire _w26006_ ;
	wire _w26005_ ;
	wire _w26004_ ;
	wire _w26003_ ;
	wire _w26002_ ;
	wire _w26001_ ;
	wire _w26000_ ;
	wire _w25999_ ;
	wire _w25998_ ;
	wire _w25997_ ;
	wire _w25996_ ;
	wire _w25995_ ;
	wire _w25994_ ;
	wire _w25993_ ;
	wire _w25992_ ;
	wire _w25991_ ;
	wire _w25990_ ;
	wire _w25989_ ;
	wire _w25988_ ;
	wire _w25987_ ;
	wire _w25986_ ;
	wire _w25985_ ;
	wire _w25984_ ;
	wire _w25983_ ;
	wire _w25982_ ;
	wire _w25981_ ;
	wire _w25980_ ;
	wire _w25979_ ;
	wire _w25978_ ;
	wire _w25977_ ;
	wire _w25976_ ;
	wire _w25975_ ;
	wire _w25974_ ;
	wire _w25973_ ;
	wire _w25972_ ;
	wire _w25971_ ;
	wire _w25970_ ;
	wire _w25969_ ;
	wire _w25968_ ;
	wire _w25967_ ;
	wire _w25966_ ;
	wire _w25965_ ;
	wire _w25964_ ;
	wire _w25963_ ;
	wire _w25962_ ;
	wire _w25961_ ;
	wire _w25960_ ;
	wire _w25959_ ;
	wire _w25958_ ;
	wire _w25957_ ;
	wire _w25956_ ;
	wire _w25955_ ;
	wire _w25954_ ;
	wire _w25953_ ;
	wire _w25952_ ;
	wire _w25951_ ;
	wire _w25950_ ;
	wire _w25949_ ;
	wire _w25948_ ;
	wire _w25947_ ;
	wire _w25946_ ;
	wire _w25945_ ;
	wire _w25944_ ;
	wire _w25943_ ;
	wire _w25942_ ;
	wire _w25941_ ;
	wire _w25940_ ;
	wire _w25939_ ;
	wire _w25938_ ;
	wire _w25937_ ;
	wire _w25936_ ;
	wire _w25935_ ;
	wire _w25934_ ;
	wire _w25933_ ;
	wire _w25932_ ;
	wire _w25931_ ;
	wire _w25930_ ;
	wire _w25929_ ;
	wire _w25928_ ;
	wire _w25927_ ;
	wire _w25926_ ;
	wire _w25925_ ;
	wire _w25924_ ;
	wire _w25923_ ;
	wire _w25922_ ;
	wire _w25921_ ;
	wire _w25920_ ;
	wire _w25919_ ;
	wire _w25918_ ;
	wire _w25917_ ;
	wire _w25916_ ;
	wire _w25915_ ;
	wire _w25914_ ;
	wire _w25913_ ;
	wire _w25912_ ;
	wire _w25911_ ;
	wire _w25910_ ;
	wire _w25909_ ;
	wire _w25908_ ;
	wire _w25907_ ;
	wire _w25906_ ;
	wire _w25905_ ;
	wire _w25904_ ;
	wire _w25903_ ;
	wire _w25902_ ;
	wire _w25901_ ;
	wire _w25900_ ;
	wire _w25899_ ;
	wire _w25898_ ;
	wire _w25897_ ;
	wire _w25896_ ;
	wire _w25895_ ;
	wire _w25894_ ;
	wire _w25893_ ;
	wire _w25892_ ;
	wire _w25891_ ;
	wire _w25890_ ;
	wire _w25889_ ;
	wire _w25888_ ;
	wire _w25887_ ;
	wire _w25886_ ;
	wire _w25885_ ;
	wire _w25884_ ;
	wire _w25883_ ;
	wire _w25882_ ;
	wire _w25881_ ;
	wire _w25880_ ;
	wire _w25879_ ;
	wire _w25878_ ;
	wire _w25877_ ;
	wire _w25876_ ;
	wire _w25875_ ;
	wire _w25874_ ;
	wire _w25873_ ;
	wire _w25872_ ;
	wire _w25871_ ;
	wire _w25870_ ;
	wire _w25869_ ;
	wire _w25868_ ;
	wire _w25867_ ;
	wire _w25866_ ;
	wire _w25865_ ;
	wire _w25864_ ;
	wire _w25863_ ;
	wire _w25862_ ;
	wire _w25861_ ;
	wire _w25860_ ;
	wire _w25859_ ;
	wire _w25858_ ;
	wire _w25857_ ;
	wire _w25856_ ;
	wire _w25855_ ;
	wire _w25854_ ;
	wire _w25853_ ;
	wire _w25852_ ;
	wire _w25851_ ;
	wire _w25850_ ;
	wire _w25849_ ;
	wire _w25848_ ;
	wire _w25847_ ;
	wire _w25846_ ;
	wire _w25845_ ;
	wire _w25844_ ;
	wire _w25843_ ;
	wire _w25842_ ;
	wire _w25841_ ;
	wire _w25840_ ;
	wire _w25839_ ;
	wire _w25838_ ;
	wire _w25837_ ;
	wire _w25836_ ;
	wire _w25835_ ;
	wire _w25834_ ;
	wire _w25833_ ;
	wire _w25832_ ;
	wire _w25831_ ;
	wire _w25830_ ;
	wire _w25829_ ;
	wire _w25828_ ;
	wire _w25827_ ;
	wire _w25826_ ;
	wire _w25825_ ;
	wire _w25824_ ;
	wire _w25823_ ;
	wire _w25822_ ;
	wire _w25821_ ;
	wire _w25820_ ;
	wire _w25819_ ;
	wire _w25818_ ;
	wire _w25817_ ;
	wire _w25816_ ;
	wire _w25815_ ;
	wire _w25814_ ;
	wire _w25813_ ;
	wire _w25812_ ;
	wire _w25811_ ;
	wire _w25810_ ;
	wire _w25809_ ;
	wire _w25808_ ;
	wire _w25807_ ;
	wire _w25806_ ;
	wire _w25805_ ;
	wire _w25804_ ;
	wire _w25803_ ;
	wire _w25802_ ;
	wire _w25801_ ;
	wire _w25800_ ;
	wire _w25799_ ;
	wire _w25798_ ;
	wire _w25797_ ;
	wire _w25796_ ;
	wire _w25795_ ;
	wire _w25794_ ;
	wire _w25793_ ;
	wire _w25792_ ;
	wire _w25791_ ;
	wire _w25790_ ;
	wire _w25789_ ;
	wire _w25788_ ;
	wire _w25787_ ;
	wire _w25786_ ;
	wire _w25785_ ;
	wire _w25784_ ;
	wire _w25783_ ;
	wire _w25782_ ;
	wire _w25781_ ;
	wire _w25780_ ;
	wire _w25779_ ;
	wire _w25778_ ;
	wire _w25777_ ;
	wire _w25776_ ;
	wire _w25775_ ;
	wire _w25774_ ;
	wire _w25773_ ;
	wire _w25772_ ;
	wire _w25771_ ;
	wire _w25770_ ;
	wire _w25769_ ;
	wire _w25768_ ;
	wire _w25767_ ;
	wire _w25766_ ;
	wire _w25765_ ;
	wire _w25764_ ;
	wire _w25763_ ;
	wire _w25762_ ;
	wire _w25761_ ;
	wire _w25760_ ;
	wire _w25759_ ;
	wire _w25758_ ;
	wire _w25757_ ;
	wire _w25756_ ;
	wire _w25755_ ;
	wire _w25754_ ;
	wire _w25753_ ;
	wire _w25752_ ;
	wire _w25751_ ;
	wire _w25750_ ;
	wire _w25749_ ;
	wire _w25748_ ;
	wire _w25747_ ;
	wire _w25746_ ;
	wire _w25745_ ;
	wire _w25744_ ;
	wire _w25743_ ;
	wire _w25742_ ;
	wire _w25741_ ;
	wire _w25740_ ;
	wire _w25739_ ;
	wire _w25738_ ;
	wire _w25737_ ;
	wire _w25736_ ;
	wire _w25735_ ;
	wire _w25734_ ;
	wire _w25733_ ;
	wire _w25732_ ;
	wire _w25731_ ;
	wire _w25730_ ;
	wire _w25729_ ;
	wire _w25728_ ;
	wire _w25727_ ;
	wire _w25726_ ;
	wire _w25725_ ;
	wire _w25724_ ;
	wire _w25723_ ;
	wire _w25722_ ;
	wire _w25721_ ;
	wire _w25720_ ;
	wire _w25719_ ;
	wire _w25718_ ;
	wire _w25717_ ;
	wire _w25716_ ;
	wire _w25715_ ;
	wire _w25714_ ;
	wire _w25713_ ;
	wire _w25712_ ;
	wire _w25711_ ;
	wire _w25710_ ;
	wire _w25709_ ;
	wire _w25708_ ;
	wire _w25707_ ;
	wire _w25706_ ;
	wire _w25705_ ;
	wire _w25704_ ;
	wire _w25703_ ;
	wire _w25702_ ;
	wire _w25701_ ;
	wire _w25700_ ;
	wire _w25699_ ;
	wire _w25698_ ;
	wire _w25697_ ;
	wire _w25696_ ;
	wire _w25695_ ;
	wire _w25694_ ;
	wire _w25693_ ;
	wire _w25692_ ;
	wire _w25691_ ;
	wire _w25690_ ;
	wire _w25689_ ;
	wire _w25688_ ;
	wire _w25687_ ;
	wire _w25686_ ;
	wire _w25685_ ;
	wire _w25684_ ;
	wire _w25683_ ;
	wire _w25682_ ;
	wire _w25681_ ;
	wire _w25680_ ;
	wire _w25679_ ;
	wire _w25678_ ;
	wire _w25677_ ;
	wire _w25676_ ;
	wire _w25675_ ;
	wire _w25674_ ;
	wire _w25673_ ;
	wire _w25672_ ;
	wire _w25671_ ;
	wire _w25670_ ;
	wire _w25669_ ;
	wire _w25668_ ;
	wire _w25667_ ;
	wire _w25666_ ;
	wire _w25665_ ;
	wire _w25664_ ;
	wire _w25663_ ;
	wire _w25662_ ;
	wire _w25661_ ;
	wire _w25660_ ;
	wire _w25659_ ;
	wire _w25658_ ;
	wire _w25657_ ;
	wire _w25656_ ;
	wire _w25655_ ;
	wire _w25654_ ;
	wire _w25653_ ;
	wire _w25652_ ;
	wire _w25651_ ;
	wire _w25650_ ;
	wire _w25649_ ;
	wire _w25648_ ;
	wire _w25647_ ;
	wire _w25646_ ;
	wire _w25645_ ;
	wire _w25644_ ;
	wire _w25643_ ;
	wire _w25642_ ;
	wire _w25641_ ;
	wire _w25640_ ;
	wire _w25639_ ;
	wire _w25638_ ;
	wire _w25637_ ;
	wire _w25636_ ;
	wire _w25635_ ;
	wire _w25634_ ;
	wire _w25633_ ;
	wire _w25632_ ;
	wire _w25631_ ;
	wire _w25630_ ;
	wire _w25629_ ;
	wire _w25628_ ;
	wire _w25627_ ;
	wire _w25626_ ;
	wire _w25625_ ;
	wire _w25624_ ;
	wire _w25623_ ;
	wire _w25622_ ;
	wire _w25621_ ;
	wire _w25620_ ;
	wire _w25619_ ;
	wire _w25618_ ;
	wire _w25617_ ;
	wire _w25616_ ;
	wire _w25615_ ;
	wire _w25614_ ;
	wire _w25613_ ;
	wire _w25612_ ;
	wire _w25611_ ;
	wire _w25610_ ;
	wire _w25609_ ;
	wire _w25608_ ;
	wire _w25607_ ;
	wire _w25606_ ;
	wire _w25605_ ;
	wire _w25604_ ;
	wire _w25603_ ;
	wire _w25602_ ;
	wire _w25601_ ;
	wire _w25600_ ;
	wire _w25599_ ;
	wire _w25598_ ;
	wire _w25597_ ;
	wire _w25596_ ;
	wire _w25595_ ;
	wire _w25594_ ;
	wire _w25593_ ;
	wire _w25592_ ;
	wire _w25591_ ;
	wire _w25590_ ;
	wire _w25589_ ;
	wire _w25588_ ;
	wire _w25587_ ;
	wire _w25586_ ;
	wire _w25585_ ;
	wire _w25584_ ;
	wire _w25583_ ;
	wire _w25582_ ;
	wire _w25581_ ;
	wire _w25580_ ;
	wire _w25579_ ;
	wire _w25578_ ;
	wire _w25577_ ;
	wire _w25576_ ;
	wire _w25575_ ;
	wire _w25574_ ;
	wire _w25573_ ;
	wire _w25572_ ;
	wire _w25571_ ;
	wire _w25570_ ;
	wire _w25569_ ;
	wire _w25568_ ;
	wire _w25567_ ;
	wire _w25566_ ;
	wire _w25565_ ;
	wire _w25564_ ;
	wire _w25563_ ;
	wire _w25562_ ;
	wire _w25561_ ;
	wire _w25560_ ;
	wire _w25559_ ;
	wire _w25558_ ;
	wire _w25557_ ;
	wire _w25556_ ;
	wire _w25555_ ;
	wire _w25554_ ;
	wire _w25553_ ;
	wire _w25552_ ;
	wire _w25551_ ;
	wire _w25550_ ;
	wire _w25549_ ;
	wire _w25548_ ;
	wire _w25547_ ;
	wire _w25546_ ;
	wire _w25545_ ;
	wire _w25544_ ;
	wire _w25543_ ;
	wire _w25542_ ;
	wire _w25541_ ;
	wire _w25540_ ;
	wire _w25539_ ;
	wire _w25538_ ;
	wire _w25537_ ;
	wire _w25536_ ;
	wire _w25535_ ;
	wire _w25534_ ;
	wire _w25533_ ;
	wire _w25532_ ;
	wire _w25531_ ;
	wire _w25530_ ;
	wire _w25529_ ;
	wire _w25528_ ;
	wire _w25527_ ;
	wire _w25526_ ;
	wire _w25525_ ;
	wire _w25524_ ;
	wire _w25523_ ;
	wire _w25522_ ;
	wire _w25521_ ;
	wire _w25520_ ;
	wire _w25519_ ;
	wire _w25518_ ;
	wire _w25517_ ;
	wire _w25516_ ;
	wire _w25515_ ;
	wire _w25514_ ;
	wire _w25513_ ;
	wire _w25512_ ;
	wire _w25511_ ;
	wire _w25510_ ;
	wire _w25509_ ;
	wire _w25508_ ;
	wire _w25507_ ;
	wire _w25506_ ;
	wire _w25505_ ;
	wire _w25504_ ;
	wire _w25503_ ;
	wire _w25502_ ;
	wire _w25501_ ;
	wire _w25500_ ;
	wire _w25499_ ;
	wire _w25498_ ;
	wire _w25497_ ;
	wire _w25496_ ;
	wire _w25495_ ;
	wire _w25494_ ;
	wire _w25493_ ;
	wire _w25492_ ;
	wire _w25491_ ;
	wire _w25490_ ;
	wire _w25489_ ;
	wire _w25488_ ;
	wire _w25487_ ;
	wire _w25486_ ;
	wire _w25485_ ;
	wire _w25484_ ;
	wire _w25483_ ;
	wire _w25482_ ;
	wire _w25481_ ;
	wire _w25480_ ;
	wire _w25479_ ;
	wire _w25478_ ;
	wire _w25477_ ;
	wire _w25476_ ;
	wire _w25475_ ;
	wire _w25474_ ;
	wire _w25473_ ;
	wire _w25472_ ;
	wire _w25471_ ;
	wire _w25470_ ;
	wire _w25469_ ;
	wire _w25468_ ;
	wire _w25467_ ;
	wire _w25466_ ;
	wire _w25465_ ;
	wire _w25464_ ;
	wire _w25463_ ;
	wire _w25462_ ;
	wire _w25461_ ;
	wire _w25460_ ;
	wire _w25459_ ;
	wire _w25458_ ;
	wire _w25457_ ;
	wire _w25456_ ;
	wire _w25455_ ;
	wire _w25454_ ;
	wire _w25453_ ;
	wire _w25452_ ;
	wire _w25451_ ;
	wire _w25450_ ;
	wire _w25449_ ;
	wire _w25448_ ;
	wire _w25447_ ;
	wire _w25446_ ;
	wire _w25445_ ;
	wire _w25444_ ;
	wire _w25443_ ;
	wire _w25442_ ;
	wire _w25441_ ;
	wire _w25440_ ;
	wire _w25439_ ;
	wire _w25438_ ;
	wire _w25437_ ;
	wire _w25436_ ;
	wire _w25435_ ;
	wire _w25434_ ;
	wire _w25433_ ;
	wire _w25432_ ;
	wire _w25431_ ;
	wire _w25430_ ;
	wire _w25429_ ;
	wire _w25428_ ;
	wire _w25427_ ;
	wire _w25426_ ;
	wire _w25425_ ;
	wire _w25424_ ;
	wire _w25423_ ;
	wire _w25422_ ;
	wire _w25421_ ;
	wire _w25420_ ;
	wire _w25419_ ;
	wire _w25418_ ;
	wire _w25417_ ;
	wire _w25416_ ;
	wire _w25415_ ;
	wire _w25414_ ;
	wire _w25413_ ;
	wire _w25412_ ;
	wire _w25411_ ;
	wire _w25410_ ;
	wire _w25409_ ;
	wire _w25408_ ;
	wire _w25407_ ;
	wire _w25406_ ;
	wire _w25405_ ;
	wire _w25404_ ;
	wire _w25403_ ;
	wire _w25402_ ;
	wire _w25401_ ;
	wire _w25400_ ;
	wire _w25399_ ;
	wire _w25398_ ;
	wire _w25397_ ;
	wire _w25396_ ;
	wire _w25395_ ;
	wire _w25394_ ;
	wire _w25393_ ;
	wire _w25392_ ;
	wire _w25391_ ;
	wire _w25390_ ;
	wire _w25389_ ;
	wire _w25388_ ;
	wire _w25387_ ;
	wire _w25386_ ;
	wire _w25385_ ;
	wire _w25384_ ;
	wire _w25383_ ;
	wire _w25382_ ;
	wire _w25381_ ;
	wire _w25380_ ;
	wire _w25379_ ;
	wire _w25378_ ;
	wire _w25377_ ;
	wire _w25376_ ;
	wire _w25375_ ;
	wire _w25374_ ;
	wire _w25373_ ;
	wire _w25372_ ;
	wire _w25371_ ;
	wire _w25370_ ;
	wire _w25369_ ;
	wire _w25368_ ;
	wire _w25367_ ;
	wire _w25366_ ;
	wire _w25365_ ;
	wire _w25364_ ;
	wire _w25363_ ;
	wire _w25362_ ;
	wire _w25361_ ;
	wire _w25360_ ;
	wire _w25359_ ;
	wire _w25358_ ;
	wire _w25357_ ;
	wire _w25356_ ;
	wire _w25355_ ;
	wire _w25354_ ;
	wire _w25353_ ;
	wire _w25352_ ;
	wire _w25351_ ;
	wire _w25350_ ;
	wire _w25349_ ;
	wire _w25348_ ;
	wire _w25347_ ;
	wire _w25346_ ;
	wire _w25345_ ;
	wire _w25344_ ;
	wire _w25343_ ;
	wire _w25342_ ;
	wire _w25341_ ;
	wire _w25340_ ;
	wire _w25339_ ;
	wire _w25338_ ;
	wire _w25337_ ;
	wire _w25336_ ;
	wire _w25335_ ;
	wire _w25334_ ;
	wire _w25333_ ;
	wire _w25332_ ;
	wire _w25331_ ;
	wire _w25330_ ;
	wire _w25329_ ;
	wire _w25328_ ;
	wire _w25327_ ;
	wire _w25326_ ;
	wire _w25325_ ;
	wire _w25324_ ;
	wire _w25323_ ;
	wire _w25322_ ;
	wire _w25321_ ;
	wire _w25320_ ;
	wire _w25319_ ;
	wire _w25318_ ;
	wire _w25317_ ;
	wire _w25316_ ;
	wire _w25315_ ;
	wire _w25314_ ;
	wire _w25313_ ;
	wire _w25312_ ;
	wire _w25311_ ;
	wire _w25310_ ;
	wire _w25309_ ;
	wire _w25308_ ;
	wire _w25307_ ;
	wire _w25306_ ;
	wire _w25305_ ;
	wire _w25304_ ;
	wire _w25303_ ;
	wire _w25302_ ;
	wire _w25301_ ;
	wire _w25300_ ;
	wire _w25299_ ;
	wire _w25298_ ;
	wire _w25297_ ;
	wire _w25296_ ;
	wire _w25295_ ;
	wire _w25294_ ;
	wire _w25293_ ;
	wire _w25292_ ;
	wire _w25291_ ;
	wire _w25290_ ;
	wire _w25289_ ;
	wire _w25288_ ;
	wire _w25287_ ;
	wire _w25286_ ;
	wire _w25285_ ;
	wire _w25284_ ;
	wire _w25283_ ;
	wire _w25282_ ;
	wire _w25281_ ;
	wire _w25280_ ;
	wire _w25279_ ;
	wire _w25278_ ;
	wire _w25277_ ;
	wire _w25276_ ;
	wire _w25275_ ;
	wire _w25274_ ;
	wire _w25273_ ;
	wire _w25272_ ;
	wire _w25271_ ;
	wire _w25270_ ;
	wire _w25269_ ;
	wire _w25268_ ;
	wire _w25267_ ;
	wire _w25266_ ;
	wire _w25265_ ;
	wire _w25264_ ;
	wire _w25263_ ;
	wire _w25262_ ;
	wire _w25261_ ;
	wire _w25260_ ;
	wire _w25259_ ;
	wire _w25258_ ;
	wire _w25257_ ;
	wire _w25256_ ;
	wire _w25255_ ;
	wire _w25254_ ;
	wire _w25253_ ;
	wire _w25252_ ;
	wire _w25251_ ;
	wire _w25250_ ;
	wire _w25249_ ;
	wire _w25248_ ;
	wire _w25247_ ;
	wire _w25246_ ;
	wire _w25245_ ;
	wire _w25244_ ;
	wire _w25243_ ;
	wire _w25242_ ;
	wire _w25241_ ;
	wire _w25240_ ;
	wire _w25239_ ;
	wire _w25238_ ;
	wire _w25237_ ;
	wire _w25236_ ;
	wire _w25235_ ;
	wire _w25234_ ;
	wire _w25233_ ;
	wire _w25232_ ;
	wire _w25231_ ;
	wire _w25230_ ;
	wire _w25229_ ;
	wire _w25228_ ;
	wire _w25227_ ;
	wire _w25226_ ;
	wire _w25225_ ;
	wire _w25224_ ;
	wire _w25223_ ;
	wire _w25222_ ;
	wire _w25221_ ;
	wire _w25220_ ;
	wire _w25219_ ;
	wire _w25218_ ;
	wire _w25217_ ;
	wire _w25216_ ;
	wire _w25215_ ;
	wire _w25214_ ;
	wire _w25213_ ;
	wire _w25212_ ;
	wire _w25211_ ;
	wire _w25210_ ;
	wire _w25209_ ;
	wire _w25208_ ;
	wire _w25207_ ;
	wire _w25206_ ;
	wire _w25205_ ;
	wire _w25204_ ;
	wire _w25203_ ;
	wire _w25202_ ;
	wire _w25201_ ;
	wire _w25200_ ;
	wire _w25199_ ;
	wire _w25198_ ;
	wire _w25197_ ;
	wire _w25196_ ;
	wire _w25195_ ;
	wire _w25194_ ;
	wire _w25193_ ;
	wire _w25192_ ;
	wire _w25191_ ;
	wire _w25190_ ;
	wire _w25189_ ;
	wire _w25188_ ;
	wire _w25187_ ;
	wire _w25186_ ;
	wire _w25185_ ;
	wire _w25184_ ;
	wire _w25183_ ;
	wire _w25182_ ;
	wire _w25181_ ;
	wire _w25180_ ;
	wire _w25179_ ;
	wire _w25178_ ;
	wire _w25177_ ;
	wire _w25176_ ;
	wire _w25175_ ;
	wire _w25174_ ;
	wire _w25173_ ;
	wire _w25172_ ;
	wire _w25171_ ;
	wire _w25170_ ;
	wire _w25169_ ;
	wire _w25168_ ;
	wire _w25167_ ;
	wire _w25166_ ;
	wire _w25165_ ;
	wire _w25164_ ;
	wire _w25163_ ;
	wire _w25162_ ;
	wire _w25161_ ;
	wire _w25160_ ;
	wire _w25159_ ;
	wire _w25158_ ;
	wire _w25157_ ;
	wire _w25156_ ;
	wire _w25155_ ;
	wire _w25154_ ;
	wire _w25153_ ;
	wire _w25152_ ;
	wire _w25151_ ;
	wire _w25150_ ;
	wire _w25149_ ;
	wire _w25148_ ;
	wire _w25147_ ;
	wire _w25146_ ;
	wire _w25145_ ;
	wire _w25144_ ;
	wire _w25143_ ;
	wire _w25142_ ;
	wire _w25141_ ;
	wire _w25140_ ;
	wire _w25139_ ;
	wire _w25138_ ;
	wire _w25137_ ;
	wire _w25136_ ;
	wire _w25135_ ;
	wire _w25134_ ;
	wire _w25133_ ;
	wire _w25132_ ;
	wire _w25131_ ;
	wire _w25130_ ;
	wire _w25129_ ;
	wire _w25128_ ;
	wire _w25127_ ;
	wire _w25126_ ;
	wire _w25125_ ;
	wire _w25124_ ;
	wire _w25123_ ;
	wire _w25122_ ;
	wire _w25121_ ;
	wire _w25120_ ;
	wire _w25119_ ;
	wire _w25118_ ;
	wire _w25117_ ;
	wire _w25116_ ;
	wire _w25115_ ;
	wire _w25114_ ;
	wire _w25113_ ;
	wire _w25112_ ;
	wire _w25111_ ;
	wire _w25110_ ;
	wire _w25109_ ;
	wire _w25108_ ;
	wire _w25107_ ;
	wire _w25106_ ;
	wire _w25105_ ;
	wire _w25104_ ;
	wire _w25103_ ;
	wire _w25102_ ;
	wire _w25101_ ;
	wire _w25100_ ;
	wire _w25099_ ;
	wire _w25098_ ;
	wire _w25097_ ;
	wire _w25096_ ;
	wire _w25095_ ;
	wire _w25094_ ;
	wire _w25093_ ;
	wire _w25092_ ;
	wire _w25091_ ;
	wire _w25090_ ;
	wire _w25089_ ;
	wire _w25088_ ;
	wire _w25087_ ;
	wire _w25086_ ;
	wire _w25085_ ;
	wire _w25084_ ;
	wire _w25083_ ;
	wire _w25082_ ;
	wire _w25081_ ;
	wire _w25080_ ;
	wire _w25079_ ;
	wire _w25078_ ;
	wire _w25077_ ;
	wire _w25076_ ;
	wire _w25075_ ;
	wire _w25074_ ;
	wire _w25073_ ;
	wire _w25072_ ;
	wire _w25071_ ;
	wire _w25070_ ;
	wire _w25069_ ;
	wire _w25068_ ;
	wire _w25067_ ;
	wire _w25066_ ;
	wire _w25065_ ;
	wire _w25064_ ;
	wire _w25063_ ;
	wire _w25062_ ;
	wire _w25061_ ;
	wire _w25060_ ;
	wire _w25059_ ;
	wire _w25058_ ;
	wire _w25057_ ;
	wire _w25056_ ;
	wire _w25055_ ;
	wire _w25054_ ;
	wire _w25053_ ;
	wire _w25052_ ;
	wire _w25051_ ;
	wire _w25050_ ;
	wire _w25049_ ;
	wire _w25048_ ;
	wire _w25047_ ;
	wire _w25046_ ;
	wire _w25045_ ;
	wire _w25044_ ;
	wire _w25043_ ;
	wire _w25042_ ;
	wire _w25041_ ;
	wire _w25040_ ;
	wire _w25039_ ;
	wire _w25038_ ;
	wire _w25037_ ;
	wire _w25036_ ;
	wire _w25035_ ;
	wire _w25034_ ;
	wire _w25033_ ;
	wire _w25032_ ;
	wire _w25031_ ;
	wire _w25030_ ;
	wire _w25029_ ;
	wire _w25028_ ;
	wire _w25027_ ;
	wire _w25026_ ;
	wire _w25025_ ;
	wire _w25024_ ;
	wire _w25023_ ;
	wire _w25022_ ;
	wire _w25021_ ;
	wire _w25020_ ;
	wire _w25019_ ;
	wire _w25018_ ;
	wire _w25017_ ;
	wire _w25016_ ;
	wire _w25015_ ;
	wire _w25014_ ;
	wire _w25013_ ;
	wire _w25012_ ;
	wire _w25011_ ;
	wire _w25010_ ;
	wire _w25009_ ;
	wire _w25008_ ;
	wire _w25007_ ;
	wire _w25006_ ;
	wire _w25005_ ;
	wire _w25004_ ;
	wire _w25003_ ;
	wire _w25002_ ;
	wire _w25001_ ;
	wire _w25000_ ;
	wire _w24999_ ;
	wire _w24998_ ;
	wire _w24997_ ;
	wire _w24996_ ;
	wire _w24995_ ;
	wire _w24994_ ;
	wire _w24993_ ;
	wire _w24992_ ;
	wire _w24991_ ;
	wire _w24990_ ;
	wire _w24989_ ;
	wire _w24988_ ;
	wire _w24987_ ;
	wire _w24986_ ;
	wire _w24985_ ;
	wire _w24984_ ;
	wire _w24983_ ;
	wire _w24982_ ;
	wire _w24981_ ;
	wire _w24980_ ;
	wire _w24979_ ;
	wire _w24978_ ;
	wire _w24977_ ;
	wire _w24976_ ;
	wire _w24975_ ;
	wire _w24974_ ;
	wire _w24973_ ;
	wire _w24972_ ;
	wire _w24971_ ;
	wire _w24970_ ;
	wire _w24969_ ;
	wire _w24968_ ;
	wire _w24967_ ;
	wire _w24966_ ;
	wire _w24965_ ;
	wire _w24964_ ;
	wire _w24963_ ;
	wire _w24962_ ;
	wire _w24961_ ;
	wire _w24960_ ;
	wire _w24959_ ;
	wire _w24958_ ;
	wire _w24957_ ;
	wire _w24956_ ;
	wire _w24955_ ;
	wire _w24954_ ;
	wire _w24953_ ;
	wire _w24952_ ;
	wire _w24951_ ;
	wire _w24950_ ;
	wire _w24949_ ;
	wire _w24948_ ;
	wire _w24947_ ;
	wire _w24946_ ;
	wire _w24945_ ;
	wire _w24944_ ;
	wire _w24943_ ;
	wire _w24942_ ;
	wire _w24941_ ;
	wire _w24940_ ;
	wire _w24939_ ;
	wire _w24938_ ;
	wire _w24937_ ;
	wire _w24936_ ;
	wire _w24935_ ;
	wire _w24934_ ;
	wire _w24933_ ;
	wire _w24932_ ;
	wire _w24931_ ;
	wire _w24930_ ;
	wire _w24929_ ;
	wire _w24928_ ;
	wire _w24927_ ;
	wire _w24926_ ;
	wire _w24925_ ;
	wire _w24924_ ;
	wire _w24923_ ;
	wire _w24922_ ;
	wire _w24921_ ;
	wire _w24920_ ;
	wire _w24919_ ;
	wire _w24918_ ;
	wire _w24917_ ;
	wire _w24916_ ;
	wire _w24915_ ;
	wire _w24914_ ;
	wire _w24913_ ;
	wire _w24912_ ;
	wire _w24911_ ;
	wire _w24910_ ;
	wire _w24909_ ;
	wire _w24908_ ;
	wire _w24907_ ;
	wire _w24906_ ;
	wire _w24905_ ;
	wire _w24904_ ;
	wire _w24903_ ;
	wire _w24902_ ;
	wire _w24901_ ;
	wire _w24900_ ;
	wire _w24899_ ;
	wire _w24898_ ;
	wire _w24897_ ;
	wire _w24896_ ;
	wire _w24895_ ;
	wire _w24894_ ;
	wire _w24893_ ;
	wire _w24892_ ;
	wire _w24891_ ;
	wire _w24890_ ;
	wire _w24889_ ;
	wire _w24888_ ;
	wire _w24887_ ;
	wire _w24886_ ;
	wire _w24885_ ;
	wire _w24884_ ;
	wire _w24883_ ;
	wire _w24882_ ;
	wire _w24881_ ;
	wire _w24880_ ;
	wire _w24879_ ;
	wire _w24878_ ;
	wire _w24877_ ;
	wire _w24876_ ;
	wire _w24875_ ;
	wire _w24874_ ;
	wire _w24873_ ;
	wire _w24872_ ;
	wire _w24871_ ;
	wire _w24870_ ;
	wire _w24869_ ;
	wire _w24868_ ;
	wire _w24867_ ;
	wire _w24866_ ;
	wire _w24865_ ;
	wire _w24864_ ;
	wire _w24863_ ;
	wire _w24862_ ;
	wire _w24861_ ;
	wire _w24860_ ;
	wire _w24859_ ;
	wire _w24858_ ;
	wire _w24857_ ;
	wire _w24856_ ;
	wire _w24855_ ;
	wire _w24854_ ;
	wire _w24853_ ;
	wire _w24852_ ;
	wire _w24851_ ;
	wire _w24850_ ;
	wire _w24849_ ;
	wire _w24848_ ;
	wire _w24847_ ;
	wire _w24846_ ;
	wire _w24845_ ;
	wire _w24844_ ;
	wire _w24843_ ;
	wire _w24842_ ;
	wire _w24841_ ;
	wire _w24840_ ;
	wire _w24839_ ;
	wire _w24838_ ;
	wire _w24837_ ;
	wire _w24836_ ;
	wire _w24835_ ;
	wire _w24834_ ;
	wire _w24833_ ;
	wire _w24832_ ;
	wire _w24831_ ;
	wire _w24830_ ;
	wire _w24829_ ;
	wire _w24828_ ;
	wire _w24827_ ;
	wire _w24826_ ;
	wire _w24825_ ;
	wire _w24824_ ;
	wire _w24823_ ;
	wire _w24822_ ;
	wire _w24821_ ;
	wire _w24820_ ;
	wire _w24819_ ;
	wire _w24818_ ;
	wire _w24817_ ;
	wire _w24816_ ;
	wire _w24815_ ;
	wire _w24814_ ;
	wire _w24813_ ;
	wire _w24812_ ;
	wire _w24811_ ;
	wire _w24810_ ;
	wire _w24809_ ;
	wire _w24808_ ;
	wire _w24807_ ;
	wire _w24806_ ;
	wire _w24805_ ;
	wire _w24804_ ;
	wire _w24803_ ;
	wire _w24802_ ;
	wire _w24801_ ;
	wire _w24800_ ;
	wire _w14319_ ;
	wire _w14318_ ;
	wire _w14317_ ;
	wire _w14316_ ;
	wire _w14315_ ;
	wire _w14314_ ;
	wire _w14313_ ;
	wire _w14312_ ;
	wire _w14311_ ;
	wire _w14310_ ;
	wire _w14309_ ;
	wire _w14308_ ;
	wire _w14307_ ;
	wire _w14306_ ;
	wire _w14305_ ;
	wire _w14304_ ;
	wire _w14303_ ;
	wire _w14302_ ;
	wire _w14301_ ;
	wire _w14300_ ;
	wire _w14299_ ;
	wire _w14298_ ;
	wire _w14297_ ;
	wire _w14296_ ;
	wire _w14295_ ;
	wire _w14294_ ;
	wire _w14293_ ;
	wire _w14292_ ;
	wire _w14291_ ;
	wire _w14290_ ;
	wire _w14289_ ;
	wire _w14288_ ;
	wire _w14287_ ;
	wire _w14286_ ;
	wire _w14285_ ;
	wire _w14284_ ;
	wire _w14283_ ;
	wire _w14282_ ;
	wire _w14281_ ;
	wire _w14280_ ;
	wire _w14279_ ;
	wire _w14278_ ;
	wire _w14277_ ;
	wire _w14276_ ;
	wire _w14275_ ;
	wire _w14274_ ;
	wire _w14273_ ;
	wire _w14272_ ;
	wire _w14271_ ;
	wire _w14270_ ;
	wire _w14269_ ;
	wire _w14268_ ;
	wire _w14267_ ;
	wire _w14266_ ;
	wire _w14265_ ;
	wire _w14264_ ;
	wire _w14263_ ;
	wire _w14262_ ;
	wire _w14261_ ;
	wire _w14260_ ;
	wire _w14259_ ;
	wire _w14258_ ;
	wire _w14257_ ;
	wire _w14256_ ;
	wire _w14255_ ;
	wire _w14254_ ;
	wire _w14253_ ;
	wire _w14252_ ;
	wire _w14251_ ;
	wire _w14250_ ;
	wire _w14249_ ;
	wire _w14248_ ;
	wire _w14247_ ;
	wire _w14246_ ;
	wire _w14245_ ;
	wire _w14244_ ;
	wire _w14243_ ;
	wire _w14242_ ;
	wire _w14241_ ;
	wire _w14240_ ;
	wire _w14239_ ;
	wire _w14238_ ;
	wire _w14237_ ;
	wire _w14236_ ;
	wire _w14235_ ;
	wire _w14234_ ;
	wire _w14233_ ;
	wire _w14232_ ;
	wire _w14231_ ;
	wire _w14230_ ;
	wire _w14229_ ;
	wire _w14228_ ;
	wire _w14227_ ;
	wire _w14226_ ;
	wire _w14225_ ;
	wire _w14224_ ;
	wire _w14223_ ;
	wire _w14222_ ;
	wire _w14221_ ;
	wire _w14220_ ;
	wire _w14219_ ;
	wire _w14218_ ;
	wire _w14217_ ;
	wire _w14216_ ;
	wire _w14215_ ;
	wire _w14214_ ;
	wire _w14213_ ;
	wire _w14212_ ;
	wire _w14211_ ;
	wire _w14210_ ;
	wire _w14209_ ;
	wire _w14208_ ;
	wire _w14207_ ;
	wire _w14206_ ;
	wire _w14205_ ;
	wire _w14204_ ;
	wire _w14203_ ;
	wire _w14202_ ;
	wire _w14201_ ;
	wire _w14200_ ;
	wire _w14199_ ;
	wire _w14198_ ;
	wire _w14197_ ;
	wire _w14196_ ;
	wire _w14195_ ;
	wire _w14194_ ;
	wire _w14193_ ;
	wire _w14192_ ;
	wire _w14191_ ;
	wire _w14190_ ;
	wire _w14189_ ;
	wire _w14188_ ;
	wire _w14187_ ;
	wire _w14186_ ;
	wire _w14185_ ;
	wire _w14184_ ;
	wire _w14183_ ;
	wire _w14182_ ;
	wire _w14181_ ;
	wire _w14180_ ;
	wire _w14179_ ;
	wire _w14178_ ;
	wire _w14177_ ;
	wire _w14176_ ;
	wire _w14175_ ;
	wire _w14174_ ;
	wire _w14173_ ;
	wire _w14172_ ;
	wire _w14171_ ;
	wire _w14170_ ;
	wire _w14169_ ;
	wire _w14168_ ;
	wire _w14167_ ;
	wire _w14166_ ;
	wire _w14165_ ;
	wire _w14164_ ;
	wire _w14163_ ;
	wire _w14162_ ;
	wire _w14161_ ;
	wire _w14160_ ;
	wire _w14159_ ;
	wire _w14158_ ;
	wire _w14157_ ;
	wire _w14156_ ;
	wire _w14155_ ;
	wire _w14154_ ;
	wire _w14153_ ;
	wire _w14152_ ;
	wire _w14151_ ;
	wire _w14150_ ;
	wire _w14149_ ;
	wire _w14148_ ;
	wire _w14147_ ;
	wire _w14146_ ;
	wire _w14145_ ;
	wire _w14144_ ;
	wire _w14143_ ;
	wire _w14142_ ;
	wire _w14141_ ;
	wire _w14140_ ;
	wire _w14139_ ;
	wire _w14138_ ;
	wire _w14137_ ;
	wire _w14136_ ;
	wire _w14135_ ;
	wire _w14134_ ;
	wire _w14133_ ;
	wire _w14132_ ;
	wire _w14131_ ;
	wire _w14130_ ;
	wire _w14129_ ;
	wire _w14128_ ;
	wire _w14127_ ;
	wire _w14126_ ;
	wire _w14125_ ;
	wire _w14124_ ;
	wire _w14123_ ;
	wire _w14122_ ;
	wire _w14121_ ;
	wire _w14120_ ;
	wire _w14119_ ;
	wire _w14118_ ;
	wire _w14117_ ;
	wire _w14116_ ;
	wire _w14115_ ;
	wire _w14114_ ;
	wire _w14113_ ;
	wire _w14112_ ;
	wire _w14111_ ;
	wire _w14110_ ;
	wire _w14109_ ;
	wire _w14108_ ;
	wire _w14107_ ;
	wire _w14106_ ;
	wire _w14105_ ;
	wire _w14104_ ;
	wire _w14103_ ;
	wire _w14102_ ;
	wire _w14101_ ;
	wire _w14100_ ;
	wire _w14099_ ;
	wire _w14098_ ;
	wire _w14097_ ;
	wire _w14096_ ;
	wire _w14095_ ;
	wire _w14094_ ;
	wire _w14093_ ;
	wire _w14092_ ;
	wire _w14091_ ;
	wire _w14090_ ;
	wire _w14089_ ;
	wire _w14088_ ;
	wire _w14087_ ;
	wire _w14086_ ;
	wire _w14085_ ;
	wire _w14084_ ;
	wire _w14083_ ;
	wire _w14082_ ;
	wire _w14081_ ;
	wire _w14080_ ;
	wire _w14079_ ;
	wire _w14078_ ;
	wire _w14077_ ;
	wire _w14076_ ;
	wire _w14075_ ;
	wire _w14074_ ;
	wire _w14073_ ;
	wire _w14072_ ;
	wire _w14071_ ;
	wire _w14070_ ;
	wire _w14069_ ;
	wire _w14068_ ;
	wire _w14067_ ;
	wire _w14066_ ;
	wire _w14065_ ;
	wire _w14064_ ;
	wire _w14063_ ;
	wire _w14062_ ;
	wire _w14061_ ;
	wire _w14060_ ;
	wire _w14059_ ;
	wire _w14058_ ;
	wire _w14057_ ;
	wire _w14056_ ;
	wire _w14055_ ;
	wire _w14054_ ;
	wire _w14053_ ;
	wire _w14052_ ;
	wire _w14051_ ;
	wire _w14050_ ;
	wire _w14049_ ;
	wire _w14048_ ;
	wire _w14047_ ;
	wire _w14046_ ;
	wire _w14045_ ;
	wire _w14044_ ;
	wire _w14043_ ;
	wire _w14042_ ;
	wire _w14041_ ;
	wire _w14040_ ;
	wire _w14039_ ;
	wire _w14038_ ;
	wire _w14037_ ;
	wire _w14036_ ;
	wire _w14035_ ;
	wire _w14034_ ;
	wire _w14033_ ;
	wire _w14032_ ;
	wire _w14031_ ;
	wire _w14030_ ;
	wire _w14029_ ;
	wire _w14028_ ;
	wire _w14027_ ;
	wire _w14026_ ;
	wire _w14025_ ;
	wire _w14024_ ;
	wire _w14023_ ;
	wire _w14022_ ;
	wire _w14021_ ;
	wire _w14020_ ;
	wire _w14019_ ;
	wire _w14018_ ;
	wire _w14017_ ;
	wire _w14016_ ;
	wire _w14015_ ;
	wire _w14014_ ;
	wire _w14013_ ;
	wire _w14012_ ;
	wire _w14011_ ;
	wire _w14010_ ;
	wire _w14009_ ;
	wire _w14008_ ;
	wire _w14007_ ;
	wire _w14006_ ;
	wire _w14005_ ;
	wire _w14004_ ;
	wire _w14003_ ;
	wire _w14002_ ;
	wire _w14001_ ;
	wire _w14000_ ;
	wire _w13999_ ;
	wire _w13998_ ;
	wire _w13997_ ;
	wire _w13996_ ;
	wire _w13995_ ;
	wire _w13994_ ;
	wire _w13993_ ;
	wire _w13992_ ;
	wire _w13991_ ;
	wire _w13990_ ;
	wire _w13989_ ;
	wire _w13988_ ;
	wire _w13987_ ;
	wire _w13986_ ;
	wire _w13985_ ;
	wire _w13984_ ;
	wire _w13983_ ;
	wire _w13982_ ;
	wire _w13981_ ;
	wire _w13980_ ;
	wire _w13979_ ;
	wire _w13978_ ;
	wire _w13977_ ;
	wire _w13976_ ;
	wire _w13975_ ;
	wire _w13974_ ;
	wire _w13973_ ;
	wire _w13972_ ;
	wire _w13971_ ;
	wire _w13970_ ;
	wire _w13969_ ;
	wire _w13968_ ;
	wire _w13967_ ;
	wire _w13966_ ;
	wire _w13965_ ;
	wire _w13964_ ;
	wire _w13963_ ;
	wire _w13962_ ;
	wire _w13961_ ;
	wire _w13960_ ;
	wire _w13959_ ;
	wire _w13958_ ;
	wire _w13957_ ;
	wire _w13956_ ;
	wire _w13955_ ;
	wire _w13954_ ;
	wire _w13953_ ;
	wire _w13952_ ;
	wire _w13951_ ;
	wire _w13950_ ;
	wire _w13949_ ;
	wire _w13948_ ;
	wire _w13947_ ;
	wire _w13946_ ;
	wire _w13945_ ;
	wire _w13944_ ;
	wire _w13943_ ;
	wire _w13942_ ;
	wire _w13941_ ;
	wire _w13940_ ;
	wire _w13939_ ;
	wire _w13938_ ;
	wire _w13937_ ;
	wire _w13936_ ;
	wire _w13935_ ;
	wire _w13934_ ;
	wire _w13933_ ;
	wire _w13932_ ;
	wire _w13931_ ;
	wire _w13930_ ;
	wire _w13929_ ;
	wire _w13928_ ;
	wire _w13927_ ;
	wire _w13926_ ;
	wire _w13925_ ;
	wire _w13924_ ;
	wire _w13923_ ;
	wire _w13922_ ;
	wire _w13921_ ;
	wire _w13920_ ;
	wire _w13919_ ;
	wire _w13918_ ;
	wire _w13917_ ;
	wire _w13916_ ;
	wire _w13915_ ;
	wire _w13914_ ;
	wire _w13913_ ;
	wire _w13912_ ;
	wire _w13911_ ;
	wire _w13910_ ;
	wire _w13909_ ;
	wire _w13908_ ;
	wire _w13907_ ;
	wire _w13906_ ;
	wire _w13905_ ;
	wire _w13904_ ;
	wire _w13903_ ;
	wire _w13902_ ;
	wire _w13901_ ;
	wire _w13900_ ;
	wire _w13899_ ;
	wire _w13898_ ;
	wire _w13897_ ;
	wire _w13896_ ;
	wire _w13895_ ;
	wire _w13894_ ;
	wire _w13893_ ;
	wire _w13892_ ;
	wire _w13891_ ;
	wire _w13890_ ;
	wire _w13889_ ;
	wire _w13888_ ;
	wire _w13887_ ;
	wire _w13886_ ;
	wire _w13885_ ;
	wire _w13884_ ;
	wire _w13883_ ;
	wire _w13882_ ;
	wire _w13881_ ;
	wire _w13880_ ;
	wire _w13879_ ;
	wire _w13878_ ;
	wire _w13877_ ;
	wire _w13876_ ;
	wire _w13875_ ;
	wire _w13874_ ;
	wire _w13873_ ;
	wire _w13872_ ;
	wire _w13871_ ;
	wire _w13870_ ;
	wire _w13869_ ;
	wire _w13868_ ;
	wire _w13867_ ;
	wire _w13866_ ;
	wire _w13865_ ;
	wire _w13864_ ;
	wire _w13863_ ;
	wire _w13862_ ;
	wire _w13861_ ;
	wire _w13860_ ;
	wire _w13859_ ;
	wire _w13858_ ;
	wire _w13857_ ;
	wire _w13856_ ;
	wire _w13855_ ;
	wire _w13854_ ;
	wire _w13853_ ;
	wire _w13852_ ;
	wire _w13851_ ;
	wire _w13850_ ;
	wire _w13849_ ;
	wire _w13848_ ;
	wire _w13847_ ;
	wire _w13846_ ;
	wire _w13845_ ;
	wire _w13844_ ;
	wire _w13843_ ;
	wire _w13842_ ;
	wire _w13841_ ;
	wire _w13840_ ;
	wire _w13839_ ;
	wire _w13838_ ;
	wire _w13837_ ;
	wire _w13836_ ;
	wire _w13835_ ;
	wire _w13834_ ;
	wire _w13833_ ;
	wire _w13832_ ;
	wire _w13831_ ;
	wire _w13830_ ;
	wire _w13829_ ;
	wire _w13828_ ;
	wire _w13827_ ;
	wire _w13826_ ;
	wire _w13825_ ;
	wire _w13824_ ;
	wire _w13823_ ;
	wire _w13822_ ;
	wire _w13821_ ;
	wire _w13820_ ;
	wire _w13819_ ;
	wire _w13818_ ;
	wire _w13817_ ;
	wire _w13816_ ;
	wire _w13815_ ;
	wire _w13814_ ;
	wire _w13813_ ;
	wire _w13812_ ;
	wire _w13811_ ;
	wire _w13810_ ;
	wire _w13809_ ;
	wire _w13808_ ;
	wire _w13807_ ;
	wire _w13806_ ;
	wire _w13805_ ;
	wire _w13804_ ;
	wire _w13803_ ;
	wire _w13802_ ;
	wire _w13801_ ;
	wire _w13800_ ;
	wire _w13799_ ;
	wire _w13798_ ;
	wire _w13797_ ;
	wire _w13796_ ;
	wire _w13795_ ;
	wire _w13794_ ;
	wire _w13793_ ;
	wire _w13792_ ;
	wire _w13791_ ;
	wire _w13790_ ;
	wire _w13789_ ;
	wire _w13788_ ;
	wire _w13787_ ;
	wire _w13786_ ;
	wire _w13785_ ;
	wire _w13784_ ;
	wire _w13783_ ;
	wire _w13782_ ;
	wire _w13781_ ;
	wire _w13780_ ;
	wire _w13779_ ;
	wire _w13778_ ;
	wire _w13777_ ;
	wire _w13776_ ;
	wire _w13775_ ;
	wire _w13774_ ;
	wire _w13773_ ;
	wire _w13772_ ;
	wire _w13771_ ;
	wire _w13770_ ;
	wire _w13769_ ;
	wire _w13768_ ;
	wire _w13767_ ;
	wire _w13766_ ;
	wire _w13765_ ;
	wire _w13764_ ;
	wire _w13763_ ;
	wire _w13762_ ;
	wire _w13761_ ;
	wire _w13760_ ;
	wire _w13759_ ;
	wire _w13758_ ;
	wire _w13757_ ;
	wire _w13756_ ;
	wire _w13755_ ;
	wire _w13754_ ;
	wire _w13753_ ;
	wire _w13752_ ;
	wire _w13751_ ;
	wire _w13750_ ;
	wire _w13749_ ;
	wire _w13748_ ;
	wire _w13747_ ;
	wire _w13746_ ;
	wire _w13745_ ;
	wire _w13744_ ;
	wire _w13743_ ;
	wire _w13742_ ;
	wire _w13741_ ;
	wire _w13740_ ;
	wire _w13739_ ;
	wire _w13738_ ;
	wire _w13737_ ;
	wire _w13736_ ;
	wire _w13735_ ;
	wire _w13734_ ;
	wire _w13733_ ;
	wire _w13732_ ;
	wire _w13731_ ;
	wire _w13730_ ;
	wire _w13729_ ;
	wire _w13728_ ;
	wire _w13727_ ;
	wire _w13726_ ;
	wire _w13725_ ;
	wire _w13724_ ;
	wire _w13723_ ;
	wire _w13722_ ;
	wire _w13721_ ;
	wire _w13720_ ;
	wire _w13719_ ;
	wire _w13718_ ;
	wire _w13717_ ;
	wire _w13716_ ;
	wire _w13715_ ;
	wire _w13714_ ;
	wire _w13713_ ;
	wire _w13712_ ;
	wire _w13711_ ;
	wire _w13710_ ;
	wire _w13709_ ;
	wire _w13708_ ;
	wire _w13707_ ;
	wire _w13706_ ;
	wire _w13705_ ;
	wire _w13704_ ;
	wire _w13703_ ;
	wire _w13702_ ;
	wire _w13701_ ;
	wire _w13700_ ;
	wire _w13699_ ;
	wire _w13698_ ;
	wire _w13697_ ;
	wire _w13696_ ;
	wire _w13695_ ;
	wire _w13694_ ;
	wire _w13693_ ;
	wire _w13692_ ;
	wire _w13691_ ;
	wire _w13690_ ;
	wire _w13689_ ;
	wire _w13688_ ;
	wire _w13687_ ;
	wire _w13686_ ;
	wire _w13685_ ;
	wire _w13684_ ;
	wire _w13683_ ;
	wire _w13682_ ;
	wire _w13681_ ;
	wire _w13680_ ;
	wire _w13679_ ;
	wire _w13678_ ;
	wire _w13677_ ;
	wire _w13676_ ;
	wire _w13675_ ;
	wire _w13674_ ;
	wire _w13673_ ;
	wire _w13672_ ;
	wire _w13671_ ;
	wire _w13670_ ;
	wire _w13669_ ;
	wire _w13668_ ;
	wire _w13667_ ;
	wire _w13666_ ;
	wire _w13665_ ;
	wire _w13664_ ;
	wire _w13663_ ;
	wire _w13662_ ;
	wire _w13661_ ;
	wire _w13660_ ;
	wire _w13659_ ;
	wire _w13658_ ;
	wire _w13657_ ;
	wire _w13656_ ;
	wire _w13655_ ;
	wire _w13654_ ;
	wire _w13653_ ;
	wire _w13652_ ;
	wire _w13651_ ;
	wire _w13650_ ;
	wire _w13649_ ;
	wire _w13648_ ;
	wire _w13647_ ;
	wire _w13646_ ;
	wire _w13645_ ;
	wire _w13644_ ;
	wire _w13643_ ;
	wire _w13642_ ;
	wire _w13641_ ;
	wire _w13640_ ;
	wire _w13639_ ;
	wire _w13638_ ;
	wire _w13637_ ;
	wire _w13636_ ;
	wire _w13635_ ;
	wire _w13634_ ;
	wire _w13633_ ;
	wire _w13632_ ;
	wire _w13631_ ;
	wire _w13630_ ;
	wire _w13629_ ;
	wire _w13628_ ;
	wire _w13627_ ;
	wire _w13626_ ;
	wire _w13625_ ;
	wire _w13624_ ;
	wire _w13623_ ;
	wire _w13622_ ;
	wire _w13621_ ;
	wire _w13620_ ;
	wire _w13619_ ;
	wire _w13618_ ;
	wire _w13617_ ;
	wire _w13616_ ;
	wire _w13615_ ;
	wire _w13614_ ;
	wire _w13613_ ;
	wire _w13612_ ;
	wire _w13611_ ;
	wire _w13610_ ;
	wire _w13609_ ;
	wire _w13608_ ;
	wire _w13607_ ;
	wire _w13606_ ;
	wire _w13605_ ;
	wire _w13604_ ;
	wire _w13603_ ;
	wire _w13602_ ;
	wire _w13601_ ;
	wire _w13600_ ;
	wire _w13599_ ;
	wire _w13598_ ;
	wire _w13597_ ;
	wire _w13596_ ;
	wire _w13595_ ;
	wire _w13594_ ;
	wire _w13593_ ;
	wire _w13592_ ;
	wire _w13591_ ;
	wire _w13590_ ;
	wire _w13589_ ;
	wire _w13588_ ;
	wire _w13587_ ;
	wire _w13586_ ;
	wire _w13585_ ;
	wire _w13584_ ;
	wire _w13583_ ;
	wire _w13582_ ;
	wire _w13581_ ;
	wire _w13580_ ;
	wire _w13579_ ;
	wire _w13578_ ;
	wire _w13577_ ;
	wire _w13576_ ;
	wire _w13575_ ;
	wire _w13574_ ;
	wire _w13573_ ;
	wire _w13572_ ;
	wire _w13571_ ;
	wire _w13570_ ;
	wire _w13569_ ;
	wire _w13568_ ;
	wire _w13567_ ;
	wire _w13566_ ;
	wire _w13565_ ;
	wire _w13564_ ;
	wire _w13563_ ;
	wire _w13562_ ;
	wire _w13561_ ;
	wire _w13560_ ;
	wire _w13559_ ;
	wire _w13558_ ;
	wire _w13557_ ;
	wire _w13556_ ;
	wire _w13555_ ;
	wire _w13554_ ;
	wire _w13553_ ;
	wire _w13552_ ;
	wire _w13551_ ;
	wire _w13550_ ;
	wire _w13549_ ;
	wire _w13548_ ;
	wire _w13547_ ;
	wire _w13546_ ;
	wire _w13545_ ;
	wire _w13544_ ;
	wire _w13543_ ;
	wire _w13542_ ;
	wire _w13541_ ;
	wire _w13540_ ;
	wire _w13539_ ;
	wire _w13538_ ;
	wire _w13537_ ;
	wire _w13536_ ;
	wire _w13535_ ;
	wire _w13534_ ;
	wire _w13533_ ;
	wire _w13532_ ;
	wire _w13531_ ;
	wire _w13530_ ;
	wire _w13529_ ;
	wire _w13528_ ;
	wire _w13527_ ;
	wire _w13526_ ;
	wire _w13525_ ;
	wire _w13524_ ;
	wire _w13523_ ;
	wire _w13522_ ;
	wire _w13521_ ;
	wire _w13520_ ;
	wire _w13519_ ;
	wire _w13518_ ;
	wire _w13517_ ;
	wire _w13516_ ;
	wire _w13515_ ;
	wire _w13514_ ;
	wire _w13513_ ;
	wire _w13512_ ;
	wire _w13511_ ;
	wire _w13510_ ;
	wire _w13509_ ;
	wire _w13508_ ;
	wire _w13507_ ;
	wire _w13506_ ;
	wire _w13505_ ;
	wire _w13504_ ;
	wire _w13503_ ;
	wire _w13502_ ;
	wire _w13501_ ;
	wire _w13500_ ;
	wire _w13499_ ;
	wire _w13498_ ;
	wire _w13497_ ;
	wire _w13496_ ;
	wire _w13495_ ;
	wire _w13494_ ;
	wire _w13493_ ;
	wire _w13492_ ;
	wire _w13491_ ;
	wire _w13490_ ;
	wire _w13489_ ;
	wire _w13488_ ;
	wire _w13487_ ;
	wire _w13486_ ;
	wire _w13485_ ;
	wire _w13484_ ;
	wire _w13483_ ;
	wire _w13482_ ;
	wire _w13481_ ;
	wire _w13480_ ;
	wire _w13479_ ;
	wire _w13478_ ;
	wire _w13477_ ;
	wire _w13476_ ;
	wire _w13475_ ;
	wire _w13474_ ;
	wire _w13473_ ;
	wire _w13472_ ;
	wire _w13471_ ;
	wire _w13470_ ;
	wire _w13469_ ;
	wire _w13468_ ;
	wire _w13467_ ;
	wire _w13466_ ;
	wire _w13465_ ;
	wire _w13464_ ;
	wire _w13463_ ;
	wire _w13462_ ;
	wire _w13461_ ;
	wire _w13460_ ;
	wire _w13459_ ;
	wire _w13458_ ;
	wire _w13457_ ;
	wire _w13456_ ;
	wire _w13455_ ;
	wire _w13454_ ;
	wire _w13453_ ;
	wire _w13452_ ;
	wire _w13451_ ;
	wire _w13450_ ;
	wire _w13449_ ;
	wire _w13448_ ;
	wire _w13447_ ;
	wire _w13446_ ;
	wire _w13445_ ;
	wire _w13444_ ;
	wire _w13443_ ;
	wire _w13442_ ;
	wire _w13441_ ;
	wire _w13440_ ;
	wire _w13439_ ;
	wire _w13438_ ;
	wire _w13437_ ;
	wire _w13436_ ;
	wire _w13435_ ;
	wire _w13434_ ;
	wire _w13433_ ;
	wire _w13432_ ;
	wire _w13431_ ;
	wire _w13430_ ;
	wire _w13429_ ;
	wire _w13428_ ;
	wire _w13427_ ;
	wire _w13426_ ;
	wire _w13425_ ;
	wire _w13424_ ;
	wire _w13423_ ;
	wire _w13422_ ;
	wire _w13421_ ;
	wire _w13420_ ;
	wire _w13419_ ;
	wire _w13418_ ;
	wire _w13417_ ;
	wire _w13416_ ;
	wire _w13415_ ;
	wire _w13414_ ;
	wire _w13413_ ;
	wire _w13412_ ;
	wire _w13411_ ;
	wire _w13410_ ;
	wire _w13409_ ;
	wire _w13408_ ;
	wire _w13407_ ;
	wire _w13406_ ;
	wire _w13405_ ;
	wire _w13404_ ;
	wire _w13403_ ;
	wire _w13402_ ;
	wire _w13401_ ;
	wire _w13400_ ;
	wire _w13399_ ;
	wire _w13398_ ;
	wire _w13397_ ;
	wire _w13396_ ;
	wire _w13395_ ;
	wire _w13394_ ;
	wire _w13393_ ;
	wire _w13392_ ;
	wire _w13391_ ;
	wire _w13390_ ;
	wire _w13389_ ;
	wire _w13388_ ;
	wire _w13387_ ;
	wire _w13386_ ;
	wire _w13385_ ;
	wire _w13384_ ;
	wire _w13383_ ;
	wire _w13382_ ;
	wire _w13381_ ;
	wire _w13380_ ;
	wire _w13379_ ;
	wire _w13378_ ;
	wire _w13377_ ;
	wire _w13376_ ;
	wire _w13375_ ;
	wire _w13374_ ;
	wire _w13373_ ;
	wire _w13372_ ;
	wire _w13371_ ;
	wire _w13370_ ;
	wire _w13369_ ;
	wire _w13368_ ;
	wire _w13367_ ;
	wire _w13366_ ;
	wire _w13365_ ;
	wire _w13364_ ;
	wire _w13363_ ;
	wire _w13362_ ;
	wire _w13361_ ;
	wire _w13360_ ;
	wire _w13359_ ;
	wire _w13358_ ;
	wire _w13357_ ;
	wire _w13356_ ;
	wire _w13355_ ;
	wire _w13354_ ;
	wire _w13353_ ;
	wire _w13352_ ;
	wire _w13351_ ;
	wire _w13350_ ;
	wire _w13349_ ;
	wire _w13348_ ;
	wire _w13347_ ;
	wire _w13346_ ;
	wire _w13345_ ;
	wire _w13344_ ;
	wire _w13343_ ;
	wire _w13342_ ;
	wire _w13341_ ;
	wire _w13340_ ;
	wire _w13339_ ;
	wire _w13338_ ;
	wire _w13337_ ;
	wire _w13336_ ;
	wire _w13335_ ;
	wire _w13334_ ;
	wire _w13333_ ;
	wire _w13332_ ;
	wire _w13331_ ;
	wire _w13330_ ;
	wire _w13329_ ;
	wire _w13328_ ;
	wire _w13327_ ;
	wire _w13326_ ;
	wire _w13325_ ;
	wire _w13324_ ;
	wire _w13323_ ;
	wire _w13322_ ;
	wire _w13321_ ;
	wire _w13320_ ;
	wire _w13319_ ;
	wire _w13318_ ;
	wire _w13317_ ;
	wire _w13316_ ;
	wire _w13315_ ;
	wire _w13314_ ;
	wire _w13313_ ;
	wire _w13312_ ;
	wire _w13311_ ;
	wire _w13310_ ;
	wire _w13309_ ;
	wire _w13308_ ;
	wire _w13307_ ;
	wire _w13306_ ;
	wire _w13305_ ;
	wire _w13304_ ;
	wire _w13303_ ;
	wire _w13302_ ;
	wire _w13301_ ;
	wire _w13300_ ;
	wire _w13299_ ;
	wire _w13298_ ;
	wire _w13297_ ;
	wire _w13296_ ;
	wire _w13295_ ;
	wire _w13294_ ;
	wire _w13293_ ;
	wire _w13292_ ;
	wire _w13291_ ;
	wire _w13290_ ;
	wire _w13289_ ;
	wire _w13288_ ;
	wire _w13287_ ;
	wire _w13286_ ;
	wire _w13285_ ;
	wire _w13284_ ;
	wire _w13283_ ;
	wire _w13282_ ;
	wire _w13281_ ;
	wire _w13280_ ;
	wire _w13279_ ;
	wire _w13278_ ;
	wire _w13277_ ;
	wire _w13276_ ;
	wire _w13275_ ;
	wire _w13274_ ;
	wire _w13273_ ;
	wire _w13272_ ;
	wire _w13271_ ;
	wire _w13270_ ;
	wire _w13269_ ;
	wire _w13268_ ;
	wire _w13267_ ;
	wire _w13266_ ;
	wire _w13265_ ;
	wire _w13264_ ;
	wire _w13263_ ;
	wire _w13262_ ;
	wire _w13261_ ;
	wire _w13260_ ;
	wire _w13259_ ;
	wire _w13258_ ;
	wire _w13257_ ;
	wire _w13256_ ;
	wire _w13255_ ;
	wire _w13254_ ;
	wire _w13253_ ;
	wire _w13252_ ;
	wire _w13251_ ;
	wire _w13250_ ;
	wire _w13249_ ;
	wire _w13248_ ;
	wire _w13247_ ;
	wire _w13246_ ;
	wire _w13245_ ;
	wire _w13244_ ;
	wire _w13243_ ;
	wire _w13242_ ;
	wire _w13241_ ;
	wire _w13240_ ;
	wire _w13239_ ;
	wire _w13238_ ;
	wire _w13237_ ;
	wire _w13236_ ;
	wire _w13235_ ;
	wire _w13234_ ;
	wire _w13233_ ;
	wire _w13232_ ;
	wire _w13231_ ;
	wire _w13230_ ;
	wire _w13229_ ;
	wire _w13228_ ;
	wire _w13227_ ;
	wire _w13226_ ;
	wire _w13225_ ;
	wire _w13224_ ;
	wire _w13223_ ;
	wire _w13222_ ;
	wire _w13221_ ;
	wire _w13220_ ;
	wire _w13219_ ;
	wire _w13218_ ;
	wire _w13217_ ;
	wire _w13216_ ;
	wire _w13215_ ;
	wire _w13214_ ;
	wire _w13213_ ;
	wire _w13212_ ;
	wire _w13211_ ;
	wire _w13210_ ;
	wire _w13209_ ;
	wire _w13208_ ;
	wire _w13207_ ;
	wire _w13206_ ;
	wire _w13205_ ;
	wire _w13204_ ;
	wire _w13203_ ;
	wire _w13202_ ;
	wire _w13201_ ;
	wire _w13200_ ;
	wire _w13199_ ;
	wire _w13198_ ;
	wire _w13197_ ;
	wire _w13196_ ;
	wire _w13195_ ;
	wire _w13194_ ;
	wire _w13193_ ;
	wire _w13192_ ;
	wire _w13191_ ;
	wire _w13190_ ;
	wire _w13189_ ;
	wire _w13188_ ;
	wire _w13187_ ;
	wire _w13186_ ;
	wire _w13185_ ;
	wire _w13184_ ;
	wire _w13183_ ;
	wire _w13182_ ;
	wire _w13181_ ;
	wire _w13180_ ;
	wire _w13179_ ;
	wire _w13178_ ;
	wire _w13177_ ;
	wire _w13176_ ;
	wire _w13175_ ;
	wire _w13174_ ;
	wire _w13173_ ;
	wire _w13172_ ;
	wire _w13171_ ;
	wire _w13170_ ;
	wire _w13169_ ;
	wire _w13168_ ;
	wire _w13167_ ;
	wire _w13166_ ;
	wire _w13165_ ;
	wire _w13164_ ;
	wire _w13163_ ;
	wire _w13162_ ;
	wire _w13161_ ;
	wire _w13160_ ;
	wire _w13159_ ;
	wire _w13158_ ;
	wire _w13157_ ;
	wire _w13156_ ;
	wire _w13155_ ;
	wire _w13154_ ;
	wire _w13153_ ;
	wire _w13152_ ;
	wire _w13151_ ;
	wire _w13150_ ;
	wire _w13149_ ;
	wire _w13148_ ;
	wire _w13147_ ;
	wire _w13146_ ;
	wire _w13145_ ;
	wire _w13144_ ;
	wire _w13143_ ;
	wire _w13142_ ;
	wire _w13141_ ;
	wire _w13140_ ;
	wire _w13139_ ;
	wire _w13138_ ;
	wire _w13137_ ;
	wire _w13136_ ;
	wire _w13135_ ;
	wire _w13134_ ;
	wire _w13133_ ;
	wire _w13132_ ;
	wire _w13131_ ;
	wire _w13130_ ;
	wire _w13129_ ;
	wire _w13128_ ;
	wire _w13127_ ;
	wire _w13126_ ;
	wire _w13125_ ;
	wire _w13124_ ;
	wire _w13123_ ;
	wire _w13122_ ;
	wire _w13121_ ;
	wire _w13120_ ;
	wire _w13119_ ;
	wire _w13118_ ;
	wire _w13117_ ;
	wire _w13116_ ;
	wire _w13115_ ;
	wire _w13114_ ;
	wire _w13113_ ;
	wire _w13112_ ;
	wire _w13111_ ;
	wire _w13110_ ;
	wire _w13109_ ;
	wire _w13108_ ;
	wire _w13107_ ;
	wire _w13106_ ;
	wire _w13105_ ;
	wire _w13104_ ;
	wire _w13103_ ;
	wire _w13102_ ;
	wire _w13101_ ;
	wire _w13100_ ;
	wire _w13099_ ;
	wire _w13098_ ;
	wire _w13097_ ;
	wire _w13096_ ;
	wire _w13095_ ;
	wire _w13094_ ;
	wire _w13093_ ;
	wire _w13092_ ;
	wire _w13091_ ;
	wire _w13090_ ;
	wire _w13089_ ;
	wire _w13088_ ;
	wire _w13087_ ;
	wire _w13086_ ;
	wire _w13085_ ;
	wire _w13084_ ;
	wire _w13083_ ;
	wire _w13082_ ;
	wire _w13081_ ;
	wire _w13080_ ;
	wire _w13079_ ;
	wire _w13078_ ;
	wire _w13077_ ;
	wire _w13076_ ;
	wire _w13075_ ;
	wire _w13074_ ;
	wire _w13073_ ;
	wire _w13072_ ;
	wire _w13071_ ;
	wire _w13070_ ;
	wire _w13069_ ;
	wire _w13068_ ;
	wire _w13067_ ;
	wire _w13066_ ;
	wire _w13065_ ;
	wire _w13064_ ;
	wire _w13063_ ;
	wire _w13062_ ;
	wire _w13061_ ;
	wire _w13060_ ;
	wire _w13059_ ;
	wire _w13058_ ;
	wire _w13057_ ;
	wire _w13056_ ;
	wire _w13055_ ;
	wire _w13054_ ;
	wire _w13053_ ;
	wire _w13052_ ;
	wire _w13051_ ;
	wire _w13050_ ;
	wire _w13049_ ;
	wire _w13048_ ;
	wire _w13047_ ;
	wire _w13046_ ;
	wire _w13045_ ;
	wire _w13044_ ;
	wire _w13043_ ;
	wire _w13042_ ;
	wire _w13041_ ;
	wire _w13040_ ;
	wire _w13039_ ;
	wire _w13038_ ;
	wire _w13037_ ;
	wire _w13036_ ;
	wire _w13035_ ;
	wire _w13034_ ;
	wire _w13033_ ;
	wire _w13032_ ;
	wire _w13031_ ;
	wire _w13030_ ;
	wire _w13029_ ;
	wire _w13028_ ;
	wire _w13027_ ;
	wire _w13026_ ;
	wire _w13025_ ;
	wire _w13024_ ;
	wire _w13023_ ;
	wire _w13022_ ;
	wire _w13021_ ;
	wire _w13020_ ;
	wire _w13019_ ;
	wire _w13018_ ;
	wire _w13017_ ;
	wire _w13016_ ;
	wire _w13015_ ;
	wire _w13014_ ;
	wire _w13013_ ;
	wire _w13012_ ;
	wire _w13011_ ;
	wire _w13010_ ;
	wire _w13009_ ;
	wire _w13008_ ;
	wire _w13007_ ;
	wire _w13006_ ;
	wire _w13005_ ;
	wire _w13004_ ;
	wire _w13003_ ;
	wire _w13002_ ;
	wire _w13001_ ;
	wire _w13000_ ;
	wire _w12999_ ;
	wire _w12998_ ;
	wire _w12997_ ;
	wire _w12996_ ;
	wire _w12995_ ;
	wire _w12994_ ;
	wire _w12993_ ;
	wire _w12992_ ;
	wire _w12991_ ;
	wire _w12990_ ;
	wire _w12989_ ;
	wire _w12988_ ;
	wire _w12987_ ;
	wire _w12986_ ;
	wire _w12985_ ;
	wire _w12984_ ;
	wire _w12983_ ;
	wire _w12982_ ;
	wire _w12981_ ;
	wire _w12980_ ;
	wire _w12979_ ;
	wire _w12978_ ;
	wire _w12977_ ;
	wire _w12976_ ;
	wire _w12975_ ;
	wire _w12974_ ;
	wire _w12973_ ;
	wire _w12972_ ;
	wire _w12971_ ;
	wire _w12970_ ;
	wire _w12969_ ;
	wire _w12968_ ;
	wire _w12967_ ;
	wire _w12966_ ;
	wire _w12965_ ;
	wire _w12964_ ;
	wire _w12963_ ;
	wire _w12962_ ;
	wire _w12961_ ;
	wire _w12960_ ;
	wire _w12959_ ;
	wire _w12958_ ;
	wire _w12957_ ;
	wire _w12956_ ;
	wire _w12955_ ;
	wire _w12954_ ;
	wire _w12953_ ;
	wire _w12952_ ;
	wire _w12951_ ;
	wire _w12950_ ;
	wire _w12949_ ;
	wire _w12948_ ;
	wire _w12947_ ;
	wire _w12946_ ;
	wire _w12945_ ;
	wire _w12944_ ;
	wire _w12943_ ;
	wire _w12942_ ;
	wire _w12941_ ;
	wire _w12940_ ;
	wire _w12939_ ;
	wire _w12938_ ;
	wire _w12937_ ;
	wire _w12936_ ;
	wire _w12935_ ;
	wire _w12934_ ;
	wire _w12933_ ;
	wire _w12932_ ;
	wire _w12931_ ;
	wire _w12930_ ;
	wire _w12929_ ;
	wire _w12928_ ;
	wire _w12927_ ;
	wire _w12926_ ;
	wire _w12925_ ;
	wire _w12924_ ;
	wire _w12923_ ;
	wire _w12922_ ;
	wire _w12921_ ;
	wire _w12920_ ;
	wire _w12919_ ;
	wire _w12918_ ;
	wire _w12917_ ;
	wire _w12916_ ;
	wire _w12915_ ;
	wire _w12914_ ;
	wire _w12913_ ;
	wire _w12912_ ;
	wire _w12911_ ;
	wire _w12910_ ;
	wire _w12909_ ;
	wire _w12908_ ;
	wire _w12907_ ;
	wire _w12906_ ;
	wire _w12905_ ;
	wire _w12904_ ;
	wire _w12903_ ;
	wire _w12902_ ;
	wire _w12901_ ;
	wire _w12900_ ;
	wire _w12899_ ;
	wire _w12898_ ;
	wire _w12897_ ;
	wire _w12896_ ;
	wire _w12895_ ;
	wire _w12894_ ;
	wire _w12893_ ;
	wire _w12892_ ;
	wire _w12891_ ;
	wire _w12890_ ;
	wire _w12889_ ;
	wire _w12888_ ;
	wire _w12887_ ;
	wire _w12886_ ;
	wire _w12885_ ;
	wire _w12884_ ;
	wire _w12883_ ;
	wire _w12882_ ;
	wire _w12881_ ;
	wire _w12880_ ;
	wire _w12879_ ;
	wire _w12878_ ;
	wire _w12877_ ;
	wire _w12876_ ;
	wire _w12875_ ;
	wire _w12874_ ;
	wire _w12873_ ;
	wire _w12872_ ;
	wire _w12871_ ;
	wire _w12870_ ;
	wire _w12869_ ;
	wire _w12868_ ;
	wire _w12867_ ;
	wire _w12866_ ;
	wire _w12865_ ;
	wire _w12864_ ;
	wire _w12863_ ;
	wire _w12862_ ;
	wire _w12861_ ;
	wire _w12860_ ;
	wire _w12859_ ;
	wire _w12858_ ;
	wire _w12857_ ;
	wire _w12856_ ;
	wire _w12855_ ;
	wire _w12854_ ;
	wire _w12853_ ;
	wire _w12852_ ;
	wire _w12851_ ;
	wire _w12850_ ;
	wire _w12849_ ;
	wire _w12848_ ;
	wire _w12847_ ;
	wire _w12846_ ;
	wire _w12845_ ;
	wire _w12844_ ;
	wire _w12843_ ;
	wire _w12842_ ;
	wire _w12841_ ;
	wire _w12840_ ;
	wire _w12839_ ;
	wire _w12838_ ;
	wire _w12837_ ;
	wire _w12836_ ;
	wire _w12835_ ;
	wire _w12834_ ;
	wire _w12833_ ;
	wire _w12832_ ;
	wire _w12831_ ;
	wire _w12830_ ;
	wire _w12829_ ;
	wire _w12828_ ;
	wire _w12827_ ;
	wire _w12826_ ;
	wire _w12825_ ;
	wire _w12824_ ;
	wire _w12823_ ;
	wire _w12822_ ;
	wire _w12821_ ;
	wire _w12820_ ;
	wire _w12819_ ;
	wire _w12818_ ;
	wire _w12817_ ;
	wire _w12816_ ;
	wire _w12815_ ;
	wire _w12814_ ;
	wire _w12813_ ;
	wire _w12812_ ;
	wire _w12811_ ;
	wire _w12810_ ;
	wire _w12809_ ;
	wire _w12808_ ;
	wire _w12807_ ;
	wire _w12806_ ;
	wire _w12805_ ;
	wire _w12804_ ;
	wire _w12803_ ;
	wire _w12802_ ;
	wire _w12801_ ;
	wire _w12800_ ;
	wire _w12799_ ;
	wire _w12798_ ;
	wire _w12797_ ;
	wire _w12796_ ;
	wire _w12795_ ;
	wire _w12794_ ;
	wire _w12793_ ;
	wire _w12792_ ;
	wire _w12791_ ;
	wire _w12790_ ;
	wire _w12789_ ;
	wire _w12788_ ;
	wire _w12787_ ;
	wire _w12786_ ;
	wire _w12785_ ;
	wire _w12784_ ;
	wire _w12783_ ;
	wire _w12782_ ;
	wire _w12781_ ;
	wire _w12780_ ;
	wire _w12779_ ;
	wire _w12778_ ;
	wire _w12777_ ;
	wire _w12776_ ;
	wire _w12775_ ;
	wire _w12774_ ;
	wire _w12773_ ;
	wire _w12772_ ;
	wire _w12771_ ;
	wire _w12770_ ;
	wire _w12769_ ;
	wire _w12768_ ;
	wire _w12767_ ;
	wire _w12766_ ;
	wire _w12765_ ;
	wire _w12764_ ;
	wire _w12763_ ;
	wire _w12762_ ;
	wire _w12761_ ;
	wire _w12760_ ;
	wire _w12759_ ;
	wire _w12758_ ;
	wire _w12757_ ;
	wire _w12756_ ;
	wire _w12755_ ;
	wire _w12754_ ;
	wire _w12753_ ;
	wire _w12752_ ;
	wire _w12751_ ;
	wire _w12750_ ;
	wire _w12749_ ;
	wire _w12748_ ;
	wire _w12747_ ;
	wire _w12746_ ;
	wire _w12745_ ;
	wire _w12744_ ;
	wire _w12743_ ;
	wire _w12742_ ;
	wire _w12741_ ;
	wire _w12740_ ;
	wire _w12739_ ;
	wire _w12738_ ;
	wire _w12737_ ;
	wire _w12736_ ;
	wire _w12735_ ;
	wire _w12734_ ;
	wire _w12733_ ;
	wire _w12732_ ;
	wire _w12731_ ;
	wire _w12730_ ;
	wire _w12729_ ;
	wire _w12728_ ;
	wire _w12727_ ;
	wire _w12726_ ;
	wire _w12725_ ;
	wire _w12724_ ;
	wire _w12723_ ;
	wire _w12722_ ;
	wire _w12721_ ;
	wire _w12720_ ;
	wire _w12719_ ;
	wire _w12718_ ;
	wire _w12717_ ;
	wire _w12716_ ;
	wire _w12715_ ;
	wire _w12714_ ;
	wire _w12713_ ;
	wire _w12712_ ;
	wire _w12711_ ;
	wire _w12710_ ;
	wire _w12709_ ;
	wire _w12708_ ;
	wire _w12707_ ;
	wire _w12706_ ;
	wire _w12705_ ;
	wire _w12704_ ;
	wire _w12703_ ;
	wire _w12702_ ;
	wire _w12701_ ;
	wire _w12700_ ;
	wire _w12699_ ;
	wire _w12698_ ;
	wire _w12697_ ;
	wire _w12696_ ;
	wire _w12695_ ;
	wire _w12694_ ;
	wire _w12693_ ;
	wire _w12692_ ;
	wire _w12691_ ;
	wire _w12690_ ;
	wire _w12689_ ;
	wire _w12688_ ;
	wire _w12687_ ;
	wire _w12686_ ;
	wire _w12685_ ;
	wire _w12684_ ;
	wire _w12683_ ;
	wire _w12682_ ;
	wire _w12681_ ;
	wire _w12680_ ;
	wire _w12679_ ;
	wire _w12678_ ;
	wire _w12677_ ;
	wire _w12676_ ;
	wire _w12675_ ;
	wire _w12674_ ;
	wire _w12673_ ;
	wire _w12672_ ;
	wire _w12671_ ;
	wire _w12670_ ;
	wire _w12669_ ;
	wire _w12668_ ;
	wire _w12667_ ;
	wire _w12666_ ;
	wire _w12665_ ;
	wire _w12664_ ;
	wire _w12663_ ;
	wire _w12662_ ;
	wire _w12661_ ;
	wire _w12660_ ;
	wire _w12659_ ;
	wire _w12658_ ;
	wire _w12657_ ;
	wire _w12656_ ;
	wire _w12655_ ;
	wire _w12654_ ;
	wire _w12653_ ;
	wire _w12652_ ;
	wire _w12651_ ;
	wire _w12650_ ;
	wire _w12649_ ;
	wire _w12648_ ;
	wire _w12647_ ;
	wire _w12646_ ;
	wire _w12645_ ;
	wire _w12644_ ;
	wire _w12643_ ;
	wire _w12642_ ;
	wire _w12641_ ;
	wire _w12640_ ;
	wire _w12639_ ;
	wire _w12638_ ;
	wire _w12637_ ;
	wire _w12636_ ;
	wire _w12635_ ;
	wire _w12634_ ;
	wire _w12633_ ;
	wire _w12632_ ;
	wire _w12631_ ;
	wire _w12630_ ;
	wire _w12629_ ;
	wire _w12628_ ;
	wire _w12627_ ;
	wire _w12626_ ;
	wire _w12625_ ;
	wire _w12624_ ;
	wire _w12623_ ;
	wire _w12622_ ;
	wire _w12621_ ;
	wire _w12620_ ;
	wire _w12619_ ;
	wire _w12618_ ;
	wire _w12617_ ;
	wire _w12616_ ;
	wire _w12615_ ;
	wire _w12614_ ;
	wire _w12613_ ;
	wire _w12612_ ;
	wire _w12611_ ;
	wire _w12610_ ;
	wire _w12609_ ;
	wire _w12608_ ;
	wire _w12607_ ;
	wire _w12606_ ;
	wire _w12605_ ;
	wire _w12604_ ;
	wire _w12603_ ;
	wire _w12602_ ;
	wire _w12601_ ;
	wire _w12600_ ;
	wire _w12599_ ;
	wire _w12598_ ;
	wire _w12597_ ;
	wire _w12596_ ;
	wire _w12595_ ;
	wire _w12594_ ;
	wire _w12593_ ;
	wire _w12592_ ;
	wire _w12591_ ;
	wire _w12590_ ;
	wire _w12589_ ;
	wire _w12588_ ;
	wire _w12587_ ;
	wire _w12586_ ;
	wire _w12585_ ;
	wire _w12584_ ;
	wire _w12583_ ;
	wire _w12582_ ;
	wire _w12581_ ;
	wire _w12580_ ;
	wire _w12579_ ;
	wire _w12578_ ;
	wire _w12577_ ;
	wire _w12576_ ;
	wire _w12575_ ;
	wire _w12574_ ;
	wire _w12573_ ;
	wire _w12572_ ;
	wire _w12571_ ;
	wire _w12570_ ;
	wire _w12569_ ;
	wire _w12568_ ;
	wire _w12567_ ;
	wire _w12566_ ;
	wire _w12565_ ;
	wire _w12564_ ;
	wire _w12563_ ;
	wire _w12562_ ;
	wire _w12561_ ;
	wire _w12560_ ;
	wire _w12559_ ;
	wire _w12558_ ;
	wire _w12557_ ;
	wire _w12556_ ;
	wire _w12555_ ;
	wire _w12554_ ;
	wire _w12553_ ;
	wire _w12552_ ;
	wire _w12551_ ;
	wire _w12550_ ;
	wire _w12549_ ;
	wire _w12548_ ;
	wire _w12547_ ;
	wire _w12546_ ;
	wire _w12545_ ;
	wire _w12544_ ;
	wire _w12543_ ;
	wire _w12542_ ;
	wire _w12541_ ;
	wire _w12540_ ;
	wire _w12539_ ;
	wire _w12538_ ;
	wire _w12537_ ;
	wire _w12536_ ;
	wire _w12535_ ;
	wire _w12534_ ;
	wire _w12533_ ;
	wire _w12532_ ;
	wire _w12531_ ;
	wire _w12530_ ;
	wire _w12529_ ;
	wire _w12528_ ;
	wire _w12527_ ;
	wire _w12526_ ;
	wire _w12525_ ;
	wire _w12524_ ;
	wire _w12523_ ;
	wire _w12522_ ;
	wire _w12521_ ;
	wire _w12520_ ;
	wire _w12519_ ;
	wire _w12518_ ;
	wire _w12517_ ;
	wire _w12516_ ;
	wire _w12515_ ;
	wire _w12514_ ;
	wire _w12513_ ;
	wire _w12512_ ;
	wire _w12511_ ;
	wire _w12510_ ;
	wire _w12509_ ;
	wire _w12508_ ;
	wire _w12507_ ;
	wire _w12506_ ;
	wire _w12505_ ;
	wire _w12504_ ;
	wire _w12503_ ;
	wire _w12502_ ;
	wire _w12501_ ;
	wire _w12500_ ;
	wire _w12499_ ;
	wire _w12498_ ;
	wire _w12497_ ;
	wire _w12496_ ;
	wire _w12495_ ;
	wire _w12494_ ;
	wire _w12493_ ;
	wire _w12492_ ;
	wire _w12491_ ;
	wire _w12490_ ;
	wire _w12489_ ;
	wire _w12488_ ;
	wire _w12487_ ;
	wire _w12486_ ;
	wire _w12485_ ;
	wire _w12484_ ;
	wire _w12483_ ;
	wire _w12482_ ;
	wire _w12481_ ;
	wire _w12480_ ;
	wire _w12479_ ;
	wire _w12478_ ;
	wire _w12477_ ;
	wire _w12476_ ;
	wire _w12475_ ;
	wire _w12474_ ;
	wire _w12473_ ;
	wire _w12472_ ;
	wire _w12471_ ;
	wire _w12470_ ;
	wire _w12469_ ;
	wire _w12468_ ;
	wire _w12467_ ;
	wire _w12466_ ;
	wire _w12465_ ;
	wire _w12464_ ;
	wire _w12463_ ;
	wire _w12462_ ;
	wire _w12461_ ;
	wire _w12460_ ;
	wire _w12459_ ;
	wire _w12458_ ;
	wire _w12457_ ;
	wire _w12456_ ;
	wire _w12455_ ;
	wire _w12454_ ;
	wire _w12453_ ;
	wire _w12452_ ;
	wire _w12451_ ;
	wire _w12450_ ;
	wire _w12449_ ;
	wire _w12448_ ;
	wire _w12447_ ;
	wire _w12446_ ;
	wire _w12445_ ;
	wire _w12444_ ;
	wire _w12443_ ;
	wire _w12442_ ;
	wire _w12441_ ;
	wire _w12440_ ;
	wire _w12439_ ;
	wire _w12438_ ;
	wire _w12437_ ;
	wire _w12436_ ;
	wire _w12435_ ;
	wire _w12434_ ;
	wire _w12433_ ;
	wire _w12432_ ;
	wire _w12431_ ;
	wire _w12430_ ;
	wire _w12429_ ;
	wire _w12428_ ;
	wire _w12427_ ;
	wire _w12426_ ;
	wire _w12425_ ;
	wire _w12424_ ;
	wire _w12423_ ;
	wire _w12422_ ;
	wire _w12421_ ;
	wire _w12420_ ;
	wire _w12419_ ;
	wire _w12418_ ;
	wire _w12417_ ;
	wire _w12416_ ;
	wire _w12415_ ;
	wire _w12414_ ;
	wire _w12413_ ;
	wire _w12412_ ;
	wire _w12411_ ;
	wire _w12410_ ;
	wire _w12409_ ;
	wire _w12408_ ;
	wire _w12407_ ;
	wire _w12406_ ;
	wire _w12405_ ;
	wire _w12404_ ;
	wire _w12403_ ;
	wire _w12402_ ;
	wire _w12401_ ;
	wire _w12400_ ;
	wire _w12399_ ;
	wire _w12398_ ;
	wire _w12397_ ;
	wire _w12396_ ;
	wire _w12395_ ;
	wire _w12394_ ;
	wire _w12393_ ;
	wire _w12392_ ;
	wire _w12391_ ;
	wire _w12390_ ;
	wire _w12389_ ;
	wire _w12388_ ;
	wire _w12387_ ;
	wire _w12386_ ;
	wire _w12385_ ;
	wire _w12384_ ;
	wire _w12383_ ;
	wire _w12382_ ;
	wire _w12381_ ;
	wire _w12380_ ;
	wire _w12379_ ;
	wire _w12378_ ;
	wire _w12377_ ;
	wire _w12376_ ;
	wire _w12375_ ;
	wire _w12374_ ;
	wire _w12373_ ;
	wire _w12372_ ;
	wire _w12371_ ;
	wire _w12370_ ;
	wire _w12369_ ;
	wire _w12368_ ;
	wire _w12367_ ;
	wire _w12366_ ;
	wire _w12365_ ;
	wire _w12364_ ;
	wire _w12363_ ;
	wire _w12362_ ;
	wire _w12361_ ;
	wire _w12360_ ;
	wire _w12359_ ;
	wire _w12358_ ;
	wire _w12357_ ;
	wire _w12356_ ;
	wire _w12355_ ;
	wire _w12354_ ;
	wire _w12353_ ;
	wire _w12352_ ;
	wire _w12351_ ;
	wire _w12350_ ;
	wire _w12349_ ;
	wire _w12348_ ;
	wire _w12347_ ;
	wire _w12346_ ;
	wire _w12345_ ;
	wire _w12344_ ;
	wire _w12343_ ;
	wire _w12342_ ;
	wire _w12341_ ;
	wire _w12340_ ;
	wire _w12339_ ;
	wire _w12338_ ;
	wire _w12337_ ;
	wire _w12336_ ;
	wire _w12335_ ;
	wire _w12334_ ;
	wire _w12333_ ;
	wire _w12332_ ;
	wire _w12331_ ;
	wire _w12330_ ;
	wire _w12329_ ;
	wire _w12328_ ;
	wire _w12327_ ;
	wire _w12326_ ;
	wire _w12325_ ;
	wire _w12324_ ;
	wire _w12323_ ;
	wire _w12322_ ;
	wire _w12321_ ;
	wire _w12320_ ;
	wire _w12319_ ;
	wire _w12318_ ;
	wire _w12317_ ;
	wire _w12316_ ;
	wire _w12315_ ;
	wire _w12314_ ;
	wire _w12313_ ;
	wire _w12312_ ;
	wire _w12311_ ;
	wire _w12310_ ;
	wire _w12309_ ;
	wire _w12308_ ;
	wire _w12307_ ;
	wire _w12306_ ;
	wire _w12305_ ;
	wire _w12304_ ;
	wire _w12303_ ;
	wire _w12302_ ;
	wire _w12301_ ;
	wire _w12300_ ;
	wire _w12299_ ;
	wire _w12298_ ;
	wire _w12297_ ;
	wire _w12296_ ;
	wire _w12295_ ;
	wire _w12294_ ;
	wire _w12293_ ;
	wire _w12292_ ;
	wire _w12291_ ;
	wire _w12290_ ;
	wire _w12289_ ;
	wire _w12288_ ;
	wire _w12287_ ;
	wire _w12286_ ;
	wire _w12285_ ;
	wire _w12284_ ;
	wire _w12283_ ;
	wire _w12282_ ;
	wire _w12281_ ;
	wire _w12280_ ;
	wire _w12279_ ;
	wire _w12278_ ;
	wire _w12277_ ;
	wire _w12276_ ;
	wire _w12275_ ;
	wire _w12274_ ;
	wire _w12273_ ;
	wire _w12272_ ;
	wire _w12271_ ;
	wire _w12270_ ;
	wire _w12269_ ;
	wire _w12268_ ;
	wire _w12267_ ;
	wire _w12266_ ;
	wire _w12265_ ;
	wire _w12264_ ;
	wire _w12263_ ;
	wire _w12262_ ;
	wire _w12261_ ;
	wire _w12260_ ;
	wire _w12259_ ;
	wire _w12258_ ;
	wire _w12257_ ;
	wire _w12256_ ;
	wire _w12255_ ;
	wire _w12254_ ;
	wire _w12253_ ;
	wire _w12252_ ;
	wire _w12251_ ;
	wire _w12250_ ;
	wire _w12249_ ;
	wire _w12248_ ;
	wire _w12247_ ;
	wire _w12246_ ;
	wire _w12245_ ;
	wire _w12244_ ;
	wire _w12243_ ;
	wire _w12242_ ;
	wire _w12241_ ;
	wire _w12240_ ;
	wire _w12239_ ;
	wire _w12238_ ;
	wire _w12237_ ;
	wire _w12236_ ;
	wire _w12235_ ;
	wire _w12234_ ;
	wire _w12233_ ;
	wire _w12232_ ;
	wire _w12231_ ;
	wire _w12230_ ;
	wire _w12229_ ;
	wire _w12228_ ;
	wire _w12227_ ;
	wire _w12226_ ;
	wire _w12225_ ;
	wire _w12224_ ;
	wire _w12223_ ;
	wire _w12222_ ;
	wire _w12221_ ;
	wire _w12220_ ;
	wire _w12219_ ;
	wire _w12218_ ;
	wire _w12217_ ;
	wire _w12216_ ;
	wire _w12215_ ;
	wire _w12214_ ;
	wire _w12213_ ;
	wire _w12212_ ;
	wire _w12211_ ;
	wire _w12210_ ;
	wire _w12209_ ;
	wire _w12208_ ;
	wire _w12207_ ;
	wire _w12206_ ;
	wire _w12205_ ;
	wire _w12204_ ;
	wire _w12203_ ;
	wire _w12202_ ;
	wire _w12201_ ;
	wire _w12200_ ;
	wire _w12199_ ;
	wire _w12198_ ;
	wire _w12197_ ;
	wire _w12196_ ;
	wire _w12195_ ;
	wire _w12194_ ;
	wire _w12193_ ;
	wire _w12192_ ;
	wire _w12191_ ;
	wire _w12190_ ;
	wire _w12189_ ;
	wire _w12188_ ;
	wire _w12187_ ;
	wire _w12186_ ;
	wire _w12185_ ;
	wire _w12184_ ;
	wire _w12183_ ;
	wire _w12182_ ;
	wire _w12181_ ;
	wire _w12180_ ;
	wire _w12179_ ;
	wire _w12178_ ;
	wire _w12177_ ;
	wire _w12176_ ;
	wire _w12175_ ;
	wire _w12174_ ;
	wire _w12173_ ;
	wire _w12172_ ;
	wire _w12171_ ;
	wire _w12170_ ;
	wire _w12169_ ;
	wire _w12168_ ;
	wire _w12167_ ;
	wire _w12166_ ;
	wire _w12165_ ;
	wire _w12164_ ;
	wire _w12163_ ;
	wire _w12162_ ;
	wire _w12161_ ;
	wire _w12160_ ;
	wire _w12159_ ;
	wire _w12158_ ;
	wire _w12157_ ;
	wire _w12156_ ;
	wire _w12155_ ;
	wire _w12154_ ;
	wire _w12153_ ;
	wire _w12152_ ;
	wire _w12151_ ;
	wire _w12150_ ;
	wire _w12149_ ;
	wire _w12148_ ;
	wire _w12147_ ;
	wire _w12146_ ;
	wire _w12145_ ;
	wire _w12144_ ;
	wire _w12143_ ;
	wire _w12142_ ;
	wire _w12141_ ;
	wire _w12140_ ;
	wire _w12139_ ;
	wire _w12138_ ;
	wire _w12137_ ;
	wire _w12136_ ;
	wire _w12135_ ;
	wire _w12134_ ;
	wire _w12133_ ;
	wire _w12132_ ;
	wire _w12131_ ;
	wire _w12130_ ;
	wire _w12129_ ;
	wire _w12128_ ;
	wire _w12127_ ;
	wire _w12126_ ;
	wire _w12125_ ;
	wire _w12124_ ;
	wire _w12123_ ;
	wire _w12122_ ;
	wire _w12121_ ;
	wire _w12120_ ;
	wire _w12119_ ;
	wire _w12118_ ;
	wire _w12117_ ;
	wire _w12116_ ;
	wire _w12115_ ;
	wire _w12114_ ;
	wire _w12113_ ;
	wire _w12112_ ;
	wire _w12111_ ;
	wire _w12110_ ;
	wire _w12109_ ;
	wire _w12108_ ;
	wire _w12107_ ;
	wire _w12106_ ;
	wire _w12105_ ;
	wire _w12104_ ;
	wire _w12103_ ;
	wire _w12102_ ;
	wire _w12101_ ;
	wire _w12100_ ;
	wire _w12099_ ;
	wire _w12098_ ;
	wire _w12097_ ;
	wire _w12096_ ;
	wire _w12095_ ;
	wire _w12094_ ;
	wire _w12093_ ;
	wire _w12092_ ;
	wire _w12091_ ;
	wire _w12090_ ;
	wire _w12089_ ;
	wire _w12088_ ;
	wire _w12087_ ;
	wire _w12086_ ;
	wire _w12085_ ;
	wire _w12084_ ;
	wire _w12083_ ;
	wire _w12082_ ;
	wire _w12081_ ;
	wire _w12080_ ;
	wire _w12079_ ;
	wire _w12078_ ;
	wire _w12077_ ;
	wire _w12076_ ;
	wire _w12075_ ;
	wire _w12074_ ;
	wire _w12073_ ;
	wire _w12072_ ;
	wire _w12071_ ;
	wire _w12070_ ;
	wire _w12069_ ;
	wire _w12068_ ;
	wire _w12067_ ;
	wire _w12066_ ;
	wire _w12065_ ;
	wire _w12064_ ;
	wire _w12063_ ;
	wire _w12062_ ;
	wire _w12061_ ;
	wire _w12060_ ;
	wire _w12059_ ;
	wire _w12058_ ;
	wire _w12057_ ;
	wire _w12056_ ;
	wire _w12055_ ;
	wire _w12054_ ;
	wire _w12053_ ;
	wire _w12052_ ;
	wire _w12051_ ;
	wire _w12050_ ;
	wire _w12049_ ;
	wire _w12048_ ;
	wire _w12047_ ;
	wire _w12046_ ;
	wire _w12045_ ;
	wire _w12044_ ;
	wire _w12043_ ;
	wire _w12042_ ;
	wire _w12041_ ;
	wire _w12040_ ;
	wire _w12039_ ;
	wire _w12038_ ;
	wire _w12037_ ;
	wire _w12036_ ;
	wire _w12035_ ;
	wire _w12034_ ;
	wire _w12033_ ;
	wire _w12032_ ;
	wire _w12031_ ;
	wire _w12030_ ;
	wire _w12029_ ;
	wire _w12028_ ;
	wire _w12027_ ;
	wire _w12026_ ;
	wire _w12025_ ;
	wire _w12024_ ;
	wire _w12023_ ;
	wire _w12022_ ;
	wire _w12021_ ;
	wire _w12020_ ;
	wire _w12019_ ;
	wire _w12018_ ;
	wire _w12017_ ;
	wire _w12016_ ;
	wire _w12015_ ;
	wire _w12014_ ;
	wire _w12013_ ;
	wire _w12012_ ;
	wire _w12011_ ;
	wire _w12010_ ;
	wire _w12009_ ;
	wire _w12008_ ;
	wire _w12007_ ;
	wire _w12006_ ;
	wire _w12005_ ;
	wire _w12004_ ;
	wire _w12003_ ;
	wire _w12002_ ;
	wire _w12001_ ;
	wire _w12000_ ;
	wire _w11999_ ;
	wire _w11998_ ;
	wire _w11997_ ;
	wire _w11996_ ;
	wire _w11995_ ;
	wire _w11994_ ;
	wire _w11993_ ;
	wire _w11992_ ;
	wire _w11991_ ;
	wire _w11990_ ;
	wire _w11989_ ;
	wire _w11988_ ;
	wire _w11987_ ;
	wire _w11986_ ;
	wire _w11985_ ;
	wire _w11984_ ;
	wire _w11983_ ;
	wire _w11982_ ;
	wire _w11981_ ;
	wire _w11980_ ;
	wire _w11979_ ;
	wire _w11978_ ;
	wire _w11977_ ;
	wire _w11976_ ;
	wire _w11975_ ;
	wire _w11974_ ;
	wire _w11973_ ;
	wire _w11972_ ;
	wire _w11971_ ;
	wire _w11970_ ;
	wire _w11969_ ;
	wire _w11968_ ;
	wire _w11967_ ;
	wire _w11966_ ;
	wire _w11965_ ;
	wire _w11964_ ;
	wire _w11963_ ;
	wire _w11962_ ;
	wire _w11961_ ;
	wire _w11960_ ;
	wire _w11959_ ;
	wire _w11958_ ;
	wire _w11957_ ;
	wire _w11956_ ;
	wire _w11955_ ;
	wire _w11954_ ;
	wire _w11953_ ;
	wire _w11952_ ;
	wire _w11951_ ;
	wire _w11950_ ;
	wire _w11949_ ;
	wire _w11948_ ;
	wire _w11947_ ;
	wire _w11946_ ;
	wire _w11945_ ;
	wire _w11944_ ;
	wire _w11943_ ;
	wire _w11942_ ;
	wire _w11941_ ;
	wire _w11940_ ;
	wire _w11939_ ;
	wire _w11938_ ;
	wire _w11937_ ;
	wire _w11936_ ;
	wire _w11935_ ;
	wire _w11934_ ;
	wire _w11933_ ;
	wire _w11932_ ;
	wire _w11931_ ;
	wire _w11930_ ;
	wire _w11929_ ;
	wire _w11928_ ;
	wire _w11927_ ;
	wire _w11926_ ;
	wire _w11925_ ;
	wire _w11924_ ;
	wire _w11923_ ;
	wire _w11922_ ;
	wire _w11921_ ;
	wire _w11920_ ;
	wire _w11919_ ;
	wire _w11918_ ;
	wire _w11917_ ;
	wire _w11916_ ;
	wire _w11915_ ;
	wire _w11914_ ;
	wire _w11913_ ;
	wire _w11912_ ;
	wire _w11911_ ;
	wire _w11910_ ;
	wire _w11909_ ;
	wire _w11908_ ;
	wire _w11907_ ;
	wire _w11906_ ;
	wire _w11905_ ;
	wire _w11904_ ;
	wire _w11903_ ;
	wire _w11902_ ;
	wire _w11901_ ;
	wire _w11900_ ;
	wire _w11899_ ;
	wire _w11898_ ;
	wire _w11897_ ;
	wire _w11896_ ;
	wire _w11895_ ;
	wire _w11894_ ;
	wire _w11893_ ;
	wire _w11892_ ;
	wire _w11891_ ;
	wire _w11890_ ;
	wire _w11889_ ;
	wire _w11888_ ;
	wire _w11887_ ;
	wire _w11886_ ;
	wire _w11885_ ;
	wire _w11884_ ;
	wire _w11883_ ;
	wire _w11882_ ;
	wire _w11881_ ;
	wire _w11880_ ;
	wire _w11879_ ;
	wire _w11878_ ;
	wire _w11877_ ;
	wire _w11876_ ;
	wire _w11875_ ;
	wire _w11874_ ;
	wire _w11873_ ;
	wire _w11872_ ;
	wire _w11871_ ;
	wire _w11870_ ;
	wire _w11869_ ;
	wire _w11868_ ;
	wire _w11867_ ;
	wire _w11866_ ;
	wire _w11865_ ;
	wire _w11864_ ;
	wire _w11863_ ;
	wire _w11862_ ;
	wire _w11861_ ;
	wire _w11860_ ;
	wire _w11859_ ;
	wire _w11858_ ;
	wire _w11857_ ;
	wire _w11856_ ;
	wire _w11855_ ;
	wire _w11854_ ;
	wire _w11853_ ;
	wire _w11852_ ;
	wire _w11851_ ;
	wire _w11850_ ;
	wire _w11849_ ;
	wire _w11848_ ;
	wire _w11847_ ;
	wire _w11846_ ;
	wire _w11845_ ;
	wire _w11844_ ;
	wire _w11843_ ;
	wire _w11842_ ;
	wire _w11841_ ;
	wire _w11840_ ;
	wire _w11839_ ;
	wire _w11838_ ;
	wire _w11837_ ;
	wire _w11836_ ;
	wire _w11835_ ;
	wire _w11834_ ;
	wire _w11833_ ;
	wire _w11832_ ;
	wire _w11831_ ;
	wire _w11830_ ;
	wire _w11829_ ;
	wire _w11828_ ;
	wire _w11827_ ;
	wire _w11826_ ;
	wire _w11825_ ;
	wire _w11824_ ;
	wire _w11823_ ;
	wire _w11822_ ;
	wire _w11821_ ;
	wire _w11820_ ;
	wire _w11819_ ;
	wire _w11818_ ;
	wire _w11817_ ;
	wire _w11816_ ;
	wire _w11815_ ;
	wire _w11814_ ;
	wire _w11813_ ;
	wire _w11812_ ;
	wire _w11811_ ;
	wire _w11810_ ;
	wire _w11809_ ;
	wire _w11808_ ;
	wire _w11807_ ;
	wire _w11806_ ;
	wire _w11805_ ;
	wire _w11804_ ;
	wire _w11803_ ;
	wire _w11802_ ;
	wire _w11801_ ;
	wire _w11800_ ;
	wire _w11799_ ;
	wire _w11798_ ;
	wire _w11797_ ;
	wire _w11796_ ;
	wire _w11795_ ;
	wire _w11794_ ;
	wire _w11793_ ;
	wire _w11792_ ;
	wire _w11791_ ;
	wire _w11790_ ;
	wire _w11789_ ;
	wire _w11788_ ;
	wire _w11787_ ;
	wire _w11786_ ;
	wire _w11785_ ;
	wire _w11784_ ;
	wire _w11783_ ;
	wire _w11782_ ;
	wire _w11781_ ;
	wire _w11780_ ;
	wire _w11779_ ;
	wire _w11778_ ;
	wire _w11777_ ;
	wire _w11776_ ;
	wire _w11775_ ;
	wire _w11774_ ;
	wire _w11773_ ;
	wire _w11772_ ;
	wire _w11771_ ;
	wire _w11770_ ;
	wire _w11769_ ;
	wire _w11768_ ;
	wire _w11767_ ;
	wire _w11766_ ;
	wire _w11765_ ;
	wire _w11764_ ;
	wire _w11763_ ;
	wire _w11762_ ;
	wire _w11761_ ;
	wire _w11760_ ;
	wire _w11759_ ;
	wire _w11758_ ;
	wire _w11757_ ;
	wire _w11756_ ;
	wire _w11755_ ;
	wire _w11754_ ;
	wire _w11753_ ;
	wire _w11752_ ;
	wire _w11751_ ;
	wire _w11750_ ;
	wire _w11749_ ;
	wire _w11748_ ;
	wire _w11747_ ;
	wire _w11746_ ;
	wire _w11745_ ;
	wire _w11744_ ;
	wire _w11743_ ;
	wire _w11742_ ;
	wire _w11741_ ;
	wire _w11740_ ;
	wire _w11739_ ;
	wire _w11738_ ;
	wire _w11737_ ;
	wire _w11736_ ;
	wire _w11735_ ;
	wire _w11734_ ;
	wire _w11733_ ;
	wire _w11732_ ;
	wire _w11731_ ;
	wire _w11730_ ;
	wire _w11729_ ;
	wire _w11728_ ;
	wire _w11727_ ;
	wire _w11726_ ;
	wire _w11725_ ;
	wire _w11724_ ;
	wire _w11723_ ;
	wire _w11722_ ;
	wire _w11721_ ;
	wire _w11720_ ;
	wire _w11719_ ;
	wire _w11718_ ;
	wire _w11717_ ;
	wire _w11716_ ;
	wire _w11715_ ;
	wire _w11714_ ;
	wire _w11713_ ;
	wire _w11712_ ;
	wire _w11711_ ;
	wire _w11710_ ;
	wire _w11709_ ;
	wire _w11708_ ;
	wire _w11707_ ;
	wire _w11706_ ;
	wire _w11705_ ;
	wire _w11704_ ;
	wire _w11703_ ;
	wire _w11702_ ;
	wire _w11701_ ;
	wire _w11700_ ;
	wire _w11699_ ;
	wire _w11698_ ;
	wire _w11697_ ;
	wire _w11696_ ;
	wire _w11695_ ;
	wire _w11694_ ;
	wire _w11693_ ;
	wire _w11692_ ;
	wire _w11691_ ;
	wire _w11690_ ;
	wire _w11689_ ;
	wire _w11688_ ;
	wire _w11687_ ;
	wire _w11686_ ;
	wire _w11685_ ;
	wire _w11684_ ;
	wire _w11683_ ;
	wire _w11682_ ;
	wire _w11681_ ;
	wire _w11680_ ;
	wire _w11679_ ;
	wire _w11678_ ;
	wire _w11677_ ;
	wire _w11676_ ;
	wire _w11675_ ;
	wire _w11674_ ;
	wire _w11673_ ;
	wire _w11672_ ;
	wire _w11671_ ;
	wire _w11670_ ;
	wire _w11669_ ;
	wire _w11668_ ;
	wire _w11667_ ;
	wire _w11666_ ;
	wire _w11665_ ;
	wire _w11664_ ;
	wire _w11663_ ;
	wire _w11662_ ;
	wire _w11661_ ;
	wire _w11660_ ;
	wire _w11659_ ;
	wire _w11658_ ;
	wire _w11657_ ;
	wire _w11656_ ;
	wire _w11655_ ;
	wire _w11654_ ;
	wire _w11653_ ;
	wire _w11652_ ;
	wire _w11651_ ;
	wire _w11650_ ;
	wire _w11649_ ;
	wire _w11648_ ;
	wire _w11647_ ;
	wire _w11646_ ;
	wire _w11645_ ;
	wire _w11644_ ;
	wire _w11643_ ;
	wire _w11642_ ;
	wire _w11641_ ;
	wire _w11640_ ;
	wire _w11639_ ;
	wire _w11638_ ;
	wire _w11637_ ;
	wire _w11636_ ;
	wire _w11635_ ;
	wire _w11634_ ;
	wire _w11633_ ;
	wire _w11632_ ;
	wire _w11631_ ;
	wire _w11630_ ;
	wire _w11629_ ;
	wire _w11628_ ;
	wire _w11627_ ;
	wire _w11626_ ;
	wire _w11625_ ;
	wire _w11624_ ;
	wire _w11623_ ;
	wire _w11622_ ;
	wire _w11621_ ;
	wire _w11620_ ;
	wire _w11619_ ;
	wire _w11618_ ;
	wire _w11617_ ;
	wire _w11616_ ;
	wire _w11615_ ;
	wire _w11614_ ;
	wire _w11613_ ;
	wire _w11612_ ;
	wire _w11611_ ;
	wire _w11610_ ;
	wire _w11609_ ;
	wire _w11608_ ;
	wire _w11607_ ;
	wire _w11606_ ;
	wire _w11605_ ;
	wire _w11604_ ;
	wire _w11603_ ;
	wire _w11602_ ;
	wire _w11601_ ;
	wire _w11600_ ;
	wire _w11599_ ;
	wire _w11598_ ;
	wire _w11597_ ;
	wire _w11596_ ;
	wire _w11595_ ;
	wire _w11594_ ;
	wire _w11593_ ;
	wire _w11592_ ;
	wire _w11591_ ;
	wire _w11590_ ;
	wire _w11589_ ;
	wire _w11588_ ;
	wire _w11587_ ;
	wire _w11586_ ;
	wire _w11585_ ;
	wire _w11584_ ;
	wire _w11583_ ;
	wire _w11582_ ;
	wire _w11581_ ;
	wire _w11580_ ;
	wire _w11579_ ;
	wire _w11578_ ;
	wire _w11577_ ;
	wire _w11576_ ;
	wire _w11575_ ;
	wire _w11574_ ;
	wire _w11573_ ;
	wire _w11572_ ;
	wire _w11571_ ;
	wire _w11570_ ;
	wire _w11569_ ;
	wire _w11568_ ;
	wire _w11567_ ;
	wire _w11566_ ;
	wire _w11565_ ;
	wire _w11564_ ;
	wire _w11563_ ;
	wire _w11562_ ;
	wire _w11561_ ;
	wire _w11560_ ;
	wire _w11559_ ;
	wire _w11558_ ;
	wire _w11557_ ;
	wire _w11556_ ;
	wire _w11555_ ;
	wire _w11554_ ;
	wire _w11553_ ;
	wire _w11552_ ;
	wire _w11551_ ;
	wire _w11550_ ;
	wire _w11549_ ;
	wire _w11548_ ;
	wire _w11547_ ;
	wire _w11546_ ;
	wire _w11545_ ;
	wire _w11544_ ;
	wire _w11543_ ;
	wire _w11542_ ;
	wire _w11541_ ;
	wire _w11540_ ;
	wire _w11539_ ;
	wire _w11538_ ;
	wire _w11537_ ;
	wire _w11536_ ;
	wire _w11535_ ;
	wire _w11534_ ;
	wire _w11533_ ;
	wire _w11532_ ;
	wire _w11531_ ;
	wire _w11530_ ;
	wire _w11529_ ;
	wire _w11528_ ;
	wire _w11527_ ;
	wire _w11526_ ;
	wire _w11525_ ;
	wire _w11524_ ;
	wire _w11523_ ;
	wire _w11522_ ;
	wire _w11521_ ;
	wire _w11520_ ;
	wire _w11519_ ;
	wire _w11518_ ;
	wire _w11517_ ;
	wire _w11516_ ;
	wire _w11515_ ;
	wire _w11514_ ;
	wire _w11513_ ;
	wire _w11512_ ;
	wire _w11511_ ;
	wire _w11510_ ;
	wire _w11509_ ;
	wire _w11508_ ;
	wire _w11507_ ;
	wire _w11506_ ;
	wire _w11505_ ;
	wire _w11504_ ;
	wire _w11503_ ;
	wire _w11502_ ;
	wire _w11501_ ;
	wire _w11500_ ;
	wire _w11499_ ;
	wire _w11498_ ;
	wire _w11497_ ;
	wire _w11496_ ;
	wire _w11495_ ;
	wire _w11494_ ;
	wire _w11493_ ;
	wire _w11492_ ;
	wire _w11491_ ;
	wire _w11490_ ;
	wire _w11489_ ;
	wire _w11488_ ;
	wire _w11487_ ;
	wire _w11486_ ;
	wire _w11485_ ;
	wire _w11484_ ;
	wire _w11483_ ;
	wire _w11482_ ;
	wire _w11481_ ;
	wire _w11480_ ;
	wire _w11479_ ;
	wire _w11478_ ;
	wire _w11477_ ;
	wire _w11476_ ;
	wire _w11475_ ;
	wire _w11474_ ;
	wire _w11473_ ;
	wire _w11472_ ;
	wire _w11471_ ;
	wire _w11470_ ;
	wire _w11469_ ;
	wire _w11468_ ;
	wire _w11467_ ;
	wire _w11466_ ;
	wire _w11465_ ;
	wire _w11464_ ;
	wire _w11463_ ;
	wire _w11462_ ;
	wire _w11461_ ;
	wire _w11460_ ;
	wire _w11459_ ;
	wire _w11458_ ;
	wire _w11457_ ;
	wire _w11456_ ;
	wire _w11455_ ;
	wire _w11454_ ;
	wire _w11453_ ;
	wire _w11452_ ;
	wire _w11451_ ;
	wire _w11450_ ;
	wire _w11449_ ;
	wire _w11448_ ;
	wire _w11447_ ;
	wire _w11446_ ;
	wire _w11445_ ;
	wire _w11444_ ;
	wire _w11443_ ;
	wire _w11442_ ;
	wire _w11441_ ;
	wire _w11440_ ;
	wire _w11439_ ;
	wire _w11438_ ;
	wire _w11437_ ;
	wire _w11436_ ;
	wire _w11435_ ;
	wire _w11434_ ;
	wire _w11433_ ;
	wire _w11432_ ;
	wire _w11431_ ;
	wire _w11430_ ;
	wire _w11429_ ;
	wire _w11428_ ;
	wire _w11427_ ;
	wire _w11426_ ;
	wire _w11425_ ;
	wire _w11424_ ;
	wire _w11423_ ;
	wire _w11422_ ;
	wire _w11421_ ;
	wire _w11420_ ;
	wire _w11419_ ;
	wire _w11418_ ;
	wire _w11417_ ;
	wire _w11416_ ;
	wire _w11415_ ;
	wire _w11414_ ;
	wire _w11413_ ;
	wire _w11412_ ;
	wire _w11411_ ;
	wire _w11410_ ;
	wire _w11409_ ;
	wire _w11408_ ;
	wire _w11407_ ;
	wire _w11406_ ;
	wire _w11405_ ;
	wire _w11404_ ;
	wire _w11403_ ;
	wire _w11402_ ;
	wire _w11401_ ;
	wire _w11400_ ;
	wire _w11399_ ;
	wire _w11398_ ;
	wire _w11397_ ;
	wire _w11396_ ;
	wire _w11395_ ;
	wire _w11394_ ;
	wire _w11393_ ;
	wire _w11392_ ;
	wire _w11391_ ;
	wire _w11390_ ;
	wire _w11389_ ;
	wire _w11388_ ;
	wire _w11387_ ;
	wire _w11386_ ;
	wire _w11385_ ;
	wire _w11384_ ;
	wire _w11383_ ;
	wire _w11382_ ;
	wire _w11381_ ;
	wire _w11380_ ;
	wire _w11379_ ;
	wire _w11378_ ;
	wire _w11377_ ;
	wire _w11376_ ;
	wire _w11375_ ;
	wire _w11374_ ;
	wire _w11373_ ;
	wire _w11372_ ;
	wire _w11371_ ;
	wire _w11370_ ;
	wire _w11369_ ;
	wire _w11368_ ;
	wire _w11367_ ;
	wire _w11366_ ;
	wire _w11365_ ;
	wire _w11364_ ;
	wire _w11363_ ;
	wire _w11362_ ;
	wire _w11361_ ;
	wire _w11360_ ;
	wire _w11359_ ;
	wire _w11358_ ;
	wire _w11357_ ;
	wire _w11356_ ;
	wire _w11355_ ;
	wire _w11354_ ;
	wire _w11353_ ;
	wire _w11352_ ;
	wire _w11351_ ;
	wire _w11350_ ;
	wire _w11349_ ;
	wire _w11348_ ;
	wire _w11347_ ;
	wire _w11346_ ;
	wire _w11345_ ;
	wire _w11344_ ;
	wire _w11343_ ;
	wire _w11342_ ;
	wire _w11341_ ;
	wire _w11340_ ;
	wire _w11339_ ;
	wire _w11338_ ;
	wire _w11337_ ;
	wire _w11336_ ;
	wire _w11335_ ;
	wire _w11334_ ;
	wire _w11333_ ;
	wire _w11332_ ;
	wire _w11331_ ;
	wire _w11330_ ;
	wire _w11329_ ;
	wire _w11328_ ;
	wire _w11327_ ;
	wire _w11326_ ;
	wire _w11325_ ;
	wire _w11324_ ;
	wire _w11323_ ;
	wire _w11322_ ;
	wire _w11321_ ;
	wire _w11320_ ;
	wire _w11319_ ;
	wire _w11318_ ;
	wire _w11317_ ;
	wire _w11316_ ;
	wire _w11315_ ;
	wire _w11314_ ;
	wire _w11313_ ;
	wire _w11312_ ;
	wire _w11311_ ;
	wire _w11310_ ;
	wire _w11309_ ;
	wire _w11308_ ;
	wire _w11307_ ;
	wire _w11306_ ;
	wire _w11305_ ;
	wire _w11304_ ;
	wire _w11303_ ;
	wire _w11302_ ;
	wire _w11301_ ;
	wire _w11300_ ;
	wire _w11299_ ;
	wire _w11298_ ;
	wire _w11297_ ;
	wire _w11296_ ;
	wire _w11295_ ;
	wire _w11294_ ;
	wire _w11293_ ;
	wire _w11292_ ;
	wire _w11291_ ;
	wire _w11290_ ;
	wire _w11289_ ;
	wire _w11288_ ;
	wire _w11287_ ;
	wire _w11286_ ;
	wire _w11285_ ;
	wire _w11284_ ;
	wire _w11283_ ;
	wire _w11282_ ;
	wire _w11281_ ;
	wire _w11280_ ;
	wire _w11279_ ;
	wire _w11278_ ;
	wire _w11277_ ;
	wire _w11276_ ;
	wire _w11275_ ;
	wire _w11274_ ;
	wire _w11273_ ;
	wire _w11272_ ;
	wire _w11271_ ;
	wire _w11270_ ;
	wire _w11269_ ;
	wire _w11268_ ;
	wire _w11267_ ;
	wire _w11266_ ;
	wire _w11265_ ;
	wire _w11264_ ;
	wire _w11263_ ;
	wire _w11262_ ;
	wire _w11261_ ;
	wire _w11260_ ;
	wire _w11259_ ;
	wire _w11258_ ;
	wire _w11257_ ;
	wire _w11256_ ;
	wire _w11255_ ;
	wire _w11254_ ;
	wire _w11253_ ;
	wire _w11252_ ;
	wire _w11251_ ;
	wire _w11250_ ;
	wire _w11249_ ;
	wire _w11248_ ;
	wire _w11247_ ;
	wire _w11246_ ;
	wire _w11245_ ;
	wire _w11244_ ;
	wire _w11243_ ;
	wire _w11242_ ;
	wire _w11241_ ;
	wire _w11240_ ;
	wire _w11239_ ;
	wire _w11238_ ;
	wire _w11237_ ;
	wire _w11236_ ;
	wire _w11235_ ;
	wire _w11234_ ;
	wire _w11233_ ;
	wire _w11232_ ;
	wire _w11231_ ;
	wire _w11230_ ;
	wire _w11229_ ;
	wire _w11228_ ;
	wire _w11227_ ;
	wire _w11226_ ;
	wire _w11225_ ;
	wire _w11224_ ;
	wire _w11223_ ;
	wire _w11222_ ;
	wire _w11221_ ;
	wire _w11220_ ;
	wire _w11219_ ;
	wire _w11218_ ;
	wire _w11217_ ;
	wire _w11216_ ;
	wire _w11215_ ;
	wire _w11214_ ;
	wire _w11213_ ;
	wire _w11212_ ;
	wire _w11211_ ;
	wire _w11210_ ;
	wire _w11209_ ;
	wire _w11208_ ;
	wire _w11207_ ;
	wire _w11206_ ;
	wire _w11205_ ;
	wire _w11204_ ;
	wire _w11203_ ;
	wire _w11202_ ;
	wire _w11201_ ;
	wire _w11200_ ;
	wire _w11199_ ;
	wire _w11198_ ;
	wire _w11197_ ;
	wire _w11196_ ;
	wire _w11195_ ;
	wire _w11194_ ;
	wire _w11193_ ;
	wire _w11192_ ;
	wire _w11191_ ;
	wire _w11190_ ;
	wire _w11189_ ;
	wire _w11188_ ;
	wire _w11187_ ;
	wire _w11186_ ;
	wire _w11185_ ;
	wire _w11184_ ;
	wire _w11183_ ;
	wire _w11182_ ;
	wire _w11181_ ;
	wire _w11180_ ;
	wire _w11179_ ;
	wire _w11178_ ;
	wire _w11177_ ;
	wire _w11176_ ;
	wire _w11175_ ;
	wire _w11174_ ;
	wire _w11173_ ;
	wire _w11172_ ;
	wire _w11171_ ;
	wire _w11170_ ;
	wire _w11169_ ;
	wire _w11168_ ;
	wire _w11167_ ;
	wire _w11166_ ;
	wire _w11165_ ;
	wire _w11164_ ;
	wire _w11163_ ;
	wire _w11162_ ;
	wire _w11161_ ;
	wire _w11160_ ;
	wire _w11159_ ;
	wire _w11158_ ;
	wire _w11157_ ;
	wire _w11156_ ;
	wire _w11155_ ;
	wire _w11154_ ;
	wire _w11153_ ;
	wire _w11152_ ;
	wire _w11151_ ;
	wire _w11150_ ;
	wire _w11149_ ;
	wire _w11148_ ;
	wire _w11147_ ;
	wire _w11146_ ;
	wire _w11145_ ;
	wire _w11144_ ;
	wire _w11143_ ;
	wire _w11142_ ;
	wire _w11141_ ;
	wire _w11140_ ;
	wire _w11139_ ;
	wire _w11138_ ;
	wire _w11137_ ;
	wire _w11136_ ;
	wire _w11135_ ;
	wire _w11134_ ;
	wire _w11133_ ;
	wire _w11132_ ;
	wire _w11131_ ;
	wire _w11130_ ;
	wire _w11129_ ;
	wire _w11128_ ;
	wire _w11127_ ;
	wire _w11126_ ;
	wire _w11125_ ;
	wire _w11124_ ;
	wire _w11123_ ;
	wire _w11122_ ;
	wire _w11121_ ;
	wire _w11120_ ;
	wire _w11119_ ;
	wire _w11118_ ;
	wire _w11117_ ;
	wire _w11116_ ;
	wire _w11115_ ;
	wire _w11114_ ;
	wire _w11113_ ;
	wire _w11112_ ;
	wire _w11111_ ;
	wire _w11110_ ;
	wire _w11109_ ;
	wire _w11108_ ;
	wire _w11107_ ;
	wire _w11106_ ;
	wire _w11105_ ;
	wire _w11104_ ;
	wire _w11103_ ;
	wire _w11102_ ;
	wire _w11101_ ;
	wire _w11100_ ;
	wire _w11099_ ;
	wire _w11098_ ;
	wire _w11097_ ;
	wire _w11096_ ;
	wire _w11095_ ;
	wire _w11094_ ;
	wire _w11093_ ;
	wire _w11092_ ;
	wire _w11091_ ;
	wire _w11090_ ;
	wire _w11089_ ;
	wire _w11088_ ;
	wire _w11087_ ;
	wire _w11086_ ;
	wire _w11085_ ;
	wire _w11084_ ;
	wire _w11083_ ;
	wire _w11082_ ;
	wire _w11081_ ;
	wire _w11080_ ;
	wire _w11079_ ;
	wire _w11078_ ;
	wire _w11077_ ;
	wire _w11076_ ;
	wire _w11075_ ;
	wire _w11074_ ;
	wire _w11073_ ;
	wire _w11072_ ;
	wire _w11071_ ;
	wire _w11070_ ;
	wire _w11069_ ;
	wire _w11068_ ;
	wire _w11067_ ;
	wire _w11066_ ;
	wire _w11065_ ;
	wire _w11064_ ;
	wire _w11063_ ;
	wire _w11062_ ;
	wire _w11061_ ;
	wire _w11060_ ;
	wire _w11059_ ;
	wire _w11058_ ;
	wire _w11057_ ;
	wire _w11056_ ;
	wire _w11055_ ;
	wire _w11054_ ;
	wire _w11053_ ;
	wire _w11052_ ;
	wire _w11051_ ;
	wire _w11050_ ;
	wire _w11049_ ;
	wire _w11048_ ;
	wire _w11047_ ;
	wire _w11046_ ;
	wire _w11045_ ;
	wire _w11044_ ;
	wire _w11043_ ;
	wire _w11042_ ;
	wire _w11041_ ;
	wire _w11040_ ;
	wire _w11039_ ;
	wire _w11038_ ;
	wire _w11037_ ;
	wire _w11036_ ;
	wire _w11035_ ;
	wire _w11034_ ;
	wire _w11033_ ;
	wire _w11032_ ;
	wire _w11031_ ;
	wire _w11030_ ;
	wire _w11029_ ;
	wire _w11028_ ;
	wire _w11027_ ;
	wire _w11026_ ;
	wire _w11025_ ;
	wire _w11024_ ;
	wire _w11023_ ;
	wire _w11022_ ;
	wire _w11021_ ;
	wire _w11020_ ;
	wire _w11019_ ;
	wire _w11018_ ;
	wire _w11017_ ;
	wire _w11016_ ;
	wire _w11015_ ;
	wire _w11014_ ;
	wire _w11013_ ;
	wire _w11012_ ;
	wire _w11011_ ;
	wire _w11010_ ;
	wire _w11009_ ;
	wire _w11008_ ;
	wire _w11007_ ;
	wire _w11006_ ;
	wire _w11005_ ;
	wire _w11004_ ;
	wire _w11003_ ;
	wire _w11002_ ;
	wire _w11001_ ;
	wire _w11000_ ;
	wire _w10999_ ;
	wire _w10998_ ;
	wire _w10997_ ;
	wire _w10996_ ;
	wire _w10995_ ;
	wire _w10994_ ;
	wire _w10993_ ;
	wire _w10992_ ;
	wire _w10991_ ;
	wire _w10990_ ;
	wire _w10989_ ;
	wire _w10988_ ;
	wire _w10987_ ;
	wire _w10986_ ;
	wire _w10985_ ;
	wire _w10984_ ;
	wire _w10983_ ;
	wire _w10982_ ;
	wire _w10981_ ;
	wire _w10980_ ;
	wire _w10979_ ;
	wire _w10978_ ;
	wire _w10977_ ;
	wire _w10976_ ;
	wire _w10975_ ;
	wire _w10974_ ;
	wire _w10973_ ;
	wire _w10972_ ;
	wire _w10971_ ;
	wire _w10970_ ;
	wire _w10969_ ;
	wire _w10968_ ;
	wire _w10967_ ;
	wire _w10966_ ;
	wire _w10965_ ;
	wire _w10964_ ;
	wire _w10963_ ;
	wire _w10962_ ;
	wire _w10961_ ;
	wire _w10960_ ;
	wire _w10959_ ;
	wire _w10958_ ;
	wire _w10957_ ;
	wire _w10956_ ;
	wire _w10955_ ;
	wire _w10954_ ;
	wire _w10953_ ;
	wire _w10952_ ;
	wire _w10951_ ;
	wire _w10950_ ;
	wire _w10949_ ;
	wire _w10948_ ;
	wire _w10947_ ;
	wire _w10946_ ;
	wire _w10945_ ;
	wire _w10944_ ;
	wire _w10943_ ;
	wire _w10942_ ;
	wire _w10941_ ;
	wire _w10940_ ;
	wire _w10939_ ;
	wire _w10938_ ;
	wire _w10937_ ;
	wire _w10936_ ;
	wire _w10935_ ;
	wire _w10934_ ;
	wire _w10933_ ;
	wire _w10932_ ;
	wire _w10931_ ;
	wire _w10930_ ;
	wire _w10929_ ;
	wire _w10928_ ;
	wire _w10927_ ;
	wire _w10926_ ;
	wire _w10925_ ;
	wire _w10924_ ;
	wire _w10923_ ;
	wire _w10922_ ;
	wire _w10921_ ;
	wire _w10920_ ;
	wire _w10919_ ;
	wire _w10918_ ;
	wire _w10917_ ;
	wire _w10916_ ;
	wire _w10915_ ;
	wire _w10914_ ;
	wire _w10913_ ;
	wire _w10912_ ;
	wire _w10911_ ;
	wire _w10910_ ;
	wire _w10909_ ;
	wire _w10908_ ;
	wire _w10907_ ;
	wire _w10906_ ;
	wire _w10905_ ;
	wire _w10904_ ;
	wire _w10903_ ;
	wire _w10902_ ;
	wire _w10901_ ;
	wire _w10900_ ;
	wire _w10899_ ;
	wire _w10898_ ;
	wire _w10897_ ;
	wire _w10896_ ;
	wire _w10895_ ;
	wire _w10894_ ;
	wire _w10893_ ;
	wire _w10892_ ;
	wire _w10891_ ;
	wire _w10890_ ;
	wire _w10889_ ;
	wire _w10888_ ;
	wire _w10887_ ;
	wire _w10886_ ;
	wire _w10885_ ;
	wire _w10884_ ;
	wire _w10883_ ;
	wire _w10882_ ;
	wire _w10881_ ;
	wire _w10880_ ;
	wire _w10879_ ;
	wire _w10878_ ;
	wire _w10877_ ;
	wire _w10876_ ;
	wire _w10875_ ;
	wire _w10874_ ;
	wire _w10873_ ;
	wire _w10872_ ;
	wire _w10871_ ;
	wire _w10870_ ;
	wire _w10869_ ;
	wire _w10868_ ;
	wire _w10867_ ;
	wire _w10866_ ;
	wire _w10865_ ;
	wire _w10864_ ;
	wire _w10863_ ;
	wire _w10862_ ;
	wire _w10861_ ;
	wire _w10860_ ;
	wire _w10859_ ;
	wire _w10858_ ;
	wire _w10857_ ;
	wire _w10856_ ;
	wire _w10855_ ;
	wire _w10854_ ;
	wire _w10853_ ;
	wire _w10852_ ;
	wire _w10851_ ;
	wire _w10850_ ;
	wire _w10849_ ;
	wire _w10848_ ;
	wire _w10847_ ;
	wire _w10846_ ;
	wire _w10845_ ;
	wire _w10844_ ;
	wire _w10843_ ;
	wire _w10842_ ;
	wire _w10841_ ;
	wire _w10840_ ;
	wire _w10839_ ;
	wire _w10838_ ;
	wire _w10837_ ;
	wire _w10836_ ;
	wire _w10835_ ;
	wire _w10834_ ;
	wire _w10833_ ;
	wire _w10832_ ;
	wire _w10831_ ;
	wire _w10830_ ;
	wire _w10829_ ;
	wire _w10828_ ;
	wire _w10827_ ;
	wire _w10826_ ;
	wire _w10825_ ;
	wire _w10824_ ;
	wire _w10823_ ;
	wire _w10822_ ;
	wire _w10821_ ;
	wire _w10820_ ;
	wire _w10819_ ;
	wire _w10818_ ;
	wire _w10817_ ;
	wire _w10816_ ;
	wire _w10815_ ;
	wire _w10814_ ;
	wire _w10813_ ;
	wire _w10812_ ;
	wire _w10811_ ;
	wire _w10810_ ;
	wire _w10809_ ;
	wire _w10808_ ;
	wire _w10807_ ;
	wire _w10806_ ;
	wire _w10805_ ;
	wire _w10804_ ;
	wire _w10803_ ;
	wire _w10802_ ;
	wire _w10801_ ;
	wire _w10800_ ;
	wire _w10799_ ;
	wire _w10798_ ;
	wire _w10797_ ;
	wire _w10796_ ;
	wire _w10795_ ;
	wire _w10794_ ;
	wire _w10793_ ;
	wire _w10792_ ;
	wire _w10791_ ;
	wire _w10790_ ;
	wire _w10789_ ;
	wire _w10788_ ;
	wire _w10787_ ;
	wire _w10786_ ;
	wire _w10785_ ;
	wire _w10784_ ;
	wire _w10783_ ;
	wire _w10782_ ;
	wire _w10781_ ;
	wire _w10780_ ;
	wire _w10779_ ;
	wire _w10778_ ;
	wire _w10777_ ;
	wire _w10776_ ;
	wire _w10775_ ;
	wire _w10774_ ;
	wire _w10773_ ;
	wire _w10772_ ;
	wire _w10771_ ;
	wire _w10770_ ;
	wire _w10769_ ;
	wire _w10768_ ;
	wire _w10767_ ;
	wire _w10766_ ;
	wire _w10765_ ;
	wire _w10764_ ;
	wire _w10763_ ;
	wire _w10762_ ;
	wire _w10761_ ;
	wire _w10760_ ;
	wire _w10759_ ;
	wire _w10758_ ;
	wire _w10757_ ;
	wire _w10756_ ;
	wire _w10755_ ;
	wire _w10754_ ;
	wire _w10753_ ;
	wire _w10752_ ;
	wire _w10751_ ;
	wire _w10750_ ;
	wire _w10749_ ;
	wire _w10748_ ;
	wire _w10747_ ;
	wire _w10746_ ;
	wire _w10745_ ;
	wire _w10744_ ;
	wire _w10743_ ;
	wire _w10742_ ;
	wire _w10741_ ;
	wire _w10740_ ;
	wire _w10739_ ;
	wire _w10738_ ;
	wire _w10737_ ;
	wire _w10736_ ;
	wire _w10735_ ;
	wire _w10734_ ;
	wire _w10733_ ;
	wire _w10732_ ;
	wire _w10731_ ;
	wire _w10730_ ;
	wire _w10729_ ;
	wire _w10728_ ;
	wire _w10727_ ;
	wire _w10726_ ;
	wire _w10725_ ;
	wire _w10724_ ;
	wire _w10723_ ;
	wire _w10722_ ;
	wire _w10721_ ;
	wire _w10720_ ;
	wire _w10719_ ;
	wire _w10718_ ;
	wire _w10717_ ;
	wire _w10716_ ;
	wire _w10715_ ;
	wire _w10714_ ;
	wire _w10713_ ;
	wire _w10712_ ;
	wire _w10711_ ;
	wire _w10710_ ;
	wire _w10709_ ;
	wire _w10708_ ;
	wire _w10707_ ;
	wire _w10706_ ;
	wire _w10705_ ;
	wire _w10704_ ;
	wire _w10703_ ;
	wire _w10702_ ;
	wire _w10701_ ;
	wire _w10700_ ;
	wire _w10699_ ;
	wire _w10698_ ;
	wire _w10697_ ;
	wire _w10696_ ;
	wire _w10695_ ;
	wire _w10694_ ;
	wire _w10693_ ;
	wire _w10692_ ;
	wire _w10691_ ;
	wire _w10690_ ;
	wire _w10689_ ;
	wire _w10688_ ;
	wire _w10687_ ;
	wire _w10686_ ;
	wire _w10685_ ;
	wire _w10684_ ;
	wire _w10683_ ;
	wire _w10682_ ;
	wire _w10681_ ;
	wire _w10680_ ;
	wire _w10679_ ;
	wire _w10678_ ;
	wire _w10677_ ;
	wire _w10676_ ;
	wire _w10675_ ;
	wire _w10674_ ;
	wire _w10673_ ;
	wire _w10672_ ;
	wire _w10671_ ;
	wire _w10670_ ;
	wire _w10669_ ;
	wire _w10668_ ;
	wire _w10667_ ;
	wire _w10666_ ;
	wire _w10665_ ;
	wire _w10664_ ;
	wire _w10663_ ;
	wire _w10662_ ;
	wire _w10661_ ;
	wire _w10660_ ;
	wire _w10659_ ;
	wire _w10658_ ;
	wire _w10657_ ;
	wire _w10656_ ;
	wire _w10655_ ;
	wire _w10654_ ;
	wire _w10653_ ;
	wire _w10652_ ;
	wire _w10651_ ;
	wire _w10650_ ;
	wire _w10649_ ;
	wire _w10648_ ;
	wire _w10647_ ;
	wire _w10646_ ;
	wire _w10645_ ;
	wire _w10644_ ;
	wire _w10643_ ;
	wire _w10642_ ;
	wire _w10641_ ;
	wire _w10640_ ;
	wire _w10639_ ;
	wire _w10638_ ;
	wire _w10637_ ;
	wire _w10636_ ;
	wire _w10635_ ;
	wire _w10634_ ;
	wire _w10633_ ;
	wire _w10632_ ;
	wire _w10631_ ;
	wire _w10630_ ;
	wire _w10629_ ;
	wire _w10628_ ;
	wire _w10627_ ;
	wire _w10626_ ;
	wire _w10625_ ;
	wire _w10624_ ;
	wire _w10623_ ;
	wire _w10622_ ;
	wire _w10621_ ;
	wire _w10620_ ;
	wire _w10619_ ;
	wire _w10618_ ;
	wire _w10617_ ;
	wire _w10616_ ;
	wire _w10615_ ;
	wire _w10614_ ;
	wire _w10613_ ;
	wire _w10612_ ;
	wire _w10611_ ;
	wire _w10610_ ;
	wire _w10609_ ;
	wire _w10608_ ;
	wire _w10607_ ;
	wire _w10606_ ;
	wire _w10605_ ;
	wire _w10604_ ;
	wire _w10603_ ;
	wire _w10602_ ;
	wire _w10601_ ;
	wire _w10600_ ;
	wire _w10599_ ;
	wire _w10598_ ;
	wire _w10597_ ;
	wire _w10596_ ;
	wire _w10595_ ;
	wire _w10594_ ;
	wire _w10593_ ;
	wire _w10592_ ;
	wire _w10591_ ;
	wire _w10590_ ;
	wire _w10589_ ;
	wire _w10588_ ;
	wire _w10587_ ;
	wire _w10586_ ;
	wire _w10585_ ;
	wire _w10584_ ;
	wire _w10583_ ;
	wire _w10582_ ;
	wire _w10581_ ;
	wire _w10580_ ;
	wire _w10579_ ;
	wire _w10578_ ;
	wire _w10577_ ;
	wire _w10576_ ;
	wire _w10575_ ;
	wire _w10574_ ;
	wire _w10573_ ;
	wire _w10572_ ;
	wire _w10571_ ;
	wire _w10570_ ;
	wire _w10569_ ;
	wire _w10568_ ;
	wire _w10567_ ;
	wire _w10566_ ;
	wire _w10565_ ;
	wire _w10564_ ;
	wire _w10563_ ;
	wire _w10562_ ;
	wire _w10561_ ;
	wire _w10560_ ;
	wire _w10559_ ;
	wire _w10558_ ;
	wire _w10557_ ;
	wire _w10556_ ;
	wire _w10555_ ;
	wire _w10554_ ;
	wire _w10553_ ;
	wire _w10552_ ;
	wire _w10551_ ;
	wire _w10550_ ;
	wire _w10549_ ;
	wire _w10548_ ;
	wire _w10547_ ;
	wire _w10546_ ;
	wire _w10545_ ;
	wire _w10544_ ;
	wire _w10543_ ;
	wire _w10542_ ;
	wire _w10541_ ;
	wire _w10540_ ;
	wire _w10539_ ;
	wire _w10538_ ;
	wire _w10537_ ;
	wire _w10536_ ;
	wire _w10535_ ;
	wire _w10534_ ;
	wire _w10533_ ;
	wire _w10532_ ;
	wire _w10531_ ;
	wire _w10530_ ;
	wire _w10529_ ;
	wire _w10528_ ;
	wire _w10527_ ;
	wire _w10526_ ;
	wire _w10525_ ;
	wire _w10524_ ;
	wire _w10523_ ;
	wire _w10522_ ;
	wire _w10521_ ;
	wire _w10520_ ;
	wire _w10519_ ;
	wire _w10518_ ;
	wire _w10517_ ;
	wire _w10516_ ;
	wire _w10515_ ;
	wire _w10514_ ;
	wire _w10513_ ;
	wire _w10512_ ;
	wire _w10511_ ;
	wire _w10510_ ;
	wire _w10509_ ;
	wire _w10508_ ;
	wire _w10507_ ;
	wire _w10506_ ;
	wire _w10505_ ;
	wire _w10504_ ;
	wire _w10503_ ;
	wire _w10502_ ;
	wire _w10501_ ;
	wire _w10500_ ;
	wire _w10499_ ;
	wire _w10498_ ;
	wire _w10497_ ;
	wire _w10496_ ;
	wire _w10495_ ;
	wire _w10494_ ;
	wire _w10493_ ;
	wire _w10492_ ;
	wire _w10491_ ;
	wire _w10490_ ;
	wire _w10489_ ;
	wire _w10488_ ;
	wire _w10487_ ;
	wire _w10486_ ;
	wire _w10485_ ;
	wire _w10484_ ;
	wire _w10483_ ;
	wire _w10482_ ;
	wire _w10481_ ;
	wire _w10480_ ;
	wire _w10479_ ;
	wire _w10478_ ;
	wire _w10477_ ;
	wire _w10476_ ;
	wire _w10475_ ;
	wire _w10474_ ;
	wire _w10473_ ;
	wire _w10472_ ;
	wire _w10471_ ;
	wire _w10470_ ;
	wire _w10469_ ;
	wire _w10468_ ;
	wire _w10467_ ;
	wire _w10466_ ;
	wire _w10465_ ;
	wire _w10464_ ;
	wire _w10463_ ;
	wire _w10462_ ;
	wire _w10461_ ;
	wire _w10460_ ;
	wire _w10459_ ;
	wire _w10458_ ;
	wire _w10457_ ;
	wire _w10456_ ;
	wire _w10455_ ;
	wire _w10454_ ;
	wire _w10453_ ;
	wire _w10452_ ;
	wire _w10451_ ;
	wire _w10450_ ;
	wire _w10449_ ;
	wire _w10448_ ;
	wire _w10447_ ;
	wire _w10446_ ;
	wire _w10445_ ;
	wire _w10444_ ;
	wire _w10443_ ;
	wire _w10442_ ;
	wire _w10441_ ;
	wire _w10440_ ;
	wire _w10439_ ;
	wire _w10438_ ;
	wire _w10437_ ;
	wire _w10436_ ;
	wire _w10435_ ;
	wire _w10434_ ;
	wire _w10433_ ;
	wire _w10432_ ;
	wire _w10431_ ;
	wire _w10430_ ;
	wire _w10429_ ;
	wire _w10428_ ;
	wire _w10427_ ;
	wire _w10426_ ;
	wire _w10425_ ;
	wire _w10424_ ;
	wire _w10423_ ;
	wire _w10422_ ;
	wire _w10421_ ;
	wire _w10420_ ;
	wire _w10419_ ;
	wire _w10418_ ;
	wire _w10417_ ;
	wire _w10416_ ;
	wire _w10415_ ;
	wire _w10414_ ;
	wire _w10413_ ;
	wire _w10412_ ;
	wire _w10411_ ;
	wire _w10410_ ;
	wire _w10409_ ;
	wire _w10408_ ;
	wire _w10407_ ;
	wire _w10406_ ;
	wire _w10405_ ;
	wire _w10404_ ;
	wire _w10403_ ;
	wire _w10402_ ;
	wire _w10401_ ;
	wire _w10400_ ;
	wire _w10399_ ;
	wire _w10398_ ;
	wire _w10397_ ;
	wire _w10396_ ;
	wire _w10395_ ;
	wire _w10394_ ;
	wire _w10393_ ;
	wire _w10392_ ;
	wire _w10391_ ;
	wire _w10390_ ;
	wire _w10389_ ;
	wire _w10388_ ;
	wire _w10387_ ;
	wire _w10386_ ;
	wire _w10385_ ;
	wire _w10384_ ;
	wire _w10383_ ;
	wire _w10382_ ;
	wire _w10381_ ;
	wire _w10380_ ;
	wire _w10379_ ;
	wire _w10378_ ;
	wire _w10377_ ;
	wire _w10376_ ;
	wire _w10375_ ;
	wire _w10374_ ;
	wire _w10373_ ;
	wire _w10372_ ;
	wire _w10371_ ;
	wire _w10370_ ;
	wire _w10369_ ;
	wire _w10368_ ;
	wire _w10367_ ;
	wire _w10366_ ;
	wire _w10365_ ;
	wire _w10364_ ;
	wire _w10363_ ;
	wire _w10362_ ;
	wire _w10361_ ;
	wire _w10360_ ;
	wire _w10359_ ;
	wire _w10358_ ;
	wire _w10357_ ;
	wire _w10356_ ;
	wire _w10355_ ;
	wire _w10354_ ;
	wire _w10353_ ;
	wire _w10352_ ;
	wire _w10351_ ;
	wire _w10350_ ;
	wire _w10349_ ;
	wire _w10348_ ;
	wire _w10347_ ;
	wire _w10346_ ;
	wire _w10345_ ;
	wire _w10344_ ;
	wire _w10343_ ;
	wire _w10342_ ;
	wire _w10341_ ;
	wire _w10340_ ;
	wire _w10339_ ;
	wire _w10338_ ;
	wire _w10337_ ;
	wire _w10336_ ;
	wire _w10335_ ;
	wire _w10334_ ;
	wire _w10333_ ;
	wire _w10332_ ;
	wire _w10331_ ;
	wire _w10330_ ;
	wire _w10329_ ;
	wire _w10328_ ;
	wire _w10327_ ;
	wire _w10326_ ;
	wire _w10325_ ;
	wire _w10324_ ;
	wire _w10323_ ;
	wire _w10322_ ;
	wire _w10321_ ;
	wire _w10320_ ;
	wire _w10319_ ;
	wire _w10318_ ;
	wire _w10317_ ;
	wire _w10316_ ;
	wire _w10315_ ;
	wire _w10314_ ;
	wire _w10313_ ;
	wire _w10312_ ;
	wire _w10311_ ;
	wire _w10310_ ;
	wire _w10309_ ;
	wire _w10308_ ;
	wire _w10307_ ;
	wire _w10306_ ;
	wire _w10305_ ;
	wire _w10304_ ;
	wire _w10303_ ;
	wire _w10302_ ;
	wire _w10301_ ;
	wire _w10300_ ;
	wire _w10299_ ;
	wire _w10298_ ;
	wire _w10297_ ;
	wire _w10296_ ;
	wire _w10295_ ;
	wire _w10294_ ;
	wire _w10293_ ;
	wire _w10292_ ;
	wire _w10291_ ;
	wire _w10290_ ;
	wire _w10289_ ;
	wire _w10288_ ;
	wire _w10287_ ;
	wire _w10286_ ;
	wire _w10285_ ;
	wire _w10284_ ;
	wire _w10283_ ;
	wire _w10282_ ;
	wire _w10281_ ;
	wire _w10280_ ;
	wire _w10279_ ;
	wire _w10278_ ;
	wire _w10277_ ;
	wire _w10276_ ;
	wire _w10275_ ;
	wire _w10274_ ;
	wire _w10273_ ;
	wire _w10272_ ;
	wire _w10271_ ;
	wire _w10270_ ;
	wire _w10269_ ;
	wire _w10268_ ;
	wire _w10267_ ;
	wire _w10266_ ;
	wire _w10265_ ;
	wire _w10264_ ;
	wire _w10263_ ;
	wire _w10262_ ;
	wire _w10261_ ;
	wire _w10260_ ;
	wire _w10259_ ;
	wire _w10258_ ;
	wire _w10257_ ;
	wire _w10256_ ;
	wire _w10255_ ;
	wire _w10254_ ;
	wire _w10253_ ;
	wire _w10252_ ;
	wire _w10251_ ;
	wire _w10250_ ;
	wire _w10249_ ;
	wire _w10248_ ;
	wire _w10247_ ;
	wire _w10246_ ;
	wire _w10245_ ;
	wire _w10244_ ;
	wire _w10243_ ;
	wire _w10242_ ;
	wire _w10241_ ;
	wire _w10240_ ;
	wire _w10239_ ;
	wire _w10238_ ;
	wire _w10237_ ;
	wire _w10236_ ;
	wire _w10235_ ;
	wire _w10234_ ;
	wire _w10233_ ;
	wire _w10232_ ;
	wire _w10231_ ;
	wire _w10230_ ;
	wire _w10229_ ;
	wire _w10228_ ;
	wire _w10227_ ;
	wire _w10226_ ;
	wire _w10225_ ;
	wire _w10224_ ;
	wire _w10223_ ;
	wire _w10222_ ;
	wire _w10221_ ;
	wire _w10220_ ;
	wire _w10219_ ;
	wire _w10218_ ;
	wire _w10217_ ;
	wire _w10216_ ;
	wire _w10215_ ;
	wire _w10214_ ;
	wire _w10213_ ;
	wire _w10212_ ;
	wire _w10211_ ;
	wire _w10210_ ;
	wire _w10209_ ;
	wire _w10208_ ;
	wire _w10207_ ;
	wire _w10206_ ;
	wire _w10205_ ;
	wire _w10204_ ;
	wire _w10203_ ;
	wire _w10202_ ;
	wire _w10201_ ;
	wire _w10200_ ;
	wire _w10199_ ;
	wire _w10198_ ;
	wire _w10197_ ;
	wire _w10196_ ;
	wire _w10195_ ;
	wire _w10194_ ;
	wire _w10193_ ;
	wire _w10192_ ;
	wire _w10191_ ;
	wire _w10190_ ;
	wire _w10189_ ;
	wire _w10188_ ;
	wire _w10187_ ;
	wire _w10186_ ;
	wire _w10185_ ;
	wire _w10184_ ;
	wire _w10183_ ;
	wire _w10182_ ;
	wire _w10181_ ;
	wire _w10180_ ;
	wire _w10179_ ;
	wire _w10178_ ;
	wire _w10177_ ;
	wire _w10176_ ;
	wire _w10175_ ;
	wire _w10174_ ;
	wire _w10173_ ;
	wire _w10172_ ;
	wire _w10171_ ;
	wire _w10170_ ;
	wire _w10169_ ;
	wire _w10168_ ;
	wire _w10167_ ;
	wire _w10166_ ;
	wire _w10165_ ;
	wire _w10164_ ;
	wire _w10163_ ;
	wire _w10162_ ;
	wire _w10161_ ;
	wire _w10160_ ;
	wire _w10159_ ;
	wire _w10158_ ;
	wire _w10157_ ;
	wire _w10156_ ;
	wire _w10155_ ;
	wire _w10154_ ;
	wire _w10153_ ;
	wire _w10152_ ;
	wire _w10151_ ;
	wire _w10150_ ;
	wire _w10149_ ;
	wire _w10148_ ;
	wire _w10147_ ;
	wire _w10146_ ;
	wire _w10145_ ;
	wire _w10144_ ;
	wire _w10143_ ;
	wire _w10142_ ;
	wire _w10141_ ;
	wire _w10140_ ;
	wire _w10139_ ;
	wire _w10138_ ;
	wire _w10137_ ;
	wire _w10136_ ;
	wire _w10135_ ;
	wire _w10134_ ;
	wire _w10133_ ;
	wire _w10132_ ;
	wire _w10131_ ;
	wire _w10130_ ;
	wire _w10129_ ;
	wire _w10128_ ;
	wire _w10127_ ;
	wire _w10126_ ;
	wire _w10125_ ;
	wire _w10124_ ;
	wire _w10123_ ;
	wire _w10122_ ;
	wire _w10121_ ;
	wire _w10120_ ;
	wire _w10119_ ;
	wire _w10118_ ;
	wire _w10117_ ;
	wire _w10116_ ;
	wire _w10115_ ;
	wire _w10114_ ;
	wire _w10113_ ;
	wire _w10112_ ;
	wire _w10111_ ;
	wire _w10110_ ;
	wire _w10109_ ;
	wire _w10108_ ;
	wire _w10107_ ;
	wire _w10106_ ;
	wire _w10105_ ;
	wire _w10104_ ;
	wire _w10103_ ;
	wire _w10102_ ;
	wire _w10101_ ;
	wire _w10100_ ;
	wire _w10099_ ;
	wire _w10098_ ;
	wire _w10097_ ;
	wire _w10096_ ;
	wire _w10095_ ;
	wire _w10094_ ;
	wire _w10093_ ;
	wire _w10092_ ;
	wire _w10091_ ;
	wire _w10090_ ;
	wire _w10089_ ;
	wire _w10088_ ;
	wire _w10087_ ;
	wire _w10086_ ;
	wire _w10085_ ;
	wire _w10084_ ;
	wire _w10083_ ;
	wire _w10082_ ;
	wire _w10081_ ;
	wire _w10080_ ;
	wire _w10079_ ;
	wire _w10078_ ;
	wire _w10077_ ;
	wire _w10076_ ;
	wire _w10075_ ;
	wire _w10074_ ;
	wire _w10073_ ;
	wire _w10072_ ;
	wire _w10071_ ;
	wire _w10070_ ;
	wire _w10069_ ;
	wire _w10068_ ;
	wire _w10067_ ;
	wire _w10066_ ;
	wire _w10065_ ;
	wire _w10064_ ;
	wire _w10063_ ;
	wire _w10062_ ;
	wire _w10061_ ;
	wire _w10060_ ;
	wire _w10059_ ;
	wire _w10058_ ;
	wire _w10057_ ;
	wire _w10056_ ;
	wire _w10055_ ;
	wire _w10054_ ;
	wire _w10053_ ;
	wire _w10052_ ;
	wire _w10051_ ;
	wire _w10050_ ;
	wire _w10049_ ;
	wire _w10048_ ;
	wire _w10047_ ;
	wire _w10046_ ;
	wire _w10045_ ;
	wire _w10044_ ;
	wire _w10043_ ;
	wire _w10042_ ;
	wire _w10041_ ;
	wire _w10040_ ;
	wire _w10039_ ;
	wire _w10038_ ;
	wire _w10037_ ;
	wire _w10036_ ;
	wire _w10035_ ;
	wire _w10034_ ;
	wire _w10033_ ;
	wire _w10032_ ;
	wire _w10031_ ;
	wire _w10030_ ;
	wire _w10029_ ;
	wire _w10028_ ;
	wire _w10027_ ;
	wire _w10026_ ;
	wire _w10025_ ;
	wire _w10024_ ;
	wire _w10023_ ;
	wire _w10022_ ;
	wire _w10021_ ;
	wire _w10020_ ;
	wire _w10019_ ;
	wire _w10018_ ;
	wire _w10017_ ;
	wire _w10016_ ;
	wire _w10015_ ;
	wire _w10014_ ;
	wire _w10013_ ;
	wire _w10012_ ;
	wire _w10011_ ;
	wire _w10010_ ;
	wire _w10009_ ;
	wire _w10008_ ;
	wire _w10007_ ;
	wire _w10006_ ;
	wire _w10005_ ;
	wire _w10004_ ;
	wire _w10003_ ;
	wire _w10002_ ;
	wire _w10001_ ;
	wire _w10000_ ;
	wire _w9999_ ;
	wire _w9998_ ;
	wire _w9997_ ;
	wire _w9996_ ;
	wire _w9995_ ;
	wire _w9994_ ;
	wire _w9993_ ;
	wire _w9992_ ;
	wire _w9991_ ;
	wire _w9990_ ;
	wire _w9989_ ;
	wire _w9988_ ;
	wire _w9987_ ;
	wire _w9986_ ;
	wire _w9985_ ;
	wire _w9984_ ;
	wire _w9983_ ;
	wire _w9982_ ;
	wire _w9981_ ;
	wire _w9980_ ;
	wire _w9979_ ;
	wire _w9978_ ;
	wire _w9977_ ;
	wire _w9976_ ;
	wire _w9975_ ;
	wire _w9974_ ;
	wire _w9973_ ;
	wire _w9972_ ;
	wire _w9971_ ;
	wire _w9970_ ;
	wire _w9969_ ;
	wire _w9968_ ;
	wire _w9967_ ;
	wire _w9966_ ;
	wire _w9965_ ;
	wire _w9964_ ;
	wire _w9963_ ;
	wire _w9962_ ;
	wire _w9961_ ;
	wire _w9960_ ;
	wire _w9959_ ;
	wire _w9958_ ;
	wire _w9957_ ;
	wire _w9956_ ;
	wire _w9955_ ;
	wire _w9954_ ;
	wire _w9953_ ;
	wire _w9952_ ;
	wire _w9951_ ;
	wire _w9950_ ;
	wire _w9949_ ;
	wire _w9948_ ;
	wire _w9947_ ;
	wire _w9946_ ;
	wire _w9945_ ;
	wire _w9944_ ;
	wire _w9943_ ;
	wire _w9942_ ;
	wire _w9941_ ;
	wire _w9940_ ;
	wire _w9939_ ;
	wire _w9938_ ;
	wire _w9937_ ;
	wire _w9936_ ;
	wire _w9935_ ;
	wire _w9934_ ;
	wire _w9933_ ;
	wire _w9932_ ;
	wire _w9931_ ;
	wire _w9930_ ;
	wire _w9929_ ;
	wire _w9928_ ;
	wire _w9927_ ;
	wire _w9926_ ;
	wire _w9925_ ;
	wire _w9924_ ;
	wire _w9923_ ;
	wire _w9922_ ;
	wire _w9921_ ;
	wire _w9920_ ;
	wire _w9919_ ;
	wire _w9918_ ;
	wire _w9917_ ;
	wire _w9916_ ;
	wire _w9915_ ;
	wire _w9914_ ;
	wire _w9913_ ;
	wire _w9912_ ;
	wire _w9911_ ;
	wire _w9910_ ;
	wire _w9909_ ;
	wire _w9908_ ;
	wire _w9907_ ;
	wire _w9906_ ;
	wire _w9905_ ;
	wire _w9904_ ;
	wire _w9903_ ;
	wire _w9902_ ;
	wire _w9901_ ;
	wire _w9900_ ;
	wire _w9899_ ;
	wire _w9898_ ;
	wire _w9897_ ;
	wire _w9896_ ;
	wire _w9895_ ;
	wire _w9894_ ;
	wire _w9893_ ;
	wire _w9892_ ;
	wire _w9891_ ;
	wire _w9890_ ;
	wire _w9889_ ;
	wire _w9888_ ;
	wire _w9887_ ;
	wire _w9886_ ;
	wire _w9885_ ;
	wire _w9884_ ;
	wire _w9883_ ;
	wire _w9882_ ;
	wire _w9881_ ;
	wire _w9880_ ;
	wire _w9879_ ;
	wire _w9878_ ;
	wire _w9877_ ;
	wire _w9876_ ;
	wire _w9875_ ;
	wire _w9874_ ;
	wire _w9873_ ;
	wire _w9872_ ;
	wire _w9871_ ;
	wire _w9870_ ;
	wire _w9869_ ;
	wire _w9868_ ;
	wire _w9867_ ;
	wire _w9866_ ;
	wire _w9865_ ;
	wire _w9864_ ;
	wire _w9863_ ;
	wire _w9862_ ;
	wire _w9861_ ;
	wire _w9860_ ;
	wire _w9859_ ;
	wire _w9858_ ;
	wire _w9857_ ;
	wire _w9856_ ;
	wire _w9855_ ;
	wire _w9854_ ;
	wire _w9853_ ;
	wire _w9852_ ;
	wire _w9851_ ;
	wire _w9850_ ;
	wire _w9849_ ;
	wire _w9848_ ;
	wire _w9847_ ;
	wire _w9846_ ;
	wire _w9845_ ;
	wire _w9844_ ;
	wire _w9843_ ;
	wire _w9842_ ;
	wire _w9841_ ;
	wire _w9840_ ;
	wire _w9839_ ;
	wire _w9838_ ;
	wire _w9837_ ;
	wire _w9836_ ;
	wire _w9835_ ;
	wire _w9834_ ;
	wire _w9833_ ;
	wire _w9832_ ;
	wire _w9831_ ;
	wire _w9830_ ;
	wire _w9829_ ;
	wire _w9828_ ;
	wire _w9827_ ;
	wire _w9826_ ;
	wire _w9825_ ;
	wire _w9824_ ;
	wire _w9823_ ;
	wire _w9822_ ;
	wire _w9821_ ;
	wire _w9820_ ;
	wire _w9819_ ;
	wire _w9818_ ;
	wire _w9817_ ;
	wire _w9816_ ;
	wire _w9815_ ;
	wire _w9814_ ;
	wire _w9813_ ;
	wire _w9812_ ;
	wire _w9811_ ;
	wire _w9810_ ;
	wire _w9809_ ;
	wire _w9808_ ;
	wire _w9807_ ;
	wire _w9806_ ;
	wire _w9805_ ;
	wire _w9804_ ;
	wire _w9803_ ;
	wire _w9802_ ;
	wire _w9801_ ;
	wire _w9800_ ;
	wire _w9799_ ;
	wire _w9798_ ;
	wire _w9797_ ;
	wire _w9796_ ;
	wire _w9795_ ;
	wire _w9794_ ;
	wire _w9793_ ;
	wire _w9792_ ;
	wire _w9791_ ;
	wire _w9790_ ;
	wire _w9789_ ;
	wire _w9788_ ;
	wire _w9787_ ;
	wire _w9786_ ;
	wire _w9785_ ;
	wire _w9784_ ;
	wire _w9783_ ;
	wire _w9782_ ;
	wire _w9781_ ;
	wire _w9780_ ;
	wire _w9779_ ;
	wire _w9778_ ;
	wire _w9777_ ;
	wire _w9776_ ;
	wire _w9775_ ;
	wire _w9774_ ;
	wire _w9773_ ;
	wire _w9772_ ;
	wire _w9771_ ;
	wire _w9770_ ;
	wire _w9769_ ;
	wire _w9768_ ;
	wire _w9767_ ;
	wire _w9766_ ;
	wire _w9765_ ;
	wire _w9764_ ;
	wire _w9763_ ;
	wire _w9762_ ;
	wire _w9761_ ;
	wire _w9760_ ;
	wire _w9759_ ;
	wire _w9758_ ;
	wire _w9757_ ;
	wire _w9756_ ;
	wire _w9755_ ;
	wire _w9754_ ;
	wire _w9753_ ;
	wire _w9752_ ;
	wire _w9751_ ;
	wire _w9750_ ;
	wire _w9749_ ;
	wire _w9748_ ;
	wire _w9747_ ;
	wire _w9746_ ;
	wire _w9745_ ;
	wire _w9744_ ;
	wire _w9743_ ;
	wire _w9742_ ;
	wire _w9741_ ;
	wire _w9740_ ;
	wire _w9739_ ;
	wire _w9738_ ;
	wire _w9737_ ;
	wire _w9736_ ;
	wire _w9735_ ;
	wire _w9734_ ;
	wire _w9733_ ;
	wire _w9732_ ;
	wire _w9731_ ;
	wire _w9730_ ;
	wire _w9729_ ;
	wire _w9728_ ;
	wire _w9727_ ;
	wire _w9726_ ;
	wire _w9725_ ;
	wire _w9724_ ;
	wire _w9723_ ;
	wire _w9722_ ;
	wire _w9721_ ;
	wire _w9720_ ;
	wire _w9719_ ;
	wire _w9718_ ;
	wire _w9717_ ;
	wire _w9716_ ;
	wire _w9715_ ;
	wire _w9714_ ;
	wire _w9713_ ;
	wire _w9712_ ;
	wire _w9711_ ;
	wire _w9710_ ;
	wire _w9709_ ;
	wire _w9708_ ;
	wire _w9707_ ;
	wire _w9706_ ;
	wire _w9705_ ;
	wire _w9704_ ;
	wire _w9703_ ;
	wire _w9702_ ;
	wire _w9701_ ;
	wire _w9700_ ;
	wire _w9699_ ;
	wire _w9698_ ;
	wire _w9697_ ;
	wire _w9696_ ;
	wire _w9695_ ;
	wire _w9694_ ;
	wire _w9693_ ;
	wire _w9692_ ;
	wire _w9691_ ;
	wire _w9690_ ;
	wire _w9689_ ;
	wire _w9688_ ;
	wire _w9687_ ;
	wire _w9686_ ;
	wire _w9685_ ;
	wire _w9684_ ;
	wire _w9683_ ;
	wire _w9682_ ;
	wire _w9681_ ;
	wire _w9680_ ;
	wire _w9679_ ;
	wire _w9678_ ;
	wire _w9677_ ;
	wire _w9676_ ;
	wire _w9675_ ;
	wire _w9674_ ;
	wire _w9673_ ;
	wire _w9672_ ;
	wire _w9671_ ;
	wire _w9670_ ;
	wire _w9669_ ;
	wire _w9668_ ;
	wire _w9667_ ;
	wire _w9666_ ;
	wire _w9665_ ;
	wire _w9664_ ;
	wire _w9663_ ;
	wire _w9662_ ;
	wire _w9661_ ;
	wire _w9660_ ;
	wire _w9659_ ;
	wire _w9658_ ;
	wire _w9657_ ;
	wire _w9656_ ;
	wire _w9655_ ;
	wire _w9654_ ;
	wire _w9653_ ;
	wire _w9652_ ;
	wire _w9651_ ;
	wire _w9650_ ;
	wire _w9649_ ;
	wire _w9648_ ;
	wire _w9647_ ;
	wire _w9646_ ;
	wire _w9645_ ;
	wire _w9644_ ;
	wire _w9643_ ;
	wire _w9642_ ;
	wire _w9641_ ;
	wire _w9640_ ;
	wire _w9639_ ;
	wire _w9638_ ;
	wire _w9637_ ;
	wire _w9636_ ;
	wire _w9635_ ;
	wire _w9634_ ;
	wire _w9633_ ;
	wire _w9632_ ;
	wire _w9631_ ;
	wire _w9630_ ;
	wire _w9629_ ;
	wire _w9628_ ;
	wire _w9627_ ;
	wire _w9626_ ;
	wire _w9625_ ;
	wire _w9624_ ;
	wire _w9623_ ;
	wire _w9622_ ;
	wire _w9621_ ;
	wire _w9620_ ;
	wire _w9619_ ;
	wire _w9618_ ;
	wire _w9617_ ;
	wire _w9616_ ;
	wire _w9615_ ;
	wire _w9614_ ;
	wire _w9613_ ;
	wire _w9612_ ;
	wire _w9611_ ;
	wire _w9610_ ;
	wire _w9609_ ;
	wire _w9608_ ;
	wire _w9607_ ;
	wire _w9606_ ;
	wire _w9605_ ;
	wire _w9604_ ;
	wire _w9603_ ;
	wire _w9602_ ;
	wire _w9601_ ;
	wire _w9600_ ;
	wire _w9599_ ;
	wire _w9598_ ;
	wire _w9597_ ;
	wire _w9596_ ;
	wire _w9595_ ;
	wire _w9594_ ;
	wire _w9593_ ;
	wire _w9592_ ;
	wire _w9591_ ;
	wire _w9590_ ;
	wire _w9589_ ;
	wire _w9588_ ;
	wire _w9587_ ;
	wire _w9586_ ;
	wire _w9585_ ;
	wire _w9584_ ;
	wire _w9583_ ;
	wire _w9582_ ;
	wire _w9581_ ;
	wire _w9580_ ;
	wire _w9579_ ;
	wire _w9578_ ;
	wire _w9577_ ;
	wire _w9576_ ;
	wire _w9575_ ;
	wire _w9574_ ;
	wire _w9573_ ;
	wire _w9572_ ;
	wire _w9571_ ;
	wire _w9570_ ;
	wire _w9569_ ;
	wire _w9568_ ;
	wire _w9567_ ;
	wire _w9566_ ;
	wire _w9565_ ;
	wire _w9564_ ;
	wire _w9563_ ;
	wire _w9562_ ;
	wire _w9561_ ;
	wire _w9560_ ;
	wire _w9559_ ;
	wire _w9558_ ;
	wire _w9557_ ;
	wire _w9556_ ;
	wire _w9555_ ;
	wire _w9554_ ;
	wire _w9553_ ;
	wire _w9552_ ;
	wire _w9551_ ;
	wire _w9550_ ;
	wire _w9549_ ;
	wire _w9548_ ;
	wire _w9547_ ;
	wire _w9546_ ;
	wire _w9545_ ;
	wire _w9544_ ;
	wire _w9543_ ;
	wire _w9542_ ;
	wire _w9541_ ;
	wire _w9540_ ;
	wire _w9539_ ;
	wire _w9538_ ;
	wire _w9537_ ;
	wire _w9536_ ;
	wire _w9535_ ;
	wire _w9534_ ;
	wire _w9533_ ;
	wire _w9532_ ;
	wire _w9531_ ;
	wire _w9530_ ;
	wire _w9529_ ;
	wire _w9528_ ;
	wire _w9527_ ;
	wire _w9526_ ;
	wire _w9525_ ;
	wire _w9524_ ;
	wire _w9523_ ;
	wire _w9522_ ;
	wire _w9521_ ;
	wire _w9520_ ;
	wire _w9519_ ;
	wire _w9518_ ;
	wire _w9517_ ;
	wire _w9516_ ;
	wire _w9515_ ;
	wire _w9514_ ;
	wire _w9513_ ;
	wire _w9512_ ;
	wire _w9511_ ;
	wire _w9510_ ;
	wire _w9509_ ;
	wire _w9508_ ;
	wire _w9507_ ;
	wire _w9506_ ;
	wire _w9505_ ;
	wire _w9504_ ;
	wire _w9503_ ;
	wire _w9502_ ;
	wire _w9501_ ;
	wire _w9500_ ;
	wire _w9499_ ;
	wire _w9498_ ;
	wire _w9497_ ;
	wire _w9496_ ;
	wire _w9495_ ;
	wire _w9494_ ;
	wire _w9493_ ;
	wire _w9492_ ;
	wire _w9491_ ;
	wire _w9490_ ;
	wire _w9489_ ;
	wire _w9488_ ;
	wire _w9487_ ;
	wire _w9486_ ;
	wire _w9485_ ;
	wire _w9484_ ;
	wire _w9483_ ;
	wire _w9482_ ;
	wire _w9481_ ;
	wire _w9480_ ;
	wire _w9479_ ;
	wire _w9478_ ;
	wire _w9477_ ;
	wire _w9476_ ;
	wire _w9475_ ;
	wire _w9474_ ;
	wire _w9473_ ;
	wire _w9472_ ;
	wire _w9471_ ;
	wire _w9470_ ;
	wire _w9469_ ;
	wire _w9468_ ;
	wire _w9467_ ;
	wire _w9466_ ;
	wire _w9465_ ;
	wire _w9464_ ;
	wire _w9463_ ;
	wire _w9462_ ;
	wire _w9461_ ;
	wire _w9460_ ;
	wire _w9459_ ;
	wire _w9458_ ;
	wire _w9457_ ;
	wire _w9456_ ;
	wire _w9455_ ;
	wire _w9454_ ;
	wire _w9453_ ;
	wire _w9452_ ;
	wire _w9451_ ;
	wire _w9450_ ;
	wire _w9449_ ;
	wire _w9448_ ;
	wire _w9447_ ;
	wire _w9446_ ;
	wire _w9445_ ;
	wire _w9444_ ;
	wire _w9443_ ;
	wire _w9442_ ;
	wire _w9441_ ;
	wire _w9440_ ;
	wire _w9439_ ;
	wire _w9438_ ;
	wire _w9437_ ;
	wire _w9436_ ;
	wire _w9435_ ;
	wire _w9434_ ;
	wire _w9433_ ;
	wire _w9432_ ;
	wire _w9431_ ;
	wire _w9430_ ;
	wire _w9429_ ;
	wire _w9428_ ;
	wire _w9427_ ;
	wire _w9426_ ;
	wire _w9425_ ;
	wire _w9424_ ;
	wire _w9423_ ;
	wire _w9422_ ;
	wire _w9421_ ;
	wire _w9420_ ;
	wire _w9419_ ;
	wire _w9418_ ;
	wire _w9417_ ;
	wire _w9416_ ;
	wire _w9415_ ;
	wire _w9414_ ;
	wire _w9413_ ;
	wire _w9412_ ;
	wire _w9411_ ;
	wire _w9410_ ;
	wire _w9409_ ;
	wire _w9408_ ;
	wire _w9407_ ;
	wire _w9406_ ;
	wire _w9405_ ;
	wire _w9404_ ;
	wire _w9403_ ;
	wire _w9402_ ;
	wire _w9401_ ;
	wire _w9400_ ;
	wire _w9399_ ;
	wire _w9398_ ;
	wire _w9397_ ;
	wire _w9396_ ;
	wire _w9395_ ;
	wire _w9394_ ;
	wire _w9393_ ;
	wire _w9392_ ;
	wire _w9391_ ;
	wire _w9390_ ;
	wire _w9389_ ;
	wire _w9388_ ;
	wire _w9387_ ;
	wire _w9386_ ;
	wire _w9385_ ;
	wire _w9384_ ;
	wire _w9383_ ;
	wire _w9382_ ;
	wire _w9381_ ;
	wire _w9380_ ;
	wire _w9379_ ;
	wire _w9378_ ;
	wire _w9377_ ;
	wire _w9376_ ;
	wire _w9375_ ;
	wire _w9374_ ;
	wire _w9373_ ;
	wire _w9372_ ;
	wire _w9371_ ;
	wire _w9370_ ;
	wire _w9369_ ;
	wire _w9368_ ;
	wire _w9367_ ;
	wire _w9366_ ;
	wire _w9365_ ;
	wire _w9364_ ;
	wire _w9363_ ;
	wire _w9362_ ;
	wire _w9361_ ;
	wire _w9360_ ;
	wire _w9359_ ;
	wire _w9358_ ;
	wire _w9357_ ;
	wire _w9356_ ;
	wire _w9355_ ;
	wire _w9354_ ;
	wire _w9353_ ;
	wire _w9352_ ;
	wire _w9351_ ;
	wire _w9350_ ;
	wire _w9349_ ;
	wire _w9348_ ;
	wire _w9347_ ;
	wire _w9346_ ;
	wire _w9345_ ;
	wire _w9344_ ;
	wire _w9343_ ;
	wire _w9342_ ;
	wire _w9341_ ;
	wire _w9340_ ;
	wire _w9339_ ;
	wire _w9338_ ;
	wire _w9337_ ;
	wire _w9336_ ;
	wire _w9335_ ;
	wire _w9334_ ;
	wire _w9333_ ;
	wire _w9332_ ;
	wire _w9331_ ;
	wire _w9330_ ;
	wire _w9329_ ;
	wire _w9328_ ;
	wire _w9327_ ;
	wire _w9326_ ;
	wire _w9325_ ;
	wire _w9324_ ;
	wire _w9323_ ;
	wire _w9322_ ;
	wire _w9321_ ;
	wire _w9320_ ;
	wire _w9319_ ;
	wire _w9318_ ;
	wire _w9317_ ;
	wire _w9316_ ;
	wire _w9315_ ;
	wire _w9314_ ;
	wire _w9313_ ;
	wire _w9312_ ;
	wire _w9311_ ;
	wire _w9310_ ;
	wire _w9309_ ;
	wire _w9308_ ;
	wire _w9307_ ;
	wire _w9306_ ;
	wire _w9305_ ;
	wire _w9304_ ;
	wire _w9303_ ;
	wire _w9302_ ;
	wire _w9301_ ;
	wire _w9300_ ;
	wire _w9299_ ;
	wire _w9298_ ;
	wire _w9297_ ;
	wire _w9296_ ;
	wire _w9295_ ;
	wire _w9294_ ;
	wire _w9293_ ;
	wire _w9292_ ;
	wire _w9291_ ;
	wire _w9290_ ;
	wire _w9289_ ;
	wire _w9288_ ;
	wire _w9287_ ;
	wire _w9286_ ;
	wire _w9285_ ;
	wire _w9284_ ;
	wire _w9283_ ;
	wire _w9282_ ;
	wire _w9281_ ;
	wire _w9280_ ;
	wire _w9279_ ;
	wire _w9278_ ;
	wire _w9277_ ;
	wire _w9276_ ;
	wire _w9275_ ;
	wire _w9274_ ;
	wire _w9273_ ;
	wire _w9272_ ;
	wire _w9271_ ;
	wire _w9270_ ;
	wire _w9269_ ;
	wire _w9268_ ;
	wire _w9267_ ;
	wire _w9266_ ;
	wire _w9265_ ;
	wire _w9264_ ;
	wire _w9263_ ;
	wire _w9262_ ;
	wire _w9261_ ;
	wire _w9260_ ;
	wire _w9259_ ;
	wire _w9258_ ;
	wire _w9257_ ;
	wire _w9256_ ;
	wire _w9255_ ;
	wire _w9254_ ;
	wire _w9253_ ;
	wire _w9252_ ;
	wire _w9251_ ;
	wire _w9250_ ;
	wire _w9249_ ;
	wire _w9248_ ;
	wire _w9247_ ;
	wire _w9246_ ;
	wire _w9245_ ;
	wire _w9244_ ;
	wire _w9243_ ;
	wire _w9242_ ;
	wire _w9241_ ;
	wire _w9240_ ;
	wire _w9239_ ;
	wire _w9238_ ;
	wire _w9237_ ;
	wire _w9236_ ;
	wire _w9235_ ;
	wire _w9234_ ;
	wire _w9233_ ;
	wire _w9232_ ;
	wire _w9231_ ;
	wire _w9230_ ;
	wire _w9229_ ;
	wire _w9228_ ;
	wire _w9227_ ;
	wire _w9226_ ;
	wire _w9225_ ;
	wire _w9224_ ;
	wire _w9223_ ;
	wire _w9222_ ;
	wire _w9221_ ;
	wire _w9220_ ;
	wire _w9219_ ;
	wire _w9218_ ;
	wire _w9217_ ;
	wire _w9216_ ;
	wire _w9215_ ;
	wire _w9214_ ;
	wire _w9213_ ;
	wire _w9212_ ;
	wire _w9211_ ;
	wire _w9210_ ;
	wire _w9209_ ;
	wire _w9208_ ;
	wire _w9207_ ;
	wire _w9206_ ;
	wire _w9205_ ;
	wire _w9204_ ;
	wire _w9203_ ;
	wire _w9202_ ;
	wire _w9201_ ;
	wire _w9200_ ;
	wire _w9199_ ;
	wire _w9198_ ;
	wire _w9197_ ;
	wire _w9196_ ;
	wire _w9195_ ;
	wire _w9194_ ;
	wire _w9193_ ;
	wire _w9192_ ;
	wire _w9191_ ;
	wire _w9190_ ;
	wire _w9189_ ;
	wire _w9188_ ;
	wire _w9187_ ;
	wire _w9186_ ;
	wire _w9185_ ;
	wire _w9184_ ;
	wire _w9183_ ;
	wire _w9182_ ;
	wire _w9181_ ;
	wire _w9180_ ;
	wire _w9179_ ;
	wire _w9178_ ;
	wire _w9177_ ;
	wire _w9176_ ;
	wire _w9175_ ;
	wire _w9174_ ;
	wire _w9173_ ;
	wire _w9172_ ;
	wire _w9171_ ;
	wire _w9170_ ;
	wire _w9169_ ;
	wire _w9168_ ;
	wire _w9167_ ;
	wire _w9166_ ;
	wire _w9165_ ;
	wire _w9164_ ;
	wire _w9163_ ;
	wire _w9162_ ;
	wire _w9161_ ;
	wire _w9160_ ;
	wire _w9159_ ;
	wire _w9158_ ;
	wire _w9157_ ;
	wire _w9156_ ;
	wire _w9155_ ;
	wire _w9154_ ;
	wire _w9153_ ;
	wire _w9152_ ;
	wire _w9151_ ;
	wire _w9150_ ;
	wire _w9149_ ;
	wire _w9148_ ;
	wire _w9147_ ;
	wire _w9146_ ;
	wire _w9145_ ;
	wire _w9144_ ;
	wire _w9143_ ;
	wire _w9142_ ;
	wire _w9141_ ;
	wire _w9140_ ;
	wire _w9139_ ;
	wire _w9138_ ;
	wire _w9137_ ;
	wire _w9136_ ;
	wire _w9135_ ;
	wire _w9134_ ;
	wire _w6403_ ;
	wire _w6402_ ;
	wire _w6401_ ;
	wire _w6400_ ;
	wire _w6399_ ;
	wire _w6398_ ;
	wire _w6397_ ;
	wire _w6396_ ;
	wire _w6395_ ;
	wire _w6394_ ;
	wire _w6393_ ;
	wire _w6392_ ;
	wire _w6391_ ;
	wire _w6390_ ;
	wire _w6389_ ;
	wire _w6388_ ;
	wire _w6387_ ;
	wire _w6386_ ;
	wire _w6385_ ;
	wire _w6384_ ;
	wire _w6383_ ;
	wire _w6382_ ;
	wire _w6381_ ;
	wire _w6380_ ;
	wire _w6379_ ;
	wire _w6378_ ;
	wire _w6377_ ;
	wire _w6376_ ;
	wire _w6375_ ;
	wire _w6374_ ;
	wire _w6373_ ;
	wire _w6372_ ;
	wire _w6371_ ;
	wire _w6370_ ;
	wire _w6369_ ;
	wire _w6368_ ;
	wire _w6367_ ;
	wire _w6366_ ;
	wire _w6365_ ;
	wire _w6364_ ;
	wire _w6363_ ;
	wire _w6362_ ;
	wire _w6361_ ;
	wire _w6360_ ;
	wire _w6359_ ;
	wire _w6358_ ;
	wire _w6357_ ;
	wire _w6356_ ;
	wire _w6355_ ;
	wire _w6354_ ;
	wire _w6353_ ;
	wire _w6352_ ;
	wire _w6351_ ;
	wire _w6350_ ;
	wire _w6349_ ;
	wire _w6348_ ;
	wire _w6347_ ;
	wire _w6346_ ;
	wire _w6345_ ;
	wire _w6344_ ;
	wire _w6343_ ;
	wire _w6342_ ;
	wire _w6341_ ;
	wire _w6340_ ;
	wire _w6339_ ;
	wire _w6338_ ;
	wire _w6337_ ;
	wire _w6336_ ;
	wire _w6335_ ;
	wire _w6334_ ;
	wire _w6333_ ;
	wire _w6332_ ;
	wire _w6331_ ;
	wire _w6330_ ;
	wire _w6329_ ;
	wire _w6328_ ;
	wire _w6327_ ;
	wire _w6326_ ;
	wire _w6325_ ;
	wire _w6324_ ;
	wire _w6323_ ;
	wire _w6322_ ;
	wire _w6321_ ;
	wire _w6320_ ;
	wire _w6319_ ;
	wire _w6318_ ;
	wire _w6317_ ;
	wire _w6316_ ;
	wire _w6315_ ;
	wire _w6314_ ;
	wire _w6313_ ;
	wire _w6312_ ;
	wire _w6311_ ;
	wire _w6310_ ;
	wire _w6309_ ;
	wire _w6308_ ;
	wire _w6307_ ;
	wire _w6306_ ;
	wire _w6305_ ;
	wire _w6304_ ;
	wire _w6303_ ;
	wire _w6302_ ;
	wire _w6301_ ;
	wire _w6300_ ;
	wire _w6299_ ;
	wire _w6298_ ;
	wire _w6297_ ;
	wire _w6296_ ;
	wire _w6295_ ;
	wire _w6294_ ;
	wire _w6293_ ;
	wire _w6292_ ;
	wire _w6291_ ;
	wire _w6290_ ;
	wire _w6289_ ;
	wire _w6288_ ;
	wire _w6287_ ;
	wire _w6286_ ;
	wire _w6285_ ;
	wire _w6284_ ;
	wire _w6283_ ;
	wire _w6282_ ;
	wire _w6281_ ;
	wire _w6280_ ;
	wire _w6279_ ;
	wire _w6278_ ;
	wire _w6277_ ;
	wire _w6276_ ;
	wire _w6275_ ;
	wire _w6274_ ;
	wire _w6273_ ;
	wire _w6272_ ;
	wire _w6271_ ;
	wire _w6270_ ;
	wire _w6269_ ;
	wire _w6268_ ;
	wire _w6267_ ;
	wire _w6266_ ;
	wire _w6265_ ;
	wire _w6264_ ;
	wire _w6263_ ;
	wire _w6262_ ;
	wire _w6261_ ;
	wire _w6260_ ;
	wire _w6259_ ;
	wire _w6258_ ;
	wire _w6257_ ;
	wire _w6256_ ;
	wire _w6255_ ;
	wire _w6254_ ;
	wire _w6253_ ;
	wire _w6252_ ;
	wire _w6251_ ;
	wire _w6250_ ;
	wire _w6249_ ;
	wire _w6248_ ;
	wire _w6247_ ;
	wire _w6246_ ;
	wire _w6245_ ;
	wire _w6244_ ;
	wire _w6243_ ;
	wire _w6242_ ;
	wire _w6241_ ;
	wire _w6240_ ;
	wire _w6239_ ;
	wire _w6238_ ;
	wire _w6237_ ;
	wire _w6236_ ;
	wire _w6235_ ;
	wire _w6234_ ;
	wire _w6233_ ;
	wire _w6232_ ;
	wire _w6231_ ;
	wire _w6230_ ;
	wire _w6229_ ;
	wire _w6228_ ;
	wire _w6227_ ;
	wire _w6226_ ;
	wire _w6225_ ;
	wire _w6224_ ;
	wire _w6223_ ;
	wire _w6222_ ;
	wire _w6221_ ;
	wire _w6220_ ;
	wire _w6219_ ;
	wire _w6218_ ;
	wire _w6217_ ;
	wire _w6216_ ;
	wire _w6215_ ;
	wire _w6214_ ;
	wire _w6213_ ;
	wire _w6212_ ;
	wire _w6211_ ;
	wire _w6210_ ;
	wire _w6209_ ;
	wire _w6208_ ;
	wire _w6207_ ;
	wire _w6206_ ;
	wire _w6205_ ;
	wire _w6204_ ;
	wire _w6203_ ;
	wire _w6202_ ;
	wire _w6201_ ;
	wire _w6200_ ;
	wire _w6199_ ;
	wire _w6198_ ;
	wire _w6197_ ;
	wire _w6196_ ;
	wire _w6195_ ;
	wire _w6194_ ;
	wire _w6193_ ;
	wire _w6192_ ;
	wire _w6191_ ;
	wire _w6190_ ;
	wire _w6189_ ;
	wire _w6188_ ;
	wire _w6187_ ;
	wire _w6186_ ;
	wire _w6185_ ;
	wire _w6184_ ;
	wire _w6183_ ;
	wire _w6182_ ;
	wire _w6181_ ;
	wire _w6180_ ;
	wire _w6179_ ;
	wire _w6178_ ;
	wire _w6177_ ;
	wire _w6176_ ;
	wire _w6175_ ;
	wire _w6174_ ;
	wire _w6173_ ;
	wire _w6172_ ;
	wire _w6171_ ;
	wire _w6170_ ;
	wire _w6169_ ;
	wire _w6168_ ;
	wire _w6167_ ;
	wire _w6166_ ;
	wire _w6165_ ;
	wire _w6164_ ;
	wire _w6163_ ;
	wire _w6162_ ;
	wire _w6161_ ;
	wire _w6160_ ;
	wire _w6159_ ;
	wire _w6158_ ;
	wire _w6157_ ;
	wire _w6156_ ;
	wire _w6155_ ;
	wire _w6154_ ;
	wire _w6153_ ;
	wire _w6152_ ;
	wire _w6151_ ;
	wire _w6150_ ;
	wire _w6149_ ;
	wire _w6148_ ;
	wire _w6147_ ;
	wire _w6146_ ;
	wire _w6145_ ;
	wire _w6144_ ;
	wire _w6143_ ;
	wire _w6142_ ;
	wire _w6141_ ;
	wire _w6140_ ;
	wire _w6139_ ;
	wire _w6138_ ;
	wire _w6137_ ;
	wire _w6136_ ;
	wire _w6135_ ;
	wire _w6134_ ;
	wire _w6133_ ;
	wire _w6132_ ;
	wire _w6131_ ;
	wire _w6130_ ;
	wire _w6129_ ;
	wire _w6128_ ;
	wire _w6127_ ;
	wire _w6126_ ;
	wire _w6125_ ;
	wire _w6124_ ;
	wire _w6123_ ;
	wire _w6122_ ;
	wire _w6121_ ;
	wire _w6120_ ;
	wire _w6119_ ;
	wire _w6118_ ;
	wire _w6117_ ;
	wire _w6116_ ;
	wire _w6115_ ;
	wire _w6114_ ;
	wire _w6113_ ;
	wire _w6112_ ;
	wire _w6111_ ;
	wire _w6110_ ;
	wire _w6109_ ;
	wire _w6108_ ;
	wire _w6107_ ;
	wire _w6106_ ;
	wire _w6105_ ;
	wire _w6104_ ;
	wire _w6103_ ;
	wire _w6102_ ;
	wire _w6101_ ;
	wire _w6100_ ;
	wire _w6099_ ;
	wire _w6098_ ;
	wire _w6097_ ;
	wire _w6096_ ;
	wire _w6095_ ;
	wire _w6094_ ;
	wire _w6093_ ;
	wire _w6092_ ;
	wire _w6091_ ;
	wire _w6090_ ;
	wire _w6089_ ;
	wire _w6088_ ;
	wire _w6087_ ;
	wire _w6086_ ;
	wire _w6085_ ;
	wire _w6084_ ;
	wire _w6083_ ;
	wire _w6082_ ;
	wire _w6081_ ;
	wire _w6080_ ;
	wire _w6079_ ;
	wire _w6078_ ;
	wire _w6077_ ;
	wire _w6076_ ;
	wire _w6075_ ;
	wire _w6074_ ;
	wire _w6073_ ;
	wire _w6072_ ;
	wire _w6071_ ;
	wire _w6070_ ;
	wire _w6069_ ;
	wire _w6068_ ;
	wire _w6067_ ;
	wire _w6066_ ;
	wire _w6065_ ;
	wire _w6064_ ;
	wire _w6063_ ;
	wire _w6062_ ;
	wire _w6061_ ;
	wire _w6060_ ;
	wire _w6059_ ;
	wire _w6058_ ;
	wire _w6057_ ;
	wire _w6056_ ;
	wire _w6055_ ;
	wire _w6054_ ;
	wire _w6053_ ;
	wire _w6052_ ;
	wire _w6051_ ;
	wire _w6050_ ;
	wire _w6049_ ;
	wire _w6048_ ;
	wire _w6047_ ;
	wire _w6046_ ;
	wire _w6045_ ;
	wire _w6044_ ;
	wire _w6043_ ;
	wire _w6042_ ;
	wire _w6041_ ;
	wire _w6040_ ;
	wire _w6039_ ;
	wire _w6038_ ;
	wire _w6037_ ;
	wire _w6036_ ;
	wire _w6035_ ;
	wire _w6034_ ;
	wire _w6033_ ;
	wire _w6032_ ;
	wire _w6031_ ;
	wire _w6030_ ;
	wire _w6029_ ;
	wire _w6028_ ;
	wire _w6027_ ;
	wire _w6026_ ;
	wire _w6025_ ;
	wire _w6024_ ;
	wire _w6023_ ;
	wire _w6022_ ;
	wire _w6021_ ;
	wire _w6020_ ;
	wire _w6019_ ;
	wire _w6018_ ;
	wire _w6017_ ;
	wire _w6016_ ;
	wire _w6015_ ;
	wire _w6014_ ;
	wire _w6013_ ;
	wire _w6012_ ;
	wire _w6011_ ;
	wire _w6010_ ;
	wire _w6009_ ;
	wire _w6008_ ;
	wire _w6007_ ;
	wire _w6006_ ;
	wire _w6005_ ;
	wire _w6004_ ;
	wire _w6003_ ;
	wire _w6002_ ;
	wire _w6001_ ;
	wire _w6000_ ;
	wire _w5999_ ;
	wire _w5998_ ;
	wire _w5997_ ;
	wire _w5996_ ;
	wire _w5995_ ;
	wire _w5994_ ;
	wire _w5993_ ;
	wire _w5992_ ;
	wire _w5991_ ;
	wire _w5990_ ;
	wire _w5989_ ;
	wire _w5988_ ;
	wire _w5987_ ;
	wire _w5986_ ;
	wire _w5985_ ;
	wire _w5984_ ;
	wire _w5983_ ;
	wire _w5982_ ;
	wire _w5981_ ;
	wire _w5980_ ;
	wire _w5979_ ;
	wire _w5978_ ;
	wire _w5977_ ;
	wire _w5976_ ;
	wire _w5975_ ;
	wire _w5974_ ;
	wire _w5973_ ;
	wire _w5972_ ;
	wire _w5971_ ;
	wire _w5970_ ;
	wire _w5969_ ;
	wire _w5968_ ;
	wire _w5967_ ;
	wire _w5966_ ;
	wire _w5965_ ;
	wire _w5964_ ;
	wire _w5963_ ;
	wire _w5962_ ;
	wire _w5961_ ;
	wire _w5960_ ;
	wire _w5959_ ;
	wire _w5958_ ;
	wire _w5957_ ;
	wire _w5956_ ;
	wire _w5955_ ;
	wire _w5954_ ;
	wire _w5953_ ;
	wire _w5952_ ;
	wire _w5951_ ;
	wire _w5950_ ;
	wire _w5949_ ;
	wire _w5948_ ;
	wire _w5947_ ;
	wire _w5946_ ;
	wire _w5945_ ;
	wire _w5944_ ;
	wire _w5943_ ;
	wire _w5942_ ;
	wire _w5941_ ;
	wire _w5940_ ;
	wire _w5939_ ;
	wire _w5938_ ;
	wire _w5937_ ;
	wire _w5936_ ;
	wire _w5935_ ;
	wire _w5934_ ;
	wire _w5933_ ;
	wire _w5932_ ;
	wire _w5931_ ;
	wire _w5930_ ;
	wire _w5929_ ;
	wire _w5928_ ;
	wire _w5927_ ;
	wire _w5926_ ;
	wire _w5925_ ;
	wire _w5924_ ;
	wire _w5923_ ;
	wire _w5922_ ;
	wire _w5921_ ;
	wire _w5920_ ;
	wire _w5919_ ;
	wire _w5918_ ;
	wire _w5917_ ;
	wire _w5916_ ;
	wire _w5915_ ;
	wire _w5914_ ;
	wire _w5913_ ;
	wire _w5912_ ;
	wire _w5911_ ;
	wire _w5910_ ;
	wire _w5909_ ;
	wire _w5908_ ;
	wire _w5907_ ;
	wire _w5906_ ;
	wire _w5905_ ;
	wire _w5904_ ;
	wire _w5903_ ;
	wire _w5902_ ;
	wire _w5901_ ;
	wire _w5900_ ;
	wire _w5899_ ;
	wire _w5898_ ;
	wire _w5897_ ;
	wire _w5896_ ;
	wire _w5895_ ;
	wire _w5894_ ;
	wire _w5893_ ;
	wire _w5892_ ;
	wire _w5891_ ;
	wire _w5890_ ;
	wire _w5889_ ;
	wire _w5888_ ;
	wire _w5887_ ;
	wire _w5886_ ;
	wire _w5885_ ;
	wire _w5884_ ;
	wire _w5883_ ;
	wire _w5882_ ;
	wire _w5881_ ;
	wire _w5880_ ;
	wire _w5879_ ;
	wire _w5878_ ;
	wire _w5877_ ;
	wire _w5876_ ;
	wire _w5875_ ;
	wire _w5874_ ;
	wire _w5873_ ;
	wire _w5872_ ;
	wire _w5871_ ;
	wire _w5870_ ;
	wire _w5869_ ;
	wire _w5868_ ;
	wire _w5867_ ;
	wire _w5866_ ;
	wire _w5865_ ;
	wire _w5864_ ;
	wire _w5863_ ;
	wire _w5862_ ;
	wire _w5861_ ;
	wire _w5860_ ;
	wire _w5859_ ;
	wire _w5858_ ;
	wire _w5857_ ;
	wire _w5856_ ;
	wire _w5855_ ;
	wire _w5854_ ;
	wire _w5853_ ;
	wire _w5852_ ;
	wire _w5851_ ;
	wire _w5850_ ;
	wire _w5849_ ;
	wire _w5848_ ;
	wire _w5847_ ;
	wire _w5846_ ;
	wire _w5845_ ;
	wire _w5844_ ;
	wire _w5843_ ;
	wire _w5842_ ;
	wire _w5841_ ;
	wire _w5840_ ;
	wire _w5839_ ;
	wire _w5838_ ;
	wire _w5837_ ;
	wire _w5836_ ;
	wire _w5835_ ;
	wire _w5834_ ;
	wire _w5833_ ;
	wire _w5832_ ;
	wire _w5831_ ;
	wire _w5830_ ;
	wire _w5829_ ;
	wire _w5828_ ;
	wire _w5827_ ;
	wire _w5826_ ;
	wire _w5825_ ;
	wire _w5824_ ;
	wire _w5823_ ;
	wire _w5822_ ;
	wire _w5821_ ;
	wire _w5820_ ;
	wire _w5819_ ;
	wire _w5818_ ;
	wire _w5817_ ;
	wire _w5816_ ;
	wire _w5815_ ;
	wire _w5814_ ;
	wire _w5813_ ;
	wire _w5812_ ;
	wire _w5811_ ;
	wire _w5810_ ;
	wire _w5809_ ;
	wire _w5808_ ;
	wire _w5807_ ;
	wire _w5806_ ;
	wire _w5805_ ;
	wire _w5804_ ;
	wire _w5803_ ;
	wire _w5802_ ;
	wire _w5801_ ;
	wire _w5800_ ;
	wire _w5799_ ;
	wire _w5798_ ;
	wire _w5797_ ;
	wire _w5796_ ;
	wire _w5795_ ;
	wire _w5794_ ;
	wire _w5793_ ;
	wire _w5792_ ;
	wire _w5791_ ;
	wire _w5790_ ;
	wire _w5789_ ;
	wire _w5788_ ;
	wire _w5787_ ;
	wire _w5786_ ;
	wire _w5785_ ;
	wire _w5784_ ;
	wire _w5783_ ;
	wire _w5782_ ;
	wire _w5781_ ;
	wire _w5780_ ;
	wire _w5779_ ;
	wire _w5778_ ;
	wire _w5777_ ;
	wire _w5776_ ;
	wire _w5775_ ;
	wire _w5774_ ;
	wire _w5773_ ;
	wire _w5772_ ;
	wire _w5771_ ;
	wire _w5770_ ;
	wire _w5769_ ;
	wire _w5768_ ;
	wire _w5767_ ;
	wire _w5766_ ;
	wire _w5765_ ;
	wire _w5764_ ;
	wire _w5763_ ;
	wire _w5762_ ;
	wire _w5761_ ;
	wire _w5760_ ;
	wire _w5759_ ;
	wire _w5758_ ;
	wire _w5757_ ;
	wire _w5756_ ;
	wire _w5755_ ;
	wire _w5754_ ;
	wire _w5753_ ;
	wire _w5752_ ;
	wire _w5751_ ;
	wire _w5750_ ;
	wire _w5749_ ;
	wire _w5748_ ;
	wire _w5747_ ;
	wire _w5746_ ;
	wire _w5745_ ;
	wire _w5744_ ;
	wire _w5743_ ;
	wire _w5742_ ;
	wire _w5741_ ;
	wire _w5740_ ;
	wire _w5739_ ;
	wire _w5738_ ;
	wire _w5737_ ;
	wire _w5736_ ;
	wire _w5735_ ;
	wire _w5734_ ;
	wire _w5733_ ;
	wire _w5732_ ;
	wire _w5731_ ;
	wire _w5730_ ;
	wire _w5729_ ;
	wire _w5728_ ;
	wire _w5727_ ;
	wire _w5726_ ;
	wire _w5725_ ;
	wire _w5724_ ;
	wire _w5723_ ;
	wire _w5722_ ;
	wire _w5721_ ;
	wire _w5720_ ;
	wire _w5719_ ;
	wire _w5718_ ;
	wire _w5717_ ;
	wire _w5716_ ;
	wire _w5715_ ;
	wire _w5714_ ;
	wire _w5713_ ;
	wire _w5712_ ;
	wire _w5711_ ;
	wire _w5710_ ;
	wire _w5709_ ;
	wire _w5708_ ;
	wire _w5707_ ;
	wire _w5706_ ;
	wire _w5705_ ;
	wire _w5704_ ;
	wire _w5703_ ;
	wire _w5702_ ;
	wire _w5701_ ;
	wire _w5700_ ;
	wire _w5699_ ;
	wire _w5698_ ;
	wire _w5697_ ;
	wire _w5696_ ;
	wire _w5695_ ;
	wire _w5694_ ;
	wire _w5693_ ;
	wire _w5692_ ;
	wire _w5691_ ;
	wire _w5690_ ;
	wire _w5689_ ;
	wire _w5688_ ;
	wire _w5687_ ;
	wire _w5686_ ;
	wire _w5685_ ;
	wire _w5684_ ;
	wire _w5683_ ;
	wire _w5682_ ;
	wire _w5681_ ;
	wire _w5680_ ;
	wire _w5679_ ;
	wire _w5678_ ;
	wire _w5677_ ;
	wire _w5676_ ;
	wire _w5675_ ;
	wire _w5674_ ;
	wire _w5673_ ;
	wire _w5672_ ;
	wire _w5671_ ;
	wire _w5670_ ;
	wire _w5669_ ;
	wire _w5668_ ;
	wire _w5667_ ;
	wire _w5666_ ;
	wire _w5665_ ;
	wire _w5664_ ;
	wire _w5663_ ;
	wire _w5662_ ;
	wire _w5661_ ;
	wire _w5660_ ;
	wire _w5659_ ;
	wire _w5658_ ;
	wire _w5657_ ;
	wire _w5656_ ;
	wire _w5655_ ;
	wire _w5654_ ;
	wire _w5653_ ;
	wire _w5652_ ;
	wire _w5651_ ;
	wire _w5650_ ;
	wire _w5649_ ;
	wire _w5648_ ;
	wire _w5647_ ;
	wire _w5646_ ;
	wire _w5645_ ;
	wire _w5644_ ;
	wire _w5643_ ;
	wire _w5642_ ;
	wire _w5641_ ;
	wire _w5640_ ;
	wire _w5639_ ;
	wire _w5638_ ;
	wire _w5637_ ;
	wire _w5636_ ;
	wire _w5635_ ;
	wire _w5634_ ;
	wire _w5633_ ;
	wire _w5632_ ;
	wire _w5631_ ;
	wire _w5630_ ;
	wire _w5629_ ;
	wire _w5628_ ;
	wire _w5627_ ;
	wire _w5626_ ;
	wire _w5625_ ;
	wire _w5624_ ;
	wire _w5623_ ;
	wire _w5622_ ;
	wire _w5621_ ;
	wire _w5620_ ;
	wire _w5619_ ;
	wire _w5618_ ;
	wire _w5617_ ;
	wire _w5616_ ;
	wire _w5615_ ;
	wire _w5614_ ;
	wire _w5613_ ;
	wire _w5612_ ;
	wire _w5611_ ;
	wire _w5610_ ;
	wire _w5609_ ;
	wire _w5608_ ;
	wire _w5607_ ;
	wire _w5606_ ;
	wire _w5605_ ;
	wire _w5604_ ;
	wire _w5603_ ;
	wire _w5602_ ;
	wire _w5601_ ;
	wire _w5600_ ;
	wire _w5599_ ;
	wire _w5598_ ;
	wire _w5597_ ;
	wire _w5596_ ;
	wire _w5595_ ;
	wire _w5594_ ;
	wire _w5593_ ;
	wire _w5592_ ;
	wire _w5591_ ;
	wire _w5590_ ;
	wire _w5589_ ;
	wire _w5588_ ;
	wire _w5587_ ;
	wire _w5586_ ;
	wire _w5585_ ;
	wire _w5584_ ;
	wire _w5583_ ;
	wire _w5582_ ;
	wire _w5581_ ;
	wire _w5580_ ;
	wire _w5579_ ;
	wire _w5578_ ;
	wire _w5577_ ;
	wire _w5576_ ;
	wire _w5575_ ;
	wire _w5574_ ;
	wire _w5573_ ;
	wire _w5572_ ;
	wire _w5571_ ;
	wire _w5570_ ;
	wire _w5569_ ;
	wire _w5568_ ;
	wire _w5567_ ;
	wire _w5566_ ;
	wire _w5565_ ;
	wire _w5564_ ;
	wire _w5563_ ;
	wire _w5562_ ;
	wire _w5561_ ;
	wire _w5560_ ;
	wire _w5559_ ;
	wire _w5558_ ;
	wire _w5557_ ;
	wire _w5556_ ;
	wire _w5555_ ;
	wire _w5554_ ;
	wire _w5553_ ;
	wire _w5552_ ;
	wire _w5551_ ;
	wire _w5550_ ;
	wire _w5549_ ;
	wire _w5548_ ;
	wire _w5547_ ;
	wire _w5546_ ;
	wire _w5545_ ;
	wire _w5544_ ;
	wire _w5543_ ;
	wire _w5542_ ;
	wire _w5541_ ;
	wire _w5540_ ;
	wire _w5539_ ;
	wire _w5538_ ;
	wire _w5537_ ;
	wire _w5536_ ;
	wire _w5535_ ;
	wire _w5534_ ;
	wire _w5533_ ;
	wire _w5532_ ;
	wire _w5531_ ;
	wire _w5530_ ;
	wire _w5529_ ;
	wire _w5528_ ;
	wire _w5527_ ;
	wire _w5526_ ;
	wire _w5525_ ;
	wire _w5524_ ;
	wire _w5523_ ;
	wire _w5522_ ;
	wire _w5521_ ;
	wire _w5520_ ;
	wire _w5519_ ;
	wire _w5518_ ;
	wire _w5517_ ;
	wire _w5516_ ;
	wire _w5515_ ;
	wire _w5514_ ;
	wire _w5513_ ;
	wire _w5512_ ;
	wire _w5511_ ;
	wire _w5510_ ;
	wire _w5509_ ;
	wire _w5508_ ;
	wire _w5507_ ;
	wire _w5506_ ;
	wire _w5505_ ;
	wire _w5504_ ;
	wire _w5503_ ;
	wire _w5502_ ;
	wire _w5501_ ;
	wire _w5500_ ;
	wire _w5499_ ;
	wire _w5498_ ;
	wire _w5497_ ;
	wire _w5496_ ;
	wire _w5495_ ;
	wire _w5494_ ;
	wire _w5493_ ;
	wire _w5492_ ;
	wire _w5491_ ;
	wire _w5490_ ;
	wire _w5489_ ;
	wire _w5488_ ;
	wire _w5487_ ;
	wire _w5486_ ;
	wire _w5485_ ;
	wire _w5484_ ;
	wire _w5483_ ;
	wire _w5482_ ;
	wire _w5481_ ;
	wire _w5480_ ;
	wire _w5479_ ;
	wire _w5478_ ;
	wire _w5477_ ;
	wire _w5476_ ;
	wire _w5475_ ;
	wire _w5474_ ;
	wire _w5473_ ;
	wire _w5472_ ;
	wire _w5471_ ;
	wire _w5470_ ;
	wire _w5469_ ;
	wire _w5468_ ;
	wire _w5467_ ;
	wire _w5466_ ;
	wire _w5465_ ;
	wire _w5464_ ;
	wire _w5463_ ;
	wire _w5462_ ;
	wire _w5461_ ;
	wire _w5460_ ;
	wire _w5459_ ;
	wire _w5458_ ;
	wire _w5457_ ;
	wire _w5456_ ;
	wire _w5455_ ;
	wire _w5454_ ;
	wire _w5453_ ;
	wire _w5452_ ;
	wire _w5451_ ;
	wire _w5450_ ;
	wire _w5449_ ;
	wire _w5448_ ;
	wire _w5447_ ;
	wire _w5446_ ;
	wire _w5445_ ;
	wire _w5444_ ;
	wire _w5443_ ;
	wire _w5442_ ;
	wire _w5441_ ;
	wire _w5440_ ;
	wire _w5439_ ;
	wire _w5438_ ;
	wire _w5437_ ;
	wire _w5436_ ;
	wire _w5435_ ;
	wire _w5434_ ;
	wire _w5433_ ;
	wire _w5432_ ;
	wire _w5431_ ;
	wire _w5430_ ;
	wire _w5429_ ;
	wire _w5428_ ;
	wire _w5427_ ;
	wire _w5426_ ;
	wire _w5425_ ;
	wire _w5424_ ;
	wire _w5423_ ;
	wire _w5422_ ;
	wire _w5421_ ;
	wire _w5420_ ;
	wire _w5419_ ;
	wire _w5418_ ;
	wire _w5417_ ;
	wire _w5416_ ;
	wire _w5415_ ;
	wire _w5414_ ;
	wire _w5413_ ;
	wire _w5412_ ;
	wire _w5411_ ;
	wire _w5410_ ;
	wire _w5409_ ;
	wire _w5408_ ;
	wire _w5407_ ;
	wire _w5406_ ;
	wire _w5405_ ;
	wire _w5404_ ;
	wire _w5403_ ;
	wire _w5402_ ;
	wire _w5401_ ;
	wire _w5400_ ;
	wire _w5399_ ;
	wire _w5398_ ;
	wire _w5397_ ;
	wire _w5396_ ;
	wire _w5395_ ;
	wire _w5394_ ;
	wire _w5393_ ;
	wire _w5392_ ;
	wire _w5391_ ;
	wire _w5390_ ;
	wire _w5389_ ;
	wire _w5388_ ;
	wire _w5387_ ;
	wire _w5386_ ;
	wire _w5385_ ;
	wire _w5384_ ;
	wire _w5383_ ;
	wire _w5382_ ;
	wire _w5381_ ;
	wire _w5380_ ;
	wire _w5379_ ;
	wire _w5378_ ;
	wire _w5377_ ;
	wire _w5376_ ;
	wire _w5375_ ;
	wire _w5374_ ;
	wire _w5373_ ;
	wire _w5372_ ;
	wire _w5371_ ;
	wire _w5370_ ;
	wire _w5369_ ;
	wire _w5368_ ;
	wire _w5367_ ;
	wire _w5366_ ;
	wire _w5365_ ;
	wire _w5364_ ;
	wire _w5363_ ;
	wire _w5362_ ;
	wire _w5361_ ;
	wire _w5360_ ;
	wire _w5359_ ;
	wire _w5358_ ;
	wire _w5357_ ;
	wire _w5356_ ;
	wire _w5355_ ;
	wire _w5354_ ;
	wire _w5353_ ;
	wire _w5352_ ;
	wire _w5351_ ;
	wire _w5350_ ;
	wire _w5349_ ;
	wire _w5348_ ;
	wire _w5347_ ;
	wire _w5346_ ;
	wire _w5345_ ;
	wire _w5344_ ;
	wire _w5343_ ;
	wire _w5342_ ;
	wire _w5341_ ;
	wire _w5340_ ;
	wire _w5339_ ;
	wire _w5338_ ;
	wire _w5337_ ;
	wire _w5336_ ;
	wire _w5335_ ;
	wire _w5334_ ;
	wire _w5333_ ;
	wire _w5332_ ;
	wire _w5331_ ;
	wire _w5330_ ;
	wire _w5329_ ;
	wire _w5328_ ;
	wire _w5327_ ;
	wire _w5326_ ;
	wire _w5325_ ;
	wire _w5324_ ;
	wire _w5323_ ;
	wire _w5322_ ;
	wire _w5321_ ;
	wire _w5320_ ;
	wire _w5319_ ;
	wire _w5318_ ;
	wire _w5317_ ;
	wire _w5316_ ;
	wire _w5315_ ;
	wire _w5314_ ;
	wire _w5313_ ;
	wire _w5312_ ;
	wire _w5311_ ;
	wire _w5310_ ;
	wire _w5309_ ;
	wire _w5308_ ;
	wire _w5307_ ;
	wire _w5306_ ;
	wire _w5305_ ;
	wire _w5304_ ;
	wire _w5303_ ;
	wire _w5302_ ;
	wire _w5301_ ;
	wire _w5300_ ;
	wire _w5299_ ;
	wire _w5298_ ;
	wire _w5297_ ;
	wire _w5296_ ;
	wire _w5295_ ;
	wire _w5294_ ;
	wire _w5293_ ;
	wire _w5292_ ;
	wire _w5291_ ;
	wire _w5290_ ;
	wire _w5289_ ;
	wire _w5288_ ;
	wire _w5287_ ;
	wire _w5286_ ;
	wire _w5285_ ;
	wire _w5284_ ;
	wire _w5283_ ;
	wire _w5282_ ;
	wire _w5281_ ;
	wire _w5280_ ;
	wire _w5279_ ;
	wire _w5278_ ;
	wire _w5277_ ;
	wire _w5276_ ;
	wire _w5275_ ;
	wire _w5274_ ;
	wire _w5273_ ;
	wire _w5272_ ;
	wire _w5271_ ;
	wire _w5270_ ;
	wire _w5269_ ;
	wire _w5268_ ;
	wire _w5267_ ;
	wire _w5266_ ;
	wire _w5265_ ;
	wire _w5264_ ;
	wire _w5263_ ;
	wire _w5262_ ;
	wire _w5261_ ;
	wire _w5260_ ;
	wire _w5259_ ;
	wire _w5258_ ;
	wire _w5257_ ;
	wire _w5256_ ;
	wire _w5255_ ;
	wire _w5254_ ;
	wire _w5253_ ;
	wire _w5252_ ;
	wire _w5251_ ;
	wire _w5250_ ;
	wire _w5249_ ;
	wire _w5248_ ;
	wire _w5247_ ;
	wire _w5246_ ;
	wire _w5245_ ;
	wire _w5244_ ;
	wire _w5243_ ;
	wire _w5242_ ;
	wire _w5241_ ;
	wire _w5240_ ;
	wire _w5239_ ;
	wire _w5238_ ;
	wire _w5237_ ;
	wire _w5236_ ;
	wire _w5235_ ;
	wire _w5234_ ;
	wire _w5233_ ;
	wire _w5232_ ;
	wire _w5231_ ;
	wire _w5230_ ;
	wire _w5229_ ;
	wire _w5228_ ;
	wire _w5227_ ;
	wire _w5226_ ;
	wire _w5225_ ;
	wire _w5224_ ;
	wire _w5223_ ;
	wire _w5222_ ;
	wire _w5221_ ;
	wire _w5220_ ;
	wire _w5219_ ;
	wire _w5218_ ;
	wire _w5217_ ;
	wire _w5216_ ;
	wire _w5215_ ;
	wire _w5214_ ;
	wire _w5213_ ;
	wire _w5212_ ;
	wire _w5211_ ;
	wire _w5210_ ;
	wire _w5209_ ;
	wire _w5208_ ;
	wire _w5207_ ;
	wire _w5206_ ;
	wire _w5205_ ;
	wire _w5204_ ;
	wire _w5203_ ;
	wire _w5202_ ;
	wire _w5201_ ;
	wire _w5200_ ;
	wire _w5199_ ;
	wire _w5198_ ;
	wire _w5197_ ;
	wire _w5196_ ;
	wire _w5195_ ;
	wire _w5194_ ;
	wire _w5193_ ;
	wire _w5192_ ;
	wire _w5191_ ;
	wire _w5190_ ;
	wire _w5189_ ;
	wire _w5188_ ;
	wire _w5187_ ;
	wire _w5186_ ;
	wire _w5185_ ;
	wire _w5184_ ;
	wire _w5183_ ;
	wire _w5182_ ;
	wire _w5181_ ;
	wire _w5180_ ;
	wire _w5179_ ;
	wire _w5178_ ;
	wire _w5177_ ;
	wire _w5176_ ;
	wire _w5175_ ;
	wire _w5174_ ;
	wire _w5173_ ;
	wire _w5172_ ;
	wire _w5171_ ;
	wire _w5170_ ;
	wire _w5169_ ;
	wire _w5168_ ;
	wire _w5167_ ;
	wire _w5166_ ;
	wire _w5165_ ;
	wire _w5164_ ;
	wire _w5163_ ;
	wire _w5162_ ;
	wire _w5161_ ;
	wire _w5160_ ;
	wire _w5159_ ;
	wire _w5158_ ;
	wire _w5157_ ;
	wire _w5156_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	wire _w7233_ ;
	wire _w7234_ ;
	wire _w7235_ ;
	wire _w7236_ ;
	wire _w7237_ ;
	wire _w7238_ ;
	wire _w7239_ ;
	wire _w7240_ ;
	wire _w7241_ ;
	wire _w7242_ ;
	wire _w7243_ ;
	wire _w7244_ ;
	wire _w7245_ ;
	wire _w7246_ ;
	wire _w7247_ ;
	wire _w7248_ ;
	wire _w7249_ ;
	wire _w7250_ ;
	wire _w7251_ ;
	wire _w7252_ ;
	wire _w7253_ ;
	wire _w7254_ ;
	wire _w7255_ ;
	wire _w7256_ ;
	wire _w7257_ ;
	wire _w7258_ ;
	wire _w7259_ ;
	wire _w7260_ ;
	wire _w7261_ ;
	wire _w7262_ ;
	wire _w7263_ ;
	wire _w7264_ ;
	wire _w7265_ ;
	wire _w7266_ ;
	wire _w7267_ ;
	wire _w7268_ ;
	wire _w7269_ ;
	wire _w7270_ ;
	wire _w7271_ ;
	wire _w7272_ ;
	wire _w7273_ ;
	wire _w7274_ ;
	wire _w7275_ ;
	wire _w7276_ ;
	wire _w7277_ ;
	wire _w7278_ ;
	wire _w7279_ ;
	wire _w7280_ ;
	wire _w7281_ ;
	wire _w7282_ ;
	wire _w7283_ ;
	wire _w7284_ ;
	wire _w7285_ ;
	wire _w7286_ ;
	wire _w7287_ ;
	wire _w7288_ ;
	wire _w7289_ ;
	wire _w7290_ ;
	wire _w7291_ ;
	wire _w7292_ ;
	wire _w7293_ ;
	wire _w7294_ ;
	wire _w7295_ ;
	wire _w7296_ ;
	wire _w7297_ ;
	wire _w7298_ ;
	wire _w7299_ ;
	wire _w7300_ ;
	wire _w7301_ ;
	wire _w7302_ ;
	wire _w7303_ ;
	wire _w7304_ ;
	wire _w7305_ ;
	wire _w7306_ ;
	wire _w7307_ ;
	wire _w7308_ ;
	wire _w7309_ ;
	wire _w7310_ ;
	wire _w7311_ ;
	wire _w7312_ ;
	wire _w7313_ ;
	wire _w7314_ ;
	wire _w7315_ ;
	wire _w7316_ ;
	wire _w7317_ ;
	wire _w7318_ ;
	wire _w7319_ ;
	wire _w7320_ ;
	wire _w7321_ ;
	wire _w7322_ ;
	wire _w7323_ ;
	wire _w7324_ ;
	wire _w7325_ ;
	wire _w7326_ ;
	wire _w7327_ ;
	wire _w7328_ ;
	wire _w7329_ ;
	wire _w7330_ ;
	wire _w7331_ ;
	wire _w7332_ ;
	wire _w7333_ ;
	wire _w7334_ ;
	wire _w7335_ ;
	wire _w7336_ ;
	wire _w7337_ ;
	wire _w7338_ ;
	wire _w7339_ ;
	wire _w7340_ ;
	wire _w7341_ ;
	wire _w7342_ ;
	wire _w7343_ ;
	wire _w7344_ ;
	wire _w7345_ ;
	wire _w7346_ ;
	wire _w7347_ ;
	wire _w7348_ ;
	wire _w7349_ ;
	wire _w7350_ ;
	wire _w7351_ ;
	wire _w7352_ ;
	wire _w7353_ ;
	wire _w7354_ ;
	wire _w7355_ ;
	wire _w7356_ ;
	wire _w7357_ ;
	wire _w7358_ ;
	wire _w7359_ ;
	wire _w7360_ ;
	wire _w7361_ ;
	wire _w7362_ ;
	wire _w7363_ ;
	wire _w7364_ ;
	wire _w7365_ ;
	wire _w7366_ ;
	wire _w7367_ ;
	wire _w7368_ ;
	wire _w7369_ ;
	wire _w7370_ ;
	wire _w7371_ ;
	wire _w7372_ ;
	wire _w7373_ ;
	wire _w7374_ ;
	wire _w7375_ ;
	wire _w7376_ ;
	wire _w7377_ ;
	wire _w7378_ ;
	wire _w7379_ ;
	wire _w7380_ ;
	wire _w7381_ ;
	wire _w7382_ ;
	wire _w7383_ ;
	wire _w7384_ ;
	wire _w7385_ ;
	wire _w7386_ ;
	wire _w7387_ ;
	wire _w7388_ ;
	wire _w7389_ ;
	wire _w7390_ ;
	wire _w7391_ ;
	wire _w7392_ ;
	wire _w7393_ ;
	wire _w7394_ ;
	wire _w7395_ ;
	wire _w7396_ ;
	wire _w7397_ ;
	wire _w7398_ ;
	wire _w7399_ ;
	wire _w7400_ ;
	wire _w7401_ ;
	wire _w7402_ ;
	wire _w7403_ ;
	wire _w7404_ ;
	wire _w7405_ ;
	wire _w7406_ ;
	wire _w7407_ ;
	wire _w7408_ ;
	wire _w7409_ ;
	wire _w7410_ ;
	wire _w7411_ ;
	wire _w7412_ ;
	wire _w7413_ ;
	wire _w7414_ ;
	wire _w7415_ ;
	wire _w7416_ ;
	wire _w7417_ ;
	wire _w7418_ ;
	wire _w7419_ ;
	wire _w7420_ ;
	wire _w7421_ ;
	wire _w7422_ ;
	wire _w7423_ ;
	wire _w7424_ ;
	wire _w7425_ ;
	wire _w7426_ ;
	wire _w7427_ ;
	wire _w7428_ ;
	wire _w7429_ ;
	wire _w7430_ ;
	wire _w7431_ ;
	wire _w7432_ ;
	wire _w7433_ ;
	wire _w7434_ ;
	wire _w7435_ ;
	wire _w7436_ ;
	wire _w7437_ ;
	wire _w7438_ ;
	wire _w7439_ ;
	wire _w7440_ ;
	wire _w7441_ ;
	wire _w7442_ ;
	wire _w7443_ ;
	wire _w7444_ ;
	wire _w7445_ ;
	wire _w7446_ ;
	wire _w7447_ ;
	wire _w7448_ ;
	wire _w7449_ ;
	wire _w7450_ ;
	wire _w7451_ ;
	wire _w7452_ ;
	wire _w7453_ ;
	wire _w7454_ ;
	wire _w7455_ ;
	wire _w7456_ ;
	wire _w7457_ ;
	wire _w7458_ ;
	wire _w7459_ ;
	wire _w7460_ ;
	wire _w7461_ ;
	wire _w7462_ ;
	wire _w7463_ ;
	wire _w7464_ ;
	wire _w7465_ ;
	wire _w7466_ ;
	wire _w7467_ ;
	wire _w7468_ ;
	wire _w7469_ ;
	wire _w7470_ ;
	wire _w7471_ ;
	wire _w7472_ ;
	wire _w7473_ ;
	wire _w7474_ ;
	wire _w7475_ ;
	wire _w7476_ ;
	wire _w7477_ ;
	wire _w7478_ ;
	wire _w7479_ ;
	wire _w7480_ ;
	wire _w7481_ ;
	wire _w7482_ ;
	wire _w7483_ ;
	wire _w7484_ ;
	wire _w7485_ ;
	wire _w7486_ ;
	wire _w7487_ ;
	wire _w7488_ ;
	wire _w7489_ ;
	wire _w7490_ ;
	wire _w7491_ ;
	wire _w7492_ ;
	wire _w7493_ ;
	wire _w7494_ ;
	wire _w7495_ ;
	wire _w7496_ ;
	wire _w7497_ ;
	wire _w7498_ ;
	wire _w7499_ ;
	wire _w7500_ ;
	wire _w7501_ ;
	wire _w7502_ ;
	wire _w7503_ ;
	wire _w7504_ ;
	wire _w7505_ ;
	wire _w7506_ ;
	wire _w7507_ ;
	wire _w7508_ ;
	wire _w7509_ ;
	wire _w7510_ ;
	wire _w7511_ ;
	wire _w7512_ ;
	wire _w7513_ ;
	wire _w7514_ ;
	wire _w7515_ ;
	wire _w7516_ ;
	wire _w7517_ ;
	wire _w7518_ ;
	wire _w7519_ ;
	wire _w7520_ ;
	wire _w7521_ ;
	wire _w7522_ ;
	wire _w7523_ ;
	wire _w7524_ ;
	wire _w7525_ ;
	wire _w7526_ ;
	wire _w7527_ ;
	wire _w7528_ ;
	wire _w7529_ ;
	wire _w7530_ ;
	wire _w7531_ ;
	wire _w7532_ ;
	wire _w7533_ ;
	wire _w7534_ ;
	wire _w7535_ ;
	wire _w7536_ ;
	wire _w7537_ ;
	wire _w7538_ ;
	wire _w7539_ ;
	wire _w7540_ ;
	wire _w7541_ ;
	wire _w7542_ ;
	wire _w7543_ ;
	wire _w7544_ ;
	wire _w7545_ ;
	wire _w7546_ ;
	wire _w7547_ ;
	wire _w7548_ ;
	wire _w7549_ ;
	wire _w7550_ ;
	wire _w7551_ ;
	wire _w7552_ ;
	wire _w7553_ ;
	wire _w7554_ ;
	wire _w7555_ ;
	wire _w7556_ ;
	wire _w7557_ ;
	wire _w7558_ ;
	wire _w7559_ ;
	wire _w7560_ ;
	wire _w7561_ ;
	wire _w7562_ ;
	wire _w7563_ ;
	wire _w7564_ ;
	wire _w7565_ ;
	wire _w7566_ ;
	wire _w7567_ ;
	wire _w7568_ ;
	wire _w7569_ ;
	wire _w7570_ ;
	wire _w7571_ ;
	wire _w7572_ ;
	wire _w7573_ ;
	wire _w7574_ ;
	wire _w7575_ ;
	wire _w7576_ ;
	wire _w7577_ ;
	wire _w7578_ ;
	wire _w7579_ ;
	wire _w7580_ ;
	wire _w7581_ ;
	wire _w7582_ ;
	wire _w7583_ ;
	wire _w7584_ ;
	wire _w7585_ ;
	wire _w7586_ ;
	wire _w7587_ ;
	wire _w7588_ ;
	wire _w7589_ ;
	wire _w7590_ ;
	wire _w7591_ ;
	wire _w7592_ ;
	wire _w7593_ ;
	wire _w7594_ ;
	wire _w7595_ ;
	wire _w7596_ ;
	wire _w7597_ ;
	wire _w7598_ ;
	wire _w7599_ ;
	wire _w7600_ ;
	wire _w7601_ ;
	wire _w7602_ ;
	wire _w7603_ ;
	wire _w7604_ ;
	wire _w7605_ ;
	wire _w7606_ ;
	wire _w7607_ ;
	wire _w7608_ ;
	wire _w7609_ ;
	wire _w7610_ ;
	wire _w7611_ ;
	wire _w7612_ ;
	wire _w7613_ ;
	wire _w7614_ ;
	wire _w7615_ ;
	wire _w7616_ ;
	wire _w7617_ ;
	wire _w7618_ ;
	wire _w7619_ ;
	wire _w7620_ ;
	wire _w7621_ ;
	wire _w7622_ ;
	wire _w7623_ ;
	wire _w7624_ ;
	wire _w7625_ ;
	wire _w7626_ ;
	wire _w7627_ ;
	wire _w7628_ ;
	wire _w7629_ ;
	wire _w7630_ ;
	wire _w7631_ ;
	wire _w7632_ ;
	wire _w7633_ ;
	wire _w7634_ ;
	wire _w7635_ ;
	wire _w7636_ ;
	wire _w7637_ ;
	wire _w7638_ ;
	wire _w7639_ ;
	wire _w7640_ ;
	wire _w7641_ ;
	wire _w7642_ ;
	wire _w7643_ ;
	wire _w7644_ ;
	wire _w7645_ ;
	wire _w7646_ ;
	wire _w7647_ ;
	wire _w7648_ ;
	wire _w7649_ ;
	wire _w7650_ ;
	wire _w7651_ ;
	wire _w7652_ ;
	wire _w7653_ ;
	wire _w7654_ ;
	wire _w7655_ ;
	wire _w7656_ ;
	wire _w7657_ ;
	wire _w7658_ ;
	wire _w7659_ ;
	wire _w7660_ ;
	wire _w7661_ ;
	wire _w7662_ ;
	wire _w7663_ ;
	wire _w7664_ ;
	wire _w7665_ ;
	wire _w7666_ ;
	wire _w7667_ ;
	wire _w7668_ ;
	wire _w7669_ ;
	wire _w7670_ ;
	wire _w7671_ ;
	wire _w7672_ ;
	wire _w7673_ ;
	wire _w7674_ ;
	wire _w7675_ ;
	wire _w7676_ ;
	wire _w7677_ ;
	wire _w7678_ ;
	wire _w7679_ ;
	wire _w7680_ ;
	wire _w7681_ ;
	wire _w7682_ ;
	wire _w7683_ ;
	wire _w7684_ ;
	wire _w7685_ ;
	wire _w7686_ ;
	wire _w7687_ ;
	wire _w7688_ ;
	wire _w7689_ ;
	wire _w7690_ ;
	wire _w7691_ ;
	wire _w7692_ ;
	wire _w7693_ ;
	wire _w7694_ ;
	wire _w7695_ ;
	wire _w7696_ ;
	wire _w7697_ ;
	wire _w7698_ ;
	wire _w7699_ ;
	wire _w7700_ ;
	wire _w7701_ ;
	wire _w7702_ ;
	wire _w7703_ ;
	wire _w7704_ ;
	wire _w7705_ ;
	wire _w7706_ ;
	wire _w7707_ ;
	wire _w7708_ ;
	wire _w7709_ ;
	wire _w7710_ ;
	wire _w7711_ ;
	wire _w7712_ ;
	wire _w7713_ ;
	wire _w7714_ ;
	wire _w7715_ ;
	wire _w7716_ ;
	wire _w7717_ ;
	wire _w7718_ ;
	wire _w7719_ ;
	wire _w7720_ ;
	wire _w7721_ ;
	wire _w7722_ ;
	wire _w7723_ ;
	wire _w7724_ ;
	wire _w7725_ ;
	wire _w7726_ ;
	wire _w7727_ ;
	wire _w7728_ ;
	wire _w7729_ ;
	wire _w7730_ ;
	wire _w7731_ ;
	wire _w7732_ ;
	wire _w7733_ ;
	wire _w7734_ ;
	wire _w7735_ ;
	wire _w7736_ ;
	wire _w7737_ ;
	wire _w7738_ ;
	wire _w7739_ ;
	wire _w7740_ ;
	wire _w7741_ ;
	wire _w7742_ ;
	wire _w7743_ ;
	wire _w7744_ ;
	wire _w7745_ ;
	wire _w7746_ ;
	wire _w7747_ ;
	wire _w7748_ ;
	wire _w7749_ ;
	wire _w7750_ ;
	wire _w7751_ ;
	wire _w7752_ ;
	wire _w7753_ ;
	wire _w7754_ ;
	wire _w7755_ ;
	wire _w7756_ ;
	wire _w7757_ ;
	wire _w7758_ ;
	wire _w7759_ ;
	wire _w7760_ ;
	wire _w7761_ ;
	wire _w7762_ ;
	wire _w7763_ ;
	wire _w7764_ ;
	wire _w7765_ ;
	wire _w7766_ ;
	wire _w7767_ ;
	wire _w7768_ ;
	wire _w7769_ ;
	wire _w7770_ ;
	wire _w7771_ ;
	wire _w7772_ ;
	wire _w7773_ ;
	wire _w7774_ ;
	wire _w7775_ ;
	wire _w7776_ ;
	wire _w7777_ ;
	wire _w7778_ ;
	wire _w7779_ ;
	wire _w7780_ ;
	wire _w7781_ ;
	wire _w7782_ ;
	wire _w7783_ ;
	wire _w7784_ ;
	wire _w7785_ ;
	wire _w7786_ ;
	wire _w7787_ ;
	wire _w7788_ ;
	wire _w7789_ ;
	wire _w7790_ ;
	wire _w7791_ ;
	wire _w7792_ ;
	wire _w7793_ ;
	wire _w7794_ ;
	wire _w7795_ ;
	wire _w7796_ ;
	wire _w7797_ ;
	wire _w7798_ ;
	wire _w7799_ ;
	wire _w7800_ ;
	wire _w7801_ ;
	wire _w7802_ ;
	wire _w7803_ ;
	wire _w7804_ ;
	wire _w7805_ ;
	wire _w7806_ ;
	wire _w7807_ ;
	wire _w7808_ ;
	wire _w7809_ ;
	wire _w7810_ ;
	wire _w7811_ ;
	wire _w7812_ ;
	wire _w7813_ ;
	wire _w7814_ ;
	wire _w7815_ ;
	wire _w7816_ ;
	wire _w7817_ ;
	wire _w7818_ ;
	wire _w7819_ ;
	wire _w7820_ ;
	wire _w7821_ ;
	wire _w7822_ ;
	wire _w7823_ ;
	wire _w7824_ ;
	wire _w7825_ ;
	wire _w7826_ ;
	wire _w7827_ ;
	wire _w7828_ ;
	wire _w7829_ ;
	wire _w7830_ ;
	wire _w7831_ ;
	wire _w7832_ ;
	wire _w7833_ ;
	wire _w7834_ ;
	wire _w7835_ ;
	wire _w7836_ ;
	wire _w7837_ ;
	wire _w7838_ ;
	wire _w7839_ ;
	wire _w7840_ ;
	wire _w7841_ ;
	wire _w7842_ ;
	wire _w7843_ ;
	wire _w7844_ ;
	wire _w7845_ ;
	wire _w7846_ ;
	wire _w7847_ ;
	wire _w7848_ ;
	wire _w7849_ ;
	wire _w7850_ ;
	wire _w7851_ ;
	wire _w7852_ ;
	wire _w7853_ ;
	wire _w7854_ ;
	wire _w7855_ ;
	wire _w7856_ ;
	wire _w7857_ ;
	wire _w7858_ ;
	wire _w7859_ ;
	wire _w7860_ ;
	wire _w7861_ ;
	wire _w7862_ ;
	wire _w7863_ ;
	wire _w7864_ ;
	wire _w7865_ ;
	wire _w7866_ ;
	wire _w7867_ ;
	wire _w7868_ ;
	wire _w7869_ ;
	wire _w7870_ ;
	wire _w7871_ ;
	wire _w7872_ ;
	wire _w7873_ ;
	wire _w7874_ ;
	wire _w7875_ ;
	wire _w7876_ ;
	wire _w7877_ ;
	wire _w7878_ ;
	wire _w7879_ ;
	wire _w7880_ ;
	wire _w7881_ ;
	wire _w7882_ ;
	wire _w7883_ ;
	wire _w7884_ ;
	wire _w7885_ ;
	wire _w7886_ ;
	wire _w7887_ ;
	wire _w7888_ ;
	wire _w7889_ ;
	wire _w7890_ ;
	wire _w7891_ ;
	wire _w7892_ ;
	wire _w7893_ ;
	wire _w7894_ ;
	wire _w7895_ ;
	wire _w7896_ ;
	wire _w7897_ ;
	wire _w7898_ ;
	wire _w7899_ ;
	wire _w7900_ ;
	wire _w7901_ ;
	wire _w7902_ ;
	wire _w7903_ ;
	wire _w7904_ ;
	wire _w7905_ ;
	wire _w7906_ ;
	wire _w7907_ ;
	wire _w7908_ ;
	wire _w7909_ ;
	wire _w7910_ ;
	wire _w7911_ ;
	wire _w7912_ ;
	wire _w7913_ ;
	wire _w7914_ ;
	wire _w7915_ ;
	wire _w7916_ ;
	wire _w7917_ ;
	wire _w7918_ ;
	wire _w7919_ ;
	wire _w7920_ ;
	wire _w7921_ ;
	wire _w7922_ ;
	wire _w7923_ ;
	wire _w7924_ ;
	wire _w7925_ ;
	wire _w7926_ ;
	wire _w7927_ ;
	wire _w7928_ ;
	wire _w7929_ ;
	wire _w7930_ ;
	wire _w7931_ ;
	wire _w7932_ ;
	wire _w7933_ ;
	wire _w7934_ ;
	wire _w7935_ ;
	wire _w7936_ ;
	wire _w7937_ ;
	wire _w7938_ ;
	wire _w7939_ ;
	wire _w7940_ ;
	wire _w7941_ ;
	wire _w7942_ ;
	wire _w7943_ ;
	wire _w7944_ ;
	wire _w7945_ ;
	wire _w7946_ ;
	wire _w7947_ ;
	wire _w7948_ ;
	wire _w7949_ ;
	wire _w7950_ ;
	wire _w7951_ ;
	wire _w7952_ ;
	wire _w7953_ ;
	wire _w7954_ ;
	wire _w7955_ ;
	wire _w7956_ ;
	wire _w7957_ ;
	wire _w7958_ ;
	wire _w7959_ ;
	wire _w7960_ ;
	wire _w7961_ ;
	wire _w7962_ ;
	wire _w7963_ ;
	wire _w7964_ ;
	wire _w7965_ ;
	wire _w7966_ ;
	wire _w7967_ ;
	wire _w7968_ ;
	wire _w7969_ ;
	wire _w7970_ ;
	wire _w7971_ ;
	wire _w7972_ ;
	wire _w7973_ ;
	wire _w7974_ ;
	wire _w7975_ ;
	wire _w7976_ ;
	wire _w7977_ ;
	wire _w7978_ ;
	wire _w7979_ ;
	wire _w7980_ ;
	wire _w7981_ ;
	wire _w7982_ ;
	wire _w7983_ ;
	wire _w7984_ ;
	wire _w7985_ ;
	wire _w7986_ ;
	wire _w7987_ ;
	wire _w7988_ ;
	wire _w7989_ ;
	wire _w7990_ ;
	wire _w7991_ ;
	wire _w7992_ ;
	wire _w7993_ ;
	wire _w7994_ ;
	wire _w7995_ ;
	wire _w7996_ ;
	wire _w7997_ ;
	wire _w7998_ ;
	wire _w7999_ ;
	wire _w8000_ ;
	wire _w8001_ ;
	wire _w8002_ ;
	wire _w8003_ ;
	wire _w8004_ ;
	wire _w8005_ ;
	wire _w8006_ ;
	wire _w8007_ ;
	wire _w8008_ ;
	wire _w8009_ ;
	wire _w8010_ ;
	wire _w8011_ ;
	wire _w8012_ ;
	wire _w8013_ ;
	wire _w8014_ ;
	wire _w8015_ ;
	wire _w8016_ ;
	wire _w8017_ ;
	wire _w8018_ ;
	wire _w8019_ ;
	wire _w8020_ ;
	wire _w8021_ ;
	wire _w8022_ ;
	wire _w8023_ ;
	wire _w8024_ ;
	wire _w8025_ ;
	wire _w8026_ ;
	wire _w8027_ ;
	wire _w8028_ ;
	wire _w8029_ ;
	wire _w8030_ ;
	wire _w8031_ ;
	wire _w8032_ ;
	wire _w8033_ ;
	wire _w8034_ ;
	wire _w8035_ ;
	wire _w8036_ ;
	wire _w8037_ ;
	wire _w8038_ ;
	wire _w8039_ ;
	wire _w8040_ ;
	wire _w8041_ ;
	wire _w8042_ ;
	wire _w8043_ ;
	wire _w8044_ ;
	wire _w8045_ ;
	wire _w8046_ ;
	wire _w8047_ ;
	wire _w8048_ ;
	wire _w8049_ ;
	wire _w8050_ ;
	wire _w8051_ ;
	wire _w8052_ ;
	wire _w8053_ ;
	wire _w8054_ ;
	wire _w8055_ ;
	wire _w8056_ ;
	wire _w8057_ ;
	wire _w8058_ ;
	wire _w8059_ ;
	wire _w8060_ ;
	wire _w8061_ ;
	wire _w8062_ ;
	wire _w8063_ ;
	wire _w8064_ ;
	wire _w8065_ ;
	wire _w8066_ ;
	wire _w8067_ ;
	wire _w8068_ ;
	wire _w8069_ ;
	wire _w8070_ ;
	wire _w8071_ ;
	wire _w8072_ ;
	wire _w8073_ ;
	wire _w8074_ ;
	wire _w8075_ ;
	wire _w8076_ ;
	wire _w8077_ ;
	wire _w8078_ ;
	wire _w8079_ ;
	wire _w8080_ ;
	wire _w8081_ ;
	wire _w8082_ ;
	wire _w8083_ ;
	wire _w8084_ ;
	wire _w8085_ ;
	wire _w8086_ ;
	wire _w8087_ ;
	wire _w8088_ ;
	wire _w8089_ ;
	wire _w8090_ ;
	wire _w8091_ ;
	wire _w8092_ ;
	wire _w8093_ ;
	wire _w8094_ ;
	wire _w8095_ ;
	wire _w8096_ ;
	wire _w8097_ ;
	wire _w8098_ ;
	wire _w8099_ ;
	wire _w8100_ ;
	wire _w8101_ ;
	wire _w8102_ ;
	wire _w8103_ ;
	wire _w8104_ ;
	wire _w8105_ ;
	wire _w8106_ ;
	wire _w8107_ ;
	wire _w8108_ ;
	wire _w8109_ ;
	wire _w8110_ ;
	wire _w8111_ ;
	wire _w8112_ ;
	wire _w8113_ ;
	wire _w8114_ ;
	wire _w8115_ ;
	wire _w8116_ ;
	wire _w8117_ ;
	wire _w8118_ ;
	wire _w8119_ ;
	wire _w8120_ ;
	wire _w8121_ ;
	wire _w8122_ ;
	wire _w8123_ ;
	wire _w8124_ ;
	wire _w8125_ ;
	wire _w8126_ ;
	wire _w8127_ ;
	wire _w8128_ ;
	wire _w8129_ ;
	wire _w8130_ ;
	wire _w8131_ ;
	wire _w8132_ ;
	wire _w8133_ ;
	wire _w8134_ ;
	wire _w8135_ ;
	wire _w8136_ ;
	wire _w8137_ ;
	wire _w8138_ ;
	wire _w8139_ ;
	wire _w8140_ ;
	wire _w8141_ ;
	wire _w8142_ ;
	wire _w8143_ ;
	wire _w8144_ ;
	wire _w8145_ ;
	wire _w8146_ ;
	wire _w8147_ ;
	wire _w8148_ ;
	wire _w8149_ ;
	wire _w8150_ ;
	wire _w8151_ ;
	wire _w8152_ ;
	wire _w8153_ ;
	wire _w8154_ ;
	wire _w8155_ ;
	wire _w8156_ ;
	wire _w8157_ ;
	wire _w8158_ ;
	wire _w8159_ ;
	wire _w8160_ ;
	wire _w8161_ ;
	wire _w8162_ ;
	wire _w8163_ ;
	wire _w8164_ ;
	wire _w8165_ ;
	wire _w8166_ ;
	wire _w8167_ ;
	wire _w8168_ ;
	wire _w8169_ ;
	wire _w8170_ ;
	wire _w8171_ ;
	wire _w8172_ ;
	wire _w8173_ ;
	wire _w8174_ ;
	wire _w8175_ ;
	wire _w8176_ ;
	wire _w8177_ ;
	wire _w8178_ ;
	wire _w8179_ ;
	wire _w8180_ ;
	wire _w8181_ ;
	wire _w8182_ ;
	wire _w8183_ ;
	wire _w8184_ ;
	wire _w8185_ ;
	wire _w8186_ ;
	wire _w8187_ ;
	wire _w8188_ ;
	wire _w8189_ ;
	wire _w8190_ ;
	wire _w8191_ ;
	wire _w8192_ ;
	wire _w8193_ ;
	wire _w8194_ ;
	wire _w8195_ ;
	wire _w8196_ ;
	wire _w8197_ ;
	wire _w8198_ ;
	wire _w8199_ ;
	wire _w8200_ ;
	wire _w8201_ ;
	wire _w8202_ ;
	wire _w8203_ ;
	wire _w8204_ ;
	wire _w8205_ ;
	wire _w8206_ ;
	wire _w8207_ ;
	wire _w8208_ ;
	wire _w8209_ ;
	wire _w8210_ ;
	wire _w8211_ ;
	wire _w8212_ ;
	wire _w8213_ ;
	wire _w8214_ ;
	wire _w8215_ ;
	wire _w8216_ ;
	wire _w8217_ ;
	wire _w8218_ ;
	wire _w8219_ ;
	wire _w8220_ ;
	wire _w8221_ ;
	wire _w8222_ ;
	wire _w8223_ ;
	wire _w8224_ ;
	wire _w8225_ ;
	wire _w8226_ ;
	wire _w8227_ ;
	wire _w8228_ ;
	wire _w8229_ ;
	wire _w8230_ ;
	wire _w8231_ ;
	wire _w8232_ ;
	wire _w8233_ ;
	wire _w8234_ ;
	wire _w8235_ ;
	wire _w8236_ ;
	wire _w8237_ ;
	wire _w8238_ ;
	wire _w8239_ ;
	wire _w8240_ ;
	wire _w8241_ ;
	wire _w8242_ ;
	wire _w8243_ ;
	wire _w8244_ ;
	wire _w8245_ ;
	wire _w8246_ ;
	wire _w8247_ ;
	wire _w8248_ ;
	wire _w8249_ ;
	wire _w8250_ ;
	wire _w8251_ ;
	wire _w8252_ ;
	wire _w8253_ ;
	wire _w8254_ ;
	wire _w8255_ ;
	wire _w8256_ ;
	wire _w8257_ ;
	wire _w8258_ ;
	wire _w8259_ ;
	wire _w8260_ ;
	wire _w8261_ ;
	wire _w8262_ ;
	wire _w8263_ ;
	wire _w8264_ ;
	wire _w8265_ ;
	wire _w8266_ ;
	wire _w8267_ ;
	wire _w8268_ ;
	wire _w8269_ ;
	wire _w8270_ ;
	wire _w8271_ ;
	wire _w8272_ ;
	wire _w8273_ ;
	wire _w8274_ ;
	wire _w8275_ ;
	wire _w8276_ ;
	wire _w8277_ ;
	wire _w8278_ ;
	wire _w8279_ ;
	wire _w8280_ ;
	wire _w8281_ ;
	wire _w8282_ ;
	wire _w8283_ ;
	wire _w8284_ ;
	wire _w8285_ ;
	wire _w8286_ ;
	wire _w8287_ ;
	wire _w8288_ ;
	wire _w8289_ ;
	wire _w8290_ ;
	wire _w8291_ ;
	wire _w8292_ ;
	wire _w8293_ ;
	wire _w8294_ ;
	wire _w8295_ ;
	wire _w8296_ ;
	wire _w8297_ ;
	wire _w8298_ ;
	wire _w8299_ ;
	wire _w8300_ ;
	wire _w8301_ ;
	wire _w8302_ ;
	wire _w8303_ ;
	wire _w8304_ ;
	wire _w8305_ ;
	wire _w8306_ ;
	wire _w8307_ ;
	wire _w8308_ ;
	wire _w8309_ ;
	wire _w8310_ ;
	wire _w8311_ ;
	wire _w8312_ ;
	wire _w8313_ ;
	wire _w8314_ ;
	wire _w8315_ ;
	wire _w8316_ ;
	wire _w8317_ ;
	wire _w8318_ ;
	wire _w8319_ ;
	wire _w8320_ ;
	wire _w8321_ ;
	wire _w8322_ ;
	wire _w8323_ ;
	wire _w8324_ ;
	wire _w8325_ ;
	wire _w8326_ ;
	wire _w8327_ ;
	wire _w8328_ ;
	wire _w8329_ ;
	wire _w8330_ ;
	wire _w8331_ ;
	wire _w8332_ ;
	wire _w8333_ ;
	wire _w8334_ ;
	wire _w8335_ ;
	wire _w8336_ ;
	wire _w8337_ ;
	wire _w8338_ ;
	wire _w8339_ ;
	wire _w8340_ ;
	wire _w8341_ ;
	wire _w8342_ ;
	wire _w8343_ ;
	wire _w8344_ ;
	wire _w8345_ ;
	wire _w8346_ ;
	wire _w8347_ ;
	wire _w8348_ ;
	wire _w8349_ ;
	wire _w8350_ ;
	wire _w8351_ ;
	wire _w8352_ ;
	wire _w8353_ ;
	wire _w8354_ ;
	wire _w8355_ ;
	wire _w8356_ ;
	wire _w8357_ ;
	wire _w8358_ ;
	wire _w8359_ ;
	wire _w8360_ ;
	wire _w8361_ ;
	wire _w8362_ ;
	wire _w8363_ ;
	wire _w8364_ ;
	wire _w8365_ ;
	wire _w8366_ ;
	wire _w8367_ ;
	wire _w8368_ ;
	wire _w8369_ ;
	wire _w8370_ ;
	wire _w8371_ ;
	wire _w8372_ ;
	wire _w8373_ ;
	wire _w8374_ ;
	wire _w8375_ ;
	wire _w8376_ ;
	wire _w8377_ ;
	wire _w8378_ ;
	wire _w8379_ ;
	wire _w8380_ ;
	wire _w8381_ ;
	wire _w8382_ ;
	wire _w8383_ ;
	wire _w8384_ ;
	wire _w8385_ ;
	wire _w8386_ ;
	wire _w8387_ ;
	wire _w8388_ ;
	wire _w8389_ ;
	wire _w8390_ ;
	wire _w8391_ ;
	wire _w8392_ ;
	wire _w8393_ ;
	wire _w8394_ ;
	wire _w8395_ ;
	wire _w8396_ ;
	wire _w8397_ ;
	wire _w8398_ ;
	wire _w8399_ ;
	wire _w8400_ ;
	wire _w8401_ ;
	wire _w8402_ ;
	wire _w8403_ ;
	wire _w8404_ ;
	wire _w8405_ ;
	wire _w8406_ ;
	wire _w8407_ ;
	wire _w8408_ ;
	wire _w8409_ ;
	wire _w8410_ ;
	wire _w8411_ ;
	wire _w8412_ ;
	wire _w8413_ ;
	wire _w8414_ ;
	wire _w8415_ ;
	wire _w8416_ ;
	wire _w8417_ ;
	wire _w8418_ ;
	wire _w8419_ ;
	wire _w8420_ ;
	wire _w8421_ ;
	wire _w8422_ ;
	wire _w8423_ ;
	wire _w8424_ ;
	wire _w8425_ ;
	wire _w8426_ ;
	wire _w8427_ ;
	wire _w8428_ ;
	wire _w8429_ ;
	wire _w8430_ ;
	wire _w8431_ ;
	wire _w8432_ ;
	wire _w8433_ ;
	wire _w8434_ ;
	wire _w8435_ ;
	wire _w8436_ ;
	wire _w8437_ ;
	wire _w8438_ ;
	wire _w8439_ ;
	wire _w8440_ ;
	wire _w8441_ ;
	wire _w8442_ ;
	wire _w8443_ ;
	wire _w8444_ ;
	wire _w8445_ ;
	wire _w8446_ ;
	wire _w8447_ ;
	wire _w8448_ ;
	wire _w8449_ ;
	wire _w8450_ ;
	wire _w8451_ ;
	wire _w8452_ ;
	wire _w8453_ ;
	wire _w8454_ ;
	wire _w8455_ ;
	wire _w8456_ ;
	wire _w8457_ ;
	wire _w8458_ ;
	wire _w8459_ ;
	wire _w8460_ ;
	wire _w8461_ ;
	wire _w8462_ ;
	wire _w8463_ ;
	wire _w8464_ ;
	wire _w8465_ ;
	wire _w8466_ ;
	wire _w8467_ ;
	wire _w8468_ ;
	wire _w8469_ ;
	wire _w8470_ ;
	wire _w8471_ ;
	wire _w8472_ ;
	wire _w8473_ ;
	wire _w8474_ ;
	wire _w8475_ ;
	wire _w8476_ ;
	wire _w8477_ ;
	wire _w8478_ ;
	wire _w8479_ ;
	wire _w8480_ ;
	wire _w8481_ ;
	wire _w8482_ ;
	wire _w8483_ ;
	wire _w8484_ ;
	wire _w8485_ ;
	wire _w8486_ ;
	wire _w8487_ ;
	wire _w8488_ ;
	wire _w8489_ ;
	wire _w8490_ ;
	wire _w8491_ ;
	wire _w8492_ ;
	wire _w8493_ ;
	wire _w8494_ ;
	wire _w8495_ ;
	wire _w8496_ ;
	wire _w8497_ ;
	wire _w8498_ ;
	wire _w8499_ ;
	wire _w8500_ ;
	wire _w8501_ ;
	wire _w8502_ ;
	wire _w8503_ ;
	wire _w8504_ ;
	wire _w8505_ ;
	wire _w8506_ ;
	wire _w8507_ ;
	wire _w8508_ ;
	wire _w8509_ ;
	wire _w8510_ ;
	wire _w8511_ ;
	wire _w8512_ ;
	wire _w8513_ ;
	wire _w8514_ ;
	wire _w8515_ ;
	wire _w8516_ ;
	wire _w8517_ ;
	wire _w8518_ ;
	wire _w8519_ ;
	wire _w8520_ ;
	wire _w8521_ ;
	wire _w8522_ ;
	wire _w8523_ ;
	wire _w8524_ ;
	wire _w8525_ ;
	wire _w8526_ ;
	wire _w8527_ ;
	wire _w8528_ ;
	wire _w8529_ ;
	wire _w8530_ ;
	wire _w8531_ ;
	wire _w8532_ ;
	wire _w8533_ ;
	wire _w8534_ ;
	wire _w8535_ ;
	wire _w8536_ ;
	wire _w8537_ ;
	wire _w8538_ ;
	wire _w8539_ ;
	wire _w8540_ ;
	wire _w8541_ ;
	wire _w8542_ ;
	wire _w8543_ ;
	wire _w8544_ ;
	wire _w8545_ ;
	wire _w8546_ ;
	wire _w8547_ ;
	wire _w8548_ ;
	wire _w8549_ ;
	wire _w8550_ ;
	wire _w8551_ ;
	wire _w8552_ ;
	wire _w8553_ ;
	wire _w8554_ ;
	wire _w8555_ ;
	wire _w8556_ ;
	wire _w8557_ ;
	wire _w8558_ ;
	wire _w8559_ ;
	wire _w8560_ ;
	wire _w8561_ ;
	wire _w8562_ ;
	wire _w8563_ ;
	wire _w8564_ ;
	wire _w8565_ ;
	wire _w8566_ ;
	wire _w8567_ ;
	wire _w8568_ ;
	wire _w8569_ ;
	wire _w8570_ ;
	wire _w8571_ ;
	wire _w8572_ ;
	wire _w8573_ ;
	wire _w8574_ ;
	wire _w8575_ ;
	wire _w8576_ ;
	wire _w8577_ ;
	wire _w8578_ ;
	wire _w8579_ ;
	wire _w8580_ ;
	wire _w8581_ ;
	wire _w8582_ ;
	wire _w8583_ ;
	wire _w8584_ ;
	wire _w8585_ ;
	wire _w8586_ ;
	wire _w8587_ ;
	wire _w8588_ ;
	wire _w8589_ ;
	wire _w8590_ ;
	wire _w8591_ ;
	wire _w8592_ ;
	wire _w8593_ ;
	wire _w8594_ ;
	wire _w8595_ ;
	wire _w8596_ ;
	wire _w8597_ ;
	wire _w8598_ ;
	wire _w8599_ ;
	wire _w8600_ ;
	wire _w8601_ ;
	wire _w8602_ ;
	wire _w8603_ ;
	wire _w8604_ ;
	wire _w8605_ ;
	wire _w8606_ ;
	wire _w8607_ ;
	wire _w8608_ ;
	wire _w8609_ ;
	wire _w8610_ ;
	wire _w8611_ ;
	wire _w8612_ ;
	wire _w8613_ ;
	wire _w8614_ ;
	wire _w8615_ ;
	wire _w8616_ ;
	wire _w8617_ ;
	wire _w8618_ ;
	wire _w8619_ ;
	wire _w8620_ ;
	wire _w8621_ ;
	wire _w8622_ ;
	wire _w8623_ ;
	wire _w8624_ ;
	wire _w8625_ ;
	wire _w8626_ ;
	wire _w8627_ ;
	wire _w8628_ ;
	wire _w8629_ ;
	wire _w8630_ ;
	wire _w8631_ ;
	wire _w8632_ ;
	wire _w8633_ ;
	wire _w8634_ ;
	wire _w8635_ ;
	wire _w8636_ ;
	wire _w8637_ ;
	wire _w8638_ ;
	wire _w8639_ ;
	wire _w8640_ ;
	wire _w8641_ ;
	wire _w8642_ ;
	wire _w8643_ ;
	wire _w8644_ ;
	wire _w8645_ ;
	wire _w8646_ ;
	wire _w8647_ ;
	wire _w8648_ ;
	wire _w8649_ ;
	wire _w8650_ ;
	wire _w8651_ ;
	wire _w8652_ ;
	wire _w8653_ ;
	wire _w8654_ ;
	wire _w8655_ ;
	wire _w8656_ ;
	wire _w8657_ ;
	wire _w8658_ ;
	wire _w8659_ ;
	wire _w8660_ ;
	wire _w8661_ ;
	wire _w8662_ ;
	wire _w8663_ ;
	wire _w8664_ ;
	wire _w8665_ ;
	wire _w8666_ ;
	wire _w8667_ ;
	wire _w8668_ ;
	wire _w8669_ ;
	wire _w8670_ ;
	wire _w8671_ ;
	wire _w8672_ ;
	wire _w8673_ ;
	wire _w8674_ ;
	wire _w8675_ ;
	wire _w8676_ ;
	wire _w8677_ ;
	wire _w8678_ ;
	wire _w8679_ ;
	wire _w8680_ ;
	wire _w8681_ ;
	wire _w8682_ ;
	wire _w8683_ ;
	wire _w8684_ ;
	wire _w8685_ ;
	wire _w8686_ ;
	wire _w8687_ ;
	wire _w8688_ ;
	wire _w8689_ ;
	wire _w8690_ ;
	wire _w8691_ ;
	wire _w8692_ ;
	wire _w8693_ ;
	wire _w8694_ ;
	wire _w8695_ ;
	wire _w8696_ ;
	wire _w8697_ ;
	wire _w8698_ ;
	wire _w8699_ ;
	wire _w8700_ ;
	wire _w8701_ ;
	wire _w8702_ ;
	wire _w8703_ ;
	wire _w8704_ ;
	wire _w8705_ ;
	wire _w8706_ ;
	wire _w8707_ ;
	wire _w8708_ ;
	wire _w8709_ ;
	wire _w8710_ ;
	wire _w8711_ ;
	wire _w8712_ ;
	wire _w8713_ ;
	wire _w8714_ ;
	wire _w8715_ ;
	wire _w8716_ ;
	wire _w8717_ ;
	wire _w8718_ ;
	wire _w8719_ ;
	wire _w8720_ ;
	wire _w8721_ ;
	wire _w8722_ ;
	wire _w8723_ ;
	wire _w8724_ ;
	wire _w8725_ ;
	wire _w8726_ ;
	wire _w8727_ ;
	wire _w8728_ ;
	wire _w8729_ ;
	wire _w8730_ ;
	wire _w8731_ ;
	wire _w8732_ ;
	wire _w8733_ ;
	wire _w8734_ ;
	wire _w8735_ ;
	wire _w8736_ ;
	wire _w8737_ ;
	wire _w8738_ ;
	wire _w8739_ ;
	wire _w8740_ ;
	wire _w8741_ ;
	wire _w8742_ ;
	wire _w8743_ ;
	wire _w8744_ ;
	wire _w8745_ ;
	wire _w8746_ ;
	wire _w8747_ ;
	wire _w8748_ ;
	wire _w8749_ ;
	wire _w8750_ ;
	wire _w8751_ ;
	wire _w8752_ ;
	wire _w8753_ ;
	wire _w8754_ ;
	wire _w8755_ ;
	wire _w8756_ ;
	wire _w8757_ ;
	wire _w8758_ ;
	wire _w8759_ ;
	wire _w8760_ ;
	wire _w8761_ ;
	wire _w8762_ ;
	wire _w8763_ ;
	wire _w8764_ ;
	wire _w8765_ ;
	wire _w8766_ ;
	wire _w8767_ ;
	wire _w8768_ ;
	wire _w8769_ ;
	wire _w8770_ ;
	wire _w8771_ ;
	wire _w8772_ ;
	wire _w8773_ ;
	wire _w8774_ ;
	wire _w8775_ ;
	wire _w8776_ ;
	wire _w8777_ ;
	wire _w8778_ ;
	wire _w8779_ ;
	wire _w8780_ ;
	wire _w8781_ ;
	wire _w8782_ ;
	wire _w8783_ ;
	wire _w8784_ ;
	wire _w8785_ ;
	wire _w8786_ ;
	wire _w8787_ ;
	wire _w8788_ ;
	wire _w8789_ ;
	wire _w8790_ ;
	wire _w8791_ ;
	wire _w8792_ ;
	wire _w8793_ ;
	wire _w8794_ ;
	wire _w8795_ ;
	wire _w8796_ ;
	wire _w8797_ ;
	wire _w8798_ ;
	wire _w8799_ ;
	wire _w8800_ ;
	wire _w8801_ ;
	wire _w8802_ ;
	wire _w8803_ ;
	wire _w8804_ ;
	wire _w8805_ ;
	wire _w8806_ ;
	wire _w8807_ ;
	wire _w8808_ ;
	wire _w8809_ ;
	wire _w8810_ ;
	wire _w8811_ ;
	wire _w8812_ ;
	wire _w8813_ ;
	wire _w8814_ ;
	wire _w8815_ ;
	wire _w8816_ ;
	wire _w8817_ ;
	wire _w8818_ ;
	wire _w8819_ ;
	wire _w8820_ ;
	wire _w8821_ ;
	wire _w8822_ ;
	wire _w8823_ ;
	wire _w8824_ ;
	wire _w8825_ ;
	wire _w8826_ ;
	wire _w8827_ ;
	wire _w8828_ ;
	wire _w8829_ ;
	wire _w8830_ ;
	wire _w8831_ ;
	wire _w8832_ ;
	wire _w8833_ ;
	wire _w8834_ ;
	wire _w8835_ ;
	wire _w8836_ ;
	wire _w8837_ ;
	wire _w8838_ ;
	wire _w8839_ ;
	wire _w8840_ ;
	wire _w8841_ ;
	wire _w8842_ ;
	wire _w8843_ ;
	wire _w8844_ ;
	wire _w8845_ ;
	wire _w8846_ ;
	wire _w8847_ ;
	wire _w8848_ ;
	wire _w8849_ ;
	wire _w8850_ ;
	wire _w8851_ ;
	wire _w8852_ ;
	wire _w8853_ ;
	wire _w8854_ ;
	wire _w8855_ ;
	wire _w8856_ ;
	wire _w8857_ ;
	wire _w8858_ ;
	wire _w8859_ ;
	wire _w8860_ ;
	wire _w8861_ ;
	wire _w8862_ ;
	wire _w8863_ ;
	wire _w8864_ ;
	wire _w8865_ ;
	wire _w8866_ ;
	wire _w8867_ ;
	wire _w8868_ ;
	wire _w8869_ ;
	wire _w8870_ ;
	wire _w8871_ ;
	wire _w8872_ ;
	wire _w8873_ ;
	wire _w8874_ ;
	wire _w8875_ ;
	wire _w8876_ ;
	wire _w8877_ ;
	wire _w8878_ ;
	wire _w8879_ ;
	wire _w8880_ ;
	wire _w8881_ ;
	wire _w8882_ ;
	wire _w8883_ ;
	wire _w8884_ ;
	wire _w8885_ ;
	wire _w8886_ ;
	wire _w8887_ ;
	wire _w8888_ ;
	wire _w8889_ ;
	wire _w8890_ ;
	wire _w8891_ ;
	wire _w8892_ ;
	wire _w8893_ ;
	wire _w8894_ ;
	wire _w8895_ ;
	wire _w8896_ ;
	wire _w8897_ ;
	wire _w8898_ ;
	wire _w8899_ ;
	wire _w8900_ ;
	wire _w8901_ ;
	wire _w8902_ ;
	wire _w8903_ ;
	wire _w8904_ ;
	wire _w8905_ ;
	wire _w8906_ ;
	wire _w8907_ ;
	wire _w8908_ ;
	wire _w8909_ ;
	wire _w8910_ ;
	wire _w8911_ ;
	wire _w8912_ ;
	wire _w8913_ ;
	wire _w8914_ ;
	wire _w8915_ ;
	wire _w8916_ ;
	wire _w8917_ ;
	wire _w8918_ ;
	wire _w8919_ ;
	wire _w8920_ ;
	wire _w8921_ ;
	wire _w8922_ ;
	wire _w8923_ ;
	wire _w8924_ ;
	wire _w8925_ ;
	wire _w8926_ ;
	wire _w8927_ ;
	wire _w8928_ ;
	wire _w8929_ ;
	wire _w8930_ ;
	wire _w8931_ ;
	wire _w8932_ ;
	wire _w8933_ ;
	wire _w8934_ ;
	wire _w8935_ ;
	wire _w8936_ ;
	wire _w8937_ ;
	wire _w8938_ ;
	wire _w8939_ ;
	wire _w8940_ ;
	wire _w8941_ ;
	wire _w8942_ ;
	wire _w8943_ ;
	wire _w8944_ ;
	wire _w8945_ ;
	wire _w8946_ ;
	wire _w8947_ ;
	wire _w8948_ ;
	wire _w8949_ ;
	wire _w8950_ ;
	wire _w8951_ ;
	wire _w8952_ ;
	wire _w8953_ ;
	wire _w8954_ ;
	wire _w8955_ ;
	wire _w8956_ ;
	wire _w8957_ ;
	wire _w8958_ ;
	wire _w8959_ ;
	wire _w8960_ ;
	wire _w8961_ ;
	wire _w8962_ ;
	wire _w8963_ ;
	wire _w8964_ ;
	wire _w8965_ ;
	wire _w8966_ ;
	wire _w8967_ ;
	wire _w8968_ ;
	wire _w8969_ ;
	wire _w8970_ ;
	wire _w8971_ ;
	wire _w8972_ ;
	wire _w8973_ ;
	wire _w8974_ ;
	wire _w8975_ ;
	wire _w8976_ ;
	wire _w8977_ ;
	wire _w8978_ ;
	wire _w8979_ ;
	wire _w8980_ ;
	wire _w8981_ ;
	wire _w8982_ ;
	wire _w8983_ ;
	wire _w8984_ ;
	wire _w8985_ ;
	wire _w8986_ ;
	wire _w8987_ ;
	wire _w8988_ ;
	wire _w8989_ ;
	wire _w8990_ ;
	wire _w8991_ ;
	wire _w8992_ ;
	wire _w8993_ ;
	wire _w8994_ ;
	wire _w8995_ ;
	wire _w8996_ ;
	wire _w8997_ ;
	wire _w8998_ ;
	wire _w8999_ ;
	wire _w9000_ ;
	wire _w9001_ ;
	wire _w9002_ ;
	wire _w9003_ ;
	wire _w9004_ ;
	wire _w9005_ ;
	wire _w9006_ ;
	wire _w9007_ ;
	wire _w9008_ ;
	wire _w9009_ ;
	wire _w9010_ ;
	wire _w9011_ ;
	wire _w9012_ ;
	wire _w9013_ ;
	wire _w9014_ ;
	wire _w9015_ ;
	wire _w9016_ ;
	wire _w9017_ ;
	wire _w9018_ ;
	wire _w9019_ ;
	wire _w9020_ ;
	wire _w9021_ ;
	wire _w9022_ ;
	wire _w9023_ ;
	wire _w9024_ ;
	wire _w9025_ ;
	wire _w9026_ ;
	wire _w9027_ ;
	wire _w9028_ ;
	wire _w9029_ ;
	wire _w9030_ ;
	wire _w9031_ ;
	wire _w9032_ ;
	wire _w9033_ ;
	wire _w9034_ ;
	wire _w9035_ ;
	wire _w9036_ ;
	wire _w9037_ ;
	wire _w9038_ ;
	wire _w9039_ ;
	wire _w9040_ ;
	wire _w9041_ ;
	wire _w9042_ ;
	wire _w9043_ ;
	wire _w9044_ ;
	wire _w9045_ ;
	wire _w9046_ ;
	wire _w9047_ ;
	wire _w9048_ ;
	wire _w9049_ ;
	wire _w9050_ ;
	wire _w9051_ ;
	wire _w9052_ ;
	wire _w9053_ ;
	wire _w9054_ ;
	wire _w9055_ ;
	wire _w9056_ ;
	wire _w9057_ ;
	wire _w9058_ ;
	wire _w9059_ ;
	wire _w9060_ ;
	wire _w9061_ ;
	wire _w9062_ ;
	wire _w9063_ ;
	wire _w9064_ ;
	wire _w9065_ ;
	wire _w9066_ ;
	wire _w9067_ ;
	wire _w9068_ ;
	wire _w9069_ ;
	wire _w9070_ ;
	wire _w9071_ ;
	wire _w9072_ ;
	wire _w9073_ ;
	wire _w9074_ ;
	wire _w9075_ ;
	wire _w9076_ ;
	wire _w9077_ ;
	wire _w9078_ ;
	wire _w9079_ ;
	wire _w9080_ ;
	wire _w9081_ ;
	wire _w9082_ ;
	wire _w9083_ ;
	wire _w9084_ ;
	wire _w9085_ ;
	wire _w9086_ ;
	wire _w9087_ ;
	wire _w9088_ ;
	wire _w9089_ ;
	wire _w9090_ ;
	wire _w9091_ ;
	wire _w9092_ ;
	wire _w9093_ ;
	wire _w9094_ ;
	wire _w9095_ ;
	wire _w9096_ ;
	wire _w9097_ ;
	wire _w9098_ ;
	wire _w9099_ ;
	wire _w9100_ ;
	wire _w9101_ ;
	wire _w9102_ ;
	wire _w9103_ ;
	wire _w9104_ ;
	wire _w9105_ ;
	wire _w9106_ ;
	wire _w9107_ ;
	wire _w9108_ ;
	wire _w9109_ ;
	wire _w9110_ ;
	wire _w9111_ ;
	wire _w9112_ ;
	wire _w9113_ ;
	wire _w9114_ ;
	wire _w9115_ ;
	wire _w9116_ ;
	wire _w9117_ ;
	wire _w9118_ ;
	wire _w9119_ ;
	wire _w9120_ ;
	wire _w9121_ ;
	wire _w9122_ ;
	wire _w9123_ ;
	wire _w9124_ ;
	wire _w9125_ ;
	wire _w9126_ ;
	wire _w9127_ ;
	wire _w9128_ ;
	wire _w9129_ ;
	wire _w9130_ ;
	wire _w9131_ ;
	wire _w9132_ ;
	wire _w9133_ ;
	wire _w14320_ ;
	wire _w14321_ ;
	wire _w14322_ ;
	wire _w14323_ ;
	wire _w14324_ ;
	wire _w14325_ ;
	wire _w14326_ ;
	wire _w14327_ ;
	wire _w14328_ ;
	wire _w14329_ ;
	wire _w14330_ ;
	wire _w14331_ ;
	wire _w14332_ ;
	wire _w14333_ ;
	wire _w14334_ ;
	wire _w14335_ ;
	wire _w14336_ ;
	wire _w14337_ ;
	wire _w14338_ ;
	wire _w14339_ ;
	wire _w14340_ ;
	wire _w14341_ ;
	wire _w14342_ ;
	wire _w14343_ ;
	wire _w14344_ ;
	wire _w14345_ ;
	wire _w14346_ ;
	wire _w14347_ ;
	wire _w14348_ ;
	wire _w14349_ ;
	wire _w14350_ ;
	wire _w14351_ ;
	wire _w14352_ ;
	wire _w14353_ ;
	wire _w14354_ ;
	wire _w14355_ ;
	wire _w14356_ ;
	wire _w14357_ ;
	wire _w14358_ ;
	wire _w14359_ ;
	wire _w14360_ ;
	wire _w14361_ ;
	wire _w14362_ ;
	wire _w14363_ ;
	wire _w14364_ ;
	wire _w14365_ ;
	wire _w14366_ ;
	wire _w14367_ ;
	wire _w14368_ ;
	wire _w14369_ ;
	wire _w14370_ ;
	wire _w14371_ ;
	wire _w14372_ ;
	wire _w14373_ ;
	wire _w14374_ ;
	wire _w14375_ ;
	wire _w14376_ ;
	wire _w14377_ ;
	wire _w14378_ ;
	wire _w14379_ ;
	wire _w14380_ ;
	wire _w14381_ ;
	wire _w14382_ ;
	wire _w14383_ ;
	wire _w14384_ ;
	wire _w14385_ ;
	wire _w14386_ ;
	wire _w14387_ ;
	wire _w14388_ ;
	wire _w14389_ ;
	wire _w14390_ ;
	wire _w14391_ ;
	wire _w14392_ ;
	wire _w14393_ ;
	wire _w14394_ ;
	wire _w14395_ ;
	wire _w14396_ ;
	wire _w14397_ ;
	wire _w14398_ ;
	wire _w14399_ ;
	wire _w14400_ ;
	wire _w14401_ ;
	wire _w14402_ ;
	wire _w14403_ ;
	wire _w14404_ ;
	wire _w14405_ ;
	wire _w14406_ ;
	wire _w14407_ ;
	wire _w14408_ ;
	wire _w14409_ ;
	wire _w14410_ ;
	wire _w14411_ ;
	wire _w14412_ ;
	wire _w14413_ ;
	wire _w14414_ ;
	wire _w14415_ ;
	wire _w14416_ ;
	wire _w14417_ ;
	wire _w14418_ ;
	wire _w14419_ ;
	wire _w14420_ ;
	wire _w14421_ ;
	wire _w14422_ ;
	wire _w14423_ ;
	wire _w14424_ ;
	wire _w14425_ ;
	wire _w14426_ ;
	wire _w14427_ ;
	wire _w14428_ ;
	wire _w14429_ ;
	wire _w14430_ ;
	wire _w14431_ ;
	wire _w14432_ ;
	wire _w14433_ ;
	wire _w14434_ ;
	wire _w14435_ ;
	wire _w14436_ ;
	wire _w14437_ ;
	wire _w14438_ ;
	wire _w14439_ ;
	wire _w14440_ ;
	wire _w14441_ ;
	wire _w14442_ ;
	wire _w14443_ ;
	wire _w14444_ ;
	wire _w14445_ ;
	wire _w14446_ ;
	wire _w14447_ ;
	wire _w14448_ ;
	wire _w14449_ ;
	wire _w14450_ ;
	wire _w14451_ ;
	wire _w14452_ ;
	wire _w14453_ ;
	wire _w14454_ ;
	wire _w14455_ ;
	wire _w14456_ ;
	wire _w14457_ ;
	wire _w14458_ ;
	wire _w14459_ ;
	wire _w14460_ ;
	wire _w14461_ ;
	wire _w14462_ ;
	wire _w14463_ ;
	wire _w14464_ ;
	wire _w14465_ ;
	wire _w14466_ ;
	wire _w14467_ ;
	wire _w14468_ ;
	wire _w14469_ ;
	wire _w14470_ ;
	wire _w14471_ ;
	wire _w14472_ ;
	wire _w14473_ ;
	wire _w14474_ ;
	wire _w14475_ ;
	wire _w14476_ ;
	wire _w14477_ ;
	wire _w14478_ ;
	wire _w14479_ ;
	wire _w14480_ ;
	wire _w14481_ ;
	wire _w14482_ ;
	wire _w14483_ ;
	wire _w14484_ ;
	wire _w14485_ ;
	wire _w14486_ ;
	wire _w14487_ ;
	wire _w14488_ ;
	wire _w14489_ ;
	wire _w14490_ ;
	wire _w14491_ ;
	wire _w14492_ ;
	wire _w14493_ ;
	wire _w14494_ ;
	wire _w14495_ ;
	wire _w14496_ ;
	wire _w14497_ ;
	wire _w14498_ ;
	wire _w14499_ ;
	wire _w14500_ ;
	wire _w14501_ ;
	wire _w14502_ ;
	wire _w14503_ ;
	wire _w14504_ ;
	wire _w14505_ ;
	wire _w14506_ ;
	wire _w14507_ ;
	wire _w14508_ ;
	wire _w14509_ ;
	wire _w14510_ ;
	wire _w14511_ ;
	wire _w14512_ ;
	wire _w14513_ ;
	wire _w14514_ ;
	wire _w14515_ ;
	wire _w14516_ ;
	wire _w14517_ ;
	wire _w14518_ ;
	wire _w14519_ ;
	wire _w14520_ ;
	wire _w14521_ ;
	wire _w14522_ ;
	wire _w14523_ ;
	wire _w14524_ ;
	wire _w14525_ ;
	wire _w14526_ ;
	wire _w14527_ ;
	wire _w14528_ ;
	wire _w14529_ ;
	wire _w14530_ ;
	wire _w14531_ ;
	wire _w14532_ ;
	wire _w14533_ ;
	wire _w14534_ ;
	wire _w14535_ ;
	wire _w14536_ ;
	wire _w14537_ ;
	wire _w14538_ ;
	wire _w14539_ ;
	wire _w14540_ ;
	wire _w14541_ ;
	wire _w14542_ ;
	wire _w14543_ ;
	wire _w14544_ ;
	wire _w14545_ ;
	wire _w14546_ ;
	wire _w14547_ ;
	wire _w14548_ ;
	wire _w14549_ ;
	wire _w14550_ ;
	wire _w14551_ ;
	wire _w14552_ ;
	wire _w14553_ ;
	wire _w14554_ ;
	wire _w14555_ ;
	wire _w14556_ ;
	wire _w14557_ ;
	wire _w14558_ ;
	wire _w14559_ ;
	wire _w14560_ ;
	wire _w14561_ ;
	wire _w14562_ ;
	wire _w14563_ ;
	wire _w14564_ ;
	wire _w14565_ ;
	wire _w14566_ ;
	wire _w14567_ ;
	wire _w14568_ ;
	wire _w14569_ ;
	wire _w14570_ ;
	wire _w14571_ ;
	wire _w14572_ ;
	wire _w14573_ ;
	wire _w14574_ ;
	wire _w14575_ ;
	wire _w14576_ ;
	wire _w14577_ ;
	wire _w14578_ ;
	wire _w14579_ ;
	wire _w14580_ ;
	wire _w14581_ ;
	wire _w14582_ ;
	wire _w14583_ ;
	wire _w14584_ ;
	wire _w14585_ ;
	wire _w14586_ ;
	wire _w14587_ ;
	wire _w14588_ ;
	wire _w14589_ ;
	wire _w14590_ ;
	wire _w14591_ ;
	wire _w14592_ ;
	wire _w14593_ ;
	wire _w14594_ ;
	wire _w14595_ ;
	wire _w14596_ ;
	wire _w14597_ ;
	wire _w14598_ ;
	wire _w14599_ ;
	wire _w14600_ ;
	wire _w14601_ ;
	wire _w14602_ ;
	wire _w14603_ ;
	wire _w14604_ ;
	wire _w14605_ ;
	wire _w14606_ ;
	wire _w14607_ ;
	wire _w14608_ ;
	wire _w14609_ ;
	wire _w14610_ ;
	wire _w14611_ ;
	wire _w14612_ ;
	wire _w14613_ ;
	wire _w14614_ ;
	wire _w14615_ ;
	wire _w14616_ ;
	wire _w14617_ ;
	wire _w14618_ ;
	wire _w14619_ ;
	wire _w14620_ ;
	wire _w14621_ ;
	wire _w14622_ ;
	wire _w14623_ ;
	wire _w14624_ ;
	wire _w14625_ ;
	wire _w14626_ ;
	wire _w14627_ ;
	wire _w14628_ ;
	wire _w14629_ ;
	wire _w14630_ ;
	wire _w14631_ ;
	wire _w14632_ ;
	wire _w14633_ ;
	wire _w14634_ ;
	wire _w14635_ ;
	wire _w14636_ ;
	wire _w14637_ ;
	wire _w14638_ ;
	wire _w14639_ ;
	wire _w14640_ ;
	wire _w14641_ ;
	wire _w14642_ ;
	wire _w14643_ ;
	wire _w14644_ ;
	wire _w14645_ ;
	wire _w14646_ ;
	wire _w14647_ ;
	wire _w14648_ ;
	wire _w14649_ ;
	wire _w14650_ ;
	wire _w14651_ ;
	wire _w14652_ ;
	wire _w14653_ ;
	wire _w14654_ ;
	wire _w14655_ ;
	wire _w14656_ ;
	wire _w14657_ ;
	wire _w14658_ ;
	wire _w14659_ ;
	wire _w14660_ ;
	wire _w14661_ ;
	wire _w14662_ ;
	wire _w14663_ ;
	wire _w14664_ ;
	wire _w14665_ ;
	wire _w14666_ ;
	wire _w14667_ ;
	wire _w14668_ ;
	wire _w14669_ ;
	wire _w14670_ ;
	wire _w14671_ ;
	wire _w14672_ ;
	wire _w14673_ ;
	wire _w14674_ ;
	wire _w14675_ ;
	wire _w14676_ ;
	wire _w14677_ ;
	wire _w14678_ ;
	wire _w14679_ ;
	wire _w14680_ ;
	wire _w14681_ ;
	wire _w14682_ ;
	wire _w14683_ ;
	wire _w14684_ ;
	wire _w14685_ ;
	wire _w14686_ ;
	wire _w14687_ ;
	wire _w14688_ ;
	wire _w14689_ ;
	wire _w14690_ ;
	wire _w14691_ ;
	wire _w14692_ ;
	wire _w14693_ ;
	wire _w14694_ ;
	wire _w14695_ ;
	wire _w14696_ ;
	wire _w14697_ ;
	wire _w14698_ ;
	wire _w14699_ ;
	wire _w14700_ ;
	wire _w14701_ ;
	wire _w14702_ ;
	wire _w14703_ ;
	wire _w14704_ ;
	wire _w14705_ ;
	wire _w14706_ ;
	wire _w14707_ ;
	wire _w14708_ ;
	wire _w14709_ ;
	wire _w14710_ ;
	wire _w14711_ ;
	wire _w14712_ ;
	wire _w14713_ ;
	wire _w14714_ ;
	wire _w14715_ ;
	wire _w14716_ ;
	wire _w14717_ ;
	wire _w14718_ ;
	wire _w14719_ ;
	wire _w14720_ ;
	wire _w14721_ ;
	wire _w14722_ ;
	wire _w14723_ ;
	wire _w14724_ ;
	wire _w14725_ ;
	wire _w14726_ ;
	wire _w14727_ ;
	wire _w14728_ ;
	wire _w14729_ ;
	wire _w14730_ ;
	wire _w14731_ ;
	wire _w14732_ ;
	wire _w14733_ ;
	wire _w14734_ ;
	wire _w14735_ ;
	wire _w14736_ ;
	wire _w14737_ ;
	wire _w14738_ ;
	wire _w14739_ ;
	wire _w14740_ ;
	wire _w14741_ ;
	wire _w14742_ ;
	wire _w14743_ ;
	wire _w14744_ ;
	wire _w14745_ ;
	wire _w14746_ ;
	wire _w14747_ ;
	wire _w14748_ ;
	wire _w14749_ ;
	wire _w14750_ ;
	wire _w14751_ ;
	wire _w14752_ ;
	wire _w14753_ ;
	wire _w14754_ ;
	wire _w14755_ ;
	wire _w14756_ ;
	wire _w14757_ ;
	wire _w14758_ ;
	wire _w14759_ ;
	wire _w14760_ ;
	wire _w14761_ ;
	wire _w14762_ ;
	wire _w14763_ ;
	wire _w14764_ ;
	wire _w14765_ ;
	wire _w14766_ ;
	wire _w14767_ ;
	wire _w14768_ ;
	wire _w14769_ ;
	wire _w14770_ ;
	wire _w14771_ ;
	wire _w14772_ ;
	wire _w14773_ ;
	wire _w14774_ ;
	wire _w14775_ ;
	wire _w14776_ ;
	wire _w14777_ ;
	wire _w14778_ ;
	wire _w14779_ ;
	wire _w14780_ ;
	wire _w14781_ ;
	wire _w14782_ ;
	wire _w14783_ ;
	wire _w14784_ ;
	wire _w14785_ ;
	wire _w14786_ ;
	wire _w14787_ ;
	wire _w14788_ ;
	wire _w14789_ ;
	wire _w14790_ ;
	wire _w14791_ ;
	wire _w14792_ ;
	wire _w14793_ ;
	wire _w14794_ ;
	wire _w14795_ ;
	wire _w14796_ ;
	wire _w14797_ ;
	wire _w14798_ ;
	wire _w14799_ ;
	wire _w14800_ ;
	wire _w14801_ ;
	wire _w14802_ ;
	wire _w14803_ ;
	wire _w14804_ ;
	wire _w14805_ ;
	wire _w14806_ ;
	wire _w14807_ ;
	wire _w14808_ ;
	wire _w14809_ ;
	wire _w14810_ ;
	wire _w14811_ ;
	wire _w14812_ ;
	wire _w14813_ ;
	wire _w14814_ ;
	wire _w14815_ ;
	wire _w14816_ ;
	wire _w14817_ ;
	wire _w14818_ ;
	wire _w14819_ ;
	wire _w14820_ ;
	wire _w14821_ ;
	wire _w14822_ ;
	wire _w14823_ ;
	wire _w14824_ ;
	wire _w14825_ ;
	wire _w14826_ ;
	wire _w14827_ ;
	wire _w14828_ ;
	wire _w14829_ ;
	wire _w14830_ ;
	wire _w14831_ ;
	wire _w14832_ ;
	wire _w14833_ ;
	wire _w14834_ ;
	wire _w14835_ ;
	wire _w14836_ ;
	wire _w14837_ ;
	wire _w14838_ ;
	wire _w14839_ ;
	wire _w14840_ ;
	wire _w14841_ ;
	wire _w14842_ ;
	wire _w14843_ ;
	wire _w14844_ ;
	wire _w14845_ ;
	wire _w14846_ ;
	wire _w14847_ ;
	wire _w14848_ ;
	wire _w14849_ ;
	wire _w14850_ ;
	wire _w14851_ ;
	wire _w14852_ ;
	wire _w14853_ ;
	wire _w14854_ ;
	wire _w14855_ ;
	wire _w14856_ ;
	wire _w14857_ ;
	wire _w14858_ ;
	wire _w14859_ ;
	wire _w14860_ ;
	wire _w14861_ ;
	wire _w14862_ ;
	wire _w14863_ ;
	wire _w14864_ ;
	wire _w14865_ ;
	wire _w14866_ ;
	wire _w14867_ ;
	wire _w14868_ ;
	wire _w14869_ ;
	wire _w14870_ ;
	wire _w14871_ ;
	wire _w14872_ ;
	wire _w14873_ ;
	wire _w14874_ ;
	wire _w14875_ ;
	wire _w14876_ ;
	wire _w14877_ ;
	wire _w14878_ ;
	wire _w14879_ ;
	wire _w14880_ ;
	wire _w14881_ ;
	wire _w14882_ ;
	wire _w14883_ ;
	wire _w14884_ ;
	wire _w14885_ ;
	wire _w14886_ ;
	wire _w14887_ ;
	wire _w14888_ ;
	wire _w14889_ ;
	wire _w14890_ ;
	wire _w14891_ ;
	wire _w14892_ ;
	wire _w14893_ ;
	wire _w14894_ ;
	wire _w14895_ ;
	wire _w14896_ ;
	wire _w14897_ ;
	wire _w14898_ ;
	wire _w14899_ ;
	wire _w14900_ ;
	wire _w14901_ ;
	wire _w14902_ ;
	wire _w14903_ ;
	wire _w14904_ ;
	wire _w14905_ ;
	wire _w14906_ ;
	wire _w14907_ ;
	wire _w14908_ ;
	wire _w14909_ ;
	wire _w14910_ ;
	wire _w14911_ ;
	wire _w14912_ ;
	wire _w14913_ ;
	wire _w14914_ ;
	wire _w14915_ ;
	wire _w14916_ ;
	wire _w14917_ ;
	wire _w14918_ ;
	wire _w14919_ ;
	wire _w14920_ ;
	wire _w14921_ ;
	wire _w14922_ ;
	wire _w14923_ ;
	wire _w14924_ ;
	wire _w14925_ ;
	wire _w14926_ ;
	wire _w14927_ ;
	wire _w14928_ ;
	wire _w14929_ ;
	wire _w14930_ ;
	wire _w14931_ ;
	wire _w14932_ ;
	wire _w14933_ ;
	wire _w14934_ ;
	wire _w14935_ ;
	wire _w14936_ ;
	wire _w14937_ ;
	wire _w14938_ ;
	wire _w14939_ ;
	wire _w14940_ ;
	wire _w14941_ ;
	wire _w14942_ ;
	wire _w14943_ ;
	wire _w14944_ ;
	wire _w14945_ ;
	wire _w14946_ ;
	wire _w14947_ ;
	wire _w14948_ ;
	wire _w14949_ ;
	wire _w14950_ ;
	wire _w14951_ ;
	wire _w14952_ ;
	wire _w14953_ ;
	wire _w14954_ ;
	wire _w14955_ ;
	wire _w14956_ ;
	wire _w14957_ ;
	wire _w14958_ ;
	wire _w14959_ ;
	wire _w14960_ ;
	wire _w14961_ ;
	wire _w14962_ ;
	wire _w14963_ ;
	wire _w14964_ ;
	wire _w14965_ ;
	wire _w14966_ ;
	wire _w14967_ ;
	wire _w14968_ ;
	wire _w14969_ ;
	wire _w14970_ ;
	wire _w14971_ ;
	wire _w14972_ ;
	wire _w14973_ ;
	wire _w14974_ ;
	wire _w14975_ ;
	wire _w14976_ ;
	wire _w14977_ ;
	wire _w14978_ ;
	wire _w14979_ ;
	wire _w14980_ ;
	wire _w14981_ ;
	wire _w14982_ ;
	wire _w14983_ ;
	wire _w14984_ ;
	wire _w14985_ ;
	wire _w14986_ ;
	wire _w14987_ ;
	wire _w14988_ ;
	wire _w14989_ ;
	wire _w14990_ ;
	wire _w14991_ ;
	wire _w14992_ ;
	wire _w14993_ ;
	wire _w14994_ ;
	wire _w14995_ ;
	wire _w14996_ ;
	wire _w14997_ ;
	wire _w14998_ ;
	wire _w14999_ ;
	wire _w15000_ ;
	wire _w15001_ ;
	wire _w15002_ ;
	wire _w15003_ ;
	wire _w15004_ ;
	wire _w15005_ ;
	wire _w15006_ ;
	wire _w15007_ ;
	wire _w15008_ ;
	wire _w15009_ ;
	wire _w15010_ ;
	wire _w15011_ ;
	wire _w15012_ ;
	wire _w15013_ ;
	wire _w15014_ ;
	wire _w15015_ ;
	wire _w15016_ ;
	wire _w15017_ ;
	wire _w15018_ ;
	wire _w15019_ ;
	wire _w15020_ ;
	wire _w15021_ ;
	wire _w15022_ ;
	wire _w15023_ ;
	wire _w15024_ ;
	wire _w15025_ ;
	wire _w15026_ ;
	wire _w15027_ ;
	wire _w15028_ ;
	wire _w15029_ ;
	wire _w15030_ ;
	wire _w15031_ ;
	wire _w15032_ ;
	wire _w15033_ ;
	wire _w15034_ ;
	wire _w15035_ ;
	wire _w15036_ ;
	wire _w15037_ ;
	wire _w15038_ ;
	wire _w15039_ ;
	wire _w15040_ ;
	wire _w15041_ ;
	wire _w15042_ ;
	wire _w15043_ ;
	wire _w15044_ ;
	wire _w15045_ ;
	wire _w15046_ ;
	wire _w15047_ ;
	wire _w15048_ ;
	wire _w15049_ ;
	wire _w15050_ ;
	wire _w15051_ ;
	wire _w15052_ ;
	wire _w15053_ ;
	wire _w15054_ ;
	wire _w15055_ ;
	wire _w15056_ ;
	wire _w15057_ ;
	wire _w15058_ ;
	wire _w15059_ ;
	wire _w15060_ ;
	wire _w15061_ ;
	wire _w15062_ ;
	wire _w15063_ ;
	wire _w15064_ ;
	wire _w15065_ ;
	wire _w15066_ ;
	wire _w15067_ ;
	wire _w15068_ ;
	wire _w15069_ ;
	wire _w15070_ ;
	wire _w15071_ ;
	wire _w15072_ ;
	wire _w15073_ ;
	wire _w15074_ ;
	wire _w15075_ ;
	wire _w15076_ ;
	wire _w15077_ ;
	wire _w15078_ ;
	wire _w15079_ ;
	wire _w15080_ ;
	wire _w15081_ ;
	wire _w15082_ ;
	wire _w15083_ ;
	wire _w15084_ ;
	wire _w15085_ ;
	wire _w15086_ ;
	wire _w15087_ ;
	wire _w15088_ ;
	wire _w15089_ ;
	wire _w15090_ ;
	wire _w15091_ ;
	wire _w15092_ ;
	wire _w15093_ ;
	wire _w15094_ ;
	wire _w15095_ ;
	wire _w15096_ ;
	wire _w15097_ ;
	wire _w15098_ ;
	wire _w15099_ ;
	wire _w15100_ ;
	wire _w15101_ ;
	wire _w15102_ ;
	wire _w15103_ ;
	wire _w15104_ ;
	wire _w15105_ ;
	wire _w15106_ ;
	wire _w15107_ ;
	wire _w15108_ ;
	wire _w15109_ ;
	wire _w15110_ ;
	wire _w15111_ ;
	wire _w15112_ ;
	wire _w15113_ ;
	wire _w15114_ ;
	wire _w15115_ ;
	wire _w15116_ ;
	wire _w15117_ ;
	wire _w15118_ ;
	wire _w15119_ ;
	wire _w15120_ ;
	wire _w15121_ ;
	wire _w15122_ ;
	wire _w15123_ ;
	wire _w15124_ ;
	wire _w15125_ ;
	wire _w15126_ ;
	wire _w15127_ ;
	wire _w15128_ ;
	wire _w15129_ ;
	wire _w15130_ ;
	wire _w15131_ ;
	wire _w15132_ ;
	wire _w15133_ ;
	wire _w15134_ ;
	wire _w15135_ ;
	wire _w15136_ ;
	wire _w15137_ ;
	wire _w15138_ ;
	wire _w15139_ ;
	wire _w15140_ ;
	wire _w15141_ ;
	wire _w15142_ ;
	wire _w15143_ ;
	wire _w15144_ ;
	wire _w15145_ ;
	wire _w15146_ ;
	wire _w15147_ ;
	wire _w15148_ ;
	wire _w15149_ ;
	wire _w15150_ ;
	wire _w15151_ ;
	wire _w15152_ ;
	wire _w15153_ ;
	wire _w15154_ ;
	wire _w15155_ ;
	wire _w15156_ ;
	wire _w15157_ ;
	wire _w15158_ ;
	wire _w15159_ ;
	wire _w15160_ ;
	wire _w15161_ ;
	wire _w15162_ ;
	wire _w15163_ ;
	wire _w15164_ ;
	wire _w15165_ ;
	wire _w15166_ ;
	wire _w15167_ ;
	wire _w15168_ ;
	wire _w15169_ ;
	wire _w15170_ ;
	wire _w15171_ ;
	wire _w15172_ ;
	wire _w15173_ ;
	wire _w15174_ ;
	wire _w15175_ ;
	wire _w15176_ ;
	wire _w15177_ ;
	wire _w15178_ ;
	wire _w15179_ ;
	wire _w15180_ ;
	wire _w15181_ ;
	wire _w15182_ ;
	wire _w15183_ ;
	wire _w15184_ ;
	wire _w15185_ ;
	wire _w15186_ ;
	wire _w15187_ ;
	wire _w15188_ ;
	wire _w15189_ ;
	wire _w15190_ ;
	wire _w15191_ ;
	wire _w15192_ ;
	wire _w15193_ ;
	wire _w15194_ ;
	wire _w15195_ ;
	wire _w15196_ ;
	wire _w15197_ ;
	wire _w15198_ ;
	wire _w15199_ ;
	wire _w15200_ ;
	wire _w15201_ ;
	wire _w15202_ ;
	wire _w15203_ ;
	wire _w15204_ ;
	wire _w15205_ ;
	wire _w15206_ ;
	wire _w15207_ ;
	wire _w15208_ ;
	wire _w15209_ ;
	wire _w15210_ ;
	wire _w15211_ ;
	wire _w15212_ ;
	wire _w15213_ ;
	wire _w15214_ ;
	wire _w15215_ ;
	wire _w15216_ ;
	wire _w15217_ ;
	wire _w15218_ ;
	wire _w15219_ ;
	wire _w15220_ ;
	wire _w15221_ ;
	wire _w15222_ ;
	wire _w15223_ ;
	wire _w15224_ ;
	wire _w15225_ ;
	wire _w15226_ ;
	wire _w15227_ ;
	wire _w15228_ ;
	wire _w15229_ ;
	wire _w15230_ ;
	wire _w15231_ ;
	wire _w15232_ ;
	wire _w15233_ ;
	wire _w15234_ ;
	wire _w15235_ ;
	wire _w15236_ ;
	wire _w15237_ ;
	wire _w15238_ ;
	wire _w15239_ ;
	wire _w15240_ ;
	wire _w15241_ ;
	wire _w15242_ ;
	wire _w15243_ ;
	wire _w15244_ ;
	wire _w15245_ ;
	wire _w15246_ ;
	wire _w15247_ ;
	wire _w15248_ ;
	wire _w15249_ ;
	wire _w15250_ ;
	wire _w15251_ ;
	wire _w15252_ ;
	wire _w15253_ ;
	wire _w15254_ ;
	wire _w15255_ ;
	wire _w15256_ ;
	wire _w15257_ ;
	wire _w15258_ ;
	wire _w15259_ ;
	wire _w15260_ ;
	wire _w15261_ ;
	wire _w15262_ ;
	wire _w15263_ ;
	wire _w15264_ ;
	wire _w15265_ ;
	wire _w15266_ ;
	wire _w15267_ ;
	wire _w15268_ ;
	wire _w15269_ ;
	wire _w15270_ ;
	wire _w15271_ ;
	wire _w15272_ ;
	wire _w15273_ ;
	wire _w15274_ ;
	wire _w15275_ ;
	wire _w15276_ ;
	wire _w15277_ ;
	wire _w15278_ ;
	wire _w15279_ ;
	wire _w15280_ ;
	wire _w15281_ ;
	wire _w15282_ ;
	wire _w15283_ ;
	wire _w15284_ ;
	wire _w15285_ ;
	wire _w15286_ ;
	wire _w15287_ ;
	wire _w15288_ ;
	wire _w15289_ ;
	wire _w15290_ ;
	wire _w15291_ ;
	wire _w15292_ ;
	wire _w15293_ ;
	wire _w15294_ ;
	wire _w15295_ ;
	wire _w15296_ ;
	wire _w15297_ ;
	wire _w15298_ ;
	wire _w15299_ ;
	wire _w15300_ ;
	wire _w15301_ ;
	wire _w15302_ ;
	wire _w15303_ ;
	wire _w15304_ ;
	wire _w15305_ ;
	wire _w15306_ ;
	wire _w15307_ ;
	wire _w15308_ ;
	wire _w15309_ ;
	wire _w15310_ ;
	wire _w15311_ ;
	wire _w15312_ ;
	wire _w15313_ ;
	wire _w15314_ ;
	wire _w15315_ ;
	wire _w15316_ ;
	wire _w15317_ ;
	wire _w15318_ ;
	wire _w15319_ ;
	wire _w15320_ ;
	wire _w15321_ ;
	wire _w15322_ ;
	wire _w15323_ ;
	wire _w15324_ ;
	wire _w15325_ ;
	wire _w15326_ ;
	wire _w15327_ ;
	wire _w15328_ ;
	wire _w15329_ ;
	wire _w15330_ ;
	wire _w15331_ ;
	wire _w15332_ ;
	wire _w15333_ ;
	wire _w15334_ ;
	wire _w15335_ ;
	wire _w15336_ ;
	wire _w15337_ ;
	wire _w15338_ ;
	wire _w15339_ ;
	wire _w15340_ ;
	wire _w15341_ ;
	wire _w15342_ ;
	wire _w15343_ ;
	wire _w15344_ ;
	wire _w15345_ ;
	wire _w15346_ ;
	wire _w15347_ ;
	wire _w15348_ ;
	wire _w15349_ ;
	wire _w15350_ ;
	wire _w15351_ ;
	wire _w15352_ ;
	wire _w15353_ ;
	wire _w15354_ ;
	wire _w15355_ ;
	wire _w15356_ ;
	wire _w15357_ ;
	wire _w15358_ ;
	wire _w15359_ ;
	wire _w15360_ ;
	wire _w15361_ ;
	wire _w15362_ ;
	wire _w15363_ ;
	wire _w15364_ ;
	wire _w15365_ ;
	wire _w15366_ ;
	wire _w15367_ ;
	wire _w15368_ ;
	wire _w15369_ ;
	wire _w15370_ ;
	wire _w15371_ ;
	wire _w15372_ ;
	wire _w15373_ ;
	wire _w15374_ ;
	wire _w15375_ ;
	wire _w15376_ ;
	wire _w15377_ ;
	wire _w15378_ ;
	wire _w15379_ ;
	wire _w15380_ ;
	wire _w15381_ ;
	wire _w15382_ ;
	wire _w15383_ ;
	wire _w15384_ ;
	wire _w15385_ ;
	wire _w15386_ ;
	wire _w15387_ ;
	wire _w15388_ ;
	wire _w15389_ ;
	wire _w15390_ ;
	wire _w15391_ ;
	wire _w15392_ ;
	wire _w15393_ ;
	wire _w15394_ ;
	wire _w15395_ ;
	wire _w15396_ ;
	wire _w15397_ ;
	wire _w15398_ ;
	wire _w15399_ ;
	wire _w15400_ ;
	wire _w15401_ ;
	wire _w15402_ ;
	wire _w15403_ ;
	wire _w15404_ ;
	wire _w15405_ ;
	wire _w15406_ ;
	wire _w15407_ ;
	wire _w15408_ ;
	wire _w15409_ ;
	wire _w15410_ ;
	wire _w15411_ ;
	wire _w15412_ ;
	wire _w15413_ ;
	wire _w15414_ ;
	wire _w15415_ ;
	wire _w15416_ ;
	wire _w15417_ ;
	wire _w15418_ ;
	wire _w15419_ ;
	wire _w15420_ ;
	wire _w15421_ ;
	wire _w15422_ ;
	wire _w15423_ ;
	wire _w15424_ ;
	wire _w15425_ ;
	wire _w15426_ ;
	wire _w15427_ ;
	wire _w15428_ ;
	wire _w15429_ ;
	wire _w15430_ ;
	wire _w15431_ ;
	wire _w15432_ ;
	wire _w15433_ ;
	wire _w15434_ ;
	wire _w15435_ ;
	wire _w15436_ ;
	wire _w15437_ ;
	wire _w15438_ ;
	wire _w15439_ ;
	wire _w15440_ ;
	wire _w15441_ ;
	wire _w15442_ ;
	wire _w15443_ ;
	wire _w15444_ ;
	wire _w15445_ ;
	wire _w15446_ ;
	wire _w15447_ ;
	wire _w15448_ ;
	wire _w15449_ ;
	wire _w15450_ ;
	wire _w15451_ ;
	wire _w15452_ ;
	wire _w15453_ ;
	wire _w15454_ ;
	wire _w15455_ ;
	wire _w15456_ ;
	wire _w15457_ ;
	wire _w15458_ ;
	wire _w15459_ ;
	wire _w15460_ ;
	wire _w15461_ ;
	wire _w15462_ ;
	wire _w15463_ ;
	wire _w15464_ ;
	wire _w15465_ ;
	wire _w15466_ ;
	wire _w15467_ ;
	wire _w15468_ ;
	wire _w15469_ ;
	wire _w15470_ ;
	wire _w15471_ ;
	wire _w15472_ ;
	wire _w15473_ ;
	wire _w15474_ ;
	wire _w15475_ ;
	wire _w15476_ ;
	wire _w15477_ ;
	wire _w15478_ ;
	wire _w15479_ ;
	wire _w15480_ ;
	wire _w15481_ ;
	wire _w15482_ ;
	wire _w15483_ ;
	wire _w15484_ ;
	wire _w15485_ ;
	wire _w15486_ ;
	wire _w15487_ ;
	wire _w15488_ ;
	wire _w15489_ ;
	wire _w15490_ ;
	wire _w15491_ ;
	wire _w15492_ ;
	wire _w15493_ ;
	wire _w15494_ ;
	wire _w15495_ ;
	wire _w15496_ ;
	wire _w15497_ ;
	wire _w15498_ ;
	wire _w15499_ ;
	wire _w15500_ ;
	wire _w15501_ ;
	wire _w15502_ ;
	wire _w15503_ ;
	wire _w15504_ ;
	wire _w15505_ ;
	wire _w15506_ ;
	wire _w15507_ ;
	wire _w15508_ ;
	wire _w15509_ ;
	wire _w15510_ ;
	wire _w15511_ ;
	wire _w15512_ ;
	wire _w15513_ ;
	wire _w15514_ ;
	wire _w15515_ ;
	wire _w15516_ ;
	wire _w15517_ ;
	wire _w15518_ ;
	wire _w15519_ ;
	wire _w15520_ ;
	wire _w15521_ ;
	wire _w15522_ ;
	wire _w15523_ ;
	wire _w15524_ ;
	wire _w15525_ ;
	wire _w15526_ ;
	wire _w15527_ ;
	wire _w15528_ ;
	wire _w15529_ ;
	wire _w15530_ ;
	wire _w15531_ ;
	wire _w15532_ ;
	wire _w15533_ ;
	wire _w15534_ ;
	wire _w15535_ ;
	wire _w15536_ ;
	wire _w15537_ ;
	wire _w15538_ ;
	wire _w15539_ ;
	wire _w15540_ ;
	wire _w15541_ ;
	wire _w15542_ ;
	wire _w15543_ ;
	wire _w15544_ ;
	wire _w15545_ ;
	wire _w15546_ ;
	wire _w15547_ ;
	wire _w15548_ ;
	wire _w15549_ ;
	wire _w15550_ ;
	wire _w15551_ ;
	wire _w15552_ ;
	wire _w15553_ ;
	wire _w15554_ ;
	wire _w15555_ ;
	wire _w15556_ ;
	wire _w15557_ ;
	wire _w15558_ ;
	wire _w15559_ ;
	wire _w15560_ ;
	wire _w15561_ ;
	wire _w15562_ ;
	wire _w15563_ ;
	wire _w15564_ ;
	wire _w15565_ ;
	wire _w15566_ ;
	wire _w15567_ ;
	wire _w15568_ ;
	wire _w15569_ ;
	wire _w15570_ ;
	wire _w15571_ ;
	wire _w15572_ ;
	wire _w15573_ ;
	wire _w15574_ ;
	wire _w15575_ ;
	wire _w15576_ ;
	wire _w15577_ ;
	wire _w15578_ ;
	wire _w15579_ ;
	wire _w15580_ ;
	wire _w15581_ ;
	wire _w15582_ ;
	wire _w15583_ ;
	wire _w15584_ ;
	wire _w15585_ ;
	wire _w15586_ ;
	wire _w15587_ ;
	wire _w15588_ ;
	wire _w15589_ ;
	wire _w15590_ ;
	wire _w15591_ ;
	wire _w15592_ ;
	wire _w15593_ ;
	wire _w15594_ ;
	wire _w15595_ ;
	wire _w15596_ ;
	wire _w15597_ ;
	wire _w15598_ ;
	wire _w15599_ ;
	wire _w15600_ ;
	wire _w15601_ ;
	wire _w15602_ ;
	wire _w15603_ ;
	wire _w15604_ ;
	wire _w15605_ ;
	wire _w15606_ ;
	wire _w15607_ ;
	wire _w15608_ ;
	wire _w15609_ ;
	wire _w15610_ ;
	wire _w15611_ ;
	wire _w15612_ ;
	wire _w15613_ ;
	wire _w15614_ ;
	wire _w15615_ ;
	wire _w15616_ ;
	wire _w15617_ ;
	wire _w15618_ ;
	wire _w15619_ ;
	wire _w15620_ ;
	wire _w15621_ ;
	wire _w15622_ ;
	wire _w15623_ ;
	wire _w15624_ ;
	wire _w15625_ ;
	wire _w15626_ ;
	wire _w15627_ ;
	wire _w15628_ ;
	wire _w15629_ ;
	wire _w15630_ ;
	wire _w15631_ ;
	wire _w15632_ ;
	wire _w15633_ ;
	wire _w15634_ ;
	wire _w15635_ ;
	wire _w15636_ ;
	wire _w15637_ ;
	wire _w15638_ ;
	wire _w15639_ ;
	wire _w15640_ ;
	wire _w15641_ ;
	wire _w15642_ ;
	wire _w15643_ ;
	wire _w15644_ ;
	wire _w15645_ ;
	wire _w15646_ ;
	wire _w15647_ ;
	wire _w15648_ ;
	wire _w15649_ ;
	wire _w15650_ ;
	wire _w15651_ ;
	wire _w15652_ ;
	wire _w15653_ ;
	wire _w15654_ ;
	wire _w15655_ ;
	wire _w15656_ ;
	wire _w15657_ ;
	wire _w15658_ ;
	wire _w15659_ ;
	wire _w15660_ ;
	wire _w15661_ ;
	wire _w15662_ ;
	wire _w15663_ ;
	wire _w15664_ ;
	wire _w15665_ ;
	wire _w15666_ ;
	wire _w15667_ ;
	wire _w15668_ ;
	wire _w15669_ ;
	wire _w15670_ ;
	wire _w15671_ ;
	wire _w15672_ ;
	wire _w15673_ ;
	wire _w15674_ ;
	wire _w15675_ ;
	wire _w15676_ ;
	wire _w15677_ ;
	wire _w15678_ ;
	wire _w15679_ ;
	wire _w15680_ ;
	wire _w15681_ ;
	wire _w15682_ ;
	wire _w15683_ ;
	wire _w15684_ ;
	wire _w15685_ ;
	wire _w15686_ ;
	wire _w15687_ ;
	wire _w15688_ ;
	wire _w15689_ ;
	wire _w15690_ ;
	wire _w15691_ ;
	wire _w15692_ ;
	wire _w15693_ ;
	wire _w15694_ ;
	wire _w15695_ ;
	wire _w15696_ ;
	wire _w15697_ ;
	wire _w15698_ ;
	wire _w15699_ ;
	wire _w15700_ ;
	wire _w15701_ ;
	wire _w15702_ ;
	wire _w15703_ ;
	wire _w15704_ ;
	wire _w15705_ ;
	wire _w15706_ ;
	wire _w15707_ ;
	wire _w15708_ ;
	wire _w15709_ ;
	wire _w15710_ ;
	wire _w15711_ ;
	wire _w15712_ ;
	wire _w15713_ ;
	wire _w15714_ ;
	wire _w15715_ ;
	wire _w15716_ ;
	wire _w15717_ ;
	wire _w15718_ ;
	wire _w15719_ ;
	wire _w15720_ ;
	wire _w15721_ ;
	wire _w15722_ ;
	wire _w15723_ ;
	wire _w15724_ ;
	wire _w15725_ ;
	wire _w15726_ ;
	wire _w15727_ ;
	wire _w15728_ ;
	wire _w15729_ ;
	wire _w15730_ ;
	wire _w15731_ ;
	wire _w15732_ ;
	wire _w15733_ ;
	wire _w15734_ ;
	wire _w15735_ ;
	wire _w15736_ ;
	wire _w15737_ ;
	wire _w15738_ ;
	wire _w15739_ ;
	wire _w15740_ ;
	wire _w15741_ ;
	wire _w15742_ ;
	wire _w15743_ ;
	wire _w15744_ ;
	wire _w15745_ ;
	wire _w15746_ ;
	wire _w15747_ ;
	wire _w15748_ ;
	wire _w15749_ ;
	wire _w15750_ ;
	wire _w15751_ ;
	wire _w15752_ ;
	wire _w15753_ ;
	wire _w15754_ ;
	wire _w15755_ ;
	wire _w15756_ ;
	wire _w15757_ ;
	wire _w15758_ ;
	wire _w15759_ ;
	wire _w15760_ ;
	wire _w15761_ ;
	wire _w15762_ ;
	wire _w15763_ ;
	wire _w15764_ ;
	wire _w15765_ ;
	wire _w15766_ ;
	wire _w15767_ ;
	wire _w15768_ ;
	wire _w15769_ ;
	wire _w15770_ ;
	wire _w15771_ ;
	wire _w15772_ ;
	wire _w15773_ ;
	wire _w15774_ ;
	wire _w15775_ ;
	wire _w15776_ ;
	wire _w15777_ ;
	wire _w15778_ ;
	wire _w15779_ ;
	wire _w15780_ ;
	wire _w15781_ ;
	wire _w15782_ ;
	wire _w15783_ ;
	wire _w15784_ ;
	wire _w15785_ ;
	wire _w15786_ ;
	wire _w15787_ ;
	wire _w15788_ ;
	wire _w15789_ ;
	wire _w15790_ ;
	wire _w15791_ ;
	wire _w15792_ ;
	wire _w15793_ ;
	wire _w15794_ ;
	wire _w15795_ ;
	wire _w15796_ ;
	wire _w15797_ ;
	wire _w15798_ ;
	wire _w15799_ ;
	wire _w15800_ ;
	wire _w15801_ ;
	wire _w15802_ ;
	wire _w15803_ ;
	wire _w15804_ ;
	wire _w15805_ ;
	wire _w15806_ ;
	wire _w15807_ ;
	wire _w15808_ ;
	wire _w15809_ ;
	wire _w15810_ ;
	wire _w15811_ ;
	wire _w15812_ ;
	wire _w15813_ ;
	wire _w15814_ ;
	wire _w15815_ ;
	wire _w15816_ ;
	wire _w15817_ ;
	wire _w15818_ ;
	wire _w15819_ ;
	wire _w15820_ ;
	wire _w15821_ ;
	wire _w15822_ ;
	wire _w15823_ ;
	wire _w15824_ ;
	wire _w15825_ ;
	wire _w15826_ ;
	wire _w15827_ ;
	wire _w15828_ ;
	wire _w15829_ ;
	wire _w15830_ ;
	wire _w15831_ ;
	wire _w15832_ ;
	wire _w15833_ ;
	wire _w15834_ ;
	wire _w15835_ ;
	wire _w15836_ ;
	wire _w15837_ ;
	wire _w15838_ ;
	wire _w15839_ ;
	wire _w15840_ ;
	wire _w15841_ ;
	wire _w15842_ ;
	wire _w15843_ ;
	wire _w15844_ ;
	wire _w15845_ ;
	wire _w15846_ ;
	wire _w15847_ ;
	wire _w15848_ ;
	wire _w15849_ ;
	wire _w15850_ ;
	wire _w15851_ ;
	wire _w15852_ ;
	wire _w15853_ ;
	wire _w15854_ ;
	wire _w15855_ ;
	wire _w15856_ ;
	wire _w15857_ ;
	wire _w15858_ ;
	wire _w15859_ ;
	wire _w15860_ ;
	wire _w15861_ ;
	wire _w15862_ ;
	wire _w15863_ ;
	wire _w15864_ ;
	wire _w15865_ ;
	wire _w15866_ ;
	wire _w15867_ ;
	wire _w15868_ ;
	wire _w15869_ ;
	wire _w15870_ ;
	wire _w15871_ ;
	wire _w15872_ ;
	wire _w15873_ ;
	wire _w15874_ ;
	wire _w15875_ ;
	wire _w15876_ ;
	wire _w15877_ ;
	wire _w15878_ ;
	wire _w15879_ ;
	wire _w15880_ ;
	wire _w15881_ ;
	wire _w15882_ ;
	wire _w15883_ ;
	wire _w15884_ ;
	wire _w15885_ ;
	wire _w15886_ ;
	wire _w15887_ ;
	wire _w15888_ ;
	wire _w15889_ ;
	wire _w15890_ ;
	wire _w15891_ ;
	wire _w15892_ ;
	wire _w15893_ ;
	wire _w15894_ ;
	wire _w15895_ ;
	wire _w15896_ ;
	wire _w15897_ ;
	wire _w15898_ ;
	wire _w15899_ ;
	wire _w15900_ ;
	wire _w15901_ ;
	wire _w15902_ ;
	wire _w15903_ ;
	wire _w15904_ ;
	wire _w15905_ ;
	wire _w15906_ ;
	wire _w15907_ ;
	wire _w15908_ ;
	wire _w15909_ ;
	wire _w15910_ ;
	wire _w15911_ ;
	wire _w15912_ ;
	wire _w15913_ ;
	wire _w15914_ ;
	wire _w15915_ ;
	wire _w15916_ ;
	wire _w15917_ ;
	wire _w15918_ ;
	wire _w15919_ ;
	wire _w15920_ ;
	wire _w15921_ ;
	wire _w15922_ ;
	wire _w15923_ ;
	wire _w15924_ ;
	wire _w15925_ ;
	wire _w15926_ ;
	wire _w15927_ ;
	wire _w15928_ ;
	wire _w15929_ ;
	wire _w15930_ ;
	wire _w15931_ ;
	wire _w15932_ ;
	wire _w15933_ ;
	wire _w15934_ ;
	wire _w15935_ ;
	wire _w15936_ ;
	wire _w15937_ ;
	wire _w15938_ ;
	wire _w15939_ ;
	wire _w15940_ ;
	wire _w15941_ ;
	wire _w15942_ ;
	wire _w15943_ ;
	wire _w15944_ ;
	wire _w15945_ ;
	wire _w15946_ ;
	wire _w15947_ ;
	wire _w15948_ ;
	wire _w15949_ ;
	wire _w15950_ ;
	wire _w15951_ ;
	wire _w15952_ ;
	wire _w15953_ ;
	wire _w15954_ ;
	wire _w15955_ ;
	wire _w15956_ ;
	wire _w15957_ ;
	wire _w15958_ ;
	wire _w15959_ ;
	wire _w15960_ ;
	wire _w15961_ ;
	wire _w15962_ ;
	wire _w15963_ ;
	wire _w15964_ ;
	wire _w15965_ ;
	wire _w15966_ ;
	wire _w15967_ ;
	wire _w15968_ ;
	wire _w15969_ ;
	wire _w15970_ ;
	wire _w15971_ ;
	wire _w15972_ ;
	wire _w15973_ ;
	wire _w15974_ ;
	wire _w15975_ ;
	wire _w15976_ ;
	wire _w15977_ ;
	wire _w15978_ ;
	wire _w15979_ ;
	wire _w15980_ ;
	wire _w15981_ ;
	wire _w15982_ ;
	wire _w15983_ ;
	wire _w15984_ ;
	wire _w15985_ ;
	wire _w15986_ ;
	wire _w15987_ ;
	wire _w15988_ ;
	wire _w15989_ ;
	wire _w15990_ ;
	wire _w15991_ ;
	wire _w15992_ ;
	wire _w15993_ ;
	wire _w15994_ ;
	wire _w15995_ ;
	wire _w15996_ ;
	wire _w15997_ ;
	wire _w15998_ ;
	wire _w15999_ ;
	wire _w16000_ ;
	wire _w16001_ ;
	wire _w16002_ ;
	wire _w16003_ ;
	wire _w16004_ ;
	wire _w16005_ ;
	wire _w16006_ ;
	wire _w16007_ ;
	wire _w16008_ ;
	wire _w16009_ ;
	wire _w16010_ ;
	wire _w16011_ ;
	wire _w16012_ ;
	wire _w16013_ ;
	wire _w16014_ ;
	wire _w16015_ ;
	wire _w16016_ ;
	wire _w16017_ ;
	wire _w16018_ ;
	wire _w16019_ ;
	wire _w16020_ ;
	wire _w16021_ ;
	wire _w16022_ ;
	wire _w16023_ ;
	wire _w16024_ ;
	wire _w16025_ ;
	wire _w16026_ ;
	wire _w16027_ ;
	wire _w16028_ ;
	wire _w16029_ ;
	wire _w16030_ ;
	wire _w16031_ ;
	wire _w16032_ ;
	wire _w16033_ ;
	wire _w16034_ ;
	wire _w16035_ ;
	wire _w16036_ ;
	wire _w16037_ ;
	wire _w16038_ ;
	wire _w16039_ ;
	wire _w16040_ ;
	wire _w16041_ ;
	wire _w16042_ ;
	wire _w16043_ ;
	wire _w16044_ ;
	wire _w16045_ ;
	wire _w16046_ ;
	wire _w16047_ ;
	wire _w16048_ ;
	wire _w16049_ ;
	wire _w16050_ ;
	wire _w16051_ ;
	wire _w16052_ ;
	wire _w16053_ ;
	wire _w16054_ ;
	wire _w16055_ ;
	wire _w16056_ ;
	wire _w16057_ ;
	wire _w16058_ ;
	wire _w16059_ ;
	wire _w16060_ ;
	wire _w16061_ ;
	wire _w16062_ ;
	wire _w16063_ ;
	wire _w16064_ ;
	wire _w16065_ ;
	wire _w16066_ ;
	wire _w16067_ ;
	wire _w16068_ ;
	wire _w16069_ ;
	wire _w16070_ ;
	wire _w16071_ ;
	wire _w16072_ ;
	wire _w16073_ ;
	wire _w16074_ ;
	wire _w16075_ ;
	wire _w16076_ ;
	wire _w16077_ ;
	wire _w16078_ ;
	wire _w16079_ ;
	wire _w16080_ ;
	wire _w16081_ ;
	wire _w16082_ ;
	wire _w16083_ ;
	wire _w16084_ ;
	wire _w16085_ ;
	wire _w16086_ ;
	wire _w16087_ ;
	wire _w16088_ ;
	wire _w16089_ ;
	wire _w16090_ ;
	wire _w16091_ ;
	wire _w16092_ ;
	wire _w16093_ ;
	wire _w16094_ ;
	wire _w16095_ ;
	wire _w16096_ ;
	wire _w16097_ ;
	wire _w16098_ ;
	wire _w16099_ ;
	wire _w16100_ ;
	wire _w16101_ ;
	wire _w16102_ ;
	wire _w16103_ ;
	wire _w16104_ ;
	wire _w16105_ ;
	wire _w16106_ ;
	wire _w16107_ ;
	wire _w16108_ ;
	wire _w16109_ ;
	wire _w16110_ ;
	wire _w16111_ ;
	wire _w16112_ ;
	wire _w16113_ ;
	wire _w16114_ ;
	wire _w16115_ ;
	wire _w16116_ ;
	wire _w16117_ ;
	wire _w16118_ ;
	wire _w16119_ ;
	wire _w16120_ ;
	wire _w16121_ ;
	wire _w16122_ ;
	wire _w16123_ ;
	wire _w16124_ ;
	wire _w16125_ ;
	wire _w16126_ ;
	wire _w16127_ ;
	wire _w16128_ ;
	wire _w16129_ ;
	wire _w16130_ ;
	wire _w16131_ ;
	wire _w16132_ ;
	wire _w16133_ ;
	wire _w16134_ ;
	wire _w16135_ ;
	wire _w16136_ ;
	wire _w16137_ ;
	wire _w16138_ ;
	wire _w16139_ ;
	wire _w16140_ ;
	wire _w16141_ ;
	wire _w16142_ ;
	wire _w16143_ ;
	wire _w16144_ ;
	wire _w16145_ ;
	wire _w16146_ ;
	wire _w16147_ ;
	wire _w16148_ ;
	wire _w16149_ ;
	wire _w16150_ ;
	wire _w16151_ ;
	wire _w16152_ ;
	wire _w16153_ ;
	wire _w16154_ ;
	wire _w16155_ ;
	wire _w16156_ ;
	wire _w16157_ ;
	wire _w16158_ ;
	wire _w16159_ ;
	wire _w16160_ ;
	wire _w16161_ ;
	wire _w16162_ ;
	wire _w16163_ ;
	wire _w16164_ ;
	wire _w16165_ ;
	wire _w16166_ ;
	wire _w16167_ ;
	wire _w16168_ ;
	wire _w16169_ ;
	wire _w16170_ ;
	wire _w16171_ ;
	wire _w16172_ ;
	wire _w16173_ ;
	wire _w16174_ ;
	wire _w16175_ ;
	wire _w16176_ ;
	wire _w16177_ ;
	wire _w16178_ ;
	wire _w16179_ ;
	wire _w16180_ ;
	wire _w16181_ ;
	wire _w16182_ ;
	wire _w16183_ ;
	wire _w16184_ ;
	wire _w16185_ ;
	wire _w16186_ ;
	wire _w16187_ ;
	wire _w16188_ ;
	wire _w16189_ ;
	wire _w16190_ ;
	wire _w16191_ ;
	wire _w16192_ ;
	wire _w16193_ ;
	wire _w16194_ ;
	wire _w16195_ ;
	wire _w16196_ ;
	wire _w16197_ ;
	wire _w16198_ ;
	wire _w16199_ ;
	wire _w16200_ ;
	wire _w16201_ ;
	wire _w16202_ ;
	wire _w16203_ ;
	wire _w16204_ ;
	wire _w16205_ ;
	wire _w16206_ ;
	wire _w16207_ ;
	wire _w16208_ ;
	wire _w16209_ ;
	wire _w16210_ ;
	wire _w16211_ ;
	wire _w16212_ ;
	wire _w16213_ ;
	wire _w16214_ ;
	wire _w16215_ ;
	wire _w16216_ ;
	wire _w16217_ ;
	wire _w16218_ ;
	wire _w16219_ ;
	wire _w16220_ ;
	wire _w16221_ ;
	wire _w16222_ ;
	wire _w16223_ ;
	wire _w16224_ ;
	wire _w16225_ ;
	wire _w16226_ ;
	wire _w16227_ ;
	wire _w16228_ ;
	wire _w16229_ ;
	wire _w16230_ ;
	wire _w16231_ ;
	wire _w16232_ ;
	wire _w16233_ ;
	wire _w16234_ ;
	wire _w16235_ ;
	wire _w16236_ ;
	wire _w16237_ ;
	wire _w16238_ ;
	wire _w16239_ ;
	wire _w16240_ ;
	wire _w16241_ ;
	wire _w16242_ ;
	wire _w16243_ ;
	wire _w16244_ ;
	wire _w16245_ ;
	wire _w16246_ ;
	wire _w16247_ ;
	wire _w16248_ ;
	wire _w16249_ ;
	wire _w16250_ ;
	wire _w16251_ ;
	wire _w16252_ ;
	wire _w16253_ ;
	wire _w16254_ ;
	wire _w16255_ ;
	wire _w16256_ ;
	wire _w16257_ ;
	wire _w16258_ ;
	wire _w16259_ ;
	wire _w16260_ ;
	wire _w16261_ ;
	wire _w16262_ ;
	wire _w16263_ ;
	wire _w16264_ ;
	wire _w16265_ ;
	wire _w16266_ ;
	wire _w16267_ ;
	wire _w16268_ ;
	wire _w16269_ ;
	wire _w16270_ ;
	wire _w16271_ ;
	wire _w16272_ ;
	wire _w16273_ ;
	wire _w16274_ ;
	wire _w16275_ ;
	wire _w16276_ ;
	wire _w16277_ ;
	wire _w16278_ ;
	wire _w16279_ ;
	wire _w16280_ ;
	wire _w16281_ ;
	wire _w16282_ ;
	wire _w16283_ ;
	wire _w16284_ ;
	wire _w16285_ ;
	wire _w16286_ ;
	wire _w16287_ ;
	wire _w16288_ ;
	wire _w16289_ ;
	wire _w16290_ ;
	wire _w16291_ ;
	wire _w16292_ ;
	wire _w16293_ ;
	wire _w16294_ ;
	wire _w16295_ ;
	wire _w16296_ ;
	wire _w16297_ ;
	wire _w16298_ ;
	wire _w16299_ ;
	wire _w16300_ ;
	wire _w16301_ ;
	wire _w16302_ ;
	wire _w16303_ ;
	wire _w16304_ ;
	wire _w16305_ ;
	wire _w16306_ ;
	wire _w16307_ ;
	wire _w16308_ ;
	wire _w16309_ ;
	wire _w16310_ ;
	wire _w16311_ ;
	wire _w16312_ ;
	wire _w16313_ ;
	wire _w16314_ ;
	wire _w16315_ ;
	wire _w16316_ ;
	wire _w16317_ ;
	wire _w16318_ ;
	wire _w16319_ ;
	wire _w16320_ ;
	wire _w16321_ ;
	wire _w16322_ ;
	wire _w16323_ ;
	wire _w16324_ ;
	wire _w16325_ ;
	wire _w16326_ ;
	wire _w16327_ ;
	wire _w16328_ ;
	wire _w16329_ ;
	wire _w16330_ ;
	wire _w16331_ ;
	wire _w16332_ ;
	wire _w16333_ ;
	wire _w16334_ ;
	wire _w16335_ ;
	wire _w16336_ ;
	wire _w16337_ ;
	wire _w16338_ ;
	wire _w16339_ ;
	wire _w16340_ ;
	wire _w16341_ ;
	wire _w16342_ ;
	wire _w16343_ ;
	wire _w16344_ ;
	wire _w16345_ ;
	wire _w16346_ ;
	wire _w16347_ ;
	wire _w16348_ ;
	wire _w16349_ ;
	wire _w16350_ ;
	wire _w16351_ ;
	wire _w16352_ ;
	wire _w16353_ ;
	wire _w16354_ ;
	wire _w16355_ ;
	wire _w16356_ ;
	wire _w16357_ ;
	wire _w16358_ ;
	wire _w16359_ ;
	wire _w16360_ ;
	wire _w16361_ ;
	wire _w16362_ ;
	wire _w16363_ ;
	wire _w16364_ ;
	wire _w16365_ ;
	wire _w16366_ ;
	wire _w16367_ ;
	wire _w16368_ ;
	wire _w16369_ ;
	wire _w16370_ ;
	wire _w16371_ ;
	wire _w16372_ ;
	wire _w16373_ ;
	wire _w16374_ ;
	wire _w16375_ ;
	wire _w16376_ ;
	wire _w16377_ ;
	wire _w16378_ ;
	wire _w16379_ ;
	wire _w16380_ ;
	wire _w16381_ ;
	wire _w16382_ ;
	wire _w16383_ ;
	wire _w16384_ ;
	wire _w16385_ ;
	wire _w16386_ ;
	wire _w16387_ ;
	wire _w16388_ ;
	wire _w16389_ ;
	wire _w16390_ ;
	wire _w16391_ ;
	wire _w16392_ ;
	wire _w16393_ ;
	wire _w16394_ ;
	wire _w16395_ ;
	wire _w16396_ ;
	wire _w16397_ ;
	wire _w16398_ ;
	wire _w16399_ ;
	wire _w16400_ ;
	wire _w16401_ ;
	wire _w16402_ ;
	wire _w16403_ ;
	wire _w16404_ ;
	wire _w16405_ ;
	wire _w16406_ ;
	wire _w16407_ ;
	wire _w16408_ ;
	wire _w16409_ ;
	wire _w16410_ ;
	wire _w16411_ ;
	wire _w16412_ ;
	wire _w16413_ ;
	wire _w16414_ ;
	wire _w16415_ ;
	wire _w16416_ ;
	wire _w16417_ ;
	wire _w16418_ ;
	wire _w16419_ ;
	wire _w16420_ ;
	wire _w16421_ ;
	wire _w16422_ ;
	wire _w16423_ ;
	wire _w16424_ ;
	wire _w16425_ ;
	wire _w16426_ ;
	wire _w16427_ ;
	wire _w16428_ ;
	wire _w16429_ ;
	wire _w16430_ ;
	wire _w16431_ ;
	wire _w16432_ ;
	wire _w16433_ ;
	wire _w16434_ ;
	wire _w16435_ ;
	wire _w16436_ ;
	wire _w16437_ ;
	wire _w16438_ ;
	wire _w16439_ ;
	wire _w16440_ ;
	wire _w16441_ ;
	wire _w16442_ ;
	wire _w16443_ ;
	wire _w16444_ ;
	wire _w16445_ ;
	wire _w16446_ ;
	wire _w16447_ ;
	wire _w16448_ ;
	wire _w16449_ ;
	wire _w16450_ ;
	wire _w16451_ ;
	wire _w16452_ ;
	wire _w16453_ ;
	wire _w16454_ ;
	wire _w16455_ ;
	wire _w16456_ ;
	wire _w16457_ ;
	wire _w16458_ ;
	wire _w16459_ ;
	wire _w16460_ ;
	wire _w16461_ ;
	wire _w16462_ ;
	wire _w16463_ ;
	wire _w16464_ ;
	wire _w16465_ ;
	wire _w16466_ ;
	wire _w16467_ ;
	wire _w16468_ ;
	wire _w16469_ ;
	wire _w16470_ ;
	wire _w16471_ ;
	wire _w16472_ ;
	wire _w16473_ ;
	wire _w16474_ ;
	wire _w16475_ ;
	wire _w16476_ ;
	wire _w16477_ ;
	wire _w16478_ ;
	wire _w16479_ ;
	wire _w16480_ ;
	wire _w16481_ ;
	wire _w16482_ ;
	wire _w16483_ ;
	wire _w16484_ ;
	wire _w16485_ ;
	wire _w16486_ ;
	wire _w16487_ ;
	wire _w16488_ ;
	wire _w16489_ ;
	wire _w16490_ ;
	wire _w16491_ ;
	wire _w16492_ ;
	wire _w16493_ ;
	wire _w16494_ ;
	wire _w16495_ ;
	wire _w16496_ ;
	wire _w16497_ ;
	wire _w16498_ ;
	wire _w16499_ ;
	wire _w16500_ ;
	wire _w16501_ ;
	wire _w16502_ ;
	wire _w16503_ ;
	wire _w16504_ ;
	wire _w16505_ ;
	wire _w16506_ ;
	wire _w16507_ ;
	wire _w16508_ ;
	wire _w16509_ ;
	wire _w16510_ ;
	wire _w16511_ ;
	wire _w16512_ ;
	wire _w16513_ ;
	wire _w16514_ ;
	wire _w16515_ ;
	wire _w16516_ ;
	wire _w16517_ ;
	wire _w16518_ ;
	wire _w16519_ ;
	wire _w16520_ ;
	wire _w16521_ ;
	wire _w16522_ ;
	wire _w16523_ ;
	wire _w16524_ ;
	wire _w16525_ ;
	wire _w16526_ ;
	wire _w16527_ ;
	wire _w16528_ ;
	wire _w16529_ ;
	wire _w16530_ ;
	wire _w16531_ ;
	wire _w16532_ ;
	wire _w16533_ ;
	wire _w16534_ ;
	wire _w16535_ ;
	wire _w16536_ ;
	wire _w16537_ ;
	wire _w16538_ ;
	wire _w16539_ ;
	wire _w16540_ ;
	wire _w16541_ ;
	wire _w16542_ ;
	wire _w16543_ ;
	wire _w16544_ ;
	wire _w16545_ ;
	wire _w16546_ ;
	wire _w16547_ ;
	wire _w16548_ ;
	wire _w16549_ ;
	wire _w16550_ ;
	wire _w16551_ ;
	wire _w16552_ ;
	wire _w16553_ ;
	wire _w16554_ ;
	wire _w16555_ ;
	wire _w16556_ ;
	wire _w16557_ ;
	wire _w16558_ ;
	wire _w16559_ ;
	wire _w16560_ ;
	wire _w16561_ ;
	wire _w16562_ ;
	wire _w16563_ ;
	wire _w16564_ ;
	wire _w16565_ ;
	wire _w16566_ ;
	wire _w16567_ ;
	wire _w16568_ ;
	wire _w16569_ ;
	wire _w16570_ ;
	wire _w16571_ ;
	wire _w16572_ ;
	wire _w16573_ ;
	wire _w16574_ ;
	wire _w16575_ ;
	wire _w16576_ ;
	wire _w16577_ ;
	wire _w16578_ ;
	wire _w16579_ ;
	wire _w16580_ ;
	wire _w16581_ ;
	wire _w16582_ ;
	wire _w16583_ ;
	wire _w16584_ ;
	wire _w16585_ ;
	wire _w16586_ ;
	wire _w16587_ ;
	wire _w16588_ ;
	wire _w16589_ ;
	wire _w16590_ ;
	wire _w16591_ ;
	wire _w16592_ ;
	wire _w16593_ ;
	wire _w16594_ ;
	wire _w16595_ ;
	wire _w16596_ ;
	wire _w16597_ ;
	wire _w16598_ ;
	wire _w16599_ ;
	wire _w16600_ ;
	wire _w16601_ ;
	wire _w16602_ ;
	wire _w16603_ ;
	wire _w16604_ ;
	wire _w16605_ ;
	wire _w16606_ ;
	wire _w16607_ ;
	wire _w16608_ ;
	wire _w16609_ ;
	wire _w16610_ ;
	wire _w16611_ ;
	wire _w16612_ ;
	wire _w16613_ ;
	wire _w16614_ ;
	wire _w16615_ ;
	wire _w16616_ ;
	wire _w16617_ ;
	wire _w16618_ ;
	wire _w16619_ ;
	wire _w16620_ ;
	wire _w16621_ ;
	wire _w16622_ ;
	wire _w16623_ ;
	wire _w16624_ ;
	wire _w16625_ ;
	wire _w16626_ ;
	wire _w16627_ ;
	wire _w16628_ ;
	wire _w16629_ ;
	wire _w16630_ ;
	wire _w16631_ ;
	wire _w16632_ ;
	wire _w16633_ ;
	wire _w16634_ ;
	wire _w16635_ ;
	wire _w16636_ ;
	wire _w16637_ ;
	wire _w16638_ ;
	wire _w16639_ ;
	wire _w16640_ ;
	wire _w16641_ ;
	wire _w16642_ ;
	wire _w16643_ ;
	wire _w16644_ ;
	wire _w16645_ ;
	wire _w16646_ ;
	wire _w16647_ ;
	wire _w16648_ ;
	wire _w16649_ ;
	wire _w16650_ ;
	wire _w16651_ ;
	wire _w16652_ ;
	wire _w16653_ ;
	wire _w16654_ ;
	wire _w16655_ ;
	wire _w16656_ ;
	wire _w16657_ ;
	wire _w16658_ ;
	wire _w16659_ ;
	wire _w16660_ ;
	wire _w16661_ ;
	wire _w16662_ ;
	wire _w16663_ ;
	wire _w16664_ ;
	wire _w16665_ ;
	wire _w16666_ ;
	wire _w16667_ ;
	wire _w16668_ ;
	wire _w16669_ ;
	wire _w16670_ ;
	wire _w16671_ ;
	wire _w16672_ ;
	wire _w16673_ ;
	wire _w16674_ ;
	wire _w16675_ ;
	wire _w16676_ ;
	wire _w16677_ ;
	wire _w16678_ ;
	wire _w16679_ ;
	wire _w16680_ ;
	wire _w16681_ ;
	wire _w16682_ ;
	wire _w16683_ ;
	wire _w16684_ ;
	wire _w16685_ ;
	wire _w16686_ ;
	wire _w16687_ ;
	wire _w16688_ ;
	wire _w16689_ ;
	wire _w16690_ ;
	wire _w16691_ ;
	wire _w16692_ ;
	wire _w16693_ ;
	wire _w16694_ ;
	wire _w16695_ ;
	wire _w16696_ ;
	wire _w16697_ ;
	wire _w16698_ ;
	wire _w16699_ ;
	wire _w16700_ ;
	wire _w16701_ ;
	wire _w16702_ ;
	wire _w16703_ ;
	wire _w16704_ ;
	wire _w16705_ ;
	wire _w16706_ ;
	wire _w16707_ ;
	wire _w16708_ ;
	wire _w16709_ ;
	wire _w16710_ ;
	wire _w16711_ ;
	wire _w16712_ ;
	wire _w16713_ ;
	wire _w16714_ ;
	wire _w16715_ ;
	wire _w16716_ ;
	wire _w16717_ ;
	wire _w16718_ ;
	wire _w16719_ ;
	wire _w16720_ ;
	wire _w16721_ ;
	wire _w16722_ ;
	wire _w16723_ ;
	wire _w16724_ ;
	wire _w16725_ ;
	wire _w16726_ ;
	wire _w16727_ ;
	wire _w16728_ ;
	wire _w16729_ ;
	wire _w16730_ ;
	wire _w16731_ ;
	wire _w16732_ ;
	wire _w16733_ ;
	wire _w16734_ ;
	wire _w16735_ ;
	wire _w16736_ ;
	wire _w16737_ ;
	wire _w16738_ ;
	wire _w16739_ ;
	wire _w16740_ ;
	wire _w16741_ ;
	wire _w16742_ ;
	wire _w16743_ ;
	wire _w16744_ ;
	wire _w16745_ ;
	wire _w16746_ ;
	wire _w16747_ ;
	wire _w16748_ ;
	wire _w16749_ ;
	wire _w16750_ ;
	wire _w16751_ ;
	wire _w16752_ ;
	wire _w16753_ ;
	wire _w16754_ ;
	wire _w16755_ ;
	wire _w16756_ ;
	wire _w16757_ ;
	wire _w16758_ ;
	wire _w16759_ ;
	wire _w16760_ ;
	wire _w16761_ ;
	wire _w16762_ ;
	wire _w16763_ ;
	wire _w16764_ ;
	wire _w16765_ ;
	wire _w16766_ ;
	wire _w16767_ ;
	wire _w16768_ ;
	wire _w16769_ ;
	wire _w16770_ ;
	wire _w16771_ ;
	wire _w16772_ ;
	wire _w16773_ ;
	wire _w16774_ ;
	wire _w16775_ ;
	wire _w16776_ ;
	wire _w16777_ ;
	wire _w16778_ ;
	wire _w16779_ ;
	wire _w16780_ ;
	wire _w16781_ ;
	wire _w16782_ ;
	wire _w16783_ ;
	wire _w16784_ ;
	wire _w16785_ ;
	wire _w16786_ ;
	wire _w16787_ ;
	wire _w16788_ ;
	wire _w16789_ ;
	wire _w16790_ ;
	wire _w16791_ ;
	wire _w16792_ ;
	wire _w16793_ ;
	wire _w16794_ ;
	wire _w16795_ ;
	wire _w16796_ ;
	wire _w16797_ ;
	wire _w16798_ ;
	wire _w16799_ ;
	wire _w16800_ ;
	wire _w16801_ ;
	wire _w16802_ ;
	wire _w16803_ ;
	wire _w16804_ ;
	wire _w16805_ ;
	wire _w16806_ ;
	wire _w16807_ ;
	wire _w16808_ ;
	wire _w16809_ ;
	wire _w16810_ ;
	wire _w16811_ ;
	wire _w16812_ ;
	wire _w16813_ ;
	wire _w16814_ ;
	wire _w16815_ ;
	wire _w16816_ ;
	wire _w16817_ ;
	wire _w16818_ ;
	wire _w16819_ ;
	wire _w16820_ ;
	wire _w16821_ ;
	wire _w16822_ ;
	wire _w16823_ ;
	wire _w16824_ ;
	wire _w16825_ ;
	wire _w16826_ ;
	wire _w16827_ ;
	wire _w16828_ ;
	wire _w16829_ ;
	wire _w16830_ ;
	wire _w16831_ ;
	wire _w16832_ ;
	wire _w16833_ ;
	wire _w16834_ ;
	wire _w16835_ ;
	wire _w16836_ ;
	wire _w16837_ ;
	wire _w16838_ ;
	wire _w16839_ ;
	wire _w16840_ ;
	wire _w16841_ ;
	wire _w16842_ ;
	wire _w16843_ ;
	wire _w16844_ ;
	wire _w16845_ ;
	wire _w16846_ ;
	wire _w16847_ ;
	wire _w16848_ ;
	wire _w16849_ ;
	wire _w16850_ ;
	wire _w16851_ ;
	wire _w16852_ ;
	wire _w16853_ ;
	wire _w16854_ ;
	wire _w16855_ ;
	wire _w16856_ ;
	wire _w16857_ ;
	wire _w16858_ ;
	wire _w16859_ ;
	wire _w16860_ ;
	wire _w16861_ ;
	wire _w16862_ ;
	wire _w16863_ ;
	wire _w16864_ ;
	wire _w16865_ ;
	wire _w16866_ ;
	wire _w16867_ ;
	wire _w16868_ ;
	wire _w16869_ ;
	wire _w16870_ ;
	wire _w16871_ ;
	wire _w16872_ ;
	wire _w16873_ ;
	wire _w16874_ ;
	wire _w16875_ ;
	wire _w16876_ ;
	wire _w16877_ ;
	wire _w16878_ ;
	wire _w16879_ ;
	wire _w16880_ ;
	wire _w16881_ ;
	wire _w16882_ ;
	wire _w16883_ ;
	wire _w16884_ ;
	wire _w16885_ ;
	wire _w16886_ ;
	wire _w16887_ ;
	wire _w16888_ ;
	wire _w16889_ ;
	wire _w16890_ ;
	wire _w16891_ ;
	wire _w16892_ ;
	wire _w16893_ ;
	wire _w16894_ ;
	wire _w16895_ ;
	wire _w16896_ ;
	wire _w16897_ ;
	wire _w16898_ ;
	wire _w16899_ ;
	wire _w16900_ ;
	wire _w16901_ ;
	wire _w16902_ ;
	wire _w16903_ ;
	wire _w16904_ ;
	wire _w16905_ ;
	wire _w16906_ ;
	wire _w16907_ ;
	wire _w16908_ ;
	wire _w16909_ ;
	wire _w16910_ ;
	wire _w16911_ ;
	wire _w16912_ ;
	wire _w16913_ ;
	wire _w16914_ ;
	wire _w16915_ ;
	wire _w16916_ ;
	wire _w16917_ ;
	wire _w16918_ ;
	wire _w16919_ ;
	wire _w16920_ ;
	wire _w16921_ ;
	wire _w16922_ ;
	wire _w16923_ ;
	wire _w16924_ ;
	wire _w16925_ ;
	wire _w16926_ ;
	wire _w16927_ ;
	wire _w16928_ ;
	wire _w16929_ ;
	wire _w16930_ ;
	wire _w16931_ ;
	wire _w16932_ ;
	wire _w16933_ ;
	wire _w16934_ ;
	wire _w16935_ ;
	wire _w16936_ ;
	wire _w16937_ ;
	wire _w16938_ ;
	wire _w16939_ ;
	wire _w16940_ ;
	wire _w16941_ ;
	wire _w16942_ ;
	wire _w16943_ ;
	wire _w16944_ ;
	wire _w16945_ ;
	wire _w16946_ ;
	wire _w16947_ ;
	wire _w16948_ ;
	wire _w16949_ ;
	wire _w16950_ ;
	wire _w16951_ ;
	wire _w16952_ ;
	wire _w16953_ ;
	wire _w16954_ ;
	wire _w16955_ ;
	wire _w16956_ ;
	wire _w16957_ ;
	wire _w16958_ ;
	wire _w16959_ ;
	wire _w16960_ ;
	wire _w16961_ ;
	wire _w16962_ ;
	wire _w16963_ ;
	wire _w16964_ ;
	wire _w16965_ ;
	wire _w16966_ ;
	wire _w16967_ ;
	wire _w16968_ ;
	wire _w16969_ ;
	wire _w16970_ ;
	wire _w16971_ ;
	wire _w16972_ ;
	wire _w16973_ ;
	wire _w16974_ ;
	wire _w16975_ ;
	wire _w16976_ ;
	wire _w16977_ ;
	wire _w16978_ ;
	wire _w16979_ ;
	wire _w16980_ ;
	wire _w16981_ ;
	wire _w16982_ ;
	wire _w16983_ ;
	wire _w16984_ ;
	wire _w16985_ ;
	wire _w16986_ ;
	wire _w16987_ ;
	wire _w16988_ ;
	wire _w16989_ ;
	wire _w16990_ ;
	wire _w16991_ ;
	wire _w16992_ ;
	wire _w16993_ ;
	wire _w16994_ ;
	wire _w16995_ ;
	wire _w16996_ ;
	wire _w16997_ ;
	wire _w16998_ ;
	wire _w16999_ ;
	wire _w17000_ ;
	wire _w17001_ ;
	wire _w17002_ ;
	wire _w17003_ ;
	wire _w17004_ ;
	wire _w17005_ ;
	wire _w17006_ ;
	wire _w17007_ ;
	wire _w17008_ ;
	wire _w17009_ ;
	wire _w17010_ ;
	wire _w17011_ ;
	wire _w17012_ ;
	wire _w17013_ ;
	wire _w17014_ ;
	wire _w17015_ ;
	wire _w17016_ ;
	wire _w17017_ ;
	wire _w17018_ ;
	wire _w17019_ ;
	wire _w17020_ ;
	wire _w17021_ ;
	wire _w17022_ ;
	wire _w17023_ ;
	wire _w17024_ ;
	wire _w17025_ ;
	wire _w17026_ ;
	wire _w17027_ ;
	wire _w17028_ ;
	wire _w17029_ ;
	wire _w17030_ ;
	wire _w17031_ ;
	wire _w17032_ ;
	wire _w17033_ ;
	wire _w17034_ ;
	wire _w17035_ ;
	wire _w17036_ ;
	wire _w17037_ ;
	wire _w17038_ ;
	wire _w17039_ ;
	wire _w17040_ ;
	wire _w17041_ ;
	wire _w17042_ ;
	wire _w17043_ ;
	wire _w17044_ ;
	wire _w17045_ ;
	wire _w17046_ ;
	wire _w17047_ ;
	wire _w17048_ ;
	wire _w17049_ ;
	wire _w17050_ ;
	wire _w17051_ ;
	wire _w17052_ ;
	wire _w17053_ ;
	wire _w17054_ ;
	wire _w17055_ ;
	wire _w17056_ ;
	wire _w17057_ ;
	wire _w17058_ ;
	wire _w17059_ ;
	wire _w17060_ ;
	wire _w17061_ ;
	wire _w17062_ ;
	wire _w17063_ ;
	wire _w17064_ ;
	wire _w17065_ ;
	wire _w17066_ ;
	wire _w17067_ ;
	wire _w17068_ ;
	wire _w17069_ ;
	wire _w17070_ ;
	wire _w17071_ ;
	wire _w17072_ ;
	wire _w17073_ ;
	wire _w17074_ ;
	wire _w17075_ ;
	wire _w17076_ ;
	wire _w17077_ ;
	wire _w17078_ ;
	wire _w17079_ ;
	wire _w17080_ ;
	wire _w17081_ ;
	wire _w17082_ ;
	wire _w17083_ ;
	wire _w17084_ ;
	wire _w17085_ ;
	wire _w17086_ ;
	wire _w17087_ ;
	wire _w17088_ ;
	wire _w17089_ ;
	wire _w17090_ ;
	wire _w17091_ ;
	wire _w17092_ ;
	wire _w17093_ ;
	wire _w17094_ ;
	wire _w17095_ ;
	wire _w17096_ ;
	wire _w17097_ ;
	wire _w17098_ ;
	wire _w17099_ ;
	wire _w17100_ ;
	wire _w17101_ ;
	wire _w17102_ ;
	wire _w17103_ ;
	wire _w17104_ ;
	wire _w17105_ ;
	wire _w17106_ ;
	wire _w17107_ ;
	wire _w17108_ ;
	wire _w17109_ ;
	wire _w17110_ ;
	wire _w17111_ ;
	wire _w17112_ ;
	wire _w17113_ ;
	wire _w17114_ ;
	wire _w17115_ ;
	wire _w17116_ ;
	wire _w17117_ ;
	wire _w17118_ ;
	wire _w17119_ ;
	wire _w17120_ ;
	wire _w17121_ ;
	wire _w17122_ ;
	wire _w17123_ ;
	wire _w17124_ ;
	wire _w17125_ ;
	wire _w17126_ ;
	wire _w17127_ ;
	wire _w17128_ ;
	wire _w17129_ ;
	wire _w17130_ ;
	wire _w17131_ ;
	wire _w17132_ ;
	wire _w17133_ ;
	wire _w17134_ ;
	wire _w17135_ ;
	wire _w17136_ ;
	wire _w17137_ ;
	wire _w17138_ ;
	wire _w17139_ ;
	wire _w17140_ ;
	wire _w17141_ ;
	wire _w17142_ ;
	wire _w17143_ ;
	wire _w17144_ ;
	wire _w17145_ ;
	wire _w17146_ ;
	wire _w17147_ ;
	wire _w17148_ ;
	wire _w17149_ ;
	wire _w17150_ ;
	wire _w17151_ ;
	wire _w17152_ ;
	wire _w17153_ ;
	wire _w17154_ ;
	wire _w17155_ ;
	wire _w17156_ ;
	wire _w17157_ ;
	wire _w17158_ ;
	wire _w17159_ ;
	wire _w17160_ ;
	wire _w17161_ ;
	wire _w17162_ ;
	wire _w17163_ ;
	wire _w17164_ ;
	wire _w17165_ ;
	wire _w17166_ ;
	wire _w17167_ ;
	wire _w17168_ ;
	wire _w17169_ ;
	wire _w17170_ ;
	wire _w17171_ ;
	wire _w17172_ ;
	wire _w17173_ ;
	wire _w17174_ ;
	wire _w17175_ ;
	wire _w17176_ ;
	wire _w17177_ ;
	wire _w17178_ ;
	wire _w17179_ ;
	wire _w17180_ ;
	wire _w17181_ ;
	wire _w17182_ ;
	wire _w17183_ ;
	wire _w17184_ ;
	wire _w17185_ ;
	wire _w17186_ ;
	wire _w17187_ ;
	wire _w17188_ ;
	wire _w17189_ ;
	wire _w17190_ ;
	wire _w17191_ ;
	wire _w17192_ ;
	wire _w17193_ ;
	wire _w17194_ ;
	wire _w17195_ ;
	wire _w17196_ ;
	wire _w17197_ ;
	wire _w17198_ ;
	wire _w17199_ ;
	wire _w17200_ ;
	wire _w17201_ ;
	wire _w17202_ ;
	wire _w17203_ ;
	wire _w17204_ ;
	wire _w17205_ ;
	wire _w17206_ ;
	wire _w17207_ ;
	wire _w17208_ ;
	wire _w17209_ ;
	wire _w17210_ ;
	wire _w17211_ ;
	wire _w17212_ ;
	wire _w17213_ ;
	wire _w17214_ ;
	wire _w17215_ ;
	wire _w17216_ ;
	wire _w17217_ ;
	wire _w17218_ ;
	wire _w17219_ ;
	wire _w17220_ ;
	wire _w17221_ ;
	wire _w17222_ ;
	wire _w17223_ ;
	wire _w17224_ ;
	wire _w17225_ ;
	wire _w17226_ ;
	wire _w17227_ ;
	wire _w17228_ ;
	wire _w17229_ ;
	wire _w17230_ ;
	wire _w17231_ ;
	wire _w17232_ ;
	wire _w17233_ ;
	wire _w17234_ ;
	wire _w17235_ ;
	wire _w17236_ ;
	wire _w17237_ ;
	wire _w17238_ ;
	wire _w17239_ ;
	wire _w17240_ ;
	wire _w17241_ ;
	wire _w17242_ ;
	wire _w17243_ ;
	wire _w17244_ ;
	wire _w17245_ ;
	wire _w17246_ ;
	wire _w17247_ ;
	wire _w17248_ ;
	wire _w17249_ ;
	wire _w17250_ ;
	wire _w17251_ ;
	wire _w17252_ ;
	wire _w17253_ ;
	wire _w17254_ ;
	wire _w17255_ ;
	wire _w17256_ ;
	wire _w17257_ ;
	wire _w17258_ ;
	wire _w17259_ ;
	wire _w17260_ ;
	wire _w17261_ ;
	wire _w17262_ ;
	wire _w17263_ ;
	wire _w17264_ ;
	wire _w17265_ ;
	wire _w17266_ ;
	wire _w17267_ ;
	wire _w17268_ ;
	wire _w17269_ ;
	wire _w17270_ ;
	wire _w17271_ ;
	wire _w17272_ ;
	wire _w17273_ ;
	wire _w17274_ ;
	wire _w17275_ ;
	wire _w17276_ ;
	wire _w17277_ ;
	wire _w17278_ ;
	wire _w17279_ ;
	wire _w17280_ ;
	wire _w17281_ ;
	wire _w17282_ ;
	wire _w17283_ ;
	wire _w17284_ ;
	wire _w17285_ ;
	wire _w17286_ ;
	wire _w17287_ ;
	wire _w17288_ ;
	wire _w17289_ ;
	wire _w17290_ ;
	wire _w17291_ ;
	wire _w17292_ ;
	wire _w17293_ ;
	wire _w17294_ ;
	wire _w17295_ ;
	wire _w17296_ ;
	wire _w17297_ ;
	wire _w17298_ ;
	wire _w17299_ ;
	wire _w17300_ ;
	wire _w17301_ ;
	wire _w17302_ ;
	wire _w17303_ ;
	wire _w17304_ ;
	wire _w17305_ ;
	wire _w17306_ ;
	wire _w17307_ ;
	wire _w17308_ ;
	wire _w17309_ ;
	wire _w17310_ ;
	wire _w17311_ ;
	wire _w17312_ ;
	wire _w17313_ ;
	wire _w17314_ ;
	wire _w17315_ ;
	wire _w17316_ ;
	wire _w17317_ ;
	wire _w17318_ ;
	wire _w17319_ ;
	wire _w17320_ ;
	wire _w17321_ ;
	wire _w17322_ ;
	wire _w17323_ ;
	wire _w17324_ ;
	wire _w17325_ ;
	wire _w17326_ ;
	wire _w17327_ ;
	wire _w17328_ ;
	wire _w17329_ ;
	wire _w17330_ ;
	wire _w17331_ ;
	wire _w17332_ ;
	wire _w17333_ ;
	wire _w17334_ ;
	wire _w17335_ ;
	wire _w17336_ ;
	wire _w17337_ ;
	wire _w17338_ ;
	wire _w17339_ ;
	wire _w17340_ ;
	wire _w17341_ ;
	wire _w17342_ ;
	wire _w17343_ ;
	wire _w17344_ ;
	wire _w17345_ ;
	wire _w17346_ ;
	wire _w17347_ ;
	wire _w17348_ ;
	wire _w17349_ ;
	wire _w17350_ ;
	wire _w17351_ ;
	wire _w17352_ ;
	wire _w17353_ ;
	wire _w17354_ ;
	wire _w17355_ ;
	wire _w17356_ ;
	wire _w17357_ ;
	wire _w17358_ ;
	wire _w17359_ ;
	wire _w17360_ ;
	wire _w17361_ ;
	wire _w17362_ ;
	wire _w17363_ ;
	wire _w17364_ ;
	wire _w17365_ ;
	wire _w17366_ ;
	wire _w17367_ ;
	wire _w17368_ ;
	wire _w17369_ ;
	wire _w17370_ ;
	wire _w17371_ ;
	wire _w17372_ ;
	wire _w17373_ ;
	wire _w17374_ ;
	wire _w17375_ ;
	wire _w17376_ ;
	wire _w17377_ ;
	wire _w17378_ ;
	wire _w17379_ ;
	wire _w17380_ ;
	wire _w17381_ ;
	wire _w17382_ ;
	wire _w17383_ ;
	wire _w17384_ ;
	wire _w17385_ ;
	wire _w17386_ ;
	wire _w17387_ ;
	wire _w17388_ ;
	wire _w17389_ ;
	wire _w17390_ ;
	wire _w17391_ ;
	wire _w17392_ ;
	wire _w17393_ ;
	wire _w17394_ ;
	wire _w17395_ ;
	wire _w17396_ ;
	wire _w17397_ ;
	wire _w17398_ ;
	wire _w17399_ ;
	wire _w17400_ ;
	wire _w17401_ ;
	wire _w17402_ ;
	wire _w17403_ ;
	wire _w17404_ ;
	wire _w17405_ ;
	wire _w17406_ ;
	wire _w17407_ ;
	wire _w17408_ ;
	wire _w17409_ ;
	wire _w17410_ ;
	wire _w17411_ ;
	wire _w17412_ ;
	wire _w17413_ ;
	wire _w17414_ ;
	wire _w17415_ ;
	wire _w17416_ ;
	wire _w17417_ ;
	wire _w17418_ ;
	wire _w17419_ ;
	wire _w17420_ ;
	wire _w17421_ ;
	wire _w17422_ ;
	wire _w17423_ ;
	wire _w17424_ ;
	wire _w17425_ ;
	wire _w17426_ ;
	wire _w17427_ ;
	wire _w17428_ ;
	wire _w17429_ ;
	wire _w17430_ ;
	wire _w17431_ ;
	wire _w17432_ ;
	wire _w17433_ ;
	wire _w17434_ ;
	wire _w17435_ ;
	wire _w17436_ ;
	wire _w17437_ ;
	wire _w17438_ ;
	wire _w17439_ ;
	wire _w17440_ ;
	wire _w17441_ ;
	wire _w17442_ ;
	wire _w17443_ ;
	wire _w17444_ ;
	wire _w17445_ ;
	wire _w17446_ ;
	wire _w17447_ ;
	wire _w17448_ ;
	wire _w17449_ ;
	wire _w17450_ ;
	wire _w17451_ ;
	wire _w17452_ ;
	wire _w17453_ ;
	wire _w17454_ ;
	wire _w17455_ ;
	wire _w17456_ ;
	wire _w17457_ ;
	wire _w17458_ ;
	wire _w17459_ ;
	wire _w17460_ ;
	wire _w17461_ ;
	wire _w17462_ ;
	wire _w17463_ ;
	wire _w17464_ ;
	wire _w17465_ ;
	wire _w17466_ ;
	wire _w17467_ ;
	wire _w17468_ ;
	wire _w17469_ ;
	wire _w17470_ ;
	wire _w17471_ ;
	wire _w17472_ ;
	wire _w17473_ ;
	wire _w17474_ ;
	wire _w17475_ ;
	wire _w17476_ ;
	wire _w17477_ ;
	wire _w17478_ ;
	wire _w17479_ ;
	wire _w17480_ ;
	wire _w17481_ ;
	wire _w17482_ ;
	wire _w17483_ ;
	wire _w17484_ ;
	wire _w17485_ ;
	wire _w17486_ ;
	wire _w17487_ ;
	wire _w17488_ ;
	wire _w17489_ ;
	wire _w17490_ ;
	wire _w17491_ ;
	wire _w17492_ ;
	wire _w17493_ ;
	wire _w17494_ ;
	wire _w17495_ ;
	wire _w17496_ ;
	wire _w17497_ ;
	wire _w17498_ ;
	wire _w17499_ ;
	wire _w17500_ ;
	wire _w17501_ ;
	wire _w17502_ ;
	wire _w17503_ ;
	wire _w17504_ ;
	wire _w17505_ ;
	wire _w17506_ ;
	wire _w17507_ ;
	wire _w17508_ ;
	wire _w17509_ ;
	wire _w17510_ ;
	wire _w17511_ ;
	wire _w17512_ ;
	wire _w17513_ ;
	wire _w17514_ ;
	wire _w17515_ ;
	wire _w17516_ ;
	wire _w17517_ ;
	wire _w17518_ ;
	wire _w17519_ ;
	wire _w17520_ ;
	wire _w17521_ ;
	wire _w17522_ ;
	wire _w17523_ ;
	wire _w17524_ ;
	wire _w17525_ ;
	wire _w17526_ ;
	wire _w17527_ ;
	wire _w17528_ ;
	wire _w17529_ ;
	wire _w17530_ ;
	wire _w17531_ ;
	wire _w17532_ ;
	wire _w17533_ ;
	wire _w17534_ ;
	wire _w17535_ ;
	wire _w17536_ ;
	wire _w17537_ ;
	wire _w17538_ ;
	wire _w17539_ ;
	wire _w17540_ ;
	wire _w17541_ ;
	wire _w17542_ ;
	wire _w17543_ ;
	wire _w17544_ ;
	wire _w17545_ ;
	wire _w17546_ ;
	wire _w17547_ ;
	wire _w17548_ ;
	wire _w17549_ ;
	wire _w17550_ ;
	wire _w17551_ ;
	wire _w17552_ ;
	wire _w17553_ ;
	wire _w17554_ ;
	wire _w17555_ ;
	wire _w17556_ ;
	wire _w17557_ ;
	wire _w17558_ ;
	wire _w17559_ ;
	wire _w17560_ ;
	wire _w17561_ ;
	wire _w17562_ ;
	wire _w17563_ ;
	wire _w17564_ ;
	wire _w17565_ ;
	wire _w17566_ ;
	wire _w17567_ ;
	wire _w17568_ ;
	wire _w17569_ ;
	wire _w17570_ ;
	wire _w17571_ ;
	wire _w17572_ ;
	wire _w17573_ ;
	wire _w17574_ ;
	wire _w17575_ ;
	wire _w17576_ ;
	wire _w17577_ ;
	wire _w17578_ ;
	wire _w17579_ ;
	wire _w17580_ ;
	wire _w17581_ ;
	wire _w17582_ ;
	wire _w17583_ ;
	wire _w17584_ ;
	wire _w17585_ ;
	wire _w17586_ ;
	wire _w17587_ ;
	wire _w17588_ ;
	wire _w17589_ ;
	wire _w17590_ ;
	wire _w17591_ ;
	wire _w17592_ ;
	wire _w17593_ ;
	wire _w17594_ ;
	wire _w17595_ ;
	wire _w17596_ ;
	wire _w17597_ ;
	wire _w17598_ ;
	wire _w17599_ ;
	wire _w17600_ ;
	wire _w17601_ ;
	wire _w17602_ ;
	wire _w17603_ ;
	wire _w17604_ ;
	wire _w17605_ ;
	wire _w17606_ ;
	wire _w17607_ ;
	wire _w17608_ ;
	wire _w17609_ ;
	wire _w17610_ ;
	wire _w17611_ ;
	wire _w17612_ ;
	wire _w17613_ ;
	wire _w17614_ ;
	wire _w17615_ ;
	wire _w17616_ ;
	wire _w17617_ ;
	wire _w17618_ ;
	wire _w17619_ ;
	wire _w17620_ ;
	wire _w17621_ ;
	wire _w17622_ ;
	wire _w17623_ ;
	wire _w17624_ ;
	wire _w17625_ ;
	wire _w17626_ ;
	wire _w17627_ ;
	wire _w17628_ ;
	wire _w17629_ ;
	wire _w17630_ ;
	wire _w17631_ ;
	wire _w17632_ ;
	wire _w17633_ ;
	wire _w17634_ ;
	wire _w17635_ ;
	wire _w17636_ ;
	wire _w17637_ ;
	wire _w17638_ ;
	wire _w17639_ ;
	wire _w17640_ ;
	wire _w17641_ ;
	wire _w17642_ ;
	wire _w17643_ ;
	wire _w17644_ ;
	wire _w17645_ ;
	wire _w17646_ ;
	wire _w17647_ ;
	wire _w17648_ ;
	wire _w17649_ ;
	wire _w17650_ ;
	wire _w17651_ ;
	wire _w17652_ ;
	wire _w17653_ ;
	wire _w17654_ ;
	wire _w17655_ ;
	wire _w17656_ ;
	wire _w17657_ ;
	wire _w17658_ ;
	wire _w17659_ ;
	wire _w17660_ ;
	wire _w17661_ ;
	wire _w17662_ ;
	wire _w17663_ ;
	wire _w17664_ ;
	wire _w17665_ ;
	wire _w17666_ ;
	wire _w17667_ ;
	wire _w17668_ ;
	wire _w17669_ ;
	wire _w17670_ ;
	wire _w17671_ ;
	wire _w17672_ ;
	wire _w17673_ ;
	wire _w17674_ ;
	wire _w17675_ ;
	wire _w17676_ ;
	wire _w17677_ ;
	wire _w17678_ ;
	wire _w17679_ ;
	wire _w17680_ ;
	wire _w17681_ ;
	wire _w17682_ ;
	wire _w17683_ ;
	wire _w17684_ ;
	wire _w17685_ ;
	wire _w17686_ ;
	wire _w17687_ ;
	wire _w17688_ ;
	wire _w17689_ ;
	wire _w17690_ ;
	wire _w17691_ ;
	wire _w17692_ ;
	wire _w17693_ ;
	wire _w17694_ ;
	wire _w17695_ ;
	wire _w17696_ ;
	wire _w17697_ ;
	wire _w17698_ ;
	wire _w17699_ ;
	wire _w17700_ ;
	wire _w17701_ ;
	wire _w17702_ ;
	wire _w17703_ ;
	wire _w17704_ ;
	wire _w17705_ ;
	wire _w17706_ ;
	wire _w17707_ ;
	wire _w17708_ ;
	wire _w17709_ ;
	wire _w17710_ ;
	wire _w17711_ ;
	wire _w17712_ ;
	wire _w17713_ ;
	wire _w17714_ ;
	wire _w17715_ ;
	wire _w17716_ ;
	wire _w17717_ ;
	wire _w17718_ ;
	wire _w17719_ ;
	wire _w17720_ ;
	wire _w17721_ ;
	wire _w17722_ ;
	wire _w17723_ ;
	wire _w17724_ ;
	wire _w17725_ ;
	wire _w17726_ ;
	wire _w17727_ ;
	wire _w17728_ ;
	wire _w17729_ ;
	wire _w17730_ ;
	wire _w17731_ ;
	wire _w17732_ ;
	wire _w17733_ ;
	wire _w17734_ ;
	wire _w17735_ ;
	wire _w17736_ ;
	wire _w17737_ ;
	wire _w17738_ ;
	wire _w17739_ ;
	wire _w17740_ ;
	wire _w17741_ ;
	wire _w17742_ ;
	wire _w17743_ ;
	wire _w17744_ ;
	wire _w17745_ ;
	wire _w17746_ ;
	wire _w17747_ ;
	wire _w17748_ ;
	wire _w17749_ ;
	wire _w17750_ ;
	wire _w17751_ ;
	wire _w17752_ ;
	wire _w17753_ ;
	wire _w17754_ ;
	wire _w17755_ ;
	wire _w17756_ ;
	wire _w17757_ ;
	wire _w17758_ ;
	wire _w17759_ ;
	wire _w17760_ ;
	wire _w17761_ ;
	wire _w17762_ ;
	wire _w17763_ ;
	wire _w17764_ ;
	wire _w17765_ ;
	wire _w17766_ ;
	wire _w17767_ ;
	wire _w17768_ ;
	wire _w17769_ ;
	wire _w17770_ ;
	wire _w17771_ ;
	wire _w17772_ ;
	wire _w17773_ ;
	wire _w17774_ ;
	wire _w17775_ ;
	wire _w17776_ ;
	wire _w17777_ ;
	wire _w17778_ ;
	wire _w17779_ ;
	wire _w17780_ ;
	wire _w17781_ ;
	wire _w17782_ ;
	wire _w17783_ ;
	wire _w17784_ ;
	wire _w17785_ ;
	wire _w17786_ ;
	wire _w17787_ ;
	wire _w17788_ ;
	wire _w17789_ ;
	wire _w17790_ ;
	wire _w17791_ ;
	wire _w17792_ ;
	wire _w17793_ ;
	wire _w17794_ ;
	wire _w17795_ ;
	wire _w17796_ ;
	wire _w17797_ ;
	wire _w17798_ ;
	wire _w17799_ ;
	wire _w17800_ ;
	wire _w17801_ ;
	wire _w17802_ ;
	wire _w17803_ ;
	wire _w17804_ ;
	wire _w17805_ ;
	wire _w17806_ ;
	wire _w17807_ ;
	wire _w17808_ ;
	wire _w17809_ ;
	wire _w17810_ ;
	wire _w17811_ ;
	wire _w17812_ ;
	wire _w17813_ ;
	wire _w17814_ ;
	wire _w17815_ ;
	wire _w17816_ ;
	wire _w17817_ ;
	wire _w17818_ ;
	wire _w17819_ ;
	wire _w17820_ ;
	wire _w17821_ ;
	wire _w17822_ ;
	wire _w17823_ ;
	wire _w17824_ ;
	wire _w17825_ ;
	wire _w17826_ ;
	wire _w17827_ ;
	wire _w17828_ ;
	wire _w17829_ ;
	wire _w17830_ ;
	wire _w17831_ ;
	wire _w17832_ ;
	wire _w17833_ ;
	wire _w17834_ ;
	wire _w17835_ ;
	wire _w17836_ ;
	wire _w17837_ ;
	wire _w17838_ ;
	wire _w17839_ ;
	wire _w17840_ ;
	wire _w17841_ ;
	wire _w17842_ ;
	wire _w17843_ ;
	wire _w17844_ ;
	wire _w17845_ ;
	wire _w17846_ ;
	wire _w17847_ ;
	wire _w17848_ ;
	wire _w17849_ ;
	wire _w17850_ ;
	wire _w17851_ ;
	wire _w17852_ ;
	wire _w17853_ ;
	wire _w17854_ ;
	wire _w17855_ ;
	wire _w17856_ ;
	wire _w17857_ ;
	wire _w17858_ ;
	wire _w17859_ ;
	wire _w17860_ ;
	wire _w17861_ ;
	wire _w17862_ ;
	wire _w17863_ ;
	wire _w17864_ ;
	wire _w17865_ ;
	wire _w17866_ ;
	wire _w17867_ ;
	wire _w17868_ ;
	wire _w17869_ ;
	wire _w17870_ ;
	wire _w17871_ ;
	wire _w17872_ ;
	wire _w17873_ ;
	wire _w17874_ ;
	wire _w17875_ ;
	wire _w17876_ ;
	wire _w17877_ ;
	wire _w17878_ ;
	wire _w17879_ ;
	wire _w17880_ ;
	wire _w17881_ ;
	wire _w17882_ ;
	wire _w17883_ ;
	wire _w17884_ ;
	wire _w17885_ ;
	wire _w17886_ ;
	wire _w17887_ ;
	wire _w17888_ ;
	wire _w17889_ ;
	wire _w17890_ ;
	wire _w17891_ ;
	wire _w17892_ ;
	wire _w17893_ ;
	wire _w17894_ ;
	wire _w17895_ ;
	wire _w17896_ ;
	wire _w17897_ ;
	wire _w17898_ ;
	wire _w17899_ ;
	wire _w17900_ ;
	wire _w17901_ ;
	wire _w17902_ ;
	wire _w17903_ ;
	wire _w17904_ ;
	wire _w17905_ ;
	wire _w17906_ ;
	wire _w17907_ ;
	wire _w17908_ ;
	wire _w17909_ ;
	wire _w17910_ ;
	wire _w17911_ ;
	wire _w17912_ ;
	wire _w17913_ ;
	wire _w17914_ ;
	wire _w17915_ ;
	wire _w17916_ ;
	wire _w17917_ ;
	wire _w17918_ ;
	wire _w17919_ ;
	wire _w17920_ ;
	wire _w17921_ ;
	wire _w17922_ ;
	wire _w17923_ ;
	wire _w17924_ ;
	wire _w17925_ ;
	wire _w17926_ ;
	wire _w17927_ ;
	wire _w17928_ ;
	wire _w17929_ ;
	wire _w17930_ ;
	wire _w17931_ ;
	wire _w17932_ ;
	wire _w17933_ ;
	wire _w17934_ ;
	wire _w17935_ ;
	wire _w17936_ ;
	wire _w17937_ ;
	wire _w17938_ ;
	wire _w17939_ ;
	wire _w17940_ ;
	wire _w17941_ ;
	wire _w17942_ ;
	wire _w17943_ ;
	wire _w17944_ ;
	wire _w17945_ ;
	wire _w17946_ ;
	wire _w17947_ ;
	wire _w17948_ ;
	wire _w17949_ ;
	wire _w17950_ ;
	wire _w17951_ ;
	wire _w17952_ ;
	wire _w17953_ ;
	wire _w17954_ ;
	wire _w17955_ ;
	wire _w17956_ ;
	wire _w17957_ ;
	wire _w17958_ ;
	wire _w17959_ ;
	wire _w17960_ ;
	wire _w17961_ ;
	wire _w17962_ ;
	wire _w17963_ ;
	wire _w17964_ ;
	wire _w17965_ ;
	wire _w17966_ ;
	wire _w17967_ ;
	wire _w17968_ ;
	wire _w17969_ ;
	wire _w17970_ ;
	wire _w17971_ ;
	wire _w17972_ ;
	wire _w17973_ ;
	wire _w17974_ ;
	wire _w17975_ ;
	wire _w17976_ ;
	wire _w17977_ ;
	wire _w17978_ ;
	wire _w17979_ ;
	wire _w17980_ ;
	wire _w17981_ ;
	wire _w17982_ ;
	wire _w17983_ ;
	wire _w17984_ ;
	wire _w17985_ ;
	wire _w17986_ ;
	wire _w17987_ ;
	wire _w17988_ ;
	wire _w17989_ ;
	wire _w17990_ ;
	wire _w17991_ ;
	wire _w17992_ ;
	wire _w17993_ ;
	wire _w17994_ ;
	wire _w17995_ ;
	wire _w17996_ ;
	wire _w17997_ ;
	wire _w17998_ ;
	wire _w17999_ ;
	wire _w18000_ ;
	wire _w18001_ ;
	wire _w18002_ ;
	wire _w18003_ ;
	wire _w18004_ ;
	wire _w18005_ ;
	wire _w18006_ ;
	wire _w18007_ ;
	wire _w18008_ ;
	wire _w18009_ ;
	wire _w18010_ ;
	wire _w18011_ ;
	wire _w18012_ ;
	wire _w18013_ ;
	wire _w18014_ ;
	wire _w18015_ ;
	wire _w18016_ ;
	wire _w18017_ ;
	wire _w18018_ ;
	wire _w18019_ ;
	wire _w18020_ ;
	wire _w18021_ ;
	wire _w18022_ ;
	wire _w18023_ ;
	wire _w18024_ ;
	wire _w18025_ ;
	wire _w18026_ ;
	wire _w18027_ ;
	wire _w18028_ ;
	wire _w18029_ ;
	wire _w18030_ ;
	wire _w18031_ ;
	wire _w18032_ ;
	wire _w18033_ ;
	wire _w18034_ ;
	wire _w18035_ ;
	wire _w18036_ ;
	wire _w18037_ ;
	wire _w18038_ ;
	wire _w18039_ ;
	wire _w18040_ ;
	wire _w18041_ ;
	wire _w18042_ ;
	wire _w18043_ ;
	wire _w18044_ ;
	wire _w18045_ ;
	wire _w18046_ ;
	wire _w18047_ ;
	wire _w18048_ ;
	wire _w18049_ ;
	wire _w18050_ ;
	wire _w18051_ ;
	wire _w18052_ ;
	wire _w18053_ ;
	wire _w18054_ ;
	wire _w18055_ ;
	wire _w18056_ ;
	wire _w18057_ ;
	wire _w18058_ ;
	wire _w18059_ ;
	wire _w18060_ ;
	wire _w18061_ ;
	wire _w18062_ ;
	wire _w18063_ ;
	wire _w18064_ ;
	wire _w18065_ ;
	wire _w18066_ ;
	wire _w18067_ ;
	wire _w18068_ ;
	wire _w18069_ ;
	wire _w18070_ ;
	wire _w18071_ ;
	wire _w18072_ ;
	wire _w18073_ ;
	wire _w18074_ ;
	wire _w18075_ ;
	wire _w18076_ ;
	wire _w18077_ ;
	wire _w18078_ ;
	wire _w18079_ ;
	wire _w18080_ ;
	wire _w18081_ ;
	wire _w18082_ ;
	wire _w18083_ ;
	wire _w18084_ ;
	wire _w18085_ ;
	wire _w18086_ ;
	wire _w18087_ ;
	wire _w18088_ ;
	wire _w18089_ ;
	wire _w18090_ ;
	wire _w18091_ ;
	wire _w18092_ ;
	wire _w18093_ ;
	wire _w18094_ ;
	wire _w18095_ ;
	wire _w18096_ ;
	wire _w18097_ ;
	wire _w18098_ ;
	wire _w18099_ ;
	wire _w18100_ ;
	wire _w18101_ ;
	wire _w18102_ ;
	wire _w18103_ ;
	wire _w18104_ ;
	wire _w18105_ ;
	wire _w18106_ ;
	wire _w18107_ ;
	wire _w18108_ ;
	wire _w18109_ ;
	wire _w18110_ ;
	wire _w18111_ ;
	wire _w18112_ ;
	wire _w18113_ ;
	wire _w18114_ ;
	wire _w18115_ ;
	wire _w18116_ ;
	wire _w18117_ ;
	wire _w18118_ ;
	wire _w18119_ ;
	wire _w18120_ ;
	wire _w18121_ ;
	wire _w18122_ ;
	wire _w18123_ ;
	wire _w18124_ ;
	wire _w18125_ ;
	wire _w18126_ ;
	wire _w18127_ ;
	wire _w18128_ ;
	wire _w18129_ ;
	wire _w18130_ ;
	wire _w18131_ ;
	wire _w18132_ ;
	wire _w18133_ ;
	wire _w18134_ ;
	wire _w18135_ ;
	wire _w18136_ ;
	wire _w18137_ ;
	wire _w18138_ ;
	wire _w18139_ ;
	wire _w18140_ ;
	wire _w18141_ ;
	wire _w18142_ ;
	wire _w18143_ ;
	wire _w18144_ ;
	wire _w18145_ ;
	wire _w18146_ ;
	wire _w18147_ ;
	wire _w18148_ ;
	wire _w18149_ ;
	wire _w18150_ ;
	wire _w18151_ ;
	wire _w18152_ ;
	wire _w18153_ ;
	wire _w18154_ ;
	wire _w18155_ ;
	wire _w18156_ ;
	wire _w18157_ ;
	wire _w18158_ ;
	wire _w18159_ ;
	wire _w18160_ ;
	wire _w18161_ ;
	wire _w18162_ ;
	wire _w18163_ ;
	wire _w18164_ ;
	wire _w18165_ ;
	wire _w18166_ ;
	wire _w18167_ ;
	wire _w18168_ ;
	wire _w18169_ ;
	wire _w18170_ ;
	wire _w18171_ ;
	wire _w18172_ ;
	wire _w18173_ ;
	wire _w18174_ ;
	wire _w18175_ ;
	wire _w18176_ ;
	wire _w18177_ ;
	wire _w18178_ ;
	wire _w18179_ ;
	wire _w18180_ ;
	wire _w18181_ ;
	wire _w18182_ ;
	wire _w18183_ ;
	wire _w18184_ ;
	wire _w18185_ ;
	wire _w18186_ ;
	wire _w18187_ ;
	wire _w18188_ ;
	wire _w18189_ ;
	wire _w18190_ ;
	wire _w18191_ ;
	wire _w18192_ ;
	wire _w18193_ ;
	wire _w18194_ ;
	wire _w18195_ ;
	wire _w18196_ ;
	wire _w18197_ ;
	wire _w18198_ ;
	wire _w18199_ ;
	wire _w18200_ ;
	wire _w18201_ ;
	wire _w18202_ ;
	wire _w18203_ ;
	wire _w18204_ ;
	wire _w18205_ ;
	wire _w18206_ ;
	wire _w18207_ ;
	wire _w18208_ ;
	wire _w18209_ ;
	wire _w18210_ ;
	wire _w18211_ ;
	wire _w18212_ ;
	wire _w18213_ ;
	wire _w18214_ ;
	wire _w18215_ ;
	wire _w18216_ ;
	wire _w18217_ ;
	wire _w18218_ ;
	wire _w18219_ ;
	wire _w18220_ ;
	wire _w18221_ ;
	wire _w18222_ ;
	wire _w18223_ ;
	wire _w18224_ ;
	wire _w18225_ ;
	wire _w18226_ ;
	wire _w18227_ ;
	wire _w18228_ ;
	wire _w18229_ ;
	wire _w18230_ ;
	wire _w18231_ ;
	wire _w18232_ ;
	wire _w18233_ ;
	wire _w18234_ ;
	wire _w18235_ ;
	wire _w18236_ ;
	wire _w18237_ ;
	wire _w18238_ ;
	wire _w18239_ ;
	wire _w18240_ ;
	wire _w18241_ ;
	wire _w18242_ ;
	wire _w18243_ ;
	wire _w18244_ ;
	wire _w18245_ ;
	wire _w18246_ ;
	wire _w18247_ ;
	wire _w18248_ ;
	wire _w18249_ ;
	wire _w18250_ ;
	wire _w18251_ ;
	wire _w18252_ ;
	wire _w18253_ ;
	wire _w18254_ ;
	wire _w18255_ ;
	wire _w18256_ ;
	wire _w18257_ ;
	wire _w18258_ ;
	wire _w18259_ ;
	wire _w18260_ ;
	wire _w18261_ ;
	wire _w18262_ ;
	wire _w18263_ ;
	wire _w18264_ ;
	wire _w18265_ ;
	wire _w18266_ ;
	wire _w18267_ ;
	wire _w18268_ ;
	wire _w18269_ ;
	wire _w18270_ ;
	wire _w18271_ ;
	wire _w18272_ ;
	wire _w18273_ ;
	wire _w18274_ ;
	wire _w18275_ ;
	wire _w18276_ ;
	wire _w18277_ ;
	wire _w18278_ ;
	wire _w18279_ ;
	wire _w18280_ ;
	wire _w18281_ ;
	wire _w18282_ ;
	wire _w18283_ ;
	wire _w18284_ ;
	wire _w18285_ ;
	wire _w18286_ ;
	wire _w18287_ ;
	wire _w18288_ ;
	wire _w18289_ ;
	wire _w18290_ ;
	wire _w18291_ ;
	wire _w18292_ ;
	wire _w18293_ ;
	wire _w18294_ ;
	wire _w18295_ ;
	wire _w18296_ ;
	wire _w18297_ ;
	wire _w18298_ ;
	wire _w18299_ ;
	wire _w18300_ ;
	wire _w18301_ ;
	wire _w18302_ ;
	wire _w18303_ ;
	wire _w18304_ ;
	wire _w18305_ ;
	wire _w18306_ ;
	wire _w18307_ ;
	wire _w18308_ ;
	wire _w18309_ ;
	wire _w18310_ ;
	wire _w18311_ ;
	wire _w18312_ ;
	wire _w18313_ ;
	wire _w18314_ ;
	wire _w18315_ ;
	wire _w18316_ ;
	wire _w18317_ ;
	wire _w18318_ ;
	wire _w18319_ ;
	wire _w18320_ ;
	wire _w18321_ ;
	wire _w18322_ ;
	wire _w18323_ ;
	wire _w18324_ ;
	wire _w18325_ ;
	wire _w18326_ ;
	wire _w18327_ ;
	wire _w18328_ ;
	wire _w18329_ ;
	wire _w18330_ ;
	wire _w18331_ ;
	wire _w18332_ ;
	wire _w18333_ ;
	wire _w18334_ ;
	wire _w18335_ ;
	wire _w18336_ ;
	wire _w18337_ ;
	wire _w18338_ ;
	wire _w18339_ ;
	wire _w18340_ ;
	wire _w18341_ ;
	wire _w18342_ ;
	wire _w18343_ ;
	wire _w18344_ ;
	wire _w18345_ ;
	wire _w18346_ ;
	wire _w18347_ ;
	wire _w18348_ ;
	wire _w18349_ ;
	wire _w18350_ ;
	wire _w18351_ ;
	wire _w18352_ ;
	wire _w18353_ ;
	wire _w18354_ ;
	wire _w18355_ ;
	wire _w18356_ ;
	wire _w18357_ ;
	wire _w18358_ ;
	wire _w18359_ ;
	wire _w18360_ ;
	wire _w18361_ ;
	wire _w18362_ ;
	wire _w18363_ ;
	wire _w18364_ ;
	wire _w18365_ ;
	wire _w18366_ ;
	wire _w18367_ ;
	wire _w18368_ ;
	wire _w18369_ ;
	wire _w18370_ ;
	wire _w18371_ ;
	wire _w18372_ ;
	wire _w18373_ ;
	wire _w18374_ ;
	wire _w18375_ ;
	wire _w18376_ ;
	wire _w18377_ ;
	wire _w18378_ ;
	wire _w18379_ ;
	wire _w18380_ ;
	wire _w18381_ ;
	wire _w18382_ ;
	wire _w18383_ ;
	wire _w18384_ ;
	wire _w18385_ ;
	wire _w18386_ ;
	wire _w18387_ ;
	wire _w18388_ ;
	wire _w18389_ ;
	wire _w18390_ ;
	wire _w18391_ ;
	wire _w18392_ ;
	wire _w18393_ ;
	wire _w18394_ ;
	wire _w18395_ ;
	wire _w18396_ ;
	wire _w18397_ ;
	wire _w18398_ ;
	wire _w18399_ ;
	wire _w18400_ ;
	wire _w18401_ ;
	wire _w18402_ ;
	wire _w18403_ ;
	wire _w18404_ ;
	wire _w18405_ ;
	wire _w18406_ ;
	wire _w18407_ ;
	wire _w18408_ ;
	wire _w18409_ ;
	wire _w18410_ ;
	wire _w18411_ ;
	wire _w18412_ ;
	wire _w18413_ ;
	wire _w18414_ ;
	wire _w18415_ ;
	wire _w18416_ ;
	wire _w18417_ ;
	wire _w18418_ ;
	wire _w18419_ ;
	wire _w18420_ ;
	wire _w18421_ ;
	wire _w18422_ ;
	wire _w18423_ ;
	wire _w18424_ ;
	wire _w18425_ ;
	wire _w18426_ ;
	wire _w18427_ ;
	wire _w18428_ ;
	wire _w18429_ ;
	wire _w18430_ ;
	wire _w18431_ ;
	wire _w18432_ ;
	wire _w18433_ ;
	wire _w18434_ ;
	wire _w18435_ ;
	wire _w18436_ ;
	wire _w18437_ ;
	wire _w18438_ ;
	wire _w18439_ ;
	wire _w18440_ ;
	wire _w18441_ ;
	wire _w18442_ ;
	wire _w18443_ ;
	wire _w18444_ ;
	wire _w18445_ ;
	wire _w18446_ ;
	wire _w18447_ ;
	wire _w18448_ ;
	wire _w18449_ ;
	wire _w18450_ ;
	wire _w18451_ ;
	wire _w18452_ ;
	wire _w18453_ ;
	wire _w18454_ ;
	wire _w18455_ ;
	wire _w18456_ ;
	wire _w18457_ ;
	wire _w18458_ ;
	wire _w18459_ ;
	wire _w18460_ ;
	wire _w18461_ ;
	wire _w18462_ ;
	wire _w18463_ ;
	wire _w18464_ ;
	wire _w18465_ ;
	wire _w18466_ ;
	wire _w18467_ ;
	wire _w18468_ ;
	wire _w18469_ ;
	wire _w18470_ ;
	wire _w18471_ ;
	wire _w18472_ ;
	wire _w18473_ ;
	wire _w18474_ ;
	wire _w18475_ ;
	wire _w18476_ ;
	wire _w18477_ ;
	wire _w18478_ ;
	wire _w18479_ ;
	wire _w18480_ ;
	wire _w18481_ ;
	wire _w18482_ ;
	wire _w18483_ ;
	wire _w18484_ ;
	wire _w18485_ ;
	wire _w18486_ ;
	wire _w18487_ ;
	wire _w18488_ ;
	wire _w18489_ ;
	wire _w18490_ ;
	wire _w18491_ ;
	wire _w18492_ ;
	wire _w18493_ ;
	wire _w18494_ ;
	wire _w18495_ ;
	wire _w18496_ ;
	wire _w18497_ ;
	wire _w18498_ ;
	wire _w18499_ ;
	wire _w18500_ ;
	wire _w18501_ ;
	wire _w18502_ ;
	wire _w18503_ ;
	wire _w18504_ ;
	wire _w18505_ ;
	wire _w18506_ ;
	wire _w18507_ ;
	wire _w18508_ ;
	wire _w18509_ ;
	wire _w18510_ ;
	wire _w18511_ ;
	wire _w18512_ ;
	wire _w18513_ ;
	wire _w18514_ ;
	wire _w18515_ ;
	wire _w18516_ ;
	wire _w18517_ ;
	wire _w18518_ ;
	wire _w18519_ ;
	wire _w18520_ ;
	wire _w18521_ ;
	wire _w18522_ ;
	wire _w18523_ ;
	wire _w18524_ ;
	wire _w18525_ ;
	wire _w18526_ ;
	wire _w18527_ ;
	wire _w18528_ ;
	wire _w18529_ ;
	wire _w18530_ ;
	wire _w18531_ ;
	wire _w18532_ ;
	wire _w18533_ ;
	wire _w18534_ ;
	wire _w18535_ ;
	wire _w18536_ ;
	wire _w18537_ ;
	wire _w18538_ ;
	wire _w18539_ ;
	wire _w18540_ ;
	wire _w18541_ ;
	wire _w18542_ ;
	wire _w18543_ ;
	wire _w18544_ ;
	wire _w18545_ ;
	wire _w18546_ ;
	wire _w18547_ ;
	wire _w18548_ ;
	wire _w18549_ ;
	wire _w18550_ ;
	wire _w18551_ ;
	wire _w18552_ ;
	wire _w18553_ ;
	wire _w18554_ ;
	wire _w18555_ ;
	wire _w18556_ ;
	wire _w18557_ ;
	wire _w18558_ ;
	wire _w18559_ ;
	wire _w18560_ ;
	wire _w18561_ ;
	wire _w18562_ ;
	wire _w18563_ ;
	wire _w18564_ ;
	wire _w18565_ ;
	wire _w18566_ ;
	wire _w18567_ ;
	wire _w18568_ ;
	wire _w18569_ ;
	wire _w18570_ ;
	wire _w18571_ ;
	wire _w18572_ ;
	wire _w18573_ ;
	wire _w18574_ ;
	wire _w18575_ ;
	wire _w18576_ ;
	wire _w18577_ ;
	wire _w18578_ ;
	wire _w18579_ ;
	wire _w18580_ ;
	wire _w18581_ ;
	wire _w18582_ ;
	wire _w18583_ ;
	wire _w18584_ ;
	wire _w18585_ ;
	wire _w18586_ ;
	wire _w18587_ ;
	wire _w18588_ ;
	wire _w18589_ ;
	wire _w18590_ ;
	wire _w18591_ ;
	wire _w18592_ ;
	wire _w18593_ ;
	wire _w18594_ ;
	wire _w18595_ ;
	wire _w18596_ ;
	wire _w18597_ ;
	wire _w18598_ ;
	wire _w18599_ ;
	wire _w18600_ ;
	wire _w18601_ ;
	wire _w18602_ ;
	wire _w18603_ ;
	wire _w18604_ ;
	wire _w18605_ ;
	wire _w18606_ ;
	wire _w18607_ ;
	wire _w18608_ ;
	wire _w18609_ ;
	wire _w18610_ ;
	wire _w18611_ ;
	wire _w18612_ ;
	wire _w18613_ ;
	wire _w18614_ ;
	wire _w18615_ ;
	wire _w18616_ ;
	wire _w18617_ ;
	wire _w18618_ ;
	wire _w18619_ ;
	wire _w18620_ ;
	wire _w18621_ ;
	wire _w18622_ ;
	wire _w18623_ ;
	wire _w18624_ ;
	wire _w18625_ ;
	wire _w18626_ ;
	wire _w18627_ ;
	wire _w18628_ ;
	wire _w18629_ ;
	wire _w18630_ ;
	wire _w18631_ ;
	wire _w18632_ ;
	wire _w18633_ ;
	wire _w18634_ ;
	wire _w18635_ ;
	wire _w18636_ ;
	wire _w18637_ ;
	wire _w18638_ ;
	wire _w18639_ ;
	wire _w18640_ ;
	wire _w18641_ ;
	wire _w18642_ ;
	wire _w18643_ ;
	wire _w18644_ ;
	wire _w18645_ ;
	wire _w18646_ ;
	wire _w18647_ ;
	wire _w18648_ ;
	wire _w18649_ ;
	wire _w18650_ ;
	wire _w18651_ ;
	wire _w18652_ ;
	wire _w18653_ ;
	wire _w18654_ ;
	wire _w18655_ ;
	wire _w18656_ ;
	wire _w18657_ ;
	wire _w18658_ ;
	wire _w18659_ ;
	wire _w18660_ ;
	wire _w18661_ ;
	wire _w18662_ ;
	wire _w18663_ ;
	wire _w18664_ ;
	wire _w18665_ ;
	wire _w18666_ ;
	wire _w18667_ ;
	wire _w18668_ ;
	wire _w18669_ ;
	wire _w18670_ ;
	wire _w18671_ ;
	wire _w18672_ ;
	wire _w18673_ ;
	wire _w18674_ ;
	wire _w18675_ ;
	wire _w18676_ ;
	wire _w18677_ ;
	wire _w18678_ ;
	wire _w18679_ ;
	wire _w18680_ ;
	wire _w18681_ ;
	wire _w18682_ ;
	wire _w18683_ ;
	wire _w18684_ ;
	wire _w18685_ ;
	wire _w18686_ ;
	wire _w18687_ ;
	wire _w18688_ ;
	wire _w18689_ ;
	wire _w18690_ ;
	wire _w18691_ ;
	wire _w18692_ ;
	wire _w18693_ ;
	wire _w18694_ ;
	wire _w18695_ ;
	wire _w18696_ ;
	wire _w18697_ ;
	wire _w18698_ ;
	wire _w18699_ ;
	wire _w18700_ ;
	wire _w18701_ ;
	wire _w18702_ ;
	wire _w18703_ ;
	wire _w18704_ ;
	wire _w18705_ ;
	wire _w18706_ ;
	wire _w18707_ ;
	wire _w18708_ ;
	wire _w18709_ ;
	wire _w18710_ ;
	wire _w18711_ ;
	wire _w18712_ ;
	wire _w18713_ ;
	wire _w18714_ ;
	wire _w18715_ ;
	wire _w18716_ ;
	wire _w18717_ ;
	wire _w18718_ ;
	wire _w18719_ ;
	wire _w18720_ ;
	wire _w18721_ ;
	wire _w18722_ ;
	wire _w18723_ ;
	wire _w18724_ ;
	wire _w18725_ ;
	wire _w18726_ ;
	wire _w18727_ ;
	wire _w18728_ ;
	wire _w18729_ ;
	wire _w18730_ ;
	wire _w18731_ ;
	wire _w18732_ ;
	wire _w18733_ ;
	wire _w18734_ ;
	wire _w18735_ ;
	wire _w18736_ ;
	wire _w18737_ ;
	wire _w18738_ ;
	wire _w18739_ ;
	wire _w18740_ ;
	wire _w18741_ ;
	wire _w18742_ ;
	wire _w18743_ ;
	wire _w18744_ ;
	wire _w18745_ ;
	wire _w18746_ ;
	wire _w18747_ ;
	wire _w18748_ ;
	wire _w18749_ ;
	wire _w18750_ ;
	wire _w18751_ ;
	wire _w18752_ ;
	wire _w18753_ ;
	wire _w18754_ ;
	wire _w18755_ ;
	wire _w18756_ ;
	wire _w18757_ ;
	wire _w18758_ ;
	wire _w18759_ ;
	wire _w18760_ ;
	wire _w18761_ ;
	wire _w18762_ ;
	wire _w18763_ ;
	wire _w18764_ ;
	wire _w18765_ ;
	wire _w18766_ ;
	wire _w18767_ ;
	wire _w18768_ ;
	wire _w18769_ ;
	wire _w18770_ ;
	wire _w18771_ ;
	wire _w18772_ ;
	wire _w18773_ ;
	wire _w18774_ ;
	wire _w18775_ ;
	wire _w18776_ ;
	wire _w18777_ ;
	wire _w18778_ ;
	wire _w18779_ ;
	wire _w18780_ ;
	wire _w18781_ ;
	wire _w18782_ ;
	wire _w18783_ ;
	wire _w18784_ ;
	wire _w18785_ ;
	wire _w18786_ ;
	wire _w18787_ ;
	wire _w18788_ ;
	wire _w18789_ ;
	wire _w18790_ ;
	wire _w18791_ ;
	wire _w18792_ ;
	wire _w18793_ ;
	wire _w18794_ ;
	wire _w18795_ ;
	wire _w18796_ ;
	wire _w18797_ ;
	wire _w18798_ ;
	wire _w18799_ ;
	wire _w18800_ ;
	wire _w18801_ ;
	wire _w18802_ ;
	wire _w18803_ ;
	wire _w18804_ ;
	wire _w18805_ ;
	wire _w18806_ ;
	wire _w18807_ ;
	wire _w18808_ ;
	wire _w18809_ ;
	wire _w18810_ ;
	wire _w18811_ ;
	wire _w18812_ ;
	wire _w18813_ ;
	wire _w18814_ ;
	wire _w18815_ ;
	wire _w18816_ ;
	wire _w18817_ ;
	wire _w18818_ ;
	wire _w18819_ ;
	wire _w18820_ ;
	wire _w18821_ ;
	wire _w18822_ ;
	wire _w18823_ ;
	wire _w18824_ ;
	wire _w18825_ ;
	wire _w18826_ ;
	wire _w18827_ ;
	wire _w18828_ ;
	wire _w18829_ ;
	wire _w18830_ ;
	wire _w18831_ ;
	wire _w18832_ ;
	wire _w18833_ ;
	wire _w18834_ ;
	wire _w18835_ ;
	wire _w18836_ ;
	wire _w18837_ ;
	wire _w18838_ ;
	wire _w18839_ ;
	wire _w18840_ ;
	wire _w18841_ ;
	wire _w18842_ ;
	wire _w18843_ ;
	wire _w18844_ ;
	wire _w18845_ ;
	wire _w18846_ ;
	wire _w18847_ ;
	wire _w18848_ ;
	wire _w18849_ ;
	wire _w18850_ ;
	wire _w18851_ ;
	wire _w18852_ ;
	wire _w18853_ ;
	wire _w18854_ ;
	wire _w18855_ ;
	wire _w18856_ ;
	wire _w18857_ ;
	wire _w18858_ ;
	wire _w18859_ ;
	wire _w18860_ ;
	wire _w18861_ ;
	wire _w18862_ ;
	wire _w18863_ ;
	wire _w18864_ ;
	wire _w18865_ ;
	wire _w18866_ ;
	wire _w18867_ ;
	wire _w18868_ ;
	wire _w18869_ ;
	wire _w18870_ ;
	wire _w18871_ ;
	wire _w18872_ ;
	wire _w18873_ ;
	wire _w18874_ ;
	wire _w18875_ ;
	wire _w18876_ ;
	wire _w18877_ ;
	wire _w18878_ ;
	wire _w18879_ ;
	wire _w18880_ ;
	wire _w18881_ ;
	wire _w18882_ ;
	wire _w18883_ ;
	wire _w18884_ ;
	wire _w18885_ ;
	wire _w18886_ ;
	wire _w18887_ ;
	wire _w18888_ ;
	wire _w18889_ ;
	wire _w18890_ ;
	wire _w18891_ ;
	wire _w18892_ ;
	wire _w18893_ ;
	wire _w18894_ ;
	wire _w18895_ ;
	wire _w18896_ ;
	wire _w18897_ ;
	wire _w18898_ ;
	wire _w18899_ ;
	wire _w18900_ ;
	wire _w18901_ ;
	wire _w18902_ ;
	wire _w18903_ ;
	wire _w18904_ ;
	wire _w18905_ ;
	wire _w18906_ ;
	wire _w18907_ ;
	wire _w18908_ ;
	wire _w18909_ ;
	wire _w18910_ ;
	wire _w18911_ ;
	wire _w18912_ ;
	wire _w18913_ ;
	wire _w18914_ ;
	wire _w18915_ ;
	wire _w18916_ ;
	wire _w18917_ ;
	wire _w18918_ ;
	wire _w18919_ ;
	wire _w18920_ ;
	wire _w18921_ ;
	wire _w18922_ ;
	wire _w18923_ ;
	wire _w18924_ ;
	wire _w18925_ ;
	wire _w18926_ ;
	wire _w18927_ ;
	wire _w18928_ ;
	wire _w18929_ ;
	wire _w18930_ ;
	wire _w18931_ ;
	wire _w18932_ ;
	wire _w18933_ ;
	wire _w18934_ ;
	wire _w18935_ ;
	wire _w18936_ ;
	wire _w18937_ ;
	wire _w18938_ ;
	wire _w18939_ ;
	wire _w18940_ ;
	wire _w18941_ ;
	wire _w18942_ ;
	wire _w18943_ ;
	wire _w18944_ ;
	wire _w18945_ ;
	wire _w18946_ ;
	wire _w18947_ ;
	wire _w18948_ ;
	wire _w18949_ ;
	wire _w18950_ ;
	wire _w18951_ ;
	wire _w18952_ ;
	wire _w18953_ ;
	wire _w18954_ ;
	wire _w18955_ ;
	wire _w18956_ ;
	wire _w18957_ ;
	wire _w18958_ ;
	wire _w18959_ ;
	wire _w18960_ ;
	wire _w18961_ ;
	wire _w18962_ ;
	wire _w18963_ ;
	wire _w18964_ ;
	wire _w18965_ ;
	wire _w18966_ ;
	wire _w18967_ ;
	wire _w18968_ ;
	wire _w18969_ ;
	wire _w18970_ ;
	wire _w18971_ ;
	wire _w18972_ ;
	wire _w18973_ ;
	wire _w18974_ ;
	wire _w18975_ ;
	wire _w18976_ ;
	wire _w18977_ ;
	wire _w18978_ ;
	wire _w18979_ ;
	wire _w18980_ ;
	wire _w18981_ ;
	wire _w18982_ ;
	wire _w18983_ ;
	wire _w18984_ ;
	wire _w18985_ ;
	wire _w18986_ ;
	wire _w18987_ ;
	wire _w18988_ ;
	wire _w18989_ ;
	wire _w18990_ ;
	wire _w18991_ ;
	wire _w18992_ ;
	wire _w18993_ ;
	wire _w18994_ ;
	wire _w18995_ ;
	wire _w18996_ ;
	wire _w18997_ ;
	wire _w18998_ ;
	wire _w18999_ ;
	wire _w19000_ ;
	wire _w19001_ ;
	wire _w19002_ ;
	wire _w19003_ ;
	wire _w19004_ ;
	wire _w19005_ ;
	wire _w19006_ ;
	wire _w19007_ ;
	wire _w19008_ ;
	wire _w19009_ ;
	wire _w19010_ ;
	wire _w19011_ ;
	wire _w19012_ ;
	wire _w19013_ ;
	wire _w19014_ ;
	wire _w19015_ ;
	wire _w19016_ ;
	wire _w19017_ ;
	wire _w19018_ ;
	wire _w19019_ ;
	wire _w19020_ ;
	wire _w19021_ ;
	wire _w19022_ ;
	wire _w19023_ ;
	wire _w19024_ ;
	wire _w19025_ ;
	wire _w19026_ ;
	wire _w19027_ ;
	wire _w19028_ ;
	wire _w19029_ ;
	wire _w19030_ ;
	wire _w19031_ ;
	wire _w19032_ ;
	wire _w19033_ ;
	wire _w19034_ ;
	wire _w19035_ ;
	wire _w19036_ ;
	wire _w19037_ ;
	wire _w19038_ ;
	wire _w19039_ ;
	wire _w19040_ ;
	wire _w19041_ ;
	wire _w19042_ ;
	wire _w19043_ ;
	wire _w19044_ ;
	wire _w19045_ ;
	wire _w19046_ ;
	wire _w19047_ ;
	wire _w19048_ ;
	wire _w19049_ ;
	wire _w19050_ ;
	wire _w19051_ ;
	wire _w19052_ ;
	wire _w19053_ ;
	wire _w19054_ ;
	wire _w19055_ ;
	wire _w19056_ ;
	wire _w19057_ ;
	wire _w19058_ ;
	wire _w19059_ ;
	wire _w19060_ ;
	wire _w19061_ ;
	wire _w19062_ ;
	wire _w19063_ ;
	wire _w19064_ ;
	wire _w19065_ ;
	wire _w19066_ ;
	wire _w19067_ ;
	wire _w19068_ ;
	wire _w19069_ ;
	wire _w19070_ ;
	wire _w19071_ ;
	wire _w19072_ ;
	wire _w19073_ ;
	wire _w19074_ ;
	wire _w19075_ ;
	wire _w19076_ ;
	wire _w19077_ ;
	wire _w19078_ ;
	wire _w19079_ ;
	wire _w19080_ ;
	wire _w19081_ ;
	wire _w19082_ ;
	wire _w19083_ ;
	wire _w19084_ ;
	wire _w19085_ ;
	wire _w19086_ ;
	wire _w19087_ ;
	wire _w19088_ ;
	wire _w19089_ ;
	wire _w19090_ ;
	wire _w19091_ ;
	wire _w19092_ ;
	wire _w19093_ ;
	wire _w19094_ ;
	wire _w19095_ ;
	wire _w19096_ ;
	wire _w19097_ ;
	wire _w19098_ ;
	wire _w19099_ ;
	wire _w19100_ ;
	wire _w19101_ ;
	wire _w19102_ ;
	wire _w19103_ ;
	wire _w19104_ ;
	wire _w19105_ ;
	wire _w19106_ ;
	wire _w19107_ ;
	wire _w19108_ ;
	wire _w19109_ ;
	wire _w19110_ ;
	wire _w19111_ ;
	wire _w19112_ ;
	wire _w19113_ ;
	wire _w19114_ ;
	wire _w19115_ ;
	wire _w19116_ ;
	wire _w19117_ ;
	wire _w19118_ ;
	wire _w19119_ ;
	wire _w19120_ ;
	wire _w19121_ ;
	wire _w19122_ ;
	wire _w19123_ ;
	wire _w19124_ ;
	wire _w19125_ ;
	wire _w19126_ ;
	wire _w19127_ ;
	wire _w19128_ ;
	wire _w19129_ ;
	wire _w19130_ ;
	wire _w19131_ ;
	wire _w19132_ ;
	wire _w19133_ ;
	wire _w19134_ ;
	wire _w19135_ ;
	wire _w19136_ ;
	wire _w19137_ ;
	wire _w19138_ ;
	wire _w19139_ ;
	wire _w19140_ ;
	wire _w19141_ ;
	wire _w19142_ ;
	wire _w19143_ ;
	wire _w19144_ ;
	wire _w19145_ ;
	wire _w19146_ ;
	wire _w19147_ ;
	wire _w19148_ ;
	wire _w19149_ ;
	wire _w19150_ ;
	wire _w19151_ ;
	wire _w19152_ ;
	wire _w19153_ ;
	wire _w19154_ ;
	wire _w19155_ ;
	wire _w19156_ ;
	wire _w19157_ ;
	wire _w19158_ ;
	wire _w19159_ ;
	wire _w19160_ ;
	wire _w19161_ ;
	wire _w19162_ ;
	wire _w19163_ ;
	wire _w19164_ ;
	wire _w19165_ ;
	wire _w19166_ ;
	wire _w19167_ ;
	wire _w19168_ ;
	wire _w19169_ ;
	wire _w19170_ ;
	wire _w19171_ ;
	wire _w19172_ ;
	wire _w19173_ ;
	wire _w19174_ ;
	wire _w19175_ ;
	wire _w19176_ ;
	wire _w19177_ ;
	wire _w19178_ ;
	wire _w19179_ ;
	wire _w19180_ ;
	wire _w19181_ ;
	wire _w19182_ ;
	wire _w19183_ ;
	wire _w19184_ ;
	wire _w19185_ ;
	wire _w19186_ ;
	wire _w19187_ ;
	wire _w19188_ ;
	wire _w19189_ ;
	wire _w19190_ ;
	wire _w19191_ ;
	wire _w19192_ ;
	wire _w19193_ ;
	wire _w19194_ ;
	wire _w19195_ ;
	wire _w19196_ ;
	wire _w19197_ ;
	wire _w19198_ ;
	wire _w19199_ ;
	wire _w19200_ ;
	wire _w19201_ ;
	wire _w19202_ ;
	wire _w19203_ ;
	wire _w19204_ ;
	wire _w19205_ ;
	wire _w19206_ ;
	wire _w19207_ ;
	wire _w19208_ ;
	wire _w19209_ ;
	wire _w19210_ ;
	wire _w19211_ ;
	wire _w19212_ ;
	wire _w19213_ ;
	wire _w19214_ ;
	wire _w19215_ ;
	wire _w19216_ ;
	wire _w19217_ ;
	wire _w19218_ ;
	wire _w19219_ ;
	wire _w19220_ ;
	wire _w19221_ ;
	wire _w19222_ ;
	wire _w19223_ ;
	wire _w19224_ ;
	wire _w19225_ ;
	wire _w19226_ ;
	wire _w19227_ ;
	wire _w19228_ ;
	wire _w19229_ ;
	wire _w19230_ ;
	wire _w19231_ ;
	wire _w19232_ ;
	wire _w19233_ ;
	wire _w19234_ ;
	wire _w19235_ ;
	wire _w19236_ ;
	wire _w19237_ ;
	wire _w19238_ ;
	wire _w19239_ ;
	wire _w19240_ ;
	wire _w19241_ ;
	wire _w19242_ ;
	wire _w19243_ ;
	wire _w19244_ ;
	wire _w19245_ ;
	wire _w19246_ ;
	wire _w19247_ ;
	wire _w19248_ ;
	wire _w19249_ ;
	wire _w19250_ ;
	wire _w19251_ ;
	wire _w19252_ ;
	wire _w19253_ ;
	wire _w19254_ ;
	wire _w19255_ ;
	wire _w19256_ ;
	wire _w19257_ ;
	wire _w19258_ ;
	wire _w19259_ ;
	wire _w19260_ ;
	wire _w19261_ ;
	wire _w19262_ ;
	wire _w19263_ ;
	wire _w19264_ ;
	wire _w19265_ ;
	wire _w19266_ ;
	wire _w19267_ ;
	wire _w19268_ ;
	wire _w19269_ ;
	wire _w19270_ ;
	wire _w19271_ ;
	wire _w19272_ ;
	wire _w19273_ ;
	wire _w19274_ ;
	wire _w19275_ ;
	wire _w19276_ ;
	wire _w19277_ ;
	wire _w19278_ ;
	wire _w19279_ ;
	wire _w19280_ ;
	wire _w19281_ ;
	wire _w19282_ ;
	wire _w19283_ ;
	wire _w19284_ ;
	wire _w19285_ ;
	wire _w19286_ ;
	wire _w19287_ ;
	wire _w19288_ ;
	wire _w19289_ ;
	wire _w19290_ ;
	wire _w19291_ ;
	wire _w19292_ ;
	wire _w19293_ ;
	wire _w19294_ ;
	wire _w19295_ ;
	wire _w19296_ ;
	wire _w19297_ ;
	wire _w19298_ ;
	wire _w19299_ ;
	wire _w19300_ ;
	wire _w19301_ ;
	wire _w19302_ ;
	wire _w19303_ ;
	wire _w19304_ ;
	wire _w19305_ ;
	wire _w19306_ ;
	wire _w19307_ ;
	wire _w19308_ ;
	wire _w19309_ ;
	wire _w19310_ ;
	wire _w19311_ ;
	wire _w19312_ ;
	wire _w19313_ ;
	wire _w19314_ ;
	wire _w19315_ ;
	wire _w19316_ ;
	wire _w19317_ ;
	wire _w19318_ ;
	wire _w19319_ ;
	wire _w19320_ ;
	wire _w19321_ ;
	wire _w19322_ ;
	wire _w19323_ ;
	wire _w19324_ ;
	wire _w19325_ ;
	wire _w19326_ ;
	wire _w19327_ ;
	wire _w19328_ ;
	wire _w19329_ ;
	wire _w19330_ ;
	wire _w19331_ ;
	wire _w19332_ ;
	wire _w19333_ ;
	wire _w19334_ ;
	wire _w19335_ ;
	wire _w19336_ ;
	wire _w19337_ ;
	wire _w19338_ ;
	wire _w19339_ ;
	wire _w19340_ ;
	wire _w19341_ ;
	wire _w19342_ ;
	wire _w19343_ ;
	wire _w19344_ ;
	wire _w19345_ ;
	wire _w19346_ ;
	wire _w19347_ ;
	wire _w19348_ ;
	wire _w19349_ ;
	wire _w19350_ ;
	wire _w19351_ ;
	wire _w19352_ ;
	wire _w19353_ ;
	wire _w19354_ ;
	wire _w19355_ ;
	wire _w19356_ ;
	wire _w19357_ ;
	wire _w19358_ ;
	wire _w19359_ ;
	wire _w19360_ ;
	wire _w19361_ ;
	wire _w19362_ ;
	wire _w19363_ ;
	wire _w19364_ ;
	wire _w19365_ ;
	wire _w19366_ ;
	wire _w19367_ ;
	wire _w19368_ ;
	wire _w19369_ ;
	wire _w19370_ ;
	wire _w19371_ ;
	wire _w19372_ ;
	wire _w19373_ ;
	wire _w19374_ ;
	wire _w19375_ ;
	wire _w19376_ ;
	wire _w19377_ ;
	wire _w19378_ ;
	wire _w19379_ ;
	wire _w19380_ ;
	wire _w19381_ ;
	wire _w19382_ ;
	wire _w19383_ ;
	wire _w19384_ ;
	wire _w19385_ ;
	wire _w19386_ ;
	wire _w19387_ ;
	wire _w19388_ ;
	wire _w19389_ ;
	wire _w19390_ ;
	wire _w19391_ ;
	wire _w19392_ ;
	wire _w19393_ ;
	wire _w19394_ ;
	wire _w19395_ ;
	wire _w19396_ ;
	wire _w19397_ ;
	wire _w19398_ ;
	wire _w19399_ ;
	wire _w19400_ ;
	wire _w19401_ ;
	wire _w19402_ ;
	wire _w19403_ ;
	wire _w19404_ ;
	wire _w19405_ ;
	wire _w19406_ ;
	wire _w19407_ ;
	wire _w19408_ ;
	wire _w19409_ ;
	wire _w19410_ ;
	wire _w19411_ ;
	wire _w19412_ ;
	wire _w19413_ ;
	wire _w19414_ ;
	wire _w19415_ ;
	wire _w19416_ ;
	wire _w19417_ ;
	wire _w19418_ ;
	wire _w19419_ ;
	wire _w19420_ ;
	wire _w19421_ ;
	wire _w19422_ ;
	wire _w19423_ ;
	wire _w19424_ ;
	wire _w19425_ ;
	wire _w19426_ ;
	wire _w19427_ ;
	wire _w19428_ ;
	wire _w19429_ ;
	wire _w19430_ ;
	wire _w19431_ ;
	wire _w19432_ ;
	wire _w19433_ ;
	wire _w19434_ ;
	wire _w19435_ ;
	wire _w19436_ ;
	wire _w19437_ ;
	wire _w19438_ ;
	wire _w19439_ ;
	wire _w19440_ ;
	wire _w19441_ ;
	wire _w19442_ ;
	wire _w19443_ ;
	wire _w19444_ ;
	wire _w19445_ ;
	wire _w19446_ ;
	wire _w19447_ ;
	wire _w19448_ ;
	wire _w19449_ ;
	wire _w19450_ ;
	wire _w19451_ ;
	wire _w19452_ ;
	wire _w19453_ ;
	wire _w19454_ ;
	wire _w19455_ ;
	wire _w19456_ ;
	wire _w19457_ ;
	wire _w19458_ ;
	wire _w19459_ ;
	wire _w19460_ ;
	wire _w19461_ ;
	wire _w19462_ ;
	wire _w19463_ ;
	wire _w19464_ ;
	wire _w19465_ ;
	wire _w19466_ ;
	wire _w19467_ ;
	wire _w19468_ ;
	wire _w19469_ ;
	wire _w19470_ ;
	wire _w19471_ ;
	wire _w19472_ ;
	wire _w19473_ ;
	wire _w19474_ ;
	wire _w19475_ ;
	wire _w19476_ ;
	wire _w19477_ ;
	wire _w19478_ ;
	wire _w19479_ ;
	wire _w19480_ ;
	wire _w19481_ ;
	wire _w19482_ ;
	wire _w19483_ ;
	wire _w19484_ ;
	wire _w19485_ ;
	wire _w19486_ ;
	wire _w19487_ ;
	wire _w19488_ ;
	wire _w19489_ ;
	wire _w19490_ ;
	wire _w19491_ ;
	wire _w19492_ ;
	wire _w19493_ ;
	wire _w19494_ ;
	wire _w19495_ ;
	wire _w19496_ ;
	wire _w19497_ ;
	wire _w19498_ ;
	wire _w19499_ ;
	wire _w19500_ ;
	wire _w19501_ ;
	wire _w19502_ ;
	wire _w19503_ ;
	wire _w19504_ ;
	wire _w19505_ ;
	wire _w19506_ ;
	wire _w19507_ ;
	wire _w19508_ ;
	wire _w19509_ ;
	wire _w19510_ ;
	wire _w19511_ ;
	wire _w19512_ ;
	wire _w19513_ ;
	wire _w19514_ ;
	wire _w19515_ ;
	wire _w19516_ ;
	wire _w19517_ ;
	wire _w19518_ ;
	wire _w19519_ ;
	wire _w19520_ ;
	wire _w19521_ ;
	wire _w19522_ ;
	wire _w19523_ ;
	wire _w19524_ ;
	wire _w19525_ ;
	wire _w19526_ ;
	wire _w19527_ ;
	wire _w19528_ ;
	wire _w19529_ ;
	wire _w19530_ ;
	wire _w19531_ ;
	wire _w19532_ ;
	wire _w19533_ ;
	wire _w19534_ ;
	wire _w19535_ ;
	wire _w19536_ ;
	wire _w19537_ ;
	wire _w19538_ ;
	wire _w19539_ ;
	wire _w19540_ ;
	wire _w19541_ ;
	wire _w19542_ ;
	wire _w19543_ ;
	wire _w19544_ ;
	wire _w19545_ ;
	wire _w19546_ ;
	wire _w19547_ ;
	wire _w19548_ ;
	wire _w19549_ ;
	wire _w19550_ ;
	wire _w19551_ ;
	wire _w19552_ ;
	wire _w19553_ ;
	wire _w19554_ ;
	wire _w19555_ ;
	wire _w19556_ ;
	wire _w19557_ ;
	wire _w19558_ ;
	wire _w19559_ ;
	wire _w19560_ ;
	wire _w19561_ ;
	wire _w19562_ ;
	wire _w19563_ ;
	wire _w19564_ ;
	wire _w19565_ ;
	wire _w19566_ ;
	wire _w19567_ ;
	wire _w19568_ ;
	wire _w19569_ ;
	wire _w19570_ ;
	wire _w19571_ ;
	wire _w19572_ ;
	wire _w19573_ ;
	wire _w19574_ ;
	wire _w19575_ ;
	wire _w19576_ ;
	wire _w19577_ ;
	wire _w19578_ ;
	wire _w19579_ ;
	wire _w19580_ ;
	wire _w19581_ ;
	wire _w19582_ ;
	wire _w19583_ ;
	wire _w19584_ ;
	wire _w19585_ ;
	wire _w19586_ ;
	wire _w19587_ ;
	wire _w19588_ ;
	wire _w19589_ ;
	wire _w19590_ ;
	wire _w19591_ ;
	wire _w19592_ ;
	wire _w19593_ ;
	wire _w19594_ ;
	wire _w19595_ ;
	wire _w19596_ ;
	wire _w19597_ ;
	wire _w19598_ ;
	wire _w19599_ ;
	wire _w19600_ ;
	wire _w19601_ ;
	wire _w19602_ ;
	wire _w19603_ ;
	wire _w19604_ ;
	wire _w19605_ ;
	wire _w19606_ ;
	wire _w19607_ ;
	wire _w19608_ ;
	wire _w19609_ ;
	wire _w19610_ ;
	wire _w19611_ ;
	wire _w19612_ ;
	wire _w19613_ ;
	wire _w19614_ ;
	wire _w19615_ ;
	wire _w19616_ ;
	wire _w19617_ ;
	wire _w19618_ ;
	wire _w19619_ ;
	wire _w19620_ ;
	wire _w19621_ ;
	wire _w19622_ ;
	wire _w19623_ ;
	wire _w19624_ ;
	wire _w19625_ ;
	wire _w19626_ ;
	wire _w19627_ ;
	wire _w19628_ ;
	wire _w19629_ ;
	wire _w19630_ ;
	wire _w19631_ ;
	wire _w19632_ ;
	wire _w19633_ ;
	wire _w19634_ ;
	wire _w19635_ ;
	wire _w19636_ ;
	wire _w19637_ ;
	wire _w19638_ ;
	wire _w19639_ ;
	wire _w19640_ ;
	wire _w19641_ ;
	wire _w19642_ ;
	wire _w19643_ ;
	wire _w19644_ ;
	wire _w19645_ ;
	wire _w19646_ ;
	wire _w19647_ ;
	wire _w19648_ ;
	wire _w19649_ ;
	wire _w19650_ ;
	wire _w19651_ ;
	wire _w19652_ ;
	wire _w19653_ ;
	wire _w19654_ ;
	wire _w19655_ ;
	wire _w19656_ ;
	wire _w19657_ ;
	wire _w19658_ ;
	wire _w19659_ ;
	wire _w19660_ ;
	wire _w19661_ ;
	wire _w19662_ ;
	wire _w19663_ ;
	wire _w19664_ ;
	wire _w19665_ ;
	wire _w19666_ ;
	wire _w19667_ ;
	wire _w19668_ ;
	wire _w19669_ ;
	wire _w19670_ ;
	wire _w19671_ ;
	wire _w19672_ ;
	wire _w19673_ ;
	wire _w19674_ ;
	wire _w19675_ ;
	wire _w19676_ ;
	wire _w19677_ ;
	wire _w19678_ ;
	wire _w19679_ ;
	wire _w19680_ ;
	wire _w19681_ ;
	wire _w19682_ ;
	wire _w19683_ ;
	wire _w19684_ ;
	wire _w19685_ ;
	wire _w19686_ ;
	wire _w19687_ ;
	wire _w19688_ ;
	wire _w19689_ ;
	wire _w19690_ ;
	wire _w19691_ ;
	wire _w19692_ ;
	wire _w19693_ ;
	wire _w19694_ ;
	wire _w19695_ ;
	wire _w19696_ ;
	wire _w19697_ ;
	wire _w19698_ ;
	wire _w19699_ ;
	wire _w19700_ ;
	wire _w19701_ ;
	wire _w19702_ ;
	wire _w19703_ ;
	wire _w19704_ ;
	wire _w19705_ ;
	wire _w19706_ ;
	wire _w19707_ ;
	wire _w19708_ ;
	wire _w19709_ ;
	wire _w19710_ ;
	wire _w19711_ ;
	wire _w19712_ ;
	wire _w19713_ ;
	wire _w19714_ ;
	wire _w19715_ ;
	wire _w19716_ ;
	wire _w19717_ ;
	wire _w19718_ ;
	wire _w19719_ ;
	wire _w19720_ ;
	wire _w19721_ ;
	wire _w19722_ ;
	wire _w19723_ ;
	wire _w19724_ ;
	wire _w19725_ ;
	wire _w19726_ ;
	wire _w19727_ ;
	wire _w19728_ ;
	wire _w19729_ ;
	wire _w19730_ ;
	wire _w19731_ ;
	wire _w19732_ ;
	wire _w19733_ ;
	wire _w19734_ ;
	wire _w19735_ ;
	wire _w19736_ ;
	wire _w19737_ ;
	wire _w19738_ ;
	wire _w19739_ ;
	wire _w19740_ ;
	wire _w19741_ ;
	wire _w19742_ ;
	wire _w19743_ ;
	wire _w19744_ ;
	wire _w19745_ ;
	wire _w19746_ ;
	wire _w19747_ ;
	wire _w19748_ ;
	wire _w19749_ ;
	wire _w19750_ ;
	wire _w19751_ ;
	wire _w19752_ ;
	wire _w19753_ ;
	wire _w19754_ ;
	wire _w19755_ ;
	wire _w19756_ ;
	wire _w19757_ ;
	wire _w19758_ ;
	wire _w19759_ ;
	wire _w19760_ ;
	wire _w19761_ ;
	wire _w19762_ ;
	wire _w19763_ ;
	wire _w19764_ ;
	wire _w19765_ ;
	wire _w19766_ ;
	wire _w19767_ ;
	wire _w19768_ ;
	wire _w19769_ ;
	wire _w19770_ ;
	wire _w19771_ ;
	wire _w19772_ ;
	wire _w19773_ ;
	wire _w19774_ ;
	wire _w19775_ ;
	wire _w19776_ ;
	wire _w19777_ ;
	wire _w19778_ ;
	wire _w19779_ ;
	wire _w19780_ ;
	wire _w19781_ ;
	wire _w19782_ ;
	wire _w19783_ ;
	wire _w19784_ ;
	wire _w19785_ ;
	wire _w19786_ ;
	wire _w19787_ ;
	wire _w19788_ ;
	wire _w19789_ ;
	wire _w19790_ ;
	wire _w19791_ ;
	wire _w19792_ ;
	wire _w19793_ ;
	wire _w19794_ ;
	wire _w19795_ ;
	wire _w19796_ ;
	wire _w19797_ ;
	wire _w19798_ ;
	wire _w19799_ ;
	wire _w19800_ ;
	wire _w19801_ ;
	wire _w19802_ ;
	wire _w19803_ ;
	wire _w19804_ ;
	wire _w19805_ ;
	wire _w19806_ ;
	wire _w19807_ ;
	wire _w19808_ ;
	wire _w19809_ ;
	wire _w19810_ ;
	wire _w19811_ ;
	wire _w19812_ ;
	wire _w19813_ ;
	wire _w19814_ ;
	wire _w19815_ ;
	wire _w19816_ ;
	wire _w19817_ ;
	wire _w19818_ ;
	wire _w19819_ ;
	wire _w19820_ ;
	wire _w19821_ ;
	wire _w19822_ ;
	wire _w19823_ ;
	wire _w19824_ ;
	wire _w19825_ ;
	wire _w19826_ ;
	wire _w19827_ ;
	wire _w19828_ ;
	wire _w19829_ ;
	wire _w19830_ ;
	wire _w19831_ ;
	wire _w19832_ ;
	wire _w19833_ ;
	wire _w19834_ ;
	wire _w19835_ ;
	wire _w19836_ ;
	wire _w19837_ ;
	wire _w19838_ ;
	wire _w19839_ ;
	wire _w19840_ ;
	wire _w19841_ ;
	wire _w19842_ ;
	wire _w19843_ ;
	wire _w19844_ ;
	wire _w19845_ ;
	wire _w19846_ ;
	wire _w19847_ ;
	wire _w19848_ ;
	wire _w19849_ ;
	wire _w19850_ ;
	wire _w19851_ ;
	wire _w19852_ ;
	wire _w19853_ ;
	wire _w19854_ ;
	wire _w19855_ ;
	wire _w19856_ ;
	wire _w19857_ ;
	wire _w19858_ ;
	wire _w19859_ ;
	wire _w19860_ ;
	wire _w19861_ ;
	wire _w19862_ ;
	wire _w19863_ ;
	wire _w19864_ ;
	wire _w19865_ ;
	wire _w19866_ ;
	wire _w19867_ ;
	wire _w19868_ ;
	wire _w19869_ ;
	wire _w19870_ ;
	wire _w19871_ ;
	wire _w19872_ ;
	wire _w19873_ ;
	wire _w19874_ ;
	wire _w19875_ ;
	wire _w19876_ ;
	wire _w19877_ ;
	wire _w19878_ ;
	wire _w19879_ ;
	wire _w19880_ ;
	wire _w19881_ ;
	wire _w19882_ ;
	wire _w19883_ ;
	wire _w19884_ ;
	wire _w19885_ ;
	wire _w19886_ ;
	wire _w19887_ ;
	wire _w19888_ ;
	wire _w19889_ ;
	wire _w19890_ ;
	wire _w19891_ ;
	wire _w19892_ ;
	wire _w19893_ ;
	wire _w19894_ ;
	wire _w19895_ ;
	wire _w19896_ ;
	wire _w19897_ ;
	wire _w19898_ ;
	wire _w19899_ ;
	wire _w19900_ ;
	wire _w19901_ ;
	wire _w19902_ ;
	wire _w19903_ ;
	wire _w19904_ ;
	wire _w19905_ ;
	wire _w19906_ ;
	wire _w19907_ ;
	wire _w19908_ ;
	wire _w19909_ ;
	wire _w19910_ ;
	wire _w19911_ ;
	wire _w19912_ ;
	wire _w19913_ ;
	wire _w19914_ ;
	wire _w19915_ ;
	wire _w19916_ ;
	wire _w19917_ ;
	wire _w19918_ ;
	wire _w19919_ ;
	wire _w19920_ ;
	wire _w19921_ ;
	wire _w19922_ ;
	wire _w19923_ ;
	wire _w19924_ ;
	wire _w19925_ ;
	wire _w19926_ ;
	wire _w19927_ ;
	wire _w19928_ ;
	wire _w19929_ ;
	wire _w19930_ ;
	wire _w19931_ ;
	wire _w19932_ ;
	wire _w19933_ ;
	wire _w19934_ ;
	wire _w19935_ ;
	wire _w19936_ ;
	wire _w19937_ ;
	wire _w19938_ ;
	wire _w19939_ ;
	wire _w19940_ ;
	wire _w19941_ ;
	wire _w19942_ ;
	wire _w19943_ ;
	wire _w19944_ ;
	wire _w19945_ ;
	wire _w19946_ ;
	wire _w19947_ ;
	wire _w19948_ ;
	wire _w19949_ ;
	wire _w19950_ ;
	wire _w19951_ ;
	wire _w19952_ ;
	wire _w19953_ ;
	wire _w19954_ ;
	wire _w19955_ ;
	wire _w19956_ ;
	wire _w19957_ ;
	wire _w19958_ ;
	wire _w19959_ ;
	wire _w19960_ ;
	wire _w19961_ ;
	wire _w19962_ ;
	wire _w19963_ ;
	wire _w19964_ ;
	wire _w19965_ ;
	wire _w19966_ ;
	wire _w19967_ ;
	wire _w19968_ ;
	wire _w19969_ ;
	wire _w19970_ ;
	wire _w19971_ ;
	wire _w19972_ ;
	wire _w19973_ ;
	wire _w19974_ ;
	wire _w19975_ ;
	wire _w19976_ ;
	wire _w19977_ ;
	wire _w19978_ ;
	wire _w19979_ ;
	wire _w19980_ ;
	wire _w19981_ ;
	wire _w19982_ ;
	wire _w19983_ ;
	wire _w19984_ ;
	wire _w19985_ ;
	wire _w19986_ ;
	wire _w19987_ ;
	wire _w19988_ ;
	wire _w19989_ ;
	wire _w19990_ ;
	wire _w19991_ ;
	wire _w19992_ ;
	wire _w19993_ ;
	wire _w19994_ ;
	wire _w19995_ ;
	wire _w19996_ ;
	wire _w19997_ ;
	wire _w19998_ ;
	wire _w19999_ ;
	wire _w20000_ ;
	wire _w20001_ ;
	wire _w20002_ ;
	wire _w20003_ ;
	wire _w20004_ ;
	wire _w20005_ ;
	wire _w20006_ ;
	wire _w20007_ ;
	wire _w20008_ ;
	wire _w20009_ ;
	wire _w20010_ ;
	wire _w20011_ ;
	wire _w20012_ ;
	wire _w20013_ ;
	wire _w20014_ ;
	wire _w20015_ ;
	wire _w20016_ ;
	wire _w20017_ ;
	wire _w20018_ ;
	wire _w20019_ ;
	wire _w20020_ ;
	wire _w20021_ ;
	wire _w20022_ ;
	wire _w20023_ ;
	wire _w20024_ ;
	wire _w20025_ ;
	wire _w20026_ ;
	wire _w20027_ ;
	wire _w20028_ ;
	wire _w20029_ ;
	wire _w20030_ ;
	wire _w20031_ ;
	wire _w20032_ ;
	wire _w20033_ ;
	wire _w20034_ ;
	wire _w20035_ ;
	wire _w20036_ ;
	wire _w20037_ ;
	wire _w20038_ ;
	wire _w20039_ ;
	wire _w20040_ ;
	wire _w20041_ ;
	wire _w20042_ ;
	wire _w20043_ ;
	wire _w20044_ ;
	wire _w20045_ ;
	wire _w20046_ ;
	wire _w20047_ ;
	wire _w20048_ ;
	wire _w20049_ ;
	wire _w20050_ ;
	wire _w20051_ ;
	wire _w20052_ ;
	wire _w20053_ ;
	wire _w20054_ ;
	wire _w20055_ ;
	wire _w20056_ ;
	wire _w20057_ ;
	wire _w20058_ ;
	wire _w20059_ ;
	wire _w20060_ ;
	wire _w20061_ ;
	wire _w20062_ ;
	wire _w20063_ ;
	wire _w20064_ ;
	wire _w20065_ ;
	wire _w20066_ ;
	wire _w20067_ ;
	wire _w20068_ ;
	wire _w20069_ ;
	wire _w20070_ ;
	wire _w20071_ ;
	wire _w20072_ ;
	wire _w20073_ ;
	wire _w20074_ ;
	wire _w20075_ ;
	wire _w20076_ ;
	wire _w20077_ ;
	wire _w20078_ ;
	wire _w20079_ ;
	wire _w20080_ ;
	wire _w20081_ ;
	wire _w20082_ ;
	wire _w20083_ ;
	wire _w20084_ ;
	wire _w20085_ ;
	wire _w20086_ ;
	wire _w20087_ ;
	wire _w20088_ ;
	wire _w20089_ ;
	wire _w20090_ ;
	wire _w20091_ ;
	wire _w20092_ ;
	wire _w20093_ ;
	wire _w20094_ ;
	wire _w20095_ ;
	wire _w20096_ ;
	wire _w20097_ ;
	wire _w20098_ ;
	wire _w20099_ ;
	wire _w20100_ ;
	wire _w20101_ ;
	wire _w20102_ ;
	wire _w20103_ ;
	wire _w20104_ ;
	wire _w20105_ ;
	wire _w20106_ ;
	wire _w20107_ ;
	wire _w20108_ ;
	wire _w20109_ ;
	wire _w20110_ ;
	wire _w20111_ ;
	wire _w20112_ ;
	wire _w20113_ ;
	wire _w20114_ ;
	wire _w20115_ ;
	wire _w20116_ ;
	wire _w20117_ ;
	wire _w20118_ ;
	wire _w20119_ ;
	wire _w20120_ ;
	wire _w20121_ ;
	wire _w20122_ ;
	wire _w20123_ ;
	wire _w20124_ ;
	wire _w20125_ ;
	wire _w20126_ ;
	wire _w20127_ ;
	wire _w20128_ ;
	wire _w20129_ ;
	wire _w20130_ ;
	wire _w20131_ ;
	wire _w20132_ ;
	wire _w20133_ ;
	wire _w20134_ ;
	wire _w20135_ ;
	wire _w20136_ ;
	wire _w20137_ ;
	wire _w20138_ ;
	wire _w20139_ ;
	wire _w20140_ ;
	wire _w20141_ ;
	wire _w20142_ ;
	wire _w20143_ ;
	wire _w20144_ ;
	wire _w20145_ ;
	wire _w20146_ ;
	wire _w20147_ ;
	wire _w20148_ ;
	wire _w20149_ ;
	wire _w20150_ ;
	wire _w20151_ ;
	wire _w20152_ ;
	wire _w20153_ ;
	wire _w20154_ ;
	wire _w20155_ ;
	wire _w20156_ ;
	wire _w20157_ ;
	wire _w20158_ ;
	wire _w20159_ ;
	wire _w20160_ ;
	wire _w20161_ ;
	wire _w20162_ ;
	wire _w20163_ ;
	wire _w20164_ ;
	wire _w20165_ ;
	wire _w20166_ ;
	wire _w20167_ ;
	wire _w20168_ ;
	wire _w20169_ ;
	wire _w20170_ ;
	wire _w20171_ ;
	wire _w20172_ ;
	wire _w20173_ ;
	wire _w20174_ ;
	wire _w20175_ ;
	wire _w20176_ ;
	wire _w20177_ ;
	wire _w20178_ ;
	wire _w20179_ ;
	wire _w20180_ ;
	wire _w20181_ ;
	wire _w20182_ ;
	wire _w20183_ ;
	wire _w20184_ ;
	wire _w20185_ ;
	wire _w20186_ ;
	wire _w20187_ ;
	wire _w20188_ ;
	wire _w20189_ ;
	wire _w20190_ ;
	wire _w20191_ ;
	wire _w20192_ ;
	wire _w20193_ ;
	wire _w20194_ ;
	wire _w20195_ ;
	wire _w20196_ ;
	wire _w20197_ ;
	wire _w20198_ ;
	wire _w20199_ ;
	wire _w20200_ ;
	wire _w20201_ ;
	wire _w20202_ ;
	wire _w20203_ ;
	wire _w20204_ ;
	wire _w20205_ ;
	wire _w20206_ ;
	wire _w20207_ ;
	wire _w20208_ ;
	wire _w20209_ ;
	wire _w20210_ ;
	wire _w20211_ ;
	wire _w20212_ ;
	wire _w20213_ ;
	wire _w20214_ ;
	wire _w20215_ ;
	wire _w20216_ ;
	wire _w20217_ ;
	wire _w20218_ ;
	wire _w20219_ ;
	wire _w20220_ ;
	wire _w20221_ ;
	wire _w20222_ ;
	wire _w20223_ ;
	wire _w20224_ ;
	wire _w20225_ ;
	wire _w20226_ ;
	wire _w20227_ ;
	wire _w20228_ ;
	wire _w20229_ ;
	wire _w20230_ ;
	wire _w20231_ ;
	wire _w20232_ ;
	wire _w20233_ ;
	wire _w20234_ ;
	wire _w20235_ ;
	wire _w20236_ ;
	wire _w20237_ ;
	wire _w20238_ ;
	wire _w20239_ ;
	wire _w20240_ ;
	wire _w20241_ ;
	wire _w20242_ ;
	wire _w20243_ ;
	wire _w20244_ ;
	wire _w20245_ ;
	wire _w20246_ ;
	wire _w20247_ ;
	wire _w20248_ ;
	wire _w20249_ ;
	wire _w20250_ ;
	wire _w20251_ ;
	wire _w20252_ ;
	wire _w20253_ ;
	wire _w20254_ ;
	wire _w20255_ ;
	wire _w20256_ ;
	wire _w20257_ ;
	wire _w20258_ ;
	wire _w20259_ ;
	wire _w20260_ ;
	wire _w20261_ ;
	wire _w20262_ ;
	wire _w20263_ ;
	wire _w20264_ ;
	wire _w20265_ ;
	wire _w20266_ ;
	wire _w20267_ ;
	wire _w20268_ ;
	wire _w20269_ ;
	wire _w20270_ ;
	wire _w20271_ ;
	wire _w20272_ ;
	wire _w20273_ ;
	wire _w20274_ ;
	wire _w20275_ ;
	wire _w20276_ ;
	wire _w20277_ ;
	wire _w20278_ ;
	wire _w20279_ ;
	wire _w20280_ ;
	wire _w20281_ ;
	wire _w20282_ ;
	wire _w20283_ ;
	wire _w20284_ ;
	wire _w20285_ ;
	wire _w20286_ ;
	wire _w20287_ ;
	wire _w20288_ ;
	wire _w20289_ ;
	wire _w20290_ ;
	wire _w20291_ ;
	wire _w20292_ ;
	wire _w20293_ ;
	wire _w20294_ ;
	wire _w20295_ ;
	wire _w20296_ ;
	wire _w20297_ ;
	wire _w20298_ ;
	wire _w20299_ ;
	wire _w20300_ ;
	wire _w20301_ ;
	wire _w20302_ ;
	wire _w20303_ ;
	wire _w20304_ ;
	wire _w20305_ ;
	wire _w20306_ ;
	wire _w20307_ ;
	wire _w20308_ ;
	wire _w20309_ ;
	wire _w20310_ ;
	wire _w20311_ ;
	wire _w20312_ ;
	wire _w20313_ ;
	wire _w20314_ ;
	wire _w20315_ ;
	wire _w20316_ ;
	wire _w20317_ ;
	wire _w20318_ ;
	wire _w20319_ ;
	wire _w20320_ ;
	wire _w20321_ ;
	wire _w20322_ ;
	wire _w20323_ ;
	wire _w20324_ ;
	wire _w20325_ ;
	wire _w20326_ ;
	wire _w20327_ ;
	wire _w20328_ ;
	wire _w20329_ ;
	wire _w20330_ ;
	wire _w20331_ ;
	wire _w20332_ ;
	wire _w20333_ ;
	wire _w20334_ ;
	wire _w20335_ ;
	wire _w20336_ ;
	wire _w20337_ ;
	wire _w20338_ ;
	wire _w20339_ ;
	wire _w20340_ ;
	wire _w20341_ ;
	wire _w20342_ ;
	wire _w20343_ ;
	wire _w20344_ ;
	wire _w20345_ ;
	wire _w20346_ ;
	wire _w20347_ ;
	wire _w20348_ ;
	wire _w20349_ ;
	wire _w20350_ ;
	wire _w20351_ ;
	wire _w20352_ ;
	wire _w20353_ ;
	wire _w20354_ ;
	wire _w20355_ ;
	wire _w20356_ ;
	wire _w20357_ ;
	wire _w20358_ ;
	wire _w20359_ ;
	wire _w20360_ ;
	wire _w20361_ ;
	wire _w20362_ ;
	wire _w20363_ ;
	wire _w20364_ ;
	wire _w20365_ ;
	wire _w20366_ ;
	wire _w20367_ ;
	wire _w20368_ ;
	wire _w20369_ ;
	wire _w20370_ ;
	wire _w20371_ ;
	wire _w20372_ ;
	wire _w20373_ ;
	wire _w20374_ ;
	wire _w20375_ ;
	wire _w20376_ ;
	wire _w20377_ ;
	wire _w20378_ ;
	wire _w20379_ ;
	wire _w20380_ ;
	wire _w20381_ ;
	wire _w20382_ ;
	wire _w20383_ ;
	wire _w20384_ ;
	wire _w20385_ ;
	wire _w20386_ ;
	wire _w20387_ ;
	wire _w20388_ ;
	wire _w20389_ ;
	wire _w20390_ ;
	wire _w20391_ ;
	wire _w20392_ ;
	wire _w20393_ ;
	wire _w20394_ ;
	wire _w20395_ ;
	wire _w20396_ ;
	wire _w20397_ ;
	wire _w20398_ ;
	wire _w20399_ ;
	wire _w20400_ ;
	wire _w20401_ ;
	wire _w20402_ ;
	wire _w20403_ ;
	wire _w20404_ ;
	wire _w20405_ ;
	wire _w20406_ ;
	wire _w20407_ ;
	wire _w20408_ ;
	wire _w20409_ ;
	wire _w20410_ ;
	wire _w20411_ ;
	wire _w20412_ ;
	wire _w20413_ ;
	wire _w20414_ ;
	wire _w20415_ ;
	wire _w20416_ ;
	wire _w20417_ ;
	wire _w20418_ ;
	wire _w20419_ ;
	wire _w20420_ ;
	wire _w20421_ ;
	wire _w20422_ ;
	wire _w20423_ ;
	wire _w20424_ ;
	wire _w20425_ ;
	wire _w20426_ ;
	wire _w20427_ ;
	wire _w20428_ ;
	wire _w20429_ ;
	wire _w20430_ ;
	wire _w20431_ ;
	wire _w20432_ ;
	wire _w20433_ ;
	wire _w20434_ ;
	wire _w20435_ ;
	wire _w20436_ ;
	wire _w20437_ ;
	wire _w20438_ ;
	wire _w20439_ ;
	wire _w20440_ ;
	wire _w20441_ ;
	wire _w20442_ ;
	wire _w20443_ ;
	wire _w20444_ ;
	wire _w20445_ ;
	wire _w20446_ ;
	wire _w20447_ ;
	wire _w20448_ ;
	wire _w20449_ ;
	wire _w20450_ ;
	wire _w20451_ ;
	wire _w20452_ ;
	wire _w20453_ ;
	wire _w20454_ ;
	wire _w20455_ ;
	wire _w20456_ ;
	wire _w20457_ ;
	wire _w20458_ ;
	wire _w20459_ ;
	wire _w20460_ ;
	wire _w20461_ ;
	wire _w20462_ ;
	wire _w20463_ ;
	wire _w20464_ ;
	wire _w20465_ ;
	wire _w20466_ ;
	wire _w20467_ ;
	wire _w20468_ ;
	wire _w20469_ ;
	wire _w20470_ ;
	wire _w20471_ ;
	wire _w20472_ ;
	wire _w20473_ ;
	wire _w20474_ ;
	wire _w20475_ ;
	wire _w20476_ ;
	wire _w20477_ ;
	wire _w20478_ ;
	wire _w20479_ ;
	wire _w20480_ ;
	wire _w20481_ ;
	wire _w20482_ ;
	wire _w20483_ ;
	wire _w20484_ ;
	wire _w20485_ ;
	wire _w20486_ ;
	wire _w20487_ ;
	wire _w20488_ ;
	wire _w20489_ ;
	wire _w20490_ ;
	wire _w20491_ ;
	wire _w20492_ ;
	wire _w20493_ ;
	wire _w20494_ ;
	wire _w20495_ ;
	wire _w20496_ ;
	wire _w20497_ ;
	wire _w20498_ ;
	wire _w20499_ ;
	wire _w20500_ ;
	wire _w20501_ ;
	wire _w20502_ ;
	wire _w20503_ ;
	wire _w20504_ ;
	wire _w20505_ ;
	wire _w20506_ ;
	wire _w20507_ ;
	wire _w20508_ ;
	wire _w20509_ ;
	wire _w20510_ ;
	wire _w20511_ ;
	wire _w20512_ ;
	wire _w20513_ ;
	wire _w20514_ ;
	wire _w20515_ ;
	wire _w20516_ ;
	wire _w20517_ ;
	wire _w20518_ ;
	wire _w20519_ ;
	wire _w20520_ ;
	wire _w20521_ ;
	wire _w20522_ ;
	wire _w20523_ ;
	wire _w20524_ ;
	wire _w20525_ ;
	wire _w20526_ ;
	wire _w20527_ ;
	wire _w20528_ ;
	wire _w20529_ ;
	wire _w20530_ ;
	wire _w20531_ ;
	wire _w20532_ ;
	wire _w20533_ ;
	wire _w20534_ ;
	wire _w20535_ ;
	wire _w20536_ ;
	wire _w20537_ ;
	wire _w20538_ ;
	wire _w20539_ ;
	wire _w20540_ ;
	wire _w20541_ ;
	wire _w20542_ ;
	wire _w20543_ ;
	wire _w20544_ ;
	wire _w20545_ ;
	wire _w20546_ ;
	wire _w20547_ ;
	wire _w20548_ ;
	wire _w20549_ ;
	wire _w20550_ ;
	wire _w20551_ ;
	wire _w20552_ ;
	wire _w20553_ ;
	wire _w20554_ ;
	wire _w20555_ ;
	wire _w20556_ ;
	wire _w20557_ ;
	wire _w20558_ ;
	wire _w20559_ ;
	wire _w20560_ ;
	wire _w20561_ ;
	wire _w20562_ ;
	wire _w20563_ ;
	wire _w20564_ ;
	wire _w20565_ ;
	wire _w20566_ ;
	wire _w20567_ ;
	wire _w20568_ ;
	wire _w20569_ ;
	wire _w20570_ ;
	wire _w20571_ ;
	wire _w20572_ ;
	wire _w20573_ ;
	wire _w20574_ ;
	wire _w20575_ ;
	wire _w20576_ ;
	wire _w20577_ ;
	wire _w20578_ ;
	wire _w20579_ ;
	wire _w20580_ ;
	wire _w20581_ ;
	wire _w20582_ ;
	wire _w20583_ ;
	wire _w20584_ ;
	wire _w20585_ ;
	wire _w20586_ ;
	wire _w20587_ ;
	wire _w20588_ ;
	wire _w20589_ ;
	wire _w20590_ ;
	wire _w20591_ ;
	wire _w20592_ ;
	wire _w20593_ ;
	wire _w20594_ ;
	wire _w20595_ ;
	wire _w20596_ ;
	wire _w20597_ ;
	wire _w20598_ ;
	wire _w20599_ ;
	wire _w20600_ ;
	wire _w20601_ ;
	wire _w20602_ ;
	wire _w20603_ ;
	wire _w20604_ ;
	wire _w20605_ ;
	wire _w20606_ ;
	wire _w20607_ ;
	wire _w20608_ ;
	wire _w20609_ ;
	wire _w20610_ ;
	wire _w20611_ ;
	wire _w20612_ ;
	wire _w20613_ ;
	wire _w20614_ ;
	wire _w20615_ ;
	wire _w20616_ ;
	wire _w20617_ ;
	wire _w20618_ ;
	wire _w20619_ ;
	wire _w20620_ ;
	wire _w20621_ ;
	wire _w20622_ ;
	wire _w20623_ ;
	wire _w20624_ ;
	wire _w20625_ ;
	wire _w20626_ ;
	wire _w20627_ ;
	wire _w20628_ ;
	wire _w20629_ ;
	wire _w20630_ ;
	wire _w20631_ ;
	wire _w20632_ ;
	wire _w20633_ ;
	wire _w20634_ ;
	wire _w20635_ ;
	wire _w20636_ ;
	wire _w20637_ ;
	wire _w20638_ ;
	wire _w20639_ ;
	wire _w20640_ ;
	wire _w20641_ ;
	wire _w20642_ ;
	wire _w20643_ ;
	wire _w20644_ ;
	wire _w20645_ ;
	wire _w20646_ ;
	wire _w20647_ ;
	wire _w20648_ ;
	wire _w20649_ ;
	wire _w20650_ ;
	wire _w20651_ ;
	wire _w20652_ ;
	wire _w20653_ ;
	wire _w20654_ ;
	wire _w20655_ ;
	wire _w20656_ ;
	wire _w20657_ ;
	wire _w20658_ ;
	wire _w20659_ ;
	wire _w20660_ ;
	wire _w20661_ ;
	wire _w20662_ ;
	wire _w20663_ ;
	wire _w20664_ ;
	wire _w20665_ ;
	wire _w20666_ ;
	wire _w20667_ ;
	wire _w20668_ ;
	wire _w20669_ ;
	wire _w20670_ ;
	wire _w20671_ ;
	wire _w20672_ ;
	wire _w20673_ ;
	wire _w20674_ ;
	wire _w20675_ ;
	wire _w20676_ ;
	wire _w20677_ ;
	wire _w20678_ ;
	wire _w20679_ ;
	wire _w20680_ ;
	wire _w20681_ ;
	wire _w20682_ ;
	wire _w20683_ ;
	wire _w20684_ ;
	wire _w20685_ ;
	wire _w20686_ ;
	wire _w20687_ ;
	wire _w20688_ ;
	wire _w20689_ ;
	wire _w20690_ ;
	wire _w20691_ ;
	wire _w20692_ ;
	wire _w20693_ ;
	wire _w20694_ ;
	wire _w20695_ ;
	wire _w20696_ ;
	wire _w20697_ ;
	wire _w20698_ ;
	wire _w20699_ ;
	wire _w20700_ ;
	wire _w20701_ ;
	wire _w20702_ ;
	wire _w20703_ ;
	wire _w20704_ ;
	wire _w20705_ ;
	wire _w20706_ ;
	wire _w20707_ ;
	wire _w20708_ ;
	wire _w20709_ ;
	wire _w20710_ ;
	wire _w20711_ ;
	wire _w20712_ ;
	wire _w20713_ ;
	wire _w20714_ ;
	wire _w20715_ ;
	wire _w20716_ ;
	wire _w20717_ ;
	wire _w20718_ ;
	wire _w20719_ ;
	wire _w20720_ ;
	wire _w20721_ ;
	wire _w20722_ ;
	wire _w20723_ ;
	wire _w20724_ ;
	wire _w20725_ ;
	wire _w20726_ ;
	wire _w20727_ ;
	wire _w20728_ ;
	wire _w20729_ ;
	wire _w20730_ ;
	wire _w20731_ ;
	wire _w20732_ ;
	wire _w20733_ ;
	wire _w20734_ ;
	wire _w20735_ ;
	wire _w20736_ ;
	wire _w20737_ ;
	wire _w20738_ ;
	wire _w20739_ ;
	wire _w20740_ ;
	wire _w20741_ ;
	wire _w20742_ ;
	wire _w20743_ ;
	wire _w20744_ ;
	wire _w20745_ ;
	wire _w20746_ ;
	wire _w20747_ ;
	wire _w20748_ ;
	wire _w20749_ ;
	wire _w20750_ ;
	wire _w20751_ ;
	wire _w20752_ ;
	wire _w20753_ ;
	wire _w20754_ ;
	wire _w20755_ ;
	wire _w20756_ ;
	wire _w20757_ ;
	wire _w20758_ ;
	wire _w20759_ ;
	wire _w20760_ ;
	wire _w20761_ ;
	wire _w20762_ ;
	wire _w20763_ ;
	wire _w20764_ ;
	wire _w20765_ ;
	wire _w20766_ ;
	wire _w20767_ ;
	wire _w20768_ ;
	wire _w20769_ ;
	wire _w20770_ ;
	wire _w20771_ ;
	wire _w20772_ ;
	wire _w20773_ ;
	wire _w20774_ ;
	wire _w20775_ ;
	wire _w20776_ ;
	wire _w20777_ ;
	wire _w20778_ ;
	wire _w20779_ ;
	wire _w20780_ ;
	wire _w20781_ ;
	wire _w20782_ ;
	wire _w20783_ ;
	wire _w20784_ ;
	wire _w20785_ ;
	wire _w20786_ ;
	wire _w20787_ ;
	wire _w20788_ ;
	wire _w20789_ ;
	wire _w20790_ ;
	wire _w20791_ ;
	wire _w20792_ ;
	wire _w20793_ ;
	wire _w20794_ ;
	wire _w20795_ ;
	wire _w20796_ ;
	wire _w20797_ ;
	wire _w20798_ ;
	wire _w20799_ ;
	wire _w20800_ ;
	wire _w20801_ ;
	wire _w20802_ ;
	wire _w20803_ ;
	wire _w20804_ ;
	wire _w20805_ ;
	wire _w20806_ ;
	wire _w20807_ ;
	wire _w20808_ ;
	wire _w20809_ ;
	wire _w20810_ ;
	wire _w20811_ ;
	wire _w20812_ ;
	wire _w20813_ ;
	wire _w20814_ ;
	wire _w20815_ ;
	wire _w20816_ ;
	wire _w20817_ ;
	wire _w20818_ ;
	wire _w20819_ ;
	wire _w20820_ ;
	wire _w20821_ ;
	wire _w20822_ ;
	wire _w20823_ ;
	wire _w20824_ ;
	wire _w20825_ ;
	wire _w20826_ ;
	wire _w20827_ ;
	wire _w20828_ ;
	wire _w20829_ ;
	wire _w20830_ ;
	wire _w20831_ ;
	wire _w20832_ ;
	wire _w20833_ ;
	wire _w20834_ ;
	wire _w20835_ ;
	wire _w20836_ ;
	wire _w20837_ ;
	wire _w20838_ ;
	wire _w20839_ ;
	wire _w20840_ ;
	wire _w20841_ ;
	wire _w20842_ ;
	wire _w20843_ ;
	wire _w20844_ ;
	wire _w20845_ ;
	wire _w20846_ ;
	wire _w20847_ ;
	wire _w20848_ ;
	wire _w20849_ ;
	wire _w20850_ ;
	wire _w20851_ ;
	wire _w20852_ ;
	wire _w20853_ ;
	wire _w20854_ ;
	wire _w20855_ ;
	wire _w20856_ ;
	wire _w20857_ ;
	wire _w20858_ ;
	wire _w20859_ ;
	wire _w20860_ ;
	wire _w20861_ ;
	wire _w20862_ ;
	wire _w20863_ ;
	wire _w20864_ ;
	wire _w20865_ ;
	wire _w20866_ ;
	wire _w20867_ ;
	wire _w20868_ ;
	wire _w20869_ ;
	wire _w20870_ ;
	wire _w20871_ ;
	wire _w20872_ ;
	wire _w20873_ ;
	wire _w20874_ ;
	wire _w20875_ ;
	wire _w20876_ ;
	wire _w20877_ ;
	wire _w20878_ ;
	wire _w20879_ ;
	wire _w20880_ ;
	wire _w20881_ ;
	wire _w20882_ ;
	wire _w20883_ ;
	wire _w20884_ ;
	wire _w20885_ ;
	wire _w20886_ ;
	wire _w20887_ ;
	wire _w20888_ ;
	wire _w20889_ ;
	wire _w20890_ ;
	wire _w20891_ ;
	wire _w20892_ ;
	wire _w20893_ ;
	wire _w20894_ ;
	wire _w20895_ ;
	wire _w20896_ ;
	wire _w20897_ ;
	wire _w20898_ ;
	wire _w20899_ ;
	wire _w20900_ ;
	wire _w20901_ ;
	wire _w20902_ ;
	wire _w20903_ ;
	wire _w20904_ ;
	wire _w20905_ ;
	wire _w20906_ ;
	wire _w20907_ ;
	wire _w20908_ ;
	wire _w20909_ ;
	wire _w20910_ ;
	wire _w20911_ ;
	wire _w20912_ ;
	wire _w20913_ ;
	wire _w20914_ ;
	wire _w20915_ ;
	wire _w20916_ ;
	wire _w20917_ ;
	wire _w20918_ ;
	wire _w20919_ ;
	wire _w20920_ ;
	wire _w20921_ ;
	wire _w20922_ ;
	wire _w20923_ ;
	wire _w20924_ ;
	wire _w20925_ ;
	wire _w20926_ ;
	wire _w20927_ ;
	wire _w20928_ ;
	wire _w20929_ ;
	wire _w20930_ ;
	wire _w20931_ ;
	wire _w20932_ ;
	wire _w20933_ ;
	wire _w20934_ ;
	wire _w20935_ ;
	wire _w20936_ ;
	wire _w20937_ ;
	wire _w20938_ ;
	wire _w20939_ ;
	wire _w20940_ ;
	wire _w20941_ ;
	wire _w20942_ ;
	wire _w20943_ ;
	wire _w20944_ ;
	wire _w20945_ ;
	wire _w20946_ ;
	wire _w20947_ ;
	wire _w20948_ ;
	wire _w20949_ ;
	wire _w20950_ ;
	wire _w20951_ ;
	wire _w20952_ ;
	wire _w20953_ ;
	wire _w20954_ ;
	wire _w20955_ ;
	wire _w20956_ ;
	wire _w20957_ ;
	wire _w20958_ ;
	wire _w20959_ ;
	wire _w20960_ ;
	wire _w20961_ ;
	wire _w20962_ ;
	wire _w20963_ ;
	wire _w20964_ ;
	wire _w20965_ ;
	wire _w20966_ ;
	wire _w20967_ ;
	wire _w20968_ ;
	wire _w20969_ ;
	wire _w20970_ ;
	wire _w20971_ ;
	wire _w20972_ ;
	wire _w20973_ ;
	wire _w20974_ ;
	wire _w20975_ ;
	wire _w20976_ ;
	wire _w20977_ ;
	wire _w20978_ ;
	wire _w20979_ ;
	wire _w20980_ ;
	wire _w20981_ ;
	wire _w20982_ ;
	wire _w20983_ ;
	wire _w20984_ ;
	wire _w20985_ ;
	wire _w20986_ ;
	wire _w20987_ ;
	wire _w20988_ ;
	wire _w20989_ ;
	wire _w20990_ ;
	wire _w20991_ ;
	wire _w20992_ ;
	wire _w20993_ ;
	wire _w20994_ ;
	wire _w20995_ ;
	wire _w20996_ ;
	wire _w20997_ ;
	wire _w20998_ ;
	wire _w20999_ ;
	wire _w21000_ ;
	wire _w21001_ ;
	wire _w21002_ ;
	wire _w21003_ ;
	wire _w21004_ ;
	wire _w21005_ ;
	wire _w21006_ ;
	wire _w21007_ ;
	wire _w21008_ ;
	wire _w21009_ ;
	wire _w21010_ ;
	wire _w21011_ ;
	wire _w21012_ ;
	wire _w21013_ ;
	wire _w21014_ ;
	wire _w21015_ ;
	wire _w21016_ ;
	wire _w21017_ ;
	wire _w21018_ ;
	wire _w21019_ ;
	wire _w21020_ ;
	wire _w21021_ ;
	wire _w21022_ ;
	wire _w21023_ ;
	wire _w21024_ ;
	wire _w21025_ ;
	wire _w21026_ ;
	wire _w21027_ ;
	wire _w21028_ ;
	wire _w21029_ ;
	wire _w21030_ ;
	wire _w21031_ ;
	wire _w21032_ ;
	wire _w21033_ ;
	wire _w21034_ ;
	wire _w21035_ ;
	wire _w21036_ ;
	wire _w21037_ ;
	wire _w21038_ ;
	wire _w21039_ ;
	wire _w21040_ ;
	wire _w21041_ ;
	wire _w21042_ ;
	wire _w21043_ ;
	wire _w21044_ ;
	wire _w21045_ ;
	wire _w21046_ ;
	wire _w21047_ ;
	wire _w21048_ ;
	wire _w21049_ ;
	wire _w21050_ ;
	wire _w21051_ ;
	wire _w21052_ ;
	wire _w21053_ ;
	wire _w21054_ ;
	wire _w21055_ ;
	wire _w21056_ ;
	wire _w21057_ ;
	wire _w21058_ ;
	wire _w21059_ ;
	wire _w21060_ ;
	wire _w21061_ ;
	wire _w21062_ ;
	wire _w21063_ ;
	wire _w21064_ ;
	wire _w21065_ ;
	wire _w21066_ ;
	wire _w21067_ ;
	wire _w21068_ ;
	wire _w21069_ ;
	wire _w21070_ ;
	wire _w21071_ ;
	wire _w21072_ ;
	wire _w21073_ ;
	wire _w21074_ ;
	wire _w21075_ ;
	wire _w21076_ ;
	wire _w21077_ ;
	wire _w21078_ ;
	wire _w21079_ ;
	wire _w21080_ ;
	wire _w21081_ ;
	wire _w21082_ ;
	wire _w21083_ ;
	wire _w21084_ ;
	wire _w21085_ ;
	wire _w21086_ ;
	wire _w21087_ ;
	wire _w21088_ ;
	wire _w21089_ ;
	wire _w21090_ ;
	wire _w21091_ ;
	wire _w21092_ ;
	wire _w21093_ ;
	wire _w21094_ ;
	wire _w21095_ ;
	wire _w21096_ ;
	wire _w21097_ ;
	wire _w21098_ ;
	wire _w21099_ ;
	wire _w21100_ ;
	wire _w21101_ ;
	wire _w21102_ ;
	wire _w21103_ ;
	wire _w21104_ ;
	wire _w21105_ ;
	wire _w21106_ ;
	wire _w21107_ ;
	wire _w21108_ ;
	wire _w21109_ ;
	wire _w21110_ ;
	wire _w21111_ ;
	wire _w21112_ ;
	wire _w21113_ ;
	wire _w21114_ ;
	wire _w21115_ ;
	wire _w21116_ ;
	wire _w21117_ ;
	wire _w21118_ ;
	wire _w21119_ ;
	wire _w21120_ ;
	wire _w21121_ ;
	wire _w21122_ ;
	wire _w21123_ ;
	wire _w21124_ ;
	wire _w21125_ ;
	wire _w21126_ ;
	wire _w21127_ ;
	wire _w21128_ ;
	wire _w21129_ ;
	wire _w21130_ ;
	wire _w21131_ ;
	wire _w21132_ ;
	wire _w21133_ ;
	wire _w21134_ ;
	wire _w21135_ ;
	wire _w21136_ ;
	wire _w21137_ ;
	wire _w21138_ ;
	wire _w21139_ ;
	wire _w21140_ ;
	wire _w21141_ ;
	wire _w21142_ ;
	wire _w21143_ ;
	wire _w21144_ ;
	wire _w21145_ ;
	wire _w21146_ ;
	wire _w21147_ ;
	wire _w21148_ ;
	wire _w21149_ ;
	wire _w21150_ ;
	wire _w21151_ ;
	wire _w21152_ ;
	wire _w21153_ ;
	wire _w21154_ ;
	wire _w21155_ ;
	wire _w21156_ ;
	wire _w21157_ ;
	wire _w21158_ ;
	wire _w21159_ ;
	wire _w21160_ ;
	wire _w21161_ ;
	wire _w21162_ ;
	wire _w21163_ ;
	wire _w21164_ ;
	wire _w21165_ ;
	wire _w21166_ ;
	wire _w21167_ ;
	wire _w21168_ ;
	wire _w21169_ ;
	wire _w21170_ ;
	wire _w21171_ ;
	wire _w21172_ ;
	wire _w21173_ ;
	wire _w21174_ ;
	wire _w21175_ ;
	wire _w21176_ ;
	wire _w21177_ ;
	wire _w21178_ ;
	wire _w21179_ ;
	wire _w21180_ ;
	wire _w21181_ ;
	wire _w21182_ ;
	wire _w21183_ ;
	wire _w21184_ ;
	wire _w21185_ ;
	wire _w21186_ ;
	wire _w21187_ ;
	wire _w21188_ ;
	wire _w21189_ ;
	wire _w21190_ ;
	wire _w21191_ ;
	wire _w21192_ ;
	wire _w21193_ ;
	wire _w21194_ ;
	wire _w21195_ ;
	wire _w21196_ ;
	wire _w21197_ ;
	wire _w21198_ ;
	wire _w21199_ ;
	wire _w21200_ ;
	wire _w21201_ ;
	wire _w21202_ ;
	wire _w21203_ ;
	wire _w21204_ ;
	wire _w21205_ ;
	wire _w21206_ ;
	wire _w21207_ ;
	wire _w21208_ ;
	wire _w21209_ ;
	wire _w21210_ ;
	wire _w21211_ ;
	wire _w21212_ ;
	wire _w21213_ ;
	wire _w21214_ ;
	wire _w21215_ ;
	wire _w21216_ ;
	wire _w21217_ ;
	wire _w21218_ ;
	wire _w21219_ ;
	wire _w21220_ ;
	wire _w21221_ ;
	wire _w21222_ ;
	wire _w21223_ ;
	wire _w21224_ ;
	wire _w21225_ ;
	wire _w21226_ ;
	wire _w21227_ ;
	wire _w21228_ ;
	wire _w21229_ ;
	wire _w21230_ ;
	wire _w21231_ ;
	wire _w21232_ ;
	wire _w21233_ ;
	wire _w21234_ ;
	wire _w21235_ ;
	wire _w21236_ ;
	wire _w21237_ ;
	wire _w21238_ ;
	wire _w21239_ ;
	wire _w21240_ ;
	wire _w21241_ ;
	wire _w21242_ ;
	wire _w21243_ ;
	wire _w21244_ ;
	wire _w21245_ ;
	wire _w21246_ ;
	wire _w21247_ ;
	wire _w21248_ ;
	wire _w21249_ ;
	wire _w21250_ ;
	wire _w21251_ ;
	wire _w21252_ ;
	wire _w21253_ ;
	wire _w21254_ ;
	wire _w21255_ ;
	wire _w21256_ ;
	wire _w21257_ ;
	wire _w21258_ ;
	wire _w21259_ ;
	wire _w21260_ ;
	wire _w21261_ ;
	wire _w21262_ ;
	wire _w21263_ ;
	wire _w21264_ ;
	wire _w21265_ ;
	wire _w21266_ ;
	wire _w21267_ ;
	wire _w21268_ ;
	wire _w21269_ ;
	wire _w21270_ ;
	wire _w21271_ ;
	wire _w21272_ ;
	wire _w21273_ ;
	wire _w21274_ ;
	wire _w21275_ ;
	wire _w21276_ ;
	wire _w21277_ ;
	wire _w21278_ ;
	wire _w21279_ ;
	wire _w21280_ ;
	wire _w21281_ ;
	wire _w21282_ ;
	wire _w21283_ ;
	wire _w21284_ ;
	wire _w21285_ ;
	wire _w21286_ ;
	wire _w21287_ ;
	wire _w21288_ ;
	wire _w21289_ ;
	wire _w21290_ ;
	wire _w21291_ ;
	wire _w21292_ ;
	wire _w21293_ ;
	wire _w21294_ ;
	wire _w21295_ ;
	wire _w21296_ ;
	wire _w21297_ ;
	wire _w21298_ ;
	wire _w21299_ ;
	wire _w21300_ ;
	wire _w21301_ ;
	wire _w21302_ ;
	wire _w21303_ ;
	wire _w21304_ ;
	wire _w21305_ ;
	wire _w21306_ ;
	wire _w21307_ ;
	wire _w21308_ ;
	wire _w21309_ ;
	wire _w21310_ ;
	wire _w21311_ ;
	wire _w21312_ ;
	wire _w21313_ ;
	wire _w21314_ ;
	wire _w21315_ ;
	wire _w21316_ ;
	wire _w21317_ ;
	wire _w21318_ ;
	wire _w21319_ ;
	wire _w21320_ ;
	wire _w21321_ ;
	wire _w21322_ ;
	wire _w21323_ ;
	wire _w21324_ ;
	wire _w21325_ ;
	wire _w21326_ ;
	wire _w21327_ ;
	wire _w21328_ ;
	wire _w21329_ ;
	wire _w21330_ ;
	wire _w21331_ ;
	wire _w21332_ ;
	wire _w21333_ ;
	wire _w21334_ ;
	wire _w21335_ ;
	wire _w21336_ ;
	wire _w21337_ ;
	wire _w21338_ ;
	wire _w21339_ ;
	wire _w21340_ ;
	wire _w21341_ ;
	wire _w21342_ ;
	wire _w21343_ ;
	wire _w21344_ ;
	wire _w21345_ ;
	wire _w21346_ ;
	wire _w21347_ ;
	wire _w21348_ ;
	wire _w21349_ ;
	wire _w21350_ ;
	wire _w21351_ ;
	wire _w21352_ ;
	wire _w21353_ ;
	wire _w21354_ ;
	wire _w21355_ ;
	wire _w21356_ ;
	wire _w21357_ ;
	wire _w21358_ ;
	wire _w21359_ ;
	wire _w21360_ ;
	wire _w21361_ ;
	wire _w21362_ ;
	wire _w21363_ ;
	wire _w21364_ ;
	wire _w21365_ ;
	wire _w21366_ ;
	wire _w21367_ ;
	wire _w21368_ ;
	wire _w21369_ ;
	wire _w21370_ ;
	wire _w21371_ ;
	wire _w21372_ ;
	wire _w21373_ ;
	wire _w21374_ ;
	wire _w21375_ ;
	wire _w21376_ ;
	wire _w21377_ ;
	wire _w21378_ ;
	wire _w21379_ ;
	wire _w21380_ ;
	wire _w21381_ ;
	wire _w21382_ ;
	wire _w21383_ ;
	wire _w21384_ ;
	wire _w21385_ ;
	wire _w21386_ ;
	wire _w21387_ ;
	wire _w21388_ ;
	wire _w21389_ ;
	wire _w21390_ ;
	wire _w21391_ ;
	wire _w21392_ ;
	wire _w21393_ ;
	wire _w21394_ ;
	wire _w21395_ ;
	wire _w21396_ ;
	wire _w21397_ ;
	wire _w21398_ ;
	wire _w21399_ ;
	wire _w21400_ ;
	wire _w21401_ ;
	wire _w21402_ ;
	wire _w21403_ ;
	wire _w21404_ ;
	wire _w21405_ ;
	wire _w21406_ ;
	wire _w21407_ ;
	wire _w21408_ ;
	wire _w21409_ ;
	wire _w21410_ ;
	wire _w21411_ ;
	wire _w21412_ ;
	wire _w21413_ ;
	wire _w21414_ ;
	wire _w21415_ ;
	wire _w21416_ ;
	wire _w21417_ ;
	wire _w21418_ ;
	wire _w21419_ ;
	wire _w21420_ ;
	wire _w21421_ ;
	wire _w21422_ ;
	wire _w21423_ ;
	wire _w21424_ ;
	wire _w21425_ ;
	wire _w21426_ ;
	wire _w21427_ ;
	wire _w21428_ ;
	wire _w21429_ ;
	wire _w21430_ ;
	wire _w21431_ ;
	wire _w21432_ ;
	wire _w21433_ ;
	wire _w21434_ ;
	wire _w21435_ ;
	wire _w21436_ ;
	wire _w21437_ ;
	wire _w21438_ ;
	wire _w21439_ ;
	wire _w21440_ ;
	wire _w21441_ ;
	wire _w21442_ ;
	wire _w21443_ ;
	wire _w21444_ ;
	wire _w21445_ ;
	wire _w21446_ ;
	wire _w21447_ ;
	wire _w21448_ ;
	wire _w21449_ ;
	wire _w21450_ ;
	wire _w21451_ ;
	wire _w21452_ ;
	wire _w21453_ ;
	wire _w21454_ ;
	wire _w21455_ ;
	wire _w21456_ ;
	wire _w21457_ ;
	wire _w21458_ ;
	wire _w21459_ ;
	wire _w21460_ ;
	wire _w21461_ ;
	wire _w21462_ ;
	wire _w21463_ ;
	wire _w21464_ ;
	wire _w21465_ ;
	wire _w21466_ ;
	wire _w21467_ ;
	wire _w21468_ ;
	wire _w21469_ ;
	wire _w21470_ ;
	wire _w21471_ ;
	wire _w21472_ ;
	wire _w21473_ ;
	wire _w21474_ ;
	wire _w21475_ ;
	wire _w21476_ ;
	wire _w21477_ ;
	wire _w21478_ ;
	wire _w21479_ ;
	wire _w21480_ ;
	wire _w21481_ ;
	wire _w21482_ ;
	wire _w21483_ ;
	wire _w21484_ ;
	wire _w21485_ ;
	wire _w21486_ ;
	wire _w21487_ ;
	wire _w21488_ ;
	wire _w21489_ ;
	wire _w21490_ ;
	wire _w21491_ ;
	wire _w21492_ ;
	wire _w21493_ ;
	wire _w21494_ ;
	wire _w21495_ ;
	wire _w21496_ ;
	wire _w21497_ ;
	wire _w21498_ ;
	wire _w21499_ ;
	wire _w21500_ ;
	wire _w21501_ ;
	wire _w21502_ ;
	wire _w21503_ ;
	wire _w21504_ ;
	wire _w21505_ ;
	wire _w21506_ ;
	wire _w21507_ ;
	wire _w21508_ ;
	wire _w21509_ ;
	wire _w21510_ ;
	wire _w21511_ ;
	wire _w21512_ ;
	wire _w21513_ ;
	wire _w21514_ ;
	wire _w21515_ ;
	wire _w21516_ ;
	wire _w21517_ ;
	wire _w21518_ ;
	wire _w21519_ ;
	wire _w21520_ ;
	wire _w21521_ ;
	wire _w21522_ ;
	wire _w21523_ ;
	wire _w21524_ ;
	wire _w21525_ ;
	wire _w21526_ ;
	wire _w21527_ ;
	wire _w21528_ ;
	wire _w21529_ ;
	wire _w21530_ ;
	wire _w21531_ ;
	wire _w21532_ ;
	wire _w21533_ ;
	wire _w21534_ ;
	wire _w21535_ ;
	wire _w21536_ ;
	wire _w21537_ ;
	wire _w21538_ ;
	wire _w21539_ ;
	wire _w21540_ ;
	wire _w21541_ ;
	wire _w21542_ ;
	wire _w21543_ ;
	wire _w21544_ ;
	wire _w21545_ ;
	wire _w21546_ ;
	wire _w21547_ ;
	wire _w21548_ ;
	wire _w21549_ ;
	wire _w21550_ ;
	wire _w21551_ ;
	wire _w21552_ ;
	wire _w21553_ ;
	wire _w21554_ ;
	wire _w21555_ ;
	wire _w21556_ ;
	wire _w21557_ ;
	wire _w21558_ ;
	wire _w21559_ ;
	wire _w21560_ ;
	wire _w21561_ ;
	wire _w21562_ ;
	wire _w21563_ ;
	wire _w21564_ ;
	wire _w21565_ ;
	wire _w21566_ ;
	wire _w21567_ ;
	wire _w21568_ ;
	wire _w21569_ ;
	wire _w21570_ ;
	wire _w21571_ ;
	wire _w21572_ ;
	wire _w21573_ ;
	wire _w21574_ ;
	wire _w21575_ ;
	wire _w21576_ ;
	wire _w21577_ ;
	wire _w21578_ ;
	wire _w21579_ ;
	wire _w21580_ ;
	wire _w21581_ ;
	wire _w21582_ ;
	wire _w21583_ ;
	wire _w21584_ ;
	wire _w21585_ ;
	wire _w21586_ ;
	wire _w21587_ ;
	wire _w21588_ ;
	wire _w21589_ ;
	wire _w21590_ ;
	wire _w21591_ ;
	wire _w21592_ ;
	wire _w21593_ ;
	wire _w21594_ ;
	wire _w21595_ ;
	wire _w21596_ ;
	wire _w21597_ ;
	wire _w21598_ ;
	wire _w21599_ ;
	wire _w21600_ ;
	wire _w21601_ ;
	wire _w21602_ ;
	wire _w21603_ ;
	wire _w21604_ ;
	wire _w21605_ ;
	wire _w21606_ ;
	wire _w21607_ ;
	wire _w21608_ ;
	wire _w21609_ ;
	wire _w21610_ ;
	wire _w21611_ ;
	wire _w21612_ ;
	wire _w21613_ ;
	wire _w21614_ ;
	wire _w21615_ ;
	wire _w21616_ ;
	wire _w21617_ ;
	wire _w21618_ ;
	wire _w21619_ ;
	wire _w21620_ ;
	wire _w21621_ ;
	wire _w21622_ ;
	wire _w21623_ ;
	wire _w21624_ ;
	wire _w21625_ ;
	wire _w21626_ ;
	wire _w21627_ ;
	wire _w21628_ ;
	wire _w21629_ ;
	wire _w21630_ ;
	wire _w21631_ ;
	wire _w21632_ ;
	wire _w21633_ ;
	wire _w21634_ ;
	wire _w21635_ ;
	wire _w21636_ ;
	wire _w21637_ ;
	wire _w21638_ ;
	wire _w21639_ ;
	wire _w21640_ ;
	wire _w21641_ ;
	wire _w21642_ ;
	wire _w21643_ ;
	wire _w21644_ ;
	wire _w21645_ ;
	wire _w21646_ ;
	wire _w21647_ ;
	wire _w21648_ ;
	wire _w21649_ ;
	wire _w21650_ ;
	wire _w21651_ ;
	wire _w21652_ ;
	wire _w21653_ ;
	wire _w21654_ ;
	wire _w21655_ ;
	wire _w21656_ ;
	wire _w21657_ ;
	wire _w21658_ ;
	wire _w21659_ ;
	wire _w21660_ ;
	wire _w21661_ ;
	wire _w21662_ ;
	wire _w21663_ ;
	wire _w21664_ ;
	wire _w21665_ ;
	wire _w21666_ ;
	wire _w21667_ ;
	wire _w21668_ ;
	wire _w21669_ ;
	wire _w21670_ ;
	wire _w21671_ ;
	wire _w21672_ ;
	wire _w21673_ ;
	wire _w21674_ ;
	wire _w21675_ ;
	wire _w21676_ ;
	wire _w21677_ ;
	wire _w21678_ ;
	wire _w21679_ ;
	wire _w21680_ ;
	wire _w21681_ ;
	wire _w21682_ ;
	wire _w21683_ ;
	wire _w21684_ ;
	wire _w21685_ ;
	wire _w21686_ ;
	wire _w21687_ ;
	wire _w21688_ ;
	wire _w21689_ ;
	wire _w21690_ ;
	wire _w21691_ ;
	wire _w21692_ ;
	wire _w21693_ ;
	wire _w21694_ ;
	wire _w21695_ ;
	wire _w21696_ ;
	wire _w21697_ ;
	wire _w21698_ ;
	wire _w21699_ ;
	wire _w21700_ ;
	wire _w21701_ ;
	wire _w21702_ ;
	wire _w21703_ ;
	wire _w21704_ ;
	wire _w21705_ ;
	wire _w21706_ ;
	wire _w21707_ ;
	wire _w21708_ ;
	wire _w21709_ ;
	wire _w21710_ ;
	wire _w21711_ ;
	wire _w21712_ ;
	wire _w21713_ ;
	wire _w21714_ ;
	wire _w21715_ ;
	wire _w21716_ ;
	wire _w21717_ ;
	wire _w21718_ ;
	wire _w21719_ ;
	wire _w21720_ ;
	wire _w21721_ ;
	wire _w21722_ ;
	wire _w21723_ ;
	wire _w21724_ ;
	wire _w21725_ ;
	wire _w21726_ ;
	wire _w21727_ ;
	wire _w21728_ ;
	wire _w21729_ ;
	wire _w21730_ ;
	wire _w21731_ ;
	wire _w21732_ ;
	wire _w21733_ ;
	wire _w21734_ ;
	wire _w21735_ ;
	wire _w21736_ ;
	wire _w21737_ ;
	wire _w21738_ ;
	wire _w21739_ ;
	wire _w21740_ ;
	wire _w21741_ ;
	wire _w21742_ ;
	wire _w21743_ ;
	wire _w21744_ ;
	wire _w21745_ ;
	wire _w21746_ ;
	wire _w21747_ ;
	wire _w21748_ ;
	wire _w21749_ ;
	wire _w21750_ ;
	wire _w21751_ ;
	wire _w21752_ ;
	wire _w21753_ ;
	wire _w21754_ ;
	wire _w21755_ ;
	wire _w21756_ ;
	wire _w21757_ ;
	wire _w21758_ ;
	wire _w21759_ ;
	wire _w21760_ ;
	wire _w21761_ ;
	wire _w21762_ ;
	wire _w21763_ ;
	wire _w21764_ ;
	wire _w21765_ ;
	wire _w21766_ ;
	wire _w21767_ ;
	wire _w21768_ ;
	wire _w21769_ ;
	wire _w21770_ ;
	wire _w21771_ ;
	wire _w21772_ ;
	wire _w21773_ ;
	wire _w21774_ ;
	wire _w21775_ ;
	wire _w21776_ ;
	wire _w21777_ ;
	wire _w21778_ ;
	wire _w21779_ ;
	wire _w21780_ ;
	wire _w21781_ ;
	wire _w21782_ ;
	wire _w21783_ ;
	wire _w21784_ ;
	wire _w21785_ ;
	wire _w21786_ ;
	wire _w21787_ ;
	wire _w21788_ ;
	wire _w21789_ ;
	wire _w21790_ ;
	wire _w21791_ ;
	wire _w21792_ ;
	wire _w21793_ ;
	wire _w21794_ ;
	wire _w21795_ ;
	wire _w21796_ ;
	wire _w21797_ ;
	wire _w21798_ ;
	wire _w21799_ ;
	wire _w21800_ ;
	wire _w21801_ ;
	wire _w21802_ ;
	wire _w21803_ ;
	wire _w21804_ ;
	wire _w21805_ ;
	wire _w21806_ ;
	wire _w21807_ ;
	wire _w21808_ ;
	wire _w21809_ ;
	wire _w21810_ ;
	wire _w21811_ ;
	wire _w21812_ ;
	wire _w21813_ ;
	wire _w21814_ ;
	wire _w21815_ ;
	wire _w21816_ ;
	wire _w21817_ ;
	wire _w21818_ ;
	wire _w21819_ ;
	wire _w21820_ ;
	wire _w21821_ ;
	wire _w21822_ ;
	wire _w21823_ ;
	wire _w21824_ ;
	wire _w21825_ ;
	wire _w21826_ ;
	wire _w21827_ ;
	wire _w21828_ ;
	wire _w21829_ ;
	wire _w21830_ ;
	wire _w21831_ ;
	wire _w21832_ ;
	wire _w21833_ ;
	wire _w21834_ ;
	wire _w21835_ ;
	wire _w21836_ ;
	wire _w21837_ ;
	wire _w21838_ ;
	wire _w21839_ ;
	wire _w21840_ ;
	wire _w21841_ ;
	wire _w21842_ ;
	wire _w21843_ ;
	wire _w21844_ ;
	wire _w21845_ ;
	wire _w21846_ ;
	wire _w21847_ ;
	wire _w21848_ ;
	wire _w21849_ ;
	wire _w21850_ ;
	wire _w21851_ ;
	wire _w21852_ ;
	wire _w21853_ ;
	wire _w21854_ ;
	wire _w21855_ ;
	wire _w21856_ ;
	wire _w21857_ ;
	wire _w21858_ ;
	wire _w21859_ ;
	wire _w21860_ ;
	wire _w21861_ ;
	wire _w21862_ ;
	wire _w21863_ ;
	wire _w21864_ ;
	wire _w21865_ ;
	wire _w21866_ ;
	wire _w21867_ ;
	wire _w21868_ ;
	wire _w21869_ ;
	wire _w21870_ ;
	wire _w21871_ ;
	wire _w21872_ ;
	wire _w21873_ ;
	wire _w21874_ ;
	wire _w21875_ ;
	wire _w21876_ ;
	wire _w21877_ ;
	wire _w21878_ ;
	wire _w21879_ ;
	wire _w21880_ ;
	wire _w21881_ ;
	wire _w21882_ ;
	wire _w21883_ ;
	wire _w21884_ ;
	wire _w21885_ ;
	wire _w21886_ ;
	wire _w21887_ ;
	wire _w21888_ ;
	wire _w21889_ ;
	wire _w21890_ ;
	wire _w21891_ ;
	wire _w21892_ ;
	wire _w21893_ ;
	wire _w21894_ ;
	wire _w21895_ ;
	wire _w21896_ ;
	wire _w21897_ ;
	wire _w21898_ ;
	wire _w21899_ ;
	wire _w21900_ ;
	wire _w21901_ ;
	wire _w21902_ ;
	wire _w21903_ ;
	wire _w21904_ ;
	wire _w21905_ ;
	wire _w21906_ ;
	wire _w21907_ ;
	wire _w21908_ ;
	wire _w21909_ ;
	wire _w21910_ ;
	wire _w21911_ ;
	wire _w21912_ ;
	wire _w21913_ ;
	wire _w21914_ ;
	wire _w21915_ ;
	wire _w21916_ ;
	wire _w21917_ ;
	wire _w21918_ ;
	wire _w21919_ ;
	wire _w21920_ ;
	wire _w21921_ ;
	wire _w21922_ ;
	wire _w21923_ ;
	wire _w21924_ ;
	wire _w21925_ ;
	wire _w21926_ ;
	wire _w21927_ ;
	wire _w21928_ ;
	wire _w21929_ ;
	wire _w21930_ ;
	wire _w21931_ ;
	wire _w21932_ ;
	wire _w21933_ ;
	wire _w21934_ ;
	wire _w21935_ ;
	wire _w21936_ ;
	wire _w21937_ ;
	wire _w21938_ ;
	wire _w21939_ ;
	wire _w21940_ ;
	wire _w21941_ ;
	wire _w21942_ ;
	wire _w21943_ ;
	wire _w21944_ ;
	wire _w21945_ ;
	wire _w21946_ ;
	wire _w21947_ ;
	wire _w21948_ ;
	wire _w21949_ ;
	wire _w21950_ ;
	wire _w21951_ ;
	wire _w21952_ ;
	wire _w21953_ ;
	wire _w21954_ ;
	wire _w21955_ ;
	wire _w21956_ ;
	wire _w21957_ ;
	wire _w21958_ ;
	wire _w21959_ ;
	wire _w21960_ ;
	wire _w21961_ ;
	wire _w21962_ ;
	wire _w21963_ ;
	wire _w21964_ ;
	wire _w21965_ ;
	wire _w21966_ ;
	wire _w21967_ ;
	wire _w21968_ ;
	wire _w21969_ ;
	wire _w21970_ ;
	wire _w21971_ ;
	wire _w21972_ ;
	wire _w21973_ ;
	wire _w21974_ ;
	wire _w21975_ ;
	wire _w21976_ ;
	wire _w21977_ ;
	wire _w21978_ ;
	wire _w21979_ ;
	wire _w21980_ ;
	wire _w21981_ ;
	wire _w21982_ ;
	wire _w21983_ ;
	wire _w21984_ ;
	wire _w21985_ ;
	wire _w21986_ ;
	wire _w21987_ ;
	wire _w21988_ ;
	wire _w21989_ ;
	wire _w21990_ ;
	wire _w21991_ ;
	wire _w21992_ ;
	wire _w21993_ ;
	wire _w21994_ ;
	wire _w21995_ ;
	wire _w21996_ ;
	wire _w21997_ ;
	wire _w21998_ ;
	wire _w21999_ ;
	wire _w22000_ ;
	wire _w22001_ ;
	wire _w22002_ ;
	wire _w22003_ ;
	wire _w22004_ ;
	wire _w22005_ ;
	wire _w22006_ ;
	wire _w22007_ ;
	wire _w22008_ ;
	wire _w22009_ ;
	wire _w22010_ ;
	wire _w22011_ ;
	wire _w22012_ ;
	wire _w22013_ ;
	wire _w22014_ ;
	wire _w22015_ ;
	wire _w22016_ ;
	wire _w22017_ ;
	wire _w22018_ ;
	wire _w22019_ ;
	wire _w22020_ ;
	wire _w22021_ ;
	wire _w22022_ ;
	wire _w22023_ ;
	wire _w22024_ ;
	wire _w22025_ ;
	wire _w22026_ ;
	wire _w22027_ ;
	wire _w22028_ ;
	wire _w22029_ ;
	wire _w22030_ ;
	wire _w22031_ ;
	wire _w22032_ ;
	wire _w22033_ ;
	wire _w22034_ ;
	wire _w22035_ ;
	wire _w22036_ ;
	wire _w22037_ ;
	wire _w22038_ ;
	wire _w22039_ ;
	wire _w22040_ ;
	wire _w22041_ ;
	wire _w22042_ ;
	wire _w22043_ ;
	wire _w22044_ ;
	wire _w22045_ ;
	wire _w22046_ ;
	wire _w22047_ ;
	wire _w22048_ ;
	wire _w22049_ ;
	wire _w22050_ ;
	wire _w22051_ ;
	wire _w22052_ ;
	wire _w22053_ ;
	wire _w22054_ ;
	wire _w22055_ ;
	wire _w22056_ ;
	wire _w22057_ ;
	wire _w22058_ ;
	wire _w22059_ ;
	wire _w22060_ ;
	wire _w22061_ ;
	wire _w22062_ ;
	wire _w22063_ ;
	wire _w22064_ ;
	wire _w22065_ ;
	wire _w22066_ ;
	wire _w22067_ ;
	wire _w22068_ ;
	wire _w22069_ ;
	wire _w22070_ ;
	wire _w22071_ ;
	wire _w22072_ ;
	wire _w22073_ ;
	wire _w22074_ ;
	wire _w22075_ ;
	wire _w22076_ ;
	wire _w22077_ ;
	wire _w22078_ ;
	wire _w22079_ ;
	wire _w22080_ ;
	wire _w22081_ ;
	wire _w22082_ ;
	wire _w22083_ ;
	wire _w22084_ ;
	wire _w22085_ ;
	wire _w22086_ ;
	wire _w22087_ ;
	wire _w22088_ ;
	wire _w22089_ ;
	wire _w22090_ ;
	wire _w22091_ ;
	wire _w22092_ ;
	wire _w22093_ ;
	wire _w22094_ ;
	wire _w22095_ ;
	wire _w22096_ ;
	wire _w22097_ ;
	wire _w22098_ ;
	wire _w22099_ ;
	wire _w22100_ ;
	wire _w22101_ ;
	wire _w22102_ ;
	wire _w22103_ ;
	wire _w22104_ ;
	wire _w22105_ ;
	wire _w22106_ ;
	wire _w22107_ ;
	wire _w22108_ ;
	wire _w22109_ ;
	wire _w22110_ ;
	wire _w22111_ ;
	wire _w22112_ ;
	wire _w22113_ ;
	wire _w22114_ ;
	wire _w22115_ ;
	wire _w22116_ ;
	wire _w22117_ ;
	wire _w22118_ ;
	wire _w22119_ ;
	wire _w22120_ ;
	wire _w22121_ ;
	wire _w22122_ ;
	wire _w22123_ ;
	wire _w22124_ ;
	wire _w22125_ ;
	wire _w22126_ ;
	wire _w22127_ ;
	wire _w22128_ ;
	wire _w22129_ ;
	wire _w22130_ ;
	wire _w22131_ ;
	wire _w22132_ ;
	wire _w22133_ ;
	wire _w22134_ ;
	wire _w22135_ ;
	wire _w22136_ ;
	wire _w22137_ ;
	wire _w22138_ ;
	wire _w22139_ ;
	wire _w22140_ ;
	wire _w22141_ ;
	wire _w22142_ ;
	wire _w22143_ ;
	wire _w22144_ ;
	wire _w22145_ ;
	wire _w22146_ ;
	wire _w22147_ ;
	wire _w22148_ ;
	wire _w22149_ ;
	wire _w22150_ ;
	wire _w22151_ ;
	wire _w22152_ ;
	wire _w22153_ ;
	wire _w22154_ ;
	wire _w22155_ ;
	wire _w22156_ ;
	wire _w22157_ ;
	wire _w22158_ ;
	wire _w22159_ ;
	wire _w22160_ ;
	wire _w22161_ ;
	wire _w22162_ ;
	wire _w22163_ ;
	wire _w22164_ ;
	wire _w22165_ ;
	wire _w22166_ ;
	wire _w22167_ ;
	wire _w22168_ ;
	wire _w22169_ ;
	wire _w22170_ ;
	wire _w22171_ ;
	wire _w22172_ ;
	wire _w22173_ ;
	wire _w22174_ ;
	wire _w22175_ ;
	wire _w22176_ ;
	wire _w22177_ ;
	wire _w22178_ ;
	wire _w22179_ ;
	wire _w22180_ ;
	wire _w22181_ ;
	wire _w22182_ ;
	wire _w22183_ ;
	wire _w22184_ ;
	wire _w22185_ ;
	wire _w22186_ ;
	wire _w22187_ ;
	wire _w22188_ ;
	wire _w22189_ ;
	wire _w22190_ ;
	wire _w22191_ ;
	wire _w22192_ ;
	wire _w22193_ ;
	wire _w22194_ ;
	wire _w22195_ ;
	wire _w22196_ ;
	wire _w22197_ ;
	wire _w22198_ ;
	wire _w22199_ ;
	wire _w22200_ ;
	wire _w22201_ ;
	wire _w22202_ ;
	wire _w22203_ ;
	wire _w22204_ ;
	wire _w22205_ ;
	wire _w22206_ ;
	wire _w22207_ ;
	wire _w22208_ ;
	wire _w22209_ ;
	wire _w22210_ ;
	wire _w22211_ ;
	wire _w22212_ ;
	wire _w22213_ ;
	wire _w22214_ ;
	wire _w22215_ ;
	wire _w22216_ ;
	wire _w22217_ ;
	wire _w22218_ ;
	wire _w22219_ ;
	wire _w22220_ ;
	wire _w22221_ ;
	wire _w22222_ ;
	wire _w22223_ ;
	wire _w22224_ ;
	wire _w22225_ ;
	wire _w22226_ ;
	wire _w22227_ ;
	wire _w22228_ ;
	wire _w22229_ ;
	wire _w22230_ ;
	wire _w22231_ ;
	wire _w22232_ ;
	wire _w22233_ ;
	wire _w22234_ ;
	wire _w22235_ ;
	wire _w22236_ ;
	wire _w22237_ ;
	wire _w22238_ ;
	wire _w22239_ ;
	wire _w22240_ ;
	wire _w22241_ ;
	wire _w22242_ ;
	wire _w22243_ ;
	wire _w22244_ ;
	wire _w22245_ ;
	wire _w22246_ ;
	wire _w22247_ ;
	wire _w22248_ ;
	wire _w22249_ ;
	wire _w22250_ ;
	wire _w22251_ ;
	wire _w22252_ ;
	wire _w22253_ ;
	wire _w22254_ ;
	wire _w22255_ ;
	wire _w22256_ ;
	wire _w22257_ ;
	wire _w22258_ ;
	wire _w22259_ ;
	wire _w22260_ ;
	wire _w22261_ ;
	wire _w22262_ ;
	wire _w22263_ ;
	wire _w22264_ ;
	wire _w22265_ ;
	wire _w22266_ ;
	wire _w22267_ ;
	wire _w22268_ ;
	wire _w22269_ ;
	wire _w22270_ ;
	wire _w22271_ ;
	wire _w22272_ ;
	wire _w22273_ ;
	wire _w22274_ ;
	wire _w22275_ ;
	wire _w22276_ ;
	wire _w22277_ ;
	wire _w22278_ ;
	wire _w22279_ ;
	wire _w22280_ ;
	wire _w22281_ ;
	wire _w22282_ ;
	wire _w22283_ ;
	wire _w22284_ ;
	wire _w22285_ ;
	wire _w22286_ ;
	wire _w22287_ ;
	wire _w22288_ ;
	wire _w22289_ ;
	wire _w22290_ ;
	wire _w22291_ ;
	wire _w22292_ ;
	wire _w22293_ ;
	wire _w22294_ ;
	wire _w22295_ ;
	wire _w22296_ ;
	wire _w22297_ ;
	wire _w22298_ ;
	wire _w22299_ ;
	wire _w22300_ ;
	wire _w22301_ ;
	wire _w22302_ ;
	wire _w22303_ ;
	wire _w22304_ ;
	wire _w22305_ ;
	wire _w22306_ ;
	wire _w22307_ ;
	wire _w22308_ ;
	wire _w22309_ ;
	wire _w22310_ ;
	wire _w22311_ ;
	wire _w22312_ ;
	wire _w22313_ ;
	wire _w22314_ ;
	wire _w22315_ ;
	wire _w22316_ ;
	wire _w22317_ ;
	wire _w22318_ ;
	wire _w22319_ ;
	wire _w22320_ ;
	wire _w22321_ ;
	wire _w22322_ ;
	wire _w22323_ ;
	wire _w22324_ ;
	wire _w22325_ ;
	wire _w22326_ ;
	wire _w22327_ ;
	wire _w22328_ ;
	wire _w22329_ ;
	wire _w22330_ ;
	wire _w22331_ ;
	wire _w22332_ ;
	wire _w22333_ ;
	wire _w22334_ ;
	wire _w22335_ ;
	wire _w22336_ ;
	wire _w22337_ ;
	wire _w22338_ ;
	wire _w22339_ ;
	wire _w22340_ ;
	wire _w22341_ ;
	wire _w22342_ ;
	wire _w22343_ ;
	wire _w22344_ ;
	wire _w22345_ ;
	wire _w22346_ ;
	wire _w22347_ ;
	wire _w22348_ ;
	wire _w22349_ ;
	wire _w22350_ ;
	wire _w22351_ ;
	wire _w22352_ ;
	wire _w22353_ ;
	wire _w22354_ ;
	wire _w22355_ ;
	wire _w22356_ ;
	wire _w22357_ ;
	wire _w22358_ ;
	wire _w22359_ ;
	wire _w22360_ ;
	wire _w22361_ ;
	wire _w22362_ ;
	wire _w22363_ ;
	wire _w22364_ ;
	wire _w22365_ ;
	wire _w22366_ ;
	wire _w22367_ ;
	wire _w22368_ ;
	wire _w22369_ ;
	wire _w22370_ ;
	wire _w22371_ ;
	wire _w22372_ ;
	wire _w22373_ ;
	wire _w22374_ ;
	wire _w22375_ ;
	wire _w22376_ ;
	wire _w22377_ ;
	wire _w22378_ ;
	wire _w22379_ ;
	wire _w22380_ ;
	wire _w22381_ ;
	wire _w22382_ ;
	wire _w22383_ ;
	wire _w22384_ ;
	wire _w22385_ ;
	wire _w22386_ ;
	wire _w22387_ ;
	wire _w22388_ ;
	wire _w22389_ ;
	wire _w22390_ ;
	wire _w22391_ ;
	wire _w22392_ ;
	wire _w22393_ ;
	wire _w22394_ ;
	wire _w22395_ ;
	wire _w22396_ ;
	wire _w22397_ ;
	wire _w22398_ ;
	wire _w22399_ ;
	wire _w22400_ ;
	wire _w22401_ ;
	wire _w22402_ ;
	wire _w22403_ ;
	wire _w22404_ ;
	wire _w22405_ ;
	wire _w22406_ ;
	wire _w22407_ ;
	wire _w22408_ ;
	wire _w22409_ ;
	wire _w22410_ ;
	wire _w22411_ ;
	wire _w22412_ ;
	wire _w22413_ ;
	wire _w22414_ ;
	wire _w22415_ ;
	wire _w22416_ ;
	wire _w22417_ ;
	wire _w22418_ ;
	wire _w22419_ ;
	wire _w22420_ ;
	wire _w22421_ ;
	wire _w22422_ ;
	wire _w22423_ ;
	wire _w22424_ ;
	wire _w22425_ ;
	wire _w22426_ ;
	wire _w22427_ ;
	wire _w22428_ ;
	wire _w22429_ ;
	wire _w22430_ ;
	wire _w22431_ ;
	wire _w22432_ ;
	wire _w22433_ ;
	wire _w22434_ ;
	wire _w22435_ ;
	wire _w22436_ ;
	wire _w22437_ ;
	wire _w22438_ ;
	wire _w22439_ ;
	wire _w22440_ ;
	wire _w22441_ ;
	wire _w22442_ ;
	wire _w22443_ ;
	wire _w22444_ ;
	wire _w22445_ ;
	wire _w22446_ ;
	wire _w22447_ ;
	wire _w22448_ ;
	wire _w22449_ ;
	wire _w22450_ ;
	wire _w22451_ ;
	wire _w22452_ ;
	wire _w22453_ ;
	wire _w22454_ ;
	wire _w22455_ ;
	wire _w22456_ ;
	wire _w22457_ ;
	wire _w22458_ ;
	wire _w22459_ ;
	wire _w22460_ ;
	wire _w22461_ ;
	wire _w22462_ ;
	wire _w22463_ ;
	wire _w22464_ ;
	wire _w22465_ ;
	wire _w22466_ ;
	wire _w22467_ ;
	wire _w22468_ ;
	wire _w22469_ ;
	wire _w22470_ ;
	wire _w22471_ ;
	wire _w22472_ ;
	wire _w22473_ ;
	wire _w22474_ ;
	wire _w22475_ ;
	wire _w22476_ ;
	wire _w22477_ ;
	wire _w22478_ ;
	wire _w22479_ ;
	wire _w22480_ ;
	wire _w22481_ ;
	wire _w22482_ ;
	wire _w22483_ ;
	wire _w22484_ ;
	wire _w22485_ ;
	wire _w22486_ ;
	wire _w22487_ ;
	wire _w22488_ ;
	wire _w22489_ ;
	wire _w22490_ ;
	wire _w22491_ ;
	wire _w22492_ ;
	wire _w22493_ ;
	wire _w22494_ ;
	wire _w22495_ ;
	wire _w22496_ ;
	wire _w22497_ ;
	wire _w22498_ ;
	wire _w22499_ ;
	wire _w22500_ ;
	wire _w22501_ ;
	wire _w22502_ ;
	wire _w22503_ ;
	wire _w22504_ ;
	wire _w22505_ ;
	wire _w22506_ ;
	wire _w22507_ ;
	wire _w22508_ ;
	wire _w22509_ ;
	wire _w22510_ ;
	wire _w22511_ ;
	wire _w22512_ ;
	wire _w22513_ ;
	wire _w22514_ ;
	wire _w22515_ ;
	wire _w22516_ ;
	wire _w22517_ ;
	wire _w22518_ ;
	wire _w22519_ ;
	wire _w22520_ ;
	wire _w22521_ ;
	wire _w22522_ ;
	wire _w22523_ ;
	wire _w22524_ ;
	wire _w22525_ ;
	wire _w22526_ ;
	wire _w22527_ ;
	wire _w22528_ ;
	wire _w22529_ ;
	wire _w22530_ ;
	wire _w22531_ ;
	wire _w22532_ ;
	wire _w22533_ ;
	wire _w22534_ ;
	wire _w22535_ ;
	wire _w22536_ ;
	wire _w22537_ ;
	wire _w22538_ ;
	wire _w22539_ ;
	wire _w22540_ ;
	wire _w22541_ ;
	wire _w22542_ ;
	wire _w22543_ ;
	wire _w22544_ ;
	wire _w22545_ ;
	wire _w22546_ ;
	wire _w22547_ ;
	wire _w22548_ ;
	wire _w22549_ ;
	wire _w22550_ ;
	wire _w22551_ ;
	wire _w22552_ ;
	wire _w22553_ ;
	wire _w22554_ ;
	wire _w22555_ ;
	wire _w22556_ ;
	wire _w22557_ ;
	wire _w22558_ ;
	wire _w22559_ ;
	wire _w22560_ ;
	wire _w22561_ ;
	wire _w22562_ ;
	wire _w22563_ ;
	wire _w22564_ ;
	wire _w22565_ ;
	wire _w22566_ ;
	wire _w22567_ ;
	wire _w22568_ ;
	wire _w22569_ ;
	wire _w22570_ ;
	wire _w22571_ ;
	wire _w22572_ ;
	wire _w22573_ ;
	wire _w22574_ ;
	wire _w22575_ ;
	wire _w22576_ ;
	wire _w22577_ ;
	wire _w22578_ ;
	wire _w22579_ ;
	wire _w22580_ ;
	wire _w22581_ ;
	wire _w22582_ ;
	wire _w22583_ ;
	wire _w22584_ ;
	wire _w22585_ ;
	wire _w22586_ ;
	wire _w22587_ ;
	wire _w22588_ ;
	wire _w22589_ ;
	wire _w22590_ ;
	wire _w22591_ ;
	wire _w22592_ ;
	wire _w22593_ ;
	wire _w22594_ ;
	wire _w22595_ ;
	wire _w22596_ ;
	wire _w22597_ ;
	wire _w22598_ ;
	wire _w22599_ ;
	wire _w22600_ ;
	wire _w22601_ ;
	wire _w22602_ ;
	wire _w22603_ ;
	wire _w22604_ ;
	wire _w22605_ ;
	wire _w22606_ ;
	wire _w22607_ ;
	wire _w22608_ ;
	wire _w22609_ ;
	wire _w22610_ ;
	wire _w22611_ ;
	wire _w22612_ ;
	wire _w22613_ ;
	wire _w22614_ ;
	wire _w22615_ ;
	wire _w22616_ ;
	wire _w22617_ ;
	wire _w22618_ ;
	wire _w22619_ ;
	wire _w22620_ ;
	wire _w22621_ ;
	wire _w22622_ ;
	wire _w22623_ ;
	wire _w22624_ ;
	wire _w22625_ ;
	wire _w22626_ ;
	wire _w22627_ ;
	wire _w22628_ ;
	wire _w22629_ ;
	wire _w22630_ ;
	wire _w22631_ ;
	wire _w22632_ ;
	wire _w22633_ ;
	wire _w22634_ ;
	wire _w22635_ ;
	wire _w22636_ ;
	wire _w22637_ ;
	wire _w22638_ ;
	wire _w22639_ ;
	wire _w22640_ ;
	wire _w22641_ ;
	wire _w22642_ ;
	wire _w22643_ ;
	wire _w22644_ ;
	wire _w22645_ ;
	wire _w22646_ ;
	wire _w22647_ ;
	wire _w22648_ ;
	wire _w22649_ ;
	wire _w22650_ ;
	wire _w22651_ ;
	wire _w22652_ ;
	wire _w22653_ ;
	wire _w22654_ ;
	wire _w22655_ ;
	wire _w22656_ ;
	wire _w22657_ ;
	wire _w22658_ ;
	wire _w22659_ ;
	wire _w22660_ ;
	wire _w22661_ ;
	wire _w22662_ ;
	wire _w22663_ ;
	wire _w22664_ ;
	wire _w22665_ ;
	wire _w22666_ ;
	wire _w22667_ ;
	wire _w22668_ ;
	wire _w22669_ ;
	wire _w22670_ ;
	wire _w22671_ ;
	wire _w22672_ ;
	wire _w22673_ ;
	wire _w22674_ ;
	wire _w22675_ ;
	wire _w22676_ ;
	wire _w22677_ ;
	wire _w22678_ ;
	wire _w22679_ ;
	wire _w22680_ ;
	wire _w22681_ ;
	wire _w22682_ ;
	wire _w22683_ ;
	wire _w22684_ ;
	wire _w22685_ ;
	wire _w22686_ ;
	wire _w22687_ ;
	wire _w22688_ ;
	wire _w22689_ ;
	wire _w22690_ ;
	wire _w22691_ ;
	wire _w22692_ ;
	wire _w22693_ ;
	wire _w22694_ ;
	wire _w22695_ ;
	wire _w22696_ ;
	wire _w22697_ ;
	wire _w22698_ ;
	wire _w22699_ ;
	wire _w22700_ ;
	wire _w22701_ ;
	wire _w22702_ ;
	wire _w22703_ ;
	wire _w22704_ ;
	wire _w22705_ ;
	wire _w22706_ ;
	wire _w22707_ ;
	wire _w22708_ ;
	wire _w22709_ ;
	wire _w22710_ ;
	wire _w22711_ ;
	wire _w22712_ ;
	wire _w22713_ ;
	wire _w22714_ ;
	wire _w22715_ ;
	wire _w22716_ ;
	wire _w22717_ ;
	wire _w22718_ ;
	wire _w22719_ ;
	wire _w22720_ ;
	wire _w22721_ ;
	wire _w22722_ ;
	wire _w22723_ ;
	wire _w22724_ ;
	wire _w22725_ ;
	wire _w22726_ ;
	wire _w22727_ ;
	wire _w22728_ ;
	wire _w22729_ ;
	wire _w22730_ ;
	wire _w22731_ ;
	wire _w22732_ ;
	wire _w22733_ ;
	wire _w22734_ ;
	wire _w22735_ ;
	wire _w22736_ ;
	wire _w22737_ ;
	wire _w22738_ ;
	wire _w22739_ ;
	wire _w22740_ ;
	wire _w22741_ ;
	wire _w22742_ ;
	wire _w22743_ ;
	wire _w22744_ ;
	wire _w22745_ ;
	wire _w22746_ ;
	wire _w22747_ ;
	wire _w22748_ ;
	wire _w22749_ ;
	wire _w22750_ ;
	wire _w22751_ ;
	wire _w22752_ ;
	wire _w22753_ ;
	wire _w22754_ ;
	wire _w22755_ ;
	wire _w22756_ ;
	wire _w22757_ ;
	wire _w22758_ ;
	wire _w22759_ ;
	wire _w22760_ ;
	wire _w22761_ ;
	wire _w22762_ ;
	wire _w22763_ ;
	wire _w22764_ ;
	wire _w22765_ ;
	wire _w22766_ ;
	wire _w22767_ ;
	wire _w22768_ ;
	wire _w22769_ ;
	wire _w22770_ ;
	wire _w22771_ ;
	wire _w22772_ ;
	wire _w22773_ ;
	wire _w22774_ ;
	wire _w22775_ ;
	wire _w22776_ ;
	wire _w22777_ ;
	wire _w22778_ ;
	wire _w22779_ ;
	wire _w22780_ ;
	wire _w22781_ ;
	wire _w22782_ ;
	wire _w22783_ ;
	wire _w22784_ ;
	wire _w22785_ ;
	wire _w22786_ ;
	wire _w22787_ ;
	wire _w22788_ ;
	wire _w22789_ ;
	wire _w22790_ ;
	wire _w22791_ ;
	wire _w22792_ ;
	wire _w22793_ ;
	wire _w22794_ ;
	wire _w22795_ ;
	wire _w22796_ ;
	wire _w22797_ ;
	wire _w22798_ ;
	wire _w22799_ ;
	wire _w22800_ ;
	wire _w22801_ ;
	wire _w22802_ ;
	wire _w22803_ ;
	wire _w22804_ ;
	wire _w22805_ ;
	wire _w22806_ ;
	wire _w22807_ ;
	wire _w22808_ ;
	wire _w22809_ ;
	wire _w22810_ ;
	wire _w22811_ ;
	wire _w22812_ ;
	wire _w22813_ ;
	wire _w22814_ ;
	wire _w22815_ ;
	wire _w22816_ ;
	wire _w22817_ ;
	wire _w22818_ ;
	wire _w22819_ ;
	wire _w22820_ ;
	wire _w22821_ ;
	wire _w22822_ ;
	wire _w22823_ ;
	wire _w22824_ ;
	wire _w22825_ ;
	wire _w22826_ ;
	wire _w22827_ ;
	wire _w22828_ ;
	wire _w22829_ ;
	wire _w22830_ ;
	wire _w22831_ ;
	wire _w22832_ ;
	wire _w22833_ ;
	wire _w22834_ ;
	wire _w22835_ ;
	wire _w22836_ ;
	wire _w22837_ ;
	wire _w22838_ ;
	wire _w22839_ ;
	wire _w22840_ ;
	wire _w22841_ ;
	wire _w22842_ ;
	wire _w22843_ ;
	wire _w22844_ ;
	wire _w22845_ ;
	wire _w22846_ ;
	wire _w22847_ ;
	wire _w22848_ ;
	wire _w22849_ ;
	wire _w22850_ ;
	wire _w22851_ ;
	wire _w22852_ ;
	wire _w22853_ ;
	wire _w22854_ ;
	wire _w22855_ ;
	wire _w22856_ ;
	wire _w22857_ ;
	wire _w22858_ ;
	wire _w22859_ ;
	wire _w22860_ ;
	wire _w22861_ ;
	wire _w22862_ ;
	wire _w22863_ ;
	wire _w22864_ ;
	wire _w22865_ ;
	wire _w22866_ ;
	wire _w22867_ ;
	wire _w22868_ ;
	wire _w22869_ ;
	wire _w22870_ ;
	wire _w22871_ ;
	wire _w22872_ ;
	wire _w22873_ ;
	wire _w22874_ ;
	wire _w22875_ ;
	wire _w22876_ ;
	wire _w22877_ ;
	wire _w22878_ ;
	wire _w22879_ ;
	wire _w22880_ ;
	wire _w22881_ ;
	wire _w22882_ ;
	wire _w22883_ ;
	wire _w22884_ ;
	wire _w22885_ ;
	wire _w22886_ ;
	wire _w22887_ ;
	wire _w22888_ ;
	wire _w22889_ ;
	wire _w22890_ ;
	wire _w22891_ ;
	wire _w22892_ ;
	wire _w22893_ ;
	wire _w22894_ ;
	wire _w22895_ ;
	wire _w22896_ ;
	wire _w22897_ ;
	wire _w22898_ ;
	wire _w22899_ ;
	wire _w22900_ ;
	wire _w22901_ ;
	wire _w22902_ ;
	wire _w22903_ ;
	wire _w22904_ ;
	wire _w22905_ ;
	wire _w22906_ ;
	wire _w22907_ ;
	wire _w22908_ ;
	wire _w22909_ ;
	wire _w22910_ ;
	wire _w22911_ ;
	wire _w22912_ ;
	wire _w22913_ ;
	wire _w22914_ ;
	wire _w22915_ ;
	wire _w22916_ ;
	wire _w22917_ ;
	wire _w22918_ ;
	wire _w22919_ ;
	wire _w22920_ ;
	wire _w22921_ ;
	wire _w22922_ ;
	wire _w22923_ ;
	wire _w22924_ ;
	wire _w22925_ ;
	wire _w22926_ ;
	wire _w22927_ ;
	wire _w22928_ ;
	wire _w22929_ ;
	wire _w22930_ ;
	wire _w22931_ ;
	wire _w22932_ ;
	wire _w22933_ ;
	wire _w22934_ ;
	wire _w22935_ ;
	wire _w22936_ ;
	wire _w22937_ ;
	wire _w22938_ ;
	wire _w22939_ ;
	wire _w22940_ ;
	wire _w22941_ ;
	wire _w22942_ ;
	wire _w22943_ ;
	wire _w22944_ ;
	wire _w22945_ ;
	wire _w22946_ ;
	wire _w22947_ ;
	wire _w22948_ ;
	wire _w22949_ ;
	wire _w22950_ ;
	wire _w22951_ ;
	wire _w22952_ ;
	wire _w22953_ ;
	wire _w22954_ ;
	wire _w22955_ ;
	wire _w22956_ ;
	wire _w22957_ ;
	wire _w22958_ ;
	wire _w22959_ ;
	wire _w22960_ ;
	wire _w22961_ ;
	wire _w22962_ ;
	wire _w22963_ ;
	wire _w22964_ ;
	wire _w22965_ ;
	wire _w22966_ ;
	wire _w22967_ ;
	wire _w22968_ ;
	wire _w22969_ ;
	wire _w22970_ ;
	wire _w22971_ ;
	wire _w22972_ ;
	wire _w22973_ ;
	wire _w22974_ ;
	wire _w22975_ ;
	wire _w22976_ ;
	wire _w22977_ ;
	wire _w22978_ ;
	wire _w22979_ ;
	wire _w22980_ ;
	wire _w22981_ ;
	wire _w22982_ ;
	wire _w22983_ ;
	wire _w22984_ ;
	wire _w22985_ ;
	wire _w22986_ ;
	wire _w22987_ ;
	wire _w22988_ ;
	wire _w22989_ ;
	wire _w22990_ ;
	wire _w22991_ ;
	wire _w22992_ ;
	wire _w22993_ ;
	wire _w22994_ ;
	wire _w22995_ ;
	wire _w22996_ ;
	wire _w22997_ ;
	wire _w22998_ ;
	wire _w22999_ ;
	wire _w23000_ ;
	wire _w23001_ ;
	wire _w23002_ ;
	wire _w23003_ ;
	wire _w23004_ ;
	wire _w23005_ ;
	wire _w23006_ ;
	wire _w23007_ ;
	wire _w23008_ ;
	wire _w23009_ ;
	wire _w23010_ ;
	wire _w23011_ ;
	wire _w23012_ ;
	wire _w23013_ ;
	wire _w23014_ ;
	wire _w23015_ ;
	wire _w23016_ ;
	wire _w23017_ ;
	wire _w23018_ ;
	wire _w23019_ ;
	wire _w23020_ ;
	wire _w23021_ ;
	wire _w23022_ ;
	wire _w23023_ ;
	wire _w23024_ ;
	wire _w23025_ ;
	wire _w23026_ ;
	wire _w23027_ ;
	wire _w23028_ ;
	wire _w23029_ ;
	wire _w23030_ ;
	wire _w23031_ ;
	wire _w23032_ ;
	wire _w23033_ ;
	wire _w23034_ ;
	wire _w23035_ ;
	wire _w23036_ ;
	wire _w23037_ ;
	wire _w23038_ ;
	wire _w23039_ ;
	wire _w23040_ ;
	wire _w23041_ ;
	wire _w23042_ ;
	wire _w23043_ ;
	wire _w23044_ ;
	wire _w23045_ ;
	wire _w23046_ ;
	wire _w23047_ ;
	wire _w23048_ ;
	wire _w23049_ ;
	wire _w23050_ ;
	wire _w23051_ ;
	wire _w23052_ ;
	wire _w23053_ ;
	wire _w23054_ ;
	wire _w23055_ ;
	wire _w23056_ ;
	wire _w23057_ ;
	wire _w23058_ ;
	wire _w23059_ ;
	wire _w23060_ ;
	wire _w23061_ ;
	wire _w23062_ ;
	wire _w23063_ ;
	wire _w23064_ ;
	wire _w23065_ ;
	wire _w23066_ ;
	wire _w23067_ ;
	wire _w23068_ ;
	wire _w23069_ ;
	wire _w23070_ ;
	wire _w23071_ ;
	wire _w23072_ ;
	wire _w23073_ ;
	wire _w23074_ ;
	wire _w23075_ ;
	wire _w23076_ ;
	wire _w23077_ ;
	wire _w23078_ ;
	wire _w23079_ ;
	wire _w23080_ ;
	wire _w23081_ ;
	wire _w23082_ ;
	wire _w23083_ ;
	wire _w23084_ ;
	wire _w23085_ ;
	wire _w23086_ ;
	wire _w23087_ ;
	wire _w23088_ ;
	wire _w23089_ ;
	wire _w23090_ ;
	wire _w23091_ ;
	wire _w23092_ ;
	wire _w23093_ ;
	wire _w23094_ ;
	wire _w23095_ ;
	wire _w23096_ ;
	wire _w23097_ ;
	wire _w23098_ ;
	wire _w23099_ ;
	wire _w23100_ ;
	wire _w23101_ ;
	wire _w23102_ ;
	wire _w23103_ ;
	wire _w23104_ ;
	wire _w23105_ ;
	wire _w23106_ ;
	wire _w23107_ ;
	wire _w23108_ ;
	wire _w23109_ ;
	wire _w23110_ ;
	wire _w23111_ ;
	wire _w23112_ ;
	wire _w23113_ ;
	wire _w23114_ ;
	wire _w23115_ ;
	wire _w23116_ ;
	wire _w23117_ ;
	wire _w23118_ ;
	wire _w23119_ ;
	wire _w23120_ ;
	wire _w23121_ ;
	wire _w23122_ ;
	wire _w23123_ ;
	wire _w23124_ ;
	wire _w23125_ ;
	wire _w23126_ ;
	wire _w23127_ ;
	wire _w23128_ ;
	wire _w23129_ ;
	wire _w23130_ ;
	wire _w23131_ ;
	wire _w23132_ ;
	wire _w23133_ ;
	wire _w23134_ ;
	wire _w23135_ ;
	wire _w23136_ ;
	wire _w23137_ ;
	wire _w23138_ ;
	wire _w23139_ ;
	wire _w23140_ ;
	wire _w23141_ ;
	wire _w23142_ ;
	wire _w23143_ ;
	wire _w23144_ ;
	wire _w23145_ ;
	wire _w23146_ ;
	wire _w23147_ ;
	wire _w23148_ ;
	wire _w23149_ ;
	wire _w23150_ ;
	wire _w23151_ ;
	wire _w23152_ ;
	wire _w23153_ ;
	wire _w23154_ ;
	wire _w23155_ ;
	wire _w23156_ ;
	wire _w23157_ ;
	wire _w23158_ ;
	wire _w23159_ ;
	wire _w23160_ ;
	wire _w23161_ ;
	wire _w23162_ ;
	wire _w23163_ ;
	wire _w23164_ ;
	wire _w23165_ ;
	wire _w23166_ ;
	wire _w23167_ ;
	wire _w23168_ ;
	wire _w23169_ ;
	wire _w23170_ ;
	wire _w23171_ ;
	wire _w23172_ ;
	wire _w23173_ ;
	wire _w23174_ ;
	wire _w23175_ ;
	wire _w23176_ ;
	wire _w23177_ ;
	wire _w23178_ ;
	wire _w23179_ ;
	wire _w23180_ ;
	wire _w23181_ ;
	wire _w23182_ ;
	wire _w23183_ ;
	wire _w23184_ ;
	wire _w23185_ ;
	wire _w23186_ ;
	wire _w23187_ ;
	wire _w23188_ ;
	wire _w23189_ ;
	wire _w23190_ ;
	wire _w23191_ ;
	wire _w23192_ ;
	wire _w23193_ ;
	wire _w23194_ ;
	wire _w23195_ ;
	wire _w23196_ ;
	wire _w23197_ ;
	wire _w23198_ ;
	wire _w23199_ ;
	wire _w23200_ ;
	wire _w23201_ ;
	wire _w23202_ ;
	wire _w23203_ ;
	wire _w23204_ ;
	wire _w23205_ ;
	wire _w23206_ ;
	wire _w23207_ ;
	wire _w23208_ ;
	wire _w23209_ ;
	wire _w23210_ ;
	wire _w23211_ ;
	wire _w23212_ ;
	wire _w23213_ ;
	wire _w23214_ ;
	wire _w23215_ ;
	wire _w23216_ ;
	wire _w23217_ ;
	wire _w23218_ ;
	wire _w23219_ ;
	wire _w23220_ ;
	wire _w23221_ ;
	wire _w23222_ ;
	wire _w23223_ ;
	wire _w23224_ ;
	wire _w23225_ ;
	wire _w23226_ ;
	wire _w23227_ ;
	wire _w23228_ ;
	wire _w23229_ ;
	wire _w23230_ ;
	wire _w23231_ ;
	wire _w23232_ ;
	wire _w23233_ ;
	wire _w23234_ ;
	wire _w23235_ ;
	wire _w23236_ ;
	wire _w23237_ ;
	wire _w23238_ ;
	wire _w23239_ ;
	wire _w23240_ ;
	wire _w23241_ ;
	wire _w23242_ ;
	wire _w23243_ ;
	wire _w23244_ ;
	wire _w23245_ ;
	wire _w23246_ ;
	wire _w23247_ ;
	wire _w23248_ ;
	wire _w23249_ ;
	wire _w23250_ ;
	wire _w23251_ ;
	wire _w23252_ ;
	wire _w23253_ ;
	wire _w23254_ ;
	wire _w23255_ ;
	wire _w23256_ ;
	wire _w23257_ ;
	wire _w23258_ ;
	wire _w23259_ ;
	wire _w23260_ ;
	wire _w23261_ ;
	wire _w23262_ ;
	wire _w23263_ ;
	wire _w23264_ ;
	wire _w23265_ ;
	wire _w23266_ ;
	wire _w23267_ ;
	wire _w23268_ ;
	wire _w23269_ ;
	wire _w23270_ ;
	wire _w23271_ ;
	wire _w23272_ ;
	wire _w23273_ ;
	wire _w23274_ ;
	wire _w23275_ ;
	wire _w23276_ ;
	wire _w23277_ ;
	wire _w23278_ ;
	wire _w23279_ ;
	wire _w23280_ ;
	wire _w23281_ ;
	wire _w23282_ ;
	wire _w23283_ ;
	wire _w23284_ ;
	wire _w23285_ ;
	wire _w23286_ ;
	wire _w23287_ ;
	wire _w23288_ ;
	wire _w23289_ ;
	wire _w23290_ ;
	wire _w23291_ ;
	wire _w23292_ ;
	wire _w23293_ ;
	wire _w23294_ ;
	wire _w23295_ ;
	wire _w23296_ ;
	wire _w23297_ ;
	wire _w23298_ ;
	wire _w23299_ ;
	wire _w23300_ ;
	wire _w23301_ ;
	wire _w23302_ ;
	wire _w23303_ ;
	wire _w23304_ ;
	wire _w23305_ ;
	wire _w23306_ ;
	wire _w23307_ ;
	wire _w23308_ ;
	wire _w23309_ ;
	wire _w23310_ ;
	wire _w23311_ ;
	wire _w23312_ ;
	wire _w23313_ ;
	wire _w23314_ ;
	wire _w23315_ ;
	wire _w23316_ ;
	wire _w23317_ ;
	wire _w23318_ ;
	wire _w23319_ ;
	wire _w23320_ ;
	wire _w23321_ ;
	wire _w23322_ ;
	wire _w23323_ ;
	wire _w23324_ ;
	wire _w23325_ ;
	wire _w23326_ ;
	wire _w23327_ ;
	wire _w23328_ ;
	wire _w23329_ ;
	wire _w23330_ ;
	wire _w23331_ ;
	wire _w23332_ ;
	wire _w23333_ ;
	wire _w23334_ ;
	wire _w23335_ ;
	wire _w23336_ ;
	wire _w23337_ ;
	wire _w23338_ ;
	wire _w23339_ ;
	wire _w23340_ ;
	wire _w23341_ ;
	wire _w23342_ ;
	wire _w23343_ ;
	wire _w23344_ ;
	wire _w23345_ ;
	wire _w23346_ ;
	wire _w23347_ ;
	wire _w23348_ ;
	wire _w23349_ ;
	wire _w23350_ ;
	wire _w23351_ ;
	wire _w23352_ ;
	wire _w23353_ ;
	wire _w23354_ ;
	wire _w23355_ ;
	wire _w23356_ ;
	wire _w23357_ ;
	wire _w23358_ ;
	wire _w23359_ ;
	wire _w23360_ ;
	wire _w23361_ ;
	wire _w23362_ ;
	wire _w23363_ ;
	wire _w23364_ ;
	wire _w23365_ ;
	wire _w23366_ ;
	wire _w23367_ ;
	wire _w23368_ ;
	wire _w23369_ ;
	wire _w23370_ ;
	wire _w23371_ ;
	wire _w23372_ ;
	wire _w23373_ ;
	wire _w23374_ ;
	wire _w23375_ ;
	wire _w23376_ ;
	wire _w23377_ ;
	wire _w23378_ ;
	wire _w23379_ ;
	wire _w23380_ ;
	wire _w23381_ ;
	wire _w23382_ ;
	wire _w23383_ ;
	wire _w23384_ ;
	wire _w23385_ ;
	wire _w23386_ ;
	wire _w23387_ ;
	wire _w23388_ ;
	wire _w23389_ ;
	wire _w23390_ ;
	wire _w23391_ ;
	wire _w23392_ ;
	wire _w23393_ ;
	wire _w23394_ ;
	wire _w23395_ ;
	wire _w23396_ ;
	wire _w23397_ ;
	wire _w23398_ ;
	wire _w23399_ ;
	wire _w23400_ ;
	wire _w23401_ ;
	wire _w23402_ ;
	wire _w23403_ ;
	wire _w23404_ ;
	wire _w23405_ ;
	wire _w23406_ ;
	wire _w23407_ ;
	wire _w23408_ ;
	wire _w23409_ ;
	wire _w23410_ ;
	wire _w23411_ ;
	wire _w23412_ ;
	wire _w23413_ ;
	wire _w23414_ ;
	wire _w23415_ ;
	wire _w23416_ ;
	wire _w23417_ ;
	wire _w23418_ ;
	wire _w23419_ ;
	wire _w23420_ ;
	wire _w23421_ ;
	wire _w23422_ ;
	wire _w23423_ ;
	wire _w23424_ ;
	wire _w23425_ ;
	wire _w23426_ ;
	wire _w23427_ ;
	wire _w23428_ ;
	wire _w23429_ ;
	wire _w23430_ ;
	wire _w23431_ ;
	wire _w23432_ ;
	wire _w23433_ ;
	wire _w23434_ ;
	wire _w23435_ ;
	wire _w23436_ ;
	wire _w23437_ ;
	wire _w23438_ ;
	wire _w23439_ ;
	wire _w23440_ ;
	wire _w23441_ ;
	wire _w23442_ ;
	wire _w23443_ ;
	wire _w23444_ ;
	wire _w23445_ ;
	wire _w23446_ ;
	wire _w23447_ ;
	wire _w23448_ ;
	wire _w23449_ ;
	wire _w23450_ ;
	wire _w23451_ ;
	wire _w23452_ ;
	wire _w23453_ ;
	wire _w23454_ ;
	wire _w23455_ ;
	wire _w23456_ ;
	wire _w23457_ ;
	wire _w23458_ ;
	wire _w23459_ ;
	wire _w23460_ ;
	wire _w23461_ ;
	wire _w23462_ ;
	wire _w23463_ ;
	wire _w23464_ ;
	wire _w23465_ ;
	wire _w23466_ ;
	wire _w23467_ ;
	wire _w23468_ ;
	wire _w23469_ ;
	wire _w23470_ ;
	wire _w23471_ ;
	wire _w23472_ ;
	wire _w23473_ ;
	wire _w23474_ ;
	wire _w23475_ ;
	wire _w23476_ ;
	wire _w23477_ ;
	wire _w23478_ ;
	wire _w23479_ ;
	wire _w23480_ ;
	wire _w23481_ ;
	wire _w23482_ ;
	wire _w23483_ ;
	wire _w23484_ ;
	wire _w23485_ ;
	wire _w23486_ ;
	wire _w23487_ ;
	wire _w23488_ ;
	wire _w23489_ ;
	wire _w23490_ ;
	wire _w23491_ ;
	wire _w23492_ ;
	wire _w23493_ ;
	wire _w23494_ ;
	wire _w23495_ ;
	wire _w23496_ ;
	wire _w23497_ ;
	wire _w23498_ ;
	wire _w23499_ ;
	wire _w23500_ ;
	wire _w23501_ ;
	wire _w23502_ ;
	wire _w23503_ ;
	wire _w23504_ ;
	wire _w23505_ ;
	wire _w23506_ ;
	wire _w23507_ ;
	wire _w23508_ ;
	wire _w23509_ ;
	wire _w23510_ ;
	wire _w23511_ ;
	wire _w23512_ ;
	wire _w23513_ ;
	wire _w23514_ ;
	wire _w23515_ ;
	wire _w23516_ ;
	wire _w23517_ ;
	wire _w23518_ ;
	wire _w23519_ ;
	wire _w23520_ ;
	wire _w23521_ ;
	wire _w23522_ ;
	wire _w23523_ ;
	wire _w23524_ ;
	wire _w23525_ ;
	wire _w23526_ ;
	wire _w23527_ ;
	wire _w23528_ ;
	wire _w23529_ ;
	wire _w23530_ ;
	wire _w23531_ ;
	wire _w23532_ ;
	wire _w23533_ ;
	wire _w23534_ ;
	wire _w23535_ ;
	wire _w23536_ ;
	wire _w23537_ ;
	wire _w23538_ ;
	wire _w23539_ ;
	wire _w23540_ ;
	wire _w23541_ ;
	wire _w23542_ ;
	wire _w23543_ ;
	wire _w23544_ ;
	wire _w23545_ ;
	wire _w23546_ ;
	wire _w23547_ ;
	wire _w23548_ ;
	wire _w23549_ ;
	wire _w23550_ ;
	wire _w23551_ ;
	wire _w23552_ ;
	wire _w23553_ ;
	wire _w23554_ ;
	wire _w23555_ ;
	wire _w23556_ ;
	wire _w23557_ ;
	wire _w23558_ ;
	wire _w23559_ ;
	wire _w23560_ ;
	wire _w23561_ ;
	wire _w23562_ ;
	wire _w23563_ ;
	wire _w23564_ ;
	wire _w23565_ ;
	wire _w23566_ ;
	wire _w23567_ ;
	wire _w23568_ ;
	wire _w23569_ ;
	wire _w23570_ ;
	wire _w23571_ ;
	wire _w23572_ ;
	wire _w23573_ ;
	wire _w23574_ ;
	wire _w23575_ ;
	wire _w23576_ ;
	wire _w23577_ ;
	wire _w23578_ ;
	wire _w23579_ ;
	wire _w23580_ ;
	wire _w23581_ ;
	wire _w23582_ ;
	wire _w23583_ ;
	wire _w23584_ ;
	wire _w23585_ ;
	wire _w23586_ ;
	wire _w23587_ ;
	wire _w23588_ ;
	wire _w23589_ ;
	wire _w23590_ ;
	wire _w23591_ ;
	wire _w23592_ ;
	wire _w23593_ ;
	wire _w23594_ ;
	wire _w23595_ ;
	wire _w23596_ ;
	wire _w23597_ ;
	wire _w23598_ ;
	wire _w23599_ ;
	wire _w23600_ ;
	wire _w23601_ ;
	wire _w23602_ ;
	wire _w23603_ ;
	wire _w23604_ ;
	wire _w23605_ ;
	wire _w23606_ ;
	wire _w23607_ ;
	wire _w23608_ ;
	wire _w23609_ ;
	wire _w23610_ ;
	wire _w23611_ ;
	wire _w23612_ ;
	wire _w23613_ ;
	wire _w23614_ ;
	wire _w23615_ ;
	wire _w23616_ ;
	wire _w23617_ ;
	wire _w23618_ ;
	wire _w23619_ ;
	wire _w23620_ ;
	wire _w23621_ ;
	wire _w23622_ ;
	wire _w23623_ ;
	wire _w23624_ ;
	wire _w23625_ ;
	wire _w23626_ ;
	wire _w23627_ ;
	wire _w23628_ ;
	wire _w23629_ ;
	wire _w23630_ ;
	wire _w23631_ ;
	wire _w23632_ ;
	wire _w23633_ ;
	wire _w23634_ ;
	wire _w23635_ ;
	wire _w23636_ ;
	wire _w23637_ ;
	wire _w23638_ ;
	wire _w23639_ ;
	wire _w23640_ ;
	wire _w23641_ ;
	wire _w23642_ ;
	wire _w23643_ ;
	wire _w23644_ ;
	wire _w23645_ ;
	wire _w23646_ ;
	wire _w23647_ ;
	wire _w23648_ ;
	wire _w23649_ ;
	wire _w23650_ ;
	wire _w23651_ ;
	wire _w23652_ ;
	wire _w23653_ ;
	wire _w23654_ ;
	wire _w23655_ ;
	wire _w23656_ ;
	wire _w23657_ ;
	wire _w23658_ ;
	wire _w23659_ ;
	wire _w23660_ ;
	wire _w23661_ ;
	wire _w23662_ ;
	wire _w23663_ ;
	wire _w23664_ ;
	wire _w23665_ ;
	wire _w23666_ ;
	wire _w23667_ ;
	wire _w23668_ ;
	wire _w23669_ ;
	wire _w23670_ ;
	wire _w23671_ ;
	wire _w23672_ ;
	wire _w23673_ ;
	wire _w23674_ ;
	wire _w23675_ ;
	wire _w23676_ ;
	wire _w23677_ ;
	wire _w23678_ ;
	wire _w23679_ ;
	wire _w23680_ ;
	wire _w23681_ ;
	wire _w23682_ ;
	wire _w23683_ ;
	wire _w23684_ ;
	wire _w23685_ ;
	wire _w23686_ ;
	wire _w23687_ ;
	wire _w23688_ ;
	wire _w23689_ ;
	wire _w23690_ ;
	wire _w23691_ ;
	wire _w23692_ ;
	wire _w23693_ ;
	wire _w23694_ ;
	wire _w23695_ ;
	wire _w23696_ ;
	wire _w23697_ ;
	wire _w23698_ ;
	wire _w23699_ ;
	wire _w23700_ ;
	wire _w23701_ ;
	wire _w23702_ ;
	wire _w23703_ ;
	wire _w23704_ ;
	wire _w23705_ ;
	wire _w23706_ ;
	wire _w23707_ ;
	wire _w23708_ ;
	wire _w23709_ ;
	wire _w23710_ ;
	wire _w23711_ ;
	wire _w23712_ ;
	wire _w23713_ ;
	wire _w23714_ ;
	wire _w23715_ ;
	wire _w23716_ ;
	wire _w23717_ ;
	wire _w23718_ ;
	wire _w23719_ ;
	wire _w23720_ ;
	wire _w23721_ ;
	wire _w23722_ ;
	wire _w23723_ ;
	wire _w23724_ ;
	wire _w23725_ ;
	wire _w23726_ ;
	wire _w23727_ ;
	wire _w23728_ ;
	wire _w23729_ ;
	wire _w23730_ ;
	wire _w23731_ ;
	wire _w23732_ ;
	wire _w23733_ ;
	wire _w23734_ ;
	wire _w23735_ ;
	wire _w23736_ ;
	wire _w23737_ ;
	wire _w23738_ ;
	wire _w23739_ ;
	wire _w23740_ ;
	wire _w23741_ ;
	wire _w23742_ ;
	wire _w23743_ ;
	wire _w23744_ ;
	wire _w23745_ ;
	wire _w23746_ ;
	wire _w23747_ ;
	wire _w23748_ ;
	wire _w23749_ ;
	wire _w23750_ ;
	wire _w23751_ ;
	wire _w23752_ ;
	wire _w23753_ ;
	wire _w23754_ ;
	wire _w23755_ ;
	wire _w23756_ ;
	wire _w23757_ ;
	wire _w23758_ ;
	wire _w23759_ ;
	wire _w23760_ ;
	wire _w23761_ ;
	wire _w23762_ ;
	wire _w23763_ ;
	wire _w23764_ ;
	wire _w23765_ ;
	wire _w23766_ ;
	wire _w23767_ ;
	wire _w23768_ ;
	wire _w23769_ ;
	wire _w23770_ ;
	wire _w23771_ ;
	wire _w23772_ ;
	wire _w23773_ ;
	wire _w23774_ ;
	wire _w23775_ ;
	wire _w23776_ ;
	wire _w23777_ ;
	wire _w23778_ ;
	wire _w23779_ ;
	wire _w23780_ ;
	wire _w23781_ ;
	wire _w23782_ ;
	wire _w23783_ ;
	wire _w23784_ ;
	wire _w23785_ ;
	wire _w23786_ ;
	wire _w23787_ ;
	wire _w23788_ ;
	wire _w23789_ ;
	wire _w23790_ ;
	wire _w23791_ ;
	wire _w23792_ ;
	wire _w23793_ ;
	wire _w23794_ ;
	wire _w23795_ ;
	wire _w23796_ ;
	wire _w23797_ ;
	wire _w23798_ ;
	wire _w23799_ ;
	wire _w23800_ ;
	wire _w23801_ ;
	wire _w23802_ ;
	wire _w23803_ ;
	wire _w23804_ ;
	wire _w23805_ ;
	wire _w23806_ ;
	wire _w23807_ ;
	wire _w23808_ ;
	wire _w23809_ ;
	wire _w23810_ ;
	wire _w23811_ ;
	wire _w23812_ ;
	wire _w23813_ ;
	wire _w23814_ ;
	wire _w23815_ ;
	wire _w23816_ ;
	wire _w23817_ ;
	wire _w23818_ ;
	wire _w23819_ ;
	wire _w23820_ ;
	wire _w23821_ ;
	wire _w23822_ ;
	wire _w23823_ ;
	wire _w23824_ ;
	wire _w23825_ ;
	wire _w23826_ ;
	wire _w23827_ ;
	wire _w23828_ ;
	wire _w23829_ ;
	wire _w23830_ ;
	wire _w23831_ ;
	wire _w23832_ ;
	wire _w23833_ ;
	wire _w23834_ ;
	wire _w23835_ ;
	wire _w23836_ ;
	wire _w23837_ ;
	wire _w23838_ ;
	wire _w23839_ ;
	wire _w23840_ ;
	wire _w23841_ ;
	wire _w23842_ ;
	wire _w23843_ ;
	wire _w23844_ ;
	wire _w23845_ ;
	wire _w23846_ ;
	wire _w23847_ ;
	wire _w23848_ ;
	wire _w23849_ ;
	wire _w23850_ ;
	wire _w23851_ ;
	wire _w23852_ ;
	wire _w23853_ ;
	wire _w23854_ ;
	wire _w23855_ ;
	wire _w23856_ ;
	wire _w23857_ ;
	wire _w23858_ ;
	wire _w23859_ ;
	wire _w23860_ ;
	wire _w23861_ ;
	wire _w23862_ ;
	wire _w23863_ ;
	wire _w23864_ ;
	wire _w23865_ ;
	wire _w23866_ ;
	wire _w23867_ ;
	wire _w23868_ ;
	wire _w23869_ ;
	wire _w23870_ ;
	wire _w23871_ ;
	wire _w23872_ ;
	wire _w23873_ ;
	wire _w23874_ ;
	wire _w23875_ ;
	wire _w23876_ ;
	wire _w23877_ ;
	wire _w23878_ ;
	wire _w23879_ ;
	wire _w23880_ ;
	wire _w23881_ ;
	wire _w23882_ ;
	wire _w23883_ ;
	wire _w23884_ ;
	wire _w23885_ ;
	wire _w23886_ ;
	wire _w23887_ ;
	wire _w23888_ ;
	wire _w23889_ ;
	wire _w23890_ ;
	wire _w23891_ ;
	wire _w23892_ ;
	wire _w23893_ ;
	wire _w23894_ ;
	wire _w23895_ ;
	wire _w23896_ ;
	wire _w23897_ ;
	wire _w23898_ ;
	wire _w23899_ ;
	wire _w23900_ ;
	wire _w23901_ ;
	wire _w23902_ ;
	wire _w23903_ ;
	wire _w23904_ ;
	wire _w23905_ ;
	wire _w23906_ ;
	wire _w23907_ ;
	wire _w23908_ ;
	wire _w23909_ ;
	wire _w23910_ ;
	wire _w23911_ ;
	wire _w23912_ ;
	wire _w23913_ ;
	wire _w23914_ ;
	wire _w23915_ ;
	wire _w23916_ ;
	wire _w23917_ ;
	wire _w23918_ ;
	wire _w23919_ ;
	wire _w23920_ ;
	wire _w23921_ ;
	wire _w23922_ ;
	wire _w23923_ ;
	wire _w23924_ ;
	wire _w23925_ ;
	wire _w23926_ ;
	wire _w23927_ ;
	wire _w23928_ ;
	wire _w23929_ ;
	wire _w23930_ ;
	wire _w23931_ ;
	wire _w23932_ ;
	wire _w23933_ ;
	wire _w23934_ ;
	wire _w23935_ ;
	wire _w23936_ ;
	wire _w23937_ ;
	wire _w23938_ ;
	wire _w23939_ ;
	wire _w23940_ ;
	wire _w23941_ ;
	wire _w23942_ ;
	wire _w23943_ ;
	wire _w23944_ ;
	wire _w23945_ ;
	wire _w23946_ ;
	wire _w23947_ ;
	wire _w23948_ ;
	wire _w23949_ ;
	wire _w23950_ ;
	wire _w23951_ ;
	wire _w23952_ ;
	wire _w23953_ ;
	wire _w23954_ ;
	wire _w23955_ ;
	wire _w23956_ ;
	wire _w23957_ ;
	wire _w23958_ ;
	wire _w23959_ ;
	wire _w23960_ ;
	wire _w23961_ ;
	wire _w23962_ ;
	wire _w23963_ ;
	wire _w23964_ ;
	wire _w23965_ ;
	wire _w23966_ ;
	wire _w23967_ ;
	wire _w23968_ ;
	wire _w23969_ ;
	wire _w23970_ ;
	wire _w23971_ ;
	wire _w23972_ ;
	wire _w23973_ ;
	wire _w23974_ ;
	wire _w23975_ ;
	wire _w23976_ ;
	wire _w23977_ ;
	wire _w23978_ ;
	wire _w23979_ ;
	wire _w23980_ ;
	wire _w23981_ ;
	wire _w23982_ ;
	wire _w23983_ ;
	wire _w23984_ ;
	wire _w23985_ ;
	wire _w23986_ ;
	wire _w23987_ ;
	wire _w23988_ ;
	wire _w23989_ ;
	wire _w23990_ ;
	wire _w23991_ ;
	wire _w23992_ ;
	wire _w23993_ ;
	wire _w23994_ ;
	wire _w23995_ ;
	wire _w23996_ ;
	wire _w23997_ ;
	wire _w23998_ ;
	wire _w23999_ ;
	wire _w24000_ ;
	wire _w24001_ ;
	wire _w24002_ ;
	wire _w24003_ ;
	wire _w24004_ ;
	wire _w24005_ ;
	wire _w24006_ ;
	wire _w24007_ ;
	wire _w24008_ ;
	wire _w24009_ ;
	wire _w24010_ ;
	wire _w24011_ ;
	wire _w24012_ ;
	wire _w24013_ ;
	wire _w24014_ ;
	wire _w24015_ ;
	wire _w24016_ ;
	wire _w24017_ ;
	wire _w24018_ ;
	wire _w24019_ ;
	wire _w24020_ ;
	wire _w24021_ ;
	wire _w24022_ ;
	wire _w24023_ ;
	wire _w24024_ ;
	wire _w24025_ ;
	wire _w24026_ ;
	wire _w24027_ ;
	wire _w24028_ ;
	wire _w24029_ ;
	wire _w24030_ ;
	wire _w24031_ ;
	wire _w24032_ ;
	wire _w24033_ ;
	wire _w24034_ ;
	wire _w24035_ ;
	wire _w24036_ ;
	wire _w24037_ ;
	wire _w24038_ ;
	wire _w24039_ ;
	wire _w24040_ ;
	wire _w24041_ ;
	wire _w24042_ ;
	wire _w24043_ ;
	wire _w24044_ ;
	wire _w24045_ ;
	wire _w24046_ ;
	wire _w24047_ ;
	wire _w24048_ ;
	wire _w24049_ ;
	wire _w24050_ ;
	wire _w24051_ ;
	wire _w24052_ ;
	wire _w24053_ ;
	wire _w24054_ ;
	wire _w24055_ ;
	wire _w24056_ ;
	wire _w24057_ ;
	wire _w24058_ ;
	wire _w24059_ ;
	wire _w24060_ ;
	wire _w24061_ ;
	wire _w24062_ ;
	wire _w24063_ ;
	wire _w24064_ ;
	wire _w24065_ ;
	wire _w24066_ ;
	wire _w24067_ ;
	wire _w24068_ ;
	wire _w24069_ ;
	wire _w24070_ ;
	wire _w24071_ ;
	wire _w24072_ ;
	wire _w24073_ ;
	wire _w24074_ ;
	wire _w24075_ ;
	wire _w24076_ ;
	wire _w24077_ ;
	wire _w24078_ ;
	wire _w24079_ ;
	wire _w24080_ ;
	wire _w24081_ ;
	wire _w24082_ ;
	wire _w24083_ ;
	wire _w24084_ ;
	wire _w24085_ ;
	wire _w24086_ ;
	wire _w24087_ ;
	wire _w24088_ ;
	wire _w24089_ ;
	wire _w24090_ ;
	wire _w24091_ ;
	wire _w24092_ ;
	wire _w24093_ ;
	wire _w24094_ ;
	wire _w24095_ ;
	wire _w24096_ ;
	wire _w24097_ ;
	wire _w24098_ ;
	wire _w24099_ ;
	wire _w24100_ ;
	wire _w24101_ ;
	wire _w24102_ ;
	wire _w24103_ ;
	wire _w24104_ ;
	wire _w24105_ ;
	wire _w24106_ ;
	wire _w24107_ ;
	wire _w24108_ ;
	wire _w24109_ ;
	wire _w24110_ ;
	wire _w24111_ ;
	wire _w24112_ ;
	wire _w24113_ ;
	wire _w24114_ ;
	wire _w24115_ ;
	wire _w24116_ ;
	wire _w24117_ ;
	wire _w24118_ ;
	wire _w24119_ ;
	wire _w24120_ ;
	wire _w24121_ ;
	wire _w24122_ ;
	wire _w24123_ ;
	wire _w24124_ ;
	wire _w24125_ ;
	wire _w24126_ ;
	wire _w24127_ ;
	wire _w24128_ ;
	wire _w24129_ ;
	wire _w24130_ ;
	wire _w24131_ ;
	wire _w24132_ ;
	wire _w24133_ ;
	wire _w24134_ ;
	wire _w24135_ ;
	wire _w24136_ ;
	wire _w24137_ ;
	wire _w24138_ ;
	wire _w24139_ ;
	wire _w24140_ ;
	wire _w24141_ ;
	wire _w24142_ ;
	wire _w24143_ ;
	wire _w24144_ ;
	wire _w24145_ ;
	wire _w24146_ ;
	wire _w24147_ ;
	wire _w24148_ ;
	wire _w24149_ ;
	wire _w24150_ ;
	wire _w24151_ ;
	wire _w24152_ ;
	wire _w24153_ ;
	wire _w24154_ ;
	wire _w24155_ ;
	wire _w24156_ ;
	wire _w24157_ ;
	wire _w24158_ ;
	wire _w24159_ ;
	wire _w24160_ ;
	wire _w24161_ ;
	wire _w24162_ ;
	wire _w24163_ ;
	wire _w24164_ ;
	wire _w24165_ ;
	wire _w24166_ ;
	wire _w24167_ ;
	wire _w24168_ ;
	wire _w24169_ ;
	wire _w24170_ ;
	wire _w24171_ ;
	wire _w24172_ ;
	wire _w24173_ ;
	wire _w24174_ ;
	wire _w24175_ ;
	wire _w24176_ ;
	wire _w24177_ ;
	wire _w24178_ ;
	wire _w24179_ ;
	wire _w24180_ ;
	wire _w24181_ ;
	wire _w24182_ ;
	wire _w24183_ ;
	wire _w24184_ ;
	wire _w24185_ ;
	wire _w24186_ ;
	wire _w24187_ ;
	wire _w24188_ ;
	wire _w24189_ ;
	wire _w24190_ ;
	wire _w24191_ ;
	wire _w24192_ ;
	wire _w24193_ ;
	wire _w24194_ ;
	wire _w24195_ ;
	wire _w24196_ ;
	wire _w24197_ ;
	wire _w24198_ ;
	wire _w24199_ ;
	wire _w24200_ ;
	wire _w24201_ ;
	wire _w24202_ ;
	wire _w24203_ ;
	wire _w24204_ ;
	wire _w24205_ ;
	wire _w24206_ ;
	wire _w24207_ ;
	wire _w24208_ ;
	wire _w24209_ ;
	wire _w24210_ ;
	wire _w24211_ ;
	wire _w24212_ ;
	wire _w24213_ ;
	wire _w24214_ ;
	wire _w24215_ ;
	wire _w24216_ ;
	wire _w24217_ ;
	wire _w24218_ ;
	wire _w24219_ ;
	wire _w24220_ ;
	wire _w24221_ ;
	wire _w24222_ ;
	wire _w24223_ ;
	wire _w24224_ ;
	wire _w24225_ ;
	wire _w24226_ ;
	wire _w24227_ ;
	wire _w24228_ ;
	wire _w24229_ ;
	wire _w24230_ ;
	wire _w24231_ ;
	wire _w24232_ ;
	wire _w24233_ ;
	wire _w24234_ ;
	wire _w24235_ ;
	wire _w24236_ ;
	wire _w24237_ ;
	wire _w24238_ ;
	wire _w24239_ ;
	wire _w24240_ ;
	wire _w24241_ ;
	wire _w24242_ ;
	wire _w24243_ ;
	wire _w24244_ ;
	wire _w24245_ ;
	wire _w24246_ ;
	wire _w24247_ ;
	wire _w24248_ ;
	wire _w24249_ ;
	wire _w24250_ ;
	wire _w24251_ ;
	wire _w24252_ ;
	wire _w24253_ ;
	wire _w24254_ ;
	wire _w24255_ ;
	wire _w24256_ ;
	wire _w24257_ ;
	wire _w24258_ ;
	wire _w24259_ ;
	wire _w24260_ ;
	wire _w24261_ ;
	wire _w24262_ ;
	wire _w24263_ ;
	wire _w24264_ ;
	wire _w24265_ ;
	wire _w24266_ ;
	wire _w24267_ ;
	wire _w24268_ ;
	wire _w24269_ ;
	wire _w24270_ ;
	wire _w24271_ ;
	wire _w24272_ ;
	wire _w24273_ ;
	wire _w24274_ ;
	wire _w24275_ ;
	wire _w24276_ ;
	wire _w24277_ ;
	wire _w24278_ ;
	wire _w24279_ ;
	wire _w24280_ ;
	wire _w24281_ ;
	wire _w24282_ ;
	wire _w24283_ ;
	wire _w24284_ ;
	wire _w24285_ ;
	wire _w24286_ ;
	wire _w24287_ ;
	wire _w24288_ ;
	wire _w24289_ ;
	wire _w24290_ ;
	wire _w24291_ ;
	wire _w24292_ ;
	wire _w24293_ ;
	wire _w24294_ ;
	wire _w24295_ ;
	wire _w24296_ ;
	wire _w24297_ ;
	wire _w24298_ ;
	wire _w24299_ ;
	wire _w24300_ ;
	wire _w24301_ ;
	wire _w24302_ ;
	wire _w24303_ ;
	wire _w24304_ ;
	wire _w24305_ ;
	wire _w24306_ ;
	wire _w24307_ ;
	wire _w24308_ ;
	wire _w24309_ ;
	wire _w24310_ ;
	wire _w24311_ ;
	wire _w24312_ ;
	wire _w24313_ ;
	wire _w24314_ ;
	wire _w24315_ ;
	wire _w24316_ ;
	wire _w24317_ ;
	wire _w24318_ ;
	wire _w24319_ ;
	wire _w24320_ ;
	wire _w24321_ ;
	wire _w24322_ ;
	wire _w24323_ ;
	wire _w24324_ ;
	wire _w24325_ ;
	wire _w24326_ ;
	wire _w24327_ ;
	wire _w24328_ ;
	wire _w24329_ ;
	wire _w24330_ ;
	wire _w24331_ ;
	wire _w24332_ ;
	wire _w24333_ ;
	wire _w24334_ ;
	wire _w24335_ ;
	wire _w24336_ ;
	wire _w24337_ ;
	wire _w24338_ ;
	wire _w24339_ ;
	wire _w24340_ ;
	wire _w24341_ ;
	wire _w24342_ ;
	wire _w24343_ ;
	wire _w24344_ ;
	wire _w24345_ ;
	wire _w24346_ ;
	wire _w24347_ ;
	wire _w24348_ ;
	wire _w24349_ ;
	wire _w24350_ ;
	wire _w24351_ ;
	wire _w24352_ ;
	wire _w24353_ ;
	wire _w24354_ ;
	wire _w24355_ ;
	wire _w24356_ ;
	wire _w24357_ ;
	wire _w24358_ ;
	wire _w24359_ ;
	wire _w24360_ ;
	wire _w24361_ ;
	wire _w24362_ ;
	wire _w24363_ ;
	wire _w24364_ ;
	wire _w24365_ ;
	wire _w24366_ ;
	wire _w24367_ ;
	wire _w24368_ ;
	wire _w24369_ ;
	wire _w24370_ ;
	wire _w24371_ ;
	wire _w24372_ ;
	wire _w24373_ ;
	wire _w24374_ ;
	wire _w24375_ ;
	wire _w24376_ ;
	wire _w24377_ ;
	wire _w24378_ ;
	wire _w24379_ ;
	wire _w24380_ ;
	wire _w24381_ ;
	wire _w24382_ ;
	wire _w24383_ ;
	wire _w24384_ ;
	wire _w24385_ ;
	wire _w24386_ ;
	wire _w24387_ ;
	wire _w24388_ ;
	wire _w24389_ ;
	wire _w24390_ ;
	wire _w24391_ ;
	wire _w24392_ ;
	wire _w24393_ ;
	wire _w24394_ ;
	wire _w24395_ ;
	wire _w24396_ ;
	wire _w24397_ ;
	wire _w24398_ ;
	wire _w24399_ ;
	wire _w24400_ ;
	wire _w24401_ ;
	wire _w24402_ ;
	wire _w24403_ ;
	wire _w24404_ ;
	wire _w24405_ ;
	wire _w24406_ ;
	wire _w24407_ ;
	wire _w24408_ ;
	wire _w24409_ ;
	wire _w24410_ ;
	wire _w24411_ ;
	wire _w24412_ ;
	wire _w24413_ ;
	wire _w24414_ ;
	wire _w24415_ ;
	wire _w24416_ ;
	wire _w24417_ ;
	wire _w24418_ ;
	wire _w24419_ ;
	wire _w24420_ ;
	wire _w24421_ ;
	wire _w24422_ ;
	wire _w24423_ ;
	wire _w24424_ ;
	wire _w24425_ ;
	wire _w24426_ ;
	wire _w24427_ ;
	wire _w24428_ ;
	wire _w24429_ ;
	wire _w24430_ ;
	wire _w24431_ ;
	wire _w24432_ ;
	wire _w24433_ ;
	wire _w24434_ ;
	wire _w24435_ ;
	wire _w24436_ ;
	wire _w24437_ ;
	wire _w24438_ ;
	wire _w24439_ ;
	wire _w24440_ ;
	wire _w24441_ ;
	wire _w24442_ ;
	wire _w24443_ ;
	wire _w24444_ ;
	wire _w24445_ ;
	wire _w24446_ ;
	wire _w24447_ ;
	wire _w24448_ ;
	wire _w24449_ ;
	wire _w24450_ ;
	wire _w24451_ ;
	wire _w24452_ ;
	wire _w24453_ ;
	wire _w24454_ ;
	wire _w24455_ ;
	wire _w24456_ ;
	wire _w24457_ ;
	wire _w24458_ ;
	wire _w24459_ ;
	wire _w24460_ ;
	wire _w24461_ ;
	wire _w24462_ ;
	wire _w24463_ ;
	wire _w24464_ ;
	wire _w24465_ ;
	wire _w24466_ ;
	wire _w24467_ ;
	wire _w24468_ ;
	wire _w24469_ ;
	wire _w24470_ ;
	wire _w24471_ ;
	wire _w24472_ ;
	wire _w24473_ ;
	wire _w24474_ ;
	wire _w24475_ ;
	wire _w24476_ ;
	wire _w24477_ ;
	wire _w24478_ ;
	wire _w24479_ ;
	wire _w24480_ ;
	wire _w24481_ ;
	wire _w24482_ ;
	wire _w24483_ ;
	wire _w24484_ ;
	wire _w24485_ ;
	wire _w24486_ ;
	wire _w24487_ ;
	wire _w24488_ ;
	wire _w24489_ ;
	wire _w24490_ ;
	wire _w24491_ ;
	wire _w24492_ ;
	wire _w24493_ ;
	wire _w24494_ ;
	wire _w24495_ ;
	wire _w24496_ ;
	wire _w24497_ ;
	wire _w24498_ ;
	wire _w24499_ ;
	wire _w24500_ ;
	wire _w24501_ ;
	wire _w24502_ ;
	wire _w24503_ ;
	wire _w24504_ ;
	wire _w24505_ ;
	wire _w24506_ ;
	wire _w24507_ ;
	wire _w24508_ ;
	wire _w24509_ ;
	wire _w24510_ ;
	wire _w24511_ ;
	wire _w24512_ ;
	wire _w24513_ ;
	wire _w24514_ ;
	wire _w24515_ ;
	wire _w24516_ ;
	wire _w24517_ ;
	wire _w24518_ ;
	wire _w24519_ ;
	wire _w24520_ ;
	wire _w24521_ ;
	wire _w24522_ ;
	wire _w24523_ ;
	wire _w24524_ ;
	wire _w24525_ ;
	wire _w24526_ ;
	wire _w24527_ ;
	wire _w24528_ ;
	wire _w24529_ ;
	wire _w24530_ ;
	wire _w24531_ ;
	wire _w24532_ ;
	wire _w24533_ ;
	wire _w24534_ ;
	wire _w24535_ ;
	wire _w24536_ ;
	wire _w24537_ ;
	wire _w24538_ ;
	wire _w24539_ ;
	wire _w24540_ ;
	wire _w24541_ ;
	wire _w24542_ ;
	wire _w24543_ ;
	wire _w24544_ ;
	wire _w24545_ ;
	wire _w24546_ ;
	wire _w24547_ ;
	wire _w24548_ ;
	wire _w24549_ ;
	wire _w24550_ ;
	wire _w24551_ ;
	wire _w24552_ ;
	wire _w24553_ ;
	wire _w24554_ ;
	wire _w24555_ ;
	wire _w24556_ ;
	wire _w24557_ ;
	wire _w24558_ ;
	wire _w24559_ ;
	wire _w24560_ ;
	wire _w24561_ ;
	wire _w24562_ ;
	wire _w24563_ ;
	wire _w24564_ ;
	wire _w24565_ ;
	wire _w24566_ ;
	wire _w24567_ ;
	wire _w24568_ ;
	wire _w24569_ ;
	wire _w24570_ ;
	wire _w24571_ ;
	wire _w24572_ ;
	wire _w24573_ ;
	wire _w24574_ ;
	wire _w24575_ ;
	wire _w24576_ ;
	wire _w24577_ ;
	wire _w24578_ ;
	wire _w24579_ ;
	wire _w24580_ ;
	wire _w24581_ ;
	wire _w24582_ ;
	wire _w24583_ ;
	wire _w24584_ ;
	wire _w24585_ ;
	wire _w24586_ ;
	wire _w24587_ ;
	wire _w24588_ ;
	wire _w24589_ ;
	wire _w24590_ ;
	wire _w24591_ ;
	wire _w24592_ ;
	wire _w24593_ ;
	wire _w24594_ ;
	wire _w24595_ ;
	wire _w24596_ ;
	wire _w24597_ ;
	wire _w24598_ ;
	wire _w24599_ ;
	wire _w24600_ ;
	wire _w24601_ ;
	wire _w24602_ ;
	wire _w24603_ ;
	wire _w24604_ ;
	wire _w24605_ ;
	wire _w24606_ ;
	wire _w24607_ ;
	wire _w24608_ ;
	wire _w24609_ ;
	wire _w24610_ ;
	wire _w24611_ ;
	wire _w24612_ ;
	wire _w24613_ ;
	wire _w24614_ ;
	wire _w24615_ ;
	wire _w24616_ ;
	wire _w24617_ ;
	wire _w24618_ ;
	wire _w24619_ ;
	wire _w24620_ ;
	wire _w24621_ ;
	wire _w24622_ ;
	wire _w24623_ ;
	wire _w24624_ ;
	wire _w24625_ ;
	wire _w24626_ ;
	wire _w24627_ ;
	wire _w24628_ ;
	wire _w24629_ ;
	wire _w24630_ ;
	wire _w24631_ ;
	wire _w24632_ ;
	wire _w24633_ ;
	wire _w24634_ ;
	wire _w24635_ ;
	wire _w24636_ ;
	wire _w24637_ ;
	wire _w24638_ ;
	wire _w24639_ ;
	wire _w24640_ ;
	wire _w24641_ ;
	wire _w24642_ ;
	wire _w24643_ ;
	wire _w24644_ ;
	wire _w24645_ ;
	wire _w24646_ ;
	wire _w24647_ ;
	wire _w24648_ ;
	wire _w24649_ ;
	wire _w24650_ ;
	wire _w24651_ ;
	wire _w24652_ ;
	wire _w24653_ ;
	wire _w24654_ ;
	wire _w24655_ ;
	wire _w24656_ ;
	wire _w24657_ ;
	wire _w24658_ ;
	wire _w24659_ ;
	wire _w24660_ ;
	wire _w24661_ ;
	wire _w24662_ ;
	wire _w24663_ ;
	wire _w24664_ ;
	wire _w24665_ ;
	wire _w24666_ ;
	wire _w24667_ ;
	wire _w24668_ ;
	wire _w24669_ ;
	wire _w24670_ ;
	wire _w24671_ ;
	wire _w24672_ ;
	wire _w24673_ ;
	wire _w24674_ ;
	wire _w24675_ ;
	wire _w24676_ ;
	wire _w24677_ ;
	wire _w24678_ ;
	wire _w24679_ ;
	wire _w24680_ ;
	wire _w24681_ ;
	wire _w24682_ ;
	wire _w24683_ ;
	wire _w24684_ ;
	wire _w24685_ ;
	wire _w24686_ ;
	wire _w24687_ ;
	wire _w24688_ ;
	wire _w24689_ ;
	wire _w24690_ ;
	wire _w24691_ ;
	wire _w24692_ ;
	wire _w24693_ ;
	wire _w24694_ ;
	wire _w24695_ ;
	wire _w24696_ ;
	wire _w24697_ ;
	wire _w24698_ ;
	wire _w24699_ ;
	wire _w24700_ ;
	wire _w24701_ ;
	wire _w24702_ ;
	wire _w24703_ ;
	wire _w24704_ ;
	wire _w24705_ ;
	wire _w24706_ ;
	wire _w24707_ ;
	wire _w24708_ ;
	wire _w24709_ ;
	wire _w24710_ ;
	wire _w24711_ ;
	wire _w24712_ ;
	wire _w24713_ ;
	wire _w24714_ ;
	wire _w24715_ ;
	wire _w24716_ ;
	wire _w24717_ ;
	wire _w24718_ ;
	wire _w24719_ ;
	wire _w24720_ ;
	wire _w24721_ ;
	wire _w24722_ ;
	wire _w24723_ ;
	wire _w24724_ ;
	wire _w24725_ ;
	wire _w24726_ ;
	wire _w24727_ ;
	wire _w24728_ ;
	wire _w24729_ ;
	wire _w24730_ ;
	wire _w24731_ ;
	wire _w24732_ ;
	wire _w24733_ ;
	wire _w24734_ ;
	wire _w24735_ ;
	wire _w24736_ ;
	wire _w24737_ ;
	wire _w24738_ ;
	wire _w24739_ ;
	wire _w24740_ ;
	wire _w24741_ ;
	wire _w24742_ ;
	wire _w24743_ ;
	wire _w24744_ ;
	wire _w24745_ ;
	wire _w24746_ ;
	wire _w24747_ ;
	wire _w24748_ ;
	wire _w24749_ ;
	wire _w24750_ ;
	wire _w24751_ ;
	wire _w24752_ ;
	wire _w24753_ ;
	wire _w24754_ ;
	wire _w24755_ ;
	wire _w24756_ ;
	wire _w24757_ ;
	wire _w24758_ ;
	wire _w24759_ ;
	wire _w24760_ ;
	wire _w24761_ ;
	wire _w24762_ ;
	wire _w24763_ ;
	wire _w24764_ ;
	wire _w24765_ ;
	wire _w24766_ ;
	wire _w24767_ ;
	wire _w24768_ ;
	wire _w24769_ ;
	wire _w24770_ ;
	wire _w24771_ ;
	wire _w24772_ ;
	wire _w24773_ ;
	wire _w24774_ ;
	wire _w24775_ ;
	wire _w24776_ ;
	wire _w24777_ ;
	wire _w24778_ ;
	wire _w24779_ ;
	wire _w24780_ ;
	wire _w24781_ ;
	wire _w24782_ ;
	wire _w24783_ ;
	wire _w24784_ ;
	wire _w24785_ ;
	wire _w24786_ ;
	wire _w24787_ ;
	wire _w24788_ ;
	wire _w24789_ ;
	wire _w24790_ ;
	wire _w24791_ ;
	wire _w24792_ ;
	wire _w24793_ ;
	wire _w24794_ ;
	wire _w24795_ ;
	wire _w24796_ ;
	wire _w24797_ ;
	wire _w24798_ ;
	wire _w24799_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\clkc_CLKOUT_reg/NET0131 ,
		\clkc_ckr_reg_DO_reg[15]/NET0131 ,
		_w4047_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\bdma_BSreq_reg/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4048_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport1_rxctl_RSreq_reg/NET0131 ,
		_w4049_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_txctl_TSreq_reg/NET0131 ,
		_w4050_
	);
	LUT2 #(
		.INIT('h4)
	) name4 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport0_rxctl_RSreq_reg/NET0131 ,
		_w4051_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w4050_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sport1_txctl_TSreq_reg/NET0131 ,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		_w4052_,
		_w4053_,
		_w4054_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		_w4049_,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\idma_DSreq_reg/NET0131 ,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		_w4048_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h4)
	) name11 (
		\idma_IDMA_boot_reg/NET0131_reg_syn_10 ,
		\idma_IDMA_boot_reg/NET0131_reg_syn_2 ,
		_w4058_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\idma_IDMA_boot_reg/NET0131_reg_syn_10 ,
		\idma_IDMA_boot_reg/NET0131_reg_syn_8 ,
		_w4059_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w4058_,
		_w4059_,
		_w4060_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		\bdma_BDMA_boot_reg/NET0131_reg_syn_10 ,
		\bdma_BDMA_boot_reg/NET0131_reg_syn_2 ,
		_w4061_
	);
	LUT2 #(
		.INIT('h8)
	) name15 (
		\bdma_BDMA_boot_reg/NET0131_reg_syn_10 ,
		\bdma_BDMA_boot_reg/NET0131_reg_syn_8 ,
		_w4062_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w4061_,
		_w4062_,
		_w4063_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		_w4060_,
		_w4063_,
		_w4064_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\bdma_BM_cyc_reg/P0001 ,
		\core_c_psq_ECYC_reg/P0001 ,
		_w4065_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_2 ,
		_w4066_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\memc_EXTC_Eg_reg/NET0131_reg_syn_10 ,
		\memc_EXTC_Eg_reg/NET0131_reg_syn_8 ,
		_w4067_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w4066_,
		_w4067_,
		_w4068_
	);
	LUT2 #(
		.INIT('h8)
	) name22 (
		\core_c_psq_PCS_reg[2]/NET0131 ,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		\core_c_psq_PCS_reg[15]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w4070_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w4069_,
		_w4070_,
		_w4071_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\clkc_Awake_reg/NET0131 ,
		\clkc_STBY_reg/NET0131 ,
		_w4072_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\clkc_STBY_reg/NET0131 ,
		\core_c_psq_TRAP_R_L_reg/NET0131 ,
		_w4073_
	);
	LUT2 #(
		.INIT('h4)
	) name27 (
		\sice_GOICE_syn_reg/P0001 ,
		_w4073_,
		_w4074_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		_w4072_,
		_w4074_,
		_w4075_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		\core_c_psq_PCS_reg[4]/NET0131 ,
		_w4075_,
		_w4076_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		\core_c_psq_PCS_reg[10]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w4077_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		\core_c_psq_MGNT_reg/NET0131 ,
		_w4078_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		\core_c_psq_PCS_reg[11]/NET0131 ,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\memc_LDaST_Eg_reg/NET0131 ,
		_w4080_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		\core_c_psq_PCS_reg[12]/NET0131 ,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		\sice_HALT_E_reg/P0001 ,
		_w4082_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_dec_IDLE_Eg_reg/P0001 ,
		_w4083_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w4082_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w4084_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name39 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4081_,
		_w4086_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		_w4085_,
		_w4086_,
		_w4087_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\core_c_psq_PCS_reg[5]/NET0131 ,
		\core_c_psq_PCS_reg[6]/NET0131 ,
		_w4088_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w4079_,
		_w4088_,
		_w4089_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w4087_,
		_w4089_,
		_w4090_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		_w4068_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w4076_,
		_w4077_,
		_w4092_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		_w4091_,
		_w4092_,
		_w4093_
	);
	LUT2 #(
		.INIT('h8)
	) name47 (
		_w4071_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		\auctl_STEAL_reg/NET0131 ,
		\clkc_STBY_reg/NET0131 ,
		_w4095_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w4094_,
		_w4095_,
		_w4096_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w4065_,
		_w4096_,
		_w4097_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w4064_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w4057_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		_w4100_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w4100_,
		_w4101_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\sice_CMRW_reg/NET0131 ,
		_w4102_
	);
	LUT2 #(
		.INIT('h8)
	) name56 (
		_w4101_,
		_w4102_,
		_w4103_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\core_c_dec_accCM_E_reg/NET0131 ,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h4)
	) name58 (
		\core_c_psq_SRST_reg/P0001 ,
		_w4064_,
		_w4105_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		_w4105_,
		_w4106_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS2or3_reg/NET0131 ,
		_w4107_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		\core_c_psq_PCS_reg[12]/NET0131 ,
		_w4107_,
		_w4108_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4108_,
		_w4109_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\core_c_psq_PCS_reg[2]/NET0131 ,
		_w4110_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w4109_,
		_w4110_,
		_w4111_
	);
	LUT2 #(
		.INIT('h4)
	) name65 (
		_w4106_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\core_c_psq_PCS_reg[11]/NET0131 ,
		_w4107_,
		_w4113_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		\sice_HALT_E_reg/P0001 ,
		_w4114_
	);
	LUT2 #(
		.INIT('h4)
	) name68 (
		_w4113_,
		_w4114_,
		_w4115_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		_w4112_,
		_w4115_,
		_w4116_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\sice_GO_NX_reg/NET0131 ,
		_w4094_,
		_w4117_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		_w4116_,
		_w4117_,
		_w4118_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		_w4104_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w4099_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w4117_,
		_w4121_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w4117_,
		_w4122_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w4121_,
		_w4122_,
		_w4123_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w4104_,
		_w4123_,
		_w4124_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w4104_,
		_w4125_
	);
	LUT2 #(
		.INIT('h1)
	) name79 (
		_w4124_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h8)
	) name80 (
		_w4120_,
		_w4126_,
		_w4127_
	);
	LUT2 #(
		.INIT('h4)
	) name81 (
		_w4099_,
		_w4119_,
		_w4128_
	);
	LUT2 #(
		.INIT('h4)
	) name82 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4105_,
		_w4129_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		\core_c_dec_IDLE_Eg_reg/P0001 ,
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		_w4130_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		_w4131_
	);
	LUT2 #(
		.INIT('h4)
	) name85 (
		\core_c_psq_CE_reg/NET0131 ,
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		_w4132_
	);
	LUT2 #(
		.INIT('h8)
	) name86 (
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		_w4132_,
		_w4133_
	);
	LUT2 #(
		.INIT('h8)
	) name87 (
		_w4131_,
		_w4133_,
		_w4134_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w4135_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w4136_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w4135_,
		_w4136_,
		_w4137_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		_w4138_,
		_w4139_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w4139_,
		_w4140_,
		_w4141_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		_w4141_,
		_w4142_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		_w4141_,
		_w4143_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		_w4144_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w4142_,
		_w4144_,
		_w4145_
	);
	LUT2 #(
		.INIT('h4)
	) name99 (
		_w4143_,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		\clkc_Cnt4096_reg/NET0131 ,
		\clkc_Cnt4096_s2_reg/NET0131 ,
		_w4147_
	);
	LUT2 #(
		.INIT('h8)
	) name101 (
		\sport0_regs_AUTO_a_reg[12]/NET0131 ,
		_w4147_,
		_w4148_
	);
	LUT2 #(
		.INIT('h1)
	) name102 (
		\bdma_RST_pin_reg/P0001 ,
		\sice_RCS_reg[1]/NET0131 ,
		_w4149_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		_w4148_,
		_w4149_,
		_w4150_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4150_,
		_w4151_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\core_eu_ec_cun_MV_reg/P0000_reg_syn_2 ,
		_w4151_,
		_w4152_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001 ,
		_w4153_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001 ,
		_w4154_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001 ,
		_w4155_
	);
	LUT2 #(
		.INIT('h8)
	) name109 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001 ,
		_w4156_
	);
	LUT2 #(
		.INIT('h8)
	) name110 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001 ,
		_w4156_,
		_w4157_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		_w4154_,
		_w4155_,
		_w4158_
	);
	LUT2 #(
		.INIT('h8)
	) name112 (
		_w4153_,
		_w4158_,
		_w4159_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		_w4157_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[1]/P0001 ,
		_w4161_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[3]/P0001 ,
		_w4162_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[4]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[5]/P0001 ,
		_w4163_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[6]/P0001 ,
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[7]/P0001 ,
		_w4164_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[8]/P0001 ,
		_w4164_,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name119 (
		_w4162_,
		_w4163_,
		_w4166_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w4161_,
		_w4166_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name121 (
		_w4165_,
		_w4167_,
		_w4168_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		\core_eu_ec_cun_updateMV_C_reg/P0001 ,
		_w4160_,
		_w4169_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		_w4168_,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		\core_eu_ec_cun_MVi_pre_C_reg/P0001 ,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h2)
	) name125 (
		_w4150_,
		_w4171_,
		_w4172_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w4172_,
		_w4173_
	);
	LUT2 #(
		.INIT('h1)
	) name127 (
		_w4152_,
		_w4173_,
		_w4174_
	);
	LUT2 #(
		.INIT('h4)
	) name128 (
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		_w4175_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		_w4176_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		_w4175_,
		_w4176_,
		_w4177_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		_w4174_,
		_w4177_,
		_w4178_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		_w4131_,
		_w4175_,
		_w4179_
	);
	LUT2 #(
		.INIT('h4)
	) name133 (
		_w4174_,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		\core_eu_ec_cun_condOK_CE_reg/P0001 ,
		_w4134_,
		_w4181_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w4146_,
		_w4181_,
		_w4182_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w4178_,
		_w4182_,
		_w4183_
	);
	LUT2 #(
		.INIT('h4)
	) name137 (
		_w4180_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h2)
	) name138 (
		\core_c_dec_Nseq_Ed_reg/P0001 ,
		_w4184_,
		_w4185_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		_w4130_,
		_w4185_,
		_w4186_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4186_,
		_w4187_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4188_
	);
	LUT2 #(
		.INIT('h1)
	) name142 (
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w4189_
	);
	LUT2 #(
		.INIT('h8)
	) name143 (
		_w4188_,
		_w4189_,
		_w4190_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001 ,
		_w4190_,
		_w4191_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w4192_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4193_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h8)
	) name148 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001 ,
		_w4194_,
		_w4195_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4196_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w4192_,
		_w4196_,
		_w4197_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001 ,
		_w4197_,
		_w4198_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w4199_
	);
	LUT2 #(
		.INIT('h8)
	) name153 (
		_w4188_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001 ,
		_w4200_,
		_w4201_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w4193_,
		_w4199_,
		_w4202_
	);
	LUT2 #(
		.INIT('h8)
	) name156 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001 ,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4204_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w4199_,
		_w4204_,
		_w4205_
	);
	LUT2 #(
		.INIT('h8)
	) name159 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001 ,
		_w4205_,
		_w4206_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w4207_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h4)
	) name162 (
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001 ,
		_w4209_,
		_w4210_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w4196_,
		_w4199_,
		_w4211_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001 ,
		_w4211_,
		_w4212_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		_w4188_,
		_w4192_,
		_w4213_
	);
	LUT2 #(
		.INIT('h8)
	) name167 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001 ,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4208_,
		_w4215_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001 ,
		_w4215_,
		_w4216_
	);
	LUT2 #(
		.INIT('h4)
	) name170 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		_w4189_,
		_w4217_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4217_,
		_w4218_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001 ,
		_w4218_,
		_w4219_
	);
	LUT2 #(
		.INIT('h8)
	) name173 (
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w4217_,
		_w4220_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001 ,
		_w4220_,
		_w4221_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		_w4193_,
		_w4207_,
		_w4222_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001 ,
		_w4222_,
		_w4223_
	);
	LUT2 #(
		.INIT('h8)
	) name177 (
		_w4192_,
		_w4204_,
		_w4224_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001 ,
		_w4224_,
		_w4225_
	);
	LUT2 #(
		.INIT('h8)
	) name179 (
		_w4196_,
		_w4207_,
		_w4226_
	);
	LUT2 #(
		.INIT('h8)
	) name180 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001 ,
		_w4226_,
		_w4227_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w4189_,
		_w4204_,
		_w4228_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001 ,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w4191_,
		_w4195_,
		_w4230_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w4198_,
		_w4201_,
		_w4231_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w4203_,
		_w4206_,
		_w4232_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w4212_,
		_w4214_,
		_w4233_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w4223_,
		_w4225_,
		_w4234_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w4227_,
		_w4229_,
		_w4235_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w4234_,
		_w4235_,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		_w4232_,
		_w4233_,
		_w4237_
	);
	LUT2 #(
		.INIT('h8)
	) name191 (
		_w4230_,
		_w4231_,
		_w4238_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w4210_,
		_w4216_,
		_w4239_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w4219_,
		_w4221_,
		_w4240_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		_w4237_,
		_w4238_,
		_w4242_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		_w4236_,
		_w4242_,
		_w4243_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w4241_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name198 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4244_,
		_w4245_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001 ,
		_w4202_,
		_w4246_
	);
	LUT2 #(
		.INIT('h8)
	) name200 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001 ,
		_w4211_,
		_w4247_
	);
	LUT2 #(
		.INIT('h8)
	) name201 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001 ,
		_w4194_,
		_w4248_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001 ,
		_w4224_,
		_w4249_
	);
	LUT2 #(
		.INIT('h8)
	) name203 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001 ,
		_w4205_,
		_w4250_
	);
	LUT2 #(
		.INIT('h8)
	) name204 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001 ,
		_w4226_,
		_w4251_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001 ,
		_w4220_,
		_w4252_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001 ,
		_w4228_,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name207 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001 ,
		_w4197_,
		_w4254_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001 ,
		_w4209_,
		_w4255_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001 ,
		_w4215_,
		_w4256_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001 ,
		_w4218_,
		_w4257_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001 ,
		_w4190_,
		_w4258_
	);
	LUT2 #(
		.INIT('h8)
	) name212 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001 ,
		_w4222_,
		_w4259_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001 ,
		_w4213_,
		_w4260_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001 ,
		_w4200_,
		_w4261_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w4246_,
		_w4247_,
		_w4262_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w4248_,
		_w4249_,
		_w4263_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		_w4250_,
		_w4251_,
		_w4264_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w4253_,
		_w4254_,
		_w4265_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w4258_,
		_w4259_,
		_w4266_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w4260_,
		_w4261_,
		_w4267_
	);
	LUT2 #(
		.INIT('h8)
	) name221 (
		_w4266_,
		_w4267_,
		_w4268_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		_w4264_,
		_w4265_,
		_w4269_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		_w4262_,
		_w4263_,
		_w4270_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w4252_,
		_w4255_,
		_w4271_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w4256_,
		_w4257_,
		_w4272_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		_w4271_,
		_w4272_,
		_w4273_
	);
	LUT2 #(
		.INIT('h8)
	) name227 (
		_w4269_,
		_w4270_,
		_w4274_
	);
	LUT2 #(
		.INIT('h8)
	) name228 (
		_w4268_,
		_w4274_,
		_w4275_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w4273_,
		_w4275_,
		_w4276_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4276_,
		_w4277_
	);
	LUT2 #(
		.INIT('h8)
	) name231 (
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		_w4174_,
		_w4278_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		\core_eu_ec_cun_TERM_E_reg[2]/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[3]/P0001 ,
		_w4279_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		_w4174_,
		_w4280_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		_w4279_,
		_w4281_
	);
	LUT2 #(
		.INIT('h4)
	) name235 (
		_w4278_,
		_w4281_,
		_w4282_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		_w4280_,
		_w4282_,
		_w4283_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		\core_c_psq_CE_reg/NET0131 ,
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		_w4284_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		_w4284_,
		_w4285_
	);
	LUT2 #(
		.INIT('h8)
	) name239 (
		_w4279_,
		_w4285_,
		_w4286_
	);
	LUT2 #(
		.INIT('h2)
	) name240 (
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		_w4138_,
		_w4287_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		_w4288_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w4287_,
		_w4288_,
		_w4289_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		_w4289_,
		_w4290_
	);
	LUT2 #(
		.INIT('h2)
	) name244 (
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		_w4289_,
		_w4291_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\core_eu_ec_cun_TERM_E_reg[2]/P0001 ,
		\core_eu_ec_cun_TERM_E_reg[3]/P0001 ,
		_w4292_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w4290_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h4)
	) name247 (
		_w4291_,
		_w4293_,
		_w4294_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		\core_eu_ec_cun_termOK_CE_reg/P0001 ,
		_w4286_,
		_w4295_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		_w4294_,
		_w4295_,
		_w4296_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		_w4283_,
		_w4296_,
		_w4297_
	);
	LUT2 #(
		.INIT('h8)
	) name251 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001 ,
		_w4190_,
		_w4298_
	);
	LUT2 #(
		.INIT('h8)
	) name252 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001 ,
		_w4194_,
		_w4299_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001 ,
		_w4197_,
		_w4300_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001 ,
		_w4200_,
		_w4301_
	);
	LUT2 #(
		.INIT('h8)
	) name255 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001 ,
		_w4202_,
		_w4302_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001 ,
		_w4205_,
		_w4303_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001 ,
		_w4209_,
		_w4304_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001 ,
		_w4211_,
		_w4305_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001 ,
		_w4213_,
		_w4306_
	);
	LUT2 #(
		.INIT('h8)
	) name260 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001 ,
		_w4215_,
		_w4307_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001 ,
		_w4218_,
		_w4308_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001 ,
		_w4220_,
		_w4309_
	);
	LUT2 #(
		.INIT('h8)
	) name263 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001 ,
		_w4222_,
		_w4310_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001 ,
		_w4224_,
		_w4311_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001 ,
		_w4226_,
		_w4312_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001 ,
		_w4228_,
		_w4313_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w4298_,
		_w4299_,
		_w4314_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w4300_,
		_w4301_,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w4302_,
		_w4303_,
		_w4316_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w4305_,
		_w4306_,
		_w4317_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		_w4310_,
		_w4311_,
		_w4318_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w4312_,
		_w4313_,
		_w4319_
	);
	LUT2 #(
		.INIT('h8)
	) name273 (
		_w4318_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w4316_,
		_w4317_,
		_w4321_
	);
	LUT2 #(
		.INIT('h8)
	) name275 (
		_w4314_,
		_w4315_,
		_w4322_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w4304_,
		_w4307_,
		_w4323_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w4308_,
		_w4309_,
		_w4324_
	);
	LUT2 #(
		.INIT('h8)
	) name278 (
		_w4323_,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h8)
	) name279 (
		_w4321_,
		_w4322_,
		_w4326_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		_w4320_,
		_w4326_,
		_w4327_
	);
	LUT2 #(
		.INIT('h8)
	) name281 (
		_w4325_,
		_w4327_,
		_w4328_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4328_,
		_w4329_
	);
	LUT2 #(
		.INIT('h8)
	) name283 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001 ,
		_w4205_,
		_w4330_
	);
	LUT2 #(
		.INIT('h8)
	) name284 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001 ,
		_w4194_,
		_w4331_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001 ,
		_w4197_,
		_w4332_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001 ,
		_w4222_,
		_w4333_
	);
	LUT2 #(
		.INIT('h8)
	) name287 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001 ,
		_w4226_,
		_w4334_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001 ,
		_w4213_,
		_w4335_
	);
	LUT2 #(
		.INIT('h8)
	) name289 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001 ,
		_w4215_,
		_w4336_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001 ,
		_w4200_,
		_w4337_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001 ,
		_w4190_,
		_w4338_
	);
	LUT2 #(
		.INIT('h8)
	) name292 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001 ,
		_w4218_,
		_w4339_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001 ,
		_w4209_,
		_w4340_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001 ,
		_w4220_,
		_w4341_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001 ,
		_w4211_,
		_w4342_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001 ,
		_w4228_,
		_w4343_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001 ,
		_w4202_,
		_w4344_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001 ,
		_w4224_,
		_w4345_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w4330_,
		_w4331_,
		_w4346_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w4332_,
		_w4333_,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w4334_,
		_w4335_,
		_w4348_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w4337_,
		_w4338_,
		_w4349_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		_w4342_,
		_w4343_,
		_w4350_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w4344_,
		_w4345_,
		_w4351_
	);
	LUT2 #(
		.INIT('h8)
	) name305 (
		_w4350_,
		_w4351_,
		_w4352_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		_w4348_,
		_w4349_,
		_w4353_
	);
	LUT2 #(
		.INIT('h8)
	) name307 (
		_w4346_,
		_w4347_,
		_w4354_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w4336_,
		_w4339_,
		_w4355_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w4340_,
		_w4341_,
		_w4356_
	);
	LUT2 #(
		.INIT('h8)
	) name310 (
		_w4355_,
		_w4356_,
		_w4357_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		_w4353_,
		_w4354_,
		_w4358_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		_w4352_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h8)
	) name313 (
		_w4357_,
		_w4359_,
		_w4360_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4360_,
		_w4361_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001 ,
		_w4226_,
		_w4362_
	);
	LUT2 #(
		.INIT('h8)
	) name316 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001 ,
		_w4222_,
		_w4363_
	);
	LUT2 #(
		.INIT('h8)
	) name317 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001 ,
		_w4211_,
		_w4364_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001 ,
		_w4213_,
		_w4365_
	);
	LUT2 #(
		.INIT('h8)
	) name319 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001 ,
		_w4228_,
		_w4366_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001 ,
		_w4197_,
		_w4367_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001 ,
		_w4209_,
		_w4368_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001 ,
		_w4194_,
		_w4369_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001 ,
		_w4200_,
		_w4370_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001 ,
		_w4215_,
		_w4371_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001 ,
		_w4218_,
		_w4372_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001 ,
		_w4220_,
		_w4373_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001 ,
		_w4224_,
		_w4374_
	);
	LUT2 #(
		.INIT('h8)
	) name328 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001 ,
		_w4190_,
		_w4375_
	);
	LUT2 #(
		.INIT('h8)
	) name329 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001 ,
		_w4202_,
		_w4376_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001 ,
		_w4205_,
		_w4377_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w4362_,
		_w4363_,
		_w4378_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w4364_,
		_w4365_,
		_w4379_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w4366_,
		_w4367_,
		_w4380_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w4369_,
		_w4370_,
		_w4381_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w4374_,
		_w4375_,
		_w4382_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w4376_,
		_w4377_,
		_w4383_
	);
	LUT2 #(
		.INIT('h8)
	) name337 (
		_w4382_,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w4380_,
		_w4381_,
		_w4385_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		_w4378_,
		_w4379_,
		_w4386_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w4368_,
		_w4371_,
		_w4387_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w4372_,
		_w4373_,
		_w4388_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		_w4387_,
		_w4388_,
		_w4389_
	);
	LUT2 #(
		.INIT('h8)
	) name343 (
		_w4385_,
		_w4386_,
		_w4390_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		_w4384_,
		_w4390_,
		_w4391_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		_w4389_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w4392_,
		_w4393_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w4392_,
		_w4394_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001 ,
		_w4228_,
		_w4395_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001 ,
		_w4213_,
		_w4396_
	);
	LUT2 #(
		.INIT('h8)
	) name350 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001 ,
		_w4211_,
		_w4397_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001 ,
		_w4194_,
		_w4398_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001 ,
		_w4222_,
		_w4399_
	);
	LUT2 #(
		.INIT('h8)
	) name353 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001 ,
		_w4197_,
		_w4400_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001 ,
		_w4220_,
		_w4401_
	);
	LUT2 #(
		.INIT('h8)
	) name355 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001 ,
		_w4205_,
		_w4402_
	);
	LUT2 #(
		.INIT('h8)
	) name356 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001 ,
		_w4226_,
		_w4403_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001 ,
		_w4209_,
		_w4404_
	);
	LUT2 #(
		.INIT('h8)
	) name358 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001 ,
		_w4215_,
		_w4405_
	);
	LUT2 #(
		.INIT('h8)
	) name359 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001 ,
		_w4218_,
		_w4406_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001 ,
		_w4224_,
		_w4407_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001 ,
		_w4202_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001 ,
		_w4190_,
		_w4409_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001 ,
		_w4200_,
		_w4410_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w4395_,
		_w4396_,
		_w4411_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w4397_,
		_w4398_,
		_w4412_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w4399_,
		_w4400_,
		_w4413_
	);
	LUT2 #(
		.INIT('h1)
	) name367 (
		_w4402_,
		_w4403_,
		_w4414_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w4407_,
		_w4408_,
		_w4415_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w4409_,
		_w4410_,
		_w4416_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		_w4415_,
		_w4416_,
		_w4417_
	);
	LUT2 #(
		.INIT('h8)
	) name371 (
		_w4413_,
		_w4414_,
		_w4418_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		_w4411_,
		_w4412_,
		_w4419_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w4401_,
		_w4404_,
		_w4420_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w4405_,
		_w4406_,
		_w4421_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		_w4420_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h8)
	) name376 (
		_w4418_,
		_w4419_,
		_w4423_
	);
	LUT2 #(
		.INIT('h8)
	) name377 (
		_w4417_,
		_w4423_,
		_w4424_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		_w4422_,
		_w4424_,
		_w4425_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001 ,
		_w4202_,
		_w4427_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001 ,
		_w4211_,
		_w4428_
	);
	LUT2 #(
		.INIT('h8)
	) name382 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001 ,
		_w4194_,
		_w4429_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001 ,
		_w4224_,
		_w4430_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001 ,
		_w4205_,
		_w4431_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001 ,
		_w4226_,
		_w4432_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001 ,
		_w4220_,
		_w4433_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001 ,
		_w4228_,
		_w4434_
	);
	LUT2 #(
		.INIT('h8)
	) name388 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001 ,
		_w4197_,
		_w4435_
	);
	LUT2 #(
		.INIT('h8)
	) name389 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001 ,
		_w4209_,
		_w4436_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001 ,
		_w4215_,
		_w4437_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001 ,
		_w4218_,
		_w4438_
	);
	LUT2 #(
		.INIT('h8)
	) name392 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001 ,
		_w4190_,
		_w4439_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001 ,
		_w4222_,
		_w4440_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001 ,
		_w4213_,
		_w4441_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001 ,
		_w4200_,
		_w4442_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w4427_,
		_w4428_,
		_w4443_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w4429_,
		_w4430_,
		_w4444_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w4431_,
		_w4432_,
		_w4445_
	);
	LUT2 #(
		.INIT('h1)
	) name399 (
		_w4434_,
		_w4435_,
		_w4446_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w4439_,
		_w4440_,
		_w4447_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w4441_,
		_w4442_,
		_w4448_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		_w4447_,
		_w4448_,
		_w4449_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		_w4445_,
		_w4446_,
		_w4450_
	);
	LUT2 #(
		.INIT('h8)
	) name404 (
		_w4443_,
		_w4444_,
		_w4451_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w4433_,
		_w4436_,
		_w4452_
	);
	LUT2 #(
		.INIT('h1)
	) name406 (
		_w4437_,
		_w4438_,
		_w4453_
	);
	LUT2 #(
		.INIT('h8)
	) name407 (
		_w4452_,
		_w4453_,
		_w4454_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		_w4450_,
		_w4451_,
		_w4455_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w4449_,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		_w4454_,
		_w4456_,
		_w4457_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h8)
	) name412 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001 ,
		_w4190_,
		_w4459_
	);
	LUT2 #(
		.INIT('h8)
	) name413 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001 ,
		_w4194_,
		_w4460_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001 ,
		_w4197_,
		_w4461_
	);
	LUT2 #(
		.INIT('h8)
	) name415 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001 ,
		_w4200_,
		_w4462_
	);
	LUT2 #(
		.INIT('h8)
	) name416 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001 ,
		_w4202_,
		_w4463_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001 ,
		_w4205_,
		_w4464_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001 ,
		_w4209_,
		_w4465_
	);
	LUT2 #(
		.INIT('h8)
	) name419 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001 ,
		_w4211_,
		_w4466_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001 ,
		_w4213_,
		_w4467_
	);
	LUT2 #(
		.INIT('h8)
	) name421 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001 ,
		_w4215_,
		_w4468_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001 ,
		_w4218_,
		_w4469_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001 ,
		_w4220_,
		_w4470_
	);
	LUT2 #(
		.INIT('h8)
	) name424 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001 ,
		_w4222_,
		_w4471_
	);
	LUT2 #(
		.INIT('h8)
	) name425 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001 ,
		_w4224_,
		_w4472_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001 ,
		_w4226_,
		_w4473_
	);
	LUT2 #(
		.INIT('h8)
	) name427 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001 ,
		_w4228_,
		_w4474_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w4459_,
		_w4460_,
		_w4475_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w4461_,
		_w4462_,
		_w4476_
	);
	LUT2 #(
		.INIT('h1)
	) name430 (
		_w4463_,
		_w4464_,
		_w4477_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w4466_,
		_w4467_,
		_w4478_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w4471_,
		_w4472_,
		_w4479_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w4473_,
		_w4474_,
		_w4480_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		_w4479_,
		_w4480_,
		_w4481_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		_w4477_,
		_w4478_,
		_w4482_
	);
	LUT2 #(
		.INIT('h8)
	) name436 (
		_w4475_,
		_w4476_,
		_w4483_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w4465_,
		_w4468_,
		_w4484_
	);
	LUT2 #(
		.INIT('h1)
	) name438 (
		_w4469_,
		_w4470_,
		_w4485_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		_w4484_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h8)
	) name440 (
		_w4482_,
		_w4483_,
		_w4487_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		_w4481_,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		_w4486_,
		_w4488_,
		_w4489_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4489_,
		_w4490_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001 ,
		_w4213_,
		_w4491_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001 ,
		_w4190_,
		_w4492_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001 ,
		_w4228_,
		_w4493_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001 ,
		_w4197_,
		_w4494_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001 ,
		_w4200_,
		_w4495_
	);
	LUT2 #(
		.INIT('h8)
	) name449 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001 ,
		_w4194_,
		_w4496_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001 ,
		_w4220_,
		_w4497_
	);
	LUT2 #(
		.INIT('h8)
	) name451 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001 ,
		_w4211_,
		_w4498_
	);
	LUT2 #(
		.INIT('h8)
	) name452 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001 ,
		_w4224_,
		_w4499_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001 ,
		_w4209_,
		_w4500_
	);
	LUT2 #(
		.INIT('h8)
	) name454 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001 ,
		_w4215_,
		_w4501_
	);
	LUT2 #(
		.INIT('h8)
	) name455 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001 ,
		_w4218_,
		_w4502_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001 ,
		_w4222_,
		_w4503_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001 ,
		_w4202_,
		_w4504_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001 ,
		_w4205_,
		_w4505_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001 ,
		_w4226_,
		_w4506_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w4491_,
		_w4492_,
		_w4507_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w4493_,
		_w4494_,
		_w4508_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w4495_,
		_w4496_,
		_w4509_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w4498_,
		_w4499_,
		_w4510_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w4503_,
		_w4504_,
		_w4511_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		_w4505_,
		_w4506_,
		_w4512_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		_w4511_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h8)
	) name467 (
		_w4509_,
		_w4510_,
		_w4514_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		_w4507_,
		_w4508_,
		_w4515_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w4497_,
		_w4500_,
		_w4516_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w4501_,
		_w4502_,
		_w4517_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		_w4516_,
		_w4517_,
		_w4518_
	);
	LUT2 #(
		.INIT('h8)
	) name472 (
		_w4514_,
		_w4515_,
		_w4519_
	);
	LUT2 #(
		.INIT('h8)
	) name473 (
		_w4513_,
		_w4519_,
		_w4520_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		_w4518_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4521_,
		_w4522_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4244_,
		_w4523_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001 ,
		_w4202_,
		_w4524_
	);
	LUT2 #(
		.INIT('h8)
	) name478 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001 ,
		_w4211_,
		_w4525_
	);
	LUT2 #(
		.INIT('h8)
	) name479 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001 ,
		_w4194_,
		_w4526_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001 ,
		_w4224_,
		_w4527_
	);
	LUT2 #(
		.INIT('h8)
	) name481 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001 ,
		_w4205_,
		_w4528_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001 ,
		_w4226_,
		_w4529_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001 ,
		_w4220_,
		_w4530_
	);
	LUT2 #(
		.INIT('h8)
	) name484 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001 ,
		_w4228_,
		_w4531_
	);
	LUT2 #(
		.INIT('h8)
	) name485 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001 ,
		_w4197_,
		_w4532_
	);
	LUT2 #(
		.INIT('h8)
	) name486 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001 ,
		_w4215_,
		_w4533_
	);
	LUT2 #(
		.INIT('h8)
	) name487 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001 ,
		_w4218_,
		_w4534_
	);
	LUT2 #(
		.INIT('h8)
	) name488 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001 ,
		_w4209_,
		_w4535_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001 ,
		_w4190_,
		_w4536_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001 ,
		_w4222_,
		_w4537_
	);
	LUT2 #(
		.INIT('h8)
	) name491 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001 ,
		_w4213_,
		_w4538_
	);
	LUT2 #(
		.INIT('h8)
	) name492 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001 ,
		_w4200_,
		_w4539_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w4524_,
		_w4525_,
		_w4540_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w4526_,
		_w4527_,
		_w4541_
	);
	LUT2 #(
		.INIT('h1)
	) name495 (
		_w4528_,
		_w4529_,
		_w4542_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w4531_,
		_w4532_,
		_w4543_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w4536_,
		_w4537_,
		_w4544_
	);
	LUT2 #(
		.INIT('h1)
	) name498 (
		_w4538_,
		_w4539_,
		_w4545_
	);
	LUT2 #(
		.INIT('h8)
	) name499 (
		_w4544_,
		_w4545_,
		_w4546_
	);
	LUT2 #(
		.INIT('h8)
	) name500 (
		_w4542_,
		_w4543_,
		_w4547_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		_w4540_,
		_w4541_,
		_w4548_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		_w4530_,
		_w4533_,
		_w4549_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w4534_,
		_w4535_,
		_w4550_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		_w4549_,
		_w4550_,
		_w4551_
	);
	LUT2 #(
		.INIT('h8)
	) name505 (
		_w4547_,
		_w4548_,
		_w4552_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		_w4546_,
		_w4552_,
		_w4553_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		_w4551_,
		_w4553_,
		_w4554_
	);
	LUT2 #(
		.INIT('h8)
	) name508 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4554_,
		_w4555_
	);
	LUT2 #(
		.INIT('h8)
	) name509 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4521_,
		_w4556_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4457_,
		_w4557_
	);
	LUT2 #(
		.INIT('h8)
	) name511 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001 ,
		_w4228_,
		_w4558_
	);
	LUT2 #(
		.INIT('h8)
	) name512 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001 ,
		_w4213_,
		_w4559_
	);
	LUT2 #(
		.INIT('h8)
	) name513 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001 ,
		_w4200_,
		_w4560_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001 ,
		_w4194_,
		_w4561_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001 ,
		_w4222_,
		_w4562_
	);
	LUT2 #(
		.INIT('h8)
	) name516 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001 ,
		_w4197_,
		_w4563_
	);
	LUT2 #(
		.INIT('h8)
	) name517 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001 ,
		_w4220_,
		_w4564_
	);
	LUT2 #(
		.INIT('h8)
	) name518 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001 ,
		_w4190_,
		_w4565_
	);
	LUT2 #(
		.INIT('h8)
	) name519 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001 ,
		_w4226_,
		_w4566_
	);
	LUT2 #(
		.INIT('h8)
	) name520 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001 ,
		_w4209_,
		_w4567_
	);
	LUT2 #(
		.INIT('h8)
	) name521 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001 ,
		_w4215_,
		_w4568_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001 ,
		_w4218_,
		_w4569_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001 ,
		_w4224_,
		_w4570_
	);
	LUT2 #(
		.INIT('h8)
	) name524 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001 ,
		_w4202_,
		_w4571_
	);
	LUT2 #(
		.INIT('h8)
	) name525 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001 ,
		_w4205_,
		_w4572_
	);
	LUT2 #(
		.INIT('h8)
	) name526 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001 ,
		_w4211_,
		_w4573_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		_w4558_,
		_w4559_,
		_w4574_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		_w4560_,
		_w4561_,
		_w4575_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		_w4562_,
		_w4563_,
		_w4576_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		_w4565_,
		_w4566_,
		_w4577_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w4570_,
		_w4571_,
		_w4578_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w4572_,
		_w4573_,
		_w4579_
	);
	LUT2 #(
		.INIT('h8)
	) name533 (
		_w4578_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		_w4576_,
		_w4577_,
		_w4581_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		_w4574_,
		_w4575_,
		_w4582_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w4564_,
		_w4567_,
		_w4583_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		_w4568_,
		_w4569_,
		_w4584_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		_w4583_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		_w4581_,
		_w4582_,
		_w4586_
	);
	LUT2 #(
		.INIT('h8)
	) name540 (
		_w4580_,
		_w4586_,
		_w4587_
	);
	LUT2 #(
		.INIT('h8)
	) name541 (
		_w4585_,
		_w4587_,
		_w4588_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4588_,
		_w4589_
	);
	LUT2 #(
		.INIT('h1)
	) name543 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4328_,
		_w4590_
	);
	LUT2 #(
		.INIT('h8)
	) name544 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4588_,
		_w4591_
	);
	LUT2 #(
		.INIT('h8)
	) name545 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001 ,
		_w4222_,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001 ,
		_w4190_,
		_w4593_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001 ,
		_w4228_,
		_w4594_
	);
	LUT2 #(
		.INIT('h8)
	) name548 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001 ,
		_w4197_,
		_w4595_
	);
	LUT2 #(
		.INIT('h8)
	) name549 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001 ,
		_w4200_,
		_w4596_
	);
	LUT2 #(
		.INIT('h8)
	) name550 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001 ,
		_w4194_,
		_w4597_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001 ,
		_w4220_,
		_w4598_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001 ,
		_w4211_,
		_w4599_
	);
	LUT2 #(
		.INIT('h8)
	) name553 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001 ,
		_w4224_,
		_w4600_
	);
	LUT2 #(
		.INIT('h8)
	) name554 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001 ,
		_w4215_,
		_w4601_
	);
	LUT2 #(
		.INIT('h8)
	) name555 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001 ,
		_w4218_,
		_w4602_
	);
	LUT2 #(
		.INIT('h8)
	) name556 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001 ,
		_w4209_,
		_w4603_
	);
	LUT2 #(
		.INIT('h8)
	) name557 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001 ,
		_w4213_,
		_w4604_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001 ,
		_w4202_,
		_w4605_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001 ,
		_w4205_,
		_w4606_
	);
	LUT2 #(
		.INIT('h8)
	) name560 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001 ,
		_w4226_,
		_w4607_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		_w4592_,
		_w4593_,
		_w4608_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w4594_,
		_w4595_,
		_w4609_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		_w4596_,
		_w4597_,
		_w4610_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w4599_,
		_w4600_,
		_w4611_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w4604_,
		_w4605_,
		_w4612_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		_w4606_,
		_w4607_,
		_w4613_
	);
	LUT2 #(
		.INIT('h8)
	) name567 (
		_w4612_,
		_w4613_,
		_w4614_
	);
	LUT2 #(
		.INIT('h8)
	) name568 (
		_w4610_,
		_w4611_,
		_w4615_
	);
	LUT2 #(
		.INIT('h8)
	) name569 (
		_w4608_,
		_w4609_,
		_w4616_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		_w4598_,
		_w4601_,
		_w4617_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w4602_,
		_w4603_,
		_w4618_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		_w4617_,
		_w4618_,
		_w4619_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w4615_,
		_w4616_,
		_w4620_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		_w4614_,
		_w4620_,
		_w4621_
	);
	LUT2 #(
		.INIT('h8)
	) name575 (
		_w4619_,
		_w4621_,
		_w4622_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4622_,
		_w4623_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4622_,
		_w4624_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		_w4623_,
		_w4624_,
		_w4625_
	);
	LUT2 #(
		.INIT('h8)
	) name579 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001 ,
		_w4228_,
		_w4626_
	);
	LUT2 #(
		.INIT('h8)
	) name580 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001 ,
		_w4205_,
		_w4627_
	);
	LUT2 #(
		.INIT('h8)
	) name581 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001 ,
		_w4211_,
		_w4628_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001 ,
		_w4194_,
		_w4629_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001 ,
		_w4200_,
		_w4630_
	);
	LUT2 #(
		.INIT('h8)
	) name584 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001 ,
		_w4197_,
		_w4631_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001 ,
		_w4220_,
		_w4632_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001 ,
		_w4213_,
		_w4633_
	);
	LUT2 #(
		.INIT('h8)
	) name587 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001 ,
		_w4226_,
		_w4634_
	);
	LUT2 #(
		.INIT('h8)
	) name588 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001 ,
		_w4209_,
		_w4635_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001 ,
		_w4215_,
		_w4636_
	);
	LUT2 #(
		.INIT('h8)
	) name590 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001 ,
		_w4218_,
		_w4637_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001 ,
		_w4224_,
		_w4638_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001 ,
		_w4202_,
		_w4639_
	);
	LUT2 #(
		.INIT('h8)
	) name593 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001 ,
		_w4190_,
		_w4640_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001 ,
		_w4222_,
		_w4641_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		_w4626_,
		_w4627_,
		_w4642_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w4628_,
		_w4629_,
		_w4643_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w4630_,
		_w4631_,
		_w4644_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		_w4633_,
		_w4634_,
		_w4645_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		_w4638_,
		_w4639_,
		_w4646_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w4640_,
		_w4641_,
		_w4647_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		_w4646_,
		_w4647_,
		_w4648_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		_w4644_,
		_w4645_,
		_w4649_
	);
	LUT2 #(
		.INIT('h8)
	) name603 (
		_w4642_,
		_w4643_,
		_w4650_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w4632_,
		_w4635_,
		_w4651_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w4636_,
		_w4637_,
		_w4652_
	);
	LUT2 #(
		.INIT('h8)
	) name606 (
		_w4651_,
		_w4652_,
		_w4653_
	);
	LUT2 #(
		.INIT('h8)
	) name607 (
		_w4649_,
		_w4650_,
		_w4654_
	);
	LUT2 #(
		.INIT('h8)
	) name608 (
		_w4648_,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		_w4653_,
		_w4655_,
		_w4656_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4656_,
		_w4657_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4554_,
		_w4658_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4489_,
		_w4659_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4276_,
		_w4660_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4656_,
		_w4661_
	);
	LUT2 #(
		.INIT('h8)
	) name615 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4425_,
		_w4662_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4360_,
		_w4663_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001 ,
		_w4228_,
		_w4664_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001 ,
		_w4213_,
		_w4665_
	);
	LUT2 #(
		.INIT('h8)
	) name619 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001 ,
		_w4200_,
		_w4666_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001 ,
		_w4194_,
		_w4667_
	);
	LUT2 #(
		.INIT('h8)
	) name621 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001 ,
		_w4222_,
		_w4668_
	);
	LUT2 #(
		.INIT('h8)
	) name622 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001 ,
		_w4197_,
		_w4669_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001 ,
		_w4220_,
		_w4670_
	);
	LUT2 #(
		.INIT('h8)
	) name624 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001 ,
		_w4190_,
		_w4671_
	);
	LUT2 #(
		.INIT('h8)
	) name625 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001 ,
		_w4226_,
		_w4672_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001 ,
		_w4209_,
		_w4673_
	);
	LUT2 #(
		.INIT('h8)
	) name627 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001 ,
		_w4215_,
		_w4674_
	);
	LUT2 #(
		.INIT('h8)
	) name628 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001 ,
		_w4218_,
		_w4675_
	);
	LUT2 #(
		.INIT('h8)
	) name629 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001 ,
		_w4224_,
		_w4676_
	);
	LUT2 #(
		.INIT('h8)
	) name630 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001 ,
		_w4202_,
		_w4677_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001 ,
		_w4205_,
		_w4678_
	);
	LUT2 #(
		.INIT('h8)
	) name632 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001 ,
		_w4211_,
		_w4679_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		_w4664_,
		_w4665_,
		_w4680_
	);
	LUT2 #(
		.INIT('h1)
	) name634 (
		_w4666_,
		_w4667_,
		_w4681_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w4668_,
		_w4669_,
		_w4682_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w4671_,
		_w4672_,
		_w4683_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		_w4676_,
		_w4677_,
		_w4684_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		_w4678_,
		_w4679_,
		_w4685_
	);
	LUT2 #(
		.INIT('h8)
	) name639 (
		_w4684_,
		_w4685_,
		_w4686_
	);
	LUT2 #(
		.INIT('h8)
	) name640 (
		_w4682_,
		_w4683_,
		_w4687_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		_w4680_,
		_w4681_,
		_w4688_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		_w4670_,
		_w4673_,
		_w4689_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w4674_,
		_w4675_,
		_w4690_
	);
	LUT2 #(
		.INIT('h8)
	) name644 (
		_w4689_,
		_w4690_,
		_w4691_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		_w4687_,
		_w4688_,
		_w4692_
	);
	LUT2 #(
		.INIT('h8)
	) name646 (
		_w4686_,
		_w4692_,
		_w4693_
	);
	LUT2 #(
		.INIT('h8)
	) name647 (
		_w4691_,
		_w4693_,
		_w4694_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w4694_,
		_w4695_
	);
	LUT2 #(
		.INIT('h8)
	) name649 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w4694_,
		_w4696_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		_w4245_,
		_w4277_,
		_w4697_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w4329_,
		_w4361_,
		_w4698_
	);
	LUT2 #(
		.INIT('h1)
	) name652 (
		_w4393_,
		_w4394_,
		_w4699_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w4426_,
		_w4458_,
		_w4700_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w4490_,
		_w4522_,
		_w4701_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		_w4523_,
		_w4555_,
		_w4702_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w4556_,
		_w4557_,
		_w4703_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w4589_,
		_w4590_,
		_w4704_
	);
	LUT2 #(
		.INIT('h1)
	) name658 (
		_w4591_,
		_w4657_,
		_w4705_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		_w4658_,
		_w4659_,
		_w4706_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		_w4660_,
		_w4661_,
		_w4707_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w4662_,
		_w4663_,
		_w4708_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w4695_,
		_w4696_,
		_w4709_
	);
	LUT2 #(
		.INIT('h8)
	) name663 (
		_w4708_,
		_w4709_,
		_w4710_
	);
	LUT2 #(
		.INIT('h8)
	) name664 (
		_w4706_,
		_w4707_,
		_w4711_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		_w4704_,
		_w4705_,
		_w4712_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		_w4702_,
		_w4703_,
		_w4713_
	);
	LUT2 #(
		.INIT('h8)
	) name667 (
		_w4700_,
		_w4701_,
		_w4714_
	);
	LUT2 #(
		.INIT('h8)
	) name668 (
		_w4698_,
		_w4699_,
		_w4715_
	);
	LUT2 #(
		.INIT('h4)
	) name669 (
		_w4625_,
		_w4697_,
		_w4716_
	);
	LUT2 #(
		.INIT('h8)
	) name670 (
		_w4715_,
		_w4716_,
		_w4717_
	);
	LUT2 #(
		.INIT('h8)
	) name671 (
		_w4713_,
		_w4714_,
		_w4718_
	);
	LUT2 #(
		.INIT('h8)
	) name672 (
		_w4711_,
		_w4712_,
		_w4719_
	);
	LUT2 #(
		.INIT('h8)
	) name673 (
		_w4710_,
		_w4719_,
		_w4720_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		_w4717_,
		_w4718_,
		_w4721_
	);
	LUT2 #(
		.INIT('h8)
	) name675 (
		_w4720_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h8)
	) name676 (
		_w4297_,
		_w4722_,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name677 (
		_w4130_,
		_w4723_,
		_w4724_
	);
	LUT2 #(
		.INIT('h2)
	) name678 (
		_w4184_,
		_w4724_,
		_w4725_
	);
	LUT2 #(
		.INIT('h8)
	) name679 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[0]/P0001 ,
		_w4726_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4588_,
		_w4727_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4728_,
		_w4729_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4622_,
		_w4730_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[11]/P0001 ,
		_w4731_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		_w4730_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h8)
	) name686 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4425_,
		_w4734_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[8]/P0001 ,
		_w4735_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w4734_,
		_w4735_,
		_w4736_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4736_,
		_w4738_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[9]/P0001 ,
		_w4739_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4554_,
		_w4740_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w4739_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4741_,
		_w4742_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[4]/P0001 ,
		_w4743_
	);
	LUT2 #(
		.INIT('h4)
	) name697 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4360_,
		_w4744_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		_w4743_,
		_w4744_,
		_w4745_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4745_,
		_w4746_
	);
	LUT2 #(
		.INIT('h8)
	) name700 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4745_,
		_w4747_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w4746_,
		_w4747_,
		_w4748_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[2]/P0001 ,
		_w4749_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4521_,
		_w4750_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w4749_,
		_w4750_,
		_w4751_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4751_,
		_w4753_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w4752_,
		_w4753_,
		_w4754_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[10]/P0001 ,
		_w4755_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4276_,
		_w4756_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		_w4755_,
		_w4756_,
		_w4757_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4757_,
		_w4758_
	);
	LUT2 #(
		.INIT('h1)
	) name712 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4244_,
		_w4759_
	);
	LUT2 #(
		.INIT('h8)
	) name713 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[5]/P0001 ,
		_w4760_
	);
	LUT2 #(
		.INIT('h1)
	) name714 (
		_w4759_,
		_w4760_,
		_w4761_
	);
	LUT2 #(
		.INIT('h8)
	) name715 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4761_,
		_w4762_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4741_,
		_w4763_
	);
	LUT2 #(
		.INIT('h8)
	) name717 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[6]/P0001 ,
		_w4764_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4392_,
		_w4765_
	);
	LUT2 #(
		.INIT('h1)
	) name719 (
		_w4764_,
		_w4765_,
		_w4766_
	);
	LUT2 #(
		.INIT('h8)
	) name720 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w4766_,
		_w4767_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4457_,
		_w4768_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[1]/P0001 ,
		_w4769_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w4768_,
		_w4769_,
		_w4770_
	);
	LUT2 #(
		.INIT('h2)
	) name724 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4770_,
		_w4771_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4770_,
		_w4772_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		_w4771_,
		_w4772_,
		_w4773_
	);
	LUT2 #(
		.INIT('h1)
	) name727 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4732_,
		_w4774_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w4766_,
		_w4775_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4328_,
		_w4776_
	);
	LUT2 #(
		.INIT('h8)
	) name730 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[3]/P0001 ,
		_w4777_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w4776_,
		_w4777_,
		_w4778_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4778_,
		_w4779_
	);
	LUT2 #(
		.INIT('h1)
	) name733 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4778_,
		_w4780_
	);
	LUT2 #(
		.INIT('h8)
	) name734 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4728_,
		_w4781_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4656_,
		_w4782_
	);
	LUT2 #(
		.INIT('h8)
	) name736 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[7]/P0001 ,
		_w4783_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		_w4782_,
		_w4783_,
		_w4784_
	);
	LUT2 #(
		.INIT('h8)
	) name738 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4784_,
		_w4785_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[13]/P0001 ,
		_w4786_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4489_,
		_w4787_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w4786_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4788_,
		_w4789_
	);
	LUT2 #(
		.INIT('h8)
	) name743 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_psq_Taddr_Eb_reg[12]/P0001 ,
		_w4790_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4694_,
		_w4791_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		_w4790_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h2)
	) name746 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w4792_,
		_w4793_
	);
	LUT2 #(
		.INIT('h4)
	) name747 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w4792_,
		_w4794_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		_w4793_,
		_w4794_,
		_w4795_
	);
	LUT2 #(
		.INIT('h1)
	) name749 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4788_,
		_w4796_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4757_,
		_w4797_
	);
	LUT2 #(
		.INIT('h1)
	) name751 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4784_,
		_w4798_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4761_,
		_w4799_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		_w4729_,
		_w4733_,
		_w4800_
	);
	LUT2 #(
		.INIT('h1)
	) name754 (
		_w4737_,
		_w4738_,
		_w4801_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w4742_,
		_w4758_,
		_w4802_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		_w4762_,
		_w4763_,
		_w4803_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w4767_,
		_w4774_,
		_w4804_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		_w4775_,
		_w4779_,
		_w4805_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w4780_,
		_w4781_,
		_w4806_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w4785_,
		_w4789_,
		_w4807_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w4796_,
		_w4797_,
		_w4808_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		_w4798_,
		_w4799_,
		_w4809_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		_w4808_,
		_w4809_,
		_w4810_
	);
	LUT2 #(
		.INIT('h8)
	) name764 (
		_w4806_,
		_w4807_,
		_w4811_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		_w4804_,
		_w4805_,
		_w4812_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		_w4802_,
		_w4803_,
		_w4813_
	);
	LUT2 #(
		.INIT('h8)
	) name767 (
		_w4800_,
		_w4801_,
		_w4814_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		_w4748_,
		_w4754_,
		_w4815_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		_w4773_,
		_w4795_,
		_w4816_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		_w4815_,
		_w4816_,
		_w4817_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		_w4813_,
		_w4814_,
		_w4818_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		_w4811_,
		_w4812_,
		_w4819_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		_w4810_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h8)
	) name774 (
		_w4817_,
		_w4818_,
		_w4821_
	);
	LUT2 #(
		.INIT('h8)
	) name775 (
		_w4297_,
		_w4821_,
		_w4822_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		_w4820_,
		_w4822_,
		_w4823_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		\core_c_dec_Nseq_Ed_reg/P0001 ,
		_w4823_,
		_w4824_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		_w4184_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		_w4130_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		\core_c_dec_Nrti_Ed_reg/P0001 ,
		\core_c_dec_RTI_Ed_reg/P0001 ,
		_w4827_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		_w4826_,
		_w4827_,
		_w4828_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w4725_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		_w4186_,
		_w4297_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w4185_,
		_w4830_,
		_w4831_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		_w4829_,
		_w4831_,
		_w4832_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w4187_,
		_w4833_
	);
	LUT2 #(
		.INIT('h4)
	) name787 (
		_w4832_,
		_w4833_,
		_w4834_
	);
	LUT2 #(
		.INIT('h2)
	) name788 (
		_w4129_,
		_w4834_,
		_w4835_
	);
	LUT2 #(
		.INIT('h4)
	) name789 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		_w4129_,
		_w4837_
	);
	LUT2 #(
		.INIT('h8)
	) name791 (
		\sice_IRR_reg[0]/P0001 ,
		_w4837_,
		_w4838_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		_w4129_,
		_w4185_,
		_w4839_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w4829_,
		_w4839_,
		_w4840_
	);
	LUT2 #(
		.INIT('h8)
	) name794 (
		_w4726_,
		_w4840_,
		_w4841_
	);
	LUT2 #(
		.INIT('h2)
	) name795 (
		_w4186_,
		_w4297_,
		_w4842_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4842_,
		_w4843_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w4844_
	);
	LUT2 #(
		.INIT('h1)
	) name798 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4845_
	);
	LUT2 #(
		.INIT('h8)
	) name799 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001 ,
		_w4845_,
		_w4846_
	);
	LUT2 #(
		.INIT('h2)
	) name800 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4847_
	);
	LUT2 #(
		.INIT('h8)
	) name801 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001 ,
		_w4847_,
		_w4848_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4849_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001 ,
		_w4849_,
		_w4850_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w4851_
	);
	LUT2 #(
		.INIT('h8)
	) name805 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001 ,
		_w4851_,
		_w4852_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		_w4846_,
		_w4848_,
		_w4853_
	);
	LUT2 #(
		.INIT('h1)
	) name807 (
		_w4850_,
		_w4852_,
		_w4854_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		_w4853_,
		_w4854_,
		_w4855_
	);
	LUT2 #(
		.INIT('h2)
	) name809 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4855_,
		_w4856_
	);
	LUT2 #(
		.INIT('h4)
	) name810 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4855_,
		_w4857_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		_w4856_,
		_w4857_,
		_w4858_
	);
	LUT2 #(
		.INIT('h8)
	) name812 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001 ,
		_w4845_,
		_w4859_
	);
	LUT2 #(
		.INIT('h8)
	) name813 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001 ,
		_w4847_,
		_w4860_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001 ,
		_w4849_,
		_w4861_
	);
	LUT2 #(
		.INIT('h8)
	) name815 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001 ,
		_w4851_,
		_w4862_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w4859_,
		_w4860_,
		_w4863_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		_w4861_,
		_w4862_,
		_w4864_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		_w4863_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4865_,
		_w4866_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4865_,
		_w4867_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w4866_,
		_w4867_,
		_w4868_
	);
	LUT2 #(
		.INIT('h8)
	) name822 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001 ,
		_w4845_,
		_w4869_
	);
	LUT2 #(
		.INIT('h8)
	) name823 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001 ,
		_w4847_,
		_w4870_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001 ,
		_w4849_,
		_w4871_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001 ,
		_w4851_,
		_w4872_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w4869_,
		_w4870_,
		_w4873_
	);
	LUT2 #(
		.INIT('h1)
	) name827 (
		_w4871_,
		_w4872_,
		_w4874_
	);
	LUT2 #(
		.INIT('h8)
	) name828 (
		_w4873_,
		_w4874_,
		_w4875_
	);
	LUT2 #(
		.INIT('h2)
	) name829 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h4)
	) name830 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4875_,
		_w4877_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		_w4876_,
		_w4877_,
		_w4878_
	);
	LUT2 #(
		.INIT('h8)
	) name832 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001 ,
		_w4845_,
		_w4879_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001 ,
		_w4847_,
		_w4880_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001 ,
		_w4849_,
		_w4881_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001 ,
		_w4851_,
		_w4882_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w4879_,
		_w4880_,
		_w4883_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w4881_,
		_w4882_,
		_w4884_
	);
	LUT2 #(
		.INIT('h8)
	) name838 (
		_w4883_,
		_w4884_,
		_w4885_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w4885_,
		_w4886_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w4885_,
		_w4887_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		_w4886_,
		_w4887_,
		_w4888_
	);
	LUT2 #(
		.INIT('h8)
	) name842 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001 ,
		_w4845_,
		_w4889_
	);
	LUT2 #(
		.INIT('h8)
	) name843 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001 ,
		_w4847_,
		_w4890_
	);
	LUT2 #(
		.INIT('h8)
	) name844 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001 ,
		_w4849_,
		_w4891_
	);
	LUT2 #(
		.INIT('h8)
	) name845 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001 ,
		_w4851_,
		_w4892_
	);
	LUT2 #(
		.INIT('h1)
	) name846 (
		_w4889_,
		_w4890_,
		_w4893_
	);
	LUT2 #(
		.INIT('h1)
	) name847 (
		_w4891_,
		_w4892_,
		_w4894_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		_w4893_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h2)
	) name849 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4895_,
		_w4896_
	);
	LUT2 #(
		.INIT('h4)
	) name850 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4895_,
		_w4897_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w4896_,
		_w4897_,
		_w4898_
	);
	LUT2 #(
		.INIT('h8)
	) name852 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001 ,
		_w4845_,
		_w4899_
	);
	LUT2 #(
		.INIT('h8)
	) name853 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001 ,
		_w4847_,
		_w4900_
	);
	LUT2 #(
		.INIT('h8)
	) name854 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001 ,
		_w4849_,
		_w4901_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001 ,
		_w4851_,
		_w4902_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w4899_,
		_w4900_,
		_w4903_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		_w4901_,
		_w4902_,
		_w4904_
	);
	LUT2 #(
		.INIT('h8)
	) name858 (
		_w4903_,
		_w4904_,
		_w4905_
	);
	LUT2 #(
		.INIT('h2)
	) name859 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4905_,
		_w4906_
	);
	LUT2 #(
		.INIT('h4)
	) name860 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4905_,
		_w4907_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		_w4906_,
		_w4907_,
		_w4908_
	);
	LUT2 #(
		.INIT('h8)
	) name862 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001 ,
		_w4851_,
		_w4909_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001 ,
		_w4849_,
		_w4910_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001 ,
		_w4847_,
		_w4911_
	);
	LUT2 #(
		.INIT('h8)
	) name865 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001 ,
		_w4845_,
		_w4912_
	);
	LUT2 #(
		.INIT('h1)
	) name866 (
		_w4909_,
		_w4910_,
		_w4913_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		_w4911_,
		_w4912_,
		_w4914_
	);
	LUT2 #(
		.INIT('h8)
	) name868 (
		_w4913_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('h2)
	) name869 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w4915_,
		_w4916_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w4915_,
		_w4917_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w4916_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h8)
	) name872 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001 ,
		_w4845_,
		_w4919_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001 ,
		_w4847_,
		_w4920_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001 ,
		_w4849_,
		_w4921_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001 ,
		_w4851_,
		_w4922_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w4919_,
		_w4920_,
		_w4923_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w4921_,
		_w4922_,
		_w4924_
	);
	LUT2 #(
		.INIT('h8)
	) name878 (
		_w4923_,
		_w4924_,
		_w4925_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4925_,
		_w4926_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4925_,
		_w4927_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w4926_,
		_w4927_,
		_w4928_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001 ,
		_w4851_,
		_w4929_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001 ,
		_w4849_,
		_w4930_
	);
	LUT2 #(
		.INIT('h8)
	) name884 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001 ,
		_w4847_,
		_w4931_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001 ,
		_w4845_,
		_w4932_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		_w4929_,
		_w4930_,
		_w4933_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w4931_,
		_w4932_,
		_w4934_
	);
	LUT2 #(
		.INIT('h8)
	) name888 (
		_w4933_,
		_w4934_,
		_w4935_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w4935_,
		_w4936_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w4935_,
		_w4937_
	);
	LUT2 #(
		.INIT('h1)
	) name891 (
		_w4936_,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001 ,
		_w4845_,
		_w4939_
	);
	LUT2 #(
		.INIT('h8)
	) name893 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001 ,
		_w4847_,
		_w4940_
	);
	LUT2 #(
		.INIT('h8)
	) name894 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001 ,
		_w4849_,
		_w4941_
	);
	LUT2 #(
		.INIT('h8)
	) name895 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001 ,
		_w4851_,
		_w4942_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w4939_,
		_w4940_,
		_w4943_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		_w4941_,
		_w4942_,
		_w4944_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		_w4943_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('h2)
	) name899 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w4945_,
		_w4946_
	);
	LUT2 #(
		.INIT('h4)
	) name900 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w4945_,
		_w4947_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w4946_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h8)
	) name902 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001 ,
		_w4845_,
		_w4949_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001 ,
		_w4847_,
		_w4950_
	);
	LUT2 #(
		.INIT('h8)
	) name904 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001 ,
		_w4849_,
		_w4951_
	);
	LUT2 #(
		.INIT('h8)
	) name905 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001 ,
		_w4851_,
		_w4952_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w4949_,
		_w4950_,
		_w4953_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w4951_,
		_w4952_,
		_w4954_
	);
	LUT2 #(
		.INIT('h8)
	) name908 (
		_w4953_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('h2)
	) name909 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4955_,
		_w4956_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4955_,
		_w4957_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w4956_,
		_w4957_,
		_w4958_
	);
	LUT2 #(
		.INIT('h8)
	) name912 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001 ,
		_w4845_,
		_w4959_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001 ,
		_w4847_,
		_w4960_
	);
	LUT2 #(
		.INIT('h8)
	) name914 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001 ,
		_w4849_,
		_w4961_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001 ,
		_w4851_,
		_w4962_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w4959_,
		_w4960_,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w4961_,
		_w4962_,
		_w4964_
	);
	LUT2 #(
		.INIT('h8)
	) name918 (
		_w4963_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h2)
	) name919 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w4965_,
		_w4966_
	);
	LUT2 #(
		.INIT('h4)
	) name920 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w4965_,
		_w4967_
	);
	LUT2 #(
		.INIT('h1)
	) name921 (
		_w4966_,
		_w4967_,
		_w4968_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001 ,
		_w4845_,
		_w4969_
	);
	LUT2 #(
		.INIT('h8)
	) name923 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001 ,
		_w4847_,
		_w4970_
	);
	LUT2 #(
		.INIT('h8)
	) name924 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001 ,
		_w4849_,
		_w4971_
	);
	LUT2 #(
		.INIT('h8)
	) name925 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001 ,
		_w4851_,
		_w4972_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		_w4969_,
		_w4970_,
		_w4973_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w4971_,
		_w4972_,
		_w4974_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		_w4973_,
		_w4974_,
		_w4975_
	);
	LUT2 #(
		.INIT('h2)
	) name929 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w4975_,
		_w4976_
	);
	LUT2 #(
		.INIT('h4)
	) name930 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w4975_,
		_w4977_
	);
	LUT2 #(
		.INIT('h1)
	) name931 (
		_w4976_,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h8)
	) name932 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001 ,
		_w4845_,
		_w4979_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001 ,
		_w4847_,
		_w4980_
	);
	LUT2 #(
		.INIT('h8)
	) name934 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001 ,
		_w4849_,
		_w4981_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001 ,
		_w4851_,
		_w4982_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w4979_,
		_w4980_,
		_w4983_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		_w4981_,
		_w4982_,
		_w4984_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		_w4983_,
		_w4984_,
		_w4985_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w4985_,
		_w4986_
	);
	LUT2 #(
		.INIT('h4)
	) name940 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w4985_,
		_w4987_
	);
	LUT2 #(
		.INIT('h1)
	) name941 (
		_w4986_,
		_w4987_,
		_w4988_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001 ,
		_w4851_,
		_w4989_
	);
	LUT2 #(
		.INIT('h8)
	) name943 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001 ,
		_w4849_,
		_w4990_
	);
	LUT2 #(
		.INIT('h8)
	) name944 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001 ,
		_w4845_,
		_w4991_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001 ,
		_w4847_,
		_w4992_
	);
	LUT2 #(
		.INIT('h1)
	) name946 (
		_w4989_,
		_w4990_,
		_w4993_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w4991_,
		_w4992_,
		_w4994_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		_w4993_,
		_w4994_,
		_w4995_
	);
	LUT2 #(
		.INIT('h2)
	) name949 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w4995_,
		_w4996_
	);
	LUT2 #(
		.INIT('h4)
	) name950 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w4995_,
		_w4997_
	);
	LUT2 #(
		.INIT('h1)
	) name951 (
		_w4996_,
		_w4997_,
		_w4998_
	);
	LUT2 #(
		.INIT('h8)
	) name952 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001 ,
		_w4845_,
		_w4999_
	);
	LUT2 #(
		.INIT('h8)
	) name953 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001 ,
		_w4847_,
		_w5000_
	);
	LUT2 #(
		.INIT('h8)
	) name954 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001 ,
		_w4849_,
		_w5001_
	);
	LUT2 #(
		.INIT('h8)
	) name955 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001 ,
		_w4851_,
		_w5002_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		_w4999_,
		_w5000_,
		_w5003_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		_w5001_,
		_w5002_,
		_w5004_
	);
	LUT2 #(
		.INIT('h8)
	) name958 (
		_w5003_,
		_w5004_,
		_w5005_
	);
	LUT2 #(
		.INIT('h2)
	) name959 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w5005_,
		_w5006_
	);
	LUT2 #(
		.INIT('h4)
	) name960 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w5005_,
		_w5007_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		_w5006_,
		_w5007_,
		_w5008_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001 ,
		_w4851_,
		_w5009_
	);
	LUT2 #(
		.INIT('h8)
	) name963 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001 ,
		_w4849_,
		_w5010_
	);
	LUT2 #(
		.INIT('h8)
	) name964 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001 ,
		_w4847_,
		_w5011_
	);
	LUT2 #(
		.INIT('h8)
	) name965 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001 ,
		_w4845_,
		_w5012_
	);
	LUT2 #(
		.INIT('h1)
	) name966 (
		_w5009_,
		_w5010_,
		_w5013_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		_w5011_,
		_w5012_,
		_w5014_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		_w5013_,
		_w5014_,
		_w5015_
	);
	LUT2 #(
		.INIT('h2)
	) name969 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name970 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w5015_,
		_w5017_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		_w5016_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001 ,
		_w4845_,
		_w5019_
	);
	LUT2 #(
		.INIT('h8)
	) name973 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001 ,
		_w4847_,
		_w5020_
	);
	LUT2 #(
		.INIT('h8)
	) name974 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001 ,
		_w4849_,
		_w5021_
	);
	LUT2 #(
		.INIT('h8)
	) name975 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001 ,
		_w4851_,
		_w5022_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w5019_,
		_w5020_,
		_w5023_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		_w5021_,
		_w5022_,
		_w5024_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h2)
	) name979 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h4)
	) name980 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w5025_,
		_w5027_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w5026_,
		_w5027_,
		_w5028_
	);
	LUT2 #(
		.INIT('h1)
	) name982 (
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w4858_,
		_w5029_
	);
	LUT2 #(
		.INIT('h1)
	) name983 (
		_w4868_,
		_w4878_,
		_w5030_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w4888_,
		_w4898_,
		_w5031_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w4908_,
		_w4918_,
		_w5032_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		_w4928_,
		_w4938_,
		_w5033_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w4948_,
		_w4958_,
		_w5034_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w4968_,
		_w4978_,
		_w5035_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w4988_,
		_w4998_,
		_w5036_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		_w5008_,
		_w5018_,
		_w5037_
	);
	LUT2 #(
		.INIT('h4)
	) name991 (
		_w5028_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		_w5035_,
		_w5036_,
		_w5039_
	);
	LUT2 #(
		.INIT('h8)
	) name993 (
		_w5033_,
		_w5034_,
		_w5040_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		_w5031_,
		_w5032_,
		_w5041_
	);
	LUT2 #(
		.INIT('h8)
	) name995 (
		_w5029_,
		_w5030_,
		_w5042_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		_w5041_,
		_w5042_,
		_w5043_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		_w5039_,
		_w5040_,
		_w5044_
	);
	LUT2 #(
		.INIT('h8)
	) name998 (
		_w5038_,
		_w5044_,
		_w5045_
	);
	LUT2 #(
		.INIT('h8)
	) name999 (
		_w5043_,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		_w4129_,
		_w4844_,
		_w5047_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w5046_,
		_w5047_,
		_w5048_
	);
	LUT2 #(
		.INIT('h4)
	) name1002 (
		_w4843_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h4)
	) name1003 (
		_w4829_,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w5050_,
		_w5051_
	);
	LUT2 #(
		.INIT('h4)
	) name1005 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4840_,
		_w5052_
	);
	LUT2 #(
		.INIT('h1)
	) name1006 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4829_,
		_w5053_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		_w4830_,
		_w5053_,
		_w5054_
	);
	LUT2 #(
		.INIT('h8)
	) name1008 (
		_w4844_,
		_w5046_,
		_w5055_
	);
	LUT2 #(
		.INIT('h2)
	) name1009 (
		_w5053_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h2)
	) name1010 (
		_w4129_,
		_w5054_,
		_w5057_
	);
	LUT2 #(
		.INIT('h4)
	) name1011 (
		_w5056_,
		_w5057_,
		_w5058_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w5052_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h1)
	) name1013 (
		_w4588_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		_w4838_,
		_w4841_,
		_w5061_
	);
	LUT2 #(
		.INIT('h4)
	) name1015 (
		_w5051_,
		_w5061_,
		_w5062_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		_w4836_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h4)
	) name1017 (
		_w5060_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h2)
	) name1018 (
		_w4128_,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		_w4048_,
		_w4056_,
		_w5066_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w5066_,
		_w5067_
	);
	LUT2 #(
		.INIT('h8)
	) name1021 (
		\idma_DSreq_reg/NET0131 ,
		_w4055_,
		_w5068_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w5068_,
		_w5069_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		_w5067_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h2)
	) name1024 (
		_w4099_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h1)
	) name1025 (
		_w4127_,
		_w5071_,
		_w5072_
	);
	LUT2 #(
		.INIT('h4)
	) name1026 (
		_w5065_,
		_w5072_,
		_w5073_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w4104_,
		_w5074_
	);
	LUT2 #(
		.INIT('h1)
	) name1028 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w4117_,
		_w5075_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w4117_,
		_w5076_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		_w5075_,
		_w5076_,
		_w5077_
	);
	LUT2 #(
		.INIT('h1)
	) name1031 (
		_w4104_,
		_w5077_,
		_w5078_
	);
	LUT2 #(
		.INIT('h1)
	) name1032 (
		_w5074_,
		_w5078_,
		_w5079_
	);
	LUT2 #(
		.INIT('h8)
	) name1033 (
		_w4120_,
		_w5079_,
		_w5080_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w4276_,
		_w5059_,
		_w5081_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		_w5082_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		\core_c_psq_EXA_reg[2]/P0001 ,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		\core_c_psq_EXA_reg[3]/P0001 ,
		_w5083_,
		_w5084_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h8)
	) name1039 (
		\core_c_psq_EXA_reg[5]/P0001 ,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('h8)
	) name1040 (
		\core_c_psq_EXA_reg[6]/P0001 ,
		_w5086_,
		_w5087_
	);
	LUT2 #(
		.INIT('h8)
	) name1041 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		_w5087_,
		_w5088_
	);
	LUT2 #(
		.INIT('h8)
	) name1042 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h8)
	) name1043 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h1)
	) name1044 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		_w5090_,
		_w5091_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		_w5090_,
		_w5092_
	);
	LUT2 #(
		.INIT('h1)
	) name1046 (
		_w5091_,
		_w5092_,
		_w5093_
	);
	LUT2 #(
		.INIT('h8)
	) name1047 (
		_w4835_,
		_w5093_,
		_w5094_
	);
	LUT2 #(
		.INIT('h8)
	) name1048 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w5095_
	);
	LUT2 #(
		.INIT('h8)
	) name1049 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w5095_,
		_w5096_
	);
	LUT2 #(
		.INIT('h8)
	) name1050 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h8)
	) name1051 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w5097_,
		_w5098_
	);
	LUT2 #(
		.INIT('h8)
	) name1052 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h8)
	) name1053 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w5099_,
		_w5100_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w5100_,
		_w5101_
	);
	LUT2 #(
		.INIT('h8)
	) name1055 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w5101_,
		_w5102_
	);
	LUT2 #(
		.INIT('h8)
	) name1056 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w5102_,
		_w5103_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w5103_,
		_w5104_
	);
	LUT2 #(
		.INIT('h8)
	) name1058 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w5103_,
		_w5105_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		_w5104_,
		_w5105_,
		_w5106_
	);
	LUT2 #(
		.INIT('h8)
	) name1060 (
		_w5050_,
		_w5106_,
		_w5107_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		_w4755_,
		_w4840_,
		_w5108_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		\sice_IRR_reg[10]/P0001 ,
		_w4837_,
		_w5109_
	);
	LUT2 #(
		.INIT('h1)
	) name1063 (
		_w5107_,
		_w5109_,
		_w5110_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w5108_,
		_w5110_,
		_w5111_
	);
	LUT2 #(
		.INIT('h4)
	) name1065 (
		_w5094_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h4)
	) name1066 (
		_w5081_,
		_w5112_,
		_w5113_
	);
	LUT2 #(
		.INIT('h2)
	) name1067 (
		_w4128_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w5066_,
		_w5115_
	);
	LUT2 #(
		.INIT('h8)
	) name1069 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w5068_,
		_w5116_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		_w5115_,
		_w5116_,
		_w5117_
	);
	LUT2 #(
		.INIT('h2)
	) name1071 (
		_w4099_,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w5080_,
		_w5118_,
		_w5119_
	);
	LUT2 #(
		.INIT('h4)
	) name1073 (
		_w5114_,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w4104_,
		_w5121_
	);
	LUT2 #(
		.INIT('h8)
	) name1075 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w4117_,
		_w5122_
	);
	LUT2 #(
		.INIT('h2)
	) name1076 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w4117_,
		_w5123_
	);
	LUT2 #(
		.INIT('h1)
	) name1077 (
		_w4104_,
		_w5122_,
		_w5124_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		_w5123_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w5121_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h8)
	) name1080 (
		_w4120_,
		_w5126_,
		_w5127_
	);
	LUT2 #(
		.INIT('h1)
	) name1081 (
		_w4622_,
		_w5059_,
		_w5128_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		_w5092_,
		_w5129_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		_w5092_,
		_w5130_
	);
	LUT2 #(
		.INIT('h1)
	) name1084 (
		_w5129_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h8)
	) name1085 (
		_w4835_,
		_w5131_,
		_w5132_
	);
	LUT2 #(
		.INIT('h1)
	) name1086 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w5105_,
		_w5133_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w5105_,
		_w5134_
	);
	LUT2 #(
		.INIT('h1)
	) name1088 (
		_w5133_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h8)
	) name1089 (
		_w5050_,
		_w5135_,
		_w5136_
	);
	LUT2 #(
		.INIT('h8)
	) name1090 (
		_w4731_,
		_w4840_,
		_w5137_
	);
	LUT2 #(
		.INIT('h8)
	) name1091 (
		\sice_IRR_reg[11]/P0001 ,
		_w4837_,
		_w5138_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w5136_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h4)
	) name1093 (
		_w5137_,
		_w5139_,
		_w5140_
	);
	LUT2 #(
		.INIT('h4)
	) name1094 (
		_w5132_,
		_w5140_,
		_w5141_
	);
	LUT2 #(
		.INIT('h4)
	) name1095 (
		_w5128_,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h2)
	) name1096 (
		_w4128_,
		_w5142_,
		_w5143_
	);
	LUT2 #(
		.INIT('h8)
	) name1097 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w5066_,
		_w5144_
	);
	LUT2 #(
		.INIT('h8)
	) name1098 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w5068_,
		_w5145_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		_w5144_,
		_w5145_,
		_w5146_
	);
	LUT2 #(
		.INIT('h2)
	) name1100 (
		_w4099_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('h1)
	) name1101 (
		_w5127_,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h4)
	) name1102 (
		_w5143_,
		_w5148_,
		_w5149_
	);
	LUT2 #(
		.INIT('h4)
	) name1103 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w4104_,
		_w5150_
	);
	LUT2 #(
		.INIT('h1)
	) name1104 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w4117_,
		_w5151_
	);
	LUT2 #(
		.INIT('h4)
	) name1105 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w4117_,
		_w5152_
	);
	LUT2 #(
		.INIT('h1)
	) name1106 (
		_w5151_,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h1)
	) name1107 (
		_w4104_,
		_w5153_,
		_w5154_
	);
	LUT2 #(
		.INIT('h1)
	) name1108 (
		_w5150_,
		_w5154_,
		_w5155_
	);
	LUT2 #(
		.INIT('h8)
	) name1109 (
		_w4120_,
		_w5155_,
		_w5156_
	);
	LUT2 #(
		.INIT('h1)
	) name1110 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_EXA_reg[1]/P0001 ,
		_w5157_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w5082_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h8)
	) name1112 (
		_w4835_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h8)
	) name1113 (
		\sice_IRR_reg[1]/P0001 ,
		_w4837_,
		_w5160_
	);
	LUT2 #(
		.INIT('h8)
	) name1114 (
		_w4769_,
		_w4840_,
		_w5161_
	);
	LUT2 #(
		.INIT('h1)
	) name1115 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w5162_
	);
	LUT2 #(
		.INIT('h1)
	) name1116 (
		_w5095_,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h8)
	) name1117 (
		_w5050_,
		_w5163_,
		_w5164_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w4457_,
		_w5059_,
		_w5165_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		_w5160_,
		_w5161_,
		_w5166_
	);
	LUT2 #(
		.INIT('h4)
	) name1120 (
		_w5164_,
		_w5166_,
		_w5167_
	);
	LUT2 #(
		.INIT('h4)
	) name1121 (
		_w5159_,
		_w5167_,
		_w5168_
	);
	LUT2 #(
		.INIT('h4)
	) name1122 (
		_w5165_,
		_w5168_,
		_w5169_
	);
	LUT2 #(
		.INIT('h2)
	) name1123 (
		_w4128_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h8)
	) name1124 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w5066_,
		_w5171_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w5068_,
		_w5172_
	);
	LUT2 #(
		.INIT('h1)
	) name1126 (
		_w5171_,
		_w5172_,
		_w5173_
	);
	LUT2 #(
		.INIT('h2)
	) name1127 (
		_w4099_,
		_w5173_,
		_w5174_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w5156_,
		_w5174_,
		_w5175_
	);
	LUT2 #(
		.INIT('h4)
	) name1129 (
		_w5170_,
		_w5175_,
		_w5176_
	);
	LUT2 #(
		.INIT('h4)
	) name1130 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w4104_,
		_w5177_
	);
	LUT2 #(
		.INIT('h1)
	) name1131 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w4117_,
		_w5178_
	);
	LUT2 #(
		.INIT('h4)
	) name1132 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w4117_,
		_w5179_
	);
	LUT2 #(
		.INIT('h1)
	) name1133 (
		_w5178_,
		_w5179_,
		_w5180_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		_w4104_,
		_w5180_,
		_w5181_
	);
	LUT2 #(
		.INIT('h1)
	) name1135 (
		_w5177_,
		_w5181_,
		_w5182_
	);
	LUT2 #(
		.INIT('h8)
	) name1136 (
		_w4120_,
		_w5182_,
		_w5183_
	);
	LUT2 #(
		.INIT('h4)
	) name1137 (
		_w4521_,
		_w5058_,
		_w5184_
	);
	LUT2 #(
		.INIT('h8)
	) name1138 (
		\sice_IRR_reg[2]/P0001 ,
		_w4837_,
		_w5185_
	);
	LUT2 #(
		.INIT('h1)
	) name1139 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w5095_,
		_w5186_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w5096_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h8)
	) name1141 (
		_w5050_,
		_w5187_,
		_w5188_
	);
	LUT2 #(
		.INIT('h2)
	) name1142 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4184_,
		_w5189_
	);
	LUT2 #(
		.INIT('h4)
	) name1143 (
		\core_c_psq_Taddr_Eb_reg[2]/P0001 ,
		_w5189_,
		_w5190_
	);
	LUT2 #(
		.INIT('h2)
	) name1144 (
		_w4521_,
		_w5189_,
		_w5191_
	);
	LUT2 #(
		.INIT('h1)
	) name1145 (
		_w5190_,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h8)
	) name1146 (
		_w4840_,
		_w5192_,
		_w5193_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		\core_c_psq_EXA_reg[2]/P0001 ,
		_w5082_,
		_w5194_
	);
	LUT2 #(
		.INIT('h1)
	) name1148 (
		_w5083_,
		_w5194_,
		_w5195_
	);
	LUT2 #(
		.INIT('h8)
	) name1149 (
		_w4835_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4105_,
		_w5197_
	);
	LUT2 #(
		.INIT('h1)
	) name1151 (
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		_w5198_
	);
	LUT2 #(
		.INIT('h1)
	) name1152 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		_w5199_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		\core_c_psq_Iact_E_reg[8]/NET0131 ,
		_w5200_
	);
	LUT2 #(
		.INIT('h8)
	) name1154 (
		_w5199_,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h8)
	) name1155 (
		_w5198_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		_w5197_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h1)
	) name1157 (
		_w5185_,
		_w5203_,
		_w5204_
	);
	LUT2 #(
		.INIT('h4)
	) name1158 (
		_w5188_,
		_w5204_,
		_w5205_
	);
	LUT2 #(
		.INIT('h4)
	) name1159 (
		_w5193_,
		_w5205_,
		_w5206_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		_w5196_,
		_w5206_,
		_w5207_
	);
	LUT2 #(
		.INIT('h4)
	) name1161 (
		_w5184_,
		_w5207_,
		_w5208_
	);
	LUT2 #(
		.INIT('h2)
	) name1162 (
		_w4128_,
		_w5208_,
		_w5209_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w5066_,
		_w5210_
	);
	LUT2 #(
		.INIT('h8)
	) name1164 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w5068_,
		_w5211_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		_w5210_,
		_w5211_,
		_w5212_
	);
	LUT2 #(
		.INIT('h2)
	) name1166 (
		_w4099_,
		_w5212_,
		_w5213_
	);
	LUT2 #(
		.INIT('h1)
	) name1167 (
		_w5183_,
		_w5213_,
		_w5214_
	);
	LUT2 #(
		.INIT('h4)
	) name1168 (
		_w5209_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h4)
	) name1169 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w4104_,
		_w5216_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w4117_,
		_w5217_
	);
	LUT2 #(
		.INIT('h4)
	) name1171 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w4117_,
		_w5218_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w5217_,
		_w5218_,
		_w5219_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		_w4104_,
		_w5219_,
		_w5220_
	);
	LUT2 #(
		.INIT('h1)
	) name1174 (
		_w5216_,
		_w5220_,
		_w5221_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		_w4120_,
		_w5221_,
		_w5222_
	);
	LUT2 #(
		.INIT('h4)
	) name1176 (
		_w4328_,
		_w5058_,
		_w5223_
	);
	LUT2 #(
		.INIT('h8)
	) name1177 (
		\sice_IRR_reg[3]/P0001 ,
		_w4837_,
		_w5224_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w5096_,
		_w5225_
	);
	LUT2 #(
		.INIT('h1)
	) name1179 (
		_w5097_,
		_w5225_,
		_w5226_
	);
	LUT2 #(
		.INIT('h8)
	) name1180 (
		_w5050_,
		_w5226_,
		_w5227_
	);
	LUT2 #(
		.INIT('h4)
	) name1181 (
		\core_c_psq_Taddr_Eb_reg[3]/P0001 ,
		_w5189_,
		_w5228_
	);
	LUT2 #(
		.INIT('h2)
	) name1182 (
		_w4328_,
		_w5189_,
		_w5229_
	);
	LUT2 #(
		.INIT('h1)
	) name1183 (
		_w5228_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h8)
	) name1184 (
		_w4840_,
		_w5230_,
		_w5231_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		\core_c_psq_EXA_reg[3]/P0001 ,
		_w5083_,
		_w5232_
	);
	LUT2 #(
		.INIT('h1)
	) name1186 (
		_w5084_,
		_w5232_,
		_w5233_
	);
	LUT2 #(
		.INIT('h8)
	) name1187 (
		_w4835_,
		_w5233_,
		_w5234_
	);
	LUT2 #(
		.INIT('h1)
	) name1188 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		_w5235_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		\core_c_psq_Iact_E_reg[9]/NET0131 ,
		_w5237_
	);
	LUT2 #(
		.INIT('h8)
	) name1191 (
		_w5236_,
		_w5237_,
		_w5238_
	);
	LUT2 #(
		.INIT('h8)
	) name1192 (
		_w5235_,
		_w5238_,
		_w5239_
	);
	LUT2 #(
		.INIT('h2)
	) name1193 (
		_w5197_,
		_w5239_,
		_w5240_
	);
	LUT2 #(
		.INIT('h1)
	) name1194 (
		_w5224_,
		_w5240_,
		_w5241_
	);
	LUT2 #(
		.INIT('h4)
	) name1195 (
		_w5227_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		_w5231_,
		_w5242_,
		_w5243_
	);
	LUT2 #(
		.INIT('h4)
	) name1197 (
		_w5234_,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h4)
	) name1198 (
		_w5223_,
		_w5244_,
		_w5245_
	);
	LUT2 #(
		.INIT('h2)
	) name1199 (
		_w4128_,
		_w5245_,
		_w5246_
	);
	LUT2 #(
		.INIT('h8)
	) name1200 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w5066_,
		_w5247_
	);
	LUT2 #(
		.INIT('h8)
	) name1201 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w5068_,
		_w5248_
	);
	LUT2 #(
		.INIT('h1)
	) name1202 (
		_w5247_,
		_w5248_,
		_w5249_
	);
	LUT2 #(
		.INIT('h2)
	) name1203 (
		_w4099_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		_w5222_,
		_w5250_,
		_w5251_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		_w5246_,
		_w5251_,
		_w5252_
	);
	LUT2 #(
		.INIT('h4)
	) name1206 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w4104_,
		_w5253_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w4117_,
		_w5254_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w4117_,
		_w5255_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w5254_,
		_w5255_,
		_w5256_
	);
	LUT2 #(
		.INIT('h1)
	) name1210 (
		_w4104_,
		_w5256_,
		_w5257_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w5253_,
		_w5257_,
		_w5258_
	);
	LUT2 #(
		.INIT('h8)
	) name1212 (
		_w4120_,
		_w5258_,
		_w5259_
	);
	LUT2 #(
		.INIT('h4)
	) name1213 (
		_w4360_,
		_w5058_,
		_w5260_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		\sice_IRR_reg[4]/P0001 ,
		_w4837_,
		_w5261_
	);
	LUT2 #(
		.INIT('h1)
	) name1215 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w5097_,
		_w5262_
	);
	LUT2 #(
		.INIT('h1)
	) name1216 (
		_w5098_,
		_w5262_,
		_w5263_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		_w5050_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h4)
	) name1218 (
		\core_c_psq_Taddr_Eb_reg[4]/P0001 ,
		_w5189_,
		_w5265_
	);
	LUT2 #(
		.INIT('h2)
	) name1219 (
		_w4360_,
		_w5189_,
		_w5266_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w5265_,
		_w5266_,
		_w5267_
	);
	LUT2 #(
		.INIT('h8)
	) name1221 (
		_w4840_,
		_w5267_,
		_w5268_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		_w5084_,
		_w5269_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w5085_,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h8)
	) name1224 (
		_w4835_,
		_w5270_,
		_w5271_
	);
	LUT2 #(
		.INIT('h1)
	) name1225 (
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[7]/NET0131 ,
		_w5272_
	);
	LUT2 #(
		.INIT('h8)
	) name1226 (
		_w5235_,
		_w5272_,
		_w5273_
	);
	LUT2 #(
		.INIT('h2)
	) name1227 (
		_w5197_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w5261_,
		_w5274_,
		_w5275_
	);
	LUT2 #(
		.INIT('h4)
	) name1229 (
		_w5264_,
		_w5275_,
		_w5276_
	);
	LUT2 #(
		.INIT('h4)
	) name1230 (
		_w5268_,
		_w5276_,
		_w5277_
	);
	LUT2 #(
		.INIT('h4)
	) name1231 (
		_w5271_,
		_w5277_,
		_w5278_
	);
	LUT2 #(
		.INIT('h4)
	) name1232 (
		_w5260_,
		_w5278_,
		_w5279_
	);
	LUT2 #(
		.INIT('h2)
	) name1233 (
		_w4128_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h8)
	) name1234 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w5066_,
		_w5281_
	);
	LUT2 #(
		.INIT('h8)
	) name1235 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w5068_,
		_w5282_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w5281_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h2)
	) name1237 (
		_w4099_,
		_w5283_,
		_w5284_
	);
	LUT2 #(
		.INIT('h1)
	) name1238 (
		_w5259_,
		_w5284_,
		_w5285_
	);
	LUT2 #(
		.INIT('h4)
	) name1239 (
		_w5280_,
		_w5285_,
		_w5286_
	);
	LUT2 #(
		.INIT('h4)
	) name1240 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w4104_,
		_w5287_
	);
	LUT2 #(
		.INIT('h1)
	) name1241 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w4117_,
		_w5288_
	);
	LUT2 #(
		.INIT('h4)
	) name1242 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w4117_,
		_w5289_
	);
	LUT2 #(
		.INIT('h1)
	) name1243 (
		_w5288_,
		_w5289_,
		_w5290_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w4104_,
		_w5290_,
		_w5291_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		_w5287_,
		_w5291_,
		_w5292_
	);
	LUT2 #(
		.INIT('h8)
	) name1246 (
		_w4120_,
		_w5292_,
		_w5293_
	);
	LUT2 #(
		.INIT('h1)
	) name1247 (
		_w4244_,
		_w5059_,
		_w5294_
	);
	LUT2 #(
		.INIT('h8)
	) name1248 (
		_w4760_,
		_w4840_,
		_w5295_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w5098_,
		_w5296_
	);
	LUT2 #(
		.INIT('h1)
	) name1250 (
		_w5099_,
		_w5296_,
		_w5297_
	);
	LUT2 #(
		.INIT('h8)
	) name1251 (
		_w5050_,
		_w5297_,
		_w5298_
	);
	LUT2 #(
		.INIT('h1)
	) name1252 (
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		_w5299_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		\core_c_psq_Iact_E_reg[3]/NET0131 ,
		_w5300_
	);
	LUT2 #(
		.INIT('h8)
	) name1254 (
		_w5299_,
		_w5300_,
		_w5301_
	);
	LUT2 #(
		.INIT('h2)
	) name1255 (
		_w5197_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h1)
	) name1256 (
		\core_c_psq_EXA_reg[5]/P0001 ,
		_w5085_,
		_w5303_
	);
	LUT2 #(
		.INIT('h1)
	) name1257 (
		_w5086_,
		_w5303_,
		_w5304_
	);
	LUT2 #(
		.INIT('h8)
	) name1258 (
		_w4835_,
		_w5304_,
		_w5305_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		\sice_IRR_reg[5]/P0001 ,
		_w4837_,
		_w5306_
	);
	LUT2 #(
		.INIT('h1)
	) name1260 (
		_w5302_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('h4)
	) name1261 (
		_w5295_,
		_w5307_,
		_w5308_
	);
	LUT2 #(
		.INIT('h4)
	) name1262 (
		_w5298_,
		_w5308_,
		_w5309_
	);
	LUT2 #(
		.INIT('h4)
	) name1263 (
		_w5305_,
		_w5309_,
		_w5310_
	);
	LUT2 #(
		.INIT('h4)
	) name1264 (
		_w5294_,
		_w5310_,
		_w5311_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		_w4128_,
		_w5311_,
		_w5312_
	);
	LUT2 #(
		.INIT('h8)
	) name1266 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w5066_,
		_w5313_
	);
	LUT2 #(
		.INIT('h8)
	) name1267 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w5068_,
		_w5314_
	);
	LUT2 #(
		.INIT('h1)
	) name1268 (
		_w5313_,
		_w5314_,
		_w5315_
	);
	LUT2 #(
		.INIT('h2)
	) name1269 (
		_w4099_,
		_w5315_,
		_w5316_
	);
	LUT2 #(
		.INIT('h1)
	) name1270 (
		_w5293_,
		_w5316_,
		_w5317_
	);
	LUT2 #(
		.INIT('h4)
	) name1271 (
		_w5312_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h4)
	) name1272 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w4104_,
		_w5319_
	);
	LUT2 #(
		.INIT('h1)
	) name1273 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w4117_,
		_w5320_
	);
	LUT2 #(
		.INIT('h4)
	) name1274 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w4117_,
		_w5321_
	);
	LUT2 #(
		.INIT('h1)
	) name1275 (
		_w5320_,
		_w5321_,
		_w5322_
	);
	LUT2 #(
		.INIT('h1)
	) name1276 (
		_w4104_,
		_w5322_,
		_w5323_
	);
	LUT2 #(
		.INIT('h1)
	) name1277 (
		_w5319_,
		_w5323_,
		_w5324_
	);
	LUT2 #(
		.INIT('h8)
	) name1278 (
		_w4120_,
		_w5324_,
		_w5325_
	);
	LUT2 #(
		.INIT('h1)
	) name1279 (
		_w4392_,
		_w5059_,
		_w5326_
	);
	LUT2 #(
		.INIT('h1)
	) name1280 (
		\core_c_psq_EXA_reg[6]/P0001 ,
		_w5086_,
		_w5327_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w5087_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h8)
	) name1282 (
		_w4835_,
		_w5328_,
		_w5329_
	);
	LUT2 #(
		.INIT('h1)
	) name1283 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w5099_,
		_w5330_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w5100_,
		_w5330_,
		_w5331_
	);
	LUT2 #(
		.INIT('h8)
	) name1285 (
		_w5050_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h8)
	) name1286 (
		_w4764_,
		_w4840_,
		_w5333_
	);
	LUT2 #(
		.INIT('h8)
	) name1287 (
		\sice_IRR_reg[6]/P0001 ,
		_w4837_,
		_w5334_
	);
	LUT2 #(
		.INIT('h1)
	) name1288 (
		_w5332_,
		_w5334_,
		_w5335_
	);
	LUT2 #(
		.INIT('h4)
	) name1289 (
		_w5333_,
		_w5335_,
		_w5336_
	);
	LUT2 #(
		.INIT('h4)
	) name1290 (
		_w5329_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h4)
	) name1291 (
		_w5326_,
		_w5337_,
		_w5338_
	);
	LUT2 #(
		.INIT('h2)
	) name1292 (
		_w4128_,
		_w5338_,
		_w5339_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w5066_,
		_w5340_
	);
	LUT2 #(
		.INIT('h8)
	) name1294 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w5068_,
		_w5341_
	);
	LUT2 #(
		.INIT('h1)
	) name1295 (
		_w5340_,
		_w5341_,
		_w5342_
	);
	LUT2 #(
		.INIT('h2)
	) name1296 (
		_w4099_,
		_w5342_,
		_w5343_
	);
	LUT2 #(
		.INIT('h1)
	) name1297 (
		_w5325_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h4)
	) name1298 (
		_w5339_,
		_w5344_,
		_w5345_
	);
	LUT2 #(
		.INIT('h4)
	) name1299 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w4104_,
		_w5346_
	);
	LUT2 #(
		.INIT('h1)
	) name1300 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w4117_,
		_w5347_
	);
	LUT2 #(
		.INIT('h4)
	) name1301 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w4117_,
		_w5348_
	);
	LUT2 #(
		.INIT('h1)
	) name1302 (
		_w5347_,
		_w5348_,
		_w5349_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		_w4104_,
		_w5349_,
		_w5350_
	);
	LUT2 #(
		.INIT('h1)
	) name1304 (
		_w5346_,
		_w5350_,
		_w5351_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		_w4120_,
		_w5351_,
		_w5352_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		_w4656_,
		_w5059_,
		_w5353_
	);
	LUT2 #(
		.INIT('h1)
	) name1307 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		_w5087_,
		_w5354_
	);
	LUT2 #(
		.INIT('h1)
	) name1308 (
		_w5088_,
		_w5354_,
		_w5355_
	);
	LUT2 #(
		.INIT('h8)
	) name1309 (
		_w4835_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h1)
	) name1310 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w5100_,
		_w5357_
	);
	LUT2 #(
		.INIT('h1)
	) name1311 (
		_w5101_,
		_w5357_,
		_w5358_
	);
	LUT2 #(
		.INIT('h8)
	) name1312 (
		_w5050_,
		_w5358_,
		_w5359_
	);
	LUT2 #(
		.INIT('h8)
	) name1313 (
		_w4783_,
		_w4840_,
		_w5360_
	);
	LUT2 #(
		.INIT('h8)
	) name1314 (
		\sice_IRR_reg[7]/P0001 ,
		_w4837_,
		_w5361_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		_w5359_,
		_w5361_,
		_w5362_
	);
	LUT2 #(
		.INIT('h4)
	) name1316 (
		_w5360_,
		_w5362_,
		_w5363_
	);
	LUT2 #(
		.INIT('h4)
	) name1317 (
		_w5356_,
		_w5363_,
		_w5364_
	);
	LUT2 #(
		.INIT('h4)
	) name1318 (
		_w5353_,
		_w5364_,
		_w5365_
	);
	LUT2 #(
		.INIT('h2)
	) name1319 (
		_w4128_,
		_w5365_,
		_w5366_
	);
	LUT2 #(
		.INIT('h8)
	) name1320 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w5066_,
		_w5367_
	);
	LUT2 #(
		.INIT('h8)
	) name1321 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w5068_,
		_w5368_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w5367_,
		_w5368_,
		_w5369_
	);
	LUT2 #(
		.INIT('h2)
	) name1323 (
		_w4099_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h1)
	) name1324 (
		_w5352_,
		_w5370_,
		_w5371_
	);
	LUT2 #(
		.INIT('h4)
	) name1325 (
		_w5366_,
		_w5371_,
		_w5372_
	);
	LUT2 #(
		.INIT('h4)
	) name1326 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w4104_,
		_w5373_
	);
	LUT2 #(
		.INIT('h1)
	) name1327 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w4117_,
		_w5374_
	);
	LUT2 #(
		.INIT('h4)
	) name1328 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w4117_,
		_w5375_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		_w5374_,
		_w5375_,
		_w5376_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w4104_,
		_w5376_,
		_w5377_
	);
	LUT2 #(
		.INIT('h1)
	) name1331 (
		_w5373_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h8)
	) name1332 (
		_w4120_,
		_w5378_,
		_w5379_
	);
	LUT2 #(
		.INIT('h1)
	) name1333 (
		_w4425_,
		_w5059_,
		_w5380_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		_w5088_,
		_w5381_
	);
	LUT2 #(
		.INIT('h1)
	) name1335 (
		_w5089_,
		_w5381_,
		_w5382_
	);
	LUT2 #(
		.INIT('h8)
	) name1336 (
		_w4835_,
		_w5382_,
		_w5383_
	);
	LUT2 #(
		.INIT('h1)
	) name1337 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w5101_,
		_w5384_
	);
	LUT2 #(
		.INIT('h1)
	) name1338 (
		_w5102_,
		_w5384_,
		_w5385_
	);
	LUT2 #(
		.INIT('h8)
	) name1339 (
		_w5050_,
		_w5385_,
		_w5386_
	);
	LUT2 #(
		.INIT('h8)
	) name1340 (
		_w4735_,
		_w4840_,
		_w5387_
	);
	LUT2 #(
		.INIT('h8)
	) name1341 (
		\sice_IRR_reg[8]/P0001 ,
		_w4837_,
		_w5388_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w5386_,
		_w5388_,
		_w5389_
	);
	LUT2 #(
		.INIT('h4)
	) name1343 (
		_w5387_,
		_w5389_,
		_w5390_
	);
	LUT2 #(
		.INIT('h4)
	) name1344 (
		_w5383_,
		_w5390_,
		_w5391_
	);
	LUT2 #(
		.INIT('h4)
	) name1345 (
		_w5380_,
		_w5391_,
		_w5392_
	);
	LUT2 #(
		.INIT('h2)
	) name1346 (
		_w4128_,
		_w5392_,
		_w5393_
	);
	LUT2 #(
		.INIT('h8)
	) name1347 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w5066_,
		_w5394_
	);
	LUT2 #(
		.INIT('h8)
	) name1348 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w5068_,
		_w5395_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		_w5394_,
		_w5395_,
		_w5396_
	);
	LUT2 #(
		.INIT('h2)
	) name1350 (
		_w4099_,
		_w5396_,
		_w5397_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		_w5379_,
		_w5397_,
		_w5398_
	);
	LUT2 #(
		.INIT('h4)
	) name1352 (
		_w5393_,
		_w5398_,
		_w5399_
	);
	LUT2 #(
		.INIT('h4)
	) name1353 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w4104_,
		_w5400_
	);
	LUT2 #(
		.INIT('h1)
	) name1354 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		_w4117_,
		_w5401_
	);
	LUT2 #(
		.INIT('h4)
	) name1355 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w4117_,
		_w5402_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		_w5401_,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h1)
	) name1357 (
		_w4104_,
		_w5403_,
		_w5404_
	);
	LUT2 #(
		.INIT('h1)
	) name1358 (
		_w5400_,
		_w5404_,
		_w5405_
	);
	LUT2 #(
		.INIT('h8)
	) name1359 (
		_w4120_,
		_w5405_,
		_w5406_
	);
	LUT2 #(
		.INIT('h1)
	) name1360 (
		_w4554_,
		_w5059_,
		_w5407_
	);
	LUT2 #(
		.INIT('h1)
	) name1361 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		_w5089_,
		_w5408_
	);
	LUT2 #(
		.INIT('h1)
	) name1362 (
		_w5090_,
		_w5408_,
		_w5409_
	);
	LUT2 #(
		.INIT('h8)
	) name1363 (
		_w4835_,
		_w5409_,
		_w5410_
	);
	LUT2 #(
		.INIT('h1)
	) name1364 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w5102_,
		_w5411_
	);
	LUT2 #(
		.INIT('h1)
	) name1365 (
		_w5103_,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		_w5050_,
		_w5412_,
		_w5413_
	);
	LUT2 #(
		.INIT('h8)
	) name1367 (
		_w4739_,
		_w4840_,
		_w5414_
	);
	LUT2 #(
		.INIT('h8)
	) name1368 (
		\sice_IRR_reg[9]/P0001 ,
		_w4837_,
		_w5415_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		_w5413_,
		_w5415_,
		_w5416_
	);
	LUT2 #(
		.INIT('h4)
	) name1370 (
		_w5414_,
		_w5416_,
		_w5417_
	);
	LUT2 #(
		.INIT('h4)
	) name1371 (
		_w5410_,
		_w5417_,
		_w5418_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w5407_,
		_w5418_,
		_w5419_
	);
	LUT2 #(
		.INIT('h2)
	) name1373 (
		_w4128_,
		_w5419_,
		_w5420_
	);
	LUT2 #(
		.INIT('h8)
	) name1374 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w5066_,
		_w5421_
	);
	LUT2 #(
		.INIT('h8)
	) name1375 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w5068_,
		_w5422_
	);
	LUT2 #(
		.INIT('h1)
	) name1376 (
		_w5421_,
		_w5422_,
		_w5423_
	);
	LUT2 #(
		.INIT('h2)
	) name1377 (
		_w4099_,
		_w5423_,
		_w5424_
	);
	LUT2 #(
		.INIT('h1)
	) name1378 (
		_w5406_,
		_w5424_,
		_w5425_
	);
	LUT2 #(
		.INIT('h4)
	) name1379 (
		_w5420_,
		_w5425_,
		_w5426_
	);
	LUT2 #(
		.INIT('h1)
	) name1380 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w5427_
	);
	LUT2 #(
		.INIT('h8)
	) name1381 (
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		_w5428_
	);
	LUT2 #(
		.INIT('h8)
	) name1382 (
		_w5427_,
		_w5428_,
		_w5429_
	);
	LUT2 #(
		.INIT('h2)
	) name1383 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w5430_
	);
	LUT2 #(
		.INIT('h4)
	) name1384 (
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		_w5431_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		_w5430_,
		_w5431_,
		_w5432_
	);
	LUT2 #(
		.INIT('h1)
	) name1386 (
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		_w5433_
	);
	LUT2 #(
		.INIT('h8)
	) name1387 (
		_w5430_,
		_w5433_,
		_w5434_
	);
	LUT2 #(
		.INIT('h2)
	) name1388 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		_w5435_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		\core_c_dec_Double_E_reg/P0001 ,
		_w5435_,
		_w5436_
	);
	LUT2 #(
		.INIT('h1)
	) name1390 (
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[1]/NET0131 ,
		_w5437_
	);
	LUT2 #(
		.INIT('h2)
	) name1391 (
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[3]/NET0131 ,
		_w5438_
	);
	LUT2 #(
		.INIT('h1)
	) name1392 (
		_w5437_,
		_w5438_,
		_w5439_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		\emc_DMcst_reg/NET0131 ,
		_w5439_,
		_w5440_
	);
	LUT2 #(
		.INIT('h2)
	) name1394 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[11]/NET0131 ,
		_w5441_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w5440_,
		_w5441_,
		_w5442_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		\emc_PMcst_reg/NET0131 ,
		_w5442_,
		_w5443_
	);
	LUT2 #(
		.INIT('h2)
	) name1397 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[7]/NET0131 ,
		_w5444_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w5443_,
		_w5444_,
		_w5445_
	);
	LUT2 #(
		.INIT('h4)
	) name1399 (
		\emc_RWcnt_reg[3]/P0001 ,
		_w5445_,
		_w5446_
	);
	LUT2 #(
		.INIT('h2)
	) name1400 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[4]/NET0131 ,
		_w5447_
	);
	LUT2 #(
		.INIT('h4)
	) name1401 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w5448_
	);
	LUT2 #(
		.INIT('h8)
	) name1402 (
		\emc_WSCRext_reg_DO_reg[2]/NET0131 ,
		_w5448_,
		_w5449_
	);
	LUT2 #(
		.INIT('h8)
	) name1403 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[6]/NET0131 ,
		_w5450_
	);
	LUT2 #(
		.INIT('h1)
	) name1404 (
		\emc_PMcst_reg/NET0131 ,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h4)
	) name1405 (
		_w5449_,
		_w5451_,
		_w5452_
	);
	LUT2 #(
		.INIT('h1)
	) name1406 (
		_w5447_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h1)
	) name1407 (
		\emc_RWcnt_reg[4]/P0001 ,
		_w5453_,
		_w5454_
	);
	LUT2 #(
		.INIT('h8)
	) name1408 (
		\emc_RWcnt_reg[4]/P0001 ,
		_w5453_,
		_w5455_
	);
	LUT2 #(
		.INIT('h1)
	) name1409 (
		_w5454_,
		_w5455_,
		_w5456_
	);
	LUT2 #(
		.INIT('h1)
	) name1410 (
		\emc_IOcst_reg/NET0131 ,
		\memc_usysr_DO_reg[15]/NET0131 ,
		_w5457_
	);
	LUT2 #(
		.INIT('h2)
	) name1411 (
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[1]/NET0131 ,
		_w5458_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		_w5457_,
		_w5458_,
		_w5459_
	);
	LUT2 #(
		.INIT('h1)
	) name1413 (
		\emc_DMcst_reg/NET0131 ,
		_w5459_,
		_w5460_
	);
	LUT2 #(
		.INIT('h2)
	) name1414 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[9]/NET0131 ,
		_w5461_
	);
	LUT2 #(
		.INIT('h1)
	) name1415 (
		_w5460_,
		_w5461_,
		_w5462_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		\emc_PMcst_reg/NET0131 ,
		_w5462_,
		_w5463_
	);
	LUT2 #(
		.INIT('h2)
	) name1417 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[5]/NET0131 ,
		_w5464_
	);
	LUT2 #(
		.INIT('h1)
	) name1418 (
		_w5463_,
		_w5464_,
		_w5465_
	);
	LUT2 #(
		.INIT('h2)
	) name1419 (
		\emc_RWcnt_reg[1]/P0001 ,
		_w5465_,
		_w5466_
	);
	LUT2 #(
		.INIT('h4)
	) name1420 (
		\emc_RWcnt_reg[1]/P0001 ,
		_w5465_,
		_w5467_
	);
	LUT2 #(
		.INIT('h1)
	) name1421 (
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[0]/NET0131 ,
		_w5468_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[2]/NET0131 ,
		_w5469_
	);
	LUT2 #(
		.INIT('h1)
	) name1423 (
		_w5468_,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		\emc_DMcst_reg/NET0131 ,
		_w5470_,
		_w5471_
	);
	LUT2 #(
		.INIT('h2)
	) name1425 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[10]/NET0131 ,
		_w5472_
	);
	LUT2 #(
		.INIT('h1)
	) name1426 (
		_w5471_,
		_w5472_,
		_w5473_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		\emc_PMcst_reg/NET0131 ,
		_w5473_,
		_w5474_
	);
	LUT2 #(
		.INIT('h2)
	) name1428 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[6]/NET0131 ,
		_w5475_
	);
	LUT2 #(
		.INIT('h1)
	) name1429 (
		_w5474_,
		_w5475_,
		_w5476_
	);
	LUT2 #(
		.INIT('h2)
	) name1430 (
		\emc_RWcnt_reg[2]/P0001 ,
		_w5476_,
		_w5477_
	);
	LUT2 #(
		.INIT('h4)
	) name1431 (
		\emc_RWcnt_reg[2]/P0001 ,
		_w5476_,
		_w5478_
	);
	LUT2 #(
		.INIT('h2)
	) name1432 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[5]/NET0131 ,
		_w5479_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		\emc_WSCRext_reg_DO_reg[3]/NET0131 ,
		_w5448_,
		_w5480_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRext_reg_DO_reg[7]/NET0131 ,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		\emc_PMcst_reg/NET0131 ,
		_w5481_,
		_w5482_
	);
	LUT2 #(
		.INIT('h4)
	) name1436 (
		_w5480_,
		_w5482_,
		_w5483_
	);
	LUT2 #(
		.INIT('h1)
	) name1437 (
		_w5479_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h4)
	) name1438 (
		\emc_RWcnt_reg[5]/P0001 ,
		_w5484_,
		_w5485_
	);
	LUT2 #(
		.INIT('h1)
	) name1439 (
		\emc_IOcst_reg/NET0131 ,
		\memc_usysr_DO_reg[14]/NET0131 ,
		_w5486_
	);
	LUT2 #(
		.INIT('h2)
	) name1440 (
		\emc_IOcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[0]/NET0131 ,
		_w5487_
	);
	LUT2 #(
		.INIT('h1)
	) name1441 (
		_w5486_,
		_w5487_,
		_w5488_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		\emc_DMcst_reg/NET0131 ,
		_w5488_,
		_w5489_
	);
	LUT2 #(
		.INIT('h2)
	) name1443 (
		\emc_DMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[8]/NET0131 ,
		_w5490_
	);
	LUT2 #(
		.INIT('h1)
	) name1444 (
		_w5489_,
		_w5490_,
		_w5491_
	);
	LUT2 #(
		.INIT('h1)
	) name1445 (
		\emc_PMcst_reg/NET0131 ,
		_w5491_,
		_w5492_
	);
	LUT2 #(
		.INIT('h2)
	) name1446 (
		\emc_PMcst_reg/NET0131 ,
		\emc_WSCRreg_DO_reg[4]/NET0131 ,
		_w5493_
	);
	LUT2 #(
		.INIT('h1)
	) name1447 (
		_w5492_,
		_w5493_,
		_w5494_
	);
	LUT2 #(
		.INIT('h4)
	) name1448 (
		\emc_RWcnt_reg[0]/P0001 ,
		_w5494_,
		_w5495_
	);
	LUT2 #(
		.INIT('h2)
	) name1449 (
		\emc_RWcnt_reg[5]/P0001 ,
		_w5484_,
		_w5496_
	);
	LUT2 #(
		.INIT('h2)
	) name1450 (
		\emc_RWcnt_reg[0]/P0001 ,
		_w5494_,
		_w5497_
	);
	LUT2 #(
		.INIT('h2)
	) name1451 (
		\emc_RWcnt_reg[3]/P0001 ,
		_w5445_,
		_w5498_
	);
	LUT2 #(
		.INIT('h1)
	) name1452 (
		_w5485_,
		_w5496_,
		_w5499_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		_w5456_,
		_w5499_,
		_w5500_
	);
	LUT2 #(
		.INIT('h4)
	) name1454 (
		_w5446_,
		_w5500_,
		_w5501_
	);
	LUT2 #(
		.INIT('h1)
	) name1455 (
		_w5466_,
		_w5467_,
		_w5502_
	);
	LUT2 #(
		.INIT('h1)
	) name1456 (
		_w5477_,
		_w5478_,
		_w5503_
	);
	LUT2 #(
		.INIT('h1)
	) name1457 (
		_w5495_,
		_w5497_,
		_w5504_
	);
	LUT2 #(
		.INIT('h4)
	) name1458 (
		_w5498_,
		_w5504_,
		_w5505_
	);
	LUT2 #(
		.INIT('h8)
	) name1459 (
		_w5502_,
		_w5503_,
		_w5506_
	);
	LUT2 #(
		.INIT('h8)
	) name1460 (
		_w5501_,
		_w5506_,
		_w5507_
	);
	LUT2 #(
		.INIT('h8)
	) name1461 (
		_w5505_,
		_w5507_,
		_w5508_
	);
	LUT2 #(
		.INIT('h4)
	) name1462 (
		_w5436_,
		_w5508_,
		_w5509_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		_w5434_,
		_w5509_,
		_w5510_
	);
	LUT2 #(
		.INIT('h1)
	) name1464 (
		\emc_DMcst_reg/NET0131 ,
		\emc_IOcst_reg/NET0131 ,
		_w5511_
	);
	LUT2 #(
		.INIT('h4)
	) name1465 (
		\emc_PMcst_reg/NET0131 ,
		_w5511_,
		_w5512_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		\core_c_psq_ECYC_reg/P0001 ,
		\emc_eRDY_reg/NET0131 ,
		_w5513_
	);
	LUT2 #(
		.INIT('h4)
	) name1467 (
		_w5512_,
		_w5513_,
		_w5514_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		\emc_ECS_reg[2]/NET0131 ,
		_w5514_,
		_w5515_
	);
	LUT2 #(
		.INIT('h4)
	) name1469 (
		\emc_ECS_reg[1]/NET0131 ,
		_w5427_,
		_w5516_
	);
	LUT2 #(
		.INIT('h4)
	) name1470 (
		_w5515_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('h8)
	) name1471 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w5518_
	);
	LUT2 #(
		.INIT('h8)
	) name1472 (
		_w5433_,
		_w5518_,
		_w5519_
	);
	LUT2 #(
		.INIT('h1)
	) name1473 (
		_w5432_,
		_w5519_,
		_w5520_
	);
	LUT2 #(
		.INIT('h1)
	) name1474 (
		_w5508_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		\emc_ECS_reg[0]/NET0131 ,
		\emc_ECS_reg[3]/NET0131 ,
		_w5522_
	);
	LUT2 #(
		.INIT('h4)
	) name1476 (
		\emc_ECS_reg[2]/NET0131 ,
		_w5522_,
		_w5523_
	);
	LUT2 #(
		.INIT('h8)
	) name1477 (
		_w5508_,
		_w5523_,
		_w5524_
	);
	LUT2 #(
		.INIT('h1)
	) name1478 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[4]/NET0131 ,
		_w5525_
	);
	LUT2 #(
		.INIT('h2)
	) name1479 (
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w5525_,
		_w5526_
	);
	LUT2 #(
		.INIT('h4)
	) name1480 (
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w5525_,
		_w5527_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		_w5526_,
		_w5527_,
		_w5528_
	);
	LUT2 #(
		.INIT('h2)
	) name1482 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[7]/NET0131 ,
		_w5529_
	);
	LUT2 #(
		.INIT('h2)
	) name1483 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w5529_,
		_w5530_
	);
	LUT2 #(
		.INIT('h4)
	) name1484 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w5529_,
		_w5531_
	);
	LUT2 #(
		.INIT('h1)
	) name1485 (
		_w5530_,
		_w5531_,
		_w5532_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w5528_,
		_w5532_,
		_w5533_
	);
	LUT2 #(
		.INIT('h8)
	) name1487 (
		_w5431_,
		_w5522_,
		_w5534_
	);
	LUT2 #(
		.INIT('h2)
	) name1488 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[4]/NET0131 ,
		_w5535_
	);
	LUT2 #(
		.INIT('h1)
	) name1489 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		_w5536_
	);
	LUT2 #(
		.INIT('h1)
	) name1490 (
		_w5535_,
		_w5536_,
		_w5537_
	);
	LUT2 #(
		.INIT('h1)
	) name1491 (
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h8)
	) name1492 (
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w5537_,
		_w5539_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		_w5538_,
		_w5539_,
		_w5540_
	);
	LUT2 #(
		.INIT('h2)
	) name1494 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		_w5541_
	);
	LUT2 #(
		.INIT('h1)
	) name1495 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[6]/NET0131 ,
		_w5542_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		_w5541_,
		_w5542_,
		_w5543_
	);
	LUT2 #(
		.INIT('h2)
	) name1497 (
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w5543_,
		_w5544_
	);
	LUT2 #(
		.INIT('h4)
	) name1498 (
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w5543_,
		_w5545_
	);
	LUT2 #(
		.INIT('h2)
	) name1499 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[6]/NET0131 ,
		_w5546_
	);
	LUT2 #(
		.INIT('h1)
	) name1500 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BCTL_reg[7]/NET0131 ,
		_w5547_
	);
	LUT2 #(
		.INIT('h1)
	) name1501 (
		_w5546_,
		_w5547_,
		_w5548_
	);
	LUT2 #(
		.INIT('h2)
	) name1502 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w5548_,
		_w5549_
	);
	LUT2 #(
		.INIT('h4)
	) name1503 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w5548_,
		_w5550_
	);
	LUT2 #(
		.INIT('h1)
	) name1504 (
		_w5544_,
		_w5545_,
		_w5551_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		_w5549_,
		_w5550_,
		_w5552_
	);
	LUT2 #(
		.INIT('h8)
	) name1506 (
		_w5551_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h4)
	) name1507 (
		_w5540_,
		_w5553_,
		_w5554_
	);
	LUT2 #(
		.INIT('h8)
	) name1508 (
		_w5533_,
		_w5534_,
		_w5555_
	);
	LUT2 #(
		.INIT('h8)
	) name1509 (
		_w5554_,
		_w5555_,
		_w5556_
	);
	LUT2 #(
		.INIT('h1)
	) name1510 (
		_w5517_,
		_w5556_,
		_w5557_
	);
	LUT2 #(
		.INIT('h4)
	) name1511 (
		_w5521_,
		_w5557_,
		_w5558_
	);
	LUT2 #(
		.INIT('h4)
	) name1512 (
		_w5524_,
		_w5558_,
		_w5559_
	);
	LUT2 #(
		.INIT('h4)
	) name1513 (
		_w5510_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		_w5431_,
		_w5518_,
		_w5561_
	);
	LUT2 #(
		.INIT('h8)
	) name1515 (
		\bdma_BSreq_reg/NET0131 ,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h8)
	) name1516 (
		_w5428_,
		_w5522_,
		_w5563_
	);
	LUT2 #(
		.INIT('h4)
	) name1517 (
		\auctl_BSack_reg/NET0131 ,
		_w5563_,
		_w5564_
	);
	LUT2 #(
		.INIT('h1)
	) name1518 (
		_w5562_,
		_w5564_,
		_w5565_
	);
	LUT2 #(
		.INIT('h4)
	) name1519 (
		\T_TMODE[1]_pad ,
		\bdma_BDMAmode_reg/NET0131 ,
		_w5566_
	);
	LUT2 #(
		.INIT('h4)
	) name1520 (
		\core_c_psq_ECYC_reg/P0001 ,
		_w5566_,
		_w5567_
	);
	LUT2 #(
		.INIT('h8)
	) name1521 (
		\T_TMODE[1]_pad ,
		\core_c_psq_ECYC_reg/P0001 ,
		_w5568_
	);
	LUT2 #(
		.INIT('h1)
	) name1522 (
		_w5567_,
		_w5568_,
		_w5569_
	);
	LUT2 #(
		.INIT('h1)
	) name1523 (
		\emc_PMcst_reg/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w5570_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		_w5427_,
		_w5570_,
		_w5571_
	);
	LUT2 #(
		.INIT('h8)
	) name1525 (
		_w5433_,
		_w5571_,
		_w5572_
	);
	LUT2 #(
		.INIT('h2)
	) name1526 (
		_w5511_,
		_w5569_,
		_w5573_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		_w5572_,
		_w5573_,
		_w5574_
	);
	LUT2 #(
		.INIT('h8)
	) name1528 (
		\T_TMODE[1]_pad ,
		\emc_ECS_reg[1]/NET0131 ,
		_w5575_
	);
	LUT2 #(
		.INIT('h8)
	) name1529 (
		_w5427_,
		_w5575_,
		_w5576_
	);
	LUT2 #(
		.INIT('h1)
	) name1530 (
		_w5519_,
		_w5523_,
		_w5577_
	);
	LUT2 #(
		.INIT('h1)
	) name1531 (
		_w5534_,
		_w5576_,
		_w5578_
	);
	LUT2 #(
		.INIT('h8)
	) name1532 (
		_w5577_,
		_w5578_,
		_w5579_
	);
	LUT2 #(
		.INIT('h8)
	) name1533 (
		_w5565_,
		_w5579_,
		_w5580_
	);
	LUT2 #(
		.INIT('h4)
	) name1534 (
		_w5574_,
		_w5580_,
		_w5581_
	);
	LUT2 #(
		.INIT('h8)
	) name1535 (
		\emc_ECS_reg[1]/NET0131 ,
		_w5523_,
		_w5582_
	);
	LUT2 #(
		.INIT('h4)
	) name1536 (
		_w5434_,
		_w5520_,
		_w5583_
	);
	LUT2 #(
		.INIT('h2)
	) name1537 (
		_w5508_,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		_w5565_,
		_w5582_,
		_w5585_
	);
	LUT2 #(
		.INIT('h4)
	) name1539 (
		_w5584_,
		_w5585_,
		_w5586_
	);
	LUT2 #(
		.INIT('h8)
	) name1540 (
		_w5581_,
		_w5586_,
		_w5587_
	);
	LUT2 #(
		.INIT('h1)
	) name1541 (
		\core_c_psq_ECYC_reg/P0001 ,
		_w5511_,
		_w5588_
	);
	LUT2 #(
		.INIT('h2)
	) name1542 (
		_w5511_,
		_w5567_,
		_w5589_
	);
	LUT2 #(
		.INIT('h2)
	) name1543 (
		_w5572_,
		_w5588_,
		_w5590_
	);
	LUT2 #(
		.INIT('h4)
	) name1544 (
		_w5589_,
		_w5590_,
		_w5591_
	);
	LUT2 #(
		.INIT('h2)
	) name1545 (
		\emc_ECS_reg[1]/NET0131 ,
		\emc_ECS_reg[2]/NET0131 ,
		_w5592_
	);
	LUT2 #(
		.INIT('h8)
	) name1546 (
		_w5430_,
		_w5592_,
		_w5593_
	);
	LUT2 #(
		.INIT('h2)
	) name1547 (
		_w5431_,
		_w5518_,
		_w5594_
	);
	LUT2 #(
		.INIT('h1)
	) name1548 (
		_w5593_,
		_w5594_,
		_w5595_
	);
	LUT2 #(
		.INIT('h8)
	) name1549 (
		_w5565_,
		_w5595_,
		_w5596_
	);
	LUT2 #(
		.INIT('h4)
	) name1550 (
		_w5591_,
		_w5596_,
		_w5597_
	);
	LUT2 #(
		.INIT('h2)
	) name1551 (
		_w5587_,
		_w5597_,
		_w5598_
	);
	LUT2 #(
		.INIT('h4)
	) name1552 (
		_w5560_,
		_w5598_,
		_w5599_
	);
	LUT2 #(
		.INIT('h1)
	) name1553 (
		_w5432_,
		_w5599_,
		_w5600_
	);
	LUT2 #(
		.INIT('h4)
	) name1554 (
		_w5429_,
		_w5600_,
		_w5601_
	);
	LUT2 #(
		.INIT('h2)
	) name1555 (
		\emc_DMcst_reg/NET0131 ,
		_w5601_,
		_w5602_
	);
	LUT2 #(
		.INIT('h8)
	) name1556 (
		\emc_WSCRreg_DO_reg[13]/NET0131 ,
		_w5602_,
		_w5603_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		_w5427_,
		_w5592_,
		_w5604_
	);
	LUT2 #(
		.INIT('h4)
	) name1558 (
		_w5560_,
		_w5597_,
		_w5605_
	);
	LUT2 #(
		.INIT('h8)
	) name1559 (
		_w5587_,
		_w5605_,
		_w5606_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w5434_,
		_w5606_,
		_w5607_
	);
	LUT2 #(
		.INIT('h4)
	) name1561 (
		_w5604_,
		_w5607_,
		_w5608_
	);
	LUT2 #(
		.INIT('h2)
	) name1562 (
		\emc_WSCRreg_DO_reg[12]/NET0131 ,
		_w5608_,
		_w5609_
	);
	LUT2 #(
		.INIT('h2)
	) name1563 (
		\emc_IOcst_reg/NET0131 ,
		_w5601_,
		_w5610_
	);
	LUT2 #(
		.INIT('h8)
	) name1564 (
		\emc_WSCRreg_DO_reg[14]/NET0131 ,
		_w5610_,
		_w5611_
	);
	LUT2 #(
		.INIT('h1)
	) name1565 (
		_w5603_,
		_w5609_,
		_w5612_
	);
	LUT2 #(
		.INIT('h4)
	) name1566 (
		_w5611_,
		_w5612_,
		_w5613_
	);
	LUT2 #(
		.INIT('h4)
	) name1567 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w4104_,
		_w5614_
	);
	LUT2 #(
		.INIT('h1)
	) name1568 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w4117_,
		_w5615_
	);
	LUT2 #(
		.INIT('h4)
	) name1569 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w4117_,
		_w5616_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		_w5615_,
		_w5616_,
		_w5617_
	);
	LUT2 #(
		.INIT('h1)
	) name1571 (
		_w4104_,
		_w5617_,
		_w5618_
	);
	LUT2 #(
		.INIT('h1)
	) name1572 (
		_w5614_,
		_w5618_,
		_w5619_
	);
	LUT2 #(
		.INIT('h8)
	) name1573 (
		_w4120_,
		_w5619_,
		_w5620_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		_w4694_,
		_w5059_,
		_w5621_
	);
	LUT2 #(
		.INIT('h8)
	) name1575 (
		\core_c_psq_EXA_reg[12]/P0001 ,
		_w5130_,
		_w5622_
	);
	LUT2 #(
		.INIT('h1)
	) name1576 (
		\core_c_psq_EXA_reg[12]/P0001 ,
		_w5130_,
		_w5623_
	);
	LUT2 #(
		.INIT('h1)
	) name1577 (
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h8)
	) name1578 (
		_w4835_,
		_w5624_,
		_w5625_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w5134_,
		_w5626_
	);
	LUT2 #(
		.INIT('h1)
	) name1580 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w5134_,
		_w5627_
	);
	LUT2 #(
		.INIT('h1)
	) name1581 (
		_w5626_,
		_w5627_,
		_w5628_
	);
	LUT2 #(
		.INIT('h8)
	) name1582 (
		_w5050_,
		_w5628_,
		_w5629_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		_w4790_,
		_w4840_,
		_w5630_
	);
	LUT2 #(
		.INIT('h8)
	) name1584 (
		\sice_IRR_reg[12]/P0001 ,
		_w4837_,
		_w5631_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		_w5629_,
		_w5631_,
		_w5632_
	);
	LUT2 #(
		.INIT('h4)
	) name1586 (
		_w5630_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h4)
	) name1587 (
		_w5625_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h4)
	) name1588 (
		_w5621_,
		_w5634_,
		_w5635_
	);
	LUT2 #(
		.INIT('h2)
	) name1589 (
		_w4128_,
		_w5635_,
		_w5636_
	);
	LUT2 #(
		.INIT('h8)
	) name1590 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w5066_,
		_w5637_
	);
	LUT2 #(
		.INIT('h8)
	) name1591 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w5068_,
		_w5638_
	);
	LUT2 #(
		.INIT('h1)
	) name1592 (
		_w5637_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('h2)
	) name1593 (
		_w4099_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h1)
	) name1594 (
		_w5620_,
		_w5640_,
		_w5641_
	);
	LUT2 #(
		.INIT('h4)
	) name1595 (
		_w5636_,
		_w5641_,
		_w5642_
	);
	LUT2 #(
		.INIT('h2)
	) name1596 (
		PM_bdry_sel_pad,
		_w5642_,
		_w5643_
	);
	LUT2 #(
		.INIT('h4)
	) name1597 (
		_w4098_,
		_w5066_,
		_w5644_
	);
	LUT2 #(
		.INIT('h8)
	) name1598 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w5644_,
		_w5645_
	);
	LUT2 #(
		.INIT('h1)
	) name1599 (
		_w4489_,
		_w5059_,
		_w5646_
	);
	LUT2 #(
		.INIT('h1)
	) name1600 (
		\core_c_psq_EXA_reg[13]/P0001 ,
		_w5622_,
		_w5647_
	);
	LUT2 #(
		.INIT('h8)
	) name1601 (
		\core_c_psq_EXA_reg[13]/P0001 ,
		_w5622_,
		_w5648_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		_w5647_,
		_w5648_,
		_w5649_
	);
	LUT2 #(
		.INIT('h8)
	) name1603 (
		_w4835_,
		_w5649_,
		_w5650_
	);
	LUT2 #(
		.INIT('h8)
	) name1604 (
		_w4786_,
		_w4840_,
		_w5651_
	);
	LUT2 #(
		.INIT('h8)
	) name1605 (
		\sice_IRR_reg[13]/P0001 ,
		_w4837_,
		_w5652_
	);
	LUT2 #(
		.INIT('h1)
	) name1606 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w5626_,
		_w5653_
	);
	LUT2 #(
		.INIT('h8)
	) name1607 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w5626_,
		_w5654_
	);
	LUT2 #(
		.INIT('h1)
	) name1608 (
		_w5653_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h8)
	) name1609 (
		_w5050_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h1)
	) name1610 (
		_w5651_,
		_w5652_,
		_w5657_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		_w5656_,
		_w5657_,
		_w5658_
	);
	LUT2 #(
		.INIT('h4)
	) name1612 (
		_w5650_,
		_w5658_,
		_w5659_
	);
	LUT2 #(
		.INIT('h4)
	) name1613 (
		_w5646_,
		_w5659_,
		_w5660_
	);
	LUT2 #(
		.INIT('h2)
	) name1614 (
		_w4128_,
		_w5660_,
		_w5661_
	);
	LUT2 #(
		.INIT('h4)
	) name1615 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w4104_,
		_w5662_
	);
	LUT2 #(
		.INIT('h8)
	) name1616 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w4117_,
		_w5663_
	);
	LUT2 #(
		.INIT('h2)
	) name1617 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w4117_,
		_w5664_
	);
	LUT2 #(
		.INIT('h1)
	) name1618 (
		_w4104_,
		_w5663_,
		_w5665_
	);
	LUT2 #(
		.INIT('h4)
	) name1619 (
		_w5664_,
		_w5665_,
		_w5666_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w5662_,
		_w5666_,
		_w5667_
	);
	LUT2 #(
		.INIT('h8)
	) name1621 (
		_w4120_,
		_w5667_,
		_w5668_
	);
	LUT2 #(
		.INIT('h8)
	) name1622 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w5068_,
		_w5669_
	);
	LUT2 #(
		.INIT('h8)
	) name1623 (
		_w4099_,
		_w5669_,
		_w5670_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w5645_,
		_w5670_,
		_w5671_
	);
	LUT2 #(
		.INIT('h4)
	) name1625 (
		_w5668_,
		_w5671_,
		_w5672_
	);
	LUT2 #(
		.INIT('h4)
	) name1626 (
		_w5661_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h4)
	) name1627 (
		_w5643_,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h2)
	) name1628 (
		\core_c_psq_PCS_reg[6]/NET0131 ,
		_w4075_,
		_w5675_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		\core_c_psq_PCS_reg[2]/NET0131 ,
		_w4107_,
		_w5676_
	);
	LUT2 #(
		.INIT('h8)
	) name1630 (
		\core_c_dec_IDLE_Eg_reg/P0001 ,
		_w4082_,
		_w5677_
	);
	LUT2 #(
		.INIT('h4)
	) name1631 (
		_w5676_,
		_w5677_,
		_w5678_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		_w5675_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		_w4104_,
		_w5679_,
		_w5680_
	);
	LUT2 #(
		.INIT('h8)
	) name1634 (
		\clkc_Cnt4096_s1_reg/NET0131 ,
		\clkc_Cnt4096_s2_reg/NET0131 ,
		_w5681_
	);
	LUT2 #(
		.INIT('h2)
	) name1635 (
		_w4115_,
		_w5681_,
		_w5682_
	);
	LUT2 #(
		.INIT('h4)
	) name1636 (
		_w5068_,
		_w5682_,
		_w5683_
	);
	LUT2 #(
		.INIT('h4)
	) name1637 (
		_w5066_,
		_w5683_,
		_w5684_
	);
	LUT2 #(
		.INIT('h4)
	) name1638 (
		\core_c_psq_MGNT_reg/NET0131 ,
		\core_c_psq_PCS_reg[10]/NET0131 ,
		_w5685_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[11]/NET0131 ,
		_w5686_
	);
	LUT2 #(
		.INIT('h2)
	) name1640 (
		_w4085_,
		_w5686_,
		_w5687_
	);
	LUT2 #(
		.INIT('h1)
	) name1641 (
		_w5685_,
		_w5687_,
		_w5688_
	);
	LUT2 #(
		.INIT('h2)
	) name1642 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w5688_,
		_w5689_
	);
	LUT2 #(
		.INIT('h4)
	) name1643 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[5]/NET0131 ,
		_w5690_
	);
	LUT2 #(
		.INIT('h4)
	) name1644 (
		\memc_STI_Cg_reg/NET0131 ,
		_w5690_,
		_w5691_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		\core_c_psq_PCS_reg[11]/NET0131 ,
		_w5691_,
		_w5692_
	);
	LUT2 #(
		.INIT('h8)
	) name1646 (
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\memc_LDaST_Eg_reg/NET0131 ,
		_w5693_
	);
	LUT2 #(
		.INIT('h8)
	) name1647 (
		_w4085_,
		_w5693_,
		_w5694_
	);
	LUT2 #(
		.INIT('h2)
	) name1648 (
		_w5692_,
		_w5694_,
		_w5695_
	);
	LUT2 #(
		.INIT('h4)
	) name1649 (
		_w5689_,
		_w5695_,
		_w5696_
	);
	LUT2 #(
		.INIT('h2)
	) name1650 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w5697_
	);
	LUT2 #(
		.INIT('h2)
	) name1651 (
		\core_c_psq_PCS_reg[10]/NET0131 ,
		_w4068_,
		_w5698_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		_w4105_,
		_w5698_,
		_w5699_
	);
	LUT2 #(
		.INIT('h1)
	) name1653 (
		_w5697_,
		_w5699_,
		_w5700_
	);
	LUT2 #(
		.INIT('h8)
	) name1654 (
		\core_c_psq_MGNT_reg/NET0131 ,
		\core_c_psq_PCS_reg[10]/NET0131 ,
		_w5701_
	);
	LUT2 #(
		.INIT('h8)
	) name1655 (
		\core_c_psq_PCS_reg[0]/NET0131 ,
		_w4105_,
		_w5702_
	);
	LUT2 #(
		.INIT('h1)
	) name1656 (
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[13]/NET0131 ,
		_w5703_
	);
	LUT2 #(
		.INIT('h2)
	) name1657 (
		_w4084_,
		_w5703_,
		_w5704_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		_w5704_,
		_w5705_
	);
	LUT2 #(
		.INIT('h4)
	) name1659 (
		_w5702_,
		_w5705_,
		_w5706_
	);
	LUT2 #(
		.INIT('h2)
	) name1660 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w5706_,
		_w5707_
	);
	LUT2 #(
		.INIT('h1)
	) name1661 (
		_w5701_,
		_w5707_,
		_w5708_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_c_psq_PCS_reg[8]/NET0131 ,
		_w5709_
	);
	LUT2 #(
		.INIT('h4)
	) name1663 (
		_w4079_,
		_w5709_,
		_w5710_
	);
	LUT2 #(
		.INIT('h4)
	) name1664 (
		_w4087_,
		_w5710_,
		_w5711_
	);
	LUT2 #(
		.INIT('h1)
	) name1665 (
		_w4068_,
		_w5711_,
		_w5712_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		_w5700_,
		_w5712_,
		_w5713_
	);
	LUT2 #(
		.INIT('h8)
	) name1667 (
		_w5696_,
		_w5713_,
		_w5714_
	);
	LUT2 #(
		.INIT('h8)
	) name1668 (
		_w5708_,
		_w5714_,
		_w5715_
	);
	LUT2 #(
		.INIT('h4)
	) name1669 (
		\sice_GO_NX_reg/NET0131 ,
		_w4096_,
		_w5716_
	);
	LUT2 #(
		.INIT('h8)
	) name1670 (
		_w4064_,
		_w5716_,
		_w5717_
	);
	LUT2 #(
		.INIT('h4)
	) name1671 (
		_w4065_,
		_w5717_,
		_w5718_
	);
	LUT2 #(
		.INIT('h8)
	) name1672 (
		_w4116_,
		_w5679_,
		_w5719_
	);
	LUT2 #(
		.INIT('h8)
	) name1673 (
		_w5715_,
		_w5719_,
		_w5720_
	);
	LUT2 #(
		.INIT('h8)
	) name1674 (
		_w5718_,
		_w5720_,
		_w5721_
	);
	LUT2 #(
		.INIT('h1)
	) name1675 (
		\T_TMODE[1]_pad ,
		_w5680_,
		_w5722_
	);
	LUT2 #(
		.INIT('h4)
	) name1676 (
		_w5684_,
		_w5722_,
		_w5723_
	);
	LUT2 #(
		.INIT('h4)
	) name1677 (
		_w5721_,
		_w5723_,
		_w5724_
	);
	LUT2 #(
		.INIT('h8)
	) name1678 (
		_w5674_,
		_w5724_,
		_w5725_
	);
	LUT2 #(
		.INIT('h1)
	) name1679 (
		PM_bdry_sel_pad,
		\bdma_BIAD_reg[12]/NET0131 ,
		_w5726_
	);
	LUT2 #(
		.INIT('h2)
	) name1680 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w5726_,
		_w5727_
	);
	LUT2 #(
		.INIT('h8)
	) name1681 (
		\bdma_BDMAmode_reg/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w5728_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		_w5729_
	);
	LUT2 #(
		.INIT('h8)
	) name1683 (
		_w5728_,
		_w5729_,
		_w5730_
	);
	LUT2 #(
		.INIT('h4)
	) name1684 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w5731_
	);
	LUT2 #(
		.INIT('h4)
	) name1685 (
		_w5727_,
		_w5731_,
		_w5732_
	);
	LUT2 #(
		.INIT('h8)
	) name1686 (
		_w5730_,
		_w5732_,
		_w5733_
	);
	LUT2 #(
		.INIT('h4)
	) name1687 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w5733_,
		_w5734_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		_w5066_,
		_w5734_,
		_w5735_
	);
	LUT2 #(
		.INIT('h2)
	) name1689 (
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w5735_,
		_w5736_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		\bdma_BRdataBUF_reg[0]/P0001 ,
		_w5735_,
		_w5737_
	);
	LUT2 #(
		.INIT('h1)
	) name1691 (
		_w5736_,
		_w5737_,
		_w5738_
	);
	LUT2 #(
		.INIT('h1)
	) name1692 (
		_w5068_,
		_w5738_,
		_w5739_
	);
	LUT2 #(
		.INIT('h8)
	) name1693 (
		\idma_DTMP_L_reg[0]/P0001 ,
		_w5068_,
		_w5740_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w5739_,
		_w5740_,
		_w5741_
	);
	LUT2 #(
		.INIT('h2)
	) name1695 (
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w5735_,
		_w5742_
	);
	LUT2 #(
		.INIT('h8)
	) name1696 (
		\bdma_BRdataBUF_reg[10]/P0001 ,
		_w5735_,
		_w5743_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		_w5742_,
		_w5743_,
		_w5744_
	);
	LUT2 #(
		.INIT('h1)
	) name1698 (
		_w5068_,
		_w5744_,
		_w5745_
	);
	LUT2 #(
		.INIT('h8)
	) name1699 (
		\idma_DTMP_H_reg[2]/P0001 ,
		_w5068_,
		_w5746_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w5745_,
		_w5746_,
		_w5747_
	);
	LUT2 #(
		.INIT('h2)
	) name1701 (
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w5735_,
		_w5748_
	);
	LUT2 #(
		.INIT('h8)
	) name1702 (
		\bdma_BRdataBUF_reg[11]/P0001 ,
		_w5735_,
		_w5749_
	);
	LUT2 #(
		.INIT('h1)
	) name1703 (
		_w5748_,
		_w5749_,
		_w5750_
	);
	LUT2 #(
		.INIT('h1)
	) name1704 (
		_w5068_,
		_w5750_,
		_w5751_
	);
	LUT2 #(
		.INIT('h8)
	) name1705 (
		\idma_DTMP_H_reg[3]/P0001 ,
		_w5068_,
		_w5752_
	);
	LUT2 #(
		.INIT('h1)
	) name1706 (
		_w5751_,
		_w5752_,
		_w5753_
	);
	LUT2 #(
		.INIT('h2)
	) name1707 (
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w5735_,
		_w5754_
	);
	LUT2 #(
		.INIT('h8)
	) name1708 (
		\bdma_BRdataBUF_reg[12]/P0001 ,
		_w5735_,
		_w5755_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w5754_,
		_w5755_,
		_w5756_
	);
	LUT2 #(
		.INIT('h1)
	) name1710 (
		_w5068_,
		_w5756_,
		_w5757_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		\idma_DTMP_H_reg[4]/P0001 ,
		_w5068_,
		_w5758_
	);
	LUT2 #(
		.INIT('h1)
	) name1712 (
		_w5757_,
		_w5758_,
		_w5759_
	);
	LUT2 #(
		.INIT('h2)
	) name1713 (
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w5735_,
		_w5760_
	);
	LUT2 #(
		.INIT('h8)
	) name1714 (
		\bdma_BRdataBUF_reg[13]/P0001 ,
		_w5735_,
		_w5761_
	);
	LUT2 #(
		.INIT('h1)
	) name1715 (
		_w5760_,
		_w5761_,
		_w5762_
	);
	LUT2 #(
		.INIT('h1)
	) name1716 (
		_w5068_,
		_w5762_,
		_w5763_
	);
	LUT2 #(
		.INIT('h8)
	) name1717 (
		\idma_DTMP_H_reg[5]/P0001 ,
		_w5068_,
		_w5764_
	);
	LUT2 #(
		.INIT('h1)
	) name1718 (
		_w5763_,
		_w5764_,
		_w5765_
	);
	LUT2 #(
		.INIT('h2)
	) name1719 (
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w5735_,
		_w5766_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		\bdma_BRdataBUF_reg[14]/P0001 ,
		_w5735_,
		_w5767_
	);
	LUT2 #(
		.INIT('h1)
	) name1721 (
		_w5766_,
		_w5767_,
		_w5768_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w5068_,
		_w5768_,
		_w5769_
	);
	LUT2 #(
		.INIT('h8)
	) name1723 (
		\idma_DTMP_H_reg[6]/P0001 ,
		_w5068_,
		_w5770_
	);
	LUT2 #(
		.INIT('h1)
	) name1724 (
		_w5769_,
		_w5770_,
		_w5771_
	);
	LUT2 #(
		.INIT('h2)
	) name1725 (
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w5735_,
		_w5772_
	);
	LUT2 #(
		.INIT('h8)
	) name1726 (
		\bdma_BRdataBUF_reg[15]/P0001 ,
		_w5735_,
		_w5773_
	);
	LUT2 #(
		.INIT('h1)
	) name1727 (
		_w5772_,
		_w5773_,
		_w5774_
	);
	LUT2 #(
		.INIT('h1)
	) name1728 (
		_w5068_,
		_w5774_,
		_w5775_
	);
	LUT2 #(
		.INIT('h8)
	) name1729 (
		\idma_DTMP_H_reg[7]/P0001 ,
		_w5068_,
		_w5776_
	);
	LUT2 #(
		.INIT('h1)
	) name1730 (
		_w5775_,
		_w5776_,
		_w5777_
	);
	LUT2 #(
		.INIT('h2)
	) name1731 (
		\sice_idr1_reg_DO_reg[4]/P0001 ,
		_w5735_,
		_w5778_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		\bdma_BRdataBUF_reg[16]/P0001 ,
		_w5735_,
		_w5779_
	);
	LUT2 #(
		.INIT('h1)
	) name1733 (
		_w5778_,
		_w5779_,
		_w5780_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w5068_,
		_w5780_,
		_w5781_
	);
	LUT2 #(
		.INIT('h8)
	) name1735 (
		\idma_DTMP_H_reg[8]/P0001 ,
		_w5068_,
		_w5782_
	);
	LUT2 #(
		.INIT('h1)
	) name1736 (
		_w5781_,
		_w5782_,
		_w5783_
	);
	LUT2 #(
		.INIT('h2)
	) name1737 (
		\sice_idr1_reg_DO_reg[5]/P0001 ,
		_w5735_,
		_w5784_
	);
	LUT2 #(
		.INIT('h8)
	) name1738 (
		\bdma_BRdataBUF_reg[17]/P0001 ,
		_w5735_,
		_w5785_
	);
	LUT2 #(
		.INIT('h1)
	) name1739 (
		_w5784_,
		_w5785_,
		_w5786_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w5068_,
		_w5786_,
		_w5787_
	);
	LUT2 #(
		.INIT('h8)
	) name1741 (
		\idma_DTMP_H_reg[9]/P0001 ,
		_w5068_,
		_w5788_
	);
	LUT2 #(
		.INIT('h1)
	) name1742 (
		_w5787_,
		_w5788_,
		_w5789_
	);
	LUT2 #(
		.INIT('h2)
	) name1743 (
		\sice_idr1_reg_DO_reg[6]/P0001 ,
		_w5735_,
		_w5790_
	);
	LUT2 #(
		.INIT('h8)
	) name1744 (
		\bdma_BRdataBUF_reg[18]/P0001 ,
		_w5735_,
		_w5791_
	);
	LUT2 #(
		.INIT('h1)
	) name1745 (
		_w5790_,
		_w5791_,
		_w5792_
	);
	LUT2 #(
		.INIT('h1)
	) name1746 (
		_w5068_,
		_w5792_,
		_w5793_
	);
	LUT2 #(
		.INIT('h8)
	) name1747 (
		\idma_DTMP_H_reg[10]/P0001 ,
		_w5068_,
		_w5794_
	);
	LUT2 #(
		.INIT('h1)
	) name1748 (
		_w5793_,
		_w5794_,
		_w5795_
	);
	LUT2 #(
		.INIT('h2)
	) name1749 (
		\sice_idr1_reg_DO_reg[7]/P0001 ,
		_w5735_,
		_w5796_
	);
	LUT2 #(
		.INIT('h8)
	) name1750 (
		\bdma_BRdataBUF_reg[19]/P0001 ,
		_w5735_,
		_w5797_
	);
	LUT2 #(
		.INIT('h1)
	) name1751 (
		_w5796_,
		_w5797_,
		_w5798_
	);
	LUT2 #(
		.INIT('h1)
	) name1752 (
		_w5068_,
		_w5798_,
		_w5799_
	);
	LUT2 #(
		.INIT('h8)
	) name1753 (
		\idma_DTMP_H_reg[11]/P0001 ,
		_w5068_,
		_w5800_
	);
	LUT2 #(
		.INIT('h1)
	) name1754 (
		_w5799_,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h2)
	) name1755 (
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w5735_,
		_w5802_
	);
	LUT2 #(
		.INIT('h8)
	) name1756 (
		\bdma_BRdataBUF_reg[1]/P0001 ,
		_w5735_,
		_w5803_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w5802_,
		_w5803_,
		_w5804_
	);
	LUT2 #(
		.INIT('h1)
	) name1758 (
		_w5068_,
		_w5804_,
		_w5805_
	);
	LUT2 #(
		.INIT('h8)
	) name1759 (
		\idma_DTMP_L_reg[1]/P0001 ,
		_w5068_,
		_w5806_
	);
	LUT2 #(
		.INIT('h1)
	) name1760 (
		_w5805_,
		_w5806_,
		_w5807_
	);
	LUT2 #(
		.INIT('h2)
	) name1761 (
		\sice_idr1_reg_DO_reg[8]/P0001 ,
		_w5735_,
		_w5808_
	);
	LUT2 #(
		.INIT('h8)
	) name1762 (
		\bdma_BRdataBUF_reg[20]/P0001 ,
		_w5735_,
		_w5809_
	);
	LUT2 #(
		.INIT('h1)
	) name1763 (
		_w5808_,
		_w5809_,
		_w5810_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		_w5068_,
		_w5810_,
		_w5811_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		\idma_DTMP_H_reg[12]/P0001 ,
		_w5068_,
		_w5812_
	);
	LUT2 #(
		.INIT('h1)
	) name1766 (
		_w5811_,
		_w5812_,
		_w5813_
	);
	LUT2 #(
		.INIT('h2)
	) name1767 (
		\sice_idr1_reg_DO_reg[9]/P0001 ,
		_w5735_,
		_w5814_
	);
	LUT2 #(
		.INIT('h8)
	) name1768 (
		\bdma_BRdataBUF_reg[21]/P0001 ,
		_w5735_,
		_w5815_
	);
	LUT2 #(
		.INIT('h1)
	) name1769 (
		_w5814_,
		_w5815_,
		_w5816_
	);
	LUT2 #(
		.INIT('h1)
	) name1770 (
		_w5068_,
		_w5816_,
		_w5817_
	);
	LUT2 #(
		.INIT('h8)
	) name1771 (
		\idma_DTMP_H_reg[13]/P0001 ,
		_w5068_,
		_w5818_
	);
	LUT2 #(
		.INIT('h1)
	) name1772 (
		_w5817_,
		_w5818_,
		_w5819_
	);
	LUT2 #(
		.INIT('h2)
	) name1773 (
		\sice_idr1_reg_DO_reg[10]/P0001 ,
		_w5735_,
		_w5820_
	);
	LUT2 #(
		.INIT('h8)
	) name1774 (
		\bdma_BRdataBUF_reg[22]/P0001 ,
		_w5735_,
		_w5821_
	);
	LUT2 #(
		.INIT('h1)
	) name1775 (
		_w5820_,
		_w5821_,
		_w5822_
	);
	LUT2 #(
		.INIT('h1)
	) name1776 (
		_w5068_,
		_w5822_,
		_w5823_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		\idma_DTMP_H_reg[14]/P0001 ,
		_w5068_,
		_w5824_
	);
	LUT2 #(
		.INIT('h1)
	) name1778 (
		_w5823_,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h2)
	) name1779 (
		\sice_idr1_reg_DO_reg[11]/P0001 ,
		_w5735_,
		_w5826_
	);
	LUT2 #(
		.INIT('h8)
	) name1780 (
		\bdma_BRdataBUF_reg[23]/P0001 ,
		_w5735_,
		_w5827_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w5826_,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h1)
	) name1782 (
		_w5068_,
		_w5828_,
		_w5829_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		\idma_DTMP_H_reg[15]/P0001 ,
		_w5068_,
		_w5830_
	);
	LUT2 #(
		.INIT('h1)
	) name1784 (
		_w5829_,
		_w5830_,
		_w5831_
	);
	LUT2 #(
		.INIT('h2)
	) name1785 (
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w5735_,
		_w5832_
	);
	LUT2 #(
		.INIT('h8)
	) name1786 (
		\bdma_BRdataBUF_reg[2]/P0001 ,
		_w5735_,
		_w5833_
	);
	LUT2 #(
		.INIT('h1)
	) name1787 (
		_w5832_,
		_w5833_,
		_w5834_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w5068_,
		_w5834_,
		_w5835_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		\idma_DTMP_L_reg[2]/P0001 ,
		_w5068_,
		_w5836_
	);
	LUT2 #(
		.INIT('h1)
	) name1790 (
		_w5835_,
		_w5836_,
		_w5837_
	);
	LUT2 #(
		.INIT('h2)
	) name1791 (
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w5735_,
		_w5838_
	);
	LUT2 #(
		.INIT('h8)
	) name1792 (
		\bdma_BRdataBUF_reg[3]/P0001 ,
		_w5735_,
		_w5839_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w5838_,
		_w5839_,
		_w5840_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		_w5068_,
		_w5840_,
		_w5841_
	);
	LUT2 #(
		.INIT('h8)
	) name1795 (
		\idma_DTMP_L_reg[3]/P0001 ,
		_w5068_,
		_w5842_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w5841_,
		_w5842_,
		_w5843_
	);
	LUT2 #(
		.INIT('h2)
	) name1797 (
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w5735_,
		_w5844_
	);
	LUT2 #(
		.INIT('h8)
	) name1798 (
		\bdma_BRdataBUF_reg[4]/P0001 ,
		_w5735_,
		_w5845_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		_w5844_,
		_w5845_,
		_w5846_
	);
	LUT2 #(
		.INIT('h1)
	) name1800 (
		_w5068_,
		_w5846_,
		_w5847_
	);
	LUT2 #(
		.INIT('h8)
	) name1801 (
		\idma_DTMP_L_reg[4]/P0001 ,
		_w5068_,
		_w5848_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		_w5847_,
		_w5848_,
		_w5849_
	);
	LUT2 #(
		.INIT('h2)
	) name1803 (
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w5735_,
		_w5850_
	);
	LUT2 #(
		.INIT('h8)
	) name1804 (
		\bdma_BRdataBUF_reg[5]/P0001 ,
		_w5735_,
		_w5851_
	);
	LUT2 #(
		.INIT('h1)
	) name1805 (
		_w5850_,
		_w5851_,
		_w5852_
	);
	LUT2 #(
		.INIT('h1)
	) name1806 (
		_w5068_,
		_w5852_,
		_w5853_
	);
	LUT2 #(
		.INIT('h8)
	) name1807 (
		\idma_DTMP_L_reg[5]/P0001 ,
		_w5068_,
		_w5854_
	);
	LUT2 #(
		.INIT('h1)
	) name1808 (
		_w5853_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h2)
	) name1809 (
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w5735_,
		_w5856_
	);
	LUT2 #(
		.INIT('h8)
	) name1810 (
		\bdma_BRdataBUF_reg[6]/P0001 ,
		_w5735_,
		_w5857_
	);
	LUT2 #(
		.INIT('h1)
	) name1811 (
		_w5856_,
		_w5857_,
		_w5858_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w5068_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('h8)
	) name1813 (
		\idma_DTMP_L_reg[6]/P0001 ,
		_w5068_,
		_w5860_
	);
	LUT2 #(
		.INIT('h1)
	) name1814 (
		_w5859_,
		_w5860_,
		_w5861_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w5735_,
		_w5862_
	);
	LUT2 #(
		.INIT('h8)
	) name1816 (
		\bdma_BRdataBUF_reg[7]/P0001 ,
		_w5735_,
		_w5863_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w5862_,
		_w5863_,
		_w5864_
	);
	LUT2 #(
		.INIT('h1)
	) name1818 (
		_w5068_,
		_w5864_,
		_w5865_
	);
	LUT2 #(
		.INIT('h8)
	) name1819 (
		\idma_DTMP_L_reg[7]/P0001 ,
		_w5068_,
		_w5866_
	);
	LUT2 #(
		.INIT('h1)
	) name1820 (
		_w5865_,
		_w5866_,
		_w5867_
	);
	LUT2 #(
		.INIT('h2)
	) name1821 (
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w5735_,
		_w5868_
	);
	LUT2 #(
		.INIT('h8)
	) name1822 (
		\bdma_BRdataBUF_reg[8]/P0001 ,
		_w5735_,
		_w5869_
	);
	LUT2 #(
		.INIT('h1)
	) name1823 (
		_w5868_,
		_w5869_,
		_w5870_
	);
	LUT2 #(
		.INIT('h1)
	) name1824 (
		_w5068_,
		_w5870_,
		_w5871_
	);
	LUT2 #(
		.INIT('h8)
	) name1825 (
		\idma_DTMP_H_reg[0]/P0001 ,
		_w5068_,
		_w5872_
	);
	LUT2 #(
		.INIT('h1)
	) name1826 (
		_w5871_,
		_w5872_,
		_w5873_
	);
	LUT2 #(
		.INIT('h2)
	) name1827 (
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w5735_,
		_w5874_
	);
	LUT2 #(
		.INIT('h8)
	) name1828 (
		\bdma_BRdataBUF_reg[9]/P0001 ,
		_w5735_,
		_w5875_
	);
	LUT2 #(
		.INIT('h1)
	) name1829 (
		_w5874_,
		_w5875_,
		_w5876_
	);
	LUT2 #(
		.INIT('h1)
	) name1830 (
		_w5068_,
		_w5876_,
		_w5877_
	);
	LUT2 #(
		.INIT('h8)
	) name1831 (
		\idma_DTMP_H_reg[1]/P0001 ,
		_w5068_,
		_w5878_
	);
	LUT2 #(
		.INIT('h1)
	) name1832 (
		_w5877_,
		_w5878_,
		_w5879_
	);
	LUT2 #(
		.INIT('h4)
	) name1833 (
		\idma_DCTL_reg[14]/NET0131 ,
		_w5068_,
		_w5880_
	);
	LUT2 #(
		.INIT('h1)
	) name1834 (
		PM_bdry_sel_pad,
		\idma_DCTL_reg[12]/NET0131 ,
		_w5881_
	);
	LUT2 #(
		.INIT('h2)
	) name1835 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w5881_,
		_w5882_
	);
	LUT2 #(
		.INIT('h2)
	) name1836 (
		\idma_WRcyc_reg/NET0131 ,
		_w5882_,
		_w5883_
	);
	LUT2 #(
		.INIT('h8)
	) name1837 (
		_w5880_,
		_w5883_,
		_w5884_
	);
	LUT2 #(
		.INIT('h1)
	) name1838 (
		_w5735_,
		_w5884_,
		_w5885_
	);
	LUT2 #(
		.INIT('h2)
	) name1839 (
		_w5679_,
		_w5885_,
		_w5886_
	);
	LUT2 #(
		.INIT('h4)
	) name1840 (
		_w5718_,
		_w5886_,
		_w5887_
	);
	LUT2 #(
		.INIT('h2)
	) name1841 (
		_w4103_,
		_w4117_,
		_w5888_
	);
	LUT2 #(
		.INIT('h2)
	) name1842 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w5679_,
		_w5889_
	);
	LUT2 #(
		.INIT('h8)
	) name1843 (
		_w5888_,
		_w5889_,
		_w5890_
	);
	LUT2 #(
		.INIT('h1)
	) name1844 (
		_w5887_,
		_w5890_,
		_w5891_
	);
	LUT2 #(
		.INIT('h4)
	) name1845 (
		PM_bdry_sel_pad,
		_w5642_,
		_w5892_
	);
	LUT2 #(
		.INIT('h1)
	) name1846 (
		_w5673_,
		_w5892_,
		_w5893_
	);
	LUT2 #(
		.INIT('h1)
	) name1847 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w5066_,
		_w5894_
	);
	LUT2 #(
		.INIT('h2)
	) name1848 (
		_w5068_,
		_w5718_,
		_w5895_
	);
	LUT2 #(
		.INIT('h4)
	) name1849 (
		\bdma_BOVL_reg[3]/NET0131 ,
		_w5066_,
		_w5896_
	);
	LUT2 #(
		.INIT('h1)
	) name1850 (
		_w5894_,
		_w5896_,
		_w5897_
	);
	LUT2 #(
		.INIT('h4)
	) name1851 (
		_w5895_,
		_w5897_,
		_w5898_
	);
	LUT2 #(
		.INIT('h8)
	) name1852 (
		\idma_DOVL_reg[3]/NET0131 ,
		_w5895_,
		_w5899_
	);
	LUT2 #(
		.INIT('h2)
	) name1853 (
		_w5724_,
		_w5898_,
		_w5900_
	);
	LUT2 #(
		.INIT('h4)
	) name1854 (
		_w5899_,
		_w5900_,
		_w5901_
	);
	LUT2 #(
		.INIT('h4)
	) name1855 (
		_w5674_,
		_w5901_,
		_w5902_
	);
	LUT2 #(
		.INIT('h4)
	) name1856 (
		_w5893_,
		_w5902_,
		_w5903_
	);
	LUT2 #(
		.INIT('h2)
	) name1857 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w5066_,
		_w5904_
	);
	LUT2 #(
		.INIT('h8)
	) name1858 (
		\bdma_BOVL_reg[2]/NET0131 ,
		_w5066_,
		_w5905_
	);
	LUT2 #(
		.INIT('h1)
	) name1859 (
		_w5904_,
		_w5905_,
		_w5906_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		_w5895_,
		_w5906_,
		_w5907_
	);
	LUT2 #(
		.INIT('h8)
	) name1861 (
		\idma_DOVL_reg[2]/NET0131 ,
		_w5895_,
		_w5908_
	);
	LUT2 #(
		.INIT('h1)
	) name1862 (
		_w5907_,
		_w5908_,
		_w5909_
	);
	LUT2 #(
		.INIT('h8)
	) name1863 (
		_w5903_,
		_w5909_,
		_w5910_
	);
	LUT2 #(
		.INIT('h2)
	) name1864 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w5066_,
		_w5911_
	);
	LUT2 #(
		.INIT('h8)
	) name1865 (
		\bdma_BOVL_reg[1]/NET0131 ,
		_w5066_,
		_w5912_
	);
	LUT2 #(
		.INIT('h1)
	) name1866 (
		_w5911_,
		_w5912_,
		_w5913_
	);
	LUT2 #(
		.INIT('h1)
	) name1867 (
		_w5895_,
		_w5913_,
		_w5914_
	);
	LUT2 #(
		.INIT('h8)
	) name1868 (
		\idma_DOVL_reg[1]/NET0131 ,
		_w5895_,
		_w5915_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w5914_,
		_w5915_,
		_w5916_
	);
	LUT2 #(
		.INIT('h8)
	) name1870 (
		_w5910_,
		_w5916_,
		_w5917_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w5066_,
		_w5918_
	);
	LUT2 #(
		.INIT('h8)
	) name1872 (
		\bdma_BOVL_reg[0]/NET0131 ,
		_w5066_,
		_w5919_
	);
	LUT2 #(
		.INIT('h1)
	) name1873 (
		_w5918_,
		_w5919_,
		_w5920_
	);
	LUT2 #(
		.INIT('h1)
	) name1874 (
		_w5895_,
		_w5920_,
		_w5921_
	);
	LUT2 #(
		.INIT('h8)
	) name1875 (
		\idma_DOVL_reg[0]/NET0131 ,
		_w5895_,
		_w5922_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		_w5921_,
		_w5922_,
		_w5923_
	);
	LUT2 #(
		.INIT('h8)
	) name1877 (
		_w5917_,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h2)
	) name1878 (
		_w5917_,
		_w5923_,
		_w5925_
	);
	LUT2 #(
		.INIT('h2)
	) name1879 (
		_w5910_,
		_w5916_,
		_w5926_
	);
	LUT2 #(
		.INIT('h8)
	) name1880 (
		_w5923_,
		_w5926_,
		_w5927_
	);
	LUT2 #(
		.INIT('h4)
	) name1881 (
		_w5923_,
		_w5926_,
		_w5928_
	);
	LUT2 #(
		.INIT('h2)
	) name1882 (
		_w5903_,
		_w5909_,
		_w5929_
	);
	LUT2 #(
		.INIT('h8)
	) name1883 (
		_w5916_,
		_w5929_,
		_w5930_
	);
	LUT2 #(
		.INIT('h8)
	) name1884 (
		_w5923_,
		_w5930_,
		_w5931_
	);
	LUT2 #(
		.INIT('h4)
	) name1885 (
		_w5923_,
		_w5930_,
		_w5932_
	);
	LUT2 #(
		.INIT('h4)
	) name1886 (
		_w5916_,
		_w5929_,
		_w5933_
	);
	LUT2 #(
		.INIT('h8)
	) name1887 (
		_w5923_,
		_w5933_,
		_w5934_
	);
	LUT2 #(
		.INIT('h4)
	) name1888 (
		_w5923_,
		_w5933_,
		_w5935_
	);
	LUT2 #(
		.INIT('h1)
	) name1889 (
		_w4055_,
		_w5716_,
		_w5936_
	);
	LUT2 #(
		.INIT('h8)
	) name1890 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w5937_
	);
	LUT2 #(
		.INIT('h8)
	) name1891 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		_w5938_
	);
	LUT2 #(
		.INIT('h8)
	) name1892 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		_w5939_
	);
	LUT2 #(
		.INIT('h8)
	) name1893 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		_w5940_
	);
	LUT2 #(
		.INIT('h8)
	) name1894 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		_w5940_,
		_w5941_
	);
	LUT2 #(
		.INIT('h8)
	) name1895 (
		_w5938_,
		_w5939_,
		_w5942_
	);
	LUT2 #(
		.INIT('h8)
	) name1896 (
		_w5937_,
		_w5942_,
		_w5943_
	);
	LUT2 #(
		.INIT('h8)
	) name1897 (
		_w5941_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h2)
	) name1898 (
		\memc_Dwrite_E_reg/NET0131 ,
		\memc_EXTC_E_reg/NET0131 ,
		_w5945_
	);
	LUT2 #(
		.INIT('h4)
	) name1899 (
		_w5944_,
		_w5945_,
		_w5946_
	);
	LUT2 #(
		.INIT('h4)
	) name1900 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w5946_,
		_w5947_
	);
	LUT2 #(
		.INIT('h1)
	) name1901 (
		_w4099_,
		_w5947_,
		_w5948_
	);
	LUT2 #(
		.INIT('h4)
	) name1902 (
		_w4117_,
		_w5948_,
		_w5949_
	);
	LUT2 #(
		.INIT('h4)
	) name1903 (
		\sice_GO_NX_reg/NET0131 ,
		_w4093_,
		_w5950_
	);
	LUT2 #(
		.INIT('h1)
	) name1904 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w5950_,
		_w5951_
	);
	LUT2 #(
		.INIT('h1)
	) name1905 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_dag_ilm2reg_IL_E_reg[0]/P0001 ,
		_w5952_
	);
	LUT2 #(
		.INIT('h1)
	) name1906 (
		\auctl_R0Sack_reg/NET0131 ,
		\auctl_R1Sack_reg/NET0131 ,
		_w5953_
	);
	LUT2 #(
		.INIT('h1)
	) name1907 (
		\auctl_T0Sack_reg/NET0131 ,
		\auctl_T1Sack_reg/NET0131 ,
		_w5954_
	);
	LUT2 #(
		.INIT('h8)
	) name1908 (
		_w5953_,
		_w5954_,
		_w5955_
	);
	LUT2 #(
		.INIT('h8)
	) name1909 (
		\core_c_dec_Post2_E_reg/P0001 ,
		_w5955_,
		_w5956_
	);
	LUT2 #(
		.INIT('h4)
	) name1910 (
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w5956_,
		_w5957_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		_w5952_,
		_w5957_,
		_w5958_
	);
	LUT2 #(
		.INIT('h1)
	) name1912 (
		\core_c_dec_MTIreg_E_reg[4]/P0001 ,
		_w5958_,
		_w5959_
	);
	LUT2 #(
		.INIT('h2)
	) name1913 (
		_w5951_,
		_w5959_,
		_w5960_
	);
	LUT2 #(
		.INIT('h4)
	) name1914 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w5961_
	);
	LUT2 #(
		.INIT('h1)
	) name1915 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w5955_,
		_w5962_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		_w5961_,
		_w5962_,
		_w5963_
	);
	LUT2 #(
		.INIT('h1)
	) name1917 (
		_w5960_,
		_w5963_,
		_w5964_
	);
	LUT2 #(
		.INIT('h8)
	) name1918 (
		\sport0_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w4050_,
		_w5965_
	);
	LUT2 #(
		.INIT('h8)
	) name1919 (
		_w4049_,
		_w4054_,
		_w5966_
	);
	LUT2 #(
		.INIT('h8)
	) name1920 (
		\sport1_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w5966_,
		_w5967_
	);
	LUT2 #(
		.INIT('h8)
	) name1921 (
		_w4052_,
		_w4053_,
		_w5968_
	);
	LUT2 #(
		.INIT('h8)
	) name1922 (
		\sport1_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w5968_,
		_w5969_
	);
	LUT2 #(
		.INIT('h4)
	) name1923 (
		_w4050_,
		_w4051_,
		_w5970_
	);
	LUT2 #(
		.INIT('h8)
	) name1924 (
		\sport0_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w5970_,
		_w5971_
	);
	LUT2 #(
		.INIT('h1)
	) name1925 (
		_w5965_,
		_w5971_,
		_w5972_
	);
	LUT2 #(
		.INIT('h4)
	) name1926 (
		_w5969_,
		_w5972_,
		_w5973_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		_w5967_,
		_w5973_,
		_w5974_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		\sport0_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w4050_,
		_w5975_
	);
	LUT2 #(
		.INIT('h8)
	) name1929 (
		\sport1_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w5966_,
		_w5976_
	);
	LUT2 #(
		.INIT('h8)
	) name1930 (
		\sport1_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w5968_,
		_w5977_
	);
	LUT2 #(
		.INIT('h8)
	) name1931 (
		\sport0_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w5970_,
		_w5978_
	);
	LUT2 #(
		.INIT('h1)
	) name1932 (
		_w5975_,
		_w5978_,
		_w5979_
	);
	LUT2 #(
		.INIT('h4)
	) name1933 (
		_w5977_,
		_w5979_,
		_w5980_
	);
	LUT2 #(
		.INIT('h4)
	) name1934 (
		_w5976_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h2)
	) name1935 (
		_w5974_,
		_w5981_,
		_w5982_
	);
	LUT2 #(
		.INIT('h8)
	) name1936 (
		\sport0_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w4050_,
		_w5983_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		\sport1_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w5966_,
		_w5984_
	);
	LUT2 #(
		.INIT('h8)
	) name1938 (
		\sport1_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w5968_,
		_w5985_
	);
	LUT2 #(
		.INIT('h8)
	) name1939 (
		\sport0_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w5970_,
		_w5986_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w5983_,
		_w5986_,
		_w5987_
	);
	LUT2 #(
		.INIT('h4)
	) name1941 (
		_w5985_,
		_w5987_,
		_w5988_
	);
	LUT2 #(
		.INIT('h4)
	) name1942 (
		_w5984_,
		_w5988_,
		_w5989_
	);
	LUT2 #(
		.INIT('h8)
	) name1943 (
		_w5982_,
		_w5989_,
		_w5990_
	);
	LUT2 #(
		.INIT('h4)
	) name1944 (
		_w5964_,
		_w5990_,
		_w5991_
	);
	LUT2 #(
		.INIT('h8)
	) name1945 (
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w5956_,
		_w5992_
	);
	LUT2 #(
		.INIT('h4)
	) name1946 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_dag_ilm2reg_IL_E_reg[0]/P0001 ,
		_w5993_
	);
	LUT2 #(
		.INIT('h8)
	) name1947 (
		_w5992_,
		_w5993_,
		_w5994_
	);
	LUT2 #(
		.INIT('h1)
	) name1948 (
		\core_c_dec_MTIreg_E_reg[7]/P0001 ,
		_w5994_,
		_w5995_
	);
	LUT2 #(
		.INIT('h2)
	) name1949 (
		_w5951_,
		_w5995_,
		_w5996_
	);
	LUT2 #(
		.INIT('h2)
	) name1950 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w5955_,
		_w5997_
	);
	LUT2 #(
		.INIT('h8)
	) name1951 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w5998_
	);
	LUT2 #(
		.INIT('h8)
	) name1952 (
		_w5997_,
		_w5998_,
		_w5999_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		_w5996_,
		_w5999_,
		_w6000_
	);
	LUT2 #(
		.INIT('h1)
	) name1954 (
		_w5974_,
		_w5981_,
		_w6001_
	);
	LUT2 #(
		.INIT('h4)
	) name1955 (
		_w5989_,
		_w6001_,
		_w6002_
	);
	LUT2 #(
		.INIT('h4)
	) name1956 (
		_w6000_,
		_w6002_,
		_w6003_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		_w5952_,
		_w5992_,
		_w6004_
	);
	LUT2 #(
		.INIT('h1)
	) name1958 (
		\core_c_dec_MTIreg_E_reg[6]/P0001 ,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h2)
	) name1959 (
		_w5951_,
		_w6005_,
		_w6006_
	);
	LUT2 #(
		.INIT('h8)
	) name1960 (
		_w5961_,
		_w5997_,
		_w6007_
	);
	LUT2 #(
		.INIT('h1)
	) name1961 (
		_w6006_,
		_w6007_,
		_w6008_
	);
	LUT2 #(
		.INIT('h8)
	) name1962 (
		_w5989_,
		_w6001_,
		_w6009_
	);
	LUT2 #(
		.INIT('h4)
	) name1963 (
		_w6008_,
		_w6009_,
		_w6010_
	);
	LUT2 #(
		.INIT('h8)
	) name1964 (
		_w5957_,
		_w5993_,
		_w6011_
	);
	LUT2 #(
		.INIT('h1)
	) name1965 (
		\core_c_dec_MTIreg_E_reg[5]/P0001 ,
		_w6011_,
		_w6012_
	);
	LUT2 #(
		.INIT('h2)
	) name1966 (
		_w5951_,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h8)
	) name1967 (
		_w5962_,
		_w5998_,
		_w6014_
	);
	LUT2 #(
		.INIT('h1)
	) name1968 (
		_w6013_,
		_w6014_,
		_w6015_
	);
	LUT2 #(
		.INIT('h2)
	) name1969 (
		_w5982_,
		_w5989_,
		_w6016_
	);
	LUT2 #(
		.INIT('h4)
	) name1970 (
		_w6015_,
		_w6016_,
		_w6017_
	);
	LUT2 #(
		.INIT('h1)
	) name1971 (
		_w5991_,
		_w6003_,
		_w6018_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		_w6010_,
		_w6017_,
		_w6019_
	);
	LUT2 #(
		.INIT('h8)
	) name1973 (
		_w6018_,
		_w6019_,
		_w6020_
	);
	LUT2 #(
		.INIT('h4)
	) name1974 (
		_w4055_,
		_w6020_,
		_w6021_
	);
	LUT2 #(
		.INIT('h2)
	) name1975 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		_w6022_
	);
	LUT2 #(
		.INIT('h8)
	) name1976 (
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6022_,
		_w6023_
	);
	LUT2 #(
		.INIT('h1)
	) name1977 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w6024_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w6025_
	);
	LUT2 #(
		.INIT('h1)
	) name1979 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6026_
	);
	LUT2 #(
		.INIT('h8)
	) name1980 (
		_w4100_,
		_w6026_,
		_w6027_
	);
	LUT2 #(
		.INIT('h8)
	) name1981 (
		_w6025_,
		_w6027_,
		_w6028_
	);
	LUT2 #(
		.INIT('h8)
	) name1982 (
		_w6024_,
		_w6028_,
		_w6029_
	);
	LUT2 #(
		.INIT('h1)
	) name1983 (
		_w6023_,
		_w6029_,
		_w6030_
	);
	LUT2 #(
		.INIT('h2)
	) name1984 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w6030_,
		_w6031_
	);
	LUT2 #(
		.INIT('h8)
	) name1985 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w6030_,
		_w6032_
	);
	LUT2 #(
		.INIT('h1)
	) name1986 (
		_w6031_,
		_w6032_,
		_w6033_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w6030_,
		_w6034_
	);
	LUT2 #(
		.INIT('h8)
	) name1988 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w6030_,
		_w6035_
	);
	LUT2 #(
		.INIT('h1)
	) name1989 (
		_w6034_,
		_w6035_,
		_w6036_
	);
	LUT2 #(
		.INIT('h8)
	) name1990 (
		_w6033_,
		_w6036_,
		_w6037_
	);
	LUT2 #(
		.INIT('h4)
	) name1991 (
		_w5964_,
		_w6037_,
		_w6038_
	);
	LUT2 #(
		.INIT('h1)
	) name1992 (
		_w6033_,
		_w6036_,
		_w6039_
	);
	LUT2 #(
		.INIT('h4)
	) name1993 (
		_w6000_,
		_w6039_,
		_w6040_
	);
	LUT2 #(
		.INIT('h4)
	) name1994 (
		_w6033_,
		_w6036_,
		_w6041_
	);
	LUT2 #(
		.INIT('h4)
	) name1995 (
		_w6008_,
		_w6041_,
		_w6042_
	);
	LUT2 #(
		.INIT('h2)
	) name1996 (
		_w6033_,
		_w6036_,
		_w6043_
	);
	LUT2 #(
		.INIT('h4)
	) name1997 (
		_w6015_,
		_w6043_,
		_w6044_
	);
	LUT2 #(
		.INIT('h1)
	) name1998 (
		_w6038_,
		_w6040_,
		_w6045_
	);
	LUT2 #(
		.INIT('h1)
	) name1999 (
		_w6042_,
		_w6044_,
		_w6046_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT2 #(
		.INIT('h8)
	) name2001 (
		_w4055_,
		_w6047_,
		_w6048_
	);
	LUT2 #(
		.INIT('h1)
	) name2002 (
		_w6021_,
		_w6048_,
		_w6049_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w6050_
	);
	LUT2 #(
		.INIT('h8)
	) name2004 (
		_w5962_,
		_w6050_,
		_w6051_
	);
	LUT2 #(
		.INIT('h4)
	) name2005 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_Post1_E_reg/P0001 ,
		_w6052_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		_w5955_,
		_w6052_,
		_w6053_
	);
	LUT2 #(
		.INIT('h4)
	) name2007 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w6053_,
		_w6054_
	);
	LUT2 #(
		.INIT('h4)
	) name2008 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w6054_,
		_w6055_
	);
	LUT2 #(
		.INIT('h1)
	) name2009 (
		\core_c_dec_MTIreg_E_reg[0]/P0001 ,
		_w6055_,
		_w6056_
	);
	LUT2 #(
		.INIT('h2)
	) name2010 (
		_w5951_,
		_w6056_,
		_w6057_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		_w6051_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h8)
	) name2012 (
		_w5974_,
		_w5981_,
		_w6059_
	);
	LUT2 #(
		.INIT('h8)
	) name2013 (
		_w5989_,
		_w6059_,
		_w6060_
	);
	LUT2 #(
		.INIT('h4)
	) name2014 (
		_w6058_,
		_w6060_,
		_w6061_
	);
	LUT2 #(
		.INIT('h2)
	) name2015 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w6062_
	);
	LUT2 #(
		.INIT('h8)
	) name2016 (
		_w5962_,
		_w6062_,
		_w6063_
	);
	LUT2 #(
		.INIT('h8)
	) name2017 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w6054_,
		_w6064_
	);
	LUT2 #(
		.INIT('h1)
	) name2018 (
		\core_c_dec_MTIreg_E_reg[1]/P0001 ,
		_w6064_,
		_w6065_
	);
	LUT2 #(
		.INIT('h2)
	) name2019 (
		_w5951_,
		_w6065_,
		_w6066_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w6063_,
		_w6066_,
		_w6067_
	);
	LUT2 #(
		.INIT('h4)
	) name2021 (
		_w5989_,
		_w6059_,
		_w6068_
	);
	LUT2 #(
		.INIT('h4)
	) name2022 (
		_w6067_,
		_w6068_,
		_w6069_
	);
	LUT2 #(
		.INIT('h8)
	) name2023 (
		_w5997_,
		_w6062_,
		_w6070_
	);
	LUT2 #(
		.INIT('h8)
	) name2024 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w6071_
	);
	LUT2 #(
		.INIT('h8)
	) name2025 (
		_w6053_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		\core_c_dec_MTIreg_E_reg[3]/P0001 ,
		_w6072_,
		_w6073_
	);
	LUT2 #(
		.INIT('h2)
	) name2027 (
		_w5951_,
		_w6073_,
		_w6074_
	);
	LUT2 #(
		.INIT('h1)
	) name2028 (
		_w6070_,
		_w6074_,
		_w6075_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		_w5974_,
		_w5981_,
		_w6076_
	);
	LUT2 #(
		.INIT('h4)
	) name2030 (
		_w5989_,
		_w6076_,
		_w6077_
	);
	LUT2 #(
		.INIT('h4)
	) name2031 (
		_w6075_,
		_w6077_,
		_w6078_
	);
	LUT2 #(
		.INIT('h8)
	) name2032 (
		_w5997_,
		_w6050_,
		_w6079_
	);
	LUT2 #(
		.INIT('h4)
	) name2033 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w6080_
	);
	LUT2 #(
		.INIT('h8)
	) name2034 (
		_w6053_,
		_w6080_,
		_w6081_
	);
	LUT2 #(
		.INIT('h1)
	) name2035 (
		\core_c_dec_MTIreg_E_reg[2]/P0001 ,
		_w6081_,
		_w6082_
	);
	LUT2 #(
		.INIT('h2)
	) name2036 (
		_w5951_,
		_w6082_,
		_w6083_
	);
	LUT2 #(
		.INIT('h1)
	) name2037 (
		_w6079_,
		_w6083_,
		_w6084_
	);
	LUT2 #(
		.INIT('h8)
	) name2038 (
		_w5989_,
		_w6076_,
		_w6085_
	);
	LUT2 #(
		.INIT('h4)
	) name2039 (
		_w6084_,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h1)
	) name2040 (
		_w4055_,
		_w6061_,
		_w6087_
	);
	LUT2 #(
		.INIT('h1)
	) name2041 (
		_w6069_,
		_w6078_,
		_w6088_
	);
	LUT2 #(
		.INIT('h4)
	) name2042 (
		_w6086_,
		_w6088_,
		_w6089_
	);
	LUT2 #(
		.INIT('h8)
	) name2043 (
		_w6087_,
		_w6089_,
		_w6090_
	);
	LUT2 #(
		.INIT('h2)
	) name2044 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w6091_
	);
	LUT2 #(
		.INIT('h4)
	) name2045 (
		_w6067_,
		_w6091_,
		_w6092_
	);
	LUT2 #(
		.INIT('h1)
	) name2046 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w6093_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w6058_,
		_w6093_,
		_w6094_
	);
	LUT2 #(
		.INIT('h4)
	) name2048 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w6095_
	);
	LUT2 #(
		.INIT('h4)
	) name2049 (
		_w6084_,
		_w6095_,
		_w6096_
	);
	LUT2 #(
		.INIT('h8)
	) name2050 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w6097_
	);
	LUT2 #(
		.INIT('h4)
	) name2051 (
		_w6075_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h1)
	) name2052 (
		_w6092_,
		_w6094_,
		_w6099_
	);
	LUT2 #(
		.INIT('h1)
	) name2053 (
		_w6096_,
		_w6098_,
		_w6100_
	);
	LUT2 #(
		.INIT('h8)
	) name2054 (
		_w6099_,
		_w6100_,
		_w6101_
	);
	LUT2 #(
		.INIT('h8)
	) name2055 (
		_w4055_,
		_w6101_,
		_w6102_
	);
	LUT2 #(
		.INIT('h1)
	) name2056 (
		_w6090_,
		_w6102_,
		_w6103_
	);
	LUT2 #(
		.INIT('h1)
	) name2057 (
		_w6049_,
		_w6103_,
		_w6104_
	);
	LUT2 #(
		.INIT('h2)
	) name2058 (
		_w5949_,
		_w6104_,
		_w6105_
	);
	LUT2 #(
		.INIT('h4)
	) name2059 (
		\core_c_dec_Post1_E_reg/P0001 ,
		_w5955_,
		_w6106_
	);
	LUT2 #(
		.INIT('h8)
	) name2060 (
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6107_
	);
	LUT2 #(
		.INIT('h2)
	) name2061 (
		_w4101_,
		_w4102_,
		_w6108_
	);
	LUT2 #(
		.INIT('h1)
	) name2062 (
		_w6107_,
		_w6108_,
		_w6109_
	);
	LUT2 #(
		.INIT('h1)
	) name2063 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w6109_,
		_w6110_
	);
	LUT2 #(
		.INIT('h1)
	) name2064 (
		_w6023_,
		_w6110_,
		_w6111_
	);
	LUT2 #(
		.INIT('h2)
	) name2065 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w6111_,
		_w6112_
	);
	LUT2 #(
		.INIT('h8)
	) name2066 (
		_w6106_,
		_w6112_,
		_w6113_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w6109_,
		_w6114_
	);
	LUT2 #(
		.INIT('h2)
	) name2068 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w6115_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w6116_
	);
	LUT2 #(
		.INIT('h2)
	) name2070 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6117_
	);
	LUT2 #(
		.INIT('h8)
	) name2071 (
		_w4100_,
		_w6117_,
		_w6118_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		_w6116_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		_w6115_,
		_w6119_,
		_w6120_
	);
	LUT2 #(
		.INIT('h1)
	) name2074 (
		_w6114_,
		_w6120_,
		_w6121_
	);
	LUT2 #(
		.INIT('h2)
	) name2075 (
		_w6049_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('h2)
	) name2076 (
		_w6111_,
		_w6122_,
		_w6123_
	);
	LUT2 #(
		.INIT('h2)
	) name2077 (
		_w6105_,
		_w6113_,
		_w6124_
	);
	LUT2 #(
		.INIT('h4)
	) name2078 (
		_w6123_,
		_w6124_,
		_w6125_
	);
	LUT2 #(
		.INIT('h1)
	) name2079 (
		_w5936_,
		_w6125_,
		_w6126_
	);
	LUT2 #(
		.INIT('h1)
	) name2080 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w6111_,
		_w6127_
	);
	LUT2 #(
		.INIT('h1)
	) name2081 (
		_w5936_,
		_w6127_,
		_w6128_
	);
	LUT2 #(
		.INIT('h1)
	) name2082 (
		_w6106_,
		_w6128_,
		_w6129_
	);
	LUT2 #(
		.INIT('h8)
	) name2083 (
		_w6103_,
		_w6129_,
		_w6130_
	);
	LUT2 #(
		.INIT('h2)
	) name2084 (
		_w5949_,
		_w6111_,
		_w6131_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		_w6049_,
		_w6131_,
		_w6132_
	);
	LUT2 #(
		.INIT('h4)
	) name2086 (
		_w6103_,
		_w6132_,
		_w6133_
	);
	LUT2 #(
		.INIT('h1)
	) name2087 (
		_w6130_,
		_w6133_,
		_w6134_
	);
	LUT2 #(
		.INIT('h4)
	) name2088 (
		_w6126_,
		_w6134_,
		_w6135_
	);
	LUT2 #(
		.INIT('h8)
	) name2089 (
		\core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 ,
		_w6058_,
		_w6136_
	);
	LUT2 #(
		.INIT('h8)
	) name2090 (
		_w6060_,
		_w6136_,
		_w6137_
	);
	LUT2 #(
		.INIT('h8)
	) name2091 (
		_w6084_,
		_w6085_,
		_w6138_
	);
	LUT2 #(
		.INIT('h8)
	) name2092 (
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w6138_,
		_w6139_
	);
	LUT2 #(
		.INIT('h8)
	) name2093 (
		_w6075_,
		_w6077_,
		_w6140_
	);
	LUT2 #(
		.INIT('h8)
	) name2094 (
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		_w6140_,
		_w6141_
	);
	LUT2 #(
		.INIT('h8)
	) name2095 (
		_w6067_,
		_w6068_,
		_w6142_
	);
	LUT2 #(
		.INIT('h8)
	) name2096 (
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w6142_,
		_w6143_
	);
	LUT2 #(
		.INIT('h1)
	) name2097 (
		_w4055_,
		_w6137_,
		_w6144_
	);
	LUT2 #(
		.INIT('h1)
	) name2098 (
		_w6139_,
		_w6141_,
		_w6145_
	);
	LUT2 #(
		.INIT('h4)
	) name2099 (
		_w6143_,
		_w6145_,
		_w6146_
	);
	LUT2 #(
		.INIT('h8)
	) name2100 (
		_w6144_,
		_w6146_,
		_w6147_
	);
	LUT2 #(
		.INIT('h8)
	) name2101 (
		_w6058_,
		_w6093_,
		_w6148_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		\core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 ,
		_w6148_,
		_w6149_
	);
	LUT2 #(
		.INIT('h8)
	) name2103 (
		_w6075_,
		_w6097_,
		_w6150_
	);
	LUT2 #(
		.INIT('h8)
	) name2104 (
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h8)
	) name2105 (
		_w6084_,
		_w6095_,
		_w6152_
	);
	LUT2 #(
		.INIT('h8)
	) name2106 (
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w6152_,
		_w6153_
	);
	LUT2 #(
		.INIT('h8)
	) name2107 (
		_w6067_,
		_w6091_,
		_w6154_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w6154_,
		_w6155_
	);
	LUT2 #(
		.INIT('h1)
	) name2109 (
		_w6149_,
		_w6151_,
		_w6156_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		_w6153_,
		_w6155_,
		_w6157_
	);
	LUT2 #(
		.INIT('h8)
	) name2111 (
		_w6156_,
		_w6157_,
		_w6158_
	);
	LUT2 #(
		.INIT('h8)
	) name2112 (
		_w4055_,
		_w6158_,
		_w6159_
	);
	LUT2 #(
		.INIT('h1)
	) name2113 (
		_w6147_,
		_w6159_,
		_w6160_
	);
	LUT2 #(
		.INIT('h4)
	) name2114 (
		_w6135_,
		_w6160_,
		_w6161_
	);
	LUT2 #(
		.INIT('h8)
	) name2115 (
		_w5936_,
		_w6104_,
		_w6162_
	);
	LUT2 #(
		.INIT('h8)
	) name2116 (
		_w6103_,
		_w6113_,
		_w6163_
	);
	LUT2 #(
		.INIT('h4)
	) name2117 (
		\core_c_dec_Post2_E_reg/P0001 ,
		_w5955_,
		_w6164_
	);
	LUT2 #(
		.INIT('h4)
	) name2118 (
		_w6121_,
		_w6164_,
		_w6165_
	);
	LUT2 #(
		.INIT('h8)
	) name2119 (
		_w6049_,
		_w6165_,
		_w6166_
	);
	LUT2 #(
		.INIT('h2)
	) name2120 (
		_w6111_,
		_w6166_,
		_w6167_
	);
	LUT2 #(
		.INIT('h2)
	) name2121 (
		_w5949_,
		_w6163_,
		_w6168_
	);
	LUT2 #(
		.INIT('h4)
	) name2122 (
		_w6167_,
		_w6168_,
		_w6169_
	);
	LUT2 #(
		.INIT('h1)
	) name2123 (
		_w5936_,
		_w6169_,
		_w6170_
	);
	LUT2 #(
		.INIT('h4)
	) name2124 (
		_w6131_,
		_w6164_,
		_w6171_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w6103_,
		_w6171_,
		_w6172_
	);
	LUT2 #(
		.INIT('h8)
	) name2126 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w6131_,
		_w6173_
	);
	LUT2 #(
		.INIT('h2)
	) name2127 (
		_w6172_,
		_w6173_,
		_w6174_
	);
	LUT2 #(
		.INIT('h1)
	) name2128 (
		_w6162_,
		_w6174_,
		_w6175_
	);
	LUT2 #(
		.INIT('h4)
	) name2129 (
		_w6170_,
		_w6175_,
		_w6176_
	);
	LUT2 #(
		.INIT('h1)
	) name2130 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		_w6177_
	);
	LUT2 #(
		.INIT('h1)
	) name2131 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w6178_
	);
	LUT2 #(
		.INIT('h4)
	) name2132 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		_w6178_,
		_w6179_
	);
	LUT2 #(
		.INIT('h1)
	) name2133 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w6180_
	);
	LUT2 #(
		.INIT('h4)
	) name2134 (
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w6180_,
		_w6181_
	);
	LUT2 #(
		.INIT('h8)
	) name2135 (
		_w6179_,
		_w6181_,
		_w6182_
	);
	LUT2 #(
		.INIT('h8)
	) name2136 (
		_w6177_,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('h1)
	) name2137 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w6184_
	);
	LUT2 #(
		.INIT('h4)
	) name2138 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		_w6184_,
		_w6185_
	);
	LUT2 #(
		.INIT('h8)
	) name2139 (
		_w6183_,
		_w6185_,
		_w6186_
	);
	LUT2 #(
		.INIT('h1)
	) name2140 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w6187_
	);
	LUT2 #(
		.INIT('h8)
	) name2141 (
		_w6186_,
		_w6187_,
		_w6188_
	);
	LUT2 #(
		.INIT('h2)
	) name2142 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		_w6188_,
		_w6189_
	);
	LUT2 #(
		.INIT('h4)
	) name2143 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		_w6184_,
		_w6190_
	);
	LUT2 #(
		.INIT('h1)
	) name2144 (
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w6191_
	);
	LUT2 #(
		.INIT('h4)
	) name2145 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		_w6179_,
		_w6192_
	);
	LUT2 #(
		.INIT('h4)
	) name2146 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w6192_,
		_w6193_
	);
	LUT2 #(
		.INIT('h8)
	) name2147 (
		_w6191_,
		_w6193_,
		_w6194_
	);
	LUT2 #(
		.INIT('h1)
	) name2148 (
		_w6190_,
		_w6194_,
		_w6195_
	);
	LUT2 #(
		.INIT('h1)
	) name2149 (
		_w6191_,
		_w6193_,
		_w6196_
	);
	LUT2 #(
		.INIT('h1)
	) name2150 (
		_w6179_,
		_w6180_,
		_w6197_
	);
	LUT2 #(
		.INIT('h8)
	) name2151 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w6198_
	);
	LUT2 #(
		.INIT('h8)
	) name2152 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w6199_
	);
	LUT2 #(
		.INIT('h8)
	) name2153 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w6200_
	);
	LUT2 #(
		.INIT('h2)
	) name2154 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		_w6178_,
		_w6201_
	);
	LUT2 #(
		.INIT('h8)
	) name2155 (
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w6202_
	);
	LUT2 #(
		.INIT('h8)
	) name2156 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w6203_
	);
	LUT2 #(
		.INIT('h2)
	) name2157 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		_w6184_,
		_w6204_
	);
	LUT2 #(
		.INIT('h1)
	) name2158 (
		_w6186_,
		_w6187_,
		_w6205_
	);
	LUT2 #(
		.INIT('h8)
	) name2159 (
		_w6183_,
		_w6184_,
		_w6206_
	);
	LUT2 #(
		.INIT('h2)
	) name2160 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		_w6206_,
		_w6207_
	);
	LUT2 #(
		.INIT('h1)
	) name2161 (
		_w6198_,
		_w6199_,
		_w6208_
	);
	LUT2 #(
		.INIT('h1)
	) name2162 (
		_w6200_,
		_w6202_,
		_w6209_
	);
	LUT2 #(
		.INIT('h4)
	) name2163 (
		_w6203_,
		_w6209_,
		_w6210_
	);
	LUT2 #(
		.INIT('h4)
	) name2164 (
		_w6201_,
		_w6208_,
		_w6211_
	);
	LUT2 #(
		.INIT('h4)
	) name2165 (
		_w6204_,
		_w6211_,
		_w6212_
	);
	LUT2 #(
		.INIT('h4)
	) name2166 (
		_w6197_,
		_w6210_,
		_w6213_
	);
	LUT2 #(
		.INIT('h8)
	) name2167 (
		_w6212_,
		_w6213_,
		_w6214_
	);
	LUT2 #(
		.INIT('h4)
	) name2168 (
		_w6196_,
		_w6214_,
		_w6215_
	);
	LUT2 #(
		.INIT('h4)
	) name2169 (
		_w6195_,
		_w6215_,
		_w6216_
	);
	LUT2 #(
		.INIT('h1)
	) name2170 (
		_w6205_,
		_w6207_,
		_w6217_
	);
	LUT2 #(
		.INIT('h8)
	) name2171 (
		_w6216_,
		_w6217_,
		_w6218_
	);
	LUT2 #(
		.INIT('h4)
	) name2172 (
		_w6189_,
		_w6218_,
		_w6219_
	);
	LUT2 #(
		.INIT('h2)
	) name2173 (
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w6219_,
		_w6220_
	);
	LUT2 #(
		.INIT('h1)
	) name2174 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		_w6221_
	);
	LUT2 #(
		.INIT('h4)
	) name2175 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w6221_,
		_w6222_
	);
	LUT2 #(
		.INIT('h4)
	) name2176 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		_w6222_,
		_w6223_
	);
	LUT2 #(
		.INIT('h8)
	) name2177 (
		_w6184_,
		_w6223_,
		_w6224_
	);
	LUT2 #(
		.INIT('h8)
	) name2178 (
		_w6177_,
		_w6224_,
		_w6225_
	);
	LUT2 #(
		.INIT('h8)
	) name2179 (
		_w6219_,
		_w6225_,
		_w6226_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		_w6181_,
		_w6226_,
		_w6227_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		_w6179_,
		_w6227_,
		_w6228_
	);
	LUT2 #(
		.INIT('h1)
	) name2182 (
		_w6220_,
		_w6228_,
		_w6229_
	);
	LUT2 #(
		.INIT('h2)
	) name2183 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		_w6229_,
		_w6230_
	);
	LUT2 #(
		.INIT('h1)
	) name2184 (
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h2)
	) name2185 (
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6232_
	);
	LUT2 #(
		.INIT('h1)
	) name2186 (
		_w6231_,
		_w6232_,
		_w6233_
	);
	LUT2 #(
		.INIT('h2)
	) name2187 (
		_w6183_,
		_w6219_,
		_w6234_
	);
	LUT2 #(
		.INIT('h2)
	) name2188 (
		_w6219_,
		_w6223_,
		_w6235_
	);
	LUT2 #(
		.INIT('h4)
	) name2189 (
		_w6190_,
		_w6219_,
		_w6236_
	);
	LUT2 #(
		.INIT('h1)
	) name2190 (
		_w6234_,
		_w6235_,
		_w6237_
	);
	LUT2 #(
		.INIT('h4)
	) name2191 (
		_w6236_,
		_w6237_,
		_w6238_
	);
	LUT2 #(
		.INIT('h8)
	) name2192 (
		\core_dag_ilm1reg_I_reg[6]/NET0131 ,
		_w6238_,
		_w6239_
	);
	LUT2 #(
		.INIT('h1)
	) name2193 (
		\core_dag_ilm1reg_M_reg[6]/NET0131 ,
		_w6239_,
		_w6240_
	);
	LUT2 #(
		.INIT('h8)
	) name2194 (
		\core_dag_ilm1reg_M_reg[6]/NET0131 ,
		_w6239_,
		_w6241_
	);
	LUT2 #(
		.INIT('h1)
	) name2195 (
		_w6240_,
		_w6241_,
		_w6242_
	);
	LUT2 #(
		.INIT('h1)
	) name2196 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6243_
	);
	LUT2 #(
		.INIT('h8)
	) name2197 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6244_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		_w6243_,
		_w6244_,
		_w6245_
	);
	LUT2 #(
		.INIT('h2)
	) name2199 (
		_w6242_,
		_w6245_,
		_w6246_
	);
	LUT2 #(
		.INIT('h4)
	) name2200 (
		_w6242_,
		_w6245_,
		_w6247_
	);
	LUT2 #(
		.INIT('h1)
	) name2201 (
		_w6246_,
		_w6247_,
		_w6248_
	);
	LUT2 #(
		.INIT('h2)
	) name2202 (
		_w6219_,
		_w6224_,
		_w6249_
	);
	LUT2 #(
		.INIT('h4)
	) name2203 (
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w6234_,
		_w6250_
	);
	LUT2 #(
		.INIT('h1)
	) name2204 (
		_w6249_,
		_w6250_,
		_w6251_
	);
	LUT2 #(
		.INIT('h8)
	) name2205 (
		\core_dag_ilm1reg_I_reg[5]/NET0131 ,
		_w6251_,
		_w6252_
	);
	LUT2 #(
		.INIT('h8)
	) name2206 (
		\core_dag_ilm1reg_M_reg[5]/NET0131 ,
		_w6252_,
		_w6253_
	);
	LUT2 #(
		.INIT('h1)
	) name2207 (
		\core_dag_ilm1reg_M_reg[5]/NET0131 ,
		_w6252_,
		_w6254_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6255_
	);
	LUT2 #(
		.INIT('h8)
	) name2209 (
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6256_
	);
	LUT2 #(
		.INIT('h1)
	) name2210 (
		_w6255_,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h1)
	) name2211 (
		_w6254_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h1)
	) name2212 (
		_w6253_,
		_w6258_,
		_w6259_
	);
	LUT2 #(
		.INIT('h4)
	) name2213 (
		_w6248_,
		_w6259_,
		_w6260_
	);
	LUT2 #(
		.INIT('h1)
	) name2214 (
		_w6194_,
		_w6219_,
		_w6261_
	);
	LUT2 #(
		.INIT('h1)
	) name2215 (
		_w6226_,
		_w6261_,
		_w6262_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		_w6262_,
		_w6263_
	);
	LUT2 #(
		.INIT('h1)
	) name2217 (
		\core_dag_ilm1reg_M_reg[7]/NET0131 ,
		_w6263_,
		_w6264_
	);
	LUT2 #(
		.INIT('h8)
	) name2218 (
		\core_dag_ilm1reg_M_reg[7]/NET0131 ,
		_w6263_,
		_w6265_
	);
	LUT2 #(
		.INIT('h1)
	) name2219 (
		_w6264_,
		_w6265_,
		_w6266_
	);
	LUT2 #(
		.INIT('h1)
	) name2220 (
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6267_
	);
	LUT2 #(
		.INIT('h8)
	) name2221 (
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6268_
	);
	LUT2 #(
		.INIT('h1)
	) name2222 (
		_w6267_,
		_w6268_,
		_w6269_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		_w6266_,
		_w6269_,
		_w6270_
	);
	LUT2 #(
		.INIT('h4)
	) name2224 (
		_w6266_,
		_w6269_,
		_w6271_
	);
	LUT2 #(
		.INIT('h1)
	) name2225 (
		_w6270_,
		_w6271_,
		_w6272_
	);
	LUT2 #(
		.INIT('h1)
	) name2226 (
		_w6240_,
		_w6245_,
		_w6273_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		_w6241_,
		_w6273_,
		_w6274_
	);
	LUT2 #(
		.INIT('h4)
	) name2228 (
		_w6272_,
		_w6274_,
		_w6275_
	);
	LUT2 #(
		.INIT('h1)
	) name2229 (
		_w6260_,
		_w6275_,
		_w6276_
	);
	LUT2 #(
		.INIT('h4)
	) name2230 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		_w6223_,
		_w6277_
	);
	LUT2 #(
		.INIT('h2)
	) name2231 (
		_w6219_,
		_w6277_,
		_w6278_
	);
	LUT2 #(
		.INIT('h8)
	) name2232 (
		_w6184_,
		_w6234_,
		_w6279_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w6278_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h8)
	) name2234 (
		\core_dag_ilm1reg_I_reg[4]/NET0131 ,
		_w6280_,
		_w6281_
	);
	LUT2 #(
		.INIT('h8)
	) name2235 (
		\core_dag_ilm1reg_M_reg[4]/NET0131 ,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h1)
	) name2236 (
		\core_dag_ilm1reg_M_reg[4]/NET0131 ,
		_w6281_,
		_w6283_
	);
	LUT2 #(
		.INIT('h1)
	) name2237 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6284_
	);
	LUT2 #(
		.INIT('h8)
	) name2238 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6285_
	);
	LUT2 #(
		.INIT('h1)
	) name2239 (
		_w6284_,
		_w6285_,
		_w6286_
	);
	LUT2 #(
		.INIT('h1)
	) name2240 (
		_w6283_,
		_w6286_,
		_w6287_
	);
	LUT2 #(
		.INIT('h1)
	) name2241 (
		_w6282_,
		_w6287_,
		_w6288_
	);
	LUT2 #(
		.INIT('h1)
	) name2242 (
		_w6253_,
		_w6254_,
		_w6289_
	);
	LUT2 #(
		.INIT('h2)
	) name2243 (
		_w6257_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h4)
	) name2244 (
		_w6257_,
		_w6289_,
		_w6291_
	);
	LUT2 #(
		.INIT('h1)
	) name2245 (
		_w6290_,
		_w6291_,
		_w6292_
	);
	LUT2 #(
		.INIT('h2)
	) name2246 (
		_w6288_,
		_w6292_,
		_w6293_
	);
	LUT2 #(
		.INIT('h2)
	) name2247 (
		_w6186_,
		_w6219_,
		_w6294_
	);
	LUT2 #(
		.INIT('h1)
	) name2248 (
		_w6235_,
		_w6294_,
		_w6295_
	);
	LUT2 #(
		.INIT('h8)
	) name2249 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		_w6295_,
		_w6296_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		\core_dag_ilm1reg_M_reg[3]/NET0131 ,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		\core_dag_ilm1reg_M_reg[3]/NET0131 ,
		_w6296_,
		_w6298_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6299_
	);
	LUT2 #(
		.INIT('h8)
	) name2253 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6300_
	);
	LUT2 #(
		.INIT('h1)
	) name2254 (
		_w6299_,
		_w6300_,
		_w6301_
	);
	LUT2 #(
		.INIT('h1)
	) name2255 (
		_w6298_,
		_w6301_,
		_w6302_
	);
	LUT2 #(
		.INIT('h1)
	) name2256 (
		_w6297_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h1)
	) name2257 (
		_w6282_,
		_w6283_,
		_w6304_
	);
	LUT2 #(
		.INIT('h2)
	) name2258 (
		_w6286_,
		_w6304_,
		_w6305_
	);
	LUT2 #(
		.INIT('h4)
	) name2259 (
		_w6286_,
		_w6304_,
		_w6306_
	);
	LUT2 #(
		.INIT('h1)
	) name2260 (
		_w6305_,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h2)
	) name2261 (
		_w6303_,
		_w6307_,
		_w6308_
	);
	LUT2 #(
		.INIT('h1)
	) name2262 (
		_w6293_,
		_w6308_,
		_w6309_
	);
	LUT2 #(
		.INIT('h1)
	) name2263 (
		_w6297_,
		_w6298_,
		_w6310_
	);
	LUT2 #(
		.INIT('h4)
	) name2264 (
		_w6301_,
		_w6310_,
		_w6311_
	);
	LUT2 #(
		.INIT('h2)
	) name2265 (
		_w6301_,
		_w6310_,
		_w6312_
	);
	LUT2 #(
		.INIT('h1)
	) name2266 (
		_w6311_,
		_w6312_,
		_w6313_
	);
	LUT2 #(
		.INIT('h2)
	) name2267 (
		_w6219_,
		_w6222_,
		_w6314_
	);
	LUT2 #(
		.INIT('h4)
	) name2268 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w6186_,
		_w6315_
	);
	LUT2 #(
		.INIT('h4)
	) name2269 (
		_w6219_,
		_w6315_,
		_w6316_
	);
	LUT2 #(
		.INIT('h1)
	) name2270 (
		_w6314_,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h8)
	) name2271 (
		\core_dag_ilm1reg_I_reg[2]/NET0131 ,
		_w6317_,
		_w6318_
	);
	LUT2 #(
		.INIT('h8)
	) name2272 (
		\core_dag_ilm1reg_M_reg[2]/NET0131 ,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		\core_dag_ilm1reg_M_reg[2]/NET0131 ,
		_w6318_,
		_w6320_
	);
	LUT2 #(
		.INIT('h1)
	) name2274 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6321_
	);
	LUT2 #(
		.INIT('h8)
	) name2275 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6322_
	);
	LUT2 #(
		.INIT('h1)
	) name2276 (
		_w6321_,
		_w6322_,
		_w6323_
	);
	LUT2 #(
		.INIT('h1)
	) name2277 (
		_w6320_,
		_w6323_,
		_w6324_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		_w6319_,
		_w6324_,
		_w6325_
	);
	LUT2 #(
		.INIT('h2)
	) name2279 (
		_w6313_,
		_w6325_,
		_w6326_
	);
	LUT2 #(
		.INIT('h4)
	) name2280 (
		_w6313_,
		_w6325_,
		_w6327_
	);
	LUT2 #(
		.INIT('h2)
	) name2281 (
		_w6188_,
		_w6218_,
		_w6328_
	);
	LUT2 #(
		.INIT('h2)
	) name2282 (
		_w6219_,
		_w6221_,
		_w6329_
	);
	LUT2 #(
		.INIT('h2)
	) name2283 (
		\core_dag_ilm1reg_I_reg[1]/NET0131 ,
		_w6328_,
		_w6330_
	);
	LUT2 #(
		.INIT('h4)
	) name2284 (
		_w6329_,
		_w6330_,
		_w6331_
	);
	LUT2 #(
		.INIT('h8)
	) name2285 (
		\core_dag_ilm1reg_M_reg[1]/NET0131 ,
		_w6331_,
		_w6332_
	);
	LUT2 #(
		.INIT('h1)
	) name2286 (
		\core_dag_ilm1reg_M_reg[1]/NET0131 ,
		_w6331_,
		_w6333_
	);
	LUT2 #(
		.INIT('h1)
	) name2287 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6334_
	);
	LUT2 #(
		.INIT('h8)
	) name2288 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6335_
	);
	LUT2 #(
		.INIT('h1)
	) name2289 (
		_w6334_,
		_w6335_,
		_w6336_
	);
	LUT2 #(
		.INIT('h1)
	) name2290 (
		_w6333_,
		_w6336_,
		_w6337_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w6332_,
		_w6337_,
		_w6338_
	);
	LUT2 #(
		.INIT('h1)
	) name2292 (
		_w6319_,
		_w6320_,
		_w6339_
	);
	LUT2 #(
		.INIT('h2)
	) name2293 (
		_w6323_,
		_w6339_,
		_w6340_
	);
	LUT2 #(
		.INIT('h4)
	) name2294 (
		_w6323_,
		_w6339_,
		_w6341_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w6340_,
		_w6341_,
		_w6342_
	);
	LUT2 #(
		.INIT('h4)
	) name2296 (
		_w6338_,
		_w6342_,
		_w6343_
	);
	LUT2 #(
		.INIT('h2)
	) name2297 (
		_w6338_,
		_w6342_,
		_w6344_
	);
	LUT2 #(
		.INIT('h8)
	) name2298 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		_w6219_,
		_w6345_
	);
	LUT2 #(
		.INIT('h8)
	) name2299 (
		_w6221_,
		_w6316_,
		_w6346_
	);
	LUT2 #(
		.INIT('h2)
	) name2300 (
		\core_dag_ilm1reg_I_reg[0]/NET0131 ,
		_w6345_,
		_w6347_
	);
	LUT2 #(
		.INIT('h4)
	) name2301 (
		_w6346_,
		_w6347_,
		_w6348_
	);
	LUT2 #(
		.INIT('h1)
	) name2302 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w6348_,
		_w6349_
	);
	LUT2 #(
		.INIT('h8)
	) name2303 (
		\core_dag_ilm1reg_M_reg[0]/NET0131 ,
		_w6348_,
		_w6350_
	);
	LUT2 #(
		.INIT('h1)
	) name2304 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6351_
	);
	LUT2 #(
		.INIT('h8)
	) name2305 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6352_
	);
	LUT2 #(
		.INIT('h1)
	) name2306 (
		_w6351_,
		_w6352_,
		_w6353_
	);
	LUT2 #(
		.INIT('h4)
	) name2307 (
		_w6350_,
		_w6353_,
		_w6354_
	);
	LUT2 #(
		.INIT('h1)
	) name2308 (
		_w6349_,
		_w6354_,
		_w6355_
	);
	LUT2 #(
		.INIT('h1)
	) name2309 (
		_w6332_,
		_w6333_,
		_w6356_
	);
	LUT2 #(
		.INIT('h2)
	) name2310 (
		_w6336_,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h4)
	) name2311 (
		_w6336_,
		_w6356_,
		_w6358_
	);
	LUT2 #(
		.INIT('h1)
	) name2312 (
		_w6357_,
		_w6358_,
		_w6359_
	);
	LUT2 #(
		.INIT('h1)
	) name2313 (
		_w6355_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h8)
	) name2314 (
		_w6355_,
		_w6359_,
		_w6361_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w6349_,
		_w6350_,
		_w6362_
	);
	LUT2 #(
		.INIT('h4)
	) name2316 (
		_w6353_,
		_w6362_,
		_w6363_
	);
	LUT2 #(
		.INIT('h2)
	) name2317 (
		_w6353_,
		_w6362_,
		_w6364_
	);
	LUT2 #(
		.INIT('h1)
	) name2318 (
		_w6363_,
		_w6364_,
		_w6365_
	);
	LUT2 #(
		.INIT('h4)
	) name2319 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6365_,
		_w6366_
	);
	LUT2 #(
		.INIT('h1)
	) name2320 (
		_w6361_,
		_w6366_,
		_w6367_
	);
	LUT2 #(
		.INIT('h1)
	) name2321 (
		_w6360_,
		_w6367_,
		_w6368_
	);
	LUT2 #(
		.INIT('h4)
	) name2322 (
		_w6344_,
		_w6368_,
		_w6369_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		_w6343_,
		_w6369_,
		_w6370_
	);
	LUT2 #(
		.INIT('h1)
	) name2324 (
		_w6327_,
		_w6370_,
		_w6371_
	);
	LUT2 #(
		.INIT('h1)
	) name2325 (
		_w6326_,
		_w6371_,
		_w6372_
	);
	LUT2 #(
		.INIT('h8)
	) name2326 (
		_w6276_,
		_w6309_,
		_w6373_
	);
	LUT2 #(
		.INIT('h4)
	) name2327 (
		_w6372_,
		_w6373_,
		_w6374_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		_w6248_,
		_w6259_,
		_w6375_
	);
	LUT2 #(
		.INIT('h4)
	) name2329 (
		_w6275_,
		_w6375_,
		_w6376_
	);
	LUT2 #(
		.INIT('h4)
	) name2330 (
		_w6288_,
		_w6292_,
		_w6377_
	);
	LUT2 #(
		.INIT('h4)
	) name2331 (
		_w6303_,
		_w6307_,
		_w6378_
	);
	LUT2 #(
		.INIT('h4)
	) name2332 (
		_w6293_,
		_w6378_,
		_w6379_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w6377_,
		_w6379_,
		_w6380_
	);
	LUT2 #(
		.INIT('h2)
	) name2334 (
		_w6276_,
		_w6380_,
		_w6381_
	);
	LUT2 #(
		.INIT('h2)
	) name2335 (
		_w6272_,
		_w6274_,
		_w6382_
	);
	LUT2 #(
		.INIT('h1)
	) name2336 (
		_w6376_,
		_w6382_,
		_w6383_
	);
	LUT2 #(
		.INIT('h4)
	) name2337 (
		_w6381_,
		_w6383_,
		_w6384_
	);
	LUT2 #(
		.INIT('h4)
	) name2338 (
		_w6374_,
		_w6384_,
		_w6385_
	);
	LUT2 #(
		.INIT('h4)
	) name2339 (
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w6226_,
		_w6386_
	);
	LUT2 #(
		.INIT('h4)
	) name2340 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h1)
	) name2341 (
		_w6193_,
		_w6219_,
		_w6388_
	);
	LUT2 #(
		.INIT('h1)
	) name2342 (
		_w6387_,
		_w6388_,
		_w6389_
	);
	LUT2 #(
		.INIT('h2)
	) name2343 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		_w6389_,
		_w6390_
	);
	LUT2 #(
		.INIT('h1)
	) name2344 (
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w6390_,
		_w6391_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w6390_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name2346 (
		_w6391_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h1)
	) name2347 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6394_
	);
	LUT2 #(
		.INIT('h8)
	) name2348 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6395_
	);
	LUT2 #(
		.INIT('h1)
	) name2349 (
		_w6394_,
		_w6395_,
		_w6396_
	);
	LUT2 #(
		.INIT('h2)
	) name2350 (
		_w6393_,
		_w6396_,
		_w6397_
	);
	LUT2 #(
		.INIT('h4)
	) name2351 (
		_w6393_,
		_w6396_,
		_w6398_
	);
	LUT2 #(
		.INIT('h1)
	) name2352 (
		_w6397_,
		_w6398_,
		_w6399_
	);
	LUT2 #(
		.INIT('h1)
	) name2353 (
		_w6182_,
		_w6219_,
		_w6400_
	);
	LUT2 #(
		.INIT('h1)
	) name2354 (
		_w6386_,
		_w6400_,
		_w6401_
	);
	LUT2 #(
		.INIT('h2)
	) name2355 (
		\core_dag_ilm1reg_I_reg[8]/NET0131 ,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w6402_,
		_w6403_
	);
	LUT2 #(
		.INIT('h1)
	) name2357 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w6402_,
		_w6404_
	);
	LUT2 #(
		.INIT('h1)
	) name2358 (
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6405_
	);
	LUT2 #(
		.INIT('h8)
	) name2359 (
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6406_
	);
	LUT2 #(
		.INIT('h1)
	) name2360 (
		_w6405_,
		_w6406_,
		_w6407_
	);
	LUT2 #(
		.INIT('h1)
	) name2361 (
		_w6404_,
		_w6407_,
		_w6408_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w6403_,
		_w6408_,
		_w6409_
	);
	LUT2 #(
		.INIT('h4)
	) name2363 (
		_w6399_,
		_w6409_,
		_w6410_
	);
	LUT2 #(
		.INIT('h1)
	) name2364 (
		_w6264_,
		_w6269_,
		_w6411_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		_w6265_,
		_w6411_,
		_w6412_
	);
	LUT2 #(
		.INIT('h1)
	) name2366 (
		_w6403_,
		_w6404_,
		_w6413_
	);
	LUT2 #(
		.INIT('h2)
	) name2367 (
		_w6407_,
		_w6413_,
		_w6414_
	);
	LUT2 #(
		.INIT('h4)
	) name2368 (
		_w6407_,
		_w6413_,
		_w6415_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		_w6414_,
		_w6415_,
		_w6416_
	);
	LUT2 #(
		.INIT('h2)
	) name2370 (
		_w6412_,
		_w6416_,
		_w6417_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w6410_,
		_w6417_,
		_w6418_
	);
	LUT2 #(
		.INIT('h4)
	) name2372 (
		_w6385_,
		_w6418_,
		_w6419_
	);
	LUT2 #(
		.INIT('h1)
	) name2373 (
		_w6391_,
		_w6396_,
		_w6420_
	);
	LUT2 #(
		.INIT('h1)
	) name2374 (
		_w6392_,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('h1)
	) name2375 (
		_w6192_,
		_w6219_,
		_w6422_
	);
	LUT2 #(
		.INIT('h1)
	) name2376 (
		_w6227_,
		_w6422_,
		_w6423_
	);
	LUT2 #(
		.INIT('h2)
	) name2377 (
		\core_dag_ilm1reg_I_reg[10]/NET0131 ,
		_w6423_,
		_w6424_
	);
	LUT2 #(
		.INIT('h1)
	) name2378 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w6424_,
		_w6425_
	);
	LUT2 #(
		.INIT('h8)
	) name2379 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w6424_,
		_w6426_
	);
	LUT2 #(
		.INIT('h1)
	) name2380 (
		_w6425_,
		_w6426_,
		_w6427_
	);
	LUT2 #(
		.INIT('h1)
	) name2381 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6428_
	);
	LUT2 #(
		.INIT('h8)
	) name2382 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6429_
	);
	LUT2 #(
		.INIT('h1)
	) name2383 (
		_w6428_,
		_w6429_,
		_w6430_
	);
	LUT2 #(
		.INIT('h2)
	) name2384 (
		_w6427_,
		_w6430_,
		_w6431_
	);
	LUT2 #(
		.INIT('h4)
	) name2385 (
		_w6427_,
		_w6430_,
		_w6432_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		_w6431_,
		_w6432_,
		_w6433_
	);
	LUT2 #(
		.INIT('h2)
	) name2387 (
		_w6421_,
		_w6433_,
		_w6434_
	);
	LUT2 #(
		.INIT('h1)
	) name2388 (
		_w6425_,
		_w6430_,
		_w6435_
	);
	LUT2 #(
		.INIT('h1)
	) name2389 (
		_w6426_,
		_w6435_,
		_w6436_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		_w6181_,
		_w6437_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		_w6225_,
		_w6437_,
		_w6438_
	);
	LUT2 #(
		.INIT('h2)
	) name2392 (
		_w6219_,
		_w6438_,
		_w6439_
	);
	LUT2 #(
		.INIT('h2)
	) name2393 (
		_w6178_,
		_w6219_,
		_w6440_
	);
	LUT2 #(
		.INIT('h4)
	) name2394 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		_w6440_,
		_w6441_
	);
	LUT2 #(
		.INIT('h1)
	) name2395 (
		_w6439_,
		_w6441_,
		_w6442_
	);
	LUT2 #(
		.INIT('h8)
	) name2396 (
		\core_dag_ilm1reg_I_reg[11]/NET0131 ,
		_w6442_,
		_w6443_
	);
	LUT2 #(
		.INIT('h8)
	) name2397 (
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w6443_,
		_w6444_
	);
	LUT2 #(
		.INIT('h1)
	) name2398 (
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w6443_,
		_w6445_
	);
	LUT2 #(
		.INIT('h1)
	) name2399 (
		_w6444_,
		_w6445_,
		_w6446_
	);
	LUT2 #(
		.INIT('h1)
	) name2400 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6447_
	);
	LUT2 #(
		.INIT('h8)
	) name2401 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6448_
	);
	LUT2 #(
		.INIT('h1)
	) name2402 (
		_w6447_,
		_w6448_,
		_w6449_
	);
	LUT2 #(
		.INIT('h2)
	) name2403 (
		_w6446_,
		_w6449_,
		_w6450_
	);
	LUT2 #(
		.INIT('h4)
	) name2404 (
		_w6446_,
		_w6449_,
		_w6451_
	);
	LUT2 #(
		.INIT('h1)
	) name2405 (
		_w6450_,
		_w6451_,
		_w6452_
	);
	LUT2 #(
		.INIT('h2)
	) name2406 (
		_w6436_,
		_w6452_,
		_w6453_
	);
	LUT2 #(
		.INIT('h1)
	) name2407 (
		_w6434_,
		_w6453_,
		_w6454_
	);
	LUT2 #(
		.INIT('h8)
	) name2408 (
		_w6419_,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('h4)
	) name2409 (
		_w6436_,
		_w6452_,
		_w6456_
	);
	LUT2 #(
		.INIT('h4)
	) name2410 (
		_w6421_,
		_w6433_,
		_w6457_
	);
	LUT2 #(
		.INIT('h2)
	) name2411 (
		_w6399_,
		_w6409_,
		_w6458_
	);
	LUT2 #(
		.INIT('h4)
	) name2412 (
		_w6412_,
		_w6416_,
		_w6459_
	);
	LUT2 #(
		.INIT('h4)
	) name2413 (
		_w6410_,
		_w6459_,
		_w6460_
	);
	LUT2 #(
		.INIT('h1)
	) name2414 (
		_w6458_,
		_w6460_,
		_w6461_
	);
	LUT2 #(
		.INIT('h4)
	) name2415 (
		_w6457_,
		_w6461_,
		_w6462_
	);
	LUT2 #(
		.INIT('h2)
	) name2416 (
		_w6454_,
		_w6462_,
		_w6463_
	);
	LUT2 #(
		.INIT('h1)
	) name2417 (
		_w6456_,
		_w6463_,
		_w6464_
	);
	LUT2 #(
		.INIT('h4)
	) name2418 (
		_w6455_,
		_w6464_,
		_w6465_
	);
	LUT2 #(
		.INIT('h8)
	) name2419 (
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w6230_,
		_w6466_
	);
	LUT2 #(
		.INIT('h1)
	) name2420 (
		_w6231_,
		_w6466_,
		_w6467_
	);
	LUT2 #(
		.INIT('h8)
	) name2421 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		_w6219_,
		_w6468_
	);
	LUT2 #(
		.INIT('h1)
	) name2422 (
		_w6439_,
		_w6440_,
		_w6469_
	);
	LUT2 #(
		.INIT('h4)
	) name2423 (
		_w6468_,
		_w6469_,
		_w6470_
	);
	LUT2 #(
		.INIT('h8)
	) name2424 (
		\core_dag_ilm1reg_I_reg[12]/NET0131 ,
		_w6470_,
		_w6471_
	);
	LUT2 #(
		.INIT('h1)
	) name2425 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w6471_,
		_w6472_
	);
	LUT2 #(
		.INIT('h8)
	) name2426 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w6471_,
		_w6473_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6474_
	);
	LUT2 #(
		.INIT('h8)
	) name2428 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6475_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w6474_,
		_w6475_,
		_w6476_
	);
	LUT2 #(
		.INIT('h4)
	) name2430 (
		_w6473_,
		_w6476_,
		_w6477_
	);
	LUT2 #(
		.INIT('h1)
	) name2431 (
		_w6472_,
		_w6477_,
		_w6478_
	);
	LUT2 #(
		.INIT('h2)
	) name2432 (
		_w6467_,
		_w6478_,
		_w6479_
	);
	LUT2 #(
		.INIT('h1)
	) name2433 (
		_w6445_,
		_w6449_,
		_w6480_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w6444_,
		_w6480_,
		_w6481_
	);
	LUT2 #(
		.INIT('h1)
	) name2435 (
		_w6472_,
		_w6473_,
		_w6482_
	);
	LUT2 #(
		.INIT('h4)
	) name2436 (
		_w6476_,
		_w6482_,
		_w6483_
	);
	LUT2 #(
		.INIT('h2)
	) name2437 (
		_w6476_,
		_w6482_,
		_w6484_
	);
	LUT2 #(
		.INIT('h1)
	) name2438 (
		_w6483_,
		_w6484_,
		_w6485_
	);
	LUT2 #(
		.INIT('h2)
	) name2439 (
		_w6481_,
		_w6485_,
		_w6486_
	);
	LUT2 #(
		.INIT('h1)
	) name2440 (
		_w6479_,
		_w6486_,
		_w6487_
	);
	LUT2 #(
		.INIT('h4)
	) name2441 (
		_w6465_,
		_w6487_,
		_w6488_
	);
	LUT2 #(
		.INIT('h4)
	) name2442 (
		_w6467_,
		_w6478_,
		_w6489_
	);
	LUT2 #(
		.INIT('h4)
	) name2443 (
		_w6481_,
		_w6485_,
		_w6490_
	);
	LUT2 #(
		.INIT('h4)
	) name2444 (
		_w6479_,
		_w6490_,
		_w6491_
	);
	LUT2 #(
		.INIT('h1)
	) name2445 (
		_w6489_,
		_w6491_,
		_w6492_
	);
	LUT2 #(
		.INIT('h4)
	) name2446 (
		_w6488_,
		_w6492_,
		_w6493_
	);
	LUT2 #(
		.INIT('h4)
	) name2447 (
		_w6233_,
		_w6493_,
		_w6494_
	);
	LUT2 #(
		.INIT('h2)
	) name2448 (
		_w6233_,
		_w6493_,
		_w6495_
	);
	LUT2 #(
		.INIT('h1)
	) name2449 (
		_w6494_,
		_w6495_,
		_w6496_
	);
	LUT2 #(
		.INIT('h2)
	) name2450 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6230_,
		_w6497_
	);
	LUT2 #(
		.INIT('h4)
	) name2451 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6230_,
		_w6498_
	);
	LUT2 #(
		.INIT('h1)
	) name2452 (
		_w6497_,
		_w6498_,
		_w6499_
	);
	LUT2 #(
		.INIT('h1)
	) name2453 (
		_w6332_,
		_w6350_,
		_w6500_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		_w6333_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h1)
	) name2455 (
		_w6319_,
		_w6501_,
		_w6502_
	);
	LUT2 #(
		.INIT('h1)
	) name2456 (
		_w6320_,
		_w6502_,
		_w6503_
	);
	LUT2 #(
		.INIT('h1)
	) name2457 (
		_w6297_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h1)
	) name2458 (
		_w6298_,
		_w6504_,
		_w6505_
	);
	LUT2 #(
		.INIT('h1)
	) name2459 (
		_w6254_,
		_w6283_,
		_w6506_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		_w6505_,
		_w6506_,
		_w6507_
	);
	LUT2 #(
		.INIT('h4)
	) name2461 (
		_w6254_,
		_w6282_,
		_w6508_
	);
	LUT2 #(
		.INIT('h1)
	) name2462 (
		_w6253_,
		_w6508_,
		_w6509_
	);
	LUT2 #(
		.INIT('h4)
	) name2463 (
		_w6507_,
		_w6509_,
		_w6510_
	);
	LUT2 #(
		.INIT('h1)
	) name2464 (
		_w6240_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('h1)
	) name2465 (
		_w6241_,
		_w6265_,
		_w6512_
	);
	LUT2 #(
		.INIT('h4)
	) name2466 (
		_w6511_,
		_w6512_,
		_w6513_
	);
	LUT2 #(
		.INIT('h1)
	) name2467 (
		_w6264_,
		_w6513_,
		_w6514_
	);
	LUT2 #(
		.INIT('h1)
	) name2468 (
		_w6391_,
		_w6404_,
		_w6515_
	);
	LUT2 #(
		.INIT('h8)
	) name2469 (
		_w6514_,
		_w6515_,
		_w6516_
	);
	LUT2 #(
		.INIT('h1)
	) name2470 (
		_w6425_,
		_w6445_,
		_w6517_
	);
	LUT2 #(
		.INIT('h8)
	) name2471 (
		_w6516_,
		_w6517_,
		_w6518_
	);
	LUT2 #(
		.INIT('h2)
	) name2472 (
		_w6426_,
		_w6445_,
		_w6519_
	);
	LUT2 #(
		.INIT('h1)
	) name2473 (
		_w6392_,
		_w6403_,
		_w6520_
	);
	LUT2 #(
		.INIT('h1)
	) name2474 (
		_w6391_,
		_w6520_,
		_w6521_
	);
	LUT2 #(
		.INIT('h8)
	) name2475 (
		_w6517_,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h1)
	) name2476 (
		_w6444_,
		_w6519_,
		_w6523_
	);
	LUT2 #(
		.INIT('h4)
	) name2477 (
		_w6522_,
		_w6523_,
		_w6524_
	);
	LUT2 #(
		.INIT('h4)
	) name2478 (
		_w6518_,
		_w6524_,
		_w6525_
	);
	LUT2 #(
		.INIT('h1)
	) name2479 (
		_w6472_,
		_w6525_,
		_w6526_
	);
	LUT2 #(
		.INIT('h1)
	) name2480 (
		_w6473_,
		_w6526_,
		_w6527_
	);
	LUT2 #(
		.INIT('h8)
	) name2481 (
		_w6499_,
		_w6527_,
		_w6528_
	);
	LUT2 #(
		.INIT('h1)
	) name2482 (
		_w6499_,
		_w6527_,
		_w6529_
	);
	LUT2 #(
		.INIT('h1)
	) name2483 (
		_w6528_,
		_w6529_,
		_w6530_
	);
	LUT2 #(
		.INIT('h1)
	) name2484 (
		_w6496_,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h1)
	) name2485 (
		_w6479_,
		_w6489_,
		_w6532_
	);
	LUT2 #(
		.INIT('h1)
	) name2486 (
		_w6465_,
		_w6486_,
		_w6533_
	);
	LUT2 #(
		.INIT('h1)
	) name2487 (
		_w6490_,
		_w6533_,
		_w6534_
	);
	LUT2 #(
		.INIT('h2)
	) name2488 (
		_w6532_,
		_w6534_,
		_w6535_
	);
	LUT2 #(
		.INIT('h4)
	) name2489 (
		_w6532_,
		_w6534_,
		_w6536_
	);
	LUT2 #(
		.INIT('h1)
	) name2490 (
		_w6535_,
		_w6536_,
		_w6537_
	);
	LUT2 #(
		.INIT('h2)
	) name2491 (
		_w6496_,
		_w6537_,
		_w6538_
	);
	LUT2 #(
		.INIT('h1)
	) name2492 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6531_,
		_w6539_
	);
	LUT2 #(
		.INIT('h4)
	) name2493 (
		_w6538_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h1)
	) name2494 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		_w6537_,
		_w6541_
	);
	LUT2 #(
		.INIT('h8)
	) name2495 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6530_,
		_w6542_
	);
	LUT2 #(
		.INIT('h4)
	) name2496 (
		_w6541_,
		_w6542_,
		_w6543_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		_w6229_,
		_w6544_
	);
	LUT2 #(
		.INIT('h1)
	) name2498 (
		_w6543_,
		_w6544_,
		_w6545_
	);
	LUT2 #(
		.INIT('h4)
	) name2499 (
		_w6540_,
		_w6545_,
		_w6546_
	);
	LUT2 #(
		.INIT('h2)
	) name2500 (
		_w6135_,
		_w6546_,
		_w6547_
	);
	LUT2 #(
		.INIT('h4)
	) name2501 (
		_w6161_,
		_w6176_,
		_w6548_
	);
	LUT2 #(
		.INIT('h4)
	) name2502 (
		_w6547_,
		_w6548_,
		_w6549_
	);
	LUT2 #(
		.INIT('h1)
	) name2503 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		_w6550_
	);
	LUT2 #(
		.INIT('h4)
	) name2504 (
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w6550_,
		_w6551_
	);
	LUT2 #(
		.INIT('h1)
	) name2505 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w6552_
	);
	LUT2 #(
		.INIT('h1)
	) name2506 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		_w6553_
	);
	LUT2 #(
		.INIT('h8)
	) name2507 (
		_w6552_,
		_w6553_,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name2508 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w6555_
	);
	LUT2 #(
		.INIT('h4)
	) name2509 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w6555_,
		_w6556_
	);
	LUT2 #(
		.INIT('h8)
	) name2510 (
		_w6554_,
		_w6556_,
		_w6557_
	);
	LUT2 #(
		.INIT('h1)
	) name2511 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w6558_
	);
	LUT2 #(
		.INIT('h4)
	) name2512 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		_w6558_,
		_w6559_
	);
	LUT2 #(
		.INIT('h8)
	) name2513 (
		_w6557_,
		_w6559_,
		_w6560_
	);
	LUT2 #(
		.INIT('h4)
	) name2514 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		_w6560_,
		_w6561_
	);
	LUT2 #(
		.INIT('h1)
	) name2515 (
		_w6551_,
		_w6561_,
		_w6562_
	);
	LUT2 #(
		.INIT('h1)
	) name2516 (
		_w6556_,
		_w6558_,
		_w6563_
	);
	LUT2 #(
		.INIT('h2)
	) name2517 (
		_w6554_,
		_w6563_,
		_w6564_
	);
	LUT2 #(
		.INIT('h4)
	) name2518 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		_w6552_,
		_w6565_
	);
	LUT2 #(
		.INIT('h2)
	) name2519 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		_w6565_,
		_w6566_
	);
	LUT2 #(
		.INIT('h4)
	) name2520 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w6558_,
		_w6567_
	);
	LUT2 #(
		.INIT('h4)
	) name2521 (
		_w6566_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h1)
	) name2522 (
		_w6564_,
		_w6568_,
		_w6569_
	);
	LUT2 #(
		.INIT('h4)
	) name2523 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w6554_,
		_w6570_
	);
	LUT2 #(
		.INIT('h1)
	) name2524 (
		_w6555_,
		_w6570_,
		_w6571_
	);
	LUT2 #(
		.INIT('h2)
	) name2525 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		_w6552_,
		_w6572_
	);
	LUT2 #(
		.INIT('h1)
	) name2526 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w6573_
	);
	LUT2 #(
		.INIT('h2)
	) name2527 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		_w6573_,
		_w6574_
	);
	LUT2 #(
		.INIT('h8)
	) name2528 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w6575_
	);
	LUT2 #(
		.INIT('h8)
	) name2529 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w6576_
	);
	LUT2 #(
		.INIT('h8)
	) name2530 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w6577_
	);
	LUT2 #(
		.INIT('h8)
	) name2531 (
		_w6557_,
		_w6558_,
		_w6578_
	);
	LUT2 #(
		.INIT('h2)
	) name2532 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		_w6578_,
		_w6579_
	);
	LUT2 #(
		.INIT('h2)
	) name2533 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		_w6560_,
		_w6580_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w6575_,
		_w6576_,
		_w6581_
	);
	LUT2 #(
		.INIT('h4)
	) name2535 (
		_w6577_,
		_w6581_,
		_w6582_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w6572_,
		_w6574_,
		_w6583_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		_w6582_,
		_w6583_,
		_w6584_
	);
	LUT2 #(
		.INIT('h4)
	) name2538 (
		_w6571_,
		_w6584_,
		_w6585_
	);
	LUT2 #(
		.INIT('h4)
	) name2539 (
		_w6569_,
		_w6585_,
		_w6586_
	);
	LUT2 #(
		.INIT('h1)
	) name2540 (
		_w6579_,
		_w6580_,
		_w6587_
	);
	LUT2 #(
		.INIT('h8)
	) name2541 (
		_w6586_,
		_w6587_,
		_w6588_
	);
	LUT2 #(
		.INIT('h8)
	) name2542 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w6589_
	);
	LUT2 #(
		.INIT('h2)
	) name2543 (
		_w6588_,
		_w6589_,
		_w6590_
	);
	LUT2 #(
		.INIT('h4)
	) name2544 (
		_w6562_,
		_w6590_,
		_w6591_
	);
	LUT2 #(
		.INIT('h8)
	) name2545 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		_w6591_,
		_w6592_
	);
	LUT2 #(
		.INIT('h8)
	) name2546 (
		\core_dag_ilm2reg_I_reg[0]/NET0131 ,
		_w6592_,
		_w6593_
	);
	LUT2 #(
		.INIT('h2)
	) name2547 (
		\core_dag_ilm2reg_I_reg[0]/NET0131 ,
		_w6592_,
		_w6594_
	);
	LUT2 #(
		.INIT('h1)
	) name2548 (
		\core_dag_ilm2reg_M_reg[0]/NET0131 ,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h8)
	) name2549 (
		\core_dag_ilm2reg_M_reg[0]/NET0131 ,
		_w6594_,
		_w6596_
	);
	LUT2 #(
		.INIT('h1)
	) name2550 (
		_w6595_,
		_w6596_,
		_w6597_
	);
	LUT2 #(
		.INIT('h2)
	) name2551 (
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w6591_,
		_w6598_
	);
	LUT2 #(
		.INIT('h4)
	) name2552 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		_w6551_,
		_w6599_
	);
	LUT2 #(
		.INIT('h8)
	) name2553 (
		_w6559_,
		_w6599_,
		_w6600_
	);
	LUT2 #(
		.INIT('h8)
	) name2554 (
		_w6555_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h8)
	) name2555 (
		_w6570_,
		_w6601_,
		_w6602_
	);
	LUT2 #(
		.INIT('h8)
	) name2556 (
		_w6591_,
		_w6602_,
		_w6603_
	);
	LUT2 #(
		.INIT('h1)
	) name2557 (
		_w6598_,
		_w6603_,
		_w6604_
	);
	LUT2 #(
		.INIT('h2)
	) name2558 (
		\core_dag_ilm2reg_I_reg[13]/NET0131 ,
		_w6604_,
		_w6605_
	);
	LUT2 #(
		.INIT('h8)
	) name2559 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h4)
	) name2560 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w6601_,
		_w6607_
	);
	LUT2 #(
		.INIT('h8)
	) name2561 (
		_w6553_,
		_w6607_,
		_w6608_
	);
	LUT2 #(
		.INIT('h2)
	) name2562 (
		_w6591_,
		_w6608_,
		_w6609_
	);
	LUT2 #(
		.INIT('h8)
	) name2563 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		_w6591_,
		_w6610_
	);
	LUT2 #(
		.INIT('h2)
	) name2564 (
		_w6552_,
		_w6591_,
		_w6611_
	);
	LUT2 #(
		.INIT('h1)
	) name2565 (
		_w6609_,
		_w6610_,
		_w6612_
	);
	LUT2 #(
		.INIT('h4)
	) name2566 (
		_w6611_,
		_w6612_,
		_w6613_
	);
	LUT2 #(
		.INIT('h8)
	) name2567 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		_w6613_,
		_w6614_
	);
	LUT2 #(
		.INIT('h8)
	) name2568 (
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w6614_,
		_w6615_
	);
	LUT2 #(
		.INIT('h1)
	) name2569 (
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w6614_,
		_w6616_
	);
	LUT2 #(
		.INIT('h4)
	) name2570 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		_w6607_,
		_w6617_
	);
	LUT2 #(
		.INIT('h2)
	) name2571 (
		_w6591_,
		_w6617_,
		_w6618_
	);
	LUT2 #(
		.INIT('h8)
	) name2572 (
		_w6553_,
		_w6611_,
		_w6619_
	);
	LUT2 #(
		.INIT('h1)
	) name2573 (
		_w6618_,
		_w6619_,
		_w6620_
	);
	LUT2 #(
		.INIT('h8)
	) name2574 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		_w6620_,
		_w6621_
	);
	LUT2 #(
		.INIT('h1)
	) name2575 (
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w6621_,
		_w6622_
	);
	LUT2 #(
		.INIT('h2)
	) name2576 (
		_w6565_,
		_w6591_,
		_w6623_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		_w6609_,
		_w6623_,
		_w6624_
	);
	LUT2 #(
		.INIT('h8)
	) name2578 (
		\core_dag_ilm2reg_I_reg[11]/NET0131 ,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w6625_,
		_w6626_
	);
	LUT2 #(
		.INIT('h1)
	) name2580 (
		_w6622_,
		_w6626_,
		_w6627_
	);
	LUT2 #(
		.INIT('h2)
	) name2581 (
		_w6591_,
		_w6607_,
		_w6628_
	);
	LUT2 #(
		.INIT('h4)
	) name2582 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w6619_,
		_w6629_
	);
	LUT2 #(
		.INIT('h1)
	) name2583 (
		_w6628_,
		_w6629_,
		_w6630_
	);
	LUT2 #(
		.INIT('h8)
	) name2584 (
		\core_dag_ilm2reg_I_reg[9]/NET0131 ,
		_w6630_,
		_w6631_
	);
	LUT2 #(
		.INIT('h1)
	) name2585 (
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w6631_,
		_w6632_
	);
	LUT2 #(
		.INIT('h4)
	) name2586 (
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w6629_,
		_w6633_
	);
	LUT2 #(
		.INIT('h2)
	) name2587 (
		_w6591_,
		_w6601_,
		_w6634_
	);
	LUT2 #(
		.INIT('h1)
	) name2588 (
		_w6633_,
		_w6634_,
		_w6635_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		\core_dag_ilm2reg_I_reg[8]/NET0131 ,
		_w6635_,
		_w6636_
	);
	LUT2 #(
		.INIT('h1)
	) name2590 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w6636_,
		_w6637_
	);
	LUT2 #(
		.INIT('h8)
	) name2591 (
		_w6556_,
		_w6619_,
		_w6638_
	);
	LUT2 #(
		.INIT('h8)
	) name2592 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		_w6591_,
		_w6639_
	);
	LUT2 #(
		.INIT('h2)
	) name2593 (
		_w6591_,
		_w6600_,
		_w6640_
	);
	LUT2 #(
		.INIT('h1)
	) name2594 (
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT2 #(
		.INIT('h4)
	) name2595 (
		_w6638_,
		_w6641_,
		_w6642_
	);
	LUT2 #(
		.INIT('h8)
	) name2596 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		_w6642_,
		_w6643_
	);
	LUT2 #(
		.INIT('h1)
	) name2597 (
		\core_dag_ilm2reg_M_reg[7]/NET0131 ,
		_w6643_,
		_w6644_
	);
	LUT2 #(
		.INIT('h8)
	) name2598 (
		\core_dag_ilm2reg_M_reg[7]/NET0131 ,
		_w6643_,
		_w6645_
	);
	LUT2 #(
		.INIT('h4)
	) name2599 (
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w6638_,
		_w6646_
	);
	LUT2 #(
		.INIT('h1)
	) name2600 (
		_w6640_,
		_w6646_,
		_w6647_
	);
	LUT2 #(
		.INIT('h8)
	) name2601 (
		\core_dag_ilm2reg_I_reg[6]/NET0131 ,
		_w6647_,
		_w6648_
	);
	LUT2 #(
		.INIT('h1)
	) name2602 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w6648_,
		_w6649_
	);
	LUT2 #(
		.INIT('h8)
	) name2603 (
		\core_dag_ilm2reg_M_reg[6]/NET0131 ,
		_w6648_,
		_w6650_
	);
	LUT2 #(
		.INIT('h2)
	) name2604 (
		_w6591_,
		_w6599_,
		_w6651_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		_w6561_,
		_w6590_,
		_w6652_
	);
	LUT2 #(
		.INIT('h1)
	) name2606 (
		_w6651_,
		_w6652_,
		_w6653_
	);
	LUT2 #(
		.INIT('h8)
	) name2607 (
		\core_dag_ilm2reg_I_reg[3]/NET0131 ,
		_w6653_,
		_w6654_
	);
	LUT2 #(
		.INIT('h1)
	) name2608 (
		\core_dag_ilm2reg_M_reg[3]/NET0131 ,
		_w6654_,
		_w6655_
	);
	LUT2 #(
		.INIT('h8)
	) name2609 (
		\core_dag_ilm2reg_M_reg[3]/NET0131 ,
		_w6654_,
		_w6656_
	);
	LUT2 #(
		.INIT('h4)
	) name2610 (
		_w6551_,
		_w6591_,
		_w6657_
	);
	LUT2 #(
		.INIT('h4)
	) name2611 (
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w6561_,
		_w6658_
	);
	LUT2 #(
		.INIT('h4)
	) name2612 (
		_w6588_,
		_w6658_,
		_w6659_
	);
	LUT2 #(
		.INIT('h1)
	) name2613 (
		_w6657_,
		_w6659_,
		_w6660_
	);
	LUT2 #(
		.INIT('h8)
	) name2614 (
		\core_dag_ilm2reg_I_reg[2]/NET0131 ,
		_w6660_,
		_w6661_
	);
	LUT2 #(
		.INIT('h1)
	) name2615 (
		\core_dag_ilm2reg_M_reg[2]/NET0131 ,
		_w6661_,
		_w6662_
	);
	LUT2 #(
		.INIT('h8)
	) name2616 (
		\core_dag_ilm2reg_M_reg[2]/NET0131 ,
		_w6661_,
		_w6663_
	);
	LUT2 #(
		.INIT('h4)
	) name2617 (
		_w6550_,
		_w6591_,
		_w6664_
	);
	LUT2 #(
		.INIT('h4)
	) name2618 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		_w6659_,
		_w6665_
	);
	LUT2 #(
		.INIT('h2)
	) name2619 (
		\core_dag_ilm2reg_I_reg[1]/NET0131 ,
		_w6665_,
		_w6666_
	);
	LUT2 #(
		.INIT('h4)
	) name2620 (
		_w6664_,
		_w6666_,
		_w6667_
	);
	LUT2 #(
		.INIT('h1)
	) name2621 (
		\core_dag_ilm2reg_M_reg[1]/NET0131 ,
		_w6667_,
		_w6668_
	);
	LUT2 #(
		.INIT('h8)
	) name2622 (
		\core_dag_ilm2reg_M_reg[1]/NET0131 ,
		_w6667_,
		_w6669_
	);
	LUT2 #(
		.INIT('h1)
	) name2623 (
		_w6596_,
		_w6669_,
		_w6670_
	);
	LUT2 #(
		.INIT('h1)
	) name2624 (
		_w6668_,
		_w6670_,
		_w6671_
	);
	LUT2 #(
		.INIT('h1)
	) name2625 (
		_w6663_,
		_w6671_,
		_w6672_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		_w6662_,
		_w6672_,
		_w6673_
	);
	LUT2 #(
		.INIT('h1)
	) name2627 (
		_w6656_,
		_w6673_,
		_w6674_
	);
	LUT2 #(
		.INIT('h1)
	) name2628 (
		_w6655_,
		_w6674_,
		_w6675_
	);
	LUT2 #(
		.INIT('h1)
	) name2629 (
		_w6578_,
		_w6591_,
		_w6676_
	);
	LUT2 #(
		.INIT('h4)
	) name2630 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		_w6599_,
		_w6677_
	);
	LUT2 #(
		.INIT('h8)
	) name2631 (
		_w6591_,
		_w6677_,
		_w6678_
	);
	LUT2 #(
		.INIT('h4)
	) name2632 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		_w6678_,
		_w6679_
	);
	LUT2 #(
		.INIT('h1)
	) name2633 (
		_w6676_,
		_w6679_,
		_w6680_
	);
	LUT2 #(
		.INIT('h2)
	) name2634 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		_w6680_,
		_w6681_
	);
	LUT2 #(
		.INIT('h1)
	) name2635 (
		\core_dag_ilm2reg_M_reg[5]/NET0131 ,
		_w6681_,
		_w6682_
	);
	LUT2 #(
		.INIT('h1)
	) name2636 (
		_w6560_,
		_w6591_,
		_w6683_
	);
	LUT2 #(
		.INIT('h1)
	) name2637 (
		_w6678_,
		_w6683_,
		_w6684_
	);
	LUT2 #(
		.INIT('h2)
	) name2638 (
		\core_dag_ilm2reg_I_reg[4]/NET0131 ,
		_w6684_,
		_w6685_
	);
	LUT2 #(
		.INIT('h1)
	) name2639 (
		\core_dag_ilm2reg_M_reg[4]/NET0131 ,
		_w6685_,
		_w6686_
	);
	LUT2 #(
		.INIT('h1)
	) name2640 (
		_w6682_,
		_w6686_,
		_w6687_
	);
	LUT2 #(
		.INIT('h8)
	) name2641 (
		_w6675_,
		_w6687_,
		_w6688_
	);
	LUT2 #(
		.INIT('h8)
	) name2642 (
		\core_dag_ilm2reg_M_reg[5]/NET0131 ,
		_w6681_,
		_w6689_
	);
	LUT2 #(
		.INIT('h8)
	) name2643 (
		\core_dag_ilm2reg_M_reg[4]/NET0131 ,
		_w6685_,
		_w6690_
	);
	LUT2 #(
		.INIT('h4)
	) name2644 (
		_w6682_,
		_w6690_,
		_w6691_
	);
	LUT2 #(
		.INIT('h1)
	) name2645 (
		_w6689_,
		_w6691_,
		_w6692_
	);
	LUT2 #(
		.INIT('h4)
	) name2646 (
		_w6688_,
		_w6692_,
		_w6693_
	);
	LUT2 #(
		.INIT('h4)
	) name2647 (
		_w6650_,
		_w6693_,
		_w6694_
	);
	LUT2 #(
		.INIT('h1)
	) name2648 (
		_w6649_,
		_w6694_,
		_w6695_
	);
	LUT2 #(
		.INIT('h1)
	) name2649 (
		_w6645_,
		_w6695_,
		_w6696_
	);
	LUT2 #(
		.INIT('h1)
	) name2650 (
		_w6644_,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h4)
	) name2651 (
		_w6637_,
		_w6697_,
		_w6698_
	);
	LUT2 #(
		.INIT('h4)
	) name2652 (
		_w6632_,
		_w6698_,
		_w6699_
	);
	LUT2 #(
		.INIT('h8)
	) name2653 (
		_w6627_,
		_w6699_,
		_w6700_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w6625_,
		_w6701_
	);
	LUT2 #(
		.INIT('h8)
	) name2655 (
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w6621_,
		_w6702_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w6636_,
		_w6703_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w6631_,
		_w6704_
	);
	LUT2 #(
		.INIT('h1)
	) name2658 (
		_w6703_,
		_w6704_,
		_w6705_
	);
	LUT2 #(
		.INIT('h1)
	) name2659 (
		_w6632_,
		_w6705_,
		_w6706_
	);
	LUT2 #(
		.INIT('h1)
	) name2660 (
		_w6702_,
		_w6706_,
		_w6707_
	);
	LUT2 #(
		.INIT('h2)
	) name2661 (
		_w6627_,
		_w6707_,
		_w6708_
	);
	LUT2 #(
		.INIT('h1)
	) name2662 (
		_w6701_,
		_w6708_,
		_w6709_
	);
	LUT2 #(
		.INIT('h4)
	) name2663 (
		_w6700_,
		_w6709_,
		_w6710_
	);
	LUT2 #(
		.INIT('h1)
	) name2664 (
		_w6616_,
		_w6710_,
		_w6711_
	);
	LUT2 #(
		.INIT('h1)
	) name2665 (
		_w6615_,
		_w6711_,
		_w6712_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		_w6606_,
		_w6712_,
		_w6713_
	);
	LUT2 #(
		.INIT('h2)
	) name2667 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6713_,
		_w6714_
	);
	LUT2 #(
		.INIT('h2)
	) name2668 (
		_w6605_,
		_w6712_,
		_w6715_
	);
	LUT2 #(
		.INIT('h1)
	) name2669 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6715_,
		_w6716_
	);
	LUT2 #(
		.INIT('h1)
	) name2670 (
		_w6714_,
		_w6716_,
		_w6717_
	);
	LUT2 #(
		.INIT('h2)
	) name2671 (
		_w6597_,
		_w6717_,
		_w6718_
	);
	LUT2 #(
		.INIT('h1)
	) name2672 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6719_
	);
	LUT2 #(
		.INIT('h8)
	) name2673 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6720_
	);
	LUT2 #(
		.INIT('h1)
	) name2674 (
		_w6719_,
		_w6720_,
		_w6721_
	);
	LUT2 #(
		.INIT('h4)
	) name2675 (
		_w6597_,
		_w6721_,
		_w6722_
	);
	LUT2 #(
		.INIT('h2)
	) name2676 (
		_w6597_,
		_w6721_,
		_w6723_
	);
	LUT2 #(
		.INIT('h1)
	) name2677 (
		_w6722_,
		_w6723_,
		_w6724_
	);
	LUT2 #(
		.INIT('h8)
	) name2678 (
		_w6713_,
		_w6724_,
		_w6725_
	);
	LUT2 #(
		.INIT('h1)
	) name2679 (
		_w6718_,
		_w6725_,
		_w6726_
	);
	LUT2 #(
		.INIT('h2)
	) name2680 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6726_,
		_w6727_
	);
	LUT2 #(
		.INIT('h1)
	) name2681 (
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w6605_,
		_w6728_
	);
	LUT2 #(
		.INIT('h2)
	) name2682 (
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6729_
	);
	LUT2 #(
		.INIT('h1)
	) name2683 (
		_w6728_,
		_w6729_,
		_w6730_
	);
	LUT2 #(
		.INIT('h1)
	) name2684 (
		_w6644_,
		_w6645_,
		_w6731_
	);
	LUT2 #(
		.INIT('h1)
	) name2685 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6732_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6733_
	);
	LUT2 #(
		.INIT('h1)
	) name2687 (
		_w6732_,
		_w6733_,
		_w6734_
	);
	LUT2 #(
		.INIT('h2)
	) name2688 (
		_w6731_,
		_w6734_,
		_w6735_
	);
	LUT2 #(
		.INIT('h4)
	) name2689 (
		_w6731_,
		_w6734_,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name2690 (
		_w6735_,
		_w6736_,
		_w6737_
	);
	LUT2 #(
		.INIT('h1)
	) name2691 (
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6738_
	);
	LUT2 #(
		.INIT('h8)
	) name2692 (
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6739_
	);
	LUT2 #(
		.INIT('h1)
	) name2693 (
		_w6738_,
		_w6739_,
		_w6740_
	);
	LUT2 #(
		.INIT('h1)
	) name2694 (
		_w6649_,
		_w6740_,
		_w6741_
	);
	LUT2 #(
		.INIT('h1)
	) name2695 (
		_w6650_,
		_w6741_,
		_w6742_
	);
	LUT2 #(
		.INIT('h4)
	) name2696 (
		_w6737_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6744_
	);
	LUT2 #(
		.INIT('h8)
	) name2698 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6745_
	);
	LUT2 #(
		.INIT('h1)
	) name2699 (
		_w6744_,
		_w6745_,
		_w6746_
	);
	LUT2 #(
		.INIT('h1)
	) name2700 (
		_w6682_,
		_w6746_,
		_w6747_
	);
	LUT2 #(
		.INIT('h1)
	) name2701 (
		_w6689_,
		_w6747_,
		_w6748_
	);
	LUT2 #(
		.INIT('h1)
	) name2702 (
		_w6649_,
		_w6650_,
		_w6749_
	);
	LUT2 #(
		.INIT('h2)
	) name2703 (
		_w6740_,
		_w6749_,
		_w6750_
	);
	LUT2 #(
		.INIT('h4)
	) name2704 (
		_w6740_,
		_w6749_,
		_w6751_
	);
	LUT2 #(
		.INIT('h1)
	) name2705 (
		_w6750_,
		_w6751_,
		_w6752_
	);
	LUT2 #(
		.INIT('h2)
	) name2706 (
		_w6748_,
		_w6752_,
		_w6753_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6754_
	);
	LUT2 #(
		.INIT('h8)
	) name2708 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6755_
	);
	LUT2 #(
		.INIT('h1)
	) name2709 (
		_w6754_,
		_w6755_,
		_w6756_
	);
	LUT2 #(
		.INIT('h1)
	) name2710 (
		_w6686_,
		_w6756_,
		_w6757_
	);
	LUT2 #(
		.INIT('h1)
	) name2711 (
		_w6690_,
		_w6757_,
		_w6758_
	);
	LUT2 #(
		.INIT('h1)
	) name2712 (
		_w6682_,
		_w6689_,
		_w6759_
	);
	LUT2 #(
		.INIT('h2)
	) name2713 (
		_w6746_,
		_w6759_,
		_w6760_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		_w6746_,
		_w6759_,
		_w6761_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w6760_,
		_w6761_,
		_w6762_
	);
	LUT2 #(
		.INIT('h4)
	) name2716 (
		_w6758_,
		_w6762_,
		_w6763_
	);
	LUT2 #(
		.INIT('h2)
	) name2717 (
		_w6758_,
		_w6762_,
		_w6764_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6765_
	);
	LUT2 #(
		.INIT('h8)
	) name2719 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6766_
	);
	LUT2 #(
		.INIT('h1)
	) name2720 (
		_w6765_,
		_w6766_,
		_w6767_
	);
	LUT2 #(
		.INIT('h1)
	) name2721 (
		_w6655_,
		_w6767_,
		_w6768_
	);
	LUT2 #(
		.INIT('h1)
	) name2722 (
		_w6656_,
		_w6768_,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		_w6686_,
		_w6690_,
		_w6770_
	);
	LUT2 #(
		.INIT('h2)
	) name2724 (
		_w6756_,
		_w6770_,
		_w6771_
	);
	LUT2 #(
		.INIT('h4)
	) name2725 (
		_w6756_,
		_w6770_,
		_w6772_
	);
	LUT2 #(
		.INIT('h1)
	) name2726 (
		_w6771_,
		_w6772_,
		_w6773_
	);
	LUT2 #(
		.INIT('h4)
	) name2727 (
		_w6769_,
		_w6773_,
		_w6774_
	);
	LUT2 #(
		.INIT('h4)
	) name2728 (
		_w6764_,
		_w6774_,
		_w6775_
	);
	LUT2 #(
		.INIT('h1)
	) name2729 (
		_w6763_,
		_w6775_,
		_w6776_
	);
	LUT2 #(
		.INIT('h1)
	) name2730 (
		_w6753_,
		_w6776_,
		_w6777_
	);
	LUT2 #(
		.INIT('h4)
	) name2731 (
		_w6748_,
		_w6752_,
		_w6778_
	);
	LUT2 #(
		.INIT('h2)
	) name2732 (
		_w6737_,
		_w6742_,
		_w6779_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		_w6778_,
		_w6779_,
		_w6780_
	);
	LUT2 #(
		.INIT('h4)
	) name2734 (
		_w6777_,
		_w6780_,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name2735 (
		_w6743_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h1)
	) name2736 (
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6783_
	);
	LUT2 #(
		.INIT('h8)
	) name2737 (
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6784_
	);
	LUT2 #(
		.INIT('h1)
	) name2738 (
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT2 #(
		.INIT('h1)
	) name2739 (
		_w6662_,
		_w6785_,
		_w6786_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		_w6663_,
		_w6786_,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name2741 (
		_w6655_,
		_w6656_,
		_w6788_
	);
	LUT2 #(
		.INIT('h2)
	) name2742 (
		_w6767_,
		_w6788_,
		_w6789_
	);
	LUT2 #(
		.INIT('h4)
	) name2743 (
		_w6767_,
		_w6788_,
		_w6790_
	);
	LUT2 #(
		.INIT('h1)
	) name2744 (
		_w6789_,
		_w6790_,
		_w6791_
	);
	LUT2 #(
		.INIT('h2)
	) name2745 (
		_w6787_,
		_w6791_,
		_w6792_
	);
	LUT2 #(
		.INIT('h4)
	) name2746 (
		_w6787_,
		_w6791_,
		_w6793_
	);
	LUT2 #(
		.INIT('h1)
	) name2747 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6794_
	);
	LUT2 #(
		.INIT('h8)
	) name2748 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6795_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		_w6794_,
		_w6795_,
		_w6796_
	);
	LUT2 #(
		.INIT('h1)
	) name2750 (
		_w6668_,
		_w6796_,
		_w6797_
	);
	LUT2 #(
		.INIT('h1)
	) name2751 (
		_w6669_,
		_w6797_,
		_w6798_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		_w6662_,
		_w6663_,
		_w6799_
	);
	LUT2 #(
		.INIT('h2)
	) name2753 (
		_w6785_,
		_w6799_,
		_w6800_
	);
	LUT2 #(
		.INIT('h4)
	) name2754 (
		_w6785_,
		_w6799_,
		_w6801_
	);
	LUT2 #(
		.INIT('h1)
	) name2755 (
		_w6800_,
		_w6801_,
		_w6802_
	);
	LUT2 #(
		.INIT('h2)
	) name2756 (
		_w6798_,
		_w6802_,
		_w6803_
	);
	LUT2 #(
		.INIT('h4)
	) name2757 (
		_w6798_,
		_w6802_,
		_w6804_
	);
	LUT2 #(
		.INIT('h4)
	) name2758 (
		_w6596_,
		_w6721_,
		_w6805_
	);
	LUT2 #(
		.INIT('h1)
	) name2759 (
		_w6595_,
		_w6805_,
		_w6806_
	);
	LUT2 #(
		.INIT('h1)
	) name2760 (
		_w6668_,
		_w6669_,
		_w6807_
	);
	LUT2 #(
		.INIT('h2)
	) name2761 (
		_w6796_,
		_w6807_,
		_w6808_
	);
	LUT2 #(
		.INIT('h4)
	) name2762 (
		_w6796_,
		_w6807_,
		_w6809_
	);
	LUT2 #(
		.INIT('h1)
	) name2763 (
		_w6808_,
		_w6809_,
		_w6810_
	);
	LUT2 #(
		.INIT('h1)
	) name2764 (
		_w6806_,
		_w6810_,
		_w6811_
	);
	LUT2 #(
		.INIT('h8)
	) name2765 (
		_w6806_,
		_w6810_,
		_w6812_
	);
	LUT2 #(
		.INIT('h4)
	) name2766 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6724_,
		_w6813_
	);
	LUT2 #(
		.INIT('h1)
	) name2767 (
		_w6812_,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h1)
	) name2768 (
		_w6811_,
		_w6814_,
		_w6815_
	);
	LUT2 #(
		.INIT('h1)
	) name2769 (
		_w6804_,
		_w6815_,
		_w6816_
	);
	LUT2 #(
		.INIT('h1)
	) name2770 (
		_w6803_,
		_w6816_,
		_w6817_
	);
	LUT2 #(
		.INIT('h1)
	) name2771 (
		_w6793_,
		_w6817_,
		_w6818_
	);
	LUT2 #(
		.INIT('h1)
	) name2772 (
		_w6792_,
		_w6818_,
		_w6819_
	);
	LUT2 #(
		.INIT('h2)
	) name2773 (
		_w6769_,
		_w6773_,
		_w6820_
	);
	LUT2 #(
		.INIT('h1)
	) name2774 (
		_w6764_,
		_w6820_,
		_w6821_
	);
	LUT2 #(
		.INIT('h4)
	) name2775 (
		_w6743_,
		_w6821_,
		_w6822_
	);
	LUT2 #(
		.INIT('h4)
	) name2776 (
		_w6753_,
		_w6822_,
		_w6823_
	);
	LUT2 #(
		.INIT('h8)
	) name2777 (
		_w6819_,
		_w6823_,
		_w6824_
	);
	LUT2 #(
		.INIT('h1)
	) name2778 (
		_w6782_,
		_w6824_,
		_w6825_
	);
	LUT2 #(
		.INIT('h1)
	) name2779 (
		_w6632_,
		_w6704_,
		_w6826_
	);
	LUT2 #(
		.INIT('h1)
	) name2780 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6827_
	);
	LUT2 #(
		.INIT('h8)
	) name2781 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6828_
	);
	LUT2 #(
		.INIT('h1)
	) name2782 (
		_w6827_,
		_w6828_,
		_w6829_
	);
	LUT2 #(
		.INIT('h2)
	) name2783 (
		_w6826_,
		_w6829_,
		_w6830_
	);
	LUT2 #(
		.INIT('h4)
	) name2784 (
		_w6826_,
		_w6829_,
		_w6831_
	);
	LUT2 #(
		.INIT('h1)
	) name2785 (
		_w6830_,
		_w6831_,
		_w6832_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6833_
	);
	LUT2 #(
		.INIT('h8)
	) name2787 (
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6834_
	);
	LUT2 #(
		.INIT('h1)
	) name2788 (
		_w6833_,
		_w6834_,
		_w6835_
	);
	LUT2 #(
		.INIT('h1)
	) name2789 (
		_w6637_,
		_w6835_,
		_w6836_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		_w6703_,
		_w6836_,
		_w6837_
	);
	LUT2 #(
		.INIT('h4)
	) name2791 (
		_w6832_,
		_w6837_,
		_w6838_
	);
	LUT2 #(
		.INIT('h1)
	) name2792 (
		_w6644_,
		_w6734_,
		_w6839_
	);
	LUT2 #(
		.INIT('h1)
	) name2793 (
		_w6645_,
		_w6839_,
		_w6840_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		_w6637_,
		_w6703_,
		_w6841_
	);
	LUT2 #(
		.INIT('h2)
	) name2795 (
		_w6835_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h4)
	) name2796 (
		_w6835_,
		_w6841_,
		_w6843_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		_w6842_,
		_w6843_,
		_w6844_
	);
	LUT2 #(
		.INIT('h2)
	) name2798 (
		_w6840_,
		_w6844_,
		_w6845_
	);
	LUT2 #(
		.INIT('h1)
	) name2799 (
		_w6838_,
		_w6845_,
		_w6846_
	);
	LUT2 #(
		.INIT('h4)
	) name2800 (
		_w6825_,
		_w6846_,
		_w6847_
	);
	LUT2 #(
		.INIT('h1)
	) name2801 (
		_w6632_,
		_w6829_,
		_w6848_
	);
	LUT2 #(
		.INIT('h1)
	) name2802 (
		_w6704_,
		_w6848_,
		_w6849_
	);
	LUT2 #(
		.INIT('h1)
	) name2803 (
		_w6622_,
		_w6702_,
		_w6850_
	);
	LUT2 #(
		.INIT('h1)
	) name2804 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6851_
	);
	LUT2 #(
		.INIT('h8)
	) name2805 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6852_
	);
	LUT2 #(
		.INIT('h1)
	) name2806 (
		_w6851_,
		_w6852_,
		_w6853_
	);
	LUT2 #(
		.INIT('h2)
	) name2807 (
		_w6850_,
		_w6853_,
		_w6854_
	);
	LUT2 #(
		.INIT('h4)
	) name2808 (
		_w6850_,
		_w6853_,
		_w6855_
	);
	LUT2 #(
		.INIT('h1)
	) name2809 (
		_w6854_,
		_w6855_,
		_w6856_
	);
	LUT2 #(
		.INIT('h2)
	) name2810 (
		_w6849_,
		_w6856_,
		_w6857_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w6622_,
		_w6853_,
		_w6858_
	);
	LUT2 #(
		.INIT('h1)
	) name2812 (
		_w6702_,
		_w6858_,
		_w6859_
	);
	LUT2 #(
		.INIT('h1)
	) name2813 (
		_w6626_,
		_w6701_,
		_w6860_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6861_
	);
	LUT2 #(
		.INIT('h8)
	) name2815 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6862_
	);
	LUT2 #(
		.INIT('h1)
	) name2816 (
		_w6861_,
		_w6862_,
		_w6863_
	);
	LUT2 #(
		.INIT('h2)
	) name2817 (
		_w6860_,
		_w6863_,
		_w6864_
	);
	LUT2 #(
		.INIT('h4)
	) name2818 (
		_w6860_,
		_w6863_,
		_w6865_
	);
	LUT2 #(
		.INIT('h1)
	) name2819 (
		_w6864_,
		_w6865_,
		_w6866_
	);
	LUT2 #(
		.INIT('h2)
	) name2820 (
		_w6859_,
		_w6866_,
		_w6867_
	);
	LUT2 #(
		.INIT('h1)
	) name2821 (
		_w6857_,
		_w6867_,
		_w6868_
	);
	LUT2 #(
		.INIT('h8)
	) name2822 (
		_w6847_,
		_w6868_,
		_w6869_
	);
	LUT2 #(
		.INIT('h4)
	) name2823 (
		_w6849_,
		_w6856_,
		_w6870_
	);
	LUT2 #(
		.INIT('h4)
	) name2824 (
		_w6867_,
		_w6870_,
		_w6871_
	);
	LUT2 #(
		.INIT('h2)
	) name2825 (
		_w6832_,
		_w6837_,
		_w6872_
	);
	LUT2 #(
		.INIT('h4)
	) name2826 (
		_w6840_,
		_w6844_,
		_w6873_
	);
	LUT2 #(
		.INIT('h4)
	) name2827 (
		_w6838_,
		_w6873_,
		_w6874_
	);
	LUT2 #(
		.INIT('h1)
	) name2828 (
		_w6872_,
		_w6874_,
		_w6875_
	);
	LUT2 #(
		.INIT('h2)
	) name2829 (
		_w6868_,
		_w6875_,
		_w6876_
	);
	LUT2 #(
		.INIT('h4)
	) name2830 (
		_w6859_,
		_w6866_,
		_w6877_
	);
	LUT2 #(
		.INIT('h1)
	) name2831 (
		_w6871_,
		_w6877_,
		_w6878_
	);
	LUT2 #(
		.INIT('h4)
	) name2832 (
		_w6876_,
		_w6878_,
		_w6879_
	);
	LUT2 #(
		.INIT('h4)
	) name2833 (
		_w6869_,
		_w6879_,
		_w6880_
	);
	LUT2 #(
		.INIT('h8)
	) name2834 (
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w6605_,
		_w6881_
	);
	LUT2 #(
		.INIT('h1)
	) name2835 (
		_w6728_,
		_w6881_,
		_w6882_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6883_
	);
	LUT2 #(
		.INIT('h8)
	) name2837 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6884_
	);
	LUT2 #(
		.INIT('h1)
	) name2838 (
		_w6883_,
		_w6884_,
		_w6885_
	);
	LUT2 #(
		.INIT('h4)
	) name2839 (
		_w6615_,
		_w6885_,
		_w6886_
	);
	LUT2 #(
		.INIT('h1)
	) name2840 (
		_w6616_,
		_w6886_,
		_w6887_
	);
	LUT2 #(
		.INIT('h2)
	) name2841 (
		_w6882_,
		_w6887_,
		_w6888_
	);
	LUT2 #(
		.INIT('h1)
	) name2842 (
		_w6626_,
		_w6863_,
		_w6889_
	);
	LUT2 #(
		.INIT('h1)
	) name2843 (
		_w6701_,
		_w6889_,
		_w6890_
	);
	LUT2 #(
		.INIT('h1)
	) name2844 (
		_w6615_,
		_w6616_,
		_w6891_
	);
	LUT2 #(
		.INIT('h4)
	) name2845 (
		_w6885_,
		_w6891_,
		_w6892_
	);
	LUT2 #(
		.INIT('h2)
	) name2846 (
		_w6885_,
		_w6891_,
		_w6893_
	);
	LUT2 #(
		.INIT('h1)
	) name2847 (
		_w6892_,
		_w6893_,
		_w6894_
	);
	LUT2 #(
		.INIT('h2)
	) name2848 (
		_w6890_,
		_w6894_,
		_w6895_
	);
	LUT2 #(
		.INIT('h1)
	) name2849 (
		_w6888_,
		_w6895_,
		_w6896_
	);
	LUT2 #(
		.INIT('h4)
	) name2850 (
		_w6880_,
		_w6896_,
		_w6897_
	);
	LUT2 #(
		.INIT('h4)
	) name2851 (
		_w6882_,
		_w6887_,
		_w6898_
	);
	LUT2 #(
		.INIT('h4)
	) name2852 (
		_w6890_,
		_w6894_,
		_w6899_
	);
	LUT2 #(
		.INIT('h4)
	) name2853 (
		_w6888_,
		_w6899_,
		_w6900_
	);
	LUT2 #(
		.INIT('h1)
	) name2854 (
		_w6898_,
		_w6900_,
		_w6901_
	);
	LUT2 #(
		.INIT('h4)
	) name2855 (
		_w6897_,
		_w6901_,
		_w6902_
	);
	LUT2 #(
		.INIT('h4)
	) name2856 (
		_w6730_,
		_w6902_,
		_w6903_
	);
	LUT2 #(
		.INIT('h2)
	) name2857 (
		_w6730_,
		_w6902_,
		_w6904_
	);
	LUT2 #(
		.INIT('h1)
	) name2858 (
		_w6903_,
		_w6904_,
		_w6905_
	);
	LUT2 #(
		.INIT('h8)
	) name2859 (
		_w6724_,
		_w6905_,
		_w6906_
	);
	LUT2 #(
		.INIT('h1)
	) name2860 (
		_w6597_,
		_w6905_,
		_w6907_
	);
	LUT2 #(
		.INIT('h1)
	) name2861 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6906_,
		_w6908_
	);
	LUT2 #(
		.INIT('h4)
	) name2862 (
		_w6907_,
		_w6908_,
		_w6909_
	);
	LUT2 #(
		.INIT('h1)
	) name2863 (
		_w6593_,
		_w6909_,
		_w6910_
	);
	LUT2 #(
		.INIT('h4)
	) name2864 (
		_w6727_,
		_w6910_,
		_w6911_
	);
	LUT2 #(
		.INIT('h2)
	) name2865 (
		_w6135_,
		_w6911_,
		_w6912_
	);
	LUT2 #(
		.INIT('h2)
	) name2866 (
		_w5066_,
		_w5718_,
		_w6913_
	);
	LUT2 #(
		.INIT('h1)
	) name2867 (
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_DM_2nd_reg/NET0131 ,
		_w6914_
	);
	LUT2 #(
		.INIT('h2)
	) name2868 (
		_w5728_,
		_w5729_,
		_w6915_
	);
	LUT2 #(
		.INIT('h1)
	) name2869 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w6914_,
		_w6916_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		_w6915_,
		_w6916_,
		_w6917_
	);
	LUT2 #(
		.INIT('h8)
	) name2871 (
		_w6913_,
		_w6917_,
		_w6918_
	);
	LUT2 #(
		.INIT('h4)
	) name2872 (
		\bdma_BCTL_reg[1]/NET0131 ,
		\bdma_DM_2nd_reg/NET0131 ,
		_w6919_
	);
	LUT2 #(
		.INIT('h2)
	) name2873 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w6919_,
		_w6920_
	);
	LUT2 #(
		.INIT('h8)
	) name2874 (
		_w6915_,
		_w6920_,
		_w6921_
	);
	LUT2 #(
		.INIT('h8)
	) name2875 (
		_w5066_,
		_w6921_,
		_w6922_
	);
	LUT2 #(
		.INIT('h4)
	) name2876 (
		_w5718_,
		_w6922_,
		_w6923_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		_w6918_,
		_w6923_,
		_w6924_
	);
	LUT2 #(
		.INIT('h8)
	) name2878 (
		\idma_DCTL_reg[14]/NET0131 ,
		_w5068_,
		_w6925_
	);
	LUT2 #(
		.INIT('h4)
	) name2879 (
		_w5717_,
		_w6925_,
		_w6926_
	);
	LUT2 #(
		.INIT('h8)
	) name2880 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w6926_,
		_w6927_
	);
	LUT2 #(
		.INIT('h4)
	) name2881 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		\core_c_psq_PCS_reg[6]/NET0131 ,
		_w6928_
	);
	LUT2 #(
		.INIT('h1)
	) name2882 (
		\core_c_psq_PCS_reg[5]/NET0131 ,
		_w6928_,
		_w6929_
	);
	LUT2 #(
		.INIT('h8)
	) name2883 (
		_w5715_,
		_w6929_,
		_w6930_
	);
	LUT2 #(
		.INIT('h1)
	) name2884 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w4117_,
		_w6931_
	);
	LUT2 #(
		.INIT('h4)
	) name2885 (
		_w4099_,
		_w5946_,
		_w6932_
	);
	LUT2 #(
		.INIT('h8)
	) name2886 (
		_w6931_,
		_w6932_,
		_w6933_
	);
	LUT2 #(
		.INIT('h2)
	) name2887 (
		_w6930_,
		_w6933_,
		_w6934_
	);
	LUT2 #(
		.INIT('h2)
	) name2888 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		_w6934_,
		_w6935_
	);
	LUT2 #(
		.INIT('h8)
	) name2889 (
		\core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 ,
		_w6058_,
		_w6936_
	);
	LUT2 #(
		.INIT('h8)
	) name2890 (
		_w6060_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w6138_,
		_w6938_
	);
	LUT2 #(
		.INIT('h8)
	) name2892 (
		\core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 ,
		_w6140_,
		_w6939_
	);
	LUT2 #(
		.INIT('h8)
	) name2893 (
		\core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 ,
		_w6142_,
		_w6940_
	);
	LUT2 #(
		.INIT('h1)
	) name2894 (
		_w4055_,
		_w6937_,
		_w6941_
	);
	LUT2 #(
		.INIT('h1)
	) name2895 (
		_w6938_,
		_w6939_,
		_w6942_
	);
	LUT2 #(
		.INIT('h4)
	) name2896 (
		_w6940_,
		_w6942_,
		_w6943_
	);
	LUT2 #(
		.INIT('h8)
	) name2897 (
		_w6941_,
		_w6943_,
		_w6944_
	);
	LUT2 #(
		.INIT('h8)
	) name2898 (
		_w6093_,
		_w6936_,
		_w6945_
	);
	LUT2 #(
		.INIT('h8)
	) name2899 (
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w6152_,
		_w6946_
	);
	LUT2 #(
		.INIT('h8)
	) name2900 (
		\core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 ,
		_w6150_,
		_w6947_
	);
	LUT2 #(
		.INIT('h8)
	) name2901 (
		\core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 ,
		_w6154_,
		_w6948_
	);
	LUT2 #(
		.INIT('h1)
	) name2902 (
		_w6945_,
		_w6946_,
		_w6949_
	);
	LUT2 #(
		.INIT('h1)
	) name2903 (
		_w6947_,
		_w6948_,
		_w6950_
	);
	LUT2 #(
		.INIT('h8)
	) name2904 (
		_w6949_,
		_w6950_,
		_w6951_
	);
	LUT2 #(
		.INIT('h8)
	) name2905 (
		_w4055_,
		_w6951_,
		_w6952_
	);
	LUT2 #(
		.INIT('h1)
	) name2906 (
		_w6944_,
		_w6952_,
		_w6953_
	);
	LUT2 #(
		.INIT('h4)
	) name2907 (
		_w6111_,
		_w6953_,
		_w6954_
	);
	LUT2 #(
		.INIT('h8)
	) name2908 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		_w6955_
	);
	LUT2 #(
		.INIT('h4)
	) name2909 (
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w6955_,
		_w6956_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w6956_,
		_w6957_
	);
	LUT2 #(
		.INIT('h8)
	) name2911 (
		_w5964_,
		_w5990_,
		_w6958_
	);
	LUT2 #(
		.INIT('h8)
	) name2912 (
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w6958_,
		_w6959_
	);
	LUT2 #(
		.INIT('h8)
	) name2913 (
		_w6000_,
		_w6002_,
		_w6960_
	);
	LUT2 #(
		.INIT('h8)
	) name2914 (
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w6960_,
		_w6961_
	);
	LUT2 #(
		.INIT('h8)
	) name2915 (
		_w6008_,
		_w6009_,
		_w6962_
	);
	LUT2 #(
		.INIT('h8)
	) name2916 (
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w6962_,
		_w6963_
	);
	LUT2 #(
		.INIT('h8)
	) name2917 (
		_w6015_,
		_w6016_,
		_w6964_
	);
	LUT2 #(
		.INIT('h8)
	) name2918 (
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		_w6964_,
		_w6965_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w6959_,
		_w6961_,
		_w6966_
	);
	LUT2 #(
		.INIT('h1)
	) name2920 (
		_w6963_,
		_w6965_,
		_w6967_
	);
	LUT2 #(
		.INIT('h8)
	) name2921 (
		_w6966_,
		_w6967_,
		_w6968_
	);
	LUT2 #(
		.INIT('h4)
	) name2922 (
		_w4055_,
		_w6968_,
		_w6969_
	);
	LUT2 #(
		.INIT('h8)
	) name2923 (
		_w6015_,
		_w6043_,
		_w6970_
	);
	LUT2 #(
		.INIT('h8)
	) name2924 (
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		_w6970_,
		_w6971_
	);
	LUT2 #(
		.INIT('h8)
	) name2925 (
		_w6000_,
		_w6039_,
		_w6972_
	);
	LUT2 #(
		.INIT('h8)
	) name2926 (
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w6972_,
		_w6973_
	);
	LUT2 #(
		.INIT('h8)
	) name2927 (
		_w6008_,
		_w6041_,
		_w6974_
	);
	LUT2 #(
		.INIT('h8)
	) name2928 (
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w6974_,
		_w6975_
	);
	LUT2 #(
		.INIT('h8)
	) name2929 (
		_w5964_,
		_w6037_,
		_w6976_
	);
	LUT2 #(
		.INIT('h8)
	) name2930 (
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w6976_,
		_w6977_
	);
	LUT2 #(
		.INIT('h1)
	) name2931 (
		_w6971_,
		_w6973_,
		_w6978_
	);
	LUT2 #(
		.INIT('h1)
	) name2932 (
		_w6975_,
		_w6977_,
		_w6979_
	);
	LUT2 #(
		.INIT('h8)
	) name2933 (
		_w6978_,
		_w6979_,
		_w6980_
	);
	LUT2 #(
		.INIT('h8)
	) name2934 (
		_w4055_,
		_w6980_,
		_w6981_
	);
	LUT2 #(
		.INIT('h1)
	) name2935 (
		_w6969_,
		_w6981_,
		_w6982_
	);
	LUT2 #(
		.INIT('h4)
	) name2936 (
		_w6121_,
		_w6982_,
		_w6983_
	);
	LUT2 #(
		.INIT('h1)
	) name2937 (
		_w6954_,
		_w6957_,
		_w6984_
	);
	LUT2 #(
		.INIT('h4)
	) name2938 (
		_w6983_,
		_w6984_,
		_w6985_
	);
	LUT2 #(
		.INIT('h2)
	) name2939 (
		_w5949_,
		_w6985_,
		_w6986_
	);
	LUT2 #(
		.INIT('h4)
	) name2940 (
		\auctl_STEAL_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w6987_
	);
	LUT2 #(
		.INIT('h8)
	) name2941 (
		\memc_STI_Cg_reg/NET0131 ,
		_w6987_,
		_w6988_
	);
	LUT2 #(
		.INIT('h8)
	) name2942 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[0]/NET0131 ,
		_w6988_,
		_w6989_
	);
	LUT2 #(
		.INIT('h1)
	) name2943 (
		_w6927_,
		_w6989_,
		_w6990_
	);
	LUT2 #(
		.INIT('h4)
	) name2944 (
		_w6935_,
		_w6990_,
		_w6991_
	);
	LUT2 #(
		.INIT('h4)
	) name2945 (
		_w6986_,
		_w6991_,
		_w6992_
	);
	LUT2 #(
		.INIT('h2)
	) name2946 (
		_w6924_,
		_w6992_,
		_w6993_
	);
	LUT2 #(
		.INIT('h2)
	) name2947 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w6924_,
		_w6994_
	);
	LUT2 #(
		.INIT('h1)
	) name2948 (
		_w6993_,
		_w6994_,
		_w6995_
	);
	LUT2 #(
		.INIT('h1)
	) name2949 (
		_w6135_,
		_w6995_,
		_w6996_
	);
	LUT2 #(
		.INIT('h1)
	) name2950 (
		_w6176_,
		_w6996_,
		_w6997_
	);
	LUT2 #(
		.INIT('h4)
	) name2951 (
		_w6912_,
		_w6997_,
		_w6998_
	);
	LUT2 #(
		.INIT('h1)
	) name2952 (
		_w6549_,
		_w6998_,
		_w6999_
	);
	LUT2 #(
		.INIT('h4)
	) name2953 (
		_w6106_,
		_w6112_,
		_w7000_
	);
	LUT2 #(
		.INIT('h2)
	) name2954 (
		_w6105_,
		_w7000_,
		_w7001_
	);
	LUT2 #(
		.INIT('h4)
	) name2955 (
		_w6167_,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('h1)
	) name2956 (
		_w5936_,
		_w7002_,
		_w7003_
	);
	LUT2 #(
		.INIT('h8)
	) name2957 (
		_w6049_,
		_w6172_,
		_w7004_
	);
	LUT2 #(
		.INIT('h1)
	) name2958 (
		_w7003_,
		_w7004_,
		_w7005_
	);
	LUT2 #(
		.INIT('h1)
	) name2959 (
		_w6999_,
		_w7005_,
		_w7006_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w6953_,
		_w6982_,
		_w7007_
	);
	LUT2 #(
		.INIT('h2)
	) name2961 (
		_w6135_,
		_w7007_,
		_w7008_
	);
	LUT2 #(
		.INIT('h1)
	) name2962 (
		\memc_DMo_oe1_reg/P0001 ,
		\memc_DMo_oe2_reg/P0001 ,
		_w7009_
	);
	LUT2 #(
		.INIT('h1)
	) name2963 (
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		_w7010_
	);
	LUT2 #(
		.INIT('h1)
	) name2964 (
		\memc_DMo_oe3_reg/P0001 ,
		\memc_DMo_oe6_reg/P0001 ,
		_w7011_
	);
	LUT2 #(
		.INIT('h8)
	) name2965 (
		_w7010_,
		_w7011_,
		_w7012_
	);
	LUT2 #(
		.INIT('h8)
	) name2966 (
		_w7009_,
		_w7012_,
		_w7013_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		\memc_DMo_oe0_reg/P0001 ,
		_w7013_,
		_w7014_
	);
	LUT2 #(
		.INIT('h2)
	) name2968 (
		\memc_DM_oe_reg/P0001 ,
		\memc_DMo_oe7_reg/P0001 ,
		_w7015_
	);
	LUT2 #(
		.INIT('h8)
	) name2969 (
		_w7014_,
		_w7015_,
		_w7016_
	);
	LUT2 #(
		.INIT('h8)
	) name2970 (
		\DM_rdm[13]_pad ,
		_w7016_,
		_w7017_
	);
	LUT2 #(
		.INIT('h1)
	) name2971 (
		\memc_DM_oe_reg/P0001 ,
		\memc_DMo_oe7_reg/P0001 ,
		_w7018_
	);
	LUT2 #(
		.INIT('h4)
	) name2972 (
		\memc_DMo_oe0_reg/P0001 ,
		_w7018_,
		_w7019_
	);
	LUT2 #(
		.INIT('h8)
	) name2973 (
		_w7012_,
		_w7019_,
		_w7020_
	);
	LUT2 #(
		.INIT('h2)
	) name2974 (
		\memc_DMo_oe1_reg/P0001 ,
		\memc_DMo_oe2_reg/P0001 ,
		_w7021_
	);
	LUT2 #(
		.INIT('h8)
	) name2975 (
		_w7020_,
		_w7021_,
		_w7022_
	);
	LUT2 #(
		.INIT('h8)
	) name2976 (
		\DM_rd1[13]_pad ,
		_w7022_,
		_w7023_
	);
	LUT2 #(
		.INIT('h8)
	) name2977 (
		_w7009_,
		_w7019_,
		_w7024_
	);
	LUT2 #(
		.INIT('h4)
	) name2978 (
		\memc_DMo_oe3_reg/P0001 ,
		_w7024_,
		_w7025_
	);
	LUT2 #(
		.INIT('h4)
	) name2979 (
		\memc_DMo_oe6_reg/P0001 ,
		_w7025_,
		_w7026_
	);
	LUT2 #(
		.INIT('h2)
	) name2980 (
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		_w7027_
	);
	LUT2 #(
		.INIT('h8)
	) name2981 (
		_w7026_,
		_w7027_,
		_w7028_
	);
	LUT2 #(
		.INIT('h8)
	) name2982 (
		\DM_rd4[13]_pad ,
		_w7028_,
		_w7029_
	);
	LUT2 #(
		.INIT('h8)
	) name2983 (
		\memc_DMo_oe6_reg/P0001 ,
		_w7010_,
		_w7030_
	);
	LUT2 #(
		.INIT('h8)
	) name2984 (
		_w7025_,
		_w7030_,
		_w7031_
	);
	LUT2 #(
		.INIT('h8)
	) name2985 (
		\DM_rd6[13]_pad ,
		_w7031_,
		_w7032_
	);
	LUT2 #(
		.INIT('h4)
	) name2986 (
		\memc_DM_oe_reg/P0001 ,
		\memc_DMo_oe7_reg/P0001 ,
		_w7033_
	);
	LUT2 #(
		.INIT('h8)
	) name2987 (
		_w7014_,
		_w7033_,
		_w7034_
	);
	LUT2 #(
		.INIT('h8)
	) name2988 (
		\DM_rd7[13]_pad ,
		_w7034_,
		_w7035_
	);
	LUT2 #(
		.INIT('h2)
	) name2989 (
		\memc_DMo_oe3_reg/P0001 ,
		\memc_DMo_oe6_reg/P0001 ,
		_w7036_
	);
	LUT2 #(
		.INIT('h8)
	) name2990 (
		_w7010_,
		_w7036_,
		_w7037_
	);
	LUT2 #(
		.INIT('h8)
	) name2991 (
		_w7024_,
		_w7037_,
		_w7038_
	);
	LUT2 #(
		.INIT('h8)
	) name2992 (
		\DM_rd3[13]_pad ,
		_w7038_,
		_w7039_
	);
	LUT2 #(
		.INIT('h4)
	) name2993 (
		\memc_DMo_oe1_reg/P0001 ,
		\memc_DMo_oe2_reg/P0001 ,
		_w7040_
	);
	LUT2 #(
		.INIT('h8)
	) name2994 (
		_w7020_,
		_w7040_,
		_w7041_
	);
	LUT2 #(
		.INIT('h4)
	) name2995 (
		\memc_DMo_oe4_reg/P0001 ,
		\memc_DMo_oe5_reg/P0001 ,
		_w7042_
	);
	LUT2 #(
		.INIT('h8)
	) name2996 (
		_w7026_,
		_w7042_,
		_w7043_
	);
	LUT2 #(
		.INIT('h1)
	) name2997 (
		_w7022_,
		_w7038_,
		_w7044_
	);
	LUT2 #(
		.INIT('h4)
	) name2998 (
		_w7041_,
		_w7044_,
		_w7045_
	);
	LUT2 #(
		.INIT('h1)
	) name2999 (
		_w7016_,
		_w7031_,
		_w7046_
	);
	LUT2 #(
		.INIT('h4)
	) name3000 (
		_w7034_,
		_w7046_,
		_w7047_
	);
	LUT2 #(
		.INIT('h4)
	) name3001 (
		_w7028_,
		_w7045_,
		_w7048_
	);
	LUT2 #(
		.INIT('h4)
	) name3002 (
		_w7043_,
		_w7048_,
		_w7049_
	);
	LUT2 #(
		.INIT('h8)
	) name3003 (
		_w7047_,
		_w7049_,
		_w7050_
	);
	LUT2 #(
		.INIT('h8)
	) name3004 (
		\memc_DMo_oe0_reg/P0001 ,
		_w7018_,
		_w7051_
	);
	LUT2 #(
		.INIT('h8)
	) name3005 (
		_w7013_,
		_w7051_,
		_w7052_
	);
	LUT2 #(
		.INIT('h1)
	) name3006 (
		_w7050_,
		_w7052_,
		_w7053_
	);
	LUT2 #(
		.INIT('h2)
	) name3007 (
		\DM_rd0[13]_pad ,
		_w7053_,
		_w7054_
	);
	LUT2 #(
		.INIT('h8)
	) name3008 (
		\DM_rd5[13]_pad ,
		_w7043_,
		_w7055_
	);
	LUT2 #(
		.INIT('h8)
	) name3009 (
		\DM_rd2[13]_pad ,
		_w7041_,
		_w7056_
	);
	LUT2 #(
		.INIT('h8)
	) name3010 (
		_w7010_,
		_w7026_,
		_w7057_
	);
	LUT2 #(
		.INIT('h1)
	) name3011 (
		_w7023_,
		_w7039_,
		_w7058_
	);
	LUT2 #(
		.INIT('h4)
	) name3012 (
		_w7056_,
		_w7058_,
		_w7059_
	);
	LUT2 #(
		.INIT('h1)
	) name3013 (
		_w7017_,
		_w7032_,
		_w7060_
	);
	LUT2 #(
		.INIT('h1)
	) name3014 (
		_w7035_,
		_w7057_,
		_w7061_
	);
	LUT2 #(
		.INIT('h8)
	) name3015 (
		_w7060_,
		_w7061_,
		_w7062_
	);
	LUT2 #(
		.INIT('h4)
	) name3016 (
		_w7029_,
		_w7059_,
		_w7063_
	);
	LUT2 #(
		.INIT('h4)
	) name3017 (
		_w7055_,
		_w7063_,
		_w7064_
	);
	LUT2 #(
		.INIT('h8)
	) name3018 (
		_w7062_,
		_w7064_,
		_w7065_
	);
	LUT2 #(
		.INIT('h4)
	) name3019 (
		_w7054_,
		_w7065_,
		_w7066_
	);
	LUT2 #(
		.INIT('h8)
	) name3020 (
		\regout_STD_C_reg[13]/P0001 ,
		_w6988_,
		_w7067_
	);
	LUT2 #(
		.INIT('h2)
	) name3021 (
		\core_c_dec_MFDAG1_Ei_reg/NET0131 ,
		_w6988_,
		_w7068_
	);
	LUT2 #(
		.INIT('h8)
	) name3022 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131 ,
		_w7069_
	);
	LUT2 #(
		.INIT('h8)
	) name3023 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[13]/NET0131 ,
		_w7070_
	);
	LUT2 #(
		.INIT('h8)
	) name3024 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w7071_
	);
	LUT2 #(
		.INIT('h8)
	) name3025 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131 ,
		_w7072_
	);
	LUT2 #(
		.INIT('h8)
	) name3026 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131 ,
		_w7073_
	);
	LUT2 #(
		.INIT('h8)
	) name3027 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131 ,
		_w7074_
	);
	LUT2 #(
		.INIT('h8)
	) name3028 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131 ,
		_w7075_
	);
	LUT2 #(
		.INIT('h1)
	) name3029 (
		_w7072_,
		_w7073_,
		_w7076_
	);
	LUT2 #(
		.INIT('h1)
	) name3030 (
		_w7074_,
		_w7075_,
		_w7077_
	);
	LUT2 #(
		.INIT('h8)
	) name3031 (
		_w7076_,
		_w7077_,
		_w7078_
	);
	LUT2 #(
		.INIT('h8)
	) name3032 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131 ,
		_w7079_
	);
	LUT2 #(
		.INIT('h8)
	) name3033 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131 ,
		_w7080_
	);
	LUT2 #(
		.INIT('h8)
	) name3034 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w7081_
	);
	LUT2 #(
		.INIT('h8)
	) name3035 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		_w7082_
	);
	LUT2 #(
		.INIT('h8)
	) name3036 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131 ,
		_w7083_
	);
	LUT2 #(
		.INIT('h1)
	) name3037 (
		_w7069_,
		_w7070_,
		_w7084_
	);
	LUT2 #(
		.INIT('h1)
	) name3038 (
		_w7071_,
		_w7079_,
		_w7085_
	);
	LUT2 #(
		.INIT('h1)
	) name3039 (
		_w7080_,
		_w7081_,
		_w7086_
	);
	LUT2 #(
		.INIT('h1)
	) name3040 (
		_w7082_,
		_w7083_,
		_w7087_
	);
	LUT2 #(
		.INIT('h8)
	) name3041 (
		_w7086_,
		_w7087_,
		_w7088_
	);
	LUT2 #(
		.INIT('h8)
	) name3042 (
		_w7084_,
		_w7085_,
		_w7089_
	);
	LUT2 #(
		.INIT('h8)
	) name3043 (
		_w7088_,
		_w7089_,
		_w7090_
	);
	LUT2 #(
		.INIT('h8)
	) name3044 (
		_w7078_,
		_w7090_,
		_w7091_
	);
	LUT2 #(
		.INIT('h2)
	) name3045 (
		_w7068_,
		_w7091_,
		_w7092_
	);
	LUT2 #(
		.INIT('h2)
	) name3046 (
		\core_c_dec_MFALU_Ei_reg/NET0131 ,
		_w6988_,
		_w7093_
	);
	LUT2 #(
		.INIT('h4)
	) name3047 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001 ,
		_w7094_
	);
	LUT2 #(
		.INIT('h8)
	) name3048 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001 ,
		_w7095_
	);
	LUT2 #(
		.INIT('h1)
	) name3049 (
		_w7094_,
		_w7095_,
		_w7096_
	);
	LUT2 #(
		.INIT('h2)
	) name3050 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w7096_,
		_w7097_
	);
	LUT2 #(
		.INIT('h4)
	) name3051 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001 ,
		_w7098_
	);
	LUT2 #(
		.INIT('h8)
	) name3052 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001 ,
		_w7099_
	);
	LUT2 #(
		.INIT('h1)
	) name3053 (
		_w7098_,
		_w7099_,
		_w7100_
	);
	LUT2 #(
		.INIT('h2)
	) name3054 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w7100_,
		_w7101_
	);
	LUT2 #(
		.INIT('h4)
	) name3055 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001 ,
		_w7102_
	);
	LUT2 #(
		.INIT('h8)
	) name3056 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001 ,
		_w7103_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w7102_,
		_w7103_,
		_w7104_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w7104_,
		_w7105_
	);
	LUT2 #(
		.INIT('h4)
	) name3059 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001 ,
		_w7106_
	);
	LUT2 #(
		.INIT('h8)
	) name3060 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001 ,
		_w7107_
	);
	LUT2 #(
		.INIT('h1)
	) name3061 (
		_w7106_,
		_w7107_,
		_w7108_
	);
	LUT2 #(
		.INIT('h2)
	) name3062 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w7108_,
		_w7109_
	);
	LUT2 #(
		.INIT('h4)
	) name3063 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001 ,
		_w7110_
	);
	LUT2 #(
		.INIT('h8)
	) name3064 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001 ,
		_w7111_
	);
	LUT2 #(
		.INIT('h1)
	) name3065 (
		_w7110_,
		_w7111_,
		_w7112_
	);
	LUT2 #(
		.INIT('h2)
	) name3066 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w7112_,
		_w7113_
	);
	LUT2 #(
		.INIT('h1)
	) name3067 (
		_w7097_,
		_w7101_,
		_w7114_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		_w7105_,
		_w7109_,
		_w7115_
	);
	LUT2 #(
		.INIT('h4)
	) name3069 (
		_w7113_,
		_w7115_,
		_w7116_
	);
	LUT2 #(
		.INIT('h8)
	) name3070 (
		_w7114_,
		_w7116_,
		_w7117_
	);
	LUT2 #(
		.INIT('h2)
	) name3071 (
		_w7093_,
		_w7117_,
		_w7118_
	);
	LUT2 #(
		.INIT('h2)
	) name3072 (
		\core_c_dec_MFSPT_Ei_reg/NET0131 ,
		_w6988_,
		_w7119_
	);
	LUT2 #(
		.INIT('h8)
	) name3073 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[13]/P0001 ,
		_w7120_
	);
	LUT2 #(
		.INIT('h8)
	) name3074 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[13]/P0001 ,
		_w7121_
	);
	LUT2 #(
		.INIT('h8)
	) name3075 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[13]/P0001 ,
		_w7122_
	);
	LUT2 #(
		.INIT('h8)
	) name3076 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[13]/P0001 ,
		_w7123_
	);
	LUT2 #(
		.INIT('h1)
	) name3077 (
		_w7120_,
		_w7121_,
		_w7124_
	);
	LUT2 #(
		.INIT('h1)
	) name3078 (
		_w7122_,
		_w7123_,
		_w7125_
	);
	LUT2 #(
		.INIT('h8)
	) name3079 (
		_w7124_,
		_w7125_,
		_w7126_
	);
	LUT2 #(
		.INIT('h2)
	) name3080 (
		_w7119_,
		_w7126_,
		_w7127_
	);
	LUT2 #(
		.INIT('h2)
	) name3081 (
		\core_c_dec_MFDAG2_Ei_reg/NET0131 ,
		_w6988_,
		_w7128_
	);
	LUT2 #(
		.INIT('h8)
	) name3082 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131 ,
		_w7129_
	);
	LUT2 #(
		.INIT('h8)
	) name3083 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w7130_
	);
	LUT2 #(
		.INIT('h8)
	) name3084 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131 ,
		_w7131_
	);
	LUT2 #(
		.INIT('h8)
	) name3085 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131 ,
		_w7132_
	);
	LUT2 #(
		.INIT('h8)
	) name3086 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131 ,
		_w7133_
	);
	LUT2 #(
		.INIT('h8)
	) name3087 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131 ,
		_w7134_
	);
	LUT2 #(
		.INIT('h1)
	) name3088 (
		_w7131_,
		_w7132_,
		_w7135_
	);
	LUT2 #(
		.INIT('h1)
	) name3089 (
		_w7133_,
		_w7134_,
		_w7136_
	);
	LUT2 #(
		.INIT('h8)
	) name3090 (
		_w7135_,
		_w7136_,
		_w7137_
	);
	LUT2 #(
		.INIT('h8)
	) name3091 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131 ,
		_w7138_
	);
	LUT2 #(
		.INIT('h8)
	) name3092 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w7139_
	);
	LUT2 #(
		.INIT('h8)
	) name3093 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		_w7140_
	);
	LUT2 #(
		.INIT('h8)
	) name3094 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131 ,
		_w7141_
	);
	LUT2 #(
		.INIT('h8)
	) name3095 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w7142_
	);
	LUT2 #(
		.INIT('h8)
	) name3096 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131 ,
		_w7143_
	);
	LUT2 #(
		.INIT('h1)
	) name3097 (
		_w7129_,
		_w7130_,
		_w7144_
	);
	LUT2 #(
		.INIT('h1)
	) name3098 (
		_w7138_,
		_w7139_,
		_w7145_
	);
	LUT2 #(
		.INIT('h1)
	) name3099 (
		_w7140_,
		_w7141_,
		_w7146_
	);
	LUT2 #(
		.INIT('h1)
	) name3100 (
		_w7142_,
		_w7143_,
		_w7147_
	);
	LUT2 #(
		.INIT('h8)
	) name3101 (
		_w7146_,
		_w7147_,
		_w7148_
	);
	LUT2 #(
		.INIT('h8)
	) name3102 (
		_w7144_,
		_w7145_,
		_w7149_
	);
	LUT2 #(
		.INIT('h8)
	) name3103 (
		_w7148_,
		_w7149_,
		_w7150_
	);
	LUT2 #(
		.INIT('h8)
	) name3104 (
		_w7137_,
		_w7150_,
		_w7151_
	);
	LUT2 #(
		.INIT('h2)
	) name3105 (
		_w7128_,
		_w7151_,
		_w7152_
	);
	LUT2 #(
		.INIT('h2)
	) name3106 (
		\core_c_dec_MFSHT_Ei_reg/NET0131 ,
		_w6988_,
		_w7153_
	);
	LUT2 #(
		.INIT('h4)
	) name3107 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 ,
		_w7154_
	);
	LUT2 #(
		.INIT('h8)
	) name3108 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 ,
		_w7155_
	);
	LUT2 #(
		.INIT('h1)
	) name3109 (
		_w7154_,
		_w7155_,
		_w7156_
	);
	LUT2 #(
		.INIT('h2)
	) name3110 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w7156_,
		_w7157_
	);
	LUT2 #(
		.INIT('h4)
	) name3111 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001 ,
		_w7158_
	);
	LUT2 #(
		.INIT('h8)
	) name3112 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001 ,
		_w7159_
	);
	LUT2 #(
		.INIT('h1)
	) name3113 (
		_w7158_,
		_w7159_,
		_w7160_
	);
	LUT2 #(
		.INIT('h2)
	) name3114 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w7160_,
		_w7161_
	);
	LUT2 #(
		.INIT('h4)
	) name3115 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 ,
		_w7162_
	);
	LUT2 #(
		.INIT('h8)
	) name3116 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 ,
		_w7163_
	);
	LUT2 #(
		.INIT('h1)
	) name3117 (
		_w7162_,
		_w7163_,
		_w7164_
	);
	LUT2 #(
		.INIT('h2)
	) name3118 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w7164_,
		_w7165_
	);
	LUT2 #(
		.INIT('h4)
	) name3119 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[4]/P0001 ,
		_w7166_
	);
	LUT2 #(
		.INIT('h8)
	) name3120 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBs_reg[4]/P0001 ,
		_w7167_
	);
	LUT2 #(
		.INIT('h1)
	) name3121 (
		_w7166_,
		_w7167_,
		_w7168_
	);
	LUT2 #(
		.INIT('h2)
	) name3122 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		_w7168_,
		_w7169_
	);
	LUT2 #(
		.INIT('h4)
	) name3123 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001 ,
		_w7170_
	);
	LUT2 #(
		.INIT('h8)
	) name3124 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001 ,
		_w7171_
	);
	LUT2 #(
		.INIT('h1)
	) name3125 (
		_w7170_,
		_w7171_,
		_w7172_
	);
	LUT2 #(
		.INIT('h2)
	) name3126 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w7172_,
		_w7173_
	);
	LUT2 #(
		.INIT('h1)
	) name3127 (
		_w7169_,
		_w7173_,
		_w7174_
	);
	LUT2 #(
		.INIT('h1)
	) name3128 (
		_w7157_,
		_w7161_,
		_w7175_
	);
	LUT2 #(
		.INIT('h4)
	) name3129 (
		_w7165_,
		_w7175_,
		_w7176_
	);
	LUT2 #(
		.INIT('h8)
	) name3130 (
		_w7174_,
		_w7176_,
		_w7177_
	);
	LUT2 #(
		.INIT('h2)
	) name3131 (
		_w7153_,
		_w7177_,
		_w7178_
	);
	LUT2 #(
		.INIT('h2)
	) name3132 (
		\core_c_dec_MFMAC_Ei_reg/NET0131 ,
		_w6988_,
		_w7179_
	);
	LUT2 #(
		.INIT('h4)
	) name3133 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001 ,
		_w7180_
	);
	LUT2 #(
		.INIT('h8)
	) name3134 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 ,
		_w7181_
	);
	LUT2 #(
		.INIT('h1)
	) name3135 (
		_w7180_,
		_w7181_,
		_w7182_
	);
	LUT2 #(
		.INIT('h2)
	) name3136 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w7182_,
		_w7183_
	);
	LUT2 #(
		.INIT('h4)
	) name3137 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001 ,
		_w7184_
	);
	LUT2 #(
		.INIT('h8)
	) name3138 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001 ,
		_w7185_
	);
	LUT2 #(
		.INIT('h1)
	) name3139 (
		_w7184_,
		_w7185_,
		_w7186_
	);
	LUT2 #(
		.INIT('h2)
	) name3140 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h4)
	) name3141 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001 ,
		_w7188_
	);
	LUT2 #(
		.INIT('h8)
	) name3142 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001 ,
		_w7189_
	);
	LUT2 #(
		.INIT('h1)
	) name3143 (
		_w7188_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h2)
	) name3144 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w7190_,
		_w7191_
	);
	LUT2 #(
		.INIT('h4)
	) name3145 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001 ,
		_w7192_
	);
	LUT2 #(
		.INIT('h8)
	) name3146 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001 ,
		_w7193_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w7192_,
		_w7193_,
		_w7194_
	);
	LUT2 #(
		.INIT('h2)
	) name3148 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w7194_,
		_w7195_
	);
	LUT2 #(
		.INIT('h4)
	) name3149 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001 ,
		_w7196_
	);
	LUT2 #(
		.INIT('h8)
	) name3150 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001 ,
		_w7197_
	);
	LUT2 #(
		.INIT('h1)
	) name3151 (
		_w7196_,
		_w7197_,
		_w7198_
	);
	LUT2 #(
		.INIT('h2)
	) name3152 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w7198_,
		_w7199_
	);
	LUT2 #(
		.INIT('h4)
	) name3153 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001 ,
		_w7200_
	);
	LUT2 #(
		.INIT('h8)
	) name3154 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 ,
		_w7201_
	);
	LUT2 #(
		.INIT('h1)
	) name3155 (
		_w7200_,
		_w7201_,
		_w7202_
	);
	LUT2 #(
		.INIT('h2)
	) name3156 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w7202_,
		_w7203_
	);
	LUT2 #(
		.INIT('h4)
	) name3157 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		_w7204_
	);
	LUT2 #(
		.INIT('h8)
	) name3158 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w7205_
	);
	LUT2 #(
		.INIT('h1)
	) name3159 (
		_w7204_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('h2)
	) name3160 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w7206_,
		_w7207_
	);
	LUT2 #(
		.INIT('h1)
	) name3161 (
		_w7183_,
		_w7187_,
		_w7208_
	);
	LUT2 #(
		.INIT('h1)
	) name3162 (
		_w7191_,
		_w7195_,
		_w7209_
	);
	LUT2 #(
		.INIT('h1)
	) name3163 (
		_w7199_,
		_w7203_,
		_w7210_
	);
	LUT2 #(
		.INIT('h4)
	) name3164 (
		_w7207_,
		_w7210_,
		_w7211_
	);
	LUT2 #(
		.INIT('h8)
	) name3165 (
		_w7208_,
		_w7209_,
		_w7212_
	);
	LUT2 #(
		.INIT('h8)
	) name3166 (
		_w7211_,
		_w7212_,
		_w7213_
	);
	LUT2 #(
		.INIT('h2)
	) name3167 (
		_w7179_,
		_w7213_,
		_w7214_
	);
	LUT2 #(
		.INIT('h2)
	) name3168 (
		\core_c_dec_MFPSQ_Ei_reg/NET0131 ,
		_w6988_,
		_w7215_
	);
	LUT2 #(
		.INIT('h1)
	) name3169 (
		\core_c_dec_imm14_E_reg/P0001 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w7216_
	);
	LUT2 #(
		.INIT('h2)
	) name3170 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w7216_,
		_w7217_
	);
	LUT2 #(
		.INIT('h8)
	) name3171 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w7218_
	);
	LUT2 #(
		.INIT('h8)
	) name3172 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w7219_
	);
	LUT2 #(
		.INIT('h2)
	) name3173 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4489_,
		_w7220_
	);
	LUT2 #(
		.INIT('h1)
	) name3174 (
		_w7218_,
		_w7219_,
		_w7221_
	);
	LUT2 #(
		.INIT('h4)
	) name3175 (
		_w7217_,
		_w7221_,
		_w7222_
	);
	LUT2 #(
		.INIT('h4)
	) name3176 (
		_w7220_,
		_w7222_,
		_w7223_
	);
	LUT2 #(
		.INIT('h2)
	) name3177 (
		_w7215_,
		_w7223_,
		_w7224_
	);
	LUT2 #(
		.INIT('h4)
	) name3178 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w7225_
	);
	LUT2 #(
		.INIT('h8)
	) name3179 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w7226_
	);
	LUT2 #(
		.INIT('h8)
	) name3180 (
		_w7225_,
		_w7226_,
		_w7227_
	);
	LUT2 #(
		.INIT('h1)
	) name3181 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w7228_
	);
	LUT2 #(
		.INIT('h8)
	) name3182 (
		_w5944_,
		_w7228_,
		_w7229_
	);
	LUT2 #(
		.INIT('h8)
	) name3183 (
		_w7227_,
		_w7229_,
		_w7230_
	);
	LUT2 #(
		.INIT('h8)
	) name3184 (
		\bdma_BCTL_reg[13]/NET0131 ,
		_w7230_,
		_w7231_
	);
	LUT2 #(
		.INIT('h2)
	) name3185 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w7232_
	);
	LUT2 #(
		.INIT('h8)
	) name3186 (
		_w7225_,
		_w7232_,
		_w7233_
	);
	LUT2 #(
		.INIT('h8)
	) name3187 (
		_w7229_,
		_w7233_,
		_w7234_
	);
	LUT2 #(
		.INIT('h8)
	) name3188 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w7234_,
		_w7235_
	);
	LUT2 #(
		.INIT('h8)
	) name3189 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w7236_
	);
	LUT2 #(
		.INIT('h4)
	) name3190 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w7237_
	);
	LUT2 #(
		.INIT('h8)
	) name3191 (
		_w7225_,
		_w7237_,
		_w7238_
	);
	LUT2 #(
		.INIT('h8)
	) name3192 (
		_w7236_,
		_w7238_,
		_w7239_
	);
	LUT2 #(
		.INIT('h8)
	) name3193 (
		\clkc_ckr_reg_DO_reg[13]/NET0131 ,
		_w7239_,
		_w7240_
	);
	LUT2 #(
		.INIT('h8)
	) name3194 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		_w7241_
	);
	LUT2 #(
		.INIT('h4)
	) name3195 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w7242_
	);
	LUT2 #(
		.INIT('h8)
	) name3196 (
		_w7241_,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h8)
	) name3197 (
		_w7228_,
		_w7243_,
		_w7244_
	);
	LUT2 #(
		.INIT('h8)
	) name3198 (
		\PIO_oe[9]_pad ,
		_w7244_,
		_w7245_
	);
	LUT2 #(
		.INIT('h4)
	) name3199 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w7246_
	);
	LUT2 #(
		.INIT('h8)
	) name3200 (
		_w7233_,
		_w7246_,
		_w7247_
	);
	LUT2 #(
		.INIT('h8)
	) name3201 (
		\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w7247_,
		_w7248_
	);
	LUT2 #(
		.INIT('h8)
	) name3202 (
		_w7243_,
		_w7246_,
		_w7249_
	);
	LUT2 #(
		.INIT('h8)
	) name3203 (
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w7249_,
		_w7250_
	);
	LUT2 #(
		.INIT('h8)
	) name3204 (
		_w7236_,
		_w7243_,
		_w7251_
	);
	LUT2 #(
		.INIT('h8)
	) name3205 (
		\emc_WSCRreg_DO_reg[13]/NET0131 ,
		_w7251_,
		_w7252_
	);
	LUT2 #(
		.INIT('h8)
	) name3206 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w7253_
	);
	LUT2 #(
		.INIT('h4)
	) name3207 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		_w7254_
	);
	LUT2 #(
		.INIT('h8)
	) name3208 (
		_w7253_,
		_w7254_,
		_w7255_
	);
	LUT2 #(
		.INIT('h8)
	) name3209 (
		_w7246_,
		_w7255_,
		_w7256_
	);
	LUT2 #(
		.INIT('h8)
	) name3210 (
		\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w7256_,
		_w7257_
	);
	LUT2 #(
		.INIT('h8)
	) name3211 (
		_w7242_,
		_w7254_,
		_w7258_
	);
	LUT2 #(
		.INIT('h8)
	) name3212 (
		_w7246_,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('h8)
	) name3213 (
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w7259_,
		_w7260_
	);
	LUT2 #(
		.INIT('h1)
	) name3214 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w7261_
	);
	LUT2 #(
		.INIT('h8)
	) name3215 (
		_w7225_,
		_w7261_,
		_w7262_
	);
	LUT2 #(
		.INIT('h8)
	) name3216 (
		_w7236_,
		_w7262_,
		_w7263_
	);
	LUT2 #(
		.INIT('h1)
	) name3217 (
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w7264_
	);
	LUT2 #(
		.INIT('h2)
	) name3218 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport1_rxctl_SLOT1_EXT_reg[3]/NET0131 ,
		_w7265_
	);
	LUT2 #(
		.INIT('h1)
	) name3219 (
		_w7264_,
		_w7265_,
		_w7266_
	);
	LUT2 #(
		.INIT('h8)
	) name3220 (
		_w7263_,
		_w7266_,
		_w7267_
	);
	LUT2 #(
		.INIT('h4)
	) name3221 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w7268_
	);
	LUT2 #(
		.INIT('h4)
	) name3222 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w7269_
	);
	LUT2 #(
		.INIT('h8)
	) name3223 (
		_w7261_,
		_w7269_,
		_w7270_
	);
	LUT2 #(
		.INIT('h8)
	) name3224 (
		_w7268_,
		_w7270_,
		_w7271_
	);
	LUT2 #(
		.INIT('h8)
	) name3225 (
		\pio_PINT_reg[9]/NET0131 ,
		_w7271_,
		_w7272_
	);
	LUT2 #(
		.INIT('h8)
	) name3226 (
		_w7246_,
		_w7262_,
		_w7273_
	);
	LUT2 #(
		.INIT('h8)
	) name3227 (
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w7273_,
		_w7274_
	);
	LUT2 #(
		.INIT('h8)
	) name3228 (
		_w7241_,
		_w7253_,
		_w7275_
	);
	LUT2 #(
		.INIT('h8)
	) name3229 (
		_w7246_,
		_w7275_,
		_w7276_
	);
	LUT2 #(
		.INIT('h1)
	) name3230 (
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w7277_
	);
	LUT2 #(
		.INIT('h2)
	) name3231 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		\sport0_rxctl_SLOT1_EXT_reg[3]/NET0131 ,
		_w7278_
	);
	LUT2 #(
		.INIT('h1)
	) name3232 (
		_w7277_,
		_w7278_,
		_w7279_
	);
	LUT2 #(
		.INIT('h8)
	) name3233 (
		_w7276_,
		_w7279_,
		_w7280_
	);
	LUT2 #(
		.INIT('h8)
	) name3234 (
		_w7238_,
		_w7246_,
		_w7281_
	);
	LUT2 #(
		.INIT('h8)
	) name3235 (
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w7281_,
		_w7282_
	);
	LUT2 #(
		.INIT('h2)
	) name3236 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w7283_
	);
	LUT2 #(
		.INIT('h8)
	) name3237 (
		_w7261_,
		_w7283_,
		_w7284_
	);
	LUT2 #(
		.INIT('h4)
	) name3238 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5944_,
		_w7285_
	);
	LUT2 #(
		.INIT('h8)
	) name3239 (
		\memc_selMIO_E_reg/P0001 ,
		_w7285_,
		_w7286_
	);
	LUT2 #(
		.INIT('h8)
	) name3240 (
		_w7284_,
		_w7286_,
		_w7287_
	);
	LUT2 #(
		.INIT('h8)
	) name3241 (
		\bdma_BWCOUNT_reg[13]/NET0131 ,
		_w7287_,
		_w7288_
	);
	LUT2 #(
		.INIT('h8)
	) name3242 (
		_w7236_,
		_w7258_,
		_w7289_
	);
	LUT2 #(
		.INIT('h8)
	) name3243 (
		\tm_TCR_TMP_reg[13]/NET0131 ,
		_w7289_,
		_w7290_
	);
	LUT2 #(
		.INIT('h8)
	) name3244 (
		_w7228_,
		_w7255_,
		_w7291_
	);
	LUT2 #(
		.INIT('h8)
	) name3245 (
		\PIO_out[9]_pad ,
		_w7291_,
		_w7292_
	);
	LUT2 #(
		.INIT('h8)
	) name3246 (
		_w7236_,
		_w7255_,
		_w7293_
	);
	LUT2 #(
		.INIT('h8)
	) name3247 (
		\tm_tpr_reg_DO_reg[13]/NET0131 ,
		_w7293_,
		_w7294_
	);
	LUT2 #(
		.INIT('h8)
	) name3248 (
		_w7227_,
		_w7246_,
		_w7295_
	);
	LUT2 #(
		.INIT('h8)
	) name3249 (
		\sport0_regs_AUTO_a_reg[13]/NET0131 ,
		_w7295_,
		_w7296_
	);
	LUT2 #(
		.INIT('h8)
	) name3250 (
		_w7228_,
		_w7275_,
		_w7297_
	);
	LUT2 #(
		.INIT('h8)
	) name3251 (
		\pio_pmask_reg_DO_reg[9]/NET0131 ,
		_w7297_,
		_w7298_
	);
	LUT2 #(
		.INIT('h8)
	) name3252 (
		_w7228_,
		_w7262_,
		_w7299_
	);
	LUT2 #(
		.INIT('h8)
	) name3253 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w7299_,
		_w7300_
	);
	LUT2 #(
		.INIT('h8)
	) name3254 (
		_w7236_,
		_w7275_,
		_w7301_
	);
	LUT2 #(
		.INIT('h8)
	) name3255 (
		\memc_usysr_DO_reg[13]/NET0131 ,
		_w7301_,
		_w7302_
	);
	LUT2 #(
		.INIT('h8)
	) name3256 (
		_w7229_,
		_w7238_,
		_w7303_
	);
	LUT2 #(
		.INIT('h8)
	) name3257 (
		\bdma_BEAD_reg[13]/NET0131 ,
		_w7303_,
		_w7304_
	);
	LUT2 #(
		.INIT('h1)
	) name3258 (
		_w7240_,
		_w7245_,
		_w7305_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w7248_,
		_w7250_,
		_w7306_
	);
	LUT2 #(
		.INIT('h1)
	) name3260 (
		_w7252_,
		_w7257_,
		_w7307_
	);
	LUT2 #(
		.INIT('h1)
	) name3261 (
		_w7260_,
		_w7267_,
		_w7308_
	);
	LUT2 #(
		.INIT('h1)
	) name3262 (
		_w7272_,
		_w7274_,
		_w7309_
	);
	LUT2 #(
		.INIT('h1)
	) name3263 (
		_w7280_,
		_w7282_,
		_w7310_
	);
	LUT2 #(
		.INIT('h1)
	) name3264 (
		_w7290_,
		_w7292_,
		_w7311_
	);
	LUT2 #(
		.INIT('h1)
	) name3265 (
		_w7294_,
		_w7296_,
		_w7312_
	);
	LUT2 #(
		.INIT('h1)
	) name3266 (
		_w7298_,
		_w7300_,
		_w7313_
	);
	LUT2 #(
		.INIT('h4)
	) name3267 (
		_w7302_,
		_w7313_,
		_w7314_
	);
	LUT2 #(
		.INIT('h8)
	) name3268 (
		_w7311_,
		_w7312_,
		_w7315_
	);
	LUT2 #(
		.INIT('h8)
	) name3269 (
		_w7309_,
		_w7310_,
		_w7316_
	);
	LUT2 #(
		.INIT('h8)
	) name3270 (
		_w7307_,
		_w7308_,
		_w7317_
	);
	LUT2 #(
		.INIT('h8)
	) name3271 (
		_w7305_,
		_w7306_,
		_w7318_
	);
	LUT2 #(
		.INIT('h8)
	) name3272 (
		_w7317_,
		_w7318_,
		_w7319_
	);
	LUT2 #(
		.INIT('h8)
	) name3273 (
		_w7315_,
		_w7316_,
		_w7320_
	);
	LUT2 #(
		.INIT('h8)
	) name3274 (
		_w7314_,
		_w7320_,
		_w7321_
	);
	LUT2 #(
		.INIT('h4)
	) name3275 (
		_w7231_,
		_w7319_,
		_w7322_
	);
	LUT2 #(
		.INIT('h1)
	) name3276 (
		_w7235_,
		_w7304_,
		_w7323_
	);
	LUT2 #(
		.INIT('h8)
	) name3277 (
		_w7322_,
		_w7323_,
		_w7324_
	);
	LUT2 #(
		.INIT('h4)
	) name3278 (
		_w7288_,
		_w7321_,
		_w7325_
	);
	LUT2 #(
		.INIT('h8)
	) name3279 (
		_w7324_,
		_w7325_,
		_w7326_
	);
	LUT2 #(
		.INIT('h2)
	) name3280 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7326_,
		_w7327_
	);
	LUT2 #(
		.INIT('h1)
	) name3281 (
		_w7092_,
		_w7127_,
		_w7328_
	);
	LUT2 #(
		.INIT('h4)
	) name3282 (
		_w7152_,
		_w7328_,
		_w7329_
	);
	LUT2 #(
		.INIT('h1)
	) name3283 (
		_w7118_,
		_w7178_,
		_w7330_
	);
	LUT2 #(
		.INIT('h4)
	) name3284 (
		_w7214_,
		_w7330_,
		_w7331_
	);
	LUT2 #(
		.INIT('h8)
	) name3285 (
		_w7329_,
		_w7331_,
		_w7332_
	);
	LUT2 #(
		.INIT('h4)
	) name3286 (
		_w7224_,
		_w7332_,
		_w7333_
	);
	LUT2 #(
		.INIT('h4)
	) name3287 (
		_w7327_,
		_w7333_,
		_w7334_
	);
	LUT2 #(
		.INIT('h4)
	) name3288 (
		_w7067_,
		_w7334_,
		_w7335_
	);
	LUT2 #(
		.INIT('h1)
	) name3289 (
		\emc_DMDoe_reg/NET0131 ,
		_w7335_,
		_w7336_
	);
	LUT2 #(
		.INIT('h8)
	) name3290 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[13]/P0001 ,
		_w7337_
	);
	LUT2 #(
		.INIT('h2)
	) name3291 (
		_w7057_,
		_w7337_,
		_w7338_
	);
	LUT2 #(
		.INIT('h4)
	) name3292 (
		_w7336_,
		_w7338_,
		_w7339_
	);
	LUT2 #(
		.INIT('h1)
	) name3293 (
		_w7066_,
		_w7339_,
		_w7340_
	);
	LUT2 #(
		.INIT('h4)
	) name3294 (
		_w6135_,
		_w7340_,
		_w7341_
	);
	LUT2 #(
		.INIT('h1)
	) name3295 (
		_w6176_,
		_w7008_,
		_w7342_
	);
	LUT2 #(
		.INIT('h4)
	) name3296 (
		_w7341_,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h8)
	) name3297 (
		\DM_rdm[0]_pad ,
		_w7016_,
		_w7344_
	);
	LUT2 #(
		.INIT('h8)
	) name3298 (
		\DM_rd1[0]_pad ,
		_w7022_,
		_w7345_
	);
	LUT2 #(
		.INIT('h8)
	) name3299 (
		\DM_rd5[0]_pad ,
		_w7043_,
		_w7346_
	);
	LUT2 #(
		.INIT('h8)
	) name3300 (
		\DM_rd6[0]_pad ,
		_w7031_,
		_w7347_
	);
	LUT2 #(
		.INIT('h8)
	) name3301 (
		\DM_rd7[0]_pad ,
		_w7034_,
		_w7348_
	);
	LUT2 #(
		.INIT('h8)
	) name3302 (
		\DM_rd3[0]_pad ,
		_w7038_,
		_w7349_
	);
	LUT2 #(
		.INIT('h2)
	) name3303 (
		\DM_rd0[0]_pad ,
		_w7053_,
		_w7350_
	);
	LUT2 #(
		.INIT('h8)
	) name3304 (
		\DM_rd4[0]_pad ,
		_w7028_,
		_w7351_
	);
	LUT2 #(
		.INIT('h8)
	) name3305 (
		\DM_rd2[0]_pad ,
		_w7041_,
		_w7352_
	);
	LUT2 #(
		.INIT('h1)
	) name3306 (
		_w7345_,
		_w7349_,
		_w7353_
	);
	LUT2 #(
		.INIT('h4)
	) name3307 (
		_w7352_,
		_w7353_,
		_w7354_
	);
	LUT2 #(
		.INIT('h1)
	) name3308 (
		_w7057_,
		_w7344_,
		_w7355_
	);
	LUT2 #(
		.INIT('h1)
	) name3309 (
		_w7347_,
		_w7348_,
		_w7356_
	);
	LUT2 #(
		.INIT('h8)
	) name3310 (
		_w7355_,
		_w7356_,
		_w7357_
	);
	LUT2 #(
		.INIT('h4)
	) name3311 (
		_w7346_,
		_w7354_,
		_w7358_
	);
	LUT2 #(
		.INIT('h4)
	) name3312 (
		_w7351_,
		_w7358_,
		_w7359_
	);
	LUT2 #(
		.INIT('h8)
	) name3313 (
		_w7357_,
		_w7359_,
		_w7360_
	);
	LUT2 #(
		.INIT('h4)
	) name3314 (
		_w7350_,
		_w7360_,
		_w7361_
	);
	LUT2 #(
		.INIT('h8)
	) name3315 (
		\regout_STD_C_reg[0]/P0001 ,
		_w6988_,
		_w7362_
	);
	LUT2 #(
		.INIT('h4)
	) name3316 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[0]/P0001 ,
		_w7363_
	);
	LUT2 #(
		.INIT('h8)
	) name3317 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBs_reg[0]/P0001 ,
		_w7364_
	);
	LUT2 #(
		.INIT('h1)
	) name3318 (
		_w7363_,
		_w7364_,
		_w7365_
	);
	LUT2 #(
		.INIT('h2)
	) name3319 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		_w7365_,
		_w7366_
	);
	LUT2 #(
		.INIT('h4)
	) name3320 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001 ,
		_w7367_
	);
	LUT2 #(
		.INIT('h8)
	) name3321 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001 ,
		_w7368_
	);
	LUT2 #(
		.INIT('h1)
	) name3322 (
		_w7367_,
		_w7368_,
		_w7369_
	);
	LUT2 #(
		.INIT('h2)
	) name3323 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w7369_,
		_w7370_
	);
	LUT2 #(
		.INIT('h4)
	) name3324 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001 ,
		_w7371_
	);
	LUT2 #(
		.INIT('h8)
	) name3325 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001 ,
		_w7372_
	);
	LUT2 #(
		.INIT('h1)
	) name3326 (
		_w7371_,
		_w7372_,
		_w7373_
	);
	LUT2 #(
		.INIT('h2)
	) name3327 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w7373_,
		_w7374_
	);
	LUT2 #(
		.INIT('h4)
	) name3328 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 ,
		_w7375_
	);
	LUT2 #(
		.INIT('h8)
	) name3329 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 ,
		_w7376_
	);
	LUT2 #(
		.INIT('h1)
	) name3330 (
		_w7375_,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('h2)
	) name3331 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w7377_,
		_w7378_
	);
	LUT2 #(
		.INIT('h4)
	) name3332 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 ,
		_w7379_
	);
	LUT2 #(
		.INIT('h8)
	) name3333 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 ,
		_w7380_
	);
	LUT2 #(
		.INIT('h1)
	) name3334 (
		_w7379_,
		_w7380_,
		_w7381_
	);
	LUT2 #(
		.INIT('h2)
	) name3335 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w7381_,
		_w7382_
	);
	LUT2 #(
		.INIT('h1)
	) name3336 (
		_w7366_,
		_w7370_,
		_w7383_
	);
	LUT2 #(
		.INIT('h1)
	) name3337 (
		_w7374_,
		_w7378_,
		_w7384_
	);
	LUT2 #(
		.INIT('h4)
	) name3338 (
		_w7382_,
		_w7384_,
		_w7385_
	);
	LUT2 #(
		.INIT('h8)
	) name3339 (
		_w7383_,
		_w7385_,
		_w7386_
	);
	LUT2 #(
		.INIT('h2)
	) name3340 (
		_w7153_,
		_w7386_,
		_w7387_
	);
	LUT2 #(
		.INIT('h8)
	) name3341 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131 ,
		_w7388_
	);
	LUT2 #(
		.INIT('h8)
	) name3342 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131 ,
		_w7389_
	);
	LUT2 #(
		.INIT('h8)
	) name3343 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131 ,
		_w7390_
	);
	LUT2 #(
		.INIT('h8)
	) name3344 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131 ,
		_w7391_
	);
	LUT2 #(
		.INIT('h8)
	) name3345 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		_w7392_
	);
	LUT2 #(
		.INIT('h8)
	) name3346 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w7393_
	);
	LUT2 #(
		.INIT('h8)
	) name3347 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131 ,
		_w7394_
	);
	LUT2 #(
		.INIT('h8)
	) name3348 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131 ,
		_w7395_
	);
	LUT2 #(
		.INIT('h8)
	) name3349 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w7396_
	);
	LUT2 #(
		.INIT('h8)
	) name3350 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w7397_
	);
	LUT2 #(
		.INIT('h8)
	) name3351 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131 ,
		_w7398_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131 ,
		_w7399_
	);
	LUT2 #(
		.INIT('h1)
	) name3353 (
		_w7388_,
		_w7389_,
		_w7400_
	);
	LUT2 #(
		.INIT('h1)
	) name3354 (
		_w7390_,
		_w7391_,
		_w7401_
	);
	LUT2 #(
		.INIT('h1)
	) name3355 (
		_w7392_,
		_w7393_,
		_w7402_
	);
	LUT2 #(
		.INIT('h1)
	) name3356 (
		_w7394_,
		_w7395_,
		_w7403_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w7396_,
		_w7397_,
		_w7404_
	);
	LUT2 #(
		.INIT('h1)
	) name3358 (
		_w7398_,
		_w7399_,
		_w7405_
	);
	LUT2 #(
		.INIT('h8)
	) name3359 (
		_w7404_,
		_w7405_,
		_w7406_
	);
	LUT2 #(
		.INIT('h8)
	) name3360 (
		_w7402_,
		_w7403_,
		_w7407_
	);
	LUT2 #(
		.INIT('h8)
	) name3361 (
		_w7400_,
		_w7401_,
		_w7408_
	);
	LUT2 #(
		.INIT('h8)
	) name3362 (
		_w7407_,
		_w7408_,
		_w7409_
	);
	LUT2 #(
		.INIT('h8)
	) name3363 (
		_w7406_,
		_w7409_,
		_w7410_
	);
	LUT2 #(
		.INIT('h2)
	) name3364 (
		_w7128_,
		_w7410_,
		_w7411_
	);
	LUT2 #(
		.INIT('h4)
	) name3365 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001 ,
		_w7412_
	);
	LUT2 #(
		.INIT('h8)
	) name3366 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001 ,
		_w7413_
	);
	LUT2 #(
		.INIT('h1)
	) name3367 (
		_w7412_,
		_w7413_,
		_w7414_
	);
	LUT2 #(
		.INIT('h2)
	) name3368 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w7414_,
		_w7415_
	);
	LUT2 #(
		.INIT('h4)
	) name3369 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001 ,
		_w7416_
	);
	LUT2 #(
		.INIT('h8)
	) name3370 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001 ,
		_w7417_
	);
	LUT2 #(
		.INIT('h1)
	) name3371 (
		_w7416_,
		_w7417_,
		_w7418_
	);
	LUT2 #(
		.INIT('h2)
	) name3372 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w7418_,
		_w7419_
	);
	LUT2 #(
		.INIT('h4)
	) name3373 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001 ,
		_w7420_
	);
	LUT2 #(
		.INIT('h8)
	) name3374 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001 ,
		_w7421_
	);
	LUT2 #(
		.INIT('h1)
	) name3375 (
		_w7420_,
		_w7421_,
		_w7422_
	);
	LUT2 #(
		.INIT('h2)
	) name3376 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w7422_,
		_w7423_
	);
	LUT2 #(
		.INIT('h4)
	) name3377 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001 ,
		_w7424_
	);
	LUT2 #(
		.INIT('h8)
	) name3378 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001 ,
		_w7425_
	);
	LUT2 #(
		.INIT('h1)
	) name3379 (
		_w7424_,
		_w7425_,
		_w7426_
	);
	LUT2 #(
		.INIT('h2)
	) name3380 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w7426_,
		_w7427_
	);
	LUT2 #(
		.INIT('h4)
	) name3381 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001 ,
		_w7428_
	);
	LUT2 #(
		.INIT('h8)
	) name3382 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001 ,
		_w7429_
	);
	LUT2 #(
		.INIT('h1)
	) name3383 (
		_w7428_,
		_w7429_,
		_w7430_
	);
	LUT2 #(
		.INIT('h2)
	) name3384 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w7430_,
		_w7431_
	);
	LUT2 #(
		.INIT('h8)
	) name3385 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w7432_
	);
	LUT2 #(
		.INIT('h1)
	) name3386 (
		_w7415_,
		_w7432_,
		_w7433_
	);
	LUT2 #(
		.INIT('h1)
	) name3387 (
		_w7419_,
		_w7423_,
		_w7434_
	);
	LUT2 #(
		.INIT('h1)
	) name3388 (
		_w7427_,
		_w7431_,
		_w7435_
	);
	LUT2 #(
		.INIT('h8)
	) name3389 (
		_w7434_,
		_w7435_,
		_w7436_
	);
	LUT2 #(
		.INIT('h8)
	) name3390 (
		_w7433_,
		_w7436_,
		_w7437_
	);
	LUT2 #(
		.INIT('h2)
	) name3391 (
		_w7093_,
		_w7437_,
		_w7438_
	);
	LUT2 #(
		.INIT('h8)
	) name3392 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[0]/P0001 ,
		_w7439_
	);
	LUT2 #(
		.INIT('h8)
	) name3393 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[0]/P0001 ,
		_w7440_
	);
	LUT2 #(
		.INIT('h8)
	) name3394 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[0]/P0001 ,
		_w7441_
	);
	LUT2 #(
		.INIT('h8)
	) name3395 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		_w7442_
	);
	LUT2 #(
		.INIT('h1)
	) name3396 (
		_w7439_,
		_w7440_,
		_w7443_
	);
	LUT2 #(
		.INIT('h1)
	) name3397 (
		_w7441_,
		_w7442_,
		_w7444_
	);
	LUT2 #(
		.INIT('h8)
	) name3398 (
		_w7443_,
		_w7444_,
		_w7445_
	);
	LUT2 #(
		.INIT('h2)
	) name3399 (
		_w7119_,
		_w7445_,
		_w7446_
	);
	LUT2 #(
		.INIT('h4)
	) name3400 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001 ,
		_w7447_
	);
	LUT2 #(
		.INIT('h8)
	) name3401 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 ,
		_w7448_
	);
	LUT2 #(
		.INIT('h1)
	) name3402 (
		_w7447_,
		_w7448_,
		_w7449_
	);
	LUT2 #(
		.INIT('h2)
	) name3403 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w7449_,
		_w7450_
	);
	LUT2 #(
		.INIT('h4)
	) name3404 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001 ,
		_w7451_
	);
	LUT2 #(
		.INIT('h8)
	) name3405 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001 ,
		_w7452_
	);
	LUT2 #(
		.INIT('h1)
	) name3406 (
		_w7451_,
		_w7452_,
		_w7453_
	);
	LUT2 #(
		.INIT('h2)
	) name3407 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w7453_,
		_w7454_
	);
	LUT2 #(
		.INIT('h4)
	) name3408 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001 ,
		_w7455_
	);
	LUT2 #(
		.INIT('h8)
	) name3409 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001 ,
		_w7456_
	);
	LUT2 #(
		.INIT('h1)
	) name3410 (
		_w7455_,
		_w7456_,
		_w7457_
	);
	LUT2 #(
		.INIT('h2)
	) name3411 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w7457_,
		_w7458_
	);
	LUT2 #(
		.INIT('h4)
	) name3412 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001 ,
		_w7459_
	);
	LUT2 #(
		.INIT('h8)
	) name3413 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001 ,
		_w7460_
	);
	LUT2 #(
		.INIT('h1)
	) name3414 (
		_w7459_,
		_w7460_,
		_w7461_
	);
	LUT2 #(
		.INIT('h2)
	) name3415 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w7461_,
		_w7462_
	);
	LUT2 #(
		.INIT('h4)
	) name3416 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001 ,
		_w7463_
	);
	LUT2 #(
		.INIT('h8)
	) name3417 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001 ,
		_w7464_
	);
	LUT2 #(
		.INIT('h1)
	) name3418 (
		_w7463_,
		_w7464_,
		_w7465_
	);
	LUT2 #(
		.INIT('h2)
	) name3419 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w7465_,
		_w7466_
	);
	LUT2 #(
		.INIT('h4)
	) name3420 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001 ,
		_w7467_
	);
	LUT2 #(
		.INIT('h8)
	) name3421 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 ,
		_w7468_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		_w7467_,
		_w7468_,
		_w7469_
	);
	LUT2 #(
		.INIT('h2)
	) name3423 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w7469_,
		_w7470_
	);
	LUT2 #(
		.INIT('h4)
	) name3424 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 ,
		_w7471_
	);
	LUT2 #(
		.INIT('h8)
	) name3425 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 ,
		_w7472_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		_w7471_,
		_w7472_,
		_w7473_
	);
	LUT2 #(
		.INIT('h2)
	) name3427 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h1)
	) name3428 (
		_w7450_,
		_w7454_,
		_w7475_
	);
	LUT2 #(
		.INIT('h1)
	) name3429 (
		_w7458_,
		_w7462_,
		_w7476_
	);
	LUT2 #(
		.INIT('h1)
	) name3430 (
		_w7466_,
		_w7470_,
		_w7477_
	);
	LUT2 #(
		.INIT('h4)
	) name3431 (
		_w7474_,
		_w7477_,
		_w7478_
	);
	LUT2 #(
		.INIT('h8)
	) name3432 (
		_w7475_,
		_w7476_,
		_w7479_
	);
	LUT2 #(
		.INIT('h8)
	) name3433 (
		_w7478_,
		_w7479_,
		_w7480_
	);
	LUT2 #(
		.INIT('h2)
	) name3434 (
		_w7179_,
		_w7480_,
		_w7481_
	);
	LUT2 #(
		.INIT('h8)
	) name3435 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 ,
		_w7482_
	);
	LUT2 #(
		.INIT('h8)
	) name3436 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 ,
		_w7483_
	);
	LUT2 #(
		.INIT('h8)
	) name3437 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131 ,
		_w7484_
	);
	LUT2 #(
		.INIT('h8)
	) name3438 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131 ,
		_w7485_
	);
	LUT2 #(
		.INIT('h8)
	) name3439 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131 ,
		_w7486_
	);
	LUT2 #(
		.INIT('h8)
	) name3440 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131 ,
		_w7487_
	);
	LUT2 #(
		.INIT('h8)
	) name3441 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 ,
		_w7488_
	);
	LUT2 #(
		.INIT('h8)
	) name3442 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w7489_
	);
	LUT2 #(
		.INIT('h8)
	) name3443 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131 ,
		_w7490_
	);
	LUT2 #(
		.INIT('h8)
	) name3444 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131 ,
		_w7491_
	);
	LUT2 #(
		.INIT('h8)
	) name3445 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131 ,
		_w7492_
	);
	LUT2 #(
		.INIT('h8)
	) name3446 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131 ,
		_w7493_
	);
	LUT2 #(
		.INIT('h1)
	) name3447 (
		_w7482_,
		_w7483_,
		_w7494_
	);
	LUT2 #(
		.INIT('h1)
	) name3448 (
		_w7484_,
		_w7485_,
		_w7495_
	);
	LUT2 #(
		.INIT('h1)
	) name3449 (
		_w7486_,
		_w7487_,
		_w7496_
	);
	LUT2 #(
		.INIT('h1)
	) name3450 (
		_w7488_,
		_w7489_,
		_w7497_
	);
	LUT2 #(
		.INIT('h1)
	) name3451 (
		_w7490_,
		_w7491_,
		_w7498_
	);
	LUT2 #(
		.INIT('h1)
	) name3452 (
		_w7492_,
		_w7493_,
		_w7499_
	);
	LUT2 #(
		.INIT('h8)
	) name3453 (
		_w7498_,
		_w7499_,
		_w7500_
	);
	LUT2 #(
		.INIT('h8)
	) name3454 (
		_w7496_,
		_w7497_,
		_w7501_
	);
	LUT2 #(
		.INIT('h8)
	) name3455 (
		_w7494_,
		_w7495_,
		_w7502_
	);
	LUT2 #(
		.INIT('h8)
	) name3456 (
		_w7501_,
		_w7502_,
		_w7503_
	);
	LUT2 #(
		.INIT('h8)
	) name3457 (
		_w7500_,
		_w7503_,
		_w7504_
	);
	LUT2 #(
		.INIT('h2)
	) name3458 (
		_w7068_,
		_w7504_,
		_w7505_
	);
	LUT2 #(
		.INIT('h8)
	) name3459 (
		\emc_WSCRreg_DO_reg[0]/NET0131 ,
		_w7251_,
		_w7506_
	);
	LUT2 #(
		.INIT('h8)
	) name3460 (
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w7259_,
		_w7507_
	);
	LUT2 #(
		.INIT('h8)
	) name3461 (
		\sport1_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w7263_,
		_w7508_
	);
	LUT2 #(
		.INIT('h8)
	) name3462 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w7287_,
		_w7509_
	);
	LUT2 #(
		.INIT('h8)
	) name3463 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w7249_,
		_w7510_
	);
	LUT2 #(
		.INIT('h8)
	) name3464 (
		\PIO_oe[0]_pad ,
		_w7244_,
		_w7511_
	);
	LUT2 #(
		.INIT('h8)
	) name3465 (
		\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w7256_,
		_w7512_
	);
	LUT2 #(
		.INIT('h8)
	) name3466 (
		_w7226_,
		_w7269_,
		_w7513_
	);
	LUT2 #(
		.INIT('h8)
	) name3467 (
		_w7268_,
		_w7513_,
		_w7514_
	);
	LUT2 #(
		.INIT('h8)
	) name3468 (
		\emc_WSCRext_reg_DO_reg[0]/NET0131 ,
		_w7514_,
		_w7515_
	);
	LUT2 #(
		.INIT('h8)
	) name3469 (
		\memc_usysr_DO_reg[0]/NET0131 ,
		_w7301_,
		_w7516_
	);
	LUT2 #(
		.INIT('h8)
	) name3470 (
		\sport0_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w7295_,
		_w7517_
	);
	LUT2 #(
		.INIT('h8)
	) name3471 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w7299_,
		_w7518_
	);
	LUT2 #(
		.INIT('h8)
	) name3472 (
		\pio_PINT_reg[0]/NET0131 ,
		_w7271_,
		_w7519_
	);
	LUT2 #(
		.INIT('h8)
	) name3473 (
		\tm_TCR_TMP_reg[0]/NET0131 ,
		_w7289_,
		_w7520_
	);
	LUT2 #(
		.INIT('h8)
	) name3474 (
		_w7237_,
		_w7268_,
		_w7521_
	);
	LUT2 #(
		.INIT('h8)
	) name3475 (
		_w7269_,
		_w7521_,
		_w7522_
	);
	LUT2 #(
		.INIT('h8)
	) name3476 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w7234_,
		_w7523_
	);
	LUT2 #(
		.INIT('h8)
	) name3477 (
		\pio_pmask_reg_DO_reg[0]/NET0131 ,
		_w7297_,
		_w7524_
	);
	LUT2 #(
		.INIT('h8)
	) name3478 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w7525_
	);
	LUT2 #(
		.INIT('h8)
	) name3479 (
		_w7226_,
		_w7525_,
		_w7526_
	);
	LUT2 #(
		.INIT('h8)
	) name3480 (
		_w7268_,
		_w7526_,
		_w7527_
	);
	LUT2 #(
		.INIT('h8)
	) name3481 (
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w7527_,
		_w7528_
	);
	LUT2 #(
		.INIT('h8)
	) name3482 (
		\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w7247_,
		_w7529_
	);
	LUT2 #(
		.INIT('h8)
	) name3483 (
		_w7232_,
		_w7269_,
		_w7530_
	);
	LUT2 #(
		.INIT('h8)
	) name3484 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\memc_selMIO_E_reg/P0001 ,
		_w7531_
	);
	LUT2 #(
		.INIT('h8)
	) name3485 (
		_w7530_,
		_w7531_,
		_w7532_
	);
	LUT2 #(
		.INIT('h8)
	) name3486 (
		\idma_DOVL_reg[0]/NET0131 ,
		_w7532_,
		_w7533_
	);
	LUT2 #(
		.INIT('h8)
	) name3487 (
		_w7286_,
		_w7530_,
		_w7534_
	);
	LUT2 #(
		.INIT('h8)
	) name3488 (
		\bdma_BOVL_reg[0]/NET0131 ,
		_w7534_,
		_w7535_
	);
	LUT2 #(
		.INIT('h8)
	) name3489 (
		\tm_tpr_reg_DO_reg[0]/NET0131 ,
		_w7293_,
		_w7536_
	);
	LUT2 #(
		.INIT('h8)
	) name3490 (
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w7273_,
		_w7537_
	);
	LUT2 #(
		.INIT('h8)
	) name3491 (
		\bdma_BEAD_reg[0]/NET0131 ,
		_w7303_,
		_w7538_
	);
	LUT2 #(
		.INIT('h8)
	) name3492 (
		\bdma_BCTL_reg[0]/NET0131 ,
		_w7230_,
		_w7539_
	);
	LUT2 #(
		.INIT('h8)
	) name3493 (
		_w7227_,
		_w7236_,
		_w7540_
	);
	LUT2 #(
		.INIT('h8)
	) name3494 (
		\tm_tsr_reg_DO_reg[0]/NET0131 ,
		_w7540_,
		_w7541_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w7281_,
		_w7542_
	);
	LUT2 #(
		.INIT('h8)
	) name3496 (
		\clkc_ckr_reg_DO_reg[0]/NET0131 ,
		_w7239_,
		_w7543_
	);
	LUT2 #(
		.INIT('h8)
	) name3497 (
		\sport0_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w7276_,
		_w7544_
	);
	LUT2 #(
		.INIT('h8)
	) name3498 (
		\PIO_out[0]_pad ,
		_w7291_,
		_w7545_
	);
	LUT2 #(
		.INIT('h1)
	) name3499 (
		_w7506_,
		_w7522_,
		_w7546_
	);
	LUT2 #(
		.INIT('h1)
	) name3500 (
		_w7507_,
		_w7508_,
		_w7547_
	);
	LUT2 #(
		.INIT('h1)
	) name3501 (
		_w7510_,
		_w7511_,
		_w7548_
	);
	LUT2 #(
		.INIT('h1)
	) name3502 (
		_w7512_,
		_w7515_,
		_w7549_
	);
	LUT2 #(
		.INIT('h1)
	) name3503 (
		_w7516_,
		_w7517_,
		_w7550_
	);
	LUT2 #(
		.INIT('h1)
	) name3504 (
		_w7518_,
		_w7519_,
		_w7551_
	);
	LUT2 #(
		.INIT('h1)
	) name3505 (
		_w7520_,
		_w7524_,
		_w7552_
	);
	LUT2 #(
		.INIT('h1)
	) name3506 (
		_w7528_,
		_w7529_,
		_w7553_
	);
	LUT2 #(
		.INIT('h1)
	) name3507 (
		_w7533_,
		_w7536_,
		_w7554_
	);
	LUT2 #(
		.INIT('h1)
	) name3508 (
		_w7537_,
		_w7541_,
		_w7555_
	);
	LUT2 #(
		.INIT('h1)
	) name3509 (
		_w7542_,
		_w7543_,
		_w7556_
	);
	LUT2 #(
		.INIT('h1)
	) name3510 (
		_w7544_,
		_w7545_,
		_w7557_
	);
	LUT2 #(
		.INIT('h8)
	) name3511 (
		_w7556_,
		_w7557_,
		_w7558_
	);
	LUT2 #(
		.INIT('h8)
	) name3512 (
		_w7554_,
		_w7555_,
		_w7559_
	);
	LUT2 #(
		.INIT('h8)
	) name3513 (
		_w7552_,
		_w7553_,
		_w7560_
	);
	LUT2 #(
		.INIT('h8)
	) name3514 (
		_w7550_,
		_w7551_,
		_w7561_
	);
	LUT2 #(
		.INIT('h8)
	) name3515 (
		_w7548_,
		_w7549_,
		_w7562_
	);
	LUT2 #(
		.INIT('h8)
	) name3516 (
		_w7546_,
		_w7547_,
		_w7563_
	);
	LUT2 #(
		.INIT('h8)
	) name3517 (
		_w7562_,
		_w7563_,
		_w7564_
	);
	LUT2 #(
		.INIT('h8)
	) name3518 (
		_w7560_,
		_w7561_,
		_w7565_
	);
	LUT2 #(
		.INIT('h8)
	) name3519 (
		_w7558_,
		_w7559_,
		_w7566_
	);
	LUT2 #(
		.INIT('h8)
	) name3520 (
		_w7565_,
		_w7566_,
		_w7567_
	);
	LUT2 #(
		.INIT('h4)
	) name3521 (
		_w7523_,
		_w7564_,
		_w7568_
	);
	LUT2 #(
		.INIT('h1)
	) name3522 (
		_w7538_,
		_w7539_,
		_w7569_
	);
	LUT2 #(
		.INIT('h8)
	) name3523 (
		_w7568_,
		_w7569_,
		_w7570_
	);
	LUT2 #(
		.INIT('h4)
	) name3524 (
		_w7509_,
		_w7567_,
		_w7571_
	);
	LUT2 #(
		.INIT('h4)
	) name3525 (
		_w7535_,
		_w7571_,
		_w7572_
	);
	LUT2 #(
		.INIT('h8)
	) name3526 (
		_w7570_,
		_w7572_,
		_w7573_
	);
	LUT2 #(
		.INIT('h2)
	) name3527 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7573_,
		_w7574_
	);
	LUT2 #(
		.INIT('h8)
	) name3528 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w7575_
	);
	LUT2 #(
		.INIT('h8)
	) name3529 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w7576_
	);
	LUT2 #(
		.INIT('h8)
	) name3530 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[0]/NET0131 ,
		_w7577_
	);
	LUT2 #(
		.INIT('h2)
	) name3531 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4588_,
		_w7578_
	);
	LUT2 #(
		.INIT('h2)
	) name3532 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w7216_,
		_w7579_
	);
	LUT2 #(
		.INIT('h8)
	) name3533 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w7580_
	);
	LUT2 #(
		.INIT('h8)
	) name3534 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		_w7581_
	);
	LUT2 #(
		.INIT('h8)
	) name3535 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w7582_
	);
	LUT2 #(
		.INIT('h8)
	) name3536 (
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\core_c_psq_ICNTL_reg_DO_reg[0]/NET0131 ,
		_w7583_
	);
	LUT2 #(
		.INIT('h8)
	) name3537 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		_w7584_
	);
	LUT2 #(
		.INIT('h1)
	) name3538 (
		_w7575_,
		_w7576_,
		_w7585_
	);
	LUT2 #(
		.INIT('h1)
	) name3539 (
		_w7577_,
		_w7580_,
		_w7586_
	);
	LUT2 #(
		.INIT('h1)
	) name3540 (
		_w7581_,
		_w7582_,
		_w7587_
	);
	LUT2 #(
		.INIT('h1)
	) name3541 (
		_w7583_,
		_w7584_,
		_w7588_
	);
	LUT2 #(
		.INIT('h8)
	) name3542 (
		_w7587_,
		_w7588_,
		_w7589_
	);
	LUT2 #(
		.INIT('h8)
	) name3543 (
		_w7585_,
		_w7586_,
		_w7590_
	);
	LUT2 #(
		.INIT('h4)
	) name3544 (
		_w7579_,
		_w7590_,
		_w7591_
	);
	LUT2 #(
		.INIT('h8)
	) name3545 (
		_w7589_,
		_w7591_,
		_w7592_
	);
	LUT2 #(
		.INIT('h4)
	) name3546 (
		_w7578_,
		_w7592_,
		_w7593_
	);
	LUT2 #(
		.INIT('h2)
	) name3547 (
		_w7215_,
		_w7593_,
		_w7594_
	);
	LUT2 #(
		.INIT('h1)
	) name3548 (
		_w7411_,
		_w7446_,
		_w7595_
	);
	LUT2 #(
		.INIT('h4)
	) name3549 (
		_w7505_,
		_w7595_,
		_w7596_
	);
	LUT2 #(
		.INIT('h1)
	) name3550 (
		_w7387_,
		_w7438_,
		_w7597_
	);
	LUT2 #(
		.INIT('h4)
	) name3551 (
		_w7481_,
		_w7597_,
		_w7598_
	);
	LUT2 #(
		.INIT('h8)
	) name3552 (
		_w7596_,
		_w7598_,
		_w7599_
	);
	LUT2 #(
		.INIT('h4)
	) name3553 (
		_w7594_,
		_w7599_,
		_w7600_
	);
	LUT2 #(
		.INIT('h4)
	) name3554 (
		_w7574_,
		_w7600_,
		_w7601_
	);
	LUT2 #(
		.INIT('h4)
	) name3555 (
		_w7362_,
		_w7601_,
		_w7602_
	);
	LUT2 #(
		.INIT('h1)
	) name3556 (
		\emc_DMDoe_reg/NET0131 ,
		_w7602_,
		_w7603_
	);
	LUT2 #(
		.INIT('h8)
	) name3557 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[0]/P0001 ,
		_w7604_
	);
	LUT2 #(
		.INIT('h2)
	) name3558 (
		_w7057_,
		_w7604_,
		_w7605_
	);
	LUT2 #(
		.INIT('h4)
	) name3559 (
		_w7603_,
		_w7605_,
		_w7606_
	);
	LUT2 #(
		.INIT('h1)
	) name3560 (
		_w7361_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h8)
	) name3561 (
		_w6135_,
		_w7607_,
		_w7608_
	);
	LUT2 #(
		.INIT('h8)
	) name3562 (
		\core_dag_ilm1reg_I_reg[0]/NET0131 ,
		_w6345_,
		_w7609_
	);
	LUT2 #(
		.INIT('h8)
	) name3563 (
		_w6497_,
		_w6527_,
		_w7610_
	);
	LUT2 #(
		.INIT('h2)
	) name3564 (
		_w6498_,
		_w6527_,
		_w7611_
	);
	LUT2 #(
		.INIT('h1)
	) name3565 (
		_w7610_,
		_w7611_,
		_w7612_
	);
	LUT2 #(
		.INIT('h4)
	) name3566 (
		_w6362_,
		_w7612_,
		_w7613_
	);
	LUT2 #(
		.INIT('h1)
	) name3567 (
		_w6365_,
		_w7612_,
		_w7614_
	);
	LUT2 #(
		.INIT('h2)
	) name3568 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w7613_,
		_w7615_
	);
	LUT2 #(
		.INIT('h4)
	) name3569 (
		_w7614_,
		_w7615_,
		_w7616_
	);
	LUT2 #(
		.INIT('h1)
	) name3570 (
		_w6362_,
		_w6496_,
		_w7617_
	);
	LUT2 #(
		.INIT('h8)
	) name3571 (
		_w6365_,
		_w6496_,
		_w7618_
	);
	LUT2 #(
		.INIT('h1)
	) name3572 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w7617_,
		_w7619_
	);
	LUT2 #(
		.INIT('h4)
	) name3573 (
		_w7618_,
		_w7619_,
		_w7620_
	);
	LUT2 #(
		.INIT('h1)
	) name3574 (
		_w7609_,
		_w7616_,
		_w7621_
	);
	LUT2 #(
		.INIT('h4)
	) name3575 (
		_w7620_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('h1)
	) name3576 (
		_w6135_,
		_w7622_,
		_w7623_
	);
	LUT2 #(
		.INIT('h2)
	) name3577 (
		_w6176_,
		_w7608_,
		_w7624_
	);
	LUT2 #(
		.INIT('h4)
	) name3578 (
		_w7623_,
		_w7624_,
		_w7625_
	);
	LUT2 #(
		.INIT('h1)
	) name3579 (
		_w7343_,
		_w7625_,
		_w7626_
	);
	LUT2 #(
		.INIT('h2)
	) name3580 (
		_w7005_,
		_w7626_,
		_w7627_
	);
	LUT2 #(
		.INIT('h1)
	) name3581 (
		_w7006_,
		_w7627_,
		_w7628_
	);
	LUT2 #(
		.INIT('h8)
	) name3582 (
		\core_dag_ilm1reg_I_reg[10]/NET0131 ,
		_w6423_,
		_w7629_
	);
	LUT2 #(
		.INIT('h4)
	) name3583 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w6496_,
		_w7630_
	);
	LUT2 #(
		.INIT('h1)
	) name3584 (
		_w7610_,
		_w7630_,
		_w7631_
	);
	LUT2 #(
		.INIT('h4)
	) name3585 (
		_w6419_,
		_w6461_,
		_w7632_
	);
	LUT2 #(
		.INIT('h1)
	) name3586 (
		_w6434_,
		_w6457_,
		_w7633_
	);
	LUT2 #(
		.INIT('h2)
	) name3587 (
		_w7632_,
		_w7633_,
		_w7634_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		_w7632_,
		_w7633_,
		_w7635_
	);
	LUT2 #(
		.INIT('h1)
	) name3589 (
		_w7634_,
		_w7635_,
		_w7636_
	);
	LUT2 #(
		.INIT('h4)
	) name3590 (
		_w7631_,
		_w7636_,
		_w7637_
	);
	LUT2 #(
		.INIT('h1)
	) name3591 (
		_w6516_,
		_w6521_,
		_w7638_
	);
	LUT2 #(
		.INIT('h2)
	) name3592 (
		_w6427_,
		_w7638_,
		_w7639_
	);
	LUT2 #(
		.INIT('h4)
	) name3593 (
		_w6427_,
		_w7638_,
		_w7640_
	);
	LUT2 #(
		.INIT('h1)
	) name3594 (
		_w7639_,
		_w7640_,
		_w7641_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		_w7631_,
		_w7641_,
		_w7642_
	);
	LUT2 #(
		.INIT('h1)
	) name3596 (
		_w7629_,
		_w7637_,
		_w7643_
	);
	LUT2 #(
		.INIT('h4)
	) name3597 (
		_w7642_,
		_w7643_,
		_w7644_
	);
	LUT2 #(
		.INIT('h4)
	) name3598 (
		_w6135_,
		_w7644_,
		_w7645_
	);
	LUT2 #(
		.INIT('h8)
	) name3599 (
		\DM_rdm[10]_pad ,
		_w7016_,
		_w7646_
	);
	LUT2 #(
		.INIT('h8)
	) name3600 (
		\DM_rd1[10]_pad ,
		_w7022_,
		_w7647_
	);
	LUT2 #(
		.INIT('h8)
	) name3601 (
		\DM_rd4[10]_pad ,
		_w7028_,
		_w7648_
	);
	LUT2 #(
		.INIT('h8)
	) name3602 (
		\DM_rd6[10]_pad ,
		_w7031_,
		_w7649_
	);
	LUT2 #(
		.INIT('h8)
	) name3603 (
		\DM_rd7[10]_pad ,
		_w7034_,
		_w7650_
	);
	LUT2 #(
		.INIT('h8)
	) name3604 (
		\DM_rd3[10]_pad ,
		_w7038_,
		_w7651_
	);
	LUT2 #(
		.INIT('h2)
	) name3605 (
		\DM_rd0[10]_pad ,
		_w7053_,
		_w7652_
	);
	LUT2 #(
		.INIT('h8)
	) name3606 (
		\DM_rd5[10]_pad ,
		_w7043_,
		_w7653_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		\DM_rd2[10]_pad ,
		_w7041_,
		_w7654_
	);
	LUT2 #(
		.INIT('h1)
	) name3608 (
		_w7647_,
		_w7651_,
		_w7655_
	);
	LUT2 #(
		.INIT('h4)
	) name3609 (
		_w7654_,
		_w7655_,
		_w7656_
	);
	LUT2 #(
		.INIT('h1)
	) name3610 (
		_w7057_,
		_w7646_,
		_w7657_
	);
	LUT2 #(
		.INIT('h1)
	) name3611 (
		_w7649_,
		_w7650_,
		_w7658_
	);
	LUT2 #(
		.INIT('h8)
	) name3612 (
		_w7657_,
		_w7658_,
		_w7659_
	);
	LUT2 #(
		.INIT('h4)
	) name3613 (
		_w7648_,
		_w7656_,
		_w7660_
	);
	LUT2 #(
		.INIT('h4)
	) name3614 (
		_w7653_,
		_w7660_,
		_w7661_
	);
	LUT2 #(
		.INIT('h8)
	) name3615 (
		_w7659_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h4)
	) name3616 (
		_w7652_,
		_w7662_,
		_w7663_
	);
	LUT2 #(
		.INIT('h8)
	) name3617 (
		\regout_STD_C_reg[10]/P0001 ,
		_w6988_,
		_w7664_
	);
	LUT2 #(
		.INIT('h8)
	) name3618 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131 ,
		_w7665_
	);
	LUT2 #(
		.INIT('h8)
	) name3619 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131 ,
		_w7666_
	);
	LUT2 #(
		.INIT('h8)
	) name3620 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131 ,
		_w7667_
	);
	LUT2 #(
		.INIT('h8)
	) name3621 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131 ,
		_w7668_
	);
	LUT2 #(
		.INIT('h8)
	) name3622 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 ,
		_w7669_
	);
	LUT2 #(
		.INIT('h8)
	) name3623 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 ,
		_w7670_
	);
	LUT2 #(
		.INIT('h8)
	) name3624 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 ,
		_w7671_
	);
	LUT2 #(
		.INIT('h8)
	) name3625 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131 ,
		_w7672_
	);
	LUT2 #(
		.INIT('h8)
	) name3626 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131 ,
		_w7673_
	);
	LUT2 #(
		.INIT('h8)
	) name3627 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w7674_
	);
	LUT2 #(
		.INIT('h8)
	) name3628 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131 ,
		_w7675_
	);
	LUT2 #(
		.INIT('h8)
	) name3629 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131 ,
		_w7676_
	);
	LUT2 #(
		.INIT('h1)
	) name3630 (
		_w7665_,
		_w7666_,
		_w7677_
	);
	LUT2 #(
		.INIT('h1)
	) name3631 (
		_w7667_,
		_w7668_,
		_w7678_
	);
	LUT2 #(
		.INIT('h1)
	) name3632 (
		_w7669_,
		_w7670_,
		_w7679_
	);
	LUT2 #(
		.INIT('h1)
	) name3633 (
		_w7671_,
		_w7672_,
		_w7680_
	);
	LUT2 #(
		.INIT('h1)
	) name3634 (
		_w7673_,
		_w7674_,
		_w7681_
	);
	LUT2 #(
		.INIT('h1)
	) name3635 (
		_w7675_,
		_w7676_,
		_w7682_
	);
	LUT2 #(
		.INIT('h8)
	) name3636 (
		_w7681_,
		_w7682_,
		_w7683_
	);
	LUT2 #(
		.INIT('h8)
	) name3637 (
		_w7679_,
		_w7680_,
		_w7684_
	);
	LUT2 #(
		.INIT('h8)
	) name3638 (
		_w7677_,
		_w7678_,
		_w7685_
	);
	LUT2 #(
		.INIT('h8)
	) name3639 (
		_w7684_,
		_w7685_,
		_w7686_
	);
	LUT2 #(
		.INIT('h8)
	) name3640 (
		_w7683_,
		_w7686_,
		_w7687_
	);
	LUT2 #(
		.INIT('h2)
	) name3641 (
		_w7068_,
		_w7687_,
		_w7688_
	);
	LUT2 #(
		.INIT('h8)
	) name3642 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w7263_,
		_w7689_
	);
	LUT2 #(
		.INIT('h8)
	) name3643 (
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		_w7689_,
		_w7690_
	);
	LUT2 #(
		.INIT('h8)
	) name3644 (
		\emc_WSCRreg_DO_reg[10]/NET0131 ,
		_w7251_,
		_w7691_
	);
	LUT2 #(
		.INIT('h8)
	) name3645 (
		\bdma_BCTL_reg[10]/NET0131 ,
		_w7230_,
		_w7692_
	);
	LUT2 #(
		.INIT('h8)
	) name3646 (
		\tm_tpr_reg_DO_reg[10]/NET0131 ,
		_w7293_,
		_w7693_
	);
	LUT2 #(
		.INIT('h8)
	) name3647 (
		\bdma_BEAD_reg[10]/NET0131 ,
		_w7303_,
		_w7694_
	);
	LUT2 #(
		.INIT('h8)
	) name3648 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		_w7287_,
		_w7695_
	);
	LUT2 #(
		.INIT('h8)
	) name3649 (
		\sport0_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w7249_,
		_w7696_
	);
	LUT2 #(
		.INIT('h8)
	) name3650 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		_w7289_,
		_w7697_
	);
	LUT2 #(
		.INIT('h8)
	) name3651 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w7234_,
		_w7698_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		\idma_DOVL_reg[10]/NET0131 ,
		_w7532_,
		_w7699_
	);
	LUT2 #(
		.INIT('h8)
	) name3653 (
		\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w7256_,
		_w7700_
	);
	LUT2 #(
		.INIT('h8)
	) name3654 (
		\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w7247_,
		_w7701_
	);
	LUT2 #(
		.INIT('h8)
	) name3655 (
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w7273_,
		_w7702_
	);
	LUT2 #(
		.INIT('h8)
	) name3656 (
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w7259_,
		_w7703_
	);
	LUT2 #(
		.INIT('h8)
	) name3657 (
		\memc_usysr_DO_reg[10]/NET0131 ,
		_w7301_,
		_w7704_
	);
	LUT2 #(
		.INIT('h8)
	) name3658 (
		\sport1_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w7281_,
		_w7705_
	);
	LUT2 #(
		.INIT('h8)
	) name3659 (
		\clkc_ckr_reg_DO_reg[10]/NET0131 ,
		_w7239_,
		_w7706_
	);
	LUT2 #(
		.INIT('h8)
	) name3660 (
		\bdma_BOVL_reg[10]/NET0131 ,
		_w7534_,
		_w7707_
	);
	LUT2 #(
		.INIT('h8)
	) name3661 (
		\sport1_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w7527_,
		_w7708_
	);
	LUT2 #(
		.INIT('h8)
	) name3662 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w7299_,
		_w7709_
	);
	LUT2 #(
		.INIT('h8)
	) name3663 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w7276_,
		_w7710_
	);
	LUT2 #(
		.INIT('h8)
	) name3664 (
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		_w7710_,
		_w7711_
	);
	LUT2 #(
		.INIT('h8)
	) name3665 (
		\sport0_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w7295_,
		_w7712_
	);
	LUT2 #(
		.INIT('h1)
	) name3666 (
		_w7691_,
		_w7693_,
		_w7713_
	);
	LUT2 #(
		.INIT('h1)
	) name3667 (
		_w7696_,
		_w7697_,
		_w7714_
	);
	LUT2 #(
		.INIT('h1)
	) name3668 (
		_w7699_,
		_w7700_,
		_w7715_
	);
	LUT2 #(
		.INIT('h1)
	) name3669 (
		_w7701_,
		_w7702_,
		_w7716_
	);
	LUT2 #(
		.INIT('h1)
	) name3670 (
		_w7703_,
		_w7704_,
		_w7717_
	);
	LUT2 #(
		.INIT('h1)
	) name3671 (
		_w7705_,
		_w7706_,
		_w7718_
	);
	LUT2 #(
		.INIT('h1)
	) name3672 (
		_w7708_,
		_w7709_,
		_w7719_
	);
	LUT2 #(
		.INIT('h4)
	) name3673 (
		_w7712_,
		_w7719_,
		_w7720_
	);
	LUT2 #(
		.INIT('h8)
	) name3674 (
		_w7717_,
		_w7718_,
		_w7721_
	);
	LUT2 #(
		.INIT('h8)
	) name3675 (
		_w7715_,
		_w7716_,
		_w7722_
	);
	LUT2 #(
		.INIT('h8)
	) name3676 (
		_w7713_,
		_w7714_,
		_w7723_
	);
	LUT2 #(
		.INIT('h1)
	) name3677 (
		_w7690_,
		_w7711_,
		_w7724_
	);
	LUT2 #(
		.INIT('h8)
	) name3678 (
		_w7723_,
		_w7724_,
		_w7725_
	);
	LUT2 #(
		.INIT('h8)
	) name3679 (
		_w7721_,
		_w7722_,
		_w7726_
	);
	LUT2 #(
		.INIT('h8)
	) name3680 (
		_w7720_,
		_w7726_,
		_w7727_
	);
	LUT2 #(
		.INIT('h4)
	) name3681 (
		_w7692_,
		_w7725_,
		_w7728_
	);
	LUT2 #(
		.INIT('h1)
	) name3682 (
		_w7694_,
		_w7698_,
		_w7729_
	);
	LUT2 #(
		.INIT('h8)
	) name3683 (
		_w7728_,
		_w7729_,
		_w7730_
	);
	LUT2 #(
		.INIT('h4)
	) name3684 (
		_w7695_,
		_w7727_,
		_w7731_
	);
	LUT2 #(
		.INIT('h4)
	) name3685 (
		_w7707_,
		_w7731_,
		_w7732_
	);
	LUT2 #(
		.INIT('h8)
	) name3686 (
		_w7730_,
		_w7732_,
		_w7733_
	);
	LUT2 #(
		.INIT('h2)
	) name3687 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w7733_,
		_w7734_
	);
	LUT2 #(
		.INIT('h4)
	) name3688 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001 ,
		_w7735_
	);
	LUT2 #(
		.INIT('h8)
	) name3689 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 ,
		_w7736_
	);
	LUT2 #(
		.INIT('h1)
	) name3690 (
		_w7735_,
		_w7736_,
		_w7737_
	);
	LUT2 #(
		.INIT('h2)
	) name3691 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w7737_,
		_w7738_
	);
	LUT2 #(
		.INIT('h4)
	) name3692 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001 ,
		_w7739_
	);
	LUT2 #(
		.INIT('h8)
	) name3693 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001 ,
		_w7740_
	);
	LUT2 #(
		.INIT('h1)
	) name3694 (
		_w7739_,
		_w7740_,
		_w7741_
	);
	LUT2 #(
		.INIT('h2)
	) name3695 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w7741_,
		_w7742_
	);
	LUT2 #(
		.INIT('h4)
	) name3696 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001 ,
		_w7743_
	);
	LUT2 #(
		.INIT('h8)
	) name3697 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001 ,
		_w7744_
	);
	LUT2 #(
		.INIT('h1)
	) name3698 (
		_w7743_,
		_w7744_,
		_w7745_
	);
	LUT2 #(
		.INIT('h2)
	) name3699 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w7745_,
		_w7746_
	);
	LUT2 #(
		.INIT('h4)
	) name3700 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001 ,
		_w7747_
	);
	LUT2 #(
		.INIT('h8)
	) name3701 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001 ,
		_w7748_
	);
	LUT2 #(
		.INIT('h1)
	) name3702 (
		_w7747_,
		_w7748_,
		_w7749_
	);
	LUT2 #(
		.INIT('h2)
	) name3703 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('h4)
	) name3704 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001 ,
		_w7751_
	);
	LUT2 #(
		.INIT('h8)
	) name3705 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 ,
		_w7752_
	);
	LUT2 #(
		.INIT('h1)
	) name3706 (
		_w7751_,
		_w7752_,
		_w7753_
	);
	LUT2 #(
		.INIT('h2)
	) name3707 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w7753_,
		_w7754_
	);
	LUT2 #(
		.INIT('h4)
	) name3708 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001 ,
		_w7755_
	);
	LUT2 #(
		.INIT('h8)
	) name3709 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001 ,
		_w7756_
	);
	LUT2 #(
		.INIT('h1)
	) name3710 (
		_w7755_,
		_w7756_,
		_w7757_
	);
	LUT2 #(
		.INIT('h2)
	) name3711 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w7757_,
		_w7758_
	);
	LUT2 #(
		.INIT('h1)
	) name3712 (
		_w7207_,
		_w7738_,
		_w7759_
	);
	LUT2 #(
		.INIT('h1)
	) name3713 (
		_w7742_,
		_w7746_,
		_w7760_
	);
	LUT2 #(
		.INIT('h1)
	) name3714 (
		_w7750_,
		_w7754_,
		_w7761_
	);
	LUT2 #(
		.INIT('h4)
	) name3715 (
		_w7758_,
		_w7761_,
		_w7762_
	);
	LUT2 #(
		.INIT('h8)
	) name3716 (
		_w7759_,
		_w7760_,
		_w7763_
	);
	LUT2 #(
		.INIT('h8)
	) name3717 (
		_w7762_,
		_w7763_,
		_w7764_
	);
	LUT2 #(
		.INIT('h2)
	) name3718 (
		_w7179_,
		_w7764_,
		_w7765_
	);
	LUT2 #(
		.INIT('h4)
	) name3719 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001 ,
		_w7766_
	);
	LUT2 #(
		.INIT('h8)
	) name3720 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001 ,
		_w7767_
	);
	LUT2 #(
		.INIT('h1)
	) name3721 (
		_w7766_,
		_w7767_,
		_w7768_
	);
	LUT2 #(
		.INIT('h2)
	) name3722 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w7768_,
		_w7769_
	);
	LUT2 #(
		.INIT('h4)
	) name3723 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001 ,
		_w7770_
	);
	LUT2 #(
		.INIT('h8)
	) name3724 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001 ,
		_w7771_
	);
	LUT2 #(
		.INIT('h1)
	) name3725 (
		_w7770_,
		_w7771_,
		_w7772_
	);
	LUT2 #(
		.INIT('h2)
	) name3726 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w7772_,
		_w7773_
	);
	LUT2 #(
		.INIT('h4)
	) name3727 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001 ,
		_w7774_
	);
	LUT2 #(
		.INIT('h8)
	) name3728 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001 ,
		_w7775_
	);
	LUT2 #(
		.INIT('h1)
	) name3729 (
		_w7774_,
		_w7775_,
		_w7776_
	);
	LUT2 #(
		.INIT('h2)
	) name3730 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w7776_,
		_w7777_
	);
	LUT2 #(
		.INIT('h4)
	) name3731 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001 ,
		_w7778_
	);
	LUT2 #(
		.INIT('h8)
	) name3732 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001 ,
		_w7779_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		_w7778_,
		_w7779_,
		_w7780_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w7780_,
		_w7781_
	);
	LUT2 #(
		.INIT('h4)
	) name3735 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001 ,
		_w7782_
	);
	LUT2 #(
		.INIT('h8)
	) name3736 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001 ,
		_w7783_
	);
	LUT2 #(
		.INIT('h1)
	) name3737 (
		_w7782_,
		_w7783_,
		_w7784_
	);
	LUT2 #(
		.INIT('h2)
	) name3738 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w7784_,
		_w7785_
	);
	LUT2 #(
		.INIT('h1)
	) name3739 (
		_w7769_,
		_w7773_,
		_w7786_
	);
	LUT2 #(
		.INIT('h1)
	) name3740 (
		_w7777_,
		_w7781_,
		_w7787_
	);
	LUT2 #(
		.INIT('h4)
	) name3741 (
		_w7785_,
		_w7787_,
		_w7788_
	);
	LUT2 #(
		.INIT('h8)
	) name3742 (
		_w7786_,
		_w7788_,
		_w7789_
	);
	LUT2 #(
		.INIT('h2)
	) name3743 (
		_w7093_,
		_w7789_,
		_w7790_
	);
	LUT2 #(
		.INIT('h2)
	) name3744 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w7216_,
		_w7791_
	);
	LUT2 #(
		.INIT('h8)
	) name3745 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w7792_
	);
	LUT2 #(
		.INIT('h8)
	) name3746 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w7793_
	);
	LUT2 #(
		.INIT('h2)
	) name3747 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4276_,
		_w7794_
	);
	LUT2 #(
		.INIT('h1)
	) name3748 (
		_w7792_,
		_w7793_,
		_w7795_
	);
	LUT2 #(
		.INIT('h4)
	) name3749 (
		_w7791_,
		_w7795_,
		_w7796_
	);
	LUT2 #(
		.INIT('h4)
	) name3750 (
		_w7794_,
		_w7796_,
		_w7797_
	);
	LUT2 #(
		.INIT('h2)
	) name3751 (
		_w7215_,
		_w7797_,
		_w7798_
	);
	LUT2 #(
		.INIT('h4)
	) name3752 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 ,
		_w7799_
	);
	LUT2 #(
		.INIT('h8)
	) name3753 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 ,
		_w7800_
	);
	LUT2 #(
		.INIT('h1)
	) name3754 (
		_w7799_,
		_w7800_,
		_w7801_
	);
	LUT2 #(
		.INIT('h2)
	) name3755 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w7801_,
		_w7802_
	);
	LUT2 #(
		.INIT('h4)
	) name3756 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001 ,
		_w7803_
	);
	LUT2 #(
		.INIT('h8)
	) name3757 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001 ,
		_w7804_
	);
	LUT2 #(
		.INIT('h1)
	) name3758 (
		_w7803_,
		_w7804_,
		_w7805_
	);
	LUT2 #(
		.INIT('h2)
	) name3759 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w7805_,
		_w7806_
	);
	LUT2 #(
		.INIT('h4)
	) name3760 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 ,
		_w7807_
	);
	LUT2 #(
		.INIT('h8)
	) name3761 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 ,
		_w7808_
	);
	LUT2 #(
		.INIT('h1)
	) name3762 (
		_w7807_,
		_w7808_,
		_w7809_
	);
	LUT2 #(
		.INIT('h2)
	) name3763 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w7809_,
		_w7810_
	);
	LUT2 #(
		.INIT('h1)
	) name3764 (
		_w7802_,
		_w7806_,
		_w7811_
	);
	LUT2 #(
		.INIT('h4)
	) name3765 (
		_w7810_,
		_w7811_,
		_w7812_
	);
	LUT2 #(
		.INIT('h8)
	) name3766 (
		_w7174_,
		_w7812_,
		_w7813_
	);
	LUT2 #(
		.INIT('h2)
	) name3767 (
		_w7153_,
		_w7813_,
		_w7814_
	);
	LUT2 #(
		.INIT('h8)
	) name3768 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[10]/P0001 ,
		_w7815_
	);
	LUT2 #(
		.INIT('h8)
	) name3769 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[10]/P0001 ,
		_w7816_
	);
	LUT2 #(
		.INIT('h8)
	) name3770 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[10]/P0001 ,
		_w7817_
	);
	LUT2 #(
		.INIT('h8)
	) name3771 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[10]/P0001 ,
		_w7818_
	);
	LUT2 #(
		.INIT('h1)
	) name3772 (
		_w7815_,
		_w7816_,
		_w7819_
	);
	LUT2 #(
		.INIT('h1)
	) name3773 (
		_w7817_,
		_w7818_,
		_w7820_
	);
	LUT2 #(
		.INIT('h8)
	) name3774 (
		_w7819_,
		_w7820_,
		_w7821_
	);
	LUT2 #(
		.INIT('h2)
	) name3775 (
		_w7119_,
		_w7821_,
		_w7822_
	);
	LUT2 #(
		.INIT('h8)
	) name3776 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		_w7823_
	);
	LUT2 #(
		.INIT('h8)
	) name3777 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131 ,
		_w7824_
	);
	LUT2 #(
		.INIT('h8)
	) name3778 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131 ,
		_w7825_
	);
	LUT2 #(
		.INIT('h8)
	) name3779 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131 ,
		_w7826_
	);
	LUT2 #(
		.INIT('h8)
	) name3780 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131 ,
		_w7827_
	);
	LUT2 #(
		.INIT('h8)
	) name3781 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131 ,
		_w7828_
	);
	LUT2 #(
		.INIT('h8)
	) name3782 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 ,
		_w7829_
	);
	LUT2 #(
		.INIT('h8)
	) name3783 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131 ,
		_w7830_
	);
	LUT2 #(
		.INIT('h8)
	) name3784 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131 ,
		_w7831_
	);
	LUT2 #(
		.INIT('h8)
	) name3785 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131 ,
		_w7832_
	);
	LUT2 #(
		.INIT('h8)
	) name3786 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 ,
		_w7833_
	);
	LUT2 #(
		.INIT('h8)
	) name3787 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w7834_
	);
	LUT2 #(
		.INIT('h1)
	) name3788 (
		_w7823_,
		_w7824_,
		_w7835_
	);
	LUT2 #(
		.INIT('h1)
	) name3789 (
		_w7825_,
		_w7826_,
		_w7836_
	);
	LUT2 #(
		.INIT('h1)
	) name3790 (
		_w7827_,
		_w7828_,
		_w7837_
	);
	LUT2 #(
		.INIT('h1)
	) name3791 (
		_w7829_,
		_w7830_,
		_w7838_
	);
	LUT2 #(
		.INIT('h1)
	) name3792 (
		_w7831_,
		_w7832_,
		_w7839_
	);
	LUT2 #(
		.INIT('h1)
	) name3793 (
		_w7833_,
		_w7834_,
		_w7840_
	);
	LUT2 #(
		.INIT('h8)
	) name3794 (
		_w7839_,
		_w7840_,
		_w7841_
	);
	LUT2 #(
		.INIT('h8)
	) name3795 (
		_w7837_,
		_w7838_,
		_w7842_
	);
	LUT2 #(
		.INIT('h8)
	) name3796 (
		_w7835_,
		_w7836_,
		_w7843_
	);
	LUT2 #(
		.INIT('h8)
	) name3797 (
		_w7842_,
		_w7843_,
		_w7844_
	);
	LUT2 #(
		.INIT('h8)
	) name3798 (
		_w7841_,
		_w7844_,
		_w7845_
	);
	LUT2 #(
		.INIT('h2)
	) name3799 (
		_w7128_,
		_w7845_,
		_w7846_
	);
	LUT2 #(
		.INIT('h1)
	) name3800 (
		_w7688_,
		_w7822_,
		_w7847_
	);
	LUT2 #(
		.INIT('h4)
	) name3801 (
		_w7846_,
		_w7847_,
		_w7848_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w7765_,
		_w7790_,
		_w7849_
	);
	LUT2 #(
		.INIT('h4)
	) name3803 (
		_w7814_,
		_w7849_,
		_w7850_
	);
	LUT2 #(
		.INIT('h8)
	) name3804 (
		_w7848_,
		_w7850_,
		_w7851_
	);
	LUT2 #(
		.INIT('h4)
	) name3805 (
		_w7798_,
		_w7851_,
		_w7852_
	);
	LUT2 #(
		.INIT('h4)
	) name3806 (
		_w7734_,
		_w7852_,
		_w7853_
	);
	LUT2 #(
		.INIT('h4)
	) name3807 (
		_w7664_,
		_w7853_,
		_w7854_
	);
	LUT2 #(
		.INIT('h1)
	) name3808 (
		\emc_DMDoe_reg/NET0131 ,
		_w7854_,
		_w7855_
	);
	LUT2 #(
		.INIT('h8)
	) name3809 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[10]/P0001 ,
		_w7856_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		_w7057_,
		_w7856_,
		_w7857_
	);
	LUT2 #(
		.INIT('h4)
	) name3811 (
		_w7855_,
		_w7857_,
		_w7858_
	);
	LUT2 #(
		.INIT('h1)
	) name3812 (
		_w7663_,
		_w7858_,
		_w7859_
	);
	LUT2 #(
		.INIT('h2)
	) name3813 (
		_w6135_,
		_w7859_,
		_w7860_
	);
	LUT2 #(
		.INIT('h2)
	) name3814 (
		_w6176_,
		_w7860_,
		_w7861_
	);
	LUT2 #(
		.INIT('h4)
	) name3815 (
		_w7645_,
		_w7861_,
		_w7862_
	);
	LUT2 #(
		.INIT('h1)
	) name3816 (
		_w6135_,
		_w6176_,
		_w7863_
	);
	LUT2 #(
		.INIT('h8)
	) name3817 (
		\DM_rdm[3]_pad ,
		_w7016_,
		_w7864_
	);
	LUT2 #(
		.INIT('h8)
	) name3818 (
		\DM_rd1[3]_pad ,
		_w7022_,
		_w7865_
	);
	LUT2 #(
		.INIT('h8)
	) name3819 (
		\DM_rd4[3]_pad ,
		_w7028_,
		_w7866_
	);
	LUT2 #(
		.INIT('h8)
	) name3820 (
		\DM_rd6[3]_pad ,
		_w7031_,
		_w7867_
	);
	LUT2 #(
		.INIT('h8)
	) name3821 (
		\DM_rd7[3]_pad ,
		_w7034_,
		_w7868_
	);
	LUT2 #(
		.INIT('h8)
	) name3822 (
		\DM_rd3[3]_pad ,
		_w7038_,
		_w7869_
	);
	LUT2 #(
		.INIT('h2)
	) name3823 (
		\DM_rd0[3]_pad ,
		_w7053_,
		_w7870_
	);
	LUT2 #(
		.INIT('h8)
	) name3824 (
		\DM_rd5[3]_pad ,
		_w7043_,
		_w7871_
	);
	LUT2 #(
		.INIT('h8)
	) name3825 (
		\DM_rd2[3]_pad ,
		_w7041_,
		_w7872_
	);
	LUT2 #(
		.INIT('h1)
	) name3826 (
		_w7865_,
		_w7869_,
		_w7873_
	);
	LUT2 #(
		.INIT('h4)
	) name3827 (
		_w7872_,
		_w7873_,
		_w7874_
	);
	LUT2 #(
		.INIT('h1)
	) name3828 (
		_w7057_,
		_w7864_,
		_w7875_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		_w7867_,
		_w7868_,
		_w7876_
	);
	LUT2 #(
		.INIT('h8)
	) name3830 (
		_w7875_,
		_w7876_,
		_w7877_
	);
	LUT2 #(
		.INIT('h4)
	) name3831 (
		_w7866_,
		_w7874_,
		_w7878_
	);
	LUT2 #(
		.INIT('h4)
	) name3832 (
		_w7871_,
		_w7878_,
		_w7879_
	);
	LUT2 #(
		.INIT('h8)
	) name3833 (
		_w7877_,
		_w7879_,
		_w7880_
	);
	LUT2 #(
		.INIT('h4)
	) name3834 (
		_w7870_,
		_w7880_,
		_w7881_
	);
	LUT2 #(
		.INIT('h8)
	) name3835 (
		\regout_STD_C_reg[3]/P0001 ,
		_w6988_,
		_w7882_
	);
	LUT2 #(
		.INIT('h4)
	) name3836 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001 ,
		_w7883_
	);
	LUT2 #(
		.INIT('h8)
	) name3837 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 ,
		_w7884_
	);
	LUT2 #(
		.INIT('h1)
	) name3838 (
		_w7883_,
		_w7884_,
		_w7885_
	);
	LUT2 #(
		.INIT('h2)
	) name3839 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w7885_,
		_w7886_
	);
	LUT2 #(
		.INIT('h4)
	) name3840 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001 ,
		_w7887_
	);
	LUT2 #(
		.INIT('h8)
	) name3841 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001 ,
		_w7888_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		_w7887_,
		_w7888_,
		_w7889_
	);
	LUT2 #(
		.INIT('h2)
	) name3843 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w7889_,
		_w7890_
	);
	LUT2 #(
		.INIT('h4)
	) name3844 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001 ,
		_w7891_
	);
	LUT2 #(
		.INIT('h8)
	) name3845 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001 ,
		_w7892_
	);
	LUT2 #(
		.INIT('h1)
	) name3846 (
		_w7891_,
		_w7892_,
		_w7893_
	);
	LUT2 #(
		.INIT('h2)
	) name3847 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w7893_,
		_w7894_
	);
	LUT2 #(
		.INIT('h4)
	) name3848 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001 ,
		_w7895_
	);
	LUT2 #(
		.INIT('h8)
	) name3849 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001 ,
		_w7896_
	);
	LUT2 #(
		.INIT('h1)
	) name3850 (
		_w7895_,
		_w7896_,
		_w7897_
	);
	LUT2 #(
		.INIT('h2)
	) name3851 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w7897_,
		_w7898_
	);
	LUT2 #(
		.INIT('h4)
	) name3852 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001 ,
		_w7899_
	);
	LUT2 #(
		.INIT('h8)
	) name3853 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001 ,
		_w7900_
	);
	LUT2 #(
		.INIT('h1)
	) name3854 (
		_w7899_,
		_w7900_,
		_w7901_
	);
	LUT2 #(
		.INIT('h2)
	) name3855 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w7901_,
		_w7902_
	);
	LUT2 #(
		.INIT('h4)
	) name3856 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 ,
		_w7903_
	);
	LUT2 #(
		.INIT('h8)
	) name3857 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 ,
		_w7904_
	);
	LUT2 #(
		.INIT('h1)
	) name3858 (
		_w7903_,
		_w7904_,
		_w7905_
	);
	LUT2 #(
		.INIT('h2)
	) name3859 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w7905_,
		_w7906_
	);
	LUT2 #(
		.INIT('h4)
	) name3860 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001 ,
		_w7907_
	);
	LUT2 #(
		.INIT('h8)
	) name3861 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 ,
		_w7908_
	);
	LUT2 #(
		.INIT('h1)
	) name3862 (
		_w7907_,
		_w7908_,
		_w7909_
	);
	LUT2 #(
		.INIT('h2)
	) name3863 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w7909_,
		_w7910_
	);
	LUT2 #(
		.INIT('h1)
	) name3864 (
		_w7886_,
		_w7890_,
		_w7911_
	);
	LUT2 #(
		.INIT('h1)
	) name3865 (
		_w7894_,
		_w7898_,
		_w7912_
	);
	LUT2 #(
		.INIT('h1)
	) name3866 (
		_w7902_,
		_w7906_,
		_w7913_
	);
	LUT2 #(
		.INIT('h4)
	) name3867 (
		_w7910_,
		_w7913_,
		_w7914_
	);
	LUT2 #(
		.INIT('h8)
	) name3868 (
		_w7911_,
		_w7912_,
		_w7915_
	);
	LUT2 #(
		.INIT('h8)
	) name3869 (
		_w7914_,
		_w7915_,
		_w7916_
	);
	LUT2 #(
		.INIT('h2)
	) name3870 (
		_w7179_,
		_w7916_,
		_w7917_
	);
	LUT2 #(
		.INIT('h8)
	) name3871 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 ,
		_w7918_
	);
	LUT2 #(
		.INIT('h8)
	) name3872 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		_w7919_
	);
	LUT2 #(
		.INIT('h8)
	) name3873 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 ,
		_w7920_
	);
	LUT2 #(
		.INIT('h8)
	) name3874 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w7921_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131 ,
		_w7922_
	);
	LUT2 #(
		.INIT('h8)
	) name3876 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131 ,
		_w7923_
	);
	LUT2 #(
		.INIT('h8)
	) name3877 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131 ,
		_w7924_
	);
	LUT2 #(
		.INIT('h8)
	) name3878 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131 ,
		_w7925_
	);
	LUT2 #(
		.INIT('h8)
	) name3879 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131 ,
		_w7926_
	);
	LUT2 #(
		.INIT('h8)
	) name3880 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131 ,
		_w7927_
	);
	LUT2 #(
		.INIT('h8)
	) name3881 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131 ,
		_w7928_
	);
	LUT2 #(
		.INIT('h8)
	) name3882 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131 ,
		_w7929_
	);
	LUT2 #(
		.INIT('h1)
	) name3883 (
		_w7918_,
		_w7919_,
		_w7930_
	);
	LUT2 #(
		.INIT('h1)
	) name3884 (
		_w7920_,
		_w7921_,
		_w7931_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		_w7922_,
		_w7923_,
		_w7932_
	);
	LUT2 #(
		.INIT('h1)
	) name3886 (
		_w7924_,
		_w7925_,
		_w7933_
	);
	LUT2 #(
		.INIT('h1)
	) name3887 (
		_w7926_,
		_w7927_,
		_w7934_
	);
	LUT2 #(
		.INIT('h1)
	) name3888 (
		_w7928_,
		_w7929_,
		_w7935_
	);
	LUT2 #(
		.INIT('h8)
	) name3889 (
		_w7934_,
		_w7935_,
		_w7936_
	);
	LUT2 #(
		.INIT('h8)
	) name3890 (
		_w7932_,
		_w7933_,
		_w7937_
	);
	LUT2 #(
		.INIT('h8)
	) name3891 (
		_w7930_,
		_w7931_,
		_w7938_
	);
	LUT2 #(
		.INIT('h8)
	) name3892 (
		_w7937_,
		_w7938_,
		_w7939_
	);
	LUT2 #(
		.INIT('h8)
	) name3893 (
		_w7936_,
		_w7939_,
		_w7940_
	);
	LUT2 #(
		.INIT('h2)
	) name3894 (
		_w7068_,
		_w7940_,
		_w7941_
	);
	LUT2 #(
		.INIT('h4)
	) name3895 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001 ,
		_w7942_
	);
	LUT2 #(
		.INIT('h8)
	) name3896 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001 ,
		_w7943_
	);
	LUT2 #(
		.INIT('h1)
	) name3897 (
		_w7942_,
		_w7943_,
		_w7944_
	);
	LUT2 #(
		.INIT('h2)
	) name3898 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w7944_,
		_w7945_
	);
	LUT2 #(
		.INIT('h4)
	) name3899 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001 ,
		_w7946_
	);
	LUT2 #(
		.INIT('h8)
	) name3900 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001 ,
		_w7947_
	);
	LUT2 #(
		.INIT('h1)
	) name3901 (
		_w7946_,
		_w7947_,
		_w7948_
	);
	LUT2 #(
		.INIT('h2)
	) name3902 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w7948_,
		_w7949_
	);
	LUT2 #(
		.INIT('h4)
	) name3903 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001 ,
		_w7950_
	);
	LUT2 #(
		.INIT('h8)
	) name3904 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001 ,
		_w7951_
	);
	LUT2 #(
		.INIT('h1)
	) name3905 (
		_w7950_,
		_w7951_,
		_w7952_
	);
	LUT2 #(
		.INIT('h2)
	) name3906 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w7952_,
		_w7953_
	);
	LUT2 #(
		.INIT('h4)
	) name3907 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001 ,
		_w7954_
	);
	LUT2 #(
		.INIT('h8)
	) name3908 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001 ,
		_w7955_
	);
	LUT2 #(
		.INIT('h1)
	) name3909 (
		_w7954_,
		_w7955_,
		_w7956_
	);
	LUT2 #(
		.INIT('h2)
	) name3910 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w7956_,
		_w7957_
	);
	LUT2 #(
		.INIT('h4)
	) name3911 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001 ,
		_w7958_
	);
	LUT2 #(
		.INIT('h8)
	) name3912 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001 ,
		_w7959_
	);
	LUT2 #(
		.INIT('h1)
	) name3913 (
		_w7958_,
		_w7959_,
		_w7960_
	);
	LUT2 #(
		.INIT('h2)
	) name3914 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w7960_,
		_w7961_
	);
	LUT2 #(
		.INIT('h8)
	) name3915 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w7962_
	);
	LUT2 #(
		.INIT('h1)
	) name3916 (
		_w7945_,
		_w7962_,
		_w7963_
	);
	LUT2 #(
		.INIT('h1)
	) name3917 (
		_w7949_,
		_w7953_,
		_w7964_
	);
	LUT2 #(
		.INIT('h1)
	) name3918 (
		_w7957_,
		_w7961_,
		_w7965_
	);
	LUT2 #(
		.INIT('h8)
	) name3919 (
		_w7964_,
		_w7965_,
		_w7966_
	);
	LUT2 #(
		.INIT('h8)
	) name3920 (
		_w7963_,
		_w7966_,
		_w7967_
	);
	LUT2 #(
		.INIT('h2)
	) name3921 (
		_w7093_,
		_w7967_,
		_w7968_
	);
	LUT2 #(
		.INIT('h8)
	) name3922 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[3]/P0001 ,
		_w7969_
	);
	LUT2 #(
		.INIT('h8)
	) name3923 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w7970_
	);
	LUT2 #(
		.INIT('h8)
	) name3924 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[3]/P0001 ,
		_w7971_
	);
	LUT2 #(
		.INIT('h8)
	) name3925 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		_w7972_
	);
	LUT2 #(
		.INIT('h1)
	) name3926 (
		_w7969_,
		_w7970_,
		_w7973_
	);
	LUT2 #(
		.INIT('h1)
	) name3927 (
		_w7971_,
		_w7972_,
		_w7974_
	);
	LUT2 #(
		.INIT('h8)
	) name3928 (
		_w7973_,
		_w7974_,
		_w7975_
	);
	LUT2 #(
		.INIT('h2)
	) name3929 (
		_w7119_,
		_w7975_,
		_w7976_
	);
	LUT2 #(
		.INIT('h4)
	) name3930 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001 ,
		_w7977_
	);
	LUT2 #(
		.INIT('h8)
	) name3931 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001 ,
		_w7978_
	);
	LUT2 #(
		.INIT('h1)
	) name3932 (
		_w7977_,
		_w7978_,
		_w7979_
	);
	LUT2 #(
		.INIT('h2)
	) name3933 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w7979_,
		_w7980_
	);
	LUT2 #(
		.INIT('h4)
	) name3934 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[3]/P0001 ,
		_w7981_
	);
	LUT2 #(
		.INIT('h8)
	) name3935 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBs_reg[3]/P0001 ,
		_w7982_
	);
	LUT2 #(
		.INIT('h1)
	) name3936 (
		_w7981_,
		_w7982_,
		_w7983_
	);
	LUT2 #(
		.INIT('h2)
	) name3937 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		_w7983_,
		_w7984_
	);
	LUT2 #(
		.INIT('h4)
	) name3938 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 ,
		_w7985_
	);
	LUT2 #(
		.INIT('h8)
	) name3939 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 ,
		_w7986_
	);
	LUT2 #(
		.INIT('h1)
	) name3940 (
		_w7985_,
		_w7986_,
		_w7987_
	);
	LUT2 #(
		.INIT('h2)
	) name3941 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w7987_,
		_w7988_
	);
	LUT2 #(
		.INIT('h4)
	) name3942 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 ,
		_w7989_
	);
	LUT2 #(
		.INIT('h8)
	) name3943 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 ,
		_w7990_
	);
	LUT2 #(
		.INIT('h1)
	) name3944 (
		_w7989_,
		_w7990_,
		_w7991_
	);
	LUT2 #(
		.INIT('h2)
	) name3945 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w7991_,
		_w7992_
	);
	LUT2 #(
		.INIT('h4)
	) name3946 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001 ,
		_w7993_
	);
	LUT2 #(
		.INIT('h8)
	) name3947 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001 ,
		_w7994_
	);
	LUT2 #(
		.INIT('h1)
	) name3948 (
		_w7993_,
		_w7994_,
		_w7995_
	);
	LUT2 #(
		.INIT('h2)
	) name3949 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w7995_,
		_w7996_
	);
	LUT2 #(
		.INIT('h1)
	) name3950 (
		_w7980_,
		_w7984_,
		_w7997_
	);
	LUT2 #(
		.INIT('h1)
	) name3951 (
		_w7988_,
		_w7992_,
		_w7998_
	);
	LUT2 #(
		.INIT('h4)
	) name3952 (
		_w7996_,
		_w7998_,
		_w7999_
	);
	LUT2 #(
		.INIT('h8)
	) name3953 (
		_w7997_,
		_w7999_,
		_w8000_
	);
	LUT2 #(
		.INIT('h2)
	) name3954 (
		_w7153_,
		_w8000_,
		_w8001_
	);
	LUT2 #(
		.INIT('h8)
	) name3955 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131 ,
		_w8002_
	);
	LUT2 #(
		.INIT('h8)
	) name3956 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w8003_
	);
	LUT2 #(
		.INIT('h8)
	) name3957 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131 ,
		_w8004_
	);
	LUT2 #(
		.INIT('h8)
	) name3958 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131 ,
		_w8005_
	);
	LUT2 #(
		.INIT('h8)
	) name3959 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		_w8006_
	);
	LUT2 #(
		.INIT('h8)
	) name3960 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w8007_
	);
	LUT2 #(
		.INIT('h8)
	) name3961 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131 ,
		_w8008_
	);
	LUT2 #(
		.INIT('h8)
	) name3962 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131 ,
		_w8009_
	);
	LUT2 #(
		.INIT('h8)
	) name3963 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w8010_
	);
	LUT2 #(
		.INIT('h8)
	) name3964 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131 ,
		_w8011_
	);
	LUT2 #(
		.INIT('h8)
	) name3965 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131 ,
		_w8012_
	);
	LUT2 #(
		.INIT('h8)
	) name3966 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131 ,
		_w8013_
	);
	LUT2 #(
		.INIT('h1)
	) name3967 (
		_w8002_,
		_w8003_,
		_w8014_
	);
	LUT2 #(
		.INIT('h1)
	) name3968 (
		_w8004_,
		_w8005_,
		_w8015_
	);
	LUT2 #(
		.INIT('h1)
	) name3969 (
		_w8006_,
		_w8007_,
		_w8016_
	);
	LUT2 #(
		.INIT('h1)
	) name3970 (
		_w8008_,
		_w8009_,
		_w8017_
	);
	LUT2 #(
		.INIT('h1)
	) name3971 (
		_w8010_,
		_w8011_,
		_w8018_
	);
	LUT2 #(
		.INIT('h1)
	) name3972 (
		_w8012_,
		_w8013_,
		_w8019_
	);
	LUT2 #(
		.INIT('h8)
	) name3973 (
		_w8018_,
		_w8019_,
		_w8020_
	);
	LUT2 #(
		.INIT('h8)
	) name3974 (
		_w8016_,
		_w8017_,
		_w8021_
	);
	LUT2 #(
		.INIT('h8)
	) name3975 (
		_w8014_,
		_w8015_,
		_w8022_
	);
	LUT2 #(
		.INIT('h8)
	) name3976 (
		_w8021_,
		_w8022_,
		_w8023_
	);
	LUT2 #(
		.INIT('h8)
	) name3977 (
		_w8020_,
		_w8023_,
		_w8024_
	);
	LUT2 #(
		.INIT('h2)
	) name3978 (
		_w7128_,
		_w8024_,
		_w8025_
	);
	LUT2 #(
		.INIT('h8)
	) name3979 (
		\idma_DOVL_reg[3]/NET0131 ,
		_w7532_,
		_w8026_
	);
	LUT2 #(
		.INIT('h8)
	) name3980 (
		\sport0_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w7295_,
		_w8027_
	);
	LUT2 #(
		.INIT('h8)
	) name3981 (
		\tm_tpr_reg_DO_reg[3]/NET0131 ,
		_w7293_,
		_w8028_
	);
	LUT2 #(
		.INIT('h8)
	) name3982 (
		\bdma_BWCOUNT_reg[3]/NET0131 ,
		_w7287_,
		_w8029_
	);
	LUT2 #(
		.INIT('h8)
	) name3983 (
		\emc_WSCRreg_DO_reg[3]/NET0131 ,
		_w7251_,
		_w8030_
	);
	LUT2 #(
		.INIT('h8)
	) name3984 (
		\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w7256_,
		_w8031_
	);
	LUT2 #(
		.INIT('h8)
	) name3985 (
		\sport1_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w7263_,
		_w8032_
	);
	LUT2 #(
		.INIT('h8)
	) name3986 (
		\tm_tsr_reg_DO_reg[3]/NET0131 ,
		_w7540_,
		_w8033_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w7249_,
		_w8034_
	);
	LUT2 #(
		.INIT('h8)
	) name3988 (
		\emc_WSCRext_reg_DO_reg[3]/NET0131 ,
		_w7514_,
		_w8035_
	);
	LUT2 #(
		.INIT('h8)
	) name3989 (
		\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w7247_,
		_w8036_
	);
	LUT2 #(
		.INIT('h8)
	) name3990 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w7281_,
		_w8037_
	);
	LUT2 #(
		.INIT('h8)
	) name3991 (
		\pio_pmask_reg_DO_reg[3]/NET0131 ,
		_w7297_,
		_w8038_
	);
	LUT2 #(
		.INIT('h8)
	) name3992 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w7234_,
		_w8039_
	);
	LUT2 #(
		.INIT('h8)
	) name3993 (
		\sport0_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w7276_,
		_w8040_
	);
	LUT2 #(
		.INIT('h8)
	) name3994 (
		\sport1_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w7527_,
		_w8041_
	);
	LUT2 #(
		.INIT('h8)
	) name3995 (
		\tm_TCR_TMP_reg[3]/NET0131 ,
		_w7289_,
		_w8042_
	);
	LUT2 #(
		.INIT('h8)
	) name3996 (
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w7259_,
		_w8043_
	);
	LUT2 #(
		.INIT('h8)
	) name3997 (
		\bdma_BOVL_reg[3]/NET0131 ,
		_w7534_,
		_w8044_
	);
	LUT2 #(
		.INIT('h8)
	) name3998 (
		\clkc_ckr_reg_DO_reg[3]/NET0131 ,
		_w7239_,
		_w8045_
	);
	LUT2 #(
		.INIT('h8)
	) name3999 (
		\memc_usysr_DO_reg[3]/NET0131 ,
		_w7301_,
		_w8046_
	);
	LUT2 #(
		.INIT('h8)
	) name4000 (
		\bdma_BEAD_reg[3]/NET0131 ,
		_w7303_,
		_w8047_
	);
	LUT2 #(
		.INIT('h8)
	) name4001 (
		\bdma_BCTL_reg[3]/NET0131 ,
		_w7230_,
		_w8048_
	);
	LUT2 #(
		.INIT('h8)
	) name4002 (
		\pio_PINT_reg[3]/NET0131 ,
		_w7271_,
		_w8049_
	);
	LUT2 #(
		.INIT('h8)
	) name4003 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w7299_,
		_w8050_
	);
	LUT2 #(
		.INIT('h8)
	) name4004 (
		\PIO_out[3]_pad ,
		_w7291_,
		_w8051_
	);
	LUT2 #(
		.INIT('h8)
	) name4005 (
		\PIO_oe[3]_pad ,
		_w7244_,
		_w8052_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w7273_,
		_w8053_
	);
	LUT2 #(
		.INIT('h1)
	) name4007 (
		_w7522_,
		_w8026_,
		_w8054_
	);
	LUT2 #(
		.INIT('h1)
	) name4008 (
		_w8027_,
		_w8028_,
		_w8055_
	);
	LUT2 #(
		.INIT('h1)
	) name4009 (
		_w8030_,
		_w8031_,
		_w8056_
	);
	LUT2 #(
		.INIT('h1)
	) name4010 (
		_w8032_,
		_w8033_,
		_w8057_
	);
	LUT2 #(
		.INIT('h1)
	) name4011 (
		_w8034_,
		_w8035_,
		_w8058_
	);
	LUT2 #(
		.INIT('h1)
	) name4012 (
		_w8036_,
		_w8037_,
		_w8059_
	);
	LUT2 #(
		.INIT('h1)
	) name4013 (
		_w8038_,
		_w8040_,
		_w8060_
	);
	LUT2 #(
		.INIT('h1)
	) name4014 (
		_w8041_,
		_w8042_,
		_w8061_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w8043_,
		_w8045_,
		_w8062_
	);
	LUT2 #(
		.INIT('h1)
	) name4016 (
		_w8046_,
		_w8049_,
		_w8063_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		_w8050_,
		_w8051_,
		_w8064_
	);
	LUT2 #(
		.INIT('h1)
	) name4018 (
		_w8052_,
		_w8053_,
		_w8065_
	);
	LUT2 #(
		.INIT('h8)
	) name4019 (
		_w8064_,
		_w8065_,
		_w8066_
	);
	LUT2 #(
		.INIT('h8)
	) name4020 (
		_w8062_,
		_w8063_,
		_w8067_
	);
	LUT2 #(
		.INIT('h8)
	) name4021 (
		_w8060_,
		_w8061_,
		_w8068_
	);
	LUT2 #(
		.INIT('h8)
	) name4022 (
		_w8058_,
		_w8059_,
		_w8069_
	);
	LUT2 #(
		.INIT('h8)
	) name4023 (
		_w8056_,
		_w8057_,
		_w8070_
	);
	LUT2 #(
		.INIT('h8)
	) name4024 (
		_w8054_,
		_w8055_,
		_w8071_
	);
	LUT2 #(
		.INIT('h8)
	) name4025 (
		_w8070_,
		_w8071_,
		_w8072_
	);
	LUT2 #(
		.INIT('h8)
	) name4026 (
		_w8068_,
		_w8069_,
		_w8073_
	);
	LUT2 #(
		.INIT('h8)
	) name4027 (
		_w8066_,
		_w8067_,
		_w8074_
	);
	LUT2 #(
		.INIT('h8)
	) name4028 (
		_w8073_,
		_w8074_,
		_w8075_
	);
	LUT2 #(
		.INIT('h4)
	) name4029 (
		_w8039_,
		_w8072_,
		_w8076_
	);
	LUT2 #(
		.INIT('h1)
	) name4030 (
		_w8047_,
		_w8048_,
		_w8077_
	);
	LUT2 #(
		.INIT('h8)
	) name4031 (
		_w8076_,
		_w8077_,
		_w8078_
	);
	LUT2 #(
		.INIT('h4)
	) name4032 (
		_w8029_,
		_w8075_,
		_w8079_
	);
	LUT2 #(
		.INIT('h4)
	) name4033 (
		_w8044_,
		_w8079_,
		_w8080_
	);
	LUT2 #(
		.INIT('h8)
	) name4034 (
		_w8078_,
		_w8080_,
		_w8081_
	);
	LUT2 #(
		.INIT('h2)
	) name4035 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w8081_,
		_w8082_
	);
	LUT2 #(
		.INIT('h8)
	) name4036 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w8083_
	);
	LUT2 #(
		.INIT('h2)
	) name4037 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w7216_,
		_w8084_
	);
	LUT2 #(
		.INIT('h8)
	) name4038 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[3]/NET0131 ,
		_w8085_
	);
	LUT2 #(
		.INIT('h2)
	) name4039 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4328_,
		_w8086_
	);
	LUT2 #(
		.INIT('h8)
	) name4040 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		_w8087_
	);
	LUT2 #(
		.INIT('h8)
	) name4041 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w8088_
	);
	LUT2 #(
		.INIT('h8)
	) name4042 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w8089_
	);
	LUT2 #(
		.INIT('h8)
	) name4043 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w8090_
	);
	LUT2 #(
		.INIT('h8)
	) name4044 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w8091_
	);
	LUT2 #(
		.INIT('h1)
	) name4045 (
		_w8083_,
		_w8085_,
		_w8092_
	);
	LUT2 #(
		.INIT('h1)
	) name4046 (
		_w8087_,
		_w8088_,
		_w8093_
	);
	LUT2 #(
		.INIT('h1)
	) name4047 (
		_w8089_,
		_w8090_,
		_w8094_
	);
	LUT2 #(
		.INIT('h4)
	) name4048 (
		_w8091_,
		_w8094_,
		_w8095_
	);
	LUT2 #(
		.INIT('h8)
	) name4049 (
		_w8092_,
		_w8093_,
		_w8096_
	);
	LUT2 #(
		.INIT('h4)
	) name4050 (
		_w8084_,
		_w8096_,
		_w8097_
	);
	LUT2 #(
		.INIT('h8)
	) name4051 (
		_w8095_,
		_w8097_,
		_w8098_
	);
	LUT2 #(
		.INIT('h4)
	) name4052 (
		_w8086_,
		_w8098_,
		_w8099_
	);
	LUT2 #(
		.INIT('h2)
	) name4053 (
		_w7215_,
		_w8099_,
		_w8100_
	);
	LUT2 #(
		.INIT('h1)
	) name4054 (
		_w7941_,
		_w7976_,
		_w8101_
	);
	LUT2 #(
		.INIT('h4)
	) name4055 (
		_w8025_,
		_w8101_,
		_w8102_
	);
	LUT2 #(
		.INIT('h1)
	) name4056 (
		_w7917_,
		_w7968_,
		_w8103_
	);
	LUT2 #(
		.INIT('h4)
	) name4057 (
		_w8001_,
		_w8103_,
		_w8104_
	);
	LUT2 #(
		.INIT('h8)
	) name4058 (
		_w8102_,
		_w8104_,
		_w8105_
	);
	LUT2 #(
		.INIT('h4)
	) name4059 (
		_w8100_,
		_w8105_,
		_w8106_
	);
	LUT2 #(
		.INIT('h4)
	) name4060 (
		_w8082_,
		_w8106_,
		_w8107_
	);
	LUT2 #(
		.INIT('h4)
	) name4061 (
		_w7882_,
		_w8107_,
		_w8108_
	);
	LUT2 #(
		.INIT('h1)
	) name4062 (
		\emc_DMDoe_reg/NET0131 ,
		_w8108_,
		_w8109_
	);
	LUT2 #(
		.INIT('h8)
	) name4063 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[3]/P0001 ,
		_w8110_
	);
	LUT2 #(
		.INIT('h2)
	) name4064 (
		_w7057_,
		_w8110_,
		_w8111_
	);
	LUT2 #(
		.INIT('h4)
	) name4065 (
		_w8109_,
		_w8111_,
		_w8112_
	);
	LUT2 #(
		.INIT('h1)
	) name4066 (
		_w7881_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h8)
	) name4067 (
		_w7863_,
		_w8113_,
		_w8114_
	);
	LUT2 #(
		.INIT('h8)
	) name4068 (
		\core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 ,
		_w6972_,
		_w8115_
	);
	LUT2 #(
		.INIT('h8)
	) name4069 (
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		_w6976_,
		_w8116_
	);
	LUT2 #(
		.INIT('h8)
	) name4070 (
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w6974_,
		_w8117_
	);
	LUT2 #(
		.INIT('h8)
	) name4071 (
		\core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 ,
		_w6970_,
		_w8118_
	);
	LUT2 #(
		.INIT('h1)
	) name4072 (
		_w8115_,
		_w8116_,
		_w8119_
	);
	LUT2 #(
		.INIT('h1)
	) name4073 (
		_w8117_,
		_w8118_,
		_w8120_
	);
	LUT2 #(
		.INIT('h8)
	) name4074 (
		_w8119_,
		_w8120_,
		_w8121_
	);
	LUT2 #(
		.INIT('h2)
	) name4075 (
		_w4055_,
		_w8121_,
		_w8122_
	);
	LUT2 #(
		.INIT('h8)
	) name4076 (
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		_w6958_,
		_w8123_
	);
	LUT2 #(
		.INIT('h8)
	) name4077 (
		\core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 ,
		_w6960_,
		_w8124_
	);
	LUT2 #(
		.INIT('h8)
	) name4078 (
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w6962_,
		_w8125_
	);
	LUT2 #(
		.INIT('h8)
	) name4079 (
		\core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 ,
		_w6964_,
		_w8126_
	);
	LUT2 #(
		.INIT('h1)
	) name4080 (
		_w8123_,
		_w8124_,
		_w8127_
	);
	LUT2 #(
		.INIT('h1)
	) name4081 (
		_w8125_,
		_w8126_,
		_w8128_
	);
	LUT2 #(
		.INIT('h8)
	) name4082 (
		_w8127_,
		_w8128_,
		_w8129_
	);
	LUT2 #(
		.INIT('h4)
	) name4083 (
		_w8122_,
		_w8129_,
		_w8130_
	);
	LUT2 #(
		.INIT('h8)
	) name4084 (
		_w6058_,
		_w6060_,
		_w8131_
	);
	LUT2 #(
		.INIT('h8)
	) name4085 (
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w8131_,
		_w8132_
	);
	LUT2 #(
		.INIT('h8)
	) name4086 (
		\core_dag_ilm1reg_I2_we_DO_reg[10]/NET0131 ,
		_w6084_,
		_w8133_
	);
	LUT2 #(
		.INIT('h8)
	) name4087 (
		_w6085_,
		_w8133_,
		_w8134_
	);
	LUT2 #(
		.INIT('h8)
	) name4088 (
		\core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 ,
		_w6067_,
		_w8135_
	);
	LUT2 #(
		.INIT('h8)
	) name4089 (
		_w6068_,
		_w8135_,
		_w8136_
	);
	LUT2 #(
		.INIT('h8)
	) name4090 (
		\core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 ,
		_w6075_,
		_w8137_
	);
	LUT2 #(
		.INIT('h8)
	) name4091 (
		_w6077_,
		_w8137_,
		_w8138_
	);
	LUT2 #(
		.INIT('h1)
	) name4092 (
		_w4055_,
		_w8132_,
		_w8139_
	);
	LUT2 #(
		.INIT('h1)
	) name4093 (
		_w8134_,
		_w8136_,
		_w8140_
	);
	LUT2 #(
		.INIT('h4)
	) name4094 (
		_w8138_,
		_w8140_,
		_w8141_
	);
	LUT2 #(
		.INIT('h8)
	) name4095 (
		_w8139_,
		_w8141_,
		_w8142_
	);
	LUT2 #(
		.INIT('h8)
	) name4096 (
		_w6097_,
		_w8137_,
		_w8143_
	);
	LUT2 #(
		.INIT('h8)
	) name4097 (
		_w6095_,
		_w8133_,
		_w8144_
	);
	LUT2 #(
		.INIT('h8)
	) name4098 (
		_w6091_,
		_w8135_,
		_w8145_
	);
	LUT2 #(
		.INIT('h8)
	) name4099 (
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w6148_,
		_w8146_
	);
	LUT2 #(
		.INIT('h1)
	) name4100 (
		_w8143_,
		_w8144_,
		_w8147_
	);
	LUT2 #(
		.INIT('h1)
	) name4101 (
		_w8145_,
		_w8146_,
		_w8148_
	);
	LUT2 #(
		.INIT('h8)
	) name4102 (
		_w8147_,
		_w8148_,
		_w8149_
	);
	LUT2 #(
		.INIT('h8)
	) name4103 (
		_w4055_,
		_w8149_,
		_w8150_
	);
	LUT2 #(
		.INIT('h1)
	) name4104 (
		_w8142_,
		_w8150_,
		_w8151_
	);
	LUT2 #(
		.INIT('h2)
	) name4105 (
		_w8130_,
		_w8151_,
		_w8152_
	);
	LUT2 #(
		.INIT('h2)
	) name4106 (
		_w6135_,
		_w6176_,
		_w8153_
	);
	LUT2 #(
		.INIT('h4)
	) name4107 (
		_w8152_,
		_w8153_,
		_w8154_
	);
	LUT2 #(
		.INIT('h1)
	) name4108 (
		_w8114_,
		_w8154_,
		_w8155_
	);
	LUT2 #(
		.INIT('h4)
	) name4109 (
		_w7862_,
		_w8155_,
		_w8156_
	);
	LUT2 #(
		.INIT('h2)
	) name4110 (
		_w7005_,
		_w8156_,
		_w8157_
	);
	LUT2 #(
		.INIT('h1)
	) name4111 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w6924_,
		_w8158_
	);
	LUT2 #(
		.INIT('h8)
	) name4112 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w6926_,
		_w8159_
	);
	LUT2 #(
		.INIT('h8)
	) name4113 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131 ,
		_w6988_,
		_w8160_
	);
	LUT2 #(
		.INIT('h1)
	) name4114 (
		_w6121_,
		_w8130_,
		_w8161_
	);
	LUT2 #(
		.INIT('h8)
	) name4115 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w6956_,
		_w8162_
	);
	LUT2 #(
		.INIT('h4)
	) name4116 (
		_w6111_,
		_w8151_,
		_w8163_
	);
	LUT2 #(
		.INIT('h1)
	) name4117 (
		_w8161_,
		_w8162_,
		_w8164_
	);
	LUT2 #(
		.INIT('h4)
	) name4118 (
		_w8163_,
		_w8164_,
		_w8165_
	);
	LUT2 #(
		.INIT('h2)
	) name4119 (
		_w5949_,
		_w8165_,
		_w8166_
	);
	LUT2 #(
		.INIT('h2)
	) name4120 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w6934_,
		_w8167_
	);
	LUT2 #(
		.INIT('h1)
	) name4121 (
		_w8159_,
		_w8160_,
		_w8168_
	);
	LUT2 #(
		.INIT('h8)
	) name4122 (
		_w6924_,
		_w8168_,
		_w8169_
	);
	LUT2 #(
		.INIT('h4)
	) name4123 (
		_w8167_,
		_w8169_,
		_w8170_
	);
	LUT2 #(
		.INIT('h4)
	) name4124 (
		_w8166_,
		_w8170_,
		_w8171_
	);
	LUT2 #(
		.INIT('h1)
	) name4125 (
		_w6176_,
		_w8158_,
		_w8172_
	);
	LUT2 #(
		.INIT('h4)
	) name4126 (
		_w8171_,
		_w8172_,
		_w8173_
	);
	LUT2 #(
		.INIT('h8)
	) name4127 (
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		_w8131_,
		_w8174_
	);
	LUT2 #(
		.INIT('h8)
	) name4128 (
		\core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 ,
		_w6140_,
		_w8175_
	);
	LUT2 #(
		.INIT('h8)
	) name4129 (
		\core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 ,
		_w6142_,
		_w8176_
	);
	LUT2 #(
		.INIT('h8)
	) name4130 (
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w6084_,
		_w8177_
	);
	LUT2 #(
		.INIT('h8)
	) name4131 (
		_w6085_,
		_w8177_,
		_w8178_
	);
	LUT2 #(
		.INIT('h1)
	) name4132 (
		_w4055_,
		_w8174_,
		_w8179_
	);
	LUT2 #(
		.INIT('h1)
	) name4133 (
		_w8175_,
		_w8176_,
		_w8180_
	);
	LUT2 #(
		.INIT('h4)
	) name4134 (
		_w8178_,
		_w8180_,
		_w8181_
	);
	LUT2 #(
		.INIT('h8)
	) name4135 (
		_w8179_,
		_w8181_,
		_w8182_
	);
	LUT2 #(
		.INIT('h8)
	) name4136 (
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w6152_,
		_w8183_
	);
	LUT2 #(
		.INIT('h8)
	) name4137 (
		\core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 ,
		_w6150_,
		_w8184_
	);
	LUT2 #(
		.INIT('h8)
	) name4138 (
		\core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 ,
		_w6154_,
		_w8185_
	);
	LUT2 #(
		.INIT('h8)
	) name4139 (
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		_w6058_,
		_w8186_
	);
	LUT2 #(
		.INIT('h8)
	) name4140 (
		_w6093_,
		_w8186_,
		_w8187_
	);
	LUT2 #(
		.INIT('h1)
	) name4141 (
		_w8183_,
		_w8184_,
		_w8188_
	);
	LUT2 #(
		.INIT('h1)
	) name4142 (
		_w8185_,
		_w8187_,
		_w8189_
	);
	LUT2 #(
		.INIT('h8)
	) name4143 (
		_w8188_,
		_w8189_,
		_w8190_
	);
	LUT2 #(
		.INIT('h8)
	) name4144 (
		_w4055_,
		_w8190_,
		_w8191_
	);
	LUT2 #(
		.INIT('h1)
	) name4145 (
		_w8182_,
		_w8191_,
		_w8192_
	);
	LUT2 #(
		.INIT('h8)
	) name4146 (
		_w6176_,
		_w8192_,
		_w8193_
	);
	LUT2 #(
		.INIT('h1)
	) name4147 (
		_w6135_,
		_w8193_,
		_w8194_
	);
	LUT2 #(
		.INIT('h4)
	) name4148 (
		_w8173_,
		_w8194_,
		_w8195_
	);
	LUT2 #(
		.INIT('h2)
	) name4149 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		_w6620_,
		_w8196_
	);
	LUT2 #(
		.INIT('h1)
	) name4150 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6905_,
		_w8197_
	);
	LUT2 #(
		.INIT('h1)
	) name4151 (
		_w6714_,
		_w8197_,
		_w8198_
	);
	LUT2 #(
		.INIT('h1)
	) name4152 (
		_w6699_,
		_w6706_,
		_w8199_
	);
	LUT2 #(
		.INIT('h1)
	) name4153 (
		_w6850_,
		_w8199_,
		_w8200_
	);
	LUT2 #(
		.INIT('h8)
	) name4154 (
		_w6850_,
		_w8199_,
		_w8201_
	);
	LUT2 #(
		.INIT('h1)
	) name4155 (
		_w8200_,
		_w8201_,
		_w8202_
	);
	LUT2 #(
		.INIT('h4)
	) name4156 (
		_w8198_,
		_w8202_,
		_w8203_
	);
	LUT2 #(
		.INIT('h4)
	) name4157 (
		_w6847_,
		_w6875_,
		_w8204_
	);
	LUT2 #(
		.INIT('h1)
	) name4158 (
		_w6857_,
		_w6870_,
		_w8205_
	);
	LUT2 #(
		.INIT('h1)
	) name4159 (
		_w8204_,
		_w8205_,
		_w8206_
	);
	LUT2 #(
		.INIT('h8)
	) name4160 (
		_w8204_,
		_w8205_,
		_w8207_
	);
	LUT2 #(
		.INIT('h1)
	) name4161 (
		_w8206_,
		_w8207_,
		_w8208_
	);
	LUT2 #(
		.INIT('h8)
	) name4162 (
		_w8198_,
		_w8208_,
		_w8209_
	);
	LUT2 #(
		.INIT('h1)
	) name4163 (
		_w8203_,
		_w8209_,
		_w8210_
	);
	LUT2 #(
		.INIT('h1)
	) name4164 (
		_w8196_,
		_w8210_,
		_w8211_
	);
	LUT2 #(
		.INIT('h1)
	) name4165 (
		_w6176_,
		_w8211_,
		_w8212_
	);
	LUT2 #(
		.INIT('h2)
	) name4166 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		_w6295_,
		_w8213_
	);
	LUT2 #(
		.INIT('h1)
	) name4167 (
		_w6310_,
		_w6503_,
		_w8214_
	);
	LUT2 #(
		.INIT('h8)
	) name4168 (
		_w6310_,
		_w6503_,
		_w8215_
	);
	LUT2 #(
		.INIT('h1)
	) name4169 (
		_w8214_,
		_w8215_,
		_w8216_
	);
	LUT2 #(
		.INIT('h8)
	) name4170 (
		_w7631_,
		_w8216_,
		_w8217_
	);
	LUT2 #(
		.INIT('h1)
	) name4171 (
		_w6326_,
		_w6327_,
		_w8218_
	);
	LUT2 #(
		.INIT('h4)
	) name4172 (
		_w6370_,
		_w8218_,
		_w8219_
	);
	LUT2 #(
		.INIT('h2)
	) name4173 (
		_w6370_,
		_w8218_,
		_w8220_
	);
	LUT2 #(
		.INIT('h1)
	) name4174 (
		_w8219_,
		_w8220_,
		_w8221_
	);
	LUT2 #(
		.INIT('h4)
	) name4175 (
		_w7631_,
		_w8221_,
		_w8222_
	);
	LUT2 #(
		.INIT('h1)
	) name4176 (
		_w8213_,
		_w8217_,
		_w8223_
	);
	LUT2 #(
		.INIT('h4)
	) name4177 (
		_w8222_,
		_w8223_,
		_w8224_
	);
	LUT2 #(
		.INIT('h2)
	) name4178 (
		_w6176_,
		_w8224_,
		_w8225_
	);
	LUT2 #(
		.INIT('h2)
	) name4179 (
		_w6135_,
		_w8212_,
		_w8226_
	);
	LUT2 #(
		.INIT('h4)
	) name4180 (
		_w8225_,
		_w8226_,
		_w8227_
	);
	LUT2 #(
		.INIT('h1)
	) name4181 (
		_w7005_,
		_w8195_,
		_w8228_
	);
	LUT2 #(
		.INIT('h4)
	) name4182 (
		_w8227_,
		_w8228_,
		_w8229_
	);
	LUT2 #(
		.INIT('h1)
	) name4183 (
		_w8157_,
		_w8229_,
		_w8230_
	);
	LUT2 #(
		.INIT('h2)
	) name4184 (
		\core_dag_ilm1reg_I_reg[11]/NET0131 ,
		_w6442_,
		_w8231_
	);
	LUT2 #(
		.INIT('h1)
	) name4185 (
		_w6453_,
		_w6456_,
		_w8232_
	);
	LUT2 #(
		.INIT('h4)
	) name4186 (
		_w6457_,
		_w7632_,
		_w8233_
	);
	LUT2 #(
		.INIT('h1)
	) name4187 (
		_w6434_,
		_w8233_,
		_w8234_
	);
	LUT2 #(
		.INIT('h1)
	) name4188 (
		_w8232_,
		_w8234_,
		_w8235_
	);
	LUT2 #(
		.INIT('h8)
	) name4189 (
		_w8232_,
		_w8234_,
		_w8236_
	);
	LUT2 #(
		.INIT('h1)
	) name4190 (
		_w8235_,
		_w8236_,
		_w8237_
	);
	LUT2 #(
		.INIT('h4)
	) name4191 (
		_w7631_,
		_w8237_,
		_w8238_
	);
	LUT2 #(
		.INIT('h1)
	) name4192 (
		_w6425_,
		_w7638_,
		_w8239_
	);
	LUT2 #(
		.INIT('h1)
	) name4193 (
		_w6426_,
		_w8239_,
		_w8240_
	);
	LUT2 #(
		.INIT('h2)
	) name4194 (
		_w6446_,
		_w8240_,
		_w8241_
	);
	LUT2 #(
		.INIT('h4)
	) name4195 (
		_w6446_,
		_w8240_,
		_w8242_
	);
	LUT2 #(
		.INIT('h1)
	) name4196 (
		_w8241_,
		_w8242_,
		_w8243_
	);
	LUT2 #(
		.INIT('h8)
	) name4197 (
		_w7631_,
		_w8243_,
		_w8244_
	);
	LUT2 #(
		.INIT('h1)
	) name4198 (
		_w8231_,
		_w8238_,
		_w8245_
	);
	LUT2 #(
		.INIT('h4)
	) name4199 (
		_w8244_,
		_w8245_,
		_w8246_
	);
	LUT2 #(
		.INIT('h4)
	) name4200 (
		_w6135_,
		_w8246_,
		_w8247_
	);
	LUT2 #(
		.INIT('h8)
	) name4201 (
		\DM_rdm[11]_pad ,
		_w7016_,
		_w8248_
	);
	LUT2 #(
		.INIT('h8)
	) name4202 (
		\DM_rd1[11]_pad ,
		_w7022_,
		_w8249_
	);
	LUT2 #(
		.INIT('h8)
	) name4203 (
		\DM_rd4[11]_pad ,
		_w7028_,
		_w8250_
	);
	LUT2 #(
		.INIT('h8)
	) name4204 (
		\DM_rd6[11]_pad ,
		_w7031_,
		_w8251_
	);
	LUT2 #(
		.INIT('h8)
	) name4205 (
		\DM_rd7[11]_pad ,
		_w7034_,
		_w8252_
	);
	LUT2 #(
		.INIT('h8)
	) name4206 (
		\DM_rd3[11]_pad ,
		_w7038_,
		_w8253_
	);
	LUT2 #(
		.INIT('h2)
	) name4207 (
		\DM_rd0[11]_pad ,
		_w7053_,
		_w8254_
	);
	LUT2 #(
		.INIT('h8)
	) name4208 (
		\DM_rd5[11]_pad ,
		_w7043_,
		_w8255_
	);
	LUT2 #(
		.INIT('h8)
	) name4209 (
		\DM_rd2[11]_pad ,
		_w7041_,
		_w8256_
	);
	LUT2 #(
		.INIT('h1)
	) name4210 (
		_w8249_,
		_w8253_,
		_w8257_
	);
	LUT2 #(
		.INIT('h4)
	) name4211 (
		_w8256_,
		_w8257_,
		_w8258_
	);
	LUT2 #(
		.INIT('h1)
	) name4212 (
		_w7057_,
		_w8248_,
		_w8259_
	);
	LUT2 #(
		.INIT('h1)
	) name4213 (
		_w8251_,
		_w8252_,
		_w8260_
	);
	LUT2 #(
		.INIT('h8)
	) name4214 (
		_w8259_,
		_w8260_,
		_w8261_
	);
	LUT2 #(
		.INIT('h4)
	) name4215 (
		_w8250_,
		_w8258_,
		_w8262_
	);
	LUT2 #(
		.INIT('h4)
	) name4216 (
		_w8255_,
		_w8262_,
		_w8263_
	);
	LUT2 #(
		.INIT('h8)
	) name4217 (
		_w8261_,
		_w8263_,
		_w8264_
	);
	LUT2 #(
		.INIT('h4)
	) name4218 (
		_w8254_,
		_w8264_,
		_w8265_
	);
	LUT2 #(
		.INIT('h8)
	) name4219 (
		\regout_STD_C_reg[11]/P0001 ,
		_w6988_,
		_w8266_
	);
	LUT2 #(
		.INIT('h8)
	) name4220 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131 ,
		_w8267_
	);
	LUT2 #(
		.INIT('h8)
	) name4221 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 ,
		_w8268_
	);
	LUT2 #(
		.INIT('h8)
	) name4222 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w8269_
	);
	LUT2 #(
		.INIT('h8)
	) name4223 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131 ,
		_w8270_
	);
	LUT2 #(
		.INIT('h8)
	) name4224 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131 ,
		_w8271_
	);
	LUT2 #(
		.INIT('h8)
	) name4225 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		_w8272_
	);
	LUT2 #(
		.INIT('h8)
	) name4226 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131 ,
		_w8273_
	);
	LUT2 #(
		.INIT('h8)
	) name4227 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131 ,
		_w8274_
	);
	LUT2 #(
		.INIT('h8)
	) name4228 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131 ,
		_w8275_
	);
	LUT2 #(
		.INIT('h8)
	) name4229 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 ,
		_w8276_
	);
	LUT2 #(
		.INIT('h8)
	) name4230 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131 ,
		_w8277_
	);
	LUT2 #(
		.INIT('h8)
	) name4231 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131 ,
		_w8278_
	);
	LUT2 #(
		.INIT('h1)
	) name4232 (
		_w8267_,
		_w8268_,
		_w8279_
	);
	LUT2 #(
		.INIT('h1)
	) name4233 (
		_w8269_,
		_w8270_,
		_w8280_
	);
	LUT2 #(
		.INIT('h1)
	) name4234 (
		_w8271_,
		_w8272_,
		_w8281_
	);
	LUT2 #(
		.INIT('h1)
	) name4235 (
		_w8273_,
		_w8274_,
		_w8282_
	);
	LUT2 #(
		.INIT('h1)
	) name4236 (
		_w8275_,
		_w8276_,
		_w8283_
	);
	LUT2 #(
		.INIT('h1)
	) name4237 (
		_w8277_,
		_w8278_,
		_w8284_
	);
	LUT2 #(
		.INIT('h8)
	) name4238 (
		_w8283_,
		_w8284_,
		_w8285_
	);
	LUT2 #(
		.INIT('h8)
	) name4239 (
		_w8281_,
		_w8282_,
		_w8286_
	);
	LUT2 #(
		.INIT('h8)
	) name4240 (
		_w8279_,
		_w8280_,
		_w8287_
	);
	LUT2 #(
		.INIT('h8)
	) name4241 (
		_w8286_,
		_w8287_,
		_w8288_
	);
	LUT2 #(
		.INIT('h8)
	) name4242 (
		_w8285_,
		_w8288_,
		_w8289_
	);
	LUT2 #(
		.INIT('h2)
	) name4243 (
		_w7128_,
		_w8289_,
		_w8290_
	);
	LUT2 #(
		.INIT('h8)
	) name4244 (
		\tm_tpr_reg_DO_reg[11]/NET0131 ,
		_w7293_,
		_w8291_
	);
	LUT2 #(
		.INIT('h8)
	) name4245 (
		\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w7247_,
		_w8292_
	);
	LUT2 #(
		.INIT('h8)
	) name4246 (
		\bdma_BCTL_reg[11]/NET0131 ,
		_w7230_,
		_w8293_
	);
	LUT2 #(
		.INIT('h8)
	) name4247 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w7299_,
		_w8294_
	);
	LUT2 #(
		.INIT('h8)
	) name4248 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w7234_,
		_w8295_
	);
	LUT2 #(
		.INIT('h8)
	) name4249 (
		\bdma_BOVL_reg[11]/NET0131 ,
		_w7534_,
		_w8296_
	);
	LUT2 #(
		.INIT('h8)
	) name4250 (
		\idma_DOVL_reg[11]/NET0131 ,
		_w7532_,
		_w8297_
	);
	LUT2 #(
		.INIT('h8)
	) name4251 (
		\bdma_BEAD_reg[11]/NET0131 ,
		_w7303_,
		_w8298_
	);
	LUT2 #(
		.INIT('h8)
	) name4252 (
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w7259_,
		_w8299_
	);
	LUT2 #(
		.INIT('h8)
	) name4253 (
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w7249_,
		_w8300_
	);
	LUT2 #(
		.INIT('h8)
	) name4254 (
		\tm_TCR_TMP_reg[11]/NET0131 ,
		_w7289_,
		_w8301_
	);
	LUT2 #(
		.INIT('h8)
	) name4255 (
		\sport0_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w7295_,
		_w8302_
	);
	LUT2 #(
		.INIT('h8)
	) name4256 (
		\emc_WSCRreg_DO_reg[11]/NET0131 ,
		_w7251_,
		_w8303_
	);
	LUT2 #(
		.INIT('h8)
	) name4257 (
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w7273_,
		_w8304_
	);
	LUT2 #(
		.INIT('h8)
	) name4258 (
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w7281_,
		_w8305_
	);
	LUT2 #(
		.INIT('h8)
	) name4259 (
		\sport1_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w7527_,
		_w8306_
	);
	LUT2 #(
		.INIT('h8)
	) name4260 (
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		_w7287_,
		_w8307_
	);
	LUT2 #(
		.INIT('h8)
	) name4261 (
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		_w7689_,
		_w8308_
	);
	LUT2 #(
		.INIT('h8)
	) name4262 (
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		_w7710_,
		_w8309_
	);
	LUT2 #(
		.INIT('h8)
	) name4263 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w7301_,
		_w8310_
	);
	LUT2 #(
		.INIT('h8)
	) name4264 (
		\clkc_ckr_reg_DO_reg[11]/NET0131 ,
		_w7239_,
		_w8311_
	);
	LUT2 #(
		.INIT('h8)
	) name4265 (
		\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w7256_,
		_w8312_
	);
	LUT2 #(
		.INIT('h1)
	) name4266 (
		_w7522_,
		_w8291_,
		_w8313_
	);
	LUT2 #(
		.INIT('h1)
	) name4267 (
		_w8292_,
		_w8294_,
		_w8314_
	);
	LUT2 #(
		.INIT('h1)
	) name4268 (
		_w8297_,
		_w8299_,
		_w8315_
	);
	LUT2 #(
		.INIT('h1)
	) name4269 (
		_w8300_,
		_w8301_,
		_w8316_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		_w8302_,
		_w8303_,
		_w8317_
	);
	LUT2 #(
		.INIT('h1)
	) name4271 (
		_w8304_,
		_w8305_,
		_w8318_
	);
	LUT2 #(
		.INIT('h1)
	) name4272 (
		_w8306_,
		_w8310_,
		_w8319_
	);
	LUT2 #(
		.INIT('h1)
	) name4273 (
		_w8311_,
		_w8312_,
		_w8320_
	);
	LUT2 #(
		.INIT('h8)
	) name4274 (
		_w8319_,
		_w8320_,
		_w8321_
	);
	LUT2 #(
		.INIT('h8)
	) name4275 (
		_w8317_,
		_w8318_,
		_w8322_
	);
	LUT2 #(
		.INIT('h8)
	) name4276 (
		_w8315_,
		_w8316_,
		_w8323_
	);
	LUT2 #(
		.INIT('h8)
	) name4277 (
		_w8313_,
		_w8314_,
		_w8324_
	);
	LUT2 #(
		.INIT('h1)
	) name4278 (
		_w8308_,
		_w8309_,
		_w8325_
	);
	LUT2 #(
		.INIT('h8)
	) name4279 (
		_w8324_,
		_w8325_,
		_w8326_
	);
	LUT2 #(
		.INIT('h8)
	) name4280 (
		_w8322_,
		_w8323_,
		_w8327_
	);
	LUT2 #(
		.INIT('h8)
	) name4281 (
		_w8321_,
		_w8327_,
		_w8328_
	);
	LUT2 #(
		.INIT('h4)
	) name4282 (
		_w8293_,
		_w8326_,
		_w8329_
	);
	LUT2 #(
		.INIT('h1)
	) name4283 (
		_w8295_,
		_w8298_,
		_w8330_
	);
	LUT2 #(
		.INIT('h8)
	) name4284 (
		_w8329_,
		_w8330_,
		_w8331_
	);
	LUT2 #(
		.INIT('h4)
	) name4285 (
		_w8296_,
		_w8328_,
		_w8332_
	);
	LUT2 #(
		.INIT('h4)
	) name4286 (
		_w8307_,
		_w8332_,
		_w8333_
	);
	LUT2 #(
		.INIT('h8)
	) name4287 (
		_w8331_,
		_w8333_,
		_w8334_
	);
	LUT2 #(
		.INIT('h2)
	) name4288 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w8334_,
		_w8335_
	);
	LUT2 #(
		.INIT('h4)
	) name4289 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001 ,
		_w8336_
	);
	LUT2 #(
		.INIT('h8)
	) name4290 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001 ,
		_w8337_
	);
	LUT2 #(
		.INIT('h1)
	) name4291 (
		_w8336_,
		_w8337_,
		_w8338_
	);
	LUT2 #(
		.INIT('h2)
	) name4292 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w8338_,
		_w8339_
	);
	LUT2 #(
		.INIT('h4)
	) name4293 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001 ,
		_w8340_
	);
	LUT2 #(
		.INIT('h8)
	) name4294 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001 ,
		_w8341_
	);
	LUT2 #(
		.INIT('h1)
	) name4295 (
		_w8340_,
		_w8341_,
		_w8342_
	);
	LUT2 #(
		.INIT('h2)
	) name4296 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w8342_,
		_w8343_
	);
	LUT2 #(
		.INIT('h4)
	) name4297 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001 ,
		_w8344_
	);
	LUT2 #(
		.INIT('h8)
	) name4298 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001 ,
		_w8345_
	);
	LUT2 #(
		.INIT('h1)
	) name4299 (
		_w8344_,
		_w8345_,
		_w8346_
	);
	LUT2 #(
		.INIT('h2)
	) name4300 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w8346_,
		_w8347_
	);
	LUT2 #(
		.INIT('h4)
	) name4301 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001 ,
		_w8348_
	);
	LUT2 #(
		.INIT('h8)
	) name4302 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001 ,
		_w8349_
	);
	LUT2 #(
		.INIT('h1)
	) name4303 (
		_w8348_,
		_w8349_,
		_w8350_
	);
	LUT2 #(
		.INIT('h2)
	) name4304 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w8350_,
		_w8351_
	);
	LUT2 #(
		.INIT('h4)
	) name4305 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001 ,
		_w8352_
	);
	LUT2 #(
		.INIT('h8)
	) name4306 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 ,
		_w8353_
	);
	LUT2 #(
		.INIT('h1)
	) name4307 (
		_w8352_,
		_w8353_,
		_w8354_
	);
	LUT2 #(
		.INIT('h2)
	) name4308 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w8354_,
		_w8355_
	);
	LUT2 #(
		.INIT('h4)
	) name4309 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001 ,
		_w8356_
	);
	LUT2 #(
		.INIT('h8)
	) name4310 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 ,
		_w8357_
	);
	LUT2 #(
		.INIT('h1)
	) name4311 (
		_w8356_,
		_w8357_,
		_w8358_
	);
	LUT2 #(
		.INIT('h2)
	) name4312 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w8358_,
		_w8359_
	);
	LUT2 #(
		.INIT('h1)
	) name4313 (
		_w7207_,
		_w8339_,
		_w8360_
	);
	LUT2 #(
		.INIT('h1)
	) name4314 (
		_w8343_,
		_w8347_,
		_w8361_
	);
	LUT2 #(
		.INIT('h1)
	) name4315 (
		_w8351_,
		_w8355_,
		_w8362_
	);
	LUT2 #(
		.INIT('h4)
	) name4316 (
		_w8359_,
		_w8362_,
		_w8363_
	);
	LUT2 #(
		.INIT('h8)
	) name4317 (
		_w8360_,
		_w8361_,
		_w8364_
	);
	LUT2 #(
		.INIT('h8)
	) name4318 (
		_w8363_,
		_w8364_,
		_w8365_
	);
	LUT2 #(
		.INIT('h2)
	) name4319 (
		_w7179_,
		_w8365_,
		_w8366_
	);
	LUT2 #(
		.INIT('h4)
	) name4320 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001 ,
		_w8367_
	);
	LUT2 #(
		.INIT('h8)
	) name4321 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001 ,
		_w8368_
	);
	LUT2 #(
		.INIT('h1)
	) name4322 (
		_w8367_,
		_w8368_,
		_w8369_
	);
	LUT2 #(
		.INIT('h2)
	) name4323 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w8369_,
		_w8370_
	);
	LUT2 #(
		.INIT('h4)
	) name4324 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001 ,
		_w8371_
	);
	LUT2 #(
		.INIT('h8)
	) name4325 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001 ,
		_w8372_
	);
	LUT2 #(
		.INIT('h1)
	) name4326 (
		_w8371_,
		_w8372_,
		_w8373_
	);
	LUT2 #(
		.INIT('h2)
	) name4327 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w8373_,
		_w8374_
	);
	LUT2 #(
		.INIT('h4)
	) name4328 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001 ,
		_w8375_
	);
	LUT2 #(
		.INIT('h8)
	) name4329 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001 ,
		_w8376_
	);
	LUT2 #(
		.INIT('h1)
	) name4330 (
		_w8375_,
		_w8376_,
		_w8377_
	);
	LUT2 #(
		.INIT('h2)
	) name4331 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w8377_,
		_w8378_
	);
	LUT2 #(
		.INIT('h4)
	) name4332 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001 ,
		_w8379_
	);
	LUT2 #(
		.INIT('h8)
	) name4333 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001 ,
		_w8380_
	);
	LUT2 #(
		.INIT('h1)
	) name4334 (
		_w8379_,
		_w8380_,
		_w8381_
	);
	LUT2 #(
		.INIT('h2)
	) name4335 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w8381_,
		_w8382_
	);
	LUT2 #(
		.INIT('h4)
	) name4336 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001 ,
		_w8383_
	);
	LUT2 #(
		.INIT('h8)
	) name4337 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001 ,
		_w8384_
	);
	LUT2 #(
		.INIT('h1)
	) name4338 (
		_w8383_,
		_w8384_,
		_w8385_
	);
	LUT2 #(
		.INIT('h2)
	) name4339 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w8385_,
		_w8386_
	);
	LUT2 #(
		.INIT('h1)
	) name4340 (
		_w8370_,
		_w8374_,
		_w8387_
	);
	LUT2 #(
		.INIT('h1)
	) name4341 (
		_w8378_,
		_w8382_,
		_w8388_
	);
	LUT2 #(
		.INIT('h4)
	) name4342 (
		_w8386_,
		_w8388_,
		_w8389_
	);
	LUT2 #(
		.INIT('h8)
	) name4343 (
		_w8387_,
		_w8389_,
		_w8390_
	);
	LUT2 #(
		.INIT('h2)
	) name4344 (
		_w7093_,
		_w8390_,
		_w8391_
	);
	LUT2 #(
		.INIT('h2)
	) name4345 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w7216_,
		_w8392_
	);
	LUT2 #(
		.INIT('h8)
	) name4346 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w8393_
	);
	LUT2 #(
		.INIT('h8)
	) name4347 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w8394_
	);
	LUT2 #(
		.INIT('h2)
	) name4348 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4622_,
		_w8395_
	);
	LUT2 #(
		.INIT('h1)
	) name4349 (
		_w8393_,
		_w8394_,
		_w8396_
	);
	LUT2 #(
		.INIT('h4)
	) name4350 (
		_w8392_,
		_w8396_,
		_w8397_
	);
	LUT2 #(
		.INIT('h4)
	) name4351 (
		_w8395_,
		_w8397_,
		_w8398_
	);
	LUT2 #(
		.INIT('h2)
	) name4352 (
		_w7215_,
		_w8398_,
		_w8399_
	);
	LUT2 #(
		.INIT('h4)
	) name4353 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 ,
		_w8400_
	);
	LUT2 #(
		.INIT('h8)
	) name4354 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 ,
		_w8401_
	);
	LUT2 #(
		.INIT('h1)
	) name4355 (
		_w8400_,
		_w8401_,
		_w8402_
	);
	LUT2 #(
		.INIT('h2)
	) name4356 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w8402_,
		_w8403_
	);
	LUT2 #(
		.INIT('h4)
	) name4357 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001 ,
		_w8404_
	);
	LUT2 #(
		.INIT('h8)
	) name4358 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001 ,
		_w8405_
	);
	LUT2 #(
		.INIT('h1)
	) name4359 (
		_w8404_,
		_w8405_,
		_w8406_
	);
	LUT2 #(
		.INIT('h2)
	) name4360 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w8406_,
		_w8407_
	);
	LUT2 #(
		.INIT('h4)
	) name4361 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 ,
		_w8408_
	);
	LUT2 #(
		.INIT('h8)
	) name4362 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 ,
		_w8409_
	);
	LUT2 #(
		.INIT('h1)
	) name4363 (
		_w8408_,
		_w8409_,
		_w8410_
	);
	LUT2 #(
		.INIT('h2)
	) name4364 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w8410_,
		_w8411_
	);
	LUT2 #(
		.INIT('h1)
	) name4365 (
		_w8403_,
		_w8407_,
		_w8412_
	);
	LUT2 #(
		.INIT('h4)
	) name4366 (
		_w8411_,
		_w8412_,
		_w8413_
	);
	LUT2 #(
		.INIT('h8)
	) name4367 (
		_w7174_,
		_w8413_,
		_w8414_
	);
	LUT2 #(
		.INIT('h2)
	) name4368 (
		_w7153_,
		_w8414_,
		_w8415_
	);
	LUT2 #(
		.INIT('h8)
	) name4369 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[11]/P0001 ,
		_w8416_
	);
	LUT2 #(
		.INIT('h8)
	) name4370 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[11]/P0001 ,
		_w8417_
	);
	LUT2 #(
		.INIT('h8)
	) name4371 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[11]/P0001 ,
		_w8418_
	);
	LUT2 #(
		.INIT('h8)
	) name4372 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[11]/P0001 ,
		_w8419_
	);
	LUT2 #(
		.INIT('h1)
	) name4373 (
		_w8416_,
		_w8417_,
		_w8420_
	);
	LUT2 #(
		.INIT('h1)
	) name4374 (
		_w8418_,
		_w8419_,
		_w8421_
	);
	LUT2 #(
		.INIT('h8)
	) name4375 (
		_w8420_,
		_w8421_,
		_w8422_
	);
	LUT2 #(
		.INIT('h2)
	) name4376 (
		_w7119_,
		_w8422_,
		_w8423_
	);
	LUT2 #(
		.INIT('h8)
	) name4377 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131 ,
		_w8424_
	);
	LUT2 #(
		.INIT('h8)
	) name4378 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 ,
		_w8425_
	);
	LUT2 #(
		.INIT('h8)
	) name4379 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 ,
		_w8426_
	);
	LUT2 #(
		.INIT('h8)
	) name4380 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131 ,
		_w8427_
	);
	LUT2 #(
		.INIT('h8)
	) name4381 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 ,
		_w8428_
	);
	LUT2 #(
		.INIT('h8)
	) name4382 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131 ,
		_w8429_
	);
	LUT2 #(
		.INIT('h8)
	) name4383 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131 ,
		_w8430_
	);
	LUT2 #(
		.INIT('h8)
	) name4384 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w8431_
	);
	LUT2 #(
		.INIT('h8)
	) name4385 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131 ,
		_w8432_
	);
	LUT2 #(
		.INIT('h8)
	) name4386 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131 ,
		_w8433_
	);
	LUT2 #(
		.INIT('h8)
	) name4387 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131 ,
		_w8434_
	);
	LUT2 #(
		.INIT('h8)
	) name4388 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131 ,
		_w8435_
	);
	LUT2 #(
		.INIT('h1)
	) name4389 (
		_w8424_,
		_w8425_,
		_w8436_
	);
	LUT2 #(
		.INIT('h1)
	) name4390 (
		_w8426_,
		_w8427_,
		_w8437_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		_w8428_,
		_w8429_,
		_w8438_
	);
	LUT2 #(
		.INIT('h1)
	) name4392 (
		_w8430_,
		_w8431_,
		_w8439_
	);
	LUT2 #(
		.INIT('h1)
	) name4393 (
		_w8432_,
		_w8433_,
		_w8440_
	);
	LUT2 #(
		.INIT('h1)
	) name4394 (
		_w8434_,
		_w8435_,
		_w8441_
	);
	LUT2 #(
		.INIT('h8)
	) name4395 (
		_w8440_,
		_w8441_,
		_w8442_
	);
	LUT2 #(
		.INIT('h8)
	) name4396 (
		_w8438_,
		_w8439_,
		_w8443_
	);
	LUT2 #(
		.INIT('h8)
	) name4397 (
		_w8436_,
		_w8437_,
		_w8444_
	);
	LUT2 #(
		.INIT('h8)
	) name4398 (
		_w8443_,
		_w8444_,
		_w8445_
	);
	LUT2 #(
		.INIT('h8)
	) name4399 (
		_w8442_,
		_w8445_,
		_w8446_
	);
	LUT2 #(
		.INIT('h2)
	) name4400 (
		_w7068_,
		_w8446_,
		_w8447_
	);
	LUT2 #(
		.INIT('h1)
	) name4401 (
		_w8290_,
		_w8423_,
		_w8448_
	);
	LUT2 #(
		.INIT('h4)
	) name4402 (
		_w8447_,
		_w8448_,
		_w8449_
	);
	LUT2 #(
		.INIT('h1)
	) name4403 (
		_w8366_,
		_w8391_,
		_w8450_
	);
	LUT2 #(
		.INIT('h4)
	) name4404 (
		_w8415_,
		_w8450_,
		_w8451_
	);
	LUT2 #(
		.INIT('h8)
	) name4405 (
		_w8449_,
		_w8451_,
		_w8452_
	);
	LUT2 #(
		.INIT('h4)
	) name4406 (
		_w8399_,
		_w8452_,
		_w8453_
	);
	LUT2 #(
		.INIT('h4)
	) name4407 (
		_w8335_,
		_w8453_,
		_w8454_
	);
	LUT2 #(
		.INIT('h4)
	) name4408 (
		_w8266_,
		_w8454_,
		_w8455_
	);
	LUT2 #(
		.INIT('h1)
	) name4409 (
		\emc_DMDoe_reg/NET0131 ,
		_w8455_,
		_w8456_
	);
	LUT2 #(
		.INIT('h8)
	) name4410 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[11]/P0001 ,
		_w8457_
	);
	LUT2 #(
		.INIT('h2)
	) name4411 (
		_w7057_,
		_w8457_,
		_w8458_
	);
	LUT2 #(
		.INIT('h4)
	) name4412 (
		_w8456_,
		_w8458_,
		_w8459_
	);
	LUT2 #(
		.INIT('h1)
	) name4413 (
		_w8265_,
		_w8459_,
		_w8460_
	);
	LUT2 #(
		.INIT('h2)
	) name4414 (
		_w6135_,
		_w8460_,
		_w8461_
	);
	LUT2 #(
		.INIT('h2)
	) name4415 (
		_w6176_,
		_w8461_,
		_w8462_
	);
	LUT2 #(
		.INIT('h4)
	) name4416 (
		_w8247_,
		_w8462_,
		_w8463_
	);
	LUT2 #(
		.INIT('h8)
	) name4417 (
		\DM_rdm[2]_pad ,
		_w7016_,
		_w8464_
	);
	LUT2 #(
		.INIT('h8)
	) name4418 (
		\DM_rd1[2]_pad ,
		_w7022_,
		_w8465_
	);
	LUT2 #(
		.INIT('h8)
	) name4419 (
		\DM_rd5[2]_pad ,
		_w7043_,
		_w8466_
	);
	LUT2 #(
		.INIT('h8)
	) name4420 (
		\DM_rd6[2]_pad ,
		_w7031_,
		_w8467_
	);
	LUT2 #(
		.INIT('h8)
	) name4421 (
		\DM_rd7[2]_pad ,
		_w7034_,
		_w8468_
	);
	LUT2 #(
		.INIT('h8)
	) name4422 (
		\DM_rd3[2]_pad ,
		_w7038_,
		_w8469_
	);
	LUT2 #(
		.INIT('h2)
	) name4423 (
		\DM_rd0[2]_pad ,
		_w7053_,
		_w8470_
	);
	LUT2 #(
		.INIT('h8)
	) name4424 (
		\DM_rd4[2]_pad ,
		_w7028_,
		_w8471_
	);
	LUT2 #(
		.INIT('h8)
	) name4425 (
		\DM_rd2[2]_pad ,
		_w7041_,
		_w8472_
	);
	LUT2 #(
		.INIT('h1)
	) name4426 (
		_w8465_,
		_w8469_,
		_w8473_
	);
	LUT2 #(
		.INIT('h4)
	) name4427 (
		_w8472_,
		_w8473_,
		_w8474_
	);
	LUT2 #(
		.INIT('h1)
	) name4428 (
		_w7057_,
		_w8464_,
		_w8475_
	);
	LUT2 #(
		.INIT('h1)
	) name4429 (
		_w8467_,
		_w8468_,
		_w8476_
	);
	LUT2 #(
		.INIT('h8)
	) name4430 (
		_w8475_,
		_w8476_,
		_w8477_
	);
	LUT2 #(
		.INIT('h4)
	) name4431 (
		_w8466_,
		_w8474_,
		_w8478_
	);
	LUT2 #(
		.INIT('h4)
	) name4432 (
		_w8471_,
		_w8478_,
		_w8479_
	);
	LUT2 #(
		.INIT('h8)
	) name4433 (
		_w8477_,
		_w8479_,
		_w8480_
	);
	LUT2 #(
		.INIT('h4)
	) name4434 (
		_w8470_,
		_w8480_,
		_w8481_
	);
	LUT2 #(
		.INIT('h8)
	) name4435 (
		\regout_STD_C_reg[2]/P0001 ,
		_w6988_,
		_w8482_
	);
	LUT2 #(
		.INIT('h4)
	) name4436 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001 ,
		_w8483_
	);
	LUT2 #(
		.INIT('h8)
	) name4437 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001 ,
		_w8484_
	);
	LUT2 #(
		.INIT('h1)
	) name4438 (
		_w8483_,
		_w8484_,
		_w8485_
	);
	LUT2 #(
		.INIT('h2)
	) name4439 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w8485_,
		_w8486_
	);
	LUT2 #(
		.INIT('h4)
	) name4440 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[2]/P0001 ,
		_w8487_
	);
	LUT2 #(
		.INIT('h8)
	) name4441 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBs_reg[2]/P0001 ,
		_w8488_
	);
	LUT2 #(
		.INIT('h1)
	) name4442 (
		_w8487_,
		_w8488_,
		_w8489_
	);
	LUT2 #(
		.INIT('h2)
	) name4443 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		_w8489_,
		_w8490_
	);
	LUT2 #(
		.INIT('h4)
	) name4444 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 ,
		_w8491_
	);
	LUT2 #(
		.INIT('h8)
	) name4445 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 ,
		_w8492_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		_w8491_,
		_w8492_,
		_w8493_
	);
	LUT2 #(
		.INIT('h2)
	) name4447 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w8493_,
		_w8494_
	);
	LUT2 #(
		.INIT('h4)
	) name4448 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 ,
		_w8495_
	);
	LUT2 #(
		.INIT('h8)
	) name4449 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 ,
		_w8496_
	);
	LUT2 #(
		.INIT('h1)
	) name4450 (
		_w8495_,
		_w8496_,
		_w8497_
	);
	LUT2 #(
		.INIT('h2)
	) name4451 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w8497_,
		_w8498_
	);
	LUT2 #(
		.INIT('h4)
	) name4452 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001 ,
		_w8499_
	);
	LUT2 #(
		.INIT('h8)
	) name4453 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001 ,
		_w8500_
	);
	LUT2 #(
		.INIT('h1)
	) name4454 (
		_w8499_,
		_w8500_,
		_w8501_
	);
	LUT2 #(
		.INIT('h2)
	) name4455 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w8501_,
		_w8502_
	);
	LUT2 #(
		.INIT('h1)
	) name4456 (
		_w8486_,
		_w8490_,
		_w8503_
	);
	LUT2 #(
		.INIT('h1)
	) name4457 (
		_w8494_,
		_w8498_,
		_w8504_
	);
	LUT2 #(
		.INIT('h4)
	) name4458 (
		_w8502_,
		_w8504_,
		_w8505_
	);
	LUT2 #(
		.INIT('h8)
	) name4459 (
		_w8503_,
		_w8505_,
		_w8506_
	);
	LUT2 #(
		.INIT('h2)
	) name4460 (
		_w7153_,
		_w8506_,
		_w8507_
	);
	LUT2 #(
		.INIT('h8)
	) name4461 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w8508_
	);
	LUT2 #(
		.INIT('h8)
	) name4462 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 ,
		_w8509_
	);
	LUT2 #(
		.INIT('h8)
	) name4463 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131 ,
		_w8510_
	);
	LUT2 #(
		.INIT('h8)
	) name4464 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131 ,
		_w8511_
	);
	LUT2 #(
		.INIT('h8)
	) name4465 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131 ,
		_w8512_
	);
	LUT2 #(
		.INIT('h8)
	) name4466 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131 ,
		_w8513_
	);
	LUT2 #(
		.INIT('h8)
	) name4467 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 ,
		_w8514_
	);
	LUT2 #(
		.INIT('h8)
	) name4468 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w8515_
	);
	LUT2 #(
		.INIT('h8)
	) name4469 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131 ,
		_w8516_
	);
	LUT2 #(
		.INIT('h8)
	) name4470 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131 ,
		_w8517_
	);
	LUT2 #(
		.INIT('h8)
	) name4471 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131 ,
		_w8518_
	);
	LUT2 #(
		.INIT('h8)
	) name4472 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131 ,
		_w8519_
	);
	LUT2 #(
		.INIT('h1)
	) name4473 (
		_w8508_,
		_w8509_,
		_w8520_
	);
	LUT2 #(
		.INIT('h1)
	) name4474 (
		_w8510_,
		_w8511_,
		_w8521_
	);
	LUT2 #(
		.INIT('h1)
	) name4475 (
		_w8512_,
		_w8513_,
		_w8522_
	);
	LUT2 #(
		.INIT('h1)
	) name4476 (
		_w8514_,
		_w8515_,
		_w8523_
	);
	LUT2 #(
		.INIT('h1)
	) name4477 (
		_w8516_,
		_w8517_,
		_w8524_
	);
	LUT2 #(
		.INIT('h1)
	) name4478 (
		_w8518_,
		_w8519_,
		_w8525_
	);
	LUT2 #(
		.INIT('h8)
	) name4479 (
		_w8524_,
		_w8525_,
		_w8526_
	);
	LUT2 #(
		.INIT('h8)
	) name4480 (
		_w8522_,
		_w8523_,
		_w8527_
	);
	LUT2 #(
		.INIT('h8)
	) name4481 (
		_w8520_,
		_w8521_,
		_w8528_
	);
	LUT2 #(
		.INIT('h8)
	) name4482 (
		_w8527_,
		_w8528_,
		_w8529_
	);
	LUT2 #(
		.INIT('h8)
	) name4483 (
		_w8526_,
		_w8529_,
		_w8530_
	);
	LUT2 #(
		.INIT('h2)
	) name4484 (
		_w7068_,
		_w8530_,
		_w8531_
	);
	LUT2 #(
		.INIT('h4)
	) name4485 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 ,
		_w8532_
	);
	LUT2 #(
		.INIT('h8)
	) name4486 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 ,
		_w8533_
	);
	LUT2 #(
		.INIT('h1)
	) name4487 (
		_w8532_,
		_w8533_,
		_w8534_
	);
	LUT2 #(
		.INIT('h2)
	) name4488 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w8534_,
		_w8535_
	);
	LUT2 #(
		.INIT('h4)
	) name4489 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001 ,
		_w8536_
	);
	LUT2 #(
		.INIT('h8)
	) name4490 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001 ,
		_w8537_
	);
	LUT2 #(
		.INIT('h1)
	) name4491 (
		_w8536_,
		_w8537_,
		_w8538_
	);
	LUT2 #(
		.INIT('h2)
	) name4492 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w8538_,
		_w8539_
	);
	LUT2 #(
		.INIT('h4)
	) name4493 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001 ,
		_w8540_
	);
	LUT2 #(
		.INIT('h8)
	) name4494 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001 ,
		_w8541_
	);
	LUT2 #(
		.INIT('h1)
	) name4495 (
		_w8540_,
		_w8541_,
		_w8542_
	);
	LUT2 #(
		.INIT('h2)
	) name4496 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w8542_,
		_w8543_
	);
	LUT2 #(
		.INIT('h4)
	) name4497 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001 ,
		_w8544_
	);
	LUT2 #(
		.INIT('h8)
	) name4498 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001 ,
		_w8545_
	);
	LUT2 #(
		.INIT('h1)
	) name4499 (
		_w8544_,
		_w8545_,
		_w8546_
	);
	LUT2 #(
		.INIT('h2)
	) name4500 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w8546_,
		_w8547_
	);
	LUT2 #(
		.INIT('h4)
	) name4501 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001 ,
		_w8548_
	);
	LUT2 #(
		.INIT('h8)
	) name4502 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001 ,
		_w8549_
	);
	LUT2 #(
		.INIT('h1)
	) name4503 (
		_w8548_,
		_w8549_,
		_w8550_
	);
	LUT2 #(
		.INIT('h2)
	) name4504 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w8550_,
		_w8551_
	);
	LUT2 #(
		.INIT('h4)
	) name4505 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001 ,
		_w8552_
	);
	LUT2 #(
		.INIT('h8)
	) name4506 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 ,
		_w8553_
	);
	LUT2 #(
		.INIT('h1)
	) name4507 (
		_w8552_,
		_w8553_,
		_w8554_
	);
	LUT2 #(
		.INIT('h2)
	) name4508 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w8554_,
		_w8555_
	);
	LUT2 #(
		.INIT('h4)
	) name4509 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001 ,
		_w8556_
	);
	LUT2 #(
		.INIT('h8)
	) name4510 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 ,
		_w8557_
	);
	LUT2 #(
		.INIT('h1)
	) name4511 (
		_w8556_,
		_w8557_,
		_w8558_
	);
	LUT2 #(
		.INIT('h2)
	) name4512 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w8558_,
		_w8559_
	);
	LUT2 #(
		.INIT('h1)
	) name4513 (
		_w8535_,
		_w8539_,
		_w8560_
	);
	LUT2 #(
		.INIT('h1)
	) name4514 (
		_w8543_,
		_w8547_,
		_w8561_
	);
	LUT2 #(
		.INIT('h1)
	) name4515 (
		_w8551_,
		_w8555_,
		_w8562_
	);
	LUT2 #(
		.INIT('h4)
	) name4516 (
		_w8559_,
		_w8562_,
		_w8563_
	);
	LUT2 #(
		.INIT('h8)
	) name4517 (
		_w8560_,
		_w8561_,
		_w8564_
	);
	LUT2 #(
		.INIT('h8)
	) name4518 (
		_w8563_,
		_w8564_,
		_w8565_
	);
	LUT2 #(
		.INIT('h2)
	) name4519 (
		_w7179_,
		_w8565_,
		_w8566_
	);
	LUT2 #(
		.INIT('h8)
	) name4520 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[2]/P0001 ,
		_w8567_
	);
	LUT2 #(
		.INIT('h8)
	) name4521 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w8568_
	);
	LUT2 #(
		.INIT('h8)
	) name4522 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[2]/P0001 ,
		_w8569_
	);
	LUT2 #(
		.INIT('h8)
	) name4523 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w8570_
	);
	LUT2 #(
		.INIT('h1)
	) name4524 (
		_w8567_,
		_w8568_,
		_w8571_
	);
	LUT2 #(
		.INIT('h1)
	) name4525 (
		_w8569_,
		_w8570_,
		_w8572_
	);
	LUT2 #(
		.INIT('h8)
	) name4526 (
		_w8571_,
		_w8572_,
		_w8573_
	);
	LUT2 #(
		.INIT('h2)
	) name4527 (
		_w7119_,
		_w8573_,
		_w8574_
	);
	LUT2 #(
		.INIT('h4)
	) name4528 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001 ,
		_w8575_
	);
	LUT2 #(
		.INIT('h8)
	) name4529 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001 ,
		_w8576_
	);
	LUT2 #(
		.INIT('h1)
	) name4530 (
		_w8575_,
		_w8576_,
		_w8577_
	);
	LUT2 #(
		.INIT('h2)
	) name4531 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w8577_,
		_w8578_
	);
	LUT2 #(
		.INIT('h4)
	) name4532 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001 ,
		_w8579_
	);
	LUT2 #(
		.INIT('h8)
	) name4533 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001 ,
		_w8580_
	);
	LUT2 #(
		.INIT('h1)
	) name4534 (
		_w8579_,
		_w8580_,
		_w8581_
	);
	LUT2 #(
		.INIT('h2)
	) name4535 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w8581_,
		_w8582_
	);
	LUT2 #(
		.INIT('h4)
	) name4536 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001 ,
		_w8583_
	);
	LUT2 #(
		.INIT('h8)
	) name4537 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001 ,
		_w8584_
	);
	LUT2 #(
		.INIT('h1)
	) name4538 (
		_w8583_,
		_w8584_,
		_w8585_
	);
	LUT2 #(
		.INIT('h2)
	) name4539 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w8585_,
		_w8586_
	);
	LUT2 #(
		.INIT('h4)
	) name4540 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001 ,
		_w8587_
	);
	LUT2 #(
		.INIT('h8)
	) name4541 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001 ,
		_w8588_
	);
	LUT2 #(
		.INIT('h1)
	) name4542 (
		_w8587_,
		_w8588_,
		_w8589_
	);
	LUT2 #(
		.INIT('h2)
	) name4543 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w8589_,
		_w8590_
	);
	LUT2 #(
		.INIT('h4)
	) name4544 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001 ,
		_w8591_
	);
	LUT2 #(
		.INIT('h8)
	) name4545 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001 ,
		_w8592_
	);
	LUT2 #(
		.INIT('h1)
	) name4546 (
		_w8591_,
		_w8592_,
		_w8593_
	);
	LUT2 #(
		.INIT('h2)
	) name4547 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w8593_,
		_w8594_
	);
	LUT2 #(
		.INIT('h8)
	) name4548 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w8595_
	);
	LUT2 #(
		.INIT('h1)
	) name4549 (
		_w8578_,
		_w8595_,
		_w8596_
	);
	LUT2 #(
		.INIT('h1)
	) name4550 (
		_w8582_,
		_w8586_,
		_w8597_
	);
	LUT2 #(
		.INIT('h1)
	) name4551 (
		_w8590_,
		_w8594_,
		_w8598_
	);
	LUT2 #(
		.INIT('h8)
	) name4552 (
		_w8597_,
		_w8598_,
		_w8599_
	);
	LUT2 #(
		.INIT('h8)
	) name4553 (
		_w8596_,
		_w8599_,
		_w8600_
	);
	LUT2 #(
		.INIT('h2)
	) name4554 (
		_w7093_,
		_w8600_,
		_w8601_
	);
	LUT2 #(
		.INIT('h8)
	) name4555 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131 ,
		_w8602_
	);
	LUT2 #(
		.INIT('h8)
	) name4556 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131 ,
		_w8603_
	);
	LUT2 #(
		.INIT('h8)
	) name4557 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131 ,
		_w8604_
	);
	LUT2 #(
		.INIT('h8)
	) name4558 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131 ,
		_w8605_
	);
	LUT2 #(
		.INIT('h8)
	) name4559 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131 ,
		_w8606_
	);
	LUT2 #(
		.INIT('h8)
	) name4560 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131 ,
		_w8607_
	);
	LUT2 #(
		.INIT('h8)
	) name4561 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131 ,
		_w8608_
	);
	LUT2 #(
		.INIT('h8)
	) name4562 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131 ,
		_w8609_
	);
	LUT2 #(
		.INIT('h8)
	) name4563 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w8610_
	);
	LUT2 #(
		.INIT('h8)
	) name4564 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w8611_
	);
	LUT2 #(
		.INIT('h8)
	) name4565 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		_w8612_
	);
	LUT2 #(
		.INIT('h8)
	) name4566 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w8613_
	);
	LUT2 #(
		.INIT('h1)
	) name4567 (
		_w8602_,
		_w8603_,
		_w8614_
	);
	LUT2 #(
		.INIT('h1)
	) name4568 (
		_w8604_,
		_w8605_,
		_w8615_
	);
	LUT2 #(
		.INIT('h1)
	) name4569 (
		_w8606_,
		_w8607_,
		_w8616_
	);
	LUT2 #(
		.INIT('h1)
	) name4570 (
		_w8608_,
		_w8609_,
		_w8617_
	);
	LUT2 #(
		.INIT('h1)
	) name4571 (
		_w8610_,
		_w8611_,
		_w8618_
	);
	LUT2 #(
		.INIT('h1)
	) name4572 (
		_w8612_,
		_w8613_,
		_w8619_
	);
	LUT2 #(
		.INIT('h8)
	) name4573 (
		_w8618_,
		_w8619_,
		_w8620_
	);
	LUT2 #(
		.INIT('h8)
	) name4574 (
		_w8616_,
		_w8617_,
		_w8621_
	);
	LUT2 #(
		.INIT('h8)
	) name4575 (
		_w8614_,
		_w8615_,
		_w8622_
	);
	LUT2 #(
		.INIT('h8)
	) name4576 (
		_w8621_,
		_w8622_,
		_w8623_
	);
	LUT2 #(
		.INIT('h8)
	) name4577 (
		_w8620_,
		_w8623_,
		_w8624_
	);
	LUT2 #(
		.INIT('h2)
	) name4578 (
		_w7128_,
		_w8624_,
		_w8625_
	);
	LUT2 #(
		.INIT('h8)
	) name4579 (
		\idma_DOVL_reg[2]/NET0131 ,
		_w7532_,
		_w8626_
	);
	LUT2 #(
		.INIT('h8)
	) name4580 (
		\sport0_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w7295_,
		_w8627_
	);
	LUT2 #(
		.INIT('h8)
	) name4581 (
		\tm_tpr_reg_DO_reg[2]/NET0131 ,
		_w7293_,
		_w8628_
	);
	LUT2 #(
		.INIT('h8)
	) name4582 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		_w7287_,
		_w8629_
	);
	LUT2 #(
		.INIT('h8)
	) name4583 (
		\emc_WSCRreg_DO_reg[2]/NET0131 ,
		_w7251_,
		_w8630_
	);
	LUT2 #(
		.INIT('h8)
	) name4584 (
		\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w7256_,
		_w8631_
	);
	LUT2 #(
		.INIT('h8)
	) name4585 (
		\sport1_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w7263_,
		_w8632_
	);
	LUT2 #(
		.INIT('h8)
	) name4586 (
		\tm_tsr_reg_DO_reg[2]/NET0131 ,
		_w7540_,
		_w8633_
	);
	LUT2 #(
		.INIT('h8)
	) name4587 (
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w7249_,
		_w8634_
	);
	LUT2 #(
		.INIT('h8)
	) name4588 (
		\emc_WSCRext_reg_DO_reg[2]/NET0131 ,
		_w7514_,
		_w8635_
	);
	LUT2 #(
		.INIT('h8)
	) name4589 (
		\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w7247_,
		_w8636_
	);
	LUT2 #(
		.INIT('h8)
	) name4590 (
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w7281_,
		_w8637_
	);
	LUT2 #(
		.INIT('h8)
	) name4591 (
		\pio_pmask_reg_DO_reg[2]/NET0131 ,
		_w7297_,
		_w8638_
	);
	LUT2 #(
		.INIT('h8)
	) name4592 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w7234_,
		_w8639_
	);
	LUT2 #(
		.INIT('h8)
	) name4593 (
		\sport0_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w7276_,
		_w8640_
	);
	LUT2 #(
		.INIT('h8)
	) name4594 (
		\sport1_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w7527_,
		_w8641_
	);
	LUT2 #(
		.INIT('h8)
	) name4595 (
		\tm_TCR_TMP_reg[2]/NET0131 ,
		_w7289_,
		_w8642_
	);
	LUT2 #(
		.INIT('h8)
	) name4596 (
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w7259_,
		_w8643_
	);
	LUT2 #(
		.INIT('h8)
	) name4597 (
		\bdma_BOVL_reg[2]/NET0131 ,
		_w7534_,
		_w8644_
	);
	LUT2 #(
		.INIT('h8)
	) name4598 (
		\clkc_ckr_reg_DO_reg[2]/NET0131 ,
		_w7239_,
		_w8645_
	);
	LUT2 #(
		.INIT('h8)
	) name4599 (
		\memc_usysr_DO_reg[2]/NET0131 ,
		_w7301_,
		_w8646_
	);
	LUT2 #(
		.INIT('h8)
	) name4600 (
		\bdma_BEAD_reg[2]/NET0131 ,
		_w7303_,
		_w8647_
	);
	LUT2 #(
		.INIT('h8)
	) name4601 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w7230_,
		_w8648_
	);
	LUT2 #(
		.INIT('h8)
	) name4602 (
		\pio_PINT_reg[2]/NET0131 ,
		_w7271_,
		_w8649_
	);
	LUT2 #(
		.INIT('h8)
	) name4603 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w7299_,
		_w8650_
	);
	LUT2 #(
		.INIT('h8)
	) name4604 (
		\PIO_out[2]_pad ,
		_w7291_,
		_w8651_
	);
	LUT2 #(
		.INIT('h8)
	) name4605 (
		\PIO_oe[2]_pad ,
		_w7244_,
		_w8652_
	);
	LUT2 #(
		.INIT('h8)
	) name4606 (
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w7273_,
		_w8653_
	);
	LUT2 #(
		.INIT('h1)
	) name4607 (
		_w7522_,
		_w8626_,
		_w8654_
	);
	LUT2 #(
		.INIT('h1)
	) name4608 (
		_w8627_,
		_w8628_,
		_w8655_
	);
	LUT2 #(
		.INIT('h1)
	) name4609 (
		_w8630_,
		_w8631_,
		_w8656_
	);
	LUT2 #(
		.INIT('h1)
	) name4610 (
		_w8632_,
		_w8633_,
		_w8657_
	);
	LUT2 #(
		.INIT('h1)
	) name4611 (
		_w8634_,
		_w8635_,
		_w8658_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		_w8636_,
		_w8637_,
		_w8659_
	);
	LUT2 #(
		.INIT('h1)
	) name4613 (
		_w8638_,
		_w8640_,
		_w8660_
	);
	LUT2 #(
		.INIT('h1)
	) name4614 (
		_w8641_,
		_w8642_,
		_w8661_
	);
	LUT2 #(
		.INIT('h1)
	) name4615 (
		_w8643_,
		_w8645_,
		_w8662_
	);
	LUT2 #(
		.INIT('h1)
	) name4616 (
		_w8646_,
		_w8649_,
		_w8663_
	);
	LUT2 #(
		.INIT('h1)
	) name4617 (
		_w8650_,
		_w8651_,
		_w8664_
	);
	LUT2 #(
		.INIT('h1)
	) name4618 (
		_w8652_,
		_w8653_,
		_w8665_
	);
	LUT2 #(
		.INIT('h8)
	) name4619 (
		_w8664_,
		_w8665_,
		_w8666_
	);
	LUT2 #(
		.INIT('h8)
	) name4620 (
		_w8662_,
		_w8663_,
		_w8667_
	);
	LUT2 #(
		.INIT('h8)
	) name4621 (
		_w8660_,
		_w8661_,
		_w8668_
	);
	LUT2 #(
		.INIT('h8)
	) name4622 (
		_w8658_,
		_w8659_,
		_w8669_
	);
	LUT2 #(
		.INIT('h8)
	) name4623 (
		_w8656_,
		_w8657_,
		_w8670_
	);
	LUT2 #(
		.INIT('h8)
	) name4624 (
		_w8654_,
		_w8655_,
		_w8671_
	);
	LUT2 #(
		.INIT('h8)
	) name4625 (
		_w8670_,
		_w8671_,
		_w8672_
	);
	LUT2 #(
		.INIT('h8)
	) name4626 (
		_w8668_,
		_w8669_,
		_w8673_
	);
	LUT2 #(
		.INIT('h8)
	) name4627 (
		_w8666_,
		_w8667_,
		_w8674_
	);
	LUT2 #(
		.INIT('h8)
	) name4628 (
		_w8673_,
		_w8674_,
		_w8675_
	);
	LUT2 #(
		.INIT('h4)
	) name4629 (
		_w8639_,
		_w8672_,
		_w8676_
	);
	LUT2 #(
		.INIT('h1)
	) name4630 (
		_w8647_,
		_w8648_,
		_w8677_
	);
	LUT2 #(
		.INIT('h8)
	) name4631 (
		_w8676_,
		_w8677_,
		_w8678_
	);
	LUT2 #(
		.INIT('h4)
	) name4632 (
		_w8629_,
		_w8675_,
		_w8679_
	);
	LUT2 #(
		.INIT('h4)
	) name4633 (
		_w8644_,
		_w8679_,
		_w8680_
	);
	LUT2 #(
		.INIT('h8)
	) name4634 (
		_w8678_,
		_w8680_,
		_w8681_
	);
	LUT2 #(
		.INIT('h2)
	) name4635 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w8681_,
		_w8682_
	);
	LUT2 #(
		.INIT('h8)
	) name4636 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w8683_
	);
	LUT2 #(
		.INIT('h8)
	) name4637 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w8684_
	);
	LUT2 #(
		.INIT('h8)
	) name4638 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w8685_
	);
	LUT2 #(
		.INIT('h2)
	) name4639 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4521_,
		_w8686_
	);
	LUT2 #(
		.INIT('h2)
	) name4640 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w7216_,
		_w8687_
	);
	LUT2 #(
		.INIT('h8)
	) name4641 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		_w8688_
	);
	LUT2 #(
		.INIT('h8)
	) name4642 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w8689_
	);
	LUT2 #(
		.INIT('h8)
	) name4643 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[2]/NET0131 ,
		_w8690_
	);
	LUT2 #(
		.INIT('h8)
	) name4644 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w8691_
	);
	LUT2 #(
		.INIT('h8)
	) name4645 (
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		_w8692_
	);
	LUT2 #(
		.INIT('h1)
	) name4646 (
		_w8683_,
		_w8684_,
		_w8693_
	);
	LUT2 #(
		.INIT('h1)
	) name4647 (
		_w8685_,
		_w8688_,
		_w8694_
	);
	LUT2 #(
		.INIT('h1)
	) name4648 (
		_w8689_,
		_w8690_,
		_w8695_
	);
	LUT2 #(
		.INIT('h1)
	) name4649 (
		_w8691_,
		_w8692_,
		_w8696_
	);
	LUT2 #(
		.INIT('h8)
	) name4650 (
		_w8695_,
		_w8696_,
		_w8697_
	);
	LUT2 #(
		.INIT('h8)
	) name4651 (
		_w8693_,
		_w8694_,
		_w8698_
	);
	LUT2 #(
		.INIT('h4)
	) name4652 (
		_w8687_,
		_w8698_,
		_w8699_
	);
	LUT2 #(
		.INIT('h8)
	) name4653 (
		_w8697_,
		_w8699_,
		_w8700_
	);
	LUT2 #(
		.INIT('h4)
	) name4654 (
		_w8686_,
		_w8700_,
		_w8701_
	);
	LUT2 #(
		.INIT('h2)
	) name4655 (
		_w7215_,
		_w8701_,
		_w8702_
	);
	LUT2 #(
		.INIT('h1)
	) name4656 (
		_w8531_,
		_w8574_,
		_w8703_
	);
	LUT2 #(
		.INIT('h4)
	) name4657 (
		_w8625_,
		_w8703_,
		_w8704_
	);
	LUT2 #(
		.INIT('h1)
	) name4658 (
		_w8507_,
		_w8566_,
		_w8705_
	);
	LUT2 #(
		.INIT('h4)
	) name4659 (
		_w8601_,
		_w8705_,
		_w8706_
	);
	LUT2 #(
		.INIT('h8)
	) name4660 (
		_w8704_,
		_w8706_,
		_w8707_
	);
	LUT2 #(
		.INIT('h4)
	) name4661 (
		_w8702_,
		_w8707_,
		_w8708_
	);
	LUT2 #(
		.INIT('h4)
	) name4662 (
		_w8682_,
		_w8708_,
		_w8709_
	);
	LUT2 #(
		.INIT('h4)
	) name4663 (
		_w8482_,
		_w8709_,
		_w8710_
	);
	LUT2 #(
		.INIT('h1)
	) name4664 (
		\emc_DMDoe_reg/NET0131 ,
		_w8710_,
		_w8711_
	);
	LUT2 #(
		.INIT('h8)
	) name4665 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[2]/P0001 ,
		_w8712_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		_w7057_,
		_w8712_,
		_w8713_
	);
	LUT2 #(
		.INIT('h4)
	) name4667 (
		_w8711_,
		_w8713_,
		_w8714_
	);
	LUT2 #(
		.INIT('h1)
	) name4668 (
		_w8481_,
		_w8714_,
		_w8715_
	);
	LUT2 #(
		.INIT('h8)
	) name4669 (
		_w7863_,
		_w8715_,
		_w8716_
	);
	LUT2 #(
		.INIT('h8)
	) name4670 (
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		_w6976_,
		_w8717_
	);
	LUT2 #(
		.INIT('h8)
	) name4671 (
		\core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 ,
		_w6970_,
		_w8718_
	);
	LUT2 #(
		.INIT('h8)
	) name4672 (
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w6974_,
		_w8719_
	);
	LUT2 #(
		.INIT('h8)
	) name4673 (
		\core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 ,
		_w6972_,
		_w8720_
	);
	LUT2 #(
		.INIT('h1)
	) name4674 (
		_w8717_,
		_w8718_,
		_w8721_
	);
	LUT2 #(
		.INIT('h1)
	) name4675 (
		_w8719_,
		_w8720_,
		_w8722_
	);
	LUT2 #(
		.INIT('h8)
	) name4676 (
		_w8721_,
		_w8722_,
		_w8723_
	);
	LUT2 #(
		.INIT('h2)
	) name4677 (
		_w4055_,
		_w8723_,
		_w8724_
	);
	LUT2 #(
		.INIT('h8)
	) name4678 (
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		_w6958_,
		_w8725_
	);
	LUT2 #(
		.INIT('h8)
	) name4679 (
		\core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 ,
		_w6964_,
		_w8726_
	);
	LUT2 #(
		.INIT('h8)
	) name4680 (
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w6962_,
		_w8727_
	);
	LUT2 #(
		.INIT('h8)
	) name4681 (
		\core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 ,
		_w6960_,
		_w8728_
	);
	LUT2 #(
		.INIT('h1)
	) name4682 (
		_w8725_,
		_w8726_,
		_w8729_
	);
	LUT2 #(
		.INIT('h1)
	) name4683 (
		_w8727_,
		_w8728_,
		_w8730_
	);
	LUT2 #(
		.INIT('h8)
	) name4684 (
		_w8729_,
		_w8730_,
		_w8731_
	);
	LUT2 #(
		.INIT('h4)
	) name4685 (
		_w8724_,
		_w8731_,
		_w8732_
	);
	LUT2 #(
		.INIT('h8)
	) name4686 (
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w8131_,
		_w8733_
	);
	LUT2 #(
		.INIT('h8)
	) name4687 (
		\core_dag_ilm1reg_I2_we_DO_reg[11]/NET0131 ,
		_w6084_,
		_w8734_
	);
	LUT2 #(
		.INIT('h8)
	) name4688 (
		_w6085_,
		_w8734_,
		_w8735_
	);
	LUT2 #(
		.INIT('h8)
	) name4689 (
		\core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 ,
		_w6067_,
		_w8736_
	);
	LUT2 #(
		.INIT('h8)
	) name4690 (
		_w6068_,
		_w8736_,
		_w8737_
	);
	LUT2 #(
		.INIT('h8)
	) name4691 (
		\core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 ,
		_w6075_,
		_w8738_
	);
	LUT2 #(
		.INIT('h8)
	) name4692 (
		_w6077_,
		_w8738_,
		_w8739_
	);
	LUT2 #(
		.INIT('h1)
	) name4693 (
		_w4055_,
		_w8733_,
		_w8740_
	);
	LUT2 #(
		.INIT('h1)
	) name4694 (
		_w8735_,
		_w8737_,
		_w8741_
	);
	LUT2 #(
		.INIT('h4)
	) name4695 (
		_w8739_,
		_w8741_,
		_w8742_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		_w8740_,
		_w8742_,
		_w8743_
	);
	LUT2 #(
		.INIT('h8)
	) name4697 (
		_w6097_,
		_w8738_,
		_w8744_
	);
	LUT2 #(
		.INIT('h8)
	) name4698 (
		_w6095_,
		_w8734_,
		_w8745_
	);
	LUT2 #(
		.INIT('h8)
	) name4699 (
		_w6091_,
		_w8736_,
		_w8746_
	);
	LUT2 #(
		.INIT('h8)
	) name4700 (
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w6148_,
		_w8747_
	);
	LUT2 #(
		.INIT('h1)
	) name4701 (
		_w8744_,
		_w8745_,
		_w8748_
	);
	LUT2 #(
		.INIT('h1)
	) name4702 (
		_w8746_,
		_w8747_,
		_w8749_
	);
	LUT2 #(
		.INIT('h8)
	) name4703 (
		_w8748_,
		_w8749_,
		_w8750_
	);
	LUT2 #(
		.INIT('h8)
	) name4704 (
		_w4055_,
		_w8750_,
		_w8751_
	);
	LUT2 #(
		.INIT('h1)
	) name4705 (
		_w8743_,
		_w8751_,
		_w8752_
	);
	LUT2 #(
		.INIT('h2)
	) name4706 (
		_w8732_,
		_w8752_,
		_w8753_
	);
	LUT2 #(
		.INIT('h2)
	) name4707 (
		_w8153_,
		_w8753_,
		_w8754_
	);
	LUT2 #(
		.INIT('h1)
	) name4708 (
		_w8716_,
		_w8754_,
		_w8755_
	);
	LUT2 #(
		.INIT('h4)
	) name4709 (
		_w8463_,
		_w8755_,
		_w8756_
	);
	LUT2 #(
		.INIT('h2)
	) name4710 (
		_w7005_,
		_w8756_,
		_w8757_
	);
	LUT2 #(
		.INIT('h8)
	) name4711 (
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w6138_,
		_w8758_
	);
	LUT2 #(
		.INIT('h8)
	) name4712 (
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w8131_,
		_w8759_
	);
	LUT2 #(
		.INIT('h8)
	) name4713 (
		\core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 ,
		_w6140_,
		_w8760_
	);
	LUT2 #(
		.INIT('h8)
	) name4714 (
		\core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 ,
		_w6142_,
		_w8761_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w4055_,
		_w8758_,
		_w8762_
	);
	LUT2 #(
		.INIT('h1)
	) name4716 (
		_w8759_,
		_w8760_,
		_w8763_
	);
	LUT2 #(
		.INIT('h4)
	) name4717 (
		_w8761_,
		_w8763_,
		_w8764_
	);
	LUT2 #(
		.INIT('h8)
	) name4718 (
		_w8762_,
		_w8764_,
		_w8765_
	);
	LUT2 #(
		.INIT('h8)
	) name4719 (
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w6084_,
		_w8766_
	);
	LUT2 #(
		.INIT('h8)
	) name4720 (
		_w6095_,
		_w8766_,
		_w8767_
	);
	LUT2 #(
		.INIT('h8)
	) name4721 (
		\core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 ,
		_w6154_,
		_w8768_
	);
	LUT2 #(
		.INIT('h8)
	) name4722 (
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w6148_,
		_w8769_
	);
	LUT2 #(
		.INIT('h8)
	) name4723 (
		\core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 ,
		_w6150_,
		_w8770_
	);
	LUT2 #(
		.INIT('h1)
	) name4724 (
		_w8767_,
		_w8768_,
		_w8771_
	);
	LUT2 #(
		.INIT('h1)
	) name4725 (
		_w8769_,
		_w8770_,
		_w8772_
	);
	LUT2 #(
		.INIT('h8)
	) name4726 (
		_w8771_,
		_w8772_,
		_w8773_
	);
	LUT2 #(
		.INIT('h8)
	) name4727 (
		_w4055_,
		_w8773_,
		_w8774_
	);
	LUT2 #(
		.INIT('h1)
	) name4728 (
		_w8765_,
		_w8774_,
		_w8775_
	);
	LUT2 #(
		.INIT('h4)
	) name4729 (
		_w6135_,
		_w8775_,
		_w8776_
	);
	LUT2 #(
		.INIT('h2)
	) name4730 (
		\core_dag_ilm1reg_I_reg[2]/NET0131 ,
		_w6317_,
		_w8777_
	);
	LUT2 #(
		.INIT('h1)
	) name4731 (
		_w6343_,
		_w6344_,
		_w8778_
	);
	LUT2 #(
		.INIT('h8)
	) name4732 (
		_w6368_,
		_w8778_,
		_w8779_
	);
	LUT2 #(
		.INIT('h1)
	) name4733 (
		_w6368_,
		_w8778_,
		_w8780_
	);
	LUT2 #(
		.INIT('h1)
	) name4734 (
		_w8779_,
		_w8780_,
		_w8781_
	);
	LUT2 #(
		.INIT('h2)
	) name4735 (
		_w6496_,
		_w8781_,
		_w8782_
	);
	LUT2 #(
		.INIT('h2)
	) name4736 (
		_w6339_,
		_w6501_,
		_w8783_
	);
	LUT2 #(
		.INIT('h4)
	) name4737 (
		_w6339_,
		_w6501_,
		_w8784_
	);
	LUT2 #(
		.INIT('h1)
	) name4738 (
		_w8783_,
		_w8784_,
		_w8785_
	);
	LUT2 #(
		.INIT('h4)
	) name4739 (
		_w6496_,
		_w8785_,
		_w8786_
	);
	LUT2 #(
		.INIT('h1)
	) name4740 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w8782_,
		_w8787_
	);
	LUT2 #(
		.INIT('h4)
	) name4741 (
		_w8786_,
		_w8787_,
		_w8788_
	);
	LUT2 #(
		.INIT('h1)
	) name4742 (
		_w7612_,
		_w8781_,
		_w8789_
	);
	LUT2 #(
		.INIT('h8)
	) name4743 (
		_w7612_,
		_w8785_,
		_w8790_
	);
	LUT2 #(
		.INIT('h2)
	) name4744 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w8789_,
		_w8791_
	);
	LUT2 #(
		.INIT('h4)
	) name4745 (
		_w8790_,
		_w8791_,
		_w8792_
	);
	LUT2 #(
		.INIT('h1)
	) name4746 (
		_w8777_,
		_w8792_,
		_w8793_
	);
	LUT2 #(
		.INIT('h4)
	) name4747 (
		_w8788_,
		_w8793_,
		_w8794_
	);
	LUT2 #(
		.INIT('h2)
	) name4748 (
		_w6135_,
		_w8794_,
		_w8795_
	);
	LUT2 #(
		.INIT('h2)
	) name4749 (
		_w6176_,
		_w8776_,
		_w8796_
	);
	LUT2 #(
		.INIT('h4)
	) name4750 (
		_w8795_,
		_w8796_,
		_w8797_
	);
	LUT2 #(
		.INIT('h2)
	) name4751 (
		\core_dag_ilm2reg_I_reg[11]/NET0131 ,
		_w6624_,
		_w8798_
	);
	LUT2 #(
		.INIT('h4)
	) name4752 (
		_w6702_,
		_w8199_,
		_w8799_
	);
	LUT2 #(
		.INIT('h1)
	) name4753 (
		_w6622_,
		_w8799_,
		_w8800_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w6860_,
		_w8800_,
		_w8801_
	);
	LUT2 #(
		.INIT('h8)
	) name4755 (
		_w6860_,
		_w8800_,
		_w8802_
	);
	LUT2 #(
		.INIT('h1)
	) name4756 (
		_w8801_,
		_w8802_,
		_w8803_
	);
	LUT2 #(
		.INIT('h4)
	) name4757 (
		_w8198_,
		_w8803_,
		_w8804_
	);
	LUT2 #(
		.INIT('h1)
	) name4758 (
		_w6867_,
		_w6877_,
		_w8805_
	);
	LUT2 #(
		.INIT('h1)
	) name4759 (
		_w6857_,
		_w8204_,
		_w8806_
	);
	LUT2 #(
		.INIT('h1)
	) name4760 (
		_w6870_,
		_w8806_,
		_w8807_
	);
	LUT2 #(
		.INIT('h2)
	) name4761 (
		_w8805_,
		_w8807_,
		_w8808_
	);
	LUT2 #(
		.INIT('h4)
	) name4762 (
		_w8805_,
		_w8807_,
		_w8809_
	);
	LUT2 #(
		.INIT('h1)
	) name4763 (
		_w8808_,
		_w8809_,
		_w8810_
	);
	LUT2 #(
		.INIT('h8)
	) name4764 (
		_w8198_,
		_w8810_,
		_w8811_
	);
	LUT2 #(
		.INIT('h1)
	) name4765 (
		_w8798_,
		_w8804_,
		_w8812_
	);
	LUT2 #(
		.INIT('h4)
	) name4766 (
		_w8811_,
		_w8812_,
		_w8813_
	);
	LUT2 #(
		.INIT('h2)
	) name4767 (
		_w6135_,
		_w8813_,
		_w8814_
	);
	LUT2 #(
		.INIT('h1)
	) name4768 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w6924_,
		_w8815_
	);
	LUT2 #(
		.INIT('h8)
	) name4769 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131 ,
		_w6988_,
		_w8816_
	);
	LUT2 #(
		.INIT('h8)
	) name4770 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w6926_,
		_w8817_
	);
	LUT2 #(
		.INIT('h4)
	) name4771 (
		_w6111_,
		_w8752_,
		_w8818_
	);
	LUT2 #(
		.INIT('h8)
	) name4772 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w6956_,
		_w8819_
	);
	LUT2 #(
		.INIT('h1)
	) name4773 (
		_w6121_,
		_w8732_,
		_w8820_
	);
	LUT2 #(
		.INIT('h1)
	) name4774 (
		_w8818_,
		_w8819_,
		_w8821_
	);
	LUT2 #(
		.INIT('h4)
	) name4775 (
		_w8820_,
		_w8821_,
		_w8822_
	);
	LUT2 #(
		.INIT('h2)
	) name4776 (
		_w5949_,
		_w8822_,
		_w8823_
	);
	LUT2 #(
		.INIT('h2)
	) name4777 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w6934_,
		_w8824_
	);
	LUT2 #(
		.INIT('h1)
	) name4778 (
		_w8816_,
		_w8817_,
		_w8825_
	);
	LUT2 #(
		.INIT('h8)
	) name4779 (
		_w6924_,
		_w8825_,
		_w8826_
	);
	LUT2 #(
		.INIT('h4)
	) name4780 (
		_w8824_,
		_w8826_,
		_w8827_
	);
	LUT2 #(
		.INIT('h4)
	) name4781 (
		_w8823_,
		_w8827_,
		_w8828_
	);
	LUT2 #(
		.INIT('h1)
	) name4782 (
		_w6135_,
		_w8815_,
		_w8829_
	);
	LUT2 #(
		.INIT('h4)
	) name4783 (
		_w8828_,
		_w8829_,
		_w8830_
	);
	LUT2 #(
		.INIT('h1)
	) name4784 (
		_w6176_,
		_w8830_,
		_w8831_
	);
	LUT2 #(
		.INIT('h4)
	) name4785 (
		_w8814_,
		_w8831_,
		_w8832_
	);
	LUT2 #(
		.INIT('h1)
	) name4786 (
		_w7005_,
		_w8797_,
		_w8833_
	);
	LUT2 #(
		.INIT('h4)
	) name4787 (
		_w8832_,
		_w8833_,
		_w8834_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		_w8757_,
		_w8834_,
		_w8835_
	);
	LUT2 #(
		.INIT('h1)
	) name4789 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w6924_,
		_w8836_
	);
	LUT2 #(
		.INIT('h8)
	) name4790 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w6926_,
		_w8837_
	);
	LUT2 #(
		.INIT('h8)
	) name4791 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131 ,
		_w6988_,
		_w8838_
	);
	LUT2 #(
		.INIT('h8)
	) name4792 (
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w6976_,
		_w8839_
	);
	LUT2 #(
		.INIT('h8)
	) name4793 (
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		_w6970_,
		_w8840_
	);
	LUT2 #(
		.INIT('h8)
	) name4794 (
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w6974_,
		_w8841_
	);
	LUT2 #(
		.INIT('h8)
	) name4795 (
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w6972_,
		_w8842_
	);
	LUT2 #(
		.INIT('h1)
	) name4796 (
		_w8839_,
		_w8840_,
		_w8843_
	);
	LUT2 #(
		.INIT('h1)
	) name4797 (
		_w8841_,
		_w8842_,
		_w8844_
	);
	LUT2 #(
		.INIT('h8)
	) name4798 (
		_w8843_,
		_w8844_,
		_w8845_
	);
	LUT2 #(
		.INIT('h2)
	) name4799 (
		_w4055_,
		_w8845_,
		_w8846_
	);
	LUT2 #(
		.INIT('h8)
	) name4800 (
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w6960_,
		_w8847_
	);
	LUT2 #(
		.INIT('h8)
	) name4801 (
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w6958_,
		_w8848_
	);
	LUT2 #(
		.INIT('h8)
	) name4802 (
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w6962_,
		_w8849_
	);
	LUT2 #(
		.INIT('h8)
	) name4803 (
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		_w6964_,
		_w8850_
	);
	LUT2 #(
		.INIT('h1)
	) name4804 (
		_w8847_,
		_w8848_,
		_w8851_
	);
	LUT2 #(
		.INIT('h1)
	) name4805 (
		_w8849_,
		_w8850_,
		_w8852_
	);
	LUT2 #(
		.INIT('h8)
	) name4806 (
		_w8851_,
		_w8852_,
		_w8853_
	);
	LUT2 #(
		.INIT('h4)
	) name4807 (
		_w8846_,
		_w8853_,
		_w8854_
	);
	LUT2 #(
		.INIT('h1)
	) name4808 (
		_w6121_,
		_w8854_,
		_w8855_
	);
	LUT2 #(
		.INIT('h8)
	) name4809 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w6956_,
		_w8856_
	);
	LUT2 #(
		.INIT('h8)
	) name4810 (
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		_w6138_,
		_w8857_
	);
	LUT2 #(
		.INIT('h8)
	) name4811 (
		\core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 ,
		_w6140_,
		_w8858_
	);
	LUT2 #(
		.INIT('h8)
	) name4812 (
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		_w6058_,
		_w8859_
	);
	LUT2 #(
		.INIT('h8)
	) name4813 (
		_w6060_,
		_w8859_,
		_w8860_
	);
	LUT2 #(
		.INIT('h8)
	) name4814 (
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w6142_,
		_w8861_
	);
	LUT2 #(
		.INIT('h1)
	) name4815 (
		_w4055_,
		_w8857_,
		_w8862_
	);
	LUT2 #(
		.INIT('h1)
	) name4816 (
		_w8858_,
		_w8860_,
		_w8863_
	);
	LUT2 #(
		.INIT('h4)
	) name4817 (
		_w8861_,
		_w8863_,
		_w8864_
	);
	LUT2 #(
		.INIT('h8)
	) name4818 (
		_w8862_,
		_w8864_,
		_w8865_
	);
	LUT2 #(
		.INIT('h8)
	) name4819 (
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		_w6148_,
		_w8866_
	);
	LUT2 #(
		.INIT('h8)
	) name4820 (
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w6154_,
		_w8867_
	);
	LUT2 #(
		.INIT('h8)
	) name4821 (
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		_w6152_,
		_w8868_
	);
	LUT2 #(
		.INIT('h8)
	) name4822 (
		\core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 ,
		_w6075_,
		_w8869_
	);
	LUT2 #(
		.INIT('h8)
	) name4823 (
		_w6097_,
		_w8869_,
		_w8870_
	);
	LUT2 #(
		.INIT('h1)
	) name4824 (
		_w8866_,
		_w8867_,
		_w8871_
	);
	LUT2 #(
		.INIT('h1)
	) name4825 (
		_w8868_,
		_w8870_,
		_w8872_
	);
	LUT2 #(
		.INIT('h8)
	) name4826 (
		_w8871_,
		_w8872_,
		_w8873_
	);
	LUT2 #(
		.INIT('h8)
	) name4827 (
		_w4055_,
		_w8873_,
		_w8874_
	);
	LUT2 #(
		.INIT('h1)
	) name4828 (
		_w8865_,
		_w8874_,
		_w8875_
	);
	LUT2 #(
		.INIT('h4)
	) name4829 (
		_w6111_,
		_w8875_,
		_w8876_
	);
	LUT2 #(
		.INIT('h1)
	) name4830 (
		_w8855_,
		_w8856_,
		_w8877_
	);
	LUT2 #(
		.INIT('h4)
	) name4831 (
		_w8876_,
		_w8877_,
		_w8878_
	);
	LUT2 #(
		.INIT('h2)
	) name4832 (
		_w5949_,
		_w8878_,
		_w8879_
	);
	LUT2 #(
		.INIT('h2)
	) name4833 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		_w6934_,
		_w8880_
	);
	LUT2 #(
		.INIT('h1)
	) name4834 (
		_w8837_,
		_w8838_,
		_w8881_
	);
	LUT2 #(
		.INIT('h8)
	) name4835 (
		_w6924_,
		_w8881_,
		_w8882_
	);
	LUT2 #(
		.INIT('h4)
	) name4836 (
		_w8880_,
		_w8882_,
		_w8883_
	);
	LUT2 #(
		.INIT('h4)
	) name4837 (
		_w8879_,
		_w8883_,
		_w8884_
	);
	LUT2 #(
		.INIT('h1)
	) name4838 (
		_w6176_,
		_w8836_,
		_w8885_
	);
	LUT2 #(
		.INIT('h4)
	) name4839 (
		_w8884_,
		_w8885_,
		_w8886_
	);
	LUT2 #(
		.INIT('h8)
	) name4840 (
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w6140_,
		_w8887_
	);
	LUT2 #(
		.INIT('h8)
	) name4841 (
		\core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 ,
		_w6058_,
		_w8888_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		_w6060_,
		_w8888_,
		_w8889_
	);
	LUT2 #(
		.INIT('h8)
	) name4843 (
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w6138_,
		_w8890_
	);
	LUT2 #(
		.INIT('h8)
	) name4844 (
		\core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 ,
		_w6067_,
		_w8891_
	);
	LUT2 #(
		.INIT('h8)
	) name4845 (
		_w6068_,
		_w8891_,
		_w8892_
	);
	LUT2 #(
		.INIT('h1)
	) name4846 (
		_w4055_,
		_w8887_,
		_w8893_
	);
	LUT2 #(
		.INIT('h1)
	) name4847 (
		_w8889_,
		_w8890_,
		_w8894_
	);
	LUT2 #(
		.INIT('h4)
	) name4848 (
		_w8892_,
		_w8894_,
		_w8895_
	);
	LUT2 #(
		.INIT('h8)
	) name4849 (
		_w8893_,
		_w8895_,
		_w8896_
	);
	LUT2 #(
		.INIT('h8)
	) name4850 (
		\core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 ,
		_w6154_,
		_w8897_
	);
	LUT2 #(
		.INIT('h8)
	) name4851 (
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w6150_,
		_w8898_
	);
	LUT2 #(
		.INIT('h8)
	) name4852 (
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w6152_,
		_w8899_
	);
	LUT2 #(
		.INIT('h8)
	) name4853 (
		_w6093_,
		_w8888_,
		_w8900_
	);
	LUT2 #(
		.INIT('h1)
	) name4854 (
		_w8897_,
		_w8898_,
		_w8901_
	);
	LUT2 #(
		.INIT('h1)
	) name4855 (
		_w8899_,
		_w8900_,
		_w8902_
	);
	LUT2 #(
		.INIT('h8)
	) name4856 (
		_w8901_,
		_w8902_,
		_w8903_
	);
	LUT2 #(
		.INIT('h8)
	) name4857 (
		_w4055_,
		_w8903_,
		_w8904_
	);
	LUT2 #(
		.INIT('h1)
	) name4858 (
		_w8896_,
		_w8904_,
		_w8905_
	);
	LUT2 #(
		.INIT('h8)
	) name4859 (
		_w6176_,
		_w8905_,
		_w8906_
	);
	LUT2 #(
		.INIT('h1)
	) name4860 (
		_w6135_,
		_w8906_,
		_w8907_
	);
	LUT2 #(
		.INIT('h4)
	) name4861 (
		_w8886_,
		_w8907_,
		_w8908_
	);
	LUT2 #(
		.INIT('h8)
	) name4862 (
		\core_dag_ilm1reg_I_reg[1]/NET0131 ,
		_w6329_,
		_w8909_
	);
	LUT2 #(
		.INIT('h2)
	) name4863 (
		_w6350_,
		_w6356_,
		_w8910_
	);
	LUT2 #(
		.INIT('h4)
	) name4864 (
		_w6350_,
		_w6356_,
		_w8911_
	);
	LUT2 #(
		.INIT('h1)
	) name4865 (
		_w8910_,
		_w8911_,
		_w8912_
	);
	LUT2 #(
		.INIT('h8)
	) name4866 (
		_w7612_,
		_w8912_,
		_w8913_
	);
	LUT2 #(
		.INIT('h1)
	) name4867 (
		_w6360_,
		_w6361_,
		_w8914_
	);
	LUT2 #(
		.INIT('h1)
	) name4868 (
		_w7612_,
		_w8914_,
		_w8915_
	);
	LUT2 #(
		.INIT('h2)
	) name4869 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w8913_,
		_w8916_
	);
	LUT2 #(
		.INIT('h4)
	) name4870 (
		_w8915_,
		_w8916_,
		_w8917_
	);
	LUT2 #(
		.INIT('h2)
	) name4871 (
		_w6365_,
		_w8914_,
		_w8918_
	);
	LUT2 #(
		.INIT('h4)
	) name4872 (
		_w6365_,
		_w8914_,
		_w8919_
	);
	LUT2 #(
		.INIT('h1)
	) name4873 (
		_w8918_,
		_w8919_,
		_w8920_
	);
	LUT2 #(
		.INIT('h8)
	) name4874 (
		_w6496_,
		_w8920_,
		_w8921_
	);
	LUT2 #(
		.INIT('h4)
	) name4875 (
		_w6496_,
		_w8912_,
		_w8922_
	);
	LUT2 #(
		.INIT('h1)
	) name4876 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w8921_,
		_w8923_
	);
	LUT2 #(
		.INIT('h4)
	) name4877 (
		_w8922_,
		_w8923_,
		_w8924_
	);
	LUT2 #(
		.INIT('h1)
	) name4878 (
		_w8909_,
		_w8917_,
		_w8925_
	);
	LUT2 #(
		.INIT('h4)
	) name4879 (
		_w8924_,
		_w8925_,
		_w8926_
	);
	LUT2 #(
		.INIT('h2)
	) name4880 (
		_w6176_,
		_w8926_,
		_w8927_
	);
	LUT2 #(
		.INIT('h4)
	) name4881 (
		_w6710_,
		_w6891_,
		_w8928_
	);
	LUT2 #(
		.INIT('h2)
	) name4882 (
		_w6710_,
		_w6891_,
		_w8929_
	);
	LUT2 #(
		.INIT('h1)
	) name4883 (
		_w8928_,
		_w8929_,
		_w8930_
	);
	LUT2 #(
		.INIT('h1)
	) name4884 (
		_w6717_,
		_w8930_,
		_w8931_
	);
	LUT2 #(
		.INIT('h1)
	) name4885 (
		_w6895_,
		_w6899_,
		_w8932_
	);
	LUT2 #(
		.INIT('h8)
	) name4886 (
		_w6880_,
		_w8932_,
		_w8933_
	);
	LUT2 #(
		.INIT('h1)
	) name4887 (
		_w6880_,
		_w8932_,
		_w8934_
	);
	LUT2 #(
		.INIT('h1)
	) name4888 (
		_w8933_,
		_w8934_,
		_w8935_
	);
	LUT2 #(
		.INIT('h8)
	) name4889 (
		_w6713_,
		_w8935_,
		_w8936_
	);
	LUT2 #(
		.INIT('h2)
	) name4890 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w8936_,
		_w8937_
	);
	LUT2 #(
		.INIT('h4)
	) name4891 (
		_w8931_,
		_w8937_,
		_w8938_
	);
	LUT2 #(
		.INIT('h2)
	) name4892 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		_w6613_,
		_w8939_
	);
	LUT2 #(
		.INIT('h8)
	) name4893 (
		_w6905_,
		_w8935_,
		_w8940_
	);
	LUT2 #(
		.INIT('h1)
	) name4894 (
		_w6905_,
		_w8930_,
		_w8941_
	);
	LUT2 #(
		.INIT('h1)
	) name4895 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w8940_,
		_w8942_
	);
	LUT2 #(
		.INIT('h4)
	) name4896 (
		_w8941_,
		_w8942_,
		_w8943_
	);
	LUT2 #(
		.INIT('h1)
	) name4897 (
		_w8939_,
		_w8943_,
		_w8944_
	);
	LUT2 #(
		.INIT('h4)
	) name4898 (
		_w8938_,
		_w8944_,
		_w8945_
	);
	LUT2 #(
		.INIT('h1)
	) name4899 (
		_w6176_,
		_w8945_,
		_w8946_
	);
	LUT2 #(
		.INIT('h2)
	) name4900 (
		_w6135_,
		_w8927_,
		_w8947_
	);
	LUT2 #(
		.INIT('h4)
	) name4901 (
		_w8946_,
		_w8947_,
		_w8948_
	);
	LUT2 #(
		.INIT('h1)
	) name4902 (
		_w7005_,
		_w8908_,
		_w8949_
	);
	LUT2 #(
		.INIT('h4)
	) name4903 (
		_w8948_,
		_w8949_,
		_w8950_
	);
	LUT2 #(
		.INIT('h2)
	) name4904 (
		\core_dag_ilm1reg_I_reg[12]/NET0131 ,
		_w6470_,
		_w8951_
	);
	LUT2 #(
		.INIT('h1)
	) name4905 (
		_w6482_,
		_w6525_,
		_w8952_
	);
	LUT2 #(
		.INIT('h8)
	) name4906 (
		_w6482_,
		_w6525_,
		_w8953_
	);
	LUT2 #(
		.INIT('h1)
	) name4907 (
		_w8952_,
		_w8953_,
		_w8954_
	);
	LUT2 #(
		.INIT('h2)
	) name4908 (
		_w7631_,
		_w8954_,
		_w8955_
	);
	LUT2 #(
		.INIT('h1)
	) name4909 (
		_w6486_,
		_w6490_,
		_w8956_
	);
	LUT2 #(
		.INIT('h2)
	) name4910 (
		_w6465_,
		_w8956_,
		_w8957_
	);
	LUT2 #(
		.INIT('h4)
	) name4911 (
		_w6465_,
		_w8956_,
		_w8958_
	);
	LUT2 #(
		.INIT('h1)
	) name4912 (
		_w8957_,
		_w8958_,
		_w8959_
	);
	LUT2 #(
		.INIT('h4)
	) name4913 (
		_w7631_,
		_w8959_,
		_w8960_
	);
	LUT2 #(
		.INIT('h1)
	) name4914 (
		_w8951_,
		_w8955_,
		_w8961_
	);
	LUT2 #(
		.INIT('h4)
	) name4915 (
		_w8960_,
		_w8961_,
		_w8962_
	);
	LUT2 #(
		.INIT('h4)
	) name4916 (
		_w6135_,
		_w8962_,
		_w8963_
	);
	LUT2 #(
		.INIT('h8)
	) name4917 (
		_w6176_,
		_w7005_,
		_w8964_
	);
	LUT2 #(
		.INIT('h8)
	) name4918 (
		\DM_rdm[12]_pad ,
		_w7016_,
		_w8965_
	);
	LUT2 #(
		.INIT('h8)
	) name4919 (
		\DM_rd1[12]_pad ,
		_w7022_,
		_w8966_
	);
	LUT2 #(
		.INIT('h8)
	) name4920 (
		\DM_rd4[12]_pad ,
		_w7028_,
		_w8967_
	);
	LUT2 #(
		.INIT('h8)
	) name4921 (
		\DM_rd6[12]_pad ,
		_w7031_,
		_w8968_
	);
	LUT2 #(
		.INIT('h8)
	) name4922 (
		\DM_rd7[12]_pad ,
		_w7034_,
		_w8969_
	);
	LUT2 #(
		.INIT('h8)
	) name4923 (
		\DM_rd3[12]_pad ,
		_w7038_,
		_w8970_
	);
	LUT2 #(
		.INIT('h2)
	) name4924 (
		\DM_rd0[12]_pad ,
		_w7053_,
		_w8971_
	);
	LUT2 #(
		.INIT('h8)
	) name4925 (
		\DM_rd5[12]_pad ,
		_w7043_,
		_w8972_
	);
	LUT2 #(
		.INIT('h8)
	) name4926 (
		\DM_rd2[12]_pad ,
		_w7041_,
		_w8973_
	);
	LUT2 #(
		.INIT('h1)
	) name4927 (
		_w8966_,
		_w8970_,
		_w8974_
	);
	LUT2 #(
		.INIT('h4)
	) name4928 (
		_w8973_,
		_w8974_,
		_w8975_
	);
	LUT2 #(
		.INIT('h1)
	) name4929 (
		_w7057_,
		_w8965_,
		_w8976_
	);
	LUT2 #(
		.INIT('h1)
	) name4930 (
		_w8968_,
		_w8969_,
		_w8977_
	);
	LUT2 #(
		.INIT('h8)
	) name4931 (
		_w8976_,
		_w8977_,
		_w8978_
	);
	LUT2 #(
		.INIT('h4)
	) name4932 (
		_w8967_,
		_w8975_,
		_w8979_
	);
	LUT2 #(
		.INIT('h4)
	) name4933 (
		_w8972_,
		_w8979_,
		_w8980_
	);
	LUT2 #(
		.INIT('h8)
	) name4934 (
		_w8978_,
		_w8980_,
		_w8981_
	);
	LUT2 #(
		.INIT('h4)
	) name4935 (
		_w8971_,
		_w8981_,
		_w8982_
	);
	LUT2 #(
		.INIT('h8)
	) name4936 (
		\regout_STD_C_reg[12]/P0001 ,
		_w6988_,
		_w8983_
	);
	LUT2 #(
		.INIT('h8)
	) name4937 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131 ,
		_w8984_
	);
	LUT2 #(
		.INIT('h8)
	) name4938 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w8985_
	);
	LUT2 #(
		.INIT('h8)
	) name4939 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		_w8986_
	);
	LUT2 #(
		.INIT('h8)
	) name4940 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131 ,
		_w8987_
	);
	LUT2 #(
		.INIT('h8)
	) name4941 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131 ,
		_w8988_
	);
	LUT2 #(
		.INIT('h8)
	) name4942 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		_w8989_
	);
	LUT2 #(
		.INIT('h8)
	) name4943 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131 ,
		_w8990_
	);
	LUT2 #(
		.INIT('h8)
	) name4944 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131 ,
		_w8991_
	);
	LUT2 #(
		.INIT('h8)
	) name4945 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131 ,
		_w8992_
	);
	LUT2 #(
		.INIT('h8)
	) name4946 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[12]/NET0131 ,
		_w8993_
	);
	LUT2 #(
		.INIT('h8)
	) name4947 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131 ,
		_w8994_
	);
	LUT2 #(
		.INIT('h8)
	) name4948 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131 ,
		_w8995_
	);
	LUT2 #(
		.INIT('h1)
	) name4949 (
		_w8984_,
		_w8985_,
		_w8996_
	);
	LUT2 #(
		.INIT('h1)
	) name4950 (
		_w8986_,
		_w8987_,
		_w8997_
	);
	LUT2 #(
		.INIT('h1)
	) name4951 (
		_w8988_,
		_w8989_,
		_w8998_
	);
	LUT2 #(
		.INIT('h1)
	) name4952 (
		_w8990_,
		_w8991_,
		_w8999_
	);
	LUT2 #(
		.INIT('h1)
	) name4953 (
		_w8992_,
		_w8993_,
		_w9000_
	);
	LUT2 #(
		.INIT('h1)
	) name4954 (
		_w8994_,
		_w8995_,
		_w9001_
	);
	LUT2 #(
		.INIT('h8)
	) name4955 (
		_w9000_,
		_w9001_,
		_w9002_
	);
	LUT2 #(
		.INIT('h8)
	) name4956 (
		_w8998_,
		_w8999_,
		_w9003_
	);
	LUT2 #(
		.INIT('h8)
	) name4957 (
		_w8996_,
		_w8997_,
		_w9004_
	);
	LUT2 #(
		.INIT('h8)
	) name4958 (
		_w9003_,
		_w9004_,
		_w9005_
	);
	LUT2 #(
		.INIT('h8)
	) name4959 (
		_w9002_,
		_w9005_,
		_w9006_
	);
	LUT2 #(
		.INIT('h2)
	) name4960 (
		_w7068_,
		_w9006_,
		_w9007_
	);
	LUT2 #(
		.INIT('h8)
	) name4961 (
		\memc_usysr_DO_reg[12]/NET0131 ,
		_w7301_,
		_w9008_
	);
	LUT2 #(
		.INIT('h8)
	) name4962 (
		\sport0_regs_AUTO_a_reg[12]/NET0131 ,
		_w7295_,
		_w9009_
	);
	LUT2 #(
		.INIT('h8)
	) name4963 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w7234_,
		_w9010_
	);
	LUT2 #(
		.INIT('h8)
	) name4964 (
		\bdma_BCTL_reg[12]/NET0131 ,
		_w7230_,
		_w9011_
	);
	LUT2 #(
		.INIT('h8)
	) name4965 (
		\emc_WSCRreg_DO_reg[12]/NET0131 ,
		_w7251_,
		_w9012_
	);
	LUT2 #(
		.INIT('h8)
	) name4966 (
		\sport1_rxctl_SLOT1_EXT_reg[2]/NET0131 ,
		_w7689_,
		_w9013_
	);
	LUT2 #(
		.INIT('h8)
	) name4967 (
		\clkc_ckr_reg_DO_reg[12]/NET0131 ,
		_w7239_,
		_w9014_
	);
	LUT2 #(
		.INIT('h8)
	) name4968 (
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w7249_,
		_w9015_
	);
	LUT2 #(
		.INIT('h8)
	) name4969 (
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w7273_,
		_w9016_
	);
	LUT2 #(
		.INIT('h8)
	) name4970 (
		\PIO_out[8]_pad ,
		_w7291_,
		_w9017_
	);
	LUT2 #(
		.INIT('h8)
	) name4971 (
		\PIO_oe[8]_pad ,
		_w7244_,
		_w9018_
	);
	LUT2 #(
		.INIT('h8)
	) name4972 (
		\tm_tpr_reg_DO_reg[12]/NET0131 ,
		_w7293_,
		_w9019_
	);
	LUT2 #(
		.INIT('h8)
	) name4973 (
		\pio_PINT_reg[8]/NET0131 ,
		_w7271_,
		_w9020_
	);
	LUT2 #(
		.INIT('h8)
	) name4974 (
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w7259_,
		_w9021_
	);
	LUT2 #(
		.INIT('h8)
	) name4975 (
		\bdma_BEAD_reg[12]/NET0131 ,
		_w7303_,
		_w9022_
	);
	LUT2 #(
		.INIT('h8)
	) name4976 (
		\pio_pmask_reg_DO_reg[8]/NET0131 ,
		_w7297_,
		_w9023_
	);
	LUT2 #(
		.INIT('h8)
	) name4977 (
		\tm_TCR_TMP_reg[12]/NET0131 ,
		_w7289_,
		_w9024_
	);
	LUT2 #(
		.INIT('h8)
	) name4978 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w7299_,
		_w9025_
	);
	LUT2 #(
		.INIT('h8)
	) name4979 (
		\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w7256_,
		_w9026_
	);
	LUT2 #(
		.INIT('h8)
	) name4980 (
		\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w7247_,
		_w9027_
	);
	LUT2 #(
		.INIT('h8)
	) name4981 (
		\sport0_rxctl_SLOT1_EXT_reg[2]/NET0131 ,
		_w7710_,
		_w9028_
	);
	LUT2 #(
		.INIT('h8)
	) name4982 (
		\bdma_BWCOUNT_reg[12]/NET0131 ,
		_w7287_,
		_w9029_
	);
	LUT2 #(
		.INIT('h8)
	) name4983 (
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w7281_,
		_w9030_
	);
	LUT2 #(
		.INIT('h1)
	) name4984 (
		_w9008_,
		_w9009_,
		_w9031_
	);
	LUT2 #(
		.INIT('h1)
	) name4985 (
		_w9012_,
		_w9014_,
		_w9032_
	);
	LUT2 #(
		.INIT('h1)
	) name4986 (
		_w9015_,
		_w9016_,
		_w9033_
	);
	LUT2 #(
		.INIT('h1)
	) name4987 (
		_w9017_,
		_w9018_,
		_w9034_
	);
	LUT2 #(
		.INIT('h1)
	) name4988 (
		_w9019_,
		_w9020_,
		_w9035_
	);
	LUT2 #(
		.INIT('h1)
	) name4989 (
		_w9021_,
		_w9023_,
		_w9036_
	);
	LUT2 #(
		.INIT('h1)
	) name4990 (
		_w9024_,
		_w9025_,
		_w9037_
	);
	LUT2 #(
		.INIT('h1)
	) name4991 (
		_w9026_,
		_w9027_,
		_w9038_
	);
	LUT2 #(
		.INIT('h4)
	) name4992 (
		_w9030_,
		_w9038_,
		_w9039_
	);
	LUT2 #(
		.INIT('h8)
	) name4993 (
		_w9036_,
		_w9037_,
		_w9040_
	);
	LUT2 #(
		.INIT('h8)
	) name4994 (
		_w9034_,
		_w9035_,
		_w9041_
	);
	LUT2 #(
		.INIT('h8)
	) name4995 (
		_w9032_,
		_w9033_,
		_w9042_
	);
	LUT2 #(
		.INIT('h4)
	) name4996 (
		_w9013_,
		_w9031_,
		_w9043_
	);
	LUT2 #(
		.INIT('h4)
	) name4997 (
		_w9028_,
		_w9043_,
		_w9044_
	);
	LUT2 #(
		.INIT('h8)
	) name4998 (
		_w9041_,
		_w9042_,
		_w9045_
	);
	LUT2 #(
		.INIT('h8)
	) name4999 (
		_w9039_,
		_w9040_,
		_w9046_
	);
	LUT2 #(
		.INIT('h8)
	) name5000 (
		_w9045_,
		_w9046_,
		_w9047_
	);
	LUT2 #(
		.INIT('h4)
	) name5001 (
		_w9010_,
		_w9044_,
		_w9048_
	);
	LUT2 #(
		.INIT('h1)
	) name5002 (
		_w9011_,
		_w9022_,
		_w9049_
	);
	LUT2 #(
		.INIT('h8)
	) name5003 (
		_w9048_,
		_w9049_,
		_w9050_
	);
	LUT2 #(
		.INIT('h4)
	) name5004 (
		_w9029_,
		_w9047_,
		_w9051_
	);
	LUT2 #(
		.INIT('h8)
	) name5005 (
		_w9050_,
		_w9051_,
		_w9052_
	);
	LUT2 #(
		.INIT('h2)
	) name5006 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w9052_,
		_w9053_
	);
	LUT2 #(
		.INIT('h4)
	) name5007 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001 ,
		_w9054_
	);
	LUT2 #(
		.INIT('h8)
	) name5008 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 ,
		_w9055_
	);
	LUT2 #(
		.INIT('h1)
	) name5009 (
		_w9054_,
		_w9055_,
		_w9056_
	);
	LUT2 #(
		.INIT('h2)
	) name5010 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w9056_,
		_w9057_
	);
	LUT2 #(
		.INIT('h4)
	) name5011 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001 ,
		_w9058_
	);
	LUT2 #(
		.INIT('h8)
	) name5012 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001 ,
		_w9059_
	);
	LUT2 #(
		.INIT('h1)
	) name5013 (
		_w9058_,
		_w9059_,
		_w9060_
	);
	LUT2 #(
		.INIT('h2)
	) name5014 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w9060_,
		_w9061_
	);
	LUT2 #(
		.INIT('h4)
	) name5015 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001 ,
		_w9062_
	);
	LUT2 #(
		.INIT('h8)
	) name5016 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001 ,
		_w9063_
	);
	LUT2 #(
		.INIT('h1)
	) name5017 (
		_w9062_,
		_w9063_,
		_w9064_
	);
	LUT2 #(
		.INIT('h2)
	) name5018 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w9064_,
		_w9065_
	);
	LUT2 #(
		.INIT('h4)
	) name5019 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001 ,
		_w9066_
	);
	LUT2 #(
		.INIT('h8)
	) name5020 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001 ,
		_w9067_
	);
	LUT2 #(
		.INIT('h1)
	) name5021 (
		_w9066_,
		_w9067_,
		_w9068_
	);
	LUT2 #(
		.INIT('h2)
	) name5022 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w9068_,
		_w9069_
	);
	LUT2 #(
		.INIT('h4)
	) name5023 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001 ,
		_w9070_
	);
	LUT2 #(
		.INIT('h8)
	) name5024 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 ,
		_w9071_
	);
	LUT2 #(
		.INIT('h1)
	) name5025 (
		_w9070_,
		_w9071_,
		_w9072_
	);
	LUT2 #(
		.INIT('h2)
	) name5026 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w9072_,
		_w9073_
	);
	LUT2 #(
		.INIT('h4)
	) name5027 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001 ,
		_w9074_
	);
	LUT2 #(
		.INIT('h8)
	) name5028 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001 ,
		_w9075_
	);
	LUT2 #(
		.INIT('h1)
	) name5029 (
		_w9074_,
		_w9075_,
		_w9076_
	);
	LUT2 #(
		.INIT('h2)
	) name5030 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w9076_,
		_w9077_
	);
	LUT2 #(
		.INIT('h1)
	) name5031 (
		_w7207_,
		_w9057_,
		_w9078_
	);
	LUT2 #(
		.INIT('h1)
	) name5032 (
		_w9061_,
		_w9065_,
		_w9079_
	);
	LUT2 #(
		.INIT('h1)
	) name5033 (
		_w9069_,
		_w9073_,
		_w9080_
	);
	LUT2 #(
		.INIT('h4)
	) name5034 (
		_w9077_,
		_w9080_,
		_w9081_
	);
	LUT2 #(
		.INIT('h8)
	) name5035 (
		_w9078_,
		_w9079_,
		_w9082_
	);
	LUT2 #(
		.INIT('h8)
	) name5036 (
		_w9081_,
		_w9082_,
		_w9083_
	);
	LUT2 #(
		.INIT('h2)
	) name5037 (
		_w7179_,
		_w9083_,
		_w9084_
	);
	LUT2 #(
		.INIT('h4)
	) name5038 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001 ,
		_w9085_
	);
	LUT2 #(
		.INIT('h8)
	) name5039 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001 ,
		_w9086_
	);
	LUT2 #(
		.INIT('h1)
	) name5040 (
		_w9085_,
		_w9086_,
		_w9087_
	);
	LUT2 #(
		.INIT('h2)
	) name5041 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w9087_,
		_w9088_
	);
	LUT2 #(
		.INIT('h4)
	) name5042 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001 ,
		_w9089_
	);
	LUT2 #(
		.INIT('h8)
	) name5043 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001 ,
		_w9090_
	);
	LUT2 #(
		.INIT('h1)
	) name5044 (
		_w9089_,
		_w9090_,
		_w9091_
	);
	LUT2 #(
		.INIT('h2)
	) name5045 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w9091_,
		_w9092_
	);
	LUT2 #(
		.INIT('h4)
	) name5046 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001 ,
		_w9093_
	);
	LUT2 #(
		.INIT('h8)
	) name5047 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001 ,
		_w9094_
	);
	LUT2 #(
		.INIT('h1)
	) name5048 (
		_w9093_,
		_w9094_,
		_w9095_
	);
	LUT2 #(
		.INIT('h2)
	) name5049 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w9095_,
		_w9096_
	);
	LUT2 #(
		.INIT('h4)
	) name5050 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001 ,
		_w9097_
	);
	LUT2 #(
		.INIT('h8)
	) name5051 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001 ,
		_w9098_
	);
	LUT2 #(
		.INIT('h1)
	) name5052 (
		_w9097_,
		_w9098_,
		_w9099_
	);
	LUT2 #(
		.INIT('h2)
	) name5053 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w9099_,
		_w9100_
	);
	LUT2 #(
		.INIT('h4)
	) name5054 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001 ,
		_w9101_
	);
	LUT2 #(
		.INIT('h8)
	) name5055 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001 ,
		_w9102_
	);
	LUT2 #(
		.INIT('h1)
	) name5056 (
		_w9101_,
		_w9102_,
		_w9103_
	);
	LUT2 #(
		.INIT('h2)
	) name5057 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w9103_,
		_w9104_
	);
	LUT2 #(
		.INIT('h1)
	) name5058 (
		_w9088_,
		_w9092_,
		_w9105_
	);
	LUT2 #(
		.INIT('h1)
	) name5059 (
		_w9096_,
		_w9100_,
		_w9106_
	);
	LUT2 #(
		.INIT('h4)
	) name5060 (
		_w9104_,
		_w9106_,
		_w9107_
	);
	LUT2 #(
		.INIT('h8)
	) name5061 (
		_w9105_,
		_w9107_,
		_w9108_
	);
	LUT2 #(
		.INIT('h2)
	) name5062 (
		_w7093_,
		_w9108_,
		_w9109_
	);
	LUT2 #(
		.INIT('h2)
	) name5063 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w7216_,
		_w9110_
	);
	LUT2 #(
		.INIT('h8)
	) name5064 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w9111_
	);
	LUT2 #(
		.INIT('h8)
	) name5065 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w9112_
	);
	LUT2 #(
		.INIT('h2)
	) name5066 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4694_,
		_w9113_
	);
	LUT2 #(
		.INIT('h1)
	) name5067 (
		_w9111_,
		_w9112_,
		_w9114_
	);
	LUT2 #(
		.INIT('h4)
	) name5068 (
		_w9110_,
		_w9114_,
		_w9115_
	);
	LUT2 #(
		.INIT('h4)
	) name5069 (
		_w9113_,
		_w9115_,
		_w9116_
	);
	LUT2 #(
		.INIT('h2)
	) name5070 (
		_w7215_,
		_w9116_,
		_w9117_
	);
	LUT2 #(
		.INIT('h4)
	) name5071 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 ,
		_w9118_
	);
	LUT2 #(
		.INIT('h8)
	) name5072 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 ,
		_w9119_
	);
	LUT2 #(
		.INIT('h1)
	) name5073 (
		_w9118_,
		_w9119_,
		_w9120_
	);
	LUT2 #(
		.INIT('h2)
	) name5074 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w9120_,
		_w9121_
	);
	LUT2 #(
		.INIT('h4)
	) name5075 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001 ,
		_w9122_
	);
	LUT2 #(
		.INIT('h8)
	) name5076 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001 ,
		_w9123_
	);
	LUT2 #(
		.INIT('h1)
	) name5077 (
		_w9122_,
		_w9123_,
		_w9124_
	);
	LUT2 #(
		.INIT('h2)
	) name5078 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w9124_,
		_w9125_
	);
	LUT2 #(
		.INIT('h4)
	) name5079 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 ,
		_w9126_
	);
	LUT2 #(
		.INIT('h8)
	) name5080 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 ,
		_w9127_
	);
	LUT2 #(
		.INIT('h1)
	) name5081 (
		_w9126_,
		_w9127_,
		_w9128_
	);
	LUT2 #(
		.INIT('h2)
	) name5082 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w9128_,
		_w9129_
	);
	LUT2 #(
		.INIT('h1)
	) name5083 (
		_w9121_,
		_w9125_,
		_w9130_
	);
	LUT2 #(
		.INIT('h4)
	) name5084 (
		_w9129_,
		_w9130_,
		_w9131_
	);
	LUT2 #(
		.INIT('h8)
	) name5085 (
		_w7174_,
		_w9131_,
		_w9132_
	);
	LUT2 #(
		.INIT('h2)
	) name5086 (
		_w7153_,
		_w9132_,
		_w9133_
	);
	LUT2 #(
		.INIT('h8)
	) name5087 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[12]/P0001 ,
		_w9134_
	);
	LUT2 #(
		.INIT('h8)
	) name5088 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[12]/P0001 ,
		_w9135_
	);
	LUT2 #(
		.INIT('h8)
	) name5089 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[12]/P0001 ,
		_w9136_
	);
	LUT2 #(
		.INIT('h8)
	) name5090 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[12]/P0001 ,
		_w9137_
	);
	LUT2 #(
		.INIT('h1)
	) name5091 (
		_w9134_,
		_w9135_,
		_w9138_
	);
	LUT2 #(
		.INIT('h1)
	) name5092 (
		_w9136_,
		_w9137_,
		_w9139_
	);
	LUT2 #(
		.INIT('h8)
	) name5093 (
		_w9138_,
		_w9139_,
		_w9140_
	);
	LUT2 #(
		.INIT('h2)
	) name5094 (
		_w7119_,
		_w9140_,
		_w9141_
	);
	LUT2 #(
		.INIT('h8)
	) name5095 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w9142_
	);
	LUT2 #(
		.INIT('h8)
	) name5096 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131 ,
		_w9143_
	);
	LUT2 #(
		.INIT('h8)
	) name5097 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131 ,
		_w9144_
	);
	LUT2 #(
		.INIT('h8)
	) name5098 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131 ,
		_w9145_
	);
	LUT2 #(
		.INIT('h8)
	) name5099 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131 ,
		_w9146_
	);
	LUT2 #(
		.INIT('h8)
	) name5100 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131 ,
		_w9147_
	);
	LUT2 #(
		.INIT('h8)
	) name5101 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		_w9148_
	);
	LUT2 #(
		.INIT('h8)
	) name5102 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131 ,
		_w9149_
	);
	LUT2 #(
		.INIT('h8)
	) name5103 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131 ,
		_w9150_
	);
	LUT2 #(
		.INIT('h8)
	) name5104 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131 ,
		_w9151_
	);
	LUT2 #(
		.INIT('h8)
	) name5105 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w9152_
	);
	LUT2 #(
		.INIT('h8)
	) name5106 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w9153_
	);
	LUT2 #(
		.INIT('h1)
	) name5107 (
		_w9142_,
		_w9143_,
		_w9154_
	);
	LUT2 #(
		.INIT('h1)
	) name5108 (
		_w9144_,
		_w9145_,
		_w9155_
	);
	LUT2 #(
		.INIT('h1)
	) name5109 (
		_w9146_,
		_w9147_,
		_w9156_
	);
	LUT2 #(
		.INIT('h1)
	) name5110 (
		_w9148_,
		_w9149_,
		_w9157_
	);
	LUT2 #(
		.INIT('h1)
	) name5111 (
		_w9150_,
		_w9151_,
		_w9158_
	);
	LUT2 #(
		.INIT('h1)
	) name5112 (
		_w9152_,
		_w9153_,
		_w9159_
	);
	LUT2 #(
		.INIT('h8)
	) name5113 (
		_w9158_,
		_w9159_,
		_w9160_
	);
	LUT2 #(
		.INIT('h8)
	) name5114 (
		_w9156_,
		_w9157_,
		_w9161_
	);
	LUT2 #(
		.INIT('h8)
	) name5115 (
		_w9154_,
		_w9155_,
		_w9162_
	);
	LUT2 #(
		.INIT('h8)
	) name5116 (
		_w9161_,
		_w9162_,
		_w9163_
	);
	LUT2 #(
		.INIT('h8)
	) name5117 (
		_w9160_,
		_w9163_,
		_w9164_
	);
	LUT2 #(
		.INIT('h2)
	) name5118 (
		_w7128_,
		_w9164_,
		_w9165_
	);
	LUT2 #(
		.INIT('h1)
	) name5119 (
		_w9007_,
		_w9141_,
		_w9166_
	);
	LUT2 #(
		.INIT('h4)
	) name5120 (
		_w9165_,
		_w9166_,
		_w9167_
	);
	LUT2 #(
		.INIT('h1)
	) name5121 (
		_w9084_,
		_w9109_,
		_w9168_
	);
	LUT2 #(
		.INIT('h4)
	) name5122 (
		_w9133_,
		_w9168_,
		_w9169_
	);
	LUT2 #(
		.INIT('h8)
	) name5123 (
		_w9167_,
		_w9169_,
		_w9170_
	);
	LUT2 #(
		.INIT('h4)
	) name5124 (
		_w9053_,
		_w9170_,
		_w9171_
	);
	LUT2 #(
		.INIT('h4)
	) name5125 (
		_w9117_,
		_w9171_,
		_w9172_
	);
	LUT2 #(
		.INIT('h4)
	) name5126 (
		_w8983_,
		_w9172_,
		_w9173_
	);
	LUT2 #(
		.INIT('h1)
	) name5127 (
		\emc_DMDoe_reg/NET0131 ,
		_w9173_,
		_w9174_
	);
	LUT2 #(
		.INIT('h8)
	) name5128 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[12]/P0001 ,
		_w9175_
	);
	LUT2 #(
		.INIT('h2)
	) name5129 (
		_w7057_,
		_w9175_,
		_w9176_
	);
	LUT2 #(
		.INIT('h4)
	) name5130 (
		_w9174_,
		_w9176_,
		_w9177_
	);
	LUT2 #(
		.INIT('h1)
	) name5131 (
		_w8982_,
		_w9177_,
		_w9178_
	);
	LUT2 #(
		.INIT('h2)
	) name5132 (
		_w6135_,
		_w9178_,
		_w9179_
	);
	LUT2 #(
		.INIT('h2)
	) name5133 (
		_w8964_,
		_w9179_,
		_w9180_
	);
	LUT2 #(
		.INIT('h4)
	) name5134 (
		_w8963_,
		_w9180_,
		_w9181_
	);
	LUT2 #(
		.INIT('h2)
	) name5135 (
		_w8854_,
		_w8875_,
		_w9182_
	);
	LUT2 #(
		.INIT('h2)
	) name5136 (
		_w8153_,
		_w9182_,
		_w9183_
	);
	LUT2 #(
		.INIT('h8)
	) name5137 (
		\DM_rdm[1]_pad ,
		_w7016_,
		_w9184_
	);
	LUT2 #(
		.INIT('h8)
	) name5138 (
		\DM_rd1[1]_pad ,
		_w7022_,
		_w9185_
	);
	LUT2 #(
		.INIT('h8)
	) name5139 (
		\DM_rd4[1]_pad ,
		_w7028_,
		_w9186_
	);
	LUT2 #(
		.INIT('h8)
	) name5140 (
		\DM_rd6[1]_pad ,
		_w7031_,
		_w9187_
	);
	LUT2 #(
		.INIT('h8)
	) name5141 (
		\DM_rd7[1]_pad ,
		_w7034_,
		_w9188_
	);
	LUT2 #(
		.INIT('h8)
	) name5142 (
		\DM_rd3[1]_pad ,
		_w7038_,
		_w9189_
	);
	LUT2 #(
		.INIT('h2)
	) name5143 (
		\DM_rd0[1]_pad ,
		_w7053_,
		_w9190_
	);
	LUT2 #(
		.INIT('h8)
	) name5144 (
		\DM_rd5[1]_pad ,
		_w7043_,
		_w9191_
	);
	LUT2 #(
		.INIT('h8)
	) name5145 (
		\DM_rd2[1]_pad ,
		_w7041_,
		_w9192_
	);
	LUT2 #(
		.INIT('h1)
	) name5146 (
		_w9185_,
		_w9189_,
		_w9193_
	);
	LUT2 #(
		.INIT('h4)
	) name5147 (
		_w9192_,
		_w9193_,
		_w9194_
	);
	LUT2 #(
		.INIT('h1)
	) name5148 (
		_w7057_,
		_w9184_,
		_w9195_
	);
	LUT2 #(
		.INIT('h1)
	) name5149 (
		_w9187_,
		_w9188_,
		_w9196_
	);
	LUT2 #(
		.INIT('h8)
	) name5150 (
		_w9195_,
		_w9196_,
		_w9197_
	);
	LUT2 #(
		.INIT('h4)
	) name5151 (
		_w9186_,
		_w9194_,
		_w9198_
	);
	LUT2 #(
		.INIT('h4)
	) name5152 (
		_w9191_,
		_w9198_,
		_w9199_
	);
	LUT2 #(
		.INIT('h8)
	) name5153 (
		_w9197_,
		_w9199_,
		_w9200_
	);
	LUT2 #(
		.INIT('h4)
	) name5154 (
		_w9190_,
		_w9200_,
		_w9201_
	);
	LUT2 #(
		.INIT('h8)
	) name5155 (
		\regout_STD_C_reg[1]/P0001 ,
		_w6988_,
		_w9202_
	);
	LUT2 #(
		.INIT('h4)
	) name5156 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001 ,
		_w9203_
	);
	LUT2 #(
		.INIT('h8)
	) name5157 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 ,
		_w9204_
	);
	LUT2 #(
		.INIT('h1)
	) name5158 (
		_w9203_,
		_w9204_,
		_w9205_
	);
	LUT2 #(
		.INIT('h2)
	) name5159 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w9205_,
		_w9206_
	);
	LUT2 #(
		.INIT('h4)
	) name5160 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001 ,
		_w9207_
	);
	LUT2 #(
		.INIT('h8)
	) name5161 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001 ,
		_w9208_
	);
	LUT2 #(
		.INIT('h1)
	) name5162 (
		_w9207_,
		_w9208_,
		_w9209_
	);
	LUT2 #(
		.INIT('h2)
	) name5163 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w9209_,
		_w9210_
	);
	LUT2 #(
		.INIT('h4)
	) name5164 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001 ,
		_w9211_
	);
	LUT2 #(
		.INIT('h8)
	) name5165 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001 ,
		_w9212_
	);
	LUT2 #(
		.INIT('h1)
	) name5166 (
		_w9211_,
		_w9212_,
		_w9213_
	);
	LUT2 #(
		.INIT('h2)
	) name5167 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w9213_,
		_w9214_
	);
	LUT2 #(
		.INIT('h4)
	) name5168 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001 ,
		_w9215_
	);
	LUT2 #(
		.INIT('h8)
	) name5169 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001 ,
		_w9216_
	);
	LUT2 #(
		.INIT('h1)
	) name5170 (
		_w9215_,
		_w9216_,
		_w9217_
	);
	LUT2 #(
		.INIT('h2)
	) name5171 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w9217_,
		_w9218_
	);
	LUT2 #(
		.INIT('h4)
	) name5172 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001 ,
		_w9219_
	);
	LUT2 #(
		.INIT('h8)
	) name5173 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001 ,
		_w9220_
	);
	LUT2 #(
		.INIT('h1)
	) name5174 (
		_w9219_,
		_w9220_,
		_w9221_
	);
	LUT2 #(
		.INIT('h2)
	) name5175 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w9221_,
		_w9222_
	);
	LUT2 #(
		.INIT('h4)
	) name5176 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001 ,
		_w9223_
	);
	LUT2 #(
		.INIT('h8)
	) name5177 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 ,
		_w9224_
	);
	LUT2 #(
		.INIT('h1)
	) name5178 (
		_w9223_,
		_w9224_,
		_w9225_
	);
	LUT2 #(
		.INIT('h2)
	) name5179 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w9225_,
		_w9226_
	);
	LUT2 #(
		.INIT('h4)
	) name5180 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 ,
		_w9227_
	);
	LUT2 #(
		.INIT('h8)
	) name5181 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 ,
		_w9228_
	);
	LUT2 #(
		.INIT('h1)
	) name5182 (
		_w9227_,
		_w9228_,
		_w9229_
	);
	LUT2 #(
		.INIT('h2)
	) name5183 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w9229_,
		_w9230_
	);
	LUT2 #(
		.INIT('h1)
	) name5184 (
		_w9206_,
		_w9210_,
		_w9231_
	);
	LUT2 #(
		.INIT('h1)
	) name5185 (
		_w9214_,
		_w9218_,
		_w9232_
	);
	LUT2 #(
		.INIT('h1)
	) name5186 (
		_w9222_,
		_w9226_,
		_w9233_
	);
	LUT2 #(
		.INIT('h4)
	) name5187 (
		_w9230_,
		_w9233_,
		_w9234_
	);
	LUT2 #(
		.INIT('h8)
	) name5188 (
		_w9231_,
		_w9232_,
		_w9235_
	);
	LUT2 #(
		.INIT('h8)
	) name5189 (
		_w9234_,
		_w9235_,
		_w9236_
	);
	LUT2 #(
		.INIT('h2)
	) name5190 (
		_w7179_,
		_w9236_,
		_w9237_
	);
	LUT2 #(
		.INIT('h8)
	) name5191 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131 ,
		_w9238_
	);
	LUT2 #(
		.INIT('h8)
	) name5192 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131 ,
		_w9239_
	);
	LUT2 #(
		.INIT('h8)
	) name5193 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131 ,
		_w9240_
	);
	LUT2 #(
		.INIT('h8)
	) name5194 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131 ,
		_w9241_
	);
	LUT2 #(
		.INIT('h8)
	) name5195 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[1]/NET0131 ,
		_w9242_
	);
	LUT2 #(
		.INIT('h8)
	) name5196 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w9243_
	);
	LUT2 #(
		.INIT('h8)
	) name5197 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131 ,
		_w9244_
	);
	LUT2 #(
		.INIT('h8)
	) name5198 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131 ,
		_w9245_
	);
	LUT2 #(
		.INIT('h8)
	) name5199 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 ,
		_w9246_
	);
	LUT2 #(
		.INIT('h8)
	) name5200 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w9247_
	);
	LUT2 #(
		.INIT('h8)
	) name5201 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131 ,
		_w9248_
	);
	LUT2 #(
		.INIT('h8)
	) name5202 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131 ,
		_w9249_
	);
	LUT2 #(
		.INIT('h1)
	) name5203 (
		_w9238_,
		_w9239_,
		_w9250_
	);
	LUT2 #(
		.INIT('h1)
	) name5204 (
		_w9240_,
		_w9241_,
		_w9251_
	);
	LUT2 #(
		.INIT('h1)
	) name5205 (
		_w9242_,
		_w9243_,
		_w9252_
	);
	LUT2 #(
		.INIT('h1)
	) name5206 (
		_w9244_,
		_w9245_,
		_w9253_
	);
	LUT2 #(
		.INIT('h1)
	) name5207 (
		_w9246_,
		_w9247_,
		_w9254_
	);
	LUT2 #(
		.INIT('h1)
	) name5208 (
		_w9248_,
		_w9249_,
		_w9255_
	);
	LUT2 #(
		.INIT('h8)
	) name5209 (
		_w9254_,
		_w9255_,
		_w9256_
	);
	LUT2 #(
		.INIT('h8)
	) name5210 (
		_w9252_,
		_w9253_,
		_w9257_
	);
	LUT2 #(
		.INIT('h8)
	) name5211 (
		_w9250_,
		_w9251_,
		_w9258_
	);
	LUT2 #(
		.INIT('h8)
	) name5212 (
		_w9257_,
		_w9258_,
		_w9259_
	);
	LUT2 #(
		.INIT('h8)
	) name5213 (
		_w9256_,
		_w9259_,
		_w9260_
	);
	LUT2 #(
		.INIT('h2)
	) name5214 (
		_w7068_,
		_w9260_,
		_w9261_
	);
	LUT2 #(
		.INIT('h4)
	) name5215 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001 ,
		_w9262_
	);
	LUT2 #(
		.INIT('h8)
	) name5216 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001 ,
		_w9263_
	);
	LUT2 #(
		.INIT('h1)
	) name5217 (
		_w9262_,
		_w9263_,
		_w9264_
	);
	LUT2 #(
		.INIT('h2)
	) name5218 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w9264_,
		_w9265_
	);
	LUT2 #(
		.INIT('h4)
	) name5219 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBr_reg[1]/P0001 ,
		_w9266_
	);
	LUT2 #(
		.INIT('h8)
	) name5220 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_SBs_reg[1]/P0001 ,
		_w9267_
	);
	LUT2 #(
		.INIT('h1)
	) name5221 (
		_w9266_,
		_w9267_,
		_w9268_
	);
	LUT2 #(
		.INIT('h2)
	) name5222 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		_w9268_,
		_w9269_
	);
	LUT2 #(
		.INIT('h4)
	) name5223 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001 ,
		_w9270_
	);
	LUT2 #(
		.INIT('h8)
	) name5224 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001 ,
		_w9271_
	);
	LUT2 #(
		.INIT('h1)
	) name5225 (
		_w9270_,
		_w9271_,
		_w9272_
	);
	LUT2 #(
		.INIT('h2)
	) name5226 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w9272_,
		_w9273_
	);
	LUT2 #(
		.INIT('h4)
	) name5227 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 ,
		_w9274_
	);
	LUT2 #(
		.INIT('h8)
	) name5228 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 ,
		_w9275_
	);
	LUT2 #(
		.INIT('h1)
	) name5229 (
		_w9274_,
		_w9275_,
		_w9276_
	);
	LUT2 #(
		.INIT('h2)
	) name5230 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w9276_,
		_w9277_
	);
	LUT2 #(
		.INIT('h4)
	) name5231 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 ,
		_w9278_
	);
	LUT2 #(
		.INIT('h8)
	) name5232 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 ,
		_w9279_
	);
	LUT2 #(
		.INIT('h1)
	) name5233 (
		_w9278_,
		_w9279_,
		_w9280_
	);
	LUT2 #(
		.INIT('h2)
	) name5234 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w9280_,
		_w9281_
	);
	LUT2 #(
		.INIT('h1)
	) name5235 (
		_w9265_,
		_w9269_,
		_w9282_
	);
	LUT2 #(
		.INIT('h1)
	) name5236 (
		_w9273_,
		_w9277_,
		_w9283_
	);
	LUT2 #(
		.INIT('h4)
	) name5237 (
		_w9281_,
		_w9283_,
		_w9284_
	);
	LUT2 #(
		.INIT('h8)
	) name5238 (
		_w9282_,
		_w9284_,
		_w9285_
	);
	LUT2 #(
		.INIT('h2)
	) name5239 (
		_w7153_,
		_w9285_,
		_w9286_
	);
	LUT2 #(
		.INIT('h8)
	) name5240 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[1]/P0001 ,
		_w9287_
	);
	LUT2 #(
		.INIT('h8)
	) name5241 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w9288_
	);
	LUT2 #(
		.INIT('h8)
	) name5242 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[1]/P0001 ,
		_w9289_
	);
	LUT2 #(
		.INIT('h8)
	) name5243 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		_w9290_
	);
	LUT2 #(
		.INIT('h1)
	) name5244 (
		_w9287_,
		_w9288_,
		_w9291_
	);
	LUT2 #(
		.INIT('h1)
	) name5245 (
		_w9289_,
		_w9290_,
		_w9292_
	);
	LUT2 #(
		.INIT('h8)
	) name5246 (
		_w9291_,
		_w9292_,
		_w9293_
	);
	LUT2 #(
		.INIT('h2)
	) name5247 (
		_w7119_,
		_w9293_,
		_w9294_
	);
	LUT2 #(
		.INIT('h4)
	) name5248 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001 ,
		_w9295_
	);
	LUT2 #(
		.INIT('h8)
	) name5249 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001 ,
		_w9296_
	);
	LUT2 #(
		.INIT('h1)
	) name5250 (
		_w9295_,
		_w9296_,
		_w9297_
	);
	LUT2 #(
		.INIT('h2)
	) name5251 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w9297_,
		_w9298_
	);
	LUT2 #(
		.INIT('h4)
	) name5252 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001 ,
		_w9299_
	);
	LUT2 #(
		.INIT('h8)
	) name5253 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001 ,
		_w9300_
	);
	LUT2 #(
		.INIT('h1)
	) name5254 (
		_w9299_,
		_w9300_,
		_w9301_
	);
	LUT2 #(
		.INIT('h2)
	) name5255 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w9301_,
		_w9302_
	);
	LUT2 #(
		.INIT('h4)
	) name5256 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001 ,
		_w9303_
	);
	LUT2 #(
		.INIT('h8)
	) name5257 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001 ,
		_w9304_
	);
	LUT2 #(
		.INIT('h1)
	) name5258 (
		_w9303_,
		_w9304_,
		_w9305_
	);
	LUT2 #(
		.INIT('h2)
	) name5259 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w9305_,
		_w9306_
	);
	LUT2 #(
		.INIT('h4)
	) name5260 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001 ,
		_w9307_
	);
	LUT2 #(
		.INIT('h8)
	) name5261 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001 ,
		_w9308_
	);
	LUT2 #(
		.INIT('h1)
	) name5262 (
		_w9307_,
		_w9308_,
		_w9309_
	);
	LUT2 #(
		.INIT('h2)
	) name5263 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w9309_,
		_w9310_
	);
	LUT2 #(
		.INIT('h4)
	) name5264 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001 ,
		_w9311_
	);
	LUT2 #(
		.INIT('h8)
	) name5265 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001 ,
		_w9312_
	);
	LUT2 #(
		.INIT('h1)
	) name5266 (
		_w9311_,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h2)
	) name5267 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w9313_,
		_w9314_
	);
	LUT2 #(
		.INIT('h8)
	) name5268 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w9315_
	);
	LUT2 #(
		.INIT('h1)
	) name5269 (
		_w9298_,
		_w9315_,
		_w9316_
	);
	LUT2 #(
		.INIT('h1)
	) name5270 (
		_w9302_,
		_w9306_,
		_w9317_
	);
	LUT2 #(
		.INIT('h1)
	) name5271 (
		_w9310_,
		_w9314_,
		_w9318_
	);
	LUT2 #(
		.INIT('h8)
	) name5272 (
		_w9317_,
		_w9318_,
		_w9319_
	);
	LUT2 #(
		.INIT('h8)
	) name5273 (
		_w9316_,
		_w9319_,
		_w9320_
	);
	LUT2 #(
		.INIT('h2)
	) name5274 (
		_w7093_,
		_w9320_,
		_w9321_
	);
	LUT2 #(
		.INIT('h8)
	) name5275 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w9322_
	);
	LUT2 #(
		.INIT('h8)
	) name5276 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w9323_
	);
	LUT2 #(
		.INIT('h8)
	) name5277 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		_w9324_
	);
	LUT2 #(
		.INIT('h8)
	) name5278 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w9325_
	);
	LUT2 #(
		.INIT('h8)
	) name5279 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131 ,
		_w9326_
	);
	LUT2 #(
		.INIT('h8)
	) name5280 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131 ,
		_w9327_
	);
	LUT2 #(
		.INIT('h8)
	) name5281 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131 ,
		_w9328_
	);
	LUT2 #(
		.INIT('h8)
	) name5282 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131 ,
		_w9329_
	);
	LUT2 #(
		.INIT('h8)
	) name5283 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131 ,
		_w9330_
	);
	LUT2 #(
		.INIT('h8)
	) name5284 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131 ,
		_w9331_
	);
	LUT2 #(
		.INIT('h8)
	) name5285 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131 ,
		_w9332_
	);
	LUT2 #(
		.INIT('h8)
	) name5286 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131 ,
		_w9333_
	);
	LUT2 #(
		.INIT('h1)
	) name5287 (
		_w9322_,
		_w9323_,
		_w9334_
	);
	LUT2 #(
		.INIT('h1)
	) name5288 (
		_w9324_,
		_w9325_,
		_w9335_
	);
	LUT2 #(
		.INIT('h1)
	) name5289 (
		_w9326_,
		_w9327_,
		_w9336_
	);
	LUT2 #(
		.INIT('h1)
	) name5290 (
		_w9328_,
		_w9329_,
		_w9337_
	);
	LUT2 #(
		.INIT('h1)
	) name5291 (
		_w9330_,
		_w9331_,
		_w9338_
	);
	LUT2 #(
		.INIT('h1)
	) name5292 (
		_w9332_,
		_w9333_,
		_w9339_
	);
	LUT2 #(
		.INIT('h8)
	) name5293 (
		_w9338_,
		_w9339_,
		_w9340_
	);
	LUT2 #(
		.INIT('h8)
	) name5294 (
		_w9336_,
		_w9337_,
		_w9341_
	);
	LUT2 #(
		.INIT('h8)
	) name5295 (
		_w9334_,
		_w9335_,
		_w9342_
	);
	LUT2 #(
		.INIT('h8)
	) name5296 (
		_w9341_,
		_w9342_,
		_w9343_
	);
	LUT2 #(
		.INIT('h8)
	) name5297 (
		_w9340_,
		_w9343_,
		_w9344_
	);
	LUT2 #(
		.INIT('h2)
	) name5298 (
		_w7128_,
		_w9344_,
		_w9345_
	);
	LUT2 #(
		.INIT('h8)
	) name5299 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w7249_,
		_w9346_
	);
	LUT2 #(
		.INIT('h8)
	) name5300 (
		\tm_tsr_reg_DO_reg[1]/NET0131 ,
		_w7540_,
		_w9347_
	);
	LUT2 #(
		.INIT('h8)
	) name5301 (
		\sport1_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w7263_,
		_w9348_
	);
	LUT2 #(
		.INIT('h8)
	) name5302 (
		\bdma_BWCOUNT_reg[1]/NET0131 ,
		_w7287_,
		_w9349_
	);
	LUT2 #(
		.INIT('h8)
	) name5303 (
		\emc_WSCRreg_DO_reg[1]/NET0131 ,
		_w7251_,
		_w9350_
	);
	LUT2 #(
		.INIT('h8)
	) name5304 (
		\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w7247_,
		_w9351_
	);
	LUT2 #(
		.INIT('h8)
	) name5305 (
		\idma_DOVL_reg[1]/NET0131 ,
		_w7532_,
		_w9352_
	);
	LUT2 #(
		.INIT('h8)
	) name5306 (
		\sport0_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w7295_,
		_w9353_
	);
	LUT2 #(
		.INIT('h8)
	) name5307 (
		\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w7256_,
		_w9354_
	);
	LUT2 #(
		.INIT('h8)
	) name5308 (
		\emc_WSCRext_reg_DO_reg[1]/NET0131 ,
		_w7514_,
		_w9355_
	);
	LUT2 #(
		.INIT('h8)
	) name5309 (
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w7259_,
		_w9356_
	);
	LUT2 #(
		.INIT('h8)
	) name5310 (
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w7527_,
		_w9357_
	);
	LUT2 #(
		.INIT('h8)
	) name5311 (
		\PIO_oe[1]_pad ,
		_w7244_,
		_w9358_
	);
	LUT2 #(
		.INIT('h8)
	) name5312 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w7234_,
		_w9359_
	);
	LUT2 #(
		.INIT('h8)
	) name5313 (
		\sport0_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w7276_,
		_w9360_
	);
	LUT2 #(
		.INIT('h8)
	) name5314 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w7299_,
		_w9361_
	);
	LUT2 #(
		.INIT('h8)
	) name5315 (
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w7273_,
		_w9362_
	);
	LUT2 #(
		.INIT('h8)
	) name5316 (
		\memc_usysr_DO_reg[1]/NET0131 ,
		_w7301_,
		_w9363_
	);
	LUT2 #(
		.INIT('h8)
	) name5317 (
		\bdma_BOVL_reg[1]/NET0131 ,
		_w7534_,
		_w9364_
	);
	LUT2 #(
		.INIT('h8)
	) name5318 (
		\tm_tpr_reg_DO_reg[1]/NET0131 ,
		_w7293_,
		_w9365_
	);
	LUT2 #(
		.INIT('h8)
	) name5319 (
		\clkc_ckr_reg_DO_reg[1]/NET0131 ,
		_w7239_,
		_w9366_
	);
	LUT2 #(
		.INIT('h8)
	) name5320 (
		\bdma_BEAD_reg[1]/NET0131 ,
		_w7303_,
		_w9367_
	);
	LUT2 #(
		.INIT('h8)
	) name5321 (
		\bdma_BCTL_reg[1]/NET0131 ,
		_w7230_,
		_w9368_
	);
	LUT2 #(
		.INIT('h8)
	) name5322 (
		\pio_PINT_reg[1]/NET0131 ,
		_w7271_,
		_w9369_
	);
	LUT2 #(
		.INIT('h8)
	) name5323 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w7281_,
		_w9370_
	);
	LUT2 #(
		.INIT('h8)
	) name5324 (
		\pio_pmask_reg_DO_reg[1]/NET0131 ,
		_w7297_,
		_w9371_
	);
	LUT2 #(
		.INIT('h8)
	) name5325 (
		\PIO_out[1]_pad ,
		_w7291_,
		_w9372_
	);
	LUT2 #(
		.INIT('h8)
	) name5326 (
		\tm_TCR_TMP_reg[1]/NET0131 ,
		_w7289_,
		_w9373_
	);
	LUT2 #(
		.INIT('h1)
	) name5327 (
		_w7522_,
		_w9346_,
		_w9374_
	);
	LUT2 #(
		.INIT('h1)
	) name5328 (
		_w9347_,
		_w9348_,
		_w9375_
	);
	LUT2 #(
		.INIT('h1)
	) name5329 (
		_w9350_,
		_w9351_,
		_w9376_
	);
	LUT2 #(
		.INIT('h1)
	) name5330 (
		_w9352_,
		_w9353_,
		_w9377_
	);
	LUT2 #(
		.INIT('h1)
	) name5331 (
		_w9354_,
		_w9355_,
		_w9378_
	);
	LUT2 #(
		.INIT('h1)
	) name5332 (
		_w9356_,
		_w9357_,
		_w9379_
	);
	LUT2 #(
		.INIT('h1)
	) name5333 (
		_w9358_,
		_w9360_,
		_w9380_
	);
	LUT2 #(
		.INIT('h1)
	) name5334 (
		_w9361_,
		_w9362_,
		_w9381_
	);
	LUT2 #(
		.INIT('h1)
	) name5335 (
		_w9363_,
		_w9365_,
		_w9382_
	);
	LUT2 #(
		.INIT('h1)
	) name5336 (
		_w9366_,
		_w9369_,
		_w9383_
	);
	LUT2 #(
		.INIT('h1)
	) name5337 (
		_w9370_,
		_w9371_,
		_w9384_
	);
	LUT2 #(
		.INIT('h1)
	) name5338 (
		_w9372_,
		_w9373_,
		_w9385_
	);
	LUT2 #(
		.INIT('h8)
	) name5339 (
		_w9384_,
		_w9385_,
		_w9386_
	);
	LUT2 #(
		.INIT('h8)
	) name5340 (
		_w9382_,
		_w9383_,
		_w9387_
	);
	LUT2 #(
		.INIT('h8)
	) name5341 (
		_w9380_,
		_w9381_,
		_w9388_
	);
	LUT2 #(
		.INIT('h8)
	) name5342 (
		_w9378_,
		_w9379_,
		_w9389_
	);
	LUT2 #(
		.INIT('h8)
	) name5343 (
		_w9376_,
		_w9377_,
		_w9390_
	);
	LUT2 #(
		.INIT('h8)
	) name5344 (
		_w9374_,
		_w9375_,
		_w9391_
	);
	LUT2 #(
		.INIT('h8)
	) name5345 (
		_w9390_,
		_w9391_,
		_w9392_
	);
	LUT2 #(
		.INIT('h8)
	) name5346 (
		_w9388_,
		_w9389_,
		_w9393_
	);
	LUT2 #(
		.INIT('h8)
	) name5347 (
		_w9386_,
		_w9387_,
		_w9394_
	);
	LUT2 #(
		.INIT('h8)
	) name5348 (
		_w9393_,
		_w9394_,
		_w9395_
	);
	LUT2 #(
		.INIT('h4)
	) name5349 (
		_w9359_,
		_w9392_,
		_w9396_
	);
	LUT2 #(
		.INIT('h1)
	) name5350 (
		_w9367_,
		_w9368_,
		_w9397_
	);
	LUT2 #(
		.INIT('h8)
	) name5351 (
		_w9396_,
		_w9397_,
		_w9398_
	);
	LUT2 #(
		.INIT('h4)
	) name5352 (
		_w9349_,
		_w9395_,
		_w9399_
	);
	LUT2 #(
		.INIT('h4)
	) name5353 (
		_w9364_,
		_w9399_,
		_w9400_
	);
	LUT2 #(
		.INIT('h8)
	) name5354 (
		_w9398_,
		_w9400_,
		_w9401_
	);
	LUT2 #(
		.INIT('h2)
	) name5355 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w9401_,
		_w9402_
	);
	LUT2 #(
		.INIT('h8)
	) name5356 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		_w9403_
	);
	LUT2 #(
		.INIT('h8)
	) name5357 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w9404_
	);
	LUT2 #(
		.INIT('h8)
	) name5358 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w9405_
	);
	LUT2 #(
		.INIT('h2)
	) name5359 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4457_,
		_w9406_
	);
	LUT2 #(
		.INIT('h2)
	) name5360 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w7216_,
		_w9407_
	);
	LUT2 #(
		.INIT('h8)
	) name5361 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w9408_
	);
	LUT2 #(
		.INIT('h8)
	) name5362 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w9409_
	);
	LUT2 #(
		.INIT('h8)
	) name5363 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[1]/NET0131 ,
		_w9410_
	);
	LUT2 #(
		.INIT('h8)
	) name5364 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w9411_
	);
	LUT2 #(
		.INIT('h8)
	) name5365 (
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\core_c_psq_ICNTL_reg_DO_reg[1]/NET0131 ,
		_w9412_
	);
	LUT2 #(
		.INIT('h1)
	) name5366 (
		_w9403_,
		_w9404_,
		_w9413_
	);
	LUT2 #(
		.INIT('h1)
	) name5367 (
		_w9405_,
		_w9408_,
		_w9414_
	);
	LUT2 #(
		.INIT('h1)
	) name5368 (
		_w9409_,
		_w9410_,
		_w9415_
	);
	LUT2 #(
		.INIT('h1)
	) name5369 (
		_w9411_,
		_w9412_,
		_w9416_
	);
	LUT2 #(
		.INIT('h8)
	) name5370 (
		_w9415_,
		_w9416_,
		_w9417_
	);
	LUT2 #(
		.INIT('h8)
	) name5371 (
		_w9413_,
		_w9414_,
		_w9418_
	);
	LUT2 #(
		.INIT('h4)
	) name5372 (
		_w9407_,
		_w9418_,
		_w9419_
	);
	LUT2 #(
		.INIT('h8)
	) name5373 (
		_w9417_,
		_w9419_,
		_w9420_
	);
	LUT2 #(
		.INIT('h4)
	) name5374 (
		_w9406_,
		_w9420_,
		_w9421_
	);
	LUT2 #(
		.INIT('h2)
	) name5375 (
		_w7215_,
		_w9421_,
		_w9422_
	);
	LUT2 #(
		.INIT('h1)
	) name5376 (
		_w9261_,
		_w9294_,
		_w9423_
	);
	LUT2 #(
		.INIT('h4)
	) name5377 (
		_w9345_,
		_w9423_,
		_w9424_
	);
	LUT2 #(
		.INIT('h1)
	) name5378 (
		_w9237_,
		_w9286_,
		_w9425_
	);
	LUT2 #(
		.INIT('h4)
	) name5379 (
		_w9321_,
		_w9425_,
		_w9426_
	);
	LUT2 #(
		.INIT('h8)
	) name5380 (
		_w9424_,
		_w9426_,
		_w9427_
	);
	LUT2 #(
		.INIT('h4)
	) name5381 (
		_w9422_,
		_w9427_,
		_w9428_
	);
	LUT2 #(
		.INIT('h4)
	) name5382 (
		_w9402_,
		_w9428_,
		_w9429_
	);
	LUT2 #(
		.INIT('h4)
	) name5383 (
		_w9202_,
		_w9429_,
		_w9430_
	);
	LUT2 #(
		.INIT('h1)
	) name5384 (
		\emc_DMDoe_reg/NET0131 ,
		_w9430_,
		_w9431_
	);
	LUT2 #(
		.INIT('h8)
	) name5385 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[1]/P0001 ,
		_w9432_
	);
	LUT2 #(
		.INIT('h2)
	) name5386 (
		_w7057_,
		_w9432_,
		_w9433_
	);
	LUT2 #(
		.INIT('h4)
	) name5387 (
		_w9431_,
		_w9433_,
		_w9434_
	);
	LUT2 #(
		.INIT('h1)
	) name5388 (
		_w9201_,
		_w9434_,
		_w9435_
	);
	LUT2 #(
		.INIT('h8)
	) name5389 (
		_w7863_,
		_w9435_,
		_w9436_
	);
	LUT2 #(
		.INIT('h1)
	) name5390 (
		_w9183_,
		_w9436_,
		_w9437_
	);
	LUT2 #(
		.INIT('h2)
	) name5391 (
		_w7005_,
		_w9437_,
		_w9438_
	);
	LUT2 #(
		.INIT('h1)
	) name5392 (
		_w9181_,
		_w9438_,
		_w9439_
	);
	LUT2 #(
		.INIT('h4)
	) name5393 (
		_w8950_,
		_w9439_,
		_w9440_
	);
	LUT2 #(
		.INIT('h1)
	) name5394 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w6924_,
		_w9441_
	);
	LUT2 #(
		.INIT('h8)
	) name5395 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131 ,
		_w6988_,
		_w9442_
	);
	LUT2 #(
		.INIT('h8)
	) name5396 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w6926_,
		_w9443_
	);
	LUT2 #(
		.INIT('h4)
	) name5397 (
		_w6111_,
		_w6160_,
		_w9444_
	);
	LUT2 #(
		.INIT('h8)
	) name5398 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w6956_,
		_w9445_
	);
	LUT2 #(
		.INIT('h8)
	) name5399 (
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w6976_,
		_w9446_
	);
	LUT2 #(
		.INIT('h8)
	) name5400 (
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		_w6970_,
		_w9447_
	);
	LUT2 #(
		.INIT('h8)
	) name5401 (
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w6974_,
		_w9448_
	);
	LUT2 #(
		.INIT('h8)
	) name5402 (
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w6972_,
		_w9449_
	);
	LUT2 #(
		.INIT('h1)
	) name5403 (
		_w9446_,
		_w9447_,
		_w9450_
	);
	LUT2 #(
		.INIT('h1)
	) name5404 (
		_w9448_,
		_w9449_,
		_w9451_
	);
	LUT2 #(
		.INIT('h8)
	) name5405 (
		_w9450_,
		_w9451_,
		_w9452_
	);
	LUT2 #(
		.INIT('h2)
	) name5406 (
		_w4055_,
		_w9452_,
		_w9453_
	);
	LUT2 #(
		.INIT('h8)
	) name5407 (
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w6960_,
		_w9454_
	);
	LUT2 #(
		.INIT('h8)
	) name5408 (
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w6958_,
		_w9455_
	);
	LUT2 #(
		.INIT('h8)
	) name5409 (
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w6962_,
		_w9456_
	);
	LUT2 #(
		.INIT('h8)
	) name5410 (
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		_w6964_,
		_w9457_
	);
	LUT2 #(
		.INIT('h1)
	) name5411 (
		_w9454_,
		_w9455_,
		_w9458_
	);
	LUT2 #(
		.INIT('h1)
	) name5412 (
		_w9456_,
		_w9457_,
		_w9459_
	);
	LUT2 #(
		.INIT('h8)
	) name5413 (
		_w9458_,
		_w9459_,
		_w9460_
	);
	LUT2 #(
		.INIT('h4)
	) name5414 (
		_w9453_,
		_w9460_,
		_w9461_
	);
	LUT2 #(
		.INIT('h1)
	) name5415 (
		_w6121_,
		_w9461_,
		_w9462_
	);
	LUT2 #(
		.INIT('h1)
	) name5416 (
		_w9444_,
		_w9445_,
		_w9463_
	);
	LUT2 #(
		.INIT('h4)
	) name5417 (
		_w9462_,
		_w9463_,
		_w9464_
	);
	LUT2 #(
		.INIT('h2)
	) name5418 (
		_w5949_,
		_w9464_,
		_w9465_
	);
	LUT2 #(
		.INIT('h2)
	) name5419 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		_w6934_,
		_w9466_
	);
	LUT2 #(
		.INIT('h1)
	) name5420 (
		_w9442_,
		_w9443_,
		_w9467_
	);
	LUT2 #(
		.INIT('h8)
	) name5421 (
		_w6924_,
		_w9467_,
		_w9468_
	);
	LUT2 #(
		.INIT('h4)
	) name5422 (
		_w9466_,
		_w9468_,
		_w9469_
	);
	LUT2 #(
		.INIT('h4)
	) name5423 (
		_w9465_,
		_w9469_,
		_w9470_
	);
	LUT2 #(
		.INIT('h1)
	) name5424 (
		_w6176_,
		_w9441_,
		_w9471_
	);
	LUT2 #(
		.INIT('h4)
	) name5425 (
		_w9470_,
		_w9471_,
		_w9472_
	);
	LUT2 #(
		.INIT('h8)
	) name5426 (
		_w6176_,
		_w6953_,
		_w9473_
	);
	LUT2 #(
		.INIT('h1)
	) name5427 (
		_w6135_,
		_w9473_,
		_w9474_
	);
	LUT2 #(
		.INIT('h4)
	) name5428 (
		_w9472_,
		_w9474_,
		_w9475_
	);
	LUT2 #(
		.INIT('h2)
	) name5429 (
		_w6176_,
		_w7622_,
		_w9476_
	);
	LUT2 #(
		.INIT('h1)
	) name5430 (
		_w6888_,
		_w6898_,
		_w9477_
	);
	LUT2 #(
		.INIT('h1)
	) name5431 (
		_w6880_,
		_w6895_,
		_w9478_
	);
	LUT2 #(
		.INIT('h1)
	) name5432 (
		_w6899_,
		_w9478_,
		_w9479_
	);
	LUT2 #(
		.INIT('h2)
	) name5433 (
		_w9477_,
		_w9479_,
		_w9480_
	);
	LUT2 #(
		.INIT('h4)
	) name5434 (
		_w9477_,
		_w9479_,
		_w9481_
	);
	LUT2 #(
		.INIT('h1)
	) name5435 (
		_w9480_,
		_w9481_,
		_w9482_
	);
	LUT2 #(
		.INIT('h2)
	) name5436 (
		_w6717_,
		_w9482_,
		_w9483_
	);
	LUT2 #(
		.INIT('h1)
	) name5437 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w6605_,
		_w9484_
	);
	LUT2 #(
		.INIT('h1)
	) name5438 (
		_w6606_,
		_w9484_,
		_w9485_
	);
	LUT2 #(
		.INIT('h4)
	) name5439 (
		_w6712_,
		_w9485_,
		_w9486_
	);
	LUT2 #(
		.INIT('h2)
	) name5440 (
		_w6712_,
		_w9485_,
		_w9487_
	);
	LUT2 #(
		.INIT('h1)
	) name5441 (
		_w9486_,
		_w9487_,
		_w9488_
	);
	LUT2 #(
		.INIT('h8)
	) name5442 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w9488_,
		_w9489_
	);
	LUT2 #(
		.INIT('h4)
	) name5443 (
		_w9483_,
		_w9489_,
		_w9490_
	);
	LUT2 #(
		.INIT('h1)
	) name5444 (
		_w6905_,
		_w9488_,
		_w9491_
	);
	LUT2 #(
		.INIT('h2)
	) name5445 (
		_w6905_,
		_w9482_,
		_w9492_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w9492_,
		_w9493_
	);
	LUT2 #(
		.INIT('h4)
	) name5447 (
		_w9491_,
		_w9493_,
		_w9494_
	);
	LUT2 #(
		.INIT('h8)
	) name5448 (
		\core_dag_ilm2reg_I_reg[13]/NET0131 ,
		_w6604_,
		_w9495_
	);
	LUT2 #(
		.INIT('h1)
	) name5449 (
		_w9494_,
		_w9495_,
		_w9496_
	);
	LUT2 #(
		.INIT('h4)
	) name5450 (
		_w9490_,
		_w9496_,
		_w9497_
	);
	LUT2 #(
		.INIT('h1)
	) name5451 (
		_w6176_,
		_w9497_,
		_w9498_
	);
	LUT2 #(
		.INIT('h2)
	) name5452 (
		_w6135_,
		_w9476_,
		_w9499_
	);
	LUT2 #(
		.INIT('h4)
	) name5453 (
		_w9498_,
		_w9499_,
		_w9500_
	);
	LUT2 #(
		.INIT('h1)
	) name5454 (
		_w7005_,
		_w9475_,
		_w9501_
	);
	LUT2 #(
		.INIT('h4)
	) name5455 (
		_w9500_,
		_w9501_,
		_w9502_
	);
	LUT2 #(
		.INIT('h4)
	) name5456 (
		_w6160_,
		_w9461_,
		_w9503_
	);
	LUT2 #(
		.INIT('h2)
	) name5457 (
		_w8153_,
		_w9503_,
		_w9504_
	);
	LUT2 #(
		.INIT('h8)
	) name5458 (
		_w7607_,
		_w7863_,
		_w9505_
	);
	LUT2 #(
		.INIT('h1)
	) name5459 (
		_w9504_,
		_w9505_,
		_w9506_
	);
	LUT2 #(
		.INIT('h2)
	) name5460 (
		_w7005_,
		_w9506_,
		_w9507_
	);
	LUT2 #(
		.INIT('h4)
	) name5461 (
		_w6135_,
		_w6546_,
		_w9508_
	);
	LUT2 #(
		.INIT('h2)
	) name5462 (
		_w6135_,
		_w7340_,
		_w9509_
	);
	LUT2 #(
		.INIT('h2)
	) name5463 (
		_w8964_,
		_w9509_,
		_w9510_
	);
	LUT2 #(
		.INIT('h4)
	) name5464 (
		_w9508_,
		_w9510_,
		_w9511_
	);
	LUT2 #(
		.INIT('h1)
	) name5465 (
		_w9507_,
		_w9511_,
		_w9512_
	);
	LUT2 #(
		.INIT('h4)
	) name5466 (
		_w9502_,
		_w9512_,
		_w9513_
	);
	LUT2 #(
		.INIT('h8)
	) name5467 (
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		_w6964_,
		_w9514_
	);
	LUT2 #(
		.INIT('h8)
	) name5468 (
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w6960_,
		_w9515_
	);
	LUT2 #(
		.INIT('h8)
	) name5469 (
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w6962_,
		_w9516_
	);
	LUT2 #(
		.INIT('h8)
	) name5470 (
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w6958_,
		_w9517_
	);
	LUT2 #(
		.INIT('h1)
	) name5471 (
		_w9514_,
		_w9515_,
		_w9518_
	);
	LUT2 #(
		.INIT('h1)
	) name5472 (
		_w9516_,
		_w9517_,
		_w9519_
	);
	LUT2 #(
		.INIT('h8)
	) name5473 (
		_w9518_,
		_w9519_,
		_w9520_
	);
	LUT2 #(
		.INIT('h4)
	) name5474 (
		_w4055_,
		_w9520_,
		_w9521_
	);
	LUT2 #(
		.INIT('h8)
	) name5475 (
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w6976_,
		_w9522_
	);
	LUT2 #(
		.INIT('h8)
	) name5476 (
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		_w6970_,
		_w9523_
	);
	LUT2 #(
		.INIT('h8)
	) name5477 (
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w6974_,
		_w9524_
	);
	LUT2 #(
		.INIT('h8)
	) name5478 (
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w6972_,
		_w9525_
	);
	LUT2 #(
		.INIT('h1)
	) name5479 (
		_w9522_,
		_w9523_,
		_w9526_
	);
	LUT2 #(
		.INIT('h1)
	) name5480 (
		_w9524_,
		_w9525_,
		_w9527_
	);
	LUT2 #(
		.INIT('h8)
	) name5481 (
		_w9526_,
		_w9527_,
		_w9528_
	);
	LUT2 #(
		.INIT('h8)
	) name5482 (
		_w4055_,
		_w9528_,
		_w9529_
	);
	LUT2 #(
		.INIT('h1)
	) name5483 (
		_w9521_,
		_w9529_,
		_w9530_
	);
	LUT2 #(
		.INIT('h1)
	) name5484 (
		_w8905_,
		_w9530_,
		_w9531_
	);
	LUT2 #(
		.INIT('h8)
	) name5485 (
		_w6135_,
		_w9531_,
		_w9532_
	);
	LUT2 #(
		.INIT('h1)
	) name5486 (
		_w6135_,
		_w9178_,
		_w9533_
	);
	LUT2 #(
		.INIT('h1)
	) name5487 (
		_w6176_,
		_w9532_,
		_w9534_
	);
	LUT2 #(
		.INIT('h4)
	) name5488 (
		_w9533_,
		_w9534_,
		_w9535_
	);
	LUT2 #(
		.INIT('h4)
	) name5489 (
		_w6135_,
		_w8926_,
		_w9536_
	);
	LUT2 #(
		.INIT('h2)
	) name5490 (
		_w6135_,
		_w9435_,
		_w9537_
	);
	LUT2 #(
		.INIT('h2)
	) name5491 (
		_w6176_,
		_w9537_,
		_w9538_
	);
	LUT2 #(
		.INIT('h4)
	) name5492 (
		_w9536_,
		_w9538_,
		_w9539_
	);
	LUT2 #(
		.INIT('h1)
	) name5493 (
		_w9535_,
		_w9539_,
		_w9540_
	);
	LUT2 #(
		.INIT('h2)
	) name5494 (
		_w7005_,
		_w9540_,
		_w9541_
	);
	LUT2 #(
		.INIT('h8)
	) name5495 (
		\core_dag_ilm2reg_I_reg[1]/NET0131 ,
		_w6664_,
		_w9542_
	);
	LUT2 #(
		.INIT('h1)
	) name5496 (
		_w6811_,
		_w6812_,
		_w9543_
	);
	LUT2 #(
		.INIT('h2)
	) name5497 (
		_w6713_,
		_w9543_,
		_w9544_
	);
	LUT2 #(
		.INIT('h2)
	) name5498 (
		_w6596_,
		_w6807_,
		_w9545_
	);
	LUT2 #(
		.INIT('h4)
	) name5499 (
		_w6596_,
		_w6807_,
		_w9546_
	);
	LUT2 #(
		.INIT('h1)
	) name5500 (
		_w9545_,
		_w9546_,
		_w9547_
	);
	LUT2 #(
		.INIT('h4)
	) name5501 (
		_w6717_,
		_w9547_,
		_w9548_
	);
	LUT2 #(
		.INIT('h2)
	) name5502 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w9544_,
		_w9549_
	);
	LUT2 #(
		.INIT('h4)
	) name5503 (
		_w9548_,
		_w9549_,
		_w9550_
	);
	LUT2 #(
		.INIT('h2)
	) name5504 (
		_w6724_,
		_w9543_,
		_w9551_
	);
	LUT2 #(
		.INIT('h4)
	) name5505 (
		_w6724_,
		_w9543_,
		_w9552_
	);
	LUT2 #(
		.INIT('h1)
	) name5506 (
		_w9551_,
		_w9552_,
		_w9553_
	);
	LUT2 #(
		.INIT('h8)
	) name5507 (
		_w6905_,
		_w9553_,
		_w9554_
	);
	LUT2 #(
		.INIT('h4)
	) name5508 (
		_w6905_,
		_w9547_,
		_w9555_
	);
	LUT2 #(
		.INIT('h1)
	) name5509 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w9554_,
		_w9556_
	);
	LUT2 #(
		.INIT('h4)
	) name5510 (
		_w9555_,
		_w9556_,
		_w9557_
	);
	LUT2 #(
		.INIT('h1)
	) name5511 (
		_w9542_,
		_w9557_,
		_w9558_
	);
	LUT2 #(
		.INIT('h4)
	) name5512 (
		_w9550_,
		_w9558_,
		_w9559_
	);
	LUT2 #(
		.INIT('h2)
	) name5513 (
		_w6135_,
		_w9559_,
		_w9560_
	);
	LUT2 #(
		.INIT('h1)
	) name5514 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w6924_,
		_w9561_
	);
	LUT2 #(
		.INIT('h2)
	) name5515 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w6934_,
		_w9562_
	);
	LUT2 #(
		.INIT('h8)
	) name5516 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w6926_,
		_w9563_
	);
	LUT2 #(
		.INIT('h8)
	) name5517 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[1]/NET0131 ,
		_w6988_,
		_w9564_
	);
	LUT2 #(
		.INIT('h4)
	) name5518 (
		_w6111_,
		_w8905_,
		_w9565_
	);
	LUT2 #(
		.INIT('h4)
	) name5519 (
		_w6121_,
		_w9530_,
		_w9566_
	);
	LUT2 #(
		.INIT('h8)
	) name5520 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w6956_,
		_w9567_
	);
	LUT2 #(
		.INIT('h1)
	) name5521 (
		_w9565_,
		_w9567_,
		_w9568_
	);
	LUT2 #(
		.INIT('h4)
	) name5522 (
		_w9566_,
		_w9568_,
		_w9569_
	);
	LUT2 #(
		.INIT('h2)
	) name5523 (
		_w5949_,
		_w9569_,
		_w9570_
	);
	LUT2 #(
		.INIT('h1)
	) name5524 (
		_w9563_,
		_w9564_,
		_w9571_
	);
	LUT2 #(
		.INIT('h8)
	) name5525 (
		_w6924_,
		_w9571_,
		_w9572_
	);
	LUT2 #(
		.INIT('h4)
	) name5526 (
		_w9562_,
		_w9572_,
		_w9573_
	);
	LUT2 #(
		.INIT('h4)
	) name5527 (
		_w9570_,
		_w9573_,
		_w9574_
	);
	LUT2 #(
		.INIT('h1)
	) name5528 (
		_w6135_,
		_w9561_,
		_w9575_
	);
	LUT2 #(
		.INIT('h4)
	) name5529 (
		_w9574_,
		_w9575_,
		_w9576_
	);
	LUT2 #(
		.INIT('h1)
	) name5530 (
		_w9560_,
		_w9576_,
		_w9577_
	);
	LUT2 #(
		.INIT('h1)
	) name5531 (
		_w6176_,
		_w9577_,
		_w9578_
	);
	LUT2 #(
		.INIT('h1)
	) name5532 (
		_w6135_,
		_w8875_,
		_w9579_
	);
	LUT2 #(
		.INIT('h8)
	) name5533 (
		_w6135_,
		_w8962_,
		_w9580_
	);
	LUT2 #(
		.INIT('h2)
	) name5534 (
		_w6176_,
		_w9579_,
		_w9581_
	);
	LUT2 #(
		.INIT('h4)
	) name5535 (
		_w9580_,
		_w9581_,
		_w9582_
	);
	LUT2 #(
		.INIT('h1)
	) name5536 (
		_w9578_,
		_w9582_,
		_w9583_
	);
	LUT2 #(
		.INIT('h1)
	) name5537 (
		_w7005_,
		_w9583_,
		_w9584_
	);
	LUT2 #(
		.INIT('h1)
	) name5538 (
		_w9541_,
		_w9584_,
		_w9585_
	);
	LUT2 #(
		.INIT('h8)
	) name5539 (
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w6960_,
		_w9586_
	);
	LUT2 #(
		.INIT('h8)
	) name5540 (
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w6958_,
		_w9587_
	);
	LUT2 #(
		.INIT('h8)
	) name5541 (
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w6962_,
		_w9588_
	);
	LUT2 #(
		.INIT('h8)
	) name5542 (
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		_w6964_,
		_w9589_
	);
	LUT2 #(
		.INIT('h1)
	) name5543 (
		_w9586_,
		_w9587_,
		_w9590_
	);
	LUT2 #(
		.INIT('h1)
	) name5544 (
		_w9588_,
		_w9589_,
		_w9591_
	);
	LUT2 #(
		.INIT('h8)
	) name5545 (
		_w9590_,
		_w9591_,
		_w9592_
	);
	LUT2 #(
		.INIT('h4)
	) name5546 (
		_w4055_,
		_w9592_,
		_w9593_
	);
	LUT2 #(
		.INIT('h8)
	) name5547 (
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w6972_,
		_w9594_
	);
	LUT2 #(
		.INIT('h8)
	) name5548 (
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w6976_,
		_w9595_
	);
	LUT2 #(
		.INIT('h8)
	) name5549 (
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w6974_,
		_w9596_
	);
	LUT2 #(
		.INIT('h8)
	) name5550 (
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		_w6970_,
		_w9597_
	);
	LUT2 #(
		.INIT('h1)
	) name5551 (
		_w9594_,
		_w9595_,
		_w9598_
	);
	LUT2 #(
		.INIT('h1)
	) name5552 (
		_w9596_,
		_w9597_,
		_w9599_
	);
	LUT2 #(
		.INIT('h8)
	) name5553 (
		_w9598_,
		_w9599_,
		_w9600_
	);
	LUT2 #(
		.INIT('h8)
	) name5554 (
		_w4055_,
		_w9600_,
		_w9601_
	);
	LUT2 #(
		.INIT('h1)
	) name5555 (
		_w9593_,
		_w9601_,
		_w9602_
	);
	LUT2 #(
		.INIT('h1)
	) name5556 (
		_w8775_,
		_w9602_,
		_w9603_
	);
	LUT2 #(
		.INIT('h8)
	) name5557 (
		_w6135_,
		_w9603_,
		_w9604_
	);
	LUT2 #(
		.INIT('h1)
	) name5558 (
		_w6135_,
		_w8460_,
		_w9605_
	);
	LUT2 #(
		.INIT('h1)
	) name5559 (
		_w6176_,
		_w9604_,
		_w9606_
	);
	LUT2 #(
		.INIT('h4)
	) name5560 (
		_w9605_,
		_w9606_,
		_w9607_
	);
	LUT2 #(
		.INIT('h4)
	) name5561 (
		_w6135_,
		_w8794_,
		_w9608_
	);
	LUT2 #(
		.INIT('h2)
	) name5562 (
		_w6135_,
		_w8715_,
		_w9609_
	);
	LUT2 #(
		.INIT('h2)
	) name5563 (
		_w6176_,
		_w9609_,
		_w9610_
	);
	LUT2 #(
		.INIT('h4)
	) name5564 (
		_w9608_,
		_w9610_,
		_w9611_
	);
	LUT2 #(
		.INIT('h1)
	) name5565 (
		_w9607_,
		_w9611_,
		_w9612_
	);
	LUT2 #(
		.INIT('h2)
	) name5566 (
		_w7005_,
		_w9612_,
		_w9613_
	);
	LUT2 #(
		.INIT('h2)
	) name5567 (
		\core_dag_ilm2reg_I_reg[2]/NET0131 ,
		_w6660_,
		_w9614_
	);
	LUT2 #(
		.INIT('h1)
	) name5568 (
		_w6803_,
		_w6804_,
		_w9615_
	);
	LUT2 #(
		.INIT('h1)
	) name5569 (
		_w6815_,
		_w9615_,
		_w9616_
	);
	LUT2 #(
		.INIT('h8)
	) name5570 (
		_w6815_,
		_w9615_,
		_w9617_
	);
	LUT2 #(
		.INIT('h1)
	) name5571 (
		_w9616_,
		_w9617_,
		_w9618_
	);
	LUT2 #(
		.INIT('h8)
	) name5572 (
		_w8198_,
		_w9618_,
		_w9619_
	);
	LUT2 #(
		.INIT('h1)
	) name5573 (
		_w6671_,
		_w6799_,
		_w9620_
	);
	LUT2 #(
		.INIT('h8)
	) name5574 (
		_w6671_,
		_w6799_,
		_w9621_
	);
	LUT2 #(
		.INIT('h1)
	) name5575 (
		_w9620_,
		_w9621_,
		_w9622_
	);
	LUT2 #(
		.INIT('h4)
	) name5576 (
		_w8198_,
		_w9622_,
		_w9623_
	);
	LUT2 #(
		.INIT('h1)
	) name5577 (
		_w9614_,
		_w9619_,
		_w9624_
	);
	LUT2 #(
		.INIT('h4)
	) name5578 (
		_w9623_,
		_w9624_,
		_w9625_
	);
	LUT2 #(
		.INIT('h2)
	) name5579 (
		_w6135_,
		_w9625_,
		_w9626_
	);
	LUT2 #(
		.INIT('h1)
	) name5580 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w6924_,
		_w9627_
	);
	LUT2 #(
		.INIT('h2)
	) name5581 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		_w6934_,
		_w9628_
	);
	LUT2 #(
		.INIT('h8)
	) name5582 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w6926_,
		_w9629_
	);
	LUT2 #(
		.INIT('h8)
	) name5583 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[2]/NET0131 ,
		_w6988_,
		_w9630_
	);
	LUT2 #(
		.INIT('h4)
	) name5584 (
		_w6111_,
		_w8775_,
		_w9631_
	);
	LUT2 #(
		.INIT('h4)
	) name5585 (
		_w6121_,
		_w9602_,
		_w9632_
	);
	LUT2 #(
		.INIT('h8)
	) name5586 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w6956_,
		_w9633_
	);
	LUT2 #(
		.INIT('h1)
	) name5587 (
		_w9631_,
		_w9633_,
		_w9634_
	);
	LUT2 #(
		.INIT('h4)
	) name5588 (
		_w9632_,
		_w9634_,
		_w9635_
	);
	LUT2 #(
		.INIT('h2)
	) name5589 (
		_w5949_,
		_w9635_,
		_w9636_
	);
	LUT2 #(
		.INIT('h1)
	) name5590 (
		_w9629_,
		_w9630_,
		_w9637_
	);
	LUT2 #(
		.INIT('h8)
	) name5591 (
		_w6924_,
		_w9637_,
		_w9638_
	);
	LUT2 #(
		.INIT('h4)
	) name5592 (
		_w9628_,
		_w9638_,
		_w9639_
	);
	LUT2 #(
		.INIT('h4)
	) name5593 (
		_w9636_,
		_w9639_,
		_w9640_
	);
	LUT2 #(
		.INIT('h1)
	) name5594 (
		_w6135_,
		_w9627_,
		_w9641_
	);
	LUT2 #(
		.INIT('h4)
	) name5595 (
		_w9640_,
		_w9641_,
		_w9642_
	);
	LUT2 #(
		.INIT('h1)
	) name5596 (
		_w9626_,
		_w9642_,
		_w9643_
	);
	LUT2 #(
		.INIT('h1)
	) name5597 (
		_w6176_,
		_w9643_,
		_w9644_
	);
	LUT2 #(
		.INIT('h8)
	) name5598 (
		_w6135_,
		_w8246_,
		_w9645_
	);
	LUT2 #(
		.INIT('h1)
	) name5599 (
		_w6135_,
		_w8752_,
		_w9646_
	);
	LUT2 #(
		.INIT('h2)
	) name5600 (
		_w6176_,
		_w9646_,
		_w9647_
	);
	LUT2 #(
		.INIT('h4)
	) name5601 (
		_w9645_,
		_w9647_,
		_w9648_
	);
	LUT2 #(
		.INIT('h1)
	) name5602 (
		_w9644_,
		_w9648_,
		_w9649_
	);
	LUT2 #(
		.INIT('h1)
	) name5603 (
		_w7005_,
		_w9649_,
		_w9650_
	);
	LUT2 #(
		.INIT('h1)
	) name5604 (
		_w9613_,
		_w9650_,
		_w9651_
	);
	LUT2 #(
		.INIT('h8)
	) name5605 (
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w6958_,
		_w9652_
	);
	LUT2 #(
		.INIT('h8)
	) name5606 (
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w6960_,
		_w9653_
	);
	LUT2 #(
		.INIT('h8)
	) name5607 (
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w6962_,
		_w9654_
	);
	LUT2 #(
		.INIT('h8)
	) name5608 (
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		_w6964_,
		_w9655_
	);
	LUT2 #(
		.INIT('h1)
	) name5609 (
		_w9652_,
		_w9653_,
		_w9656_
	);
	LUT2 #(
		.INIT('h1)
	) name5610 (
		_w9654_,
		_w9655_,
		_w9657_
	);
	LUT2 #(
		.INIT('h8)
	) name5611 (
		_w9656_,
		_w9657_,
		_w9658_
	);
	LUT2 #(
		.INIT('h4)
	) name5612 (
		_w4055_,
		_w9658_,
		_w9659_
	);
	LUT2 #(
		.INIT('h8)
	) name5613 (
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w6976_,
		_w9660_
	);
	LUT2 #(
		.INIT('h8)
	) name5614 (
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		_w6970_,
		_w9661_
	);
	LUT2 #(
		.INIT('h8)
	) name5615 (
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w6974_,
		_w9662_
	);
	LUT2 #(
		.INIT('h8)
	) name5616 (
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w6972_,
		_w9663_
	);
	LUT2 #(
		.INIT('h1)
	) name5617 (
		_w9660_,
		_w9661_,
		_w9664_
	);
	LUT2 #(
		.INIT('h1)
	) name5618 (
		_w9662_,
		_w9663_,
		_w9665_
	);
	LUT2 #(
		.INIT('h8)
	) name5619 (
		_w9664_,
		_w9665_,
		_w9666_
	);
	LUT2 #(
		.INIT('h8)
	) name5620 (
		_w4055_,
		_w9666_,
		_w9667_
	);
	LUT2 #(
		.INIT('h1)
	) name5621 (
		_w9659_,
		_w9667_,
		_w9668_
	);
	LUT2 #(
		.INIT('h1)
	) name5622 (
		_w8192_,
		_w9668_,
		_w9669_
	);
	LUT2 #(
		.INIT('h2)
	) name5623 (
		_w6135_,
		_w9669_,
		_w9670_
	);
	LUT2 #(
		.INIT('h4)
	) name5624 (
		_w6135_,
		_w7859_,
		_w9671_
	);
	LUT2 #(
		.INIT('h1)
	) name5625 (
		_w6176_,
		_w9670_,
		_w9672_
	);
	LUT2 #(
		.INIT('h4)
	) name5626 (
		_w9671_,
		_w9672_,
		_w9673_
	);
	LUT2 #(
		.INIT('h8)
	) name5627 (
		_w6135_,
		_w8113_,
		_w9674_
	);
	LUT2 #(
		.INIT('h1)
	) name5628 (
		_w6135_,
		_w8224_,
		_w9675_
	);
	LUT2 #(
		.INIT('h2)
	) name5629 (
		_w6176_,
		_w9674_,
		_w9676_
	);
	LUT2 #(
		.INIT('h4)
	) name5630 (
		_w9675_,
		_w9676_,
		_w9677_
	);
	LUT2 #(
		.INIT('h1)
	) name5631 (
		_w9673_,
		_w9677_,
		_w9678_
	);
	LUT2 #(
		.INIT('h2)
	) name5632 (
		_w7005_,
		_w9678_,
		_w9679_
	);
	LUT2 #(
		.INIT('h4)
	) name5633 (
		_w6135_,
		_w8151_,
		_w9680_
	);
	LUT2 #(
		.INIT('h2)
	) name5634 (
		_w6135_,
		_w7644_,
		_w9681_
	);
	LUT2 #(
		.INIT('h2)
	) name5635 (
		_w6176_,
		_w9680_,
		_w9682_
	);
	LUT2 #(
		.INIT('h4)
	) name5636 (
		_w9681_,
		_w9682_,
		_w9683_
	);
	LUT2 #(
		.INIT('h2)
	) name5637 (
		\core_dag_ilm2reg_I_reg[3]/NET0131 ,
		_w6653_,
		_w9684_
	);
	LUT2 #(
		.INIT('h1)
	) name5638 (
		_w6792_,
		_w6793_,
		_w9685_
	);
	LUT2 #(
		.INIT('h1)
	) name5639 (
		_w6817_,
		_w9685_,
		_w9686_
	);
	LUT2 #(
		.INIT('h8)
	) name5640 (
		_w6817_,
		_w9685_,
		_w9687_
	);
	LUT2 #(
		.INIT('h1)
	) name5641 (
		_w9686_,
		_w9687_,
		_w9688_
	);
	LUT2 #(
		.INIT('h8)
	) name5642 (
		_w8198_,
		_w9688_,
		_w9689_
	);
	LUT2 #(
		.INIT('h1)
	) name5643 (
		_w6673_,
		_w6788_,
		_w9690_
	);
	LUT2 #(
		.INIT('h8)
	) name5644 (
		_w6673_,
		_w6788_,
		_w9691_
	);
	LUT2 #(
		.INIT('h1)
	) name5645 (
		_w9690_,
		_w9691_,
		_w9692_
	);
	LUT2 #(
		.INIT('h4)
	) name5646 (
		_w8198_,
		_w9692_,
		_w9693_
	);
	LUT2 #(
		.INIT('h1)
	) name5647 (
		_w9684_,
		_w9689_,
		_w9694_
	);
	LUT2 #(
		.INIT('h4)
	) name5648 (
		_w9693_,
		_w9694_,
		_w9695_
	);
	LUT2 #(
		.INIT('h2)
	) name5649 (
		_w6135_,
		_w9695_,
		_w9696_
	);
	LUT2 #(
		.INIT('h8)
	) name5650 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w6926_,
		_w9697_
	);
	LUT2 #(
		.INIT('h2)
	) name5651 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w6934_,
		_w9698_
	);
	LUT2 #(
		.INIT('h4)
	) name5652 (
		_w6111_,
		_w8192_,
		_w9699_
	);
	LUT2 #(
		.INIT('h8)
	) name5653 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w6956_,
		_w9700_
	);
	LUT2 #(
		.INIT('h4)
	) name5654 (
		_w6121_,
		_w9668_,
		_w9701_
	);
	LUT2 #(
		.INIT('h1)
	) name5655 (
		_w9699_,
		_w9700_,
		_w9702_
	);
	LUT2 #(
		.INIT('h4)
	) name5656 (
		_w9701_,
		_w9702_,
		_w9703_
	);
	LUT2 #(
		.INIT('h2)
	) name5657 (
		_w5949_,
		_w9703_,
		_w9704_
	);
	LUT2 #(
		.INIT('h8)
	) name5658 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[3]/NET0131 ,
		_w6988_,
		_w9705_
	);
	LUT2 #(
		.INIT('h1)
	) name5659 (
		_w9697_,
		_w9705_,
		_w9706_
	);
	LUT2 #(
		.INIT('h4)
	) name5660 (
		_w9698_,
		_w9706_,
		_w9707_
	);
	LUT2 #(
		.INIT('h4)
	) name5661 (
		_w9704_,
		_w9707_,
		_w9708_
	);
	LUT2 #(
		.INIT('h2)
	) name5662 (
		_w6924_,
		_w9708_,
		_w9709_
	);
	LUT2 #(
		.INIT('h2)
	) name5663 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w6924_,
		_w9710_
	);
	LUT2 #(
		.INIT('h1)
	) name5664 (
		_w9709_,
		_w9710_,
		_w9711_
	);
	LUT2 #(
		.INIT('h1)
	) name5665 (
		_w6135_,
		_w9711_,
		_w9712_
	);
	LUT2 #(
		.INIT('h1)
	) name5666 (
		_w6176_,
		_w9712_,
		_w9713_
	);
	LUT2 #(
		.INIT('h4)
	) name5667 (
		_w9696_,
		_w9713_,
		_w9714_
	);
	LUT2 #(
		.INIT('h1)
	) name5668 (
		_w9683_,
		_w9714_,
		_w9715_
	);
	LUT2 #(
		.INIT('h1)
	) name5669 (
		_w7005_,
		_w9715_,
		_w9716_
	);
	LUT2 #(
		.INIT('h1)
	) name5670 (
		_w9679_,
		_w9716_,
		_w9717_
	);
	LUT2 #(
		.INIT('h8)
	) name5671 (
		\core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 ,
		_w6058_,
		_w9718_
	);
	LUT2 #(
		.INIT('h8)
	) name5672 (
		_w6060_,
		_w9718_,
		_w9719_
	);
	LUT2 #(
		.INIT('h8)
	) name5673 (
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w6138_,
		_w9720_
	);
	LUT2 #(
		.INIT('h8)
	) name5674 (
		\core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 ,
		_w6142_,
		_w9721_
	);
	LUT2 #(
		.INIT('h8)
	) name5675 (
		\core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 ,
		_w6140_,
		_w9722_
	);
	LUT2 #(
		.INIT('h1)
	) name5676 (
		_w4055_,
		_w9719_,
		_w9723_
	);
	LUT2 #(
		.INIT('h1)
	) name5677 (
		_w9720_,
		_w9721_,
		_w9724_
	);
	LUT2 #(
		.INIT('h4)
	) name5678 (
		_w9722_,
		_w9724_,
		_w9725_
	);
	LUT2 #(
		.INIT('h8)
	) name5679 (
		_w9723_,
		_w9725_,
		_w9726_
	);
	LUT2 #(
		.INIT('h8)
	) name5680 (
		_w6093_,
		_w9718_,
		_w9727_
	);
	LUT2 #(
		.INIT('h8)
	) name5681 (
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w6152_,
		_w9728_
	);
	LUT2 #(
		.INIT('h8)
	) name5682 (
		\core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 ,
		_w6150_,
		_w9729_
	);
	LUT2 #(
		.INIT('h8)
	) name5683 (
		\core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 ,
		_w6154_,
		_w9730_
	);
	LUT2 #(
		.INIT('h1)
	) name5684 (
		_w9727_,
		_w9728_,
		_w9731_
	);
	LUT2 #(
		.INIT('h1)
	) name5685 (
		_w9729_,
		_w9730_,
		_w9732_
	);
	LUT2 #(
		.INIT('h8)
	) name5686 (
		_w9731_,
		_w9732_,
		_w9733_
	);
	LUT2 #(
		.INIT('h8)
	) name5687 (
		_w4055_,
		_w9733_,
		_w9734_
	);
	LUT2 #(
		.INIT('h1)
	) name5688 (
		_w9726_,
		_w9734_,
		_w9735_
	);
	LUT2 #(
		.INIT('h4)
	) name5689 (
		_w6135_,
		_w9735_,
		_w9736_
	);
	LUT2 #(
		.INIT('h8)
	) name5690 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		_w6389_,
		_w9737_
	);
	LUT2 #(
		.INIT('h1)
	) name5691 (
		_w6410_,
		_w6458_,
		_w9738_
	);
	LUT2 #(
		.INIT('h1)
	) name5692 (
		_w6385_,
		_w6417_,
		_w9739_
	);
	LUT2 #(
		.INIT('h1)
	) name5693 (
		_w6459_,
		_w9739_,
		_w9740_
	);
	LUT2 #(
		.INIT('h2)
	) name5694 (
		_w9738_,
		_w9740_,
		_w9741_
	);
	LUT2 #(
		.INIT('h4)
	) name5695 (
		_w9738_,
		_w9740_,
		_w9742_
	);
	LUT2 #(
		.INIT('h1)
	) name5696 (
		_w9741_,
		_w9742_,
		_w9743_
	);
	LUT2 #(
		.INIT('h1)
	) name5697 (
		_w7631_,
		_w9743_,
		_w9744_
	);
	LUT2 #(
		.INIT('h1)
	) name5698 (
		_w6403_,
		_w6514_,
		_w9745_
	);
	LUT2 #(
		.INIT('h1)
	) name5699 (
		_w6404_,
		_w9745_,
		_w9746_
	);
	LUT2 #(
		.INIT('h2)
	) name5700 (
		_w6393_,
		_w9746_,
		_w9747_
	);
	LUT2 #(
		.INIT('h4)
	) name5701 (
		_w6393_,
		_w9746_,
		_w9748_
	);
	LUT2 #(
		.INIT('h1)
	) name5702 (
		_w9747_,
		_w9748_,
		_w9749_
	);
	LUT2 #(
		.INIT('h8)
	) name5703 (
		_w7631_,
		_w9749_,
		_w9750_
	);
	LUT2 #(
		.INIT('h1)
	) name5704 (
		_w9744_,
		_w9750_,
		_w9751_
	);
	LUT2 #(
		.INIT('h1)
	) name5705 (
		_w9737_,
		_w9751_,
		_w9752_
	);
	LUT2 #(
		.INIT('h2)
	) name5706 (
		_w6135_,
		_w9752_,
		_w9753_
	);
	LUT2 #(
		.INIT('h2)
	) name5707 (
		_w6176_,
		_w9736_,
		_w9754_
	);
	LUT2 #(
		.INIT('h4)
	) name5708 (
		_w9753_,
		_w9754_,
		_w9755_
	);
	LUT2 #(
		.INIT('h8)
	) name5709 (
		\core_dag_ilm2reg_I_reg[4]/NET0131 ,
		_w6684_,
		_w9756_
	);
	LUT2 #(
		.INIT('h1)
	) name5710 (
		_w6675_,
		_w6770_,
		_w9757_
	);
	LUT2 #(
		.INIT('h8)
	) name5711 (
		_w6675_,
		_w6770_,
		_w9758_
	);
	LUT2 #(
		.INIT('h1)
	) name5712 (
		_w9757_,
		_w9758_,
		_w9759_
	);
	LUT2 #(
		.INIT('h4)
	) name5713 (
		_w8198_,
		_w9759_,
		_w9760_
	);
	LUT2 #(
		.INIT('h1)
	) name5714 (
		_w6774_,
		_w6820_,
		_w9761_
	);
	LUT2 #(
		.INIT('h1)
	) name5715 (
		_w6819_,
		_w9761_,
		_w9762_
	);
	LUT2 #(
		.INIT('h8)
	) name5716 (
		_w6819_,
		_w9761_,
		_w9763_
	);
	LUT2 #(
		.INIT('h1)
	) name5717 (
		_w9762_,
		_w9763_,
		_w9764_
	);
	LUT2 #(
		.INIT('h8)
	) name5718 (
		_w8198_,
		_w9764_,
		_w9765_
	);
	LUT2 #(
		.INIT('h1)
	) name5719 (
		_w9756_,
		_w9760_,
		_w9766_
	);
	LUT2 #(
		.INIT('h4)
	) name5720 (
		_w9765_,
		_w9766_,
		_w9767_
	);
	LUT2 #(
		.INIT('h2)
	) name5721 (
		_w6135_,
		_w9767_,
		_w9768_
	);
	LUT2 #(
		.INIT('h8)
	) name5722 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w6926_,
		_w9769_
	);
	LUT2 #(
		.INIT('h2)
	) name5723 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w6934_,
		_w9770_
	);
	LUT2 #(
		.INIT('h8)
	) name5724 (
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		_w6058_,
		_w9771_
	);
	LUT2 #(
		.INIT('h8)
	) name5725 (
		_w6060_,
		_w9771_,
		_w9772_
	);
	LUT2 #(
		.INIT('h8)
	) name5726 (
		\core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 ,
		_w6140_,
		_w9773_
	);
	LUT2 #(
		.INIT('h8)
	) name5727 (
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w6138_,
		_w9774_
	);
	LUT2 #(
		.INIT('h8)
	) name5728 (
		\core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 ,
		_w6142_,
		_w9775_
	);
	LUT2 #(
		.INIT('h1)
	) name5729 (
		_w4055_,
		_w9772_,
		_w9776_
	);
	LUT2 #(
		.INIT('h1)
	) name5730 (
		_w9773_,
		_w9774_,
		_w9777_
	);
	LUT2 #(
		.INIT('h4)
	) name5731 (
		_w9775_,
		_w9777_,
		_w9778_
	);
	LUT2 #(
		.INIT('h8)
	) name5732 (
		_w9776_,
		_w9778_,
		_w9779_
	);
	LUT2 #(
		.INIT('h8)
	) name5733 (
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		_w6148_,
		_w9780_
	);
	LUT2 #(
		.INIT('h8)
	) name5734 (
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w6152_,
		_w9781_
	);
	LUT2 #(
		.INIT('h8)
	) name5735 (
		\core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 ,
		_w6150_,
		_w9782_
	);
	LUT2 #(
		.INIT('h8)
	) name5736 (
		\core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 ,
		_w6154_,
		_w9783_
	);
	LUT2 #(
		.INIT('h1)
	) name5737 (
		_w9780_,
		_w9781_,
		_w9784_
	);
	LUT2 #(
		.INIT('h1)
	) name5738 (
		_w9782_,
		_w9783_,
		_w9785_
	);
	LUT2 #(
		.INIT('h8)
	) name5739 (
		_w9784_,
		_w9785_,
		_w9786_
	);
	LUT2 #(
		.INIT('h8)
	) name5740 (
		_w4055_,
		_w9786_,
		_w9787_
	);
	LUT2 #(
		.INIT('h1)
	) name5741 (
		_w9779_,
		_w9787_,
		_w9788_
	);
	LUT2 #(
		.INIT('h4)
	) name5742 (
		_w6111_,
		_w9788_,
		_w9789_
	);
	LUT2 #(
		.INIT('h8)
	) name5743 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w6956_,
		_w9790_
	);
	LUT2 #(
		.INIT('h8)
	) name5744 (
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w6960_,
		_w9791_
	);
	LUT2 #(
		.INIT('h8)
	) name5745 (
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		_w6964_,
		_w9792_
	);
	LUT2 #(
		.INIT('h8)
	) name5746 (
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w6962_,
		_w9793_
	);
	LUT2 #(
		.INIT('h8)
	) name5747 (
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w6958_,
		_w9794_
	);
	LUT2 #(
		.INIT('h1)
	) name5748 (
		_w9791_,
		_w9792_,
		_w9795_
	);
	LUT2 #(
		.INIT('h1)
	) name5749 (
		_w9793_,
		_w9794_,
		_w9796_
	);
	LUT2 #(
		.INIT('h8)
	) name5750 (
		_w9795_,
		_w9796_,
		_w9797_
	);
	LUT2 #(
		.INIT('h4)
	) name5751 (
		_w4055_,
		_w9797_,
		_w9798_
	);
	LUT2 #(
		.INIT('h8)
	) name5752 (
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w6972_,
		_w9799_
	);
	LUT2 #(
		.INIT('h8)
	) name5753 (
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w6976_,
		_w9800_
	);
	LUT2 #(
		.INIT('h8)
	) name5754 (
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w6974_,
		_w9801_
	);
	LUT2 #(
		.INIT('h8)
	) name5755 (
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		_w6970_,
		_w9802_
	);
	LUT2 #(
		.INIT('h1)
	) name5756 (
		_w9799_,
		_w9800_,
		_w9803_
	);
	LUT2 #(
		.INIT('h1)
	) name5757 (
		_w9801_,
		_w9802_,
		_w9804_
	);
	LUT2 #(
		.INIT('h8)
	) name5758 (
		_w9803_,
		_w9804_,
		_w9805_
	);
	LUT2 #(
		.INIT('h8)
	) name5759 (
		_w4055_,
		_w9805_,
		_w9806_
	);
	LUT2 #(
		.INIT('h1)
	) name5760 (
		_w9798_,
		_w9806_,
		_w9807_
	);
	LUT2 #(
		.INIT('h4)
	) name5761 (
		_w6121_,
		_w9807_,
		_w9808_
	);
	LUT2 #(
		.INIT('h1)
	) name5762 (
		_w9789_,
		_w9790_,
		_w9809_
	);
	LUT2 #(
		.INIT('h4)
	) name5763 (
		_w9808_,
		_w9809_,
		_w9810_
	);
	LUT2 #(
		.INIT('h2)
	) name5764 (
		_w5949_,
		_w9810_,
		_w9811_
	);
	LUT2 #(
		.INIT('h8)
	) name5765 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[4]/NET0131 ,
		_w6988_,
		_w9812_
	);
	LUT2 #(
		.INIT('h1)
	) name5766 (
		_w9769_,
		_w9812_,
		_w9813_
	);
	LUT2 #(
		.INIT('h4)
	) name5767 (
		_w9770_,
		_w9813_,
		_w9814_
	);
	LUT2 #(
		.INIT('h4)
	) name5768 (
		_w9811_,
		_w9814_,
		_w9815_
	);
	LUT2 #(
		.INIT('h2)
	) name5769 (
		_w6924_,
		_w9815_,
		_w9816_
	);
	LUT2 #(
		.INIT('h2)
	) name5770 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w6924_,
		_w9817_
	);
	LUT2 #(
		.INIT('h1)
	) name5771 (
		_w9816_,
		_w9817_,
		_w9818_
	);
	LUT2 #(
		.INIT('h1)
	) name5772 (
		_w6135_,
		_w9818_,
		_w9819_
	);
	LUT2 #(
		.INIT('h1)
	) name5773 (
		_w6176_,
		_w9819_,
		_w9820_
	);
	LUT2 #(
		.INIT('h4)
	) name5774 (
		_w9768_,
		_w9820_,
		_w9821_
	);
	LUT2 #(
		.INIT('h1)
	) name5775 (
		_w9755_,
		_w9821_,
		_w9822_
	);
	LUT2 #(
		.INIT('h1)
	) name5776 (
		_w7005_,
		_w9822_,
		_w9823_
	);
	LUT2 #(
		.INIT('h8)
	) name5777 (
		\DM_rdm[4]_pad ,
		_w7016_,
		_w9824_
	);
	LUT2 #(
		.INIT('h8)
	) name5778 (
		\DM_rd1[4]_pad ,
		_w7022_,
		_w9825_
	);
	LUT2 #(
		.INIT('h8)
	) name5779 (
		\DM_rd4[4]_pad ,
		_w7028_,
		_w9826_
	);
	LUT2 #(
		.INIT('h8)
	) name5780 (
		\DM_rd6[4]_pad ,
		_w7031_,
		_w9827_
	);
	LUT2 #(
		.INIT('h8)
	) name5781 (
		\DM_rd7[4]_pad ,
		_w7034_,
		_w9828_
	);
	LUT2 #(
		.INIT('h8)
	) name5782 (
		\DM_rd3[4]_pad ,
		_w7038_,
		_w9829_
	);
	LUT2 #(
		.INIT('h2)
	) name5783 (
		\DM_rd0[4]_pad ,
		_w7053_,
		_w9830_
	);
	LUT2 #(
		.INIT('h8)
	) name5784 (
		\DM_rd5[4]_pad ,
		_w7043_,
		_w9831_
	);
	LUT2 #(
		.INIT('h8)
	) name5785 (
		\DM_rd2[4]_pad ,
		_w7041_,
		_w9832_
	);
	LUT2 #(
		.INIT('h1)
	) name5786 (
		_w9825_,
		_w9829_,
		_w9833_
	);
	LUT2 #(
		.INIT('h4)
	) name5787 (
		_w9832_,
		_w9833_,
		_w9834_
	);
	LUT2 #(
		.INIT('h1)
	) name5788 (
		_w7057_,
		_w9824_,
		_w9835_
	);
	LUT2 #(
		.INIT('h1)
	) name5789 (
		_w9827_,
		_w9828_,
		_w9836_
	);
	LUT2 #(
		.INIT('h8)
	) name5790 (
		_w9835_,
		_w9836_,
		_w9837_
	);
	LUT2 #(
		.INIT('h4)
	) name5791 (
		_w9826_,
		_w9834_,
		_w9838_
	);
	LUT2 #(
		.INIT('h4)
	) name5792 (
		_w9831_,
		_w9838_,
		_w9839_
	);
	LUT2 #(
		.INIT('h8)
	) name5793 (
		_w9837_,
		_w9839_,
		_w9840_
	);
	LUT2 #(
		.INIT('h4)
	) name5794 (
		_w9830_,
		_w9840_,
		_w9841_
	);
	LUT2 #(
		.INIT('h8)
	) name5795 (
		\regout_STD_C_reg[4]/P0001 ,
		_w6988_,
		_w9842_
	);
	LUT2 #(
		.INIT('h4)
	) name5796 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001 ,
		_w9843_
	);
	LUT2 #(
		.INIT('h8)
	) name5797 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 ,
		_w9844_
	);
	LUT2 #(
		.INIT('h1)
	) name5798 (
		_w9843_,
		_w9844_,
		_w9845_
	);
	LUT2 #(
		.INIT('h2)
	) name5799 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w9845_,
		_w9846_
	);
	LUT2 #(
		.INIT('h4)
	) name5800 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001 ,
		_w9847_
	);
	LUT2 #(
		.INIT('h8)
	) name5801 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001 ,
		_w9848_
	);
	LUT2 #(
		.INIT('h1)
	) name5802 (
		_w9847_,
		_w9848_,
		_w9849_
	);
	LUT2 #(
		.INIT('h2)
	) name5803 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w9849_,
		_w9850_
	);
	LUT2 #(
		.INIT('h4)
	) name5804 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001 ,
		_w9851_
	);
	LUT2 #(
		.INIT('h8)
	) name5805 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001 ,
		_w9852_
	);
	LUT2 #(
		.INIT('h1)
	) name5806 (
		_w9851_,
		_w9852_,
		_w9853_
	);
	LUT2 #(
		.INIT('h2)
	) name5807 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w9853_,
		_w9854_
	);
	LUT2 #(
		.INIT('h4)
	) name5808 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001 ,
		_w9855_
	);
	LUT2 #(
		.INIT('h8)
	) name5809 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001 ,
		_w9856_
	);
	LUT2 #(
		.INIT('h1)
	) name5810 (
		_w9855_,
		_w9856_,
		_w9857_
	);
	LUT2 #(
		.INIT('h2)
	) name5811 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w9857_,
		_w9858_
	);
	LUT2 #(
		.INIT('h4)
	) name5812 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001 ,
		_w9859_
	);
	LUT2 #(
		.INIT('h8)
	) name5813 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001 ,
		_w9860_
	);
	LUT2 #(
		.INIT('h1)
	) name5814 (
		_w9859_,
		_w9860_,
		_w9861_
	);
	LUT2 #(
		.INIT('h2)
	) name5815 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w9861_,
		_w9862_
	);
	LUT2 #(
		.INIT('h4)
	) name5816 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 ,
		_w9863_
	);
	LUT2 #(
		.INIT('h8)
	) name5817 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 ,
		_w9864_
	);
	LUT2 #(
		.INIT('h1)
	) name5818 (
		_w9863_,
		_w9864_,
		_w9865_
	);
	LUT2 #(
		.INIT('h2)
	) name5819 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w9865_,
		_w9866_
	);
	LUT2 #(
		.INIT('h4)
	) name5820 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001 ,
		_w9867_
	);
	LUT2 #(
		.INIT('h8)
	) name5821 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 ,
		_w9868_
	);
	LUT2 #(
		.INIT('h1)
	) name5822 (
		_w9867_,
		_w9868_,
		_w9869_
	);
	LUT2 #(
		.INIT('h2)
	) name5823 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w9869_,
		_w9870_
	);
	LUT2 #(
		.INIT('h1)
	) name5824 (
		_w9846_,
		_w9850_,
		_w9871_
	);
	LUT2 #(
		.INIT('h1)
	) name5825 (
		_w9854_,
		_w9858_,
		_w9872_
	);
	LUT2 #(
		.INIT('h1)
	) name5826 (
		_w9862_,
		_w9866_,
		_w9873_
	);
	LUT2 #(
		.INIT('h4)
	) name5827 (
		_w9870_,
		_w9873_,
		_w9874_
	);
	LUT2 #(
		.INIT('h8)
	) name5828 (
		_w9871_,
		_w9872_,
		_w9875_
	);
	LUT2 #(
		.INIT('h8)
	) name5829 (
		_w9874_,
		_w9875_,
		_w9876_
	);
	LUT2 #(
		.INIT('h2)
	) name5830 (
		_w7179_,
		_w9876_,
		_w9877_
	);
	LUT2 #(
		.INIT('h8)
	) name5831 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131 ,
		_w9878_
	);
	LUT2 #(
		.INIT('h8)
	) name5832 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131 ,
		_w9879_
	);
	LUT2 #(
		.INIT('h8)
	) name5833 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131 ,
		_w9880_
	);
	LUT2 #(
		.INIT('h8)
	) name5834 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131 ,
		_w9881_
	);
	LUT2 #(
		.INIT('h8)
	) name5835 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131 ,
		_w9882_
	);
	LUT2 #(
		.INIT('h8)
	) name5836 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131 ,
		_w9883_
	);
	LUT2 #(
		.INIT('h8)
	) name5837 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131 ,
		_w9884_
	);
	LUT2 #(
		.INIT('h8)
	) name5838 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131 ,
		_w9885_
	);
	LUT2 #(
		.INIT('h8)
	) name5839 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 ,
		_w9886_
	);
	LUT2 #(
		.INIT('h8)
	) name5840 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		_w9887_
	);
	LUT2 #(
		.INIT('h8)
	) name5841 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 ,
		_w9888_
	);
	LUT2 #(
		.INIT('h8)
	) name5842 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w9889_
	);
	LUT2 #(
		.INIT('h1)
	) name5843 (
		_w9878_,
		_w9879_,
		_w9890_
	);
	LUT2 #(
		.INIT('h1)
	) name5844 (
		_w9880_,
		_w9881_,
		_w9891_
	);
	LUT2 #(
		.INIT('h1)
	) name5845 (
		_w9882_,
		_w9883_,
		_w9892_
	);
	LUT2 #(
		.INIT('h1)
	) name5846 (
		_w9884_,
		_w9885_,
		_w9893_
	);
	LUT2 #(
		.INIT('h1)
	) name5847 (
		_w9886_,
		_w9887_,
		_w9894_
	);
	LUT2 #(
		.INIT('h1)
	) name5848 (
		_w9888_,
		_w9889_,
		_w9895_
	);
	LUT2 #(
		.INIT('h8)
	) name5849 (
		_w9894_,
		_w9895_,
		_w9896_
	);
	LUT2 #(
		.INIT('h8)
	) name5850 (
		_w9892_,
		_w9893_,
		_w9897_
	);
	LUT2 #(
		.INIT('h8)
	) name5851 (
		_w9890_,
		_w9891_,
		_w9898_
	);
	LUT2 #(
		.INIT('h8)
	) name5852 (
		_w9897_,
		_w9898_,
		_w9899_
	);
	LUT2 #(
		.INIT('h8)
	) name5853 (
		_w9896_,
		_w9899_,
		_w9900_
	);
	LUT2 #(
		.INIT('h2)
	) name5854 (
		_w7068_,
		_w9900_,
		_w9901_
	);
	LUT2 #(
		.INIT('h4)
	) name5855 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001 ,
		_w9902_
	);
	LUT2 #(
		.INIT('h8)
	) name5856 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001 ,
		_w9903_
	);
	LUT2 #(
		.INIT('h1)
	) name5857 (
		_w9902_,
		_w9903_,
		_w9904_
	);
	LUT2 #(
		.INIT('h2)
	) name5858 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w9904_,
		_w9905_
	);
	LUT2 #(
		.INIT('h4)
	) name5859 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001 ,
		_w9906_
	);
	LUT2 #(
		.INIT('h8)
	) name5860 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001 ,
		_w9907_
	);
	LUT2 #(
		.INIT('h1)
	) name5861 (
		_w9906_,
		_w9907_,
		_w9908_
	);
	LUT2 #(
		.INIT('h2)
	) name5862 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w9908_,
		_w9909_
	);
	LUT2 #(
		.INIT('h4)
	) name5863 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001 ,
		_w9910_
	);
	LUT2 #(
		.INIT('h8)
	) name5864 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001 ,
		_w9911_
	);
	LUT2 #(
		.INIT('h1)
	) name5865 (
		_w9910_,
		_w9911_,
		_w9912_
	);
	LUT2 #(
		.INIT('h2)
	) name5866 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w9912_,
		_w9913_
	);
	LUT2 #(
		.INIT('h4)
	) name5867 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001 ,
		_w9914_
	);
	LUT2 #(
		.INIT('h8)
	) name5868 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001 ,
		_w9915_
	);
	LUT2 #(
		.INIT('h1)
	) name5869 (
		_w9914_,
		_w9915_,
		_w9916_
	);
	LUT2 #(
		.INIT('h2)
	) name5870 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w9916_,
		_w9917_
	);
	LUT2 #(
		.INIT('h4)
	) name5871 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001 ,
		_w9918_
	);
	LUT2 #(
		.INIT('h8)
	) name5872 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001 ,
		_w9919_
	);
	LUT2 #(
		.INIT('h1)
	) name5873 (
		_w9918_,
		_w9919_,
		_w9920_
	);
	LUT2 #(
		.INIT('h2)
	) name5874 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w9920_,
		_w9921_
	);
	LUT2 #(
		.INIT('h8)
	) name5875 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w9922_
	);
	LUT2 #(
		.INIT('h1)
	) name5876 (
		_w9905_,
		_w9922_,
		_w9923_
	);
	LUT2 #(
		.INIT('h1)
	) name5877 (
		_w9909_,
		_w9913_,
		_w9924_
	);
	LUT2 #(
		.INIT('h1)
	) name5878 (
		_w9917_,
		_w9921_,
		_w9925_
	);
	LUT2 #(
		.INIT('h8)
	) name5879 (
		_w9924_,
		_w9925_,
		_w9926_
	);
	LUT2 #(
		.INIT('h8)
	) name5880 (
		_w9923_,
		_w9926_,
		_w9927_
	);
	LUT2 #(
		.INIT('h2)
	) name5881 (
		_w7093_,
		_w9927_,
		_w9928_
	);
	LUT2 #(
		.INIT('h8)
	) name5882 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[4]/P0001 ,
		_w9929_
	);
	LUT2 #(
		.INIT('h8)
	) name5883 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[4]/P0001 ,
		_w9930_
	);
	LUT2 #(
		.INIT('h8)
	) name5884 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[4]/P0001 ,
		_w9931_
	);
	LUT2 #(
		.INIT('h8)
	) name5885 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w9932_
	);
	LUT2 #(
		.INIT('h1)
	) name5886 (
		_w9929_,
		_w9930_,
		_w9933_
	);
	LUT2 #(
		.INIT('h1)
	) name5887 (
		_w9931_,
		_w9932_,
		_w9934_
	);
	LUT2 #(
		.INIT('h8)
	) name5888 (
		_w9933_,
		_w9934_,
		_w9935_
	);
	LUT2 #(
		.INIT('h2)
	) name5889 (
		_w7119_,
		_w9935_,
		_w9936_
	);
	LUT2 #(
		.INIT('h4)
	) name5890 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001 ,
		_w9937_
	);
	LUT2 #(
		.INIT('h8)
	) name5891 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001 ,
		_w9938_
	);
	LUT2 #(
		.INIT('h1)
	) name5892 (
		_w9937_,
		_w9938_,
		_w9939_
	);
	LUT2 #(
		.INIT('h2)
	) name5893 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w9939_,
		_w9940_
	);
	LUT2 #(
		.INIT('h4)
	) name5894 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001 ,
		_w9941_
	);
	LUT2 #(
		.INIT('h8)
	) name5895 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001 ,
		_w9942_
	);
	LUT2 #(
		.INIT('h1)
	) name5896 (
		_w9941_,
		_w9942_,
		_w9943_
	);
	LUT2 #(
		.INIT('h2)
	) name5897 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w9943_,
		_w9944_
	);
	LUT2 #(
		.INIT('h4)
	) name5898 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 ,
		_w9945_
	);
	LUT2 #(
		.INIT('h8)
	) name5899 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 ,
		_w9946_
	);
	LUT2 #(
		.INIT('h1)
	) name5900 (
		_w9945_,
		_w9946_,
		_w9947_
	);
	LUT2 #(
		.INIT('h2)
	) name5901 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w9947_,
		_w9948_
	);
	LUT2 #(
		.INIT('h4)
	) name5902 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 ,
		_w9949_
	);
	LUT2 #(
		.INIT('h8)
	) name5903 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 ,
		_w9950_
	);
	LUT2 #(
		.INIT('h1)
	) name5904 (
		_w9949_,
		_w9950_,
		_w9951_
	);
	LUT2 #(
		.INIT('h2)
	) name5905 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w9951_,
		_w9952_
	);
	LUT2 #(
		.INIT('h1)
	) name5906 (
		_w7169_,
		_w9940_,
		_w9953_
	);
	LUT2 #(
		.INIT('h1)
	) name5907 (
		_w9944_,
		_w9948_,
		_w9954_
	);
	LUT2 #(
		.INIT('h4)
	) name5908 (
		_w9952_,
		_w9954_,
		_w9955_
	);
	LUT2 #(
		.INIT('h8)
	) name5909 (
		_w9953_,
		_w9955_,
		_w9956_
	);
	LUT2 #(
		.INIT('h2)
	) name5910 (
		_w7153_,
		_w9956_,
		_w9957_
	);
	LUT2 #(
		.INIT('h8)
	) name5911 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w9958_
	);
	LUT2 #(
		.INIT('h8)
	) name5912 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w9959_
	);
	LUT2 #(
		.INIT('h8)
	) name5913 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131 ,
		_w9960_
	);
	LUT2 #(
		.INIT('h8)
	) name5914 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131 ,
		_w9961_
	);
	LUT2 #(
		.INIT('h8)
	) name5915 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131 ,
		_w9962_
	);
	LUT2 #(
		.INIT('h8)
	) name5916 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131 ,
		_w9963_
	);
	LUT2 #(
		.INIT('h8)
	) name5917 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		_w9964_
	);
	LUT2 #(
		.INIT('h8)
	) name5918 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w9965_
	);
	LUT2 #(
		.INIT('h8)
	) name5919 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131 ,
		_w9966_
	);
	LUT2 #(
		.INIT('h8)
	) name5920 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131 ,
		_w9967_
	);
	LUT2 #(
		.INIT('h8)
	) name5921 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131 ,
		_w9968_
	);
	LUT2 #(
		.INIT('h8)
	) name5922 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131 ,
		_w9969_
	);
	LUT2 #(
		.INIT('h1)
	) name5923 (
		_w9958_,
		_w9959_,
		_w9970_
	);
	LUT2 #(
		.INIT('h1)
	) name5924 (
		_w9960_,
		_w9961_,
		_w9971_
	);
	LUT2 #(
		.INIT('h1)
	) name5925 (
		_w9962_,
		_w9963_,
		_w9972_
	);
	LUT2 #(
		.INIT('h1)
	) name5926 (
		_w9964_,
		_w9965_,
		_w9973_
	);
	LUT2 #(
		.INIT('h1)
	) name5927 (
		_w9966_,
		_w9967_,
		_w9974_
	);
	LUT2 #(
		.INIT('h1)
	) name5928 (
		_w9968_,
		_w9969_,
		_w9975_
	);
	LUT2 #(
		.INIT('h8)
	) name5929 (
		_w9974_,
		_w9975_,
		_w9976_
	);
	LUT2 #(
		.INIT('h8)
	) name5930 (
		_w9972_,
		_w9973_,
		_w9977_
	);
	LUT2 #(
		.INIT('h8)
	) name5931 (
		_w9970_,
		_w9971_,
		_w9978_
	);
	LUT2 #(
		.INIT('h8)
	) name5932 (
		_w9977_,
		_w9978_,
		_w9979_
	);
	LUT2 #(
		.INIT('h8)
	) name5933 (
		_w9976_,
		_w9979_,
		_w9980_
	);
	LUT2 #(
		.INIT('h2)
	) name5934 (
		_w7128_,
		_w9980_,
		_w9981_
	);
	LUT2 #(
		.INIT('h8)
	) name5935 (
		\idma_DOVL_reg[4]/NET0131 ,
		_w7532_,
		_w9982_
	);
	LUT2 #(
		.INIT('h8)
	) name5936 (
		\sport0_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w7295_,
		_w9983_
	);
	LUT2 #(
		.INIT('h8)
	) name5937 (
		\tm_tpr_reg_DO_reg[4]/NET0131 ,
		_w7293_,
		_w9984_
	);
	LUT2 #(
		.INIT('h8)
	) name5938 (
		\bdma_BWCOUNT_reg[4]/NET0131 ,
		_w7287_,
		_w9985_
	);
	LUT2 #(
		.INIT('h8)
	) name5939 (
		\emc_WSCRreg_DO_reg[4]/NET0131 ,
		_w7251_,
		_w9986_
	);
	LUT2 #(
		.INIT('h8)
	) name5940 (
		\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w7256_,
		_w9987_
	);
	LUT2 #(
		.INIT('h8)
	) name5941 (
		\sport1_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w7263_,
		_w9988_
	);
	LUT2 #(
		.INIT('h8)
	) name5942 (
		\tm_tsr_reg_DO_reg[4]/NET0131 ,
		_w7540_,
		_w9989_
	);
	LUT2 #(
		.INIT('h8)
	) name5943 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w7249_,
		_w9990_
	);
	LUT2 #(
		.INIT('h8)
	) name5944 (
		\emc_WSCRext_reg_DO_reg[4]/NET0131 ,
		_w7514_,
		_w9991_
	);
	LUT2 #(
		.INIT('h8)
	) name5945 (
		\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w7247_,
		_w9992_
	);
	LUT2 #(
		.INIT('h8)
	) name5946 (
		\sport1_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w7281_,
		_w9993_
	);
	LUT2 #(
		.INIT('h8)
	) name5947 (
		\pio_pmask_reg_DO_reg[4]/NET0131 ,
		_w7297_,
		_w9994_
	);
	LUT2 #(
		.INIT('h8)
	) name5948 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w7234_,
		_w9995_
	);
	LUT2 #(
		.INIT('h8)
	) name5949 (
		\sport0_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w7276_,
		_w9996_
	);
	LUT2 #(
		.INIT('h8)
	) name5950 (
		\sport1_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w7527_,
		_w9997_
	);
	LUT2 #(
		.INIT('h8)
	) name5951 (
		\tm_TCR_TMP_reg[4]/NET0131 ,
		_w7289_,
		_w9998_
	);
	LUT2 #(
		.INIT('h8)
	) name5952 (
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w7259_,
		_w9999_
	);
	LUT2 #(
		.INIT('h8)
	) name5953 (
		\bdma_BOVL_reg[4]/NET0131 ,
		_w7534_,
		_w10000_
	);
	LUT2 #(
		.INIT('h8)
	) name5954 (
		\clkc_ckr_reg_DO_reg[4]/NET0131 ,
		_w7239_,
		_w10001_
	);
	LUT2 #(
		.INIT('h8)
	) name5955 (
		\memc_usysr_DO_reg[4]/NET0131 ,
		_w7301_,
		_w10002_
	);
	LUT2 #(
		.INIT('h8)
	) name5956 (
		\bdma_BEAD_reg[4]/NET0131 ,
		_w7303_,
		_w10003_
	);
	LUT2 #(
		.INIT('h8)
	) name5957 (
		\bdma_BCTL_reg[4]/NET0131 ,
		_w7230_,
		_w10004_
	);
	LUT2 #(
		.INIT('h8)
	) name5958 (
		\pio_PINT_reg[4]/NET0131 ,
		_w7271_,
		_w10005_
	);
	LUT2 #(
		.INIT('h8)
	) name5959 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w7299_,
		_w10006_
	);
	LUT2 #(
		.INIT('h8)
	) name5960 (
		\PIO_out[4]_pad ,
		_w7291_,
		_w10007_
	);
	LUT2 #(
		.INIT('h8)
	) name5961 (
		\PIO_oe[4]_pad ,
		_w7244_,
		_w10008_
	);
	LUT2 #(
		.INIT('h8)
	) name5962 (
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w7273_,
		_w10009_
	);
	LUT2 #(
		.INIT('h1)
	) name5963 (
		_w7522_,
		_w9982_,
		_w10010_
	);
	LUT2 #(
		.INIT('h1)
	) name5964 (
		_w9983_,
		_w9984_,
		_w10011_
	);
	LUT2 #(
		.INIT('h1)
	) name5965 (
		_w9986_,
		_w9987_,
		_w10012_
	);
	LUT2 #(
		.INIT('h1)
	) name5966 (
		_w9988_,
		_w9989_,
		_w10013_
	);
	LUT2 #(
		.INIT('h1)
	) name5967 (
		_w9990_,
		_w9991_,
		_w10014_
	);
	LUT2 #(
		.INIT('h1)
	) name5968 (
		_w9992_,
		_w9993_,
		_w10015_
	);
	LUT2 #(
		.INIT('h1)
	) name5969 (
		_w9994_,
		_w9996_,
		_w10016_
	);
	LUT2 #(
		.INIT('h1)
	) name5970 (
		_w9997_,
		_w9998_,
		_w10017_
	);
	LUT2 #(
		.INIT('h1)
	) name5971 (
		_w9999_,
		_w10001_,
		_w10018_
	);
	LUT2 #(
		.INIT('h1)
	) name5972 (
		_w10002_,
		_w10005_,
		_w10019_
	);
	LUT2 #(
		.INIT('h1)
	) name5973 (
		_w10006_,
		_w10007_,
		_w10020_
	);
	LUT2 #(
		.INIT('h1)
	) name5974 (
		_w10008_,
		_w10009_,
		_w10021_
	);
	LUT2 #(
		.INIT('h8)
	) name5975 (
		_w10020_,
		_w10021_,
		_w10022_
	);
	LUT2 #(
		.INIT('h8)
	) name5976 (
		_w10018_,
		_w10019_,
		_w10023_
	);
	LUT2 #(
		.INIT('h8)
	) name5977 (
		_w10016_,
		_w10017_,
		_w10024_
	);
	LUT2 #(
		.INIT('h8)
	) name5978 (
		_w10014_,
		_w10015_,
		_w10025_
	);
	LUT2 #(
		.INIT('h8)
	) name5979 (
		_w10012_,
		_w10013_,
		_w10026_
	);
	LUT2 #(
		.INIT('h8)
	) name5980 (
		_w10010_,
		_w10011_,
		_w10027_
	);
	LUT2 #(
		.INIT('h8)
	) name5981 (
		_w10026_,
		_w10027_,
		_w10028_
	);
	LUT2 #(
		.INIT('h8)
	) name5982 (
		_w10024_,
		_w10025_,
		_w10029_
	);
	LUT2 #(
		.INIT('h8)
	) name5983 (
		_w10022_,
		_w10023_,
		_w10030_
	);
	LUT2 #(
		.INIT('h8)
	) name5984 (
		_w10029_,
		_w10030_,
		_w10031_
	);
	LUT2 #(
		.INIT('h4)
	) name5985 (
		_w9995_,
		_w10028_,
		_w10032_
	);
	LUT2 #(
		.INIT('h1)
	) name5986 (
		_w10003_,
		_w10004_,
		_w10033_
	);
	LUT2 #(
		.INIT('h8)
	) name5987 (
		_w10032_,
		_w10033_,
		_w10034_
	);
	LUT2 #(
		.INIT('h4)
	) name5988 (
		_w9985_,
		_w10031_,
		_w10035_
	);
	LUT2 #(
		.INIT('h4)
	) name5989 (
		_w10000_,
		_w10035_,
		_w10036_
	);
	LUT2 #(
		.INIT('h8)
	) name5990 (
		_w10034_,
		_w10036_,
		_w10037_
	);
	LUT2 #(
		.INIT('h2)
	) name5991 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w10037_,
		_w10038_
	);
	LUT2 #(
		.INIT('h8)
	) name5992 (
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w10039_
	);
	LUT2 #(
		.INIT('h2)
	) name5993 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7216_,
		_w10040_
	);
	LUT2 #(
		.INIT('h8)
	) name5994 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w10041_
	);
	LUT2 #(
		.INIT('h2)
	) name5995 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4360_,
		_w10042_
	);
	LUT2 #(
		.INIT('h8)
	) name5996 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w10043_
	);
	LUT2 #(
		.INIT('h8)
	) name5997 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w10044_
	);
	LUT2 #(
		.INIT('h8)
	) name5998 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		_w10045_
	);
	LUT2 #(
		.INIT('h8)
	) name5999 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w10046_
	);
	LUT2 #(
		.INIT('h8)
	) name6000 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[4]/NET0131 ,
		_w10047_
	);
	LUT2 #(
		.INIT('h1)
	) name6001 (
		_w10039_,
		_w10041_,
		_w10048_
	);
	LUT2 #(
		.INIT('h1)
	) name6002 (
		_w10043_,
		_w10044_,
		_w10049_
	);
	LUT2 #(
		.INIT('h1)
	) name6003 (
		_w10045_,
		_w10046_,
		_w10050_
	);
	LUT2 #(
		.INIT('h4)
	) name6004 (
		_w10047_,
		_w10050_,
		_w10051_
	);
	LUT2 #(
		.INIT('h8)
	) name6005 (
		_w10048_,
		_w10049_,
		_w10052_
	);
	LUT2 #(
		.INIT('h4)
	) name6006 (
		_w10040_,
		_w10052_,
		_w10053_
	);
	LUT2 #(
		.INIT('h8)
	) name6007 (
		_w10051_,
		_w10053_,
		_w10054_
	);
	LUT2 #(
		.INIT('h4)
	) name6008 (
		_w10042_,
		_w10054_,
		_w10055_
	);
	LUT2 #(
		.INIT('h2)
	) name6009 (
		_w7215_,
		_w10055_,
		_w10056_
	);
	LUT2 #(
		.INIT('h1)
	) name6010 (
		_w9901_,
		_w9936_,
		_w10057_
	);
	LUT2 #(
		.INIT('h4)
	) name6011 (
		_w9981_,
		_w10057_,
		_w10058_
	);
	LUT2 #(
		.INIT('h1)
	) name6012 (
		_w9877_,
		_w9928_,
		_w10059_
	);
	LUT2 #(
		.INIT('h4)
	) name6013 (
		_w9957_,
		_w10059_,
		_w10060_
	);
	LUT2 #(
		.INIT('h8)
	) name6014 (
		_w10058_,
		_w10060_,
		_w10061_
	);
	LUT2 #(
		.INIT('h4)
	) name6015 (
		_w10056_,
		_w10061_,
		_w10062_
	);
	LUT2 #(
		.INIT('h4)
	) name6016 (
		_w10038_,
		_w10062_,
		_w10063_
	);
	LUT2 #(
		.INIT('h4)
	) name6017 (
		_w9842_,
		_w10063_,
		_w10064_
	);
	LUT2 #(
		.INIT('h1)
	) name6018 (
		\emc_DMDoe_reg/NET0131 ,
		_w10064_,
		_w10065_
	);
	LUT2 #(
		.INIT('h8)
	) name6019 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[4]/P0001 ,
		_w10066_
	);
	LUT2 #(
		.INIT('h2)
	) name6020 (
		_w7057_,
		_w10066_,
		_w10067_
	);
	LUT2 #(
		.INIT('h4)
	) name6021 (
		_w10065_,
		_w10067_,
		_w10068_
	);
	LUT2 #(
		.INIT('h1)
	) name6022 (
		_w9841_,
		_w10068_,
		_w10069_
	);
	LUT2 #(
		.INIT('h2)
	) name6023 (
		_w6176_,
		_w10069_,
		_w10070_
	);
	LUT2 #(
		.INIT('h1)
	) name6024 (
		_w9788_,
		_w9807_,
		_w10071_
	);
	LUT2 #(
		.INIT('h4)
	) name6025 (
		_w6176_,
		_w10071_,
		_w10072_
	);
	LUT2 #(
		.INIT('h2)
	) name6026 (
		_w6135_,
		_w10070_,
		_w10073_
	);
	LUT2 #(
		.INIT('h4)
	) name6027 (
		_w10072_,
		_w10073_,
		_w10074_
	);
	LUT2 #(
		.INIT('h8)
	) name6028 (
		\DM_rdm[9]_pad ,
		_w7016_,
		_w10075_
	);
	LUT2 #(
		.INIT('h8)
	) name6029 (
		\DM_rd1[9]_pad ,
		_w7022_,
		_w10076_
	);
	LUT2 #(
		.INIT('h8)
	) name6030 (
		\DM_rd5[9]_pad ,
		_w7043_,
		_w10077_
	);
	LUT2 #(
		.INIT('h8)
	) name6031 (
		\DM_rd6[9]_pad ,
		_w7031_,
		_w10078_
	);
	LUT2 #(
		.INIT('h8)
	) name6032 (
		\DM_rd7[9]_pad ,
		_w7034_,
		_w10079_
	);
	LUT2 #(
		.INIT('h8)
	) name6033 (
		\DM_rd3[9]_pad ,
		_w7038_,
		_w10080_
	);
	LUT2 #(
		.INIT('h2)
	) name6034 (
		\DM_rd0[9]_pad ,
		_w7053_,
		_w10081_
	);
	LUT2 #(
		.INIT('h8)
	) name6035 (
		\DM_rd4[9]_pad ,
		_w7028_,
		_w10082_
	);
	LUT2 #(
		.INIT('h8)
	) name6036 (
		\DM_rd2[9]_pad ,
		_w7041_,
		_w10083_
	);
	LUT2 #(
		.INIT('h1)
	) name6037 (
		_w10076_,
		_w10080_,
		_w10084_
	);
	LUT2 #(
		.INIT('h4)
	) name6038 (
		_w10083_,
		_w10084_,
		_w10085_
	);
	LUT2 #(
		.INIT('h1)
	) name6039 (
		_w7057_,
		_w10075_,
		_w10086_
	);
	LUT2 #(
		.INIT('h1)
	) name6040 (
		_w10078_,
		_w10079_,
		_w10087_
	);
	LUT2 #(
		.INIT('h8)
	) name6041 (
		_w10086_,
		_w10087_,
		_w10088_
	);
	LUT2 #(
		.INIT('h4)
	) name6042 (
		_w10077_,
		_w10085_,
		_w10089_
	);
	LUT2 #(
		.INIT('h4)
	) name6043 (
		_w10082_,
		_w10089_,
		_w10090_
	);
	LUT2 #(
		.INIT('h8)
	) name6044 (
		_w10088_,
		_w10090_,
		_w10091_
	);
	LUT2 #(
		.INIT('h4)
	) name6045 (
		_w10081_,
		_w10091_,
		_w10092_
	);
	LUT2 #(
		.INIT('h8)
	) name6046 (
		\regout_STD_C_reg[9]/P0001 ,
		_w6988_,
		_w10093_
	);
	LUT2 #(
		.INIT('h4)
	) name6047 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001 ,
		_w10094_
	);
	LUT2 #(
		.INIT('h8)
	) name6048 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 ,
		_w10095_
	);
	LUT2 #(
		.INIT('h1)
	) name6049 (
		_w10094_,
		_w10095_,
		_w10096_
	);
	LUT2 #(
		.INIT('h2)
	) name6050 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w10096_,
		_w10097_
	);
	LUT2 #(
		.INIT('h4)
	) name6051 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001 ,
		_w10098_
	);
	LUT2 #(
		.INIT('h8)
	) name6052 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001 ,
		_w10099_
	);
	LUT2 #(
		.INIT('h1)
	) name6053 (
		_w10098_,
		_w10099_,
		_w10100_
	);
	LUT2 #(
		.INIT('h2)
	) name6054 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w10100_,
		_w10101_
	);
	LUT2 #(
		.INIT('h4)
	) name6055 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001 ,
		_w10102_
	);
	LUT2 #(
		.INIT('h8)
	) name6056 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001 ,
		_w10103_
	);
	LUT2 #(
		.INIT('h1)
	) name6057 (
		_w10102_,
		_w10103_,
		_w10104_
	);
	LUT2 #(
		.INIT('h2)
	) name6058 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w10104_,
		_w10105_
	);
	LUT2 #(
		.INIT('h4)
	) name6059 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001 ,
		_w10106_
	);
	LUT2 #(
		.INIT('h8)
	) name6060 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001 ,
		_w10107_
	);
	LUT2 #(
		.INIT('h1)
	) name6061 (
		_w10106_,
		_w10107_,
		_w10108_
	);
	LUT2 #(
		.INIT('h2)
	) name6062 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w10108_,
		_w10109_
	);
	LUT2 #(
		.INIT('h4)
	) name6063 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001 ,
		_w10110_
	);
	LUT2 #(
		.INIT('h8)
	) name6064 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 ,
		_w10111_
	);
	LUT2 #(
		.INIT('h1)
	) name6065 (
		_w10110_,
		_w10111_,
		_w10112_
	);
	LUT2 #(
		.INIT('h2)
	) name6066 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w10112_,
		_w10113_
	);
	LUT2 #(
		.INIT('h4)
	) name6067 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001 ,
		_w10114_
	);
	LUT2 #(
		.INIT('h8)
	) name6068 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001 ,
		_w10115_
	);
	LUT2 #(
		.INIT('h1)
	) name6069 (
		_w10114_,
		_w10115_,
		_w10116_
	);
	LUT2 #(
		.INIT('h2)
	) name6070 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w10116_,
		_w10117_
	);
	LUT2 #(
		.INIT('h1)
	) name6071 (
		_w7207_,
		_w10097_,
		_w10118_
	);
	LUT2 #(
		.INIT('h1)
	) name6072 (
		_w10101_,
		_w10105_,
		_w10119_
	);
	LUT2 #(
		.INIT('h1)
	) name6073 (
		_w10109_,
		_w10113_,
		_w10120_
	);
	LUT2 #(
		.INIT('h4)
	) name6074 (
		_w10117_,
		_w10120_,
		_w10121_
	);
	LUT2 #(
		.INIT('h8)
	) name6075 (
		_w10118_,
		_w10119_,
		_w10122_
	);
	LUT2 #(
		.INIT('h8)
	) name6076 (
		_w10121_,
		_w10122_,
		_w10123_
	);
	LUT2 #(
		.INIT('h2)
	) name6077 (
		_w7179_,
		_w10123_,
		_w10124_
	);
	LUT2 #(
		.INIT('h8)
	) name6078 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131 ,
		_w10125_
	);
	LUT2 #(
		.INIT('h8)
	) name6079 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131 ,
		_w10126_
	);
	LUT2 #(
		.INIT('h8)
	) name6080 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131 ,
		_w10127_
	);
	LUT2 #(
		.INIT('h8)
	) name6081 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131 ,
		_w10128_
	);
	LUT2 #(
		.INIT('h8)
	) name6082 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 ,
		_w10129_
	);
	LUT2 #(
		.INIT('h8)
	) name6083 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131 ,
		_w10130_
	);
	LUT2 #(
		.INIT('h8)
	) name6084 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w10131_
	);
	LUT2 #(
		.INIT('h8)
	) name6085 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131 ,
		_w10132_
	);
	LUT2 #(
		.INIT('h8)
	) name6086 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 ,
		_w10133_
	);
	LUT2 #(
		.INIT('h8)
	) name6087 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 ,
		_w10134_
	);
	LUT2 #(
		.INIT('h8)
	) name6088 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131 ,
		_w10135_
	);
	LUT2 #(
		.INIT('h8)
	) name6089 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131 ,
		_w10136_
	);
	LUT2 #(
		.INIT('h1)
	) name6090 (
		_w10125_,
		_w10126_,
		_w10137_
	);
	LUT2 #(
		.INIT('h1)
	) name6091 (
		_w10127_,
		_w10128_,
		_w10138_
	);
	LUT2 #(
		.INIT('h1)
	) name6092 (
		_w10129_,
		_w10130_,
		_w10139_
	);
	LUT2 #(
		.INIT('h1)
	) name6093 (
		_w10131_,
		_w10132_,
		_w10140_
	);
	LUT2 #(
		.INIT('h1)
	) name6094 (
		_w10133_,
		_w10134_,
		_w10141_
	);
	LUT2 #(
		.INIT('h1)
	) name6095 (
		_w10135_,
		_w10136_,
		_w10142_
	);
	LUT2 #(
		.INIT('h8)
	) name6096 (
		_w10141_,
		_w10142_,
		_w10143_
	);
	LUT2 #(
		.INIT('h8)
	) name6097 (
		_w10139_,
		_w10140_,
		_w10144_
	);
	LUT2 #(
		.INIT('h8)
	) name6098 (
		_w10137_,
		_w10138_,
		_w10145_
	);
	LUT2 #(
		.INIT('h8)
	) name6099 (
		_w10144_,
		_w10145_,
		_w10146_
	);
	LUT2 #(
		.INIT('h8)
	) name6100 (
		_w10143_,
		_w10146_,
		_w10147_
	);
	LUT2 #(
		.INIT('h2)
	) name6101 (
		_w7068_,
		_w10147_,
		_w10148_
	);
	LUT2 #(
		.INIT('h8)
	) name6102 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131 ,
		_w10149_
	);
	LUT2 #(
		.INIT('h8)
	) name6103 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131 ,
		_w10150_
	);
	LUT2 #(
		.INIT('h8)
	) name6104 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131 ,
		_w10151_
	);
	LUT2 #(
		.INIT('h8)
	) name6105 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w10152_
	);
	LUT2 #(
		.INIT('h8)
	) name6106 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w10153_
	);
	LUT2 #(
		.INIT('h8)
	) name6107 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w10154_
	);
	LUT2 #(
		.INIT('h8)
	) name6108 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131 ,
		_w10155_
	);
	LUT2 #(
		.INIT('h8)
	) name6109 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131 ,
		_w10156_
	);
	LUT2 #(
		.INIT('h8)
	) name6110 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131 ,
		_w10157_
	);
	LUT2 #(
		.INIT('h8)
	) name6111 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131 ,
		_w10158_
	);
	LUT2 #(
		.INIT('h8)
	) name6112 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131 ,
		_w10159_
	);
	LUT2 #(
		.INIT('h8)
	) name6113 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w10160_
	);
	LUT2 #(
		.INIT('h1)
	) name6114 (
		_w10149_,
		_w10150_,
		_w10161_
	);
	LUT2 #(
		.INIT('h1)
	) name6115 (
		_w10151_,
		_w10152_,
		_w10162_
	);
	LUT2 #(
		.INIT('h1)
	) name6116 (
		_w10153_,
		_w10154_,
		_w10163_
	);
	LUT2 #(
		.INIT('h1)
	) name6117 (
		_w10155_,
		_w10156_,
		_w10164_
	);
	LUT2 #(
		.INIT('h1)
	) name6118 (
		_w10157_,
		_w10158_,
		_w10165_
	);
	LUT2 #(
		.INIT('h1)
	) name6119 (
		_w10159_,
		_w10160_,
		_w10166_
	);
	LUT2 #(
		.INIT('h8)
	) name6120 (
		_w10165_,
		_w10166_,
		_w10167_
	);
	LUT2 #(
		.INIT('h8)
	) name6121 (
		_w10163_,
		_w10164_,
		_w10168_
	);
	LUT2 #(
		.INIT('h8)
	) name6122 (
		_w10161_,
		_w10162_,
		_w10169_
	);
	LUT2 #(
		.INIT('h8)
	) name6123 (
		_w10168_,
		_w10169_,
		_w10170_
	);
	LUT2 #(
		.INIT('h8)
	) name6124 (
		_w10167_,
		_w10170_,
		_w10171_
	);
	LUT2 #(
		.INIT('h2)
	) name6125 (
		_w7128_,
		_w10171_,
		_w10172_
	);
	LUT2 #(
		.INIT('h4)
	) name6126 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001 ,
		_w10173_
	);
	LUT2 #(
		.INIT('h8)
	) name6127 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001 ,
		_w10174_
	);
	LUT2 #(
		.INIT('h1)
	) name6128 (
		_w10173_,
		_w10174_,
		_w10175_
	);
	LUT2 #(
		.INIT('h2)
	) name6129 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w10175_,
		_w10176_
	);
	LUT2 #(
		.INIT('h4)
	) name6130 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001 ,
		_w10177_
	);
	LUT2 #(
		.INIT('h8)
	) name6131 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001 ,
		_w10178_
	);
	LUT2 #(
		.INIT('h1)
	) name6132 (
		_w10177_,
		_w10178_,
		_w10179_
	);
	LUT2 #(
		.INIT('h2)
	) name6133 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w10179_,
		_w10180_
	);
	LUT2 #(
		.INIT('h4)
	) name6134 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001 ,
		_w10181_
	);
	LUT2 #(
		.INIT('h8)
	) name6135 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001 ,
		_w10182_
	);
	LUT2 #(
		.INIT('h1)
	) name6136 (
		_w10181_,
		_w10182_,
		_w10183_
	);
	LUT2 #(
		.INIT('h2)
	) name6137 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w10183_,
		_w10184_
	);
	LUT2 #(
		.INIT('h4)
	) name6138 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001 ,
		_w10185_
	);
	LUT2 #(
		.INIT('h8)
	) name6139 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001 ,
		_w10186_
	);
	LUT2 #(
		.INIT('h1)
	) name6140 (
		_w10185_,
		_w10186_,
		_w10187_
	);
	LUT2 #(
		.INIT('h2)
	) name6141 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w10187_,
		_w10188_
	);
	LUT2 #(
		.INIT('h4)
	) name6142 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001 ,
		_w10189_
	);
	LUT2 #(
		.INIT('h8)
	) name6143 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001 ,
		_w10190_
	);
	LUT2 #(
		.INIT('h1)
	) name6144 (
		_w10189_,
		_w10190_,
		_w10191_
	);
	LUT2 #(
		.INIT('h2)
	) name6145 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w10191_,
		_w10192_
	);
	LUT2 #(
		.INIT('h1)
	) name6146 (
		_w10176_,
		_w10180_,
		_w10193_
	);
	LUT2 #(
		.INIT('h1)
	) name6147 (
		_w10184_,
		_w10188_,
		_w10194_
	);
	LUT2 #(
		.INIT('h4)
	) name6148 (
		_w10192_,
		_w10194_,
		_w10195_
	);
	LUT2 #(
		.INIT('h8)
	) name6149 (
		_w10193_,
		_w10195_,
		_w10196_
	);
	LUT2 #(
		.INIT('h2)
	) name6150 (
		_w7093_,
		_w10196_,
		_w10197_
	);
	LUT2 #(
		.INIT('h8)
	) name6151 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[9]/P0001 ,
		_w10198_
	);
	LUT2 #(
		.INIT('h8)
	) name6152 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[9]/P0001 ,
		_w10199_
	);
	LUT2 #(
		.INIT('h8)
	) name6153 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[9]/P0001 ,
		_w10200_
	);
	LUT2 #(
		.INIT('h8)
	) name6154 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w10201_
	);
	LUT2 #(
		.INIT('h1)
	) name6155 (
		_w10198_,
		_w10199_,
		_w10202_
	);
	LUT2 #(
		.INIT('h1)
	) name6156 (
		_w10200_,
		_w10201_,
		_w10203_
	);
	LUT2 #(
		.INIT('h8)
	) name6157 (
		_w10202_,
		_w10203_,
		_w10204_
	);
	LUT2 #(
		.INIT('h2)
	) name6158 (
		_w7119_,
		_w10204_,
		_w10205_
	);
	LUT2 #(
		.INIT('h8)
	) name6159 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w10206_
	);
	LUT2 #(
		.INIT('h2)
	) name6160 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4554_,
		_w10207_
	);
	LUT2 #(
		.INIT('h8)
	) name6161 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w10208_
	);
	LUT2 #(
		.INIT('h2)
	) name6162 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w7216_,
		_w10209_
	);
	LUT2 #(
		.INIT('h8)
	) name6163 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w10210_
	);
	LUT2 #(
		.INIT('h1)
	) name6164 (
		_w10206_,
		_w10208_,
		_w10211_
	);
	LUT2 #(
		.INIT('h4)
	) name6165 (
		_w10210_,
		_w10211_,
		_w10212_
	);
	LUT2 #(
		.INIT('h4)
	) name6166 (
		_w10209_,
		_w10212_,
		_w10213_
	);
	LUT2 #(
		.INIT('h4)
	) name6167 (
		_w10207_,
		_w10213_,
		_w10214_
	);
	LUT2 #(
		.INIT('h2)
	) name6168 (
		_w7215_,
		_w10214_,
		_w10215_
	);
	LUT2 #(
		.INIT('h4)
	) name6169 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 ,
		_w10216_
	);
	LUT2 #(
		.INIT('h8)
	) name6170 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 ,
		_w10217_
	);
	LUT2 #(
		.INIT('h1)
	) name6171 (
		_w10216_,
		_w10217_,
		_w10218_
	);
	LUT2 #(
		.INIT('h2)
	) name6172 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w10218_,
		_w10219_
	);
	LUT2 #(
		.INIT('h4)
	) name6173 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001 ,
		_w10220_
	);
	LUT2 #(
		.INIT('h8)
	) name6174 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001 ,
		_w10221_
	);
	LUT2 #(
		.INIT('h1)
	) name6175 (
		_w10220_,
		_w10221_,
		_w10222_
	);
	LUT2 #(
		.INIT('h2)
	) name6176 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w10222_,
		_w10223_
	);
	LUT2 #(
		.INIT('h4)
	) name6177 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 ,
		_w10224_
	);
	LUT2 #(
		.INIT('h8)
	) name6178 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 ,
		_w10225_
	);
	LUT2 #(
		.INIT('h1)
	) name6179 (
		_w10224_,
		_w10225_,
		_w10226_
	);
	LUT2 #(
		.INIT('h2)
	) name6180 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w10226_,
		_w10227_
	);
	LUT2 #(
		.INIT('h1)
	) name6181 (
		_w10219_,
		_w10223_,
		_w10228_
	);
	LUT2 #(
		.INIT('h4)
	) name6182 (
		_w10227_,
		_w10228_,
		_w10229_
	);
	LUT2 #(
		.INIT('h8)
	) name6183 (
		_w7174_,
		_w10229_,
		_w10230_
	);
	LUT2 #(
		.INIT('h2)
	) name6184 (
		_w7153_,
		_w10230_,
		_w10231_
	);
	LUT2 #(
		.INIT('h8)
	) name6185 (
		\tm_tpr_reg_DO_reg[9]/NET0131 ,
		_w7293_,
		_w10232_
	);
	LUT2 #(
		.INIT('h8)
	) name6186 (
		\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w7256_,
		_w10233_
	);
	LUT2 #(
		.INIT('h8)
	) name6187 (
		\bdma_BCTL_reg[9]/NET0131 ,
		_w7230_,
		_w10234_
	);
	LUT2 #(
		.INIT('h8)
	) name6188 (
		\idma_DOVL_reg[9]/NET0131 ,
		_w7532_,
		_w10235_
	);
	LUT2 #(
		.INIT('h8)
	) name6189 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w7234_,
		_w10236_
	);
	LUT2 #(
		.INIT('h8)
	) name6190 (
		\bdma_BOVL_reg[9]/NET0131 ,
		_w7534_,
		_w10237_
	);
	LUT2 #(
		.INIT('h8)
	) name6191 (
		\emc_WSCRreg_DO_reg[9]/NET0131 ,
		_w7251_,
		_w10238_
	);
	LUT2 #(
		.INIT('h8)
	) name6192 (
		\bdma_BEAD_reg[9]/NET0131 ,
		_w7303_,
		_w10239_
	);
	LUT2 #(
		.INIT('h8)
	) name6193 (
		\ITFS1_pad ,
		_w7281_,
		_w10240_
	);
	LUT2 #(
		.INIT('h8)
	) name6194 (
		\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w7247_,
		_w10241_
	);
	LUT2 #(
		.INIT('h8)
	) name6195 (
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w7289_,
		_w10242_
	);
	LUT2 #(
		.INIT('h8)
	) name6196 (
		\sport0_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w7295_,
		_w10243_
	);
	LUT2 #(
		.INIT('h8)
	) name6197 (
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w7273_,
		_w10244_
	);
	LUT2 #(
		.INIT('h8)
	) name6198 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w7299_,
		_w10245_
	);
	LUT2 #(
		.INIT('h8)
	) name6199 (
		\ITFS0_pad ,
		_w7249_,
		_w10246_
	);
	LUT2 #(
		.INIT('h8)
	) name6200 (
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w7259_,
		_w10247_
	);
	LUT2 #(
		.INIT('h8)
	) name6201 (
		\bdma_BWCOUNT_reg[9]/NET0131 ,
		_w7287_,
		_w10248_
	);
	LUT2 #(
		.INIT('h8)
	) name6202 (
		\sport0_txctl_Wcnt_reg[1]/NET0131 ,
		_w7710_,
		_w10249_
	);
	LUT2 #(
		.INIT('h8)
	) name6203 (
		\sport1_txctl_Wcnt_reg[1]/NET0131 ,
		_w7689_,
		_w10250_
	);
	LUT2 #(
		.INIT('h8)
	) name6204 (
		\memc_usysr_DO_reg[9]/NET0131 ,
		_w7301_,
		_w10251_
	);
	LUT2 #(
		.INIT('h8)
	) name6205 (
		\clkc_ckr_reg_DO_reg[9]/NET0131 ,
		_w7239_,
		_w10252_
	);
	LUT2 #(
		.INIT('h8)
	) name6206 (
		\sport1_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w7527_,
		_w10253_
	);
	LUT2 #(
		.INIT('h1)
	) name6207 (
		_w7522_,
		_w10232_,
		_w10254_
	);
	LUT2 #(
		.INIT('h1)
	) name6208 (
		_w10233_,
		_w10235_,
		_w10255_
	);
	LUT2 #(
		.INIT('h1)
	) name6209 (
		_w10238_,
		_w10240_,
		_w10256_
	);
	LUT2 #(
		.INIT('h1)
	) name6210 (
		_w10241_,
		_w10242_,
		_w10257_
	);
	LUT2 #(
		.INIT('h1)
	) name6211 (
		_w10243_,
		_w10244_,
		_w10258_
	);
	LUT2 #(
		.INIT('h1)
	) name6212 (
		_w10245_,
		_w10246_,
		_w10259_
	);
	LUT2 #(
		.INIT('h1)
	) name6213 (
		_w10247_,
		_w10251_,
		_w10260_
	);
	LUT2 #(
		.INIT('h1)
	) name6214 (
		_w10252_,
		_w10253_,
		_w10261_
	);
	LUT2 #(
		.INIT('h8)
	) name6215 (
		_w10260_,
		_w10261_,
		_w10262_
	);
	LUT2 #(
		.INIT('h8)
	) name6216 (
		_w10258_,
		_w10259_,
		_w10263_
	);
	LUT2 #(
		.INIT('h8)
	) name6217 (
		_w10256_,
		_w10257_,
		_w10264_
	);
	LUT2 #(
		.INIT('h8)
	) name6218 (
		_w10254_,
		_w10255_,
		_w10265_
	);
	LUT2 #(
		.INIT('h1)
	) name6219 (
		_w10249_,
		_w10250_,
		_w10266_
	);
	LUT2 #(
		.INIT('h8)
	) name6220 (
		_w10265_,
		_w10266_,
		_w10267_
	);
	LUT2 #(
		.INIT('h8)
	) name6221 (
		_w10263_,
		_w10264_,
		_w10268_
	);
	LUT2 #(
		.INIT('h8)
	) name6222 (
		_w10262_,
		_w10268_,
		_w10269_
	);
	LUT2 #(
		.INIT('h4)
	) name6223 (
		_w10234_,
		_w10267_,
		_w10270_
	);
	LUT2 #(
		.INIT('h1)
	) name6224 (
		_w10236_,
		_w10239_,
		_w10271_
	);
	LUT2 #(
		.INIT('h8)
	) name6225 (
		_w10270_,
		_w10271_,
		_w10272_
	);
	LUT2 #(
		.INIT('h4)
	) name6226 (
		_w10237_,
		_w10269_,
		_w10273_
	);
	LUT2 #(
		.INIT('h4)
	) name6227 (
		_w10248_,
		_w10273_,
		_w10274_
	);
	LUT2 #(
		.INIT('h8)
	) name6228 (
		_w10272_,
		_w10274_,
		_w10275_
	);
	LUT2 #(
		.INIT('h2)
	) name6229 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w10275_,
		_w10276_
	);
	LUT2 #(
		.INIT('h1)
	) name6230 (
		_w10148_,
		_w10205_,
		_w10277_
	);
	LUT2 #(
		.INIT('h4)
	) name6231 (
		_w10172_,
		_w10277_,
		_w10278_
	);
	LUT2 #(
		.INIT('h1)
	) name6232 (
		_w10124_,
		_w10197_,
		_w10279_
	);
	LUT2 #(
		.INIT('h4)
	) name6233 (
		_w10231_,
		_w10279_,
		_w10280_
	);
	LUT2 #(
		.INIT('h8)
	) name6234 (
		_w10278_,
		_w10280_,
		_w10281_
	);
	LUT2 #(
		.INIT('h4)
	) name6235 (
		_w10215_,
		_w10281_,
		_w10282_
	);
	LUT2 #(
		.INIT('h4)
	) name6236 (
		_w10276_,
		_w10282_,
		_w10283_
	);
	LUT2 #(
		.INIT('h4)
	) name6237 (
		_w10093_,
		_w10283_,
		_w10284_
	);
	LUT2 #(
		.INIT('h1)
	) name6238 (
		\emc_DMDoe_reg/NET0131 ,
		_w10284_,
		_w10285_
	);
	LUT2 #(
		.INIT('h8)
	) name6239 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[9]/P0001 ,
		_w10286_
	);
	LUT2 #(
		.INIT('h2)
	) name6240 (
		_w7057_,
		_w10286_,
		_w10287_
	);
	LUT2 #(
		.INIT('h4)
	) name6241 (
		_w10285_,
		_w10287_,
		_w10288_
	);
	LUT2 #(
		.INIT('h1)
	) name6242 (
		_w10092_,
		_w10288_,
		_w10289_
	);
	LUT2 #(
		.INIT('h1)
	) name6243 (
		_w6176_,
		_w10289_,
		_w10290_
	);
	LUT2 #(
		.INIT('h2)
	) name6244 (
		\core_dag_ilm1reg_I_reg[4]/NET0131 ,
		_w6280_,
		_w10291_
	);
	LUT2 #(
		.INIT('h1)
	) name6245 (
		_w6308_,
		_w6378_,
		_w10292_
	);
	LUT2 #(
		.INIT('h4)
	) name6246 (
		_w6372_,
		_w10292_,
		_w10293_
	);
	LUT2 #(
		.INIT('h2)
	) name6247 (
		_w6372_,
		_w10292_,
		_w10294_
	);
	LUT2 #(
		.INIT('h1)
	) name6248 (
		_w10293_,
		_w10294_,
		_w10295_
	);
	LUT2 #(
		.INIT('h4)
	) name6249 (
		_w7631_,
		_w10295_,
		_w10296_
	);
	LUT2 #(
		.INIT('h1)
	) name6250 (
		_w6304_,
		_w6505_,
		_w10297_
	);
	LUT2 #(
		.INIT('h8)
	) name6251 (
		_w6304_,
		_w6505_,
		_w10298_
	);
	LUT2 #(
		.INIT('h1)
	) name6252 (
		_w10297_,
		_w10298_,
		_w10299_
	);
	LUT2 #(
		.INIT('h8)
	) name6253 (
		_w7631_,
		_w10299_,
		_w10300_
	);
	LUT2 #(
		.INIT('h1)
	) name6254 (
		_w10291_,
		_w10296_,
		_w10301_
	);
	LUT2 #(
		.INIT('h4)
	) name6255 (
		_w10300_,
		_w10301_,
		_w10302_
	);
	LUT2 #(
		.INIT('h8)
	) name6256 (
		_w6176_,
		_w10302_,
		_w10303_
	);
	LUT2 #(
		.INIT('h1)
	) name6257 (
		_w6135_,
		_w10290_,
		_w10304_
	);
	LUT2 #(
		.INIT('h4)
	) name6258 (
		_w10303_,
		_w10304_,
		_w10305_
	);
	LUT2 #(
		.INIT('h2)
	) name6259 (
		_w7005_,
		_w10074_,
		_w10306_
	);
	LUT2 #(
		.INIT('h4)
	) name6260 (
		_w10305_,
		_w10306_,
		_w10307_
	);
	LUT2 #(
		.INIT('h1)
	) name6261 (
		_w9823_,
		_w10307_,
		_w10308_
	);
	LUT2 #(
		.INIT('h8)
	) name6262 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		_w6680_,
		_w10309_
	);
	LUT2 #(
		.INIT('h1)
	) name6263 (
		_w6675_,
		_w6690_,
		_w10310_
	);
	LUT2 #(
		.INIT('h1)
	) name6264 (
		_w6686_,
		_w10310_,
		_w10311_
	);
	LUT2 #(
		.INIT('h1)
	) name6265 (
		_w6759_,
		_w10311_,
		_w10312_
	);
	LUT2 #(
		.INIT('h8)
	) name6266 (
		_w6759_,
		_w10311_,
		_w10313_
	);
	LUT2 #(
		.INIT('h1)
	) name6267 (
		_w10312_,
		_w10313_,
		_w10314_
	);
	LUT2 #(
		.INIT('h4)
	) name6268 (
		_w8198_,
		_w10314_,
		_w10315_
	);
	LUT2 #(
		.INIT('h1)
	) name6269 (
		_w6763_,
		_w6764_,
		_w10316_
	);
	LUT2 #(
		.INIT('h1)
	) name6270 (
		_w6774_,
		_w6819_,
		_w10317_
	);
	LUT2 #(
		.INIT('h1)
	) name6271 (
		_w6820_,
		_w10317_,
		_w10318_
	);
	LUT2 #(
		.INIT('h1)
	) name6272 (
		_w10316_,
		_w10318_,
		_w10319_
	);
	LUT2 #(
		.INIT('h8)
	) name6273 (
		_w10316_,
		_w10318_,
		_w10320_
	);
	LUT2 #(
		.INIT('h1)
	) name6274 (
		_w10319_,
		_w10320_,
		_w10321_
	);
	LUT2 #(
		.INIT('h8)
	) name6275 (
		_w8198_,
		_w10321_,
		_w10322_
	);
	LUT2 #(
		.INIT('h1)
	) name6276 (
		_w10309_,
		_w10315_,
		_w10323_
	);
	LUT2 #(
		.INIT('h4)
	) name6277 (
		_w10322_,
		_w10323_,
		_w10324_
	);
	LUT2 #(
		.INIT('h4)
	) name6278 (
		_w6176_,
		_w10324_,
		_w10325_
	);
	LUT2 #(
		.INIT('h8)
	) name6279 (
		\core_dag_ilm1reg_I_reg[8]/NET0131 ,
		_w6401_,
		_w10326_
	);
	LUT2 #(
		.INIT('h4)
	) name6280 (
		_w6413_,
		_w6514_,
		_w10327_
	);
	LUT2 #(
		.INIT('h2)
	) name6281 (
		_w6413_,
		_w6514_,
		_w10328_
	);
	LUT2 #(
		.INIT('h1)
	) name6282 (
		_w10327_,
		_w10328_,
		_w10329_
	);
	LUT2 #(
		.INIT('h8)
	) name6283 (
		_w7612_,
		_w10329_,
		_w10330_
	);
	LUT2 #(
		.INIT('h1)
	) name6284 (
		_w6417_,
		_w6459_,
		_w10331_
	);
	LUT2 #(
		.INIT('h4)
	) name6285 (
		_w6385_,
		_w10331_,
		_w10332_
	);
	LUT2 #(
		.INIT('h2)
	) name6286 (
		_w6385_,
		_w10331_,
		_w10333_
	);
	LUT2 #(
		.INIT('h1)
	) name6287 (
		_w10332_,
		_w10333_,
		_w10334_
	);
	LUT2 #(
		.INIT('h1)
	) name6288 (
		_w7612_,
		_w10334_,
		_w10335_
	);
	LUT2 #(
		.INIT('h2)
	) name6289 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w10330_,
		_w10336_
	);
	LUT2 #(
		.INIT('h4)
	) name6290 (
		_w10335_,
		_w10336_,
		_w10337_
	);
	LUT2 #(
		.INIT('h4)
	) name6291 (
		_w6496_,
		_w10329_,
		_w10338_
	);
	LUT2 #(
		.INIT('h2)
	) name6292 (
		_w6496_,
		_w10334_,
		_w10339_
	);
	LUT2 #(
		.INIT('h1)
	) name6293 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w10338_,
		_w10340_
	);
	LUT2 #(
		.INIT('h4)
	) name6294 (
		_w10339_,
		_w10340_,
		_w10341_
	);
	LUT2 #(
		.INIT('h1)
	) name6295 (
		_w10326_,
		_w10337_,
		_w10342_
	);
	LUT2 #(
		.INIT('h4)
	) name6296 (
		_w10341_,
		_w10342_,
		_w10343_
	);
	LUT2 #(
		.INIT('h8)
	) name6297 (
		_w6176_,
		_w10343_,
		_w10344_
	);
	LUT2 #(
		.INIT('h1)
	) name6298 (
		_w10325_,
		_w10344_,
		_w10345_
	);
	LUT2 #(
		.INIT('h2)
	) name6299 (
		_w6135_,
		_w10345_,
		_w10346_
	);
	LUT2 #(
		.INIT('h1)
	) name6300 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w6924_,
		_w10347_
	);
	LUT2 #(
		.INIT('h8)
	) name6301 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w6926_,
		_w10348_
	);
	LUT2 #(
		.INIT('h8)
	) name6302 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131 ,
		_w6988_,
		_w10349_
	);
	LUT2 #(
		.INIT('h8)
	) name6303 (
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w6976_,
		_w10350_
	);
	LUT2 #(
		.INIT('h8)
	) name6304 (
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w6972_,
		_w10351_
	);
	LUT2 #(
		.INIT('h8)
	) name6305 (
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w6974_,
		_w10352_
	);
	LUT2 #(
		.INIT('h8)
	) name6306 (
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		_w6970_,
		_w10353_
	);
	LUT2 #(
		.INIT('h1)
	) name6307 (
		_w10350_,
		_w10351_,
		_w10354_
	);
	LUT2 #(
		.INIT('h1)
	) name6308 (
		_w10352_,
		_w10353_,
		_w10355_
	);
	LUT2 #(
		.INIT('h8)
	) name6309 (
		_w10354_,
		_w10355_,
		_w10356_
	);
	LUT2 #(
		.INIT('h2)
	) name6310 (
		_w4055_,
		_w10356_,
		_w10357_
	);
	LUT2 #(
		.INIT('h8)
	) name6311 (
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w6960_,
		_w10358_
	);
	LUT2 #(
		.INIT('h8)
	) name6312 (
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w6958_,
		_w10359_
	);
	LUT2 #(
		.INIT('h8)
	) name6313 (
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w6962_,
		_w10360_
	);
	LUT2 #(
		.INIT('h8)
	) name6314 (
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		_w6964_,
		_w10361_
	);
	LUT2 #(
		.INIT('h1)
	) name6315 (
		_w10358_,
		_w10359_,
		_w10362_
	);
	LUT2 #(
		.INIT('h1)
	) name6316 (
		_w10360_,
		_w10361_,
		_w10363_
	);
	LUT2 #(
		.INIT('h8)
	) name6317 (
		_w10362_,
		_w10363_,
		_w10364_
	);
	LUT2 #(
		.INIT('h4)
	) name6318 (
		_w10357_,
		_w10364_,
		_w10365_
	);
	LUT2 #(
		.INIT('h1)
	) name6319 (
		_w6121_,
		_w10365_,
		_w10366_
	);
	LUT2 #(
		.INIT('h8)
	) name6320 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w6956_,
		_w10367_
	);
	LUT2 #(
		.INIT('h8)
	) name6321 (
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		_w6142_,
		_w10368_
	);
	LUT2 #(
		.INIT('h8)
	) name6322 (
		\core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 ,
		_w6058_,
		_w10369_
	);
	LUT2 #(
		.INIT('h8)
	) name6323 (
		_w6060_,
		_w10369_,
		_w10370_
	);
	LUT2 #(
		.INIT('h8)
	) name6324 (
		\core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 ,
		_w6084_,
		_w10371_
	);
	LUT2 #(
		.INIT('h8)
	) name6325 (
		_w6085_,
		_w10371_,
		_w10372_
	);
	LUT2 #(
		.INIT('h8)
	) name6326 (
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w6140_,
		_w10373_
	);
	LUT2 #(
		.INIT('h1)
	) name6327 (
		_w4055_,
		_w10368_,
		_w10374_
	);
	LUT2 #(
		.INIT('h1)
	) name6328 (
		_w10370_,
		_w10372_,
		_w10375_
	);
	LUT2 #(
		.INIT('h4)
	) name6329 (
		_w10373_,
		_w10375_,
		_w10376_
	);
	LUT2 #(
		.INIT('h8)
	) name6330 (
		_w10374_,
		_w10376_,
		_w10377_
	);
	LUT2 #(
		.INIT('h8)
	) name6331 (
		_w6095_,
		_w10371_,
		_w10378_
	);
	LUT2 #(
		.INIT('h8)
	) name6332 (
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w6150_,
		_w10379_
	);
	LUT2 #(
		.INIT('h8)
	) name6333 (
		\core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 ,
		_w6148_,
		_w10380_
	);
	LUT2 #(
		.INIT('h8)
	) name6334 (
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		_w6154_,
		_w10381_
	);
	LUT2 #(
		.INIT('h1)
	) name6335 (
		_w10378_,
		_w10379_,
		_w10382_
	);
	LUT2 #(
		.INIT('h1)
	) name6336 (
		_w10380_,
		_w10381_,
		_w10383_
	);
	LUT2 #(
		.INIT('h8)
	) name6337 (
		_w10382_,
		_w10383_,
		_w10384_
	);
	LUT2 #(
		.INIT('h8)
	) name6338 (
		_w4055_,
		_w10384_,
		_w10385_
	);
	LUT2 #(
		.INIT('h1)
	) name6339 (
		_w10377_,
		_w10385_,
		_w10386_
	);
	LUT2 #(
		.INIT('h4)
	) name6340 (
		_w6111_,
		_w10386_,
		_w10387_
	);
	LUT2 #(
		.INIT('h1)
	) name6341 (
		_w10366_,
		_w10367_,
		_w10388_
	);
	LUT2 #(
		.INIT('h4)
	) name6342 (
		_w10387_,
		_w10388_,
		_w10389_
	);
	LUT2 #(
		.INIT('h2)
	) name6343 (
		_w5949_,
		_w10389_,
		_w10390_
	);
	LUT2 #(
		.INIT('h2)
	) name6344 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		_w6934_,
		_w10391_
	);
	LUT2 #(
		.INIT('h1)
	) name6345 (
		_w10348_,
		_w10349_,
		_w10392_
	);
	LUT2 #(
		.INIT('h8)
	) name6346 (
		_w6924_,
		_w10392_,
		_w10393_
	);
	LUT2 #(
		.INIT('h4)
	) name6347 (
		_w10391_,
		_w10393_,
		_w10394_
	);
	LUT2 #(
		.INIT('h4)
	) name6348 (
		_w10390_,
		_w10394_,
		_w10395_
	);
	LUT2 #(
		.INIT('h1)
	) name6349 (
		_w6176_,
		_w10347_,
		_w10396_
	);
	LUT2 #(
		.INIT('h4)
	) name6350 (
		_w10395_,
		_w10396_,
		_w10397_
	);
	LUT2 #(
		.INIT('h8)
	) name6351 (
		\core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 ,
		_w6084_,
		_w10398_
	);
	LUT2 #(
		.INIT('h8)
	) name6352 (
		_w6085_,
		_w10398_,
		_w10399_
	);
	LUT2 #(
		.INIT('h8)
	) name6353 (
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		_w6140_,
		_w10400_
	);
	LUT2 #(
		.INIT('h8)
	) name6354 (
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		_w8131_,
		_w10401_
	);
	LUT2 #(
		.INIT('h8)
	) name6355 (
		\core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 ,
		_w6067_,
		_w10402_
	);
	LUT2 #(
		.INIT('h8)
	) name6356 (
		_w6068_,
		_w10402_,
		_w10403_
	);
	LUT2 #(
		.INIT('h1)
	) name6357 (
		_w4055_,
		_w10399_,
		_w10404_
	);
	LUT2 #(
		.INIT('h1)
	) name6358 (
		_w10400_,
		_w10401_,
		_w10405_
	);
	LUT2 #(
		.INIT('h4)
	) name6359 (
		_w10403_,
		_w10405_,
		_w10406_
	);
	LUT2 #(
		.INIT('h8)
	) name6360 (
		_w10404_,
		_w10406_,
		_w10407_
	);
	LUT2 #(
		.INIT('h8)
	) name6361 (
		_w6091_,
		_w10402_,
		_w10408_
	);
	LUT2 #(
		.INIT('h8)
	) name6362 (
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		_w6150_,
		_w10409_
	);
	LUT2 #(
		.INIT('h8)
	) name6363 (
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		_w6148_,
		_w10410_
	);
	LUT2 #(
		.INIT('h8)
	) name6364 (
		\core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 ,
		_w6152_,
		_w10411_
	);
	LUT2 #(
		.INIT('h1)
	) name6365 (
		_w10408_,
		_w10409_,
		_w10412_
	);
	LUT2 #(
		.INIT('h1)
	) name6366 (
		_w10410_,
		_w10411_,
		_w10413_
	);
	LUT2 #(
		.INIT('h8)
	) name6367 (
		_w10412_,
		_w10413_,
		_w10414_
	);
	LUT2 #(
		.INIT('h8)
	) name6368 (
		_w4055_,
		_w10414_,
		_w10415_
	);
	LUT2 #(
		.INIT('h1)
	) name6369 (
		_w10407_,
		_w10415_,
		_w10416_
	);
	LUT2 #(
		.INIT('h8)
	) name6370 (
		_w6176_,
		_w10416_,
		_w10417_
	);
	LUT2 #(
		.INIT('h1)
	) name6371 (
		_w6135_,
		_w10417_,
		_w10418_
	);
	LUT2 #(
		.INIT('h4)
	) name6372 (
		_w10397_,
		_w10418_,
		_w10419_
	);
	LUT2 #(
		.INIT('h1)
	) name6373 (
		_w7005_,
		_w10419_,
		_w10420_
	);
	LUT2 #(
		.INIT('h4)
	) name6374 (
		_w10346_,
		_w10420_,
		_w10421_
	);
	LUT2 #(
		.INIT('h2)
	) name6375 (
		_w10365_,
		_w10386_,
		_w10422_
	);
	LUT2 #(
		.INIT('h2)
	) name6376 (
		_w8153_,
		_w10422_,
		_w10423_
	);
	LUT2 #(
		.INIT('h8)
	) name6377 (
		\DM_rdm[8]_pad ,
		_w7016_,
		_w10424_
	);
	LUT2 #(
		.INIT('h8)
	) name6378 (
		\DM_rd1[8]_pad ,
		_w7022_,
		_w10425_
	);
	LUT2 #(
		.INIT('h8)
	) name6379 (
		\DM_rd4[8]_pad ,
		_w7028_,
		_w10426_
	);
	LUT2 #(
		.INIT('h8)
	) name6380 (
		\DM_rd6[8]_pad ,
		_w7031_,
		_w10427_
	);
	LUT2 #(
		.INIT('h8)
	) name6381 (
		\DM_rd7[8]_pad ,
		_w7034_,
		_w10428_
	);
	LUT2 #(
		.INIT('h8)
	) name6382 (
		\DM_rd3[8]_pad ,
		_w7038_,
		_w10429_
	);
	LUT2 #(
		.INIT('h2)
	) name6383 (
		\DM_rd0[8]_pad ,
		_w7053_,
		_w10430_
	);
	LUT2 #(
		.INIT('h8)
	) name6384 (
		\DM_rd5[8]_pad ,
		_w7043_,
		_w10431_
	);
	LUT2 #(
		.INIT('h8)
	) name6385 (
		\DM_rd2[8]_pad ,
		_w7041_,
		_w10432_
	);
	LUT2 #(
		.INIT('h1)
	) name6386 (
		_w10425_,
		_w10429_,
		_w10433_
	);
	LUT2 #(
		.INIT('h4)
	) name6387 (
		_w10432_,
		_w10433_,
		_w10434_
	);
	LUT2 #(
		.INIT('h1)
	) name6388 (
		_w7057_,
		_w10424_,
		_w10435_
	);
	LUT2 #(
		.INIT('h1)
	) name6389 (
		_w10427_,
		_w10428_,
		_w10436_
	);
	LUT2 #(
		.INIT('h8)
	) name6390 (
		_w10435_,
		_w10436_,
		_w10437_
	);
	LUT2 #(
		.INIT('h4)
	) name6391 (
		_w10426_,
		_w10434_,
		_w10438_
	);
	LUT2 #(
		.INIT('h4)
	) name6392 (
		_w10431_,
		_w10438_,
		_w10439_
	);
	LUT2 #(
		.INIT('h8)
	) name6393 (
		_w10437_,
		_w10439_,
		_w10440_
	);
	LUT2 #(
		.INIT('h4)
	) name6394 (
		_w10430_,
		_w10440_,
		_w10441_
	);
	LUT2 #(
		.INIT('h8)
	) name6395 (
		\regout_STD_C_reg[8]/P0001 ,
		_w6988_,
		_w10442_
	);
	LUT2 #(
		.INIT('h4)
	) name6396 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001 ,
		_w10443_
	);
	LUT2 #(
		.INIT('h8)
	) name6397 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001 ,
		_w10444_
	);
	LUT2 #(
		.INIT('h1)
	) name6398 (
		_w10443_,
		_w10444_,
		_w10445_
	);
	LUT2 #(
		.INIT('h2)
	) name6399 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w10445_,
		_w10446_
	);
	LUT2 #(
		.INIT('h4)
	) name6400 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001 ,
		_w10447_
	);
	LUT2 #(
		.INIT('h8)
	) name6401 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001 ,
		_w10448_
	);
	LUT2 #(
		.INIT('h1)
	) name6402 (
		_w10447_,
		_w10448_,
		_w10449_
	);
	LUT2 #(
		.INIT('h2)
	) name6403 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w10449_,
		_w10450_
	);
	LUT2 #(
		.INIT('h4)
	) name6404 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001 ,
		_w10451_
	);
	LUT2 #(
		.INIT('h8)
	) name6405 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001 ,
		_w10452_
	);
	LUT2 #(
		.INIT('h1)
	) name6406 (
		_w10451_,
		_w10452_,
		_w10453_
	);
	LUT2 #(
		.INIT('h2)
	) name6407 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w10453_,
		_w10454_
	);
	LUT2 #(
		.INIT('h4)
	) name6408 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001 ,
		_w10455_
	);
	LUT2 #(
		.INIT('h8)
	) name6409 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001 ,
		_w10456_
	);
	LUT2 #(
		.INIT('h1)
	) name6410 (
		_w10455_,
		_w10456_,
		_w10457_
	);
	LUT2 #(
		.INIT('h2)
	) name6411 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w10457_,
		_w10458_
	);
	LUT2 #(
		.INIT('h4)
	) name6412 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001 ,
		_w10459_
	);
	LUT2 #(
		.INIT('h8)
	) name6413 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001 ,
		_w10460_
	);
	LUT2 #(
		.INIT('h1)
	) name6414 (
		_w10459_,
		_w10460_,
		_w10461_
	);
	LUT2 #(
		.INIT('h2)
	) name6415 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w10461_,
		_w10462_
	);
	LUT2 #(
		.INIT('h1)
	) name6416 (
		_w10446_,
		_w10450_,
		_w10463_
	);
	LUT2 #(
		.INIT('h1)
	) name6417 (
		_w10454_,
		_w10458_,
		_w10464_
	);
	LUT2 #(
		.INIT('h4)
	) name6418 (
		_w10462_,
		_w10464_,
		_w10465_
	);
	LUT2 #(
		.INIT('h8)
	) name6419 (
		_w10463_,
		_w10465_,
		_w10466_
	);
	LUT2 #(
		.INIT('h2)
	) name6420 (
		_w7093_,
		_w10466_,
		_w10467_
	);
	LUT2 #(
		.INIT('h8)
	) name6421 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w10468_
	);
	LUT2 #(
		.INIT('h8)
	) name6422 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131 ,
		_w10469_
	);
	LUT2 #(
		.INIT('h8)
	) name6423 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 ,
		_w10470_
	);
	LUT2 #(
		.INIT('h8)
	) name6424 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 ,
		_w10471_
	);
	LUT2 #(
		.INIT('h8)
	) name6425 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131 ,
		_w10472_
	);
	LUT2 #(
		.INIT('h8)
	) name6426 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131 ,
		_w10473_
	);
	LUT2 #(
		.INIT('h8)
	) name6427 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131 ,
		_w10474_
	);
	LUT2 #(
		.INIT('h8)
	) name6428 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		_w10475_
	);
	LUT2 #(
		.INIT('h8)
	) name6429 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131 ,
		_w10476_
	);
	LUT2 #(
		.INIT('h8)
	) name6430 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131 ,
		_w10477_
	);
	LUT2 #(
		.INIT('h8)
	) name6431 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131 ,
		_w10478_
	);
	LUT2 #(
		.INIT('h8)
	) name6432 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131 ,
		_w10479_
	);
	LUT2 #(
		.INIT('h1)
	) name6433 (
		_w10468_,
		_w10469_,
		_w10480_
	);
	LUT2 #(
		.INIT('h1)
	) name6434 (
		_w10470_,
		_w10471_,
		_w10481_
	);
	LUT2 #(
		.INIT('h1)
	) name6435 (
		_w10472_,
		_w10473_,
		_w10482_
	);
	LUT2 #(
		.INIT('h1)
	) name6436 (
		_w10474_,
		_w10475_,
		_w10483_
	);
	LUT2 #(
		.INIT('h1)
	) name6437 (
		_w10476_,
		_w10477_,
		_w10484_
	);
	LUT2 #(
		.INIT('h1)
	) name6438 (
		_w10478_,
		_w10479_,
		_w10485_
	);
	LUT2 #(
		.INIT('h8)
	) name6439 (
		_w10484_,
		_w10485_,
		_w10486_
	);
	LUT2 #(
		.INIT('h8)
	) name6440 (
		_w10482_,
		_w10483_,
		_w10487_
	);
	LUT2 #(
		.INIT('h8)
	) name6441 (
		_w10480_,
		_w10481_,
		_w10488_
	);
	LUT2 #(
		.INIT('h8)
	) name6442 (
		_w10487_,
		_w10488_,
		_w10489_
	);
	LUT2 #(
		.INIT('h8)
	) name6443 (
		_w10486_,
		_w10489_,
		_w10490_
	);
	LUT2 #(
		.INIT('h2)
	) name6444 (
		_w7128_,
		_w10490_,
		_w10491_
	);
	LUT2 #(
		.INIT('h8)
	) name6445 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131 ,
		_w10492_
	);
	LUT2 #(
		.INIT('h8)
	) name6446 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131 ,
		_w10493_
	);
	LUT2 #(
		.INIT('h8)
	) name6447 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131 ,
		_w10494_
	);
	LUT2 #(
		.INIT('h8)
	) name6448 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		_w10495_
	);
	LUT2 #(
		.INIT('h8)
	) name6449 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		_w10496_
	);
	LUT2 #(
		.INIT('h8)
	) name6450 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131 ,
		_w10497_
	);
	LUT2 #(
		.INIT('h8)
	) name6451 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131 ,
		_w10498_
	);
	LUT2 #(
		.INIT('h8)
	) name6452 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131 ,
		_w10499_
	);
	LUT2 #(
		.INIT('h8)
	) name6453 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131 ,
		_w10500_
	);
	LUT2 #(
		.INIT('h8)
	) name6454 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[8]/NET0131 ,
		_w10501_
	);
	LUT2 #(
		.INIT('h8)
	) name6455 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[8]/NET0131 ,
		_w10502_
	);
	LUT2 #(
		.INIT('h8)
	) name6456 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131 ,
		_w10503_
	);
	LUT2 #(
		.INIT('h1)
	) name6457 (
		_w10492_,
		_w10493_,
		_w10504_
	);
	LUT2 #(
		.INIT('h1)
	) name6458 (
		_w10494_,
		_w10495_,
		_w10505_
	);
	LUT2 #(
		.INIT('h1)
	) name6459 (
		_w10496_,
		_w10497_,
		_w10506_
	);
	LUT2 #(
		.INIT('h1)
	) name6460 (
		_w10498_,
		_w10499_,
		_w10507_
	);
	LUT2 #(
		.INIT('h1)
	) name6461 (
		_w10500_,
		_w10501_,
		_w10508_
	);
	LUT2 #(
		.INIT('h1)
	) name6462 (
		_w10502_,
		_w10503_,
		_w10509_
	);
	LUT2 #(
		.INIT('h8)
	) name6463 (
		_w10508_,
		_w10509_,
		_w10510_
	);
	LUT2 #(
		.INIT('h8)
	) name6464 (
		_w10506_,
		_w10507_,
		_w10511_
	);
	LUT2 #(
		.INIT('h8)
	) name6465 (
		_w10504_,
		_w10505_,
		_w10512_
	);
	LUT2 #(
		.INIT('h8)
	) name6466 (
		_w10511_,
		_w10512_,
		_w10513_
	);
	LUT2 #(
		.INIT('h8)
	) name6467 (
		_w10510_,
		_w10513_,
		_w10514_
	);
	LUT2 #(
		.INIT('h2)
	) name6468 (
		_w7068_,
		_w10514_,
		_w10515_
	);
	LUT2 #(
		.INIT('h4)
	) name6469 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001 ,
		_w10516_
	);
	LUT2 #(
		.INIT('h8)
	) name6470 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001 ,
		_w10517_
	);
	LUT2 #(
		.INIT('h1)
	) name6471 (
		_w10516_,
		_w10517_,
		_w10518_
	);
	LUT2 #(
		.INIT('h2)
	) name6472 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w10518_,
		_w10519_
	);
	LUT2 #(
		.INIT('h4)
	) name6473 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001 ,
		_w10520_
	);
	LUT2 #(
		.INIT('h8)
	) name6474 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001 ,
		_w10521_
	);
	LUT2 #(
		.INIT('h1)
	) name6475 (
		_w10520_,
		_w10521_,
		_w10522_
	);
	LUT2 #(
		.INIT('h2)
	) name6476 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w10522_,
		_w10523_
	);
	LUT2 #(
		.INIT('h4)
	) name6477 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001 ,
		_w10524_
	);
	LUT2 #(
		.INIT('h8)
	) name6478 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001 ,
		_w10525_
	);
	LUT2 #(
		.INIT('h1)
	) name6479 (
		_w10524_,
		_w10525_,
		_w10526_
	);
	LUT2 #(
		.INIT('h2)
	) name6480 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w10526_,
		_w10527_
	);
	LUT2 #(
		.INIT('h4)
	) name6481 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001 ,
		_w10528_
	);
	LUT2 #(
		.INIT('h8)
	) name6482 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001 ,
		_w10529_
	);
	LUT2 #(
		.INIT('h1)
	) name6483 (
		_w10528_,
		_w10529_,
		_w10530_
	);
	LUT2 #(
		.INIT('h2)
	) name6484 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w10530_,
		_w10531_
	);
	LUT2 #(
		.INIT('h4)
	) name6485 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001 ,
		_w10532_
	);
	LUT2 #(
		.INIT('h8)
	) name6486 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 ,
		_w10533_
	);
	LUT2 #(
		.INIT('h1)
	) name6487 (
		_w10532_,
		_w10533_,
		_w10534_
	);
	LUT2 #(
		.INIT('h2)
	) name6488 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w10534_,
		_w10535_
	);
	LUT2 #(
		.INIT('h4)
	) name6489 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001 ,
		_w10536_
	);
	LUT2 #(
		.INIT('h8)
	) name6490 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 ,
		_w10537_
	);
	LUT2 #(
		.INIT('h1)
	) name6491 (
		_w10536_,
		_w10537_,
		_w10538_
	);
	LUT2 #(
		.INIT('h2)
	) name6492 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w10538_,
		_w10539_
	);
	LUT2 #(
		.INIT('h1)
	) name6493 (
		_w7207_,
		_w10519_,
		_w10540_
	);
	LUT2 #(
		.INIT('h1)
	) name6494 (
		_w10523_,
		_w10527_,
		_w10541_
	);
	LUT2 #(
		.INIT('h1)
	) name6495 (
		_w10531_,
		_w10535_,
		_w10542_
	);
	LUT2 #(
		.INIT('h4)
	) name6496 (
		_w10539_,
		_w10542_,
		_w10543_
	);
	LUT2 #(
		.INIT('h8)
	) name6497 (
		_w10540_,
		_w10541_,
		_w10544_
	);
	LUT2 #(
		.INIT('h8)
	) name6498 (
		_w10543_,
		_w10544_,
		_w10545_
	);
	LUT2 #(
		.INIT('h2)
	) name6499 (
		_w7179_,
		_w10545_,
		_w10546_
	);
	LUT2 #(
		.INIT('h8)
	) name6500 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[8]/P0001 ,
		_w10547_
	);
	LUT2 #(
		.INIT('h8)
	) name6501 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w10548_
	);
	LUT2 #(
		.INIT('h8)
	) name6502 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[8]/P0001 ,
		_w10549_
	);
	LUT2 #(
		.INIT('h8)
	) name6503 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[8]/P0001 ,
		_w10550_
	);
	LUT2 #(
		.INIT('h1)
	) name6504 (
		_w10547_,
		_w10548_,
		_w10551_
	);
	LUT2 #(
		.INIT('h1)
	) name6505 (
		_w10549_,
		_w10550_,
		_w10552_
	);
	LUT2 #(
		.INIT('h8)
	) name6506 (
		_w10551_,
		_w10552_,
		_w10553_
	);
	LUT2 #(
		.INIT('h2)
	) name6507 (
		_w7119_,
		_w10553_,
		_w10554_
	);
	LUT2 #(
		.INIT('h8)
	) name6508 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w10555_
	);
	LUT2 #(
		.INIT('h2)
	) name6509 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4425_,
		_w10556_
	);
	LUT2 #(
		.INIT('h8)
	) name6510 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w10557_
	);
	LUT2 #(
		.INIT('h2)
	) name6511 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w7216_,
		_w10558_
	);
	LUT2 #(
		.INIT('h8)
	) name6512 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w10559_
	);
	LUT2 #(
		.INIT('h1)
	) name6513 (
		_w10555_,
		_w10557_,
		_w10560_
	);
	LUT2 #(
		.INIT('h4)
	) name6514 (
		_w10559_,
		_w10560_,
		_w10561_
	);
	LUT2 #(
		.INIT('h4)
	) name6515 (
		_w10558_,
		_w10561_,
		_w10562_
	);
	LUT2 #(
		.INIT('h4)
	) name6516 (
		_w10556_,
		_w10562_,
		_w10563_
	);
	LUT2 #(
		.INIT('h2)
	) name6517 (
		_w7215_,
		_w10563_,
		_w10564_
	);
	LUT2 #(
		.INIT('h4)
	) name6518 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 ,
		_w10565_
	);
	LUT2 #(
		.INIT('h8)
	) name6519 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 ,
		_w10566_
	);
	LUT2 #(
		.INIT('h1)
	) name6520 (
		_w10565_,
		_w10566_,
		_w10567_
	);
	LUT2 #(
		.INIT('h2)
	) name6521 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w10567_,
		_w10568_
	);
	LUT2 #(
		.INIT('h4)
	) name6522 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001 ,
		_w10569_
	);
	LUT2 #(
		.INIT('h8)
	) name6523 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001 ,
		_w10570_
	);
	LUT2 #(
		.INIT('h1)
	) name6524 (
		_w10569_,
		_w10570_,
		_w10571_
	);
	LUT2 #(
		.INIT('h2)
	) name6525 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w10571_,
		_w10572_
	);
	LUT2 #(
		.INIT('h4)
	) name6526 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 ,
		_w10573_
	);
	LUT2 #(
		.INIT('h8)
	) name6527 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 ,
		_w10574_
	);
	LUT2 #(
		.INIT('h1)
	) name6528 (
		_w10573_,
		_w10574_,
		_w10575_
	);
	LUT2 #(
		.INIT('h2)
	) name6529 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w10575_,
		_w10576_
	);
	LUT2 #(
		.INIT('h1)
	) name6530 (
		_w10568_,
		_w10572_,
		_w10577_
	);
	LUT2 #(
		.INIT('h4)
	) name6531 (
		_w10576_,
		_w10577_,
		_w10578_
	);
	LUT2 #(
		.INIT('h8)
	) name6532 (
		_w7174_,
		_w10578_,
		_w10579_
	);
	LUT2 #(
		.INIT('h2)
	) name6533 (
		_w7153_,
		_w10579_,
		_w10580_
	);
	LUT2 #(
		.INIT('h8)
	) name6534 (
		\tm_tpr_reg_DO_reg[8]/NET0131 ,
		_w7293_,
		_w10581_
	);
	LUT2 #(
		.INIT('h8)
	) name6535 (
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w7273_,
		_w10582_
	);
	LUT2 #(
		.INIT('h8)
	) name6536 (
		\bdma_BCTL_reg[8]/NET0131 ,
		_w7230_,
		_w10583_
	);
	LUT2 #(
		.INIT('h8)
	) name6537 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w7299_,
		_w10584_
	);
	LUT2 #(
		.INIT('h8)
	) name6538 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w7234_,
		_w10585_
	);
	LUT2 #(
		.INIT('h8)
	) name6539 (
		\bdma_BOVL_reg[8]/NET0131 ,
		_w7534_,
		_w10586_
	);
	LUT2 #(
		.INIT('h8)
	) name6540 (
		\idma_DOVL_reg[8]/NET0131 ,
		_w7532_,
		_w10587_
	);
	LUT2 #(
		.INIT('h8)
	) name6541 (
		\bdma_BEAD_reg[8]/NET0131 ,
		_w7303_,
		_w10588_
	);
	LUT2 #(
		.INIT('h8)
	) name6542 (
		\IRFS0_pad ,
		_w7249_,
		_w10589_
	);
	LUT2 #(
		.INIT('h8)
	) name6543 (
		\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w7256_,
		_w10590_
	);
	LUT2 #(
		.INIT('h8)
	) name6544 (
		\tm_TCR_TMP_reg[8]/NET0131 ,
		_w7289_,
		_w10591_
	);
	LUT2 #(
		.INIT('h8)
	) name6545 (
		\sport0_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w7295_,
		_w10592_
	);
	LUT2 #(
		.INIT('h8)
	) name6546 (
		\emc_WSCRreg_DO_reg[8]/NET0131 ,
		_w7251_,
		_w10593_
	);
	LUT2 #(
		.INIT('h8)
	) name6547 (
		\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w7247_,
		_w10594_
	);
	LUT2 #(
		.INIT('h8)
	) name6548 (
		\sport1_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w7527_,
		_w10595_
	);
	LUT2 #(
		.INIT('h8)
	) name6549 (
		\IRFS1_pad ,
		_w7281_,
		_w10596_
	);
	LUT2 #(
		.INIT('h8)
	) name6550 (
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		_w7287_,
		_w10597_
	);
	LUT2 #(
		.INIT('h8)
	) name6551 (
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		_w7689_,
		_w10598_
	);
	LUT2 #(
		.INIT('h8)
	) name6552 (
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		_w7710_,
		_w10599_
	);
	LUT2 #(
		.INIT('h8)
	) name6553 (
		\memc_usysr_DO_reg[8]/NET0131 ,
		_w7301_,
		_w10600_
	);
	LUT2 #(
		.INIT('h8)
	) name6554 (
		\clkc_ckr_reg_DO_reg[8]/NET0131 ,
		_w7239_,
		_w10601_
	);
	LUT2 #(
		.INIT('h8)
	) name6555 (
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w7259_,
		_w10602_
	);
	LUT2 #(
		.INIT('h1)
	) name6556 (
		_w7522_,
		_w10581_,
		_w10603_
	);
	LUT2 #(
		.INIT('h1)
	) name6557 (
		_w10582_,
		_w10584_,
		_w10604_
	);
	LUT2 #(
		.INIT('h1)
	) name6558 (
		_w10587_,
		_w10589_,
		_w10605_
	);
	LUT2 #(
		.INIT('h1)
	) name6559 (
		_w10590_,
		_w10591_,
		_w10606_
	);
	LUT2 #(
		.INIT('h1)
	) name6560 (
		_w10592_,
		_w10593_,
		_w10607_
	);
	LUT2 #(
		.INIT('h1)
	) name6561 (
		_w10594_,
		_w10595_,
		_w10608_
	);
	LUT2 #(
		.INIT('h1)
	) name6562 (
		_w10596_,
		_w10600_,
		_w10609_
	);
	LUT2 #(
		.INIT('h1)
	) name6563 (
		_w10601_,
		_w10602_,
		_w10610_
	);
	LUT2 #(
		.INIT('h8)
	) name6564 (
		_w10609_,
		_w10610_,
		_w10611_
	);
	LUT2 #(
		.INIT('h8)
	) name6565 (
		_w10607_,
		_w10608_,
		_w10612_
	);
	LUT2 #(
		.INIT('h8)
	) name6566 (
		_w10605_,
		_w10606_,
		_w10613_
	);
	LUT2 #(
		.INIT('h8)
	) name6567 (
		_w10603_,
		_w10604_,
		_w10614_
	);
	LUT2 #(
		.INIT('h1)
	) name6568 (
		_w10598_,
		_w10599_,
		_w10615_
	);
	LUT2 #(
		.INIT('h8)
	) name6569 (
		_w10614_,
		_w10615_,
		_w10616_
	);
	LUT2 #(
		.INIT('h8)
	) name6570 (
		_w10612_,
		_w10613_,
		_w10617_
	);
	LUT2 #(
		.INIT('h8)
	) name6571 (
		_w10611_,
		_w10617_,
		_w10618_
	);
	LUT2 #(
		.INIT('h4)
	) name6572 (
		_w10583_,
		_w10616_,
		_w10619_
	);
	LUT2 #(
		.INIT('h1)
	) name6573 (
		_w10585_,
		_w10588_,
		_w10620_
	);
	LUT2 #(
		.INIT('h8)
	) name6574 (
		_w10619_,
		_w10620_,
		_w10621_
	);
	LUT2 #(
		.INIT('h4)
	) name6575 (
		_w10586_,
		_w10618_,
		_w10622_
	);
	LUT2 #(
		.INIT('h4)
	) name6576 (
		_w10597_,
		_w10622_,
		_w10623_
	);
	LUT2 #(
		.INIT('h8)
	) name6577 (
		_w10621_,
		_w10623_,
		_w10624_
	);
	LUT2 #(
		.INIT('h2)
	) name6578 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w10624_,
		_w10625_
	);
	LUT2 #(
		.INIT('h1)
	) name6579 (
		_w10491_,
		_w10554_,
		_w10626_
	);
	LUT2 #(
		.INIT('h4)
	) name6580 (
		_w10515_,
		_w10626_,
		_w10627_
	);
	LUT2 #(
		.INIT('h1)
	) name6581 (
		_w10467_,
		_w10546_,
		_w10628_
	);
	LUT2 #(
		.INIT('h4)
	) name6582 (
		_w10580_,
		_w10628_,
		_w10629_
	);
	LUT2 #(
		.INIT('h8)
	) name6583 (
		_w10627_,
		_w10629_,
		_w10630_
	);
	LUT2 #(
		.INIT('h4)
	) name6584 (
		_w10564_,
		_w10630_,
		_w10631_
	);
	LUT2 #(
		.INIT('h4)
	) name6585 (
		_w10625_,
		_w10631_,
		_w10632_
	);
	LUT2 #(
		.INIT('h4)
	) name6586 (
		_w10442_,
		_w10632_,
		_w10633_
	);
	LUT2 #(
		.INIT('h1)
	) name6587 (
		\emc_DMDoe_reg/NET0131 ,
		_w10633_,
		_w10634_
	);
	LUT2 #(
		.INIT('h8)
	) name6588 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[8]/P0001 ,
		_w10635_
	);
	LUT2 #(
		.INIT('h2)
	) name6589 (
		_w7057_,
		_w10635_,
		_w10636_
	);
	LUT2 #(
		.INIT('h4)
	) name6590 (
		_w10634_,
		_w10636_,
		_w10637_
	);
	LUT2 #(
		.INIT('h1)
	) name6591 (
		_w10441_,
		_w10637_,
		_w10638_
	);
	LUT2 #(
		.INIT('h8)
	) name6592 (
		_w7863_,
		_w10638_,
		_w10639_
	);
	LUT2 #(
		.INIT('h1)
	) name6593 (
		_w10423_,
		_w10639_,
		_w10640_
	);
	LUT2 #(
		.INIT('h2)
	) name6594 (
		_w7005_,
		_w10640_,
		_w10641_
	);
	LUT2 #(
		.INIT('h2)
	) name6595 (
		\core_dag_ilm1reg_I_reg[5]/NET0131 ,
		_w6251_,
		_w10642_
	);
	LUT2 #(
		.INIT('h1)
	) name6596 (
		_w6293_,
		_w6377_,
		_w10643_
	);
	LUT2 #(
		.INIT('h1)
	) name6597 (
		_w6308_,
		_w6372_,
		_w10644_
	);
	LUT2 #(
		.INIT('h1)
	) name6598 (
		_w6378_,
		_w10644_,
		_w10645_
	);
	LUT2 #(
		.INIT('h8)
	) name6599 (
		_w10643_,
		_w10645_,
		_w10646_
	);
	LUT2 #(
		.INIT('h1)
	) name6600 (
		_w10643_,
		_w10645_,
		_w10647_
	);
	LUT2 #(
		.INIT('h1)
	) name6601 (
		_w10646_,
		_w10647_,
		_w10648_
	);
	LUT2 #(
		.INIT('h4)
	) name6602 (
		_w7612_,
		_w10648_,
		_w10649_
	);
	LUT2 #(
		.INIT('h1)
	) name6603 (
		_w6282_,
		_w6505_,
		_w10650_
	);
	LUT2 #(
		.INIT('h1)
	) name6604 (
		_w6283_,
		_w10650_,
		_w10651_
	);
	LUT2 #(
		.INIT('h4)
	) name6605 (
		_w6289_,
		_w10651_,
		_w10652_
	);
	LUT2 #(
		.INIT('h2)
	) name6606 (
		_w6289_,
		_w10651_,
		_w10653_
	);
	LUT2 #(
		.INIT('h1)
	) name6607 (
		_w10652_,
		_w10653_,
		_w10654_
	);
	LUT2 #(
		.INIT('h8)
	) name6608 (
		_w7612_,
		_w10654_,
		_w10655_
	);
	LUT2 #(
		.INIT('h2)
	) name6609 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w10649_,
		_w10656_
	);
	LUT2 #(
		.INIT('h4)
	) name6610 (
		_w10655_,
		_w10656_,
		_w10657_
	);
	LUT2 #(
		.INIT('h8)
	) name6611 (
		_w6496_,
		_w10648_,
		_w10658_
	);
	LUT2 #(
		.INIT('h4)
	) name6612 (
		_w6496_,
		_w10654_,
		_w10659_
	);
	LUT2 #(
		.INIT('h1)
	) name6613 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w10658_,
		_w10660_
	);
	LUT2 #(
		.INIT('h4)
	) name6614 (
		_w10659_,
		_w10660_,
		_w10661_
	);
	LUT2 #(
		.INIT('h1)
	) name6615 (
		_w10642_,
		_w10657_,
		_w10662_
	);
	LUT2 #(
		.INIT('h4)
	) name6616 (
		_w10661_,
		_w10662_,
		_w10663_
	);
	LUT2 #(
		.INIT('h4)
	) name6617 (
		_w6135_,
		_w10663_,
		_w10664_
	);
	LUT2 #(
		.INIT('h8)
	) name6618 (
		\DM_rdm[5]_pad ,
		_w7016_,
		_w10665_
	);
	LUT2 #(
		.INIT('h8)
	) name6619 (
		\DM_rd1[5]_pad ,
		_w7022_,
		_w10666_
	);
	LUT2 #(
		.INIT('h8)
	) name6620 (
		\DM_rd4[5]_pad ,
		_w7028_,
		_w10667_
	);
	LUT2 #(
		.INIT('h8)
	) name6621 (
		\DM_rd6[5]_pad ,
		_w7031_,
		_w10668_
	);
	LUT2 #(
		.INIT('h8)
	) name6622 (
		\DM_rd7[5]_pad ,
		_w7034_,
		_w10669_
	);
	LUT2 #(
		.INIT('h8)
	) name6623 (
		\DM_rd3[5]_pad ,
		_w7038_,
		_w10670_
	);
	LUT2 #(
		.INIT('h2)
	) name6624 (
		\DM_rd0[5]_pad ,
		_w7053_,
		_w10671_
	);
	LUT2 #(
		.INIT('h8)
	) name6625 (
		\DM_rd5[5]_pad ,
		_w7043_,
		_w10672_
	);
	LUT2 #(
		.INIT('h8)
	) name6626 (
		\DM_rd2[5]_pad ,
		_w7041_,
		_w10673_
	);
	LUT2 #(
		.INIT('h1)
	) name6627 (
		_w10666_,
		_w10670_,
		_w10674_
	);
	LUT2 #(
		.INIT('h4)
	) name6628 (
		_w10673_,
		_w10674_,
		_w10675_
	);
	LUT2 #(
		.INIT('h1)
	) name6629 (
		_w7057_,
		_w10665_,
		_w10676_
	);
	LUT2 #(
		.INIT('h1)
	) name6630 (
		_w10668_,
		_w10669_,
		_w10677_
	);
	LUT2 #(
		.INIT('h8)
	) name6631 (
		_w10676_,
		_w10677_,
		_w10678_
	);
	LUT2 #(
		.INIT('h4)
	) name6632 (
		_w10667_,
		_w10675_,
		_w10679_
	);
	LUT2 #(
		.INIT('h4)
	) name6633 (
		_w10672_,
		_w10679_,
		_w10680_
	);
	LUT2 #(
		.INIT('h8)
	) name6634 (
		_w10678_,
		_w10680_,
		_w10681_
	);
	LUT2 #(
		.INIT('h4)
	) name6635 (
		_w10671_,
		_w10681_,
		_w10682_
	);
	LUT2 #(
		.INIT('h8)
	) name6636 (
		\regout_STD_C_reg[5]/P0001 ,
		_w6988_,
		_w10683_
	);
	LUT2 #(
		.INIT('h4)
	) name6637 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001 ,
		_w10684_
	);
	LUT2 #(
		.INIT('h8)
	) name6638 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001 ,
		_w10685_
	);
	LUT2 #(
		.INIT('h1)
	) name6639 (
		_w10684_,
		_w10685_,
		_w10686_
	);
	LUT2 #(
		.INIT('h2)
	) name6640 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w10686_,
		_w10687_
	);
	LUT2 #(
		.INIT('h4)
	) name6641 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001 ,
		_w10688_
	);
	LUT2 #(
		.INIT('h8)
	) name6642 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001 ,
		_w10689_
	);
	LUT2 #(
		.INIT('h1)
	) name6643 (
		_w10688_,
		_w10689_,
		_w10690_
	);
	LUT2 #(
		.INIT('h2)
	) name6644 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w10690_,
		_w10691_
	);
	LUT2 #(
		.INIT('h4)
	) name6645 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001 ,
		_w10692_
	);
	LUT2 #(
		.INIT('h8)
	) name6646 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001 ,
		_w10693_
	);
	LUT2 #(
		.INIT('h1)
	) name6647 (
		_w10692_,
		_w10693_,
		_w10694_
	);
	LUT2 #(
		.INIT('h2)
	) name6648 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w10694_,
		_w10695_
	);
	LUT2 #(
		.INIT('h4)
	) name6649 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001 ,
		_w10696_
	);
	LUT2 #(
		.INIT('h8)
	) name6650 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001 ,
		_w10697_
	);
	LUT2 #(
		.INIT('h1)
	) name6651 (
		_w10696_,
		_w10697_,
		_w10698_
	);
	LUT2 #(
		.INIT('h2)
	) name6652 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w10698_,
		_w10699_
	);
	LUT2 #(
		.INIT('h4)
	) name6653 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001 ,
		_w10700_
	);
	LUT2 #(
		.INIT('h8)
	) name6654 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001 ,
		_w10701_
	);
	LUT2 #(
		.INIT('h1)
	) name6655 (
		_w10700_,
		_w10701_,
		_w10702_
	);
	LUT2 #(
		.INIT('h2)
	) name6656 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w10702_,
		_w10703_
	);
	LUT2 #(
		.INIT('h8)
	) name6657 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w10704_
	);
	LUT2 #(
		.INIT('h1)
	) name6658 (
		_w10687_,
		_w10704_,
		_w10705_
	);
	LUT2 #(
		.INIT('h1)
	) name6659 (
		_w10691_,
		_w10695_,
		_w10706_
	);
	LUT2 #(
		.INIT('h1)
	) name6660 (
		_w10699_,
		_w10703_,
		_w10707_
	);
	LUT2 #(
		.INIT('h8)
	) name6661 (
		_w10706_,
		_w10707_,
		_w10708_
	);
	LUT2 #(
		.INIT('h8)
	) name6662 (
		_w10705_,
		_w10708_,
		_w10709_
	);
	LUT2 #(
		.INIT('h2)
	) name6663 (
		_w7093_,
		_w10709_,
		_w10710_
	);
	LUT2 #(
		.INIT('h8)
	) name6664 (
		\idma_DOVL_reg[5]/NET0131 ,
		_w7532_,
		_w10711_
	);
	LUT2 #(
		.INIT('h8)
	) name6665 (
		\sport0_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w7295_,
		_w10712_
	);
	LUT2 #(
		.INIT('h8)
	) name6666 (
		\tm_tpr_reg_DO_reg[5]/NET0131 ,
		_w7293_,
		_w10713_
	);
	LUT2 #(
		.INIT('h4)
	) name6667 (
		\bdma_BDMA_boot_reg/NET0131_reg_syn_10 ,
		\bdma_BWCOUNT_reg[5]/NET0131_reg_syn_2 ,
		_w10714_
	);
	LUT2 #(
		.INIT('h8)
	) name6668 (
		\bdma_BDMA_boot_reg/NET0131_reg_syn_10 ,
		\bdma_BWCOUNT_reg[5]/NET0131_reg_syn_8 ,
		_w10715_
	);
	LUT2 #(
		.INIT('h1)
	) name6669 (
		_w10714_,
		_w10715_,
		_w10716_
	);
	LUT2 #(
		.INIT('h2)
	) name6670 (
		_w7287_,
		_w10716_,
		_w10717_
	);
	LUT2 #(
		.INIT('h8)
	) name6671 (
		\emc_WSCRreg_DO_reg[5]/NET0131 ,
		_w7251_,
		_w10718_
	);
	LUT2 #(
		.INIT('h8)
	) name6672 (
		\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w7256_,
		_w10719_
	);
	LUT2 #(
		.INIT('h8)
	) name6673 (
		\sport1_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w7263_,
		_w10720_
	);
	LUT2 #(
		.INIT('h8)
	) name6674 (
		\tm_tsr_reg_DO_reg[5]/NET0131 ,
		_w7540_,
		_w10721_
	);
	LUT2 #(
		.INIT('h8)
	) name6675 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w7249_,
		_w10722_
	);
	LUT2 #(
		.INIT('h8)
	) name6676 (
		\emc_WSCRext_reg_DO_reg[5]/NET0131 ,
		_w7514_,
		_w10723_
	);
	LUT2 #(
		.INIT('h8)
	) name6677 (
		\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w7247_,
		_w10724_
	);
	LUT2 #(
		.INIT('h8)
	) name6678 (
		\sport1_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w7281_,
		_w10725_
	);
	LUT2 #(
		.INIT('h8)
	) name6679 (
		\pio_pmask_reg_DO_reg[5]/NET0131 ,
		_w7297_,
		_w10726_
	);
	LUT2 #(
		.INIT('h8)
	) name6680 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w7234_,
		_w10727_
	);
	LUT2 #(
		.INIT('h8)
	) name6681 (
		\sport0_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w7276_,
		_w10728_
	);
	LUT2 #(
		.INIT('h8)
	) name6682 (
		\sport1_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w7527_,
		_w10729_
	);
	LUT2 #(
		.INIT('h8)
	) name6683 (
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w7289_,
		_w10730_
	);
	LUT2 #(
		.INIT('h8)
	) name6684 (
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w7259_,
		_w10731_
	);
	LUT2 #(
		.INIT('h8)
	) name6685 (
		\bdma_BOVL_reg[5]/NET0131 ,
		_w7534_,
		_w10732_
	);
	LUT2 #(
		.INIT('h8)
	) name6686 (
		\clkc_ckr_reg_DO_reg[5]/NET0131 ,
		_w7239_,
		_w10733_
	);
	LUT2 #(
		.INIT('h8)
	) name6687 (
		\memc_usysr_DO_reg[5]/NET0131 ,
		_w7301_,
		_w10734_
	);
	LUT2 #(
		.INIT('h8)
	) name6688 (
		\bdma_BEAD_reg[5]/NET0131 ,
		_w7303_,
		_w10735_
	);
	LUT2 #(
		.INIT('h8)
	) name6689 (
		\bdma_BCTL_reg[5]/NET0131 ,
		_w7230_,
		_w10736_
	);
	LUT2 #(
		.INIT('h8)
	) name6690 (
		\pio_PINT_reg[5]/NET0131 ,
		_w7271_,
		_w10737_
	);
	LUT2 #(
		.INIT('h8)
	) name6691 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w7299_,
		_w10738_
	);
	LUT2 #(
		.INIT('h8)
	) name6692 (
		\PIO_out[5]_pad ,
		_w7291_,
		_w10739_
	);
	LUT2 #(
		.INIT('h8)
	) name6693 (
		\PIO_oe[5]_pad ,
		_w7244_,
		_w10740_
	);
	LUT2 #(
		.INIT('h8)
	) name6694 (
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w7273_,
		_w10741_
	);
	LUT2 #(
		.INIT('h1)
	) name6695 (
		_w7522_,
		_w10711_,
		_w10742_
	);
	LUT2 #(
		.INIT('h1)
	) name6696 (
		_w10712_,
		_w10713_,
		_w10743_
	);
	LUT2 #(
		.INIT('h1)
	) name6697 (
		_w10718_,
		_w10719_,
		_w10744_
	);
	LUT2 #(
		.INIT('h1)
	) name6698 (
		_w10720_,
		_w10721_,
		_w10745_
	);
	LUT2 #(
		.INIT('h1)
	) name6699 (
		_w10722_,
		_w10723_,
		_w10746_
	);
	LUT2 #(
		.INIT('h1)
	) name6700 (
		_w10724_,
		_w10725_,
		_w10747_
	);
	LUT2 #(
		.INIT('h1)
	) name6701 (
		_w10726_,
		_w10728_,
		_w10748_
	);
	LUT2 #(
		.INIT('h1)
	) name6702 (
		_w10729_,
		_w10730_,
		_w10749_
	);
	LUT2 #(
		.INIT('h1)
	) name6703 (
		_w10731_,
		_w10733_,
		_w10750_
	);
	LUT2 #(
		.INIT('h1)
	) name6704 (
		_w10734_,
		_w10737_,
		_w10751_
	);
	LUT2 #(
		.INIT('h1)
	) name6705 (
		_w10738_,
		_w10739_,
		_w10752_
	);
	LUT2 #(
		.INIT('h1)
	) name6706 (
		_w10740_,
		_w10741_,
		_w10753_
	);
	LUT2 #(
		.INIT('h8)
	) name6707 (
		_w10752_,
		_w10753_,
		_w10754_
	);
	LUT2 #(
		.INIT('h8)
	) name6708 (
		_w10750_,
		_w10751_,
		_w10755_
	);
	LUT2 #(
		.INIT('h8)
	) name6709 (
		_w10748_,
		_w10749_,
		_w10756_
	);
	LUT2 #(
		.INIT('h8)
	) name6710 (
		_w10746_,
		_w10747_,
		_w10757_
	);
	LUT2 #(
		.INIT('h8)
	) name6711 (
		_w10744_,
		_w10745_,
		_w10758_
	);
	LUT2 #(
		.INIT('h8)
	) name6712 (
		_w10742_,
		_w10743_,
		_w10759_
	);
	LUT2 #(
		.INIT('h8)
	) name6713 (
		_w10758_,
		_w10759_,
		_w10760_
	);
	LUT2 #(
		.INIT('h8)
	) name6714 (
		_w10756_,
		_w10757_,
		_w10761_
	);
	LUT2 #(
		.INIT('h8)
	) name6715 (
		_w10754_,
		_w10755_,
		_w10762_
	);
	LUT2 #(
		.INIT('h8)
	) name6716 (
		_w10761_,
		_w10762_,
		_w10763_
	);
	LUT2 #(
		.INIT('h4)
	) name6717 (
		_w10727_,
		_w10760_,
		_w10764_
	);
	LUT2 #(
		.INIT('h1)
	) name6718 (
		_w10735_,
		_w10736_,
		_w10765_
	);
	LUT2 #(
		.INIT('h8)
	) name6719 (
		_w10764_,
		_w10765_,
		_w10766_
	);
	LUT2 #(
		.INIT('h4)
	) name6720 (
		_w10717_,
		_w10763_,
		_w10767_
	);
	LUT2 #(
		.INIT('h4)
	) name6721 (
		_w10732_,
		_w10767_,
		_w10768_
	);
	LUT2 #(
		.INIT('h8)
	) name6722 (
		_w10766_,
		_w10768_,
		_w10769_
	);
	LUT2 #(
		.INIT('h2)
	) name6723 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w10769_,
		_w10770_
	);
	LUT2 #(
		.INIT('h8)
	) name6724 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w10771_
	);
	LUT2 #(
		.INIT('h2)
	) name6725 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4244_,
		_w10772_
	);
	LUT2 #(
		.INIT('h2)
	) name6726 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w7216_,
		_w10773_
	);
	LUT2 #(
		.INIT('h8)
	) name6727 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w10774_
	);
	LUT2 #(
		.INIT('h8)
	) name6728 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w10775_
	);
	LUT2 #(
		.INIT('h8)
	) name6729 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w10776_
	);
	LUT2 #(
		.INIT('h8)
	) name6730 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[5]/NET0131 ,
		_w10777_
	);
	LUT2 #(
		.INIT('h8)
	) name6731 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w10778_
	);
	LUT2 #(
		.INIT('h1)
	) name6732 (
		_w10771_,
		_w10774_,
		_w10779_
	);
	LUT2 #(
		.INIT('h1)
	) name6733 (
		_w10775_,
		_w10776_,
		_w10780_
	);
	LUT2 #(
		.INIT('h1)
	) name6734 (
		_w10777_,
		_w10778_,
		_w10781_
	);
	LUT2 #(
		.INIT('h8)
	) name6735 (
		_w10780_,
		_w10781_,
		_w10782_
	);
	LUT2 #(
		.INIT('h4)
	) name6736 (
		_w10773_,
		_w10779_,
		_w10783_
	);
	LUT2 #(
		.INIT('h8)
	) name6737 (
		_w10782_,
		_w10783_,
		_w10784_
	);
	LUT2 #(
		.INIT('h4)
	) name6738 (
		_w10772_,
		_w10784_,
		_w10785_
	);
	LUT2 #(
		.INIT('h2)
	) name6739 (
		_w7215_,
		_w10785_,
		_w10786_
	);
	LUT2 #(
		.INIT('h4)
	) name6740 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001 ,
		_w10787_
	);
	LUT2 #(
		.INIT('h8)
	) name6741 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001 ,
		_w10788_
	);
	LUT2 #(
		.INIT('h1)
	) name6742 (
		_w10787_,
		_w10788_,
		_w10789_
	);
	LUT2 #(
		.INIT('h2)
	) name6743 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w10789_,
		_w10790_
	);
	LUT2 #(
		.INIT('h4)
	) name6744 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001 ,
		_w10791_
	);
	LUT2 #(
		.INIT('h8)
	) name6745 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001 ,
		_w10792_
	);
	LUT2 #(
		.INIT('h1)
	) name6746 (
		_w10791_,
		_w10792_,
		_w10793_
	);
	LUT2 #(
		.INIT('h2)
	) name6747 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w10793_,
		_w10794_
	);
	LUT2 #(
		.INIT('h4)
	) name6748 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 ,
		_w10795_
	);
	LUT2 #(
		.INIT('h8)
	) name6749 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 ,
		_w10796_
	);
	LUT2 #(
		.INIT('h1)
	) name6750 (
		_w10795_,
		_w10796_,
		_w10797_
	);
	LUT2 #(
		.INIT('h2)
	) name6751 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w10797_,
		_w10798_
	);
	LUT2 #(
		.INIT('h4)
	) name6752 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 ,
		_w10799_
	);
	LUT2 #(
		.INIT('h8)
	) name6753 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 ,
		_w10800_
	);
	LUT2 #(
		.INIT('h1)
	) name6754 (
		_w10799_,
		_w10800_,
		_w10801_
	);
	LUT2 #(
		.INIT('h2)
	) name6755 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w10801_,
		_w10802_
	);
	LUT2 #(
		.INIT('h1)
	) name6756 (
		_w7169_,
		_w10790_,
		_w10803_
	);
	LUT2 #(
		.INIT('h1)
	) name6757 (
		_w10794_,
		_w10798_,
		_w10804_
	);
	LUT2 #(
		.INIT('h4)
	) name6758 (
		_w10802_,
		_w10804_,
		_w10805_
	);
	LUT2 #(
		.INIT('h8)
	) name6759 (
		_w10803_,
		_w10805_,
		_w10806_
	);
	LUT2 #(
		.INIT('h2)
	) name6760 (
		_w7153_,
		_w10806_,
		_w10807_
	);
	LUT2 #(
		.INIT('h8)
	) name6761 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131 ,
		_w10808_
	);
	LUT2 #(
		.INIT('h8)
	) name6762 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131 ,
		_w10809_
	);
	LUT2 #(
		.INIT('h8)
	) name6763 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131 ,
		_w10810_
	);
	LUT2 #(
		.INIT('h8)
	) name6764 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131 ,
		_w10811_
	);
	LUT2 #(
		.INIT('h8)
	) name6765 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131 ,
		_w10812_
	);
	LUT2 #(
		.INIT('h8)
	) name6766 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131 ,
		_w10813_
	);
	LUT2 #(
		.INIT('h8)
	) name6767 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131 ,
		_w10814_
	);
	LUT2 #(
		.INIT('h8)
	) name6768 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131 ,
		_w10815_
	);
	LUT2 #(
		.INIT('h8)
	) name6769 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w10816_
	);
	LUT2 #(
		.INIT('h8)
	) name6770 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[5]/NET0131 ,
		_w10817_
	);
	LUT2 #(
		.INIT('h8)
	) name6771 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		_w10818_
	);
	LUT2 #(
		.INIT('h8)
	) name6772 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 ,
		_w10819_
	);
	LUT2 #(
		.INIT('h1)
	) name6773 (
		_w10808_,
		_w10809_,
		_w10820_
	);
	LUT2 #(
		.INIT('h1)
	) name6774 (
		_w10810_,
		_w10811_,
		_w10821_
	);
	LUT2 #(
		.INIT('h1)
	) name6775 (
		_w10812_,
		_w10813_,
		_w10822_
	);
	LUT2 #(
		.INIT('h1)
	) name6776 (
		_w10814_,
		_w10815_,
		_w10823_
	);
	LUT2 #(
		.INIT('h1)
	) name6777 (
		_w10816_,
		_w10817_,
		_w10824_
	);
	LUT2 #(
		.INIT('h1)
	) name6778 (
		_w10818_,
		_w10819_,
		_w10825_
	);
	LUT2 #(
		.INIT('h8)
	) name6779 (
		_w10824_,
		_w10825_,
		_w10826_
	);
	LUT2 #(
		.INIT('h8)
	) name6780 (
		_w10822_,
		_w10823_,
		_w10827_
	);
	LUT2 #(
		.INIT('h8)
	) name6781 (
		_w10820_,
		_w10821_,
		_w10828_
	);
	LUT2 #(
		.INIT('h8)
	) name6782 (
		_w10827_,
		_w10828_,
		_w10829_
	);
	LUT2 #(
		.INIT('h8)
	) name6783 (
		_w10826_,
		_w10829_,
		_w10830_
	);
	LUT2 #(
		.INIT('h2)
	) name6784 (
		_w7068_,
		_w10830_,
		_w10831_
	);
	LUT2 #(
		.INIT('h8)
	) name6785 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w10832_
	);
	LUT2 #(
		.INIT('h8)
	) name6786 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131 ,
		_w10833_
	);
	LUT2 #(
		.INIT('h8)
	) name6787 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131 ,
		_w10834_
	);
	LUT2 #(
		.INIT('h8)
	) name6788 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131 ,
		_w10835_
	);
	LUT2 #(
		.INIT('h8)
	) name6789 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131 ,
		_w10836_
	);
	LUT2 #(
		.INIT('h8)
	) name6790 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131 ,
		_w10837_
	);
	LUT2 #(
		.INIT('h8)
	) name6791 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w10838_
	);
	LUT2 #(
		.INIT('h8)
	) name6792 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		_w10839_
	);
	LUT2 #(
		.INIT('h8)
	) name6793 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w10840_
	);
	LUT2 #(
		.INIT('h8)
	) name6794 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131 ,
		_w10841_
	);
	LUT2 #(
		.INIT('h8)
	) name6795 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131 ,
		_w10842_
	);
	LUT2 #(
		.INIT('h8)
	) name6796 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131 ,
		_w10843_
	);
	LUT2 #(
		.INIT('h1)
	) name6797 (
		_w10832_,
		_w10833_,
		_w10844_
	);
	LUT2 #(
		.INIT('h1)
	) name6798 (
		_w10834_,
		_w10835_,
		_w10845_
	);
	LUT2 #(
		.INIT('h1)
	) name6799 (
		_w10836_,
		_w10837_,
		_w10846_
	);
	LUT2 #(
		.INIT('h1)
	) name6800 (
		_w10838_,
		_w10839_,
		_w10847_
	);
	LUT2 #(
		.INIT('h1)
	) name6801 (
		_w10840_,
		_w10841_,
		_w10848_
	);
	LUT2 #(
		.INIT('h1)
	) name6802 (
		_w10842_,
		_w10843_,
		_w10849_
	);
	LUT2 #(
		.INIT('h8)
	) name6803 (
		_w10848_,
		_w10849_,
		_w10850_
	);
	LUT2 #(
		.INIT('h8)
	) name6804 (
		_w10846_,
		_w10847_,
		_w10851_
	);
	LUT2 #(
		.INIT('h8)
	) name6805 (
		_w10844_,
		_w10845_,
		_w10852_
	);
	LUT2 #(
		.INIT('h8)
	) name6806 (
		_w10851_,
		_w10852_,
		_w10853_
	);
	LUT2 #(
		.INIT('h8)
	) name6807 (
		_w10850_,
		_w10853_,
		_w10854_
	);
	LUT2 #(
		.INIT('h2)
	) name6808 (
		_w7128_,
		_w10854_,
		_w10855_
	);
	LUT2 #(
		.INIT('h4)
	) name6809 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001 ,
		_w10856_
	);
	LUT2 #(
		.INIT('h8)
	) name6810 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 ,
		_w10857_
	);
	LUT2 #(
		.INIT('h1)
	) name6811 (
		_w10856_,
		_w10857_,
		_w10858_
	);
	LUT2 #(
		.INIT('h2)
	) name6812 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w10858_,
		_w10859_
	);
	LUT2 #(
		.INIT('h4)
	) name6813 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001 ,
		_w10860_
	);
	LUT2 #(
		.INIT('h8)
	) name6814 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001 ,
		_w10861_
	);
	LUT2 #(
		.INIT('h1)
	) name6815 (
		_w10860_,
		_w10861_,
		_w10862_
	);
	LUT2 #(
		.INIT('h2)
	) name6816 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w10862_,
		_w10863_
	);
	LUT2 #(
		.INIT('h4)
	) name6817 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001 ,
		_w10864_
	);
	LUT2 #(
		.INIT('h8)
	) name6818 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001 ,
		_w10865_
	);
	LUT2 #(
		.INIT('h1)
	) name6819 (
		_w10864_,
		_w10865_,
		_w10866_
	);
	LUT2 #(
		.INIT('h2)
	) name6820 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w10866_,
		_w10867_
	);
	LUT2 #(
		.INIT('h4)
	) name6821 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001 ,
		_w10868_
	);
	LUT2 #(
		.INIT('h8)
	) name6822 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001 ,
		_w10869_
	);
	LUT2 #(
		.INIT('h1)
	) name6823 (
		_w10868_,
		_w10869_,
		_w10870_
	);
	LUT2 #(
		.INIT('h2)
	) name6824 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w10870_,
		_w10871_
	);
	LUT2 #(
		.INIT('h4)
	) name6825 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001 ,
		_w10872_
	);
	LUT2 #(
		.INIT('h8)
	) name6826 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001 ,
		_w10873_
	);
	LUT2 #(
		.INIT('h1)
	) name6827 (
		_w10872_,
		_w10873_,
		_w10874_
	);
	LUT2 #(
		.INIT('h2)
	) name6828 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w10874_,
		_w10875_
	);
	LUT2 #(
		.INIT('h4)
	) name6829 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001 ,
		_w10876_
	);
	LUT2 #(
		.INIT('h8)
	) name6830 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 ,
		_w10877_
	);
	LUT2 #(
		.INIT('h1)
	) name6831 (
		_w10876_,
		_w10877_,
		_w10878_
	);
	LUT2 #(
		.INIT('h2)
	) name6832 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w10878_,
		_w10879_
	);
	LUT2 #(
		.INIT('h4)
	) name6833 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 ,
		_w10880_
	);
	LUT2 #(
		.INIT('h8)
	) name6834 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 ,
		_w10881_
	);
	LUT2 #(
		.INIT('h1)
	) name6835 (
		_w10880_,
		_w10881_,
		_w10882_
	);
	LUT2 #(
		.INIT('h2)
	) name6836 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w10882_,
		_w10883_
	);
	LUT2 #(
		.INIT('h1)
	) name6837 (
		_w10859_,
		_w10863_,
		_w10884_
	);
	LUT2 #(
		.INIT('h1)
	) name6838 (
		_w10867_,
		_w10871_,
		_w10885_
	);
	LUT2 #(
		.INIT('h1)
	) name6839 (
		_w10875_,
		_w10879_,
		_w10886_
	);
	LUT2 #(
		.INIT('h4)
	) name6840 (
		_w10883_,
		_w10886_,
		_w10887_
	);
	LUT2 #(
		.INIT('h8)
	) name6841 (
		_w10884_,
		_w10885_,
		_w10888_
	);
	LUT2 #(
		.INIT('h8)
	) name6842 (
		_w10887_,
		_w10888_,
		_w10889_
	);
	LUT2 #(
		.INIT('h2)
	) name6843 (
		_w7179_,
		_w10889_,
		_w10890_
	);
	LUT2 #(
		.INIT('h8)
	) name6844 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[5]/P0001 ,
		_w10891_
	);
	LUT2 #(
		.INIT('h8)
	) name6845 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w10892_
	);
	LUT2 #(
		.INIT('h8)
	) name6846 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[5]/P0001 ,
		_w10893_
	);
	LUT2 #(
		.INIT('h8)
	) name6847 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w10894_
	);
	LUT2 #(
		.INIT('h1)
	) name6848 (
		_w10891_,
		_w10892_,
		_w10895_
	);
	LUT2 #(
		.INIT('h1)
	) name6849 (
		_w10893_,
		_w10894_,
		_w10896_
	);
	LUT2 #(
		.INIT('h8)
	) name6850 (
		_w10895_,
		_w10896_,
		_w10897_
	);
	LUT2 #(
		.INIT('h2)
	) name6851 (
		_w7119_,
		_w10897_,
		_w10898_
	);
	LUT2 #(
		.INIT('h1)
	) name6852 (
		_w10831_,
		_w10898_,
		_w10899_
	);
	LUT2 #(
		.INIT('h4)
	) name6853 (
		_w10855_,
		_w10899_,
		_w10900_
	);
	LUT2 #(
		.INIT('h1)
	) name6854 (
		_w10710_,
		_w10807_,
		_w10901_
	);
	LUT2 #(
		.INIT('h4)
	) name6855 (
		_w10890_,
		_w10901_,
		_w10902_
	);
	LUT2 #(
		.INIT('h8)
	) name6856 (
		_w10900_,
		_w10902_,
		_w10903_
	);
	LUT2 #(
		.INIT('h4)
	) name6857 (
		_w10786_,
		_w10903_,
		_w10904_
	);
	LUT2 #(
		.INIT('h4)
	) name6858 (
		_w10770_,
		_w10904_,
		_w10905_
	);
	LUT2 #(
		.INIT('h4)
	) name6859 (
		_w10683_,
		_w10905_,
		_w10906_
	);
	LUT2 #(
		.INIT('h1)
	) name6860 (
		\emc_DMDoe_reg/NET0131 ,
		_w10906_,
		_w10907_
	);
	LUT2 #(
		.INIT('h8)
	) name6861 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[5]/P0001 ,
		_w10908_
	);
	LUT2 #(
		.INIT('h2)
	) name6862 (
		_w7057_,
		_w10908_,
		_w10909_
	);
	LUT2 #(
		.INIT('h4)
	) name6863 (
		_w10907_,
		_w10909_,
		_w10910_
	);
	LUT2 #(
		.INIT('h1)
	) name6864 (
		_w10682_,
		_w10910_,
		_w10911_
	);
	LUT2 #(
		.INIT('h2)
	) name6865 (
		_w6135_,
		_w10911_,
		_w10912_
	);
	LUT2 #(
		.INIT('h2)
	) name6866 (
		_w8964_,
		_w10912_,
		_w10913_
	);
	LUT2 #(
		.INIT('h4)
	) name6867 (
		_w10664_,
		_w10913_,
		_w10914_
	);
	LUT2 #(
		.INIT('h1)
	) name6868 (
		_w10641_,
		_w10914_,
		_w10915_
	);
	LUT2 #(
		.INIT('h4)
	) name6869 (
		_w10421_,
		_w10915_,
		_w10916_
	);
	LUT2 #(
		.INIT('h2)
	) name6870 (
		\core_dag_ilm2reg_I_reg[6]/NET0131 ,
		_w6647_,
		_w10917_
	);
	LUT2 #(
		.INIT('h1)
	) name6871 (
		_w6753_,
		_w6778_,
		_w10918_
	);
	LUT2 #(
		.INIT('h8)
	) name6872 (
		_w6819_,
		_w6821_,
		_w10919_
	);
	LUT2 #(
		.INIT('h2)
	) name6873 (
		_w6776_,
		_w10919_,
		_w10920_
	);
	LUT2 #(
		.INIT('h1)
	) name6874 (
		_w10918_,
		_w10920_,
		_w10921_
	);
	LUT2 #(
		.INIT('h8)
	) name6875 (
		_w10918_,
		_w10920_,
		_w10922_
	);
	LUT2 #(
		.INIT('h1)
	) name6876 (
		_w10921_,
		_w10922_,
		_w10923_
	);
	LUT2 #(
		.INIT('h8)
	) name6877 (
		_w8198_,
		_w10923_,
		_w10924_
	);
	LUT2 #(
		.INIT('h1)
	) name6878 (
		_w6693_,
		_w6749_,
		_w10925_
	);
	LUT2 #(
		.INIT('h8)
	) name6879 (
		_w6693_,
		_w6749_,
		_w10926_
	);
	LUT2 #(
		.INIT('h1)
	) name6880 (
		_w10925_,
		_w10926_,
		_w10927_
	);
	LUT2 #(
		.INIT('h4)
	) name6881 (
		_w8198_,
		_w10927_,
		_w10928_
	);
	LUT2 #(
		.INIT('h1)
	) name6882 (
		_w10924_,
		_w10928_,
		_w10929_
	);
	LUT2 #(
		.INIT('h1)
	) name6883 (
		_w10917_,
		_w10929_,
		_w10930_
	);
	LUT2 #(
		.INIT('h4)
	) name6884 (
		_w6176_,
		_w10930_,
		_w10931_
	);
	LUT2 #(
		.INIT('h8)
	) name6885 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		_w6262_,
		_w10932_
	);
	LUT2 #(
		.INIT('h1)
	) name6886 (
		_w6275_,
		_w6382_,
		_w10933_
	);
	LUT2 #(
		.INIT('h2)
	) name6887 (
		_w6309_,
		_w6372_,
		_w10934_
	);
	LUT2 #(
		.INIT('h2)
	) name6888 (
		_w6380_,
		_w10934_,
		_w10935_
	);
	LUT2 #(
		.INIT('h1)
	) name6889 (
		_w6260_,
		_w10935_,
		_w10936_
	);
	LUT2 #(
		.INIT('h1)
	) name6890 (
		_w6375_,
		_w10936_,
		_w10937_
	);
	LUT2 #(
		.INIT('h8)
	) name6891 (
		_w10933_,
		_w10937_,
		_w10938_
	);
	LUT2 #(
		.INIT('h1)
	) name6892 (
		_w10933_,
		_w10937_,
		_w10939_
	);
	LUT2 #(
		.INIT('h1)
	) name6893 (
		_w10938_,
		_w10939_,
		_w10940_
	);
	LUT2 #(
		.INIT('h4)
	) name6894 (
		_w7612_,
		_w10940_,
		_w10941_
	);
	LUT2 #(
		.INIT('h1)
	) name6895 (
		_w6241_,
		_w6511_,
		_w10942_
	);
	LUT2 #(
		.INIT('h2)
	) name6896 (
		_w6266_,
		_w10942_,
		_w10943_
	);
	LUT2 #(
		.INIT('h4)
	) name6897 (
		_w6266_,
		_w10942_,
		_w10944_
	);
	LUT2 #(
		.INIT('h1)
	) name6898 (
		_w10943_,
		_w10944_,
		_w10945_
	);
	LUT2 #(
		.INIT('h2)
	) name6899 (
		_w7612_,
		_w10945_,
		_w10946_
	);
	LUT2 #(
		.INIT('h2)
	) name6900 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w10941_,
		_w10947_
	);
	LUT2 #(
		.INIT('h4)
	) name6901 (
		_w10946_,
		_w10947_,
		_w10948_
	);
	LUT2 #(
		.INIT('h8)
	) name6902 (
		_w6496_,
		_w10940_,
		_w10949_
	);
	LUT2 #(
		.INIT('h1)
	) name6903 (
		_w6496_,
		_w10945_,
		_w10950_
	);
	LUT2 #(
		.INIT('h1)
	) name6904 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w10949_,
		_w10951_
	);
	LUT2 #(
		.INIT('h4)
	) name6905 (
		_w10950_,
		_w10951_,
		_w10952_
	);
	LUT2 #(
		.INIT('h1)
	) name6906 (
		_w10932_,
		_w10948_,
		_w10953_
	);
	LUT2 #(
		.INIT('h4)
	) name6907 (
		_w10952_,
		_w10953_,
		_w10954_
	);
	LUT2 #(
		.INIT('h8)
	) name6908 (
		_w6176_,
		_w10954_,
		_w10955_
	);
	LUT2 #(
		.INIT('h1)
	) name6909 (
		_w10931_,
		_w10955_,
		_w10956_
	);
	LUT2 #(
		.INIT('h2)
	) name6910 (
		_w6135_,
		_w10956_,
		_w10957_
	);
	LUT2 #(
		.INIT('h1)
	) name6911 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w6924_,
		_w10958_
	);
	LUT2 #(
		.INIT('h8)
	) name6912 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w6926_,
		_w10959_
	);
	LUT2 #(
		.INIT('h8)
	) name6913 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131 ,
		_w6988_,
		_w10960_
	);
	LUT2 #(
		.INIT('h8)
	) name6914 (
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w6976_,
		_w10961_
	);
	LUT2 #(
		.INIT('h8)
	) name6915 (
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w6972_,
		_w10962_
	);
	LUT2 #(
		.INIT('h8)
	) name6916 (
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w6974_,
		_w10963_
	);
	LUT2 #(
		.INIT('h8)
	) name6917 (
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		_w6970_,
		_w10964_
	);
	LUT2 #(
		.INIT('h1)
	) name6918 (
		_w10961_,
		_w10962_,
		_w10965_
	);
	LUT2 #(
		.INIT('h1)
	) name6919 (
		_w10963_,
		_w10964_,
		_w10966_
	);
	LUT2 #(
		.INIT('h8)
	) name6920 (
		_w10965_,
		_w10966_,
		_w10967_
	);
	LUT2 #(
		.INIT('h2)
	) name6921 (
		_w4055_,
		_w10967_,
		_w10968_
	);
	LUT2 #(
		.INIT('h8)
	) name6922 (
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w6958_,
		_w10969_
	);
	LUT2 #(
		.INIT('h8)
	) name6923 (
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w6960_,
		_w10970_
	);
	LUT2 #(
		.INIT('h8)
	) name6924 (
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w6962_,
		_w10971_
	);
	LUT2 #(
		.INIT('h8)
	) name6925 (
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		_w6964_,
		_w10972_
	);
	LUT2 #(
		.INIT('h1)
	) name6926 (
		_w10969_,
		_w10970_,
		_w10973_
	);
	LUT2 #(
		.INIT('h1)
	) name6927 (
		_w10971_,
		_w10972_,
		_w10974_
	);
	LUT2 #(
		.INIT('h8)
	) name6928 (
		_w10973_,
		_w10974_,
		_w10975_
	);
	LUT2 #(
		.INIT('h4)
	) name6929 (
		_w10968_,
		_w10975_,
		_w10976_
	);
	LUT2 #(
		.INIT('h1)
	) name6930 (
		_w6121_,
		_w10976_,
		_w10977_
	);
	LUT2 #(
		.INIT('h8)
	) name6931 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w6956_,
		_w10978_
	);
	LUT2 #(
		.INIT('h8)
	) name6932 (
		\core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 ,
		_w6084_,
		_w10979_
	);
	LUT2 #(
		.INIT('h8)
	) name6933 (
		_w6085_,
		_w10979_,
		_w10980_
	);
	LUT2 #(
		.INIT('h8)
	) name6934 (
		\core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 ,
		_w6142_,
		_w10981_
	);
	LUT2 #(
		.INIT('h8)
	) name6935 (
		\core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 ,
		_w6140_,
		_w10982_
	);
	LUT2 #(
		.INIT('h8)
	) name6936 (
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		_w8131_,
		_w10983_
	);
	LUT2 #(
		.INIT('h1)
	) name6937 (
		_w4055_,
		_w10980_,
		_w10984_
	);
	LUT2 #(
		.INIT('h1)
	) name6938 (
		_w10981_,
		_w10982_,
		_w10985_
	);
	LUT2 #(
		.INIT('h4)
	) name6939 (
		_w10983_,
		_w10985_,
		_w10986_
	);
	LUT2 #(
		.INIT('h8)
	) name6940 (
		_w10984_,
		_w10986_,
		_w10987_
	);
	LUT2 #(
		.INIT('h8)
	) name6941 (
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		_w6148_,
		_w10988_
	);
	LUT2 #(
		.INIT('h8)
	) name6942 (
		\core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 ,
		_w6154_,
		_w10989_
	);
	LUT2 #(
		.INIT('h8)
	) name6943 (
		\core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 ,
		_w6150_,
		_w10990_
	);
	LUT2 #(
		.INIT('h8)
	) name6944 (
		_w6095_,
		_w10979_,
		_w10991_
	);
	LUT2 #(
		.INIT('h1)
	) name6945 (
		_w10988_,
		_w10989_,
		_w10992_
	);
	LUT2 #(
		.INIT('h1)
	) name6946 (
		_w10990_,
		_w10991_,
		_w10993_
	);
	LUT2 #(
		.INIT('h8)
	) name6947 (
		_w10992_,
		_w10993_,
		_w10994_
	);
	LUT2 #(
		.INIT('h8)
	) name6948 (
		_w4055_,
		_w10994_,
		_w10995_
	);
	LUT2 #(
		.INIT('h1)
	) name6949 (
		_w10987_,
		_w10995_,
		_w10996_
	);
	LUT2 #(
		.INIT('h4)
	) name6950 (
		_w6111_,
		_w10996_,
		_w10997_
	);
	LUT2 #(
		.INIT('h1)
	) name6951 (
		_w10977_,
		_w10978_,
		_w10998_
	);
	LUT2 #(
		.INIT('h4)
	) name6952 (
		_w10997_,
		_w10998_,
		_w10999_
	);
	LUT2 #(
		.INIT('h2)
	) name6953 (
		_w5949_,
		_w10999_,
		_w11000_
	);
	LUT2 #(
		.INIT('h2)
	) name6954 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		_w6934_,
		_w11001_
	);
	LUT2 #(
		.INIT('h1)
	) name6955 (
		_w10959_,
		_w10960_,
		_w11002_
	);
	LUT2 #(
		.INIT('h8)
	) name6956 (
		_w6924_,
		_w11002_,
		_w11003_
	);
	LUT2 #(
		.INIT('h4)
	) name6957 (
		_w11001_,
		_w11003_,
		_w11004_
	);
	LUT2 #(
		.INIT('h4)
	) name6958 (
		_w11000_,
		_w11004_,
		_w11005_
	);
	LUT2 #(
		.INIT('h1)
	) name6959 (
		_w6176_,
		_w10958_,
		_w11006_
	);
	LUT2 #(
		.INIT('h4)
	) name6960 (
		_w11005_,
		_w11006_,
		_w11007_
	);
	LUT2 #(
		.INIT('h8)
	) name6961 (
		\core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 ,
		_w6084_,
		_w11008_
	);
	LUT2 #(
		.INIT('h8)
	) name6962 (
		_w6085_,
		_w11008_,
		_w11009_
	);
	LUT2 #(
		.INIT('h8)
	) name6963 (
		\core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 ,
		_w6140_,
		_w11010_
	);
	LUT2 #(
		.INIT('h8)
	) name6964 (
		\core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 ,
		_w6142_,
		_w11011_
	);
	LUT2 #(
		.INIT('h8)
	) name6965 (
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		_w8131_,
		_w11012_
	);
	LUT2 #(
		.INIT('h1)
	) name6966 (
		_w4055_,
		_w11009_,
		_w11013_
	);
	LUT2 #(
		.INIT('h1)
	) name6967 (
		_w11010_,
		_w11011_,
		_w11014_
	);
	LUT2 #(
		.INIT('h4)
	) name6968 (
		_w11012_,
		_w11014_,
		_w11015_
	);
	LUT2 #(
		.INIT('h8)
	) name6969 (
		_w11013_,
		_w11015_,
		_w11016_
	);
	LUT2 #(
		.INIT('h8)
	) name6970 (
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		_w6148_,
		_w11017_
	);
	LUT2 #(
		.INIT('h8)
	) name6971 (
		\core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 ,
		_w6154_,
		_w11018_
	);
	LUT2 #(
		.INIT('h8)
	) name6972 (
		\core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 ,
		_w6150_,
		_w11019_
	);
	LUT2 #(
		.INIT('h8)
	) name6973 (
		_w6095_,
		_w11008_,
		_w11020_
	);
	LUT2 #(
		.INIT('h1)
	) name6974 (
		_w11017_,
		_w11018_,
		_w11021_
	);
	LUT2 #(
		.INIT('h1)
	) name6975 (
		_w11019_,
		_w11020_,
		_w11022_
	);
	LUT2 #(
		.INIT('h8)
	) name6976 (
		_w11021_,
		_w11022_,
		_w11023_
	);
	LUT2 #(
		.INIT('h8)
	) name6977 (
		_w4055_,
		_w11023_,
		_w11024_
	);
	LUT2 #(
		.INIT('h1)
	) name6978 (
		_w11016_,
		_w11024_,
		_w11025_
	);
	LUT2 #(
		.INIT('h8)
	) name6979 (
		_w6176_,
		_w11025_,
		_w11026_
	);
	LUT2 #(
		.INIT('h1)
	) name6980 (
		_w6135_,
		_w11026_,
		_w11027_
	);
	LUT2 #(
		.INIT('h4)
	) name6981 (
		_w11007_,
		_w11027_,
		_w11028_
	);
	LUT2 #(
		.INIT('h1)
	) name6982 (
		_w7005_,
		_w11028_,
		_w11029_
	);
	LUT2 #(
		.INIT('h4)
	) name6983 (
		_w10957_,
		_w11029_,
		_w11030_
	);
	LUT2 #(
		.INIT('h2)
	) name6984 (
		_w10976_,
		_w10996_,
		_w11031_
	);
	LUT2 #(
		.INIT('h2)
	) name6985 (
		_w8153_,
		_w11031_,
		_w11032_
	);
	LUT2 #(
		.INIT('h8)
	) name6986 (
		\DM_rdm[7]_pad ,
		_w7016_,
		_w11033_
	);
	LUT2 #(
		.INIT('h8)
	) name6987 (
		\DM_rd1[7]_pad ,
		_w7022_,
		_w11034_
	);
	LUT2 #(
		.INIT('h8)
	) name6988 (
		\DM_rd4[7]_pad ,
		_w7028_,
		_w11035_
	);
	LUT2 #(
		.INIT('h8)
	) name6989 (
		\DM_rd6[7]_pad ,
		_w7031_,
		_w11036_
	);
	LUT2 #(
		.INIT('h8)
	) name6990 (
		\DM_rd7[7]_pad ,
		_w7034_,
		_w11037_
	);
	LUT2 #(
		.INIT('h8)
	) name6991 (
		\DM_rd3[7]_pad ,
		_w7038_,
		_w11038_
	);
	LUT2 #(
		.INIT('h2)
	) name6992 (
		\DM_rd0[7]_pad ,
		_w7053_,
		_w11039_
	);
	LUT2 #(
		.INIT('h8)
	) name6993 (
		\DM_rd5[7]_pad ,
		_w7043_,
		_w11040_
	);
	LUT2 #(
		.INIT('h8)
	) name6994 (
		\DM_rd2[7]_pad ,
		_w7041_,
		_w11041_
	);
	LUT2 #(
		.INIT('h1)
	) name6995 (
		_w11034_,
		_w11038_,
		_w11042_
	);
	LUT2 #(
		.INIT('h4)
	) name6996 (
		_w11041_,
		_w11042_,
		_w11043_
	);
	LUT2 #(
		.INIT('h1)
	) name6997 (
		_w7057_,
		_w11033_,
		_w11044_
	);
	LUT2 #(
		.INIT('h1)
	) name6998 (
		_w11036_,
		_w11037_,
		_w11045_
	);
	LUT2 #(
		.INIT('h8)
	) name6999 (
		_w11044_,
		_w11045_,
		_w11046_
	);
	LUT2 #(
		.INIT('h4)
	) name7000 (
		_w11035_,
		_w11043_,
		_w11047_
	);
	LUT2 #(
		.INIT('h4)
	) name7001 (
		_w11040_,
		_w11047_,
		_w11048_
	);
	LUT2 #(
		.INIT('h8)
	) name7002 (
		_w11046_,
		_w11048_,
		_w11049_
	);
	LUT2 #(
		.INIT('h4)
	) name7003 (
		_w11039_,
		_w11049_,
		_w11050_
	);
	LUT2 #(
		.INIT('h8)
	) name7004 (
		\regout_STD_C_reg[7]/P0001 ,
		_w6988_,
		_w11051_
	);
	LUT2 #(
		.INIT('h4)
	) name7005 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001 ,
		_w11052_
	);
	LUT2 #(
		.INIT('h8)
	) name7006 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001 ,
		_w11053_
	);
	LUT2 #(
		.INIT('h1)
	) name7007 (
		_w11052_,
		_w11053_,
		_w11054_
	);
	LUT2 #(
		.INIT('h2)
	) name7008 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w11054_,
		_w11055_
	);
	LUT2 #(
		.INIT('h4)
	) name7009 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001 ,
		_w11056_
	);
	LUT2 #(
		.INIT('h8)
	) name7010 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001 ,
		_w11057_
	);
	LUT2 #(
		.INIT('h1)
	) name7011 (
		_w11056_,
		_w11057_,
		_w11058_
	);
	LUT2 #(
		.INIT('h2)
	) name7012 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w11058_,
		_w11059_
	);
	LUT2 #(
		.INIT('h4)
	) name7013 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001 ,
		_w11060_
	);
	LUT2 #(
		.INIT('h8)
	) name7014 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001 ,
		_w11061_
	);
	LUT2 #(
		.INIT('h1)
	) name7015 (
		_w11060_,
		_w11061_,
		_w11062_
	);
	LUT2 #(
		.INIT('h2)
	) name7016 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w11062_,
		_w11063_
	);
	LUT2 #(
		.INIT('h4)
	) name7017 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001 ,
		_w11064_
	);
	LUT2 #(
		.INIT('h8)
	) name7018 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001 ,
		_w11065_
	);
	LUT2 #(
		.INIT('h1)
	) name7019 (
		_w11064_,
		_w11065_,
		_w11066_
	);
	LUT2 #(
		.INIT('h2)
	) name7020 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w11066_,
		_w11067_
	);
	LUT2 #(
		.INIT('h4)
	) name7021 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001 ,
		_w11068_
	);
	LUT2 #(
		.INIT('h8)
	) name7022 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001 ,
		_w11069_
	);
	LUT2 #(
		.INIT('h1)
	) name7023 (
		_w11068_,
		_w11069_,
		_w11070_
	);
	LUT2 #(
		.INIT('h2)
	) name7024 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w11070_,
		_w11071_
	);
	LUT2 #(
		.INIT('h8)
	) name7025 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w11072_
	);
	LUT2 #(
		.INIT('h1)
	) name7026 (
		_w11055_,
		_w11072_,
		_w11073_
	);
	LUT2 #(
		.INIT('h1)
	) name7027 (
		_w11059_,
		_w11063_,
		_w11074_
	);
	LUT2 #(
		.INIT('h1)
	) name7028 (
		_w11067_,
		_w11071_,
		_w11075_
	);
	LUT2 #(
		.INIT('h8)
	) name7029 (
		_w11074_,
		_w11075_,
		_w11076_
	);
	LUT2 #(
		.INIT('h8)
	) name7030 (
		_w11073_,
		_w11076_,
		_w11077_
	);
	LUT2 #(
		.INIT('h2)
	) name7031 (
		_w7093_,
		_w11077_,
		_w11078_
	);
	LUT2 #(
		.INIT('h8)
	) name7032 (
		\sport1_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w7263_,
		_w11079_
	);
	LUT2 #(
		.INIT('h8)
	) name7033 (
		\emc_WSCRext_reg_DO_reg[7]/NET0131 ,
		_w7514_,
		_w11080_
	);
	LUT2 #(
		.INIT('h8)
	) name7034 (
		\tm_tpr_reg_DO_reg[7]/NET0131 ,
		_w7293_,
		_w11081_
	);
	LUT2 #(
		.INIT('h8)
	) name7035 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		_w7287_,
		_w11082_
	);
	LUT2 #(
		.INIT('h8)
	) name7036 (
		\emc_WSCRreg_DO_reg[7]/NET0131 ,
		_w7251_,
		_w11083_
	);
	LUT2 #(
		.INIT('h8)
	) name7037 (
		\tm_TCR_TMP_reg[7]/NET0131 ,
		_w7289_,
		_w11084_
	);
	LUT2 #(
		.INIT('h8)
	) name7038 (
		\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w7256_,
		_w11085_
	);
	LUT2 #(
		.INIT('h8)
	) name7039 (
		\sport0_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w7295_,
		_w11086_
	);
	LUT2 #(
		.INIT('h8)
	) name7040 (
		\idma_DOVL_reg[7]/NET0131 ,
		_w7532_,
		_w11087_
	);
	LUT2 #(
		.INIT('h8)
	) name7041 (
		\tm_tsr_reg_DO_reg[7]/NET0131 ,
		_w7540_,
		_w11088_
	);
	LUT2 #(
		.INIT('h8)
	) name7042 (
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w7273_,
		_w11089_
	);
	LUT2 #(
		.INIT('h8)
	) name7043 (
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w7259_,
		_w11090_
	);
	LUT2 #(
		.INIT('h8)
	) name7044 (
		\pio_pmask_reg_DO_reg[7]/NET0131 ,
		_w7297_,
		_w11091_
	);
	LUT2 #(
		.INIT('h8)
	) name7045 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w7234_,
		_w11092_
	);
	LUT2 #(
		.INIT('h8)
	) name7046 (
		\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w7247_,
		_w11093_
	);
	LUT2 #(
		.INIT('h8)
	) name7047 (
		\sport0_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w7276_,
		_w11094_
	);
	LUT2 #(
		.INIT('h8)
	) name7048 (
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w7249_,
		_w11095_
	);
	LUT2 #(
		.INIT('h8)
	) name7049 (
		\sport1_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w7527_,
		_w11096_
	);
	LUT2 #(
		.INIT('h8)
	) name7050 (
		\bdma_BOVL_reg[7]/NET0131 ,
		_w7534_,
		_w11097_
	);
	LUT2 #(
		.INIT('h8)
	) name7051 (
		\clkc_ckr_reg_DO_reg[7]/NET0131 ,
		_w7239_,
		_w11098_
	);
	LUT2 #(
		.INIT('h8)
	) name7052 (
		\memc_usysr_DO_reg[7]/NET0131 ,
		_w7301_,
		_w11099_
	);
	LUT2 #(
		.INIT('h8)
	) name7053 (
		\bdma_BEAD_reg[7]/NET0131 ,
		_w7303_,
		_w11100_
	);
	LUT2 #(
		.INIT('h8)
	) name7054 (
		\bdma_BCTL_reg[7]/NET0131 ,
		_w7230_,
		_w11101_
	);
	LUT2 #(
		.INIT('h8)
	) name7055 (
		\pio_PINT_reg[7]/NET0131 ,
		_w7271_,
		_w11102_
	);
	LUT2 #(
		.INIT('h8)
	) name7056 (
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w7281_,
		_w11103_
	);
	LUT2 #(
		.INIT('h8)
	) name7057 (
		\PIO_out[7]_pad ,
		_w7291_,
		_w11104_
	);
	LUT2 #(
		.INIT('h8)
	) name7058 (
		\PIO_oe[7]_pad ,
		_w7244_,
		_w11105_
	);
	LUT2 #(
		.INIT('h8)
	) name7059 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w7299_,
		_w11106_
	);
	LUT2 #(
		.INIT('h1)
	) name7060 (
		_w7522_,
		_w11079_,
		_w11107_
	);
	LUT2 #(
		.INIT('h1)
	) name7061 (
		_w11080_,
		_w11081_,
		_w11108_
	);
	LUT2 #(
		.INIT('h1)
	) name7062 (
		_w11083_,
		_w11084_,
		_w11109_
	);
	LUT2 #(
		.INIT('h1)
	) name7063 (
		_w11085_,
		_w11086_,
		_w11110_
	);
	LUT2 #(
		.INIT('h1)
	) name7064 (
		_w11087_,
		_w11088_,
		_w11111_
	);
	LUT2 #(
		.INIT('h1)
	) name7065 (
		_w11089_,
		_w11090_,
		_w11112_
	);
	LUT2 #(
		.INIT('h1)
	) name7066 (
		_w11091_,
		_w11093_,
		_w11113_
	);
	LUT2 #(
		.INIT('h1)
	) name7067 (
		_w11094_,
		_w11095_,
		_w11114_
	);
	LUT2 #(
		.INIT('h1)
	) name7068 (
		_w11096_,
		_w11098_,
		_w11115_
	);
	LUT2 #(
		.INIT('h1)
	) name7069 (
		_w11099_,
		_w11102_,
		_w11116_
	);
	LUT2 #(
		.INIT('h1)
	) name7070 (
		_w11103_,
		_w11104_,
		_w11117_
	);
	LUT2 #(
		.INIT('h1)
	) name7071 (
		_w11105_,
		_w11106_,
		_w11118_
	);
	LUT2 #(
		.INIT('h8)
	) name7072 (
		_w11117_,
		_w11118_,
		_w11119_
	);
	LUT2 #(
		.INIT('h8)
	) name7073 (
		_w11115_,
		_w11116_,
		_w11120_
	);
	LUT2 #(
		.INIT('h8)
	) name7074 (
		_w11113_,
		_w11114_,
		_w11121_
	);
	LUT2 #(
		.INIT('h8)
	) name7075 (
		_w11111_,
		_w11112_,
		_w11122_
	);
	LUT2 #(
		.INIT('h8)
	) name7076 (
		_w11109_,
		_w11110_,
		_w11123_
	);
	LUT2 #(
		.INIT('h8)
	) name7077 (
		_w11107_,
		_w11108_,
		_w11124_
	);
	LUT2 #(
		.INIT('h8)
	) name7078 (
		_w11123_,
		_w11124_,
		_w11125_
	);
	LUT2 #(
		.INIT('h8)
	) name7079 (
		_w11121_,
		_w11122_,
		_w11126_
	);
	LUT2 #(
		.INIT('h8)
	) name7080 (
		_w11119_,
		_w11120_,
		_w11127_
	);
	LUT2 #(
		.INIT('h8)
	) name7081 (
		_w11126_,
		_w11127_,
		_w11128_
	);
	LUT2 #(
		.INIT('h4)
	) name7082 (
		_w11092_,
		_w11125_,
		_w11129_
	);
	LUT2 #(
		.INIT('h1)
	) name7083 (
		_w11100_,
		_w11101_,
		_w11130_
	);
	LUT2 #(
		.INIT('h8)
	) name7084 (
		_w11129_,
		_w11130_,
		_w11131_
	);
	LUT2 #(
		.INIT('h4)
	) name7085 (
		_w11082_,
		_w11128_,
		_w11132_
	);
	LUT2 #(
		.INIT('h4)
	) name7086 (
		_w11097_,
		_w11132_,
		_w11133_
	);
	LUT2 #(
		.INIT('h8)
	) name7087 (
		_w11131_,
		_w11133_,
		_w11134_
	);
	LUT2 #(
		.INIT('h2)
	) name7088 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w11134_,
		_w11135_
	);
	LUT2 #(
		.INIT('h8)
	) name7089 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w11136_
	);
	LUT2 #(
		.INIT('h2)
	) name7090 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7216_,
		_w11137_
	);
	LUT2 #(
		.INIT('h8)
	) name7091 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w11138_
	);
	LUT2 #(
		.INIT('h8)
	) name7092 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[7]/NET0131 ,
		_w11139_
	);
	LUT2 #(
		.INIT('h2)
	) name7093 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4656_,
		_w11140_
	);
	LUT2 #(
		.INIT('h8)
	) name7094 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w11141_
	);
	LUT2 #(
		.INIT('h8)
	) name7095 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w11142_
	);
	LUT2 #(
		.INIT('h1)
	) name7096 (
		_w11136_,
		_w11138_,
		_w11143_
	);
	LUT2 #(
		.INIT('h1)
	) name7097 (
		_w11139_,
		_w11141_,
		_w11144_
	);
	LUT2 #(
		.INIT('h4)
	) name7098 (
		_w11142_,
		_w11144_,
		_w11145_
	);
	LUT2 #(
		.INIT('h4)
	) name7099 (
		_w11137_,
		_w11143_,
		_w11146_
	);
	LUT2 #(
		.INIT('h8)
	) name7100 (
		_w11145_,
		_w11146_,
		_w11147_
	);
	LUT2 #(
		.INIT('h4)
	) name7101 (
		_w11140_,
		_w11147_,
		_w11148_
	);
	LUT2 #(
		.INIT('h2)
	) name7102 (
		_w7215_,
		_w11148_,
		_w11149_
	);
	LUT2 #(
		.INIT('h8)
	) name7103 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131 ,
		_w11150_
	);
	LUT2 #(
		.INIT('h8)
	) name7104 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131 ,
		_w11151_
	);
	LUT2 #(
		.INIT('h8)
	) name7105 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131 ,
		_w11152_
	);
	LUT2 #(
		.INIT('h8)
	) name7106 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131 ,
		_w11153_
	);
	LUT2 #(
		.INIT('h8)
	) name7107 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 ,
		_w11154_
	);
	LUT2 #(
		.INIT('h8)
	) name7108 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131 ,
		_w11155_
	);
	LUT2 #(
		.INIT('h8)
	) name7109 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 ,
		_w11156_
	);
	LUT2 #(
		.INIT('h8)
	) name7110 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131 ,
		_w11157_
	);
	LUT2 #(
		.INIT('h8)
	) name7111 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		_w11158_
	);
	LUT2 #(
		.INIT('h8)
	) name7112 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 ,
		_w11159_
	);
	LUT2 #(
		.INIT('h8)
	) name7113 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131 ,
		_w11160_
	);
	LUT2 #(
		.INIT('h8)
	) name7114 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131 ,
		_w11161_
	);
	LUT2 #(
		.INIT('h1)
	) name7115 (
		_w11150_,
		_w11151_,
		_w11162_
	);
	LUT2 #(
		.INIT('h1)
	) name7116 (
		_w11152_,
		_w11153_,
		_w11163_
	);
	LUT2 #(
		.INIT('h1)
	) name7117 (
		_w11154_,
		_w11155_,
		_w11164_
	);
	LUT2 #(
		.INIT('h1)
	) name7118 (
		_w11156_,
		_w11157_,
		_w11165_
	);
	LUT2 #(
		.INIT('h1)
	) name7119 (
		_w11158_,
		_w11159_,
		_w11166_
	);
	LUT2 #(
		.INIT('h1)
	) name7120 (
		_w11160_,
		_w11161_,
		_w11167_
	);
	LUT2 #(
		.INIT('h8)
	) name7121 (
		_w11166_,
		_w11167_,
		_w11168_
	);
	LUT2 #(
		.INIT('h8)
	) name7122 (
		_w11164_,
		_w11165_,
		_w11169_
	);
	LUT2 #(
		.INIT('h8)
	) name7123 (
		_w11162_,
		_w11163_,
		_w11170_
	);
	LUT2 #(
		.INIT('h8)
	) name7124 (
		_w11169_,
		_w11170_,
		_w11171_
	);
	LUT2 #(
		.INIT('h8)
	) name7125 (
		_w11168_,
		_w11171_,
		_w11172_
	);
	LUT2 #(
		.INIT('h2)
	) name7126 (
		_w7068_,
		_w11172_,
		_w11173_
	);
	LUT2 #(
		.INIT('h4)
	) name7127 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001 ,
		_w11174_
	);
	LUT2 #(
		.INIT('h8)
	) name7128 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001 ,
		_w11175_
	);
	LUT2 #(
		.INIT('h1)
	) name7129 (
		_w11174_,
		_w11175_,
		_w11176_
	);
	LUT2 #(
		.INIT('h2)
	) name7130 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w11176_,
		_w11177_
	);
	LUT2 #(
		.INIT('h4)
	) name7131 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001 ,
		_w11178_
	);
	LUT2 #(
		.INIT('h8)
	) name7132 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001 ,
		_w11179_
	);
	LUT2 #(
		.INIT('h1)
	) name7133 (
		_w11178_,
		_w11179_,
		_w11180_
	);
	LUT2 #(
		.INIT('h2)
	) name7134 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w11180_,
		_w11181_
	);
	LUT2 #(
		.INIT('h4)
	) name7135 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001 ,
		_w11182_
	);
	LUT2 #(
		.INIT('h8)
	) name7136 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001 ,
		_w11183_
	);
	LUT2 #(
		.INIT('h1)
	) name7137 (
		_w11182_,
		_w11183_,
		_w11184_
	);
	LUT2 #(
		.INIT('h2)
	) name7138 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w11184_,
		_w11185_
	);
	LUT2 #(
		.INIT('h4)
	) name7139 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001 ,
		_w11186_
	);
	LUT2 #(
		.INIT('h8)
	) name7140 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001 ,
		_w11187_
	);
	LUT2 #(
		.INIT('h1)
	) name7141 (
		_w11186_,
		_w11187_,
		_w11188_
	);
	LUT2 #(
		.INIT('h2)
	) name7142 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w11188_,
		_w11189_
	);
	LUT2 #(
		.INIT('h4)
	) name7143 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001 ,
		_w11190_
	);
	LUT2 #(
		.INIT('h8)
	) name7144 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 ,
		_w11191_
	);
	LUT2 #(
		.INIT('h1)
	) name7145 (
		_w11190_,
		_w11191_,
		_w11192_
	);
	LUT2 #(
		.INIT('h2)
	) name7146 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w11192_,
		_w11193_
	);
	LUT2 #(
		.INIT('h4)
	) name7147 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001 ,
		_w11194_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 ,
		_w11195_
	);
	LUT2 #(
		.INIT('h1)
	) name7149 (
		_w11194_,
		_w11195_,
		_w11196_
	);
	LUT2 #(
		.INIT('h2)
	) name7150 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w11196_,
		_w11197_
	);
	LUT2 #(
		.INIT('h1)
	) name7151 (
		_w7207_,
		_w11177_,
		_w11198_
	);
	LUT2 #(
		.INIT('h1)
	) name7152 (
		_w11181_,
		_w11185_,
		_w11199_
	);
	LUT2 #(
		.INIT('h1)
	) name7153 (
		_w11189_,
		_w11193_,
		_w11200_
	);
	LUT2 #(
		.INIT('h4)
	) name7154 (
		_w11197_,
		_w11200_,
		_w11201_
	);
	LUT2 #(
		.INIT('h8)
	) name7155 (
		_w11198_,
		_w11199_,
		_w11202_
	);
	LUT2 #(
		.INIT('h8)
	) name7156 (
		_w11201_,
		_w11202_,
		_w11203_
	);
	LUT2 #(
		.INIT('h2)
	) name7157 (
		_w7179_,
		_w11203_,
		_w11204_
	);
	LUT2 #(
		.INIT('h8)
	) name7158 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131 ,
		_w11205_
	);
	LUT2 #(
		.INIT('h8)
	) name7159 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131 ,
		_w11206_
	);
	LUT2 #(
		.INIT('h8)
	) name7160 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131 ,
		_w11207_
	);
	LUT2 #(
		.INIT('h8)
	) name7161 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w11208_
	);
	LUT2 #(
		.INIT('h8)
	) name7162 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 ,
		_w11209_
	);
	LUT2 #(
		.INIT('h8)
	) name7163 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131 ,
		_w11210_
	);
	LUT2 #(
		.INIT('h8)
	) name7164 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131 ,
		_w11211_
	);
	LUT2 #(
		.INIT('h8)
	) name7165 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131 ,
		_w11212_
	);
	LUT2 #(
		.INIT('h8)
	) name7166 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131 ,
		_w11213_
	);
	LUT2 #(
		.INIT('h8)
	) name7167 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w11214_
	);
	LUT2 #(
		.INIT('h8)
	) name7168 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 ,
		_w11215_
	);
	LUT2 #(
		.INIT('h8)
	) name7169 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131 ,
		_w11216_
	);
	LUT2 #(
		.INIT('h1)
	) name7170 (
		_w11205_,
		_w11206_,
		_w11217_
	);
	LUT2 #(
		.INIT('h1)
	) name7171 (
		_w11207_,
		_w11208_,
		_w11218_
	);
	LUT2 #(
		.INIT('h1)
	) name7172 (
		_w11209_,
		_w11210_,
		_w11219_
	);
	LUT2 #(
		.INIT('h1)
	) name7173 (
		_w11211_,
		_w11212_,
		_w11220_
	);
	LUT2 #(
		.INIT('h1)
	) name7174 (
		_w11213_,
		_w11214_,
		_w11221_
	);
	LUT2 #(
		.INIT('h1)
	) name7175 (
		_w11215_,
		_w11216_,
		_w11222_
	);
	LUT2 #(
		.INIT('h8)
	) name7176 (
		_w11221_,
		_w11222_,
		_w11223_
	);
	LUT2 #(
		.INIT('h8)
	) name7177 (
		_w11219_,
		_w11220_,
		_w11224_
	);
	LUT2 #(
		.INIT('h8)
	) name7178 (
		_w11217_,
		_w11218_,
		_w11225_
	);
	LUT2 #(
		.INIT('h8)
	) name7179 (
		_w11224_,
		_w11225_,
		_w11226_
	);
	LUT2 #(
		.INIT('h8)
	) name7180 (
		_w11223_,
		_w11226_,
		_w11227_
	);
	LUT2 #(
		.INIT('h2)
	) name7181 (
		_w7128_,
		_w11227_,
		_w11228_
	);
	LUT2 #(
		.INIT('h4)
	) name7182 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 ,
		_w11229_
	);
	LUT2 #(
		.INIT('h8)
	) name7183 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 ,
		_w11230_
	);
	LUT2 #(
		.INIT('h1)
	) name7184 (
		_w11229_,
		_w11230_,
		_w11231_
	);
	LUT2 #(
		.INIT('h2)
	) name7185 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w11231_,
		_w11232_
	);
	LUT2 #(
		.INIT('h4)
	) name7186 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001 ,
		_w11233_
	);
	LUT2 #(
		.INIT('h8)
	) name7187 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001 ,
		_w11234_
	);
	LUT2 #(
		.INIT('h1)
	) name7188 (
		_w11233_,
		_w11234_,
		_w11235_
	);
	LUT2 #(
		.INIT('h2)
	) name7189 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w11235_,
		_w11236_
	);
	LUT2 #(
		.INIT('h4)
	) name7190 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 ,
		_w11237_
	);
	LUT2 #(
		.INIT('h8)
	) name7191 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 ,
		_w11238_
	);
	LUT2 #(
		.INIT('h1)
	) name7192 (
		_w11237_,
		_w11238_,
		_w11239_
	);
	LUT2 #(
		.INIT('h2)
	) name7193 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w11239_,
		_w11240_
	);
	LUT2 #(
		.INIT('h1)
	) name7194 (
		_w11232_,
		_w11236_,
		_w11241_
	);
	LUT2 #(
		.INIT('h4)
	) name7195 (
		_w11240_,
		_w11241_,
		_w11242_
	);
	LUT2 #(
		.INIT('h8)
	) name7196 (
		_w7174_,
		_w11242_,
		_w11243_
	);
	LUT2 #(
		.INIT('h2)
	) name7197 (
		_w7153_,
		_w11243_,
		_w11244_
	);
	LUT2 #(
		.INIT('h8)
	) name7198 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[7]/P0001 ,
		_w11245_
	);
	LUT2 #(
		.INIT('h8)
	) name7199 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[7]/P0001 ,
		_w11246_
	);
	LUT2 #(
		.INIT('h8)
	) name7200 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[7]/P0001 ,
		_w11247_
	);
	LUT2 #(
		.INIT('h8)
	) name7201 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w11248_
	);
	LUT2 #(
		.INIT('h1)
	) name7202 (
		_w11245_,
		_w11246_,
		_w11249_
	);
	LUT2 #(
		.INIT('h1)
	) name7203 (
		_w11247_,
		_w11248_,
		_w11250_
	);
	LUT2 #(
		.INIT('h8)
	) name7204 (
		_w11249_,
		_w11250_,
		_w11251_
	);
	LUT2 #(
		.INIT('h2)
	) name7205 (
		_w7119_,
		_w11251_,
		_w11252_
	);
	LUT2 #(
		.INIT('h1)
	) name7206 (
		_w11173_,
		_w11252_,
		_w11253_
	);
	LUT2 #(
		.INIT('h4)
	) name7207 (
		_w11228_,
		_w11253_,
		_w11254_
	);
	LUT2 #(
		.INIT('h1)
	) name7208 (
		_w11078_,
		_w11204_,
		_w11255_
	);
	LUT2 #(
		.INIT('h4)
	) name7209 (
		_w11244_,
		_w11255_,
		_w11256_
	);
	LUT2 #(
		.INIT('h8)
	) name7210 (
		_w11254_,
		_w11256_,
		_w11257_
	);
	LUT2 #(
		.INIT('h4)
	) name7211 (
		_w11149_,
		_w11257_,
		_w11258_
	);
	LUT2 #(
		.INIT('h4)
	) name7212 (
		_w11135_,
		_w11258_,
		_w11259_
	);
	LUT2 #(
		.INIT('h4)
	) name7213 (
		_w11051_,
		_w11259_,
		_w11260_
	);
	LUT2 #(
		.INIT('h1)
	) name7214 (
		\emc_DMDoe_reg/NET0131 ,
		_w11260_,
		_w11261_
	);
	LUT2 #(
		.INIT('h8)
	) name7215 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[7]/P0001 ,
		_w11262_
	);
	LUT2 #(
		.INIT('h2)
	) name7216 (
		_w7057_,
		_w11262_,
		_w11263_
	);
	LUT2 #(
		.INIT('h4)
	) name7217 (
		_w11261_,
		_w11263_,
		_w11264_
	);
	LUT2 #(
		.INIT('h1)
	) name7218 (
		_w11050_,
		_w11264_,
		_w11265_
	);
	LUT2 #(
		.INIT('h8)
	) name7219 (
		_w7863_,
		_w11265_,
		_w11266_
	);
	LUT2 #(
		.INIT('h1)
	) name7220 (
		_w11032_,
		_w11266_,
		_w11267_
	);
	LUT2 #(
		.INIT('h2)
	) name7221 (
		_w7005_,
		_w11267_,
		_w11268_
	);
	LUT2 #(
		.INIT('h2)
	) name7222 (
		\core_dag_ilm1reg_I_reg[6]/NET0131 ,
		_w6238_,
		_w11269_
	);
	LUT2 #(
		.INIT('h1)
	) name7223 (
		_w6242_,
		_w6510_,
		_w11270_
	);
	LUT2 #(
		.INIT('h8)
	) name7224 (
		_w6242_,
		_w6510_,
		_w11271_
	);
	LUT2 #(
		.INIT('h1)
	) name7225 (
		_w11270_,
		_w11271_,
		_w11272_
	);
	LUT2 #(
		.INIT('h2)
	) name7226 (
		_w7631_,
		_w11272_,
		_w11273_
	);
	LUT2 #(
		.INIT('h1)
	) name7227 (
		_w6260_,
		_w6375_,
		_w11274_
	);
	LUT2 #(
		.INIT('h4)
	) name7228 (
		_w10935_,
		_w11274_,
		_w11275_
	);
	LUT2 #(
		.INIT('h2)
	) name7229 (
		_w10935_,
		_w11274_,
		_w11276_
	);
	LUT2 #(
		.INIT('h1)
	) name7230 (
		_w11275_,
		_w11276_,
		_w11277_
	);
	LUT2 #(
		.INIT('h4)
	) name7231 (
		_w7631_,
		_w11277_,
		_w11278_
	);
	LUT2 #(
		.INIT('h1)
	) name7232 (
		_w11269_,
		_w11273_,
		_w11279_
	);
	LUT2 #(
		.INIT('h4)
	) name7233 (
		_w11278_,
		_w11279_,
		_w11280_
	);
	LUT2 #(
		.INIT('h4)
	) name7234 (
		_w6135_,
		_w11280_,
		_w11281_
	);
	LUT2 #(
		.INIT('h8)
	) name7235 (
		\DM_rdm[6]_pad ,
		_w7016_,
		_w11282_
	);
	LUT2 #(
		.INIT('h8)
	) name7236 (
		\DM_rd1[6]_pad ,
		_w7022_,
		_w11283_
	);
	LUT2 #(
		.INIT('h8)
	) name7237 (
		\DM_rd4[6]_pad ,
		_w7028_,
		_w11284_
	);
	LUT2 #(
		.INIT('h8)
	) name7238 (
		\DM_rd6[6]_pad ,
		_w7031_,
		_w11285_
	);
	LUT2 #(
		.INIT('h8)
	) name7239 (
		\DM_rd7[6]_pad ,
		_w7034_,
		_w11286_
	);
	LUT2 #(
		.INIT('h8)
	) name7240 (
		\DM_rd3[6]_pad ,
		_w7038_,
		_w11287_
	);
	LUT2 #(
		.INIT('h2)
	) name7241 (
		\DM_rd0[6]_pad ,
		_w7053_,
		_w11288_
	);
	LUT2 #(
		.INIT('h8)
	) name7242 (
		\DM_rd5[6]_pad ,
		_w7043_,
		_w11289_
	);
	LUT2 #(
		.INIT('h8)
	) name7243 (
		\DM_rd2[6]_pad ,
		_w7041_,
		_w11290_
	);
	LUT2 #(
		.INIT('h1)
	) name7244 (
		_w11283_,
		_w11287_,
		_w11291_
	);
	LUT2 #(
		.INIT('h4)
	) name7245 (
		_w11290_,
		_w11291_,
		_w11292_
	);
	LUT2 #(
		.INIT('h1)
	) name7246 (
		_w7057_,
		_w11282_,
		_w11293_
	);
	LUT2 #(
		.INIT('h1)
	) name7247 (
		_w11285_,
		_w11286_,
		_w11294_
	);
	LUT2 #(
		.INIT('h8)
	) name7248 (
		_w11293_,
		_w11294_,
		_w11295_
	);
	LUT2 #(
		.INIT('h4)
	) name7249 (
		_w11284_,
		_w11292_,
		_w11296_
	);
	LUT2 #(
		.INIT('h4)
	) name7250 (
		_w11289_,
		_w11296_,
		_w11297_
	);
	LUT2 #(
		.INIT('h8)
	) name7251 (
		_w11295_,
		_w11297_,
		_w11298_
	);
	LUT2 #(
		.INIT('h4)
	) name7252 (
		_w11288_,
		_w11298_,
		_w11299_
	);
	LUT2 #(
		.INIT('h8)
	) name7253 (
		\regout_STD_C_reg[6]/P0001 ,
		_w6988_,
		_w11300_
	);
	LUT2 #(
		.INIT('h4)
	) name7254 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001 ,
		_w11301_
	);
	LUT2 #(
		.INIT('h8)
	) name7255 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001 ,
		_w11302_
	);
	LUT2 #(
		.INIT('h1)
	) name7256 (
		_w11301_,
		_w11302_,
		_w11303_
	);
	LUT2 #(
		.INIT('h2)
	) name7257 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w11303_,
		_w11304_
	);
	LUT2 #(
		.INIT('h4)
	) name7258 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001 ,
		_w11305_
	);
	LUT2 #(
		.INIT('h8)
	) name7259 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001 ,
		_w11306_
	);
	LUT2 #(
		.INIT('h1)
	) name7260 (
		_w11305_,
		_w11306_,
		_w11307_
	);
	LUT2 #(
		.INIT('h2)
	) name7261 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w11307_,
		_w11308_
	);
	LUT2 #(
		.INIT('h4)
	) name7262 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 ,
		_w11309_
	);
	LUT2 #(
		.INIT('h8)
	) name7263 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 ,
		_w11310_
	);
	LUT2 #(
		.INIT('h1)
	) name7264 (
		_w11309_,
		_w11310_,
		_w11311_
	);
	LUT2 #(
		.INIT('h2)
	) name7265 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w11311_,
		_w11312_
	);
	LUT2 #(
		.INIT('h4)
	) name7266 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 ,
		_w11313_
	);
	LUT2 #(
		.INIT('h8)
	) name7267 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 ,
		_w11314_
	);
	LUT2 #(
		.INIT('h1)
	) name7268 (
		_w11313_,
		_w11314_,
		_w11315_
	);
	LUT2 #(
		.INIT('h2)
	) name7269 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w11315_,
		_w11316_
	);
	LUT2 #(
		.INIT('h1)
	) name7270 (
		_w7169_,
		_w11304_,
		_w11317_
	);
	LUT2 #(
		.INIT('h1)
	) name7271 (
		_w11308_,
		_w11312_,
		_w11318_
	);
	LUT2 #(
		.INIT('h4)
	) name7272 (
		_w11316_,
		_w11318_,
		_w11319_
	);
	LUT2 #(
		.INIT('h8)
	) name7273 (
		_w11317_,
		_w11319_,
		_w11320_
	);
	LUT2 #(
		.INIT('h2)
	) name7274 (
		_w7153_,
		_w11320_,
		_w11321_
	);
	LUT2 #(
		.INIT('h2)
	) name7275 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		_w4174_,
		_w11322_
	);
	LUT2 #(
		.INIT('h4)
	) name7276 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001 ,
		_w11323_
	);
	LUT2 #(
		.INIT('h8)
	) name7277 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001 ,
		_w11324_
	);
	LUT2 #(
		.INIT('h1)
	) name7278 (
		_w11323_,
		_w11324_,
		_w11325_
	);
	LUT2 #(
		.INIT('h2)
	) name7279 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w11325_,
		_w11326_
	);
	LUT2 #(
		.INIT('h4)
	) name7280 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001 ,
		_w11327_
	);
	LUT2 #(
		.INIT('h8)
	) name7281 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001 ,
		_w11328_
	);
	LUT2 #(
		.INIT('h1)
	) name7282 (
		_w11327_,
		_w11328_,
		_w11329_
	);
	LUT2 #(
		.INIT('h2)
	) name7283 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w11329_,
		_w11330_
	);
	LUT2 #(
		.INIT('h4)
	) name7284 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001 ,
		_w11331_
	);
	LUT2 #(
		.INIT('h8)
	) name7285 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001 ,
		_w11332_
	);
	LUT2 #(
		.INIT('h1)
	) name7286 (
		_w11331_,
		_w11332_,
		_w11333_
	);
	LUT2 #(
		.INIT('h2)
	) name7287 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w11333_,
		_w11334_
	);
	LUT2 #(
		.INIT('h4)
	) name7288 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001 ,
		_w11335_
	);
	LUT2 #(
		.INIT('h8)
	) name7289 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001 ,
		_w11336_
	);
	LUT2 #(
		.INIT('h1)
	) name7290 (
		_w11335_,
		_w11336_,
		_w11337_
	);
	LUT2 #(
		.INIT('h2)
	) name7291 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w11337_,
		_w11338_
	);
	LUT2 #(
		.INIT('h4)
	) name7292 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001 ,
		_w11339_
	);
	LUT2 #(
		.INIT('h8)
	) name7293 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001 ,
		_w11340_
	);
	LUT2 #(
		.INIT('h1)
	) name7294 (
		_w11339_,
		_w11340_,
		_w11341_
	);
	LUT2 #(
		.INIT('h2)
	) name7295 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w11341_,
		_w11342_
	);
	LUT2 #(
		.INIT('h1)
	) name7296 (
		_w11326_,
		_w11330_,
		_w11343_
	);
	LUT2 #(
		.INIT('h1)
	) name7297 (
		_w11334_,
		_w11338_,
		_w11344_
	);
	LUT2 #(
		.INIT('h4)
	) name7298 (
		_w11342_,
		_w11344_,
		_w11345_
	);
	LUT2 #(
		.INIT('h8)
	) name7299 (
		_w11343_,
		_w11345_,
		_w11346_
	);
	LUT2 #(
		.INIT('h4)
	) name7300 (
		_w11322_,
		_w11346_,
		_w11347_
	);
	LUT2 #(
		.INIT('h2)
	) name7301 (
		_w7093_,
		_w11347_,
		_w11348_
	);
	LUT2 #(
		.INIT('h8)
	) name7302 (
		\sport1_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w7263_,
		_w11349_
	);
	LUT2 #(
		.INIT('h8)
	) name7303 (
		\emc_WSCRext_reg_DO_reg[6]/NET0131 ,
		_w7514_,
		_w11350_
	);
	LUT2 #(
		.INIT('h8)
	) name7304 (
		\tm_tpr_reg_DO_reg[6]/NET0131 ,
		_w7293_,
		_w11351_
	);
	LUT2 #(
		.INIT('h8)
	) name7305 (
		\bdma_BWCOUNT_reg[6]/NET0131 ,
		_w7287_,
		_w11352_
	);
	LUT2 #(
		.INIT('h8)
	) name7306 (
		\emc_WSCRreg_DO_reg[6]/NET0131 ,
		_w7251_,
		_w11353_
	);
	LUT2 #(
		.INIT('h8)
	) name7307 (
		\tm_TCR_TMP_reg[6]/NET0131 ,
		_w7289_,
		_w11354_
	);
	LUT2 #(
		.INIT('h8)
	) name7308 (
		\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w7256_,
		_w11355_
	);
	LUT2 #(
		.INIT('h8)
	) name7309 (
		\sport0_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w7295_,
		_w11356_
	);
	LUT2 #(
		.INIT('h8)
	) name7310 (
		\idma_DOVL_reg[6]/NET0131 ,
		_w7532_,
		_w11357_
	);
	LUT2 #(
		.INIT('h8)
	) name7311 (
		\tm_tsr_reg_DO_reg[6]/NET0131 ,
		_w7540_,
		_w11358_
	);
	LUT2 #(
		.INIT('h8)
	) name7312 (
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w7273_,
		_w11359_
	);
	LUT2 #(
		.INIT('h8)
	) name7313 (
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w7259_,
		_w11360_
	);
	LUT2 #(
		.INIT('h8)
	) name7314 (
		\pio_pmask_reg_DO_reg[6]/NET0131 ,
		_w7297_,
		_w11361_
	);
	LUT2 #(
		.INIT('h8)
	) name7315 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w7234_,
		_w11362_
	);
	LUT2 #(
		.INIT('h8)
	) name7316 (
		\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w7247_,
		_w11363_
	);
	LUT2 #(
		.INIT('h8)
	) name7317 (
		\sport0_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w7276_,
		_w11364_
	);
	LUT2 #(
		.INIT('h8)
	) name7318 (
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w7249_,
		_w11365_
	);
	LUT2 #(
		.INIT('h8)
	) name7319 (
		\sport1_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w7527_,
		_w11366_
	);
	LUT2 #(
		.INIT('h8)
	) name7320 (
		\bdma_BOVL_reg[6]/NET0131 ,
		_w7534_,
		_w11367_
	);
	LUT2 #(
		.INIT('h8)
	) name7321 (
		\clkc_ckr_reg_DO_reg[6]/NET0131 ,
		_w7239_,
		_w11368_
	);
	LUT2 #(
		.INIT('h8)
	) name7322 (
		\memc_usysr_DO_reg[6]/NET0131 ,
		_w7301_,
		_w11369_
	);
	LUT2 #(
		.INIT('h8)
	) name7323 (
		\bdma_BEAD_reg[6]/NET0131 ,
		_w7303_,
		_w11370_
	);
	LUT2 #(
		.INIT('h8)
	) name7324 (
		\bdma_BCTL_reg[6]/NET0131 ,
		_w7230_,
		_w11371_
	);
	LUT2 #(
		.INIT('h8)
	) name7325 (
		\pio_PINT_reg[6]/NET0131 ,
		_w7271_,
		_w11372_
	);
	LUT2 #(
		.INIT('h8)
	) name7326 (
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w7281_,
		_w11373_
	);
	LUT2 #(
		.INIT('h8)
	) name7327 (
		\PIO_out[6]_pad ,
		_w7291_,
		_w11374_
	);
	LUT2 #(
		.INIT('h8)
	) name7328 (
		\PIO_oe[6]_pad ,
		_w7244_,
		_w11375_
	);
	LUT2 #(
		.INIT('h8)
	) name7329 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w7299_,
		_w11376_
	);
	LUT2 #(
		.INIT('h1)
	) name7330 (
		_w7522_,
		_w11349_,
		_w11377_
	);
	LUT2 #(
		.INIT('h1)
	) name7331 (
		_w11350_,
		_w11351_,
		_w11378_
	);
	LUT2 #(
		.INIT('h1)
	) name7332 (
		_w11353_,
		_w11354_,
		_w11379_
	);
	LUT2 #(
		.INIT('h1)
	) name7333 (
		_w11355_,
		_w11356_,
		_w11380_
	);
	LUT2 #(
		.INIT('h1)
	) name7334 (
		_w11357_,
		_w11358_,
		_w11381_
	);
	LUT2 #(
		.INIT('h1)
	) name7335 (
		_w11359_,
		_w11360_,
		_w11382_
	);
	LUT2 #(
		.INIT('h1)
	) name7336 (
		_w11361_,
		_w11363_,
		_w11383_
	);
	LUT2 #(
		.INIT('h1)
	) name7337 (
		_w11364_,
		_w11365_,
		_w11384_
	);
	LUT2 #(
		.INIT('h1)
	) name7338 (
		_w11366_,
		_w11368_,
		_w11385_
	);
	LUT2 #(
		.INIT('h1)
	) name7339 (
		_w11369_,
		_w11372_,
		_w11386_
	);
	LUT2 #(
		.INIT('h1)
	) name7340 (
		_w11373_,
		_w11374_,
		_w11387_
	);
	LUT2 #(
		.INIT('h1)
	) name7341 (
		_w11375_,
		_w11376_,
		_w11388_
	);
	LUT2 #(
		.INIT('h8)
	) name7342 (
		_w11387_,
		_w11388_,
		_w11389_
	);
	LUT2 #(
		.INIT('h8)
	) name7343 (
		_w11385_,
		_w11386_,
		_w11390_
	);
	LUT2 #(
		.INIT('h8)
	) name7344 (
		_w11383_,
		_w11384_,
		_w11391_
	);
	LUT2 #(
		.INIT('h8)
	) name7345 (
		_w11381_,
		_w11382_,
		_w11392_
	);
	LUT2 #(
		.INIT('h8)
	) name7346 (
		_w11379_,
		_w11380_,
		_w11393_
	);
	LUT2 #(
		.INIT('h8)
	) name7347 (
		_w11377_,
		_w11378_,
		_w11394_
	);
	LUT2 #(
		.INIT('h8)
	) name7348 (
		_w11393_,
		_w11394_,
		_w11395_
	);
	LUT2 #(
		.INIT('h8)
	) name7349 (
		_w11391_,
		_w11392_,
		_w11396_
	);
	LUT2 #(
		.INIT('h8)
	) name7350 (
		_w11389_,
		_w11390_,
		_w11397_
	);
	LUT2 #(
		.INIT('h8)
	) name7351 (
		_w11396_,
		_w11397_,
		_w11398_
	);
	LUT2 #(
		.INIT('h4)
	) name7352 (
		_w11362_,
		_w11395_,
		_w11399_
	);
	LUT2 #(
		.INIT('h1)
	) name7353 (
		_w11370_,
		_w11371_,
		_w11400_
	);
	LUT2 #(
		.INIT('h8)
	) name7354 (
		_w11399_,
		_w11400_,
		_w11401_
	);
	LUT2 #(
		.INIT('h4)
	) name7355 (
		_w11352_,
		_w11398_,
		_w11402_
	);
	LUT2 #(
		.INIT('h4)
	) name7356 (
		_w11367_,
		_w11402_,
		_w11403_
	);
	LUT2 #(
		.INIT('h8)
	) name7357 (
		_w11401_,
		_w11403_,
		_w11404_
	);
	LUT2 #(
		.INIT('h2)
	) name7358 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w11404_,
		_w11405_
	);
	LUT2 #(
		.INIT('h8)
	) name7359 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w11406_
	);
	LUT2 #(
		.INIT('h2)
	) name7360 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4392_,
		_w11407_
	);
	LUT2 #(
		.INIT('h2)
	) name7361 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w7216_,
		_w11408_
	);
	LUT2 #(
		.INIT('h8)
	) name7362 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w11409_
	);
	LUT2 #(
		.INIT('h8)
	) name7363 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w11410_
	);
	LUT2 #(
		.INIT('h8)
	) name7364 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w11411_
	);
	LUT2 #(
		.INIT('h8)
	) name7365 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		\core_c_psq_SSTAT_reg[6]/NET0131 ,
		_w11412_
	);
	LUT2 #(
		.INIT('h8)
	) name7366 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		_w11413_
	);
	LUT2 #(
		.INIT('h1)
	) name7367 (
		_w11406_,
		_w11409_,
		_w11414_
	);
	LUT2 #(
		.INIT('h1)
	) name7368 (
		_w11410_,
		_w11411_,
		_w11415_
	);
	LUT2 #(
		.INIT('h1)
	) name7369 (
		_w11412_,
		_w11413_,
		_w11416_
	);
	LUT2 #(
		.INIT('h8)
	) name7370 (
		_w11415_,
		_w11416_,
		_w11417_
	);
	LUT2 #(
		.INIT('h4)
	) name7371 (
		_w11408_,
		_w11414_,
		_w11418_
	);
	LUT2 #(
		.INIT('h8)
	) name7372 (
		_w11417_,
		_w11418_,
		_w11419_
	);
	LUT2 #(
		.INIT('h4)
	) name7373 (
		_w11407_,
		_w11419_,
		_w11420_
	);
	LUT2 #(
		.INIT('h2)
	) name7374 (
		_w7215_,
		_w11420_,
		_w11421_
	);
	LUT2 #(
		.INIT('h4)
	) name7375 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 ,
		_w11422_
	);
	LUT2 #(
		.INIT('h8)
	) name7376 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001 ,
		_w11423_
	);
	LUT2 #(
		.INIT('h1)
	) name7377 (
		_w11422_,
		_w11423_,
		_w11424_
	);
	LUT2 #(
		.INIT('h2)
	) name7378 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w11424_,
		_w11425_
	);
	LUT2 #(
		.INIT('h4)
	) name7379 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001 ,
		_w11426_
	);
	LUT2 #(
		.INIT('h8)
	) name7380 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001 ,
		_w11427_
	);
	LUT2 #(
		.INIT('h1)
	) name7381 (
		_w11426_,
		_w11427_,
		_w11428_
	);
	LUT2 #(
		.INIT('h2)
	) name7382 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w11428_,
		_w11429_
	);
	LUT2 #(
		.INIT('h4)
	) name7383 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001 ,
		_w11430_
	);
	LUT2 #(
		.INIT('h8)
	) name7384 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001 ,
		_w11431_
	);
	LUT2 #(
		.INIT('h1)
	) name7385 (
		_w11430_,
		_w11431_,
		_w11432_
	);
	LUT2 #(
		.INIT('h2)
	) name7386 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w11432_,
		_w11433_
	);
	LUT2 #(
		.INIT('h4)
	) name7387 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001 ,
		_w11434_
	);
	LUT2 #(
		.INIT('h8)
	) name7388 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001 ,
		_w11435_
	);
	LUT2 #(
		.INIT('h1)
	) name7389 (
		_w11434_,
		_w11435_,
		_w11436_
	);
	LUT2 #(
		.INIT('h2)
	) name7390 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w11436_,
		_w11437_
	);
	LUT2 #(
		.INIT('h4)
	) name7391 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001 ,
		_w11438_
	);
	LUT2 #(
		.INIT('h8)
	) name7392 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001 ,
		_w11439_
	);
	LUT2 #(
		.INIT('h1)
	) name7393 (
		_w11438_,
		_w11439_,
		_w11440_
	);
	LUT2 #(
		.INIT('h2)
	) name7394 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w11440_,
		_w11441_
	);
	LUT2 #(
		.INIT('h4)
	) name7395 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001 ,
		_w11442_
	);
	LUT2 #(
		.INIT('h8)
	) name7396 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 ,
		_w11443_
	);
	LUT2 #(
		.INIT('h1)
	) name7397 (
		_w11442_,
		_w11443_,
		_w11444_
	);
	LUT2 #(
		.INIT('h2)
	) name7398 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w11444_,
		_w11445_
	);
	LUT2 #(
		.INIT('h4)
	) name7399 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001 ,
		_w11446_
	);
	LUT2 #(
		.INIT('h8)
	) name7400 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 ,
		_w11447_
	);
	LUT2 #(
		.INIT('h1)
	) name7401 (
		_w11446_,
		_w11447_,
		_w11448_
	);
	LUT2 #(
		.INIT('h2)
	) name7402 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w11448_,
		_w11449_
	);
	LUT2 #(
		.INIT('h1)
	) name7403 (
		_w11425_,
		_w11429_,
		_w11450_
	);
	LUT2 #(
		.INIT('h1)
	) name7404 (
		_w11433_,
		_w11437_,
		_w11451_
	);
	LUT2 #(
		.INIT('h1)
	) name7405 (
		_w11441_,
		_w11445_,
		_w11452_
	);
	LUT2 #(
		.INIT('h4)
	) name7406 (
		_w11449_,
		_w11452_,
		_w11453_
	);
	LUT2 #(
		.INIT('h8)
	) name7407 (
		_w11450_,
		_w11451_,
		_w11454_
	);
	LUT2 #(
		.INIT('h8)
	) name7408 (
		_w11453_,
		_w11454_,
		_w11455_
	);
	LUT2 #(
		.INIT('h2)
	) name7409 (
		_w7179_,
		_w11455_,
		_w11456_
	);
	LUT2 #(
		.INIT('h8)
	) name7410 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 ,
		_w11457_
	);
	LUT2 #(
		.INIT('h8)
	) name7411 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		_w11458_
	);
	LUT2 #(
		.INIT('h8)
	) name7412 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 ,
		_w11459_
	);
	LUT2 #(
		.INIT('h8)
	) name7413 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 ,
		_w11460_
	);
	LUT2 #(
		.INIT('h8)
	) name7414 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131 ,
		_w11461_
	);
	LUT2 #(
		.INIT('h8)
	) name7415 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131 ,
		_w11462_
	);
	LUT2 #(
		.INIT('h8)
	) name7416 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		\core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131 ,
		_w11463_
	);
	LUT2 #(
		.INIT('h8)
	) name7417 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131 ,
		_w11464_
	);
	LUT2 #(
		.INIT('h8)
	) name7418 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131 ,
		_w11465_
	);
	LUT2 #(
		.INIT('h8)
	) name7419 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		\core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131 ,
		_w11466_
	);
	LUT2 #(
		.INIT('h8)
	) name7420 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		\core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131 ,
		_w11467_
	);
	LUT2 #(
		.INIT('h8)
	) name7421 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		\core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131 ,
		_w11468_
	);
	LUT2 #(
		.INIT('h1)
	) name7422 (
		_w11457_,
		_w11458_,
		_w11469_
	);
	LUT2 #(
		.INIT('h1)
	) name7423 (
		_w11459_,
		_w11460_,
		_w11470_
	);
	LUT2 #(
		.INIT('h1)
	) name7424 (
		_w11461_,
		_w11462_,
		_w11471_
	);
	LUT2 #(
		.INIT('h1)
	) name7425 (
		_w11463_,
		_w11464_,
		_w11472_
	);
	LUT2 #(
		.INIT('h1)
	) name7426 (
		_w11465_,
		_w11466_,
		_w11473_
	);
	LUT2 #(
		.INIT('h1)
	) name7427 (
		_w11467_,
		_w11468_,
		_w11474_
	);
	LUT2 #(
		.INIT('h8)
	) name7428 (
		_w11473_,
		_w11474_,
		_w11475_
	);
	LUT2 #(
		.INIT('h8)
	) name7429 (
		_w11471_,
		_w11472_,
		_w11476_
	);
	LUT2 #(
		.INIT('h8)
	) name7430 (
		_w11469_,
		_w11470_,
		_w11477_
	);
	LUT2 #(
		.INIT('h8)
	) name7431 (
		_w11476_,
		_w11477_,
		_w11478_
	);
	LUT2 #(
		.INIT('h8)
	) name7432 (
		_w11475_,
		_w11478_,
		_w11479_
	);
	LUT2 #(
		.INIT('h2)
	) name7433 (
		_w7068_,
		_w11479_,
		_w11480_
	);
	LUT2 #(
		.INIT('h8)
	) name7434 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131 ,
		_w11481_
	);
	LUT2 #(
		.INIT('h8)
	) name7435 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131 ,
		_w11482_
	);
	LUT2 #(
		.INIT('h8)
	) name7436 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131 ,
		_w11483_
	);
	LUT2 #(
		.INIT('h8)
	) name7437 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131 ,
		_w11484_
	);
	LUT2 #(
		.INIT('h8)
	) name7438 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131 ,
		_w11485_
	);
	LUT2 #(
		.INIT('h8)
	) name7439 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131 ,
		_w11486_
	);
	LUT2 #(
		.INIT('h8)
	) name7440 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131 ,
		_w11487_
	);
	LUT2 #(
		.INIT('h8)
	) name7441 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131 ,
		_w11488_
	);
	LUT2 #(
		.INIT('h8)
	) name7442 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w11489_
	);
	LUT2 #(
		.INIT('h8)
	) name7443 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w11490_
	);
	LUT2 #(
		.INIT('h8)
	) name7444 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		_w11491_
	);
	LUT2 #(
		.INIT('h8)
	) name7445 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w11492_
	);
	LUT2 #(
		.INIT('h1)
	) name7446 (
		_w11481_,
		_w11482_,
		_w11493_
	);
	LUT2 #(
		.INIT('h1)
	) name7447 (
		_w11483_,
		_w11484_,
		_w11494_
	);
	LUT2 #(
		.INIT('h1)
	) name7448 (
		_w11485_,
		_w11486_,
		_w11495_
	);
	LUT2 #(
		.INIT('h1)
	) name7449 (
		_w11487_,
		_w11488_,
		_w11496_
	);
	LUT2 #(
		.INIT('h1)
	) name7450 (
		_w11489_,
		_w11490_,
		_w11497_
	);
	LUT2 #(
		.INIT('h1)
	) name7451 (
		_w11491_,
		_w11492_,
		_w11498_
	);
	LUT2 #(
		.INIT('h8)
	) name7452 (
		_w11497_,
		_w11498_,
		_w11499_
	);
	LUT2 #(
		.INIT('h8)
	) name7453 (
		_w11495_,
		_w11496_,
		_w11500_
	);
	LUT2 #(
		.INIT('h8)
	) name7454 (
		_w11493_,
		_w11494_,
		_w11501_
	);
	LUT2 #(
		.INIT('h8)
	) name7455 (
		_w11500_,
		_w11501_,
		_w11502_
	);
	LUT2 #(
		.INIT('h8)
	) name7456 (
		_w11499_,
		_w11502_,
		_w11503_
	);
	LUT2 #(
		.INIT('h2)
	) name7457 (
		_w7128_,
		_w11503_,
		_w11504_
	);
	LUT2 #(
		.INIT('h8)
	) name7458 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[6]/P0001 ,
		_w11505_
	);
	LUT2 #(
		.INIT('h8)
	) name7459 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w11506_
	);
	LUT2 #(
		.INIT('h8)
	) name7460 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[6]/P0001 ,
		_w11507_
	);
	LUT2 #(
		.INIT('h8)
	) name7461 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w11508_
	);
	LUT2 #(
		.INIT('h1)
	) name7462 (
		_w11505_,
		_w11506_,
		_w11509_
	);
	LUT2 #(
		.INIT('h1)
	) name7463 (
		_w11507_,
		_w11508_,
		_w11510_
	);
	LUT2 #(
		.INIT('h8)
	) name7464 (
		_w11509_,
		_w11510_,
		_w11511_
	);
	LUT2 #(
		.INIT('h2)
	) name7465 (
		_w7119_,
		_w11511_,
		_w11512_
	);
	LUT2 #(
		.INIT('h1)
	) name7466 (
		_w11480_,
		_w11512_,
		_w11513_
	);
	LUT2 #(
		.INIT('h4)
	) name7467 (
		_w11504_,
		_w11513_,
		_w11514_
	);
	LUT2 #(
		.INIT('h1)
	) name7468 (
		_w11321_,
		_w11456_,
		_w11515_
	);
	LUT2 #(
		.INIT('h8)
	) name7469 (
		_w11514_,
		_w11515_,
		_w11516_
	);
	LUT2 #(
		.INIT('h4)
	) name7470 (
		_w11421_,
		_w11516_,
		_w11517_
	);
	LUT2 #(
		.INIT('h4)
	) name7471 (
		_w11405_,
		_w11517_,
		_w11518_
	);
	LUT2 #(
		.INIT('h4)
	) name7472 (
		_w11348_,
		_w11518_,
		_w11519_
	);
	LUT2 #(
		.INIT('h4)
	) name7473 (
		_w11300_,
		_w11519_,
		_w11520_
	);
	LUT2 #(
		.INIT('h1)
	) name7474 (
		\emc_DMDoe_reg/NET0131 ,
		_w11520_,
		_w11521_
	);
	LUT2 #(
		.INIT('h8)
	) name7475 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[6]/P0001 ,
		_w11522_
	);
	LUT2 #(
		.INIT('h2)
	) name7476 (
		_w7057_,
		_w11522_,
		_w11523_
	);
	LUT2 #(
		.INIT('h4)
	) name7477 (
		_w11521_,
		_w11523_,
		_w11524_
	);
	LUT2 #(
		.INIT('h1)
	) name7478 (
		_w11299_,
		_w11524_,
		_w11525_
	);
	LUT2 #(
		.INIT('h2)
	) name7479 (
		_w6135_,
		_w11525_,
		_w11526_
	);
	LUT2 #(
		.INIT('h2)
	) name7480 (
		_w8964_,
		_w11526_,
		_w11527_
	);
	LUT2 #(
		.INIT('h4)
	) name7481 (
		_w11281_,
		_w11527_,
		_w11528_
	);
	LUT2 #(
		.INIT('h1)
	) name7482 (
		_w11268_,
		_w11528_,
		_w11529_
	);
	LUT2 #(
		.INIT('h4)
	) name7483 (
		_w11030_,
		_w11529_,
		_w11530_
	);
	LUT2 #(
		.INIT('h1)
	) name7484 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w6924_,
		_w11531_
	);
	LUT2 #(
		.INIT('h8)
	) name7485 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131 ,
		_w6988_,
		_w11532_
	);
	LUT2 #(
		.INIT('h8)
	) name7486 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w6926_,
		_w11533_
	);
	LUT2 #(
		.INIT('h8)
	) name7487 (
		\core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 ,
		_w6972_,
		_w11534_
	);
	LUT2 #(
		.INIT('h8)
	) name7488 (
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w6976_,
		_w11535_
	);
	LUT2 #(
		.INIT('h8)
	) name7489 (
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w6974_,
		_w11536_
	);
	LUT2 #(
		.INIT('h8)
	) name7490 (
		\core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 ,
		_w6970_,
		_w11537_
	);
	LUT2 #(
		.INIT('h1)
	) name7491 (
		_w11534_,
		_w11535_,
		_w11538_
	);
	LUT2 #(
		.INIT('h1)
	) name7492 (
		_w11536_,
		_w11537_,
		_w11539_
	);
	LUT2 #(
		.INIT('h8)
	) name7493 (
		_w11538_,
		_w11539_,
		_w11540_
	);
	LUT2 #(
		.INIT('h2)
	) name7494 (
		_w4055_,
		_w11540_,
		_w11541_
	);
	LUT2 #(
		.INIT('h8)
	) name7495 (
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w6958_,
		_w11542_
	);
	LUT2 #(
		.INIT('h8)
	) name7496 (
		\core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 ,
		_w6960_,
		_w11543_
	);
	LUT2 #(
		.INIT('h8)
	) name7497 (
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w6962_,
		_w11544_
	);
	LUT2 #(
		.INIT('h8)
	) name7498 (
		\core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 ,
		_w6964_,
		_w11545_
	);
	LUT2 #(
		.INIT('h1)
	) name7499 (
		_w11542_,
		_w11543_,
		_w11546_
	);
	LUT2 #(
		.INIT('h1)
	) name7500 (
		_w11544_,
		_w11545_,
		_w11547_
	);
	LUT2 #(
		.INIT('h8)
	) name7501 (
		_w11546_,
		_w11547_,
		_w11548_
	);
	LUT2 #(
		.INIT('h4)
	) name7502 (
		_w11541_,
		_w11548_,
		_w11549_
	);
	LUT2 #(
		.INIT('h1)
	) name7503 (
		_w6121_,
		_w11549_,
		_w11550_
	);
	LUT2 #(
		.INIT('h8)
	) name7504 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w6956_,
		_w11551_
	);
	LUT2 #(
		.INIT('h4)
	) name7505 (
		_w6111_,
		_w11025_,
		_w11552_
	);
	LUT2 #(
		.INIT('h1)
	) name7506 (
		_w11550_,
		_w11551_,
		_w11553_
	);
	LUT2 #(
		.INIT('h4)
	) name7507 (
		_w11552_,
		_w11553_,
		_w11554_
	);
	LUT2 #(
		.INIT('h2)
	) name7508 (
		_w5949_,
		_w11554_,
		_w11555_
	);
	LUT2 #(
		.INIT('h2)
	) name7509 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		_w6934_,
		_w11556_
	);
	LUT2 #(
		.INIT('h1)
	) name7510 (
		_w11532_,
		_w11533_,
		_w11557_
	);
	LUT2 #(
		.INIT('h8)
	) name7511 (
		_w6924_,
		_w11557_,
		_w11558_
	);
	LUT2 #(
		.INIT('h4)
	) name7512 (
		_w11556_,
		_w11558_,
		_w11559_
	);
	LUT2 #(
		.INIT('h4)
	) name7513 (
		_w11555_,
		_w11559_,
		_w11560_
	);
	LUT2 #(
		.INIT('h1)
	) name7514 (
		_w6176_,
		_w11531_,
		_w11561_
	);
	LUT2 #(
		.INIT('h4)
	) name7515 (
		_w11560_,
		_w11561_,
		_w11562_
	);
	LUT2 #(
		.INIT('h8)
	) name7516 (
		_w6176_,
		_w10996_,
		_w11563_
	);
	LUT2 #(
		.INIT('h1)
	) name7517 (
		_w6135_,
		_w11563_,
		_w11564_
	);
	LUT2 #(
		.INIT('h4)
	) name7518 (
		_w11562_,
		_w11564_,
		_w11565_
	);
	LUT2 #(
		.INIT('h2)
	) name7519 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		_w6642_,
		_w11566_
	);
	LUT2 #(
		.INIT('h1)
	) name7520 (
		_w6695_,
		_w6731_,
		_w11567_
	);
	LUT2 #(
		.INIT('h8)
	) name7521 (
		_w6695_,
		_w6731_,
		_w11568_
	);
	LUT2 #(
		.INIT('h1)
	) name7522 (
		_w11567_,
		_w11568_,
		_w11569_
	);
	LUT2 #(
		.INIT('h4)
	) name7523 (
		_w8198_,
		_w11569_,
		_w11570_
	);
	LUT2 #(
		.INIT('h1)
	) name7524 (
		_w6743_,
		_w6779_,
		_w11571_
	);
	LUT2 #(
		.INIT('h4)
	) name7525 (
		_w6778_,
		_w10920_,
		_w11572_
	);
	LUT2 #(
		.INIT('h1)
	) name7526 (
		_w6753_,
		_w11572_,
		_w11573_
	);
	LUT2 #(
		.INIT('h1)
	) name7527 (
		_w11571_,
		_w11573_,
		_w11574_
	);
	LUT2 #(
		.INIT('h8)
	) name7528 (
		_w11571_,
		_w11573_,
		_w11575_
	);
	LUT2 #(
		.INIT('h1)
	) name7529 (
		_w11574_,
		_w11575_,
		_w11576_
	);
	LUT2 #(
		.INIT('h8)
	) name7530 (
		_w8198_,
		_w11576_,
		_w11577_
	);
	LUT2 #(
		.INIT('h1)
	) name7531 (
		_w11566_,
		_w11570_,
		_w11578_
	);
	LUT2 #(
		.INIT('h4)
	) name7532 (
		_w11577_,
		_w11578_,
		_w11579_
	);
	LUT2 #(
		.INIT('h1)
	) name7533 (
		_w6176_,
		_w11579_,
		_w11580_
	);
	LUT2 #(
		.INIT('h2)
	) name7534 (
		_w6176_,
		_w11280_,
		_w11581_
	);
	LUT2 #(
		.INIT('h2)
	) name7535 (
		_w6135_,
		_w11580_,
		_w11582_
	);
	LUT2 #(
		.INIT('h4)
	) name7536 (
		_w11581_,
		_w11582_,
		_w11583_
	);
	LUT2 #(
		.INIT('h1)
	) name7537 (
		_w7005_,
		_w11565_,
		_w11584_
	);
	LUT2 #(
		.INIT('h4)
	) name7538 (
		_w11583_,
		_w11584_,
		_w11585_
	);
	LUT2 #(
		.INIT('h2)
	) name7539 (
		_w6176_,
		_w11265_,
		_w11586_
	);
	LUT2 #(
		.INIT('h4)
	) name7540 (
		_w11025_,
		_w11549_,
		_w11587_
	);
	LUT2 #(
		.INIT('h4)
	) name7541 (
		_w6176_,
		_w11587_,
		_w11588_
	);
	LUT2 #(
		.INIT('h1)
	) name7542 (
		_w11586_,
		_w11588_,
		_w11589_
	);
	LUT2 #(
		.INIT('h2)
	) name7543 (
		_w6135_,
		_w11589_,
		_w11590_
	);
	LUT2 #(
		.INIT('h1)
	) name7544 (
		_w6176_,
		_w11525_,
		_w11591_
	);
	LUT2 #(
		.INIT('h1)
	) name7545 (
		_w10955_,
		_w11591_,
		_w11592_
	);
	LUT2 #(
		.INIT('h1)
	) name7546 (
		_w6135_,
		_w11592_,
		_w11593_
	);
	LUT2 #(
		.INIT('h2)
	) name7547 (
		_w7005_,
		_w11590_,
		_w11594_
	);
	LUT2 #(
		.INIT('h4)
	) name7548 (
		_w11593_,
		_w11594_,
		_w11595_
	);
	LUT2 #(
		.INIT('h1)
	) name7549 (
		_w11585_,
		_w11595_,
		_w11596_
	);
	LUT2 #(
		.INIT('h1)
	) name7550 (
		_w6176_,
		_w10911_,
		_w11597_
	);
	LUT2 #(
		.INIT('h1)
	) name7551 (
		_w10344_,
		_w11597_,
		_w11598_
	);
	LUT2 #(
		.INIT('h2)
	) name7552 (
		_w7005_,
		_w11598_,
		_w11599_
	);
	LUT2 #(
		.INIT('h8)
	) name7553 (
		_w6176_,
		_w10386_,
		_w11600_
	);
	LUT2 #(
		.INIT('h8)
	) name7554 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w6926_,
		_w11601_
	);
	LUT2 #(
		.INIT('h2)
	) name7555 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		_w6934_,
		_w11602_
	);
	LUT2 #(
		.INIT('h8)
	) name7556 (
		\core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 ,
		_w6972_,
		_w11603_
	);
	LUT2 #(
		.INIT('h8)
	) name7557 (
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		_w6976_,
		_w11604_
	);
	LUT2 #(
		.INIT('h8)
	) name7558 (
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w6974_,
		_w11605_
	);
	LUT2 #(
		.INIT('h8)
	) name7559 (
		\core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 ,
		_w6970_,
		_w11606_
	);
	LUT2 #(
		.INIT('h1)
	) name7560 (
		_w11603_,
		_w11604_,
		_w11607_
	);
	LUT2 #(
		.INIT('h1)
	) name7561 (
		_w11605_,
		_w11606_,
		_w11608_
	);
	LUT2 #(
		.INIT('h8)
	) name7562 (
		_w11607_,
		_w11608_,
		_w11609_
	);
	LUT2 #(
		.INIT('h2)
	) name7563 (
		_w4055_,
		_w11609_,
		_w11610_
	);
	LUT2 #(
		.INIT('h8)
	) name7564 (
		\core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 ,
		_w6960_,
		_w11611_
	);
	LUT2 #(
		.INIT('h8)
	) name7565 (
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		_w6958_,
		_w11612_
	);
	LUT2 #(
		.INIT('h8)
	) name7566 (
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w6962_,
		_w11613_
	);
	LUT2 #(
		.INIT('h8)
	) name7567 (
		\core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 ,
		_w6964_,
		_w11614_
	);
	LUT2 #(
		.INIT('h1)
	) name7568 (
		_w11611_,
		_w11612_,
		_w11615_
	);
	LUT2 #(
		.INIT('h1)
	) name7569 (
		_w11613_,
		_w11614_,
		_w11616_
	);
	LUT2 #(
		.INIT('h8)
	) name7570 (
		_w11615_,
		_w11616_,
		_w11617_
	);
	LUT2 #(
		.INIT('h4)
	) name7571 (
		_w11610_,
		_w11617_,
		_w11618_
	);
	LUT2 #(
		.INIT('h1)
	) name7572 (
		_w6121_,
		_w11618_,
		_w11619_
	);
	LUT2 #(
		.INIT('h8)
	) name7573 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w6956_,
		_w11620_
	);
	LUT2 #(
		.INIT('h4)
	) name7574 (
		_w6111_,
		_w10416_,
		_w11621_
	);
	LUT2 #(
		.INIT('h1)
	) name7575 (
		_w11619_,
		_w11620_,
		_w11622_
	);
	LUT2 #(
		.INIT('h4)
	) name7576 (
		_w11621_,
		_w11622_,
		_w11623_
	);
	LUT2 #(
		.INIT('h2)
	) name7577 (
		_w5949_,
		_w11623_,
		_w11624_
	);
	LUT2 #(
		.INIT('h8)
	) name7578 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131 ,
		_w6988_,
		_w11625_
	);
	LUT2 #(
		.INIT('h1)
	) name7579 (
		_w11601_,
		_w11625_,
		_w11626_
	);
	LUT2 #(
		.INIT('h4)
	) name7580 (
		_w11602_,
		_w11626_,
		_w11627_
	);
	LUT2 #(
		.INIT('h4)
	) name7581 (
		_w11624_,
		_w11627_,
		_w11628_
	);
	LUT2 #(
		.INIT('h2)
	) name7582 (
		_w6924_,
		_w11628_,
		_w11629_
	);
	LUT2 #(
		.INIT('h2)
	) name7583 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w6924_,
		_w11630_
	);
	LUT2 #(
		.INIT('h1)
	) name7584 (
		_w11629_,
		_w11630_,
		_w11631_
	);
	LUT2 #(
		.INIT('h1)
	) name7585 (
		_w6176_,
		_w11631_,
		_w11632_
	);
	LUT2 #(
		.INIT('h1)
	) name7586 (
		_w7005_,
		_w11600_,
		_w11633_
	);
	LUT2 #(
		.INIT('h4)
	) name7587 (
		_w11632_,
		_w11633_,
		_w11634_
	);
	LUT2 #(
		.INIT('h1)
	) name7588 (
		_w11599_,
		_w11634_,
		_w11635_
	);
	LUT2 #(
		.INIT('h1)
	) name7589 (
		_w6135_,
		_w11635_,
		_w11636_
	);
	LUT2 #(
		.INIT('h2)
	) name7590 (
		_w6176_,
		_w10638_,
		_w11637_
	);
	LUT2 #(
		.INIT('h4)
	) name7591 (
		_w10416_,
		_w11618_,
		_w11638_
	);
	LUT2 #(
		.INIT('h4)
	) name7592 (
		_w6176_,
		_w11638_,
		_w11639_
	);
	LUT2 #(
		.INIT('h1)
	) name7593 (
		_w11637_,
		_w11639_,
		_w11640_
	);
	LUT2 #(
		.INIT('h2)
	) name7594 (
		_w7005_,
		_w11640_,
		_w11641_
	);
	LUT2 #(
		.INIT('h2)
	) name7595 (
		_w6176_,
		_w10663_,
		_w11642_
	);
	LUT2 #(
		.INIT('h2)
	) name7596 (
		\core_dag_ilm2reg_I_reg[8]/NET0131 ,
		_w6635_,
		_w11643_
	);
	LUT2 #(
		.INIT('h1)
	) name7597 (
		_w6697_,
		_w6841_,
		_w11644_
	);
	LUT2 #(
		.INIT('h8)
	) name7598 (
		_w6697_,
		_w6841_,
		_w11645_
	);
	LUT2 #(
		.INIT('h1)
	) name7599 (
		_w11644_,
		_w11645_,
		_w11646_
	);
	LUT2 #(
		.INIT('h4)
	) name7600 (
		_w8198_,
		_w11646_,
		_w11647_
	);
	LUT2 #(
		.INIT('h1)
	) name7601 (
		_w6845_,
		_w6873_,
		_w11648_
	);
	LUT2 #(
		.INIT('h2)
	) name7602 (
		_w6825_,
		_w11648_,
		_w11649_
	);
	LUT2 #(
		.INIT('h4)
	) name7603 (
		_w6825_,
		_w11648_,
		_w11650_
	);
	LUT2 #(
		.INIT('h1)
	) name7604 (
		_w11649_,
		_w11650_,
		_w11651_
	);
	LUT2 #(
		.INIT('h8)
	) name7605 (
		_w8198_,
		_w11651_,
		_w11652_
	);
	LUT2 #(
		.INIT('h1)
	) name7606 (
		_w11643_,
		_w11647_,
		_w11653_
	);
	LUT2 #(
		.INIT('h4)
	) name7607 (
		_w11652_,
		_w11653_,
		_w11654_
	);
	LUT2 #(
		.INIT('h1)
	) name7608 (
		_w6176_,
		_w11654_,
		_w11655_
	);
	LUT2 #(
		.INIT('h1)
	) name7609 (
		_w7005_,
		_w11642_,
		_w11656_
	);
	LUT2 #(
		.INIT('h4)
	) name7610 (
		_w11655_,
		_w11656_,
		_w11657_
	);
	LUT2 #(
		.INIT('h1)
	) name7611 (
		_w11641_,
		_w11657_,
		_w11658_
	);
	LUT2 #(
		.INIT('h2)
	) name7612 (
		_w6135_,
		_w11658_,
		_w11659_
	);
	LUT2 #(
		.INIT('h1)
	) name7613 (
		_w11636_,
		_w11659_,
		_w11660_
	);
	LUT2 #(
		.INIT('h8)
	) name7614 (
		_w7863_,
		_w10069_,
		_w11661_
	);
	LUT2 #(
		.INIT('h8)
	) name7615 (
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w6970_,
		_w11662_
	);
	LUT2 #(
		.INIT('h8)
	) name7616 (
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w6972_,
		_w11663_
	);
	LUT2 #(
		.INIT('h8)
	) name7617 (
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w6974_,
		_w11664_
	);
	LUT2 #(
		.INIT('h8)
	) name7618 (
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w6976_,
		_w11665_
	);
	LUT2 #(
		.INIT('h1)
	) name7619 (
		_w11662_,
		_w11663_,
		_w11666_
	);
	LUT2 #(
		.INIT('h1)
	) name7620 (
		_w11664_,
		_w11665_,
		_w11667_
	);
	LUT2 #(
		.INIT('h8)
	) name7621 (
		_w11666_,
		_w11667_,
		_w11668_
	);
	LUT2 #(
		.INIT('h2)
	) name7622 (
		_w4055_,
		_w11668_,
		_w11669_
	);
	LUT2 #(
		.INIT('h8)
	) name7623 (
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w6958_,
		_w11670_
	);
	LUT2 #(
		.INIT('h8)
	) name7624 (
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w6960_,
		_w11671_
	);
	LUT2 #(
		.INIT('h8)
	) name7625 (
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w6962_,
		_w11672_
	);
	LUT2 #(
		.INIT('h8)
	) name7626 (
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w6964_,
		_w11673_
	);
	LUT2 #(
		.INIT('h1)
	) name7627 (
		_w11670_,
		_w11671_,
		_w11674_
	);
	LUT2 #(
		.INIT('h1)
	) name7628 (
		_w11672_,
		_w11673_,
		_w11675_
	);
	LUT2 #(
		.INIT('h8)
	) name7629 (
		_w11674_,
		_w11675_,
		_w11676_
	);
	LUT2 #(
		.INIT('h4)
	) name7630 (
		_w11669_,
		_w11676_,
		_w11677_
	);
	LUT2 #(
		.INIT('h4)
	) name7631 (
		_w9735_,
		_w11677_,
		_w11678_
	);
	LUT2 #(
		.INIT('h2)
	) name7632 (
		_w8153_,
		_w11678_,
		_w11679_
	);
	LUT2 #(
		.INIT('h4)
	) name7633 (
		_w6135_,
		_w9752_,
		_w11680_
	);
	LUT2 #(
		.INIT('h2)
	) name7634 (
		_w6135_,
		_w10289_,
		_w11681_
	);
	LUT2 #(
		.INIT('h2)
	) name7635 (
		_w6176_,
		_w11681_,
		_w11682_
	);
	LUT2 #(
		.INIT('h4)
	) name7636 (
		_w11680_,
		_w11682_,
		_w11683_
	);
	LUT2 #(
		.INIT('h1)
	) name7637 (
		_w11661_,
		_w11679_,
		_w11684_
	);
	LUT2 #(
		.INIT('h4)
	) name7638 (
		_w11683_,
		_w11684_,
		_w11685_
	);
	LUT2 #(
		.INIT('h2)
	) name7639 (
		_w7005_,
		_w11685_,
		_w11686_
	);
	LUT2 #(
		.INIT('h8)
	) name7640 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131 ,
		_w6988_,
		_w11687_
	);
	LUT2 #(
		.INIT('h8)
	) name7641 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w6926_,
		_w11688_
	);
	LUT2 #(
		.INIT('h2)
	) name7642 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		_w6934_,
		_w11689_
	);
	LUT2 #(
		.INIT('h4)
	) name7643 (
		_w6111_,
		_w9735_,
		_w11690_
	);
	LUT2 #(
		.INIT('h1)
	) name7644 (
		_w6121_,
		_w11677_,
		_w11691_
	);
	LUT2 #(
		.INIT('h8)
	) name7645 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		_w6956_,
		_w11692_
	);
	LUT2 #(
		.INIT('h1)
	) name7646 (
		_w11690_,
		_w11692_,
		_w11693_
	);
	LUT2 #(
		.INIT('h4)
	) name7647 (
		_w11691_,
		_w11693_,
		_w11694_
	);
	LUT2 #(
		.INIT('h2)
	) name7648 (
		_w5949_,
		_w11694_,
		_w11695_
	);
	LUT2 #(
		.INIT('h1)
	) name7649 (
		_w11687_,
		_w11688_,
		_w11696_
	);
	LUT2 #(
		.INIT('h4)
	) name7650 (
		_w11689_,
		_w11696_,
		_w11697_
	);
	LUT2 #(
		.INIT('h4)
	) name7651 (
		_w11695_,
		_w11697_,
		_w11698_
	);
	LUT2 #(
		.INIT('h2)
	) name7652 (
		_w6924_,
		_w11698_,
		_w11699_
	);
	LUT2 #(
		.INIT('h2)
	) name7653 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w6924_,
		_w11700_
	);
	LUT2 #(
		.INIT('h1)
	) name7654 (
		_w6176_,
		_w11700_,
		_w11701_
	);
	LUT2 #(
		.INIT('h4)
	) name7655 (
		_w11699_,
		_w11701_,
		_w11702_
	);
	LUT2 #(
		.INIT('h2)
	) name7656 (
		_w6176_,
		_w9788_,
		_w11703_
	);
	LUT2 #(
		.INIT('h1)
	) name7657 (
		_w6135_,
		_w11703_,
		_w11704_
	);
	LUT2 #(
		.INIT('h4)
	) name7658 (
		_w11702_,
		_w11704_,
		_w11705_
	);
	LUT2 #(
		.INIT('h2)
	) name7659 (
		\core_dag_ilm2reg_I_reg[9]/NET0131 ,
		_w6630_,
		_w11706_
	);
	LUT2 #(
		.INIT('h1)
	) name7660 (
		_w6838_,
		_w6872_,
		_w11707_
	);
	LUT2 #(
		.INIT('h1)
	) name7661 (
		_w6825_,
		_w6845_,
		_w11708_
	);
	LUT2 #(
		.INIT('h1)
	) name7662 (
		_w6873_,
		_w11708_,
		_w11709_
	);
	LUT2 #(
		.INIT('h2)
	) name7663 (
		_w11707_,
		_w11709_,
		_w11710_
	);
	LUT2 #(
		.INIT('h4)
	) name7664 (
		_w11707_,
		_w11709_,
		_w11711_
	);
	LUT2 #(
		.INIT('h1)
	) name7665 (
		_w11710_,
		_w11711_,
		_w11712_
	);
	LUT2 #(
		.INIT('h8)
	) name7666 (
		_w8198_,
		_w11712_,
		_w11713_
	);
	LUT2 #(
		.INIT('h1)
	) name7667 (
		_w6698_,
		_w6703_,
		_w11714_
	);
	LUT2 #(
		.INIT('h2)
	) name7668 (
		_w6826_,
		_w11714_,
		_w11715_
	);
	LUT2 #(
		.INIT('h4)
	) name7669 (
		_w6826_,
		_w11714_,
		_w11716_
	);
	LUT2 #(
		.INIT('h1)
	) name7670 (
		_w11715_,
		_w11716_,
		_w11717_
	);
	LUT2 #(
		.INIT('h4)
	) name7671 (
		_w8198_,
		_w11717_,
		_w11718_
	);
	LUT2 #(
		.INIT('h1)
	) name7672 (
		_w11706_,
		_w11713_,
		_w11719_
	);
	LUT2 #(
		.INIT('h4)
	) name7673 (
		_w11718_,
		_w11719_,
		_w11720_
	);
	LUT2 #(
		.INIT('h4)
	) name7674 (
		_w6176_,
		_w11720_,
		_w11721_
	);
	LUT2 #(
		.INIT('h2)
	) name7675 (
		_w6135_,
		_w11721_,
		_w11722_
	);
	LUT2 #(
		.INIT('h4)
	) name7676 (
		_w10303_,
		_w11722_,
		_w11723_
	);
	LUT2 #(
		.INIT('h1)
	) name7677 (
		_w11705_,
		_w11723_,
		_w11724_
	);
	LUT2 #(
		.INIT('h1)
	) name7678 (
		_w7005_,
		_w11724_,
		_w11725_
	);
	LUT2 #(
		.INIT('h1)
	) name7679 (
		_w11686_,
		_w11725_,
		_w11726_
	);
	LUT2 #(
		.INIT('h1)
	) name7680 (
		_w9440_,
		_w9513_,
		_w11727_
	);
	LUT2 #(
		.INIT('h1)
	) name7681 (
		_w10916_,
		_w11530_,
		_w11728_
	);
	LUT2 #(
		.INIT('h4)
	) name7682 (
		_w11596_,
		_w11728_,
		_w11729_
	);
	LUT2 #(
		.INIT('h4)
	) name7683 (
		_w8230_,
		_w11727_,
		_w11730_
	);
	LUT2 #(
		.INIT('h4)
	) name7684 (
		_w8835_,
		_w11660_,
		_w11731_
	);
	LUT2 #(
		.INIT('h4)
	) name7685 (
		_w11726_,
		_w11731_,
		_w11732_
	);
	LUT2 #(
		.INIT('h8)
	) name7686 (
		_w11729_,
		_w11730_,
		_w11733_
	);
	LUT2 #(
		.INIT('h8)
	) name7687 (
		_w11732_,
		_w11733_,
		_w11734_
	);
	LUT2 #(
		.INIT('h1)
	) name7688 (
		_w9513_,
		_w11734_,
		_w11735_
	);
	LUT2 #(
		.INIT('h8)
	) name7689 (
		\memc_Dwrite_C_reg/NET0131 ,
		_w5950_,
		_w11736_
	);
	LUT2 #(
		.INIT('h4)
	) name7690 (
		_w5950_,
		_w6932_,
		_w11737_
	);
	LUT2 #(
		.INIT('h1)
	) name7691 (
		_w11736_,
		_w11737_,
		_w11738_
	);
	LUT2 #(
		.INIT('h8)
	) name7692 (
		\memc_Dread_E_reg/NET0131 ,
		_w4117_,
		_w11739_
	);
	LUT2 #(
		.INIT('h1)
	) name7693 (
		\core_c_dec_Long_Cg_reg/P0001 ,
		\core_c_dec_Prderr_Cg_reg/NET0131 ,
		_w11740_
	);
	LUT2 #(
		.INIT('h8)
	) name7694 (
		_w5053_,
		_w11740_,
		_w11741_
	);
	LUT2 #(
		.INIT('h4)
	) name7695 (
		_w4117_,
		_w11741_,
		_w11742_
	);
	LUT2 #(
		.INIT('h4)
	) name7696 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w6120_,
		_w11743_
	);
	LUT2 #(
		.INIT('h4)
	) name7697 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w6108_,
		_w11744_
	);
	LUT2 #(
		.INIT('h8)
	) name7698 (
		_w6026_,
		_w6955_,
		_w11745_
	);
	LUT2 #(
		.INIT('h1)
	) name7699 (
		_w6023_,
		_w11745_,
		_w11746_
	);
	LUT2 #(
		.INIT('h4)
	) name7700 (
		_w11744_,
		_w11746_,
		_w11747_
	);
	LUT2 #(
		.INIT('h4)
	) name7701 (
		_w11743_,
		_w11747_,
		_w11748_
	);
	LUT2 #(
		.INIT('h2)
	) name7702 (
		_w11742_,
		_w11748_,
		_w11749_
	);
	LUT2 #(
		.INIT('h8)
	) name7703 (
		_w5948_,
		_w11749_,
		_w11750_
	);
	LUT2 #(
		.INIT('h1)
	) name7704 (
		_w11739_,
		_w11750_,
		_w11751_
	);
	LUT2 #(
		.INIT('h8)
	) name7705 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_RDcyc_reg/NET0131 ,
		_w11752_
	);
	LUT2 #(
		.INIT('h8)
	) name7706 (
		_w5068_,
		_w11752_,
		_w11753_
	);
	LUT2 #(
		.INIT('h1)
	) name7707 (
		_w4050_,
		_w5968_,
		_w11754_
	);
	LUT2 #(
		.INIT('h4)
	) name7708 (
		_w11753_,
		_w11754_,
		_w11755_
	);
	LUT2 #(
		.INIT('h4)
	) name7709 (
		_w6922_,
		_w11755_,
		_w11756_
	);
	LUT2 #(
		.INIT('h1)
	) name7710 (
		_w5718_,
		_w11756_,
		_w11757_
	);
	LUT2 #(
		.INIT('h2)
	) name7711 (
		_w11751_,
		_w11757_,
		_w11758_
	);
	LUT2 #(
		.INIT('h1)
	) name7712 (
		_w5966_,
		_w5970_,
		_w11759_
	);
	LUT2 #(
		.INIT('h1)
	) name7713 (
		_w5718_,
		_w11759_,
		_w11760_
	);
	LUT2 #(
		.INIT('h2)
	) name7714 (
		\idma_WRcyc_reg/NET0131 ,
		_w5718_,
		_w11761_
	);
	LUT2 #(
		.INIT('h8)
	) name7715 (
		_w6925_,
		_w11761_,
		_w11762_
	);
	LUT2 #(
		.INIT('h1)
	) name7716 (
		_w6918_,
		_w11762_,
		_w11763_
	);
	LUT2 #(
		.INIT('h4)
	) name7717 (
		_w11760_,
		_w11763_,
		_w11764_
	);
	LUT2 #(
		.INIT('h8)
	) name7718 (
		_w11738_,
		_w11764_,
		_w11765_
	);
	LUT2 #(
		.INIT('h8)
	) name7719 (
		_w11758_,
		_w11765_,
		_w11766_
	);
	LUT2 #(
		.INIT('h2)
	) name7720 (
		_w11735_,
		_w11766_,
		_w11767_
	);
	LUT2 #(
		.INIT('h8)
	) name7721 (
		\idma_DTMP_H_reg[0]/P0001 ,
		_w11762_,
		_w11768_
	);
	LUT2 #(
		.INIT('h1)
	) name7722 (
		_w4097_,
		_w11759_,
		_w11769_
	);
	LUT2 #(
		.INIT('h2)
	) name7723 (
		_w11763_,
		_w11769_,
		_w11770_
	);
	LUT2 #(
		.INIT('h4)
	) name7724 (
		_w7602_,
		_w11770_,
		_w11771_
	);
	LUT2 #(
		.INIT('h4)
	) name7725 (
		_w4097_,
		_w5966_,
		_w11772_
	);
	LUT2 #(
		.INIT('h8)
	) name7726 (
		\sport1_rxctl_RX_reg[0]/P0001 ,
		_w11772_,
		_w11773_
	);
	LUT2 #(
		.INIT('h4)
	) name7727 (
		_w4097_,
		_w5970_,
		_w11774_
	);
	LUT2 #(
		.INIT('h8)
	) name7728 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		_w11774_,
		_w11775_
	);
	LUT2 #(
		.INIT('h8)
	) name7729 (
		\bdma_BRdataBUF_reg[0]/P0001 ,
		_w6918_,
		_w11776_
	);
	LUT2 #(
		.INIT('h1)
	) name7730 (
		_w11773_,
		_w11775_,
		_w11777_
	);
	LUT2 #(
		.INIT('h4)
	) name7731 (
		_w11768_,
		_w11777_,
		_w11778_
	);
	LUT2 #(
		.INIT('h4)
	) name7732 (
		_w11776_,
		_w11778_,
		_w11779_
	);
	LUT2 #(
		.INIT('h4)
	) name7733 (
		_w11771_,
		_w11779_,
		_w11780_
	);
	LUT2 #(
		.INIT('h8)
	) name7734 (
		\idma_DTMP_H_reg[10]/P0001 ,
		_w11762_,
		_w11781_
	);
	LUT2 #(
		.INIT('h4)
	) name7735 (
		_w7854_,
		_w11770_,
		_w11782_
	);
	LUT2 #(
		.INIT('h8)
	) name7736 (
		\sport0_rxctl_RX_reg[10]/P0001 ,
		_w11774_,
		_w11783_
	);
	LUT2 #(
		.INIT('h8)
	) name7737 (
		\sport1_rxctl_RX_reg[10]/P0001 ,
		_w11772_,
		_w11784_
	);
	LUT2 #(
		.INIT('h8)
	) name7738 (
		\bdma_BRdataBUF_reg[10]/P0001 ,
		_w6918_,
		_w11785_
	);
	LUT2 #(
		.INIT('h1)
	) name7739 (
		_w11783_,
		_w11784_,
		_w11786_
	);
	LUT2 #(
		.INIT('h4)
	) name7740 (
		_w11781_,
		_w11786_,
		_w11787_
	);
	LUT2 #(
		.INIT('h4)
	) name7741 (
		_w11785_,
		_w11787_,
		_w11788_
	);
	LUT2 #(
		.INIT('h4)
	) name7742 (
		_w11782_,
		_w11788_,
		_w11789_
	);
	LUT2 #(
		.INIT('h8)
	) name7743 (
		\idma_DTMP_H_reg[11]/P0001 ,
		_w11762_,
		_w11790_
	);
	LUT2 #(
		.INIT('h4)
	) name7744 (
		_w8455_,
		_w11770_,
		_w11791_
	);
	LUT2 #(
		.INIT('h8)
	) name7745 (
		\sport1_rxctl_RX_reg[11]/P0001 ,
		_w11772_,
		_w11792_
	);
	LUT2 #(
		.INIT('h8)
	) name7746 (
		\sport0_rxctl_RX_reg[11]/P0001 ,
		_w11774_,
		_w11793_
	);
	LUT2 #(
		.INIT('h8)
	) name7747 (
		\bdma_BRdataBUF_reg[11]/P0001 ,
		_w6918_,
		_w11794_
	);
	LUT2 #(
		.INIT('h1)
	) name7748 (
		_w11792_,
		_w11793_,
		_w11795_
	);
	LUT2 #(
		.INIT('h4)
	) name7749 (
		_w11790_,
		_w11795_,
		_w11796_
	);
	LUT2 #(
		.INIT('h4)
	) name7750 (
		_w11794_,
		_w11796_,
		_w11797_
	);
	LUT2 #(
		.INIT('h4)
	) name7751 (
		_w11791_,
		_w11797_,
		_w11798_
	);
	LUT2 #(
		.INIT('h8)
	) name7752 (
		\idma_DTMP_H_reg[12]/P0001 ,
		_w11762_,
		_w11799_
	);
	LUT2 #(
		.INIT('h4)
	) name7753 (
		_w9173_,
		_w11770_,
		_w11800_
	);
	LUT2 #(
		.INIT('h8)
	) name7754 (
		\sport0_rxctl_RX_reg[12]/P0001 ,
		_w11774_,
		_w11801_
	);
	LUT2 #(
		.INIT('h8)
	) name7755 (
		\sport1_rxctl_RX_reg[12]/P0001 ,
		_w11772_,
		_w11802_
	);
	LUT2 #(
		.INIT('h8)
	) name7756 (
		\bdma_BRdataBUF_reg[12]/P0001 ,
		_w6918_,
		_w11803_
	);
	LUT2 #(
		.INIT('h1)
	) name7757 (
		_w11801_,
		_w11802_,
		_w11804_
	);
	LUT2 #(
		.INIT('h4)
	) name7758 (
		_w11799_,
		_w11804_,
		_w11805_
	);
	LUT2 #(
		.INIT('h4)
	) name7759 (
		_w11803_,
		_w11805_,
		_w11806_
	);
	LUT2 #(
		.INIT('h4)
	) name7760 (
		_w11800_,
		_w11806_,
		_w11807_
	);
	LUT2 #(
		.INIT('h8)
	) name7761 (
		\idma_DTMP_H_reg[13]/P0001 ,
		_w11762_,
		_w11808_
	);
	LUT2 #(
		.INIT('h4)
	) name7762 (
		_w7335_,
		_w11770_,
		_w11809_
	);
	LUT2 #(
		.INIT('h8)
	) name7763 (
		\sport0_rxctl_RX_reg[13]/P0001 ,
		_w11774_,
		_w11810_
	);
	LUT2 #(
		.INIT('h8)
	) name7764 (
		\sport1_rxctl_RX_reg[13]/P0001 ,
		_w11772_,
		_w11811_
	);
	LUT2 #(
		.INIT('h8)
	) name7765 (
		\bdma_BRdataBUF_reg[13]/P0001 ,
		_w6918_,
		_w11812_
	);
	LUT2 #(
		.INIT('h1)
	) name7766 (
		_w11810_,
		_w11811_,
		_w11813_
	);
	LUT2 #(
		.INIT('h4)
	) name7767 (
		_w11808_,
		_w11813_,
		_w11814_
	);
	LUT2 #(
		.INIT('h4)
	) name7768 (
		_w11812_,
		_w11814_,
		_w11815_
	);
	LUT2 #(
		.INIT('h4)
	) name7769 (
		_w11809_,
		_w11815_,
		_w11816_
	);
	LUT2 #(
		.INIT('h8)
	) name7770 (
		\idma_DTMP_H_reg[14]/P0001 ,
		_w11762_,
		_w11817_
	);
	LUT2 #(
		.INIT('h8)
	) name7771 (
		\regout_STD_C_reg[14]/P0001 ,
		_w6988_,
		_w11818_
	);
	LUT2 #(
		.INIT('h4)
	) name7772 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001 ,
		_w11819_
	);
	LUT2 #(
		.INIT('h8)
	) name7773 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001 ,
		_w11820_
	);
	LUT2 #(
		.INIT('h1)
	) name7774 (
		_w11819_,
		_w11820_,
		_w11821_
	);
	LUT2 #(
		.INIT('h2)
	) name7775 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w11821_,
		_w11822_
	);
	LUT2 #(
		.INIT('h4)
	) name7776 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001 ,
		_w11823_
	);
	LUT2 #(
		.INIT('h8)
	) name7777 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001 ,
		_w11824_
	);
	LUT2 #(
		.INIT('h1)
	) name7778 (
		_w11823_,
		_w11824_,
		_w11825_
	);
	LUT2 #(
		.INIT('h2)
	) name7779 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w11825_,
		_w11826_
	);
	LUT2 #(
		.INIT('h4)
	) name7780 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001 ,
		_w11827_
	);
	LUT2 #(
		.INIT('h8)
	) name7781 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001 ,
		_w11828_
	);
	LUT2 #(
		.INIT('h1)
	) name7782 (
		_w11827_,
		_w11828_,
		_w11829_
	);
	LUT2 #(
		.INIT('h2)
	) name7783 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w11829_,
		_w11830_
	);
	LUT2 #(
		.INIT('h4)
	) name7784 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001 ,
		_w11831_
	);
	LUT2 #(
		.INIT('h8)
	) name7785 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001 ,
		_w11832_
	);
	LUT2 #(
		.INIT('h1)
	) name7786 (
		_w11831_,
		_w11832_,
		_w11833_
	);
	LUT2 #(
		.INIT('h2)
	) name7787 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w11833_,
		_w11834_
	);
	LUT2 #(
		.INIT('h4)
	) name7788 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001 ,
		_w11835_
	);
	LUT2 #(
		.INIT('h8)
	) name7789 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001 ,
		_w11836_
	);
	LUT2 #(
		.INIT('h1)
	) name7790 (
		_w11835_,
		_w11836_,
		_w11837_
	);
	LUT2 #(
		.INIT('h2)
	) name7791 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w11837_,
		_w11838_
	);
	LUT2 #(
		.INIT('h1)
	) name7792 (
		_w11822_,
		_w11826_,
		_w11839_
	);
	LUT2 #(
		.INIT('h1)
	) name7793 (
		_w11830_,
		_w11834_,
		_w11840_
	);
	LUT2 #(
		.INIT('h4)
	) name7794 (
		_w11838_,
		_w11840_,
		_w11841_
	);
	LUT2 #(
		.INIT('h8)
	) name7795 (
		_w11839_,
		_w11841_,
		_w11842_
	);
	LUT2 #(
		.INIT('h2)
	) name7796 (
		_w7093_,
		_w11842_,
		_w11843_
	);
	LUT2 #(
		.INIT('h4)
	) name7797 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 ,
		_w11844_
	);
	LUT2 #(
		.INIT('h8)
	) name7798 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 ,
		_w11845_
	);
	LUT2 #(
		.INIT('h1)
	) name7799 (
		_w11844_,
		_w11845_,
		_w11846_
	);
	LUT2 #(
		.INIT('h2)
	) name7800 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w11846_,
		_w11847_
	);
	LUT2 #(
		.INIT('h4)
	) name7801 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001 ,
		_w11848_
	);
	LUT2 #(
		.INIT('h8)
	) name7802 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001 ,
		_w11849_
	);
	LUT2 #(
		.INIT('h1)
	) name7803 (
		_w11848_,
		_w11849_,
		_w11850_
	);
	LUT2 #(
		.INIT('h2)
	) name7804 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w11850_,
		_w11851_
	);
	LUT2 #(
		.INIT('h4)
	) name7805 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 ,
		_w11852_
	);
	LUT2 #(
		.INIT('h8)
	) name7806 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 ,
		_w11853_
	);
	LUT2 #(
		.INIT('h1)
	) name7807 (
		_w11852_,
		_w11853_,
		_w11854_
	);
	LUT2 #(
		.INIT('h2)
	) name7808 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w11854_,
		_w11855_
	);
	LUT2 #(
		.INIT('h1)
	) name7809 (
		_w11847_,
		_w11851_,
		_w11856_
	);
	LUT2 #(
		.INIT('h4)
	) name7810 (
		_w11855_,
		_w11856_,
		_w11857_
	);
	LUT2 #(
		.INIT('h8)
	) name7811 (
		_w7174_,
		_w11857_,
		_w11858_
	);
	LUT2 #(
		.INIT('h2)
	) name7812 (
		_w7153_,
		_w11858_,
		_w11859_
	);
	LUT2 #(
		.INIT('h4)
	) name7813 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001 ,
		_w11860_
	);
	LUT2 #(
		.INIT('h8)
	) name7814 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001 ,
		_w11861_
	);
	LUT2 #(
		.INIT('h1)
	) name7815 (
		_w11860_,
		_w11861_,
		_w11862_
	);
	LUT2 #(
		.INIT('h2)
	) name7816 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w11862_,
		_w11863_
	);
	LUT2 #(
		.INIT('h4)
	) name7817 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001 ,
		_w11864_
	);
	LUT2 #(
		.INIT('h8)
	) name7818 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001 ,
		_w11865_
	);
	LUT2 #(
		.INIT('h1)
	) name7819 (
		_w11864_,
		_w11865_,
		_w11866_
	);
	LUT2 #(
		.INIT('h2)
	) name7820 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w11866_,
		_w11867_
	);
	LUT2 #(
		.INIT('h4)
	) name7821 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001 ,
		_w11868_
	);
	LUT2 #(
		.INIT('h8)
	) name7822 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001 ,
		_w11869_
	);
	LUT2 #(
		.INIT('h1)
	) name7823 (
		_w11868_,
		_w11869_,
		_w11870_
	);
	LUT2 #(
		.INIT('h2)
	) name7824 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w11870_,
		_w11871_
	);
	LUT2 #(
		.INIT('h4)
	) name7825 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001 ,
		_w11872_
	);
	LUT2 #(
		.INIT('h8)
	) name7826 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001 ,
		_w11873_
	);
	LUT2 #(
		.INIT('h1)
	) name7827 (
		_w11872_,
		_w11873_,
		_w11874_
	);
	LUT2 #(
		.INIT('h2)
	) name7828 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w11874_,
		_w11875_
	);
	LUT2 #(
		.INIT('h4)
	) name7829 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001 ,
		_w11876_
	);
	LUT2 #(
		.INIT('h8)
	) name7830 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 ,
		_w11877_
	);
	LUT2 #(
		.INIT('h1)
	) name7831 (
		_w11876_,
		_w11877_,
		_w11878_
	);
	LUT2 #(
		.INIT('h2)
	) name7832 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w11878_,
		_w11879_
	);
	LUT2 #(
		.INIT('h4)
	) name7833 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001 ,
		_w11880_
	);
	LUT2 #(
		.INIT('h8)
	) name7834 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 ,
		_w11881_
	);
	LUT2 #(
		.INIT('h1)
	) name7835 (
		_w11880_,
		_w11881_,
		_w11882_
	);
	LUT2 #(
		.INIT('h2)
	) name7836 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w11882_,
		_w11883_
	);
	LUT2 #(
		.INIT('h1)
	) name7837 (
		_w7207_,
		_w11863_,
		_w11884_
	);
	LUT2 #(
		.INIT('h1)
	) name7838 (
		_w11867_,
		_w11871_,
		_w11885_
	);
	LUT2 #(
		.INIT('h1)
	) name7839 (
		_w11875_,
		_w11879_,
		_w11886_
	);
	LUT2 #(
		.INIT('h4)
	) name7840 (
		_w11883_,
		_w11886_,
		_w11887_
	);
	LUT2 #(
		.INIT('h8)
	) name7841 (
		_w11884_,
		_w11885_,
		_w11888_
	);
	LUT2 #(
		.INIT('h8)
	) name7842 (
		_w11887_,
		_w11888_,
		_w11889_
	);
	LUT2 #(
		.INIT('h2)
	) name7843 (
		_w7179_,
		_w11889_,
		_w11890_
	);
	LUT2 #(
		.INIT('h8)
	) name7844 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[14]/P0001 ,
		_w11891_
	);
	LUT2 #(
		.INIT('h8)
	) name7845 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[14]/P0001 ,
		_w11892_
	);
	LUT2 #(
		.INIT('h8)
	) name7846 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[14]/P0001 ,
		_w11893_
	);
	LUT2 #(
		.INIT('h8)
	) name7847 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[14]/P0001 ,
		_w11894_
	);
	LUT2 #(
		.INIT('h1)
	) name7848 (
		_w11891_,
		_w11892_,
		_w11895_
	);
	LUT2 #(
		.INIT('h1)
	) name7849 (
		_w11893_,
		_w11894_,
		_w11896_
	);
	LUT2 #(
		.INIT('h8)
	) name7850 (
		_w11895_,
		_w11896_,
		_w11897_
	);
	LUT2 #(
		.INIT('h2)
	) name7851 (
		_w7119_,
		_w11897_,
		_w11898_
	);
	LUT2 #(
		.INIT('h8)
	) name7852 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		\core_c_dec_imm14_E_reg/P0001 ,
		_w11899_
	);
	LUT2 #(
		.INIT('h8)
	) name7853 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w11900_
	);
	LUT2 #(
		.INIT('h8)
	) name7854 (
		\core_c_dec_IRE_reg[18]/NET0131 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w11901_
	);
	LUT2 #(
		.INIT('h1)
	) name7855 (
		_w11899_,
		_w11900_,
		_w11902_
	);
	LUT2 #(
		.INIT('h4)
	) name7856 (
		_w11901_,
		_w11902_,
		_w11903_
	);
	LUT2 #(
		.INIT('h2)
	) name7857 (
		_w7215_,
		_w11903_,
		_w11904_
	);
	LUT2 #(
		.INIT('h2)
	) name7858 (
		_w7068_,
		_w7078_,
		_w11905_
	);
	LUT2 #(
		.INIT('h2)
	) name7859 (
		_w7128_,
		_w7137_,
		_w11906_
	);
	LUT2 #(
		.INIT('h1)
	) name7860 (
		_w11905_,
		_w11906_,
		_w11907_
	);
	LUT2 #(
		.INIT('h8)
	) name7861 (
		\PIO_out[10]_pad ,
		_w7291_,
		_w11908_
	);
	LUT2 #(
		.INIT('h8)
	) name7862 (
		\pio_PINT_reg[10]/NET0131 ,
		_w7271_,
		_w11909_
	);
	LUT2 #(
		.INIT('h8)
	) name7863 (
		\ISCLK0_pad ,
		_w7249_,
		_w11910_
	);
	LUT2 #(
		.INIT('h8)
	) name7864 (
		\bdma_BCTL_reg[14]/NET0131 ,
		_w7230_,
		_w11911_
	);
	LUT2 #(
		.INIT('h8)
	) name7865 (
		\clkc_ckr_reg_DO_reg[14]/NET0131 ,
		_w7239_,
		_w11912_
	);
	LUT2 #(
		.INIT('h8)
	) name7866 (
		\idma_DCTL_reg[14]/NET0131 ,
		_w7299_,
		_w11913_
	);
	LUT2 #(
		.INIT('h8)
	) name7867 (
		\emc_WSCRreg_DO_reg[14]/NET0131 ,
		_w7251_,
		_w11914_
	);
	LUT2 #(
		.INIT('h8)
	) name7868 (
		\PIO_oe[10]_pad ,
		_w7244_,
		_w11915_
	);
	LUT2 #(
		.INIT('h8)
	) name7869 (
		\tm_TCR_TMP_reg[14]/NET0131 ,
		_w7289_,
		_w11916_
	);
	LUT2 #(
		.INIT('h8)
	) name7870 (
		\sport0_regs_AUTO_a_reg[14]/NET0131 ,
		_w7295_,
		_w11917_
	);
	LUT2 #(
		.INIT('h8)
	) name7871 (
		\ISCLK1_pad ,
		_w7281_,
		_w11918_
	);
	LUT2 #(
		.INIT('h8)
	) name7872 (
		\tm_tpr_reg_DO_reg[14]/NET0131 ,
		_w7293_,
		_w11919_
	);
	LUT2 #(
		.INIT('h8)
	) name7873 (
		\pio_pmask_reg_DO_reg[10]/NET0131 ,
		_w7297_,
		_w11920_
	);
	LUT2 #(
		.INIT('h8)
	) name7874 (
		\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w7247_,
		_w11921_
	);
	LUT2 #(
		.INIT('h8)
	) name7875 (
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w7273_,
		_w11922_
	);
	LUT2 #(
		.INIT('h8)
	) name7876 (
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w7259_,
		_w11923_
	);
	LUT2 #(
		.INIT('h8)
	) name7877 (
		PM_bdry_sel_pad,
		_w7522_,
		_w11924_
	);
	LUT2 #(
		.INIT('h8)
	) name7878 (
		\memc_usysr_DO_reg[14]/NET0131 ,
		_w7301_,
		_w11925_
	);
	LUT2 #(
		.INIT('h8)
	) name7879 (
		\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w7256_,
		_w11926_
	);
	LUT2 #(
		.INIT('h1)
	) name7880 (
		_w7689_,
		_w7710_,
		_w11927_
	);
	LUT2 #(
		.INIT('h1)
	) name7881 (
		_w11908_,
		_w11909_,
		_w11928_
	);
	LUT2 #(
		.INIT('h1)
	) name7882 (
		_w11910_,
		_w11912_,
		_w11929_
	);
	LUT2 #(
		.INIT('h1)
	) name7883 (
		_w11913_,
		_w11914_,
		_w11930_
	);
	LUT2 #(
		.INIT('h1)
	) name7884 (
		_w11915_,
		_w11916_,
		_w11931_
	);
	LUT2 #(
		.INIT('h1)
	) name7885 (
		_w11917_,
		_w11918_,
		_w11932_
	);
	LUT2 #(
		.INIT('h1)
	) name7886 (
		_w11919_,
		_w11920_,
		_w11933_
	);
	LUT2 #(
		.INIT('h1)
	) name7887 (
		_w11921_,
		_w11922_,
		_w11934_
	);
	LUT2 #(
		.INIT('h1)
	) name7888 (
		_w11923_,
		_w11924_,
		_w11935_
	);
	LUT2 #(
		.INIT('h1)
	) name7889 (
		_w11925_,
		_w11926_,
		_w11936_
	);
	LUT2 #(
		.INIT('h8)
	) name7890 (
		_w11935_,
		_w11936_,
		_w11937_
	);
	LUT2 #(
		.INIT('h8)
	) name7891 (
		_w11933_,
		_w11934_,
		_w11938_
	);
	LUT2 #(
		.INIT('h8)
	) name7892 (
		_w11931_,
		_w11932_,
		_w11939_
	);
	LUT2 #(
		.INIT('h8)
	) name7893 (
		_w11929_,
		_w11930_,
		_w11940_
	);
	LUT2 #(
		.INIT('h8)
	) name7894 (
		_w11927_,
		_w11928_,
		_w11941_
	);
	LUT2 #(
		.INIT('h8)
	) name7895 (
		_w11940_,
		_w11941_,
		_w11942_
	);
	LUT2 #(
		.INIT('h8)
	) name7896 (
		_w11938_,
		_w11939_,
		_w11943_
	);
	LUT2 #(
		.INIT('h8)
	) name7897 (
		_w11937_,
		_w11943_,
		_w11944_
	);
	LUT2 #(
		.INIT('h4)
	) name7898 (
		_w11911_,
		_w11942_,
		_w11945_
	);
	LUT2 #(
		.INIT('h8)
	) name7899 (
		_w11944_,
		_w11945_,
		_w11946_
	);
	LUT2 #(
		.INIT('h2)
	) name7900 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w11946_,
		_w11947_
	);
	LUT2 #(
		.INIT('h1)
	) name7901 (
		_w11898_,
		_w11904_,
		_w11948_
	);
	LUT2 #(
		.INIT('h8)
	) name7902 (
		_w11907_,
		_w11948_,
		_w11949_
	);
	LUT2 #(
		.INIT('h4)
	) name7903 (
		_w11843_,
		_w11949_,
		_w11950_
	);
	LUT2 #(
		.INIT('h1)
	) name7904 (
		_w11859_,
		_w11890_,
		_w11951_
	);
	LUT2 #(
		.INIT('h8)
	) name7905 (
		_w11950_,
		_w11951_,
		_w11952_
	);
	LUT2 #(
		.INIT('h4)
	) name7906 (
		_w11947_,
		_w11952_,
		_w11953_
	);
	LUT2 #(
		.INIT('h4)
	) name7907 (
		_w11818_,
		_w11953_,
		_w11954_
	);
	LUT2 #(
		.INIT('h2)
	) name7908 (
		_w11770_,
		_w11954_,
		_w11955_
	);
	LUT2 #(
		.INIT('h8)
	) name7909 (
		\sport0_rxctl_RX_reg[14]/P0001 ,
		_w11774_,
		_w11956_
	);
	LUT2 #(
		.INIT('h8)
	) name7910 (
		\sport1_rxctl_RX_reg[14]/P0001 ,
		_w11772_,
		_w11957_
	);
	LUT2 #(
		.INIT('h8)
	) name7911 (
		\bdma_BRdataBUF_reg[14]/P0001 ,
		_w6918_,
		_w11958_
	);
	LUT2 #(
		.INIT('h1)
	) name7912 (
		_w11956_,
		_w11957_,
		_w11959_
	);
	LUT2 #(
		.INIT('h4)
	) name7913 (
		_w11817_,
		_w11959_,
		_w11960_
	);
	LUT2 #(
		.INIT('h4)
	) name7914 (
		_w11958_,
		_w11960_,
		_w11961_
	);
	LUT2 #(
		.INIT('h4)
	) name7915 (
		_w11955_,
		_w11961_,
		_w11962_
	);
	LUT2 #(
		.INIT('h8)
	) name7916 (
		\idma_DTMP_H_reg[15]/P0001 ,
		_w11762_,
		_w11963_
	);
	LUT2 #(
		.INIT('h8)
	) name7917 (
		\regout_STD_C_reg[15]/P0001 ,
		_w6988_,
		_w11964_
	);
	LUT2 #(
		.INIT('h4)
	) name7918 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001 ,
		_w11965_
	);
	LUT2 #(
		.INIT('h8)
	) name7919 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001 ,
		_w11966_
	);
	LUT2 #(
		.INIT('h1)
	) name7920 (
		_w11965_,
		_w11966_,
		_w11967_
	);
	LUT2 #(
		.INIT('h2)
	) name7921 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w11967_,
		_w11968_
	);
	LUT2 #(
		.INIT('h4)
	) name7922 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001 ,
		_w11969_
	);
	LUT2 #(
		.INIT('h8)
	) name7923 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001 ,
		_w11970_
	);
	LUT2 #(
		.INIT('h1)
	) name7924 (
		_w11969_,
		_w11970_,
		_w11971_
	);
	LUT2 #(
		.INIT('h2)
	) name7925 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w11971_,
		_w11972_
	);
	LUT2 #(
		.INIT('h4)
	) name7926 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001 ,
		_w11973_
	);
	LUT2 #(
		.INIT('h8)
	) name7927 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001 ,
		_w11974_
	);
	LUT2 #(
		.INIT('h1)
	) name7928 (
		_w11973_,
		_w11974_,
		_w11975_
	);
	LUT2 #(
		.INIT('h2)
	) name7929 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w11975_,
		_w11976_
	);
	LUT2 #(
		.INIT('h4)
	) name7930 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001 ,
		_w11977_
	);
	LUT2 #(
		.INIT('h8)
	) name7931 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001 ,
		_w11978_
	);
	LUT2 #(
		.INIT('h1)
	) name7932 (
		_w11977_,
		_w11978_,
		_w11979_
	);
	LUT2 #(
		.INIT('h2)
	) name7933 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w11979_,
		_w11980_
	);
	LUT2 #(
		.INIT('h4)
	) name7934 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001 ,
		_w11981_
	);
	LUT2 #(
		.INIT('h8)
	) name7935 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001 ,
		_w11982_
	);
	LUT2 #(
		.INIT('h1)
	) name7936 (
		_w11981_,
		_w11982_,
		_w11983_
	);
	LUT2 #(
		.INIT('h2)
	) name7937 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w11983_,
		_w11984_
	);
	LUT2 #(
		.INIT('h1)
	) name7938 (
		_w11968_,
		_w11972_,
		_w11985_
	);
	LUT2 #(
		.INIT('h1)
	) name7939 (
		_w11976_,
		_w11980_,
		_w11986_
	);
	LUT2 #(
		.INIT('h4)
	) name7940 (
		_w11984_,
		_w11986_,
		_w11987_
	);
	LUT2 #(
		.INIT('h8)
	) name7941 (
		_w11985_,
		_w11987_,
		_w11988_
	);
	LUT2 #(
		.INIT('h2)
	) name7942 (
		_w7093_,
		_w11988_,
		_w11989_
	);
	LUT2 #(
		.INIT('h4)
	) name7943 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 ,
		_w11990_
	);
	LUT2 #(
		.INIT('h8)
	) name7944 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 ,
		_w11991_
	);
	LUT2 #(
		.INIT('h1)
	) name7945 (
		_w11990_,
		_w11991_,
		_w11992_
	);
	LUT2 #(
		.INIT('h2)
	) name7946 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w11992_,
		_w11993_
	);
	LUT2 #(
		.INIT('h4)
	) name7947 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001 ,
		_w11994_
	);
	LUT2 #(
		.INIT('h8)
	) name7948 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001 ,
		_w11995_
	);
	LUT2 #(
		.INIT('h1)
	) name7949 (
		_w11994_,
		_w11995_,
		_w11996_
	);
	LUT2 #(
		.INIT('h2)
	) name7950 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w11996_,
		_w11997_
	);
	LUT2 #(
		.INIT('h4)
	) name7951 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 ,
		_w11998_
	);
	LUT2 #(
		.INIT('h8)
	) name7952 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 ,
		_w11999_
	);
	LUT2 #(
		.INIT('h1)
	) name7953 (
		_w11998_,
		_w11999_,
		_w12000_
	);
	LUT2 #(
		.INIT('h2)
	) name7954 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w12000_,
		_w12001_
	);
	LUT2 #(
		.INIT('h1)
	) name7955 (
		_w11993_,
		_w11997_,
		_w12002_
	);
	LUT2 #(
		.INIT('h4)
	) name7956 (
		_w12001_,
		_w12002_,
		_w12003_
	);
	LUT2 #(
		.INIT('h8)
	) name7957 (
		_w7174_,
		_w12003_,
		_w12004_
	);
	LUT2 #(
		.INIT('h2)
	) name7958 (
		_w7153_,
		_w12004_,
		_w12005_
	);
	LUT2 #(
		.INIT('h4)
	) name7959 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001 ,
		_w12006_
	);
	LUT2 #(
		.INIT('h8)
	) name7960 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001 ,
		_w12007_
	);
	LUT2 #(
		.INIT('h1)
	) name7961 (
		_w12006_,
		_w12007_,
		_w12008_
	);
	LUT2 #(
		.INIT('h2)
	) name7962 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w12008_,
		_w12009_
	);
	LUT2 #(
		.INIT('h4)
	) name7963 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001 ,
		_w12010_
	);
	LUT2 #(
		.INIT('h8)
	) name7964 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001 ,
		_w12011_
	);
	LUT2 #(
		.INIT('h1)
	) name7965 (
		_w12010_,
		_w12011_,
		_w12012_
	);
	LUT2 #(
		.INIT('h2)
	) name7966 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w12012_,
		_w12013_
	);
	LUT2 #(
		.INIT('h4)
	) name7967 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001 ,
		_w12014_
	);
	LUT2 #(
		.INIT('h8)
	) name7968 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001 ,
		_w12015_
	);
	LUT2 #(
		.INIT('h1)
	) name7969 (
		_w12014_,
		_w12015_,
		_w12016_
	);
	LUT2 #(
		.INIT('h2)
	) name7970 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w12016_,
		_w12017_
	);
	LUT2 #(
		.INIT('h4)
	) name7971 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001 ,
		_w12018_
	);
	LUT2 #(
		.INIT('h8)
	) name7972 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001 ,
		_w12019_
	);
	LUT2 #(
		.INIT('h1)
	) name7973 (
		_w12018_,
		_w12019_,
		_w12020_
	);
	LUT2 #(
		.INIT('h2)
	) name7974 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w12020_,
		_w12021_
	);
	LUT2 #(
		.INIT('h4)
	) name7975 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001 ,
		_w12022_
	);
	LUT2 #(
		.INIT('h8)
	) name7976 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 ,
		_w12023_
	);
	LUT2 #(
		.INIT('h1)
	) name7977 (
		_w12022_,
		_w12023_,
		_w12024_
	);
	LUT2 #(
		.INIT('h2)
	) name7978 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w12024_,
		_w12025_
	);
	LUT2 #(
		.INIT('h4)
	) name7979 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 ,
		_w12026_
	);
	LUT2 #(
		.INIT('h8)
	) name7980 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 ,
		_w12027_
	);
	LUT2 #(
		.INIT('h1)
	) name7981 (
		_w12026_,
		_w12027_,
		_w12028_
	);
	LUT2 #(
		.INIT('h2)
	) name7982 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w12028_,
		_w12029_
	);
	LUT2 #(
		.INIT('h1)
	) name7983 (
		_w7207_,
		_w12009_,
		_w12030_
	);
	LUT2 #(
		.INIT('h1)
	) name7984 (
		_w12013_,
		_w12017_,
		_w12031_
	);
	LUT2 #(
		.INIT('h1)
	) name7985 (
		_w12021_,
		_w12025_,
		_w12032_
	);
	LUT2 #(
		.INIT('h4)
	) name7986 (
		_w12029_,
		_w12032_,
		_w12033_
	);
	LUT2 #(
		.INIT('h8)
	) name7987 (
		_w12030_,
		_w12031_,
		_w12034_
	);
	LUT2 #(
		.INIT('h8)
	) name7988 (
		_w12033_,
		_w12034_,
		_w12035_
	);
	LUT2 #(
		.INIT('h2)
	) name7989 (
		_w7179_,
		_w12035_,
		_w12036_
	);
	LUT2 #(
		.INIT('h8)
	) name7990 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		\sport1_txctl_TX_reg[15]/P0001 ,
		_w12037_
	);
	LUT2 #(
		.INIT('h8)
	) name7991 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		\sport1_rxctl_RX_reg[15]/P0001 ,
		_w12038_
	);
	LUT2 #(
		.INIT('h8)
	) name7992 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w12039_
	);
	LUT2 #(
		.INIT('h8)
	) name7993 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		\sport0_rxctl_RX_reg[15]/P0001 ,
		_w12040_
	);
	LUT2 #(
		.INIT('h1)
	) name7994 (
		_w12037_,
		_w12038_,
		_w12041_
	);
	LUT2 #(
		.INIT('h1)
	) name7995 (
		_w12039_,
		_w12040_,
		_w12042_
	);
	LUT2 #(
		.INIT('h8)
	) name7996 (
		_w12041_,
		_w12042_,
		_w12043_
	);
	LUT2 #(
		.INIT('h2)
	) name7997 (
		_w7119_,
		_w12043_,
		_w12044_
	);
	LUT2 #(
		.INIT('h8)
	) name7998 (
		\core_c_dec_IRE_reg[19]/NET0131 ,
		\core_c_dec_imm16_E_reg/P0001 ,
		_w12045_
	);
	LUT2 #(
		.INIT('h8)
	) name7999 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w12046_
	);
	LUT2 #(
		.INIT('h1)
	) name8000 (
		_w11899_,
		_w12045_,
		_w12047_
	);
	LUT2 #(
		.INIT('h4)
	) name8001 (
		_w12046_,
		_w12047_,
		_w12048_
	);
	LUT2 #(
		.INIT('h2)
	) name8002 (
		_w7215_,
		_w12048_,
		_w12049_
	);
	LUT2 #(
		.INIT('h8)
	) name8003 (
		\tm_tsr_reg_DO_reg[8]/NET0131 ,
		_w7540_,
		_w12050_
	);
	LUT2 #(
		.INIT('h8)
	) name8004 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w7263_,
		_w12051_
	);
	LUT2 #(
		.INIT('h8)
	) name8005 (
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w7281_,
		_w12052_
	);
	LUT2 #(
		.INIT('h8)
	) name8006 (
		\bdma_BCTL_reg[15]/NET0131 ,
		_w7230_,
		_w12053_
	);
	LUT2 #(
		.INIT('h8)
	) name8007 (
		\PIO_oe[11]_pad ,
		_w7244_,
		_w12054_
	);
	LUT2 #(
		.INIT('h8)
	) name8008 (
		\tm_tpr_reg_DO_reg[15]/NET0131 ,
		_w7293_,
		_w12055_
	);
	LUT2 #(
		.INIT('h8)
	) name8009 (
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w7295_,
		_w12056_
	);
	LUT2 #(
		.INIT('h8)
	) name8010 (
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w7259_,
		_w12057_
	);
	LUT2 #(
		.INIT('h8)
	) name8011 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w7276_,
		_w12058_
	);
	LUT2 #(
		.INIT('h8)
	) name8012 (
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w7249_,
		_w12059_
	);
	LUT2 #(
		.INIT('h8)
	) name8013 (
		\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w7247_,
		_w12060_
	);
	LUT2 #(
		.INIT('h8)
	) name8014 (
		\pio_PINT_reg[11]/NET0131 ,
		_w7271_,
		_w12061_
	);
	LUT2 #(
		.INIT('h8)
	) name8015 (
		\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w7256_,
		_w12062_
	);
	LUT2 #(
		.INIT('h8)
	) name8016 (
		\pio_pmask_reg_DO_reg[11]/NET0131 ,
		_w7297_,
		_w12063_
	);
	LUT2 #(
		.INIT('h8)
	) name8017 (
		\sice_ICYC_en_reg/NET0131 ,
		_w7522_,
		_w12064_
	);
	LUT2 #(
		.INIT('h8)
	) name8018 (
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w7273_,
		_w12065_
	);
	LUT2 #(
		.INIT('h8)
	) name8019 (
		\memc_usysr_DO_reg[15]/NET0131 ,
		_w7301_,
		_w12066_
	);
	LUT2 #(
		.INIT('h8)
	) name8020 (
		\tm_TCR_TMP_reg[15]/NET0131 ,
		_w7289_,
		_w12067_
	);
	LUT2 #(
		.INIT('h8)
	) name8021 (
		\clkc_ckr_reg_DO_reg[15]/NET0131 ,
		_w7239_,
		_w12068_
	);
	LUT2 #(
		.INIT('h8)
	) name8022 (
		\PIO_out[11]_pad ,
		_w7291_,
		_w12069_
	);
	LUT2 #(
		.INIT('h1)
	) name8023 (
		_w12050_,
		_w12051_,
		_w12070_
	);
	LUT2 #(
		.INIT('h1)
	) name8024 (
		_w12052_,
		_w12054_,
		_w12071_
	);
	LUT2 #(
		.INIT('h1)
	) name8025 (
		_w12055_,
		_w12056_,
		_w12072_
	);
	LUT2 #(
		.INIT('h1)
	) name8026 (
		_w12057_,
		_w12058_,
		_w12073_
	);
	LUT2 #(
		.INIT('h1)
	) name8027 (
		_w12059_,
		_w12060_,
		_w12074_
	);
	LUT2 #(
		.INIT('h1)
	) name8028 (
		_w12061_,
		_w12062_,
		_w12075_
	);
	LUT2 #(
		.INIT('h1)
	) name8029 (
		_w12063_,
		_w12064_,
		_w12076_
	);
	LUT2 #(
		.INIT('h1)
	) name8030 (
		_w12065_,
		_w12066_,
		_w12077_
	);
	LUT2 #(
		.INIT('h1)
	) name8031 (
		_w12067_,
		_w12068_,
		_w12078_
	);
	LUT2 #(
		.INIT('h4)
	) name8032 (
		_w12069_,
		_w12078_,
		_w12079_
	);
	LUT2 #(
		.INIT('h8)
	) name8033 (
		_w12076_,
		_w12077_,
		_w12080_
	);
	LUT2 #(
		.INIT('h8)
	) name8034 (
		_w12074_,
		_w12075_,
		_w12081_
	);
	LUT2 #(
		.INIT('h8)
	) name8035 (
		_w12072_,
		_w12073_,
		_w12082_
	);
	LUT2 #(
		.INIT('h8)
	) name8036 (
		_w12070_,
		_w12071_,
		_w12083_
	);
	LUT2 #(
		.INIT('h8)
	) name8037 (
		_w12082_,
		_w12083_,
		_w12084_
	);
	LUT2 #(
		.INIT('h8)
	) name8038 (
		_w12080_,
		_w12081_,
		_w12085_
	);
	LUT2 #(
		.INIT('h8)
	) name8039 (
		_w12079_,
		_w12085_,
		_w12086_
	);
	LUT2 #(
		.INIT('h4)
	) name8040 (
		_w12053_,
		_w12084_,
		_w12087_
	);
	LUT2 #(
		.INIT('h8)
	) name8041 (
		_w12086_,
		_w12087_,
		_w12088_
	);
	LUT2 #(
		.INIT('h2)
	) name8042 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w12088_,
		_w12089_
	);
	LUT2 #(
		.INIT('h1)
	) name8043 (
		_w12044_,
		_w12049_,
		_w12090_
	);
	LUT2 #(
		.INIT('h8)
	) name8044 (
		_w11907_,
		_w12090_,
		_w12091_
	);
	LUT2 #(
		.INIT('h4)
	) name8045 (
		_w11989_,
		_w12091_,
		_w12092_
	);
	LUT2 #(
		.INIT('h1)
	) name8046 (
		_w12005_,
		_w12036_,
		_w12093_
	);
	LUT2 #(
		.INIT('h8)
	) name8047 (
		_w12092_,
		_w12093_,
		_w12094_
	);
	LUT2 #(
		.INIT('h4)
	) name8048 (
		_w12089_,
		_w12094_,
		_w12095_
	);
	LUT2 #(
		.INIT('h4)
	) name8049 (
		_w11964_,
		_w12095_,
		_w12096_
	);
	LUT2 #(
		.INIT('h2)
	) name8050 (
		_w11770_,
		_w12096_,
		_w12097_
	);
	LUT2 #(
		.INIT('h8)
	) name8051 (
		\sport0_rxctl_RX_reg[15]/P0001 ,
		_w11774_,
		_w12098_
	);
	LUT2 #(
		.INIT('h8)
	) name8052 (
		\sport1_rxctl_RX_reg[15]/P0001 ,
		_w11772_,
		_w12099_
	);
	LUT2 #(
		.INIT('h8)
	) name8053 (
		\bdma_BRdataBUF_reg[15]/P0001 ,
		_w6918_,
		_w12100_
	);
	LUT2 #(
		.INIT('h1)
	) name8054 (
		_w12098_,
		_w12099_,
		_w12101_
	);
	LUT2 #(
		.INIT('h4)
	) name8055 (
		_w11963_,
		_w12101_,
		_w12102_
	);
	LUT2 #(
		.INIT('h4)
	) name8056 (
		_w12100_,
		_w12102_,
		_w12103_
	);
	LUT2 #(
		.INIT('h4)
	) name8057 (
		_w12097_,
		_w12103_,
		_w12104_
	);
	LUT2 #(
		.INIT('h8)
	) name8058 (
		\idma_DTMP_H_reg[1]/P0001 ,
		_w11762_,
		_w12105_
	);
	LUT2 #(
		.INIT('h4)
	) name8059 (
		_w9430_,
		_w11770_,
		_w12106_
	);
	LUT2 #(
		.INIT('h8)
	) name8060 (
		\sport1_rxctl_RX_reg[1]/P0001 ,
		_w11772_,
		_w12107_
	);
	LUT2 #(
		.INIT('h8)
	) name8061 (
		\sport0_rxctl_RX_reg[1]/P0001 ,
		_w11774_,
		_w12108_
	);
	LUT2 #(
		.INIT('h8)
	) name8062 (
		\bdma_BRdataBUF_reg[1]/P0001 ,
		_w6918_,
		_w12109_
	);
	LUT2 #(
		.INIT('h1)
	) name8063 (
		_w12107_,
		_w12108_,
		_w12110_
	);
	LUT2 #(
		.INIT('h4)
	) name8064 (
		_w12105_,
		_w12110_,
		_w12111_
	);
	LUT2 #(
		.INIT('h4)
	) name8065 (
		_w12109_,
		_w12111_,
		_w12112_
	);
	LUT2 #(
		.INIT('h4)
	) name8066 (
		_w12106_,
		_w12112_,
		_w12113_
	);
	LUT2 #(
		.INIT('h8)
	) name8067 (
		\idma_DTMP_H_reg[2]/P0001 ,
		_w11762_,
		_w12114_
	);
	LUT2 #(
		.INIT('h4)
	) name8068 (
		_w8710_,
		_w11770_,
		_w12115_
	);
	LUT2 #(
		.INIT('h8)
	) name8069 (
		\sport1_rxctl_RX_reg[2]/P0001 ,
		_w11772_,
		_w12116_
	);
	LUT2 #(
		.INIT('h8)
	) name8070 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w11774_,
		_w12117_
	);
	LUT2 #(
		.INIT('h8)
	) name8071 (
		\bdma_BRdataBUF_reg[2]/P0001 ,
		_w6918_,
		_w12118_
	);
	LUT2 #(
		.INIT('h1)
	) name8072 (
		_w12116_,
		_w12117_,
		_w12119_
	);
	LUT2 #(
		.INIT('h4)
	) name8073 (
		_w12114_,
		_w12119_,
		_w12120_
	);
	LUT2 #(
		.INIT('h4)
	) name8074 (
		_w12118_,
		_w12120_,
		_w12121_
	);
	LUT2 #(
		.INIT('h4)
	) name8075 (
		_w12115_,
		_w12121_,
		_w12122_
	);
	LUT2 #(
		.INIT('h8)
	) name8076 (
		\idma_DTMP_H_reg[3]/P0001 ,
		_w11762_,
		_w12123_
	);
	LUT2 #(
		.INIT('h4)
	) name8077 (
		_w8108_,
		_w11770_,
		_w12124_
	);
	LUT2 #(
		.INIT('h8)
	) name8078 (
		\sport1_rxctl_RX_reg[3]/P0001 ,
		_w11772_,
		_w12125_
	);
	LUT2 #(
		.INIT('h8)
	) name8079 (
		\sport0_rxctl_RX_reg[3]/P0001 ,
		_w11774_,
		_w12126_
	);
	LUT2 #(
		.INIT('h8)
	) name8080 (
		\bdma_BRdataBUF_reg[3]/P0001 ,
		_w6918_,
		_w12127_
	);
	LUT2 #(
		.INIT('h1)
	) name8081 (
		_w12125_,
		_w12126_,
		_w12128_
	);
	LUT2 #(
		.INIT('h4)
	) name8082 (
		_w12123_,
		_w12128_,
		_w12129_
	);
	LUT2 #(
		.INIT('h4)
	) name8083 (
		_w12127_,
		_w12129_,
		_w12130_
	);
	LUT2 #(
		.INIT('h4)
	) name8084 (
		_w12124_,
		_w12130_,
		_w12131_
	);
	LUT2 #(
		.INIT('h8)
	) name8085 (
		\idma_DTMP_H_reg[4]/P0001 ,
		_w11762_,
		_w12132_
	);
	LUT2 #(
		.INIT('h4)
	) name8086 (
		_w10064_,
		_w11770_,
		_w12133_
	);
	LUT2 #(
		.INIT('h8)
	) name8087 (
		\sport1_rxctl_RX_reg[4]/P0001 ,
		_w11772_,
		_w12134_
	);
	LUT2 #(
		.INIT('h8)
	) name8088 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w11774_,
		_w12135_
	);
	LUT2 #(
		.INIT('h8)
	) name8089 (
		\bdma_BRdataBUF_reg[4]/P0001 ,
		_w6918_,
		_w12136_
	);
	LUT2 #(
		.INIT('h1)
	) name8090 (
		_w12134_,
		_w12135_,
		_w12137_
	);
	LUT2 #(
		.INIT('h4)
	) name8091 (
		_w12132_,
		_w12137_,
		_w12138_
	);
	LUT2 #(
		.INIT('h4)
	) name8092 (
		_w12136_,
		_w12138_,
		_w12139_
	);
	LUT2 #(
		.INIT('h4)
	) name8093 (
		_w12133_,
		_w12139_,
		_w12140_
	);
	LUT2 #(
		.INIT('h8)
	) name8094 (
		\idma_DTMP_H_reg[5]/P0001 ,
		_w11762_,
		_w12141_
	);
	LUT2 #(
		.INIT('h4)
	) name8095 (
		_w10906_,
		_w11770_,
		_w12142_
	);
	LUT2 #(
		.INIT('h8)
	) name8096 (
		\sport1_rxctl_RX_reg[5]/P0001 ,
		_w11772_,
		_w12143_
	);
	LUT2 #(
		.INIT('h8)
	) name8097 (
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w11774_,
		_w12144_
	);
	LUT2 #(
		.INIT('h8)
	) name8098 (
		\bdma_BRdataBUF_reg[5]/P0001 ,
		_w6918_,
		_w12145_
	);
	LUT2 #(
		.INIT('h1)
	) name8099 (
		_w12143_,
		_w12144_,
		_w12146_
	);
	LUT2 #(
		.INIT('h4)
	) name8100 (
		_w12141_,
		_w12146_,
		_w12147_
	);
	LUT2 #(
		.INIT('h4)
	) name8101 (
		_w12145_,
		_w12147_,
		_w12148_
	);
	LUT2 #(
		.INIT('h4)
	) name8102 (
		_w12142_,
		_w12148_,
		_w12149_
	);
	LUT2 #(
		.INIT('h8)
	) name8103 (
		\idma_DTMP_H_reg[6]/P0001 ,
		_w11762_,
		_w12150_
	);
	LUT2 #(
		.INIT('h4)
	) name8104 (
		_w11520_,
		_w11770_,
		_w12151_
	);
	LUT2 #(
		.INIT('h8)
	) name8105 (
		\sport1_rxctl_RX_reg[6]/P0001 ,
		_w11772_,
		_w12152_
	);
	LUT2 #(
		.INIT('h8)
	) name8106 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w11774_,
		_w12153_
	);
	LUT2 #(
		.INIT('h8)
	) name8107 (
		\bdma_BRdataBUF_reg[6]/P0001 ,
		_w6918_,
		_w12154_
	);
	LUT2 #(
		.INIT('h1)
	) name8108 (
		_w12152_,
		_w12153_,
		_w12155_
	);
	LUT2 #(
		.INIT('h4)
	) name8109 (
		_w12150_,
		_w12155_,
		_w12156_
	);
	LUT2 #(
		.INIT('h4)
	) name8110 (
		_w12154_,
		_w12156_,
		_w12157_
	);
	LUT2 #(
		.INIT('h4)
	) name8111 (
		_w12151_,
		_w12157_,
		_w12158_
	);
	LUT2 #(
		.INIT('h8)
	) name8112 (
		\bdma_BRdataBUF_reg[7]/P0001 ,
		_w6918_,
		_w12159_
	);
	LUT2 #(
		.INIT('h8)
	) name8113 (
		\sport1_rxctl_RX_reg[7]/P0001 ,
		_w11772_,
		_w12160_
	);
	LUT2 #(
		.INIT('h8)
	) name8114 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w11774_,
		_w12161_
	);
	LUT2 #(
		.INIT('h8)
	) name8115 (
		\idma_DTMP_H_reg[7]/P0001 ,
		_w11762_,
		_w12162_
	);
	LUT2 #(
		.INIT('h4)
	) name8116 (
		_w11260_,
		_w11770_,
		_w12163_
	);
	LUT2 #(
		.INIT('h1)
	) name8117 (
		_w12160_,
		_w12161_,
		_w12164_
	);
	LUT2 #(
		.INIT('h4)
	) name8118 (
		_w12159_,
		_w12164_,
		_w12165_
	);
	LUT2 #(
		.INIT('h4)
	) name8119 (
		_w12162_,
		_w12165_,
		_w12166_
	);
	LUT2 #(
		.INIT('h4)
	) name8120 (
		_w12163_,
		_w12166_,
		_w12167_
	);
	LUT2 #(
		.INIT('h8)
	) name8121 (
		\idma_DTMP_H_reg[8]/P0001 ,
		_w11762_,
		_w12168_
	);
	LUT2 #(
		.INIT('h4)
	) name8122 (
		_w10633_,
		_w11770_,
		_w12169_
	);
	LUT2 #(
		.INIT('h8)
	) name8123 (
		\sport1_rxctl_RX_reg[8]/P0001 ,
		_w11772_,
		_w12170_
	);
	LUT2 #(
		.INIT('h8)
	) name8124 (
		\sport0_rxctl_RX_reg[8]/P0001 ,
		_w11774_,
		_w12171_
	);
	LUT2 #(
		.INIT('h8)
	) name8125 (
		\bdma_BRdataBUF_reg[8]/P0001 ,
		_w6918_,
		_w12172_
	);
	LUT2 #(
		.INIT('h1)
	) name8126 (
		_w12170_,
		_w12171_,
		_w12173_
	);
	LUT2 #(
		.INIT('h4)
	) name8127 (
		_w12168_,
		_w12173_,
		_w12174_
	);
	LUT2 #(
		.INIT('h4)
	) name8128 (
		_w12172_,
		_w12174_,
		_w12175_
	);
	LUT2 #(
		.INIT('h4)
	) name8129 (
		_w12169_,
		_w12175_,
		_w12176_
	);
	LUT2 #(
		.INIT('h8)
	) name8130 (
		\idma_DTMP_H_reg[9]/P0001 ,
		_w11762_,
		_w12177_
	);
	LUT2 #(
		.INIT('h4)
	) name8131 (
		_w10284_,
		_w11770_,
		_w12178_
	);
	LUT2 #(
		.INIT('h8)
	) name8132 (
		\sport0_rxctl_RX_reg[9]/P0001 ,
		_w11774_,
		_w12179_
	);
	LUT2 #(
		.INIT('h8)
	) name8133 (
		\sport1_rxctl_RX_reg[9]/P0001 ,
		_w11772_,
		_w12180_
	);
	LUT2 #(
		.INIT('h8)
	) name8134 (
		\bdma_BRdataBUF_reg[9]/P0001 ,
		_w6918_,
		_w12181_
	);
	LUT2 #(
		.INIT('h1)
	) name8135 (
		_w12179_,
		_w12180_,
		_w12182_
	);
	LUT2 #(
		.INIT('h4)
	) name8136 (
		_w12177_,
		_w12182_,
		_w12183_
	);
	LUT2 #(
		.INIT('h4)
	) name8137 (
		_w12181_,
		_w12183_,
		_w12184_
	);
	LUT2 #(
		.INIT('h4)
	) name8138 (
		_w12178_,
		_w12184_,
		_w12185_
	);
	LUT2 #(
		.INIT('h2)
	) name8139 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		_w5066_,
		_w12186_
	);
	LUT2 #(
		.INIT('h8)
	) name8140 (
		\bdma_BOVL_reg[6]/NET0131 ,
		_w5066_,
		_w12187_
	);
	LUT2 #(
		.INIT('h1)
	) name8141 (
		_w12186_,
		_w12187_,
		_w12188_
	);
	LUT2 #(
		.INIT('h1)
	) name8142 (
		_w5895_,
		_w12188_,
		_w12189_
	);
	LUT2 #(
		.INIT('h8)
	) name8143 (
		\idma_DOVL_reg[6]/NET0131 ,
		_w5895_,
		_w12190_
	);
	LUT2 #(
		.INIT('h1)
	) name8144 (
		_w12189_,
		_w12190_,
		_w12191_
	);
	LUT2 #(
		.INIT('h2)
	) name8145 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		_w5066_,
		_w12192_
	);
	LUT2 #(
		.INIT('h8)
	) name8146 (
		\bdma_BOVL_reg[7]/NET0131 ,
		_w5066_,
		_w12193_
	);
	LUT2 #(
		.INIT('h1)
	) name8147 (
		_w12192_,
		_w12193_,
		_w12194_
	);
	LUT2 #(
		.INIT('h1)
	) name8148 (
		_w5895_,
		_w12194_,
		_w12195_
	);
	LUT2 #(
		.INIT('h8)
	) name8149 (
		\idma_DOVL_reg[7]/NET0131 ,
		_w5895_,
		_w12196_
	);
	LUT2 #(
		.INIT('h1)
	) name8150 (
		_w12195_,
		_w12196_,
		_w12197_
	);
	LUT2 #(
		.INIT('h8)
	) name8151 (
		_w12191_,
		_w12197_,
		_w12198_
	);
	LUT2 #(
		.INIT('h2)
	) name8152 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		_w5066_,
		_w12199_
	);
	LUT2 #(
		.INIT('h8)
	) name8153 (
		\bdma_BOVL_reg[4]/NET0131 ,
		_w5066_,
		_w12200_
	);
	LUT2 #(
		.INIT('h1)
	) name8154 (
		_w12199_,
		_w12200_,
		_w12201_
	);
	LUT2 #(
		.INIT('h1)
	) name8155 (
		_w5895_,
		_w12201_,
		_w12202_
	);
	LUT2 #(
		.INIT('h8)
	) name8156 (
		\idma_DOVL_reg[4]/NET0131 ,
		_w5895_,
		_w12203_
	);
	LUT2 #(
		.INIT('h1)
	) name8157 (
		_w12202_,
		_w12203_,
		_w12204_
	);
	LUT2 #(
		.INIT('h8)
	) name8158 (
		_w12198_,
		_w12204_,
		_w12205_
	);
	LUT2 #(
		.INIT('h2)
	) name8159 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		_w5066_,
		_w12206_
	);
	LUT2 #(
		.INIT('h8)
	) name8160 (
		\bdma_BOVL_reg[5]/NET0131 ,
		_w5066_,
		_w12207_
	);
	LUT2 #(
		.INIT('h1)
	) name8161 (
		_w12206_,
		_w12207_,
		_w12208_
	);
	LUT2 #(
		.INIT('h1)
	) name8162 (
		_w5895_,
		_w12208_,
		_w12209_
	);
	LUT2 #(
		.INIT('h8)
	) name8163 (
		\idma_DOVL_reg[5]/NET0131 ,
		_w5895_,
		_w12210_
	);
	LUT2 #(
		.INIT('h1)
	) name8164 (
		_w12209_,
		_w12210_,
		_w12211_
	);
	LUT2 #(
		.INIT('h8)
	) name8165 (
		_w9513_,
		_w12211_,
		_w12212_
	);
	LUT2 #(
		.INIT('h8)
	) name8166 (
		_w12205_,
		_w12212_,
		_w12213_
	);
	LUT2 #(
		.INIT('h4)
	) name8167 (
		_w11766_,
		_w12213_,
		_w12214_
	);
	LUT2 #(
		.INIT('h2)
	) name8168 (
		_w12198_,
		_w12204_,
		_w12215_
	);
	LUT2 #(
		.INIT('h8)
	) name8169 (
		_w12212_,
		_w12215_,
		_w12216_
	);
	LUT2 #(
		.INIT('h4)
	) name8170 (
		_w11766_,
		_w12216_,
		_w12217_
	);
	LUT2 #(
		.INIT('h2)
	) name8171 (
		_w9513_,
		_w12211_,
		_w12218_
	);
	LUT2 #(
		.INIT('h8)
	) name8172 (
		_w12205_,
		_w12218_,
		_w12219_
	);
	LUT2 #(
		.INIT('h4)
	) name8173 (
		_w11766_,
		_w12219_,
		_w12220_
	);
	LUT2 #(
		.INIT('h8)
	) name8174 (
		_w12215_,
		_w12218_,
		_w12221_
	);
	LUT2 #(
		.INIT('h4)
	) name8175 (
		_w11766_,
		_w12221_,
		_w12222_
	);
	LUT2 #(
		.INIT('h4)
	) name8176 (
		_w12191_,
		_w12197_,
		_w12223_
	);
	LUT2 #(
		.INIT('h8)
	) name8177 (
		_w12204_,
		_w12223_,
		_w12224_
	);
	LUT2 #(
		.INIT('h8)
	) name8178 (
		_w12212_,
		_w12224_,
		_w12225_
	);
	LUT2 #(
		.INIT('h4)
	) name8179 (
		_w11766_,
		_w12225_,
		_w12226_
	);
	LUT2 #(
		.INIT('h4)
	) name8180 (
		_w12204_,
		_w12223_,
		_w12227_
	);
	LUT2 #(
		.INIT('h8)
	) name8181 (
		_w12212_,
		_w12227_,
		_w12228_
	);
	LUT2 #(
		.INIT('h4)
	) name8182 (
		_w11766_,
		_w12228_,
		_w12229_
	);
	LUT2 #(
		.INIT('h8)
	) name8183 (
		_w12218_,
		_w12224_,
		_w12230_
	);
	LUT2 #(
		.INIT('h4)
	) name8184 (
		_w11766_,
		_w12230_,
		_w12231_
	);
	LUT2 #(
		.INIT('h8)
	) name8185 (
		_w12218_,
		_w12227_,
		_w12232_
	);
	LUT2 #(
		.INIT('h4)
	) name8186 (
		_w11766_,
		_w12232_,
		_w12233_
	);
	LUT2 #(
		.INIT('h8)
	) name8187 (
		T_ICE_RSTn_pad,
		T_RSTn_pad,
		_w12234_
	);
	LUT2 #(
		.INIT('h8)
	) name8188 (
		\clkc_DSPoff_reg/NET0131 ,
		_w12234_,
		_w12235_
	);
	LUT2 #(
		.INIT('h8)
	) name8189 (
		\clkc_SlowDn_reg/NET0131 ,
		_w12234_,
		_w12236_
	);
	LUT2 #(
		.INIT('h4)
	) name8190 (
		T_CLKI_PLL_pad,
		T_Sel_PLL_pad,
		_w12237_
	);
	LUT2 #(
		.INIT('h1)
	) name8191 (
		T_CLKI_OSC_pad,
		T_Sel_PLL_pad,
		_w12238_
	);
	LUT2 #(
		.INIT('h8)
	) name8192 (
		\clkc_OSCoff_reg/NET0131 ,
		_w12234_,
		_w12239_
	);
	LUT2 #(
		.INIT('h1)
	) name8193 (
		_w12237_,
		_w12238_,
		_w12240_
	);
	LUT2 #(
		.INIT('h4)
	) name8194 (
		_w12239_,
		_w12240_,
		_w12241_
	);
	LUT2 #(
		.INIT('h4)
	) name8195 (
		_w12236_,
		_w12241_,
		_w12242_
	);
	LUT2 #(
		.INIT('h8)
	) name8196 (
		\clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131 ,
		_w12236_,
		_w12243_
	);
	LUT2 #(
		.INIT('h1)
	) name8197 (
		_w12242_,
		_w12243_,
		_w12244_
	);
	LUT2 #(
		.INIT('h4)
	) name8198 (
		_w12235_,
		_w12244_,
		_w12245_
	);
	LUT2 #(
		.INIT('h8)
	) name8199 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		_w5602_,
		_w12246_
	);
	LUT2 #(
		.INIT('h8)
	) name8200 (
		\emc_ECS_reg[3]/NET0131 ,
		_w5592_,
		_w12247_
	);
	LUT2 #(
		.INIT('h8)
	) name8201 (
		\emc_ECMcs_reg/NET0131 ,
		_w12247_,
		_w12248_
	);
	LUT2 #(
		.INIT('h8)
	) name8202 (
		\sice_idr1_reg_DO_reg[4]/P0001 ,
		_w12248_,
		_w12249_
	);
	LUT2 #(
		.INIT('h2)
	) name8203 (
		\emc_ECMcs_reg/NET0131 ,
		_w12247_,
		_w12250_
	);
	LUT2 #(
		.INIT('h8)
	) name8204 (
		\emc_ECMA_reg[0]/P0001 ,
		_w12250_,
		_w12251_
	);
	LUT2 #(
		.INIT('h2)
	) name8205 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		_w5608_,
		_w12252_
	);
	LUT2 #(
		.INIT('h8)
	) name8206 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w5610_,
		_w12253_
	);
	LUT2 #(
		.INIT('h1)
	) name8207 (
		_w12249_,
		_w12251_,
		_w12254_
	);
	LUT2 #(
		.INIT('h4)
	) name8208 (
		_w12246_,
		_w12254_,
		_w12255_
	);
	LUT2 #(
		.INIT('h1)
	) name8209 (
		_w12252_,
		_w12253_,
		_w12256_
	);
	LUT2 #(
		.INIT('h8)
	) name8210 (
		_w12255_,
		_w12256_,
		_w12257_
	);
	LUT2 #(
		.INIT('h1)
	) name8211 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12257_,
		_w12258_
	);
	LUT2 #(
		.INIT('h8)
	) name8212 (
		\bdma_BEAD_reg[0]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12259_
	);
	LUT2 #(
		.INIT('h1)
	) name8213 (
		_w12258_,
		_w12259_,
		_w12260_
	);
	LUT2 #(
		.INIT('h8)
	) name8214 (
		\bdma_BEAD_reg[10]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12261_
	);
	LUT2 #(
		.INIT('h8)
	) name8215 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w5602_,
		_w12262_
	);
	LUT2 #(
		.INIT('h2)
	) name8216 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w5608_,
		_w12263_
	);
	LUT2 #(
		.INIT('h8)
	) name8217 (
		\emc_ECMA_reg[10]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w12264_
	);
	LUT2 #(
		.INIT('h8)
	) name8218 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w5610_,
		_w12265_
	);
	LUT2 #(
		.INIT('h1)
	) name8219 (
		_w12262_,
		_w12264_,
		_w12266_
	);
	LUT2 #(
		.INIT('h1)
	) name8220 (
		_w12263_,
		_w12265_,
		_w12267_
	);
	LUT2 #(
		.INIT('h8)
	) name8221 (
		_w12266_,
		_w12267_,
		_w12268_
	);
	LUT2 #(
		.INIT('h1)
	) name8222 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12268_,
		_w12269_
	);
	LUT2 #(
		.INIT('h1)
	) name8223 (
		_w12261_,
		_w12269_,
		_w12270_
	);
	LUT2 #(
		.INIT('h8)
	) name8224 (
		\bdma_BEAD_reg[12]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12271_
	);
	LUT2 #(
		.INIT('h8)
	) name8225 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		_w5602_,
		_w12272_
	);
	LUT2 #(
		.INIT('h1)
	) name8226 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w5673_,
		_w12273_
	);
	LUT2 #(
		.INIT('h8)
	) name8227 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w12274_
	);
	LUT2 #(
		.INIT('h2)
	) name8228 (
		_w5642_,
		_w12274_,
		_w12275_
	);
	LUT2 #(
		.INIT('h8)
	) name8229 (
		_w12273_,
		_w12275_,
		_w12276_
	);
	LUT2 #(
		.INIT('h1)
	) name8230 (
		\emc_ECMA_reg[12]/P0001 ,
		_w12276_,
		_w12277_
	);
	LUT2 #(
		.INIT('h4)
	) name8231 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w12276_,
		_w12278_
	);
	LUT2 #(
		.INIT('h1)
	) name8232 (
		PM_bdry_sel_pad,
		_w12277_,
		_w12279_
	);
	LUT2 #(
		.INIT('h4)
	) name8233 (
		_w12278_,
		_w12279_,
		_w12280_
	);
	LUT2 #(
		.INIT('h4)
	) name8234 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w5673_,
		_w12281_
	);
	LUT2 #(
		.INIT('h1)
	) name8235 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w12282_
	);
	LUT2 #(
		.INIT('h4)
	) name8236 (
		\emc_ECMA_reg[12]/P0001 ,
		_w12282_,
		_w12283_
	);
	LUT2 #(
		.INIT('h4)
	) name8237 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w5643_,
		_w12284_
	);
	LUT2 #(
		.INIT('h2)
	) name8238 (
		_w12281_,
		_w12283_,
		_w12285_
	);
	LUT2 #(
		.INIT('h8)
	) name8239 (
		_w12284_,
		_w12285_,
		_w12286_
	);
	LUT2 #(
		.INIT('h1)
	) name8240 (
		_w12280_,
		_w12286_,
		_w12287_
	);
	LUT2 #(
		.INIT('h2)
	) name8241 (
		\emc_ECMcs_reg/NET0131 ,
		_w12287_,
		_w12288_
	);
	LUT2 #(
		.INIT('h1)
	) name8242 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		_w12289_
	);
	LUT2 #(
		.INIT('h2)
	) name8243 (
		PM_bdry_sel_pad,
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w12290_
	);
	LUT2 #(
		.INIT('h1)
	) name8244 (
		_w12289_,
		_w12290_,
		_w12291_
	);
	LUT2 #(
		.INIT('h4)
	) name8245 (
		_w5608_,
		_w12291_,
		_w12292_
	);
	LUT2 #(
		.INIT('h1)
	) name8246 (
		_w12272_,
		_w12292_,
		_w12293_
	);
	LUT2 #(
		.INIT('h4)
	) name8247 (
		_w12288_,
		_w12293_,
		_w12294_
	);
	LUT2 #(
		.INIT('h1)
	) name8248 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12294_,
		_w12295_
	);
	LUT2 #(
		.INIT('h1)
	) name8249 (
		_w12271_,
		_w12295_,
		_w12296_
	);
	LUT2 #(
		.INIT('h8)
	) name8250 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		_w5602_,
		_w12297_
	);
	LUT2 #(
		.INIT('h8)
	) name8251 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w5673_,
		_w12298_
	);
	LUT2 #(
		.INIT('h4)
	) name8252 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w12298_,
		_w12299_
	);
	LUT2 #(
		.INIT('h8)
	) name8253 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w12281_,
		_w12300_
	);
	LUT2 #(
		.INIT('h1)
	) name8254 (
		_w12299_,
		_w12300_,
		_w12301_
	);
	LUT2 #(
		.INIT('h2)
	) name8255 (
		_w12284_,
		_w12301_,
		_w12302_
	);
	LUT2 #(
		.INIT('h4)
	) name8256 (
		PM_bdry_sel_pad,
		_w12273_,
		_w12303_
	);
	LUT2 #(
		.INIT('h4)
	) name8257 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w5642_,
		_w12304_
	);
	LUT2 #(
		.INIT('h8)
	) name8258 (
		_w12303_,
		_w12304_,
		_w12305_
	);
	LUT2 #(
		.INIT('h1)
	) name8259 (
		_w12302_,
		_w12305_,
		_w12306_
	);
	LUT2 #(
		.INIT('h2)
	) name8260 (
		\emc_ECMcs_reg/NET0131 ,
		_w12306_,
		_w12307_
	);
	LUT2 #(
		.INIT('h1)
	) name8261 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w12308_
	);
	LUT2 #(
		.INIT('h2)
	) name8262 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		_w12309_
	);
	LUT2 #(
		.INIT('h1)
	) name8263 (
		_w12308_,
		_w12309_,
		_w12310_
	);
	LUT2 #(
		.INIT('h4)
	) name8264 (
		_w5608_,
		_w12310_,
		_w12311_
	);
	LUT2 #(
		.INIT('h1)
	) name8265 (
		_w12297_,
		_w12311_,
		_w12312_
	);
	LUT2 #(
		.INIT('h4)
	) name8266 (
		_w12307_,
		_w12312_,
		_w12313_
	);
	LUT2 #(
		.INIT('h1)
	) name8267 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12313_,
		_w12314_
	);
	LUT2 #(
		.INIT('h8)
	) name8268 (
		\bdma_BEAD_reg[13]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12315_
	);
	LUT2 #(
		.INIT('h1)
	) name8269 (
		_w12314_,
		_w12315_,
		_w12316_
	);
	LUT2 #(
		.INIT('h8)
	) name8270 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		_w5602_,
		_w12317_
	);
	LUT2 #(
		.INIT('h1)
	) name8271 (
		_w12281_,
		_w12299_,
		_w12318_
	);
	LUT2 #(
		.INIT('h2)
	) name8272 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w12318_,
		_w12319_
	);
	LUT2 #(
		.INIT('h2)
	) name8273 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w12320_
	);
	LUT2 #(
		.INIT('h8)
	) name8274 (
		_w12298_,
		_w12320_,
		_w12321_
	);
	LUT2 #(
		.INIT('h1)
	) name8275 (
		_w12319_,
		_w12321_,
		_w12322_
	);
	LUT2 #(
		.INIT('h2)
	) name8276 (
		_w12284_,
		_w12322_,
		_w12323_
	);
	LUT2 #(
		.INIT('h2)
	) name8277 (
		_w12275_,
		_w12282_,
		_w12324_
	);
	LUT2 #(
		.INIT('h8)
	) name8278 (
		_w12303_,
		_w12324_,
		_w12325_
	);
	LUT2 #(
		.INIT('h1)
	) name8279 (
		_w12323_,
		_w12325_,
		_w12326_
	);
	LUT2 #(
		.INIT('h2)
	) name8280 (
		\emc_ECMcs_reg/NET0131 ,
		_w12326_,
		_w12327_
	);
	LUT2 #(
		.INIT('h1)
	) name8281 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		_w12328_
	);
	LUT2 #(
		.INIT('h2)
	) name8282 (
		PM_bdry_sel_pad,
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w12329_
	);
	LUT2 #(
		.INIT('h1)
	) name8283 (
		_w12328_,
		_w12329_,
		_w12330_
	);
	LUT2 #(
		.INIT('h4)
	) name8284 (
		_w5608_,
		_w12330_,
		_w12331_
	);
	LUT2 #(
		.INIT('h1)
	) name8285 (
		_w12317_,
		_w12331_,
		_w12332_
	);
	LUT2 #(
		.INIT('h4)
	) name8286 (
		_w12327_,
		_w12332_,
		_w12333_
	);
	LUT2 #(
		.INIT('h1)
	) name8287 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12333_,
		_w12334_
	);
	LUT2 #(
		.INIT('h8)
	) name8288 (
		\bdma_BCTL_reg[8]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12335_
	);
	LUT2 #(
		.INIT('h1)
	) name8289 (
		_w12334_,
		_w12335_,
		_w12336_
	);
	LUT2 #(
		.INIT('h8)
	) name8290 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w5602_,
		_w12337_
	);
	LUT2 #(
		.INIT('h8)
	) name8291 (
		\sice_idr1_reg_DO_reg[5]/P0001 ,
		_w12248_,
		_w12338_
	);
	LUT2 #(
		.INIT('h8)
	) name8292 (
		\emc_ECMA_reg[1]/P0001 ,
		_w12250_,
		_w12339_
	);
	LUT2 #(
		.INIT('h2)
	) name8293 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		_w5608_,
		_w12340_
	);
	LUT2 #(
		.INIT('h8)
	) name8294 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w5610_,
		_w12341_
	);
	LUT2 #(
		.INIT('h1)
	) name8295 (
		_w12338_,
		_w12339_,
		_w12342_
	);
	LUT2 #(
		.INIT('h4)
	) name8296 (
		_w12337_,
		_w12342_,
		_w12343_
	);
	LUT2 #(
		.INIT('h1)
	) name8297 (
		_w12340_,
		_w12341_,
		_w12344_
	);
	LUT2 #(
		.INIT('h8)
	) name8298 (
		_w12343_,
		_w12344_,
		_w12345_
	);
	LUT2 #(
		.INIT('h1)
	) name8299 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12345_,
		_w12346_
	);
	LUT2 #(
		.INIT('h8)
	) name8300 (
		\bdma_BEAD_reg[1]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12347_
	);
	LUT2 #(
		.INIT('h1)
	) name8301 (
		_w12346_,
		_w12347_,
		_w12348_
	);
	LUT2 #(
		.INIT('h8)
	) name8302 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		_w5602_,
		_w12349_
	);
	LUT2 #(
		.INIT('h8)
	) name8303 (
		\sice_idr1_reg_DO_reg[6]/P0001 ,
		_w12248_,
		_w12350_
	);
	LUT2 #(
		.INIT('h8)
	) name8304 (
		\emc_ECMA_reg[2]/P0001 ,
		_w12250_,
		_w12351_
	);
	LUT2 #(
		.INIT('h2)
	) name8305 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		_w5608_,
		_w12352_
	);
	LUT2 #(
		.INIT('h8)
	) name8306 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w5610_,
		_w12353_
	);
	LUT2 #(
		.INIT('h1)
	) name8307 (
		_w12350_,
		_w12351_,
		_w12354_
	);
	LUT2 #(
		.INIT('h4)
	) name8308 (
		_w12349_,
		_w12354_,
		_w12355_
	);
	LUT2 #(
		.INIT('h1)
	) name8309 (
		_w12352_,
		_w12353_,
		_w12356_
	);
	LUT2 #(
		.INIT('h8)
	) name8310 (
		_w12355_,
		_w12356_,
		_w12357_
	);
	LUT2 #(
		.INIT('h1)
	) name8311 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12357_,
		_w12358_
	);
	LUT2 #(
		.INIT('h8)
	) name8312 (
		\bdma_BEAD_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12359_
	);
	LUT2 #(
		.INIT('h1)
	) name8313 (
		_w12358_,
		_w12359_,
		_w12360_
	);
	LUT2 #(
		.INIT('h8)
	) name8314 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w5602_,
		_w12361_
	);
	LUT2 #(
		.INIT('h8)
	) name8315 (
		\sice_idr1_reg_DO_reg[7]/P0001 ,
		_w12248_,
		_w12362_
	);
	LUT2 #(
		.INIT('h8)
	) name8316 (
		\emc_ECMA_reg[3]/P0001 ,
		_w12250_,
		_w12363_
	);
	LUT2 #(
		.INIT('h2)
	) name8317 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		_w5608_,
		_w12364_
	);
	LUT2 #(
		.INIT('h8)
	) name8318 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w5610_,
		_w12365_
	);
	LUT2 #(
		.INIT('h1)
	) name8319 (
		_w12362_,
		_w12363_,
		_w12366_
	);
	LUT2 #(
		.INIT('h4)
	) name8320 (
		_w12361_,
		_w12366_,
		_w12367_
	);
	LUT2 #(
		.INIT('h1)
	) name8321 (
		_w12364_,
		_w12365_,
		_w12368_
	);
	LUT2 #(
		.INIT('h8)
	) name8322 (
		_w12367_,
		_w12368_,
		_w12369_
	);
	LUT2 #(
		.INIT('h1)
	) name8323 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12369_,
		_w12370_
	);
	LUT2 #(
		.INIT('h8)
	) name8324 (
		\bdma_BEAD_reg[3]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12371_
	);
	LUT2 #(
		.INIT('h1)
	) name8325 (
		_w12370_,
		_w12371_,
		_w12372_
	);
	LUT2 #(
		.INIT('h8)
	) name8326 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5602_,
		_w12373_
	);
	LUT2 #(
		.INIT('h8)
	) name8327 (
		\sice_idr1_reg_DO_reg[8]/P0001 ,
		_w12248_,
		_w12374_
	);
	LUT2 #(
		.INIT('h8)
	) name8328 (
		\emc_ECMA_reg[4]/P0001 ,
		_w12250_,
		_w12375_
	);
	LUT2 #(
		.INIT('h2)
	) name8329 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		_w5608_,
		_w12376_
	);
	LUT2 #(
		.INIT('h8)
	) name8330 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w5610_,
		_w12377_
	);
	LUT2 #(
		.INIT('h1)
	) name8331 (
		_w12374_,
		_w12375_,
		_w12378_
	);
	LUT2 #(
		.INIT('h4)
	) name8332 (
		_w12373_,
		_w12378_,
		_w12379_
	);
	LUT2 #(
		.INIT('h1)
	) name8333 (
		_w12376_,
		_w12377_,
		_w12380_
	);
	LUT2 #(
		.INIT('h8)
	) name8334 (
		_w12379_,
		_w12380_,
		_w12381_
	);
	LUT2 #(
		.INIT('h1)
	) name8335 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12381_,
		_w12382_
	);
	LUT2 #(
		.INIT('h8)
	) name8336 (
		\bdma_BEAD_reg[4]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12383_
	);
	LUT2 #(
		.INIT('h1)
	) name8337 (
		_w12382_,
		_w12383_,
		_w12384_
	);
	LUT2 #(
		.INIT('h8)
	) name8338 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		_w5602_,
		_w12385_
	);
	LUT2 #(
		.INIT('h8)
	) name8339 (
		\sice_idr1_reg_DO_reg[9]/P0001 ,
		_w12248_,
		_w12386_
	);
	LUT2 #(
		.INIT('h8)
	) name8340 (
		\emc_ECMA_reg[5]/P0001 ,
		_w12250_,
		_w12387_
	);
	LUT2 #(
		.INIT('h2)
	) name8341 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		_w5608_,
		_w12388_
	);
	LUT2 #(
		.INIT('h8)
	) name8342 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w5610_,
		_w12389_
	);
	LUT2 #(
		.INIT('h1)
	) name8343 (
		_w12386_,
		_w12387_,
		_w12390_
	);
	LUT2 #(
		.INIT('h4)
	) name8344 (
		_w12385_,
		_w12390_,
		_w12391_
	);
	LUT2 #(
		.INIT('h1)
	) name8345 (
		_w12388_,
		_w12389_,
		_w12392_
	);
	LUT2 #(
		.INIT('h8)
	) name8346 (
		_w12391_,
		_w12392_,
		_w12393_
	);
	LUT2 #(
		.INIT('h1)
	) name8347 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12393_,
		_w12394_
	);
	LUT2 #(
		.INIT('h8)
	) name8348 (
		\bdma_BEAD_reg[5]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12395_
	);
	LUT2 #(
		.INIT('h1)
	) name8349 (
		_w12394_,
		_w12395_,
		_w12396_
	);
	LUT2 #(
		.INIT('h8)
	) name8350 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		_w5602_,
		_w12397_
	);
	LUT2 #(
		.INIT('h8)
	) name8351 (
		\sice_idr1_reg_DO_reg[10]/P0001 ,
		_w12248_,
		_w12398_
	);
	LUT2 #(
		.INIT('h8)
	) name8352 (
		\emc_ECMA_reg[6]/P0001 ,
		_w12250_,
		_w12399_
	);
	LUT2 #(
		.INIT('h2)
	) name8353 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		_w5608_,
		_w12400_
	);
	LUT2 #(
		.INIT('h8)
	) name8354 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w5610_,
		_w12401_
	);
	LUT2 #(
		.INIT('h1)
	) name8355 (
		_w12398_,
		_w12399_,
		_w12402_
	);
	LUT2 #(
		.INIT('h4)
	) name8356 (
		_w12397_,
		_w12402_,
		_w12403_
	);
	LUT2 #(
		.INIT('h1)
	) name8357 (
		_w12400_,
		_w12401_,
		_w12404_
	);
	LUT2 #(
		.INIT('h8)
	) name8358 (
		_w12403_,
		_w12404_,
		_w12405_
	);
	LUT2 #(
		.INIT('h1)
	) name8359 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12405_,
		_w12406_
	);
	LUT2 #(
		.INIT('h8)
	) name8360 (
		\bdma_BEAD_reg[6]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12407_
	);
	LUT2 #(
		.INIT('h1)
	) name8361 (
		_w12406_,
		_w12407_,
		_w12408_
	);
	LUT2 #(
		.INIT('h8)
	) name8362 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		_w5602_,
		_w12409_
	);
	LUT2 #(
		.INIT('h8)
	) name8363 (
		\sice_idr1_reg_DO_reg[11]/P0001 ,
		_w12248_,
		_w12410_
	);
	LUT2 #(
		.INIT('h8)
	) name8364 (
		\emc_ECMA_reg[7]/P0001 ,
		_w12250_,
		_w12411_
	);
	LUT2 #(
		.INIT('h2)
	) name8365 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		_w5608_,
		_w12412_
	);
	LUT2 #(
		.INIT('h8)
	) name8366 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w5610_,
		_w12413_
	);
	LUT2 #(
		.INIT('h1)
	) name8367 (
		_w12410_,
		_w12411_,
		_w12414_
	);
	LUT2 #(
		.INIT('h4)
	) name8368 (
		_w12409_,
		_w12414_,
		_w12415_
	);
	LUT2 #(
		.INIT('h1)
	) name8369 (
		_w12412_,
		_w12413_,
		_w12416_
	);
	LUT2 #(
		.INIT('h8)
	) name8370 (
		_w12415_,
		_w12416_,
		_w12417_
	);
	LUT2 #(
		.INIT('h1)
	) name8371 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12417_,
		_w12418_
	);
	LUT2 #(
		.INIT('h8)
	) name8372 (
		\bdma_BEAD_reg[7]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12419_
	);
	LUT2 #(
		.INIT('h1)
	) name8373 (
		_w12418_,
		_w12419_,
		_w12420_
	);
	LUT2 #(
		.INIT('h8)
	) name8374 (
		\bdma_BEAD_reg[8]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12421_
	);
	LUT2 #(
		.INIT('h8)
	) name8375 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		_w5602_,
		_w12422_
	);
	LUT2 #(
		.INIT('h2)
	) name8376 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		_w5608_,
		_w12423_
	);
	LUT2 #(
		.INIT('h8)
	) name8377 (
		\emc_ECMA_reg[8]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w12424_
	);
	LUT2 #(
		.INIT('h8)
	) name8378 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w5610_,
		_w12425_
	);
	LUT2 #(
		.INIT('h1)
	) name8379 (
		_w12422_,
		_w12424_,
		_w12426_
	);
	LUT2 #(
		.INIT('h1)
	) name8380 (
		_w12423_,
		_w12425_,
		_w12427_
	);
	LUT2 #(
		.INIT('h8)
	) name8381 (
		_w12426_,
		_w12427_,
		_w12428_
	);
	LUT2 #(
		.INIT('h1)
	) name8382 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12428_,
		_w12429_
	);
	LUT2 #(
		.INIT('h1)
	) name8383 (
		_w12421_,
		_w12429_,
		_w12430_
	);
	LUT2 #(
		.INIT('h8)
	) name8384 (
		\bdma_BEAD_reg[9]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12431_
	);
	LUT2 #(
		.INIT('h8)
	) name8385 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		_w5602_,
		_w12432_
	);
	LUT2 #(
		.INIT('h2)
	) name8386 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		_w5608_,
		_w12433_
	);
	LUT2 #(
		.INIT('h8)
	) name8387 (
		\emc_ECMA_reg[9]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w12434_
	);
	LUT2 #(
		.INIT('h8)
	) name8388 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w5610_,
		_w12435_
	);
	LUT2 #(
		.INIT('h1)
	) name8389 (
		_w12432_,
		_w12434_,
		_w12436_
	);
	LUT2 #(
		.INIT('h1)
	) name8390 (
		_w12433_,
		_w12435_,
		_w12437_
	);
	LUT2 #(
		.INIT('h8)
	) name8391 (
		_w12436_,
		_w12437_,
		_w12438_
	);
	LUT2 #(
		.INIT('h1)
	) name8392 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12438_,
		_w12439_
	);
	LUT2 #(
		.INIT('h1)
	) name8393 (
		_w12431_,
		_w12439_,
		_w12440_
	);
	LUT2 #(
		.INIT('h1)
	) name8394 (
		_w5602_,
		_w5610_,
		_w12441_
	);
	LUT2 #(
		.INIT('h2)
	) name8395 (
		\core_c_dec_accCM_E_reg/NET0131 ,
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w12442_
	);
	LUT2 #(
		.INIT('h8)
	) name8396 (
		_w12247_,
		_w12442_,
		_w12443_
	);
	LUT2 #(
		.INIT('h4)
	) name8397 (
		\emc_ECS_reg[1]/NET0131 ,
		_w5523_,
		_w12444_
	);
	LUT2 #(
		.INIT('h1)
	) name8398 (
		\bdma_BM_cyc_reg/P0001 ,
		_w5519_,
		_w12445_
	);
	LUT2 #(
		.INIT('h4)
	) name8399 (
		_w12443_,
		_w12445_,
		_w12446_
	);
	LUT2 #(
		.INIT('h4)
	) name8400 (
		_w12444_,
		_w12446_,
		_w12447_
	);
	LUT2 #(
		.INIT('h8)
	) name8401 (
		_w5608_,
		_w12447_,
		_w12448_
	);
	LUT2 #(
		.INIT('h8)
	) name8402 (
		_w12441_,
		_w12448_,
		_w12449_
	);
	LUT2 #(
		.INIT('h1)
	) name8403 (
		\core_c_psq_MGNT_reg/NET0131 ,
		_w12449_,
		_w12450_
	);
	LUT2 #(
		.INIT('h4)
	) name8404 (
		\core_c_psq_MGNT_reg/NET0131 ,
		\emc_ED_oei_reg/P0001 ,
		_w12451_
	);
	LUT2 #(
		.INIT('h2)
	) name8405 (
		\emc_selPMDi_reg/P0001 ,
		_w5608_,
		_w12452_
	);
	LUT2 #(
		.INIT('h2)
	) name8406 (
		\emc_selDMDi_reg/P0001 ,
		_w12441_,
		_w12453_
	);
	LUT2 #(
		.INIT('h1)
	) name8407 (
		_w12452_,
		_w12453_,
		_w12454_
	);
	LUT2 #(
		.INIT('h8)
	) name8408 (
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w12454_,
		_w12455_
	);
	LUT2 #(
		.INIT('h4)
	) name8409 (
		_w12452_,
		_w12453_,
		_w12456_
	);
	LUT2 #(
		.INIT('h8)
	) name8410 (
		_w7607_,
		_w12456_,
		_w12457_
	);
	LUT2 #(
		.INIT('h8)
	) name8411 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[0]/P0001 ,
		_w12458_
	);
	LUT2 #(
		.INIT('h1)
	) name8412 (
		\memc_PMo_oe2_reg/P0001 ,
		\memc_PMo_oe3_reg/P0001 ,
		_w12459_
	);
	LUT2 #(
		.INIT('h1)
	) name8413 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		_w12460_
	);
	LUT2 #(
		.INIT('h4)
	) name8414 (
		\memc_PMo_oe6_reg/P0001 ,
		_w12460_,
		_w12461_
	);
	LUT2 #(
		.INIT('h4)
	) name8415 (
		\memc_PMo_oe7_reg/P0001 ,
		_w12461_,
		_w12462_
	);
	LUT2 #(
		.INIT('h1)
	) name8416 (
		\memc_PMo_oe0_reg/P0001 ,
		\memc_PMo_oe1_reg/P0001 ,
		_w12463_
	);
	LUT2 #(
		.INIT('h8)
	) name8417 (
		_w12462_,
		_w12463_,
		_w12464_
	);
	LUT2 #(
		.INIT('h8)
	) name8418 (
		_w12459_,
		_w12464_,
		_w12465_
	);
	LUT2 #(
		.INIT('h2)
	) name8419 (
		\core_c_dec_pMFSHT_Ei_reg/NET0131 ,
		_w6988_,
		_w12466_
	);
	LUT2 #(
		.INIT('h4)
	) name8420 (
		_w7386_,
		_w12466_,
		_w12467_
	);
	LUT2 #(
		.INIT('h2)
	) name8421 (
		\core_c_dec_pMFALU_Ei_reg/NET0131 ,
		_w6988_,
		_w12468_
	);
	LUT2 #(
		.INIT('h4)
	) name8422 (
		_w7437_,
		_w12468_,
		_w12469_
	);
	LUT2 #(
		.INIT('h2)
	) name8423 (
		\core_c_dec_pMFMAC_Ei_reg/NET0131 ,
		_w6988_,
		_w12470_
	);
	LUT2 #(
		.INIT('h4)
	) name8424 (
		_w7480_,
		_w12470_,
		_w12471_
	);
	LUT2 #(
		.INIT('h1)
	) name8425 (
		_w12467_,
		_w12469_,
		_w12472_
	);
	LUT2 #(
		.INIT('h4)
	) name8426 (
		_w12471_,
		_w12472_,
		_w12473_
	);
	LUT2 #(
		.INIT('h1)
	) name8427 (
		\emc_PMDoe_reg/NET0131 ,
		_w12473_,
		_w12474_
	);
	LUT2 #(
		.INIT('h4)
	) name8428 (
		_w12458_,
		_w12465_,
		_w12475_
	);
	LUT2 #(
		.INIT('h4)
	) name8429 (
		_w12474_,
		_w12475_,
		_w12476_
	);
	LUT2 #(
		.INIT('h2)
	) name8430 (
		\memc_PMo_oe2_reg/P0001 ,
		\memc_PMo_oe3_reg/P0001 ,
		_w12477_
	);
	LUT2 #(
		.INIT('h8)
	) name8431 (
		_w12464_,
		_w12477_,
		_w12478_
	);
	LUT2 #(
		.INIT('h8)
	) name8432 (
		\PM_rd2[0]_pad ,
		_w12478_,
		_w12479_
	);
	LUT2 #(
		.INIT('h8)
	) name8433 (
		_w12459_,
		_w12463_,
		_w12480_
	);
	LUT2 #(
		.INIT('h4)
	) name8434 (
		\memc_PMo_oe7_reg/P0001 ,
		_w12480_,
		_w12481_
	);
	LUT2 #(
		.INIT('h8)
	) name8435 (
		\memc_PMo_oe6_reg/P0001 ,
		_w12460_,
		_w12482_
	);
	LUT2 #(
		.INIT('h8)
	) name8436 (
		_w12481_,
		_w12482_,
		_w12483_
	);
	LUT2 #(
		.INIT('h8)
	) name8437 (
		\memc_PMo_oe7_reg/P0001 ,
		_w12461_,
		_w12484_
	);
	LUT2 #(
		.INIT('h8)
	) name8438 (
		_w12480_,
		_w12484_,
		_w12485_
	);
	LUT2 #(
		.INIT('h4)
	) name8439 (
		\memc_PMo_oe6_reg/P0001 ,
		_w12481_,
		_w12486_
	);
	LUT2 #(
		.INIT('h2)
	) name8440 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		_w12487_
	);
	LUT2 #(
		.INIT('h8)
	) name8441 (
		_w12486_,
		_w12487_,
		_w12488_
	);
	LUT2 #(
		.INIT('h8)
	) name8442 (
		_w12459_,
		_w12462_,
		_w12489_
	);
	LUT2 #(
		.INIT('h4)
	) name8443 (
		\memc_PMo_oe0_reg/P0001 ,
		\memc_PMo_oe1_reg/P0001 ,
		_w12490_
	);
	LUT2 #(
		.INIT('h8)
	) name8444 (
		_w12489_,
		_w12490_,
		_w12491_
	);
	LUT2 #(
		.INIT('h4)
	) name8445 (
		\memc_PMo_oe2_reg/P0001 ,
		\memc_PMo_oe3_reg/P0001 ,
		_w12492_
	);
	LUT2 #(
		.INIT('h8)
	) name8446 (
		_w12464_,
		_w12492_,
		_w12493_
	);
	LUT2 #(
		.INIT('h4)
	) name8447 (
		\memc_PMo_oe4_reg/P0001 ,
		\memc_PMo_oe5_reg/P0001 ,
		_w12494_
	);
	LUT2 #(
		.INIT('h8)
	) name8448 (
		_w12486_,
		_w12494_,
		_w12495_
	);
	LUT2 #(
		.INIT('h1)
	) name8449 (
		_w12483_,
		_w12485_,
		_w12496_
	);
	LUT2 #(
		.INIT('h4)
	) name8450 (
		_w12478_,
		_w12496_,
		_w12497_
	);
	LUT2 #(
		.INIT('h1)
	) name8451 (
		_w12488_,
		_w12491_,
		_w12498_
	);
	LUT2 #(
		.INIT('h1)
	) name8452 (
		_w12493_,
		_w12495_,
		_w12499_
	);
	LUT2 #(
		.INIT('h8)
	) name8453 (
		_w12498_,
		_w12499_,
		_w12500_
	);
	LUT2 #(
		.INIT('h8)
	) name8454 (
		_w12497_,
		_w12500_,
		_w12501_
	);
	LUT2 #(
		.INIT('h2)
	) name8455 (
		\memc_PMo_oe0_reg/P0001 ,
		\memc_PMo_oe1_reg/P0001 ,
		_w12502_
	);
	LUT2 #(
		.INIT('h8)
	) name8456 (
		_w12489_,
		_w12502_,
		_w12503_
	);
	LUT2 #(
		.INIT('h1)
	) name8457 (
		_w12501_,
		_w12503_,
		_w12504_
	);
	LUT2 #(
		.INIT('h2)
	) name8458 (
		\PM_rd0[0]_pad ,
		_w12504_,
		_w12505_
	);
	LUT2 #(
		.INIT('h8)
	) name8459 (
		\PM_rd4[0]_pad ,
		_w12488_,
		_w12506_
	);
	LUT2 #(
		.INIT('h8)
	) name8460 (
		\PM_rd6[0]_pad ,
		_w12483_,
		_w12507_
	);
	LUT2 #(
		.INIT('h8)
	) name8461 (
		\PM_rd7[0]_pad ,
		_w12485_,
		_w12508_
	);
	LUT2 #(
		.INIT('h8)
	) name8462 (
		\PM_rd3[0]_pad ,
		_w12493_,
		_w12509_
	);
	LUT2 #(
		.INIT('h8)
	) name8463 (
		\PM_rd1[0]_pad ,
		_w12491_,
		_w12510_
	);
	LUT2 #(
		.INIT('h8)
	) name8464 (
		\PM_rd5[0]_pad ,
		_w12495_,
		_w12511_
	);
	LUT2 #(
		.INIT('h1)
	) name8465 (
		_w12465_,
		_w12507_,
		_w12512_
	);
	LUT2 #(
		.INIT('h4)
	) name8466 (
		_w12508_,
		_w12512_,
		_w12513_
	);
	LUT2 #(
		.INIT('h1)
	) name8467 (
		_w12479_,
		_w12506_,
		_w12514_
	);
	LUT2 #(
		.INIT('h1)
	) name8468 (
		_w12509_,
		_w12510_,
		_w12515_
	);
	LUT2 #(
		.INIT('h4)
	) name8469 (
		_w12511_,
		_w12515_,
		_w12516_
	);
	LUT2 #(
		.INIT('h8)
	) name8470 (
		_w12513_,
		_w12514_,
		_w12517_
	);
	LUT2 #(
		.INIT('h8)
	) name8471 (
		_w12516_,
		_w12517_,
		_w12518_
	);
	LUT2 #(
		.INIT('h4)
	) name8472 (
		_w12505_,
		_w12518_,
		_w12519_
	);
	LUT2 #(
		.INIT('h1)
	) name8473 (
		_w12476_,
		_w12519_,
		_w12520_
	);
	LUT2 #(
		.INIT('h8)
	) name8474 (
		_w12452_,
		_w12520_,
		_w12521_
	);
	LUT2 #(
		.INIT('h1)
	) name8475 (
		_w12455_,
		_w12521_,
		_w12522_
	);
	LUT2 #(
		.INIT('h4)
	) name8476 (
		_w12457_,
		_w12522_,
		_w12523_
	);
	LUT2 #(
		.INIT('h2)
	) name8477 (
		_w12451_,
		_w12523_,
		_w12524_
	);
	LUT2 #(
		.INIT('h8)
	) name8478 (
		\bdma_BCTL_reg[2]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12525_
	);
	LUT2 #(
		.INIT('h8)
	) name8479 (
		\bdma_BWdataBUF_reg[0]/P0001 ,
		_w12525_,
		_w12526_
	);
	LUT2 #(
		.INIT('h1)
	) name8480 (
		_w12524_,
		_w12526_,
		_w12527_
	);
	LUT2 #(
		.INIT('h8)
	) name8481 (
		\bdma_BCTL_reg[11]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12528_
	);
	LUT2 #(
		.INIT('h8)
	) name8482 (
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w12454_,
		_w12529_
	);
	LUT2 #(
		.INIT('h8)
	) name8483 (
		_w7859_,
		_w12456_,
		_w12530_
	);
	LUT2 #(
		.INIT('h8)
	) name8484 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[10]/P0001 ,
		_w12531_
	);
	LUT2 #(
		.INIT('h4)
	) name8485 (
		_w7764_,
		_w12470_,
		_w12532_
	);
	LUT2 #(
		.INIT('h4)
	) name8486 (
		_w7813_,
		_w12466_,
		_w12533_
	);
	LUT2 #(
		.INIT('h4)
	) name8487 (
		_w7789_,
		_w12468_,
		_w12534_
	);
	LUT2 #(
		.INIT('h1)
	) name8488 (
		_w12532_,
		_w12533_,
		_w12535_
	);
	LUT2 #(
		.INIT('h4)
	) name8489 (
		_w12534_,
		_w12535_,
		_w12536_
	);
	LUT2 #(
		.INIT('h1)
	) name8490 (
		\emc_PMDoe_reg/NET0131 ,
		_w12536_,
		_w12537_
	);
	LUT2 #(
		.INIT('h2)
	) name8491 (
		_w12465_,
		_w12531_,
		_w12538_
	);
	LUT2 #(
		.INIT('h4)
	) name8492 (
		_w12537_,
		_w12538_,
		_w12539_
	);
	LUT2 #(
		.INIT('h8)
	) name8493 (
		\PM_rd2[10]_pad ,
		_w12478_,
		_w12540_
	);
	LUT2 #(
		.INIT('h2)
	) name8494 (
		\PM_rd0[10]_pad ,
		_w12504_,
		_w12541_
	);
	LUT2 #(
		.INIT('h8)
	) name8495 (
		\PM_rd4[10]_pad ,
		_w12488_,
		_w12542_
	);
	LUT2 #(
		.INIT('h8)
	) name8496 (
		\PM_rd6[10]_pad ,
		_w12483_,
		_w12543_
	);
	LUT2 #(
		.INIT('h8)
	) name8497 (
		\PM_rd7[10]_pad ,
		_w12485_,
		_w12544_
	);
	LUT2 #(
		.INIT('h8)
	) name8498 (
		\PM_rd3[10]_pad ,
		_w12493_,
		_w12545_
	);
	LUT2 #(
		.INIT('h8)
	) name8499 (
		\PM_rd1[10]_pad ,
		_w12491_,
		_w12546_
	);
	LUT2 #(
		.INIT('h8)
	) name8500 (
		\PM_rd5[10]_pad ,
		_w12495_,
		_w12547_
	);
	LUT2 #(
		.INIT('h1)
	) name8501 (
		_w12465_,
		_w12543_,
		_w12548_
	);
	LUT2 #(
		.INIT('h4)
	) name8502 (
		_w12544_,
		_w12548_,
		_w12549_
	);
	LUT2 #(
		.INIT('h1)
	) name8503 (
		_w12540_,
		_w12542_,
		_w12550_
	);
	LUT2 #(
		.INIT('h1)
	) name8504 (
		_w12545_,
		_w12546_,
		_w12551_
	);
	LUT2 #(
		.INIT('h4)
	) name8505 (
		_w12547_,
		_w12551_,
		_w12552_
	);
	LUT2 #(
		.INIT('h8)
	) name8506 (
		_w12549_,
		_w12550_,
		_w12553_
	);
	LUT2 #(
		.INIT('h8)
	) name8507 (
		_w12552_,
		_w12553_,
		_w12554_
	);
	LUT2 #(
		.INIT('h4)
	) name8508 (
		_w12541_,
		_w12554_,
		_w12555_
	);
	LUT2 #(
		.INIT('h1)
	) name8509 (
		_w12539_,
		_w12555_,
		_w12556_
	);
	LUT2 #(
		.INIT('h8)
	) name8510 (
		_w12452_,
		_w12556_,
		_w12557_
	);
	LUT2 #(
		.INIT('h1)
	) name8511 (
		_w12529_,
		_w12557_,
		_w12558_
	);
	LUT2 #(
		.INIT('h4)
	) name8512 (
		_w12530_,
		_w12558_,
		_w12559_
	);
	LUT2 #(
		.INIT('h2)
	) name8513 (
		_w12451_,
		_w12559_,
		_w12560_
	);
	LUT2 #(
		.INIT('h1)
	) name8514 (
		_w12528_,
		_w12560_,
		_w12561_
	);
	LUT2 #(
		.INIT('h8)
	) name8515 (
		\bdma_BCTL_reg[12]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12562_
	);
	LUT2 #(
		.INIT('h8)
	) name8516 (
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w12454_,
		_w12563_
	);
	LUT2 #(
		.INIT('h8)
	) name8517 (
		_w8460_,
		_w12456_,
		_w12564_
	);
	LUT2 #(
		.INIT('h8)
	) name8518 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[11]/P0001 ,
		_w12565_
	);
	LUT2 #(
		.INIT('h4)
	) name8519 (
		_w8365_,
		_w12470_,
		_w12566_
	);
	LUT2 #(
		.INIT('h4)
	) name8520 (
		_w8414_,
		_w12466_,
		_w12567_
	);
	LUT2 #(
		.INIT('h4)
	) name8521 (
		_w8390_,
		_w12468_,
		_w12568_
	);
	LUT2 #(
		.INIT('h1)
	) name8522 (
		_w12566_,
		_w12567_,
		_w12569_
	);
	LUT2 #(
		.INIT('h4)
	) name8523 (
		_w12568_,
		_w12569_,
		_w12570_
	);
	LUT2 #(
		.INIT('h1)
	) name8524 (
		\emc_PMDoe_reg/NET0131 ,
		_w12570_,
		_w12571_
	);
	LUT2 #(
		.INIT('h2)
	) name8525 (
		_w12465_,
		_w12565_,
		_w12572_
	);
	LUT2 #(
		.INIT('h4)
	) name8526 (
		_w12571_,
		_w12572_,
		_w12573_
	);
	LUT2 #(
		.INIT('h8)
	) name8527 (
		\PM_rd2[11]_pad ,
		_w12478_,
		_w12574_
	);
	LUT2 #(
		.INIT('h2)
	) name8528 (
		\PM_rd0[11]_pad ,
		_w12504_,
		_w12575_
	);
	LUT2 #(
		.INIT('h8)
	) name8529 (
		\PM_rd4[11]_pad ,
		_w12488_,
		_w12576_
	);
	LUT2 #(
		.INIT('h8)
	) name8530 (
		\PM_rd6[11]_pad ,
		_w12483_,
		_w12577_
	);
	LUT2 #(
		.INIT('h8)
	) name8531 (
		\PM_rd7[11]_pad ,
		_w12485_,
		_w12578_
	);
	LUT2 #(
		.INIT('h8)
	) name8532 (
		\PM_rd3[11]_pad ,
		_w12493_,
		_w12579_
	);
	LUT2 #(
		.INIT('h8)
	) name8533 (
		\PM_rd1[11]_pad ,
		_w12491_,
		_w12580_
	);
	LUT2 #(
		.INIT('h8)
	) name8534 (
		\PM_rd5[11]_pad ,
		_w12495_,
		_w12581_
	);
	LUT2 #(
		.INIT('h1)
	) name8535 (
		_w12465_,
		_w12577_,
		_w12582_
	);
	LUT2 #(
		.INIT('h4)
	) name8536 (
		_w12578_,
		_w12582_,
		_w12583_
	);
	LUT2 #(
		.INIT('h1)
	) name8537 (
		_w12574_,
		_w12576_,
		_w12584_
	);
	LUT2 #(
		.INIT('h1)
	) name8538 (
		_w12579_,
		_w12580_,
		_w12585_
	);
	LUT2 #(
		.INIT('h4)
	) name8539 (
		_w12581_,
		_w12585_,
		_w12586_
	);
	LUT2 #(
		.INIT('h8)
	) name8540 (
		_w12583_,
		_w12584_,
		_w12587_
	);
	LUT2 #(
		.INIT('h8)
	) name8541 (
		_w12586_,
		_w12587_,
		_w12588_
	);
	LUT2 #(
		.INIT('h4)
	) name8542 (
		_w12575_,
		_w12588_,
		_w12589_
	);
	LUT2 #(
		.INIT('h1)
	) name8543 (
		_w12573_,
		_w12589_,
		_w12590_
	);
	LUT2 #(
		.INIT('h8)
	) name8544 (
		_w12452_,
		_w12590_,
		_w12591_
	);
	LUT2 #(
		.INIT('h1)
	) name8545 (
		_w12563_,
		_w12591_,
		_w12592_
	);
	LUT2 #(
		.INIT('h4)
	) name8546 (
		_w12564_,
		_w12592_,
		_w12593_
	);
	LUT2 #(
		.INIT('h2)
	) name8547 (
		_w12451_,
		_w12593_,
		_w12594_
	);
	LUT2 #(
		.INIT('h1)
	) name8548 (
		_w12562_,
		_w12594_,
		_w12595_
	);
	LUT2 #(
		.INIT('h8)
	) name8549 (
		\bdma_BCTL_reg[13]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12596_
	);
	LUT2 #(
		.INIT('h8)
	) name8550 (
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w12454_,
		_w12597_
	);
	LUT2 #(
		.INIT('h8)
	) name8551 (
		_w9178_,
		_w12456_,
		_w12598_
	);
	LUT2 #(
		.INIT('h8)
	) name8552 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[12]/P0001 ,
		_w12599_
	);
	LUT2 #(
		.INIT('h4)
	) name8553 (
		_w9083_,
		_w12470_,
		_w12600_
	);
	LUT2 #(
		.INIT('h4)
	) name8554 (
		_w9132_,
		_w12466_,
		_w12601_
	);
	LUT2 #(
		.INIT('h4)
	) name8555 (
		_w9108_,
		_w12468_,
		_w12602_
	);
	LUT2 #(
		.INIT('h1)
	) name8556 (
		_w12600_,
		_w12601_,
		_w12603_
	);
	LUT2 #(
		.INIT('h4)
	) name8557 (
		_w12602_,
		_w12603_,
		_w12604_
	);
	LUT2 #(
		.INIT('h1)
	) name8558 (
		\emc_PMDoe_reg/NET0131 ,
		_w12604_,
		_w12605_
	);
	LUT2 #(
		.INIT('h2)
	) name8559 (
		_w12465_,
		_w12599_,
		_w12606_
	);
	LUT2 #(
		.INIT('h4)
	) name8560 (
		_w12605_,
		_w12606_,
		_w12607_
	);
	LUT2 #(
		.INIT('h8)
	) name8561 (
		\PM_rd2[12]_pad ,
		_w12478_,
		_w12608_
	);
	LUT2 #(
		.INIT('h2)
	) name8562 (
		\PM_rd0[12]_pad ,
		_w12504_,
		_w12609_
	);
	LUT2 #(
		.INIT('h8)
	) name8563 (
		\PM_rd4[12]_pad ,
		_w12488_,
		_w12610_
	);
	LUT2 #(
		.INIT('h8)
	) name8564 (
		\PM_rd6[12]_pad ,
		_w12483_,
		_w12611_
	);
	LUT2 #(
		.INIT('h8)
	) name8565 (
		\PM_rd7[12]_pad ,
		_w12485_,
		_w12612_
	);
	LUT2 #(
		.INIT('h8)
	) name8566 (
		\PM_rd3[12]_pad ,
		_w12493_,
		_w12613_
	);
	LUT2 #(
		.INIT('h8)
	) name8567 (
		\PM_rd1[12]_pad ,
		_w12491_,
		_w12614_
	);
	LUT2 #(
		.INIT('h8)
	) name8568 (
		\PM_rd5[12]_pad ,
		_w12495_,
		_w12615_
	);
	LUT2 #(
		.INIT('h1)
	) name8569 (
		_w12465_,
		_w12611_,
		_w12616_
	);
	LUT2 #(
		.INIT('h4)
	) name8570 (
		_w12612_,
		_w12616_,
		_w12617_
	);
	LUT2 #(
		.INIT('h1)
	) name8571 (
		_w12608_,
		_w12610_,
		_w12618_
	);
	LUT2 #(
		.INIT('h1)
	) name8572 (
		_w12613_,
		_w12614_,
		_w12619_
	);
	LUT2 #(
		.INIT('h4)
	) name8573 (
		_w12615_,
		_w12619_,
		_w12620_
	);
	LUT2 #(
		.INIT('h8)
	) name8574 (
		_w12617_,
		_w12618_,
		_w12621_
	);
	LUT2 #(
		.INIT('h8)
	) name8575 (
		_w12620_,
		_w12621_,
		_w12622_
	);
	LUT2 #(
		.INIT('h4)
	) name8576 (
		_w12609_,
		_w12622_,
		_w12623_
	);
	LUT2 #(
		.INIT('h1)
	) name8577 (
		_w12607_,
		_w12623_,
		_w12624_
	);
	LUT2 #(
		.INIT('h8)
	) name8578 (
		_w12452_,
		_w12624_,
		_w12625_
	);
	LUT2 #(
		.INIT('h1)
	) name8579 (
		_w12597_,
		_w12625_,
		_w12626_
	);
	LUT2 #(
		.INIT('h4)
	) name8580 (
		_w12598_,
		_w12626_,
		_w12627_
	);
	LUT2 #(
		.INIT('h2)
	) name8581 (
		_w12451_,
		_w12627_,
		_w12628_
	);
	LUT2 #(
		.INIT('h1)
	) name8582 (
		_w12596_,
		_w12628_,
		_w12629_
	);
	LUT2 #(
		.INIT('h8)
	) name8583 (
		\bdma_BCTL_reg[14]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12630_
	);
	LUT2 #(
		.INIT('h8)
	) name8584 (
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w12454_,
		_w12631_
	);
	LUT2 #(
		.INIT('h8)
	) name8585 (
		_w7340_,
		_w12456_,
		_w12632_
	);
	LUT2 #(
		.INIT('h8)
	) name8586 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[13]/P0001 ,
		_w12633_
	);
	LUT2 #(
		.INIT('h4)
	) name8587 (
		_w7213_,
		_w12470_,
		_w12634_
	);
	LUT2 #(
		.INIT('h4)
	) name8588 (
		_w7177_,
		_w12466_,
		_w12635_
	);
	LUT2 #(
		.INIT('h4)
	) name8589 (
		_w7117_,
		_w12468_,
		_w12636_
	);
	LUT2 #(
		.INIT('h1)
	) name8590 (
		_w12634_,
		_w12635_,
		_w12637_
	);
	LUT2 #(
		.INIT('h4)
	) name8591 (
		_w12636_,
		_w12637_,
		_w12638_
	);
	LUT2 #(
		.INIT('h1)
	) name8592 (
		\emc_PMDoe_reg/NET0131 ,
		_w12638_,
		_w12639_
	);
	LUT2 #(
		.INIT('h2)
	) name8593 (
		_w12465_,
		_w12633_,
		_w12640_
	);
	LUT2 #(
		.INIT('h4)
	) name8594 (
		_w12639_,
		_w12640_,
		_w12641_
	);
	LUT2 #(
		.INIT('h8)
	) name8595 (
		\PM_rd2[13]_pad ,
		_w12478_,
		_w12642_
	);
	LUT2 #(
		.INIT('h2)
	) name8596 (
		\PM_rd0[13]_pad ,
		_w12504_,
		_w12643_
	);
	LUT2 #(
		.INIT('h8)
	) name8597 (
		\PM_rd4[13]_pad ,
		_w12488_,
		_w12644_
	);
	LUT2 #(
		.INIT('h8)
	) name8598 (
		\PM_rd6[13]_pad ,
		_w12483_,
		_w12645_
	);
	LUT2 #(
		.INIT('h8)
	) name8599 (
		\PM_rd7[13]_pad ,
		_w12485_,
		_w12646_
	);
	LUT2 #(
		.INIT('h8)
	) name8600 (
		\PM_rd3[13]_pad ,
		_w12493_,
		_w12647_
	);
	LUT2 #(
		.INIT('h8)
	) name8601 (
		\PM_rd1[13]_pad ,
		_w12491_,
		_w12648_
	);
	LUT2 #(
		.INIT('h8)
	) name8602 (
		\PM_rd5[13]_pad ,
		_w12495_,
		_w12649_
	);
	LUT2 #(
		.INIT('h1)
	) name8603 (
		_w12465_,
		_w12645_,
		_w12650_
	);
	LUT2 #(
		.INIT('h4)
	) name8604 (
		_w12646_,
		_w12650_,
		_w12651_
	);
	LUT2 #(
		.INIT('h1)
	) name8605 (
		_w12642_,
		_w12644_,
		_w12652_
	);
	LUT2 #(
		.INIT('h1)
	) name8606 (
		_w12647_,
		_w12648_,
		_w12653_
	);
	LUT2 #(
		.INIT('h4)
	) name8607 (
		_w12649_,
		_w12653_,
		_w12654_
	);
	LUT2 #(
		.INIT('h8)
	) name8608 (
		_w12651_,
		_w12652_,
		_w12655_
	);
	LUT2 #(
		.INIT('h8)
	) name8609 (
		_w12654_,
		_w12655_,
		_w12656_
	);
	LUT2 #(
		.INIT('h4)
	) name8610 (
		_w12643_,
		_w12656_,
		_w12657_
	);
	LUT2 #(
		.INIT('h1)
	) name8611 (
		_w12641_,
		_w12657_,
		_w12658_
	);
	LUT2 #(
		.INIT('h8)
	) name8612 (
		_w12452_,
		_w12658_,
		_w12659_
	);
	LUT2 #(
		.INIT('h1)
	) name8613 (
		_w12631_,
		_w12659_,
		_w12660_
	);
	LUT2 #(
		.INIT('h4)
	) name8614 (
		_w12632_,
		_w12660_,
		_w12661_
	);
	LUT2 #(
		.INIT('h2)
	) name8615 (
		_w12451_,
		_w12661_,
		_w12662_
	);
	LUT2 #(
		.INIT('h1)
	) name8616 (
		_w12630_,
		_w12662_,
		_w12663_
	);
	LUT2 #(
		.INIT('h8)
	) name8617 (
		\bdma_BCTL_reg[15]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w12664_
	);
	LUT2 #(
		.INIT('h8)
	) name8618 (
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w12454_,
		_w12665_
	);
	LUT2 #(
		.INIT('h8)
	) name8619 (
		\DM_rdm[14]_pad ,
		_w7016_,
		_w12666_
	);
	LUT2 #(
		.INIT('h8)
	) name8620 (
		\DM_rd1[14]_pad ,
		_w7022_,
		_w12667_
	);
	LUT2 #(
		.INIT('h8)
	) name8621 (
		\DM_rd4[14]_pad ,
		_w7028_,
		_w12668_
	);
	LUT2 #(
		.INIT('h8)
	) name8622 (
		\DM_rd6[14]_pad ,
		_w7031_,
		_w12669_
	);
	LUT2 #(
		.INIT('h8)
	) name8623 (
		\DM_rd7[14]_pad ,
		_w7034_,
		_w12670_
	);
	LUT2 #(
		.INIT('h8)
	) name8624 (
		\DM_rd3[14]_pad ,
		_w7038_,
		_w12671_
	);
	LUT2 #(
		.INIT('h2)
	) name8625 (
		\DM_rd0[14]_pad ,
		_w7053_,
		_w12672_
	);
	LUT2 #(
		.INIT('h8)
	) name8626 (
		\DM_rd5[14]_pad ,
		_w7043_,
		_w12673_
	);
	LUT2 #(
		.INIT('h8)
	) name8627 (
		\DM_rd2[14]_pad ,
		_w7041_,
		_w12674_
	);
	LUT2 #(
		.INIT('h1)
	) name8628 (
		_w12667_,
		_w12671_,
		_w12675_
	);
	LUT2 #(
		.INIT('h4)
	) name8629 (
		_w12674_,
		_w12675_,
		_w12676_
	);
	LUT2 #(
		.INIT('h1)
	) name8630 (
		_w7057_,
		_w12666_,
		_w12677_
	);
	LUT2 #(
		.INIT('h1)
	) name8631 (
		_w12669_,
		_w12670_,
		_w12678_
	);
	LUT2 #(
		.INIT('h8)
	) name8632 (
		_w12677_,
		_w12678_,
		_w12679_
	);
	LUT2 #(
		.INIT('h4)
	) name8633 (
		_w12668_,
		_w12676_,
		_w12680_
	);
	LUT2 #(
		.INIT('h4)
	) name8634 (
		_w12673_,
		_w12680_,
		_w12681_
	);
	LUT2 #(
		.INIT('h8)
	) name8635 (
		_w12679_,
		_w12681_,
		_w12682_
	);
	LUT2 #(
		.INIT('h4)
	) name8636 (
		_w12672_,
		_w12682_,
		_w12683_
	);
	LUT2 #(
		.INIT('h1)
	) name8637 (
		\emc_DMDoe_reg/NET0131 ,
		_w11954_,
		_w12684_
	);
	LUT2 #(
		.INIT('h8)
	) name8638 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[14]/P0001 ,
		_w12685_
	);
	LUT2 #(
		.INIT('h2)
	) name8639 (
		_w7057_,
		_w12685_,
		_w12686_
	);
	LUT2 #(
		.INIT('h4)
	) name8640 (
		_w12684_,
		_w12686_,
		_w12687_
	);
	LUT2 #(
		.INIT('h1)
	) name8641 (
		_w12683_,
		_w12687_,
		_w12688_
	);
	LUT2 #(
		.INIT('h8)
	) name8642 (
		_w12456_,
		_w12688_,
		_w12689_
	);
	LUT2 #(
		.INIT('h8)
	) name8643 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[14]/P0001 ,
		_w12690_
	);
	LUT2 #(
		.INIT('h4)
	) name8644 (
		_w11842_,
		_w12468_,
		_w12691_
	);
	LUT2 #(
		.INIT('h4)
	) name8645 (
		_w11858_,
		_w12466_,
		_w12692_
	);
	LUT2 #(
		.INIT('h4)
	) name8646 (
		_w11889_,
		_w12470_,
		_w12693_
	);
	LUT2 #(
		.INIT('h1)
	) name8647 (
		_w12691_,
		_w12692_,
		_w12694_
	);
	LUT2 #(
		.INIT('h4)
	) name8648 (
		_w12693_,
		_w12694_,
		_w12695_
	);
	LUT2 #(
		.INIT('h1)
	) name8649 (
		\emc_PMDoe_reg/NET0131 ,
		_w12695_,
		_w12696_
	);
	LUT2 #(
		.INIT('h2)
	) name8650 (
		_w12465_,
		_w12690_,
		_w12697_
	);
	LUT2 #(
		.INIT('h4)
	) name8651 (
		_w12696_,
		_w12697_,
		_w12698_
	);
	LUT2 #(
		.INIT('h8)
	) name8652 (
		\PM_rd2[14]_pad ,
		_w12478_,
		_w12699_
	);
	LUT2 #(
		.INIT('h2)
	) name8653 (
		\PM_rd0[14]_pad ,
		_w12504_,
		_w12700_
	);
	LUT2 #(
		.INIT('h8)
	) name8654 (
		\PM_rd4[14]_pad ,
		_w12488_,
		_w12701_
	);
	LUT2 #(
		.INIT('h8)
	) name8655 (
		\PM_rd6[14]_pad ,
		_w12483_,
		_w12702_
	);
	LUT2 #(
		.INIT('h8)
	) name8656 (
		\PM_rd7[14]_pad ,
		_w12485_,
		_w12703_
	);
	LUT2 #(
		.INIT('h8)
	) name8657 (
		\PM_rd3[14]_pad ,
		_w12493_,
		_w12704_
	);
	LUT2 #(
		.INIT('h8)
	) name8658 (
		\PM_rd1[14]_pad ,
		_w12491_,
		_w12705_
	);
	LUT2 #(
		.INIT('h8)
	) name8659 (
		\PM_rd5[14]_pad ,
		_w12495_,
		_w12706_
	);
	LUT2 #(
		.INIT('h1)
	) name8660 (
		_w12465_,
		_w12702_,
		_w12707_
	);
	LUT2 #(
		.INIT('h4)
	) name8661 (
		_w12703_,
		_w12707_,
		_w12708_
	);
	LUT2 #(
		.INIT('h1)
	) name8662 (
		_w12699_,
		_w12701_,
		_w12709_
	);
	LUT2 #(
		.INIT('h1)
	) name8663 (
		_w12704_,
		_w12705_,
		_w12710_
	);
	LUT2 #(
		.INIT('h4)
	) name8664 (
		_w12706_,
		_w12710_,
		_w12711_
	);
	LUT2 #(
		.INIT('h8)
	) name8665 (
		_w12708_,
		_w12709_,
		_w12712_
	);
	LUT2 #(
		.INIT('h8)
	) name8666 (
		_w12711_,
		_w12712_,
		_w12713_
	);
	LUT2 #(
		.INIT('h4)
	) name8667 (
		_w12700_,
		_w12713_,
		_w12714_
	);
	LUT2 #(
		.INIT('h1)
	) name8668 (
		_w12698_,
		_w12714_,
		_w12715_
	);
	LUT2 #(
		.INIT('h8)
	) name8669 (
		_w12452_,
		_w12715_,
		_w12716_
	);
	LUT2 #(
		.INIT('h1)
	) name8670 (
		_w12665_,
		_w12716_,
		_w12717_
	);
	LUT2 #(
		.INIT('h4)
	) name8671 (
		_w12689_,
		_w12717_,
		_w12718_
	);
	LUT2 #(
		.INIT('h2)
	) name8672 (
		_w12451_,
		_w12718_,
		_w12719_
	);
	LUT2 #(
		.INIT('h1)
	) name8673 (
		_w12664_,
		_w12719_,
		_w12720_
	);
	LUT2 #(
		.INIT('h8)
	) name8674 (
		\DM_rdm[15]_pad ,
		_w7016_,
		_w12721_
	);
	LUT2 #(
		.INIT('h8)
	) name8675 (
		\DM_rd1[15]_pad ,
		_w7022_,
		_w12722_
	);
	LUT2 #(
		.INIT('h8)
	) name8676 (
		\DM_rd4[15]_pad ,
		_w7028_,
		_w12723_
	);
	LUT2 #(
		.INIT('h8)
	) name8677 (
		\DM_rd6[15]_pad ,
		_w7031_,
		_w12724_
	);
	LUT2 #(
		.INIT('h8)
	) name8678 (
		\DM_rd7[15]_pad ,
		_w7034_,
		_w12725_
	);
	LUT2 #(
		.INIT('h8)
	) name8679 (
		\DM_rd3[15]_pad ,
		_w7038_,
		_w12726_
	);
	LUT2 #(
		.INIT('h2)
	) name8680 (
		\DM_rd0[15]_pad ,
		_w7053_,
		_w12727_
	);
	LUT2 #(
		.INIT('h8)
	) name8681 (
		\DM_rd5[15]_pad ,
		_w7043_,
		_w12728_
	);
	LUT2 #(
		.INIT('h8)
	) name8682 (
		\DM_rd2[15]_pad ,
		_w7041_,
		_w12729_
	);
	LUT2 #(
		.INIT('h1)
	) name8683 (
		_w12722_,
		_w12726_,
		_w12730_
	);
	LUT2 #(
		.INIT('h4)
	) name8684 (
		_w12729_,
		_w12730_,
		_w12731_
	);
	LUT2 #(
		.INIT('h1)
	) name8685 (
		_w7057_,
		_w12721_,
		_w12732_
	);
	LUT2 #(
		.INIT('h1)
	) name8686 (
		_w12724_,
		_w12725_,
		_w12733_
	);
	LUT2 #(
		.INIT('h8)
	) name8687 (
		_w12732_,
		_w12733_,
		_w12734_
	);
	LUT2 #(
		.INIT('h4)
	) name8688 (
		_w12723_,
		_w12731_,
		_w12735_
	);
	LUT2 #(
		.INIT('h4)
	) name8689 (
		_w12728_,
		_w12735_,
		_w12736_
	);
	LUT2 #(
		.INIT('h8)
	) name8690 (
		_w12734_,
		_w12736_,
		_w12737_
	);
	LUT2 #(
		.INIT('h4)
	) name8691 (
		_w12727_,
		_w12737_,
		_w12738_
	);
	LUT2 #(
		.INIT('h1)
	) name8692 (
		\emc_DMDoe_reg/NET0131 ,
		_w12096_,
		_w12739_
	);
	LUT2 #(
		.INIT('h8)
	) name8693 (
		\emc_DMDoe_reg/NET0131 ,
		\emc_DMDreg_reg[15]/P0001 ,
		_w12740_
	);
	LUT2 #(
		.INIT('h2)
	) name8694 (
		_w7057_,
		_w12740_,
		_w12741_
	);
	LUT2 #(
		.INIT('h4)
	) name8695 (
		_w12739_,
		_w12741_,
		_w12742_
	);
	LUT2 #(
		.INIT('h1)
	) name8696 (
		_w12738_,
		_w12742_,
		_w12743_
	);
	LUT2 #(
		.INIT('h8)
	) name8697 (
		_w12456_,
		_w12743_,
		_w12744_
	);
	LUT2 #(
		.INIT('h8)
	) name8698 (
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w12454_,
		_w12745_
	);
	LUT2 #(
		.INIT('h8)
	) name8699 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[15]/P0001 ,
		_w12746_
	);
	LUT2 #(
		.INIT('h4)
	) name8700 (
		_w11988_,
		_w12468_,
		_w12747_
	);
	LUT2 #(
		.INIT('h4)
	) name8701 (
		_w12004_,
		_w12466_,
		_w12748_
	);
	LUT2 #(
		.INIT('h4)
	) name8702 (
		_w12035_,
		_w12470_,
		_w12749_
	);
	LUT2 #(
		.INIT('h1)
	) name8703 (
		_w12747_,
		_w12748_,
		_w12750_
	);
	LUT2 #(
		.INIT('h4)
	) name8704 (
		_w12749_,
		_w12750_,
		_w12751_
	);
	LUT2 #(
		.INIT('h1)
	) name8705 (
		\emc_PMDoe_reg/NET0131 ,
		_w12751_,
		_w12752_
	);
	LUT2 #(
		.INIT('h2)
	) name8706 (
		_w12465_,
		_w12746_,
		_w12753_
	);
	LUT2 #(
		.INIT('h4)
	) name8707 (
		_w12752_,
		_w12753_,
		_w12754_
	);
	LUT2 #(
		.INIT('h8)
	) name8708 (
		\PM_rd2[15]_pad ,
		_w12478_,
		_w12755_
	);
	LUT2 #(
		.INIT('h2)
	) name8709 (
		\PM_rd0[15]_pad ,
		_w12504_,
		_w12756_
	);
	LUT2 #(
		.INIT('h8)
	) name8710 (
		\PM_rd4[15]_pad ,
		_w12488_,
		_w12757_
	);
	LUT2 #(
		.INIT('h8)
	) name8711 (
		\PM_rd6[15]_pad ,
		_w12483_,
		_w12758_
	);
	LUT2 #(
		.INIT('h8)
	) name8712 (
		\PM_rd7[15]_pad ,
		_w12485_,
		_w12759_
	);
	LUT2 #(
		.INIT('h8)
	) name8713 (
		\PM_rd3[15]_pad ,
		_w12493_,
		_w12760_
	);
	LUT2 #(
		.INIT('h8)
	) name8714 (
		\PM_rd1[15]_pad ,
		_w12491_,
		_w12761_
	);
	LUT2 #(
		.INIT('h8)
	) name8715 (
		\PM_rd5[15]_pad ,
		_w12495_,
		_w12762_
	);
	LUT2 #(
		.INIT('h1)
	) name8716 (
		_w12465_,
		_w12758_,
		_w12763_
	);
	LUT2 #(
		.INIT('h4)
	) name8717 (
		_w12759_,
		_w12763_,
		_w12764_
	);
	LUT2 #(
		.INIT('h1)
	) name8718 (
		_w12755_,
		_w12757_,
		_w12765_
	);
	LUT2 #(
		.INIT('h1)
	) name8719 (
		_w12760_,
		_w12761_,
		_w12766_
	);
	LUT2 #(
		.INIT('h4)
	) name8720 (
		_w12762_,
		_w12766_,
		_w12767_
	);
	LUT2 #(
		.INIT('h8)
	) name8721 (
		_w12764_,
		_w12765_,
		_w12768_
	);
	LUT2 #(
		.INIT('h8)
	) name8722 (
		_w12767_,
		_w12768_,
		_w12769_
	);
	LUT2 #(
		.INIT('h4)
	) name8723 (
		_w12756_,
		_w12769_,
		_w12770_
	);
	LUT2 #(
		.INIT('h1)
	) name8724 (
		_w12754_,
		_w12770_,
		_w12771_
	);
	LUT2 #(
		.INIT('h8)
	) name8725 (
		_w12452_,
		_w12771_,
		_w12772_
	);
	LUT2 #(
		.INIT('h1)
	) name8726 (
		_w12744_,
		_w12772_,
		_w12773_
	);
	LUT2 #(
		.INIT('h4)
	) name8727 (
		_w12745_,
		_w12773_,
		_w12774_
	);
	LUT2 #(
		.INIT('h8)
	) name8728 (
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w12454_,
		_w12775_
	);
	LUT2 #(
		.INIT('h8)
	) name8729 (
		_w9435_,
		_w12456_,
		_w12776_
	);
	LUT2 #(
		.INIT('h8)
	) name8730 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[1]/P0001 ,
		_w12777_
	);
	LUT2 #(
		.INIT('h4)
	) name8731 (
		_w9285_,
		_w12466_,
		_w12778_
	);
	LUT2 #(
		.INIT('h4)
	) name8732 (
		_w9320_,
		_w12468_,
		_w12779_
	);
	LUT2 #(
		.INIT('h4)
	) name8733 (
		_w9236_,
		_w12470_,
		_w12780_
	);
	LUT2 #(
		.INIT('h1)
	) name8734 (
		_w12778_,
		_w12779_,
		_w12781_
	);
	LUT2 #(
		.INIT('h4)
	) name8735 (
		_w12780_,
		_w12781_,
		_w12782_
	);
	LUT2 #(
		.INIT('h1)
	) name8736 (
		\emc_PMDoe_reg/NET0131 ,
		_w12782_,
		_w12783_
	);
	LUT2 #(
		.INIT('h2)
	) name8737 (
		_w12465_,
		_w12777_,
		_w12784_
	);
	LUT2 #(
		.INIT('h4)
	) name8738 (
		_w12783_,
		_w12784_,
		_w12785_
	);
	LUT2 #(
		.INIT('h8)
	) name8739 (
		\PM_rd2[1]_pad ,
		_w12478_,
		_w12786_
	);
	LUT2 #(
		.INIT('h2)
	) name8740 (
		\PM_rd0[1]_pad ,
		_w12504_,
		_w12787_
	);
	LUT2 #(
		.INIT('h8)
	) name8741 (
		\PM_rd4[1]_pad ,
		_w12488_,
		_w12788_
	);
	LUT2 #(
		.INIT('h8)
	) name8742 (
		\PM_rd6[1]_pad ,
		_w12483_,
		_w12789_
	);
	LUT2 #(
		.INIT('h8)
	) name8743 (
		\PM_rd7[1]_pad ,
		_w12485_,
		_w12790_
	);
	LUT2 #(
		.INIT('h8)
	) name8744 (
		\PM_rd3[1]_pad ,
		_w12493_,
		_w12791_
	);
	LUT2 #(
		.INIT('h8)
	) name8745 (
		\PM_rd1[1]_pad ,
		_w12491_,
		_w12792_
	);
	LUT2 #(
		.INIT('h8)
	) name8746 (
		\PM_rd5[1]_pad ,
		_w12495_,
		_w12793_
	);
	LUT2 #(
		.INIT('h1)
	) name8747 (
		_w12465_,
		_w12789_,
		_w12794_
	);
	LUT2 #(
		.INIT('h4)
	) name8748 (
		_w12790_,
		_w12794_,
		_w12795_
	);
	LUT2 #(
		.INIT('h1)
	) name8749 (
		_w12786_,
		_w12788_,
		_w12796_
	);
	LUT2 #(
		.INIT('h1)
	) name8750 (
		_w12791_,
		_w12792_,
		_w12797_
	);
	LUT2 #(
		.INIT('h4)
	) name8751 (
		_w12793_,
		_w12797_,
		_w12798_
	);
	LUT2 #(
		.INIT('h8)
	) name8752 (
		_w12795_,
		_w12796_,
		_w12799_
	);
	LUT2 #(
		.INIT('h8)
	) name8753 (
		_w12798_,
		_w12799_,
		_w12800_
	);
	LUT2 #(
		.INIT('h4)
	) name8754 (
		_w12787_,
		_w12800_,
		_w12801_
	);
	LUT2 #(
		.INIT('h1)
	) name8755 (
		_w12785_,
		_w12801_,
		_w12802_
	);
	LUT2 #(
		.INIT('h8)
	) name8756 (
		_w12452_,
		_w12802_,
		_w12803_
	);
	LUT2 #(
		.INIT('h1)
	) name8757 (
		_w12775_,
		_w12803_,
		_w12804_
	);
	LUT2 #(
		.INIT('h4)
	) name8758 (
		_w12776_,
		_w12804_,
		_w12805_
	);
	LUT2 #(
		.INIT('h2)
	) name8759 (
		_w12451_,
		_w12805_,
		_w12806_
	);
	LUT2 #(
		.INIT('h8)
	) name8760 (
		\bdma_BWdataBUF_reg[1]/P0001 ,
		_w12525_,
		_w12807_
	);
	LUT2 #(
		.INIT('h1)
	) name8761 (
		_w12806_,
		_w12807_,
		_w12808_
	);
	LUT2 #(
		.INIT('h8)
	) name8762 (
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w12454_,
		_w12809_
	);
	LUT2 #(
		.INIT('h8)
	) name8763 (
		_w8715_,
		_w12456_,
		_w12810_
	);
	LUT2 #(
		.INIT('h8)
	) name8764 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[2]/P0001 ,
		_w12811_
	);
	LUT2 #(
		.INIT('h4)
	) name8765 (
		_w8565_,
		_w12470_,
		_w12812_
	);
	LUT2 #(
		.INIT('h4)
	) name8766 (
		_w8600_,
		_w12468_,
		_w12813_
	);
	LUT2 #(
		.INIT('h4)
	) name8767 (
		_w8506_,
		_w12466_,
		_w12814_
	);
	LUT2 #(
		.INIT('h1)
	) name8768 (
		_w12812_,
		_w12813_,
		_w12815_
	);
	LUT2 #(
		.INIT('h4)
	) name8769 (
		_w12814_,
		_w12815_,
		_w12816_
	);
	LUT2 #(
		.INIT('h1)
	) name8770 (
		\emc_PMDoe_reg/NET0131 ,
		_w12816_,
		_w12817_
	);
	LUT2 #(
		.INIT('h2)
	) name8771 (
		_w12465_,
		_w12811_,
		_w12818_
	);
	LUT2 #(
		.INIT('h4)
	) name8772 (
		_w12817_,
		_w12818_,
		_w12819_
	);
	LUT2 #(
		.INIT('h8)
	) name8773 (
		\PM_rd2[2]_pad ,
		_w12478_,
		_w12820_
	);
	LUT2 #(
		.INIT('h2)
	) name8774 (
		\PM_rd0[2]_pad ,
		_w12504_,
		_w12821_
	);
	LUT2 #(
		.INIT('h8)
	) name8775 (
		\PM_rd4[2]_pad ,
		_w12488_,
		_w12822_
	);
	LUT2 #(
		.INIT('h8)
	) name8776 (
		\PM_rd6[2]_pad ,
		_w12483_,
		_w12823_
	);
	LUT2 #(
		.INIT('h8)
	) name8777 (
		\PM_rd7[2]_pad ,
		_w12485_,
		_w12824_
	);
	LUT2 #(
		.INIT('h8)
	) name8778 (
		\PM_rd3[2]_pad ,
		_w12493_,
		_w12825_
	);
	LUT2 #(
		.INIT('h8)
	) name8779 (
		\PM_rd1[2]_pad ,
		_w12491_,
		_w12826_
	);
	LUT2 #(
		.INIT('h8)
	) name8780 (
		\PM_rd5[2]_pad ,
		_w12495_,
		_w12827_
	);
	LUT2 #(
		.INIT('h1)
	) name8781 (
		_w12465_,
		_w12823_,
		_w12828_
	);
	LUT2 #(
		.INIT('h4)
	) name8782 (
		_w12824_,
		_w12828_,
		_w12829_
	);
	LUT2 #(
		.INIT('h1)
	) name8783 (
		_w12820_,
		_w12822_,
		_w12830_
	);
	LUT2 #(
		.INIT('h1)
	) name8784 (
		_w12825_,
		_w12826_,
		_w12831_
	);
	LUT2 #(
		.INIT('h4)
	) name8785 (
		_w12827_,
		_w12831_,
		_w12832_
	);
	LUT2 #(
		.INIT('h8)
	) name8786 (
		_w12829_,
		_w12830_,
		_w12833_
	);
	LUT2 #(
		.INIT('h8)
	) name8787 (
		_w12832_,
		_w12833_,
		_w12834_
	);
	LUT2 #(
		.INIT('h4)
	) name8788 (
		_w12821_,
		_w12834_,
		_w12835_
	);
	LUT2 #(
		.INIT('h1)
	) name8789 (
		_w12819_,
		_w12835_,
		_w12836_
	);
	LUT2 #(
		.INIT('h8)
	) name8790 (
		_w12452_,
		_w12836_,
		_w12837_
	);
	LUT2 #(
		.INIT('h1)
	) name8791 (
		_w12809_,
		_w12837_,
		_w12838_
	);
	LUT2 #(
		.INIT('h4)
	) name8792 (
		_w12810_,
		_w12838_,
		_w12839_
	);
	LUT2 #(
		.INIT('h2)
	) name8793 (
		_w12451_,
		_w12839_,
		_w12840_
	);
	LUT2 #(
		.INIT('h8)
	) name8794 (
		\bdma_BWdataBUF_reg[2]/P0001 ,
		_w12525_,
		_w12841_
	);
	LUT2 #(
		.INIT('h1)
	) name8795 (
		_w12840_,
		_w12841_,
		_w12842_
	);
	LUT2 #(
		.INIT('h8)
	) name8796 (
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w12454_,
		_w12843_
	);
	LUT2 #(
		.INIT('h8)
	) name8797 (
		_w8113_,
		_w12456_,
		_w12844_
	);
	LUT2 #(
		.INIT('h8)
	) name8798 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[3]/P0001 ,
		_w12845_
	);
	LUT2 #(
		.INIT('h4)
	) name8799 (
		_w8000_,
		_w12466_,
		_w12846_
	);
	LUT2 #(
		.INIT('h4)
	) name8800 (
		_w7967_,
		_w12468_,
		_w12847_
	);
	LUT2 #(
		.INIT('h4)
	) name8801 (
		_w7916_,
		_w12470_,
		_w12848_
	);
	LUT2 #(
		.INIT('h1)
	) name8802 (
		_w12846_,
		_w12847_,
		_w12849_
	);
	LUT2 #(
		.INIT('h4)
	) name8803 (
		_w12848_,
		_w12849_,
		_w12850_
	);
	LUT2 #(
		.INIT('h1)
	) name8804 (
		\emc_PMDoe_reg/NET0131 ,
		_w12850_,
		_w12851_
	);
	LUT2 #(
		.INIT('h2)
	) name8805 (
		_w12465_,
		_w12845_,
		_w12852_
	);
	LUT2 #(
		.INIT('h4)
	) name8806 (
		_w12851_,
		_w12852_,
		_w12853_
	);
	LUT2 #(
		.INIT('h8)
	) name8807 (
		\PM_rd2[3]_pad ,
		_w12478_,
		_w12854_
	);
	LUT2 #(
		.INIT('h2)
	) name8808 (
		\PM_rd0[3]_pad ,
		_w12504_,
		_w12855_
	);
	LUT2 #(
		.INIT('h8)
	) name8809 (
		\PM_rd4[3]_pad ,
		_w12488_,
		_w12856_
	);
	LUT2 #(
		.INIT('h8)
	) name8810 (
		\PM_rd6[3]_pad ,
		_w12483_,
		_w12857_
	);
	LUT2 #(
		.INIT('h8)
	) name8811 (
		\PM_rd7[3]_pad ,
		_w12485_,
		_w12858_
	);
	LUT2 #(
		.INIT('h8)
	) name8812 (
		\PM_rd3[3]_pad ,
		_w12493_,
		_w12859_
	);
	LUT2 #(
		.INIT('h8)
	) name8813 (
		\PM_rd1[3]_pad ,
		_w12491_,
		_w12860_
	);
	LUT2 #(
		.INIT('h8)
	) name8814 (
		\PM_rd5[3]_pad ,
		_w12495_,
		_w12861_
	);
	LUT2 #(
		.INIT('h1)
	) name8815 (
		_w12465_,
		_w12857_,
		_w12862_
	);
	LUT2 #(
		.INIT('h4)
	) name8816 (
		_w12858_,
		_w12862_,
		_w12863_
	);
	LUT2 #(
		.INIT('h1)
	) name8817 (
		_w12854_,
		_w12856_,
		_w12864_
	);
	LUT2 #(
		.INIT('h1)
	) name8818 (
		_w12859_,
		_w12860_,
		_w12865_
	);
	LUT2 #(
		.INIT('h4)
	) name8819 (
		_w12861_,
		_w12865_,
		_w12866_
	);
	LUT2 #(
		.INIT('h8)
	) name8820 (
		_w12863_,
		_w12864_,
		_w12867_
	);
	LUT2 #(
		.INIT('h8)
	) name8821 (
		_w12866_,
		_w12867_,
		_w12868_
	);
	LUT2 #(
		.INIT('h4)
	) name8822 (
		_w12855_,
		_w12868_,
		_w12869_
	);
	LUT2 #(
		.INIT('h1)
	) name8823 (
		_w12853_,
		_w12869_,
		_w12870_
	);
	LUT2 #(
		.INIT('h8)
	) name8824 (
		_w12452_,
		_w12870_,
		_w12871_
	);
	LUT2 #(
		.INIT('h1)
	) name8825 (
		_w12843_,
		_w12871_,
		_w12872_
	);
	LUT2 #(
		.INIT('h4)
	) name8826 (
		_w12844_,
		_w12872_,
		_w12873_
	);
	LUT2 #(
		.INIT('h2)
	) name8827 (
		_w12451_,
		_w12873_,
		_w12874_
	);
	LUT2 #(
		.INIT('h8)
	) name8828 (
		\bdma_BWdataBUF_reg[3]/P0001 ,
		_w12525_,
		_w12875_
	);
	LUT2 #(
		.INIT('h1)
	) name8829 (
		_w12874_,
		_w12875_,
		_w12876_
	);
	LUT2 #(
		.INIT('h8)
	) name8830 (
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w12454_,
		_w12877_
	);
	LUT2 #(
		.INIT('h8)
	) name8831 (
		_w10069_,
		_w12456_,
		_w12878_
	);
	LUT2 #(
		.INIT('h8)
	) name8832 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[4]/P0001 ,
		_w12879_
	);
	LUT2 #(
		.INIT('h4)
	) name8833 (
		_w9927_,
		_w12468_,
		_w12880_
	);
	LUT2 #(
		.INIT('h4)
	) name8834 (
		_w9956_,
		_w12466_,
		_w12881_
	);
	LUT2 #(
		.INIT('h4)
	) name8835 (
		_w9876_,
		_w12470_,
		_w12882_
	);
	LUT2 #(
		.INIT('h1)
	) name8836 (
		_w12880_,
		_w12881_,
		_w12883_
	);
	LUT2 #(
		.INIT('h4)
	) name8837 (
		_w12882_,
		_w12883_,
		_w12884_
	);
	LUT2 #(
		.INIT('h1)
	) name8838 (
		\emc_PMDoe_reg/NET0131 ,
		_w12884_,
		_w12885_
	);
	LUT2 #(
		.INIT('h2)
	) name8839 (
		_w12465_,
		_w12879_,
		_w12886_
	);
	LUT2 #(
		.INIT('h4)
	) name8840 (
		_w12885_,
		_w12886_,
		_w12887_
	);
	LUT2 #(
		.INIT('h8)
	) name8841 (
		\PM_rd2[4]_pad ,
		_w12478_,
		_w12888_
	);
	LUT2 #(
		.INIT('h2)
	) name8842 (
		\PM_rd0[4]_pad ,
		_w12504_,
		_w12889_
	);
	LUT2 #(
		.INIT('h8)
	) name8843 (
		\PM_rd4[4]_pad ,
		_w12488_,
		_w12890_
	);
	LUT2 #(
		.INIT('h8)
	) name8844 (
		\PM_rd6[4]_pad ,
		_w12483_,
		_w12891_
	);
	LUT2 #(
		.INIT('h8)
	) name8845 (
		\PM_rd7[4]_pad ,
		_w12485_,
		_w12892_
	);
	LUT2 #(
		.INIT('h8)
	) name8846 (
		\PM_rd3[4]_pad ,
		_w12493_,
		_w12893_
	);
	LUT2 #(
		.INIT('h8)
	) name8847 (
		\PM_rd1[4]_pad ,
		_w12491_,
		_w12894_
	);
	LUT2 #(
		.INIT('h8)
	) name8848 (
		\PM_rd5[4]_pad ,
		_w12495_,
		_w12895_
	);
	LUT2 #(
		.INIT('h1)
	) name8849 (
		_w12465_,
		_w12891_,
		_w12896_
	);
	LUT2 #(
		.INIT('h4)
	) name8850 (
		_w12892_,
		_w12896_,
		_w12897_
	);
	LUT2 #(
		.INIT('h1)
	) name8851 (
		_w12888_,
		_w12890_,
		_w12898_
	);
	LUT2 #(
		.INIT('h1)
	) name8852 (
		_w12893_,
		_w12894_,
		_w12899_
	);
	LUT2 #(
		.INIT('h4)
	) name8853 (
		_w12895_,
		_w12899_,
		_w12900_
	);
	LUT2 #(
		.INIT('h8)
	) name8854 (
		_w12897_,
		_w12898_,
		_w12901_
	);
	LUT2 #(
		.INIT('h8)
	) name8855 (
		_w12900_,
		_w12901_,
		_w12902_
	);
	LUT2 #(
		.INIT('h4)
	) name8856 (
		_w12889_,
		_w12902_,
		_w12903_
	);
	LUT2 #(
		.INIT('h1)
	) name8857 (
		_w12887_,
		_w12903_,
		_w12904_
	);
	LUT2 #(
		.INIT('h8)
	) name8858 (
		_w12452_,
		_w12904_,
		_w12905_
	);
	LUT2 #(
		.INIT('h1)
	) name8859 (
		_w12877_,
		_w12905_,
		_w12906_
	);
	LUT2 #(
		.INIT('h4)
	) name8860 (
		_w12878_,
		_w12906_,
		_w12907_
	);
	LUT2 #(
		.INIT('h2)
	) name8861 (
		_w12451_,
		_w12907_,
		_w12908_
	);
	LUT2 #(
		.INIT('h8)
	) name8862 (
		\bdma_BWdataBUF_reg[4]/P0001 ,
		_w12525_,
		_w12909_
	);
	LUT2 #(
		.INIT('h1)
	) name8863 (
		_w12908_,
		_w12909_,
		_w12910_
	);
	LUT2 #(
		.INIT('h8)
	) name8864 (
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w12454_,
		_w12911_
	);
	LUT2 #(
		.INIT('h8)
	) name8865 (
		_w10911_,
		_w12456_,
		_w12912_
	);
	LUT2 #(
		.INIT('h8)
	) name8866 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[5]/P0001 ,
		_w12913_
	);
	LUT2 #(
		.INIT('h4)
	) name8867 (
		_w10709_,
		_w12468_,
		_w12914_
	);
	LUT2 #(
		.INIT('h4)
	) name8868 (
		_w10806_,
		_w12466_,
		_w12915_
	);
	LUT2 #(
		.INIT('h4)
	) name8869 (
		_w10889_,
		_w12470_,
		_w12916_
	);
	LUT2 #(
		.INIT('h1)
	) name8870 (
		_w12914_,
		_w12915_,
		_w12917_
	);
	LUT2 #(
		.INIT('h4)
	) name8871 (
		_w12916_,
		_w12917_,
		_w12918_
	);
	LUT2 #(
		.INIT('h1)
	) name8872 (
		\emc_PMDoe_reg/NET0131 ,
		_w12918_,
		_w12919_
	);
	LUT2 #(
		.INIT('h2)
	) name8873 (
		_w12465_,
		_w12913_,
		_w12920_
	);
	LUT2 #(
		.INIT('h4)
	) name8874 (
		_w12919_,
		_w12920_,
		_w12921_
	);
	LUT2 #(
		.INIT('h8)
	) name8875 (
		\PM_rd2[5]_pad ,
		_w12478_,
		_w12922_
	);
	LUT2 #(
		.INIT('h2)
	) name8876 (
		\PM_rd0[5]_pad ,
		_w12504_,
		_w12923_
	);
	LUT2 #(
		.INIT('h8)
	) name8877 (
		\PM_rd4[5]_pad ,
		_w12488_,
		_w12924_
	);
	LUT2 #(
		.INIT('h8)
	) name8878 (
		\PM_rd6[5]_pad ,
		_w12483_,
		_w12925_
	);
	LUT2 #(
		.INIT('h8)
	) name8879 (
		\PM_rd7[5]_pad ,
		_w12485_,
		_w12926_
	);
	LUT2 #(
		.INIT('h8)
	) name8880 (
		\PM_rd3[5]_pad ,
		_w12493_,
		_w12927_
	);
	LUT2 #(
		.INIT('h8)
	) name8881 (
		\PM_rd1[5]_pad ,
		_w12491_,
		_w12928_
	);
	LUT2 #(
		.INIT('h8)
	) name8882 (
		\PM_rd5[5]_pad ,
		_w12495_,
		_w12929_
	);
	LUT2 #(
		.INIT('h1)
	) name8883 (
		_w12465_,
		_w12925_,
		_w12930_
	);
	LUT2 #(
		.INIT('h4)
	) name8884 (
		_w12926_,
		_w12930_,
		_w12931_
	);
	LUT2 #(
		.INIT('h1)
	) name8885 (
		_w12922_,
		_w12924_,
		_w12932_
	);
	LUT2 #(
		.INIT('h1)
	) name8886 (
		_w12927_,
		_w12928_,
		_w12933_
	);
	LUT2 #(
		.INIT('h4)
	) name8887 (
		_w12929_,
		_w12933_,
		_w12934_
	);
	LUT2 #(
		.INIT('h8)
	) name8888 (
		_w12931_,
		_w12932_,
		_w12935_
	);
	LUT2 #(
		.INIT('h8)
	) name8889 (
		_w12934_,
		_w12935_,
		_w12936_
	);
	LUT2 #(
		.INIT('h4)
	) name8890 (
		_w12923_,
		_w12936_,
		_w12937_
	);
	LUT2 #(
		.INIT('h1)
	) name8891 (
		_w12921_,
		_w12937_,
		_w12938_
	);
	LUT2 #(
		.INIT('h8)
	) name8892 (
		_w12452_,
		_w12938_,
		_w12939_
	);
	LUT2 #(
		.INIT('h1)
	) name8893 (
		_w12911_,
		_w12939_,
		_w12940_
	);
	LUT2 #(
		.INIT('h4)
	) name8894 (
		_w12912_,
		_w12940_,
		_w12941_
	);
	LUT2 #(
		.INIT('h2)
	) name8895 (
		_w12451_,
		_w12941_,
		_w12942_
	);
	LUT2 #(
		.INIT('h8)
	) name8896 (
		\bdma_BWdataBUF_reg[5]/P0001 ,
		_w12525_,
		_w12943_
	);
	LUT2 #(
		.INIT('h1)
	) name8897 (
		_w12942_,
		_w12943_,
		_w12944_
	);
	LUT2 #(
		.INIT('h8)
	) name8898 (
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w12454_,
		_w12945_
	);
	LUT2 #(
		.INIT('h8)
	) name8899 (
		_w11525_,
		_w12456_,
		_w12946_
	);
	LUT2 #(
		.INIT('h8)
	) name8900 (
		\PM_rd6[6]_pad ,
		_w12483_,
		_w12947_
	);
	LUT2 #(
		.INIT('h8)
	) name8901 (
		\PM_rd3[6]_pad ,
		_w12493_,
		_w12948_
	);
	LUT2 #(
		.INIT('h2)
	) name8902 (
		\PM_rd0[6]_pad ,
		_w12504_,
		_w12949_
	);
	LUT2 #(
		.INIT('h8)
	) name8903 (
		\PM_rd4[6]_pad ,
		_w12488_,
		_w12950_
	);
	LUT2 #(
		.INIT('h8)
	) name8904 (
		\PM_rd5[6]_pad ,
		_w12495_,
		_w12951_
	);
	LUT2 #(
		.INIT('h8)
	) name8905 (
		\PM_rd7[6]_pad ,
		_w12485_,
		_w12952_
	);
	LUT2 #(
		.INIT('h8)
	) name8906 (
		\PM_rd2[6]_pad ,
		_w12478_,
		_w12953_
	);
	LUT2 #(
		.INIT('h8)
	) name8907 (
		\PM_rd1[6]_pad ,
		_w12491_,
		_w12954_
	);
	LUT2 #(
		.INIT('h1)
	) name8908 (
		_w12465_,
		_w12947_,
		_w12955_
	);
	LUT2 #(
		.INIT('h4)
	) name8909 (
		_w12952_,
		_w12955_,
		_w12956_
	);
	LUT2 #(
		.INIT('h1)
	) name8910 (
		_w12948_,
		_w12950_,
		_w12957_
	);
	LUT2 #(
		.INIT('h1)
	) name8911 (
		_w12951_,
		_w12953_,
		_w12958_
	);
	LUT2 #(
		.INIT('h4)
	) name8912 (
		_w12954_,
		_w12958_,
		_w12959_
	);
	LUT2 #(
		.INIT('h8)
	) name8913 (
		_w12956_,
		_w12957_,
		_w12960_
	);
	LUT2 #(
		.INIT('h8)
	) name8914 (
		_w12959_,
		_w12960_,
		_w12961_
	);
	LUT2 #(
		.INIT('h4)
	) name8915 (
		_w12949_,
		_w12961_,
		_w12962_
	);
	LUT2 #(
		.INIT('h8)
	) name8916 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[6]/P0001 ,
		_w12963_
	);
	LUT2 #(
		.INIT('h4)
	) name8917 (
		_w11455_,
		_w12470_,
		_w12964_
	);
	LUT2 #(
		.INIT('h4)
	) name8918 (
		_w11347_,
		_w12468_,
		_w12965_
	);
	LUT2 #(
		.INIT('h4)
	) name8919 (
		_w11320_,
		_w12466_,
		_w12966_
	);
	LUT2 #(
		.INIT('h1)
	) name8920 (
		_w12964_,
		_w12966_,
		_w12967_
	);
	LUT2 #(
		.INIT('h4)
	) name8921 (
		_w12965_,
		_w12967_,
		_w12968_
	);
	LUT2 #(
		.INIT('h1)
	) name8922 (
		\emc_PMDoe_reg/NET0131 ,
		_w12968_,
		_w12969_
	);
	LUT2 #(
		.INIT('h2)
	) name8923 (
		_w12465_,
		_w12963_,
		_w12970_
	);
	LUT2 #(
		.INIT('h4)
	) name8924 (
		_w12969_,
		_w12970_,
		_w12971_
	);
	LUT2 #(
		.INIT('h1)
	) name8925 (
		_w12962_,
		_w12971_,
		_w12972_
	);
	LUT2 #(
		.INIT('h8)
	) name8926 (
		_w12452_,
		_w12972_,
		_w12973_
	);
	LUT2 #(
		.INIT('h1)
	) name8927 (
		_w12945_,
		_w12973_,
		_w12974_
	);
	LUT2 #(
		.INIT('h4)
	) name8928 (
		_w12946_,
		_w12974_,
		_w12975_
	);
	LUT2 #(
		.INIT('h2)
	) name8929 (
		_w12451_,
		_w12975_,
		_w12976_
	);
	LUT2 #(
		.INIT('h8)
	) name8930 (
		\bdma_BWdataBUF_reg[6]/P0001 ,
		_w12525_,
		_w12977_
	);
	LUT2 #(
		.INIT('h1)
	) name8931 (
		_w12976_,
		_w12977_,
		_w12978_
	);
	LUT2 #(
		.INIT('h8)
	) name8932 (
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w12454_,
		_w12979_
	);
	LUT2 #(
		.INIT('h8)
	) name8933 (
		_w11265_,
		_w12456_,
		_w12980_
	);
	LUT2 #(
		.INIT('h8)
	) name8934 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[7]/P0001 ,
		_w12981_
	);
	LUT2 #(
		.INIT('h4)
	) name8935 (
		_w11077_,
		_w12468_,
		_w12982_
	);
	LUT2 #(
		.INIT('h4)
	) name8936 (
		_w11243_,
		_w12466_,
		_w12983_
	);
	LUT2 #(
		.INIT('h4)
	) name8937 (
		_w11203_,
		_w12470_,
		_w12984_
	);
	LUT2 #(
		.INIT('h1)
	) name8938 (
		_w12982_,
		_w12983_,
		_w12985_
	);
	LUT2 #(
		.INIT('h4)
	) name8939 (
		_w12984_,
		_w12985_,
		_w12986_
	);
	LUT2 #(
		.INIT('h1)
	) name8940 (
		\emc_PMDoe_reg/NET0131 ,
		_w12986_,
		_w12987_
	);
	LUT2 #(
		.INIT('h2)
	) name8941 (
		_w12465_,
		_w12981_,
		_w12988_
	);
	LUT2 #(
		.INIT('h4)
	) name8942 (
		_w12987_,
		_w12988_,
		_w12989_
	);
	LUT2 #(
		.INIT('h8)
	) name8943 (
		\PM_rd2[7]_pad ,
		_w12478_,
		_w12990_
	);
	LUT2 #(
		.INIT('h2)
	) name8944 (
		\PM_rd0[7]_pad ,
		_w12504_,
		_w12991_
	);
	LUT2 #(
		.INIT('h8)
	) name8945 (
		\PM_rd4[7]_pad ,
		_w12488_,
		_w12992_
	);
	LUT2 #(
		.INIT('h8)
	) name8946 (
		\PM_rd6[7]_pad ,
		_w12483_,
		_w12993_
	);
	LUT2 #(
		.INIT('h8)
	) name8947 (
		\PM_rd7[7]_pad ,
		_w12485_,
		_w12994_
	);
	LUT2 #(
		.INIT('h8)
	) name8948 (
		\PM_rd3[7]_pad ,
		_w12493_,
		_w12995_
	);
	LUT2 #(
		.INIT('h8)
	) name8949 (
		\PM_rd1[7]_pad ,
		_w12491_,
		_w12996_
	);
	LUT2 #(
		.INIT('h8)
	) name8950 (
		\PM_rd5[7]_pad ,
		_w12495_,
		_w12997_
	);
	LUT2 #(
		.INIT('h1)
	) name8951 (
		_w12465_,
		_w12993_,
		_w12998_
	);
	LUT2 #(
		.INIT('h4)
	) name8952 (
		_w12994_,
		_w12998_,
		_w12999_
	);
	LUT2 #(
		.INIT('h1)
	) name8953 (
		_w12990_,
		_w12992_,
		_w13000_
	);
	LUT2 #(
		.INIT('h1)
	) name8954 (
		_w12995_,
		_w12996_,
		_w13001_
	);
	LUT2 #(
		.INIT('h4)
	) name8955 (
		_w12997_,
		_w13001_,
		_w13002_
	);
	LUT2 #(
		.INIT('h8)
	) name8956 (
		_w12999_,
		_w13000_,
		_w13003_
	);
	LUT2 #(
		.INIT('h8)
	) name8957 (
		_w13002_,
		_w13003_,
		_w13004_
	);
	LUT2 #(
		.INIT('h4)
	) name8958 (
		_w12991_,
		_w13004_,
		_w13005_
	);
	LUT2 #(
		.INIT('h1)
	) name8959 (
		_w12989_,
		_w13005_,
		_w13006_
	);
	LUT2 #(
		.INIT('h8)
	) name8960 (
		_w12452_,
		_w13006_,
		_w13007_
	);
	LUT2 #(
		.INIT('h1)
	) name8961 (
		_w12979_,
		_w13007_,
		_w13008_
	);
	LUT2 #(
		.INIT('h4)
	) name8962 (
		_w12980_,
		_w13008_,
		_w13009_
	);
	LUT2 #(
		.INIT('h2)
	) name8963 (
		_w12451_,
		_w13009_,
		_w13010_
	);
	LUT2 #(
		.INIT('h8)
	) name8964 (
		\bdma_BWdataBUF_reg[7]/P0001 ,
		_w12525_,
		_w13011_
	);
	LUT2 #(
		.INIT('h1)
	) name8965 (
		_w13010_,
		_w13011_,
		_w13012_
	);
	LUT2 #(
		.INIT('h8)
	) name8966 (
		\bdma_BCTL_reg[9]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w13013_
	);
	LUT2 #(
		.INIT('h8)
	) name8967 (
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w12454_,
		_w13014_
	);
	LUT2 #(
		.INIT('h8)
	) name8968 (
		_w10638_,
		_w12456_,
		_w13015_
	);
	LUT2 #(
		.INIT('h8)
	) name8969 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[8]/P0001 ,
		_w13016_
	);
	LUT2 #(
		.INIT('h4)
	) name8970 (
		_w10545_,
		_w12470_,
		_w13017_
	);
	LUT2 #(
		.INIT('h4)
	) name8971 (
		_w10579_,
		_w12466_,
		_w13018_
	);
	LUT2 #(
		.INIT('h4)
	) name8972 (
		_w10466_,
		_w12468_,
		_w13019_
	);
	LUT2 #(
		.INIT('h1)
	) name8973 (
		_w13017_,
		_w13018_,
		_w13020_
	);
	LUT2 #(
		.INIT('h4)
	) name8974 (
		_w13019_,
		_w13020_,
		_w13021_
	);
	LUT2 #(
		.INIT('h1)
	) name8975 (
		\emc_PMDoe_reg/NET0131 ,
		_w13021_,
		_w13022_
	);
	LUT2 #(
		.INIT('h2)
	) name8976 (
		_w12465_,
		_w13016_,
		_w13023_
	);
	LUT2 #(
		.INIT('h4)
	) name8977 (
		_w13022_,
		_w13023_,
		_w13024_
	);
	LUT2 #(
		.INIT('h8)
	) name8978 (
		\PM_rd2[8]_pad ,
		_w12478_,
		_w13025_
	);
	LUT2 #(
		.INIT('h2)
	) name8979 (
		\PM_rd0[8]_pad ,
		_w12504_,
		_w13026_
	);
	LUT2 #(
		.INIT('h8)
	) name8980 (
		\PM_rd4[8]_pad ,
		_w12488_,
		_w13027_
	);
	LUT2 #(
		.INIT('h8)
	) name8981 (
		\PM_rd6[8]_pad ,
		_w12483_,
		_w13028_
	);
	LUT2 #(
		.INIT('h8)
	) name8982 (
		\PM_rd7[8]_pad ,
		_w12485_,
		_w13029_
	);
	LUT2 #(
		.INIT('h8)
	) name8983 (
		\PM_rd3[8]_pad ,
		_w12493_,
		_w13030_
	);
	LUT2 #(
		.INIT('h8)
	) name8984 (
		\PM_rd1[8]_pad ,
		_w12491_,
		_w13031_
	);
	LUT2 #(
		.INIT('h8)
	) name8985 (
		\PM_rd5[8]_pad ,
		_w12495_,
		_w13032_
	);
	LUT2 #(
		.INIT('h1)
	) name8986 (
		_w12465_,
		_w13028_,
		_w13033_
	);
	LUT2 #(
		.INIT('h4)
	) name8987 (
		_w13029_,
		_w13033_,
		_w13034_
	);
	LUT2 #(
		.INIT('h1)
	) name8988 (
		_w13025_,
		_w13027_,
		_w13035_
	);
	LUT2 #(
		.INIT('h1)
	) name8989 (
		_w13030_,
		_w13031_,
		_w13036_
	);
	LUT2 #(
		.INIT('h4)
	) name8990 (
		_w13032_,
		_w13036_,
		_w13037_
	);
	LUT2 #(
		.INIT('h8)
	) name8991 (
		_w13034_,
		_w13035_,
		_w13038_
	);
	LUT2 #(
		.INIT('h8)
	) name8992 (
		_w13037_,
		_w13038_,
		_w13039_
	);
	LUT2 #(
		.INIT('h4)
	) name8993 (
		_w13026_,
		_w13039_,
		_w13040_
	);
	LUT2 #(
		.INIT('h1)
	) name8994 (
		_w13024_,
		_w13040_,
		_w13041_
	);
	LUT2 #(
		.INIT('h8)
	) name8995 (
		_w12452_,
		_w13041_,
		_w13042_
	);
	LUT2 #(
		.INIT('h1)
	) name8996 (
		_w13014_,
		_w13042_,
		_w13043_
	);
	LUT2 #(
		.INIT('h4)
	) name8997 (
		_w13015_,
		_w13043_,
		_w13044_
	);
	LUT2 #(
		.INIT('h2)
	) name8998 (
		_w12451_,
		_w13044_,
		_w13045_
	);
	LUT2 #(
		.INIT('h1)
	) name8999 (
		_w13013_,
		_w13045_,
		_w13046_
	);
	LUT2 #(
		.INIT('h8)
	) name9000 (
		\bdma_BCTL_reg[10]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w13047_
	);
	LUT2 #(
		.INIT('h8)
	) name9001 (
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w12454_,
		_w13048_
	);
	LUT2 #(
		.INIT('h8)
	) name9002 (
		_w10289_,
		_w12456_,
		_w13049_
	);
	LUT2 #(
		.INIT('h8)
	) name9003 (
		\emc_PMDoe_reg/NET0131 ,
		\emc_PMDreg_reg[9]/P0001 ,
		_w13050_
	);
	LUT2 #(
		.INIT('h4)
	) name9004 (
		_w10123_,
		_w12470_,
		_w13051_
	);
	LUT2 #(
		.INIT('h4)
	) name9005 (
		_w10230_,
		_w12466_,
		_w13052_
	);
	LUT2 #(
		.INIT('h4)
	) name9006 (
		_w10196_,
		_w12468_,
		_w13053_
	);
	LUT2 #(
		.INIT('h1)
	) name9007 (
		_w13051_,
		_w13052_,
		_w13054_
	);
	LUT2 #(
		.INIT('h4)
	) name9008 (
		_w13053_,
		_w13054_,
		_w13055_
	);
	LUT2 #(
		.INIT('h1)
	) name9009 (
		\emc_PMDoe_reg/NET0131 ,
		_w13055_,
		_w13056_
	);
	LUT2 #(
		.INIT('h2)
	) name9010 (
		_w12465_,
		_w13050_,
		_w13057_
	);
	LUT2 #(
		.INIT('h4)
	) name9011 (
		_w13056_,
		_w13057_,
		_w13058_
	);
	LUT2 #(
		.INIT('h8)
	) name9012 (
		\PM_rd2[9]_pad ,
		_w12478_,
		_w13059_
	);
	LUT2 #(
		.INIT('h2)
	) name9013 (
		\PM_rd0[9]_pad ,
		_w12504_,
		_w13060_
	);
	LUT2 #(
		.INIT('h8)
	) name9014 (
		\PM_rd4[9]_pad ,
		_w12488_,
		_w13061_
	);
	LUT2 #(
		.INIT('h8)
	) name9015 (
		\PM_rd6[9]_pad ,
		_w12483_,
		_w13062_
	);
	LUT2 #(
		.INIT('h8)
	) name9016 (
		\PM_rd7[9]_pad ,
		_w12485_,
		_w13063_
	);
	LUT2 #(
		.INIT('h8)
	) name9017 (
		\PM_rd3[9]_pad ,
		_w12493_,
		_w13064_
	);
	LUT2 #(
		.INIT('h8)
	) name9018 (
		\PM_rd1[9]_pad ,
		_w12491_,
		_w13065_
	);
	LUT2 #(
		.INIT('h8)
	) name9019 (
		\PM_rd5[9]_pad ,
		_w12495_,
		_w13066_
	);
	LUT2 #(
		.INIT('h1)
	) name9020 (
		_w12465_,
		_w13062_,
		_w13067_
	);
	LUT2 #(
		.INIT('h4)
	) name9021 (
		_w13063_,
		_w13067_,
		_w13068_
	);
	LUT2 #(
		.INIT('h1)
	) name9022 (
		_w13059_,
		_w13061_,
		_w13069_
	);
	LUT2 #(
		.INIT('h1)
	) name9023 (
		_w13064_,
		_w13065_,
		_w13070_
	);
	LUT2 #(
		.INIT('h4)
	) name9024 (
		_w13066_,
		_w13070_,
		_w13071_
	);
	LUT2 #(
		.INIT('h8)
	) name9025 (
		_w13068_,
		_w13069_,
		_w13072_
	);
	LUT2 #(
		.INIT('h8)
	) name9026 (
		_w13071_,
		_w13072_,
		_w13073_
	);
	LUT2 #(
		.INIT('h4)
	) name9027 (
		_w13060_,
		_w13073_,
		_w13074_
	);
	LUT2 #(
		.INIT('h1)
	) name9028 (
		_w13058_,
		_w13074_,
		_w13075_
	);
	LUT2 #(
		.INIT('h8)
	) name9029 (
		_w12452_,
		_w13075_,
		_w13076_
	);
	LUT2 #(
		.INIT('h1)
	) name9030 (
		_w13048_,
		_w13076_,
		_w13077_
	);
	LUT2 #(
		.INIT('h4)
	) name9031 (
		_w13049_,
		_w13077_,
		_w13078_
	);
	LUT2 #(
		.INIT('h2)
	) name9032 (
		_w12451_,
		_w13078_,
		_w13079_
	);
	LUT2 #(
		.INIT('h1)
	) name9033 (
		_w13047_,
		_w13079_,
		_w13080_
	);
	LUT2 #(
		.INIT('h1)
	) name9034 (
		\bdma_BM_cyc_reg/P0001 ,
		_w12451_,
		_w13081_
	);
	LUT2 #(
		.INIT('h1)
	) name9035 (
		_w12451_,
		_w12525_,
		_w13082_
	);
	LUT2 #(
		.INIT('h1)
	) name9036 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PCrd_1st_reg/NET0131 ,
		_w13083_
	);
	LUT2 #(
		.INIT('h1)
	) name9037 (
		\idma_DTMP_H_reg[0]/P0001 ,
		_w13083_,
		_w13084_
	);
	LUT2 #(
		.INIT('h4)
	) name9038 (
		\idma_DTMP_L_reg[0]/P0001 ,
		_w13083_,
		_w13085_
	);
	LUT2 #(
		.INIT('h1)
	) name9039 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13084_,
		_w13086_
	);
	LUT2 #(
		.INIT('h4)
	) name9040 (
		_w13085_,
		_w13086_,
		_w13087_
	);
	LUT2 #(
		.INIT('h2)
	) name9041 (
		\idma_DTMP_H_reg[10]/P0001 ,
		_w13083_,
		_w13088_
	);
	LUT2 #(
		.INIT('h1)
	) name9042 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13088_,
		_w13089_
	);
	LUT2 #(
		.INIT('h1)
	) name9043 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13083_,
		_w13090_
	);
	LUT2 #(
		.INIT('h8)
	) name9044 (
		\idma_DTMP_H_reg[11]/P0001 ,
		_w13090_,
		_w13091_
	);
	LUT2 #(
		.INIT('h8)
	) name9045 (
		\idma_DTMP_H_reg[12]/P0001 ,
		_w13090_,
		_w13092_
	);
	LUT2 #(
		.INIT('h2)
	) name9046 (
		\idma_DTMP_H_reg[13]/P0001 ,
		_w13083_,
		_w13093_
	);
	LUT2 #(
		.INIT('h1)
	) name9047 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13093_,
		_w13094_
	);
	LUT2 #(
		.INIT('h8)
	) name9048 (
		\idma_DTMP_H_reg[14]/P0001 ,
		_w13090_,
		_w13095_
	);
	LUT2 #(
		.INIT('h2)
	) name9049 (
		\idma_DTMP_H_reg[15]/P0001 ,
		_w13083_,
		_w13096_
	);
	LUT2 #(
		.INIT('h1)
	) name9050 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13096_,
		_w13097_
	);
	LUT2 #(
		.INIT('h1)
	) name9051 (
		\idma_DTMP_H_reg[1]/P0001 ,
		_w13083_,
		_w13098_
	);
	LUT2 #(
		.INIT('h4)
	) name9052 (
		\idma_DTMP_L_reg[1]/P0001 ,
		_w13083_,
		_w13099_
	);
	LUT2 #(
		.INIT('h1)
	) name9053 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13098_,
		_w13100_
	);
	LUT2 #(
		.INIT('h4)
	) name9054 (
		_w13099_,
		_w13100_,
		_w13101_
	);
	LUT2 #(
		.INIT('h8)
	) name9055 (
		\idma_DTMP_L_reg[2]/P0001 ,
		_w13083_,
		_w13102_
	);
	LUT2 #(
		.INIT('h2)
	) name9056 (
		\idma_DTMP_H_reg[2]/P0001 ,
		_w13083_,
		_w13103_
	);
	LUT2 #(
		.INIT('h1)
	) name9057 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13102_,
		_w13104_
	);
	LUT2 #(
		.INIT('h4)
	) name9058 (
		_w13103_,
		_w13104_,
		_w13105_
	);
	LUT2 #(
		.INIT('h1)
	) name9059 (
		\idma_DTMP_H_reg[3]/P0001 ,
		_w13083_,
		_w13106_
	);
	LUT2 #(
		.INIT('h4)
	) name9060 (
		\idma_DTMP_L_reg[3]/P0001 ,
		_w13083_,
		_w13107_
	);
	LUT2 #(
		.INIT('h1)
	) name9061 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13106_,
		_w13108_
	);
	LUT2 #(
		.INIT('h4)
	) name9062 (
		_w13107_,
		_w13108_,
		_w13109_
	);
	LUT2 #(
		.INIT('h1)
	) name9063 (
		\idma_DTMP_H_reg[4]/P0001 ,
		_w13083_,
		_w13110_
	);
	LUT2 #(
		.INIT('h4)
	) name9064 (
		\idma_DTMP_L_reg[4]/P0001 ,
		_w13083_,
		_w13111_
	);
	LUT2 #(
		.INIT('h1)
	) name9065 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13110_,
		_w13112_
	);
	LUT2 #(
		.INIT('h4)
	) name9066 (
		_w13111_,
		_w13112_,
		_w13113_
	);
	LUT2 #(
		.INIT('h8)
	) name9067 (
		\idma_DTMP_L_reg[5]/P0001 ,
		_w13083_,
		_w13114_
	);
	LUT2 #(
		.INIT('h2)
	) name9068 (
		\idma_DTMP_H_reg[5]/P0001 ,
		_w13083_,
		_w13115_
	);
	LUT2 #(
		.INIT('h1)
	) name9069 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13114_,
		_w13116_
	);
	LUT2 #(
		.INIT('h4)
	) name9070 (
		_w13115_,
		_w13116_,
		_w13117_
	);
	LUT2 #(
		.INIT('h1)
	) name9071 (
		\idma_DTMP_H_reg[6]/P0001 ,
		_w13083_,
		_w13118_
	);
	LUT2 #(
		.INIT('h4)
	) name9072 (
		\idma_DTMP_L_reg[6]/P0001 ,
		_w13083_,
		_w13119_
	);
	LUT2 #(
		.INIT('h1)
	) name9073 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13118_,
		_w13120_
	);
	LUT2 #(
		.INIT('h4)
	) name9074 (
		_w13119_,
		_w13120_,
		_w13121_
	);
	LUT2 #(
		.INIT('h8)
	) name9075 (
		\idma_DTMP_L_reg[7]/P0001 ,
		_w13083_,
		_w13122_
	);
	LUT2 #(
		.INIT('h2)
	) name9076 (
		\idma_DTMP_H_reg[7]/P0001 ,
		_w13083_,
		_w13123_
	);
	LUT2 #(
		.INIT('h1)
	) name9077 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w13122_,
		_w13124_
	);
	LUT2 #(
		.INIT('h4)
	) name9078 (
		_w13123_,
		_w13124_,
		_w13125_
	);
	LUT2 #(
		.INIT('h8)
	) name9079 (
		\idma_DTMP_H_reg[8]/P0001 ,
		_w13090_,
		_w13126_
	);
	LUT2 #(
		.INIT('h8)
	) name9080 (
		\idma_DTMP_H_reg[9]/P0001 ,
		_w13090_,
		_w13127_
	);
	LUT2 #(
		.INIT('h1)
	) name9081 (
		\idma_RDCMD_reg/P0001 ,
		\idma_RDcyc_reg/NET0131 ,
		_w13128_
	);
	LUT2 #(
		.INIT('h4)
	) name9082 (
		T_IMS_pad,
		\sice_OE_reg/P0001 ,
		_w13129_
	);
	LUT2 #(
		.INIT('h4)
	) name9083 (
		\memc_EXTC_E_reg/NET0131 ,
		\memc_Pwrite_E_reg/NET0131 ,
		_w13130_
	);
	LUT2 #(
		.INIT('h4)
	) name9084 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w13130_,
		_w13131_
	);
	LUT2 #(
		.INIT('h1)
	) name9085 (
		_w4099_,
		_w13131_,
		_w13132_
	);
	LUT2 #(
		.INIT('h4)
	) name9086 (
		_w4117_,
		_w13132_,
		_w13133_
	);
	LUT2 #(
		.INIT('h2)
	) name9087 (
		_w6020_,
		_w13133_,
		_w13134_
	);
	LUT2 #(
		.INIT('h8)
	) name9088 (
		_w6047_,
		_w13133_,
		_w13135_
	);
	LUT2 #(
		.INIT('h1)
	) name9089 (
		_w5936_,
		_w13133_,
		_w13136_
	);
	LUT2 #(
		.INIT('h1)
	) name9090 (
		_w13135_,
		_w13136_,
		_w13137_
	);
	LUT2 #(
		.INIT('h8)
	) name9091 (
		_w6164_,
		_w13137_,
		_w13138_
	);
	LUT2 #(
		.INIT('h4)
	) name9092 (
		_w13134_,
		_w13138_,
		_w13139_
	);
	LUT2 #(
		.INIT('h8)
	) name9093 (
		_w6980_,
		_w13135_,
		_w13140_
	);
	LUT2 #(
		.INIT('h8)
	) name9094 (
		_w6911_,
		_w13137_,
		_w13141_
	);
	LUT2 #(
		.INIT('h1)
	) name9095 (
		_w13134_,
		_w13136_,
		_w13142_
	);
	LUT2 #(
		.INIT('h4)
	) name9096 (
		_w13140_,
		_w13142_,
		_w13143_
	);
	LUT2 #(
		.INIT('h4)
	) name9097 (
		_w13141_,
		_w13143_,
		_w13144_
	);
	LUT2 #(
		.INIT('h2)
	) name9098 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w13145_
	);
	LUT2 #(
		.INIT('h8)
	) name9099 (
		_w5730_,
		_w13145_,
		_w13146_
	);
	LUT2 #(
		.INIT('h8)
	) name9100 (
		_w5727_,
		_w13146_,
		_w13147_
	);
	LUT2 #(
		.INIT('h4)
	) name9101 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w13147_,
		_w13148_
	);
	LUT2 #(
		.INIT('h1)
	) name9102 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w13149_
	);
	LUT2 #(
		.INIT('h8)
	) name9103 (
		_w5730_,
		_w13149_,
		_w13150_
	);
	LUT2 #(
		.INIT('h8)
	) name9104 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w13150_,
		_w13151_
	);
	LUT2 #(
		.INIT('h8)
	) name9105 (
		_w5727_,
		_w13151_,
		_w13152_
	);
	LUT2 #(
		.INIT('h1)
	) name9106 (
		_w13148_,
		_w13152_,
		_w13153_
	);
	LUT2 #(
		.INIT('h2)
	) name9107 (
		_w6913_,
		_w13153_,
		_w13154_
	);
	LUT2 #(
		.INIT('h8)
	) name9108 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w13154_,
		_w13155_
	);
	LUT2 #(
		.INIT('h4)
	) name9109 (
		_w4099_,
		_w13130_,
		_w13156_
	);
	LUT2 #(
		.INIT('h8)
	) name9110 (
		_w6931_,
		_w13156_,
		_w13157_
	);
	LUT2 #(
		.INIT('h2)
	) name9111 (
		_w6930_,
		_w13157_,
		_w13158_
	);
	LUT2 #(
		.INIT('h2)
	) name9112 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		_w13158_,
		_w13159_
	);
	LUT2 #(
		.INIT('h4)
	) name9113 (
		_w5717_,
		_w5880_,
		_w13160_
	);
	LUT2 #(
		.INIT('h8)
	) name9114 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w13160_,
		_w13161_
	);
	LUT2 #(
		.INIT('h1)
	) name9115 (
		_w6989_,
		_w13161_,
		_w13162_
	);
	LUT2 #(
		.INIT('h4)
	) name9116 (
		_w13159_,
		_w13162_,
		_w13163_
	);
	LUT2 #(
		.INIT('h1)
	) name9117 (
		_w13154_,
		_w13163_,
		_w13164_
	);
	LUT2 #(
		.INIT('h1)
	) name9118 (
		_w13137_,
		_w13155_,
		_w13165_
	);
	LUT2 #(
		.INIT('h4)
	) name9119 (
		_w13164_,
		_w13165_,
		_w13166_
	);
	LUT2 #(
		.INIT('h8)
	) name9120 (
		_w6968_,
		_w13137_,
		_w13167_
	);
	LUT2 #(
		.INIT('h1)
	) name9121 (
		_w13142_,
		_w13167_,
		_w13168_
	);
	LUT2 #(
		.INIT('h4)
	) name9122 (
		_w13166_,
		_w13168_,
		_w13169_
	);
	LUT2 #(
		.INIT('h1)
	) name9123 (
		_w13144_,
		_w13169_,
		_w13170_
	);
	LUT2 #(
		.INIT('h1)
	) name9124 (
		_w13139_,
		_w13170_,
		_w13171_
	);
	LUT2 #(
		.INIT('h8)
	) name9125 (
		_w7607_,
		_w13139_,
		_w13172_
	);
	LUT2 #(
		.INIT('h1)
	) name9126 (
		_w13171_,
		_w13172_,
		_w13173_
	);
	LUT2 #(
		.INIT('h8)
	) name9127 (
		_w8121_,
		_w13135_,
		_w13174_
	);
	LUT2 #(
		.INIT('h8)
	) name9128 (
		_w8211_,
		_w13137_,
		_w13175_
	);
	LUT2 #(
		.INIT('h2)
	) name9129 (
		_w13142_,
		_w13174_,
		_w13176_
	);
	LUT2 #(
		.INIT('h4)
	) name9130 (
		_w13175_,
		_w13176_,
		_w13177_
	);
	LUT2 #(
		.INIT('h8)
	) name9131 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w13154_,
		_w13178_
	);
	LUT2 #(
		.INIT('h2)
	) name9132 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w13158_,
		_w13179_
	);
	LUT2 #(
		.INIT('h8)
	) name9133 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w13160_,
		_w13180_
	);
	LUT2 #(
		.INIT('h1)
	) name9134 (
		_w8160_,
		_w13180_,
		_w13181_
	);
	LUT2 #(
		.INIT('h4)
	) name9135 (
		_w13179_,
		_w13181_,
		_w13182_
	);
	LUT2 #(
		.INIT('h1)
	) name9136 (
		_w13154_,
		_w13182_,
		_w13183_
	);
	LUT2 #(
		.INIT('h1)
	) name9137 (
		_w13137_,
		_w13178_,
		_w13184_
	);
	LUT2 #(
		.INIT('h4)
	) name9138 (
		_w13183_,
		_w13184_,
		_w13185_
	);
	LUT2 #(
		.INIT('h8)
	) name9139 (
		_w8129_,
		_w13137_,
		_w13186_
	);
	LUT2 #(
		.INIT('h1)
	) name9140 (
		_w13142_,
		_w13186_,
		_w13187_
	);
	LUT2 #(
		.INIT('h4)
	) name9141 (
		_w13185_,
		_w13187_,
		_w13188_
	);
	LUT2 #(
		.INIT('h1)
	) name9142 (
		_w13177_,
		_w13188_,
		_w13189_
	);
	LUT2 #(
		.INIT('h1)
	) name9143 (
		_w13139_,
		_w13189_,
		_w13190_
	);
	LUT2 #(
		.INIT('h8)
	) name9144 (
		_w7859_,
		_w13139_,
		_w13191_
	);
	LUT2 #(
		.INIT('h1)
	) name9145 (
		_w13190_,
		_w13191_,
		_w13192_
	);
	LUT2 #(
		.INIT('h8)
	) name9146 (
		_w8723_,
		_w13135_,
		_w13193_
	);
	LUT2 #(
		.INIT('h8)
	) name9147 (
		_w8813_,
		_w13137_,
		_w13194_
	);
	LUT2 #(
		.INIT('h2)
	) name9148 (
		_w13142_,
		_w13193_,
		_w13195_
	);
	LUT2 #(
		.INIT('h4)
	) name9149 (
		_w13194_,
		_w13195_,
		_w13196_
	);
	LUT2 #(
		.INIT('h8)
	) name9150 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w13154_,
		_w13197_
	);
	LUT2 #(
		.INIT('h2)
	) name9151 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		_w13158_,
		_w13198_
	);
	LUT2 #(
		.INIT('h8)
	) name9152 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w13160_,
		_w13199_
	);
	LUT2 #(
		.INIT('h1)
	) name9153 (
		_w8816_,
		_w13199_,
		_w13200_
	);
	LUT2 #(
		.INIT('h4)
	) name9154 (
		_w13198_,
		_w13200_,
		_w13201_
	);
	LUT2 #(
		.INIT('h1)
	) name9155 (
		_w13154_,
		_w13201_,
		_w13202_
	);
	LUT2 #(
		.INIT('h1)
	) name9156 (
		_w13137_,
		_w13197_,
		_w13203_
	);
	LUT2 #(
		.INIT('h4)
	) name9157 (
		_w13202_,
		_w13203_,
		_w13204_
	);
	LUT2 #(
		.INIT('h8)
	) name9158 (
		_w8731_,
		_w13137_,
		_w13205_
	);
	LUT2 #(
		.INIT('h1)
	) name9159 (
		_w13142_,
		_w13205_,
		_w13206_
	);
	LUT2 #(
		.INIT('h4)
	) name9160 (
		_w13204_,
		_w13206_,
		_w13207_
	);
	LUT2 #(
		.INIT('h1)
	) name9161 (
		_w13196_,
		_w13207_,
		_w13208_
	);
	LUT2 #(
		.INIT('h1)
	) name9162 (
		_w13139_,
		_w13208_,
		_w13209_
	);
	LUT2 #(
		.INIT('h8)
	) name9163 (
		_w8460_,
		_w13139_,
		_w13210_
	);
	LUT2 #(
		.INIT('h1)
	) name9164 (
		_w13209_,
		_w13210_,
		_w13211_
	);
	LUT2 #(
		.INIT('h8)
	) name9165 (
		_w9528_,
		_w13135_,
		_w13212_
	);
	LUT2 #(
		.INIT('h8)
	) name9166 (
		_w9559_,
		_w13137_,
		_w13213_
	);
	LUT2 #(
		.INIT('h2)
	) name9167 (
		_w13142_,
		_w13212_,
		_w13214_
	);
	LUT2 #(
		.INIT('h4)
	) name9168 (
		_w13213_,
		_w13214_,
		_w13215_
	);
	LUT2 #(
		.INIT('h8)
	) name9169 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w13154_,
		_w13216_
	);
	LUT2 #(
		.INIT('h2)
	) name9170 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		_w13158_,
		_w13217_
	);
	LUT2 #(
		.INIT('h8)
	) name9171 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w13160_,
		_w13218_
	);
	LUT2 #(
		.INIT('h1)
	) name9172 (
		_w9564_,
		_w13218_,
		_w13219_
	);
	LUT2 #(
		.INIT('h4)
	) name9173 (
		_w13217_,
		_w13219_,
		_w13220_
	);
	LUT2 #(
		.INIT('h1)
	) name9174 (
		_w13154_,
		_w13220_,
		_w13221_
	);
	LUT2 #(
		.INIT('h1)
	) name9175 (
		_w13137_,
		_w13216_,
		_w13222_
	);
	LUT2 #(
		.INIT('h4)
	) name9176 (
		_w13221_,
		_w13222_,
		_w13223_
	);
	LUT2 #(
		.INIT('h8)
	) name9177 (
		_w9520_,
		_w13137_,
		_w13224_
	);
	LUT2 #(
		.INIT('h1)
	) name9178 (
		_w13142_,
		_w13224_,
		_w13225_
	);
	LUT2 #(
		.INIT('h4)
	) name9179 (
		_w13223_,
		_w13225_,
		_w13226_
	);
	LUT2 #(
		.INIT('h1)
	) name9180 (
		_w13215_,
		_w13226_,
		_w13227_
	);
	LUT2 #(
		.INIT('h1)
	) name9181 (
		_w13139_,
		_w13227_,
		_w13228_
	);
	LUT2 #(
		.INIT('h8)
	) name9182 (
		_w9435_,
		_w13139_,
		_w13229_
	);
	LUT2 #(
		.INIT('h1)
	) name9183 (
		_w13228_,
		_w13229_,
		_w13230_
	);
	LUT2 #(
		.INIT('h8)
	) name9184 (
		_w9600_,
		_w13135_,
		_w13231_
	);
	LUT2 #(
		.INIT('h8)
	) name9185 (
		_w9625_,
		_w13137_,
		_w13232_
	);
	LUT2 #(
		.INIT('h2)
	) name9186 (
		_w13142_,
		_w13231_,
		_w13233_
	);
	LUT2 #(
		.INIT('h4)
	) name9187 (
		_w13232_,
		_w13233_,
		_w13234_
	);
	LUT2 #(
		.INIT('h8)
	) name9188 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w13154_,
		_w13235_
	);
	LUT2 #(
		.INIT('h2)
	) name9189 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		_w13158_,
		_w13236_
	);
	LUT2 #(
		.INIT('h8)
	) name9190 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w13160_,
		_w13237_
	);
	LUT2 #(
		.INIT('h1)
	) name9191 (
		_w9630_,
		_w13237_,
		_w13238_
	);
	LUT2 #(
		.INIT('h4)
	) name9192 (
		_w13236_,
		_w13238_,
		_w13239_
	);
	LUT2 #(
		.INIT('h1)
	) name9193 (
		_w13154_,
		_w13239_,
		_w13240_
	);
	LUT2 #(
		.INIT('h1)
	) name9194 (
		_w13137_,
		_w13235_,
		_w13241_
	);
	LUT2 #(
		.INIT('h4)
	) name9195 (
		_w13240_,
		_w13241_,
		_w13242_
	);
	LUT2 #(
		.INIT('h8)
	) name9196 (
		_w9592_,
		_w13137_,
		_w13243_
	);
	LUT2 #(
		.INIT('h1)
	) name9197 (
		_w13142_,
		_w13243_,
		_w13244_
	);
	LUT2 #(
		.INIT('h4)
	) name9198 (
		_w13242_,
		_w13244_,
		_w13245_
	);
	LUT2 #(
		.INIT('h1)
	) name9199 (
		_w13234_,
		_w13245_,
		_w13246_
	);
	LUT2 #(
		.INIT('h1)
	) name9200 (
		_w13139_,
		_w13246_,
		_w13247_
	);
	LUT2 #(
		.INIT('h8)
	) name9201 (
		_w8715_,
		_w13139_,
		_w13248_
	);
	LUT2 #(
		.INIT('h1)
	) name9202 (
		_w13247_,
		_w13248_,
		_w13249_
	);
	LUT2 #(
		.INIT('h8)
	) name9203 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w13154_,
		_w13250_
	);
	LUT2 #(
		.INIT('h2)
	) name9204 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		_w13158_,
		_w13251_
	);
	LUT2 #(
		.INIT('h8)
	) name9205 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w13160_,
		_w13252_
	);
	LUT2 #(
		.INIT('h1)
	) name9206 (
		_w9705_,
		_w13252_,
		_w13253_
	);
	LUT2 #(
		.INIT('h4)
	) name9207 (
		_w13251_,
		_w13253_,
		_w13254_
	);
	LUT2 #(
		.INIT('h1)
	) name9208 (
		_w13154_,
		_w13254_,
		_w13255_
	);
	LUT2 #(
		.INIT('h2)
	) name9209 (
		_w13136_,
		_w13250_,
		_w13256_
	);
	LUT2 #(
		.INIT('h4)
	) name9210 (
		_w13255_,
		_w13256_,
		_w13257_
	);
	LUT2 #(
		.INIT('h4)
	) name9211 (
		_w9666_,
		_w13135_,
		_w13258_
	);
	LUT2 #(
		.INIT('h4)
	) name9212 (
		_w9658_,
		_w13134_,
		_w13259_
	);
	LUT2 #(
		.INIT('h2)
	) name9213 (
		_w6164_,
		_w8113_,
		_w13260_
	);
	LUT2 #(
		.INIT('h4)
	) name9214 (
		_w6164_,
		_w9695_,
		_w13261_
	);
	LUT2 #(
		.INIT('h1)
	) name9215 (
		_w13260_,
		_w13261_,
		_w13262_
	);
	LUT2 #(
		.INIT('h4)
	) name9216 (
		_w13134_,
		_w13262_,
		_w13263_
	);
	LUT2 #(
		.INIT('h1)
	) name9217 (
		_w13259_,
		_w13263_,
		_w13264_
	);
	LUT2 #(
		.INIT('h1)
	) name9218 (
		_w13135_,
		_w13264_,
		_w13265_
	);
	LUT2 #(
		.INIT('h1)
	) name9219 (
		_w13136_,
		_w13258_,
		_w13266_
	);
	LUT2 #(
		.INIT('h4)
	) name9220 (
		_w13265_,
		_w13266_,
		_w13267_
	);
	LUT2 #(
		.INIT('h1)
	) name9221 (
		_w13257_,
		_w13267_,
		_w13268_
	);
	LUT2 #(
		.INIT('h4)
	) name9222 (
		_w10069_,
		_w13139_,
		_w13269_
	);
	LUT2 #(
		.INIT('h8)
	) name9223 (
		_w9797_,
		_w13134_,
		_w13270_
	);
	LUT2 #(
		.INIT('h4)
	) name9224 (
		_w6164_,
		_w9767_,
		_w13271_
	);
	LUT2 #(
		.INIT('h4)
	) name9225 (
		_w13134_,
		_w13271_,
		_w13272_
	);
	LUT2 #(
		.INIT('h1)
	) name9226 (
		_w13135_,
		_w13270_,
		_w13273_
	);
	LUT2 #(
		.INIT('h4)
	) name9227 (
		_w13272_,
		_w13273_,
		_w13274_
	);
	LUT2 #(
		.INIT('h4)
	) name9228 (
		_w9805_,
		_w13135_,
		_w13275_
	);
	LUT2 #(
		.INIT('h1)
	) name9229 (
		_w13136_,
		_w13275_,
		_w13276_
	);
	LUT2 #(
		.INIT('h4)
	) name9230 (
		_w13274_,
		_w13276_,
		_w13277_
	);
	LUT2 #(
		.INIT('h8)
	) name9231 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w13154_,
		_w13278_
	);
	LUT2 #(
		.INIT('h2)
	) name9232 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		_w13158_,
		_w13279_
	);
	LUT2 #(
		.INIT('h8)
	) name9233 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w13160_,
		_w13280_
	);
	LUT2 #(
		.INIT('h1)
	) name9234 (
		_w9812_,
		_w13280_,
		_w13281_
	);
	LUT2 #(
		.INIT('h4)
	) name9235 (
		_w13279_,
		_w13281_,
		_w13282_
	);
	LUT2 #(
		.INIT('h1)
	) name9236 (
		_w13154_,
		_w13282_,
		_w13283_
	);
	LUT2 #(
		.INIT('h2)
	) name9237 (
		_w13136_,
		_w13278_,
		_w13284_
	);
	LUT2 #(
		.INIT('h4)
	) name9238 (
		_w13283_,
		_w13284_,
		_w13285_
	);
	LUT2 #(
		.INIT('h1)
	) name9239 (
		_w13269_,
		_w13285_,
		_w13286_
	);
	LUT2 #(
		.INIT('h4)
	) name9240 (
		_w13277_,
		_w13286_,
		_w13287_
	);
	LUT2 #(
		.INIT('h4)
	) name9241 (
		_w10911_,
		_w13139_,
		_w13288_
	);
	LUT2 #(
		.INIT('h8)
	) name9242 (
		_w10364_,
		_w13134_,
		_w13289_
	);
	LUT2 #(
		.INIT('h4)
	) name9243 (
		_w6164_,
		_w10324_,
		_w13290_
	);
	LUT2 #(
		.INIT('h4)
	) name9244 (
		_w13134_,
		_w13290_,
		_w13291_
	);
	LUT2 #(
		.INIT('h1)
	) name9245 (
		_w13135_,
		_w13289_,
		_w13292_
	);
	LUT2 #(
		.INIT('h4)
	) name9246 (
		_w13291_,
		_w13292_,
		_w13293_
	);
	LUT2 #(
		.INIT('h4)
	) name9247 (
		_w10356_,
		_w13135_,
		_w13294_
	);
	LUT2 #(
		.INIT('h1)
	) name9248 (
		_w13136_,
		_w13294_,
		_w13295_
	);
	LUT2 #(
		.INIT('h4)
	) name9249 (
		_w13293_,
		_w13295_,
		_w13296_
	);
	LUT2 #(
		.INIT('h8)
	) name9250 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w13154_,
		_w13297_
	);
	LUT2 #(
		.INIT('h2)
	) name9251 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		_w13158_,
		_w13298_
	);
	LUT2 #(
		.INIT('h8)
	) name9252 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w13160_,
		_w13299_
	);
	LUT2 #(
		.INIT('h1)
	) name9253 (
		_w10349_,
		_w13299_,
		_w13300_
	);
	LUT2 #(
		.INIT('h4)
	) name9254 (
		_w13298_,
		_w13300_,
		_w13301_
	);
	LUT2 #(
		.INIT('h1)
	) name9255 (
		_w13154_,
		_w13301_,
		_w13302_
	);
	LUT2 #(
		.INIT('h2)
	) name9256 (
		_w13136_,
		_w13297_,
		_w13303_
	);
	LUT2 #(
		.INIT('h4)
	) name9257 (
		_w13302_,
		_w13303_,
		_w13304_
	);
	LUT2 #(
		.INIT('h1)
	) name9258 (
		_w13288_,
		_w13304_,
		_w13305_
	);
	LUT2 #(
		.INIT('h4)
	) name9259 (
		_w13296_,
		_w13305_,
		_w13306_
	);
	LUT2 #(
		.INIT('h4)
	) name9260 (
		_w11525_,
		_w13139_,
		_w13307_
	);
	LUT2 #(
		.INIT('h8)
	) name9261 (
		_w10975_,
		_w13134_,
		_w13308_
	);
	LUT2 #(
		.INIT('h4)
	) name9262 (
		_w6164_,
		_w10930_,
		_w13309_
	);
	LUT2 #(
		.INIT('h4)
	) name9263 (
		_w13134_,
		_w13309_,
		_w13310_
	);
	LUT2 #(
		.INIT('h1)
	) name9264 (
		_w13135_,
		_w13308_,
		_w13311_
	);
	LUT2 #(
		.INIT('h4)
	) name9265 (
		_w13310_,
		_w13311_,
		_w13312_
	);
	LUT2 #(
		.INIT('h4)
	) name9266 (
		_w10967_,
		_w13135_,
		_w13313_
	);
	LUT2 #(
		.INIT('h1)
	) name9267 (
		_w13136_,
		_w13313_,
		_w13314_
	);
	LUT2 #(
		.INIT('h4)
	) name9268 (
		_w13312_,
		_w13314_,
		_w13315_
	);
	LUT2 #(
		.INIT('h8)
	) name9269 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w13154_,
		_w13316_
	);
	LUT2 #(
		.INIT('h2)
	) name9270 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		_w13158_,
		_w13317_
	);
	LUT2 #(
		.INIT('h8)
	) name9271 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w13160_,
		_w13318_
	);
	LUT2 #(
		.INIT('h1)
	) name9272 (
		_w10960_,
		_w13318_,
		_w13319_
	);
	LUT2 #(
		.INIT('h4)
	) name9273 (
		_w13317_,
		_w13319_,
		_w13320_
	);
	LUT2 #(
		.INIT('h1)
	) name9274 (
		_w13154_,
		_w13320_,
		_w13321_
	);
	LUT2 #(
		.INIT('h2)
	) name9275 (
		_w13136_,
		_w13316_,
		_w13322_
	);
	LUT2 #(
		.INIT('h4)
	) name9276 (
		_w13321_,
		_w13322_,
		_w13323_
	);
	LUT2 #(
		.INIT('h1)
	) name9277 (
		_w13307_,
		_w13323_,
		_w13324_
	);
	LUT2 #(
		.INIT('h4)
	) name9278 (
		_w13315_,
		_w13324_,
		_w13325_
	);
	LUT2 #(
		.INIT('h4)
	) name9279 (
		_w11265_,
		_w13139_,
		_w13326_
	);
	LUT2 #(
		.INIT('h8)
	) name9280 (
		_w11548_,
		_w13134_,
		_w13327_
	);
	LUT2 #(
		.INIT('h4)
	) name9281 (
		_w6164_,
		_w11579_,
		_w13328_
	);
	LUT2 #(
		.INIT('h4)
	) name9282 (
		_w13134_,
		_w13328_,
		_w13329_
	);
	LUT2 #(
		.INIT('h1)
	) name9283 (
		_w13135_,
		_w13327_,
		_w13330_
	);
	LUT2 #(
		.INIT('h4)
	) name9284 (
		_w13329_,
		_w13330_,
		_w13331_
	);
	LUT2 #(
		.INIT('h4)
	) name9285 (
		_w11540_,
		_w13135_,
		_w13332_
	);
	LUT2 #(
		.INIT('h1)
	) name9286 (
		_w13136_,
		_w13332_,
		_w13333_
	);
	LUT2 #(
		.INIT('h4)
	) name9287 (
		_w13331_,
		_w13333_,
		_w13334_
	);
	LUT2 #(
		.INIT('h8)
	) name9288 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w13154_,
		_w13335_
	);
	LUT2 #(
		.INIT('h2)
	) name9289 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		_w13158_,
		_w13336_
	);
	LUT2 #(
		.INIT('h8)
	) name9290 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w13160_,
		_w13337_
	);
	LUT2 #(
		.INIT('h1)
	) name9291 (
		_w11532_,
		_w13337_,
		_w13338_
	);
	LUT2 #(
		.INIT('h4)
	) name9292 (
		_w13336_,
		_w13338_,
		_w13339_
	);
	LUT2 #(
		.INIT('h1)
	) name9293 (
		_w13154_,
		_w13339_,
		_w13340_
	);
	LUT2 #(
		.INIT('h2)
	) name9294 (
		_w13136_,
		_w13335_,
		_w13341_
	);
	LUT2 #(
		.INIT('h4)
	) name9295 (
		_w13340_,
		_w13341_,
		_w13342_
	);
	LUT2 #(
		.INIT('h1)
	) name9296 (
		_w13326_,
		_w13342_,
		_w13343_
	);
	LUT2 #(
		.INIT('h4)
	) name9297 (
		_w13334_,
		_w13343_,
		_w13344_
	);
	LUT2 #(
		.INIT('h4)
	) name9298 (
		_w10638_,
		_w13139_,
		_w13345_
	);
	LUT2 #(
		.INIT('h8)
	) name9299 (
		_w11617_,
		_w13134_,
		_w13346_
	);
	LUT2 #(
		.INIT('h4)
	) name9300 (
		_w6164_,
		_w11654_,
		_w13347_
	);
	LUT2 #(
		.INIT('h4)
	) name9301 (
		_w13134_,
		_w13347_,
		_w13348_
	);
	LUT2 #(
		.INIT('h1)
	) name9302 (
		_w13135_,
		_w13346_,
		_w13349_
	);
	LUT2 #(
		.INIT('h4)
	) name9303 (
		_w13348_,
		_w13349_,
		_w13350_
	);
	LUT2 #(
		.INIT('h4)
	) name9304 (
		_w11609_,
		_w13135_,
		_w13351_
	);
	LUT2 #(
		.INIT('h1)
	) name9305 (
		_w13136_,
		_w13351_,
		_w13352_
	);
	LUT2 #(
		.INIT('h4)
	) name9306 (
		_w13350_,
		_w13352_,
		_w13353_
	);
	LUT2 #(
		.INIT('h8)
	) name9307 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w13154_,
		_w13354_
	);
	LUT2 #(
		.INIT('h2)
	) name9308 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		_w13158_,
		_w13355_
	);
	LUT2 #(
		.INIT('h8)
	) name9309 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w13160_,
		_w13356_
	);
	LUT2 #(
		.INIT('h1)
	) name9310 (
		_w11625_,
		_w13356_,
		_w13357_
	);
	LUT2 #(
		.INIT('h4)
	) name9311 (
		_w13355_,
		_w13357_,
		_w13358_
	);
	LUT2 #(
		.INIT('h1)
	) name9312 (
		_w13154_,
		_w13358_,
		_w13359_
	);
	LUT2 #(
		.INIT('h2)
	) name9313 (
		_w13136_,
		_w13354_,
		_w13360_
	);
	LUT2 #(
		.INIT('h4)
	) name9314 (
		_w13359_,
		_w13360_,
		_w13361_
	);
	LUT2 #(
		.INIT('h1)
	) name9315 (
		_w13345_,
		_w13361_,
		_w13362_
	);
	LUT2 #(
		.INIT('h4)
	) name9316 (
		_w13353_,
		_w13362_,
		_w13363_
	);
	LUT2 #(
		.INIT('h4)
	) name9317 (
		_w10289_,
		_w13139_,
		_w13364_
	);
	LUT2 #(
		.INIT('h8)
	) name9318 (
		_w11676_,
		_w13134_,
		_w13365_
	);
	LUT2 #(
		.INIT('h4)
	) name9319 (
		_w6164_,
		_w11720_,
		_w13366_
	);
	LUT2 #(
		.INIT('h4)
	) name9320 (
		_w13134_,
		_w13366_,
		_w13367_
	);
	LUT2 #(
		.INIT('h1)
	) name9321 (
		_w13135_,
		_w13365_,
		_w13368_
	);
	LUT2 #(
		.INIT('h4)
	) name9322 (
		_w13367_,
		_w13368_,
		_w13369_
	);
	LUT2 #(
		.INIT('h4)
	) name9323 (
		_w11668_,
		_w13135_,
		_w13370_
	);
	LUT2 #(
		.INIT('h1)
	) name9324 (
		_w13136_,
		_w13370_,
		_w13371_
	);
	LUT2 #(
		.INIT('h4)
	) name9325 (
		_w13369_,
		_w13371_,
		_w13372_
	);
	LUT2 #(
		.INIT('h8)
	) name9326 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w13154_,
		_w13373_
	);
	LUT2 #(
		.INIT('h2)
	) name9327 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		_w13158_,
		_w13374_
	);
	LUT2 #(
		.INIT('h8)
	) name9328 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w13160_,
		_w13375_
	);
	LUT2 #(
		.INIT('h1)
	) name9329 (
		_w11687_,
		_w13375_,
		_w13376_
	);
	LUT2 #(
		.INIT('h4)
	) name9330 (
		_w13374_,
		_w13376_,
		_w13377_
	);
	LUT2 #(
		.INIT('h1)
	) name9331 (
		_w13154_,
		_w13377_,
		_w13378_
	);
	LUT2 #(
		.INIT('h2)
	) name9332 (
		_w13136_,
		_w13373_,
		_w13379_
	);
	LUT2 #(
		.INIT('h4)
	) name9333 (
		_w13378_,
		_w13379_,
		_w13380_
	);
	LUT2 #(
		.INIT('h1)
	) name9334 (
		_w13364_,
		_w13380_,
		_w13381_
	);
	LUT2 #(
		.INIT('h4)
	) name9335 (
		_w13372_,
		_w13381_,
		_w13382_
	);
	LUT2 #(
		.INIT('h8)
	) name9336 (
		_w5880_,
		_w5882_,
		_w13383_
	);
	LUT2 #(
		.INIT('h8)
	) name9337 (
		_w11761_,
		_w13383_,
		_w13384_
	);
	LUT2 #(
		.INIT('h8)
	) name9338 (
		_w6913_,
		_w13148_,
		_w13385_
	);
	LUT2 #(
		.INIT('h4)
	) name9339 (
		_w7362_,
		_w12473_,
		_w13386_
	);
	LUT2 #(
		.INIT('h4)
	) name9340 (
		_w13385_,
		_w13386_,
		_w13387_
	);
	LUT2 #(
		.INIT('h4)
	) name9341 (
		\bdma_BRdataBUF_reg[8]/P0001 ,
		_w13385_,
		_w13388_
	);
	LUT2 #(
		.INIT('h1)
	) name9342 (
		_w13387_,
		_w13388_,
		_w13389_
	);
	LUT2 #(
		.INIT('h1)
	) name9343 (
		_w13384_,
		_w13389_,
		_w13390_
	);
	LUT2 #(
		.INIT('h4)
	) name9344 (
		\idma_DTMP_H_reg[0]/P0001 ,
		_w13384_,
		_w13391_
	);
	LUT2 #(
		.INIT('h1)
	) name9345 (
		_w13390_,
		_w13391_,
		_w13392_
	);
	LUT2 #(
		.INIT('h4)
	) name9346 (
		_w7664_,
		_w12536_,
		_w13393_
	);
	LUT2 #(
		.INIT('h4)
	) name9347 (
		_w13385_,
		_w13393_,
		_w13394_
	);
	LUT2 #(
		.INIT('h4)
	) name9348 (
		\bdma_BRdataBUF_reg[18]/P0001 ,
		_w13385_,
		_w13395_
	);
	LUT2 #(
		.INIT('h1)
	) name9349 (
		_w13394_,
		_w13395_,
		_w13396_
	);
	LUT2 #(
		.INIT('h1)
	) name9350 (
		_w13384_,
		_w13396_,
		_w13397_
	);
	LUT2 #(
		.INIT('h4)
	) name9351 (
		\idma_DTMP_H_reg[10]/P0001 ,
		_w13384_,
		_w13398_
	);
	LUT2 #(
		.INIT('h1)
	) name9352 (
		_w13397_,
		_w13398_,
		_w13399_
	);
	LUT2 #(
		.INIT('h4)
	) name9353 (
		_w8266_,
		_w12570_,
		_w13400_
	);
	LUT2 #(
		.INIT('h4)
	) name9354 (
		_w13385_,
		_w13400_,
		_w13401_
	);
	LUT2 #(
		.INIT('h4)
	) name9355 (
		\bdma_BRdataBUF_reg[19]/P0001 ,
		_w13385_,
		_w13402_
	);
	LUT2 #(
		.INIT('h1)
	) name9356 (
		_w13401_,
		_w13402_,
		_w13403_
	);
	LUT2 #(
		.INIT('h1)
	) name9357 (
		_w13384_,
		_w13403_,
		_w13404_
	);
	LUT2 #(
		.INIT('h4)
	) name9358 (
		\idma_DTMP_H_reg[11]/P0001 ,
		_w13384_,
		_w13405_
	);
	LUT2 #(
		.INIT('h1)
	) name9359 (
		_w13404_,
		_w13405_,
		_w13406_
	);
	LUT2 #(
		.INIT('h4)
	) name9360 (
		_w8983_,
		_w12604_,
		_w13407_
	);
	LUT2 #(
		.INIT('h4)
	) name9361 (
		_w13385_,
		_w13407_,
		_w13408_
	);
	LUT2 #(
		.INIT('h4)
	) name9362 (
		\bdma_BRdataBUF_reg[20]/P0001 ,
		_w13385_,
		_w13409_
	);
	LUT2 #(
		.INIT('h1)
	) name9363 (
		_w13408_,
		_w13409_,
		_w13410_
	);
	LUT2 #(
		.INIT('h1)
	) name9364 (
		_w13384_,
		_w13410_,
		_w13411_
	);
	LUT2 #(
		.INIT('h4)
	) name9365 (
		\idma_DTMP_H_reg[12]/P0001 ,
		_w13384_,
		_w13412_
	);
	LUT2 #(
		.INIT('h1)
	) name9366 (
		_w13411_,
		_w13412_,
		_w13413_
	);
	LUT2 #(
		.INIT('h4)
	) name9367 (
		_w7067_,
		_w12638_,
		_w13414_
	);
	LUT2 #(
		.INIT('h4)
	) name9368 (
		_w13385_,
		_w13414_,
		_w13415_
	);
	LUT2 #(
		.INIT('h4)
	) name9369 (
		\bdma_BRdataBUF_reg[21]/P0001 ,
		_w13385_,
		_w13416_
	);
	LUT2 #(
		.INIT('h1)
	) name9370 (
		_w13415_,
		_w13416_,
		_w13417_
	);
	LUT2 #(
		.INIT('h1)
	) name9371 (
		_w13384_,
		_w13417_,
		_w13418_
	);
	LUT2 #(
		.INIT('h4)
	) name9372 (
		\idma_DTMP_H_reg[13]/P0001 ,
		_w13384_,
		_w13419_
	);
	LUT2 #(
		.INIT('h1)
	) name9373 (
		_w13418_,
		_w13419_,
		_w13420_
	);
	LUT2 #(
		.INIT('h4)
	) name9374 (
		_w11818_,
		_w12695_,
		_w13421_
	);
	LUT2 #(
		.INIT('h4)
	) name9375 (
		_w13385_,
		_w13421_,
		_w13422_
	);
	LUT2 #(
		.INIT('h4)
	) name9376 (
		\bdma_BRdataBUF_reg[22]/P0001 ,
		_w13385_,
		_w13423_
	);
	LUT2 #(
		.INIT('h1)
	) name9377 (
		_w13422_,
		_w13423_,
		_w13424_
	);
	LUT2 #(
		.INIT('h1)
	) name9378 (
		_w13384_,
		_w13424_,
		_w13425_
	);
	LUT2 #(
		.INIT('h4)
	) name9379 (
		\idma_DTMP_H_reg[14]/P0001 ,
		_w13384_,
		_w13426_
	);
	LUT2 #(
		.INIT('h1)
	) name9380 (
		_w13425_,
		_w13426_,
		_w13427_
	);
	LUT2 #(
		.INIT('h4)
	) name9381 (
		_w11964_,
		_w12751_,
		_w13428_
	);
	LUT2 #(
		.INIT('h4)
	) name9382 (
		_w13385_,
		_w13428_,
		_w13429_
	);
	LUT2 #(
		.INIT('h4)
	) name9383 (
		\bdma_BRdataBUF_reg[23]/P0001 ,
		_w13385_,
		_w13430_
	);
	LUT2 #(
		.INIT('h1)
	) name9384 (
		_w13429_,
		_w13430_,
		_w13431_
	);
	LUT2 #(
		.INIT('h1)
	) name9385 (
		_w13384_,
		_w13431_,
		_w13432_
	);
	LUT2 #(
		.INIT('h4)
	) name9386 (
		\idma_DTMP_H_reg[15]/P0001 ,
		_w13384_,
		_w13433_
	);
	LUT2 #(
		.INIT('h1)
	) name9387 (
		_w13432_,
		_w13433_,
		_w13434_
	);
	LUT2 #(
		.INIT('h4)
	) name9388 (
		_w9202_,
		_w12782_,
		_w13435_
	);
	LUT2 #(
		.INIT('h4)
	) name9389 (
		_w13385_,
		_w13435_,
		_w13436_
	);
	LUT2 #(
		.INIT('h4)
	) name9390 (
		\bdma_BRdataBUF_reg[9]/P0001 ,
		_w13385_,
		_w13437_
	);
	LUT2 #(
		.INIT('h1)
	) name9391 (
		_w13436_,
		_w13437_,
		_w13438_
	);
	LUT2 #(
		.INIT('h1)
	) name9392 (
		_w13384_,
		_w13438_,
		_w13439_
	);
	LUT2 #(
		.INIT('h4)
	) name9393 (
		\idma_DTMP_H_reg[1]/P0001 ,
		_w13384_,
		_w13440_
	);
	LUT2 #(
		.INIT('h1)
	) name9394 (
		_w13439_,
		_w13440_,
		_w13441_
	);
	LUT2 #(
		.INIT('h4)
	) name9395 (
		_w8482_,
		_w12816_,
		_w13442_
	);
	LUT2 #(
		.INIT('h4)
	) name9396 (
		_w13385_,
		_w13442_,
		_w13443_
	);
	LUT2 #(
		.INIT('h4)
	) name9397 (
		\bdma_BRdataBUF_reg[10]/P0001 ,
		_w13385_,
		_w13444_
	);
	LUT2 #(
		.INIT('h1)
	) name9398 (
		_w13443_,
		_w13444_,
		_w13445_
	);
	LUT2 #(
		.INIT('h1)
	) name9399 (
		_w13384_,
		_w13445_,
		_w13446_
	);
	LUT2 #(
		.INIT('h4)
	) name9400 (
		\idma_DTMP_H_reg[2]/P0001 ,
		_w13384_,
		_w13447_
	);
	LUT2 #(
		.INIT('h1)
	) name9401 (
		_w13446_,
		_w13447_,
		_w13448_
	);
	LUT2 #(
		.INIT('h4)
	) name9402 (
		_w7882_,
		_w12850_,
		_w13449_
	);
	LUT2 #(
		.INIT('h4)
	) name9403 (
		_w13385_,
		_w13449_,
		_w13450_
	);
	LUT2 #(
		.INIT('h4)
	) name9404 (
		\bdma_BRdataBUF_reg[11]/P0001 ,
		_w13385_,
		_w13451_
	);
	LUT2 #(
		.INIT('h1)
	) name9405 (
		_w13450_,
		_w13451_,
		_w13452_
	);
	LUT2 #(
		.INIT('h1)
	) name9406 (
		_w13384_,
		_w13452_,
		_w13453_
	);
	LUT2 #(
		.INIT('h4)
	) name9407 (
		\idma_DTMP_H_reg[3]/P0001 ,
		_w13384_,
		_w13454_
	);
	LUT2 #(
		.INIT('h1)
	) name9408 (
		_w13453_,
		_w13454_,
		_w13455_
	);
	LUT2 #(
		.INIT('h4)
	) name9409 (
		_w9842_,
		_w12884_,
		_w13456_
	);
	LUT2 #(
		.INIT('h4)
	) name9410 (
		_w13385_,
		_w13456_,
		_w13457_
	);
	LUT2 #(
		.INIT('h4)
	) name9411 (
		\bdma_BRdataBUF_reg[12]/P0001 ,
		_w13385_,
		_w13458_
	);
	LUT2 #(
		.INIT('h1)
	) name9412 (
		_w13457_,
		_w13458_,
		_w13459_
	);
	LUT2 #(
		.INIT('h1)
	) name9413 (
		_w13384_,
		_w13459_,
		_w13460_
	);
	LUT2 #(
		.INIT('h4)
	) name9414 (
		\idma_DTMP_H_reg[4]/P0001 ,
		_w13384_,
		_w13461_
	);
	LUT2 #(
		.INIT('h1)
	) name9415 (
		_w13460_,
		_w13461_,
		_w13462_
	);
	LUT2 #(
		.INIT('h4)
	) name9416 (
		_w10683_,
		_w12918_,
		_w13463_
	);
	LUT2 #(
		.INIT('h4)
	) name9417 (
		_w13385_,
		_w13463_,
		_w13464_
	);
	LUT2 #(
		.INIT('h4)
	) name9418 (
		\bdma_BRdataBUF_reg[13]/P0001 ,
		_w13385_,
		_w13465_
	);
	LUT2 #(
		.INIT('h1)
	) name9419 (
		_w13464_,
		_w13465_,
		_w13466_
	);
	LUT2 #(
		.INIT('h1)
	) name9420 (
		_w13384_,
		_w13466_,
		_w13467_
	);
	LUT2 #(
		.INIT('h4)
	) name9421 (
		\idma_DTMP_H_reg[5]/P0001 ,
		_w13384_,
		_w13468_
	);
	LUT2 #(
		.INIT('h1)
	) name9422 (
		_w13467_,
		_w13468_,
		_w13469_
	);
	LUT2 #(
		.INIT('h4)
	) name9423 (
		_w11300_,
		_w12968_,
		_w13470_
	);
	LUT2 #(
		.INIT('h4)
	) name9424 (
		_w13385_,
		_w13470_,
		_w13471_
	);
	LUT2 #(
		.INIT('h4)
	) name9425 (
		\bdma_BRdataBUF_reg[14]/P0001 ,
		_w13385_,
		_w13472_
	);
	LUT2 #(
		.INIT('h1)
	) name9426 (
		_w13471_,
		_w13472_,
		_w13473_
	);
	LUT2 #(
		.INIT('h1)
	) name9427 (
		_w13384_,
		_w13473_,
		_w13474_
	);
	LUT2 #(
		.INIT('h4)
	) name9428 (
		\idma_DTMP_H_reg[6]/P0001 ,
		_w13384_,
		_w13475_
	);
	LUT2 #(
		.INIT('h1)
	) name9429 (
		_w13474_,
		_w13475_,
		_w13476_
	);
	LUT2 #(
		.INIT('h4)
	) name9430 (
		_w11051_,
		_w12986_,
		_w13477_
	);
	LUT2 #(
		.INIT('h4)
	) name9431 (
		_w13385_,
		_w13477_,
		_w13478_
	);
	LUT2 #(
		.INIT('h4)
	) name9432 (
		\bdma_BRdataBUF_reg[15]/P0001 ,
		_w13385_,
		_w13479_
	);
	LUT2 #(
		.INIT('h1)
	) name9433 (
		_w13478_,
		_w13479_,
		_w13480_
	);
	LUT2 #(
		.INIT('h1)
	) name9434 (
		_w13384_,
		_w13480_,
		_w13481_
	);
	LUT2 #(
		.INIT('h4)
	) name9435 (
		\idma_DTMP_H_reg[7]/P0001 ,
		_w13384_,
		_w13482_
	);
	LUT2 #(
		.INIT('h1)
	) name9436 (
		_w13481_,
		_w13482_,
		_w13483_
	);
	LUT2 #(
		.INIT('h4)
	) name9437 (
		_w10442_,
		_w13021_,
		_w13484_
	);
	LUT2 #(
		.INIT('h4)
	) name9438 (
		_w13385_,
		_w13484_,
		_w13485_
	);
	LUT2 #(
		.INIT('h4)
	) name9439 (
		\bdma_BRdataBUF_reg[16]/P0001 ,
		_w13385_,
		_w13486_
	);
	LUT2 #(
		.INIT('h1)
	) name9440 (
		_w13485_,
		_w13486_,
		_w13487_
	);
	LUT2 #(
		.INIT('h1)
	) name9441 (
		_w13384_,
		_w13487_,
		_w13488_
	);
	LUT2 #(
		.INIT('h4)
	) name9442 (
		\idma_DTMP_H_reg[8]/P0001 ,
		_w13384_,
		_w13489_
	);
	LUT2 #(
		.INIT('h1)
	) name9443 (
		_w13488_,
		_w13489_,
		_w13490_
	);
	LUT2 #(
		.INIT('h4)
	) name9444 (
		_w10093_,
		_w13055_,
		_w13491_
	);
	LUT2 #(
		.INIT('h4)
	) name9445 (
		_w13385_,
		_w13491_,
		_w13492_
	);
	LUT2 #(
		.INIT('h4)
	) name9446 (
		\bdma_BRdataBUF_reg[17]/P0001 ,
		_w13385_,
		_w13493_
	);
	LUT2 #(
		.INIT('h1)
	) name9447 (
		_w13492_,
		_w13493_,
		_w13494_
	);
	LUT2 #(
		.INIT('h1)
	) name9448 (
		_w13384_,
		_w13494_,
		_w13495_
	);
	LUT2 #(
		.INIT('h4)
	) name9449 (
		\idma_DTMP_H_reg[9]/P0001 ,
		_w13384_,
		_w13496_
	);
	LUT2 #(
		.INIT('h1)
	) name9450 (
		_w13495_,
		_w13496_,
		_w13497_
	);
	LUT2 #(
		.INIT('h8)
	) name9451 (
		_w9178_,
		_w13139_,
		_w13498_
	);
	LUT2 #(
		.INIT('h8)
	) name9452 (
		_w5936_,
		_w13134_,
		_w13499_
	);
	LUT2 #(
		.INIT('h4)
	) name9453 (
		_w8853_,
		_w13499_,
		_w13500_
	);
	LUT2 #(
		.INIT('h4)
	) name9454 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w13154_,
		_w13501_
	);
	LUT2 #(
		.INIT('h2)
	) name9455 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w13158_,
		_w13502_
	);
	LUT2 #(
		.INIT('h8)
	) name9456 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w13160_,
		_w13503_
	);
	LUT2 #(
		.INIT('h1)
	) name9457 (
		_w8838_,
		_w13503_,
		_w13504_
	);
	LUT2 #(
		.INIT('h4)
	) name9458 (
		_w13154_,
		_w13504_,
		_w13505_
	);
	LUT2 #(
		.INIT('h4)
	) name9459 (
		_w13502_,
		_w13505_,
		_w13506_
	);
	LUT2 #(
		.INIT('h2)
	) name9460 (
		_w13136_,
		_w13501_,
		_w13507_
	);
	LUT2 #(
		.INIT('h4)
	) name9461 (
		_w13506_,
		_w13507_,
		_w13508_
	);
	LUT2 #(
		.INIT('h8)
	) name9462 (
		_w8945_,
		_w13137_,
		_w13509_
	);
	LUT2 #(
		.INIT('h4)
	) name9463 (
		_w13138_,
		_w13142_,
		_w13510_
	);
	LUT2 #(
		.INIT('h2)
	) name9464 (
		_w8845_,
		_w13137_,
		_w13511_
	);
	LUT2 #(
		.INIT('h2)
	) name9465 (
		_w13510_,
		_w13511_,
		_w13512_
	);
	LUT2 #(
		.INIT('h4)
	) name9466 (
		_w13509_,
		_w13512_,
		_w13513_
	);
	LUT2 #(
		.INIT('h1)
	) name9467 (
		_w13500_,
		_w13508_,
		_w13514_
	);
	LUT2 #(
		.INIT('h4)
	) name9468 (
		_w13498_,
		_w13514_,
		_w13515_
	);
	LUT2 #(
		.INIT('h4)
	) name9469 (
		_w13513_,
		_w13515_,
		_w13516_
	);
	LUT2 #(
		.INIT('h4)
	) name9470 (
		PM_bdry_sel_pad,
		_w13516_,
		_w13517_
	);
	LUT2 #(
		.INIT('h8)
	) name9471 (
		_w7340_,
		_w13139_,
		_w13518_
	);
	LUT2 #(
		.INIT('h4)
	) name9472 (
		_w9460_,
		_w13499_,
		_w13519_
	);
	LUT2 #(
		.INIT('h4)
	) name9473 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w13154_,
		_w13520_
	);
	LUT2 #(
		.INIT('h2)
	) name9474 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		_w13158_,
		_w13521_
	);
	LUT2 #(
		.INIT('h8)
	) name9475 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w13160_,
		_w13522_
	);
	LUT2 #(
		.INIT('h1)
	) name9476 (
		_w9442_,
		_w13522_,
		_w13523_
	);
	LUT2 #(
		.INIT('h4)
	) name9477 (
		_w13154_,
		_w13523_,
		_w13524_
	);
	LUT2 #(
		.INIT('h4)
	) name9478 (
		_w13521_,
		_w13524_,
		_w13525_
	);
	LUT2 #(
		.INIT('h2)
	) name9479 (
		_w13136_,
		_w13520_,
		_w13526_
	);
	LUT2 #(
		.INIT('h4)
	) name9480 (
		_w13525_,
		_w13526_,
		_w13527_
	);
	LUT2 #(
		.INIT('h8)
	) name9481 (
		_w9497_,
		_w13137_,
		_w13528_
	);
	LUT2 #(
		.INIT('h2)
	) name9482 (
		_w9452_,
		_w13137_,
		_w13529_
	);
	LUT2 #(
		.INIT('h2)
	) name9483 (
		_w13510_,
		_w13529_,
		_w13530_
	);
	LUT2 #(
		.INIT('h4)
	) name9484 (
		_w13528_,
		_w13530_,
		_w13531_
	);
	LUT2 #(
		.INIT('h1)
	) name9485 (
		_w13519_,
		_w13527_,
		_w13532_
	);
	LUT2 #(
		.INIT('h4)
	) name9486 (
		_w13518_,
		_w13532_,
		_w13533_
	);
	LUT2 #(
		.INIT('h4)
	) name9487 (
		_w13531_,
		_w13533_,
		_w13534_
	);
	LUT2 #(
		.INIT('h1)
	) name9488 (
		_w13517_,
		_w13534_,
		_w13535_
	);
	LUT2 #(
		.INIT('h2)
	) name9489 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w5066_,
		_w13536_
	);
	LUT2 #(
		.INIT('h8)
	) name9490 (
		\bdma_BOVL_reg[9]/NET0131 ,
		_w5066_,
		_w13537_
	);
	LUT2 #(
		.INIT('h1)
	) name9491 (
		_w13536_,
		_w13537_,
		_w13538_
	);
	LUT2 #(
		.INIT('h1)
	) name9492 (
		_w5895_,
		_w13538_,
		_w13539_
	);
	LUT2 #(
		.INIT('h8)
	) name9493 (
		\idma_DOVL_reg[9]/NET0131 ,
		_w5895_,
		_w13540_
	);
	LUT2 #(
		.INIT('h1)
	) name9494 (
		_w13539_,
		_w13540_,
		_w13541_
	);
	LUT2 #(
		.INIT('h8)
	) name9495 (
		_w13535_,
		_w13541_,
		_w13542_
	);
	LUT2 #(
		.INIT('h2)
	) name9496 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w5066_,
		_w13543_
	);
	LUT2 #(
		.INIT('h8)
	) name9497 (
		\bdma_BOVL_reg[11]/NET0131 ,
		_w5066_,
		_w13544_
	);
	LUT2 #(
		.INIT('h1)
	) name9498 (
		_w13543_,
		_w13544_,
		_w13545_
	);
	LUT2 #(
		.INIT('h1)
	) name9499 (
		_w5895_,
		_w13545_,
		_w13546_
	);
	LUT2 #(
		.INIT('h8)
	) name9500 (
		\idma_DOVL_reg[11]/NET0131 ,
		_w5895_,
		_w13547_
	);
	LUT2 #(
		.INIT('h1)
	) name9501 (
		_w13546_,
		_w13547_,
		_w13548_
	);
	LUT2 #(
		.INIT('h2)
	) name9502 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		_w5066_,
		_w13549_
	);
	LUT2 #(
		.INIT('h8)
	) name9503 (
		\bdma_BOVL_reg[10]/NET0131 ,
		_w5066_,
		_w13550_
	);
	LUT2 #(
		.INIT('h1)
	) name9504 (
		_w13549_,
		_w13550_,
		_w13551_
	);
	LUT2 #(
		.INIT('h1)
	) name9505 (
		_w5895_,
		_w13551_,
		_w13552_
	);
	LUT2 #(
		.INIT('h8)
	) name9506 (
		\idma_DOVL_reg[10]/NET0131 ,
		_w5895_,
		_w13553_
	);
	LUT2 #(
		.INIT('h1)
	) name9507 (
		_w13552_,
		_w13553_,
		_w13554_
	);
	LUT2 #(
		.INIT('h8)
	) name9508 (
		_w13548_,
		_w13554_,
		_w13555_
	);
	LUT2 #(
		.INIT('h2)
	) name9509 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		_w5066_,
		_w13556_
	);
	LUT2 #(
		.INIT('h8)
	) name9510 (
		\bdma_BOVL_reg[8]/NET0131 ,
		_w5066_,
		_w13557_
	);
	LUT2 #(
		.INIT('h1)
	) name9511 (
		_w13556_,
		_w13557_,
		_w13558_
	);
	LUT2 #(
		.INIT('h1)
	) name9512 (
		_w5895_,
		_w13558_,
		_w13559_
	);
	LUT2 #(
		.INIT('h8)
	) name9513 (
		\idma_DOVL_reg[8]/NET0131 ,
		_w5895_,
		_w13560_
	);
	LUT2 #(
		.INIT('h1)
	) name9514 (
		_w13559_,
		_w13560_,
		_w13561_
	);
	LUT2 #(
		.INIT('h8)
	) name9515 (
		_w13555_,
		_w13561_,
		_w13562_
	);
	LUT2 #(
		.INIT('h8)
	) name9516 (
		_w13542_,
		_w13562_,
		_w13563_
	);
	LUT2 #(
		.INIT('h1)
	) name9517 (
		_w13384_,
		_w13385_,
		_w13564_
	);
	LUT2 #(
		.INIT('h8)
	) name9518 (
		\memc_Pwrite_C_reg/NET0131 ,
		_w5950_,
		_w13565_
	);
	LUT2 #(
		.INIT('h4)
	) name9519 (
		_w5950_,
		_w13156_,
		_w13566_
	);
	LUT2 #(
		.INIT('h1)
	) name9520 (
		_w13565_,
		_w13566_,
		_w13567_
	);
	LUT2 #(
		.INIT('h8)
	) name9521 (
		_w5066_,
		_w13152_,
		_w13568_
	);
	LUT2 #(
		.INIT('h4)
	) name9522 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_RDcyc_reg/NET0131 ,
		_w13569_
	);
	LUT2 #(
		.INIT('h8)
	) name9523 (
		_w5882_,
		_w13569_,
		_w13570_
	);
	LUT2 #(
		.INIT('h8)
	) name9524 (
		_w5068_,
		_w13570_,
		_w13571_
	);
	LUT2 #(
		.INIT('h1)
	) name9525 (
		_w13568_,
		_w13571_,
		_w13572_
	);
	LUT2 #(
		.INIT('h1)
	) name9526 (
		_w5718_,
		_w13572_,
		_w13573_
	);
	LUT2 #(
		.INIT('h8)
	) name9527 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w6119_,
		_w13574_
	);
	LUT2 #(
		.INIT('h4)
	) name9528 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w13574_,
		_w13575_
	);
	LUT2 #(
		.INIT('h4)
	) name9529 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		\core_c_dec_IR_reg[22]/NET0131 ,
		_w13576_
	);
	LUT2 #(
		.INIT('h8)
	) name9530 (
		_w6026_,
		_w13576_,
		_w13577_
	);
	LUT2 #(
		.INIT('h4)
	) name9531 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w13577_,
		_w13578_
	);
	LUT2 #(
		.INIT('h1)
	) name9532 (
		_w6023_,
		_w13578_,
		_w13579_
	);
	LUT2 #(
		.INIT('h4)
	) name9533 (
		_w13575_,
		_w13579_,
		_w13580_
	);
	LUT2 #(
		.INIT('h2)
	) name9534 (
		_w11742_,
		_w13580_,
		_w13581_
	);
	LUT2 #(
		.INIT('h8)
	) name9535 (
		_w13132_,
		_w13581_,
		_w13582_
	);
	LUT2 #(
		.INIT('h8)
	) name9536 (
		\memc_Pread_E_reg/NET0131 ,
		_w4117_,
		_w13583_
	);
	LUT2 #(
		.INIT('h1)
	) name9537 (
		_w13573_,
		_w13583_,
		_w13584_
	);
	LUT2 #(
		.INIT('h4)
	) name9538 (
		_w13582_,
		_w13584_,
		_w13585_
	);
	LUT2 #(
		.INIT('h8)
	) name9539 (
		_w13564_,
		_w13567_,
		_w13586_
	);
	LUT2 #(
		.INIT('h8)
	) name9540 (
		_w13585_,
		_w13586_,
		_w13587_
	);
	LUT2 #(
		.INIT('h2)
	) name9541 (
		_w13563_,
		_w13587_,
		_w13588_
	);
	LUT2 #(
		.INIT('h2)
	) name9542 (
		_w13555_,
		_w13561_,
		_w13589_
	);
	LUT2 #(
		.INIT('h8)
	) name9543 (
		_w13542_,
		_w13589_,
		_w13590_
	);
	LUT2 #(
		.INIT('h4)
	) name9544 (
		_w13587_,
		_w13590_,
		_w13591_
	);
	LUT2 #(
		.INIT('h2)
	) name9545 (
		_w13535_,
		_w13541_,
		_w13592_
	);
	LUT2 #(
		.INIT('h8)
	) name9546 (
		_w13562_,
		_w13592_,
		_w13593_
	);
	LUT2 #(
		.INIT('h4)
	) name9547 (
		_w13587_,
		_w13593_,
		_w13594_
	);
	LUT2 #(
		.INIT('h8)
	) name9548 (
		_w13589_,
		_w13592_,
		_w13595_
	);
	LUT2 #(
		.INIT('h4)
	) name9549 (
		_w13587_,
		_w13595_,
		_w13596_
	);
	LUT2 #(
		.INIT('h8)
	) name9550 (
		_w13535_,
		_w13548_,
		_w13597_
	);
	LUT2 #(
		.INIT('h4)
	) name9551 (
		_w13554_,
		_w13597_,
		_w13598_
	);
	LUT2 #(
		.INIT('h8)
	) name9552 (
		_w13561_,
		_w13598_,
		_w13599_
	);
	LUT2 #(
		.INIT('h8)
	) name9553 (
		_w13541_,
		_w13599_,
		_w13600_
	);
	LUT2 #(
		.INIT('h4)
	) name9554 (
		_w13587_,
		_w13600_,
		_w13601_
	);
	LUT2 #(
		.INIT('h4)
	) name9555 (
		_w13561_,
		_w13598_,
		_w13602_
	);
	LUT2 #(
		.INIT('h8)
	) name9556 (
		_w13541_,
		_w13602_,
		_w13603_
	);
	LUT2 #(
		.INIT('h4)
	) name9557 (
		_w13587_,
		_w13603_,
		_w13604_
	);
	LUT2 #(
		.INIT('h4)
	) name9558 (
		_w13541_,
		_w13599_,
		_w13605_
	);
	LUT2 #(
		.INIT('h4)
	) name9559 (
		_w13587_,
		_w13605_,
		_w13606_
	);
	LUT2 #(
		.INIT('h4)
	) name9560 (
		_w13541_,
		_w13602_,
		_w13607_
	);
	LUT2 #(
		.INIT('h4)
	) name9561 (
		_w13587_,
		_w13607_,
		_w13608_
	);
	LUT2 #(
		.INIT('h4)
	) name9562 (
		\sport0_cfg_FSi_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w13609_
	);
	LUT2 #(
		.INIT('h8)
	) name9563 (
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w13610_
	);
	LUT2 #(
		.INIT('h2)
	) name9564 (
		\sport0_cfg_FSi_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w13611_
	);
	LUT2 #(
		.INIT('h1)
	) name9565 (
		_w13609_,
		_w13610_,
		_w13612_
	);
	LUT2 #(
		.INIT('h4)
	) name9566 (
		_w13611_,
		_w13612_,
		_w13613_
	);
	LUT2 #(
		.INIT('h4)
	) name9567 (
		\sport1_cfg_FSi_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w13614_
	);
	LUT2 #(
		.INIT('h8)
	) name9568 (
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w13615_
	);
	LUT2 #(
		.INIT('h2)
	) name9569 (
		\sport1_cfg_FSi_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w13616_
	);
	LUT2 #(
		.INIT('h1)
	) name9570 (
		_w13614_,
		_w13615_,
		_w13617_
	);
	LUT2 #(
		.INIT('h4)
	) name9571 (
		_w13616_,
		_w13617_,
		_w13618_
	);
	LUT2 #(
		.INIT('h2)
	) name9572 (
		\sport0_cfg_SCLKi_h_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w13619_
	);
	LUT2 #(
		.INIT('h4)
	) name9573 (
		\sport0_cfg_SCLKi_h_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w13620_
	);
	LUT2 #(
		.INIT('h1)
	) name9574 (
		_w13619_,
		_w13620_,
		_w13621_
	);
	LUT2 #(
		.INIT('h2)
	) name9575 (
		\sport1_cfg_SCLKi_h_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w13622_
	);
	LUT2 #(
		.INIT('h4)
	) name9576 (
		\sport1_cfg_SCLKi_h_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w13623_
	);
	LUT2 #(
		.INIT('h1)
	) name9577 (
		_w13622_,
		_w13623_,
		_w13624_
	);
	LUT2 #(
		.INIT('h1)
	) name9578 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w13625_
	);
	LUT2 #(
		.INIT('h8)
	) name9579 (
		\sport0_txctl_TXSHT_reg[0]/P0001 ,
		_w13625_,
		_w13626_
	);
	LUT2 #(
		.INIT('h2)
	) name9580 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w13627_
	);
	LUT2 #(
		.INIT('h8)
	) name9581 (
		\sport0_txctl_TXSHT_reg[2]/P0001 ,
		_w13627_,
		_w13628_
	);
	LUT2 #(
		.INIT('h1)
	) name9582 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w13626_,
		_w13629_
	);
	LUT2 #(
		.INIT('h4)
	) name9583 (
		_w13628_,
		_w13629_,
		_w13630_
	);
	LUT2 #(
		.INIT('h8)
	) name9584 (
		\sport0_txctl_TXSHT_reg[1]/P0001 ,
		_w13625_,
		_w13631_
	);
	LUT2 #(
		.INIT('h8)
	) name9585 (
		\sport0_txctl_TXSHT_reg[3]/P0001 ,
		_w13627_,
		_w13632_
	);
	LUT2 #(
		.INIT('h2)
	) name9586 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w13631_,
		_w13633_
	);
	LUT2 #(
		.INIT('h4)
	) name9587 (
		_w13632_,
		_w13633_,
		_w13634_
	);
	LUT2 #(
		.INIT('h1)
	) name9588 (
		_w13630_,
		_w13634_,
		_w13635_
	);
	LUT2 #(
		.INIT('h8)
	) name9589 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w13636_
	);
	LUT2 #(
		.INIT('h1)
	) name9590 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[6]/P0001 ,
		_w13637_
	);
	LUT2 #(
		.INIT('h2)
	) name9591 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[7]/P0001 ,
		_w13638_
	);
	LUT2 #(
		.INIT('h2)
	) name9592 (
		_w13636_,
		_w13637_,
		_w13639_
	);
	LUT2 #(
		.INIT('h4)
	) name9593 (
		_w13638_,
		_w13639_,
		_w13640_
	);
	LUT2 #(
		.INIT('h4)
	) name9594 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w13641_
	);
	LUT2 #(
		.INIT('h1)
	) name9595 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[4]/P0001 ,
		_w13642_
	);
	LUT2 #(
		.INIT('h2)
	) name9596 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[5]/P0001 ,
		_w13643_
	);
	LUT2 #(
		.INIT('h2)
	) name9597 (
		_w13641_,
		_w13642_,
		_w13644_
	);
	LUT2 #(
		.INIT('h4)
	) name9598 (
		_w13643_,
		_w13644_,
		_w13645_
	);
	LUT2 #(
		.INIT('h1)
	) name9599 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w13640_,
		_w13646_
	);
	LUT2 #(
		.INIT('h4)
	) name9600 (
		_w13645_,
		_w13646_,
		_w13647_
	);
	LUT2 #(
		.INIT('h4)
	) name9601 (
		_w13635_,
		_w13647_,
		_w13648_
	);
	LUT2 #(
		.INIT('h8)
	) name9602 (
		\sport0_txctl_TXSHT_reg[13]/P0001 ,
		_w13641_,
		_w13649_
	);
	LUT2 #(
		.INIT('h8)
	) name9603 (
		\sport0_txctl_TXSHT_reg[11]/P0001 ,
		_w13627_,
		_w13650_
	);
	LUT2 #(
		.INIT('h8)
	) name9604 (
		\sport0_txctl_TXSHT_reg[9]/P0001 ,
		_w13625_,
		_w13651_
	);
	LUT2 #(
		.INIT('h2)
	) name9605 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w13649_,
		_w13652_
	);
	LUT2 #(
		.INIT('h1)
	) name9606 (
		_w13650_,
		_w13651_,
		_w13653_
	);
	LUT2 #(
		.INIT('h8)
	) name9607 (
		_w13652_,
		_w13653_,
		_w13654_
	);
	LUT2 #(
		.INIT('h8)
	) name9608 (
		\sport0_txctl_TXSHT_reg[8]/P0001 ,
		_w13625_,
		_w13655_
	);
	LUT2 #(
		.INIT('h8)
	) name9609 (
		\sport0_txctl_TXSHT_reg[12]/P0001 ,
		_w13641_,
		_w13656_
	);
	LUT2 #(
		.INIT('h8)
	) name9610 (
		\sport0_txctl_TXSHT_reg[10]/P0001 ,
		_w13627_,
		_w13657_
	);
	LUT2 #(
		.INIT('h1)
	) name9611 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w13655_,
		_w13658_
	);
	LUT2 #(
		.INIT('h1)
	) name9612 (
		_w13656_,
		_w13657_,
		_w13659_
	);
	LUT2 #(
		.INIT('h8)
	) name9613 (
		_w13658_,
		_w13659_,
		_w13660_
	);
	LUT2 #(
		.INIT('h1)
	) name9614 (
		_w13654_,
		_w13660_,
		_w13661_
	);
	LUT2 #(
		.INIT('h1)
	) name9615 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[14]/P0001 ,
		_w13662_
	);
	LUT2 #(
		.INIT('h2)
	) name9616 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport0_txctl_TXSHT_reg[15]/P0001 ,
		_w13663_
	);
	LUT2 #(
		.INIT('h2)
	) name9617 (
		_w13636_,
		_w13662_,
		_w13664_
	);
	LUT2 #(
		.INIT('h4)
	) name9618 (
		_w13663_,
		_w13664_,
		_w13665_
	);
	LUT2 #(
		.INIT('h2)
	) name9619 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w13665_,
		_w13666_
	);
	LUT2 #(
		.INIT('h4)
	) name9620 (
		_w13661_,
		_w13666_,
		_w13667_
	);
	LUT2 #(
		.INIT('h1)
	) name9621 (
		_w13648_,
		_w13667_,
		_w13668_
	);
	LUT2 #(
		.INIT('h1)
	) name9622 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w13668_,
		_w13669_
	);
	LUT2 #(
		.INIT('h2)
	) name9623 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport0_txctl_TXSHT_reg[15]/P0001 ,
		_w13670_
	);
	LUT2 #(
		.INIT('h1)
	) name9624 (
		_w13669_,
		_w13670_,
		_w13671_
	);
	LUT2 #(
		.INIT('h4)
	) name9625 (
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w13671_,
		_w13672_
	);
	LUT2 #(
		.INIT('h2)
	) name9626 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		\sport1_txctl_TXSHT_reg[15]/P0001 ,
		_w13673_
	);
	LUT2 #(
		.INIT('h2)
	) name9627 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w13674_
	);
	LUT2 #(
		.INIT('h2)
	) name9628 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[3]/P0001 ,
		_w13675_
	);
	LUT2 #(
		.INIT('h1)
	) name9629 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[2]/P0001 ,
		_w13676_
	);
	LUT2 #(
		.INIT('h2)
	) name9630 (
		_w13674_,
		_w13675_,
		_w13677_
	);
	LUT2 #(
		.INIT('h4)
	) name9631 (
		_w13676_,
		_w13677_,
		_w13678_
	);
	LUT2 #(
		.INIT('h8)
	) name9632 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w13679_
	);
	LUT2 #(
		.INIT('h1)
	) name9633 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[6]/P0001 ,
		_w13680_
	);
	LUT2 #(
		.INIT('h2)
	) name9634 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[7]/P0001 ,
		_w13681_
	);
	LUT2 #(
		.INIT('h2)
	) name9635 (
		_w13679_,
		_w13680_,
		_w13682_
	);
	LUT2 #(
		.INIT('h4)
	) name9636 (
		_w13681_,
		_w13682_,
		_w13683_
	);
	LUT2 #(
		.INIT('h4)
	) name9637 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w13684_
	);
	LUT2 #(
		.INIT('h1)
	) name9638 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[4]/P0001 ,
		_w13685_
	);
	LUT2 #(
		.INIT('h2)
	) name9639 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[5]/P0001 ,
		_w13686_
	);
	LUT2 #(
		.INIT('h2)
	) name9640 (
		_w13684_,
		_w13685_,
		_w13687_
	);
	LUT2 #(
		.INIT('h4)
	) name9641 (
		_w13686_,
		_w13687_,
		_w13688_
	);
	LUT2 #(
		.INIT('h1)
	) name9642 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w13689_
	);
	LUT2 #(
		.INIT('h1)
	) name9643 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[0]/P0001 ,
		_w13690_
	);
	LUT2 #(
		.INIT('h2)
	) name9644 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[1]/P0001 ,
		_w13691_
	);
	LUT2 #(
		.INIT('h2)
	) name9645 (
		_w13689_,
		_w13690_,
		_w13692_
	);
	LUT2 #(
		.INIT('h4)
	) name9646 (
		_w13691_,
		_w13692_,
		_w13693_
	);
	LUT2 #(
		.INIT('h1)
	) name9647 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w13678_,
		_w13694_
	);
	LUT2 #(
		.INIT('h1)
	) name9648 (
		_w13683_,
		_w13688_,
		_w13695_
	);
	LUT2 #(
		.INIT('h4)
	) name9649 (
		_w13693_,
		_w13695_,
		_w13696_
	);
	LUT2 #(
		.INIT('h8)
	) name9650 (
		_w13694_,
		_w13696_,
		_w13697_
	);
	LUT2 #(
		.INIT('h1)
	) name9651 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[14]/P0001 ,
		_w13698_
	);
	LUT2 #(
		.INIT('h2)
	) name9652 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[15]/P0001 ,
		_w13699_
	);
	LUT2 #(
		.INIT('h2)
	) name9653 (
		_w13679_,
		_w13698_,
		_w13700_
	);
	LUT2 #(
		.INIT('h4)
	) name9654 (
		_w13699_,
		_w13700_,
		_w13701_
	);
	LUT2 #(
		.INIT('h1)
	) name9655 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[8]/P0001 ,
		_w13702_
	);
	LUT2 #(
		.INIT('h2)
	) name9656 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[9]/P0001 ,
		_w13703_
	);
	LUT2 #(
		.INIT('h2)
	) name9657 (
		_w13689_,
		_w13702_,
		_w13704_
	);
	LUT2 #(
		.INIT('h4)
	) name9658 (
		_w13703_,
		_w13704_,
		_w13705_
	);
	LUT2 #(
		.INIT('h1)
	) name9659 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[10]/P0001 ,
		_w13706_
	);
	LUT2 #(
		.INIT('h2)
	) name9660 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[11]/P0001 ,
		_w13707_
	);
	LUT2 #(
		.INIT('h2)
	) name9661 (
		_w13674_,
		_w13706_,
		_w13708_
	);
	LUT2 #(
		.INIT('h4)
	) name9662 (
		_w13707_,
		_w13708_,
		_w13709_
	);
	LUT2 #(
		.INIT('h1)
	) name9663 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[12]/P0001 ,
		_w13710_
	);
	LUT2 #(
		.INIT('h2)
	) name9664 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		\sport1_txctl_TXSHT_reg[13]/P0001 ,
		_w13711_
	);
	LUT2 #(
		.INIT('h2)
	) name9665 (
		_w13684_,
		_w13710_,
		_w13712_
	);
	LUT2 #(
		.INIT('h4)
	) name9666 (
		_w13711_,
		_w13712_,
		_w13713_
	);
	LUT2 #(
		.INIT('h2)
	) name9667 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w13701_,
		_w13714_
	);
	LUT2 #(
		.INIT('h1)
	) name9668 (
		_w13705_,
		_w13709_,
		_w13715_
	);
	LUT2 #(
		.INIT('h4)
	) name9669 (
		_w13713_,
		_w13715_,
		_w13716_
	);
	LUT2 #(
		.INIT('h8)
	) name9670 (
		_w13714_,
		_w13716_,
		_w13717_
	);
	LUT2 #(
		.INIT('h1)
	) name9671 (
		_w13697_,
		_w13717_,
		_w13718_
	);
	LUT2 #(
		.INIT('h1)
	) name9672 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w13718_,
		_w13719_
	);
	LUT2 #(
		.INIT('h1)
	) name9673 (
		_w13673_,
		_w13719_,
		_w13720_
	);
	LUT2 #(
		.INIT('h4)
	) name9674 (
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w13720_,
		_w13721_
	);
	LUT2 #(
		.INIT('h2)
	) name9675 (
		\sport0_cfg_FSi_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w13722_
	);
	LUT2 #(
		.INIT('h4)
	) name9676 (
		\sport0_cfg_FSi_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w13723_
	);
	LUT2 #(
		.INIT('h1)
	) name9677 (
		_w13610_,
		_w13722_,
		_w13724_
	);
	LUT2 #(
		.INIT('h4)
	) name9678 (
		_w13723_,
		_w13724_,
		_w13725_
	);
	LUT2 #(
		.INIT('h2)
	) name9679 (
		\sport1_cfg_FSi_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w13726_
	);
	LUT2 #(
		.INIT('h4)
	) name9680 (
		\sport1_cfg_FSi_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w13727_
	);
	LUT2 #(
		.INIT('h1)
	) name9681 (
		_w13615_,
		_w13726_,
		_w13728_
	);
	LUT2 #(
		.INIT('h4)
	) name9682 (
		_w13727_,
		_w13728_,
		_w13729_
	);
	LUT2 #(
		.INIT('h4)
	) name9683 (
		\bdma_BM_cyc_reg/P0001 ,
		\emc_WRn_h_reg/P0001 ,
		_w13730_
	);
	LUT2 #(
		.INIT('h8)
	) name9684 (
		\bdma_BM_cyc_reg/P0001 ,
		\bdma_BWRn_reg/NET0131 ,
		_w13731_
	);
	LUT2 #(
		.INIT('h1)
	) name9685 (
		_w13730_,
		_w13731_,
		_w13732_
	);
	LUT2 #(
		.INIT('h1)
	) name9686 (
		T_BMODE_pad,
		T_MMAP_pad,
		_w13733_
	);
	LUT2 #(
		.INIT('h8)
	) name9687 (
		\bdma_RST_pin_reg/P0001 ,
		_w13733_,
		_w13734_
	);
	LUT2 #(
		.INIT('h1)
	) name9688 (
		\bdma_BWCOUNT_reg[3]/NET0131 ,
		\bdma_BWCOUNT_reg[4]/NET0131 ,
		_w13735_
	);
	LUT2 #(
		.INIT('h1)
	) name9689 (
		\bdma_BWCOUNT_reg[1]/NET0131 ,
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		_w13736_
	);
	LUT2 #(
		.INIT('h4)
	) name9690 (
		\bdma_BWCOUNT_reg[6]/NET0131 ,
		_w13736_,
		_w13737_
	);
	LUT2 #(
		.INIT('h8)
	) name9691 (
		_w13735_,
		_w13737_,
		_w13738_
	);
	LUT2 #(
		.INIT('h8)
	) name9692 (
		_w10716_,
		_w13738_,
		_w13739_
	);
	LUT2 #(
		.INIT('h1)
	) name9693 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		_w13740_
	);
	LUT2 #(
		.INIT('h1)
	) name9694 (
		\bdma_BWCOUNT_reg[12]/NET0131 ,
		\bdma_BWCOUNT_reg[13]/NET0131 ,
		_w13741_
	);
	LUT2 #(
		.INIT('h1)
	) name9695 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		_w13742_
	);
	LUT2 #(
		.INIT('h4)
	) name9696 (
		\bdma_BWCOUNT_reg[9]/NET0131 ,
		_w13742_,
		_w13743_
	);
	LUT2 #(
		.INIT('h8)
	) name9697 (
		_w13740_,
		_w13741_,
		_w13744_
	);
	LUT2 #(
		.INIT('h8)
	) name9698 (
		_w13743_,
		_w13744_,
		_w13745_
	);
	LUT2 #(
		.INIT('h8)
	) name9699 (
		_w13739_,
		_w13745_,
		_w13746_
	);
	LUT2 #(
		.INIT('h1)
	) name9700 (
		_w5733_,
		_w13147_,
		_w13747_
	);
	LUT2 #(
		.INIT('h1)
	) name9701 (
		_w5561_,
		_w5563_,
		_w13748_
	);
	LUT2 #(
		.INIT('h8)
	) name9702 (
		_w5560_,
		_w5597_,
		_w13749_
	);
	LUT2 #(
		.INIT('h8)
	) name9703 (
		_w5587_,
		_w13749_,
		_w13750_
	);
	LUT2 #(
		.INIT('h4)
	) name9704 (
		_w13748_,
		_w13750_,
		_w13751_
	);
	LUT2 #(
		.INIT('h4)
	) name9705 (
		_w13747_,
		_w13751_,
		_w13752_
	);
	LUT2 #(
		.INIT('h8)
	) name9706 (
		_w6915_,
		_w13751_,
		_w13753_
	);
	LUT2 #(
		.INIT('h4)
	) name9707 (
		_w6914_,
		_w13753_,
		_w13754_
	);
	LUT2 #(
		.INIT('h1)
	) name9708 (
		_w13752_,
		_w13754_,
		_w13755_
	);
	LUT2 #(
		.INIT('h8)
	) name9709 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w13746_,
		_w13756_
	);
	LUT2 #(
		.INIT('h4)
	) name9710 (
		_w13755_,
		_w13756_,
		_w13757_
	);
	LUT2 #(
		.INIT('h1)
	) name9711 (
		_w4063_,
		_w13757_,
		_w13758_
	);
	LUT2 #(
		.INIT('h1)
	) name9712 (
		_w13734_,
		_w13758_,
		_w13759_
	);
	LUT2 #(
		.INIT('h2)
	) name9713 (
		\memc_Dwrite_E_reg/NET0131 ,
		_w5950_,
		_w13760_
	);
	LUT2 #(
		.INIT('h4)
	) name9714 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w13760_,
		_w13761_
	);
	LUT2 #(
		.INIT('h8)
	) name9715 (
		_w7285_,
		_w13761_,
		_w13762_
	);
	LUT2 #(
		.INIT('h8)
	) name9716 (
		_w7284_,
		_w13762_,
		_w13763_
	);
	LUT2 #(
		.INIT('h1)
	) name9717 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w13755_,
		_w13764_
	);
	LUT2 #(
		.INIT('h4)
	) name9718 (
		\bdma_BWCOUNT_reg[1]/NET0131 ,
		_w13764_,
		_w13765_
	);
	LUT2 #(
		.INIT('h4)
	) name9719 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		_w13765_,
		_w13766_
	);
	LUT2 #(
		.INIT('h8)
	) name9720 (
		_w13735_,
		_w13766_,
		_w13767_
	);
	LUT2 #(
		.INIT('h1)
	) name9721 (
		_w10716_,
		_w13767_,
		_w13768_
	);
	LUT2 #(
		.INIT('h8)
	) name9722 (
		_w10716_,
		_w13767_,
		_w13769_
	);
	LUT2 #(
		.INIT('h1)
	) name9723 (
		_w13763_,
		_w13768_,
		_w13770_
	);
	LUT2 #(
		.INIT('h4)
	) name9724 (
		_w13769_,
		_w13770_,
		_w13771_
	);
	LUT2 #(
		.INIT('h4)
	) name9725 (
		_w10911_,
		_w13763_,
		_w13772_
	);
	LUT2 #(
		.INIT('h1)
	) name9726 (
		_w13771_,
		_w13772_,
		_w13773_
	);
	LUT2 #(
		.INIT('h1)
	) name9727 (
		_w13734_,
		_w13773_,
		_w13774_
	);
	LUT2 #(
		.INIT('h8)
	) name9728 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w13775_
	);
	LUT2 #(
		.INIT('h4)
	) name9729 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w13775_,
		_w13776_
	);
	LUT2 #(
		.INIT('h8)
	) name9730 (
		\core_c_dec_MTCNTR_Eg_reg/P0001 ,
		\core_c_psq_CNTRval_reg/NET0131 ,
		_w13777_
	);
	LUT2 #(
		.INIT('h4)
	) name9731 (
		_w5950_,
		_w13777_,
		_w13778_
	);
	LUT2 #(
		.INIT('h4)
	) name9732 (
		_w13776_,
		_w13778_,
		_w13779_
	);
	LUT2 #(
		.INIT('h8)
	) name9733 (
		_w13775_,
		_w13779_,
		_w13780_
	);
	LUT2 #(
		.INIT('h2)
	) name9734 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001 ,
		_w13780_,
		_w13781_
	);
	LUT2 #(
		.INIT('h8)
	) name9735 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w13780_,
		_w13782_
	);
	LUT2 #(
		.INIT('h1)
	) name9736 (
		_w13781_,
		_w13782_,
		_w13783_
	);
	LUT2 #(
		.INIT('h1)
	) name9737 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w13784_
	);
	LUT2 #(
		.INIT('h8)
	) name9738 (
		_w13778_,
		_w13784_,
		_w13785_
	);
	LUT2 #(
		.INIT('h2)
	) name9739 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001 ,
		_w13785_,
		_w13786_
	);
	LUT2 #(
		.INIT('h8)
	) name9740 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w13785_,
		_w13787_
	);
	LUT2 #(
		.INIT('h1)
	) name9741 (
		_w13786_,
		_w13787_,
		_w13788_
	);
	LUT2 #(
		.INIT('h2)
	) name9742 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w13789_
	);
	LUT2 #(
		.INIT('h8)
	) name9743 (
		_w13778_,
		_w13789_,
		_w13790_
	);
	LUT2 #(
		.INIT('h2)
	) name9744 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001 ,
		_w13790_,
		_w13791_
	);
	LUT2 #(
		.INIT('h8)
	) name9745 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w13790_,
		_w13792_
	);
	LUT2 #(
		.INIT('h1)
	) name9746 (
		_w13791_,
		_w13792_,
		_w13793_
	);
	LUT2 #(
		.INIT('h4)
	) name9747 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		\core_c_psq_cntstk_ptr_reg[1]/NET0131 ,
		_w13794_
	);
	LUT2 #(
		.INIT('h8)
	) name9748 (
		_w13778_,
		_w13794_,
		_w13795_
	);
	LUT2 #(
		.INIT('h2)
	) name9749 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001 ,
		_w13795_,
		_w13796_
	);
	LUT2 #(
		.INIT('h8)
	) name9750 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w13795_,
		_w13797_
	);
	LUT2 #(
		.INIT('h1)
	) name9751 (
		_w13796_,
		_w13797_,
		_w13798_
	);
	LUT2 #(
		.INIT('h1)
	) name9752 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w13799_
	);
	LUT2 #(
		.INIT('h4)
	) name9753 (
		\core_c_dec_updAF_E_reg/P0001 ,
		_w13799_,
		_w13800_
	);
	LUT2 #(
		.INIT('h1)
	) name9754 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w5950_,
		_w13801_
	);
	LUT2 #(
		.INIT('h8)
	) name9755 (
		\core_c_dec_Usecond_E_reg/P0001 ,
		_w4184_,
		_w13802_
	);
	LUT2 #(
		.INIT('h1)
	) name9756 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w13802_,
		_w13803_
	);
	LUT2 #(
		.INIT('h8)
	) name9757 (
		_w13801_,
		_w13803_,
		_w13804_
	);
	LUT2 #(
		.INIT('h4)
	) name9758 (
		_w13800_,
		_w13804_,
		_w13805_
	);
	LUT2 #(
		.INIT('h1)
	) name9759 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w13799_,
		_w13806_
	);
	LUT2 #(
		.INIT('h8)
	) name9760 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		_w13807_
	);
	LUT2 #(
		.INIT('h8)
	) name9761 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w13808_
	);
	LUT2 #(
		.INIT('h4)
	) name9762 (
		_w13807_,
		_w13808_,
		_w13809_
	);
	LUT2 #(
		.INIT('h8)
	) name9763 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w13807_,
		_w13810_
	);
	LUT2 #(
		.INIT('h8)
	) name9764 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		_w13810_,
		_w13811_
	);
	LUT2 #(
		.INIT('h2)
	) name9765 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w13812_
	);
	LUT2 #(
		.INIT('h8)
	) name9766 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w13812_,
		_w13813_
	);
	LUT2 #(
		.INIT('h4)
	) name9767 (
		_w7206_,
		_w13813_,
		_w13814_
	);
	LUT2 #(
		.INIT('h1)
	) name9768 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w13815_
	);
	LUT2 #(
		.INIT('h8)
	) name9769 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w13815_,
		_w13816_
	);
	LUT2 #(
		.INIT('h4)
	) name9770 (
		_w11983_,
		_w13816_,
		_w13817_
	);
	LUT2 #(
		.INIT('h8)
	) name9771 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w13818_
	);
	LUT2 #(
		.INIT('h4)
	) name9772 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w13818_,
		_w13819_
	);
	LUT2 #(
		.INIT('h4)
	) name9773 (
		_w12024_,
		_w13819_,
		_w13820_
	);
	LUT2 #(
		.INIT('h4)
	) name9774 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w13812_,
		_w13821_
	);
	LUT2 #(
		.INIT('h4)
	) name9775 (
		_w12028_,
		_w13821_,
		_w13822_
	);
	LUT2 #(
		.INIT('h8)
	) name9776 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w13823_
	);
	LUT2 #(
		.INIT('h4)
	) name9777 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11992_,
		_w13824_
	);
	LUT2 #(
		.INIT('h8)
	) name9778 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w12000_,
		_w13825_
	);
	LUT2 #(
		.INIT('h2)
	) name9779 (
		_w13823_,
		_w13824_,
		_w13826_
	);
	LUT2 #(
		.INIT('h4)
	) name9780 (
		_w13825_,
		_w13826_,
		_w13827_
	);
	LUT2 #(
		.INIT('h1)
	) name9781 (
		_w13814_,
		_w13817_,
		_w13828_
	);
	LUT2 #(
		.INIT('h1)
	) name9782 (
		_w13820_,
		_w13822_,
		_w13829_
	);
	LUT2 #(
		.INIT('h8)
	) name9783 (
		_w13828_,
		_w13829_,
		_w13830_
	);
	LUT2 #(
		.INIT('h4)
	) name9784 (
		_w13827_,
		_w13830_,
		_w13831_
	);
	LUT2 #(
		.INIT('h1)
	) name9785 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w13832_
	);
	LUT2 #(
		.INIT('h4)
	) name9786 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11967_,
		_w13833_
	);
	LUT2 #(
		.INIT('h8)
	) name9787 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11971_,
		_w13834_
	);
	LUT2 #(
		.INIT('h2)
	) name9788 (
		_w13832_,
		_w13833_,
		_w13835_
	);
	LUT2 #(
		.INIT('h4)
	) name9789 (
		_w13834_,
		_w13835_,
		_w13836_
	);
	LUT2 #(
		.INIT('h2)
	) name9790 (
		_w13831_,
		_w13836_,
		_w13837_
	);
	LUT2 #(
		.INIT('h2)
	) name9791 (
		_w13811_,
		_w13837_,
		_w13838_
	);
	LUT2 #(
		.INIT('h1)
	) name9792 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		\core_c_dec_DIVQ_E_reg/P0001 ,
		_w13839_
	);
	LUT2 #(
		.INIT('h4)
	) name9793 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w13839_,
		_w13840_
	);
	LUT2 #(
		.INIT('h2)
	) name9794 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w13841_
	);
	LUT2 #(
		.INIT('h1)
	) name9795 (
		_w13840_,
		_w13841_,
		_w13842_
	);
	LUT2 #(
		.INIT('h1)
	) name9796 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		_w13843_
	);
	LUT2 #(
		.INIT('h8)
	) name9797 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		_w13843_,
		_w13844_
	);
	LUT2 #(
		.INIT('h4)
	) name9798 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w13845_
	);
	LUT2 #(
		.INIT('h4)
	) name9799 (
		_w13844_,
		_w13845_,
		_w13846_
	);
	LUT2 #(
		.INIT('h2)
	) name9800 (
		_w13842_,
		_w13846_,
		_w13847_
	);
	LUT2 #(
		.INIT('h4)
	) name9801 (
		_w13838_,
		_w13847_,
		_w13848_
	);
	LUT2 #(
		.INIT('h1)
	) name9802 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		_w13849_
	);
	LUT2 #(
		.INIT('h4)
	) name9803 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		_w13849_,
		_w13850_
	);
	LUT2 #(
		.INIT('h2)
	) name9804 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w13850_,
		_w13851_
	);
	LUT2 #(
		.INIT('h1)
	) name9805 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		_w13851_,
		_w13852_
	);
	LUT2 #(
		.INIT('h1)
	) name9806 (
		_w13840_,
		_w13852_,
		_w13853_
	);
	LUT2 #(
		.INIT('h4)
	) name9807 (
		_w10191_,
		_w13816_,
		_w13854_
	);
	LUT2 #(
		.INIT('h4)
	) name9808 (
		_w10112_,
		_w13819_,
		_w13855_
	);
	LUT2 #(
		.INIT('h4)
	) name9809 (
		_w10096_,
		_w13821_,
		_w13856_
	);
	LUT2 #(
		.INIT('h4)
	) name9810 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10218_,
		_w13857_
	);
	LUT2 #(
		.INIT('h8)
	) name9811 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10226_,
		_w13858_
	);
	LUT2 #(
		.INIT('h2)
	) name9812 (
		_w13823_,
		_w13857_,
		_w13859_
	);
	LUT2 #(
		.INIT('h4)
	) name9813 (
		_w13858_,
		_w13859_,
		_w13860_
	);
	LUT2 #(
		.INIT('h1)
	) name9814 (
		_w13814_,
		_w13854_,
		_w13861_
	);
	LUT2 #(
		.INIT('h1)
	) name9815 (
		_w13855_,
		_w13856_,
		_w13862_
	);
	LUT2 #(
		.INIT('h8)
	) name9816 (
		_w13861_,
		_w13862_,
		_w13863_
	);
	LUT2 #(
		.INIT('h4)
	) name9817 (
		_w13860_,
		_w13863_,
		_w13864_
	);
	LUT2 #(
		.INIT('h4)
	) name9818 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10187_,
		_w13865_
	);
	LUT2 #(
		.INIT('h8)
	) name9819 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10179_,
		_w13866_
	);
	LUT2 #(
		.INIT('h2)
	) name9820 (
		_w13832_,
		_w13865_,
		_w13867_
	);
	LUT2 #(
		.INIT('h4)
	) name9821 (
		_w13866_,
		_w13867_,
		_w13868_
	);
	LUT2 #(
		.INIT('h2)
	) name9822 (
		_w13864_,
		_w13868_,
		_w13869_
	);
	LUT2 #(
		.INIT('h2)
	) name9823 (
		_w13853_,
		_w13869_,
		_w13870_
	);
	LUT2 #(
		.INIT('h2)
	) name9824 (
		_w13848_,
		_w13870_,
		_w13871_
	);
	LUT2 #(
		.INIT('h4)
	) name9825 (
		_w13848_,
		_w13870_,
		_w13872_
	);
	LUT2 #(
		.INIT('h1)
	) name9826 (
		_w13871_,
		_w13872_,
		_w13873_
	);
	LUT2 #(
		.INIT('h2)
	) name9827 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[2]/NET0131 ,
		\core_eu_ea_alu_ea_dec_AMF_E_reg[3]/NET0131 ,
		_w13874_
	);
	LUT2 #(
		.INIT('h1)
	) name9828 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w13875_
	);
	LUT2 #(
		.INIT('h1)
	) name9829 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w13876_
	);
	LUT2 #(
		.INIT('h8)
	) name9830 (
		_w13875_,
		_w13876_,
		_w13877_
	);
	LUT2 #(
		.INIT('h2)
	) name9831 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w13877_,
		_w13878_
	);
	LUT2 #(
		.INIT('h4)
	) name9832 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001 ,
		_w13878_,
		_w13879_
	);
	LUT2 #(
		.INIT('h1)
	) name9833 (
		_w13810_,
		_w13840_,
		_w13880_
	);
	LUT2 #(
		.INIT('h2)
	) name9834 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w13881_
	);
	LUT2 #(
		.INIT('h4)
	) name9835 (
		_w10175_,
		_w13881_,
		_w13882_
	);
	LUT2 #(
		.INIT('h4)
	) name9836 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w10183_,
		_w13883_
	);
	LUT2 #(
		.INIT('h1)
	) name9837 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001 ,
		_w13884_
	);
	LUT2 #(
		.INIT('h2)
	) name9838 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001 ,
		_w13885_
	);
	LUT2 #(
		.INIT('h1)
	) name9839 (
		_w13884_,
		_w13885_,
		_w13886_
	);
	LUT2 #(
		.INIT('h2)
	) name9840 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w13886_,
		_w13887_
	);
	LUT2 #(
		.INIT('h1)
	) name9841 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w13883_,
		_w13888_
	);
	LUT2 #(
		.INIT('h4)
	) name9842 (
		_w13887_,
		_w13888_,
		_w13889_
	);
	LUT2 #(
		.INIT('h1)
	) name9843 (
		_w13878_,
		_w13882_,
		_w13890_
	);
	LUT2 #(
		.INIT('h4)
	) name9844 (
		_w13889_,
		_w13890_,
		_w13891_
	);
	LUT2 #(
		.INIT('h4)
	) name9845 (
		_w13879_,
		_w13880_,
		_w13892_
	);
	LUT2 #(
		.INIT('h4)
	) name9846 (
		_w13891_,
		_w13892_,
		_w13893_
	);
	LUT2 #(
		.INIT('h4)
	) name9847 (
		_w13874_,
		_w13893_,
		_w13894_
	);
	LUT2 #(
		.INIT('h1)
	) name9848 (
		_w13840_,
		_w13874_,
		_w13895_
	);
	LUT2 #(
		.INIT('h1)
	) name9849 (
		_w13893_,
		_w13895_,
		_w13896_
	);
	LUT2 #(
		.INIT('h1)
	) name9850 (
		_w13894_,
		_w13896_,
		_w13897_
	);
	LUT2 #(
		.INIT('h4)
	) name9851 (
		_w13873_,
		_w13897_,
		_w13898_
	);
	LUT2 #(
		.INIT('h4)
	) name9852 (
		_w10461_,
		_w13816_,
		_w13899_
	);
	LUT2 #(
		.INIT('h4)
	) name9853 (
		_w10534_,
		_w13819_,
		_w13900_
	);
	LUT2 #(
		.INIT('h4)
	) name9854 (
		_w10538_,
		_w13821_,
		_w13901_
	);
	LUT2 #(
		.INIT('h4)
	) name9855 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10567_,
		_w13902_
	);
	LUT2 #(
		.INIT('h8)
	) name9856 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10575_,
		_w13903_
	);
	LUT2 #(
		.INIT('h2)
	) name9857 (
		_w13823_,
		_w13902_,
		_w13904_
	);
	LUT2 #(
		.INIT('h4)
	) name9858 (
		_w13903_,
		_w13904_,
		_w13905_
	);
	LUT2 #(
		.INIT('h1)
	) name9859 (
		_w13814_,
		_w13899_,
		_w13906_
	);
	LUT2 #(
		.INIT('h1)
	) name9860 (
		_w13900_,
		_w13901_,
		_w13907_
	);
	LUT2 #(
		.INIT('h8)
	) name9861 (
		_w13906_,
		_w13907_,
		_w13908_
	);
	LUT2 #(
		.INIT('h4)
	) name9862 (
		_w13905_,
		_w13908_,
		_w13909_
	);
	LUT2 #(
		.INIT('h4)
	) name9863 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10449_,
		_w13910_
	);
	LUT2 #(
		.INIT('h8)
	) name9864 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10457_,
		_w13911_
	);
	LUT2 #(
		.INIT('h2)
	) name9865 (
		_w13832_,
		_w13910_,
		_w13912_
	);
	LUT2 #(
		.INIT('h4)
	) name9866 (
		_w13911_,
		_w13912_,
		_w13913_
	);
	LUT2 #(
		.INIT('h2)
	) name9867 (
		_w13909_,
		_w13913_,
		_w13914_
	);
	LUT2 #(
		.INIT('h2)
	) name9868 (
		_w13853_,
		_w13914_,
		_w13915_
	);
	LUT2 #(
		.INIT('h2)
	) name9869 (
		_w13848_,
		_w13915_,
		_w13916_
	);
	LUT2 #(
		.INIT('h4)
	) name9870 (
		_w13848_,
		_w13915_,
		_w13917_
	);
	LUT2 #(
		.INIT('h1)
	) name9871 (
		_w13916_,
		_w13917_,
		_w13918_
	);
	LUT2 #(
		.INIT('h4)
	) name9872 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001 ,
		_w13878_,
		_w13919_
	);
	LUT2 #(
		.INIT('h4)
	) name9873 (
		_w10445_,
		_w13881_,
		_w13920_
	);
	LUT2 #(
		.INIT('h4)
	) name9874 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w10453_,
		_w13921_
	);
	LUT2 #(
		.INIT('h1)
	) name9875 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001 ,
		_w13922_
	);
	LUT2 #(
		.INIT('h2)
	) name9876 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001 ,
		_w13923_
	);
	LUT2 #(
		.INIT('h1)
	) name9877 (
		_w13922_,
		_w13923_,
		_w13924_
	);
	LUT2 #(
		.INIT('h2)
	) name9878 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w13924_,
		_w13925_
	);
	LUT2 #(
		.INIT('h1)
	) name9879 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w13921_,
		_w13926_
	);
	LUT2 #(
		.INIT('h4)
	) name9880 (
		_w13925_,
		_w13926_,
		_w13927_
	);
	LUT2 #(
		.INIT('h1)
	) name9881 (
		_w13878_,
		_w13920_,
		_w13928_
	);
	LUT2 #(
		.INIT('h4)
	) name9882 (
		_w13927_,
		_w13928_,
		_w13929_
	);
	LUT2 #(
		.INIT('h2)
	) name9883 (
		_w13880_,
		_w13919_,
		_w13930_
	);
	LUT2 #(
		.INIT('h4)
	) name9884 (
		_w13929_,
		_w13930_,
		_w13931_
	);
	LUT2 #(
		.INIT('h2)
	) name9885 (
		_w13895_,
		_w13931_,
		_w13932_
	);
	LUT2 #(
		.INIT('h8)
	) name9886 (
		_w13874_,
		_w13931_,
		_w13933_
	);
	LUT2 #(
		.INIT('h1)
	) name9887 (
		_w13932_,
		_w13933_,
		_w13934_
	);
	LUT2 #(
		.INIT('h1)
	) name9888 (
		_w13918_,
		_w13934_,
		_w13935_
	);
	LUT2 #(
		.INIT('h4)
	) name9889 (
		_w11192_,
		_w13819_,
		_w13936_
	);
	LUT2 #(
		.INIT('h4)
	) name9890 (
		_w11196_,
		_w13821_,
		_w13937_
	);
	LUT2 #(
		.INIT('h4)
	) name9891 (
		_w11062_,
		_w13816_,
		_w13938_
	);
	LUT2 #(
		.INIT('h4)
	) name9892 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11231_,
		_w13939_
	);
	LUT2 #(
		.INIT('h8)
	) name9893 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11239_,
		_w13940_
	);
	LUT2 #(
		.INIT('h2)
	) name9894 (
		_w13823_,
		_w13939_,
		_w13941_
	);
	LUT2 #(
		.INIT('h4)
	) name9895 (
		_w13940_,
		_w13941_,
		_w13942_
	);
	LUT2 #(
		.INIT('h1)
	) name9896 (
		_w13814_,
		_w13936_,
		_w13943_
	);
	LUT2 #(
		.INIT('h1)
	) name9897 (
		_w13937_,
		_w13938_,
		_w13944_
	);
	LUT2 #(
		.INIT('h8)
	) name9898 (
		_w13943_,
		_w13944_,
		_w13945_
	);
	LUT2 #(
		.INIT('h4)
	) name9899 (
		_w13942_,
		_w13945_,
		_w13946_
	);
	LUT2 #(
		.INIT('h4)
	) name9900 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11070_,
		_w13947_
	);
	LUT2 #(
		.INIT('h8)
	) name9901 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11066_,
		_w13948_
	);
	LUT2 #(
		.INIT('h2)
	) name9902 (
		_w13832_,
		_w13947_,
		_w13949_
	);
	LUT2 #(
		.INIT('h4)
	) name9903 (
		_w13948_,
		_w13949_,
		_w13950_
	);
	LUT2 #(
		.INIT('h2)
	) name9904 (
		_w13946_,
		_w13950_,
		_w13951_
	);
	LUT2 #(
		.INIT('h2)
	) name9905 (
		_w13853_,
		_w13951_,
		_w13952_
	);
	LUT2 #(
		.INIT('h4)
	) name9906 (
		_w13848_,
		_w13952_,
		_w13953_
	);
	LUT2 #(
		.INIT('h2)
	) name9907 (
		_w13848_,
		_w13952_,
		_w13954_
	);
	LUT2 #(
		.INIT('h1)
	) name9908 (
		_w13953_,
		_w13954_,
		_w13955_
	);
	LUT2 #(
		.INIT('h4)
	) name9909 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001 ,
		_w13878_,
		_w13956_
	);
	LUT2 #(
		.INIT('h4)
	) name9910 (
		_w11058_,
		_w13881_,
		_w13957_
	);
	LUT2 #(
		.INIT('h4)
	) name9911 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11054_,
		_w13958_
	);
	LUT2 #(
		.INIT('h1)
	) name9912 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001 ,
		_w13959_
	);
	LUT2 #(
		.INIT('h2)
	) name9913 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001 ,
		_w13960_
	);
	LUT2 #(
		.INIT('h1)
	) name9914 (
		_w13959_,
		_w13960_,
		_w13961_
	);
	LUT2 #(
		.INIT('h2)
	) name9915 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w13961_,
		_w13962_
	);
	LUT2 #(
		.INIT('h1)
	) name9916 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w13958_,
		_w13963_
	);
	LUT2 #(
		.INIT('h4)
	) name9917 (
		_w13962_,
		_w13963_,
		_w13964_
	);
	LUT2 #(
		.INIT('h1)
	) name9918 (
		_w13878_,
		_w13957_,
		_w13965_
	);
	LUT2 #(
		.INIT('h4)
	) name9919 (
		_w13964_,
		_w13965_,
		_w13966_
	);
	LUT2 #(
		.INIT('h2)
	) name9920 (
		_w13880_,
		_w13956_,
		_w13967_
	);
	LUT2 #(
		.INIT('h4)
	) name9921 (
		_w13966_,
		_w13967_,
		_w13968_
	);
	LUT2 #(
		.INIT('h2)
	) name9922 (
		_w13895_,
		_w13968_,
		_w13969_
	);
	LUT2 #(
		.INIT('h8)
	) name9923 (
		_w13874_,
		_w13968_,
		_w13970_
	);
	LUT2 #(
		.INIT('h1)
	) name9924 (
		_w13969_,
		_w13970_,
		_w13971_
	);
	LUT2 #(
		.INIT('h1)
	) name9925 (
		_w13955_,
		_w13971_,
		_w13972_
	);
	LUT2 #(
		.INIT('h4)
	) name9926 (
		_w11424_,
		_w13813_,
		_w13973_
	);
	LUT2 #(
		.INIT('h4)
	) name9927 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11315_,
		_w13974_
	);
	LUT2 #(
		.INIT('h8)
	) name9928 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11311_,
		_w13975_
	);
	LUT2 #(
		.INIT('h2)
	) name9929 (
		_w13823_,
		_w13974_,
		_w13976_
	);
	LUT2 #(
		.INIT('h4)
	) name9930 (
		_w13975_,
		_w13976_,
		_w13977_
	);
	LUT2 #(
		.INIT('h4)
	) name9931 (
		_w11341_,
		_w13816_,
		_w13978_
	);
	LUT2 #(
		.INIT('h4)
	) name9932 (
		_w11444_,
		_w13819_,
		_w13979_
	);
	LUT2 #(
		.INIT('h4)
	) name9933 (
		_w11448_,
		_w13821_,
		_w13980_
	);
	LUT2 #(
		.INIT('h1)
	) name9934 (
		_w13973_,
		_w13978_,
		_w13981_
	);
	LUT2 #(
		.INIT('h1)
	) name9935 (
		_w13979_,
		_w13980_,
		_w13982_
	);
	LUT2 #(
		.INIT('h8)
	) name9936 (
		_w13981_,
		_w13982_,
		_w13983_
	);
	LUT2 #(
		.INIT('h4)
	) name9937 (
		_w13977_,
		_w13983_,
		_w13984_
	);
	LUT2 #(
		.INIT('h4)
	) name9938 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11325_,
		_w13985_
	);
	LUT2 #(
		.INIT('h8)
	) name9939 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11337_,
		_w13986_
	);
	LUT2 #(
		.INIT('h2)
	) name9940 (
		_w13832_,
		_w13985_,
		_w13987_
	);
	LUT2 #(
		.INIT('h4)
	) name9941 (
		_w13986_,
		_w13987_,
		_w13988_
	);
	LUT2 #(
		.INIT('h2)
	) name9942 (
		_w13984_,
		_w13988_,
		_w13989_
	);
	LUT2 #(
		.INIT('h2)
	) name9943 (
		_w13853_,
		_w13989_,
		_w13990_
	);
	LUT2 #(
		.INIT('h2)
	) name9944 (
		_w13848_,
		_w13990_,
		_w13991_
	);
	LUT2 #(
		.INIT('h4)
	) name9945 (
		_w13848_,
		_w13990_,
		_w13992_
	);
	LUT2 #(
		.INIT('h1)
	) name9946 (
		_w13991_,
		_w13992_,
		_w13993_
	);
	LUT2 #(
		.INIT('h4)
	) name9947 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001 ,
		_w13878_,
		_w13994_
	);
	LUT2 #(
		.INIT('h4)
	) name9948 (
		_w11333_,
		_w13881_,
		_w13995_
	);
	LUT2 #(
		.INIT('h4)
	) name9949 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11329_,
		_w13996_
	);
	LUT2 #(
		.INIT('h1)
	) name9950 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001 ,
		_w13997_
	);
	LUT2 #(
		.INIT('h2)
	) name9951 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001 ,
		_w13998_
	);
	LUT2 #(
		.INIT('h1)
	) name9952 (
		_w13997_,
		_w13998_,
		_w13999_
	);
	LUT2 #(
		.INIT('h2)
	) name9953 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w13999_,
		_w14000_
	);
	LUT2 #(
		.INIT('h1)
	) name9954 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w13996_,
		_w14001_
	);
	LUT2 #(
		.INIT('h4)
	) name9955 (
		_w14000_,
		_w14001_,
		_w14002_
	);
	LUT2 #(
		.INIT('h1)
	) name9956 (
		_w13878_,
		_w13995_,
		_w14003_
	);
	LUT2 #(
		.INIT('h4)
	) name9957 (
		_w14002_,
		_w14003_,
		_w14004_
	);
	LUT2 #(
		.INIT('h2)
	) name9958 (
		_w13880_,
		_w13994_,
		_w14005_
	);
	LUT2 #(
		.INIT('h4)
	) name9959 (
		_w14004_,
		_w14005_,
		_w14006_
	);
	LUT2 #(
		.INIT('h2)
	) name9960 (
		_w13895_,
		_w14006_,
		_w14007_
	);
	LUT2 #(
		.INIT('h8)
	) name9961 (
		_w13874_,
		_w14006_,
		_w14008_
	);
	LUT2 #(
		.INIT('h1)
	) name9962 (
		_w14007_,
		_w14008_,
		_w14009_
	);
	LUT2 #(
		.INIT('h1)
	) name9963 (
		_w13993_,
		_w14009_,
		_w14010_
	);
	LUT2 #(
		.INIT('h4)
	) name9964 (
		_w10878_,
		_w13819_,
		_w14011_
	);
	LUT2 #(
		.INIT('h4)
	) name9965 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10801_,
		_w14012_
	);
	LUT2 #(
		.INIT('h8)
	) name9966 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10797_,
		_w14013_
	);
	LUT2 #(
		.INIT('h2)
	) name9967 (
		_w13823_,
		_w14012_,
		_w14014_
	);
	LUT2 #(
		.INIT('h4)
	) name9968 (
		_w14013_,
		_w14014_,
		_w14015_
	);
	LUT2 #(
		.INIT('h4)
	) name9969 (
		_w10858_,
		_w13821_,
		_w14016_
	);
	LUT2 #(
		.INIT('h4)
	) name9970 (
		_w10882_,
		_w13813_,
		_w14017_
	);
	LUT2 #(
		.INIT('h4)
	) name9971 (
		_w10694_,
		_w13816_,
		_w14018_
	);
	LUT2 #(
		.INIT('h1)
	) name9972 (
		_w14011_,
		_w14016_,
		_w14019_
	);
	LUT2 #(
		.INIT('h1)
	) name9973 (
		_w14017_,
		_w14018_,
		_w14020_
	);
	LUT2 #(
		.INIT('h8)
	) name9974 (
		_w14019_,
		_w14020_,
		_w14021_
	);
	LUT2 #(
		.INIT('h4)
	) name9975 (
		_w14015_,
		_w14021_,
		_w14022_
	);
	LUT2 #(
		.INIT('h4)
	) name9976 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10702_,
		_w14023_
	);
	LUT2 #(
		.INIT('h8)
	) name9977 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w10698_,
		_w14024_
	);
	LUT2 #(
		.INIT('h2)
	) name9978 (
		_w13832_,
		_w14023_,
		_w14025_
	);
	LUT2 #(
		.INIT('h4)
	) name9979 (
		_w14024_,
		_w14025_,
		_w14026_
	);
	LUT2 #(
		.INIT('h2)
	) name9980 (
		_w14022_,
		_w14026_,
		_w14027_
	);
	LUT2 #(
		.INIT('h2)
	) name9981 (
		_w13853_,
		_w14027_,
		_w14028_
	);
	LUT2 #(
		.INIT('h4)
	) name9982 (
		_w13848_,
		_w14028_,
		_w14029_
	);
	LUT2 #(
		.INIT('h2)
	) name9983 (
		_w13848_,
		_w14028_,
		_w14030_
	);
	LUT2 #(
		.INIT('h1)
	) name9984 (
		_w14029_,
		_w14030_,
		_w14031_
	);
	LUT2 #(
		.INIT('h4)
	) name9985 (
		_w13874_,
		_w13880_,
		_w14032_
	);
	LUT2 #(
		.INIT('h4)
	) name9986 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14033_
	);
	LUT2 #(
		.INIT('h1)
	) name9987 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001 ,
		_w14034_
	);
	LUT2 #(
		.INIT('h2)
	) name9988 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001 ,
		_w14035_
	);
	LUT2 #(
		.INIT('h2)
	) name9989 (
		_w14033_,
		_w14034_,
		_w14036_
	);
	LUT2 #(
		.INIT('h4)
	) name9990 (
		_w14035_,
		_w14036_,
		_w14037_
	);
	LUT2 #(
		.INIT('h4)
	) name9991 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w10686_,
		_w14038_
	);
	LUT2 #(
		.INIT('h8)
	) name9992 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w10690_,
		_w14039_
	);
	LUT2 #(
		.INIT('h1)
	) name9993 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14038_,
		_w14040_
	);
	LUT2 #(
		.INIT('h4)
	) name9994 (
		_w14039_,
		_w14040_,
		_w14041_
	);
	LUT2 #(
		.INIT('h1)
	) name9995 (
		_w14037_,
		_w14041_,
		_w14042_
	);
	LUT2 #(
		.INIT('h1)
	) name9996 (
		_w13878_,
		_w14042_,
		_w14043_
	);
	LUT2 #(
		.INIT('h8)
	) name9997 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001 ,
		_w13878_,
		_w14044_
	);
	LUT2 #(
		.INIT('h1)
	) name9998 (
		_w14043_,
		_w14044_,
		_w14045_
	);
	LUT2 #(
		.INIT('h2)
	) name9999 (
		_w14032_,
		_w14045_,
		_w14046_
	);
	LUT2 #(
		.INIT('h8)
	) name10000 (
		_w13874_,
		_w14045_,
		_w14047_
	);
	LUT2 #(
		.INIT('h1)
	) name10001 (
		_w13840_,
		_w14046_,
		_w14048_
	);
	LUT2 #(
		.INIT('h4)
	) name10002 (
		_w14047_,
		_w14048_,
		_w14049_
	);
	LUT2 #(
		.INIT('h2)
	) name10003 (
		_w14031_,
		_w14049_,
		_w14050_
	);
	LUT2 #(
		.INIT('h1)
	) name10004 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7960_,
		_w14051_
	);
	LUT2 #(
		.INIT('h2)
	) name10005 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7956_,
		_w14052_
	);
	LUT2 #(
		.INIT('h2)
	) name10006 (
		_w13832_,
		_w14051_,
		_w14053_
	);
	LUT2 #(
		.INIT('h4)
	) name10007 (
		_w14052_,
		_w14053_,
		_w14054_
	);
	LUT2 #(
		.INIT('h4)
	) name10008 (
		_w7905_,
		_w13813_,
		_w14055_
	);
	LUT2 #(
		.INIT('h4)
	) name10009 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7987_,
		_w14056_
	);
	LUT2 #(
		.INIT('h8)
	) name10010 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7991_,
		_w14057_
	);
	LUT2 #(
		.INIT('h2)
	) name10011 (
		_w13823_,
		_w14056_,
		_w14058_
	);
	LUT2 #(
		.INIT('h4)
	) name10012 (
		_w14057_,
		_w14058_,
		_w14059_
	);
	LUT2 #(
		.INIT('h4)
	) name10013 (
		_w7909_,
		_w13819_,
		_w14060_
	);
	LUT2 #(
		.INIT('h4)
	) name10014 (
		_w7885_,
		_w13821_,
		_w14061_
	);
	LUT2 #(
		.INIT('h4)
	) name10015 (
		_w7952_,
		_w13816_,
		_w14062_
	);
	LUT2 #(
		.INIT('h1)
	) name10016 (
		_w14055_,
		_w14060_,
		_w14063_
	);
	LUT2 #(
		.INIT('h1)
	) name10017 (
		_w14061_,
		_w14062_,
		_w14064_
	);
	LUT2 #(
		.INIT('h8)
	) name10018 (
		_w14063_,
		_w14064_,
		_w14065_
	);
	LUT2 #(
		.INIT('h4)
	) name10019 (
		_w14059_,
		_w14065_,
		_w14066_
	);
	LUT2 #(
		.INIT('h4)
	) name10020 (
		_w13832_,
		_w14066_,
		_w14067_
	);
	LUT2 #(
		.INIT('h2)
	) name10021 (
		_w13853_,
		_w14054_,
		_w14068_
	);
	LUT2 #(
		.INIT('h4)
	) name10022 (
		_w14067_,
		_w14068_,
		_w14069_
	);
	LUT2 #(
		.INIT('h8)
	) name10023 (
		_w13848_,
		_w14069_,
		_w14070_
	);
	LUT2 #(
		.INIT('h1)
	) name10024 (
		_w13848_,
		_w14069_,
		_w14071_
	);
	LUT2 #(
		.INIT('h1)
	) name10025 (
		_w14070_,
		_w14071_,
		_w14072_
	);
	LUT2 #(
		.INIT('h1)
	) name10026 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001 ,
		_w14073_
	);
	LUT2 #(
		.INIT('h2)
	) name10027 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001 ,
		_w14074_
	);
	LUT2 #(
		.INIT('h2)
	) name10028 (
		_w14033_,
		_w14073_,
		_w14075_
	);
	LUT2 #(
		.INIT('h4)
	) name10029 (
		_w14074_,
		_w14075_,
		_w14076_
	);
	LUT2 #(
		.INIT('h4)
	) name10030 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7944_,
		_w14077_
	);
	LUT2 #(
		.INIT('h8)
	) name10031 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7948_,
		_w14078_
	);
	LUT2 #(
		.INIT('h1)
	) name10032 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14077_,
		_w14079_
	);
	LUT2 #(
		.INIT('h4)
	) name10033 (
		_w14078_,
		_w14079_,
		_w14080_
	);
	LUT2 #(
		.INIT('h1)
	) name10034 (
		_w14076_,
		_w14080_,
		_w14081_
	);
	LUT2 #(
		.INIT('h1)
	) name10035 (
		_w13878_,
		_w14081_,
		_w14082_
	);
	LUT2 #(
		.INIT('h8)
	) name10036 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001 ,
		_w13878_,
		_w14083_
	);
	LUT2 #(
		.INIT('h1)
	) name10037 (
		_w14082_,
		_w14083_,
		_w14084_
	);
	LUT2 #(
		.INIT('h2)
	) name10038 (
		_w14032_,
		_w14084_,
		_w14085_
	);
	LUT2 #(
		.INIT('h8)
	) name10039 (
		_w13874_,
		_w14084_,
		_w14086_
	);
	LUT2 #(
		.INIT('h1)
	) name10040 (
		_w13840_,
		_w14085_,
		_w14087_
	);
	LUT2 #(
		.INIT('h4)
	) name10041 (
		_w14086_,
		_w14087_,
		_w14088_
	);
	LUT2 #(
		.INIT('h8)
	) name10042 (
		_w14072_,
		_w14088_,
		_w14089_
	);
	LUT2 #(
		.INIT('h4)
	) name10043 (
		_w9865_,
		_w13813_,
		_w14090_
	);
	LUT2 #(
		.INIT('h4)
	) name10044 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9951_,
		_w14091_
	);
	LUT2 #(
		.INIT('h8)
	) name10045 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9947_,
		_w14092_
	);
	LUT2 #(
		.INIT('h2)
	) name10046 (
		_w13823_,
		_w14091_,
		_w14093_
	);
	LUT2 #(
		.INIT('h4)
	) name10047 (
		_w14092_,
		_w14093_,
		_w14094_
	);
	LUT2 #(
		.INIT('h4)
	) name10048 (
		_w9869_,
		_w13819_,
		_w14095_
	);
	LUT2 #(
		.INIT('h4)
	) name10049 (
		_w9845_,
		_w13821_,
		_w14096_
	);
	LUT2 #(
		.INIT('h4)
	) name10050 (
		_w9912_,
		_w13816_,
		_w14097_
	);
	LUT2 #(
		.INIT('h1)
	) name10051 (
		_w14090_,
		_w14095_,
		_w14098_
	);
	LUT2 #(
		.INIT('h1)
	) name10052 (
		_w14096_,
		_w14097_,
		_w14099_
	);
	LUT2 #(
		.INIT('h8)
	) name10053 (
		_w14098_,
		_w14099_,
		_w14100_
	);
	LUT2 #(
		.INIT('h4)
	) name10054 (
		_w14094_,
		_w14100_,
		_w14101_
	);
	LUT2 #(
		.INIT('h4)
	) name10055 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9920_,
		_w14102_
	);
	LUT2 #(
		.INIT('h8)
	) name10056 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9916_,
		_w14103_
	);
	LUT2 #(
		.INIT('h2)
	) name10057 (
		_w13832_,
		_w14102_,
		_w14104_
	);
	LUT2 #(
		.INIT('h4)
	) name10058 (
		_w14103_,
		_w14104_,
		_w14105_
	);
	LUT2 #(
		.INIT('h2)
	) name10059 (
		_w14101_,
		_w14105_,
		_w14106_
	);
	LUT2 #(
		.INIT('h2)
	) name10060 (
		_w13853_,
		_w14106_,
		_w14107_
	);
	LUT2 #(
		.INIT('h2)
	) name10061 (
		_w13848_,
		_w14107_,
		_w14108_
	);
	LUT2 #(
		.INIT('h4)
	) name10062 (
		_w13848_,
		_w14107_,
		_w14109_
	);
	LUT2 #(
		.INIT('h1)
	) name10063 (
		_w14108_,
		_w14109_,
		_w14110_
	);
	LUT2 #(
		.INIT('h4)
	) name10064 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001 ,
		_w13878_,
		_w14111_
	);
	LUT2 #(
		.INIT('h4)
	) name10065 (
		_w9908_,
		_w13881_,
		_w14112_
	);
	LUT2 #(
		.INIT('h4)
	) name10066 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9904_,
		_w14113_
	);
	LUT2 #(
		.INIT('h1)
	) name10067 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001 ,
		_w14114_
	);
	LUT2 #(
		.INIT('h2)
	) name10068 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001 ,
		_w14115_
	);
	LUT2 #(
		.INIT('h1)
	) name10069 (
		_w14114_,
		_w14115_,
		_w14116_
	);
	LUT2 #(
		.INIT('h2)
	) name10070 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14116_,
		_w14117_
	);
	LUT2 #(
		.INIT('h1)
	) name10071 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w14113_,
		_w14118_
	);
	LUT2 #(
		.INIT('h4)
	) name10072 (
		_w14117_,
		_w14118_,
		_w14119_
	);
	LUT2 #(
		.INIT('h1)
	) name10073 (
		_w13878_,
		_w14112_,
		_w14120_
	);
	LUT2 #(
		.INIT('h4)
	) name10074 (
		_w14119_,
		_w14120_,
		_w14121_
	);
	LUT2 #(
		.INIT('h2)
	) name10075 (
		_w13880_,
		_w14111_,
		_w14122_
	);
	LUT2 #(
		.INIT('h4)
	) name10076 (
		_w14121_,
		_w14122_,
		_w14123_
	);
	LUT2 #(
		.INIT('h2)
	) name10077 (
		_w13895_,
		_w14123_,
		_w14124_
	);
	LUT2 #(
		.INIT('h8)
	) name10078 (
		_w13874_,
		_w14123_,
		_w14125_
	);
	LUT2 #(
		.INIT('h1)
	) name10079 (
		_w14124_,
		_w14125_,
		_w14126_
	);
	LUT2 #(
		.INIT('h8)
	) name10080 (
		_w14110_,
		_w14126_,
		_w14127_
	);
	LUT2 #(
		.INIT('h4)
	) name10081 (
		_w14089_,
		_w14127_,
		_w14128_
	);
	LUT2 #(
		.INIT('h4)
	) name10082 (
		_w8534_,
		_w13813_,
		_w14129_
	);
	LUT2 #(
		.INIT('h4)
	) name10083 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w8493_,
		_w14130_
	);
	LUT2 #(
		.INIT('h8)
	) name10084 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w8497_,
		_w14131_
	);
	LUT2 #(
		.INIT('h2)
	) name10085 (
		_w13823_,
		_w14130_,
		_w14132_
	);
	LUT2 #(
		.INIT('h4)
	) name10086 (
		_w14131_,
		_w14132_,
		_w14133_
	);
	LUT2 #(
		.INIT('h4)
	) name10087 (
		_w8585_,
		_w13816_,
		_w14134_
	);
	LUT2 #(
		.INIT('h4)
	) name10088 (
		_w8554_,
		_w13819_,
		_w14135_
	);
	LUT2 #(
		.INIT('h4)
	) name10089 (
		_w8558_,
		_w13821_,
		_w14136_
	);
	LUT2 #(
		.INIT('h1)
	) name10090 (
		_w14129_,
		_w14134_,
		_w14137_
	);
	LUT2 #(
		.INIT('h1)
	) name10091 (
		_w14135_,
		_w14136_,
		_w14138_
	);
	LUT2 #(
		.INIT('h8)
	) name10092 (
		_w14137_,
		_w14138_,
		_w14139_
	);
	LUT2 #(
		.INIT('h4)
	) name10093 (
		_w14133_,
		_w14139_,
		_w14140_
	);
	LUT2 #(
		.INIT('h4)
	) name10094 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w8593_,
		_w14141_
	);
	LUT2 #(
		.INIT('h8)
	) name10095 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w8589_,
		_w14142_
	);
	LUT2 #(
		.INIT('h2)
	) name10096 (
		_w13832_,
		_w14141_,
		_w14143_
	);
	LUT2 #(
		.INIT('h4)
	) name10097 (
		_w14142_,
		_w14143_,
		_w14144_
	);
	LUT2 #(
		.INIT('h2)
	) name10098 (
		_w14140_,
		_w14144_,
		_w14145_
	);
	LUT2 #(
		.INIT('h2)
	) name10099 (
		_w13853_,
		_w14145_,
		_w14146_
	);
	LUT2 #(
		.INIT('h2)
	) name10100 (
		_w13848_,
		_w14146_,
		_w14147_
	);
	LUT2 #(
		.INIT('h4)
	) name10101 (
		_w13848_,
		_w14146_,
		_w14148_
	);
	LUT2 #(
		.INIT('h1)
	) name10102 (
		_w14147_,
		_w14148_,
		_w14149_
	);
	LUT2 #(
		.INIT('h4)
	) name10103 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001 ,
		_w13878_,
		_w14150_
	);
	LUT2 #(
		.INIT('h4)
	) name10104 (
		_w8581_,
		_w13881_,
		_w14151_
	);
	LUT2 #(
		.INIT('h4)
	) name10105 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w8577_,
		_w14152_
	);
	LUT2 #(
		.INIT('h1)
	) name10106 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001 ,
		_w14153_
	);
	LUT2 #(
		.INIT('h2)
	) name10107 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001 ,
		_w14154_
	);
	LUT2 #(
		.INIT('h1)
	) name10108 (
		_w14153_,
		_w14154_,
		_w14155_
	);
	LUT2 #(
		.INIT('h2)
	) name10109 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14155_,
		_w14156_
	);
	LUT2 #(
		.INIT('h1)
	) name10110 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w14152_,
		_w14157_
	);
	LUT2 #(
		.INIT('h4)
	) name10111 (
		_w14156_,
		_w14157_,
		_w14158_
	);
	LUT2 #(
		.INIT('h1)
	) name10112 (
		_w13878_,
		_w14151_,
		_w14159_
	);
	LUT2 #(
		.INIT('h4)
	) name10113 (
		_w14158_,
		_w14159_,
		_w14160_
	);
	LUT2 #(
		.INIT('h2)
	) name10114 (
		_w13880_,
		_w14150_,
		_w14161_
	);
	LUT2 #(
		.INIT('h4)
	) name10115 (
		_w14160_,
		_w14161_,
		_w14162_
	);
	LUT2 #(
		.INIT('h2)
	) name10116 (
		_w13895_,
		_w14162_,
		_w14163_
	);
	LUT2 #(
		.INIT('h8)
	) name10117 (
		_w13874_,
		_w14162_,
		_w14164_
	);
	LUT2 #(
		.INIT('h1)
	) name10118 (
		_w14163_,
		_w14164_,
		_w14165_
	);
	LUT2 #(
		.INIT('h1)
	) name10119 (
		_w14149_,
		_w14165_,
		_w14166_
	);
	LUT2 #(
		.INIT('h4)
	) name10120 (
		_w9229_,
		_w13813_,
		_w14167_
	);
	LUT2 #(
		.INIT('h4)
	) name10121 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9276_,
		_w14168_
	);
	LUT2 #(
		.INIT('h8)
	) name10122 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9280_,
		_w14169_
	);
	LUT2 #(
		.INIT('h2)
	) name10123 (
		_w13823_,
		_w14168_,
		_w14170_
	);
	LUT2 #(
		.INIT('h4)
	) name10124 (
		_w14169_,
		_w14170_,
		_w14171_
	);
	LUT2 #(
		.INIT('h4)
	) name10125 (
		_w9297_,
		_w13816_,
		_w14172_
	);
	LUT2 #(
		.INIT('h4)
	) name10126 (
		_w9225_,
		_w13819_,
		_w14173_
	);
	LUT2 #(
		.INIT('h4)
	) name10127 (
		_w9205_,
		_w13821_,
		_w14174_
	);
	LUT2 #(
		.INIT('h1)
	) name10128 (
		_w14167_,
		_w14172_,
		_w14175_
	);
	LUT2 #(
		.INIT('h1)
	) name10129 (
		_w14173_,
		_w14174_,
		_w14176_
	);
	LUT2 #(
		.INIT('h8)
	) name10130 (
		_w14175_,
		_w14176_,
		_w14177_
	);
	LUT2 #(
		.INIT('h4)
	) name10131 (
		_w14171_,
		_w14177_,
		_w14178_
	);
	LUT2 #(
		.INIT('h4)
	) name10132 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9309_,
		_w14179_
	);
	LUT2 #(
		.INIT('h8)
	) name10133 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9313_,
		_w14180_
	);
	LUT2 #(
		.INIT('h2)
	) name10134 (
		_w13832_,
		_w14179_,
		_w14181_
	);
	LUT2 #(
		.INIT('h4)
	) name10135 (
		_w14180_,
		_w14181_,
		_w14182_
	);
	LUT2 #(
		.INIT('h2)
	) name10136 (
		_w14178_,
		_w14182_,
		_w14183_
	);
	LUT2 #(
		.INIT('h2)
	) name10137 (
		_w13853_,
		_w14183_,
		_w14184_
	);
	LUT2 #(
		.INIT('h2)
	) name10138 (
		_w13848_,
		_w14184_,
		_w14185_
	);
	LUT2 #(
		.INIT('h4)
	) name10139 (
		_w13848_,
		_w14184_,
		_w14186_
	);
	LUT2 #(
		.INIT('h1)
	) name10140 (
		_w14185_,
		_w14186_,
		_w14187_
	);
	LUT2 #(
		.INIT('h4)
	) name10141 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001 ,
		_w13878_,
		_w14188_
	);
	LUT2 #(
		.INIT('h4)
	) name10142 (
		_w9301_,
		_w13881_,
		_w14189_
	);
	LUT2 #(
		.INIT('h4)
	) name10143 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9305_,
		_w14190_
	);
	LUT2 #(
		.INIT('h1)
	) name10144 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001 ,
		_w14191_
	);
	LUT2 #(
		.INIT('h2)
	) name10145 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001 ,
		_w14192_
	);
	LUT2 #(
		.INIT('h1)
	) name10146 (
		_w14191_,
		_w14192_,
		_w14193_
	);
	LUT2 #(
		.INIT('h2)
	) name10147 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14193_,
		_w14194_
	);
	LUT2 #(
		.INIT('h1)
	) name10148 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w14190_,
		_w14195_
	);
	LUT2 #(
		.INIT('h4)
	) name10149 (
		_w14194_,
		_w14195_,
		_w14196_
	);
	LUT2 #(
		.INIT('h1)
	) name10150 (
		_w13878_,
		_w14189_,
		_w14197_
	);
	LUT2 #(
		.INIT('h4)
	) name10151 (
		_w14196_,
		_w14197_,
		_w14198_
	);
	LUT2 #(
		.INIT('h2)
	) name10152 (
		_w13880_,
		_w14188_,
		_w14199_
	);
	LUT2 #(
		.INIT('h4)
	) name10153 (
		_w14198_,
		_w14199_,
		_w14200_
	);
	LUT2 #(
		.INIT('h2)
	) name10154 (
		_w13895_,
		_w14200_,
		_w14201_
	);
	LUT2 #(
		.INIT('h8)
	) name10155 (
		_w13874_,
		_w14200_,
		_w14202_
	);
	LUT2 #(
		.INIT('h1)
	) name10156 (
		_w14201_,
		_w14202_,
		_w14203_
	);
	LUT2 #(
		.INIT('h8)
	) name10157 (
		_w14187_,
		_w14203_,
		_w14204_
	);
	LUT2 #(
		.INIT('h4)
	) name10158 (
		_w7449_,
		_w13821_,
		_w14205_
	);
	LUT2 #(
		.INIT('h4)
	) name10159 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7381_,
		_w14206_
	);
	LUT2 #(
		.INIT('h8)
	) name10160 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7377_,
		_w14207_
	);
	LUT2 #(
		.INIT('h2)
	) name10161 (
		_w13823_,
		_w14206_,
		_w14208_
	);
	LUT2 #(
		.INIT('h4)
	) name10162 (
		_w14207_,
		_w14208_,
		_w14209_
	);
	LUT2 #(
		.INIT('h4)
	) name10163 (
		_w7469_,
		_w13819_,
		_w14210_
	);
	LUT2 #(
		.INIT('h4)
	) name10164 (
		_w7473_,
		_w13813_,
		_w14211_
	);
	LUT2 #(
		.INIT('h4)
	) name10165 (
		_w7422_,
		_w13816_,
		_w14212_
	);
	LUT2 #(
		.INIT('h1)
	) name10166 (
		_w14205_,
		_w14210_,
		_w14213_
	);
	LUT2 #(
		.INIT('h1)
	) name10167 (
		_w14211_,
		_w14212_,
		_w14214_
	);
	LUT2 #(
		.INIT('h8)
	) name10168 (
		_w14213_,
		_w14214_,
		_w14215_
	);
	LUT2 #(
		.INIT('h4)
	) name10169 (
		_w14209_,
		_w14215_,
		_w14216_
	);
	LUT2 #(
		.INIT('h1)
	) name10170 (
		_w13832_,
		_w14216_,
		_w14217_
	);
	LUT2 #(
		.INIT('h4)
	) name10171 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7430_,
		_w14218_
	);
	LUT2 #(
		.INIT('h8)
	) name10172 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7426_,
		_w14219_
	);
	LUT2 #(
		.INIT('h2)
	) name10173 (
		_w13832_,
		_w14218_,
		_w14220_
	);
	LUT2 #(
		.INIT('h4)
	) name10174 (
		_w14219_,
		_w14220_,
		_w14221_
	);
	LUT2 #(
		.INIT('h1)
	) name10175 (
		_w14217_,
		_w14221_,
		_w14222_
	);
	LUT2 #(
		.INIT('h2)
	) name10176 (
		_w13853_,
		_w14222_,
		_w14223_
	);
	LUT2 #(
		.INIT('h2)
	) name10177 (
		_w13848_,
		_w14223_,
		_w14224_
	);
	LUT2 #(
		.INIT('h4)
	) name10178 (
		_w13848_,
		_w14223_,
		_w14225_
	);
	LUT2 #(
		.INIT('h1)
	) name10179 (
		_w14224_,
		_w14225_,
		_w14226_
	);
	LUT2 #(
		.INIT('h4)
	) name10180 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001 ,
		_w13878_,
		_w14227_
	);
	LUT2 #(
		.INIT('h4)
	) name10181 (
		_w7418_,
		_w13881_,
		_w14228_
	);
	LUT2 #(
		.INIT('h4)
	) name10182 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w7414_,
		_w14229_
	);
	LUT2 #(
		.INIT('h1)
	) name10183 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001 ,
		_w14230_
	);
	LUT2 #(
		.INIT('h2)
	) name10184 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001 ,
		_w14231_
	);
	LUT2 #(
		.INIT('h1)
	) name10185 (
		_w14230_,
		_w14231_,
		_w14232_
	);
	LUT2 #(
		.INIT('h2)
	) name10186 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14232_,
		_w14233_
	);
	LUT2 #(
		.INIT('h1)
	) name10187 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w14229_,
		_w14234_
	);
	LUT2 #(
		.INIT('h4)
	) name10188 (
		_w14233_,
		_w14234_,
		_w14235_
	);
	LUT2 #(
		.INIT('h1)
	) name10189 (
		_w13878_,
		_w14228_,
		_w14236_
	);
	LUT2 #(
		.INIT('h4)
	) name10190 (
		_w14235_,
		_w14236_,
		_w14237_
	);
	LUT2 #(
		.INIT('h2)
	) name10191 (
		_w13880_,
		_w14227_,
		_w14238_
	);
	LUT2 #(
		.INIT('h4)
	) name10192 (
		_w14237_,
		_w14238_,
		_w14239_
	);
	LUT2 #(
		.INIT('h2)
	) name10193 (
		_w13895_,
		_w14239_,
		_w14240_
	);
	LUT2 #(
		.INIT('h8)
	) name10194 (
		_w13874_,
		_w14239_,
		_w14241_
	);
	LUT2 #(
		.INIT('h1)
	) name10195 (
		_w14240_,
		_w14241_,
		_w14242_
	);
	LUT2 #(
		.INIT('h1)
	) name10196 (
		_w14226_,
		_w14242_,
		_w14243_
	);
	LUT2 #(
		.INIT('h1)
	) name10197 (
		_w14187_,
		_w14203_,
		_w14244_
	);
	LUT2 #(
		.INIT('h8)
	) name10198 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w14245_
	);
	LUT2 #(
		.INIT('h1)
	) name10199 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[0]/NET0131 ,
		_w14245_,
		_w14246_
	);
	LUT2 #(
		.INIT('h1)
	) name10200 (
		_w13807_,
		_w13808_,
		_w14247_
	);
	LUT2 #(
		.INIT('h4)
	) name10201 (
		_w14246_,
		_w14247_,
		_w14248_
	);
	LUT2 #(
		.INIT('h8)
	) name10202 (
		_w13807_,
		_w13874_,
		_w14249_
	);
	LUT2 #(
		.INIT('h2)
	) name10203 (
		_w13842_,
		_w14249_,
		_w14250_
	);
	LUT2 #(
		.INIT('h4)
	) name10204 (
		_w14248_,
		_w14250_,
		_w14251_
	);
	LUT2 #(
		.INIT('h4)
	) name10205 (
		_w13838_,
		_w14251_,
		_w14252_
	);
	LUT2 #(
		.INIT('h1)
	) name10206 (
		_w14244_,
		_w14252_,
		_w14253_
	);
	LUT2 #(
		.INIT('h8)
	) name10207 (
		_w14226_,
		_w14242_,
		_w14254_
	);
	LUT2 #(
		.INIT('h1)
	) name10208 (
		_w14253_,
		_w14254_,
		_w14255_
	);
	LUT2 #(
		.INIT('h1)
	) name10209 (
		_w14243_,
		_w14255_,
		_w14256_
	);
	LUT2 #(
		.INIT('h1)
	) name10210 (
		_w14204_,
		_w14256_,
		_w14257_
	);
	LUT2 #(
		.INIT('h1)
	) name10211 (
		_w14166_,
		_w14257_,
		_w14258_
	);
	LUT2 #(
		.INIT('h4)
	) name10212 (
		_w14089_,
		_w14258_,
		_w14259_
	);
	LUT2 #(
		.INIT('h1)
	) name10213 (
		_w14072_,
		_w14088_,
		_w14260_
	);
	LUT2 #(
		.INIT('h4)
	) name10214 (
		_w14031_,
		_w14049_,
		_w14261_
	);
	LUT2 #(
		.INIT('h8)
	) name10215 (
		_w14149_,
		_w14165_,
		_w14262_
	);
	LUT2 #(
		.INIT('h4)
	) name10216 (
		_w14261_,
		_w14262_,
		_w14263_
	);
	LUT2 #(
		.INIT('h1)
	) name10217 (
		_w14260_,
		_w14263_,
		_w14264_
	);
	LUT2 #(
		.INIT('h4)
	) name10218 (
		_w14259_,
		_w14264_,
		_w14265_
	);
	LUT2 #(
		.INIT('h1)
	) name10219 (
		_w14110_,
		_w14126_,
		_w14266_
	);
	LUT2 #(
		.INIT('h1)
	) name10220 (
		_w14261_,
		_w14266_,
		_w14267_
	);
	LUT2 #(
		.INIT('h4)
	) name10221 (
		_w14265_,
		_w14267_,
		_w14268_
	);
	LUT2 #(
		.INIT('h1)
	) name10222 (
		_w14050_,
		_w14128_,
		_w14269_
	);
	LUT2 #(
		.INIT('h4)
	) name10223 (
		_w14268_,
		_w14269_,
		_w14270_
	);
	LUT2 #(
		.INIT('h1)
	) name10224 (
		_w13972_,
		_w14010_,
		_w14271_
	);
	LUT2 #(
		.INIT('h4)
	) name10225 (
		_w14270_,
		_w14271_,
		_w14272_
	);
	LUT2 #(
		.INIT('h8)
	) name10226 (
		_w13955_,
		_w13971_,
		_w14273_
	);
	LUT2 #(
		.INIT('h8)
	) name10227 (
		_w13993_,
		_w14009_,
		_w14274_
	);
	LUT2 #(
		.INIT('h4)
	) name10228 (
		_w13972_,
		_w14274_,
		_w14275_
	);
	LUT2 #(
		.INIT('h1)
	) name10229 (
		_w14273_,
		_w14275_,
		_w14276_
	);
	LUT2 #(
		.INIT('h4)
	) name10230 (
		_w14272_,
		_w14276_,
		_w14277_
	);
	LUT2 #(
		.INIT('h1)
	) name10231 (
		_w13898_,
		_w13935_,
		_w14278_
	);
	LUT2 #(
		.INIT('h4)
	) name10232 (
		_w14277_,
		_w14278_,
		_w14279_
	);
	LUT2 #(
		.INIT('h4)
	) name10233 (
		_w8354_,
		_w13819_,
		_w14280_
	);
	LUT2 #(
		.INIT('h4)
	) name10234 (
		_w8358_,
		_w13821_,
		_w14281_
	);
	LUT2 #(
		.INIT('h4)
	) name10235 (
		_w8385_,
		_w13816_,
		_w14282_
	);
	LUT2 #(
		.INIT('h4)
	) name10236 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w8402_,
		_w14283_
	);
	LUT2 #(
		.INIT('h8)
	) name10237 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w8410_,
		_w14284_
	);
	LUT2 #(
		.INIT('h2)
	) name10238 (
		_w13823_,
		_w14283_,
		_w14285_
	);
	LUT2 #(
		.INIT('h4)
	) name10239 (
		_w14284_,
		_w14285_,
		_w14286_
	);
	LUT2 #(
		.INIT('h1)
	) name10240 (
		_w13814_,
		_w14280_,
		_w14287_
	);
	LUT2 #(
		.INIT('h1)
	) name10241 (
		_w14281_,
		_w14282_,
		_w14288_
	);
	LUT2 #(
		.INIT('h8)
	) name10242 (
		_w14287_,
		_w14288_,
		_w14289_
	);
	LUT2 #(
		.INIT('h4)
	) name10243 (
		_w14286_,
		_w14289_,
		_w14290_
	);
	LUT2 #(
		.INIT('h4)
	) name10244 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w8369_,
		_w14291_
	);
	LUT2 #(
		.INIT('h8)
	) name10245 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w8373_,
		_w14292_
	);
	LUT2 #(
		.INIT('h2)
	) name10246 (
		_w13832_,
		_w14291_,
		_w14293_
	);
	LUT2 #(
		.INIT('h4)
	) name10247 (
		_w14292_,
		_w14293_,
		_w14294_
	);
	LUT2 #(
		.INIT('h2)
	) name10248 (
		_w14290_,
		_w14294_,
		_w14295_
	);
	LUT2 #(
		.INIT('h2)
	) name10249 (
		_w13853_,
		_w14295_,
		_w14296_
	);
	LUT2 #(
		.INIT('h4)
	) name10250 (
		_w13848_,
		_w14296_,
		_w14297_
	);
	LUT2 #(
		.INIT('h2)
	) name10251 (
		_w13848_,
		_w14296_,
		_w14298_
	);
	LUT2 #(
		.INIT('h1)
	) name10252 (
		_w14297_,
		_w14298_,
		_w14299_
	);
	LUT2 #(
		.INIT('h4)
	) name10253 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001 ,
		_w13878_,
		_w14300_
	);
	LUT2 #(
		.INIT('h4)
	) name10254 (
		_w8381_,
		_w13881_,
		_w14301_
	);
	LUT2 #(
		.INIT('h4)
	) name10255 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w8377_,
		_w14302_
	);
	LUT2 #(
		.INIT('h1)
	) name10256 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001 ,
		_w14303_
	);
	LUT2 #(
		.INIT('h2)
	) name10257 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001 ,
		_w14304_
	);
	LUT2 #(
		.INIT('h1)
	) name10258 (
		_w14303_,
		_w14304_,
		_w14305_
	);
	LUT2 #(
		.INIT('h2)
	) name10259 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14305_,
		_w14306_
	);
	LUT2 #(
		.INIT('h1)
	) name10260 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w14302_,
		_w14307_
	);
	LUT2 #(
		.INIT('h4)
	) name10261 (
		_w14306_,
		_w14307_,
		_w14308_
	);
	LUT2 #(
		.INIT('h1)
	) name10262 (
		_w13878_,
		_w14301_,
		_w14309_
	);
	LUT2 #(
		.INIT('h4)
	) name10263 (
		_w14308_,
		_w14309_,
		_w14310_
	);
	LUT2 #(
		.INIT('h2)
	) name10264 (
		_w13880_,
		_w14300_,
		_w14311_
	);
	LUT2 #(
		.INIT('h4)
	) name10265 (
		_w14310_,
		_w14311_,
		_w14312_
	);
	LUT2 #(
		.INIT('h4)
	) name10266 (
		_w13874_,
		_w14312_,
		_w14313_
	);
	LUT2 #(
		.INIT('h1)
	) name10267 (
		_w13895_,
		_w14312_,
		_w14314_
	);
	LUT2 #(
		.INIT('h1)
	) name10268 (
		_w14313_,
		_w14314_,
		_w14315_
	);
	LUT2 #(
		.INIT('h4)
	) name10269 (
		_w14299_,
		_w14315_,
		_w14316_
	);
	LUT2 #(
		.INIT('h8)
	) name10270 (
		_w13918_,
		_w13934_,
		_w14317_
	);
	LUT2 #(
		.INIT('h4)
	) name10271 (
		_w14316_,
		_w14317_,
		_w14318_
	);
	LUT2 #(
		.INIT('h2)
	) name10272 (
		_w13873_,
		_w13897_,
		_w14319_
	);
	LUT2 #(
		.INIT('h1)
	) name10273 (
		_w14318_,
		_w14319_,
		_w14320_
	);
	LUT2 #(
		.INIT('h4)
	) name10274 (
		_w14279_,
		_w14320_,
		_w14321_
	);
	LUT2 #(
		.INIT('h4)
	) name10275 (
		_w7753_,
		_w13819_,
		_w14322_
	);
	LUT2 #(
		.INIT('h4)
	) name10276 (
		_w7737_,
		_w13821_,
		_w14323_
	);
	LUT2 #(
		.INIT('h4)
	) name10277 (
		_w7784_,
		_w13816_,
		_w14324_
	);
	LUT2 #(
		.INIT('h4)
	) name10278 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7801_,
		_w14325_
	);
	LUT2 #(
		.INIT('h8)
	) name10279 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7809_,
		_w14326_
	);
	LUT2 #(
		.INIT('h2)
	) name10280 (
		_w13823_,
		_w14325_,
		_w14327_
	);
	LUT2 #(
		.INIT('h4)
	) name10281 (
		_w14326_,
		_w14327_,
		_w14328_
	);
	LUT2 #(
		.INIT('h1)
	) name10282 (
		_w13814_,
		_w14322_,
		_w14329_
	);
	LUT2 #(
		.INIT('h1)
	) name10283 (
		_w14323_,
		_w14324_,
		_w14330_
	);
	LUT2 #(
		.INIT('h8)
	) name10284 (
		_w14329_,
		_w14330_,
		_w14331_
	);
	LUT2 #(
		.INIT('h4)
	) name10285 (
		_w14328_,
		_w14331_,
		_w14332_
	);
	LUT2 #(
		.INIT('h4)
	) name10286 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7768_,
		_w14333_
	);
	LUT2 #(
		.INIT('h8)
	) name10287 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7780_,
		_w14334_
	);
	LUT2 #(
		.INIT('h2)
	) name10288 (
		_w13832_,
		_w14333_,
		_w14335_
	);
	LUT2 #(
		.INIT('h4)
	) name10289 (
		_w14334_,
		_w14335_,
		_w14336_
	);
	LUT2 #(
		.INIT('h2)
	) name10290 (
		_w14332_,
		_w14336_,
		_w14337_
	);
	LUT2 #(
		.INIT('h2)
	) name10291 (
		_w13853_,
		_w14337_,
		_w14338_
	);
	LUT2 #(
		.INIT('h2)
	) name10292 (
		_w13848_,
		_w14338_,
		_w14339_
	);
	LUT2 #(
		.INIT('h4)
	) name10293 (
		_w13848_,
		_w14338_,
		_w14340_
	);
	LUT2 #(
		.INIT('h1)
	) name10294 (
		_w14339_,
		_w14340_,
		_w14341_
	);
	LUT2 #(
		.INIT('h4)
	) name10295 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001 ,
		_w13878_,
		_w14342_
	);
	LUT2 #(
		.INIT('h4)
	) name10296 (
		_w7772_,
		_w13881_,
		_w14343_
	);
	LUT2 #(
		.INIT('h4)
	) name10297 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w7776_,
		_w14344_
	);
	LUT2 #(
		.INIT('h1)
	) name10298 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001 ,
		_w14345_
	);
	LUT2 #(
		.INIT('h2)
	) name10299 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001 ,
		_w14346_
	);
	LUT2 #(
		.INIT('h1)
	) name10300 (
		_w14345_,
		_w14346_,
		_w14347_
	);
	LUT2 #(
		.INIT('h2)
	) name10301 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14347_,
		_w14348_
	);
	LUT2 #(
		.INIT('h1)
	) name10302 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w14344_,
		_w14349_
	);
	LUT2 #(
		.INIT('h4)
	) name10303 (
		_w14348_,
		_w14349_,
		_w14350_
	);
	LUT2 #(
		.INIT('h1)
	) name10304 (
		_w13878_,
		_w14343_,
		_w14351_
	);
	LUT2 #(
		.INIT('h4)
	) name10305 (
		_w14350_,
		_w14351_,
		_w14352_
	);
	LUT2 #(
		.INIT('h2)
	) name10306 (
		_w13880_,
		_w14342_,
		_w14353_
	);
	LUT2 #(
		.INIT('h4)
	) name10307 (
		_w14352_,
		_w14353_,
		_w14354_
	);
	LUT2 #(
		.INIT('h4)
	) name10308 (
		_w13874_,
		_w14354_,
		_w14355_
	);
	LUT2 #(
		.INIT('h1)
	) name10309 (
		_w13895_,
		_w14354_,
		_w14356_
	);
	LUT2 #(
		.INIT('h1)
	) name10310 (
		_w14355_,
		_w14356_,
		_w14357_
	);
	LUT2 #(
		.INIT('h4)
	) name10311 (
		_w14341_,
		_w14357_,
		_w14358_
	);
	LUT2 #(
		.INIT('h1)
	) name10312 (
		_w14316_,
		_w14358_,
		_w14359_
	);
	LUT2 #(
		.INIT('h4)
	) name10313 (
		_w14321_,
		_w14359_,
		_w14360_
	);
	LUT2 #(
		.INIT('h2)
	) name10314 (
		_w14299_,
		_w14315_,
		_w14361_
	);
	LUT2 #(
		.INIT('h2)
	) name10315 (
		_w14341_,
		_w14357_,
		_w14362_
	);
	LUT2 #(
		.INIT('h4)
	) name10316 (
		_w13898_,
		_w14362_,
		_w14363_
	);
	LUT2 #(
		.INIT('h1)
	) name10317 (
		_w14361_,
		_w14363_,
		_w14364_
	);
	LUT2 #(
		.INIT('h4)
	) name10318 (
		_w14360_,
		_w14364_,
		_w14365_
	);
	LUT2 #(
		.INIT('h1)
	) name10319 (
		_w13809_,
		_w14365_,
		_w14366_
	);
	LUT2 #(
		.INIT('h4)
	) name10320 (
		_w9072_,
		_w13819_,
		_w14367_
	);
	LUT2 #(
		.INIT('h4)
	) name10321 (
		_w9056_,
		_w13821_,
		_w14368_
	);
	LUT2 #(
		.INIT('h4)
	) name10322 (
		_w9103_,
		_w13816_,
		_w14369_
	);
	LUT2 #(
		.INIT('h4)
	) name10323 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9120_,
		_w14370_
	);
	LUT2 #(
		.INIT('h8)
	) name10324 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9128_,
		_w14371_
	);
	LUT2 #(
		.INIT('h2)
	) name10325 (
		_w13823_,
		_w14370_,
		_w14372_
	);
	LUT2 #(
		.INIT('h4)
	) name10326 (
		_w14371_,
		_w14372_,
		_w14373_
	);
	LUT2 #(
		.INIT('h1)
	) name10327 (
		_w13814_,
		_w14367_,
		_w14374_
	);
	LUT2 #(
		.INIT('h1)
	) name10328 (
		_w14368_,
		_w14369_,
		_w14375_
	);
	LUT2 #(
		.INIT('h8)
	) name10329 (
		_w14374_,
		_w14375_,
		_w14376_
	);
	LUT2 #(
		.INIT('h4)
	) name10330 (
		_w14373_,
		_w14376_,
		_w14377_
	);
	LUT2 #(
		.INIT('h4)
	) name10331 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9091_,
		_w14378_
	);
	LUT2 #(
		.INIT('h8)
	) name10332 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w9099_,
		_w14379_
	);
	LUT2 #(
		.INIT('h2)
	) name10333 (
		_w13832_,
		_w14378_,
		_w14380_
	);
	LUT2 #(
		.INIT('h4)
	) name10334 (
		_w14379_,
		_w14380_,
		_w14381_
	);
	LUT2 #(
		.INIT('h2)
	) name10335 (
		_w14377_,
		_w14381_,
		_w14382_
	);
	LUT2 #(
		.INIT('h2)
	) name10336 (
		_w13853_,
		_w14382_,
		_w14383_
	);
	LUT2 #(
		.INIT('h2)
	) name10337 (
		_w13848_,
		_w14383_,
		_w14384_
	);
	LUT2 #(
		.INIT('h4)
	) name10338 (
		_w13848_,
		_w14383_,
		_w14385_
	);
	LUT2 #(
		.INIT('h1)
	) name10339 (
		_w14384_,
		_w14385_,
		_w14386_
	);
	LUT2 #(
		.INIT('h4)
	) name10340 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001 ,
		_w13878_,
		_w14387_
	);
	LUT2 #(
		.INIT('h4)
	) name10341 (
		_w9087_,
		_w13881_,
		_w14388_
	);
	LUT2 #(
		.INIT('h4)
	) name10342 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w9095_,
		_w14389_
	);
	LUT2 #(
		.INIT('h1)
	) name10343 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001 ,
		_w14390_
	);
	LUT2 #(
		.INIT('h2)
	) name10344 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001 ,
		_w14391_
	);
	LUT2 #(
		.INIT('h1)
	) name10345 (
		_w14390_,
		_w14391_,
		_w14392_
	);
	LUT2 #(
		.INIT('h2)
	) name10346 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14392_,
		_w14393_
	);
	LUT2 #(
		.INIT('h1)
	) name10347 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w14389_,
		_w14394_
	);
	LUT2 #(
		.INIT('h4)
	) name10348 (
		_w14393_,
		_w14394_,
		_w14395_
	);
	LUT2 #(
		.INIT('h1)
	) name10349 (
		_w13878_,
		_w14388_,
		_w14396_
	);
	LUT2 #(
		.INIT('h4)
	) name10350 (
		_w14395_,
		_w14396_,
		_w14397_
	);
	LUT2 #(
		.INIT('h2)
	) name10351 (
		_w13880_,
		_w14387_,
		_w14398_
	);
	LUT2 #(
		.INIT('h4)
	) name10352 (
		_w14397_,
		_w14398_,
		_w14399_
	);
	LUT2 #(
		.INIT('h2)
	) name10353 (
		_w13895_,
		_w14399_,
		_w14400_
	);
	LUT2 #(
		.INIT('h8)
	) name10354 (
		_w13874_,
		_w14399_,
		_w14401_
	);
	LUT2 #(
		.INIT('h1)
	) name10355 (
		_w14400_,
		_w14401_,
		_w14402_
	);
	LUT2 #(
		.INIT('h8)
	) name10356 (
		_w14386_,
		_w14402_,
		_w14403_
	);
	LUT2 #(
		.INIT('h8)
	) name10357 (
		_w13808_,
		_w13843_,
		_w14404_
	);
	LUT2 #(
		.INIT('h4)
	) name10358 (
		_w14403_,
		_w14404_,
		_w14405_
	);
	LUT2 #(
		.INIT('h4)
	) name10359 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[1]/NET0131 ,
		_w13808_,
		_w14406_
	);
	LUT2 #(
		.INIT('h2)
	) name10360 (
		_w14403_,
		_w14406_,
		_w14407_
	);
	LUT2 #(
		.INIT('h1)
	) name10361 (
		_w14386_,
		_w14402_,
		_w14408_
	);
	LUT2 #(
		.INIT('h1)
	) name10362 (
		_w14405_,
		_w14408_,
		_w14409_
	);
	LUT2 #(
		.INIT('h4)
	) name10363 (
		_w14407_,
		_w14409_,
		_w14410_
	);
	LUT2 #(
		.INIT('h2)
	) name10364 (
		_w14366_,
		_w14410_,
		_w14411_
	);
	LUT2 #(
		.INIT('h4)
	) name10365 (
		_w14366_,
		_w14410_,
		_w14412_
	);
	LUT2 #(
		.INIT('h1)
	) name10366 (
		_w14411_,
		_w14412_,
		_w14413_
	);
	LUT2 #(
		.INIT('h4)
	) name10367 (
		_w13806_,
		_w14413_,
		_w14414_
	);
	LUT2 #(
		.INIT('h2)
	) name10368 (
		_w14361_,
		_w14406_,
		_w14415_
	);
	LUT2 #(
		.INIT('h4)
	) name10369 (
		_w14361_,
		_w14404_,
		_w14416_
	);
	LUT2 #(
		.INIT('h1)
	) name10370 (
		_w14316_,
		_w14415_,
		_w14417_
	);
	LUT2 #(
		.INIT('h4)
	) name10371 (
		_w14416_,
		_w14417_,
		_w14418_
	);
	LUT2 #(
		.INIT('h2)
	) name10372 (
		_w14321_,
		_w14362_,
		_w14419_
	);
	LUT2 #(
		.INIT('h1)
	) name10373 (
		_w13809_,
		_w14358_,
		_w14420_
	);
	LUT2 #(
		.INIT('h4)
	) name10374 (
		_w14419_,
		_w14420_,
		_w14421_
	);
	LUT2 #(
		.INIT('h4)
	) name10375 (
		_w14418_,
		_w14421_,
		_w14422_
	);
	LUT2 #(
		.INIT('h2)
	) name10376 (
		_w14418_,
		_w14421_,
		_w14423_
	);
	LUT2 #(
		.INIT('h1)
	) name10377 (
		_w14422_,
		_w14423_,
		_w14424_
	);
	LUT2 #(
		.INIT('h8)
	) name10378 (
		_w13806_,
		_w14424_,
		_w14425_
	);
	LUT2 #(
		.INIT('h1)
	) name10379 (
		_w14414_,
		_w14425_,
		_w14426_
	);
	LUT2 #(
		.INIT('h2)
	) name10380 (
		_w13805_,
		_w14426_,
		_w14427_
	);
	LUT2 #(
		.INIT('h1)
	) name10381 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001 ,
		_w13805_,
		_w14428_
	);
	LUT2 #(
		.INIT('h1)
	) name10382 (
		_w14427_,
		_w14428_,
		_w14429_
	);
	LUT2 #(
		.INIT('h1)
	) name10383 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7096_,
		_w14430_
	);
	LUT2 #(
		.INIT('h2)
	) name10384 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7100_,
		_w14431_
	);
	LUT2 #(
		.INIT('h2)
	) name10385 (
		_w13832_,
		_w14430_,
		_w14432_
	);
	LUT2 #(
		.INIT('h4)
	) name10386 (
		_w14431_,
		_w14432_,
		_w14433_
	);
	LUT2 #(
		.INIT('h4)
	) name10387 (
		_w7182_,
		_w13819_,
		_w14434_
	);
	LUT2 #(
		.INIT('h4)
	) name10388 (
		_w7202_,
		_w13821_,
		_w14435_
	);
	LUT2 #(
		.INIT('h4)
	) name10389 (
		_w7112_,
		_w13816_,
		_w14436_
	);
	LUT2 #(
		.INIT('h4)
	) name10390 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7164_,
		_w14437_
	);
	LUT2 #(
		.INIT('h8)
	) name10391 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w7156_,
		_w14438_
	);
	LUT2 #(
		.INIT('h2)
	) name10392 (
		_w13823_,
		_w14437_,
		_w14439_
	);
	LUT2 #(
		.INIT('h4)
	) name10393 (
		_w14438_,
		_w14439_,
		_w14440_
	);
	LUT2 #(
		.INIT('h1)
	) name10394 (
		_w13814_,
		_w14434_,
		_w14441_
	);
	LUT2 #(
		.INIT('h1)
	) name10395 (
		_w14435_,
		_w14436_,
		_w14442_
	);
	LUT2 #(
		.INIT('h8)
	) name10396 (
		_w14441_,
		_w14442_,
		_w14443_
	);
	LUT2 #(
		.INIT('h4)
	) name10397 (
		_w14440_,
		_w14443_,
		_w14444_
	);
	LUT2 #(
		.INIT('h4)
	) name10398 (
		_w13832_,
		_w14444_,
		_w14445_
	);
	LUT2 #(
		.INIT('h2)
	) name10399 (
		_w13853_,
		_w14433_,
		_w14446_
	);
	LUT2 #(
		.INIT('h4)
	) name10400 (
		_w14445_,
		_w14446_,
		_w14447_
	);
	LUT2 #(
		.INIT('h8)
	) name10401 (
		_w13848_,
		_w14447_,
		_w14448_
	);
	LUT2 #(
		.INIT('h1)
	) name10402 (
		_w13848_,
		_w14447_,
		_w14449_
	);
	LUT2 #(
		.INIT('h1)
	) name10403 (
		_w14448_,
		_w14449_,
		_w14450_
	);
	LUT2 #(
		.INIT('h1)
	) name10404 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001 ,
		_w14451_
	);
	LUT2 #(
		.INIT('h2)
	) name10405 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001 ,
		_w14452_
	);
	LUT2 #(
		.INIT('h2)
	) name10406 (
		_w14033_,
		_w14451_,
		_w14453_
	);
	LUT2 #(
		.INIT('h4)
	) name10407 (
		_w14452_,
		_w14453_,
		_w14454_
	);
	LUT2 #(
		.INIT('h4)
	) name10408 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7104_,
		_w14455_
	);
	LUT2 #(
		.INIT('h8)
	) name10409 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7108_,
		_w14456_
	);
	LUT2 #(
		.INIT('h1)
	) name10410 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14455_,
		_w14457_
	);
	LUT2 #(
		.INIT('h4)
	) name10411 (
		_w14456_,
		_w14457_,
		_w14458_
	);
	LUT2 #(
		.INIT('h1)
	) name10412 (
		_w14454_,
		_w14458_,
		_w14459_
	);
	LUT2 #(
		.INIT('h1)
	) name10413 (
		_w13878_,
		_w14459_,
		_w14460_
	);
	LUT2 #(
		.INIT('h8)
	) name10414 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001 ,
		_w13878_,
		_w14461_
	);
	LUT2 #(
		.INIT('h1)
	) name10415 (
		_w14460_,
		_w14461_,
		_w14462_
	);
	LUT2 #(
		.INIT('h2)
	) name10416 (
		_w14032_,
		_w14462_,
		_w14463_
	);
	LUT2 #(
		.INIT('h8)
	) name10417 (
		_w13874_,
		_w14462_,
		_w14464_
	);
	LUT2 #(
		.INIT('h1)
	) name10418 (
		_w13840_,
		_w14463_,
		_w14465_
	);
	LUT2 #(
		.INIT('h4)
	) name10419 (
		_w14464_,
		_w14465_,
		_w14466_
	);
	LUT2 #(
		.INIT('h8)
	) name10420 (
		_w14450_,
		_w14466_,
		_w14467_
	);
	LUT2 #(
		.INIT('h1)
	) name10421 (
		_w14408_,
		_w14467_,
		_w14468_
	);
	LUT2 #(
		.INIT('h4)
	) name10422 (
		_w14365_,
		_w14468_,
		_w14469_
	);
	LUT2 #(
		.INIT('h1)
	) name10423 (
		_w14450_,
		_w14466_,
		_w14470_
	);
	LUT2 #(
		.INIT('h4)
	) name10424 (
		_w13837_,
		_w13853_,
		_w14471_
	);
	LUT2 #(
		.INIT('h2)
	) name10425 (
		_w13848_,
		_w14471_,
		_w14472_
	);
	LUT2 #(
		.INIT('h4)
	) name10426 (
		_w13848_,
		_w14471_,
		_w14473_
	);
	LUT2 #(
		.INIT('h1)
	) name10427 (
		_w14472_,
		_w14473_,
		_w14474_
	);
	LUT2 #(
		.INIT('h4)
	) name10428 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11975_,
		_w14475_
	);
	LUT2 #(
		.INIT('h8)
	) name10429 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11979_,
		_w14476_
	);
	LUT2 #(
		.INIT('h1)
	) name10430 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14475_,
		_w14477_
	);
	LUT2 #(
		.INIT('h4)
	) name10431 (
		_w14476_,
		_w14477_,
		_w14478_
	);
	LUT2 #(
		.INIT('h1)
	) name10432 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001 ,
		_w14479_
	);
	LUT2 #(
		.INIT('h2)
	) name10433 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001 ,
		_w14480_
	);
	LUT2 #(
		.INIT('h2)
	) name10434 (
		_w14033_,
		_w14479_,
		_w14481_
	);
	LUT2 #(
		.INIT('h4)
	) name10435 (
		_w14480_,
		_w14481_,
		_w14482_
	);
	LUT2 #(
		.INIT('h1)
	) name10436 (
		_w13878_,
		_w14482_,
		_w14483_
	);
	LUT2 #(
		.INIT('h4)
	) name10437 (
		_w14478_,
		_w14483_,
		_w14484_
	);
	LUT2 #(
		.INIT('h4)
	) name10438 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001 ,
		_w13878_,
		_w14485_
	);
	LUT2 #(
		.INIT('h1)
	) name10439 (
		_w14484_,
		_w14485_,
		_w14486_
	);
	LUT2 #(
		.INIT('h8)
	) name10440 (
		_w13880_,
		_w14486_,
		_w14487_
	);
	LUT2 #(
		.INIT('h4)
	) name10441 (
		_w13874_,
		_w14487_,
		_w14488_
	);
	LUT2 #(
		.INIT('h1)
	) name10442 (
		_w13895_,
		_w14487_,
		_w14489_
	);
	LUT2 #(
		.INIT('h1)
	) name10443 (
		_w14488_,
		_w14489_,
		_w14490_
	);
	LUT2 #(
		.INIT('h4)
	) name10444 (
		_w14474_,
		_w14490_,
		_w14491_
	);
	LUT2 #(
		.INIT('h2)
	) name10445 (
		_w14403_,
		_w14491_,
		_w14492_
	);
	LUT2 #(
		.INIT('h1)
	) name10446 (
		_w14470_,
		_w14492_,
		_w14493_
	);
	LUT2 #(
		.INIT('h4)
	) name10447 (
		_w14469_,
		_w14493_,
		_w14494_
	);
	LUT2 #(
		.INIT('h1)
	) name10448 (
		_w13809_,
		_w14494_,
		_w14495_
	);
	LUT2 #(
		.INIT('h4)
	) name10449 (
		_w11837_,
		_w13816_,
		_w14496_
	);
	LUT2 #(
		.INIT('h4)
	) name10450 (
		_w11878_,
		_w13819_,
		_w14497_
	);
	LUT2 #(
		.INIT('h4)
	) name10451 (
		_w11882_,
		_w13821_,
		_w14498_
	);
	LUT2 #(
		.INIT('h4)
	) name10452 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11846_,
		_w14499_
	);
	LUT2 #(
		.INIT('h8)
	) name10453 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11854_,
		_w14500_
	);
	LUT2 #(
		.INIT('h2)
	) name10454 (
		_w13823_,
		_w14499_,
		_w14501_
	);
	LUT2 #(
		.INIT('h4)
	) name10455 (
		_w14500_,
		_w14501_,
		_w14502_
	);
	LUT2 #(
		.INIT('h1)
	) name10456 (
		_w13814_,
		_w14496_,
		_w14503_
	);
	LUT2 #(
		.INIT('h1)
	) name10457 (
		_w14497_,
		_w14498_,
		_w14504_
	);
	LUT2 #(
		.INIT('h8)
	) name10458 (
		_w14503_,
		_w14504_,
		_w14505_
	);
	LUT2 #(
		.INIT('h4)
	) name10459 (
		_w14502_,
		_w14505_,
		_w14506_
	);
	LUT2 #(
		.INIT('h4)
	) name10460 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11821_,
		_w14507_
	);
	LUT2 #(
		.INIT('h8)
	) name10461 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w11825_,
		_w14508_
	);
	LUT2 #(
		.INIT('h2)
	) name10462 (
		_w13832_,
		_w14507_,
		_w14509_
	);
	LUT2 #(
		.INIT('h4)
	) name10463 (
		_w14508_,
		_w14509_,
		_w14510_
	);
	LUT2 #(
		.INIT('h2)
	) name10464 (
		_w14506_,
		_w14510_,
		_w14511_
	);
	LUT2 #(
		.INIT('h2)
	) name10465 (
		_w13853_,
		_w14511_,
		_w14512_
	);
	LUT2 #(
		.INIT('h2)
	) name10466 (
		_w13848_,
		_w14512_,
		_w14513_
	);
	LUT2 #(
		.INIT('h4)
	) name10467 (
		_w13848_,
		_w14512_,
		_w14514_
	);
	LUT2 #(
		.INIT('h1)
	) name10468 (
		_w14513_,
		_w14514_,
		_w14515_
	);
	LUT2 #(
		.INIT('h4)
	) name10469 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001 ,
		_w13878_,
		_w14516_
	);
	LUT2 #(
		.INIT('h4)
	) name10470 (
		_w11833_,
		_w13881_,
		_w14517_
	);
	LUT2 #(
		.INIT('h4)
	) name10471 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w11829_,
		_w14518_
	);
	LUT2 #(
		.INIT('h1)
	) name10472 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001 ,
		_w14519_
	);
	LUT2 #(
		.INIT('h2)
	) name10473 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001 ,
		_w14520_
	);
	LUT2 #(
		.INIT('h1)
	) name10474 (
		_w14519_,
		_w14520_,
		_w14521_
	);
	LUT2 #(
		.INIT('h2)
	) name10475 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w14521_,
		_w14522_
	);
	LUT2 #(
		.INIT('h1)
	) name10476 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w14518_,
		_w14523_
	);
	LUT2 #(
		.INIT('h4)
	) name10477 (
		_w14522_,
		_w14523_,
		_w14524_
	);
	LUT2 #(
		.INIT('h1)
	) name10478 (
		_w13878_,
		_w14517_,
		_w14525_
	);
	LUT2 #(
		.INIT('h4)
	) name10479 (
		_w14524_,
		_w14525_,
		_w14526_
	);
	LUT2 #(
		.INIT('h2)
	) name10480 (
		_w13880_,
		_w14516_,
		_w14527_
	);
	LUT2 #(
		.INIT('h4)
	) name10481 (
		_w14526_,
		_w14527_,
		_w14528_
	);
	LUT2 #(
		.INIT('h2)
	) name10482 (
		_w13895_,
		_w14528_,
		_w14529_
	);
	LUT2 #(
		.INIT('h8)
	) name10483 (
		_w13874_,
		_w14528_,
		_w14530_
	);
	LUT2 #(
		.INIT('h1)
	) name10484 (
		_w14529_,
		_w14530_,
		_w14531_
	);
	LUT2 #(
		.INIT('h8)
	) name10485 (
		_w14515_,
		_w14531_,
		_w14532_
	);
	LUT2 #(
		.INIT('h8)
	) name10486 (
		_w14406_,
		_w14532_,
		_w14533_
	);
	LUT2 #(
		.INIT('h1)
	) name10487 (
		_w14515_,
		_w14531_,
		_w14534_
	);
	LUT2 #(
		.INIT('h1)
	) name10488 (
		_w14404_,
		_w14532_,
		_w14535_
	);
	LUT2 #(
		.INIT('h4)
	) name10489 (
		_w14534_,
		_w14535_,
		_w14536_
	);
	LUT2 #(
		.INIT('h1)
	) name10490 (
		_w14533_,
		_w14536_,
		_w14537_
	);
	LUT2 #(
		.INIT('h2)
	) name10491 (
		_w14495_,
		_w14537_,
		_w14538_
	);
	LUT2 #(
		.INIT('h4)
	) name10492 (
		_w14495_,
		_w14537_,
		_w14539_
	);
	LUT2 #(
		.INIT('h1)
	) name10493 (
		_w14538_,
		_w14539_,
		_w14540_
	);
	LUT2 #(
		.INIT('h1)
	) name10494 (
		_w13806_,
		_w14540_,
		_w14541_
	);
	LUT2 #(
		.INIT('h2)
	) name10495 (
		_w14404_,
		_w14470_,
		_w14542_
	);
	LUT2 #(
		.INIT('h4)
	) name10496 (
		_w14406_,
		_w14470_,
		_w14543_
	);
	LUT2 #(
		.INIT('h1)
	) name10497 (
		_w14467_,
		_w14542_,
		_w14544_
	);
	LUT2 #(
		.INIT('h4)
	) name10498 (
		_w14543_,
		_w14544_,
		_w14545_
	);
	LUT2 #(
		.INIT('h2)
	) name10499 (
		_w14365_,
		_w14403_,
		_w14546_
	);
	LUT2 #(
		.INIT('h1)
	) name10500 (
		_w13809_,
		_w14408_,
		_w14547_
	);
	LUT2 #(
		.INIT('h4)
	) name10501 (
		_w14546_,
		_w14547_,
		_w14548_
	);
	LUT2 #(
		.INIT('h4)
	) name10502 (
		_w14545_,
		_w14548_,
		_w14549_
	);
	LUT2 #(
		.INIT('h2)
	) name10503 (
		_w14545_,
		_w14548_,
		_w14550_
	);
	LUT2 #(
		.INIT('h1)
	) name10504 (
		_w14549_,
		_w14550_,
		_w14551_
	);
	LUT2 #(
		.INIT('h8)
	) name10505 (
		_w13806_,
		_w14551_,
		_w14552_
	);
	LUT2 #(
		.INIT('h1)
	) name10506 (
		_w14541_,
		_w14552_,
		_w14553_
	);
	LUT2 #(
		.INIT('h2)
	) name10507 (
		_w13805_,
		_w14553_,
		_w14554_
	);
	LUT2 #(
		.INIT('h1)
	) name10508 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001 ,
		_w13805_,
		_w14555_
	);
	LUT2 #(
		.INIT('h1)
	) name10509 (
		_w14554_,
		_w14555_,
		_w14556_
	);
	LUT2 #(
		.INIT('h1)
	) name10510 (
		_w13809_,
		_w14252_,
		_w14557_
	);
	LUT2 #(
		.INIT('h2)
	) name10511 (
		_w14254_,
		_w14406_,
		_w14558_
	);
	LUT2 #(
		.INIT('h4)
	) name10512 (
		_w14254_,
		_w14404_,
		_w14559_
	);
	LUT2 #(
		.INIT('h1)
	) name10513 (
		_w14243_,
		_w14558_,
		_w14560_
	);
	LUT2 #(
		.INIT('h4)
	) name10514 (
		_w14559_,
		_w14560_,
		_w14561_
	);
	LUT2 #(
		.INIT('h2)
	) name10515 (
		_w14557_,
		_w14561_,
		_w14562_
	);
	LUT2 #(
		.INIT('h4)
	) name10516 (
		_w14557_,
		_w14561_,
		_w14563_
	);
	LUT2 #(
		.INIT('h1)
	) name10517 (
		_w14562_,
		_w14563_,
		_w14564_
	);
	LUT2 #(
		.INIT('h2)
	) name10518 (
		_w13806_,
		_w14564_,
		_w14565_
	);
	LUT2 #(
		.INIT('h1)
	) name10519 (
		_w13809_,
		_w14255_,
		_w14566_
	);
	LUT2 #(
		.INIT('h8)
	) name10520 (
		_w14204_,
		_w14406_,
		_w14567_
	);
	LUT2 #(
		.INIT('h1)
	) name10521 (
		_w14204_,
		_w14404_,
		_w14568_
	);
	LUT2 #(
		.INIT('h4)
	) name10522 (
		_w14244_,
		_w14568_,
		_w14569_
	);
	LUT2 #(
		.INIT('h1)
	) name10523 (
		_w14567_,
		_w14569_,
		_w14570_
	);
	LUT2 #(
		.INIT('h2)
	) name10524 (
		_w14566_,
		_w14570_,
		_w14571_
	);
	LUT2 #(
		.INIT('h4)
	) name10525 (
		_w14566_,
		_w14570_,
		_w14572_
	);
	LUT2 #(
		.INIT('h1)
	) name10526 (
		_w14571_,
		_w14572_,
		_w14573_
	);
	LUT2 #(
		.INIT('h4)
	) name10527 (
		_w13806_,
		_w14573_,
		_w14574_
	);
	LUT2 #(
		.INIT('h1)
	) name10528 (
		_w14565_,
		_w14574_,
		_w14575_
	);
	LUT2 #(
		.INIT('h2)
	) name10529 (
		_w13805_,
		_w14575_,
		_w14576_
	);
	LUT2 #(
		.INIT('h2)
	) name10530 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001 ,
		_w13805_,
		_w14577_
	);
	LUT2 #(
		.INIT('h1)
	) name10531 (
		_w14576_,
		_w14577_,
		_w14578_
	);
	LUT2 #(
		.INIT('h1)
	) name10532 (
		_w13809_,
		_w14257_,
		_w14579_
	);
	LUT2 #(
		.INIT('h2)
	) name10533 (
		_w14262_,
		_w14406_,
		_w14580_
	);
	LUT2 #(
		.INIT('h4)
	) name10534 (
		_w14262_,
		_w14404_,
		_w14581_
	);
	LUT2 #(
		.INIT('h1)
	) name10535 (
		_w14166_,
		_w14580_,
		_w14582_
	);
	LUT2 #(
		.INIT('h4)
	) name10536 (
		_w14581_,
		_w14582_,
		_w14583_
	);
	LUT2 #(
		.INIT('h2)
	) name10537 (
		_w14579_,
		_w14583_,
		_w14584_
	);
	LUT2 #(
		.INIT('h4)
	) name10538 (
		_w14579_,
		_w14583_,
		_w14585_
	);
	LUT2 #(
		.INIT('h1)
	) name10539 (
		_w14584_,
		_w14585_,
		_w14586_
	);
	LUT2 #(
		.INIT('h1)
	) name10540 (
		_w13806_,
		_w14586_,
		_w14587_
	);
	LUT2 #(
		.INIT('h8)
	) name10541 (
		_w13806_,
		_w14573_,
		_w14588_
	);
	LUT2 #(
		.INIT('h1)
	) name10542 (
		_w14587_,
		_w14588_,
		_w14589_
	);
	LUT2 #(
		.INIT('h2)
	) name10543 (
		_w13805_,
		_w14589_,
		_w14590_
	);
	LUT2 #(
		.INIT('h2)
	) name10544 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001 ,
		_w13805_,
		_w14591_
	);
	LUT2 #(
		.INIT('h1)
	) name10545 (
		_w14590_,
		_w14591_,
		_w14592_
	);
	LUT2 #(
		.INIT('h1)
	) name10546 (
		_w13809_,
		_w14265_,
		_w14593_
	);
	LUT2 #(
		.INIT('h2)
	) name10547 (
		_w14127_,
		_w14406_,
		_w14594_
	);
	LUT2 #(
		.INIT('h4)
	) name10548 (
		_w14127_,
		_w14404_,
		_w14595_
	);
	LUT2 #(
		.INIT('h1)
	) name10549 (
		_w14266_,
		_w14594_,
		_w14596_
	);
	LUT2 #(
		.INIT('h4)
	) name10550 (
		_w14595_,
		_w14596_,
		_w14597_
	);
	LUT2 #(
		.INIT('h2)
	) name10551 (
		_w14593_,
		_w14597_,
		_w14598_
	);
	LUT2 #(
		.INIT('h4)
	) name10552 (
		_w14593_,
		_w14597_,
		_w14599_
	);
	LUT2 #(
		.INIT('h1)
	) name10553 (
		_w14598_,
		_w14599_,
		_w14600_
	);
	LUT2 #(
		.INIT('h1)
	) name10554 (
		_w13806_,
		_w14600_,
		_w14601_
	);
	LUT2 #(
		.INIT('h1)
	) name10555 (
		_w14258_,
		_w14262_,
		_w14602_
	);
	LUT2 #(
		.INIT('h1)
	) name10556 (
		_w13809_,
		_w14602_,
		_w14603_
	);
	LUT2 #(
		.INIT('h2)
	) name10557 (
		_w14260_,
		_w14406_,
		_w14604_
	);
	LUT2 #(
		.INIT('h4)
	) name10558 (
		_w14260_,
		_w14404_,
		_w14605_
	);
	LUT2 #(
		.INIT('h1)
	) name10559 (
		_w14089_,
		_w14604_,
		_w14606_
	);
	LUT2 #(
		.INIT('h4)
	) name10560 (
		_w14605_,
		_w14606_,
		_w14607_
	);
	LUT2 #(
		.INIT('h2)
	) name10561 (
		_w14603_,
		_w14607_,
		_w14608_
	);
	LUT2 #(
		.INIT('h4)
	) name10562 (
		_w14603_,
		_w14607_,
		_w14609_
	);
	LUT2 #(
		.INIT('h1)
	) name10563 (
		_w14608_,
		_w14609_,
		_w14610_
	);
	LUT2 #(
		.INIT('h2)
	) name10564 (
		_w13806_,
		_w14610_,
		_w14611_
	);
	LUT2 #(
		.INIT('h1)
	) name10565 (
		_w14601_,
		_w14611_,
		_w14612_
	);
	LUT2 #(
		.INIT('h2)
	) name10566 (
		_w13805_,
		_w14612_,
		_w14613_
	);
	LUT2 #(
		.INIT('h2)
	) name10567 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001 ,
		_w13805_,
		_w14614_
	);
	LUT2 #(
		.INIT('h1)
	) name10568 (
		_w14613_,
		_w14614_,
		_w14615_
	);
	LUT2 #(
		.INIT('h1)
	) name10569 (
		_w13809_,
		_w14270_,
		_w14616_
	);
	LUT2 #(
		.INIT('h2)
	) name10570 (
		_w14274_,
		_w14406_,
		_w14617_
	);
	LUT2 #(
		.INIT('h4)
	) name10571 (
		_w14274_,
		_w14404_,
		_w14618_
	);
	LUT2 #(
		.INIT('h1)
	) name10572 (
		_w14010_,
		_w14617_,
		_w14619_
	);
	LUT2 #(
		.INIT('h4)
	) name10573 (
		_w14618_,
		_w14619_,
		_w14620_
	);
	LUT2 #(
		.INIT('h2)
	) name10574 (
		_w14616_,
		_w14620_,
		_w14621_
	);
	LUT2 #(
		.INIT('h4)
	) name10575 (
		_w14616_,
		_w14620_,
		_w14622_
	);
	LUT2 #(
		.INIT('h1)
	) name10576 (
		_w14621_,
		_w14622_,
		_w14623_
	);
	LUT2 #(
		.INIT('h1)
	) name10577 (
		_w13806_,
		_w14623_,
		_w14624_
	);
	LUT2 #(
		.INIT('h2)
	) name10578 (
		_w14050_,
		_w14406_,
		_w14625_
	);
	LUT2 #(
		.INIT('h4)
	) name10579 (
		_w14050_,
		_w14404_,
		_w14626_
	);
	LUT2 #(
		.INIT('h1)
	) name10580 (
		_w14261_,
		_w14625_,
		_w14627_
	);
	LUT2 #(
		.INIT('h4)
	) name10581 (
		_w14626_,
		_w14627_,
		_w14628_
	);
	LUT2 #(
		.INIT('h4)
	) name10582 (
		_w14127_,
		_w14265_,
		_w14629_
	);
	LUT2 #(
		.INIT('h1)
	) name10583 (
		_w13809_,
		_w14266_,
		_w14630_
	);
	LUT2 #(
		.INIT('h4)
	) name10584 (
		_w14629_,
		_w14630_,
		_w14631_
	);
	LUT2 #(
		.INIT('h4)
	) name10585 (
		_w14628_,
		_w14631_,
		_w14632_
	);
	LUT2 #(
		.INIT('h2)
	) name10586 (
		_w14628_,
		_w14631_,
		_w14633_
	);
	LUT2 #(
		.INIT('h1)
	) name10587 (
		_w14632_,
		_w14633_,
		_w14634_
	);
	LUT2 #(
		.INIT('h2)
	) name10588 (
		_w13806_,
		_w14634_,
		_w14635_
	);
	LUT2 #(
		.INIT('h1)
	) name10589 (
		_w14624_,
		_w14635_,
		_w14636_
	);
	LUT2 #(
		.INIT('h2)
	) name10590 (
		_w13805_,
		_w14636_,
		_w14637_
	);
	LUT2 #(
		.INIT('h2)
	) name10591 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001 ,
		_w13805_,
		_w14638_
	);
	LUT2 #(
		.INIT('h1)
	) name10592 (
		_w14637_,
		_w14638_,
		_w14639_
	);
	LUT2 #(
		.INIT('h2)
	) name10593 (
		_w14319_,
		_w14406_,
		_w14640_
	);
	LUT2 #(
		.INIT('h4)
	) name10594 (
		_w14319_,
		_w14404_,
		_w14641_
	);
	LUT2 #(
		.INIT('h1)
	) name10595 (
		_w13898_,
		_w14640_,
		_w14642_
	);
	LUT2 #(
		.INIT('h4)
	) name10596 (
		_w14641_,
		_w14642_,
		_w14643_
	);
	LUT2 #(
		.INIT('h2)
	) name10597 (
		_w14277_,
		_w14317_,
		_w14644_
	);
	LUT2 #(
		.INIT('h1)
	) name10598 (
		_w13809_,
		_w13935_,
		_w14645_
	);
	LUT2 #(
		.INIT('h4)
	) name10599 (
		_w14644_,
		_w14645_,
		_w14646_
	);
	LUT2 #(
		.INIT('h4)
	) name10600 (
		_w14643_,
		_w14646_,
		_w14647_
	);
	LUT2 #(
		.INIT('h2)
	) name10601 (
		_w14643_,
		_w14646_,
		_w14648_
	);
	LUT2 #(
		.INIT('h1)
	) name10602 (
		_w14647_,
		_w14648_,
		_w14649_
	);
	LUT2 #(
		.INIT('h1)
	) name10603 (
		_w13806_,
		_w14649_,
		_w14650_
	);
	LUT2 #(
		.INIT('h1)
	) name10604 (
		_w13809_,
		_w14277_,
		_w14651_
	);
	LUT2 #(
		.INIT('h2)
	) name10605 (
		_w14317_,
		_w14406_,
		_w14652_
	);
	LUT2 #(
		.INIT('h4)
	) name10606 (
		_w14317_,
		_w14404_,
		_w14653_
	);
	LUT2 #(
		.INIT('h1)
	) name10607 (
		_w13935_,
		_w14652_,
		_w14654_
	);
	LUT2 #(
		.INIT('h4)
	) name10608 (
		_w14653_,
		_w14654_,
		_w14655_
	);
	LUT2 #(
		.INIT('h2)
	) name10609 (
		_w14651_,
		_w14655_,
		_w14656_
	);
	LUT2 #(
		.INIT('h4)
	) name10610 (
		_w14651_,
		_w14655_,
		_w14657_
	);
	LUT2 #(
		.INIT('h1)
	) name10611 (
		_w14656_,
		_w14657_,
		_w14658_
	);
	LUT2 #(
		.INIT('h2)
	) name10612 (
		_w13806_,
		_w14658_,
		_w14659_
	);
	LUT2 #(
		.INIT('h1)
	) name10613 (
		_w14650_,
		_w14659_,
		_w14660_
	);
	LUT2 #(
		.INIT('h2)
	) name10614 (
		_w13805_,
		_w14660_,
		_w14661_
	);
	LUT2 #(
		.INIT('h2)
	) name10615 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001 ,
		_w13805_,
		_w14662_
	);
	LUT2 #(
		.INIT('h1)
	) name10616 (
		_w14661_,
		_w14662_,
		_w14663_
	);
	LUT2 #(
		.INIT('h2)
	) name10617 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w5950_,
		_w14664_
	);
	LUT2 #(
		.INIT('h4)
	) name10618 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w14664_,
		_w14665_
	);
	LUT2 #(
		.INIT('h4)
	) name10619 (
		_w13802_,
		_w14665_,
		_w14666_
	);
	LUT2 #(
		.INIT('h4)
	) name10620 (
		_w13800_,
		_w14666_,
		_w14667_
	);
	LUT2 #(
		.INIT('h4)
	) name10621 (
		_w14426_,
		_w14667_,
		_w14668_
	);
	LUT2 #(
		.INIT('h1)
	) name10622 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001 ,
		_w14667_,
		_w14669_
	);
	LUT2 #(
		.INIT('h1)
	) name10623 (
		_w14668_,
		_w14669_,
		_w14670_
	);
	LUT2 #(
		.INIT('h4)
	) name10624 (
		_w14553_,
		_w14667_,
		_w14671_
	);
	LUT2 #(
		.INIT('h1)
	) name10625 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001 ,
		_w14667_,
		_w14672_
	);
	LUT2 #(
		.INIT('h1)
	) name10626 (
		_w14671_,
		_w14672_,
		_w14673_
	);
	LUT2 #(
		.INIT('h4)
	) name10627 (
		_w14575_,
		_w14667_,
		_w14674_
	);
	LUT2 #(
		.INIT('h2)
	) name10628 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001 ,
		_w14667_,
		_w14675_
	);
	LUT2 #(
		.INIT('h1)
	) name10629 (
		_w14674_,
		_w14675_,
		_w14676_
	);
	LUT2 #(
		.INIT('h4)
	) name10630 (
		_w14589_,
		_w14667_,
		_w14677_
	);
	LUT2 #(
		.INIT('h2)
	) name10631 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001 ,
		_w14667_,
		_w14678_
	);
	LUT2 #(
		.INIT('h1)
	) name10632 (
		_w14677_,
		_w14678_,
		_w14679_
	);
	LUT2 #(
		.INIT('h4)
	) name10633 (
		_w14612_,
		_w14667_,
		_w14680_
	);
	LUT2 #(
		.INIT('h2)
	) name10634 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001 ,
		_w14667_,
		_w14681_
	);
	LUT2 #(
		.INIT('h1)
	) name10635 (
		_w14680_,
		_w14681_,
		_w14682_
	);
	LUT2 #(
		.INIT('h4)
	) name10636 (
		_w14636_,
		_w14667_,
		_w14683_
	);
	LUT2 #(
		.INIT('h2)
	) name10637 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001 ,
		_w14667_,
		_w14684_
	);
	LUT2 #(
		.INIT('h1)
	) name10638 (
		_w14683_,
		_w14684_,
		_w14685_
	);
	LUT2 #(
		.INIT('h4)
	) name10639 (
		_w14660_,
		_w14667_,
		_w14686_
	);
	LUT2 #(
		.INIT('h2)
	) name10640 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001 ,
		_w14667_,
		_w14687_
	);
	LUT2 #(
		.INIT('h1)
	) name10641 (
		_w14686_,
		_w14687_,
		_w14688_
	);
	LUT2 #(
		.INIT('h8)
	) name10642 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w11525_,
		_w14689_
	);
	LUT2 #(
		.INIT('h2)
	) name10643 (
		\core_c_dec_RTI_Ed_reg/P0001 ,
		_w4184_,
		_w14690_
	);
	LUT2 #(
		.INIT('h8)
	) name10644 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w14691_
	);
	LUT2 #(
		.INIT('h1)
	) name10645 (
		_w14690_,
		_w14691_,
		_w14692_
	);
	LUT2 #(
		.INIT('h1)
	) name10646 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w14690_,
		_w14693_
	);
	LUT2 #(
		.INIT('h8)
	) name10647 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		_w14694_
	);
	LUT2 #(
		.INIT('h8)
	) name10648 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w14694_,
		_w14695_
	);
	LUT2 #(
		.INIT('h1)
	) name10649 (
		_w14693_,
		_w14695_,
		_w14696_
	);
	LUT2 #(
		.INIT('h4)
	) name10650 (
		_w14692_,
		_w14696_,
		_w14697_
	);
	LUT2 #(
		.INIT('h2)
	) name10651 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		_w14698_
	);
	LUT2 #(
		.INIT('h8)
	) name10652 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w14698_,
		_w14699_
	);
	LUT2 #(
		.INIT('h8)
	) name10653 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001 ,
		_w14699_,
		_w14700_
	);
	LUT2 #(
		.INIT('h1)
	) name10654 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		_w14701_
	);
	LUT2 #(
		.INIT('h4)
	) name10655 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w14701_,
		_w14702_
	);
	LUT2 #(
		.INIT('h8)
	) name10656 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001 ,
		_w14702_,
		_w14703_
	);
	LUT2 #(
		.INIT('h4)
	) name10657 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w14694_,
		_w14704_
	);
	LUT2 #(
		.INIT('h8)
	) name10658 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001 ,
		_w14704_,
		_w14705_
	);
	LUT2 #(
		.INIT('h8)
	) name10659 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w14701_,
		_w14706_
	);
	LUT2 #(
		.INIT('h8)
	) name10660 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001 ,
		_w14706_,
		_w14707_
	);
	LUT2 #(
		.INIT('h4)
	) name10661 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w14698_,
		_w14708_
	);
	LUT2 #(
		.INIT('h8)
	) name10662 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001 ,
		_w14708_,
		_w14709_
	);
	LUT2 #(
		.INIT('h4)
	) name10663 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		\core_c_psq_ststk_ptr_reg[1]/NET0131 ,
		_w14710_
	);
	LUT2 #(
		.INIT('h8)
	) name10664 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w14710_,
		_w14711_
	);
	LUT2 #(
		.INIT('h8)
	) name10665 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001 ,
		_w14711_,
		_w14712_
	);
	LUT2 #(
		.INIT('h4)
	) name10666 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w14710_,
		_w14713_
	);
	LUT2 #(
		.INIT('h8)
	) name10667 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001 ,
		_w14713_,
		_w14714_
	);
	LUT2 #(
		.INIT('h1)
	) name10668 (
		_w14700_,
		_w14703_,
		_w14715_
	);
	LUT2 #(
		.INIT('h1)
	) name10669 (
		_w14705_,
		_w14707_,
		_w14716_
	);
	LUT2 #(
		.INIT('h1)
	) name10670 (
		_w14709_,
		_w14712_,
		_w14717_
	);
	LUT2 #(
		.INIT('h4)
	) name10671 (
		_w14714_,
		_w14717_,
		_w14718_
	);
	LUT2 #(
		.INIT('h8)
	) name10672 (
		_w14715_,
		_w14716_,
		_w14719_
	);
	LUT2 #(
		.INIT('h8)
	) name10673 (
		_w14718_,
		_w14719_,
		_w14720_
	);
	LUT2 #(
		.INIT('h2)
	) name10674 (
		_w14697_,
		_w14720_,
		_w14721_
	);
	LUT2 #(
		.INIT('h1)
	) name10675 (
		_w14689_,
		_w14721_,
		_w14722_
	);
	LUT2 #(
		.INIT('h1)
	) name10676 (
		_w5950_,
		_w14722_,
		_w14723_
	);
	LUT2 #(
		.INIT('h8)
	) name10677 (
		\core_eu_ec_cun_MVi_pre_C_reg/P0001 ,
		_w5950_,
		_w14724_
	);
	LUT2 #(
		.INIT('h1)
	) name10678 (
		_w14723_,
		_w14724_,
		_w14725_
	);
	LUT2 #(
		.INIT('h4)
	) name10679 (
		\core_eu_em_mac_em_reg_Sq_E_reg/P0001 ,
		_w4117_,
		_w14726_
	);
	LUT2 #(
		.INIT('h8)
	) name10680 (
		_w6022_,
		_w6026_,
		_w14727_
	);
	LUT2 #(
		.INIT('h4)
	) name10681 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w14727_,
		_w14728_
	);
	LUT2 #(
		.INIT('h1)
	) name10682 (
		_w4117_,
		_w14728_,
		_w14729_
	);
	LUT2 #(
		.INIT('h1)
	) name10683 (
		_w4121_,
		_w14726_,
		_w14730_
	);
	LUT2 #(
		.INIT('h4)
	) name10684 (
		_w14729_,
		_w14730_,
		_w14731_
	);
	LUT2 #(
		.INIT('h1)
	) name10685 (
		\memc_Dread_E_reg/NET0131 ,
		\memc_IOcmd_E_reg/NET0131 ,
		_w14732_
	);
	LUT2 #(
		.INIT('h4)
	) name10686 (
		\emc_EXTC_Eg_syn_reg/P0001 ,
		_w4068_,
		_w14733_
	);
	LUT2 #(
		.INIT('h2)
	) name10687 (
		_w5508_,
		_w14733_,
		_w14734_
	);
	LUT2 #(
		.INIT('h2)
	) name10688 (
		_w5432_,
		_w14732_,
		_w14735_
	);
	LUT2 #(
		.INIT('h8)
	) name10689 (
		_w14734_,
		_w14735_,
		_w14736_
	);
	LUT2 #(
		.INIT('h4)
	) name10690 (
		_w12441_,
		_w14736_,
		_w14737_
	);
	LUT2 #(
		.INIT('h2)
	) name10691 (
		\emc_DMDreg_reg[8]/P0001 ,
		_w14737_,
		_w14738_
	);
	LUT2 #(
		.INIT('h8)
	) name10692 (
		\T_ED[8]_pad ,
		_w14737_,
		_w14739_
	);
	LUT2 #(
		.INIT('h1)
	) name10693 (
		_w14738_,
		_w14739_,
		_w14740_
	);
	LUT2 #(
		.INIT('h2)
	) name10694 (
		\emc_DMDreg_reg[9]/P0001 ,
		_w14737_,
		_w14741_
	);
	LUT2 #(
		.INIT('h8)
	) name10695 (
		\T_ED[9]_pad ,
		_w14737_,
		_w14742_
	);
	LUT2 #(
		.INIT('h1)
	) name10696 (
		_w14741_,
		_w14742_,
		_w14743_
	);
	LUT2 #(
		.INIT('h8)
	) name10697 (
		\memc_Pread_E_reg/NET0131 ,
		_w5434_,
		_w14744_
	);
	LUT2 #(
		.INIT('h8)
	) name10698 (
		_w14734_,
		_w14744_,
		_w14745_
	);
	LUT2 #(
		.INIT('h2)
	) name10699 (
		\emc_PMDreg_reg[8]/P0001 ,
		_w14745_,
		_w14746_
	);
	LUT2 #(
		.INIT('h8)
	) name10700 (
		\T_ED[8]_pad ,
		_w14745_,
		_w14747_
	);
	LUT2 #(
		.INIT('h1)
	) name10701 (
		_w14746_,
		_w14747_,
		_w14748_
	);
	LUT2 #(
		.INIT('h2)
	) name10702 (
		\emc_PMDreg_reg[9]/P0001 ,
		_w14745_,
		_w14749_
	);
	LUT2 #(
		.INIT('h8)
	) name10703 (
		\T_ED[9]_pad ,
		_w14745_,
		_w14750_
	);
	LUT2 #(
		.INIT('h1)
	) name10704 (
		_w14749_,
		_w14750_,
		_w14751_
	);
	LUT2 #(
		.INIT('h8)
	) name10705 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w13804_,
		_w14752_
	);
	LUT2 #(
		.INIT('h4)
	) name10706 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14753_
	);
	LUT2 #(
		.INIT('h1)
	) name10707 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 ,
		_w14754_
	);
	LUT2 #(
		.INIT('h8)
	) name10708 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 ,
		_w14755_
	);
	LUT2 #(
		.INIT('h1)
	) name10709 (
		_w14754_,
		_w14755_,
		_w14756_
	);
	LUT2 #(
		.INIT('h4)
	) name10710 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w14756_,
		_w14757_
	);
	LUT2 #(
		.INIT('h8)
	) name10711 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14757_,
		_w14758_
	);
	LUT2 #(
		.INIT('h8)
	) name10712 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w14756_,
		_w14759_
	);
	LUT2 #(
		.INIT('h4)
	) name10713 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14759_,
		_w14760_
	);
	LUT2 #(
		.INIT('h1)
	) name10714 (
		_w14758_,
		_w14760_,
		_w14761_
	);
	LUT2 #(
		.INIT('h1)
	) name10715 (
		_w14753_,
		_w14761_,
		_w14762_
	);
	LUT2 #(
		.INIT('h4)
	) name10716 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14757_,
		_w14763_
	);
	LUT2 #(
		.INIT('h8)
	) name10717 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14759_,
		_w14764_
	);
	LUT2 #(
		.INIT('h1)
	) name10718 (
		_w14763_,
		_w14764_,
		_w14765_
	);
	LUT2 #(
		.INIT('h2)
	) name10719 (
		_w14753_,
		_w14765_,
		_w14766_
	);
	LUT2 #(
		.INIT('h1)
	) name10720 (
		_w14762_,
		_w14766_,
		_w14767_
	);
	LUT2 #(
		.INIT('h8)
	) name10721 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w14754_,
		_w14768_
	);
	LUT2 #(
		.INIT('h1)
	) name10722 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14768_,
		_w14769_
	);
	LUT2 #(
		.INIT('h4)
	) name10723 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w14755_,
		_w14770_
	);
	LUT2 #(
		.INIT('h2)
	) name10724 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14770_,
		_w14771_
	);
	LUT2 #(
		.INIT('h1)
	) name10725 (
		_w14769_,
		_w14771_,
		_w14772_
	);
	LUT2 #(
		.INIT('h4)
	) name10726 (
		_w14753_,
		_w14772_,
		_w14773_
	);
	LUT2 #(
		.INIT('h2)
	) name10727 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14768_,
		_w14774_
	);
	LUT2 #(
		.INIT('h1)
	) name10728 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14770_,
		_w14775_
	);
	LUT2 #(
		.INIT('h1)
	) name10729 (
		_w14774_,
		_w14775_,
		_w14776_
	);
	LUT2 #(
		.INIT('h8)
	) name10730 (
		_w14753_,
		_w14776_,
		_w14777_
	);
	LUT2 #(
		.INIT('h1)
	) name10731 (
		_w14773_,
		_w14777_,
		_w14778_
	);
	LUT2 #(
		.INIT('h8)
	) name10732 (
		_w14767_,
		_w14778_,
		_w14779_
	);
	LUT2 #(
		.INIT('h1)
	) name10733 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 ,
		_w14780_
	);
	LUT2 #(
		.INIT('h8)
	) name10734 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 ,
		_w14781_
	);
	LUT2 #(
		.INIT('h1)
	) name10735 (
		_w14780_,
		_w14781_,
		_w14782_
	);
	LUT2 #(
		.INIT('h4)
	) name10736 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w14782_,
		_w14783_
	);
	LUT2 #(
		.INIT('h8)
	) name10737 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14783_,
		_w14784_
	);
	LUT2 #(
		.INIT('h8)
	) name10738 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w14782_,
		_w14785_
	);
	LUT2 #(
		.INIT('h4)
	) name10739 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14785_,
		_w14786_
	);
	LUT2 #(
		.INIT('h1)
	) name10740 (
		_w14784_,
		_w14786_,
		_w14787_
	);
	LUT2 #(
		.INIT('h1)
	) name10741 (
		_w14753_,
		_w14787_,
		_w14788_
	);
	LUT2 #(
		.INIT('h4)
	) name10742 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14783_,
		_w14789_
	);
	LUT2 #(
		.INIT('h8)
	) name10743 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14785_,
		_w14790_
	);
	LUT2 #(
		.INIT('h1)
	) name10744 (
		_w14789_,
		_w14790_,
		_w14791_
	);
	LUT2 #(
		.INIT('h2)
	) name10745 (
		_w14753_,
		_w14791_,
		_w14792_
	);
	LUT2 #(
		.INIT('h1)
	) name10746 (
		_w14788_,
		_w14792_,
		_w14793_
	);
	LUT2 #(
		.INIT('h8)
	) name10747 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w14780_,
		_w14794_
	);
	LUT2 #(
		.INIT('h1)
	) name10748 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14794_,
		_w14795_
	);
	LUT2 #(
		.INIT('h4)
	) name10749 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w14781_,
		_w14796_
	);
	LUT2 #(
		.INIT('h2)
	) name10750 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14796_,
		_w14797_
	);
	LUT2 #(
		.INIT('h1)
	) name10751 (
		_w14795_,
		_w14797_,
		_w14798_
	);
	LUT2 #(
		.INIT('h4)
	) name10752 (
		_w14753_,
		_w14798_,
		_w14799_
	);
	LUT2 #(
		.INIT('h2)
	) name10753 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14794_,
		_w14800_
	);
	LUT2 #(
		.INIT('h1)
	) name10754 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14796_,
		_w14801_
	);
	LUT2 #(
		.INIT('h1)
	) name10755 (
		_w14800_,
		_w14801_,
		_w14802_
	);
	LUT2 #(
		.INIT('h8)
	) name10756 (
		_w14753_,
		_w14802_,
		_w14803_
	);
	LUT2 #(
		.INIT('h1)
	) name10757 (
		_w14799_,
		_w14803_,
		_w14804_
	);
	LUT2 #(
		.INIT('h8)
	) name10758 (
		_w14793_,
		_w14804_,
		_w14805_
	);
	LUT2 #(
		.INIT('h8)
	) name10759 (
		_w14779_,
		_w14805_,
		_w14806_
	);
	LUT2 #(
		.INIT('h8)
	) name10760 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 ,
		_w14807_
	);
	LUT2 #(
		.INIT('h1)
	) name10761 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 ,
		_w14808_
	);
	LUT2 #(
		.INIT('h1)
	) name10762 (
		_w14807_,
		_w14808_,
		_w14809_
	);
	LUT2 #(
		.INIT('h4)
	) name10763 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w14809_,
		_w14810_
	);
	LUT2 #(
		.INIT('h8)
	) name10764 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14810_,
		_w14811_
	);
	LUT2 #(
		.INIT('h8)
	) name10765 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w14809_,
		_w14812_
	);
	LUT2 #(
		.INIT('h4)
	) name10766 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14812_,
		_w14813_
	);
	LUT2 #(
		.INIT('h1)
	) name10767 (
		_w14811_,
		_w14813_,
		_w14814_
	);
	LUT2 #(
		.INIT('h1)
	) name10768 (
		_w14753_,
		_w14814_,
		_w14815_
	);
	LUT2 #(
		.INIT('h8)
	) name10769 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14812_,
		_w14816_
	);
	LUT2 #(
		.INIT('h4)
	) name10770 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14810_,
		_w14817_
	);
	LUT2 #(
		.INIT('h1)
	) name10771 (
		_w14816_,
		_w14817_,
		_w14818_
	);
	LUT2 #(
		.INIT('h2)
	) name10772 (
		_w14753_,
		_w14818_,
		_w14819_
	);
	LUT2 #(
		.INIT('h1)
	) name10773 (
		_w14815_,
		_w14819_,
		_w14820_
	);
	LUT2 #(
		.INIT('h8)
	) name10774 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w14808_,
		_w14821_
	);
	LUT2 #(
		.INIT('h1)
	) name10775 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14821_,
		_w14822_
	);
	LUT2 #(
		.INIT('h4)
	) name10776 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w14807_,
		_w14823_
	);
	LUT2 #(
		.INIT('h2)
	) name10777 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14823_,
		_w14824_
	);
	LUT2 #(
		.INIT('h1)
	) name10778 (
		_w14822_,
		_w14824_,
		_w14825_
	);
	LUT2 #(
		.INIT('h4)
	) name10779 (
		_w14753_,
		_w14825_,
		_w14826_
	);
	LUT2 #(
		.INIT('h1)
	) name10780 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14823_,
		_w14827_
	);
	LUT2 #(
		.INIT('h2)
	) name10781 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14821_,
		_w14828_
	);
	LUT2 #(
		.INIT('h1)
	) name10782 (
		_w14827_,
		_w14828_,
		_w14829_
	);
	LUT2 #(
		.INIT('h8)
	) name10783 (
		_w14753_,
		_w14829_,
		_w14830_
	);
	LUT2 #(
		.INIT('h1)
	) name10784 (
		_w14826_,
		_w14830_,
		_w14831_
	);
	LUT2 #(
		.INIT('h8)
	) name10785 (
		_w14820_,
		_w14831_,
		_w14832_
	);
	LUT2 #(
		.INIT('h8)
	) name10786 (
		_w14806_,
		_w14832_,
		_w14833_
	);
	LUT2 #(
		.INIT('h8)
	) name10787 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w14834_
	);
	LUT2 #(
		.INIT('h4)
	) name10788 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14834_,
		_w14835_
	);
	LUT2 #(
		.INIT('h2)
	) name10789 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w14836_
	);
	LUT2 #(
		.INIT('h8)
	) name10790 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14836_,
		_w14837_
	);
	LUT2 #(
		.INIT('h1)
	) name10791 (
		_w14835_,
		_w14837_,
		_w14838_
	);
	LUT2 #(
		.INIT('h1)
	) name10792 (
		_w14753_,
		_w14838_,
		_w14839_
	);
	LUT2 #(
		.INIT('h8)
	) name10793 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14834_,
		_w14840_
	);
	LUT2 #(
		.INIT('h4)
	) name10794 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14836_,
		_w14841_
	);
	LUT2 #(
		.INIT('h1)
	) name10795 (
		_w14840_,
		_w14841_,
		_w14842_
	);
	LUT2 #(
		.INIT('h2)
	) name10796 (
		_w14753_,
		_w14842_,
		_w14843_
	);
	LUT2 #(
		.INIT('h1)
	) name10797 (
		_w14839_,
		_w14843_,
		_w14844_
	);
	LUT2 #(
		.INIT('h1)
	) name10798 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		_w14845_
	);
	LUT2 #(
		.INIT('h8)
	) name10799 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w14845_,
		_w14846_
	);
	LUT2 #(
		.INIT('h4)
	) name10800 (
		_w14753_,
		_w14846_,
		_w14847_
	);
	LUT2 #(
		.INIT('h2)
	) name10801 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		_w14848_
	);
	LUT2 #(
		.INIT('h8)
	) name10802 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w14848_,
		_w14849_
	);
	LUT2 #(
		.INIT('h8)
	) name10803 (
		_w14753_,
		_w14849_,
		_w14850_
	);
	LUT2 #(
		.INIT('h1)
	) name10804 (
		_w14847_,
		_w14850_,
		_w14851_
	);
	LUT2 #(
		.INIT('h8)
	) name10805 (
		_w14844_,
		_w14851_,
		_w14852_
	);
	LUT2 #(
		.INIT('h8)
	) name10806 (
		_w14833_,
		_w14852_,
		_w14853_
	);
	LUT2 #(
		.INIT('h1)
	) name10807 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		_w14854_
	);
	LUT2 #(
		.INIT('h8)
	) name10808 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		_w14855_
	);
	LUT2 #(
		.INIT('h1)
	) name10809 (
		_w14854_,
		_w14855_,
		_w14856_
	);
	LUT2 #(
		.INIT('h4)
	) name10810 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w14856_,
		_w14857_
	);
	LUT2 #(
		.INIT('h8)
	) name10811 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14857_,
		_w14858_
	);
	LUT2 #(
		.INIT('h8)
	) name10812 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w14856_,
		_w14859_
	);
	LUT2 #(
		.INIT('h4)
	) name10813 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14859_,
		_w14860_
	);
	LUT2 #(
		.INIT('h1)
	) name10814 (
		_w14858_,
		_w14860_,
		_w14861_
	);
	LUT2 #(
		.INIT('h1)
	) name10815 (
		_w14753_,
		_w14861_,
		_w14862_
	);
	LUT2 #(
		.INIT('h4)
	) name10816 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14857_,
		_w14863_
	);
	LUT2 #(
		.INIT('h8)
	) name10817 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14859_,
		_w14864_
	);
	LUT2 #(
		.INIT('h1)
	) name10818 (
		_w14863_,
		_w14864_,
		_w14865_
	);
	LUT2 #(
		.INIT('h2)
	) name10819 (
		_w14753_,
		_w14865_,
		_w14866_
	);
	LUT2 #(
		.INIT('h1)
	) name10820 (
		_w14862_,
		_w14866_,
		_w14867_
	);
	LUT2 #(
		.INIT('h8)
	) name10821 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w14854_,
		_w14868_
	);
	LUT2 #(
		.INIT('h1)
	) name10822 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14868_,
		_w14869_
	);
	LUT2 #(
		.INIT('h4)
	) name10823 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w14855_,
		_w14870_
	);
	LUT2 #(
		.INIT('h2)
	) name10824 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14870_,
		_w14871_
	);
	LUT2 #(
		.INIT('h1)
	) name10825 (
		_w14869_,
		_w14871_,
		_w14872_
	);
	LUT2 #(
		.INIT('h4)
	) name10826 (
		_w14753_,
		_w14872_,
		_w14873_
	);
	LUT2 #(
		.INIT('h2)
	) name10827 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14868_,
		_w14874_
	);
	LUT2 #(
		.INIT('h1)
	) name10828 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14870_,
		_w14875_
	);
	LUT2 #(
		.INIT('h1)
	) name10829 (
		_w14874_,
		_w14875_,
		_w14876_
	);
	LUT2 #(
		.INIT('h8)
	) name10830 (
		_w14753_,
		_w14876_,
		_w14877_
	);
	LUT2 #(
		.INIT('h1)
	) name10831 (
		_w14873_,
		_w14877_,
		_w14878_
	);
	LUT2 #(
		.INIT('h8)
	) name10832 (
		_w14867_,
		_w14878_,
		_w14879_
	);
	LUT2 #(
		.INIT('h1)
	) name10833 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w14880_
	);
	LUT2 #(
		.INIT('h8)
	) name10834 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w14881_
	);
	LUT2 #(
		.INIT('h1)
	) name10835 (
		_w14880_,
		_w14881_,
		_w14882_
	);
	LUT2 #(
		.INIT('h4)
	) name10836 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		_w14882_,
		_w14883_
	);
	LUT2 #(
		.INIT('h8)
	) name10837 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14883_,
		_w14884_
	);
	LUT2 #(
		.INIT('h8)
	) name10838 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		_w14882_,
		_w14885_
	);
	LUT2 #(
		.INIT('h4)
	) name10839 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14885_,
		_w14886_
	);
	LUT2 #(
		.INIT('h1)
	) name10840 (
		_w14884_,
		_w14886_,
		_w14887_
	);
	LUT2 #(
		.INIT('h1)
	) name10841 (
		_w14753_,
		_w14887_,
		_w14888_
	);
	LUT2 #(
		.INIT('h4)
	) name10842 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14883_,
		_w14889_
	);
	LUT2 #(
		.INIT('h8)
	) name10843 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14885_,
		_w14890_
	);
	LUT2 #(
		.INIT('h1)
	) name10844 (
		_w14889_,
		_w14890_,
		_w14891_
	);
	LUT2 #(
		.INIT('h2)
	) name10845 (
		_w14753_,
		_w14891_,
		_w14892_
	);
	LUT2 #(
		.INIT('h1)
	) name10846 (
		_w14888_,
		_w14892_,
		_w14893_
	);
	LUT2 #(
		.INIT('h8)
	) name10847 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		_w14880_,
		_w14894_
	);
	LUT2 #(
		.INIT('h1)
	) name10848 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14894_,
		_w14895_
	);
	LUT2 #(
		.INIT('h4)
	) name10849 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		_w14881_,
		_w14896_
	);
	LUT2 #(
		.INIT('h2)
	) name10850 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14896_,
		_w14897_
	);
	LUT2 #(
		.INIT('h1)
	) name10851 (
		_w14895_,
		_w14897_,
		_w14898_
	);
	LUT2 #(
		.INIT('h4)
	) name10852 (
		_w14753_,
		_w14898_,
		_w14899_
	);
	LUT2 #(
		.INIT('h2)
	) name10853 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14894_,
		_w14900_
	);
	LUT2 #(
		.INIT('h1)
	) name10854 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14896_,
		_w14901_
	);
	LUT2 #(
		.INIT('h1)
	) name10855 (
		_w14900_,
		_w14901_,
		_w14902_
	);
	LUT2 #(
		.INIT('h8)
	) name10856 (
		_w14753_,
		_w14902_,
		_w14903_
	);
	LUT2 #(
		.INIT('h1)
	) name10857 (
		_w14899_,
		_w14903_,
		_w14904_
	);
	LUT2 #(
		.INIT('h8)
	) name10858 (
		_w14893_,
		_w14904_,
		_w14905_
	);
	LUT2 #(
		.INIT('h8)
	) name10859 (
		_w14879_,
		_w14905_,
		_w14906_
	);
	LUT2 #(
		.INIT('h8)
	) name10860 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 ,
		_w14907_
	);
	LUT2 #(
		.INIT('h1)
	) name10861 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 ,
		_w14908_
	);
	LUT2 #(
		.INIT('h1)
	) name10862 (
		_w14907_,
		_w14908_,
		_w14909_
	);
	LUT2 #(
		.INIT('h4)
	) name10863 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w14909_,
		_w14910_
	);
	LUT2 #(
		.INIT('h8)
	) name10864 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14910_,
		_w14911_
	);
	LUT2 #(
		.INIT('h8)
	) name10865 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w14909_,
		_w14912_
	);
	LUT2 #(
		.INIT('h4)
	) name10866 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14912_,
		_w14913_
	);
	LUT2 #(
		.INIT('h1)
	) name10867 (
		_w14911_,
		_w14913_,
		_w14914_
	);
	LUT2 #(
		.INIT('h1)
	) name10868 (
		_w14753_,
		_w14914_,
		_w14915_
	);
	LUT2 #(
		.INIT('h8)
	) name10869 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14912_,
		_w14916_
	);
	LUT2 #(
		.INIT('h4)
	) name10870 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14910_,
		_w14917_
	);
	LUT2 #(
		.INIT('h1)
	) name10871 (
		_w14916_,
		_w14917_,
		_w14918_
	);
	LUT2 #(
		.INIT('h2)
	) name10872 (
		_w14753_,
		_w14918_,
		_w14919_
	);
	LUT2 #(
		.INIT('h1)
	) name10873 (
		_w14915_,
		_w14919_,
		_w14920_
	);
	LUT2 #(
		.INIT('h8)
	) name10874 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w14908_,
		_w14921_
	);
	LUT2 #(
		.INIT('h1)
	) name10875 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14921_,
		_w14922_
	);
	LUT2 #(
		.INIT('h4)
	) name10876 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w14907_,
		_w14923_
	);
	LUT2 #(
		.INIT('h2)
	) name10877 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14923_,
		_w14924_
	);
	LUT2 #(
		.INIT('h1)
	) name10878 (
		_w14922_,
		_w14924_,
		_w14925_
	);
	LUT2 #(
		.INIT('h4)
	) name10879 (
		_w14753_,
		_w14925_,
		_w14926_
	);
	LUT2 #(
		.INIT('h1)
	) name10880 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14923_,
		_w14927_
	);
	LUT2 #(
		.INIT('h2)
	) name10881 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14921_,
		_w14928_
	);
	LUT2 #(
		.INIT('h1)
	) name10882 (
		_w14927_,
		_w14928_,
		_w14929_
	);
	LUT2 #(
		.INIT('h8)
	) name10883 (
		_w14753_,
		_w14929_,
		_w14930_
	);
	LUT2 #(
		.INIT('h1)
	) name10884 (
		_w14926_,
		_w14930_,
		_w14931_
	);
	LUT2 #(
		.INIT('h8)
	) name10885 (
		_w14920_,
		_w14931_,
		_w14932_
	);
	LUT2 #(
		.INIT('h8)
	) name10886 (
		_w14906_,
		_w14932_,
		_w14933_
	);
	LUT2 #(
		.INIT('h2)
	) name10887 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w7473_,
		_w14934_
	);
	LUT2 #(
		.INIT('h2)
	) name10888 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14934_,
		_w14935_
	);
	LUT2 #(
		.INIT('h2)
	) name10889 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w9229_,
		_w14936_
	);
	LUT2 #(
		.INIT('h1)
	) name10890 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14936_,
		_w14937_
	);
	LUT2 #(
		.INIT('h1)
	) name10891 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w14935_,
		_w14938_
	);
	LUT2 #(
		.INIT('h4)
	) name10892 (
		_w14937_,
		_w14938_,
		_w14939_
	);
	LUT2 #(
		.INIT('h1)
	) name10893 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 ,
		_w14940_
	);
	LUT2 #(
		.INIT('h8)
	) name10894 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 ,
		_w14941_
	);
	LUT2 #(
		.INIT('h1)
	) name10895 (
		_w14940_,
		_w14941_,
		_w14942_
	);
	LUT2 #(
		.INIT('h4)
	) name10896 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w14942_,
		_w14943_
	);
	LUT2 #(
		.INIT('h8)
	) name10897 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14943_,
		_w14944_
	);
	LUT2 #(
		.INIT('h8)
	) name10898 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w14942_,
		_w14945_
	);
	LUT2 #(
		.INIT('h4)
	) name10899 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14945_,
		_w14946_
	);
	LUT2 #(
		.INIT('h1)
	) name10900 (
		_w14944_,
		_w14946_,
		_w14947_
	);
	LUT2 #(
		.INIT('h1)
	) name10901 (
		_w14753_,
		_w14947_,
		_w14948_
	);
	LUT2 #(
		.INIT('h4)
	) name10902 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14943_,
		_w14949_
	);
	LUT2 #(
		.INIT('h8)
	) name10903 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14945_,
		_w14950_
	);
	LUT2 #(
		.INIT('h1)
	) name10904 (
		_w14949_,
		_w14950_,
		_w14951_
	);
	LUT2 #(
		.INIT('h2)
	) name10905 (
		_w14753_,
		_w14951_,
		_w14952_
	);
	LUT2 #(
		.INIT('h1)
	) name10906 (
		_w14948_,
		_w14952_,
		_w14953_
	);
	LUT2 #(
		.INIT('h8)
	) name10907 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w14940_,
		_w14954_
	);
	LUT2 #(
		.INIT('h1)
	) name10908 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14954_,
		_w14955_
	);
	LUT2 #(
		.INIT('h4)
	) name10909 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w14941_,
		_w14956_
	);
	LUT2 #(
		.INIT('h2)
	) name10910 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14956_,
		_w14957_
	);
	LUT2 #(
		.INIT('h1)
	) name10911 (
		_w14955_,
		_w14957_,
		_w14958_
	);
	LUT2 #(
		.INIT('h4)
	) name10912 (
		_w14753_,
		_w14958_,
		_w14959_
	);
	LUT2 #(
		.INIT('h2)
	) name10913 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14954_,
		_w14960_
	);
	LUT2 #(
		.INIT('h1)
	) name10914 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14956_,
		_w14961_
	);
	LUT2 #(
		.INIT('h1)
	) name10915 (
		_w14960_,
		_w14961_,
		_w14962_
	);
	LUT2 #(
		.INIT('h8)
	) name10916 (
		_w14753_,
		_w14962_,
		_w14963_
	);
	LUT2 #(
		.INIT('h1)
	) name10917 (
		_w14959_,
		_w14963_,
		_w14964_
	);
	LUT2 #(
		.INIT('h8)
	) name10918 (
		_w14953_,
		_w14964_,
		_w14965_
	);
	LUT2 #(
		.INIT('h8)
	) name10919 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w14966_
	);
	LUT2 #(
		.INIT('h8)
	) name10920 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14966_,
		_w14967_
	);
	LUT2 #(
		.INIT('h4)
	) name10921 (
		_w14753_,
		_w14967_,
		_w14968_
	);
	LUT2 #(
		.INIT('h4)
	) name10922 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w14966_,
		_w14969_
	);
	LUT2 #(
		.INIT('h8)
	) name10923 (
		_w14753_,
		_w14969_,
		_w14970_
	);
	LUT2 #(
		.INIT('h1)
	) name10924 (
		_w14968_,
		_w14970_,
		_w14971_
	);
	LUT2 #(
		.INIT('h8)
	) name10925 (
		_w14965_,
		_w14971_,
		_w14972_
	);
	LUT2 #(
		.INIT('h4)
	) name10926 (
		_w14939_,
		_w14972_,
		_w14973_
	);
	LUT2 #(
		.INIT('h2)
	) name10927 (
		_w14939_,
		_w14972_,
		_w14974_
	);
	LUT2 #(
		.INIT('h1)
	) name10928 (
		_w14973_,
		_w14974_,
		_w14975_
	);
	LUT2 #(
		.INIT('h1)
	) name10929 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14967_,
		_w14976_
	);
	LUT2 #(
		.INIT('h2)
	) name10930 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14969_,
		_w14977_
	);
	LUT2 #(
		.INIT('h1)
	) name10931 (
		_w14976_,
		_w14977_,
		_w14978_
	);
	LUT2 #(
		.INIT('h2)
	) name10932 (
		_w14965_,
		_w14978_,
		_w14979_
	);
	LUT2 #(
		.INIT('h4)
	) name10933 (
		_w14965_,
		_w14978_,
		_w14980_
	);
	LUT2 #(
		.INIT('h2)
	) name10934 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w12028_,
		_w14981_
	);
	LUT2 #(
		.INIT('h2)
	) name10935 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14981_,
		_w14982_
	);
	LUT2 #(
		.INIT('h1)
	) name10936 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14934_,
		_w14983_
	);
	LUT2 #(
		.INIT('h1)
	) name10937 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w14982_,
		_w14984_
	);
	LUT2 #(
		.INIT('h4)
	) name10938 (
		_w14983_,
		_w14984_,
		_w14985_
	);
	LUT2 #(
		.INIT('h1)
	) name10939 (
		_w14980_,
		_w14985_,
		_w14986_
	);
	LUT2 #(
		.INIT('h1)
	) name10940 (
		_w14979_,
		_w14986_,
		_w14987_
	);
	LUT2 #(
		.INIT('h1)
	) name10941 (
		_w14975_,
		_w14987_,
		_w14988_
	);
	LUT2 #(
		.INIT('h1)
	) name10942 (
		_w14933_,
		_w14988_,
		_w14989_
	);
	LUT2 #(
		.INIT('h1)
	) name10943 (
		_w14879_,
		_w14905_,
		_w14990_
	);
	LUT2 #(
		.INIT('h4)
	) name10944 (
		_w14932_,
		_w14990_,
		_w14991_
	);
	LUT2 #(
		.INIT('h1)
	) name10945 (
		_w14933_,
		_w14991_,
		_w14992_
	);
	LUT2 #(
		.INIT('h2)
	) name10946 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14993_
	);
	LUT2 #(
		.INIT('h4)
	) name10947 (
		_w8534_,
		_w14993_,
		_w14994_
	);
	LUT2 #(
		.INIT('h8)
	) name10948 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14936_,
		_w14995_
	);
	LUT2 #(
		.INIT('h1)
	) name10949 (
		_w14994_,
		_w14995_,
		_w14996_
	);
	LUT2 #(
		.INIT('h1)
	) name10950 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w14996_,
		_w14997_
	);
	LUT2 #(
		.INIT('h2)
	) name10951 (
		_w14972_,
		_w14997_,
		_w14998_
	);
	LUT2 #(
		.INIT('h4)
	) name10952 (
		_w14972_,
		_w14997_,
		_w14999_
	);
	LUT2 #(
		.INIT('h1)
	) name10953 (
		_w14998_,
		_w14999_,
		_w15000_
	);
	LUT2 #(
		.INIT('h1)
	) name10954 (
		_w14974_,
		_w15000_,
		_w15001_
	);
	LUT2 #(
		.INIT('h2)
	) name10955 (
		_w14974_,
		_w14997_,
		_w15002_
	);
	LUT2 #(
		.INIT('h1)
	) name10956 (
		_w15001_,
		_w15002_,
		_w15003_
	);
	LUT2 #(
		.INIT('h2)
	) name10957 (
		_w14992_,
		_w15003_,
		_w15004_
	);
	LUT2 #(
		.INIT('h4)
	) name10958 (
		_w14992_,
		_w15003_,
		_w15005_
	);
	LUT2 #(
		.INIT('h1)
	) name10959 (
		_w15004_,
		_w15005_,
		_w15006_
	);
	LUT2 #(
		.INIT('h1)
	) name10960 (
		_w14989_,
		_w15006_,
		_w15007_
	);
	LUT2 #(
		.INIT('h8)
	) name10961 (
		_w14989_,
		_w15006_,
		_w15008_
	);
	LUT2 #(
		.INIT('h1)
	) name10962 (
		_w15007_,
		_w15008_,
		_w15009_
	);
	LUT2 #(
		.INIT('h1)
	) name10963 (
		_w14979_,
		_w14980_,
		_w15010_
	);
	LUT2 #(
		.INIT('h2)
	) name10964 (
		_w14985_,
		_w15010_,
		_w15011_
	);
	LUT2 #(
		.INIT('h4)
	) name10965 (
		_w14985_,
		_w15010_,
		_w15012_
	);
	LUT2 #(
		.INIT('h1)
	) name10966 (
		_w15011_,
		_w15012_,
		_w15013_
	);
	LUT2 #(
		.INIT('h1)
	) name10967 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14967_,
		_w15014_
	);
	LUT2 #(
		.INIT('h2)
	) name10968 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14969_,
		_w15015_
	);
	LUT2 #(
		.INIT('h1)
	) name10969 (
		_w15014_,
		_w15015_,
		_w15016_
	);
	LUT2 #(
		.INIT('h4)
	) name10970 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14958_,
		_w15017_
	);
	LUT2 #(
		.INIT('h8)
	) name10971 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14962_,
		_w15018_
	);
	LUT2 #(
		.INIT('h1)
	) name10972 (
		_w15017_,
		_w15018_,
		_w15019_
	);
	LUT2 #(
		.INIT('h8)
	) name10973 (
		_w14953_,
		_w15019_,
		_w15020_
	);
	LUT2 #(
		.INIT('h4)
	) name10974 (
		_w15016_,
		_w15020_,
		_w15021_
	);
	LUT2 #(
		.INIT('h2)
	) name10975 (
		_w15016_,
		_w15020_,
		_w15022_
	);
	LUT2 #(
		.INIT('h2)
	) name10976 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w11882_,
		_w15023_
	);
	LUT2 #(
		.INIT('h2)
	) name10977 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15023_,
		_w15024_
	);
	LUT2 #(
		.INIT('h1)
	) name10978 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w14981_,
		_w15025_
	);
	LUT2 #(
		.INIT('h1)
	) name10979 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15024_,
		_w15026_
	);
	LUT2 #(
		.INIT('h4)
	) name10980 (
		_w15025_,
		_w15026_,
		_w15027_
	);
	LUT2 #(
		.INIT('h1)
	) name10981 (
		_w15022_,
		_w15027_,
		_w15028_
	);
	LUT2 #(
		.INIT('h1)
	) name10982 (
		_w15021_,
		_w15028_,
		_w15029_
	);
	LUT2 #(
		.INIT('h2)
	) name10983 (
		_w15013_,
		_w15029_,
		_w15030_
	);
	LUT2 #(
		.INIT('h1)
	) name10984 (
		_w14933_,
		_w15030_,
		_w15031_
	);
	LUT2 #(
		.INIT('h8)
	) name10985 (
		_w14975_,
		_w14987_,
		_w15032_
	);
	LUT2 #(
		.INIT('h1)
	) name10986 (
		_w14988_,
		_w15032_,
		_w15033_
	);
	LUT2 #(
		.INIT('h8)
	) name10987 (
		_w14992_,
		_w15033_,
		_w15034_
	);
	LUT2 #(
		.INIT('h1)
	) name10988 (
		_w14992_,
		_w15033_,
		_w15035_
	);
	LUT2 #(
		.INIT('h1)
	) name10989 (
		_w15034_,
		_w15035_,
		_w15036_
	);
	LUT2 #(
		.INIT('h4)
	) name10990 (
		_w15031_,
		_w15036_,
		_w15037_
	);
	LUT2 #(
		.INIT('h1)
	) name10991 (
		_w14991_,
		_w15032_,
		_w15038_
	);
	LUT2 #(
		.INIT('h4)
	) name10992 (
		_w15036_,
		_w15038_,
		_w15039_
	);
	LUT2 #(
		.INIT('h1)
	) name10993 (
		_w15037_,
		_w15039_,
		_w15040_
	);
	LUT2 #(
		.INIT('h2)
	) name10994 (
		_w15009_,
		_w15040_,
		_w15041_
	);
	LUT2 #(
		.INIT('h1)
	) name10995 (
		_w14853_,
		_w15041_,
		_w15042_
	);
	LUT2 #(
		.INIT('h1)
	) name10996 (
		_w14933_,
		_w15001_,
		_w15043_
	);
	LUT2 #(
		.INIT('h8)
	) name10997 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15044_
	);
	LUT2 #(
		.INIT('h4)
	) name10998 (
		_w8534_,
		_w15044_,
		_w15045_
	);
	LUT2 #(
		.INIT('h2)
	) name10999 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w7905_,
		_w15046_
	);
	LUT2 #(
		.INIT('h4)
	) name11000 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15046_,
		_w15047_
	);
	LUT2 #(
		.INIT('h1)
	) name11001 (
		_w15045_,
		_w15047_,
		_w15048_
	);
	LUT2 #(
		.INIT('h1)
	) name11002 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15048_,
		_w15049_
	);
	LUT2 #(
		.INIT('h2)
	) name11003 (
		_w14972_,
		_w15049_,
		_w15050_
	);
	LUT2 #(
		.INIT('h4)
	) name11004 (
		_w14972_,
		_w15049_,
		_w15051_
	);
	LUT2 #(
		.INIT('h1)
	) name11005 (
		_w15050_,
		_w15051_,
		_w15052_
	);
	LUT2 #(
		.INIT('h1)
	) name11006 (
		_w14999_,
		_w15052_,
		_w15053_
	);
	LUT2 #(
		.INIT('h8)
	) name11007 (
		_w14999_,
		_w15048_,
		_w15054_
	);
	LUT2 #(
		.INIT('h1)
	) name11008 (
		_w15053_,
		_w15054_,
		_w15055_
	);
	LUT2 #(
		.INIT('h2)
	) name11009 (
		_w14992_,
		_w15055_,
		_w15056_
	);
	LUT2 #(
		.INIT('h4)
	) name11010 (
		_w14992_,
		_w15055_,
		_w15057_
	);
	LUT2 #(
		.INIT('h1)
	) name11011 (
		_w15056_,
		_w15057_,
		_w15058_
	);
	LUT2 #(
		.INIT('h1)
	) name11012 (
		_w15043_,
		_w15058_,
		_w15059_
	);
	LUT2 #(
		.INIT('h8)
	) name11013 (
		_w15043_,
		_w15058_,
		_w15060_
	);
	LUT2 #(
		.INIT('h1)
	) name11014 (
		_w15059_,
		_w15060_,
		_w15061_
	);
	LUT2 #(
		.INIT('h1)
	) name11015 (
		_w14991_,
		_w15002_,
		_w15062_
	);
	LUT2 #(
		.INIT('h8)
	) name11016 (
		_w15006_,
		_w15062_,
		_w15063_
	);
	LUT2 #(
		.INIT('h1)
	) name11017 (
		_w15007_,
		_w15063_,
		_w15064_
	);
	LUT2 #(
		.INIT('h2)
	) name11018 (
		_w15061_,
		_w15064_,
		_w15065_
	);
	LUT2 #(
		.INIT('h4)
	) name11019 (
		_w15061_,
		_w15064_,
		_w15066_
	);
	LUT2 #(
		.INIT('h1)
	) name11020 (
		_w15065_,
		_w15066_,
		_w15067_
	);
	LUT2 #(
		.INIT('h2)
	) name11021 (
		_w14853_,
		_w15067_,
		_w15068_
	);
	LUT2 #(
		.INIT('h4)
	) name11022 (
		_w14853_,
		_w15067_,
		_w15069_
	);
	LUT2 #(
		.INIT('h1)
	) name11023 (
		_w15068_,
		_w15069_,
		_w15070_
	);
	LUT2 #(
		.INIT('h4)
	) name11024 (
		_w15042_,
		_w15070_,
		_w15071_
	);
	LUT2 #(
		.INIT('h4)
	) name11025 (
		_w15041_,
		_w15069_,
		_w15072_
	);
	LUT2 #(
		.INIT('h1)
	) name11026 (
		_w15071_,
		_w15072_,
		_w15073_
	);
	LUT2 #(
		.INIT('h2)
	) name11027 (
		_w15031_,
		_w15036_,
		_w15074_
	);
	LUT2 #(
		.INIT('h1)
	) name11028 (
		_w15037_,
		_w15074_,
		_w15075_
	);
	LUT2 #(
		.INIT('h1)
	) name11029 (
		_w15021_,
		_w15022_,
		_w15076_
	);
	LUT2 #(
		.INIT('h2)
	) name11030 (
		_w15027_,
		_w15076_,
		_w15077_
	);
	LUT2 #(
		.INIT('h4)
	) name11031 (
		_w15027_,
		_w15076_,
		_w15078_
	);
	LUT2 #(
		.INIT('h1)
	) name11032 (
		_w15077_,
		_w15078_,
		_w15079_
	);
	LUT2 #(
		.INIT('h1)
	) name11033 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14967_,
		_w15080_
	);
	LUT2 #(
		.INIT('h2)
	) name11034 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14969_,
		_w15081_
	);
	LUT2 #(
		.INIT('h1)
	) name11035 (
		_w15080_,
		_w15081_,
		_w15082_
	);
	LUT2 #(
		.INIT('h1)
	) name11036 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14947_,
		_w15083_
	);
	LUT2 #(
		.INIT('h2)
	) name11037 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14951_,
		_w15084_
	);
	LUT2 #(
		.INIT('h4)
	) name11038 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14958_,
		_w15085_
	);
	LUT2 #(
		.INIT('h8)
	) name11039 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14962_,
		_w15086_
	);
	LUT2 #(
		.INIT('h1)
	) name11040 (
		_w15085_,
		_w15086_,
		_w15087_
	);
	LUT2 #(
		.INIT('h4)
	) name11041 (
		_w15083_,
		_w15087_,
		_w15088_
	);
	LUT2 #(
		.INIT('h4)
	) name11042 (
		_w15084_,
		_w15088_,
		_w15089_
	);
	LUT2 #(
		.INIT('h4)
	) name11043 (
		_w15082_,
		_w15089_,
		_w15090_
	);
	LUT2 #(
		.INIT('h2)
	) name11044 (
		_w15082_,
		_w15089_,
		_w15091_
	);
	LUT2 #(
		.INIT('h2)
	) name11045 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w7202_,
		_w15092_
	);
	LUT2 #(
		.INIT('h2)
	) name11046 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15092_,
		_w15093_
	);
	LUT2 #(
		.INIT('h1)
	) name11047 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15023_,
		_w15094_
	);
	LUT2 #(
		.INIT('h1)
	) name11048 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15093_,
		_w15095_
	);
	LUT2 #(
		.INIT('h4)
	) name11049 (
		_w15094_,
		_w15095_,
		_w15096_
	);
	LUT2 #(
		.INIT('h1)
	) name11050 (
		_w15091_,
		_w15096_,
		_w15097_
	);
	LUT2 #(
		.INIT('h1)
	) name11051 (
		_w15090_,
		_w15097_,
		_w15098_
	);
	LUT2 #(
		.INIT('h2)
	) name11052 (
		_w15079_,
		_w15098_,
		_w15099_
	);
	LUT2 #(
		.INIT('h1)
	) name11053 (
		_w14933_,
		_w15099_,
		_w15100_
	);
	LUT2 #(
		.INIT('h4)
	) name11054 (
		_w15013_,
		_w15029_,
		_w15101_
	);
	LUT2 #(
		.INIT('h1)
	) name11055 (
		_w15030_,
		_w15101_,
		_w15102_
	);
	LUT2 #(
		.INIT('h2)
	) name11056 (
		_w14992_,
		_w15102_,
		_w15103_
	);
	LUT2 #(
		.INIT('h4)
	) name11057 (
		_w14992_,
		_w15102_,
		_w15104_
	);
	LUT2 #(
		.INIT('h1)
	) name11058 (
		_w15103_,
		_w15104_,
		_w15105_
	);
	LUT2 #(
		.INIT('h1)
	) name11059 (
		_w15100_,
		_w15105_,
		_w15106_
	);
	LUT2 #(
		.INIT('h1)
	) name11060 (
		_w14991_,
		_w15101_,
		_w15107_
	);
	LUT2 #(
		.INIT('h8)
	) name11061 (
		_w15105_,
		_w15107_,
		_w15108_
	);
	LUT2 #(
		.INIT('h1)
	) name11062 (
		_w15106_,
		_w15108_,
		_w15109_
	);
	LUT2 #(
		.INIT('h2)
	) name11063 (
		_w15075_,
		_w15109_,
		_w15110_
	);
	LUT2 #(
		.INIT('h1)
	) name11064 (
		_w14853_,
		_w15110_,
		_w15111_
	);
	LUT2 #(
		.INIT('h4)
	) name11065 (
		_w15009_,
		_w15040_,
		_w15112_
	);
	LUT2 #(
		.INIT('h1)
	) name11066 (
		_w15041_,
		_w15112_,
		_w15113_
	);
	LUT2 #(
		.INIT('h8)
	) name11067 (
		_w14853_,
		_w15113_,
		_w15114_
	);
	LUT2 #(
		.INIT('h1)
	) name11068 (
		_w14853_,
		_w15113_,
		_w15115_
	);
	LUT2 #(
		.INIT('h1)
	) name11069 (
		_w15114_,
		_w15115_,
		_w15116_
	);
	LUT2 #(
		.INIT('h1)
	) name11070 (
		_w15111_,
		_w15116_,
		_w15117_
	);
	LUT2 #(
		.INIT('h4)
	) name11071 (
		_w15112_,
		_w15116_,
		_w15118_
	);
	LUT2 #(
		.INIT('h1)
	) name11072 (
		_w15117_,
		_w15118_,
		_w15119_
	);
	LUT2 #(
		.INIT('h2)
	) name11073 (
		_w15073_,
		_w15119_,
		_w15120_
	);
	LUT2 #(
		.INIT('h4)
	) name11074 (
		_w15073_,
		_w15119_,
		_w15121_
	);
	LUT2 #(
		.INIT('h1)
	) name11075 (
		_w15120_,
		_w15121_,
		_w15122_
	);
	LUT2 #(
		.INIT('h8)
	) name11076 (
		_w15100_,
		_w15105_,
		_w15123_
	);
	LUT2 #(
		.INIT('h1)
	) name11077 (
		_w15106_,
		_w15123_,
		_w15124_
	);
	LUT2 #(
		.INIT('h4)
	) name11078 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14925_,
		_w15125_
	);
	LUT2 #(
		.INIT('h8)
	) name11079 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14929_,
		_w15126_
	);
	LUT2 #(
		.INIT('h1)
	) name11080 (
		_w15125_,
		_w15126_,
		_w15127_
	);
	LUT2 #(
		.INIT('h8)
	) name11081 (
		_w14920_,
		_w15127_,
		_w15128_
	);
	LUT2 #(
		.INIT('h1)
	) name11082 (
		_w14906_,
		_w15128_,
		_w15129_
	);
	LUT2 #(
		.INIT('h1)
	) name11083 (
		_w14990_,
		_w15129_,
		_w15130_
	);
	LUT2 #(
		.INIT('h1)
	) name11084 (
		_w14906_,
		_w14990_,
		_w15131_
	);
	LUT2 #(
		.INIT('h4)
	) name11085 (
		_w14932_,
		_w15131_,
		_w15132_
	);
	LUT2 #(
		.INIT('h2)
	) name11086 (
		_w14932_,
		_w15131_,
		_w15133_
	);
	LUT2 #(
		.INIT('h1)
	) name11087 (
		_w15132_,
		_w15133_,
		_w15134_
	);
	LUT2 #(
		.INIT('h2)
	) name11088 (
		_w15130_,
		_w15134_,
		_w15135_
	);
	LUT2 #(
		.INIT('h1)
	) name11089 (
		_w15090_,
		_w15091_,
		_w15136_
	);
	LUT2 #(
		.INIT('h2)
	) name11090 (
		_w15096_,
		_w15136_,
		_w15137_
	);
	LUT2 #(
		.INIT('h4)
	) name11091 (
		_w15096_,
		_w15136_,
		_w15138_
	);
	LUT2 #(
		.INIT('h1)
	) name11092 (
		_w15137_,
		_w15138_,
		_w15139_
	);
	LUT2 #(
		.INIT('h2)
	) name11093 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w9056_,
		_w15140_
	);
	LUT2 #(
		.INIT('h2)
	) name11094 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15140_,
		_w15141_
	);
	LUT2 #(
		.INIT('h1)
	) name11095 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15092_,
		_w15142_
	);
	LUT2 #(
		.INIT('h1)
	) name11096 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15141_,
		_w15143_
	);
	LUT2 #(
		.INIT('h4)
	) name11097 (
		_w15142_,
		_w15143_,
		_w15144_
	);
	LUT2 #(
		.INIT('h1)
	) name11098 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14947_,
		_w15145_
	);
	LUT2 #(
		.INIT('h2)
	) name11099 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14951_,
		_w15146_
	);
	LUT2 #(
		.INIT('h4)
	) name11100 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14958_,
		_w15147_
	);
	LUT2 #(
		.INIT('h8)
	) name11101 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14962_,
		_w15148_
	);
	LUT2 #(
		.INIT('h1)
	) name11102 (
		_w15147_,
		_w15148_,
		_w15149_
	);
	LUT2 #(
		.INIT('h4)
	) name11103 (
		_w15145_,
		_w15149_,
		_w15150_
	);
	LUT2 #(
		.INIT('h4)
	) name11104 (
		_w15146_,
		_w15150_,
		_w15151_
	);
	LUT2 #(
		.INIT('h2)
	) name11105 (
		_w15144_,
		_w15151_,
		_w15152_
	);
	LUT2 #(
		.INIT('h4)
	) name11106 (
		_w15144_,
		_w15151_,
		_w15153_
	);
	LUT2 #(
		.INIT('h4)
	) name11107 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14967_,
		_w15154_
	);
	LUT2 #(
		.INIT('h8)
	) name11108 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14969_,
		_w15155_
	);
	LUT2 #(
		.INIT('h1)
	) name11109 (
		_w15154_,
		_w15155_,
		_w15156_
	);
	LUT2 #(
		.INIT('h1)
	) name11110 (
		_w15153_,
		_w15156_,
		_w15157_
	);
	LUT2 #(
		.INIT('h1)
	) name11111 (
		_w15152_,
		_w15157_,
		_w15158_
	);
	LUT2 #(
		.INIT('h8)
	) name11112 (
		_w15139_,
		_w15158_,
		_w15159_
	);
	LUT2 #(
		.INIT('h1)
	) name11113 (
		_w15135_,
		_w15159_,
		_w15160_
	);
	LUT2 #(
		.INIT('h4)
	) name11114 (
		_w15079_,
		_w15098_,
		_w15161_
	);
	LUT2 #(
		.INIT('h1)
	) name11115 (
		_w15099_,
		_w15161_,
		_w15162_
	);
	LUT2 #(
		.INIT('h2)
	) name11116 (
		_w14992_,
		_w15162_,
		_w15163_
	);
	LUT2 #(
		.INIT('h4)
	) name11117 (
		_w14992_,
		_w15162_,
		_w15164_
	);
	LUT2 #(
		.INIT('h1)
	) name11118 (
		_w15163_,
		_w15164_,
		_w15165_
	);
	LUT2 #(
		.INIT('h1)
	) name11119 (
		_w15160_,
		_w15165_,
		_w15166_
	);
	LUT2 #(
		.INIT('h1)
	) name11120 (
		_w14991_,
		_w15161_,
		_w15167_
	);
	LUT2 #(
		.INIT('h8)
	) name11121 (
		_w15165_,
		_w15167_,
		_w15168_
	);
	LUT2 #(
		.INIT('h1)
	) name11122 (
		_w15166_,
		_w15168_,
		_w15169_
	);
	LUT2 #(
		.INIT('h2)
	) name11123 (
		_w15124_,
		_w15169_,
		_w15170_
	);
	LUT2 #(
		.INIT('h1)
	) name11124 (
		_w14853_,
		_w15170_,
		_w15171_
	);
	LUT2 #(
		.INIT('h4)
	) name11125 (
		_w15075_,
		_w15109_,
		_w15172_
	);
	LUT2 #(
		.INIT('h1)
	) name11126 (
		_w15110_,
		_w15172_,
		_w15173_
	);
	LUT2 #(
		.INIT('h8)
	) name11127 (
		_w14853_,
		_w15173_,
		_w15174_
	);
	LUT2 #(
		.INIT('h1)
	) name11128 (
		_w14853_,
		_w15173_,
		_w15175_
	);
	LUT2 #(
		.INIT('h1)
	) name11129 (
		_w15174_,
		_w15175_,
		_w15176_
	);
	LUT2 #(
		.INIT('h1)
	) name11130 (
		_w15171_,
		_w15176_,
		_w15177_
	);
	LUT2 #(
		.INIT('h4)
	) name11131 (
		_w15172_,
		_w15176_,
		_w15178_
	);
	LUT2 #(
		.INIT('h1)
	) name11132 (
		_w15177_,
		_w15178_,
		_w15179_
	);
	LUT2 #(
		.INIT('h8)
	) name11133 (
		_w15111_,
		_w15113_,
		_w15180_
	);
	LUT2 #(
		.INIT('h1)
	) name11134 (
		_w15117_,
		_w15180_,
		_w15181_
	);
	LUT2 #(
		.INIT('h2)
	) name11135 (
		_w15179_,
		_w15181_,
		_w15182_
	);
	LUT2 #(
		.INIT('h4)
	) name11136 (
		_w15179_,
		_w15181_,
		_w15183_
	);
	LUT2 #(
		.INIT('h8)
	) name11137 (
		_w15160_,
		_w15165_,
		_w15184_
	);
	LUT2 #(
		.INIT('h1)
	) name11138 (
		_w15166_,
		_w15184_,
		_w15185_
	);
	LUT2 #(
		.INIT('h1)
	) name11139 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14914_,
		_w15186_
	);
	LUT2 #(
		.INIT('h2)
	) name11140 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14918_,
		_w15187_
	);
	LUT2 #(
		.INIT('h4)
	) name11141 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14925_,
		_w15188_
	);
	LUT2 #(
		.INIT('h8)
	) name11142 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14929_,
		_w15189_
	);
	LUT2 #(
		.INIT('h1)
	) name11143 (
		_w15188_,
		_w15189_,
		_w15190_
	);
	LUT2 #(
		.INIT('h4)
	) name11144 (
		_w15186_,
		_w15190_,
		_w15191_
	);
	LUT2 #(
		.INIT('h4)
	) name11145 (
		_w15187_,
		_w15191_,
		_w15192_
	);
	LUT2 #(
		.INIT('h1)
	) name11146 (
		_w14906_,
		_w15192_,
		_w15193_
	);
	LUT2 #(
		.INIT('h1)
	) name11147 (
		_w14990_,
		_w15193_,
		_w15194_
	);
	LUT2 #(
		.INIT('h4)
	) name11148 (
		_w15128_,
		_w15131_,
		_w15195_
	);
	LUT2 #(
		.INIT('h2)
	) name11149 (
		_w15128_,
		_w15131_,
		_w15196_
	);
	LUT2 #(
		.INIT('h1)
	) name11150 (
		_w15195_,
		_w15196_,
		_w15197_
	);
	LUT2 #(
		.INIT('h2)
	) name11151 (
		_w15194_,
		_w15197_,
		_w15198_
	);
	LUT2 #(
		.INIT('h1)
	) name11152 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14967_,
		_w15199_
	);
	LUT2 #(
		.INIT('h2)
	) name11153 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14969_,
		_w15200_
	);
	LUT2 #(
		.INIT('h1)
	) name11154 (
		_w15199_,
		_w15200_,
		_w15201_
	);
	LUT2 #(
		.INIT('h1)
	) name11155 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14947_,
		_w15202_
	);
	LUT2 #(
		.INIT('h2)
	) name11156 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14951_,
		_w15203_
	);
	LUT2 #(
		.INIT('h4)
	) name11157 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14958_,
		_w15204_
	);
	LUT2 #(
		.INIT('h8)
	) name11158 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14962_,
		_w15205_
	);
	LUT2 #(
		.INIT('h1)
	) name11159 (
		_w15204_,
		_w15205_,
		_w15206_
	);
	LUT2 #(
		.INIT('h4)
	) name11160 (
		_w15202_,
		_w15206_,
		_w15207_
	);
	LUT2 #(
		.INIT('h4)
	) name11161 (
		_w15203_,
		_w15207_,
		_w15208_
	);
	LUT2 #(
		.INIT('h2)
	) name11162 (
		_w15201_,
		_w15208_,
		_w15209_
	);
	LUT2 #(
		.INIT('h4)
	) name11163 (
		_w15201_,
		_w15208_,
		_w15210_
	);
	LUT2 #(
		.INIT('h2)
	) name11164 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w8358_,
		_w15211_
	);
	LUT2 #(
		.INIT('h2)
	) name11165 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15211_,
		_w15212_
	);
	LUT2 #(
		.INIT('h1)
	) name11166 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15140_,
		_w15213_
	);
	LUT2 #(
		.INIT('h1)
	) name11167 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15212_,
		_w15214_
	);
	LUT2 #(
		.INIT('h4)
	) name11168 (
		_w15213_,
		_w15214_,
		_w15215_
	);
	LUT2 #(
		.INIT('h4)
	) name11169 (
		_w15210_,
		_w15215_,
		_w15216_
	);
	LUT2 #(
		.INIT('h1)
	) name11170 (
		_w15209_,
		_w15216_,
		_w15217_
	);
	LUT2 #(
		.INIT('h1)
	) name11171 (
		_w15152_,
		_w15153_,
		_w15218_
	);
	LUT2 #(
		.INIT('h4)
	) name11172 (
		_w15156_,
		_w15218_,
		_w15219_
	);
	LUT2 #(
		.INIT('h2)
	) name11173 (
		_w15156_,
		_w15218_,
		_w15220_
	);
	LUT2 #(
		.INIT('h1)
	) name11174 (
		_w15219_,
		_w15220_,
		_w15221_
	);
	LUT2 #(
		.INIT('h2)
	) name11175 (
		_w15217_,
		_w15221_,
		_w15222_
	);
	LUT2 #(
		.INIT('h1)
	) name11176 (
		_w15198_,
		_w15222_,
		_w15223_
	);
	LUT2 #(
		.INIT('h4)
	) name11177 (
		_w15130_,
		_w15134_,
		_w15224_
	);
	LUT2 #(
		.INIT('h1)
	) name11178 (
		_w15135_,
		_w15224_,
		_w15225_
	);
	LUT2 #(
		.INIT('h1)
	) name11179 (
		_w15139_,
		_w15158_,
		_w15226_
	);
	LUT2 #(
		.INIT('h1)
	) name11180 (
		_w15159_,
		_w15226_,
		_w15227_
	);
	LUT2 #(
		.INIT('h8)
	) name11181 (
		_w15225_,
		_w15227_,
		_w15228_
	);
	LUT2 #(
		.INIT('h1)
	) name11182 (
		_w15225_,
		_w15227_,
		_w15229_
	);
	LUT2 #(
		.INIT('h1)
	) name11183 (
		_w15228_,
		_w15229_,
		_w15230_
	);
	LUT2 #(
		.INIT('h4)
	) name11184 (
		_w15223_,
		_w15230_,
		_w15231_
	);
	LUT2 #(
		.INIT('h1)
	) name11185 (
		_w15224_,
		_w15226_,
		_w15232_
	);
	LUT2 #(
		.INIT('h4)
	) name11186 (
		_w15230_,
		_w15232_,
		_w15233_
	);
	LUT2 #(
		.INIT('h1)
	) name11187 (
		_w15231_,
		_w15233_,
		_w15234_
	);
	LUT2 #(
		.INIT('h2)
	) name11188 (
		_w15185_,
		_w15234_,
		_w15235_
	);
	LUT2 #(
		.INIT('h1)
	) name11189 (
		_w14853_,
		_w15235_,
		_w15236_
	);
	LUT2 #(
		.INIT('h4)
	) name11190 (
		_w15124_,
		_w15169_,
		_w15237_
	);
	LUT2 #(
		.INIT('h1)
	) name11191 (
		_w15170_,
		_w15237_,
		_w15238_
	);
	LUT2 #(
		.INIT('h8)
	) name11192 (
		_w14853_,
		_w15238_,
		_w15239_
	);
	LUT2 #(
		.INIT('h1)
	) name11193 (
		_w14853_,
		_w15238_,
		_w15240_
	);
	LUT2 #(
		.INIT('h1)
	) name11194 (
		_w15239_,
		_w15240_,
		_w15241_
	);
	LUT2 #(
		.INIT('h1)
	) name11195 (
		_w15236_,
		_w15241_,
		_w15242_
	);
	LUT2 #(
		.INIT('h8)
	) name11196 (
		_w15236_,
		_w15238_,
		_w15243_
	);
	LUT2 #(
		.INIT('h1)
	) name11197 (
		_w15242_,
		_w15243_,
		_w15244_
	);
	LUT2 #(
		.INIT('h8)
	) name11198 (
		_w15171_,
		_w15173_,
		_w15245_
	);
	LUT2 #(
		.INIT('h1)
	) name11199 (
		_w15177_,
		_w15245_,
		_w15246_
	);
	LUT2 #(
		.INIT('h1)
	) name11200 (
		_w15244_,
		_w15246_,
		_w15247_
	);
	LUT2 #(
		.INIT('h2)
	) name11201 (
		_w15223_,
		_w15230_,
		_w15248_
	);
	LUT2 #(
		.INIT('h1)
	) name11202 (
		_w15231_,
		_w15248_,
		_w15249_
	);
	LUT2 #(
		.INIT('h1)
	) name11203 (
		_w15209_,
		_w15210_,
		_w15250_
	);
	LUT2 #(
		.INIT('h8)
	) name11204 (
		_w15215_,
		_w15250_,
		_w15251_
	);
	LUT2 #(
		.INIT('h1)
	) name11205 (
		_w15215_,
		_w15250_,
		_w15252_
	);
	LUT2 #(
		.INIT('h1)
	) name11206 (
		_w15251_,
		_w15252_,
		_w15253_
	);
	LUT2 #(
		.INIT('h2)
	) name11207 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w7737_,
		_w15254_
	);
	LUT2 #(
		.INIT('h2)
	) name11208 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15254_,
		_w15255_
	);
	LUT2 #(
		.INIT('h1)
	) name11209 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15211_,
		_w15256_
	);
	LUT2 #(
		.INIT('h1)
	) name11210 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15255_,
		_w15257_
	);
	LUT2 #(
		.INIT('h4)
	) name11211 (
		_w15256_,
		_w15257_,
		_w15258_
	);
	LUT2 #(
		.INIT('h1)
	) name11212 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14947_,
		_w15259_
	);
	LUT2 #(
		.INIT('h2)
	) name11213 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14951_,
		_w15260_
	);
	LUT2 #(
		.INIT('h4)
	) name11214 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14958_,
		_w15261_
	);
	LUT2 #(
		.INIT('h8)
	) name11215 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14962_,
		_w15262_
	);
	LUT2 #(
		.INIT('h1)
	) name11216 (
		_w15261_,
		_w15262_,
		_w15263_
	);
	LUT2 #(
		.INIT('h4)
	) name11217 (
		_w15259_,
		_w15263_,
		_w15264_
	);
	LUT2 #(
		.INIT('h4)
	) name11218 (
		_w15260_,
		_w15264_,
		_w15265_
	);
	LUT2 #(
		.INIT('h2)
	) name11219 (
		_w15258_,
		_w15265_,
		_w15266_
	);
	LUT2 #(
		.INIT('h4)
	) name11220 (
		_w15258_,
		_w15265_,
		_w15267_
	);
	LUT2 #(
		.INIT('h4)
	) name11221 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14967_,
		_w15268_
	);
	LUT2 #(
		.INIT('h8)
	) name11222 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14969_,
		_w15269_
	);
	LUT2 #(
		.INIT('h1)
	) name11223 (
		_w15268_,
		_w15269_,
		_w15270_
	);
	LUT2 #(
		.INIT('h1)
	) name11224 (
		_w15267_,
		_w15270_,
		_w15271_
	);
	LUT2 #(
		.INIT('h1)
	) name11225 (
		_w15266_,
		_w15271_,
		_w15272_
	);
	LUT2 #(
		.INIT('h4)
	) name11226 (
		_w15253_,
		_w15272_,
		_w15273_
	);
	LUT2 #(
		.INIT('h1)
	) name11227 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14914_,
		_w15274_
	);
	LUT2 #(
		.INIT('h2)
	) name11228 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14918_,
		_w15275_
	);
	LUT2 #(
		.INIT('h4)
	) name11229 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14925_,
		_w15276_
	);
	LUT2 #(
		.INIT('h8)
	) name11230 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14929_,
		_w15277_
	);
	LUT2 #(
		.INIT('h1)
	) name11231 (
		_w15276_,
		_w15277_,
		_w15278_
	);
	LUT2 #(
		.INIT('h4)
	) name11232 (
		_w15274_,
		_w15278_,
		_w15279_
	);
	LUT2 #(
		.INIT('h4)
	) name11233 (
		_w15275_,
		_w15279_,
		_w15280_
	);
	LUT2 #(
		.INIT('h8)
	) name11234 (
		_w14879_,
		_w15280_,
		_w15281_
	);
	LUT2 #(
		.INIT('h4)
	) name11235 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14898_,
		_w15282_
	);
	LUT2 #(
		.INIT('h8)
	) name11236 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14902_,
		_w15283_
	);
	LUT2 #(
		.INIT('h1)
	) name11237 (
		_w15282_,
		_w15283_,
		_w15284_
	);
	LUT2 #(
		.INIT('h8)
	) name11238 (
		_w14893_,
		_w15284_,
		_w15285_
	);
	LUT2 #(
		.INIT('h1)
	) name11239 (
		_w15281_,
		_w15285_,
		_w15286_
	);
	LUT2 #(
		.INIT('h1)
	) name11240 (
		_w14879_,
		_w15280_,
		_w15287_
	);
	LUT2 #(
		.INIT('h1)
	) name11241 (
		_w15286_,
		_w15287_,
		_w15288_
	);
	LUT2 #(
		.INIT('h2)
	) name11242 (
		_w15131_,
		_w15192_,
		_w15289_
	);
	LUT2 #(
		.INIT('h4)
	) name11243 (
		_w15131_,
		_w15192_,
		_w15290_
	);
	LUT2 #(
		.INIT('h1)
	) name11244 (
		_w15289_,
		_w15290_,
		_w15291_
	);
	LUT2 #(
		.INIT('h2)
	) name11245 (
		_w15288_,
		_w15291_,
		_w15292_
	);
	LUT2 #(
		.INIT('h1)
	) name11246 (
		_w15273_,
		_w15292_,
		_w15293_
	);
	LUT2 #(
		.INIT('h4)
	) name11247 (
		_w15194_,
		_w15197_,
		_w15294_
	);
	LUT2 #(
		.INIT('h1)
	) name11248 (
		_w15198_,
		_w15294_,
		_w15295_
	);
	LUT2 #(
		.INIT('h4)
	) name11249 (
		_w15217_,
		_w15221_,
		_w15296_
	);
	LUT2 #(
		.INIT('h1)
	) name11250 (
		_w15222_,
		_w15296_,
		_w15297_
	);
	LUT2 #(
		.INIT('h8)
	) name11251 (
		_w15295_,
		_w15297_,
		_w15298_
	);
	LUT2 #(
		.INIT('h1)
	) name11252 (
		_w15295_,
		_w15297_,
		_w15299_
	);
	LUT2 #(
		.INIT('h1)
	) name11253 (
		_w15298_,
		_w15299_,
		_w15300_
	);
	LUT2 #(
		.INIT('h4)
	) name11254 (
		_w15293_,
		_w15300_,
		_w15301_
	);
	LUT2 #(
		.INIT('h1)
	) name11255 (
		_w15294_,
		_w15296_,
		_w15302_
	);
	LUT2 #(
		.INIT('h4)
	) name11256 (
		_w15300_,
		_w15302_,
		_w15303_
	);
	LUT2 #(
		.INIT('h1)
	) name11257 (
		_w15301_,
		_w15303_,
		_w15304_
	);
	LUT2 #(
		.INIT('h2)
	) name11258 (
		_w15249_,
		_w15304_,
		_w15305_
	);
	LUT2 #(
		.INIT('h1)
	) name11259 (
		_w14853_,
		_w15305_,
		_w15306_
	);
	LUT2 #(
		.INIT('h4)
	) name11260 (
		_w15185_,
		_w15234_,
		_w15307_
	);
	LUT2 #(
		.INIT('h1)
	) name11261 (
		_w15235_,
		_w15307_,
		_w15308_
	);
	LUT2 #(
		.INIT('h8)
	) name11262 (
		_w14853_,
		_w15308_,
		_w15309_
	);
	LUT2 #(
		.INIT('h1)
	) name11263 (
		_w14853_,
		_w15308_,
		_w15310_
	);
	LUT2 #(
		.INIT('h1)
	) name11264 (
		_w15309_,
		_w15310_,
		_w15311_
	);
	LUT2 #(
		.INIT('h1)
	) name11265 (
		_w15306_,
		_w15311_,
		_w15312_
	);
	LUT2 #(
		.INIT('h4)
	) name11266 (
		_w15307_,
		_w15311_,
		_w15313_
	);
	LUT2 #(
		.INIT('h1)
	) name11267 (
		_w15312_,
		_w15313_,
		_w15314_
	);
	LUT2 #(
		.INIT('h4)
	) name11268 (
		_w15237_,
		_w15241_,
		_w15315_
	);
	LUT2 #(
		.INIT('h1)
	) name11269 (
		_w15242_,
		_w15315_,
		_w15316_
	);
	LUT2 #(
		.INIT('h2)
	) name11270 (
		_w15246_,
		_w15316_,
		_w15317_
	);
	LUT2 #(
		.INIT('h2)
	) name11271 (
		_w15314_,
		_w15317_,
		_w15318_
	);
	LUT2 #(
		.INIT('h1)
	) name11272 (
		_w15247_,
		_w15318_,
		_w15319_
	);
	LUT2 #(
		.INIT('h4)
	) name11273 (
		_w8354_,
		_w14993_,
		_w15320_
	);
	LUT2 #(
		.INIT('h2)
	) name11274 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w7753_,
		_w15321_
	);
	LUT2 #(
		.INIT('h8)
	) name11275 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15321_,
		_w15322_
	);
	LUT2 #(
		.INIT('h1)
	) name11276 (
		_w15320_,
		_w15322_,
		_w15323_
	);
	LUT2 #(
		.INIT('h1)
	) name11277 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15323_,
		_w15324_
	);
	LUT2 #(
		.INIT('h1)
	) name11278 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14838_,
		_w15325_
	);
	LUT2 #(
		.INIT('h2)
	) name11279 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14842_,
		_w15326_
	);
	LUT2 #(
		.INIT('h4)
	) name11280 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14846_,
		_w15327_
	);
	LUT2 #(
		.INIT('h8)
	) name11281 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14849_,
		_w15328_
	);
	LUT2 #(
		.INIT('h1)
	) name11282 (
		_w15327_,
		_w15328_,
		_w15329_
	);
	LUT2 #(
		.INIT('h4)
	) name11283 (
		_w15325_,
		_w15329_,
		_w15330_
	);
	LUT2 #(
		.INIT('h4)
	) name11284 (
		_w15326_,
		_w15330_,
		_w15331_
	);
	LUT2 #(
		.INIT('h4)
	) name11285 (
		_w15324_,
		_w15331_,
		_w15332_
	);
	LUT2 #(
		.INIT('h2)
	) name11286 (
		_w15324_,
		_w15331_,
		_w15333_
	);
	LUT2 #(
		.INIT('h2)
	) name11287 (
		_w14887_,
		_w15333_,
		_w15334_
	);
	LUT2 #(
		.INIT('h1)
	) name11288 (
		_w15332_,
		_w15334_,
		_w15335_
	);
	LUT2 #(
		.INIT('h4)
	) name11289 (
		_w9072_,
		_w14993_,
		_w15336_
	);
	LUT2 #(
		.INIT('h4)
	) name11290 (
		_w8354_,
		_w15044_,
		_w15337_
	);
	LUT2 #(
		.INIT('h1)
	) name11291 (
		_w15336_,
		_w15337_,
		_w15338_
	);
	LUT2 #(
		.INIT('h1)
	) name11292 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15338_,
		_w15339_
	);
	LUT2 #(
		.INIT('h1)
	) name11293 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14838_,
		_w15340_
	);
	LUT2 #(
		.INIT('h2)
	) name11294 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14842_,
		_w15341_
	);
	LUT2 #(
		.INIT('h4)
	) name11295 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14846_,
		_w15342_
	);
	LUT2 #(
		.INIT('h8)
	) name11296 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14849_,
		_w15343_
	);
	LUT2 #(
		.INIT('h1)
	) name11297 (
		_w15342_,
		_w15343_,
		_w15344_
	);
	LUT2 #(
		.INIT('h4)
	) name11298 (
		_w15340_,
		_w15344_,
		_w15345_
	);
	LUT2 #(
		.INIT('h4)
	) name11299 (
		_w15341_,
		_w15345_,
		_w15346_
	);
	LUT2 #(
		.INIT('h2)
	) name11300 (
		_w15339_,
		_w15346_,
		_w15347_
	);
	LUT2 #(
		.INIT('h4)
	) name11301 (
		_w15339_,
		_w15346_,
		_w15348_
	);
	LUT2 #(
		.INIT('h1)
	) name11302 (
		_w15347_,
		_w15348_,
		_w15349_
	);
	LUT2 #(
		.INIT('h8)
	) name11303 (
		_w14898_,
		_w15349_,
		_w15350_
	);
	LUT2 #(
		.INIT('h1)
	) name11304 (
		_w14898_,
		_w15349_,
		_w15351_
	);
	LUT2 #(
		.INIT('h1)
	) name11305 (
		_w15350_,
		_w15351_,
		_w15352_
	);
	LUT2 #(
		.INIT('h1)
	) name11306 (
		_w15335_,
		_w15352_,
		_w15353_
	);
	LUT2 #(
		.INIT('h1)
	) name11307 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14787_,
		_w15354_
	);
	LUT2 #(
		.INIT('h2)
	) name11308 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14791_,
		_w15355_
	);
	LUT2 #(
		.INIT('h4)
	) name11309 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14798_,
		_w15356_
	);
	LUT2 #(
		.INIT('h8)
	) name11310 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14802_,
		_w15357_
	);
	LUT2 #(
		.INIT('h1)
	) name11311 (
		_w15356_,
		_w15357_,
		_w15358_
	);
	LUT2 #(
		.INIT('h4)
	) name11312 (
		_w15354_,
		_w15358_,
		_w15359_
	);
	LUT2 #(
		.INIT('h4)
	) name11313 (
		_w15355_,
		_w15359_,
		_w15360_
	);
	LUT2 #(
		.INIT('h1)
	) name11314 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14761_,
		_w15361_
	);
	LUT2 #(
		.INIT('h2)
	) name11315 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14765_,
		_w15362_
	);
	LUT2 #(
		.INIT('h4)
	) name11316 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14772_,
		_w15363_
	);
	LUT2 #(
		.INIT('h8)
	) name11317 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14776_,
		_w15364_
	);
	LUT2 #(
		.INIT('h1)
	) name11318 (
		_w15363_,
		_w15364_,
		_w15365_
	);
	LUT2 #(
		.INIT('h4)
	) name11319 (
		_w15361_,
		_w15365_,
		_w15366_
	);
	LUT2 #(
		.INIT('h4)
	) name11320 (
		_w15362_,
		_w15366_,
		_w15367_
	);
	LUT2 #(
		.INIT('h1)
	) name11321 (
		_w15360_,
		_w15367_,
		_w15368_
	);
	LUT2 #(
		.INIT('h8)
	) name11322 (
		_w15360_,
		_w15367_,
		_w15369_
	);
	LUT2 #(
		.INIT('h1)
	) name11323 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14814_,
		_w15370_
	);
	LUT2 #(
		.INIT('h2)
	) name11324 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14818_,
		_w15371_
	);
	LUT2 #(
		.INIT('h4)
	) name11325 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14825_,
		_w15372_
	);
	LUT2 #(
		.INIT('h8)
	) name11326 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14829_,
		_w15373_
	);
	LUT2 #(
		.INIT('h1)
	) name11327 (
		_w15372_,
		_w15373_,
		_w15374_
	);
	LUT2 #(
		.INIT('h4)
	) name11328 (
		_w15370_,
		_w15374_,
		_w15375_
	);
	LUT2 #(
		.INIT('h4)
	) name11329 (
		_w15371_,
		_w15375_,
		_w15376_
	);
	LUT2 #(
		.INIT('h1)
	) name11330 (
		_w15369_,
		_w15376_,
		_w15377_
	);
	LUT2 #(
		.INIT('h1)
	) name11331 (
		_w15368_,
		_w15377_,
		_w15378_
	);
	LUT2 #(
		.INIT('h1)
	) name11332 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14787_,
		_w15379_
	);
	LUT2 #(
		.INIT('h2)
	) name11333 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14791_,
		_w15380_
	);
	LUT2 #(
		.INIT('h4)
	) name11334 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14798_,
		_w15381_
	);
	LUT2 #(
		.INIT('h8)
	) name11335 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14802_,
		_w15382_
	);
	LUT2 #(
		.INIT('h1)
	) name11336 (
		_w15381_,
		_w15382_,
		_w15383_
	);
	LUT2 #(
		.INIT('h4)
	) name11337 (
		_w15379_,
		_w15383_,
		_w15384_
	);
	LUT2 #(
		.INIT('h4)
	) name11338 (
		_w15380_,
		_w15384_,
		_w15385_
	);
	LUT2 #(
		.INIT('h1)
	) name11339 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14761_,
		_w15386_
	);
	LUT2 #(
		.INIT('h2)
	) name11340 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14765_,
		_w15387_
	);
	LUT2 #(
		.INIT('h4)
	) name11341 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14772_,
		_w15388_
	);
	LUT2 #(
		.INIT('h8)
	) name11342 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14776_,
		_w15389_
	);
	LUT2 #(
		.INIT('h1)
	) name11343 (
		_w15388_,
		_w15389_,
		_w15390_
	);
	LUT2 #(
		.INIT('h4)
	) name11344 (
		_w15386_,
		_w15390_,
		_w15391_
	);
	LUT2 #(
		.INIT('h4)
	) name11345 (
		_w15387_,
		_w15391_,
		_w15392_
	);
	LUT2 #(
		.INIT('h8)
	) name11346 (
		_w15385_,
		_w15392_,
		_w15393_
	);
	LUT2 #(
		.INIT('h1)
	) name11347 (
		_w15385_,
		_w15392_,
		_w15394_
	);
	LUT2 #(
		.INIT('h1)
	) name11348 (
		_w15393_,
		_w15394_,
		_w15395_
	);
	LUT2 #(
		.INIT('h1)
	) name11349 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14814_,
		_w15396_
	);
	LUT2 #(
		.INIT('h2)
	) name11350 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14818_,
		_w15397_
	);
	LUT2 #(
		.INIT('h4)
	) name11351 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14825_,
		_w15398_
	);
	LUT2 #(
		.INIT('h8)
	) name11352 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14829_,
		_w15399_
	);
	LUT2 #(
		.INIT('h1)
	) name11353 (
		_w15398_,
		_w15399_,
		_w15400_
	);
	LUT2 #(
		.INIT('h4)
	) name11354 (
		_w15396_,
		_w15400_,
		_w15401_
	);
	LUT2 #(
		.INIT('h4)
	) name11355 (
		_w15397_,
		_w15401_,
		_w15402_
	);
	LUT2 #(
		.INIT('h4)
	) name11356 (
		_w15395_,
		_w15402_,
		_w15403_
	);
	LUT2 #(
		.INIT('h2)
	) name11357 (
		_w15395_,
		_w15402_,
		_w15404_
	);
	LUT2 #(
		.INIT('h1)
	) name11358 (
		_w15403_,
		_w15404_,
		_w15405_
	);
	LUT2 #(
		.INIT('h2)
	) name11359 (
		_w15378_,
		_w15405_,
		_w15406_
	);
	LUT2 #(
		.INIT('h1)
	) name11360 (
		_w15353_,
		_w15406_,
		_w15407_
	);
	LUT2 #(
		.INIT('h1)
	) name11361 (
		_w15393_,
		_w15402_,
		_w15408_
	);
	LUT2 #(
		.INIT('h1)
	) name11362 (
		_w15394_,
		_w15408_,
		_w15409_
	);
	LUT2 #(
		.INIT('h1)
	) name11363 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14761_,
		_w15410_
	);
	LUT2 #(
		.INIT('h2)
	) name11364 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14765_,
		_w15411_
	);
	LUT2 #(
		.INIT('h4)
	) name11365 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14772_,
		_w15412_
	);
	LUT2 #(
		.INIT('h8)
	) name11366 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14776_,
		_w15413_
	);
	LUT2 #(
		.INIT('h1)
	) name11367 (
		_w15412_,
		_w15413_,
		_w15414_
	);
	LUT2 #(
		.INIT('h4)
	) name11368 (
		_w15410_,
		_w15414_,
		_w15415_
	);
	LUT2 #(
		.INIT('h4)
	) name11369 (
		_w15411_,
		_w15415_,
		_w15416_
	);
	LUT2 #(
		.INIT('h1)
	) name11370 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14787_,
		_w15417_
	);
	LUT2 #(
		.INIT('h2)
	) name11371 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14791_,
		_w15418_
	);
	LUT2 #(
		.INIT('h4)
	) name11372 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14798_,
		_w15419_
	);
	LUT2 #(
		.INIT('h8)
	) name11373 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14802_,
		_w15420_
	);
	LUT2 #(
		.INIT('h1)
	) name11374 (
		_w15419_,
		_w15420_,
		_w15421_
	);
	LUT2 #(
		.INIT('h4)
	) name11375 (
		_w15417_,
		_w15421_,
		_w15422_
	);
	LUT2 #(
		.INIT('h4)
	) name11376 (
		_w15418_,
		_w15422_,
		_w15423_
	);
	LUT2 #(
		.INIT('h8)
	) name11377 (
		_w15416_,
		_w15423_,
		_w15424_
	);
	LUT2 #(
		.INIT('h1)
	) name11378 (
		_w15416_,
		_w15423_,
		_w15425_
	);
	LUT2 #(
		.INIT('h1)
	) name11379 (
		_w15424_,
		_w15425_,
		_w15426_
	);
	LUT2 #(
		.INIT('h1)
	) name11380 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14814_,
		_w15427_
	);
	LUT2 #(
		.INIT('h2)
	) name11381 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14818_,
		_w15428_
	);
	LUT2 #(
		.INIT('h4)
	) name11382 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14825_,
		_w15429_
	);
	LUT2 #(
		.INIT('h8)
	) name11383 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14829_,
		_w15430_
	);
	LUT2 #(
		.INIT('h1)
	) name11384 (
		_w15429_,
		_w15430_,
		_w15431_
	);
	LUT2 #(
		.INIT('h4)
	) name11385 (
		_w15427_,
		_w15431_,
		_w15432_
	);
	LUT2 #(
		.INIT('h4)
	) name11386 (
		_w15428_,
		_w15432_,
		_w15433_
	);
	LUT2 #(
		.INIT('h4)
	) name11387 (
		_w15426_,
		_w15433_,
		_w15434_
	);
	LUT2 #(
		.INIT('h2)
	) name11388 (
		_w15426_,
		_w15433_,
		_w15435_
	);
	LUT2 #(
		.INIT('h1)
	) name11389 (
		_w15434_,
		_w15435_,
		_w15436_
	);
	LUT2 #(
		.INIT('h2)
	) name11390 (
		_w15409_,
		_w15436_,
		_w15437_
	);
	LUT2 #(
		.INIT('h4)
	) name11391 (
		_w15409_,
		_w15436_,
		_w15438_
	);
	LUT2 #(
		.INIT('h1)
	) name11392 (
		_w15437_,
		_w15438_,
		_w15439_
	);
	LUT2 #(
		.INIT('h1)
	) name11393 (
		_w14898_,
		_w15347_,
		_w15440_
	);
	LUT2 #(
		.INIT('h1)
	) name11394 (
		_w15348_,
		_w15440_,
		_w15441_
	);
	LUT2 #(
		.INIT('h4)
	) name11395 (
		_w7182_,
		_w14993_,
		_w15442_
	);
	LUT2 #(
		.INIT('h4)
	) name11396 (
		_w9072_,
		_w15044_,
		_w15443_
	);
	LUT2 #(
		.INIT('h1)
	) name11397 (
		_w15442_,
		_w15443_,
		_w15444_
	);
	LUT2 #(
		.INIT('h1)
	) name11398 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15444_,
		_w15445_
	);
	LUT2 #(
		.INIT('h1)
	) name11399 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14838_,
		_w15446_
	);
	LUT2 #(
		.INIT('h2)
	) name11400 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14842_,
		_w15447_
	);
	LUT2 #(
		.INIT('h4)
	) name11401 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14846_,
		_w15448_
	);
	LUT2 #(
		.INIT('h8)
	) name11402 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14849_,
		_w15449_
	);
	LUT2 #(
		.INIT('h1)
	) name11403 (
		_w15448_,
		_w15449_,
		_w15450_
	);
	LUT2 #(
		.INIT('h4)
	) name11404 (
		_w15446_,
		_w15450_,
		_w15451_
	);
	LUT2 #(
		.INIT('h4)
	) name11405 (
		_w15447_,
		_w15451_,
		_w15452_
	);
	LUT2 #(
		.INIT('h2)
	) name11406 (
		_w15445_,
		_w15452_,
		_w15453_
	);
	LUT2 #(
		.INIT('h4)
	) name11407 (
		_w15445_,
		_w15452_,
		_w15454_
	);
	LUT2 #(
		.INIT('h1)
	) name11408 (
		_w15453_,
		_w15454_,
		_w15455_
	);
	LUT2 #(
		.INIT('h2)
	) name11409 (
		_w14914_,
		_w15455_,
		_w15456_
	);
	LUT2 #(
		.INIT('h4)
	) name11410 (
		_w14914_,
		_w15455_,
		_w15457_
	);
	LUT2 #(
		.INIT('h1)
	) name11411 (
		_w15456_,
		_w15457_,
		_w15458_
	);
	LUT2 #(
		.INIT('h1)
	) name11412 (
		_w15441_,
		_w15458_,
		_w15459_
	);
	LUT2 #(
		.INIT('h8)
	) name11413 (
		_w15441_,
		_w15458_,
		_w15460_
	);
	LUT2 #(
		.INIT('h1)
	) name11414 (
		_w15459_,
		_w15460_,
		_w15461_
	);
	LUT2 #(
		.INIT('h8)
	) name11415 (
		_w15439_,
		_w15461_,
		_w15462_
	);
	LUT2 #(
		.INIT('h1)
	) name11416 (
		_w15439_,
		_w15461_,
		_w15463_
	);
	LUT2 #(
		.INIT('h1)
	) name11417 (
		_w15462_,
		_w15463_,
		_w15464_
	);
	LUT2 #(
		.INIT('h4)
	) name11418 (
		_w15407_,
		_w15464_,
		_w15465_
	);
	LUT2 #(
		.INIT('h2)
	) name11419 (
		_w15407_,
		_w15464_,
		_w15466_
	);
	LUT2 #(
		.INIT('h1)
	) name11420 (
		_w15465_,
		_w15466_,
		_w15467_
	);
	LUT2 #(
		.INIT('h1)
	) name11421 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14787_,
		_w15468_
	);
	LUT2 #(
		.INIT('h2)
	) name11422 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14791_,
		_w15469_
	);
	LUT2 #(
		.INIT('h4)
	) name11423 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14798_,
		_w15470_
	);
	LUT2 #(
		.INIT('h8)
	) name11424 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14802_,
		_w15471_
	);
	LUT2 #(
		.INIT('h1)
	) name11425 (
		_w15470_,
		_w15471_,
		_w15472_
	);
	LUT2 #(
		.INIT('h4)
	) name11426 (
		_w15468_,
		_w15472_,
		_w15473_
	);
	LUT2 #(
		.INIT('h4)
	) name11427 (
		_w15469_,
		_w15473_,
		_w15474_
	);
	LUT2 #(
		.INIT('h1)
	) name11428 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14761_,
		_w15475_
	);
	LUT2 #(
		.INIT('h2)
	) name11429 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14765_,
		_w15476_
	);
	LUT2 #(
		.INIT('h4)
	) name11430 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14772_,
		_w15477_
	);
	LUT2 #(
		.INIT('h8)
	) name11431 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14776_,
		_w15478_
	);
	LUT2 #(
		.INIT('h1)
	) name11432 (
		_w15477_,
		_w15478_,
		_w15479_
	);
	LUT2 #(
		.INIT('h4)
	) name11433 (
		_w15475_,
		_w15479_,
		_w15480_
	);
	LUT2 #(
		.INIT('h4)
	) name11434 (
		_w15476_,
		_w15480_,
		_w15481_
	);
	LUT2 #(
		.INIT('h1)
	) name11435 (
		_w15474_,
		_w15481_,
		_w15482_
	);
	LUT2 #(
		.INIT('h8)
	) name11436 (
		_w15474_,
		_w15481_,
		_w15483_
	);
	LUT2 #(
		.INIT('h1)
	) name11437 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14814_,
		_w15484_
	);
	LUT2 #(
		.INIT('h2)
	) name11438 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14818_,
		_w15485_
	);
	LUT2 #(
		.INIT('h4)
	) name11439 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14825_,
		_w15486_
	);
	LUT2 #(
		.INIT('h8)
	) name11440 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14829_,
		_w15487_
	);
	LUT2 #(
		.INIT('h1)
	) name11441 (
		_w15486_,
		_w15487_,
		_w15488_
	);
	LUT2 #(
		.INIT('h4)
	) name11442 (
		_w15484_,
		_w15488_,
		_w15489_
	);
	LUT2 #(
		.INIT('h4)
	) name11443 (
		_w15485_,
		_w15489_,
		_w15490_
	);
	LUT2 #(
		.INIT('h1)
	) name11444 (
		_w15483_,
		_w15490_,
		_w15491_
	);
	LUT2 #(
		.INIT('h1)
	) name11445 (
		_w15482_,
		_w15491_,
		_w15492_
	);
	LUT2 #(
		.INIT('h1)
	) name11446 (
		_w15368_,
		_w15369_,
		_w15493_
	);
	LUT2 #(
		.INIT('h2)
	) name11447 (
		_w15376_,
		_w15493_,
		_w15494_
	);
	LUT2 #(
		.INIT('h4)
	) name11448 (
		_w15376_,
		_w15493_,
		_w15495_
	);
	LUT2 #(
		.INIT('h1)
	) name11449 (
		_w15494_,
		_w15495_,
		_w15496_
	);
	LUT2 #(
		.INIT('h2)
	) name11450 (
		_w15492_,
		_w15496_,
		_w15497_
	);
	LUT2 #(
		.INIT('h4)
	) name11451 (
		_w10112_,
		_w15044_,
		_w15498_
	);
	LUT2 #(
		.INIT('h4)
	) name11452 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15321_,
		_w15499_
	);
	LUT2 #(
		.INIT('h1)
	) name11453 (
		_w15498_,
		_w15499_,
		_w15500_
	);
	LUT2 #(
		.INIT('h1)
	) name11454 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15500_,
		_w15501_
	);
	LUT2 #(
		.INIT('h1)
	) name11455 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14838_,
		_w15502_
	);
	LUT2 #(
		.INIT('h2)
	) name11456 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14842_,
		_w15503_
	);
	LUT2 #(
		.INIT('h4)
	) name11457 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14846_,
		_w15504_
	);
	LUT2 #(
		.INIT('h8)
	) name11458 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14849_,
		_w15505_
	);
	LUT2 #(
		.INIT('h1)
	) name11459 (
		_w15504_,
		_w15505_,
		_w15506_
	);
	LUT2 #(
		.INIT('h4)
	) name11460 (
		_w15502_,
		_w15506_,
		_w15507_
	);
	LUT2 #(
		.INIT('h4)
	) name11461 (
		_w15503_,
		_w15507_,
		_w15508_
	);
	LUT2 #(
		.INIT('h4)
	) name11462 (
		_w15501_,
		_w15508_,
		_w15509_
	);
	LUT2 #(
		.INIT('h2)
	) name11463 (
		_w15501_,
		_w15508_,
		_w15510_
	);
	LUT2 #(
		.INIT('h1)
	) name11464 (
		_w14872_,
		_w15510_,
		_w15511_
	);
	LUT2 #(
		.INIT('h1)
	) name11465 (
		_w15509_,
		_w15511_,
		_w15512_
	);
	LUT2 #(
		.INIT('h1)
	) name11466 (
		_w15332_,
		_w15333_,
		_w15513_
	);
	LUT2 #(
		.INIT('h2)
	) name11467 (
		_w14887_,
		_w15513_,
		_w15514_
	);
	LUT2 #(
		.INIT('h4)
	) name11468 (
		_w14887_,
		_w15513_,
		_w15515_
	);
	LUT2 #(
		.INIT('h1)
	) name11469 (
		_w15514_,
		_w15515_,
		_w15516_
	);
	LUT2 #(
		.INIT('h1)
	) name11470 (
		_w15512_,
		_w15516_,
		_w15517_
	);
	LUT2 #(
		.INIT('h1)
	) name11471 (
		_w15497_,
		_w15517_,
		_w15518_
	);
	LUT2 #(
		.INIT('h4)
	) name11472 (
		_w15378_,
		_w15405_,
		_w15519_
	);
	LUT2 #(
		.INIT('h1)
	) name11473 (
		_w15406_,
		_w15519_,
		_w15520_
	);
	LUT2 #(
		.INIT('h8)
	) name11474 (
		_w15335_,
		_w15352_,
		_w15521_
	);
	LUT2 #(
		.INIT('h1)
	) name11475 (
		_w15353_,
		_w15521_,
		_w15522_
	);
	LUT2 #(
		.INIT('h8)
	) name11476 (
		_w15520_,
		_w15522_,
		_w15523_
	);
	LUT2 #(
		.INIT('h1)
	) name11477 (
		_w15520_,
		_w15522_,
		_w15524_
	);
	LUT2 #(
		.INIT('h1)
	) name11478 (
		_w15523_,
		_w15524_,
		_w15525_
	);
	LUT2 #(
		.INIT('h8)
	) name11479 (
		_w15518_,
		_w15525_,
		_w15526_
	);
	LUT2 #(
		.INIT('h1)
	) name11480 (
		_w15519_,
		_w15521_,
		_w15527_
	);
	LUT2 #(
		.INIT('h1)
	) name11481 (
		_w15525_,
		_w15527_,
		_w15528_
	);
	LUT2 #(
		.INIT('h1)
	) name11482 (
		_w15526_,
		_w15528_,
		_w15529_
	);
	LUT2 #(
		.INIT('h8)
	) name11483 (
		_w15467_,
		_w15529_,
		_w15530_
	);
	LUT2 #(
		.INIT('h2)
	) name11484 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14891_,
		_w15531_
	);
	LUT2 #(
		.INIT('h1)
	) name11485 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14887_,
		_w15532_
	);
	LUT2 #(
		.INIT('h1)
	) name11486 (
		_w15531_,
		_w15532_,
		_w15533_
	);
	LUT2 #(
		.INIT('h1)
	) name11487 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14861_,
		_w15534_
	);
	LUT2 #(
		.INIT('h2)
	) name11488 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14865_,
		_w15535_
	);
	LUT2 #(
		.INIT('h4)
	) name11489 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14872_,
		_w15536_
	);
	LUT2 #(
		.INIT('h8)
	) name11490 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14876_,
		_w15537_
	);
	LUT2 #(
		.INIT('h1)
	) name11491 (
		_w15536_,
		_w15537_,
		_w15538_
	);
	LUT2 #(
		.INIT('h4)
	) name11492 (
		_w15534_,
		_w15538_,
		_w15539_
	);
	LUT2 #(
		.INIT('h4)
	) name11493 (
		_w15535_,
		_w15539_,
		_w15540_
	);
	LUT2 #(
		.INIT('h1)
	) name11494 (
		_w15533_,
		_w15540_,
		_w15541_
	);
	LUT2 #(
		.INIT('h1)
	) name11495 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14887_,
		_w15542_
	);
	LUT2 #(
		.INIT('h2)
	) name11496 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14891_,
		_w15543_
	);
	LUT2 #(
		.INIT('h4)
	) name11497 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14898_,
		_w15544_
	);
	LUT2 #(
		.INIT('h8)
	) name11498 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14902_,
		_w15545_
	);
	LUT2 #(
		.INIT('h1)
	) name11499 (
		_w15544_,
		_w15545_,
		_w15546_
	);
	LUT2 #(
		.INIT('h4)
	) name11500 (
		_w15542_,
		_w15546_,
		_w15547_
	);
	LUT2 #(
		.INIT('h4)
	) name11501 (
		_w15543_,
		_w15547_,
		_w15548_
	);
	LUT2 #(
		.INIT('h1)
	) name11502 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14861_,
		_w15549_
	);
	LUT2 #(
		.INIT('h2)
	) name11503 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14865_,
		_w15550_
	);
	LUT2 #(
		.INIT('h4)
	) name11504 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14872_,
		_w15551_
	);
	LUT2 #(
		.INIT('h8)
	) name11505 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14876_,
		_w15552_
	);
	LUT2 #(
		.INIT('h1)
	) name11506 (
		_w15551_,
		_w15552_,
		_w15553_
	);
	LUT2 #(
		.INIT('h4)
	) name11507 (
		_w15549_,
		_w15553_,
		_w15554_
	);
	LUT2 #(
		.INIT('h4)
	) name11508 (
		_w15550_,
		_w15554_,
		_w15555_
	);
	LUT2 #(
		.INIT('h1)
	) name11509 (
		_w15548_,
		_w15555_,
		_w15556_
	);
	LUT2 #(
		.INIT('h8)
	) name11510 (
		_w15548_,
		_w15555_,
		_w15557_
	);
	LUT2 #(
		.INIT('h1)
	) name11511 (
		_w15556_,
		_w15557_,
		_w15558_
	);
	LUT2 #(
		.INIT('h8)
	) name11512 (
		_w15541_,
		_w15558_,
		_w15559_
	);
	LUT2 #(
		.INIT('h1)
	) name11513 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14914_,
		_w15560_
	);
	LUT2 #(
		.INIT('h2)
	) name11514 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14918_,
		_w15561_
	);
	LUT2 #(
		.INIT('h1)
	) name11515 (
		_w15560_,
		_w15561_,
		_w15562_
	);
	LUT2 #(
		.INIT('h1)
	) name11516 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14887_,
		_w15563_
	);
	LUT2 #(
		.INIT('h2)
	) name11517 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14891_,
		_w15564_
	);
	LUT2 #(
		.INIT('h4)
	) name11518 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14898_,
		_w15565_
	);
	LUT2 #(
		.INIT('h8)
	) name11519 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14902_,
		_w15566_
	);
	LUT2 #(
		.INIT('h1)
	) name11520 (
		_w15565_,
		_w15566_,
		_w15567_
	);
	LUT2 #(
		.INIT('h4)
	) name11521 (
		_w15563_,
		_w15567_,
		_w15568_
	);
	LUT2 #(
		.INIT('h4)
	) name11522 (
		_w15564_,
		_w15568_,
		_w15569_
	);
	LUT2 #(
		.INIT('h8)
	) name11523 (
		_w15562_,
		_w15569_,
		_w15570_
	);
	LUT2 #(
		.INIT('h1)
	) name11524 (
		_w15562_,
		_w15569_,
		_w15571_
	);
	LUT2 #(
		.INIT('h1)
	) name11525 (
		_w15570_,
		_w15571_,
		_w15572_
	);
	LUT2 #(
		.INIT('h1)
	) name11526 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14861_,
		_w15573_
	);
	LUT2 #(
		.INIT('h2)
	) name11527 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14865_,
		_w15574_
	);
	LUT2 #(
		.INIT('h4)
	) name11528 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14872_,
		_w15575_
	);
	LUT2 #(
		.INIT('h8)
	) name11529 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14876_,
		_w15576_
	);
	LUT2 #(
		.INIT('h1)
	) name11530 (
		_w15575_,
		_w15576_,
		_w15577_
	);
	LUT2 #(
		.INIT('h4)
	) name11531 (
		_w15573_,
		_w15577_,
		_w15578_
	);
	LUT2 #(
		.INIT('h4)
	) name11532 (
		_w15574_,
		_w15578_,
		_w15579_
	);
	LUT2 #(
		.INIT('h4)
	) name11533 (
		_w15572_,
		_w15579_,
		_w15580_
	);
	LUT2 #(
		.INIT('h2)
	) name11534 (
		_w15572_,
		_w15579_,
		_w15581_
	);
	LUT2 #(
		.INIT('h1)
	) name11535 (
		_w15580_,
		_w15581_,
		_w15582_
	);
	LUT2 #(
		.INIT('h8)
	) name11536 (
		_w15556_,
		_w15582_,
		_w15583_
	);
	LUT2 #(
		.INIT('h1)
	) name11537 (
		_w15556_,
		_w15582_,
		_w15584_
	);
	LUT2 #(
		.INIT('h1)
	) name11538 (
		_w15583_,
		_w15584_,
		_w15585_
	);
	LUT2 #(
		.INIT('h1)
	) name11539 (
		_w15559_,
		_w15585_,
		_w15586_
	);
	LUT2 #(
		.INIT('h1)
	) name11540 (
		_w15530_,
		_w15586_,
		_w15587_
	);
	LUT2 #(
		.INIT('h1)
	) name11541 (
		_w15437_,
		_w15459_,
		_w15588_
	);
	LUT2 #(
		.INIT('h1)
	) name11542 (
		_w15424_,
		_w15433_,
		_w15589_
	);
	LUT2 #(
		.INIT('h1)
	) name11543 (
		_w15425_,
		_w15589_,
		_w15590_
	);
	LUT2 #(
		.INIT('h1)
	) name11544 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14787_,
		_w15591_
	);
	LUT2 #(
		.INIT('h2)
	) name11545 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14791_,
		_w15592_
	);
	LUT2 #(
		.INIT('h4)
	) name11546 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14798_,
		_w15593_
	);
	LUT2 #(
		.INIT('h8)
	) name11547 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14802_,
		_w15594_
	);
	LUT2 #(
		.INIT('h1)
	) name11548 (
		_w15593_,
		_w15594_,
		_w15595_
	);
	LUT2 #(
		.INIT('h4)
	) name11549 (
		_w15591_,
		_w15595_,
		_w15596_
	);
	LUT2 #(
		.INIT('h4)
	) name11550 (
		_w15592_,
		_w15596_,
		_w15597_
	);
	LUT2 #(
		.INIT('h1)
	) name11551 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14761_,
		_w15598_
	);
	LUT2 #(
		.INIT('h2)
	) name11552 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14765_,
		_w15599_
	);
	LUT2 #(
		.INIT('h4)
	) name11553 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14772_,
		_w15600_
	);
	LUT2 #(
		.INIT('h8)
	) name11554 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14776_,
		_w15601_
	);
	LUT2 #(
		.INIT('h1)
	) name11555 (
		_w15600_,
		_w15601_,
		_w15602_
	);
	LUT2 #(
		.INIT('h4)
	) name11556 (
		_w15598_,
		_w15602_,
		_w15603_
	);
	LUT2 #(
		.INIT('h4)
	) name11557 (
		_w15599_,
		_w15603_,
		_w15604_
	);
	LUT2 #(
		.INIT('h8)
	) name11558 (
		_w15597_,
		_w15604_,
		_w15605_
	);
	LUT2 #(
		.INIT('h1)
	) name11559 (
		_w15597_,
		_w15604_,
		_w15606_
	);
	LUT2 #(
		.INIT('h1)
	) name11560 (
		_w15605_,
		_w15606_,
		_w15607_
	);
	LUT2 #(
		.INIT('h1)
	) name11561 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14814_,
		_w15608_
	);
	LUT2 #(
		.INIT('h2)
	) name11562 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14818_,
		_w15609_
	);
	LUT2 #(
		.INIT('h4)
	) name11563 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14825_,
		_w15610_
	);
	LUT2 #(
		.INIT('h8)
	) name11564 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14829_,
		_w15611_
	);
	LUT2 #(
		.INIT('h1)
	) name11565 (
		_w15610_,
		_w15611_,
		_w15612_
	);
	LUT2 #(
		.INIT('h4)
	) name11566 (
		_w15608_,
		_w15612_,
		_w15613_
	);
	LUT2 #(
		.INIT('h4)
	) name11567 (
		_w15609_,
		_w15613_,
		_w15614_
	);
	LUT2 #(
		.INIT('h4)
	) name11568 (
		_w15607_,
		_w15614_,
		_w15615_
	);
	LUT2 #(
		.INIT('h2)
	) name11569 (
		_w15607_,
		_w15614_,
		_w15616_
	);
	LUT2 #(
		.INIT('h1)
	) name11570 (
		_w15615_,
		_w15616_,
		_w15617_
	);
	LUT2 #(
		.INIT('h2)
	) name11571 (
		_w15590_,
		_w15617_,
		_w15618_
	);
	LUT2 #(
		.INIT('h4)
	) name11572 (
		_w15590_,
		_w15617_,
		_w15619_
	);
	LUT2 #(
		.INIT('h1)
	) name11573 (
		_w15618_,
		_w15619_,
		_w15620_
	);
	LUT2 #(
		.INIT('h4)
	) name11574 (
		_w11878_,
		_w14993_,
		_w15621_
	);
	LUT2 #(
		.INIT('h4)
	) name11575 (
		_w7182_,
		_w15044_,
		_w15622_
	);
	LUT2 #(
		.INIT('h1)
	) name11576 (
		_w15621_,
		_w15622_,
		_w15623_
	);
	LUT2 #(
		.INIT('h1)
	) name11577 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15623_,
		_w15624_
	);
	LUT2 #(
		.INIT('h1)
	) name11578 (
		_w14925_,
		_w15624_,
		_w15625_
	);
	LUT2 #(
		.INIT('h8)
	) name11579 (
		_w14925_,
		_w15624_,
		_w15626_
	);
	LUT2 #(
		.INIT('h1)
	) name11580 (
		_w15625_,
		_w15626_,
		_w15627_
	);
	LUT2 #(
		.INIT('h1)
	) name11581 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14838_,
		_w15628_
	);
	LUT2 #(
		.INIT('h2)
	) name11582 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14842_,
		_w15629_
	);
	LUT2 #(
		.INIT('h4)
	) name11583 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14846_,
		_w15630_
	);
	LUT2 #(
		.INIT('h8)
	) name11584 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14849_,
		_w15631_
	);
	LUT2 #(
		.INIT('h1)
	) name11585 (
		_w15630_,
		_w15631_,
		_w15632_
	);
	LUT2 #(
		.INIT('h4)
	) name11586 (
		_w15628_,
		_w15632_,
		_w15633_
	);
	LUT2 #(
		.INIT('h4)
	) name11587 (
		_w15629_,
		_w15633_,
		_w15634_
	);
	LUT2 #(
		.INIT('h4)
	) name11588 (
		_w15627_,
		_w15634_,
		_w15635_
	);
	LUT2 #(
		.INIT('h2)
	) name11589 (
		_w15627_,
		_w15634_,
		_w15636_
	);
	LUT2 #(
		.INIT('h1)
	) name11590 (
		_w15635_,
		_w15636_,
		_w15637_
	);
	LUT2 #(
		.INIT('h2)
	) name11591 (
		_w14914_,
		_w15453_,
		_w15638_
	);
	LUT2 #(
		.INIT('h1)
	) name11592 (
		_w15454_,
		_w15638_,
		_w15639_
	);
	LUT2 #(
		.INIT('h1)
	) name11593 (
		_w15637_,
		_w15639_,
		_w15640_
	);
	LUT2 #(
		.INIT('h8)
	) name11594 (
		_w15637_,
		_w15639_,
		_w15641_
	);
	LUT2 #(
		.INIT('h1)
	) name11595 (
		_w15640_,
		_w15641_,
		_w15642_
	);
	LUT2 #(
		.INIT('h8)
	) name11596 (
		_w15620_,
		_w15642_,
		_w15643_
	);
	LUT2 #(
		.INIT('h1)
	) name11597 (
		_w15620_,
		_w15642_,
		_w15644_
	);
	LUT2 #(
		.INIT('h1)
	) name11598 (
		_w15643_,
		_w15644_,
		_w15645_
	);
	LUT2 #(
		.INIT('h4)
	) name11599 (
		_w15588_,
		_w15645_,
		_w15646_
	);
	LUT2 #(
		.INIT('h2)
	) name11600 (
		_w15588_,
		_w15645_,
		_w15647_
	);
	LUT2 #(
		.INIT('h1)
	) name11601 (
		_w15646_,
		_w15647_,
		_w15648_
	);
	LUT2 #(
		.INIT('h1)
	) name11602 (
		_w15438_,
		_w15460_,
		_w15649_
	);
	LUT2 #(
		.INIT('h4)
	) name11603 (
		_w15464_,
		_w15649_,
		_w15650_
	);
	LUT2 #(
		.INIT('h1)
	) name11604 (
		_w15465_,
		_w15650_,
		_w15651_
	);
	LUT2 #(
		.INIT('h2)
	) name11605 (
		_w15648_,
		_w15651_,
		_w15652_
	);
	LUT2 #(
		.INIT('h4)
	) name11606 (
		_w15648_,
		_w15651_,
		_w15653_
	);
	LUT2 #(
		.INIT('h1)
	) name11607 (
		_w15652_,
		_w15653_,
		_w15654_
	);
	LUT2 #(
		.INIT('h1)
	) name11608 (
		_w15570_,
		_w15579_,
		_w15655_
	);
	LUT2 #(
		.INIT('h1)
	) name11609 (
		_w15571_,
		_w15655_,
		_w15656_
	);
	LUT2 #(
		.INIT('h1)
	) name11610 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14861_,
		_w15657_
	);
	LUT2 #(
		.INIT('h2)
	) name11611 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14865_,
		_w15658_
	);
	LUT2 #(
		.INIT('h4)
	) name11612 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14872_,
		_w15659_
	);
	LUT2 #(
		.INIT('h8)
	) name11613 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14876_,
		_w15660_
	);
	LUT2 #(
		.INIT('h1)
	) name11614 (
		_w15659_,
		_w15660_,
		_w15661_
	);
	LUT2 #(
		.INIT('h4)
	) name11615 (
		_w15657_,
		_w15661_,
		_w15662_
	);
	LUT2 #(
		.INIT('h4)
	) name11616 (
		_w15658_,
		_w15662_,
		_w15663_
	);
	LUT2 #(
		.INIT('h1)
	) name11617 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14914_,
		_w15664_
	);
	LUT2 #(
		.INIT('h2)
	) name11618 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14918_,
		_w15665_
	);
	LUT2 #(
		.INIT('h4)
	) name11619 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14925_,
		_w15666_
	);
	LUT2 #(
		.INIT('h8)
	) name11620 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14929_,
		_w15667_
	);
	LUT2 #(
		.INIT('h1)
	) name11621 (
		_w15666_,
		_w15667_,
		_w15668_
	);
	LUT2 #(
		.INIT('h4)
	) name11622 (
		_w15664_,
		_w15668_,
		_w15669_
	);
	LUT2 #(
		.INIT('h4)
	) name11623 (
		_w15665_,
		_w15669_,
		_w15670_
	);
	LUT2 #(
		.INIT('h8)
	) name11624 (
		_w15663_,
		_w15670_,
		_w15671_
	);
	LUT2 #(
		.INIT('h1)
	) name11625 (
		_w15663_,
		_w15670_,
		_w15672_
	);
	LUT2 #(
		.INIT('h1)
	) name11626 (
		_w15671_,
		_w15672_,
		_w15673_
	);
	LUT2 #(
		.INIT('h1)
	) name11627 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14887_,
		_w15674_
	);
	LUT2 #(
		.INIT('h2)
	) name11628 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14891_,
		_w15675_
	);
	LUT2 #(
		.INIT('h4)
	) name11629 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14898_,
		_w15676_
	);
	LUT2 #(
		.INIT('h8)
	) name11630 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14902_,
		_w15677_
	);
	LUT2 #(
		.INIT('h1)
	) name11631 (
		_w15676_,
		_w15677_,
		_w15678_
	);
	LUT2 #(
		.INIT('h4)
	) name11632 (
		_w15674_,
		_w15678_,
		_w15679_
	);
	LUT2 #(
		.INIT('h4)
	) name11633 (
		_w15675_,
		_w15679_,
		_w15680_
	);
	LUT2 #(
		.INIT('h4)
	) name11634 (
		_w15673_,
		_w15680_,
		_w15681_
	);
	LUT2 #(
		.INIT('h2)
	) name11635 (
		_w15673_,
		_w15680_,
		_w15682_
	);
	LUT2 #(
		.INIT('h1)
	) name11636 (
		_w15681_,
		_w15682_,
		_w15683_
	);
	LUT2 #(
		.INIT('h2)
	) name11637 (
		_w15656_,
		_w15683_,
		_w15684_
	);
	LUT2 #(
		.INIT('h4)
	) name11638 (
		_w15656_,
		_w15683_,
		_w15685_
	);
	LUT2 #(
		.INIT('h1)
	) name11639 (
		_w15684_,
		_w15685_,
		_w15686_
	);
	LUT2 #(
		.INIT('h1)
	) name11640 (
		_w15583_,
		_w15686_,
		_w15687_
	);
	LUT2 #(
		.INIT('h8)
	) name11641 (
		_w15583_,
		_w15686_,
		_w15688_
	);
	LUT2 #(
		.INIT('h1)
	) name11642 (
		_w15687_,
		_w15688_,
		_w15689_
	);
	LUT2 #(
		.INIT('h8)
	) name11643 (
		_w15654_,
		_w15689_,
		_w15690_
	);
	LUT2 #(
		.INIT('h1)
	) name11644 (
		_w15654_,
		_w15689_,
		_w15691_
	);
	LUT2 #(
		.INIT('h1)
	) name11645 (
		_w15690_,
		_w15691_,
		_w15692_
	);
	LUT2 #(
		.INIT('h2)
	) name11646 (
		_w15587_,
		_w15692_,
		_w15693_
	);
	LUT2 #(
		.INIT('h4)
	) name11647 (
		_w15587_,
		_w15692_,
		_w15694_
	);
	LUT2 #(
		.INIT('h1)
	) name11648 (
		_w15693_,
		_w15694_,
		_w15695_
	);
	LUT2 #(
		.INIT('h1)
	) name11649 (
		_w15541_,
		_w15558_,
		_w15696_
	);
	LUT2 #(
		.INIT('h1)
	) name11650 (
		_w15559_,
		_w15696_,
		_w15697_
	);
	LUT2 #(
		.INIT('h1)
	) name11651 (
		_w15518_,
		_w15525_,
		_w15698_
	);
	LUT2 #(
		.INIT('h1)
	) name11652 (
		_w15526_,
		_w15698_,
		_w15699_
	);
	LUT2 #(
		.INIT('h1)
	) name11653 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14761_,
		_w15700_
	);
	LUT2 #(
		.INIT('h2)
	) name11654 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14765_,
		_w15701_
	);
	LUT2 #(
		.INIT('h4)
	) name11655 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14772_,
		_w15702_
	);
	LUT2 #(
		.INIT('h8)
	) name11656 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14776_,
		_w15703_
	);
	LUT2 #(
		.INIT('h1)
	) name11657 (
		_w15702_,
		_w15703_,
		_w15704_
	);
	LUT2 #(
		.INIT('h4)
	) name11658 (
		_w15700_,
		_w15704_,
		_w15705_
	);
	LUT2 #(
		.INIT('h4)
	) name11659 (
		_w15701_,
		_w15705_,
		_w15706_
	);
	LUT2 #(
		.INIT('h1)
	) name11660 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14787_,
		_w15707_
	);
	LUT2 #(
		.INIT('h2)
	) name11661 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14791_,
		_w15708_
	);
	LUT2 #(
		.INIT('h4)
	) name11662 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14798_,
		_w15709_
	);
	LUT2 #(
		.INIT('h8)
	) name11663 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14802_,
		_w15710_
	);
	LUT2 #(
		.INIT('h1)
	) name11664 (
		_w15709_,
		_w15710_,
		_w15711_
	);
	LUT2 #(
		.INIT('h4)
	) name11665 (
		_w15707_,
		_w15711_,
		_w15712_
	);
	LUT2 #(
		.INIT('h4)
	) name11666 (
		_w15708_,
		_w15712_,
		_w15713_
	);
	LUT2 #(
		.INIT('h1)
	) name11667 (
		_w15706_,
		_w15713_,
		_w15714_
	);
	LUT2 #(
		.INIT('h8)
	) name11668 (
		_w15706_,
		_w15713_,
		_w15715_
	);
	LUT2 #(
		.INIT('h1)
	) name11669 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14814_,
		_w15716_
	);
	LUT2 #(
		.INIT('h2)
	) name11670 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14818_,
		_w15717_
	);
	LUT2 #(
		.INIT('h4)
	) name11671 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14825_,
		_w15718_
	);
	LUT2 #(
		.INIT('h8)
	) name11672 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14829_,
		_w15719_
	);
	LUT2 #(
		.INIT('h1)
	) name11673 (
		_w15718_,
		_w15719_,
		_w15720_
	);
	LUT2 #(
		.INIT('h4)
	) name11674 (
		_w15716_,
		_w15720_,
		_w15721_
	);
	LUT2 #(
		.INIT('h4)
	) name11675 (
		_w15717_,
		_w15721_,
		_w15722_
	);
	LUT2 #(
		.INIT('h1)
	) name11676 (
		_w15715_,
		_w15722_,
		_w15723_
	);
	LUT2 #(
		.INIT('h1)
	) name11677 (
		_w15714_,
		_w15723_,
		_w15724_
	);
	LUT2 #(
		.INIT('h1)
	) name11678 (
		_w15482_,
		_w15483_,
		_w15725_
	);
	LUT2 #(
		.INIT('h2)
	) name11679 (
		_w15490_,
		_w15725_,
		_w15726_
	);
	LUT2 #(
		.INIT('h4)
	) name11680 (
		_w15490_,
		_w15725_,
		_w15727_
	);
	LUT2 #(
		.INIT('h1)
	) name11681 (
		_w15726_,
		_w15727_,
		_w15728_
	);
	LUT2 #(
		.INIT('h2)
	) name11682 (
		_w15724_,
		_w15728_,
		_w15729_
	);
	LUT2 #(
		.INIT('h4)
	) name11683 (
		_w10112_,
		_w14993_,
		_w15730_
	);
	LUT2 #(
		.INIT('h4)
	) name11684 (
		_w10534_,
		_w15044_,
		_w15731_
	);
	LUT2 #(
		.INIT('h1)
	) name11685 (
		_w15730_,
		_w15731_,
		_w15732_
	);
	LUT2 #(
		.INIT('h1)
	) name11686 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15732_,
		_w15733_
	);
	LUT2 #(
		.INIT('h1)
	) name11687 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14838_,
		_w15734_
	);
	LUT2 #(
		.INIT('h2)
	) name11688 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14842_,
		_w15735_
	);
	LUT2 #(
		.INIT('h4)
	) name11689 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14846_,
		_w15736_
	);
	LUT2 #(
		.INIT('h8)
	) name11690 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14849_,
		_w15737_
	);
	LUT2 #(
		.INIT('h1)
	) name11691 (
		_w15736_,
		_w15737_,
		_w15738_
	);
	LUT2 #(
		.INIT('h4)
	) name11692 (
		_w15734_,
		_w15738_,
		_w15739_
	);
	LUT2 #(
		.INIT('h4)
	) name11693 (
		_w15735_,
		_w15739_,
		_w15740_
	);
	LUT2 #(
		.INIT('h4)
	) name11694 (
		_w15733_,
		_w15740_,
		_w15741_
	);
	LUT2 #(
		.INIT('h2)
	) name11695 (
		_w15733_,
		_w15740_,
		_w15742_
	);
	LUT2 #(
		.INIT('h2)
	) name11696 (
		_w14861_,
		_w15742_,
		_w15743_
	);
	LUT2 #(
		.INIT('h1)
	) name11697 (
		_w15741_,
		_w15743_,
		_w15744_
	);
	LUT2 #(
		.INIT('h1)
	) name11698 (
		_w15509_,
		_w15510_,
		_w15745_
	);
	LUT2 #(
		.INIT('h8)
	) name11699 (
		_w14872_,
		_w15745_,
		_w15746_
	);
	LUT2 #(
		.INIT('h1)
	) name11700 (
		_w14872_,
		_w15745_,
		_w15747_
	);
	LUT2 #(
		.INIT('h1)
	) name11701 (
		_w15746_,
		_w15747_,
		_w15748_
	);
	LUT2 #(
		.INIT('h1)
	) name11702 (
		_w15744_,
		_w15748_,
		_w15749_
	);
	LUT2 #(
		.INIT('h1)
	) name11703 (
		_w15729_,
		_w15749_,
		_w15750_
	);
	LUT2 #(
		.INIT('h4)
	) name11704 (
		_w15492_,
		_w15496_,
		_w15751_
	);
	LUT2 #(
		.INIT('h1)
	) name11705 (
		_w15497_,
		_w15751_,
		_w15752_
	);
	LUT2 #(
		.INIT('h8)
	) name11706 (
		_w15512_,
		_w15516_,
		_w15753_
	);
	LUT2 #(
		.INIT('h1)
	) name11707 (
		_w15517_,
		_w15753_,
		_w15754_
	);
	LUT2 #(
		.INIT('h8)
	) name11708 (
		_w15752_,
		_w15754_,
		_w15755_
	);
	LUT2 #(
		.INIT('h1)
	) name11709 (
		_w15752_,
		_w15754_,
		_w15756_
	);
	LUT2 #(
		.INIT('h1)
	) name11710 (
		_w15755_,
		_w15756_,
		_w15757_
	);
	LUT2 #(
		.INIT('h4)
	) name11711 (
		_w15750_,
		_w15757_,
		_w15758_
	);
	LUT2 #(
		.INIT('h1)
	) name11712 (
		_w15751_,
		_w15753_,
		_w15759_
	);
	LUT2 #(
		.INIT('h4)
	) name11713 (
		_w15757_,
		_w15759_,
		_w15760_
	);
	LUT2 #(
		.INIT('h1)
	) name11714 (
		_w15758_,
		_w15760_,
		_w15761_
	);
	LUT2 #(
		.INIT('h1)
	) name11715 (
		_w15699_,
		_w15761_,
		_w15762_
	);
	LUT2 #(
		.INIT('h2)
	) name11716 (
		_w15697_,
		_w15762_,
		_w15763_
	);
	LUT2 #(
		.INIT('h1)
	) name11717 (
		_w15467_,
		_w15529_,
		_w15764_
	);
	LUT2 #(
		.INIT('h1)
	) name11718 (
		_w15530_,
		_w15764_,
		_w15765_
	);
	LUT2 #(
		.INIT('h8)
	) name11719 (
		_w15559_,
		_w15582_,
		_w15766_
	);
	LUT2 #(
		.INIT('h1)
	) name11720 (
		_w15586_,
		_w15766_,
		_w15767_
	);
	LUT2 #(
		.INIT('h8)
	) name11721 (
		_w15765_,
		_w15767_,
		_w15768_
	);
	LUT2 #(
		.INIT('h1)
	) name11722 (
		_w15765_,
		_w15767_,
		_w15769_
	);
	LUT2 #(
		.INIT('h1)
	) name11723 (
		_w15768_,
		_w15769_,
		_w15770_
	);
	LUT2 #(
		.INIT('h4)
	) name11724 (
		_w15763_,
		_w15770_,
		_w15771_
	);
	LUT2 #(
		.INIT('h1)
	) name11725 (
		_w15764_,
		_w15766_,
		_w15772_
	);
	LUT2 #(
		.INIT('h4)
	) name11726 (
		_w15770_,
		_w15772_,
		_w15773_
	);
	LUT2 #(
		.INIT('h1)
	) name11727 (
		_w15771_,
		_w15773_,
		_w15774_
	);
	LUT2 #(
		.INIT('h2)
	) name11728 (
		_w15695_,
		_w15774_,
		_w15775_
	);
	LUT2 #(
		.INIT('h1)
	) name11729 (
		_w15652_,
		_w15687_,
		_w15776_
	);
	LUT2 #(
		.INIT('h4)
	) name11730 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 ,
		_w15777_
	);
	LUT2 #(
		.INIT('h2)
	) name11731 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14951_,
		_w15778_
	);
	LUT2 #(
		.INIT('h1)
	) name11732 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14947_,
		_w15779_
	);
	LUT2 #(
		.INIT('h1)
	) name11733 (
		_w15778_,
		_w15779_,
		_w15780_
	);
	LUT2 #(
		.INIT('h2)
	) name11734 (
		_w15777_,
		_w15780_,
		_w15781_
	);
	LUT2 #(
		.INIT('h4)
	) name11735 (
		_w15777_,
		_w15780_,
		_w15782_
	);
	LUT2 #(
		.INIT('h1)
	) name11736 (
		_w15781_,
		_w15782_,
		_w15783_
	);
	LUT2 #(
		.INIT('h1)
	) name11737 (
		_w15671_,
		_w15680_,
		_w15784_
	);
	LUT2 #(
		.INIT('h1)
	) name11738 (
		_w15672_,
		_w15784_,
		_w15785_
	);
	LUT2 #(
		.INIT('h1)
	) name11739 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14887_,
		_w15786_
	);
	LUT2 #(
		.INIT('h2)
	) name11740 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14891_,
		_w15787_
	);
	LUT2 #(
		.INIT('h4)
	) name11741 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14898_,
		_w15788_
	);
	LUT2 #(
		.INIT('h8)
	) name11742 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14902_,
		_w15789_
	);
	LUT2 #(
		.INIT('h1)
	) name11743 (
		_w15788_,
		_w15789_,
		_w15790_
	);
	LUT2 #(
		.INIT('h4)
	) name11744 (
		_w15786_,
		_w15790_,
		_w15791_
	);
	LUT2 #(
		.INIT('h4)
	) name11745 (
		_w15787_,
		_w15791_,
		_w15792_
	);
	LUT2 #(
		.INIT('h1)
	) name11746 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14861_,
		_w15793_
	);
	LUT2 #(
		.INIT('h2)
	) name11747 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14865_,
		_w15794_
	);
	LUT2 #(
		.INIT('h4)
	) name11748 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14872_,
		_w15795_
	);
	LUT2 #(
		.INIT('h8)
	) name11749 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14876_,
		_w15796_
	);
	LUT2 #(
		.INIT('h1)
	) name11750 (
		_w15795_,
		_w15796_,
		_w15797_
	);
	LUT2 #(
		.INIT('h4)
	) name11751 (
		_w15793_,
		_w15797_,
		_w15798_
	);
	LUT2 #(
		.INIT('h4)
	) name11752 (
		_w15794_,
		_w15798_,
		_w15799_
	);
	LUT2 #(
		.INIT('h8)
	) name11753 (
		_w15792_,
		_w15799_,
		_w15800_
	);
	LUT2 #(
		.INIT('h1)
	) name11754 (
		_w15792_,
		_w15799_,
		_w15801_
	);
	LUT2 #(
		.INIT('h1)
	) name11755 (
		_w15800_,
		_w15801_,
		_w15802_
	);
	LUT2 #(
		.INIT('h1)
	) name11756 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14914_,
		_w15803_
	);
	LUT2 #(
		.INIT('h2)
	) name11757 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14918_,
		_w15804_
	);
	LUT2 #(
		.INIT('h4)
	) name11758 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14925_,
		_w15805_
	);
	LUT2 #(
		.INIT('h8)
	) name11759 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14929_,
		_w15806_
	);
	LUT2 #(
		.INIT('h1)
	) name11760 (
		_w15805_,
		_w15806_,
		_w15807_
	);
	LUT2 #(
		.INIT('h4)
	) name11761 (
		_w15803_,
		_w15807_,
		_w15808_
	);
	LUT2 #(
		.INIT('h4)
	) name11762 (
		_w15804_,
		_w15808_,
		_w15809_
	);
	LUT2 #(
		.INIT('h4)
	) name11763 (
		_w15802_,
		_w15809_,
		_w15810_
	);
	LUT2 #(
		.INIT('h2)
	) name11764 (
		_w15802_,
		_w15809_,
		_w15811_
	);
	LUT2 #(
		.INIT('h1)
	) name11765 (
		_w15810_,
		_w15811_,
		_w15812_
	);
	LUT2 #(
		.INIT('h4)
	) name11766 (
		_w15785_,
		_w15812_,
		_w15813_
	);
	LUT2 #(
		.INIT('h2)
	) name11767 (
		_w15785_,
		_w15812_,
		_w15814_
	);
	LUT2 #(
		.INIT('h1)
	) name11768 (
		_w15813_,
		_w15814_,
		_w15815_
	);
	LUT2 #(
		.INIT('h8)
	) name11769 (
		_w15783_,
		_w15815_,
		_w15816_
	);
	LUT2 #(
		.INIT('h1)
	) name11770 (
		_w15783_,
		_w15815_,
		_w15817_
	);
	LUT2 #(
		.INIT('h1)
	) name11771 (
		_w15816_,
		_w15817_,
		_w15818_
	);
	LUT2 #(
		.INIT('h1)
	) name11772 (
		_w15685_,
		_w15818_,
		_w15819_
	);
	LUT2 #(
		.INIT('h8)
	) name11773 (
		_w15685_,
		_w15818_,
		_w15820_
	);
	LUT2 #(
		.INIT('h1)
	) name11774 (
		_w15819_,
		_w15820_,
		_w15821_
	);
	LUT2 #(
		.INIT('h1)
	) name11775 (
		_w15618_,
		_w15640_,
		_w15822_
	);
	LUT2 #(
		.INIT('h1)
	) name11776 (
		_w15605_,
		_w15614_,
		_w15823_
	);
	LUT2 #(
		.INIT('h1)
	) name11777 (
		_w15606_,
		_w15823_,
		_w15824_
	);
	LUT2 #(
		.INIT('h1)
	) name11778 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14787_,
		_w15825_
	);
	LUT2 #(
		.INIT('h2)
	) name11779 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14791_,
		_w15826_
	);
	LUT2 #(
		.INIT('h4)
	) name11780 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14798_,
		_w15827_
	);
	LUT2 #(
		.INIT('h8)
	) name11781 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14802_,
		_w15828_
	);
	LUT2 #(
		.INIT('h1)
	) name11782 (
		_w15827_,
		_w15828_,
		_w15829_
	);
	LUT2 #(
		.INIT('h4)
	) name11783 (
		_w15825_,
		_w15829_,
		_w15830_
	);
	LUT2 #(
		.INIT('h4)
	) name11784 (
		_w15826_,
		_w15830_,
		_w15831_
	);
	LUT2 #(
		.INIT('h1)
	) name11785 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14761_,
		_w15832_
	);
	LUT2 #(
		.INIT('h2)
	) name11786 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14765_,
		_w15833_
	);
	LUT2 #(
		.INIT('h4)
	) name11787 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14772_,
		_w15834_
	);
	LUT2 #(
		.INIT('h8)
	) name11788 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14776_,
		_w15835_
	);
	LUT2 #(
		.INIT('h1)
	) name11789 (
		_w15834_,
		_w15835_,
		_w15836_
	);
	LUT2 #(
		.INIT('h4)
	) name11790 (
		_w15832_,
		_w15836_,
		_w15837_
	);
	LUT2 #(
		.INIT('h4)
	) name11791 (
		_w15833_,
		_w15837_,
		_w15838_
	);
	LUT2 #(
		.INIT('h8)
	) name11792 (
		_w15831_,
		_w15838_,
		_w15839_
	);
	LUT2 #(
		.INIT('h1)
	) name11793 (
		_w15831_,
		_w15838_,
		_w15840_
	);
	LUT2 #(
		.INIT('h1)
	) name11794 (
		_w15839_,
		_w15840_,
		_w15841_
	);
	LUT2 #(
		.INIT('h1)
	) name11795 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14814_,
		_w15842_
	);
	LUT2 #(
		.INIT('h2)
	) name11796 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14818_,
		_w15843_
	);
	LUT2 #(
		.INIT('h4)
	) name11797 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14825_,
		_w15844_
	);
	LUT2 #(
		.INIT('h8)
	) name11798 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14829_,
		_w15845_
	);
	LUT2 #(
		.INIT('h1)
	) name11799 (
		_w15844_,
		_w15845_,
		_w15846_
	);
	LUT2 #(
		.INIT('h4)
	) name11800 (
		_w15842_,
		_w15846_,
		_w15847_
	);
	LUT2 #(
		.INIT('h4)
	) name11801 (
		_w15843_,
		_w15847_,
		_w15848_
	);
	LUT2 #(
		.INIT('h4)
	) name11802 (
		_w15841_,
		_w15848_,
		_w15849_
	);
	LUT2 #(
		.INIT('h2)
	) name11803 (
		_w15841_,
		_w15848_,
		_w15850_
	);
	LUT2 #(
		.INIT('h1)
	) name11804 (
		_w15849_,
		_w15850_,
		_w15851_
	);
	LUT2 #(
		.INIT('h2)
	) name11805 (
		_w15824_,
		_w15851_,
		_w15852_
	);
	LUT2 #(
		.INIT('h4)
	) name11806 (
		_w15824_,
		_w15851_,
		_w15853_
	);
	LUT2 #(
		.INIT('h1)
	) name11807 (
		_w15852_,
		_w15853_,
		_w15854_
	);
	LUT2 #(
		.INIT('h1)
	) name11808 (
		_w15625_,
		_w15634_,
		_w15855_
	);
	LUT2 #(
		.INIT('h1)
	) name11809 (
		_w15626_,
		_w15855_,
		_w15856_
	);
	LUT2 #(
		.INIT('h4)
	) name11810 (
		_w12024_,
		_w14993_,
		_w15857_
	);
	LUT2 #(
		.INIT('h4)
	) name11811 (
		_w11878_,
		_w15044_,
		_w15858_
	);
	LUT2 #(
		.INIT('h1)
	) name11812 (
		_w15857_,
		_w15858_,
		_w15859_
	);
	LUT2 #(
		.INIT('h1)
	) name11813 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15859_,
		_w15860_
	);
	LUT2 #(
		.INIT('h1)
	) name11814 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14838_,
		_w15861_
	);
	LUT2 #(
		.INIT('h2)
	) name11815 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14842_,
		_w15862_
	);
	LUT2 #(
		.INIT('h4)
	) name11816 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14846_,
		_w15863_
	);
	LUT2 #(
		.INIT('h8)
	) name11817 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14849_,
		_w15864_
	);
	LUT2 #(
		.INIT('h1)
	) name11818 (
		_w15863_,
		_w15864_,
		_w15865_
	);
	LUT2 #(
		.INIT('h4)
	) name11819 (
		_w15861_,
		_w15865_,
		_w15866_
	);
	LUT2 #(
		.INIT('h4)
	) name11820 (
		_w15862_,
		_w15866_,
		_w15867_
	);
	LUT2 #(
		.INIT('h4)
	) name11821 (
		_w15860_,
		_w15867_,
		_w15868_
	);
	LUT2 #(
		.INIT('h2)
	) name11822 (
		_w15860_,
		_w15867_,
		_w15869_
	);
	LUT2 #(
		.INIT('h1)
	) name11823 (
		_w15868_,
		_w15869_,
		_w15870_
	);
	LUT2 #(
		.INIT('h8)
	) name11824 (
		_w14947_,
		_w15870_,
		_w15871_
	);
	LUT2 #(
		.INIT('h1)
	) name11825 (
		_w14947_,
		_w15870_,
		_w15872_
	);
	LUT2 #(
		.INIT('h1)
	) name11826 (
		_w15871_,
		_w15872_,
		_w15873_
	);
	LUT2 #(
		.INIT('h8)
	) name11827 (
		_w15856_,
		_w15873_,
		_w15874_
	);
	LUT2 #(
		.INIT('h1)
	) name11828 (
		_w15856_,
		_w15873_,
		_w15875_
	);
	LUT2 #(
		.INIT('h1)
	) name11829 (
		_w15874_,
		_w15875_,
		_w15876_
	);
	LUT2 #(
		.INIT('h8)
	) name11830 (
		_w15854_,
		_w15876_,
		_w15877_
	);
	LUT2 #(
		.INIT('h1)
	) name11831 (
		_w15854_,
		_w15876_,
		_w15878_
	);
	LUT2 #(
		.INIT('h1)
	) name11832 (
		_w15877_,
		_w15878_,
		_w15879_
	);
	LUT2 #(
		.INIT('h4)
	) name11833 (
		_w15822_,
		_w15879_,
		_w15880_
	);
	LUT2 #(
		.INIT('h2)
	) name11834 (
		_w15822_,
		_w15879_,
		_w15881_
	);
	LUT2 #(
		.INIT('h1)
	) name11835 (
		_w15880_,
		_w15881_,
		_w15882_
	);
	LUT2 #(
		.INIT('h1)
	) name11836 (
		_w15619_,
		_w15641_,
		_w15883_
	);
	LUT2 #(
		.INIT('h4)
	) name11837 (
		_w15645_,
		_w15883_,
		_w15884_
	);
	LUT2 #(
		.INIT('h1)
	) name11838 (
		_w15646_,
		_w15884_,
		_w15885_
	);
	LUT2 #(
		.INIT('h2)
	) name11839 (
		_w15882_,
		_w15885_,
		_w15886_
	);
	LUT2 #(
		.INIT('h4)
	) name11840 (
		_w15882_,
		_w15885_,
		_w15887_
	);
	LUT2 #(
		.INIT('h1)
	) name11841 (
		_w15886_,
		_w15887_,
		_w15888_
	);
	LUT2 #(
		.INIT('h8)
	) name11842 (
		_w15821_,
		_w15888_,
		_w15889_
	);
	LUT2 #(
		.INIT('h1)
	) name11843 (
		_w15821_,
		_w15888_,
		_w15890_
	);
	LUT2 #(
		.INIT('h1)
	) name11844 (
		_w15889_,
		_w15890_,
		_w15891_
	);
	LUT2 #(
		.INIT('h4)
	) name11845 (
		_w15776_,
		_w15891_,
		_w15892_
	);
	LUT2 #(
		.INIT('h2)
	) name11846 (
		_w15776_,
		_w15891_,
		_w15893_
	);
	LUT2 #(
		.INIT('h1)
	) name11847 (
		_w15892_,
		_w15893_,
		_w15894_
	);
	LUT2 #(
		.INIT('h1)
	) name11848 (
		_w15653_,
		_w15688_,
		_w15895_
	);
	LUT2 #(
		.INIT('h4)
	) name11849 (
		_w15692_,
		_w15895_,
		_w15896_
	);
	LUT2 #(
		.INIT('h1)
	) name11850 (
		_w15694_,
		_w15896_,
		_w15897_
	);
	LUT2 #(
		.INIT('h2)
	) name11851 (
		_w15894_,
		_w15897_,
		_w15898_
	);
	LUT2 #(
		.INIT('h1)
	) name11852 (
		_w15775_,
		_w15898_,
		_w15899_
	);
	LUT2 #(
		.INIT('h8)
	) name11853 (
		_w15533_,
		_w15540_,
		_w15900_
	);
	LUT2 #(
		.INIT('h1)
	) name11854 (
		_w15541_,
		_w15900_,
		_w15901_
	);
	LUT2 #(
		.INIT('h2)
	) name11855 (
		_w15750_,
		_w15757_,
		_w15902_
	);
	LUT2 #(
		.INIT('h1)
	) name11856 (
		_w15758_,
		_w15902_,
		_w15903_
	);
	LUT2 #(
		.INIT('h1)
	) name11857 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14761_,
		_w15904_
	);
	LUT2 #(
		.INIT('h2)
	) name11858 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14765_,
		_w15905_
	);
	LUT2 #(
		.INIT('h4)
	) name11859 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14772_,
		_w15906_
	);
	LUT2 #(
		.INIT('h8)
	) name11860 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14776_,
		_w15907_
	);
	LUT2 #(
		.INIT('h1)
	) name11861 (
		_w15906_,
		_w15907_,
		_w15908_
	);
	LUT2 #(
		.INIT('h4)
	) name11862 (
		_w15904_,
		_w15908_,
		_w15909_
	);
	LUT2 #(
		.INIT('h4)
	) name11863 (
		_w15905_,
		_w15909_,
		_w15910_
	);
	LUT2 #(
		.INIT('h1)
	) name11864 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14787_,
		_w15911_
	);
	LUT2 #(
		.INIT('h2)
	) name11865 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14791_,
		_w15912_
	);
	LUT2 #(
		.INIT('h4)
	) name11866 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14798_,
		_w15913_
	);
	LUT2 #(
		.INIT('h8)
	) name11867 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14802_,
		_w15914_
	);
	LUT2 #(
		.INIT('h1)
	) name11868 (
		_w15913_,
		_w15914_,
		_w15915_
	);
	LUT2 #(
		.INIT('h4)
	) name11869 (
		_w15911_,
		_w15915_,
		_w15916_
	);
	LUT2 #(
		.INIT('h4)
	) name11870 (
		_w15912_,
		_w15916_,
		_w15917_
	);
	LUT2 #(
		.INIT('h1)
	) name11871 (
		_w15910_,
		_w15917_,
		_w15918_
	);
	LUT2 #(
		.INIT('h8)
	) name11872 (
		_w15910_,
		_w15917_,
		_w15919_
	);
	LUT2 #(
		.INIT('h1)
	) name11873 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14814_,
		_w15920_
	);
	LUT2 #(
		.INIT('h2)
	) name11874 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14818_,
		_w15921_
	);
	LUT2 #(
		.INIT('h4)
	) name11875 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14825_,
		_w15922_
	);
	LUT2 #(
		.INIT('h8)
	) name11876 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14829_,
		_w15923_
	);
	LUT2 #(
		.INIT('h1)
	) name11877 (
		_w15922_,
		_w15923_,
		_w15924_
	);
	LUT2 #(
		.INIT('h4)
	) name11878 (
		_w15920_,
		_w15924_,
		_w15925_
	);
	LUT2 #(
		.INIT('h4)
	) name11879 (
		_w15921_,
		_w15925_,
		_w15926_
	);
	LUT2 #(
		.INIT('h1)
	) name11880 (
		_w15919_,
		_w15926_,
		_w15927_
	);
	LUT2 #(
		.INIT('h1)
	) name11881 (
		_w15918_,
		_w15927_,
		_w15928_
	);
	LUT2 #(
		.INIT('h1)
	) name11882 (
		_w15714_,
		_w15715_,
		_w15929_
	);
	LUT2 #(
		.INIT('h2)
	) name11883 (
		_w15722_,
		_w15929_,
		_w15930_
	);
	LUT2 #(
		.INIT('h4)
	) name11884 (
		_w15722_,
		_w15929_,
		_w15931_
	);
	LUT2 #(
		.INIT('h1)
	) name11885 (
		_w15930_,
		_w15931_,
		_w15932_
	);
	LUT2 #(
		.INIT('h2)
	) name11886 (
		_w15928_,
		_w15932_,
		_w15933_
	);
	LUT2 #(
		.INIT('h1)
	) name11887 (
		_w15741_,
		_w15742_,
		_w15934_
	);
	LUT2 #(
		.INIT('h2)
	) name11888 (
		_w14861_,
		_w15934_,
		_w15935_
	);
	LUT2 #(
		.INIT('h4)
	) name11889 (
		_w14861_,
		_w15934_,
		_w15936_
	);
	LUT2 #(
		.INIT('h1)
	) name11890 (
		_w15935_,
		_w15936_,
		_w15937_
	);
	LUT2 #(
		.INIT('h1)
	) name11891 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14838_,
		_w15938_
	);
	LUT2 #(
		.INIT('h2)
	) name11892 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14842_,
		_w15939_
	);
	LUT2 #(
		.INIT('h4)
	) name11893 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14846_,
		_w15940_
	);
	LUT2 #(
		.INIT('h8)
	) name11894 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14849_,
		_w15941_
	);
	LUT2 #(
		.INIT('h1)
	) name11895 (
		_w15940_,
		_w15941_,
		_w15942_
	);
	LUT2 #(
		.INIT('h4)
	) name11896 (
		_w15938_,
		_w15942_,
		_w15943_
	);
	LUT2 #(
		.INIT('h4)
	) name11897 (
		_w15939_,
		_w15943_,
		_w15944_
	);
	LUT2 #(
		.INIT('h4)
	) name11898 (
		_w14825_,
		_w15944_,
		_w15945_
	);
	LUT2 #(
		.INIT('h4)
	) name11899 (
		_w10534_,
		_w14993_,
		_w15946_
	);
	LUT2 #(
		.INIT('h4)
	) name11900 (
		_w11192_,
		_w15044_,
		_w15947_
	);
	LUT2 #(
		.INIT('h1)
	) name11901 (
		_w15946_,
		_w15947_,
		_w15948_
	);
	LUT2 #(
		.INIT('h1)
	) name11902 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w15948_,
		_w15949_
	);
	LUT2 #(
		.INIT('h2)
	) name11903 (
		_w14825_,
		_w15944_,
		_w15950_
	);
	LUT2 #(
		.INIT('h1)
	) name11904 (
		_w15949_,
		_w15950_,
		_w15951_
	);
	LUT2 #(
		.INIT('h1)
	) name11905 (
		_w15945_,
		_w15951_,
		_w15952_
	);
	LUT2 #(
		.INIT('h1)
	) name11906 (
		_w15937_,
		_w15952_,
		_w15953_
	);
	LUT2 #(
		.INIT('h1)
	) name11907 (
		_w15933_,
		_w15953_,
		_w15954_
	);
	LUT2 #(
		.INIT('h4)
	) name11908 (
		_w15724_,
		_w15728_,
		_w15955_
	);
	LUT2 #(
		.INIT('h1)
	) name11909 (
		_w15729_,
		_w15955_,
		_w15956_
	);
	LUT2 #(
		.INIT('h8)
	) name11910 (
		_w15744_,
		_w15748_,
		_w15957_
	);
	LUT2 #(
		.INIT('h1)
	) name11911 (
		_w15749_,
		_w15957_,
		_w15958_
	);
	LUT2 #(
		.INIT('h8)
	) name11912 (
		_w15956_,
		_w15958_,
		_w15959_
	);
	LUT2 #(
		.INIT('h1)
	) name11913 (
		_w15956_,
		_w15958_,
		_w15960_
	);
	LUT2 #(
		.INIT('h1)
	) name11914 (
		_w15959_,
		_w15960_,
		_w15961_
	);
	LUT2 #(
		.INIT('h4)
	) name11915 (
		_w15954_,
		_w15961_,
		_w15962_
	);
	LUT2 #(
		.INIT('h1)
	) name11916 (
		_w15955_,
		_w15957_,
		_w15963_
	);
	LUT2 #(
		.INIT('h4)
	) name11917 (
		_w15961_,
		_w15963_,
		_w15964_
	);
	LUT2 #(
		.INIT('h1)
	) name11918 (
		_w15962_,
		_w15964_,
		_w15965_
	);
	LUT2 #(
		.INIT('h2)
	) name11919 (
		_w15903_,
		_w15965_,
		_w15966_
	);
	LUT2 #(
		.INIT('h2)
	) name11920 (
		_w15901_,
		_w15966_,
		_w15967_
	);
	LUT2 #(
		.INIT('h8)
	) name11921 (
		_w15699_,
		_w15761_,
		_w15968_
	);
	LUT2 #(
		.INIT('h1)
	) name11922 (
		_w15762_,
		_w15968_,
		_w15969_
	);
	LUT2 #(
		.INIT('h2)
	) name11923 (
		_w15697_,
		_w15969_,
		_w15970_
	);
	LUT2 #(
		.INIT('h4)
	) name11924 (
		_w15697_,
		_w15969_,
		_w15971_
	);
	LUT2 #(
		.INIT('h1)
	) name11925 (
		_w15970_,
		_w15971_,
		_w15972_
	);
	LUT2 #(
		.INIT('h1)
	) name11926 (
		_w15967_,
		_w15972_,
		_w15973_
	);
	LUT2 #(
		.INIT('h4)
	) name11927 (
		_w15968_,
		_w15972_,
		_w15974_
	);
	LUT2 #(
		.INIT('h1)
	) name11928 (
		_w15973_,
		_w15974_,
		_w15975_
	);
	LUT2 #(
		.INIT('h2)
	) name11929 (
		_w15763_,
		_w15770_,
		_w15976_
	);
	LUT2 #(
		.INIT('h1)
	) name11930 (
		_w15771_,
		_w15976_,
		_w15977_
	);
	LUT2 #(
		.INIT('h4)
	) name11931 (
		_w15975_,
		_w15977_,
		_w15978_
	);
	LUT2 #(
		.INIT('h2)
	) name11932 (
		_w15954_,
		_w15961_,
		_w15979_
	);
	LUT2 #(
		.INIT('h1)
	) name11933 (
		_w15962_,
		_w15979_,
		_w15980_
	);
	LUT2 #(
		.INIT('h1)
	) name11934 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14814_,
		_w15981_
	);
	LUT2 #(
		.INIT('h2)
	) name11935 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14818_,
		_w15982_
	);
	LUT2 #(
		.INIT('h1)
	) name11936 (
		_w15981_,
		_w15982_,
		_w15983_
	);
	LUT2 #(
		.INIT('h1)
	) name11937 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14761_,
		_w15984_
	);
	LUT2 #(
		.INIT('h2)
	) name11938 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14765_,
		_w15985_
	);
	LUT2 #(
		.INIT('h4)
	) name11939 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14772_,
		_w15986_
	);
	LUT2 #(
		.INIT('h8)
	) name11940 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14776_,
		_w15987_
	);
	LUT2 #(
		.INIT('h1)
	) name11941 (
		_w15986_,
		_w15987_,
		_w15988_
	);
	LUT2 #(
		.INIT('h4)
	) name11942 (
		_w15984_,
		_w15988_,
		_w15989_
	);
	LUT2 #(
		.INIT('h4)
	) name11943 (
		_w15985_,
		_w15989_,
		_w15990_
	);
	LUT2 #(
		.INIT('h1)
	) name11944 (
		_w15983_,
		_w15990_,
		_w15991_
	);
	LUT2 #(
		.INIT('h8)
	) name11945 (
		_w15983_,
		_w15990_,
		_w15992_
	);
	LUT2 #(
		.INIT('h1)
	) name11946 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14787_,
		_w15993_
	);
	LUT2 #(
		.INIT('h2)
	) name11947 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14791_,
		_w15994_
	);
	LUT2 #(
		.INIT('h4)
	) name11948 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14798_,
		_w15995_
	);
	LUT2 #(
		.INIT('h8)
	) name11949 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14802_,
		_w15996_
	);
	LUT2 #(
		.INIT('h1)
	) name11950 (
		_w15995_,
		_w15996_,
		_w15997_
	);
	LUT2 #(
		.INIT('h4)
	) name11951 (
		_w15993_,
		_w15997_,
		_w15998_
	);
	LUT2 #(
		.INIT('h4)
	) name11952 (
		_w15994_,
		_w15998_,
		_w15999_
	);
	LUT2 #(
		.INIT('h1)
	) name11953 (
		_w15992_,
		_w15999_,
		_w16000_
	);
	LUT2 #(
		.INIT('h1)
	) name11954 (
		_w15991_,
		_w16000_,
		_w16001_
	);
	LUT2 #(
		.INIT('h1)
	) name11955 (
		_w15918_,
		_w15919_,
		_w16002_
	);
	LUT2 #(
		.INIT('h2)
	) name11956 (
		_w15926_,
		_w16002_,
		_w16003_
	);
	LUT2 #(
		.INIT('h4)
	) name11957 (
		_w15926_,
		_w16002_,
		_w16004_
	);
	LUT2 #(
		.INIT('h1)
	) name11958 (
		_w16003_,
		_w16004_,
		_w16005_
	);
	LUT2 #(
		.INIT('h2)
	) name11959 (
		_w16001_,
		_w16005_,
		_w16006_
	);
	LUT2 #(
		.INIT('h1)
	) name11960 (
		_w15945_,
		_w15950_,
		_w16007_
	);
	LUT2 #(
		.INIT('h8)
	) name11961 (
		_w15949_,
		_w16007_,
		_w16008_
	);
	LUT2 #(
		.INIT('h1)
	) name11962 (
		_w15949_,
		_w16007_,
		_w16009_
	);
	LUT2 #(
		.INIT('h1)
	) name11963 (
		_w16008_,
		_w16009_,
		_w16010_
	);
	LUT2 #(
		.INIT('h4)
	) name11964 (
		_w11192_,
		_w14993_,
		_w16011_
	);
	LUT2 #(
		.INIT('h4)
	) name11965 (
		_w11444_,
		_w15044_,
		_w16012_
	);
	LUT2 #(
		.INIT('h1)
	) name11966 (
		_w16011_,
		_w16012_,
		_w16013_
	);
	LUT2 #(
		.INIT('h1)
	) name11967 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16013_,
		_w16014_
	);
	LUT2 #(
		.INIT('h4)
	) name11968 (
		_w14814_,
		_w16014_,
		_w16015_
	);
	LUT2 #(
		.INIT('h2)
	) name11969 (
		_w14814_,
		_w16014_,
		_w16016_
	);
	LUT2 #(
		.INIT('h1)
	) name11970 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14838_,
		_w16017_
	);
	LUT2 #(
		.INIT('h2)
	) name11971 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14842_,
		_w16018_
	);
	LUT2 #(
		.INIT('h4)
	) name11972 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14846_,
		_w16019_
	);
	LUT2 #(
		.INIT('h8)
	) name11973 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14849_,
		_w16020_
	);
	LUT2 #(
		.INIT('h1)
	) name11974 (
		_w16019_,
		_w16020_,
		_w16021_
	);
	LUT2 #(
		.INIT('h4)
	) name11975 (
		_w16017_,
		_w16021_,
		_w16022_
	);
	LUT2 #(
		.INIT('h4)
	) name11976 (
		_w16018_,
		_w16022_,
		_w16023_
	);
	LUT2 #(
		.INIT('h1)
	) name11977 (
		_w16016_,
		_w16023_,
		_w16024_
	);
	LUT2 #(
		.INIT('h1)
	) name11978 (
		_w16015_,
		_w16024_,
		_w16025_
	);
	LUT2 #(
		.INIT('h4)
	) name11979 (
		_w16010_,
		_w16025_,
		_w16026_
	);
	LUT2 #(
		.INIT('h1)
	) name11980 (
		_w16006_,
		_w16026_,
		_w16027_
	);
	LUT2 #(
		.INIT('h4)
	) name11981 (
		_w15928_,
		_w15932_,
		_w16028_
	);
	LUT2 #(
		.INIT('h1)
	) name11982 (
		_w15933_,
		_w16028_,
		_w16029_
	);
	LUT2 #(
		.INIT('h8)
	) name11983 (
		_w15937_,
		_w15952_,
		_w16030_
	);
	LUT2 #(
		.INIT('h1)
	) name11984 (
		_w15953_,
		_w16030_,
		_w16031_
	);
	LUT2 #(
		.INIT('h8)
	) name11985 (
		_w16029_,
		_w16031_,
		_w16032_
	);
	LUT2 #(
		.INIT('h1)
	) name11986 (
		_w16029_,
		_w16031_,
		_w16033_
	);
	LUT2 #(
		.INIT('h1)
	) name11987 (
		_w16032_,
		_w16033_,
		_w16034_
	);
	LUT2 #(
		.INIT('h4)
	) name11988 (
		_w16027_,
		_w16034_,
		_w16035_
	);
	LUT2 #(
		.INIT('h1)
	) name11989 (
		_w16028_,
		_w16030_,
		_w16036_
	);
	LUT2 #(
		.INIT('h4)
	) name11990 (
		_w16034_,
		_w16036_,
		_w16037_
	);
	LUT2 #(
		.INIT('h1)
	) name11991 (
		_w16035_,
		_w16037_,
		_w16038_
	);
	LUT2 #(
		.INIT('h2)
	) name11992 (
		_w15980_,
		_w16038_,
		_w16039_
	);
	LUT2 #(
		.INIT('h1)
	) name11993 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14861_,
		_w16040_
	);
	LUT2 #(
		.INIT('h2)
	) name11994 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14865_,
		_w16041_
	);
	LUT2 #(
		.INIT('h4)
	) name11995 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14872_,
		_w16042_
	);
	LUT2 #(
		.INIT('h8)
	) name11996 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14876_,
		_w16043_
	);
	LUT2 #(
		.INIT('h1)
	) name11997 (
		_w16042_,
		_w16043_,
		_w16044_
	);
	LUT2 #(
		.INIT('h4)
	) name11998 (
		_w16040_,
		_w16044_,
		_w16045_
	);
	LUT2 #(
		.INIT('h4)
	) name11999 (
		_w16041_,
		_w16045_,
		_w16046_
	);
	LUT2 #(
		.INIT('h1)
	) name12000 (
		_w16039_,
		_w16046_,
		_w16047_
	);
	LUT2 #(
		.INIT('h4)
	) name12001 (
		_w15903_,
		_w15965_,
		_w16048_
	);
	LUT2 #(
		.INIT('h1)
	) name12002 (
		_w15966_,
		_w16048_,
		_w16049_
	);
	LUT2 #(
		.INIT('h1)
	) name12003 (
		_w15901_,
		_w16049_,
		_w16050_
	);
	LUT2 #(
		.INIT('h8)
	) name12004 (
		_w15901_,
		_w16049_,
		_w16051_
	);
	LUT2 #(
		.INIT('h1)
	) name12005 (
		_w16050_,
		_w16051_,
		_w16052_
	);
	LUT2 #(
		.INIT('h4)
	) name12006 (
		_w16047_,
		_w16052_,
		_w16053_
	);
	LUT2 #(
		.INIT('h1)
	) name12007 (
		_w16048_,
		_w16052_,
		_w16054_
	);
	LUT2 #(
		.INIT('h1)
	) name12008 (
		_w16053_,
		_w16054_,
		_w16055_
	);
	LUT2 #(
		.INIT('h8)
	) name12009 (
		_w15967_,
		_w15972_,
		_w16056_
	);
	LUT2 #(
		.INIT('h1)
	) name12010 (
		_w15973_,
		_w16056_,
		_w16057_
	);
	LUT2 #(
		.INIT('h4)
	) name12011 (
		_w16055_,
		_w16057_,
		_w16058_
	);
	LUT2 #(
		.INIT('h1)
	) name12012 (
		_w15978_,
		_w16058_,
		_w16059_
	);
	LUT2 #(
		.INIT('h1)
	) name12013 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14787_,
		_w16060_
	);
	LUT2 #(
		.INIT('h2)
	) name12014 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14791_,
		_w16061_
	);
	LUT2 #(
		.INIT('h4)
	) name12015 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14798_,
		_w16062_
	);
	LUT2 #(
		.INIT('h8)
	) name12016 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14802_,
		_w16063_
	);
	LUT2 #(
		.INIT('h1)
	) name12017 (
		_w16062_,
		_w16063_,
		_w16064_
	);
	LUT2 #(
		.INIT('h4)
	) name12018 (
		_w16060_,
		_w16064_,
		_w16065_
	);
	LUT2 #(
		.INIT('h4)
	) name12019 (
		_w16061_,
		_w16065_,
		_w16066_
	);
	LUT2 #(
		.INIT('h1)
	) name12020 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14761_,
		_w16067_
	);
	LUT2 #(
		.INIT('h2)
	) name12021 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14765_,
		_w16068_
	);
	LUT2 #(
		.INIT('h4)
	) name12022 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14772_,
		_w16069_
	);
	LUT2 #(
		.INIT('h8)
	) name12023 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14776_,
		_w16070_
	);
	LUT2 #(
		.INIT('h1)
	) name12024 (
		_w16069_,
		_w16070_,
		_w16071_
	);
	LUT2 #(
		.INIT('h4)
	) name12025 (
		_w16067_,
		_w16071_,
		_w16072_
	);
	LUT2 #(
		.INIT('h4)
	) name12026 (
		_w16068_,
		_w16072_,
		_w16073_
	);
	LUT2 #(
		.INIT('h1)
	) name12027 (
		_w16066_,
		_w16073_,
		_w16074_
	);
	LUT2 #(
		.INIT('h1)
	) name12028 (
		_w15991_,
		_w15992_,
		_w16075_
	);
	LUT2 #(
		.INIT('h2)
	) name12029 (
		_w15999_,
		_w16075_,
		_w16076_
	);
	LUT2 #(
		.INIT('h4)
	) name12030 (
		_w15999_,
		_w16075_,
		_w16077_
	);
	LUT2 #(
		.INIT('h1)
	) name12031 (
		_w16076_,
		_w16077_,
		_w16078_
	);
	LUT2 #(
		.INIT('h1)
	) name12032 (
		_w16074_,
		_w16078_,
		_w16079_
	);
	LUT2 #(
		.INIT('h4)
	) name12033 (
		_w11444_,
		_w14993_,
		_w16080_
	);
	LUT2 #(
		.INIT('h4)
	) name12034 (
		_w10878_,
		_w15044_,
		_w16081_
	);
	LUT2 #(
		.INIT('h1)
	) name12035 (
		_w16080_,
		_w16081_,
		_w16082_
	);
	LUT2 #(
		.INIT('h1)
	) name12036 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16082_,
		_w16083_
	);
	LUT2 #(
		.INIT('h1)
	) name12037 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14838_,
		_w16084_
	);
	LUT2 #(
		.INIT('h2)
	) name12038 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14842_,
		_w16085_
	);
	LUT2 #(
		.INIT('h4)
	) name12039 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14846_,
		_w16086_
	);
	LUT2 #(
		.INIT('h8)
	) name12040 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14849_,
		_w16087_
	);
	LUT2 #(
		.INIT('h1)
	) name12041 (
		_w16086_,
		_w16087_,
		_w16088_
	);
	LUT2 #(
		.INIT('h4)
	) name12042 (
		_w16084_,
		_w16088_,
		_w16089_
	);
	LUT2 #(
		.INIT('h4)
	) name12043 (
		_w16085_,
		_w16089_,
		_w16090_
	);
	LUT2 #(
		.INIT('h4)
	) name12044 (
		_w16083_,
		_w16090_,
		_w16091_
	);
	LUT2 #(
		.INIT('h2)
	) name12045 (
		_w16083_,
		_w16090_,
		_w16092_
	);
	LUT2 #(
		.INIT('h1)
	) name12046 (
		_w14798_,
		_w16092_,
		_w16093_
	);
	LUT2 #(
		.INIT('h1)
	) name12047 (
		_w16091_,
		_w16093_,
		_w16094_
	);
	LUT2 #(
		.INIT('h1)
	) name12048 (
		_w16015_,
		_w16016_,
		_w16095_
	);
	LUT2 #(
		.INIT('h8)
	) name12049 (
		_w16023_,
		_w16095_,
		_w16096_
	);
	LUT2 #(
		.INIT('h1)
	) name12050 (
		_w16023_,
		_w16095_,
		_w16097_
	);
	LUT2 #(
		.INIT('h1)
	) name12051 (
		_w16096_,
		_w16097_,
		_w16098_
	);
	LUT2 #(
		.INIT('h4)
	) name12052 (
		_w16094_,
		_w16098_,
		_w16099_
	);
	LUT2 #(
		.INIT('h1)
	) name12053 (
		_w16079_,
		_w16099_,
		_w16100_
	);
	LUT2 #(
		.INIT('h4)
	) name12054 (
		_w16001_,
		_w16005_,
		_w16101_
	);
	LUT2 #(
		.INIT('h1)
	) name12055 (
		_w16006_,
		_w16101_,
		_w16102_
	);
	LUT2 #(
		.INIT('h2)
	) name12056 (
		_w16010_,
		_w16025_,
		_w16103_
	);
	LUT2 #(
		.INIT('h1)
	) name12057 (
		_w16026_,
		_w16103_,
		_w16104_
	);
	LUT2 #(
		.INIT('h2)
	) name12058 (
		_w16102_,
		_w16104_,
		_w16105_
	);
	LUT2 #(
		.INIT('h4)
	) name12059 (
		_w16102_,
		_w16104_,
		_w16106_
	);
	LUT2 #(
		.INIT('h1)
	) name12060 (
		_w16105_,
		_w16106_,
		_w16107_
	);
	LUT2 #(
		.INIT('h1)
	) name12061 (
		_w16100_,
		_w16107_,
		_w16108_
	);
	LUT2 #(
		.INIT('h8)
	) name12062 (
		_w16100_,
		_w16107_,
		_w16109_
	);
	LUT2 #(
		.INIT('h1)
	) name12063 (
		_w16108_,
		_w16109_,
		_w16110_
	);
	LUT2 #(
		.INIT('h2)
	) name12064 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14791_,
		_w16111_
	);
	LUT2 #(
		.INIT('h1)
	) name12065 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14787_,
		_w16112_
	);
	LUT2 #(
		.INIT('h1)
	) name12066 (
		_w16111_,
		_w16112_,
		_w16113_
	);
	LUT2 #(
		.INIT('h1)
	) name12067 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14761_,
		_w16114_
	);
	LUT2 #(
		.INIT('h2)
	) name12068 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14765_,
		_w16115_
	);
	LUT2 #(
		.INIT('h4)
	) name12069 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14772_,
		_w16116_
	);
	LUT2 #(
		.INIT('h8)
	) name12070 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14776_,
		_w16117_
	);
	LUT2 #(
		.INIT('h1)
	) name12071 (
		_w16116_,
		_w16117_,
		_w16118_
	);
	LUT2 #(
		.INIT('h4)
	) name12072 (
		_w16114_,
		_w16118_,
		_w16119_
	);
	LUT2 #(
		.INIT('h4)
	) name12073 (
		_w16115_,
		_w16119_,
		_w16120_
	);
	LUT2 #(
		.INIT('h1)
	) name12074 (
		_w16113_,
		_w16120_,
		_w16121_
	);
	LUT2 #(
		.INIT('h8)
	) name12075 (
		_w16066_,
		_w16073_,
		_w16122_
	);
	LUT2 #(
		.INIT('h1)
	) name12076 (
		_w16074_,
		_w16122_,
		_w16123_
	);
	LUT2 #(
		.INIT('h1)
	) name12077 (
		_w16121_,
		_w16123_,
		_w16124_
	);
	LUT2 #(
		.INIT('h4)
	) name12078 (
		_w10878_,
		_w14993_,
		_w16125_
	);
	LUT2 #(
		.INIT('h4)
	) name12079 (
		_w9869_,
		_w15044_,
		_w16126_
	);
	LUT2 #(
		.INIT('h1)
	) name12080 (
		_w16125_,
		_w16126_,
		_w16127_
	);
	LUT2 #(
		.INIT('h1)
	) name12081 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16127_,
		_w16128_
	);
	LUT2 #(
		.INIT('h4)
	) name12082 (
		_w14787_,
		_w16128_,
		_w16129_
	);
	LUT2 #(
		.INIT('h2)
	) name12083 (
		_w14787_,
		_w16128_,
		_w16130_
	);
	LUT2 #(
		.INIT('h1)
	) name12084 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14838_,
		_w16131_
	);
	LUT2 #(
		.INIT('h2)
	) name12085 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14842_,
		_w16132_
	);
	LUT2 #(
		.INIT('h4)
	) name12086 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14846_,
		_w16133_
	);
	LUT2 #(
		.INIT('h8)
	) name12087 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14849_,
		_w16134_
	);
	LUT2 #(
		.INIT('h1)
	) name12088 (
		_w16133_,
		_w16134_,
		_w16135_
	);
	LUT2 #(
		.INIT('h4)
	) name12089 (
		_w16131_,
		_w16135_,
		_w16136_
	);
	LUT2 #(
		.INIT('h4)
	) name12090 (
		_w16132_,
		_w16136_,
		_w16137_
	);
	LUT2 #(
		.INIT('h1)
	) name12091 (
		_w16130_,
		_w16137_,
		_w16138_
	);
	LUT2 #(
		.INIT('h1)
	) name12092 (
		_w16129_,
		_w16138_,
		_w16139_
	);
	LUT2 #(
		.INIT('h1)
	) name12093 (
		_w16091_,
		_w16092_,
		_w16140_
	);
	LUT2 #(
		.INIT('h2)
	) name12094 (
		_w14798_,
		_w16140_,
		_w16141_
	);
	LUT2 #(
		.INIT('h4)
	) name12095 (
		_w14798_,
		_w16140_,
		_w16142_
	);
	LUT2 #(
		.INIT('h1)
	) name12096 (
		_w16141_,
		_w16142_,
		_w16143_
	);
	LUT2 #(
		.INIT('h8)
	) name12097 (
		_w16139_,
		_w16143_,
		_w16144_
	);
	LUT2 #(
		.INIT('h1)
	) name12098 (
		_w16124_,
		_w16144_,
		_w16145_
	);
	LUT2 #(
		.INIT('h8)
	) name12099 (
		_w16074_,
		_w16078_,
		_w16146_
	);
	LUT2 #(
		.INIT('h1)
	) name12100 (
		_w16079_,
		_w16146_,
		_w16147_
	);
	LUT2 #(
		.INIT('h2)
	) name12101 (
		_w16094_,
		_w16098_,
		_w16148_
	);
	LUT2 #(
		.INIT('h1)
	) name12102 (
		_w16099_,
		_w16148_,
		_w16149_
	);
	LUT2 #(
		.INIT('h8)
	) name12103 (
		_w16147_,
		_w16149_,
		_w16150_
	);
	LUT2 #(
		.INIT('h1)
	) name12104 (
		_w16147_,
		_w16149_,
		_w16151_
	);
	LUT2 #(
		.INIT('h1)
	) name12105 (
		_w16150_,
		_w16151_,
		_w16152_
	);
	LUT2 #(
		.INIT('h4)
	) name12106 (
		_w16145_,
		_w16152_,
		_w16153_
	);
	LUT2 #(
		.INIT('h1)
	) name12107 (
		_w16146_,
		_w16148_,
		_w16154_
	);
	LUT2 #(
		.INIT('h4)
	) name12108 (
		_w16152_,
		_w16154_,
		_w16155_
	);
	LUT2 #(
		.INIT('h1)
	) name12109 (
		_w16153_,
		_w16155_,
		_w16156_
	);
	LUT2 #(
		.INIT('h4)
	) name12110 (
		_w16110_,
		_w16156_,
		_w16157_
	);
	LUT2 #(
		.INIT('h2)
	) name12111 (
		_w16110_,
		_w16156_,
		_w16158_
	);
	LUT2 #(
		.INIT('h1)
	) name12112 (
		_w16157_,
		_w16158_,
		_w16159_
	);
	LUT2 #(
		.INIT('h2)
	) name12113 (
		_w16145_,
		_w16152_,
		_w16160_
	);
	LUT2 #(
		.INIT('h1)
	) name12114 (
		_w16153_,
		_w16160_,
		_w16161_
	);
	LUT2 #(
		.INIT('h4)
	) name12115 (
		_w9869_,
		_w14993_,
		_w16162_
	);
	LUT2 #(
		.INIT('h4)
	) name12116 (
		_w7909_,
		_w15044_,
		_w16163_
	);
	LUT2 #(
		.INIT('h1)
	) name12117 (
		_w16162_,
		_w16163_,
		_w16164_
	);
	LUT2 #(
		.INIT('h1)
	) name12118 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16164_,
		_w16165_
	);
	LUT2 #(
		.INIT('h2)
	) name12119 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14842_,
		_w16166_
	);
	LUT2 #(
		.INIT('h1)
	) name12120 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14838_,
		_w16167_
	);
	LUT2 #(
		.INIT('h8)
	) name12121 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14849_,
		_w16168_
	);
	LUT2 #(
		.INIT('h4)
	) name12122 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14846_,
		_w16169_
	);
	LUT2 #(
		.INIT('h1)
	) name12123 (
		_w16168_,
		_w16169_,
		_w16170_
	);
	LUT2 #(
		.INIT('h4)
	) name12124 (
		_w16166_,
		_w16170_,
		_w16171_
	);
	LUT2 #(
		.INIT('h4)
	) name12125 (
		_w16167_,
		_w16171_,
		_w16172_
	);
	LUT2 #(
		.INIT('h4)
	) name12126 (
		_w16165_,
		_w16172_,
		_w16173_
	);
	LUT2 #(
		.INIT('h2)
	) name12127 (
		_w16165_,
		_w16172_,
		_w16174_
	);
	LUT2 #(
		.INIT('h1)
	) name12128 (
		_w14772_,
		_w16174_,
		_w16175_
	);
	LUT2 #(
		.INIT('h1)
	) name12129 (
		_w16173_,
		_w16175_,
		_w16176_
	);
	LUT2 #(
		.INIT('h1)
	) name12130 (
		_w16129_,
		_w16130_,
		_w16177_
	);
	LUT2 #(
		.INIT('h4)
	) name12131 (
		_w16137_,
		_w16177_,
		_w16178_
	);
	LUT2 #(
		.INIT('h2)
	) name12132 (
		_w16137_,
		_w16177_,
		_w16179_
	);
	LUT2 #(
		.INIT('h1)
	) name12133 (
		_w16178_,
		_w16179_,
		_w16180_
	);
	LUT2 #(
		.INIT('h1)
	) name12134 (
		_w16176_,
		_w16180_,
		_w16181_
	);
	LUT2 #(
		.INIT('h8)
	) name12135 (
		_w16113_,
		_w16120_,
		_w16182_
	);
	LUT2 #(
		.INIT('h1)
	) name12136 (
		_w16121_,
		_w16182_,
		_w16183_
	);
	LUT2 #(
		.INIT('h4)
	) name12137 (
		_w16181_,
		_w16183_,
		_w16184_
	);
	LUT2 #(
		.INIT('h1)
	) name12138 (
		_w16139_,
		_w16143_,
		_w16185_
	);
	LUT2 #(
		.INIT('h1)
	) name12139 (
		_w16144_,
		_w16185_,
		_w16186_
	);
	LUT2 #(
		.INIT('h8)
	) name12140 (
		_w16121_,
		_w16123_,
		_w16187_
	);
	LUT2 #(
		.INIT('h1)
	) name12141 (
		_w16124_,
		_w16187_,
		_w16188_
	);
	LUT2 #(
		.INIT('h8)
	) name12142 (
		_w16186_,
		_w16188_,
		_w16189_
	);
	LUT2 #(
		.INIT('h1)
	) name12143 (
		_w16186_,
		_w16188_,
		_w16190_
	);
	LUT2 #(
		.INIT('h1)
	) name12144 (
		_w16189_,
		_w16190_,
		_w16191_
	);
	LUT2 #(
		.INIT('h4)
	) name12145 (
		_w16184_,
		_w16191_,
		_w16192_
	);
	LUT2 #(
		.INIT('h1)
	) name12146 (
		_w16185_,
		_w16187_,
		_w16193_
	);
	LUT2 #(
		.INIT('h4)
	) name12147 (
		_w16191_,
		_w16193_,
		_w16194_
	);
	LUT2 #(
		.INIT('h1)
	) name12148 (
		_w16192_,
		_w16194_,
		_w16195_
	);
	LUT2 #(
		.INIT('h4)
	) name12149 (
		_w16161_,
		_w16195_,
		_w16196_
	);
	LUT2 #(
		.INIT('h2)
	) name12150 (
		_w16161_,
		_w16195_,
		_w16197_
	);
	LUT2 #(
		.INIT('h4)
	) name12151 (
		_w7909_,
		_w14993_,
		_w16198_
	);
	LUT2 #(
		.INIT('h2)
	) name12152 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w8554_,
		_w16199_
	);
	LUT2 #(
		.INIT('h8)
	) name12153 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16199_,
		_w16200_
	);
	LUT2 #(
		.INIT('h1)
	) name12154 (
		_w16198_,
		_w16200_,
		_w16201_
	);
	LUT2 #(
		.INIT('h1)
	) name12155 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16201_,
		_w16202_
	);
	LUT2 #(
		.INIT('h1)
	) name12156 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14838_,
		_w16203_
	);
	LUT2 #(
		.INIT('h2)
	) name12157 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14842_,
		_w16204_
	);
	LUT2 #(
		.INIT('h4)
	) name12158 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14846_,
		_w16205_
	);
	LUT2 #(
		.INIT('h8)
	) name12159 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14849_,
		_w16206_
	);
	LUT2 #(
		.INIT('h1)
	) name12160 (
		_w16205_,
		_w16206_,
		_w16207_
	);
	LUT2 #(
		.INIT('h4)
	) name12161 (
		_w16203_,
		_w16207_,
		_w16208_
	);
	LUT2 #(
		.INIT('h4)
	) name12162 (
		_w16204_,
		_w16208_,
		_w16209_
	);
	LUT2 #(
		.INIT('h4)
	) name12163 (
		_w16202_,
		_w16209_,
		_w16210_
	);
	LUT2 #(
		.INIT('h2)
	) name12164 (
		_w16202_,
		_w16209_,
		_w16211_
	);
	LUT2 #(
		.INIT('h2)
	) name12165 (
		_w14761_,
		_w16211_,
		_w16212_
	);
	LUT2 #(
		.INIT('h1)
	) name12166 (
		_w16210_,
		_w16212_,
		_w16213_
	);
	LUT2 #(
		.INIT('h1)
	) name12167 (
		_w16173_,
		_w16174_,
		_w16214_
	);
	LUT2 #(
		.INIT('h2)
	) name12168 (
		_w14772_,
		_w16214_,
		_w16215_
	);
	LUT2 #(
		.INIT('h4)
	) name12169 (
		_w14772_,
		_w16214_,
		_w16216_
	);
	LUT2 #(
		.INIT('h1)
	) name12170 (
		_w16215_,
		_w16216_,
		_w16217_
	);
	LUT2 #(
		.INIT('h4)
	) name12171 (
		_w16213_,
		_w16217_,
		_w16218_
	);
	LUT2 #(
		.INIT('h1)
	) name12172 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14761_,
		_w16219_
	);
	LUT2 #(
		.INIT('h2)
	) name12173 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14765_,
		_w16220_
	);
	LUT2 #(
		.INIT('h4)
	) name12174 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14772_,
		_w16221_
	);
	LUT2 #(
		.INIT('h8)
	) name12175 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14776_,
		_w16222_
	);
	LUT2 #(
		.INIT('h1)
	) name12176 (
		_w16221_,
		_w16222_,
		_w16223_
	);
	LUT2 #(
		.INIT('h4)
	) name12177 (
		_w16219_,
		_w16223_,
		_w16224_
	);
	LUT2 #(
		.INIT('h4)
	) name12178 (
		_w16220_,
		_w16224_,
		_w16225_
	);
	LUT2 #(
		.INIT('h1)
	) name12179 (
		_w16218_,
		_w16225_,
		_w16226_
	);
	LUT2 #(
		.INIT('h8)
	) name12180 (
		_w16176_,
		_w16180_,
		_w16227_
	);
	LUT2 #(
		.INIT('h1)
	) name12181 (
		_w16181_,
		_w16227_,
		_w16228_
	);
	LUT2 #(
		.INIT('h8)
	) name12182 (
		_w16183_,
		_w16228_,
		_w16229_
	);
	LUT2 #(
		.INIT('h1)
	) name12183 (
		_w16183_,
		_w16228_,
		_w16230_
	);
	LUT2 #(
		.INIT('h1)
	) name12184 (
		_w16229_,
		_w16230_,
		_w16231_
	);
	LUT2 #(
		.INIT('h4)
	) name12185 (
		_w16226_,
		_w16231_,
		_w16232_
	);
	LUT2 #(
		.INIT('h1)
	) name12186 (
		_w16227_,
		_w16231_,
		_w16233_
	);
	LUT2 #(
		.INIT('h1)
	) name12187 (
		_w16232_,
		_w16233_,
		_w16234_
	);
	LUT2 #(
		.INIT('h2)
	) name12188 (
		_w16184_,
		_w16191_,
		_w16235_
	);
	LUT2 #(
		.INIT('h1)
	) name12189 (
		_w16192_,
		_w16235_,
		_w16236_
	);
	LUT2 #(
		.INIT('h2)
	) name12190 (
		_w16234_,
		_w16236_,
		_w16237_
	);
	LUT2 #(
		.INIT('h4)
	) name12191 (
		_w16234_,
		_w16236_,
		_w16238_
	);
	LUT2 #(
		.INIT('h1)
	) name12192 (
		_w16237_,
		_w16238_,
		_w16239_
	);
	LUT2 #(
		.INIT('h2)
	) name12193 (
		_w16226_,
		_w16231_,
		_w16240_
	);
	LUT2 #(
		.INIT('h1)
	) name12194 (
		_w16232_,
		_w16240_,
		_w16241_
	);
	LUT2 #(
		.INIT('h4)
	) name12195 (
		_w9225_,
		_w15044_,
		_w16242_
	);
	LUT2 #(
		.INIT('h4)
	) name12196 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16199_,
		_w16243_
	);
	LUT2 #(
		.INIT('h1)
	) name12197 (
		_w16242_,
		_w16243_,
		_w16244_
	);
	LUT2 #(
		.INIT('h1)
	) name12198 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16244_,
		_w16245_
	);
	LUT2 #(
		.INIT('h1)
	) name12199 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14838_,
		_w16246_
	);
	LUT2 #(
		.INIT('h2)
	) name12200 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14842_,
		_w16247_
	);
	LUT2 #(
		.INIT('h4)
	) name12201 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14846_,
		_w16248_
	);
	LUT2 #(
		.INIT('h8)
	) name12202 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14849_,
		_w16249_
	);
	LUT2 #(
		.INIT('h1)
	) name12203 (
		_w16248_,
		_w16249_,
		_w16250_
	);
	LUT2 #(
		.INIT('h4)
	) name12204 (
		_w16246_,
		_w16250_,
		_w16251_
	);
	LUT2 #(
		.INIT('h4)
	) name12205 (
		_w16247_,
		_w16251_,
		_w16252_
	);
	LUT2 #(
		.INIT('h2)
	) name12206 (
		_w16245_,
		_w16252_,
		_w16253_
	);
	LUT2 #(
		.INIT('h4)
	) name12207 (
		_w16245_,
		_w16252_,
		_w16254_
	);
	LUT2 #(
		.INIT('h2)
	) name12208 (
		_w14846_,
		_w16254_,
		_w16255_
	);
	LUT2 #(
		.INIT('h1)
	) name12209 (
		_w16253_,
		_w16255_,
		_w16256_
	);
	LUT2 #(
		.INIT('h1)
	) name12210 (
		_w16210_,
		_w16211_,
		_w16257_
	);
	LUT2 #(
		.INIT('h8)
	) name12211 (
		_w14761_,
		_w16257_,
		_w16258_
	);
	LUT2 #(
		.INIT('h1)
	) name12212 (
		_w14761_,
		_w16257_,
		_w16259_
	);
	LUT2 #(
		.INIT('h1)
	) name12213 (
		_w16258_,
		_w16259_,
		_w16260_
	);
	LUT2 #(
		.INIT('h8)
	) name12214 (
		_w16256_,
		_w16260_,
		_w16261_
	);
	LUT2 #(
		.INIT('h2)
	) name12215 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14765_,
		_w16262_
	);
	LUT2 #(
		.INIT('h1)
	) name12216 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14761_,
		_w16263_
	);
	LUT2 #(
		.INIT('h1)
	) name12217 (
		_w16262_,
		_w16263_,
		_w16264_
	);
	LUT2 #(
		.INIT('h1)
	) name12218 (
		_w16261_,
		_w16264_,
		_w16265_
	);
	LUT2 #(
		.INIT('h2)
	) name12219 (
		_w16213_,
		_w16217_,
		_w16266_
	);
	LUT2 #(
		.INIT('h1)
	) name12220 (
		_w16218_,
		_w16266_,
		_w16267_
	);
	LUT2 #(
		.INIT('h2)
	) name12221 (
		_w16225_,
		_w16267_,
		_w16268_
	);
	LUT2 #(
		.INIT('h4)
	) name12222 (
		_w16225_,
		_w16267_,
		_w16269_
	);
	LUT2 #(
		.INIT('h1)
	) name12223 (
		_w16268_,
		_w16269_,
		_w16270_
	);
	LUT2 #(
		.INIT('h4)
	) name12224 (
		_w16265_,
		_w16270_,
		_w16271_
	);
	LUT2 #(
		.INIT('h1)
	) name12225 (
		_w16266_,
		_w16270_,
		_w16272_
	);
	LUT2 #(
		.INIT('h1)
	) name12226 (
		_w16271_,
		_w16272_,
		_w16273_
	);
	LUT2 #(
		.INIT('h4)
	) name12227 (
		_w16241_,
		_w16273_,
		_w16274_
	);
	LUT2 #(
		.INIT('h2)
	) name12228 (
		_w16241_,
		_w16273_,
		_w16275_
	);
	LUT2 #(
		.INIT('h1)
	) name12229 (
		_w16274_,
		_w16275_,
		_w16276_
	);
	LUT2 #(
		.INIT('h1)
	) name12230 (
		_w16253_,
		_w16254_,
		_w16277_
	);
	LUT2 #(
		.INIT('h8)
	) name12231 (
		_w14846_,
		_w16277_,
		_w16278_
	);
	LUT2 #(
		.INIT('h1)
	) name12232 (
		_w14846_,
		_w16277_,
		_w16279_
	);
	LUT2 #(
		.INIT('h1)
	) name12233 (
		_w16278_,
		_w16279_,
		_w16280_
	);
	LUT2 #(
		.INIT('h8)
	) name12234 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14842_,
		_w16281_
	);
	LUT2 #(
		.INIT('h1)
	) name12235 (
		_w14838_,
		_w16281_,
		_w16282_
	);
	LUT2 #(
		.INIT('h4)
	) name12236 (
		_w7469_,
		_w15044_,
		_w16283_
	);
	LUT2 #(
		.INIT('h4)
	) name12237 (
		_w9225_,
		_w14993_,
		_w16284_
	);
	LUT2 #(
		.INIT('h1)
	) name12238 (
		_w16283_,
		_w16284_,
		_w16285_
	);
	LUT2 #(
		.INIT('h1)
	) name12239 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16285_,
		_w16286_
	);
	LUT2 #(
		.INIT('h2)
	) name12240 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14842_,
		_w16287_
	);
	LUT2 #(
		.INIT('h2)
	) name12241 (
		_w14838_,
		_w16287_,
		_w16288_
	);
	LUT2 #(
		.INIT('h2)
	) name12242 (
		_w16286_,
		_w16288_,
		_w16289_
	);
	LUT2 #(
		.INIT('h1)
	) name12243 (
		_w16282_,
		_w16289_,
		_w16290_
	);
	LUT2 #(
		.INIT('h2)
	) name12244 (
		_w16280_,
		_w16290_,
		_w16291_
	);
	LUT2 #(
		.INIT('h1)
	) name12245 (
		_w16256_,
		_w16260_,
		_w16292_
	);
	LUT2 #(
		.INIT('h1)
	) name12246 (
		_w16261_,
		_w16292_,
		_w16293_
	);
	LUT2 #(
		.INIT('h4)
	) name12247 (
		_w16264_,
		_w16293_,
		_w16294_
	);
	LUT2 #(
		.INIT('h2)
	) name12248 (
		_w16264_,
		_w16293_,
		_w16295_
	);
	LUT2 #(
		.INIT('h1)
	) name12249 (
		_w16294_,
		_w16295_,
		_w16296_
	);
	LUT2 #(
		.INIT('h8)
	) name12250 (
		_w16291_,
		_w16296_,
		_w16297_
	);
	LUT2 #(
		.INIT('h8)
	) name12251 (
		_w16264_,
		_w16292_,
		_w16298_
	);
	LUT2 #(
		.INIT('h2)
	) name12252 (
		_w16265_,
		_w16270_,
		_w16299_
	);
	LUT2 #(
		.INIT('h1)
	) name12253 (
		_w16271_,
		_w16298_,
		_w16300_
	);
	LUT2 #(
		.INIT('h4)
	) name12254 (
		_w16299_,
		_w16300_,
		_w16301_
	);
	LUT2 #(
		.INIT('h2)
	) name12255 (
		_w16297_,
		_w16301_,
		_w16302_
	);
	LUT2 #(
		.INIT('h8)
	) name12256 (
		_w16270_,
		_w16298_,
		_w16303_
	);
	LUT2 #(
		.INIT('h1)
	) name12257 (
		_w16302_,
		_w16303_,
		_w16304_
	);
	LUT2 #(
		.INIT('h2)
	) name12258 (
		_w16276_,
		_w16304_,
		_w16305_
	);
	LUT2 #(
		.INIT('h1)
	) name12259 (
		_w16274_,
		_w16305_,
		_w16306_
	);
	LUT2 #(
		.INIT('h2)
	) name12260 (
		_w16239_,
		_w16306_,
		_w16307_
	);
	LUT2 #(
		.INIT('h1)
	) name12261 (
		_w16237_,
		_w16307_,
		_w16308_
	);
	LUT2 #(
		.INIT('h1)
	) name12262 (
		_w16197_,
		_w16308_,
		_w16309_
	);
	LUT2 #(
		.INIT('h1)
	) name12263 (
		_w16196_,
		_w16309_,
		_w16310_
	);
	LUT2 #(
		.INIT('h2)
	) name12264 (
		_w16159_,
		_w16310_,
		_w16311_
	);
	LUT2 #(
		.INIT('h1)
	) name12265 (
		_w16157_,
		_w16311_,
		_w16312_
	);
	LUT2 #(
		.INIT('h2)
	) name12266 (
		_w16027_,
		_w16034_,
		_w16313_
	);
	LUT2 #(
		.INIT('h1)
	) name12267 (
		_w16035_,
		_w16313_,
		_w16314_
	);
	LUT2 #(
		.INIT('h1)
	) name12268 (
		_w16101_,
		_w16103_,
		_w16315_
	);
	LUT2 #(
		.INIT('h8)
	) name12269 (
		_w16107_,
		_w16315_,
		_w16316_
	);
	LUT2 #(
		.INIT('h1)
	) name12270 (
		_w16108_,
		_w16316_,
		_w16317_
	);
	LUT2 #(
		.INIT('h2)
	) name12271 (
		_w16314_,
		_w16317_,
		_w16318_
	);
	LUT2 #(
		.INIT('h4)
	) name12272 (
		_w16314_,
		_w16317_,
		_w16319_
	);
	LUT2 #(
		.INIT('h1)
	) name12273 (
		_w16318_,
		_w16319_,
		_w16320_
	);
	LUT2 #(
		.INIT('h2)
	) name12274 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14865_,
		_w16321_
	);
	LUT2 #(
		.INIT('h1)
	) name12275 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14861_,
		_w16322_
	);
	LUT2 #(
		.INIT('h1)
	) name12276 (
		_w16321_,
		_w16322_,
		_w16323_
	);
	LUT2 #(
		.INIT('h4)
	) name12277 (
		_w16320_,
		_w16323_,
		_w16324_
	);
	LUT2 #(
		.INIT('h2)
	) name12278 (
		_w16320_,
		_w16323_,
		_w16325_
	);
	LUT2 #(
		.INIT('h1)
	) name12279 (
		_w16324_,
		_w16325_,
		_w16326_
	);
	LUT2 #(
		.INIT('h4)
	) name12280 (
		_w16312_,
		_w16326_,
		_w16327_
	);
	LUT2 #(
		.INIT('h1)
	) name12281 (
		_w16318_,
		_w16323_,
		_w16328_
	);
	LUT2 #(
		.INIT('h4)
	) name12282 (
		_w15980_,
		_w16038_,
		_w16329_
	);
	LUT2 #(
		.INIT('h1)
	) name12283 (
		_w16039_,
		_w16329_,
		_w16330_
	);
	LUT2 #(
		.INIT('h2)
	) name12284 (
		_w16046_,
		_w16330_,
		_w16331_
	);
	LUT2 #(
		.INIT('h4)
	) name12285 (
		_w16046_,
		_w16330_,
		_w16332_
	);
	LUT2 #(
		.INIT('h1)
	) name12286 (
		_w16331_,
		_w16332_,
		_w16333_
	);
	LUT2 #(
		.INIT('h4)
	) name12287 (
		_w16328_,
		_w16333_,
		_w16334_
	);
	LUT2 #(
		.INIT('h1)
	) name12288 (
		_w16329_,
		_w16333_,
		_w16335_
	);
	LUT2 #(
		.INIT('h1)
	) name12289 (
		_w16334_,
		_w16335_,
		_w16336_
	);
	LUT2 #(
		.INIT('h2)
	) name12290 (
		_w16047_,
		_w16052_,
		_w16337_
	);
	LUT2 #(
		.INIT('h1)
	) name12291 (
		_w16053_,
		_w16337_,
		_w16338_
	);
	LUT2 #(
		.INIT('h4)
	) name12292 (
		_w16336_,
		_w16338_,
		_w16339_
	);
	LUT2 #(
		.INIT('h8)
	) name12293 (
		_w16319_,
		_w16323_,
		_w16340_
	);
	LUT2 #(
		.INIT('h2)
	) name12294 (
		_w16328_,
		_w16333_,
		_w16341_
	);
	LUT2 #(
		.INIT('h1)
	) name12295 (
		_w16334_,
		_w16340_,
		_w16342_
	);
	LUT2 #(
		.INIT('h4)
	) name12296 (
		_w16341_,
		_w16342_,
		_w16343_
	);
	LUT2 #(
		.INIT('h1)
	) name12297 (
		_w16339_,
		_w16343_,
		_w16344_
	);
	LUT2 #(
		.INIT('h8)
	) name12298 (
		_w16327_,
		_w16344_,
		_w16345_
	);
	LUT2 #(
		.INIT('h2)
	) name12299 (
		_w16336_,
		_w16338_,
		_w16346_
	);
	LUT2 #(
		.INIT('h8)
	) name12300 (
		_w16333_,
		_w16340_,
		_w16347_
	);
	LUT2 #(
		.INIT('h4)
	) name12301 (
		_w16339_,
		_w16347_,
		_w16348_
	);
	LUT2 #(
		.INIT('h1)
	) name12302 (
		_w16346_,
		_w16348_,
		_w16349_
	);
	LUT2 #(
		.INIT('h4)
	) name12303 (
		_w16345_,
		_w16349_,
		_w16350_
	);
	LUT2 #(
		.INIT('h8)
	) name12304 (
		_w15899_,
		_w16059_,
		_w16351_
	);
	LUT2 #(
		.INIT('h4)
	) name12305 (
		_w16350_,
		_w16351_,
		_w16352_
	);
	LUT2 #(
		.INIT('h4)
	) name12306 (
		_w15695_,
		_w15774_,
		_w16353_
	);
	LUT2 #(
		.INIT('h4)
	) name12307 (
		_w15898_,
		_w16353_,
		_w16354_
	);
	LUT2 #(
		.INIT('h2)
	) name12308 (
		_w15975_,
		_w15977_,
		_w16355_
	);
	LUT2 #(
		.INIT('h2)
	) name12309 (
		_w16055_,
		_w16057_,
		_w16356_
	);
	LUT2 #(
		.INIT('h4)
	) name12310 (
		_w15978_,
		_w16356_,
		_w16357_
	);
	LUT2 #(
		.INIT('h1)
	) name12311 (
		_w16355_,
		_w16357_,
		_w16358_
	);
	LUT2 #(
		.INIT('h2)
	) name12312 (
		_w15899_,
		_w16358_,
		_w16359_
	);
	LUT2 #(
		.INIT('h4)
	) name12313 (
		_w15894_,
		_w15897_,
		_w16360_
	);
	LUT2 #(
		.INIT('h1)
	) name12314 (
		_w16354_,
		_w16360_,
		_w16361_
	);
	LUT2 #(
		.INIT('h4)
	) name12315 (
		_w16359_,
		_w16361_,
		_w16362_
	);
	LUT2 #(
		.INIT('h4)
	) name12316 (
		_w16352_,
		_w16362_,
		_w16363_
	);
	LUT2 #(
		.INIT('h1)
	) name12317 (
		_w14779_,
		_w14805_,
		_w16364_
	);
	LUT2 #(
		.INIT('h1)
	) name12318 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14814_,
		_w16365_
	);
	LUT2 #(
		.INIT('h2)
	) name12319 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14818_,
		_w16366_
	);
	LUT2 #(
		.INIT('h4)
	) name12320 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14825_,
		_w16367_
	);
	LUT2 #(
		.INIT('h8)
	) name12321 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14829_,
		_w16368_
	);
	LUT2 #(
		.INIT('h1)
	) name12322 (
		_w16367_,
		_w16368_,
		_w16369_
	);
	LUT2 #(
		.INIT('h4)
	) name12323 (
		_w16365_,
		_w16369_,
		_w16370_
	);
	LUT2 #(
		.INIT('h4)
	) name12324 (
		_w16366_,
		_w16370_,
		_w16371_
	);
	LUT2 #(
		.INIT('h1)
	) name12325 (
		_w14806_,
		_w16371_,
		_w16372_
	);
	LUT2 #(
		.INIT('h1)
	) name12326 (
		_w16364_,
		_w16372_,
		_w16373_
	);
	LUT2 #(
		.INIT('h1)
	) name12327 (
		_w14806_,
		_w16364_,
		_w16374_
	);
	LUT2 #(
		.INIT('h4)
	) name12328 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14825_,
		_w16375_
	);
	LUT2 #(
		.INIT('h8)
	) name12329 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14829_,
		_w16376_
	);
	LUT2 #(
		.INIT('h1)
	) name12330 (
		_w16375_,
		_w16376_,
		_w16377_
	);
	LUT2 #(
		.INIT('h8)
	) name12331 (
		_w14820_,
		_w16377_,
		_w16378_
	);
	LUT2 #(
		.INIT('h2)
	) name12332 (
		_w16374_,
		_w16378_,
		_w16379_
	);
	LUT2 #(
		.INIT('h4)
	) name12333 (
		_w16374_,
		_w16378_,
		_w16380_
	);
	LUT2 #(
		.INIT('h1)
	) name12334 (
		_w16379_,
		_w16380_,
		_w16381_
	);
	LUT2 #(
		.INIT('h2)
	) name12335 (
		_w16373_,
		_w16381_,
		_w16382_
	);
	LUT2 #(
		.INIT('h1)
	) name12336 (
		_w14852_,
		_w16382_,
		_w16383_
	);
	LUT2 #(
		.INIT('h1)
	) name12337 (
		_w14806_,
		_w16378_,
		_w16384_
	);
	LUT2 #(
		.INIT('h1)
	) name12338 (
		_w16364_,
		_w16384_,
		_w16385_
	);
	LUT2 #(
		.INIT('h4)
	) name12339 (
		_w14832_,
		_w16374_,
		_w16386_
	);
	LUT2 #(
		.INIT('h2)
	) name12340 (
		_w14832_,
		_w16374_,
		_w16387_
	);
	LUT2 #(
		.INIT('h1)
	) name12341 (
		_w16386_,
		_w16387_,
		_w16388_
	);
	LUT2 #(
		.INIT('h4)
	) name12342 (
		_w16385_,
		_w16388_,
		_w16389_
	);
	LUT2 #(
		.INIT('h2)
	) name12343 (
		_w16385_,
		_w16388_,
		_w16390_
	);
	LUT2 #(
		.INIT('h1)
	) name12344 (
		_w16389_,
		_w16390_,
		_w16391_
	);
	LUT2 #(
		.INIT('h4)
	) name12345 (
		_w14852_,
		_w16391_,
		_w16392_
	);
	LUT2 #(
		.INIT('h2)
	) name12346 (
		_w14852_,
		_w16391_,
		_w16393_
	);
	LUT2 #(
		.INIT('h1)
	) name12347 (
		_w16392_,
		_w16393_,
		_w16394_
	);
	LUT2 #(
		.INIT('h4)
	) name12348 (
		_w16383_,
		_w16394_,
		_w16395_
	);
	LUT2 #(
		.INIT('h4)
	) name12349 (
		_w16382_,
		_w16392_,
		_w16396_
	);
	LUT2 #(
		.INIT('h1)
	) name12350 (
		_w16395_,
		_w16396_,
		_w16397_
	);
	LUT2 #(
		.INIT('h4)
	) name12351 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14798_,
		_w16398_
	);
	LUT2 #(
		.INIT('h8)
	) name12352 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14802_,
		_w16399_
	);
	LUT2 #(
		.INIT('h1)
	) name12353 (
		_w16398_,
		_w16399_,
		_w16400_
	);
	LUT2 #(
		.INIT('h8)
	) name12354 (
		_w14793_,
		_w16400_,
		_w16401_
	);
	LUT2 #(
		.INIT('h8)
	) name12355 (
		_w14779_,
		_w16401_,
		_w16402_
	);
	LUT2 #(
		.INIT('h1)
	) name12356 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14814_,
		_w16403_
	);
	LUT2 #(
		.INIT('h2)
	) name12357 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14818_,
		_w16404_
	);
	LUT2 #(
		.INIT('h4)
	) name12358 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14825_,
		_w16405_
	);
	LUT2 #(
		.INIT('h8)
	) name12359 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14829_,
		_w16406_
	);
	LUT2 #(
		.INIT('h1)
	) name12360 (
		_w16405_,
		_w16406_,
		_w16407_
	);
	LUT2 #(
		.INIT('h4)
	) name12361 (
		_w16403_,
		_w16407_,
		_w16408_
	);
	LUT2 #(
		.INIT('h4)
	) name12362 (
		_w16404_,
		_w16408_,
		_w16409_
	);
	LUT2 #(
		.INIT('h1)
	) name12363 (
		_w16402_,
		_w16409_,
		_w16410_
	);
	LUT2 #(
		.INIT('h1)
	) name12364 (
		_w14779_,
		_w16401_,
		_w16411_
	);
	LUT2 #(
		.INIT('h1)
	) name12365 (
		_w16410_,
		_w16411_,
		_w16412_
	);
	LUT2 #(
		.INIT('h4)
	) name12366 (
		_w16371_,
		_w16374_,
		_w16413_
	);
	LUT2 #(
		.INIT('h2)
	) name12367 (
		_w16371_,
		_w16374_,
		_w16414_
	);
	LUT2 #(
		.INIT('h1)
	) name12368 (
		_w16413_,
		_w16414_,
		_w16415_
	);
	LUT2 #(
		.INIT('h2)
	) name12369 (
		_w16412_,
		_w16415_,
		_w16416_
	);
	LUT2 #(
		.INIT('h1)
	) name12370 (
		_w14852_,
		_w16416_,
		_w16417_
	);
	LUT2 #(
		.INIT('h4)
	) name12371 (
		_w16373_,
		_w16381_,
		_w16418_
	);
	LUT2 #(
		.INIT('h1)
	) name12372 (
		_w16382_,
		_w16418_,
		_w16419_
	);
	LUT2 #(
		.INIT('h2)
	) name12373 (
		_w14852_,
		_w16419_,
		_w16420_
	);
	LUT2 #(
		.INIT('h2)
	) name12374 (
		_w16383_,
		_w16418_,
		_w16421_
	);
	LUT2 #(
		.INIT('h1)
	) name12375 (
		_w16420_,
		_w16421_,
		_w16422_
	);
	LUT2 #(
		.INIT('h4)
	) name12376 (
		_w16417_,
		_w16422_,
		_w16423_
	);
	LUT2 #(
		.INIT('h1)
	) name12377 (
		_w16418_,
		_w16422_,
		_w16424_
	);
	LUT2 #(
		.INIT('h1)
	) name12378 (
		_w16423_,
		_w16424_,
		_w16425_
	);
	LUT2 #(
		.INIT('h2)
	) name12379 (
		_w16397_,
		_w16425_,
		_w16426_
	);
	LUT2 #(
		.INIT('h2)
	) name12380 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14865_,
		_w16427_
	);
	LUT2 #(
		.INIT('h1)
	) name12381 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14861_,
		_w16428_
	);
	LUT2 #(
		.INIT('h4)
	) name12382 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14872_,
		_w16429_
	);
	LUT2 #(
		.INIT('h8)
	) name12383 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14876_,
		_w16430_
	);
	LUT2 #(
		.INIT('h1)
	) name12384 (
		_w16429_,
		_w16430_,
		_w16431_
	);
	LUT2 #(
		.INIT('h4)
	) name12385 (
		_w16427_,
		_w16431_,
		_w16432_
	);
	LUT2 #(
		.INIT('h4)
	) name12386 (
		_w16428_,
		_w16432_,
		_w16433_
	);
	LUT2 #(
		.INIT('h1)
	) name12387 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14887_,
		_w16434_
	);
	LUT2 #(
		.INIT('h2)
	) name12388 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14891_,
		_w16435_
	);
	LUT2 #(
		.INIT('h4)
	) name12389 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14898_,
		_w16436_
	);
	LUT2 #(
		.INIT('h8)
	) name12390 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14902_,
		_w16437_
	);
	LUT2 #(
		.INIT('h1)
	) name12391 (
		_w16436_,
		_w16437_,
		_w16438_
	);
	LUT2 #(
		.INIT('h4)
	) name12392 (
		_w16434_,
		_w16438_,
		_w16439_
	);
	LUT2 #(
		.INIT('h4)
	) name12393 (
		_w16435_,
		_w16439_,
		_w16440_
	);
	LUT2 #(
		.INIT('h8)
	) name12394 (
		_w16433_,
		_w16440_,
		_w16441_
	);
	LUT2 #(
		.INIT('h1)
	) name12395 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14914_,
		_w16442_
	);
	LUT2 #(
		.INIT('h2)
	) name12396 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14918_,
		_w16443_
	);
	LUT2 #(
		.INIT('h4)
	) name12397 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14925_,
		_w16444_
	);
	LUT2 #(
		.INIT('h8)
	) name12398 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14929_,
		_w16445_
	);
	LUT2 #(
		.INIT('h1)
	) name12399 (
		_w16444_,
		_w16445_,
		_w16446_
	);
	LUT2 #(
		.INIT('h4)
	) name12400 (
		_w16442_,
		_w16446_,
		_w16447_
	);
	LUT2 #(
		.INIT('h4)
	) name12401 (
		_w16443_,
		_w16447_,
		_w16448_
	);
	LUT2 #(
		.INIT('h1)
	) name12402 (
		_w16441_,
		_w16448_,
		_w16449_
	);
	LUT2 #(
		.INIT('h1)
	) name12403 (
		_w16433_,
		_w16440_,
		_w16450_
	);
	LUT2 #(
		.INIT('h1)
	) name12404 (
		_w16449_,
		_w16450_,
		_w16451_
	);
	LUT2 #(
		.INIT('h1)
	) name12405 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14861_,
		_w16452_
	);
	LUT2 #(
		.INIT('h2)
	) name12406 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14865_,
		_w16453_
	);
	LUT2 #(
		.INIT('h4)
	) name12407 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14872_,
		_w16454_
	);
	LUT2 #(
		.INIT('h8)
	) name12408 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14876_,
		_w16455_
	);
	LUT2 #(
		.INIT('h1)
	) name12409 (
		_w16454_,
		_w16455_,
		_w16456_
	);
	LUT2 #(
		.INIT('h4)
	) name12410 (
		_w16452_,
		_w16456_,
		_w16457_
	);
	LUT2 #(
		.INIT('h4)
	) name12411 (
		_w16453_,
		_w16457_,
		_w16458_
	);
	LUT2 #(
		.INIT('h1)
	) name12412 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14887_,
		_w16459_
	);
	LUT2 #(
		.INIT('h2)
	) name12413 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14891_,
		_w16460_
	);
	LUT2 #(
		.INIT('h4)
	) name12414 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14898_,
		_w16461_
	);
	LUT2 #(
		.INIT('h8)
	) name12415 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14902_,
		_w16462_
	);
	LUT2 #(
		.INIT('h1)
	) name12416 (
		_w16461_,
		_w16462_,
		_w16463_
	);
	LUT2 #(
		.INIT('h4)
	) name12417 (
		_w16459_,
		_w16463_,
		_w16464_
	);
	LUT2 #(
		.INIT('h4)
	) name12418 (
		_w16460_,
		_w16464_,
		_w16465_
	);
	LUT2 #(
		.INIT('h8)
	) name12419 (
		_w16458_,
		_w16465_,
		_w16466_
	);
	LUT2 #(
		.INIT('h1)
	) name12420 (
		_w16458_,
		_w16465_,
		_w16467_
	);
	LUT2 #(
		.INIT('h1)
	) name12421 (
		_w16466_,
		_w16467_,
		_w16468_
	);
	LUT2 #(
		.INIT('h1)
	) name12422 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14914_,
		_w16469_
	);
	LUT2 #(
		.INIT('h2)
	) name12423 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14918_,
		_w16470_
	);
	LUT2 #(
		.INIT('h4)
	) name12424 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14925_,
		_w16471_
	);
	LUT2 #(
		.INIT('h8)
	) name12425 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14929_,
		_w16472_
	);
	LUT2 #(
		.INIT('h1)
	) name12426 (
		_w16471_,
		_w16472_,
		_w16473_
	);
	LUT2 #(
		.INIT('h4)
	) name12427 (
		_w16469_,
		_w16473_,
		_w16474_
	);
	LUT2 #(
		.INIT('h4)
	) name12428 (
		_w16470_,
		_w16474_,
		_w16475_
	);
	LUT2 #(
		.INIT('h4)
	) name12429 (
		_w16468_,
		_w16475_,
		_w16476_
	);
	LUT2 #(
		.INIT('h2)
	) name12430 (
		_w16468_,
		_w16475_,
		_w16477_
	);
	LUT2 #(
		.INIT('h1)
	) name12431 (
		_w16476_,
		_w16477_,
		_w16478_
	);
	LUT2 #(
		.INIT('h2)
	) name12432 (
		_w16451_,
		_w16478_,
		_w16479_
	);
	LUT2 #(
		.INIT('h1)
	) name12433 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14967_,
		_w16480_
	);
	LUT2 #(
		.INIT('h2)
	) name12434 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14969_,
		_w16481_
	);
	LUT2 #(
		.INIT('h1)
	) name12435 (
		_w16480_,
		_w16481_,
		_w16482_
	);
	LUT2 #(
		.INIT('h1)
	) name12436 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14947_,
		_w16483_
	);
	LUT2 #(
		.INIT('h2)
	) name12437 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14951_,
		_w16484_
	);
	LUT2 #(
		.INIT('h4)
	) name12438 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14958_,
		_w16485_
	);
	LUT2 #(
		.INIT('h8)
	) name12439 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14962_,
		_w16486_
	);
	LUT2 #(
		.INIT('h1)
	) name12440 (
		_w16485_,
		_w16486_,
		_w16487_
	);
	LUT2 #(
		.INIT('h4)
	) name12441 (
		_w16483_,
		_w16487_,
		_w16488_
	);
	LUT2 #(
		.INIT('h4)
	) name12442 (
		_w16484_,
		_w16488_,
		_w16489_
	);
	LUT2 #(
		.INIT('h4)
	) name12443 (
		_w16482_,
		_w16489_,
		_w16490_
	);
	LUT2 #(
		.INIT('h2)
	) name12444 (
		_w16482_,
		_w16489_,
		_w16491_
	);
	LUT2 #(
		.INIT('h1)
	) name12445 (
		_w16490_,
		_w16491_,
		_w16492_
	);
	LUT2 #(
		.INIT('h2)
	) name12446 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w11448_,
		_w16493_
	);
	LUT2 #(
		.INIT('h2)
	) name12447 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16493_,
		_w16494_
	);
	LUT2 #(
		.INIT('h2)
	) name12448 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w11196_,
		_w16495_
	);
	LUT2 #(
		.INIT('h1)
	) name12449 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16495_,
		_w16496_
	);
	LUT2 #(
		.INIT('h1)
	) name12450 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16494_,
		_w16497_
	);
	LUT2 #(
		.INIT('h4)
	) name12451 (
		_w16496_,
		_w16497_,
		_w16498_
	);
	LUT2 #(
		.INIT('h4)
	) name12452 (
		_w16492_,
		_w16498_,
		_w16499_
	);
	LUT2 #(
		.INIT('h2)
	) name12453 (
		_w16492_,
		_w16498_,
		_w16500_
	);
	LUT2 #(
		.INIT('h1)
	) name12454 (
		_w16499_,
		_w16500_,
		_w16501_
	);
	LUT2 #(
		.INIT('h1)
	) name12455 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14967_,
		_w16502_
	);
	LUT2 #(
		.INIT('h2)
	) name12456 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14969_,
		_w16503_
	);
	LUT2 #(
		.INIT('h1)
	) name12457 (
		_w16502_,
		_w16503_,
		_w16504_
	);
	LUT2 #(
		.INIT('h1)
	) name12458 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14947_,
		_w16505_
	);
	LUT2 #(
		.INIT('h2)
	) name12459 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14951_,
		_w16506_
	);
	LUT2 #(
		.INIT('h4)
	) name12460 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14958_,
		_w16507_
	);
	LUT2 #(
		.INIT('h8)
	) name12461 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14962_,
		_w16508_
	);
	LUT2 #(
		.INIT('h1)
	) name12462 (
		_w16507_,
		_w16508_,
		_w16509_
	);
	LUT2 #(
		.INIT('h4)
	) name12463 (
		_w16505_,
		_w16509_,
		_w16510_
	);
	LUT2 #(
		.INIT('h4)
	) name12464 (
		_w16506_,
		_w16510_,
		_w16511_
	);
	LUT2 #(
		.INIT('h4)
	) name12465 (
		_w16504_,
		_w16511_,
		_w16512_
	);
	LUT2 #(
		.INIT('h2)
	) name12466 (
		_w16504_,
		_w16511_,
		_w16513_
	);
	LUT2 #(
		.INIT('h2)
	) name12467 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w10858_,
		_w16514_
	);
	LUT2 #(
		.INIT('h2)
	) name12468 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16514_,
		_w16515_
	);
	LUT2 #(
		.INIT('h1)
	) name12469 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16493_,
		_w16516_
	);
	LUT2 #(
		.INIT('h1)
	) name12470 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16515_,
		_w16517_
	);
	LUT2 #(
		.INIT('h4)
	) name12471 (
		_w16516_,
		_w16517_,
		_w16518_
	);
	LUT2 #(
		.INIT('h1)
	) name12472 (
		_w16513_,
		_w16518_,
		_w16519_
	);
	LUT2 #(
		.INIT('h1)
	) name12473 (
		_w16512_,
		_w16519_,
		_w16520_
	);
	LUT2 #(
		.INIT('h2)
	) name12474 (
		_w16501_,
		_w16520_,
		_w16521_
	);
	LUT2 #(
		.INIT('h1)
	) name12475 (
		_w16479_,
		_w16521_,
		_w16522_
	);
	LUT2 #(
		.INIT('h4)
	) name12476 (
		_w16490_,
		_w16498_,
		_w16523_
	);
	LUT2 #(
		.INIT('h1)
	) name12477 (
		_w16491_,
		_w16523_,
		_w16524_
	);
	LUT2 #(
		.INIT('h2)
	) name12478 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16495_,
		_w16525_
	);
	LUT2 #(
		.INIT('h2)
	) name12479 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w10538_,
		_w16526_
	);
	LUT2 #(
		.INIT('h1)
	) name12480 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16526_,
		_w16527_
	);
	LUT2 #(
		.INIT('h1)
	) name12481 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16525_,
		_w16528_
	);
	LUT2 #(
		.INIT('h4)
	) name12482 (
		_w16527_,
		_w16528_,
		_w16529_
	);
	LUT2 #(
		.INIT('h1)
	) name12483 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14947_,
		_w16530_
	);
	LUT2 #(
		.INIT('h2)
	) name12484 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14951_,
		_w16531_
	);
	LUT2 #(
		.INIT('h4)
	) name12485 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14958_,
		_w16532_
	);
	LUT2 #(
		.INIT('h8)
	) name12486 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14962_,
		_w16533_
	);
	LUT2 #(
		.INIT('h1)
	) name12487 (
		_w16532_,
		_w16533_,
		_w16534_
	);
	LUT2 #(
		.INIT('h4)
	) name12488 (
		_w16530_,
		_w16534_,
		_w16535_
	);
	LUT2 #(
		.INIT('h4)
	) name12489 (
		_w16531_,
		_w16535_,
		_w16536_
	);
	LUT2 #(
		.INIT('h2)
	) name12490 (
		_w16529_,
		_w16536_,
		_w16537_
	);
	LUT2 #(
		.INIT('h4)
	) name12491 (
		_w16529_,
		_w16536_,
		_w16538_
	);
	LUT2 #(
		.INIT('h1)
	) name12492 (
		_w16537_,
		_w16538_,
		_w16539_
	);
	LUT2 #(
		.INIT('h4)
	) name12493 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14967_,
		_w16540_
	);
	LUT2 #(
		.INIT('h8)
	) name12494 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14969_,
		_w16541_
	);
	LUT2 #(
		.INIT('h1)
	) name12495 (
		_w16540_,
		_w16541_,
		_w16542_
	);
	LUT2 #(
		.INIT('h8)
	) name12496 (
		_w16539_,
		_w16542_,
		_w16543_
	);
	LUT2 #(
		.INIT('h1)
	) name12497 (
		_w16539_,
		_w16542_,
		_w16544_
	);
	LUT2 #(
		.INIT('h1)
	) name12498 (
		_w16543_,
		_w16544_,
		_w16545_
	);
	LUT2 #(
		.INIT('h8)
	) name12499 (
		_w16524_,
		_w16545_,
		_w16546_
	);
	LUT2 #(
		.INIT('h1)
	) name12500 (
		_w16524_,
		_w16545_,
		_w16547_
	);
	LUT2 #(
		.INIT('h1)
	) name12501 (
		_w16546_,
		_w16547_,
		_w16548_
	);
	LUT2 #(
		.INIT('h1)
	) name12502 (
		_w16466_,
		_w16475_,
		_w16549_
	);
	LUT2 #(
		.INIT('h1)
	) name12503 (
		_w16467_,
		_w16549_,
		_w16550_
	);
	LUT2 #(
		.INIT('h1)
	) name12504 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14887_,
		_w16551_
	);
	LUT2 #(
		.INIT('h2)
	) name12505 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14891_,
		_w16552_
	);
	LUT2 #(
		.INIT('h4)
	) name12506 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14898_,
		_w16553_
	);
	LUT2 #(
		.INIT('h8)
	) name12507 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14902_,
		_w16554_
	);
	LUT2 #(
		.INIT('h1)
	) name12508 (
		_w16553_,
		_w16554_,
		_w16555_
	);
	LUT2 #(
		.INIT('h4)
	) name12509 (
		_w16551_,
		_w16555_,
		_w16556_
	);
	LUT2 #(
		.INIT('h4)
	) name12510 (
		_w16552_,
		_w16556_,
		_w16557_
	);
	LUT2 #(
		.INIT('h1)
	) name12511 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14861_,
		_w16558_
	);
	LUT2 #(
		.INIT('h2)
	) name12512 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14865_,
		_w16559_
	);
	LUT2 #(
		.INIT('h4)
	) name12513 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14872_,
		_w16560_
	);
	LUT2 #(
		.INIT('h8)
	) name12514 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14876_,
		_w16561_
	);
	LUT2 #(
		.INIT('h1)
	) name12515 (
		_w16560_,
		_w16561_,
		_w16562_
	);
	LUT2 #(
		.INIT('h4)
	) name12516 (
		_w16558_,
		_w16562_,
		_w16563_
	);
	LUT2 #(
		.INIT('h4)
	) name12517 (
		_w16559_,
		_w16563_,
		_w16564_
	);
	LUT2 #(
		.INIT('h8)
	) name12518 (
		_w16557_,
		_w16564_,
		_w16565_
	);
	LUT2 #(
		.INIT('h1)
	) name12519 (
		_w16557_,
		_w16564_,
		_w16566_
	);
	LUT2 #(
		.INIT('h1)
	) name12520 (
		_w16565_,
		_w16566_,
		_w16567_
	);
	LUT2 #(
		.INIT('h1)
	) name12521 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14914_,
		_w16568_
	);
	LUT2 #(
		.INIT('h2)
	) name12522 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14918_,
		_w16569_
	);
	LUT2 #(
		.INIT('h4)
	) name12523 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14925_,
		_w16570_
	);
	LUT2 #(
		.INIT('h8)
	) name12524 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14929_,
		_w16571_
	);
	LUT2 #(
		.INIT('h1)
	) name12525 (
		_w16570_,
		_w16571_,
		_w16572_
	);
	LUT2 #(
		.INIT('h4)
	) name12526 (
		_w16568_,
		_w16572_,
		_w16573_
	);
	LUT2 #(
		.INIT('h4)
	) name12527 (
		_w16569_,
		_w16573_,
		_w16574_
	);
	LUT2 #(
		.INIT('h4)
	) name12528 (
		_w16567_,
		_w16574_,
		_w16575_
	);
	LUT2 #(
		.INIT('h2)
	) name12529 (
		_w16567_,
		_w16574_,
		_w16576_
	);
	LUT2 #(
		.INIT('h1)
	) name12530 (
		_w16575_,
		_w16576_,
		_w16577_
	);
	LUT2 #(
		.INIT('h2)
	) name12531 (
		_w16550_,
		_w16577_,
		_w16578_
	);
	LUT2 #(
		.INIT('h4)
	) name12532 (
		_w16550_,
		_w16577_,
		_w16579_
	);
	LUT2 #(
		.INIT('h1)
	) name12533 (
		_w16578_,
		_w16579_,
		_w16580_
	);
	LUT2 #(
		.INIT('h2)
	) name12534 (
		_w16548_,
		_w16580_,
		_w16581_
	);
	LUT2 #(
		.INIT('h4)
	) name12535 (
		_w16548_,
		_w16580_,
		_w16582_
	);
	LUT2 #(
		.INIT('h1)
	) name12536 (
		_w16581_,
		_w16582_,
		_w16583_
	);
	LUT2 #(
		.INIT('h1)
	) name12537 (
		_w16522_,
		_w16583_,
		_w16584_
	);
	LUT2 #(
		.INIT('h8)
	) name12538 (
		_w16522_,
		_w16583_,
		_w16585_
	);
	LUT2 #(
		.INIT('h1)
	) name12539 (
		_w16584_,
		_w16585_,
		_w16586_
	);
	LUT2 #(
		.INIT('h1)
	) name12540 (
		_w16512_,
		_w16513_,
		_w16587_
	);
	LUT2 #(
		.INIT('h2)
	) name12541 (
		_w16518_,
		_w16587_,
		_w16588_
	);
	LUT2 #(
		.INIT('h4)
	) name12542 (
		_w16518_,
		_w16587_,
		_w16589_
	);
	LUT2 #(
		.INIT('h1)
	) name12543 (
		_w16588_,
		_w16589_,
		_w16590_
	);
	LUT2 #(
		.INIT('h2)
	) name12544 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w9845_,
		_w16591_
	);
	LUT2 #(
		.INIT('h2)
	) name12545 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16591_,
		_w16592_
	);
	LUT2 #(
		.INIT('h1)
	) name12546 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16514_,
		_w16593_
	);
	LUT2 #(
		.INIT('h1)
	) name12547 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16592_,
		_w16594_
	);
	LUT2 #(
		.INIT('h4)
	) name12548 (
		_w16593_,
		_w16594_,
		_w16595_
	);
	LUT2 #(
		.INIT('h1)
	) name12549 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14947_,
		_w16596_
	);
	LUT2 #(
		.INIT('h2)
	) name12550 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14951_,
		_w16597_
	);
	LUT2 #(
		.INIT('h4)
	) name12551 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14958_,
		_w16598_
	);
	LUT2 #(
		.INIT('h8)
	) name12552 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14962_,
		_w16599_
	);
	LUT2 #(
		.INIT('h1)
	) name12553 (
		_w16598_,
		_w16599_,
		_w16600_
	);
	LUT2 #(
		.INIT('h4)
	) name12554 (
		_w16596_,
		_w16600_,
		_w16601_
	);
	LUT2 #(
		.INIT('h4)
	) name12555 (
		_w16597_,
		_w16601_,
		_w16602_
	);
	LUT2 #(
		.INIT('h2)
	) name12556 (
		_w16595_,
		_w16602_,
		_w16603_
	);
	LUT2 #(
		.INIT('h4)
	) name12557 (
		_w16595_,
		_w16602_,
		_w16604_
	);
	LUT2 #(
		.INIT('h4)
	) name12558 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14967_,
		_w16605_
	);
	LUT2 #(
		.INIT('h8)
	) name12559 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14969_,
		_w16606_
	);
	LUT2 #(
		.INIT('h1)
	) name12560 (
		_w16605_,
		_w16606_,
		_w16607_
	);
	LUT2 #(
		.INIT('h1)
	) name12561 (
		_w16604_,
		_w16607_,
		_w16608_
	);
	LUT2 #(
		.INIT('h1)
	) name12562 (
		_w16603_,
		_w16608_,
		_w16609_
	);
	LUT2 #(
		.INIT('h8)
	) name12563 (
		_w16590_,
		_w16609_,
		_w16610_
	);
	LUT2 #(
		.INIT('h1)
	) name12564 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14887_,
		_w16611_
	);
	LUT2 #(
		.INIT('h2)
	) name12565 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14891_,
		_w16612_
	);
	LUT2 #(
		.INIT('h4)
	) name12566 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14898_,
		_w16613_
	);
	LUT2 #(
		.INIT('h8)
	) name12567 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14902_,
		_w16614_
	);
	LUT2 #(
		.INIT('h1)
	) name12568 (
		_w16613_,
		_w16614_,
		_w16615_
	);
	LUT2 #(
		.INIT('h4)
	) name12569 (
		_w16611_,
		_w16615_,
		_w16616_
	);
	LUT2 #(
		.INIT('h4)
	) name12570 (
		_w16612_,
		_w16616_,
		_w16617_
	);
	LUT2 #(
		.INIT('h1)
	) name12571 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14861_,
		_w16618_
	);
	LUT2 #(
		.INIT('h2)
	) name12572 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14865_,
		_w16619_
	);
	LUT2 #(
		.INIT('h4)
	) name12573 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14872_,
		_w16620_
	);
	LUT2 #(
		.INIT('h8)
	) name12574 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14876_,
		_w16621_
	);
	LUT2 #(
		.INIT('h1)
	) name12575 (
		_w16620_,
		_w16621_,
		_w16622_
	);
	LUT2 #(
		.INIT('h4)
	) name12576 (
		_w16618_,
		_w16622_,
		_w16623_
	);
	LUT2 #(
		.INIT('h4)
	) name12577 (
		_w16619_,
		_w16623_,
		_w16624_
	);
	LUT2 #(
		.INIT('h8)
	) name12578 (
		_w16617_,
		_w16624_,
		_w16625_
	);
	LUT2 #(
		.INIT('h1)
	) name12579 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14914_,
		_w16626_
	);
	LUT2 #(
		.INIT('h2)
	) name12580 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14918_,
		_w16627_
	);
	LUT2 #(
		.INIT('h4)
	) name12581 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14925_,
		_w16628_
	);
	LUT2 #(
		.INIT('h8)
	) name12582 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14929_,
		_w16629_
	);
	LUT2 #(
		.INIT('h1)
	) name12583 (
		_w16628_,
		_w16629_,
		_w16630_
	);
	LUT2 #(
		.INIT('h4)
	) name12584 (
		_w16626_,
		_w16630_,
		_w16631_
	);
	LUT2 #(
		.INIT('h4)
	) name12585 (
		_w16627_,
		_w16631_,
		_w16632_
	);
	LUT2 #(
		.INIT('h1)
	) name12586 (
		_w16625_,
		_w16632_,
		_w16633_
	);
	LUT2 #(
		.INIT('h1)
	) name12587 (
		_w16617_,
		_w16624_,
		_w16634_
	);
	LUT2 #(
		.INIT('h1)
	) name12588 (
		_w16633_,
		_w16634_,
		_w16635_
	);
	LUT2 #(
		.INIT('h1)
	) name12589 (
		_w16441_,
		_w16450_,
		_w16636_
	);
	LUT2 #(
		.INIT('h2)
	) name12590 (
		_w16448_,
		_w16636_,
		_w16637_
	);
	LUT2 #(
		.INIT('h4)
	) name12591 (
		_w16448_,
		_w16636_,
		_w16638_
	);
	LUT2 #(
		.INIT('h1)
	) name12592 (
		_w16637_,
		_w16638_,
		_w16639_
	);
	LUT2 #(
		.INIT('h2)
	) name12593 (
		_w16635_,
		_w16639_,
		_w16640_
	);
	LUT2 #(
		.INIT('h1)
	) name12594 (
		_w16610_,
		_w16640_,
		_w16641_
	);
	LUT2 #(
		.INIT('h4)
	) name12595 (
		_w16451_,
		_w16478_,
		_w16642_
	);
	LUT2 #(
		.INIT('h1)
	) name12596 (
		_w16479_,
		_w16642_,
		_w16643_
	);
	LUT2 #(
		.INIT('h4)
	) name12597 (
		_w16501_,
		_w16520_,
		_w16644_
	);
	LUT2 #(
		.INIT('h1)
	) name12598 (
		_w16521_,
		_w16644_,
		_w16645_
	);
	LUT2 #(
		.INIT('h8)
	) name12599 (
		_w16643_,
		_w16645_,
		_w16646_
	);
	LUT2 #(
		.INIT('h1)
	) name12600 (
		_w16643_,
		_w16645_,
		_w16647_
	);
	LUT2 #(
		.INIT('h1)
	) name12601 (
		_w16646_,
		_w16647_,
		_w16648_
	);
	LUT2 #(
		.INIT('h4)
	) name12602 (
		_w16641_,
		_w16648_,
		_w16649_
	);
	LUT2 #(
		.INIT('h1)
	) name12603 (
		_w16642_,
		_w16644_,
		_w16650_
	);
	LUT2 #(
		.INIT('h4)
	) name12604 (
		_w16648_,
		_w16650_,
		_w16651_
	);
	LUT2 #(
		.INIT('h1)
	) name12605 (
		_w16649_,
		_w16651_,
		_w16652_
	);
	LUT2 #(
		.INIT('h2)
	) name12606 (
		_w16586_,
		_w16652_,
		_w16653_
	);
	LUT2 #(
		.INIT('h1)
	) name12607 (
		_w16426_,
		_w16653_,
		_w16654_
	);
	LUT2 #(
		.INIT('h1)
	) name12608 (
		_w16546_,
		_w16578_,
		_w16655_
	);
	LUT2 #(
		.INIT('h1)
	) name12609 (
		_w16565_,
		_w16574_,
		_w16656_
	);
	LUT2 #(
		.INIT('h1)
	) name12610 (
		_w16566_,
		_w16656_,
		_w16657_
	);
	LUT2 #(
		.INIT('h4)
	) name12611 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14872_,
		_w16658_
	);
	LUT2 #(
		.INIT('h8)
	) name12612 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14876_,
		_w16659_
	);
	LUT2 #(
		.INIT('h1)
	) name12613 (
		_w16658_,
		_w16659_,
		_w16660_
	);
	LUT2 #(
		.INIT('h8)
	) name12614 (
		_w14867_,
		_w16660_,
		_w16661_
	);
	LUT2 #(
		.INIT('h1)
	) name12615 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14887_,
		_w16662_
	);
	LUT2 #(
		.INIT('h2)
	) name12616 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14891_,
		_w16663_
	);
	LUT2 #(
		.INIT('h4)
	) name12617 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14898_,
		_w16664_
	);
	LUT2 #(
		.INIT('h8)
	) name12618 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14902_,
		_w16665_
	);
	LUT2 #(
		.INIT('h1)
	) name12619 (
		_w16664_,
		_w16665_,
		_w16666_
	);
	LUT2 #(
		.INIT('h4)
	) name12620 (
		_w16662_,
		_w16666_,
		_w16667_
	);
	LUT2 #(
		.INIT('h4)
	) name12621 (
		_w16663_,
		_w16667_,
		_w16668_
	);
	LUT2 #(
		.INIT('h8)
	) name12622 (
		_w16661_,
		_w16668_,
		_w16669_
	);
	LUT2 #(
		.INIT('h1)
	) name12623 (
		_w16661_,
		_w16668_,
		_w16670_
	);
	LUT2 #(
		.INIT('h1)
	) name12624 (
		_w16669_,
		_w16670_,
		_w16671_
	);
	LUT2 #(
		.INIT('h1)
	) name12625 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14914_,
		_w16672_
	);
	LUT2 #(
		.INIT('h2)
	) name12626 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14918_,
		_w16673_
	);
	LUT2 #(
		.INIT('h4)
	) name12627 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14925_,
		_w16674_
	);
	LUT2 #(
		.INIT('h8)
	) name12628 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14929_,
		_w16675_
	);
	LUT2 #(
		.INIT('h1)
	) name12629 (
		_w16674_,
		_w16675_,
		_w16676_
	);
	LUT2 #(
		.INIT('h4)
	) name12630 (
		_w16672_,
		_w16676_,
		_w16677_
	);
	LUT2 #(
		.INIT('h4)
	) name12631 (
		_w16673_,
		_w16677_,
		_w16678_
	);
	LUT2 #(
		.INIT('h4)
	) name12632 (
		_w16671_,
		_w16678_,
		_w16679_
	);
	LUT2 #(
		.INIT('h2)
	) name12633 (
		_w16671_,
		_w16678_,
		_w16680_
	);
	LUT2 #(
		.INIT('h1)
	) name12634 (
		_w16679_,
		_w16680_,
		_w16681_
	);
	LUT2 #(
		.INIT('h4)
	) name12635 (
		_w16657_,
		_w16681_,
		_w16682_
	);
	LUT2 #(
		.INIT('h2)
	) name12636 (
		_w16657_,
		_w16681_,
		_w16683_
	);
	LUT2 #(
		.INIT('h1)
	) name12637 (
		_w16682_,
		_w16683_,
		_w16684_
	);
	LUT2 #(
		.INIT('h1)
	) name12638 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14967_,
		_w16685_
	);
	LUT2 #(
		.INIT('h2)
	) name12639 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14969_,
		_w16686_
	);
	LUT2 #(
		.INIT('h1)
	) name12640 (
		_w16685_,
		_w16686_,
		_w16687_
	);
	LUT2 #(
		.INIT('h1)
	) name12641 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14947_,
		_w16688_
	);
	LUT2 #(
		.INIT('h2)
	) name12642 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14951_,
		_w16689_
	);
	LUT2 #(
		.INIT('h4)
	) name12643 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14958_,
		_w16690_
	);
	LUT2 #(
		.INIT('h8)
	) name12644 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14962_,
		_w16691_
	);
	LUT2 #(
		.INIT('h1)
	) name12645 (
		_w16690_,
		_w16691_,
		_w16692_
	);
	LUT2 #(
		.INIT('h4)
	) name12646 (
		_w16688_,
		_w16692_,
		_w16693_
	);
	LUT2 #(
		.INIT('h4)
	) name12647 (
		_w16689_,
		_w16693_,
		_w16694_
	);
	LUT2 #(
		.INIT('h4)
	) name12648 (
		_w16687_,
		_w16694_,
		_w16695_
	);
	LUT2 #(
		.INIT('h2)
	) name12649 (
		_w16687_,
		_w16694_,
		_w16696_
	);
	LUT2 #(
		.INIT('h1)
	) name12650 (
		_w16695_,
		_w16696_,
		_w16697_
	);
	LUT2 #(
		.INIT('h2)
	) name12651 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16526_,
		_w16698_
	);
	LUT2 #(
		.INIT('h2)
	) name12652 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w10096_,
		_w16699_
	);
	LUT2 #(
		.INIT('h1)
	) name12653 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16699_,
		_w16700_
	);
	LUT2 #(
		.INIT('h1)
	) name12654 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16698_,
		_w16701_
	);
	LUT2 #(
		.INIT('h4)
	) name12655 (
		_w16700_,
		_w16701_,
		_w16702_
	);
	LUT2 #(
		.INIT('h8)
	) name12656 (
		_w16697_,
		_w16702_,
		_w16703_
	);
	LUT2 #(
		.INIT('h1)
	) name12657 (
		_w16697_,
		_w16702_,
		_w16704_
	);
	LUT2 #(
		.INIT('h1)
	) name12658 (
		_w16703_,
		_w16704_,
		_w16705_
	);
	LUT2 #(
		.INIT('h1)
	) name12659 (
		_w16538_,
		_w16542_,
		_w16706_
	);
	LUT2 #(
		.INIT('h1)
	) name12660 (
		_w16537_,
		_w16706_,
		_w16707_
	);
	LUT2 #(
		.INIT('h2)
	) name12661 (
		_w16705_,
		_w16707_,
		_w16708_
	);
	LUT2 #(
		.INIT('h4)
	) name12662 (
		_w16705_,
		_w16707_,
		_w16709_
	);
	LUT2 #(
		.INIT('h1)
	) name12663 (
		_w16708_,
		_w16709_,
		_w16710_
	);
	LUT2 #(
		.INIT('h8)
	) name12664 (
		_w16684_,
		_w16710_,
		_w16711_
	);
	LUT2 #(
		.INIT('h1)
	) name12665 (
		_w16684_,
		_w16710_,
		_w16712_
	);
	LUT2 #(
		.INIT('h1)
	) name12666 (
		_w16711_,
		_w16712_,
		_w16713_
	);
	LUT2 #(
		.INIT('h4)
	) name12667 (
		_w16655_,
		_w16713_,
		_w16714_
	);
	LUT2 #(
		.INIT('h2)
	) name12668 (
		_w16655_,
		_w16713_,
		_w16715_
	);
	LUT2 #(
		.INIT('h1)
	) name12669 (
		_w16714_,
		_w16715_,
		_w16716_
	);
	LUT2 #(
		.INIT('h1)
	) name12670 (
		_w16547_,
		_w16579_,
		_w16717_
	);
	LUT2 #(
		.INIT('h8)
	) name12671 (
		_w16583_,
		_w16717_,
		_w16718_
	);
	LUT2 #(
		.INIT('h1)
	) name12672 (
		_w16584_,
		_w16718_,
		_w16719_
	);
	LUT2 #(
		.INIT('h4)
	) name12673 (
		_w16716_,
		_w16719_,
		_w16720_
	);
	LUT2 #(
		.INIT('h2)
	) name12674 (
		_w16716_,
		_w16719_,
		_w16721_
	);
	LUT2 #(
		.INIT('h1)
	) name12675 (
		_w16720_,
		_w16721_,
		_w16722_
	);
	LUT2 #(
		.INIT('h1)
	) name12676 (
		_w16389_,
		_w16394_,
		_w16723_
	);
	LUT2 #(
		.INIT('h1)
	) name12677 (
		_w16395_,
		_w16723_,
		_w16724_
	);
	LUT2 #(
		.INIT('h4)
	) name12678 (
		_w14832_,
		_w16364_,
		_w16725_
	);
	LUT2 #(
		.INIT('h1)
	) name12679 (
		_w14833_,
		_w16725_,
		_w16726_
	);
	LUT2 #(
		.INIT('h4)
	) name12680 (
		_w14852_,
		_w16390_,
		_w16727_
	);
	LUT2 #(
		.INIT('h2)
	) name12681 (
		_w16726_,
		_w16727_,
		_w16728_
	);
	LUT2 #(
		.INIT('h4)
	) name12682 (
		_w16726_,
		_w16727_,
		_w16729_
	);
	LUT2 #(
		.INIT('h1)
	) name12683 (
		_w16728_,
		_w16729_,
		_w16730_
	);
	LUT2 #(
		.INIT('h2)
	) name12684 (
		_w16724_,
		_w16730_,
		_w16731_
	);
	LUT2 #(
		.INIT('h4)
	) name12685 (
		_w16724_,
		_w16730_,
		_w16732_
	);
	LUT2 #(
		.INIT('h1)
	) name12686 (
		_w16731_,
		_w16732_,
		_w16733_
	);
	LUT2 #(
		.INIT('h8)
	) name12687 (
		_w16722_,
		_w16733_,
		_w16734_
	);
	LUT2 #(
		.INIT('h1)
	) name12688 (
		_w16722_,
		_w16733_,
		_w16735_
	);
	LUT2 #(
		.INIT('h1)
	) name12689 (
		_w16734_,
		_w16735_,
		_w16736_
	);
	LUT2 #(
		.INIT('h4)
	) name12690 (
		_w16654_,
		_w16736_,
		_w16737_
	);
	LUT2 #(
		.INIT('h2)
	) name12691 (
		_w16654_,
		_w16736_,
		_w16738_
	);
	LUT2 #(
		.INIT('h1)
	) name12692 (
		_w16737_,
		_w16738_,
		_w16739_
	);
	LUT2 #(
		.INIT('h8)
	) name12693 (
		_w16417_,
		_w16419_,
		_w16740_
	);
	LUT2 #(
		.INIT('h1)
	) name12694 (
		_w16423_,
		_w16740_,
		_w16741_
	);
	LUT2 #(
		.INIT('h1)
	) name12695 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14787_,
		_w16742_
	);
	LUT2 #(
		.INIT('h2)
	) name12696 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14791_,
		_w16743_
	);
	LUT2 #(
		.INIT('h4)
	) name12697 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14798_,
		_w16744_
	);
	LUT2 #(
		.INIT('h8)
	) name12698 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14802_,
		_w16745_
	);
	LUT2 #(
		.INIT('h1)
	) name12699 (
		_w16744_,
		_w16745_,
		_w16746_
	);
	LUT2 #(
		.INIT('h4)
	) name12700 (
		_w16742_,
		_w16746_,
		_w16747_
	);
	LUT2 #(
		.INIT('h4)
	) name12701 (
		_w16743_,
		_w16747_,
		_w16748_
	);
	LUT2 #(
		.INIT('h8)
	) name12702 (
		_w14779_,
		_w16748_,
		_w16749_
	);
	LUT2 #(
		.INIT('h1)
	) name12703 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14814_,
		_w16750_
	);
	LUT2 #(
		.INIT('h2)
	) name12704 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14818_,
		_w16751_
	);
	LUT2 #(
		.INIT('h4)
	) name12705 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14825_,
		_w16752_
	);
	LUT2 #(
		.INIT('h8)
	) name12706 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14829_,
		_w16753_
	);
	LUT2 #(
		.INIT('h1)
	) name12707 (
		_w16752_,
		_w16753_,
		_w16754_
	);
	LUT2 #(
		.INIT('h4)
	) name12708 (
		_w16750_,
		_w16754_,
		_w16755_
	);
	LUT2 #(
		.INIT('h4)
	) name12709 (
		_w16751_,
		_w16755_,
		_w16756_
	);
	LUT2 #(
		.INIT('h1)
	) name12710 (
		_w16749_,
		_w16756_,
		_w16757_
	);
	LUT2 #(
		.INIT('h1)
	) name12711 (
		_w14779_,
		_w16748_,
		_w16758_
	);
	LUT2 #(
		.INIT('h1)
	) name12712 (
		_w16757_,
		_w16758_,
		_w16759_
	);
	LUT2 #(
		.INIT('h1)
	) name12713 (
		_w16402_,
		_w16411_,
		_w16760_
	);
	LUT2 #(
		.INIT('h2)
	) name12714 (
		_w16409_,
		_w16760_,
		_w16761_
	);
	LUT2 #(
		.INIT('h4)
	) name12715 (
		_w16409_,
		_w16760_,
		_w16762_
	);
	LUT2 #(
		.INIT('h1)
	) name12716 (
		_w16761_,
		_w16762_,
		_w16763_
	);
	LUT2 #(
		.INIT('h2)
	) name12717 (
		_w16759_,
		_w16763_,
		_w16764_
	);
	LUT2 #(
		.INIT('h1)
	) name12718 (
		_w14852_,
		_w16764_,
		_w16765_
	);
	LUT2 #(
		.INIT('h4)
	) name12719 (
		_w16412_,
		_w16415_,
		_w16766_
	);
	LUT2 #(
		.INIT('h1)
	) name12720 (
		_w16416_,
		_w16766_,
		_w16767_
	);
	LUT2 #(
		.INIT('h4)
	) name12721 (
		_w14852_,
		_w16767_,
		_w16768_
	);
	LUT2 #(
		.INIT('h2)
	) name12722 (
		_w14852_,
		_w16767_,
		_w16769_
	);
	LUT2 #(
		.INIT('h1)
	) name12723 (
		_w16768_,
		_w16769_,
		_w16770_
	);
	LUT2 #(
		.INIT('h4)
	) name12724 (
		_w16765_,
		_w16770_,
		_w16771_
	);
	LUT2 #(
		.INIT('h1)
	) name12725 (
		_w16766_,
		_w16770_,
		_w16772_
	);
	LUT2 #(
		.INIT('h1)
	) name12726 (
		_w16771_,
		_w16772_,
		_w16773_
	);
	LUT2 #(
		.INIT('h2)
	) name12727 (
		_w16741_,
		_w16773_,
		_w16774_
	);
	LUT2 #(
		.INIT('h2)
	) name12728 (
		_w16641_,
		_w16648_,
		_w16775_
	);
	LUT2 #(
		.INIT('h1)
	) name12729 (
		_w16649_,
		_w16775_,
		_w16776_
	);
	LUT2 #(
		.INIT('h1)
	) name12730 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14967_,
		_w16777_
	);
	LUT2 #(
		.INIT('h2)
	) name12731 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14969_,
		_w16778_
	);
	LUT2 #(
		.INIT('h1)
	) name12732 (
		_w16777_,
		_w16778_,
		_w16779_
	);
	LUT2 #(
		.INIT('h1)
	) name12733 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14947_,
		_w16780_
	);
	LUT2 #(
		.INIT('h2)
	) name12734 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14951_,
		_w16781_
	);
	LUT2 #(
		.INIT('h4)
	) name12735 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14958_,
		_w16782_
	);
	LUT2 #(
		.INIT('h8)
	) name12736 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14962_,
		_w16783_
	);
	LUT2 #(
		.INIT('h1)
	) name12737 (
		_w16782_,
		_w16783_,
		_w16784_
	);
	LUT2 #(
		.INIT('h4)
	) name12738 (
		_w16780_,
		_w16784_,
		_w16785_
	);
	LUT2 #(
		.INIT('h4)
	) name12739 (
		_w16781_,
		_w16785_,
		_w16786_
	);
	LUT2 #(
		.INIT('h4)
	) name12740 (
		_w16779_,
		_w16786_,
		_w16787_
	);
	LUT2 #(
		.INIT('h2)
	) name12741 (
		_w16779_,
		_w16786_,
		_w16788_
	);
	LUT2 #(
		.INIT('h2)
	) name12742 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w7885_,
		_w16789_
	);
	LUT2 #(
		.INIT('h2)
	) name12743 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16789_,
		_w16790_
	);
	LUT2 #(
		.INIT('h1)
	) name12744 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16591_,
		_w16791_
	);
	LUT2 #(
		.INIT('h1)
	) name12745 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16790_,
		_w16792_
	);
	LUT2 #(
		.INIT('h4)
	) name12746 (
		_w16791_,
		_w16792_,
		_w16793_
	);
	LUT2 #(
		.INIT('h1)
	) name12747 (
		_w16788_,
		_w16793_,
		_w16794_
	);
	LUT2 #(
		.INIT('h1)
	) name12748 (
		_w16787_,
		_w16794_,
		_w16795_
	);
	LUT2 #(
		.INIT('h1)
	) name12749 (
		_w16603_,
		_w16604_,
		_w16796_
	);
	LUT2 #(
		.INIT('h4)
	) name12750 (
		_w16607_,
		_w16796_,
		_w16797_
	);
	LUT2 #(
		.INIT('h2)
	) name12751 (
		_w16607_,
		_w16796_,
		_w16798_
	);
	LUT2 #(
		.INIT('h1)
	) name12752 (
		_w16797_,
		_w16798_,
		_w16799_
	);
	LUT2 #(
		.INIT('h1)
	) name12753 (
		_w16795_,
		_w16799_,
		_w16800_
	);
	LUT2 #(
		.INIT('h1)
	) name12754 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14861_,
		_w16801_
	);
	LUT2 #(
		.INIT('h2)
	) name12755 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14865_,
		_w16802_
	);
	LUT2 #(
		.INIT('h4)
	) name12756 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14872_,
		_w16803_
	);
	LUT2 #(
		.INIT('h8)
	) name12757 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14876_,
		_w16804_
	);
	LUT2 #(
		.INIT('h1)
	) name12758 (
		_w16803_,
		_w16804_,
		_w16805_
	);
	LUT2 #(
		.INIT('h4)
	) name12759 (
		_w16801_,
		_w16805_,
		_w16806_
	);
	LUT2 #(
		.INIT('h4)
	) name12760 (
		_w16802_,
		_w16806_,
		_w16807_
	);
	LUT2 #(
		.INIT('h1)
	) name12761 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14887_,
		_w16808_
	);
	LUT2 #(
		.INIT('h2)
	) name12762 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14891_,
		_w16809_
	);
	LUT2 #(
		.INIT('h4)
	) name12763 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14898_,
		_w16810_
	);
	LUT2 #(
		.INIT('h8)
	) name12764 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14902_,
		_w16811_
	);
	LUT2 #(
		.INIT('h1)
	) name12765 (
		_w16810_,
		_w16811_,
		_w16812_
	);
	LUT2 #(
		.INIT('h4)
	) name12766 (
		_w16808_,
		_w16812_,
		_w16813_
	);
	LUT2 #(
		.INIT('h4)
	) name12767 (
		_w16809_,
		_w16813_,
		_w16814_
	);
	LUT2 #(
		.INIT('h8)
	) name12768 (
		_w16807_,
		_w16814_,
		_w16815_
	);
	LUT2 #(
		.INIT('h1)
	) name12769 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14914_,
		_w16816_
	);
	LUT2 #(
		.INIT('h2)
	) name12770 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14918_,
		_w16817_
	);
	LUT2 #(
		.INIT('h4)
	) name12771 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14925_,
		_w16818_
	);
	LUT2 #(
		.INIT('h8)
	) name12772 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14929_,
		_w16819_
	);
	LUT2 #(
		.INIT('h1)
	) name12773 (
		_w16818_,
		_w16819_,
		_w16820_
	);
	LUT2 #(
		.INIT('h4)
	) name12774 (
		_w16816_,
		_w16820_,
		_w16821_
	);
	LUT2 #(
		.INIT('h4)
	) name12775 (
		_w16817_,
		_w16821_,
		_w16822_
	);
	LUT2 #(
		.INIT('h1)
	) name12776 (
		_w16815_,
		_w16822_,
		_w16823_
	);
	LUT2 #(
		.INIT('h1)
	) name12777 (
		_w16807_,
		_w16814_,
		_w16824_
	);
	LUT2 #(
		.INIT('h1)
	) name12778 (
		_w16823_,
		_w16824_,
		_w16825_
	);
	LUT2 #(
		.INIT('h1)
	) name12779 (
		_w16625_,
		_w16634_,
		_w16826_
	);
	LUT2 #(
		.INIT('h2)
	) name12780 (
		_w16632_,
		_w16826_,
		_w16827_
	);
	LUT2 #(
		.INIT('h4)
	) name12781 (
		_w16632_,
		_w16826_,
		_w16828_
	);
	LUT2 #(
		.INIT('h1)
	) name12782 (
		_w16827_,
		_w16828_,
		_w16829_
	);
	LUT2 #(
		.INIT('h2)
	) name12783 (
		_w16825_,
		_w16829_,
		_w16830_
	);
	LUT2 #(
		.INIT('h1)
	) name12784 (
		_w16800_,
		_w16830_,
		_w16831_
	);
	LUT2 #(
		.INIT('h4)
	) name12785 (
		_w16635_,
		_w16639_,
		_w16832_
	);
	LUT2 #(
		.INIT('h1)
	) name12786 (
		_w16640_,
		_w16832_,
		_w16833_
	);
	LUT2 #(
		.INIT('h1)
	) name12787 (
		_w16590_,
		_w16609_,
		_w16834_
	);
	LUT2 #(
		.INIT('h1)
	) name12788 (
		_w16610_,
		_w16834_,
		_w16835_
	);
	LUT2 #(
		.INIT('h2)
	) name12789 (
		_w16833_,
		_w16835_,
		_w16836_
	);
	LUT2 #(
		.INIT('h4)
	) name12790 (
		_w16833_,
		_w16835_,
		_w16837_
	);
	LUT2 #(
		.INIT('h1)
	) name12791 (
		_w16836_,
		_w16837_,
		_w16838_
	);
	LUT2 #(
		.INIT('h1)
	) name12792 (
		_w16831_,
		_w16838_,
		_w16839_
	);
	LUT2 #(
		.INIT('h1)
	) name12793 (
		_w16832_,
		_w16834_,
		_w16840_
	);
	LUT2 #(
		.INIT('h8)
	) name12794 (
		_w16838_,
		_w16840_,
		_w16841_
	);
	LUT2 #(
		.INIT('h1)
	) name12795 (
		_w16839_,
		_w16841_,
		_w16842_
	);
	LUT2 #(
		.INIT('h2)
	) name12796 (
		_w16776_,
		_w16842_,
		_w16843_
	);
	LUT2 #(
		.INIT('h1)
	) name12797 (
		_w16774_,
		_w16843_,
		_w16844_
	);
	LUT2 #(
		.INIT('h4)
	) name12798 (
		_w16397_,
		_w16425_,
		_w16845_
	);
	LUT2 #(
		.INIT('h1)
	) name12799 (
		_w16426_,
		_w16845_,
		_w16846_
	);
	LUT2 #(
		.INIT('h4)
	) name12800 (
		_w16586_,
		_w16652_,
		_w16847_
	);
	LUT2 #(
		.INIT('h1)
	) name12801 (
		_w16653_,
		_w16847_,
		_w16848_
	);
	LUT2 #(
		.INIT('h8)
	) name12802 (
		_w16846_,
		_w16848_,
		_w16849_
	);
	LUT2 #(
		.INIT('h1)
	) name12803 (
		_w16846_,
		_w16848_,
		_w16850_
	);
	LUT2 #(
		.INIT('h1)
	) name12804 (
		_w16849_,
		_w16850_,
		_w16851_
	);
	LUT2 #(
		.INIT('h8)
	) name12805 (
		_w16844_,
		_w16851_,
		_w16852_
	);
	LUT2 #(
		.INIT('h1)
	) name12806 (
		_w16845_,
		_w16847_,
		_w16853_
	);
	LUT2 #(
		.INIT('h1)
	) name12807 (
		_w16851_,
		_w16853_,
		_w16854_
	);
	LUT2 #(
		.INIT('h1)
	) name12808 (
		_w16852_,
		_w16854_,
		_w16855_
	);
	LUT2 #(
		.INIT('h8)
	) name12809 (
		_w16739_,
		_w16855_,
		_w16856_
	);
	LUT2 #(
		.INIT('h1)
	) name12810 (
		_w16844_,
		_w16851_,
		_w16857_
	);
	LUT2 #(
		.INIT('h1)
	) name12811 (
		_w16852_,
		_w16857_,
		_w16858_
	);
	LUT2 #(
		.INIT('h8)
	) name12812 (
		_w16831_,
		_w16838_,
		_w16859_
	);
	LUT2 #(
		.INIT('h1)
	) name12813 (
		_w16839_,
		_w16859_,
		_w16860_
	);
	LUT2 #(
		.INIT('h1)
	) name12814 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14861_,
		_w16861_
	);
	LUT2 #(
		.INIT('h2)
	) name12815 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14865_,
		_w16862_
	);
	LUT2 #(
		.INIT('h4)
	) name12816 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14872_,
		_w16863_
	);
	LUT2 #(
		.INIT('h8)
	) name12817 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14876_,
		_w16864_
	);
	LUT2 #(
		.INIT('h1)
	) name12818 (
		_w16863_,
		_w16864_,
		_w16865_
	);
	LUT2 #(
		.INIT('h4)
	) name12819 (
		_w16861_,
		_w16865_,
		_w16866_
	);
	LUT2 #(
		.INIT('h4)
	) name12820 (
		_w16862_,
		_w16866_,
		_w16867_
	);
	LUT2 #(
		.INIT('h1)
	) name12821 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14887_,
		_w16868_
	);
	LUT2 #(
		.INIT('h2)
	) name12822 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14891_,
		_w16869_
	);
	LUT2 #(
		.INIT('h4)
	) name12823 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14898_,
		_w16870_
	);
	LUT2 #(
		.INIT('h8)
	) name12824 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14902_,
		_w16871_
	);
	LUT2 #(
		.INIT('h1)
	) name12825 (
		_w16870_,
		_w16871_,
		_w16872_
	);
	LUT2 #(
		.INIT('h4)
	) name12826 (
		_w16868_,
		_w16872_,
		_w16873_
	);
	LUT2 #(
		.INIT('h4)
	) name12827 (
		_w16869_,
		_w16873_,
		_w16874_
	);
	LUT2 #(
		.INIT('h8)
	) name12828 (
		_w16867_,
		_w16874_,
		_w16875_
	);
	LUT2 #(
		.INIT('h1)
	) name12829 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14914_,
		_w16876_
	);
	LUT2 #(
		.INIT('h2)
	) name12830 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14918_,
		_w16877_
	);
	LUT2 #(
		.INIT('h4)
	) name12831 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14925_,
		_w16878_
	);
	LUT2 #(
		.INIT('h8)
	) name12832 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14929_,
		_w16879_
	);
	LUT2 #(
		.INIT('h1)
	) name12833 (
		_w16878_,
		_w16879_,
		_w16880_
	);
	LUT2 #(
		.INIT('h4)
	) name12834 (
		_w16876_,
		_w16880_,
		_w16881_
	);
	LUT2 #(
		.INIT('h4)
	) name12835 (
		_w16877_,
		_w16881_,
		_w16882_
	);
	LUT2 #(
		.INIT('h1)
	) name12836 (
		_w16875_,
		_w16882_,
		_w16883_
	);
	LUT2 #(
		.INIT('h1)
	) name12837 (
		_w16867_,
		_w16874_,
		_w16884_
	);
	LUT2 #(
		.INIT('h1)
	) name12838 (
		_w16883_,
		_w16884_,
		_w16885_
	);
	LUT2 #(
		.INIT('h1)
	) name12839 (
		_w16815_,
		_w16824_,
		_w16886_
	);
	LUT2 #(
		.INIT('h2)
	) name12840 (
		_w16822_,
		_w16886_,
		_w16887_
	);
	LUT2 #(
		.INIT('h4)
	) name12841 (
		_w16822_,
		_w16886_,
		_w16888_
	);
	LUT2 #(
		.INIT('h1)
	) name12842 (
		_w16887_,
		_w16888_,
		_w16889_
	);
	LUT2 #(
		.INIT('h2)
	) name12843 (
		_w16885_,
		_w16889_,
		_w16890_
	);
	LUT2 #(
		.INIT('h1)
	) name12844 (
		_w16787_,
		_w16788_,
		_w16891_
	);
	LUT2 #(
		.INIT('h2)
	) name12845 (
		_w16793_,
		_w16891_,
		_w16892_
	);
	LUT2 #(
		.INIT('h4)
	) name12846 (
		_w16793_,
		_w16891_,
		_w16893_
	);
	LUT2 #(
		.INIT('h1)
	) name12847 (
		_w16892_,
		_w16893_,
		_w16894_
	);
	LUT2 #(
		.INIT('h2)
	) name12848 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w8558_,
		_w16895_
	);
	LUT2 #(
		.INIT('h2)
	) name12849 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16895_,
		_w16896_
	);
	LUT2 #(
		.INIT('h1)
	) name12850 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16789_,
		_w16897_
	);
	LUT2 #(
		.INIT('h1)
	) name12851 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w16896_,
		_w16898_
	);
	LUT2 #(
		.INIT('h4)
	) name12852 (
		_w16897_,
		_w16898_,
		_w16899_
	);
	LUT2 #(
		.INIT('h1)
	) name12853 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14947_,
		_w16900_
	);
	LUT2 #(
		.INIT('h2)
	) name12854 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14951_,
		_w16901_
	);
	LUT2 #(
		.INIT('h4)
	) name12855 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14958_,
		_w16902_
	);
	LUT2 #(
		.INIT('h8)
	) name12856 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14962_,
		_w16903_
	);
	LUT2 #(
		.INIT('h1)
	) name12857 (
		_w16902_,
		_w16903_,
		_w16904_
	);
	LUT2 #(
		.INIT('h4)
	) name12858 (
		_w16900_,
		_w16904_,
		_w16905_
	);
	LUT2 #(
		.INIT('h4)
	) name12859 (
		_w16901_,
		_w16905_,
		_w16906_
	);
	LUT2 #(
		.INIT('h2)
	) name12860 (
		_w16899_,
		_w16906_,
		_w16907_
	);
	LUT2 #(
		.INIT('h4)
	) name12861 (
		_w16899_,
		_w16906_,
		_w16908_
	);
	LUT2 #(
		.INIT('h4)
	) name12862 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14967_,
		_w16909_
	);
	LUT2 #(
		.INIT('h8)
	) name12863 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14969_,
		_w16910_
	);
	LUT2 #(
		.INIT('h1)
	) name12864 (
		_w16909_,
		_w16910_,
		_w16911_
	);
	LUT2 #(
		.INIT('h1)
	) name12865 (
		_w16908_,
		_w16911_,
		_w16912_
	);
	LUT2 #(
		.INIT('h1)
	) name12866 (
		_w16907_,
		_w16912_,
		_w16913_
	);
	LUT2 #(
		.INIT('h8)
	) name12867 (
		_w16894_,
		_w16913_,
		_w16914_
	);
	LUT2 #(
		.INIT('h1)
	) name12868 (
		_w16890_,
		_w16914_,
		_w16915_
	);
	LUT2 #(
		.INIT('h4)
	) name12869 (
		_w16825_,
		_w16829_,
		_w16916_
	);
	LUT2 #(
		.INIT('h1)
	) name12870 (
		_w16830_,
		_w16916_,
		_w16917_
	);
	LUT2 #(
		.INIT('h8)
	) name12871 (
		_w16795_,
		_w16799_,
		_w16918_
	);
	LUT2 #(
		.INIT('h1)
	) name12872 (
		_w16800_,
		_w16918_,
		_w16919_
	);
	LUT2 #(
		.INIT('h2)
	) name12873 (
		_w16917_,
		_w16919_,
		_w16920_
	);
	LUT2 #(
		.INIT('h4)
	) name12874 (
		_w16917_,
		_w16919_,
		_w16921_
	);
	LUT2 #(
		.INIT('h1)
	) name12875 (
		_w16920_,
		_w16921_,
		_w16922_
	);
	LUT2 #(
		.INIT('h2)
	) name12876 (
		_w16915_,
		_w16922_,
		_w16923_
	);
	LUT2 #(
		.INIT('h1)
	) name12877 (
		_w16916_,
		_w16918_,
		_w16924_
	);
	LUT2 #(
		.INIT('h2)
	) name12878 (
		_w16922_,
		_w16924_,
		_w16925_
	);
	LUT2 #(
		.INIT('h1)
	) name12879 (
		_w16923_,
		_w16925_,
		_w16926_
	);
	LUT2 #(
		.INIT('h8)
	) name12880 (
		_w16860_,
		_w16926_,
		_w16927_
	);
	LUT2 #(
		.INIT('h1)
	) name12881 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14814_,
		_w16928_
	);
	LUT2 #(
		.INIT('h2)
	) name12882 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14818_,
		_w16929_
	);
	LUT2 #(
		.INIT('h4)
	) name12883 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14825_,
		_w16930_
	);
	LUT2 #(
		.INIT('h8)
	) name12884 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14829_,
		_w16931_
	);
	LUT2 #(
		.INIT('h1)
	) name12885 (
		_w16930_,
		_w16931_,
		_w16932_
	);
	LUT2 #(
		.INIT('h4)
	) name12886 (
		_w16928_,
		_w16932_,
		_w16933_
	);
	LUT2 #(
		.INIT('h4)
	) name12887 (
		_w16929_,
		_w16933_,
		_w16934_
	);
	LUT2 #(
		.INIT('h1)
	) name12888 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14787_,
		_w16935_
	);
	LUT2 #(
		.INIT('h2)
	) name12889 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14791_,
		_w16936_
	);
	LUT2 #(
		.INIT('h4)
	) name12890 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14798_,
		_w16937_
	);
	LUT2 #(
		.INIT('h8)
	) name12891 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14802_,
		_w16938_
	);
	LUT2 #(
		.INIT('h1)
	) name12892 (
		_w16937_,
		_w16938_,
		_w16939_
	);
	LUT2 #(
		.INIT('h4)
	) name12893 (
		_w16935_,
		_w16939_,
		_w16940_
	);
	LUT2 #(
		.INIT('h4)
	) name12894 (
		_w16936_,
		_w16940_,
		_w16941_
	);
	LUT2 #(
		.INIT('h8)
	) name12895 (
		_w16934_,
		_w16941_,
		_w16942_
	);
	LUT2 #(
		.INIT('h4)
	) name12896 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14772_,
		_w16943_
	);
	LUT2 #(
		.INIT('h8)
	) name12897 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14776_,
		_w16944_
	);
	LUT2 #(
		.INIT('h1)
	) name12898 (
		_w16943_,
		_w16944_,
		_w16945_
	);
	LUT2 #(
		.INIT('h8)
	) name12899 (
		_w14767_,
		_w16945_,
		_w16946_
	);
	LUT2 #(
		.INIT('h1)
	) name12900 (
		_w16942_,
		_w16946_,
		_w16947_
	);
	LUT2 #(
		.INIT('h1)
	) name12901 (
		_w16934_,
		_w16941_,
		_w16948_
	);
	LUT2 #(
		.INIT('h1)
	) name12902 (
		_w16947_,
		_w16948_,
		_w16949_
	);
	LUT2 #(
		.INIT('h1)
	) name12903 (
		_w16749_,
		_w16758_,
		_w16950_
	);
	LUT2 #(
		.INIT('h2)
	) name12904 (
		_w16756_,
		_w16950_,
		_w16951_
	);
	LUT2 #(
		.INIT('h4)
	) name12905 (
		_w16756_,
		_w16950_,
		_w16952_
	);
	LUT2 #(
		.INIT('h1)
	) name12906 (
		_w16951_,
		_w16952_,
		_w16953_
	);
	LUT2 #(
		.INIT('h2)
	) name12907 (
		_w16949_,
		_w16953_,
		_w16954_
	);
	LUT2 #(
		.INIT('h1)
	) name12908 (
		_w14852_,
		_w16954_,
		_w16955_
	);
	LUT2 #(
		.INIT('h4)
	) name12909 (
		_w16759_,
		_w16763_,
		_w16956_
	);
	LUT2 #(
		.INIT('h1)
	) name12910 (
		_w16764_,
		_w16956_,
		_w16957_
	);
	LUT2 #(
		.INIT('h2)
	) name12911 (
		_w14852_,
		_w16957_,
		_w16958_
	);
	LUT2 #(
		.INIT('h2)
	) name12912 (
		_w16765_,
		_w16956_,
		_w16959_
	);
	LUT2 #(
		.INIT('h1)
	) name12913 (
		_w16958_,
		_w16959_,
		_w16960_
	);
	LUT2 #(
		.INIT('h4)
	) name12914 (
		_w16955_,
		_w16960_,
		_w16961_
	);
	LUT2 #(
		.INIT('h1)
	) name12915 (
		_w16956_,
		_w16960_,
		_w16962_
	);
	LUT2 #(
		.INIT('h1)
	) name12916 (
		_w16961_,
		_w16962_,
		_w16963_
	);
	LUT2 #(
		.INIT('h4)
	) name12917 (
		_w16764_,
		_w16768_,
		_w16964_
	);
	LUT2 #(
		.INIT('h1)
	) name12918 (
		_w16771_,
		_w16964_,
		_w16965_
	);
	LUT2 #(
		.INIT('h4)
	) name12919 (
		_w16963_,
		_w16965_,
		_w16966_
	);
	LUT2 #(
		.INIT('h1)
	) name12920 (
		_w16927_,
		_w16966_,
		_w16967_
	);
	LUT2 #(
		.INIT('h4)
	) name12921 (
		_w16741_,
		_w16773_,
		_w16968_
	);
	LUT2 #(
		.INIT('h1)
	) name12922 (
		_w16774_,
		_w16968_,
		_w16969_
	);
	LUT2 #(
		.INIT('h4)
	) name12923 (
		_w16776_,
		_w16842_,
		_w16970_
	);
	LUT2 #(
		.INIT('h1)
	) name12924 (
		_w16843_,
		_w16970_,
		_w16971_
	);
	LUT2 #(
		.INIT('h8)
	) name12925 (
		_w16969_,
		_w16971_,
		_w16972_
	);
	LUT2 #(
		.INIT('h1)
	) name12926 (
		_w16969_,
		_w16971_,
		_w16973_
	);
	LUT2 #(
		.INIT('h1)
	) name12927 (
		_w16972_,
		_w16973_,
		_w16974_
	);
	LUT2 #(
		.INIT('h4)
	) name12928 (
		_w16967_,
		_w16974_,
		_w16975_
	);
	LUT2 #(
		.INIT('h1)
	) name12929 (
		_w16968_,
		_w16970_,
		_w16976_
	);
	LUT2 #(
		.INIT('h4)
	) name12930 (
		_w16974_,
		_w16976_,
		_w16977_
	);
	LUT2 #(
		.INIT('h1)
	) name12931 (
		_w16975_,
		_w16977_,
		_w16978_
	);
	LUT2 #(
		.INIT('h1)
	) name12932 (
		_w16858_,
		_w16978_,
		_w16979_
	);
	LUT2 #(
		.INIT('h1)
	) name12933 (
		_w16856_,
		_w16979_,
		_w16980_
	);
	LUT2 #(
		.INIT('h1)
	) name12934 (
		_w16683_,
		_w16709_,
		_w16981_
	);
	LUT2 #(
		.INIT('h1)
	) name12935 (
		_w16669_,
		_w16678_,
		_w16982_
	);
	LUT2 #(
		.INIT('h1)
	) name12936 (
		_w16670_,
		_w16982_,
		_w16983_
	);
	LUT2 #(
		.INIT('h1)
	) name12937 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14914_,
		_w16984_
	);
	LUT2 #(
		.INIT('h2)
	) name12938 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14918_,
		_w16985_
	);
	LUT2 #(
		.INIT('h4)
	) name12939 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14925_,
		_w16986_
	);
	LUT2 #(
		.INIT('h8)
	) name12940 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14929_,
		_w16987_
	);
	LUT2 #(
		.INIT('h1)
	) name12941 (
		_w16986_,
		_w16987_,
		_w16988_
	);
	LUT2 #(
		.INIT('h4)
	) name12942 (
		_w16984_,
		_w16988_,
		_w16989_
	);
	LUT2 #(
		.INIT('h4)
	) name12943 (
		_w16985_,
		_w16989_,
		_w16990_
	);
	LUT2 #(
		.INIT('h8)
	) name12944 (
		_w14879_,
		_w16990_,
		_w16991_
	);
	LUT2 #(
		.INIT('h1)
	) name12945 (
		_w14879_,
		_w16990_,
		_w16992_
	);
	LUT2 #(
		.INIT('h1)
	) name12946 (
		_w16991_,
		_w16992_,
		_w16993_
	);
	LUT2 #(
		.INIT('h2)
	) name12947 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14891_,
		_w16994_
	);
	LUT2 #(
		.INIT('h1)
	) name12948 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14887_,
		_w16995_
	);
	LUT2 #(
		.INIT('h4)
	) name12949 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14898_,
		_w16996_
	);
	LUT2 #(
		.INIT('h8)
	) name12950 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14902_,
		_w16997_
	);
	LUT2 #(
		.INIT('h1)
	) name12951 (
		_w16996_,
		_w16997_,
		_w16998_
	);
	LUT2 #(
		.INIT('h4)
	) name12952 (
		_w16994_,
		_w16998_,
		_w16999_
	);
	LUT2 #(
		.INIT('h4)
	) name12953 (
		_w16995_,
		_w16999_,
		_w17000_
	);
	LUT2 #(
		.INIT('h4)
	) name12954 (
		_w16993_,
		_w17000_,
		_w17001_
	);
	LUT2 #(
		.INIT('h2)
	) name12955 (
		_w16993_,
		_w17000_,
		_w17002_
	);
	LUT2 #(
		.INIT('h1)
	) name12956 (
		_w17001_,
		_w17002_,
		_w17003_
	);
	LUT2 #(
		.INIT('h2)
	) name12957 (
		_w16983_,
		_w17003_,
		_w17004_
	);
	LUT2 #(
		.INIT('h4)
	) name12958 (
		_w16983_,
		_w17003_,
		_w17005_
	);
	LUT2 #(
		.INIT('h1)
	) name12959 (
		_w17004_,
		_w17005_,
		_w17006_
	);
	LUT2 #(
		.INIT('h1)
	) name12960 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14967_,
		_w17007_
	);
	LUT2 #(
		.INIT('h2)
	) name12961 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14969_,
		_w17008_
	);
	LUT2 #(
		.INIT('h1)
	) name12962 (
		_w17007_,
		_w17008_,
		_w17009_
	);
	LUT2 #(
		.INIT('h1)
	) name12963 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14947_,
		_w17010_
	);
	LUT2 #(
		.INIT('h2)
	) name12964 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14951_,
		_w17011_
	);
	LUT2 #(
		.INIT('h4)
	) name12965 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14958_,
		_w17012_
	);
	LUT2 #(
		.INIT('h8)
	) name12966 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14962_,
		_w17013_
	);
	LUT2 #(
		.INIT('h1)
	) name12967 (
		_w17012_,
		_w17013_,
		_w17014_
	);
	LUT2 #(
		.INIT('h4)
	) name12968 (
		_w17010_,
		_w17014_,
		_w17015_
	);
	LUT2 #(
		.INIT('h4)
	) name12969 (
		_w17011_,
		_w17015_,
		_w17016_
	);
	LUT2 #(
		.INIT('h2)
	) name12970 (
		_w17009_,
		_w17016_,
		_w17017_
	);
	LUT2 #(
		.INIT('h4)
	) name12971 (
		_w17009_,
		_w17016_,
		_w17018_
	);
	LUT2 #(
		.INIT('h1)
	) name12972 (
		_w17017_,
		_w17018_,
		_w17019_
	);
	LUT2 #(
		.INIT('h2)
	) name12973 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16699_,
		_w17020_
	);
	LUT2 #(
		.INIT('h1)
	) name12974 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15254_,
		_w17021_
	);
	LUT2 #(
		.INIT('h1)
	) name12975 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w17020_,
		_w17022_
	);
	LUT2 #(
		.INIT('h4)
	) name12976 (
		_w17021_,
		_w17022_,
		_w17023_
	);
	LUT2 #(
		.INIT('h4)
	) name12977 (
		_w17019_,
		_w17023_,
		_w17024_
	);
	LUT2 #(
		.INIT('h2)
	) name12978 (
		_w17019_,
		_w17023_,
		_w17025_
	);
	LUT2 #(
		.INIT('h1)
	) name12979 (
		_w17024_,
		_w17025_,
		_w17026_
	);
	LUT2 #(
		.INIT('h1)
	) name12980 (
		_w16696_,
		_w16702_,
		_w17027_
	);
	LUT2 #(
		.INIT('h1)
	) name12981 (
		_w16695_,
		_w17027_,
		_w17028_
	);
	LUT2 #(
		.INIT('h2)
	) name12982 (
		_w17026_,
		_w17028_,
		_w17029_
	);
	LUT2 #(
		.INIT('h4)
	) name12983 (
		_w17026_,
		_w17028_,
		_w17030_
	);
	LUT2 #(
		.INIT('h1)
	) name12984 (
		_w17029_,
		_w17030_,
		_w17031_
	);
	LUT2 #(
		.INIT('h8)
	) name12985 (
		_w17006_,
		_w17031_,
		_w17032_
	);
	LUT2 #(
		.INIT('h1)
	) name12986 (
		_w17006_,
		_w17031_,
		_w17033_
	);
	LUT2 #(
		.INIT('h1)
	) name12987 (
		_w17032_,
		_w17033_,
		_w17034_
	);
	LUT2 #(
		.INIT('h4)
	) name12988 (
		_w16981_,
		_w17034_,
		_w17035_
	);
	LUT2 #(
		.INIT('h2)
	) name12989 (
		_w16981_,
		_w17034_,
		_w17036_
	);
	LUT2 #(
		.INIT('h1)
	) name12990 (
		_w17035_,
		_w17036_,
		_w17037_
	);
	LUT2 #(
		.INIT('h1)
	) name12991 (
		_w16682_,
		_w16708_,
		_w17038_
	);
	LUT2 #(
		.INIT('h4)
	) name12992 (
		_w16713_,
		_w17038_,
		_w17039_
	);
	LUT2 #(
		.INIT('h1)
	) name12993 (
		_w16714_,
		_w17039_,
		_w17040_
	);
	LUT2 #(
		.INIT('h2)
	) name12994 (
		_w17037_,
		_w17040_,
		_w17041_
	);
	LUT2 #(
		.INIT('h1)
	) name12995 (
		_w14853_,
		_w17041_,
		_w17042_
	);
	LUT2 #(
		.INIT('h1)
	) name12996 (
		_w17004_,
		_w17029_,
		_w17043_
	);
	LUT2 #(
		.INIT('h1)
	) name12997 (
		_w16991_,
		_w17000_,
		_w17044_
	);
	LUT2 #(
		.INIT('h1)
	) name12998 (
		_w16992_,
		_w17044_,
		_w17045_
	);
	LUT2 #(
		.INIT('h1)
	) name12999 (
		_w15281_,
		_w15287_,
		_w17046_
	);
	LUT2 #(
		.INIT('h2)
	) name13000 (
		_w15285_,
		_w17046_,
		_w17047_
	);
	LUT2 #(
		.INIT('h4)
	) name13001 (
		_w15285_,
		_w17046_,
		_w17048_
	);
	LUT2 #(
		.INIT('h1)
	) name13002 (
		_w17047_,
		_w17048_,
		_w17049_
	);
	LUT2 #(
		.INIT('h4)
	) name13003 (
		_w17045_,
		_w17049_,
		_w17050_
	);
	LUT2 #(
		.INIT('h2)
	) name13004 (
		_w17045_,
		_w17049_,
		_w17051_
	);
	LUT2 #(
		.INIT('h1)
	) name13005 (
		_w17050_,
		_w17051_,
		_w17052_
	);
	LUT2 #(
		.INIT('h1)
	) name13006 (
		_w15266_,
		_w15267_,
		_w17053_
	);
	LUT2 #(
		.INIT('h4)
	) name13007 (
		_w15270_,
		_w17053_,
		_w17054_
	);
	LUT2 #(
		.INIT('h2)
	) name13008 (
		_w15270_,
		_w17053_,
		_w17055_
	);
	LUT2 #(
		.INIT('h1)
	) name13009 (
		_w17054_,
		_w17055_,
		_w17056_
	);
	LUT2 #(
		.INIT('h4)
	) name13010 (
		_w17018_,
		_w17023_,
		_w17057_
	);
	LUT2 #(
		.INIT('h1)
	) name13011 (
		_w17017_,
		_w17057_,
		_w17058_
	);
	LUT2 #(
		.INIT('h2)
	) name13012 (
		_w17056_,
		_w17058_,
		_w17059_
	);
	LUT2 #(
		.INIT('h4)
	) name13013 (
		_w17056_,
		_w17058_,
		_w17060_
	);
	LUT2 #(
		.INIT('h1)
	) name13014 (
		_w17059_,
		_w17060_,
		_w17061_
	);
	LUT2 #(
		.INIT('h8)
	) name13015 (
		_w17052_,
		_w17061_,
		_w17062_
	);
	LUT2 #(
		.INIT('h1)
	) name13016 (
		_w17052_,
		_w17061_,
		_w17063_
	);
	LUT2 #(
		.INIT('h1)
	) name13017 (
		_w17062_,
		_w17063_,
		_w17064_
	);
	LUT2 #(
		.INIT('h2)
	) name13018 (
		_w17043_,
		_w17064_,
		_w17065_
	);
	LUT2 #(
		.INIT('h4)
	) name13019 (
		_w17043_,
		_w17064_,
		_w17066_
	);
	LUT2 #(
		.INIT('h1)
	) name13020 (
		_w17065_,
		_w17066_,
		_w17067_
	);
	LUT2 #(
		.INIT('h1)
	) name13021 (
		_w17005_,
		_w17030_,
		_w17068_
	);
	LUT2 #(
		.INIT('h4)
	) name13022 (
		_w17034_,
		_w17068_,
		_w17069_
	);
	LUT2 #(
		.INIT('h1)
	) name13023 (
		_w17035_,
		_w17069_,
		_w17070_
	);
	LUT2 #(
		.INIT('h2)
	) name13024 (
		_w17067_,
		_w17070_,
		_w17071_
	);
	LUT2 #(
		.INIT('h4)
	) name13025 (
		_w17067_,
		_w17070_,
		_w17072_
	);
	LUT2 #(
		.INIT('h1)
	) name13026 (
		_w17071_,
		_w17072_,
		_w17073_
	);
	LUT2 #(
		.INIT('h8)
	) name13027 (
		_w14853_,
		_w17073_,
		_w17074_
	);
	LUT2 #(
		.INIT('h1)
	) name13028 (
		_w14853_,
		_w17073_,
		_w17075_
	);
	LUT2 #(
		.INIT('h1)
	) name13029 (
		_w17074_,
		_w17075_,
		_w17076_
	);
	LUT2 #(
		.INIT('h1)
	) name13030 (
		_w17042_,
		_w17076_,
		_w17077_
	);
	LUT2 #(
		.INIT('h8)
	) name13031 (
		_w17042_,
		_w17073_,
		_w17078_
	);
	LUT2 #(
		.INIT('h1)
	) name13032 (
		_w17077_,
		_w17078_,
		_w17079_
	);
	LUT2 #(
		.INIT('h1)
	) name13033 (
		_w16721_,
		_w16732_,
		_w17080_
	);
	LUT2 #(
		.INIT('h4)
	) name13034 (
		_w17037_,
		_w17040_,
		_w17081_
	);
	LUT2 #(
		.INIT('h1)
	) name13035 (
		_w17041_,
		_w17081_,
		_w17082_
	);
	LUT2 #(
		.INIT('h8)
	) name13036 (
		_w14853_,
		_w17082_,
		_w17083_
	);
	LUT2 #(
		.INIT('h1)
	) name13037 (
		_w14853_,
		_w17082_,
		_w17084_
	);
	LUT2 #(
		.INIT('h1)
	) name13038 (
		_w17083_,
		_w17084_,
		_w17085_
	);
	LUT2 #(
		.INIT('h1)
	) name13039 (
		_w17080_,
		_w17085_,
		_w17086_
	);
	LUT2 #(
		.INIT('h8)
	) name13040 (
		_w17080_,
		_w17085_,
		_w17087_
	);
	LUT2 #(
		.INIT('h1)
	) name13041 (
		_w17086_,
		_w17087_,
		_w17088_
	);
	LUT2 #(
		.INIT('h1)
	) name13042 (
		_w16720_,
		_w16731_,
		_w17089_
	);
	LUT2 #(
		.INIT('h4)
	) name13043 (
		_w16736_,
		_w17089_,
		_w17090_
	);
	LUT2 #(
		.INIT('h1)
	) name13044 (
		_w16737_,
		_w17090_,
		_w17091_
	);
	LUT2 #(
		.INIT('h2)
	) name13045 (
		_w17088_,
		_w17091_,
		_w17092_
	);
	LUT2 #(
		.INIT('h1)
	) name13046 (
		_w17079_,
		_w17092_,
		_w17093_
	);
	LUT2 #(
		.INIT('h4)
	) name13047 (
		_w17081_,
		_w17085_,
		_w17094_
	);
	LUT2 #(
		.INIT('h1)
	) name13048 (
		_w17086_,
		_w17094_,
		_w17095_
	);
	LUT2 #(
		.INIT('h8)
	) name13049 (
		_w17091_,
		_w17095_,
		_w17096_
	);
	LUT2 #(
		.INIT('h1)
	) name13050 (
		_w17093_,
		_w17096_,
		_w17097_
	);
	LUT2 #(
		.INIT('h2)
	) name13051 (
		_w16980_,
		_w17097_,
		_w17098_
	);
	LUT2 #(
		.INIT('h1)
	) name13052 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14787_,
		_w17099_
	);
	LUT2 #(
		.INIT('h2)
	) name13053 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14791_,
		_w17100_
	);
	LUT2 #(
		.INIT('h4)
	) name13054 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14798_,
		_w17101_
	);
	LUT2 #(
		.INIT('h8)
	) name13055 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14802_,
		_w17102_
	);
	LUT2 #(
		.INIT('h1)
	) name13056 (
		_w17101_,
		_w17102_,
		_w17103_
	);
	LUT2 #(
		.INIT('h4)
	) name13057 (
		_w17099_,
		_w17103_,
		_w17104_
	);
	LUT2 #(
		.INIT('h4)
	) name13058 (
		_w17100_,
		_w17104_,
		_w17105_
	);
	LUT2 #(
		.INIT('h1)
	) name13059 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14761_,
		_w17106_
	);
	LUT2 #(
		.INIT('h2)
	) name13060 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14765_,
		_w17107_
	);
	LUT2 #(
		.INIT('h4)
	) name13061 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14772_,
		_w17108_
	);
	LUT2 #(
		.INIT('h8)
	) name13062 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14776_,
		_w17109_
	);
	LUT2 #(
		.INIT('h1)
	) name13063 (
		_w17108_,
		_w17109_,
		_w17110_
	);
	LUT2 #(
		.INIT('h4)
	) name13064 (
		_w17106_,
		_w17110_,
		_w17111_
	);
	LUT2 #(
		.INIT('h4)
	) name13065 (
		_w17107_,
		_w17111_,
		_w17112_
	);
	LUT2 #(
		.INIT('h8)
	) name13066 (
		_w17105_,
		_w17112_,
		_w17113_
	);
	LUT2 #(
		.INIT('h1)
	) name13067 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14814_,
		_w17114_
	);
	LUT2 #(
		.INIT('h2)
	) name13068 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14818_,
		_w17115_
	);
	LUT2 #(
		.INIT('h4)
	) name13069 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14825_,
		_w17116_
	);
	LUT2 #(
		.INIT('h8)
	) name13070 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14829_,
		_w17117_
	);
	LUT2 #(
		.INIT('h1)
	) name13071 (
		_w17116_,
		_w17117_,
		_w17118_
	);
	LUT2 #(
		.INIT('h4)
	) name13072 (
		_w17114_,
		_w17118_,
		_w17119_
	);
	LUT2 #(
		.INIT('h4)
	) name13073 (
		_w17115_,
		_w17119_,
		_w17120_
	);
	LUT2 #(
		.INIT('h1)
	) name13074 (
		_w17113_,
		_w17120_,
		_w17121_
	);
	LUT2 #(
		.INIT('h1)
	) name13075 (
		_w17105_,
		_w17112_,
		_w17122_
	);
	LUT2 #(
		.INIT('h1)
	) name13076 (
		_w17121_,
		_w17122_,
		_w17123_
	);
	LUT2 #(
		.INIT('h1)
	) name13077 (
		_w16942_,
		_w16948_,
		_w17124_
	);
	LUT2 #(
		.INIT('h2)
	) name13078 (
		_w16946_,
		_w17124_,
		_w17125_
	);
	LUT2 #(
		.INIT('h4)
	) name13079 (
		_w16946_,
		_w17124_,
		_w17126_
	);
	LUT2 #(
		.INIT('h1)
	) name13080 (
		_w17125_,
		_w17126_,
		_w17127_
	);
	LUT2 #(
		.INIT('h2)
	) name13081 (
		_w17123_,
		_w17127_,
		_w17128_
	);
	LUT2 #(
		.INIT('h1)
	) name13082 (
		_w14852_,
		_w17128_,
		_w17129_
	);
	LUT2 #(
		.INIT('h4)
	) name13083 (
		_w16949_,
		_w16953_,
		_w17130_
	);
	LUT2 #(
		.INIT('h1)
	) name13084 (
		_w16954_,
		_w17130_,
		_w17131_
	);
	LUT2 #(
		.INIT('h4)
	) name13085 (
		_w14852_,
		_w17131_,
		_w17132_
	);
	LUT2 #(
		.INIT('h2)
	) name13086 (
		_w14852_,
		_w17131_,
		_w17133_
	);
	LUT2 #(
		.INIT('h1)
	) name13087 (
		_w17132_,
		_w17133_,
		_w17134_
	);
	LUT2 #(
		.INIT('h4)
	) name13088 (
		_w17129_,
		_w17134_,
		_w17135_
	);
	LUT2 #(
		.INIT('h4)
	) name13089 (
		_w17128_,
		_w17132_,
		_w17136_
	);
	LUT2 #(
		.INIT('h1)
	) name13090 (
		_w17135_,
		_w17136_,
		_w17137_
	);
	LUT2 #(
		.INIT('h1)
	) name13091 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14787_,
		_w17138_
	);
	LUT2 #(
		.INIT('h2)
	) name13092 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14791_,
		_w17139_
	);
	LUT2 #(
		.INIT('h4)
	) name13093 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14798_,
		_w17140_
	);
	LUT2 #(
		.INIT('h8)
	) name13094 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14802_,
		_w17141_
	);
	LUT2 #(
		.INIT('h1)
	) name13095 (
		_w17140_,
		_w17141_,
		_w17142_
	);
	LUT2 #(
		.INIT('h4)
	) name13096 (
		_w17138_,
		_w17142_,
		_w17143_
	);
	LUT2 #(
		.INIT('h4)
	) name13097 (
		_w17139_,
		_w17143_,
		_w17144_
	);
	LUT2 #(
		.INIT('h1)
	) name13098 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14761_,
		_w17145_
	);
	LUT2 #(
		.INIT('h2)
	) name13099 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14765_,
		_w17146_
	);
	LUT2 #(
		.INIT('h4)
	) name13100 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14772_,
		_w17147_
	);
	LUT2 #(
		.INIT('h8)
	) name13101 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14776_,
		_w17148_
	);
	LUT2 #(
		.INIT('h1)
	) name13102 (
		_w17147_,
		_w17148_,
		_w17149_
	);
	LUT2 #(
		.INIT('h4)
	) name13103 (
		_w17145_,
		_w17149_,
		_w17150_
	);
	LUT2 #(
		.INIT('h4)
	) name13104 (
		_w17146_,
		_w17150_,
		_w17151_
	);
	LUT2 #(
		.INIT('h8)
	) name13105 (
		_w17144_,
		_w17151_,
		_w17152_
	);
	LUT2 #(
		.INIT('h1)
	) name13106 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14814_,
		_w17153_
	);
	LUT2 #(
		.INIT('h2)
	) name13107 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14818_,
		_w17154_
	);
	LUT2 #(
		.INIT('h4)
	) name13108 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14825_,
		_w17155_
	);
	LUT2 #(
		.INIT('h8)
	) name13109 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14829_,
		_w17156_
	);
	LUT2 #(
		.INIT('h1)
	) name13110 (
		_w17155_,
		_w17156_,
		_w17157_
	);
	LUT2 #(
		.INIT('h4)
	) name13111 (
		_w17153_,
		_w17157_,
		_w17158_
	);
	LUT2 #(
		.INIT('h4)
	) name13112 (
		_w17154_,
		_w17158_,
		_w17159_
	);
	LUT2 #(
		.INIT('h1)
	) name13113 (
		_w17152_,
		_w17159_,
		_w17160_
	);
	LUT2 #(
		.INIT('h1)
	) name13114 (
		_w17144_,
		_w17151_,
		_w17161_
	);
	LUT2 #(
		.INIT('h1)
	) name13115 (
		_w17160_,
		_w17161_,
		_w17162_
	);
	LUT2 #(
		.INIT('h1)
	) name13116 (
		_w17113_,
		_w17122_,
		_w17163_
	);
	LUT2 #(
		.INIT('h2)
	) name13117 (
		_w17120_,
		_w17163_,
		_w17164_
	);
	LUT2 #(
		.INIT('h4)
	) name13118 (
		_w17120_,
		_w17163_,
		_w17165_
	);
	LUT2 #(
		.INIT('h1)
	) name13119 (
		_w17164_,
		_w17165_,
		_w17166_
	);
	LUT2 #(
		.INIT('h2)
	) name13120 (
		_w17162_,
		_w17166_,
		_w17167_
	);
	LUT2 #(
		.INIT('h4)
	) name13121 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14846_,
		_w17168_
	);
	LUT2 #(
		.INIT('h8)
	) name13122 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14849_,
		_w17169_
	);
	LUT2 #(
		.INIT('h1)
	) name13123 (
		_w17168_,
		_w17169_,
		_w17170_
	);
	LUT2 #(
		.INIT('h8)
	) name13124 (
		_w14844_,
		_w17170_,
		_w17171_
	);
	LUT2 #(
		.INIT('h2)
	) name13125 (
		_w14967_,
		_w17171_,
		_w17172_
	);
	LUT2 #(
		.INIT('h2)
	) name13126 (
		_w14852_,
		_w17172_,
		_w17173_
	);
	LUT2 #(
		.INIT('h1)
	) name13127 (
		_w17167_,
		_w17173_,
		_w17174_
	);
	LUT2 #(
		.INIT('h4)
	) name13128 (
		_w17123_,
		_w17127_,
		_w17175_
	);
	LUT2 #(
		.INIT('h1)
	) name13129 (
		_w17128_,
		_w17175_,
		_w17176_
	);
	LUT2 #(
		.INIT('h2)
	) name13130 (
		_w14852_,
		_w17176_,
		_w17177_
	);
	LUT2 #(
		.INIT('h4)
	) name13131 (
		_w14852_,
		_w17176_,
		_w17178_
	);
	LUT2 #(
		.INIT('h1)
	) name13132 (
		_w17177_,
		_w17178_,
		_w17179_
	);
	LUT2 #(
		.INIT('h8)
	) name13133 (
		_w17174_,
		_w17179_,
		_w17180_
	);
	LUT2 #(
		.INIT('h8)
	) name13134 (
		_w14852_,
		_w17175_,
		_w17181_
	);
	LUT2 #(
		.INIT('h1)
	) name13135 (
		_w17180_,
		_w17181_,
		_w17182_
	);
	LUT2 #(
		.INIT('h8)
	) name13136 (
		_w17137_,
		_w17182_,
		_w17183_
	);
	LUT2 #(
		.INIT('h1)
	) name13137 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14861_,
		_w17184_
	);
	LUT2 #(
		.INIT('h2)
	) name13138 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14865_,
		_w17185_
	);
	LUT2 #(
		.INIT('h4)
	) name13139 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14872_,
		_w17186_
	);
	LUT2 #(
		.INIT('h8)
	) name13140 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14876_,
		_w17187_
	);
	LUT2 #(
		.INIT('h1)
	) name13141 (
		_w17186_,
		_w17187_,
		_w17188_
	);
	LUT2 #(
		.INIT('h4)
	) name13142 (
		_w17184_,
		_w17188_,
		_w17189_
	);
	LUT2 #(
		.INIT('h4)
	) name13143 (
		_w17185_,
		_w17189_,
		_w17190_
	);
	LUT2 #(
		.INIT('h1)
	) name13144 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14914_,
		_w17191_
	);
	LUT2 #(
		.INIT('h2)
	) name13145 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14918_,
		_w17192_
	);
	LUT2 #(
		.INIT('h4)
	) name13146 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14925_,
		_w17193_
	);
	LUT2 #(
		.INIT('h8)
	) name13147 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14929_,
		_w17194_
	);
	LUT2 #(
		.INIT('h1)
	) name13148 (
		_w17193_,
		_w17194_,
		_w17195_
	);
	LUT2 #(
		.INIT('h4)
	) name13149 (
		_w17191_,
		_w17195_,
		_w17196_
	);
	LUT2 #(
		.INIT('h4)
	) name13150 (
		_w17192_,
		_w17196_,
		_w17197_
	);
	LUT2 #(
		.INIT('h8)
	) name13151 (
		_w17190_,
		_w17197_,
		_w17198_
	);
	LUT2 #(
		.INIT('h1)
	) name13152 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14887_,
		_w17199_
	);
	LUT2 #(
		.INIT('h2)
	) name13153 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14891_,
		_w17200_
	);
	LUT2 #(
		.INIT('h4)
	) name13154 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14898_,
		_w17201_
	);
	LUT2 #(
		.INIT('h8)
	) name13155 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14902_,
		_w17202_
	);
	LUT2 #(
		.INIT('h1)
	) name13156 (
		_w17201_,
		_w17202_,
		_w17203_
	);
	LUT2 #(
		.INIT('h4)
	) name13157 (
		_w17199_,
		_w17203_,
		_w17204_
	);
	LUT2 #(
		.INIT('h4)
	) name13158 (
		_w17200_,
		_w17204_,
		_w17205_
	);
	LUT2 #(
		.INIT('h1)
	) name13159 (
		_w17198_,
		_w17205_,
		_w17206_
	);
	LUT2 #(
		.INIT('h1)
	) name13160 (
		_w17190_,
		_w17197_,
		_w17207_
	);
	LUT2 #(
		.INIT('h1)
	) name13161 (
		_w17206_,
		_w17207_,
		_w17208_
	);
	LUT2 #(
		.INIT('h1)
	) name13162 (
		_w16875_,
		_w16884_,
		_w17209_
	);
	LUT2 #(
		.INIT('h2)
	) name13163 (
		_w16882_,
		_w17209_,
		_w17210_
	);
	LUT2 #(
		.INIT('h4)
	) name13164 (
		_w16882_,
		_w17209_,
		_w17211_
	);
	LUT2 #(
		.INIT('h1)
	) name13165 (
		_w17210_,
		_w17211_,
		_w17212_
	);
	LUT2 #(
		.INIT('h2)
	) name13166 (
		_w17208_,
		_w17212_,
		_w17213_
	);
	LUT2 #(
		.INIT('h1)
	) name13167 (
		_w16907_,
		_w16908_,
		_w17214_
	);
	LUT2 #(
		.INIT('h4)
	) name13168 (
		_w16911_,
		_w17214_,
		_w17215_
	);
	LUT2 #(
		.INIT('h2)
	) name13169 (
		_w16911_,
		_w17214_,
		_w17216_
	);
	LUT2 #(
		.INIT('h1)
	) name13170 (
		_w17215_,
		_w17216_,
		_w17217_
	);
	LUT2 #(
		.INIT('h2)
	) name13171 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w9205_,
		_w17218_
	);
	LUT2 #(
		.INIT('h2)
	) name13172 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17218_,
		_w17219_
	);
	LUT2 #(
		.INIT('h1)
	) name13173 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w16895_,
		_w17220_
	);
	LUT2 #(
		.INIT('h1)
	) name13174 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w17219_,
		_w17221_
	);
	LUT2 #(
		.INIT('h4)
	) name13175 (
		_w17220_,
		_w17221_,
		_w17222_
	);
	LUT2 #(
		.INIT('h1)
	) name13176 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14947_,
		_w17223_
	);
	LUT2 #(
		.INIT('h2)
	) name13177 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14951_,
		_w17224_
	);
	LUT2 #(
		.INIT('h4)
	) name13178 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14958_,
		_w17225_
	);
	LUT2 #(
		.INIT('h8)
	) name13179 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14962_,
		_w17226_
	);
	LUT2 #(
		.INIT('h1)
	) name13180 (
		_w17225_,
		_w17226_,
		_w17227_
	);
	LUT2 #(
		.INIT('h4)
	) name13181 (
		_w17223_,
		_w17227_,
		_w17228_
	);
	LUT2 #(
		.INIT('h4)
	) name13182 (
		_w17224_,
		_w17228_,
		_w17229_
	);
	LUT2 #(
		.INIT('h2)
	) name13183 (
		_w17222_,
		_w17229_,
		_w17230_
	);
	LUT2 #(
		.INIT('h4)
	) name13184 (
		_w17222_,
		_w17229_,
		_w17231_
	);
	LUT2 #(
		.INIT('h4)
	) name13185 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14967_,
		_w17232_
	);
	LUT2 #(
		.INIT('h8)
	) name13186 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14969_,
		_w17233_
	);
	LUT2 #(
		.INIT('h1)
	) name13187 (
		_w17232_,
		_w17233_,
		_w17234_
	);
	LUT2 #(
		.INIT('h1)
	) name13188 (
		_w17231_,
		_w17234_,
		_w17235_
	);
	LUT2 #(
		.INIT('h1)
	) name13189 (
		_w17230_,
		_w17235_,
		_w17236_
	);
	LUT2 #(
		.INIT('h4)
	) name13190 (
		_w17217_,
		_w17236_,
		_w17237_
	);
	LUT2 #(
		.INIT('h1)
	) name13191 (
		_w17213_,
		_w17237_,
		_w17238_
	);
	LUT2 #(
		.INIT('h4)
	) name13192 (
		_w16885_,
		_w16889_,
		_w17239_
	);
	LUT2 #(
		.INIT('h1)
	) name13193 (
		_w16890_,
		_w17239_,
		_w17240_
	);
	LUT2 #(
		.INIT('h1)
	) name13194 (
		_w16894_,
		_w16913_,
		_w17241_
	);
	LUT2 #(
		.INIT('h1)
	) name13195 (
		_w16914_,
		_w17241_,
		_w17242_
	);
	LUT2 #(
		.INIT('h8)
	) name13196 (
		_w17240_,
		_w17242_,
		_w17243_
	);
	LUT2 #(
		.INIT('h1)
	) name13197 (
		_w17240_,
		_w17242_,
		_w17244_
	);
	LUT2 #(
		.INIT('h1)
	) name13198 (
		_w17243_,
		_w17244_,
		_w17245_
	);
	LUT2 #(
		.INIT('h4)
	) name13199 (
		_w17238_,
		_w17245_,
		_w17246_
	);
	LUT2 #(
		.INIT('h2)
	) name13200 (
		_w17238_,
		_w17245_,
		_w17247_
	);
	LUT2 #(
		.INIT('h1)
	) name13201 (
		_w17246_,
		_w17247_,
		_w17248_
	);
	LUT2 #(
		.INIT('h1)
	) name13202 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14887_,
		_w17249_
	);
	LUT2 #(
		.INIT('h2)
	) name13203 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14891_,
		_w17250_
	);
	LUT2 #(
		.INIT('h4)
	) name13204 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14898_,
		_w17251_
	);
	LUT2 #(
		.INIT('h8)
	) name13205 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14902_,
		_w17252_
	);
	LUT2 #(
		.INIT('h1)
	) name13206 (
		_w17251_,
		_w17252_,
		_w17253_
	);
	LUT2 #(
		.INIT('h4)
	) name13207 (
		_w17249_,
		_w17253_,
		_w17254_
	);
	LUT2 #(
		.INIT('h4)
	) name13208 (
		_w17250_,
		_w17254_,
		_w17255_
	);
	LUT2 #(
		.INIT('h1)
	) name13209 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14861_,
		_w17256_
	);
	LUT2 #(
		.INIT('h2)
	) name13210 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14865_,
		_w17257_
	);
	LUT2 #(
		.INIT('h4)
	) name13211 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14872_,
		_w17258_
	);
	LUT2 #(
		.INIT('h8)
	) name13212 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14876_,
		_w17259_
	);
	LUT2 #(
		.INIT('h1)
	) name13213 (
		_w17258_,
		_w17259_,
		_w17260_
	);
	LUT2 #(
		.INIT('h4)
	) name13214 (
		_w17256_,
		_w17260_,
		_w17261_
	);
	LUT2 #(
		.INIT('h4)
	) name13215 (
		_w17257_,
		_w17261_,
		_w17262_
	);
	LUT2 #(
		.INIT('h8)
	) name13216 (
		_w17255_,
		_w17262_,
		_w17263_
	);
	LUT2 #(
		.INIT('h1)
	) name13217 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14914_,
		_w17264_
	);
	LUT2 #(
		.INIT('h2)
	) name13218 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14918_,
		_w17265_
	);
	LUT2 #(
		.INIT('h4)
	) name13219 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14925_,
		_w17266_
	);
	LUT2 #(
		.INIT('h8)
	) name13220 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14929_,
		_w17267_
	);
	LUT2 #(
		.INIT('h1)
	) name13221 (
		_w17266_,
		_w17267_,
		_w17268_
	);
	LUT2 #(
		.INIT('h4)
	) name13222 (
		_w17264_,
		_w17268_,
		_w17269_
	);
	LUT2 #(
		.INIT('h4)
	) name13223 (
		_w17265_,
		_w17269_,
		_w17270_
	);
	LUT2 #(
		.INIT('h1)
	) name13224 (
		_w17263_,
		_w17270_,
		_w17271_
	);
	LUT2 #(
		.INIT('h1)
	) name13225 (
		_w17255_,
		_w17262_,
		_w17272_
	);
	LUT2 #(
		.INIT('h1)
	) name13226 (
		_w17271_,
		_w17272_,
		_w17273_
	);
	LUT2 #(
		.INIT('h1)
	) name13227 (
		_w17198_,
		_w17207_,
		_w17274_
	);
	LUT2 #(
		.INIT('h2)
	) name13228 (
		_w17205_,
		_w17274_,
		_w17275_
	);
	LUT2 #(
		.INIT('h4)
	) name13229 (
		_w17205_,
		_w17274_,
		_w17276_
	);
	LUT2 #(
		.INIT('h1)
	) name13230 (
		_w17275_,
		_w17276_,
		_w17277_
	);
	LUT2 #(
		.INIT('h2)
	) name13231 (
		_w17273_,
		_w17277_,
		_w17278_
	);
	LUT2 #(
		.INIT('h1)
	) name13232 (
		_w17230_,
		_w17231_,
		_w17279_
	);
	LUT2 #(
		.INIT('h4)
	) name13233 (
		_w17234_,
		_w17279_,
		_w17280_
	);
	LUT2 #(
		.INIT('h2)
	) name13234 (
		_w17234_,
		_w17279_,
		_w17281_
	);
	LUT2 #(
		.INIT('h1)
	) name13235 (
		_w17280_,
		_w17281_,
		_w17282_
	);
	LUT2 #(
		.INIT('h2)
	) name13236 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w7449_,
		_w17283_
	);
	LUT2 #(
		.INIT('h2)
	) name13237 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17283_,
		_w17284_
	);
	LUT2 #(
		.INIT('h1)
	) name13238 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17218_,
		_w17285_
	);
	LUT2 #(
		.INIT('h1)
	) name13239 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w17284_,
		_w17286_
	);
	LUT2 #(
		.INIT('h4)
	) name13240 (
		_w17285_,
		_w17286_,
		_w17287_
	);
	LUT2 #(
		.INIT('h1)
	) name13241 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14947_,
		_w17288_
	);
	LUT2 #(
		.INIT('h2)
	) name13242 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14951_,
		_w17289_
	);
	LUT2 #(
		.INIT('h4)
	) name13243 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14958_,
		_w17290_
	);
	LUT2 #(
		.INIT('h8)
	) name13244 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14962_,
		_w17291_
	);
	LUT2 #(
		.INIT('h1)
	) name13245 (
		_w17290_,
		_w17291_,
		_w17292_
	);
	LUT2 #(
		.INIT('h4)
	) name13246 (
		_w17288_,
		_w17292_,
		_w17293_
	);
	LUT2 #(
		.INIT('h4)
	) name13247 (
		_w17289_,
		_w17293_,
		_w17294_
	);
	LUT2 #(
		.INIT('h2)
	) name13248 (
		_w17287_,
		_w17294_,
		_w17295_
	);
	LUT2 #(
		.INIT('h4)
	) name13249 (
		_w17287_,
		_w17294_,
		_w17296_
	);
	LUT2 #(
		.INIT('h4)
	) name13250 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14967_,
		_w17297_
	);
	LUT2 #(
		.INIT('h8)
	) name13251 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14969_,
		_w17298_
	);
	LUT2 #(
		.INIT('h1)
	) name13252 (
		_w17297_,
		_w17298_,
		_w17299_
	);
	LUT2 #(
		.INIT('h1)
	) name13253 (
		_w17296_,
		_w17299_,
		_w17300_
	);
	LUT2 #(
		.INIT('h1)
	) name13254 (
		_w17295_,
		_w17300_,
		_w17301_
	);
	LUT2 #(
		.INIT('h4)
	) name13255 (
		_w17282_,
		_w17301_,
		_w17302_
	);
	LUT2 #(
		.INIT('h1)
	) name13256 (
		_w17278_,
		_w17302_,
		_w17303_
	);
	LUT2 #(
		.INIT('h4)
	) name13257 (
		_w17208_,
		_w17212_,
		_w17304_
	);
	LUT2 #(
		.INIT('h1)
	) name13258 (
		_w17213_,
		_w17304_,
		_w17305_
	);
	LUT2 #(
		.INIT('h2)
	) name13259 (
		_w17217_,
		_w17236_,
		_w17306_
	);
	LUT2 #(
		.INIT('h1)
	) name13260 (
		_w17237_,
		_w17306_,
		_w17307_
	);
	LUT2 #(
		.INIT('h8)
	) name13261 (
		_w17305_,
		_w17307_,
		_w17308_
	);
	LUT2 #(
		.INIT('h1)
	) name13262 (
		_w17305_,
		_w17307_,
		_w17309_
	);
	LUT2 #(
		.INIT('h1)
	) name13263 (
		_w17308_,
		_w17309_,
		_w17310_
	);
	LUT2 #(
		.INIT('h4)
	) name13264 (
		_w17303_,
		_w17310_,
		_w17311_
	);
	LUT2 #(
		.INIT('h1)
	) name13265 (
		_w17304_,
		_w17306_,
		_w17312_
	);
	LUT2 #(
		.INIT('h4)
	) name13266 (
		_w17310_,
		_w17312_,
		_w17313_
	);
	LUT2 #(
		.INIT('h1)
	) name13267 (
		_w17311_,
		_w17313_,
		_w17314_
	);
	LUT2 #(
		.INIT('h2)
	) name13268 (
		_w17248_,
		_w17314_,
		_w17315_
	);
	LUT2 #(
		.INIT('h1)
	) name13269 (
		_w17183_,
		_w17315_,
		_w17316_
	);
	LUT2 #(
		.INIT('h4)
	) name13270 (
		_w16915_,
		_w16922_,
		_w17317_
	);
	LUT2 #(
		.INIT('h1)
	) name13271 (
		_w16923_,
		_w17317_,
		_w17318_
	);
	LUT2 #(
		.INIT('h1)
	) name13272 (
		_w17239_,
		_w17241_,
		_w17319_
	);
	LUT2 #(
		.INIT('h4)
	) name13273 (
		_w17245_,
		_w17319_,
		_w17320_
	);
	LUT2 #(
		.INIT('h1)
	) name13274 (
		_w17246_,
		_w17320_,
		_w17321_
	);
	LUT2 #(
		.INIT('h1)
	) name13275 (
		_w17318_,
		_w17321_,
		_w17322_
	);
	LUT2 #(
		.INIT('h8)
	) name13276 (
		_w17318_,
		_w17321_,
		_w17323_
	);
	LUT2 #(
		.INIT('h1)
	) name13277 (
		_w17322_,
		_w17323_,
		_w17324_
	);
	LUT2 #(
		.INIT('h8)
	) name13278 (
		_w16955_,
		_w16957_,
		_w17325_
	);
	LUT2 #(
		.INIT('h1)
	) name13279 (
		_w16961_,
		_w17325_,
		_w17326_
	);
	LUT2 #(
		.INIT('h1)
	) name13280 (
		_w17130_,
		_w17134_,
		_w17327_
	);
	LUT2 #(
		.INIT('h1)
	) name13281 (
		_w17135_,
		_w17327_,
		_w17328_
	);
	LUT2 #(
		.INIT('h4)
	) name13282 (
		_w17326_,
		_w17328_,
		_w17329_
	);
	LUT2 #(
		.INIT('h2)
	) name13283 (
		_w17326_,
		_w17328_,
		_w17330_
	);
	LUT2 #(
		.INIT('h1)
	) name13284 (
		_w17329_,
		_w17330_,
		_w17331_
	);
	LUT2 #(
		.INIT('h8)
	) name13285 (
		_w17324_,
		_w17331_,
		_w17332_
	);
	LUT2 #(
		.INIT('h1)
	) name13286 (
		_w17324_,
		_w17331_,
		_w17333_
	);
	LUT2 #(
		.INIT('h1)
	) name13287 (
		_w17332_,
		_w17333_,
		_w17334_
	);
	LUT2 #(
		.INIT('h1)
	) name13288 (
		_w17316_,
		_w17334_,
		_w17335_
	);
	LUT2 #(
		.INIT('h8)
	) name13289 (
		_w17316_,
		_w17334_,
		_w17336_
	);
	LUT2 #(
		.INIT('h1)
	) name13290 (
		_w17335_,
		_w17336_,
		_w17337_
	);
	LUT2 #(
		.INIT('h2)
	) name13291 (
		_w17303_,
		_w17310_,
		_w17338_
	);
	LUT2 #(
		.INIT('h1)
	) name13292 (
		_w17311_,
		_w17338_,
		_w17339_
	);
	LUT2 #(
		.INIT('h8)
	) name13293 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 ,
		_w17340_
	);
	LUT2 #(
		.INIT('h1)
	) name13294 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w17341_
	);
	LUT2 #(
		.INIT('h8)
	) name13295 (
		_w17283_,
		_w17341_,
		_w17342_
	);
	LUT2 #(
		.INIT('h1)
	) name13296 (
		_w17340_,
		_w17342_,
		_w17343_
	);
	LUT2 #(
		.INIT('h2)
	) name13297 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14951_,
		_w17344_
	);
	LUT2 #(
		.INIT('h1)
	) name13298 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w14947_,
		_w17345_
	);
	LUT2 #(
		.INIT('h4)
	) name13299 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14958_,
		_w17346_
	);
	LUT2 #(
		.INIT('h8)
	) name13300 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w14962_,
		_w17347_
	);
	LUT2 #(
		.INIT('h1)
	) name13301 (
		_w17346_,
		_w17347_,
		_w17348_
	);
	LUT2 #(
		.INIT('h4)
	) name13302 (
		_w17344_,
		_w17348_,
		_w17349_
	);
	LUT2 #(
		.INIT('h4)
	) name13303 (
		_w17345_,
		_w17349_,
		_w17350_
	);
	LUT2 #(
		.INIT('h1)
	) name13304 (
		_w17343_,
		_w17350_,
		_w17351_
	);
	LUT2 #(
		.INIT('h1)
	) name13305 (
		_w17295_,
		_w17296_,
		_w17352_
	);
	LUT2 #(
		.INIT('h4)
	) name13306 (
		_w17299_,
		_w17352_,
		_w17353_
	);
	LUT2 #(
		.INIT('h2)
	) name13307 (
		_w17299_,
		_w17352_,
		_w17354_
	);
	LUT2 #(
		.INIT('h1)
	) name13308 (
		_w17353_,
		_w17354_,
		_w17355_
	);
	LUT2 #(
		.INIT('h1)
	) name13309 (
		_w17351_,
		_w17355_,
		_w17356_
	);
	LUT2 #(
		.INIT('h1)
	) name13310 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14887_,
		_w17357_
	);
	LUT2 #(
		.INIT('h2)
	) name13311 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w14891_,
		_w17358_
	);
	LUT2 #(
		.INIT('h4)
	) name13312 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14898_,
		_w17359_
	);
	LUT2 #(
		.INIT('h8)
	) name13313 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w14902_,
		_w17360_
	);
	LUT2 #(
		.INIT('h1)
	) name13314 (
		_w17359_,
		_w17360_,
		_w17361_
	);
	LUT2 #(
		.INIT('h4)
	) name13315 (
		_w17357_,
		_w17361_,
		_w17362_
	);
	LUT2 #(
		.INIT('h4)
	) name13316 (
		_w17358_,
		_w17362_,
		_w17363_
	);
	LUT2 #(
		.INIT('h1)
	) name13317 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14861_,
		_w17364_
	);
	LUT2 #(
		.INIT('h2)
	) name13318 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w14865_,
		_w17365_
	);
	LUT2 #(
		.INIT('h4)
	) name13319 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14872_,
		_w17366_
	);
	LUT2 #(
		.INIT('h8)
	) name13320 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w14876_,
		_w17367_
	);
	LUT2 #(
		.INIT('h1)
	) name13321 (
		_w17366_,
		_w17367_,
		_w17368_
	);
	LUT2 #(
		.INIT('h4)
	) name13322 (
		_w17364_,
		_w17368_,
		_w17369_
	);
	LUT2 #(
		.INIT('h4)
	) name13323 (
		_w17365_,
		_w17369_,
		_w17370_
	);
	LUT2 #(
		.INIT('h8)
	) name13324 (
		_w17363_,
		_w17370_,
		_w17371_
	);
	LUT2 #(
		.INIT('h1)
	) name13325 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14914_,
		_w17372_
	);
	LUT2 #(
		.INIT('h2)
	) name13326 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w14918_,
		_w17373_
	);
	LUT2 #(
		.INIT('h4)
	) name13327 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14925_,
		_w17374_
	);
	LUT2 #(
		.INIT('h8)
	) name13328 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w14929_,
		_w17375_
	);
	LUT2 #(
		.INIT('h1)
	) name13329 (
		_w17374_,
		_w17375_,
		_w17376_
	);
	LUT2 #(
		.INIT('h4)
	) name13330 (
		_w17372_,
		_w17376_,
		_w17377_
	);
	LUT2 #(
		.INIT('h4)
	) name13331 (
		_w17373_,
		_w17377_,
		_w17378_
	);
	LUT2 #(
		.INIT('h1)
	) name13332 (
		_w17371_,
		_w17378_,
		_w17379_
	);
	LUT2 #(
		.INIT('h1)
	) name13333 (
		_w17363_,
		_w17370_,
		_w17380_
	);
	LUT2 #(
		.INIT('h1)
	) name13334 (
		_w17379_,
		_w17380_,
		_w17381_
	);
	LUT2 #(
		.INIT('h1)
	) name13335 (
		_w17263_,
		_w17272_,
		_w17382_
	);
	LUT2 #(
		.INIT('h2)
	) name13336 (
		_w17270_,
		_w17382_,
		_w17383_
	);
	LUT2 #(
		.INIT('h4)
	) name13337 (
		_w17270_,
		_w17382_,
		_w17384_
	);
	LUT2 #(
		.INIT('h1)
	) name13338 (
		_w17383_,
		_w17384_,
		_w17385_
	);
	LUT2 #(
		.INIT('h2)
	) name13339 (
		_w17381_,
		_w17385_,
		_w17386_
	);
	LUT2 #(
		.INIT('h1)
	) name13340 (
		_w17356_,
		_w17386_,
		_w17387_
	);
	LUT2 #(
		.INIT('h4)
	) name13341 (
		_w17273_,
		_w17277_,
		_w17388_
	);
	LUT2 #(
		.INIT('h1)
	) name13342 (
		_w17278_,
		_w17388_,
		_w17389_
	);
	LUT2 #(
		.INIT('h2)
	) name13343 (
		_w17282_,
		_w17301_,
		_w17390_
	);
	LUT2 #(
		.INIT('h1)
	) name13344 (
		_w17302_,
		_w17390_,
		_w17391_
	);
	LUT2 #(
		.INIT('h2)
	) name13345 (
		_w17389_,
		_w17391_,
		_w17392_
	);
	LUT2 #(
		.INIT('h4)
	) name13346 (
		_w17389_,
		_w17391_,
		_w17393_
	);
	LUT2 #(
		.INIT('h1)
	) name13347 (
		_w17392_,
		_w17393_,
		_w17394_
	);
	LUT2 #(
		.INIT('h2)
	) name13348 (
		_w17387_,
		_w17394_,
		_w17395_
	);
	LUT2 #(
		.INIT('h1)
	) name13349 (
		_w17388_,
		_w17390_,
		_w17396_
	);
	LUT2 #(
		.INIT('h2)
	) name13350 (
		_w17394_,
		_w17396_,
		_w17397_
	);
	LUT2 #(
		.INIT('h1)
	) name13351 (
		_w17395_,
		_w17397_,
		_w17398_
	);
	LUT2 #(
		.INIT('h8)
	) name13352 (
		_w17339_,
		_w17398_,
		_w17399_
	);
	LUT2 #(
		.INIT('h1)
	) name13353 (
		_w17174_,
		_w17179_,
		_w17400_
	);
	LUT2 #(
		.INIT('h1)
	) name13354 (
		_w17180_,
		_w17400_,
		_w17401_
	);
	LUT2 #(
		.INIT('h1)
	) name13355 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14787_,
		_w17402_
	);
	LUT2 #(
		.INIT('h2)
	) name13356 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w14791_,
		_w17403_
	);
	LUT2 #(
		.INIT('h4)
	) name13357 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14798_,
		_w17404_
	);
	LUT2 #(
		.INIT('h8)
	) name13358 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w14802_,
		_w17405_
	);
	LUT2 #(
		.INIT('h1)
	) name13359 (
		_w17404_,
		_w17405_,
		_w17406_
	);
	LUT2 #(
		.INIT('h4)
	) name13360 (
		_w17402_,
		_w17406_,
		_w17407_
	);
	LUT2 #(
		.INIT('h4)
	) name13361 (
		_w17403_,
		_w17407_,
		_w17408_
	);
	LUT2 #(
		.INIT('h1)
	) name13362 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14761_,
		_w17409_
	);
	LUT2 #(
		.INIT('h2)
	) name13363 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w14765_,
		_w17410_
	);
	LUT2 #(
		.INIT('h4)
	) name13364 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14772_,
		_w17411_
	);
	LUT2 #(
		.INIT('h8)
	) name13365 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w14776_,
		_w17412_
	);
	LUT2 #(
		.INIT('h1)
	) name13366 (
		_w17411_,
		_w17412_,
		_w17413_
	);
	LUT2 #(
		.INIT('h4)
	) name13367 (
		_w17409_,
		_w17413_,
		_w17414_
	);
	LUT2 #(
		.INIT('h4)
	) name13368 (
		_w17410_,
		_w17414_,
		_w17415_
	);
	LUT2 #(
		.INIT('h8)
	) name13369 (
		_w17408_,
		_w17415_,
		_w17416_
	);
	LUT2 #(
		.INIT('h1)
	) name13370 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14814_,
		_w17417_
	);
	LUT2 #(
		.INIT('h2)
	) name13371 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w14818_,
		_w17418_
	);
	LUT2 #(
		.INIT('h4)
	) name13372 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14825_,
		_w17419_
	);
	LUT2 #(
		.INIT('h8)
	) name13373 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w14829_,
		_w17420_
	);
	LUT2 #(
		.INIT('h1)
	) name13374 (
		_w17419_,
		_w17420_,
		_w17421_
	);
	LUT2 #(
		.INIT('h4)
	) name13375 (
		_w17417_,
		_w17421_,
		_w17422_
	);
	LUT2 #(
		.INIT('h4)
	) name13376 (
		_w17418_,
		_w17422_,
		_w17423_
	);
	LUT2 #(
		.INIT('h1)
	) name13377 (
		_w17416_,
		_w17423_,
		_w17424_
	);
	LUT2 #(
		.INIT('h1)
	) name13378 (
		_w17408_,
		_w17415_,
		_w17425_
	);
	LUT2 #(
		.INIT('h1)
	) name13379 (
		_w17424_,
		_w17425_,
		_w17426_
	);
	LUT2 #(
		.INIT('h1)
	) name13380 (
		_w17152_,
		_w17161_,
		_w17427_
	);
	LUT2 #(
		.INIT('h2)
	) name13381 (
		_w17159_,
		_w17427_,
		_w17428_
	);
	LUT2 #(
		.INIT('h4)
	) name13382 (
		_w17159_,
		_w17427_,
		_w17429_
	);
	LUT2 #(
		.INIT('h1)
	) name13383 (
		_w17428_,
		_w17429_,
		_w17430_
	);
	LUT2 #(
		.INIT('h2)
	) name13384 (
		_w17426_,
		_w17430_,
		_w17431_
	);
	LUT2 #(
		.INIT('h4)
	) name13385 (
		_w14967_,
		_w17171_,
		_w17432_
	);
	LUT2 #(
		.INIT('h1)
	) name13386 (
		_w17172_,
		_w17432_,
		_w17433_
	);
	LUT2 #(
		.INIT('h1)
	) name13387 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14838_,
		_w17434_
	);
	LUT2 #(
		.INIT('h2)
	) name13388 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w14842_,
		_w17435_
	);
	LUT2 #(
		.INIT('h4)
	) name13389 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14846_,
		_w17436_
	);
	LUT2 #(
		.INIT('h8)
	) name13390 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w14849_,
		_w17437_
	);
	LUT2 #(
		.INIT('h1)
	) name13391 (
		_w17436_,
		_w17437_,
		_w17438_
	);
	LUT2 #(
		.INIT('h4)
	) name13392 (
		_w17434_,
		_w17438_,
		_w17439_
	);
	LUT2 #(
		.INIT('h4)
	) name13393 (
		_w17435_,
		_w17439_,
		_w17440_
	);
	LUT2 #(
		.INIT('h2)
	) name13394 (
		_w14958_,
		_w17440_,
		_w17441_
	);
	LUT2 #(
		.INIT('h4)
	) name13395 (
		_w14958_,
		_w17440_,
		_w17442_
	);
	LUT2 #(
		.INIT('h2)
	) name13396 (
		\core_c_dec_MACop_E_reg/P0001 ,
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w17443_
	);
	LUT2 #(
		.INIT('h8)
	) name13397 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17443_,
		_w17444_
	);
	LUT2 #(
		.INIT('h4)
	) name13398 (
		_w12024_,
		_w17444_,
		_w17445_
	);
	LUT2 #(
		.INIT('h4)
	) name13399 (
		_w17442_,
		_w17445_,
		_w17446_
	);
	LUT2 #(
		.INIT('h1)
	) name13400 (
		_w17441_,
		_w17446_,
		_w17447_
	);
	LUT2 #(
		.INIT('h4)
	) name13401 (
		_w17433_,
		_w17447_,
		_w17448_
	);
	LUT2 #(
		.INIT('h1)
	) name13402 (
		_w17431_,
		_w17448_,
		_w17449_
	);
	LUT2 #(
		.INIT('h4)
	) name13403 (
		_w17162_,
		_w17166_,
		_w17450_
	);
	LUT2 #(
		.INIT('h1)
	) name13404 (
		_w17167_,
		_w17450_,
		_w17451_
	);
	LUT2 #(
		.INIT('h4)
	) name13405 (
		_w14852_,
		_w17172_,
		_w17452_
	);
	LUT2 #(
		.INIT('h1)
	) name13406 (
		_w17173_,
		_w17452_,
		_w17453_
	);
	LUT2 #(
		.INIT('h8)
	) name13407 (
		_w17451_,
		_w17453_,
		_w17454_
	);
	LUT2 #(
		.INIT('h1)
	) name13408 (
		_w17451_,
		_w17453_,
		_w17455_
	);
	LUT2 #(
		.INIT('h1)
	) name13409 (
		_w17454_,
		_w17455_,
		_w17456_
	);
	LUT2 #(
		.INIT('h8)
	) name13410 (
		_w17449_,
		_w17456_,
		_w17457_
	);
	LUT2 #(
		.INIT('h1)
	) name13411 (
		_w17450_,
		_w17452_,
		_w17458_
	);
	LUT2 #(
		.INIT('h1)
	) name13412 (
		_w17456_,
		_w17458_,
		_w17459_
	);
	LUT2 #(
		.INIT('h1)
	) name13413 (
		_w17457_,
		_w17459_,
		_w17460_
	);
	LUT2 #(
		.INIT('h4)
	) name13414 (
		_w17401_,
		_w17460_,
		_w17461_
	);
	LUT2 #(
		.INIT('h1)
	) name13415 (
		_w17399_,
		_w17461_,
		_w17462_
	);
	LUT2 #(
		.INIT('h4)
	) name13416 (
		_w17248_,
		_w17314_,
		_w17463_
	);
	LUT2 #(
		.INIT('h1)
	) name13417 (
		_w17315_,
		_w17463_,
		_w17464_
	);
	LUT2 #(
		.INIT('h1)
	) name13418 (
		_w17137_,
		_w17182_,
		_w17465_
	);
	LUT2 #(
		.INIT('h1)
	) name13419 (
		_w17183_,
		_w17465_,
		_w17466_
	);
	LUT2 #(
		.INIT('h2)
	) name13420 (
		_w17464_,
		_w17466_,
		_w17467_
	);
	LUT2 #(
		.INIT('h4)
	) name13421 (
		_w17464_,
		_w17466_,
		_w17468_
	);
	LUT2 #(
		.INIT('h1)
	) name13422 (
		_w17467_,
		_w17468_,
		_w17469_
	);
	LUT2 #(
		.INIT('h1)
	) name13423 (
		_w17462_,
		_w17469_,
		_w17470_
	);
	LUT2 #(
		.INIT('h1)
	) name13424 (
		_w17463_,
		_w17465_,
		_w17471_
	);
	LUT2 #(
		.INIT('h8)
	) name13425 (
		_w17469_,
		_w17471_,
		_w17472_
	);
	LUT2 #(
		.INIT('h1)
	) name13426 (
		_w17470_,
		_w17472_,
		_w17473_
	);
	LUT2 #(
		.INIT('h1)
	) name13427 (
		_w17337_,
		_w17473_,
		_w17474_
	);
	LUT2 #(
		.INIT('h8)
	) name13428 (
		_w17462_,
		_w17469_,
		_w17475_
	);
	LUT2 #(
		.INIT('h1)
	) name13429 (
		_w17470_,
		_w17475_,
		_w17476_
	);
	LUT2 #(
		.INIT('h1)
	) name13430 (
		_w17449_,
		_w17456_,
		_w17477_
	);
	LUT2 #(
		.INIT('h1)
	) name13431 (
		_w17457_,
		_w17477_,
		_w17478_
	);
	LUT2 #(
		.INIT('h1)
	) name13432 (
		_w14947_,
		_w15868_,
		_w17479_
	);
	LUT2 #(
		.INIT('h1)
	) name13433 (
		_w15869_,
		_w17479_,
		_w17480_
	);
	LUT2 #(
		.INIT('h1)
	) name13434 (
		_w17441_,
		_w17442_,
		_w17481_
	);
	LUT2 #(
		.INIT('h8)
	) name13435 (
		_w17445_,
		_w17481_,
		_w17482_
	);
	LUT2 #(
		.INIT('h1)
	) name13436 (
		_w17445_,
		_w17481_,
		_w17483_
	);
	LUT2 #(
		.INIT('h1)
	) name13437 (
		_w17482_,
		_w17483_,
		_w17484_
	);
	LUT2 #(
		.INIT('h2)
	) name13438 (
		_w17480_,
		_w17484_,
		_w17485_
	);
	LUT2 #(
		.INIT('h1)
	) name13439 (
		_w15839_,
		_w15848_,
		_w17486_
	);
	LUT2 #(
		.INIT('h1)
	) name13440 (
		_w15840_,
		_w17486_,
		_w17487_
	);
	LUT2 #(
		.INIT('h1)
	) name13441 (
		_w17416_,
		_w17425_,
		_w17488_
	);
	LUT2 #(
		.INIT('h2)
	) name13442 (
		_w17423_,
		_w17488_,
		_w17489_
	);
	LUT2 #(
		.INIT('h4)
	) name13443 (
		_w17423_,
		_w17488_,
		_w17490_
	);
	LUT2 #(
		.INIT('h1)
	) name13444 (
		_w17489_,
		_w17490_,
		_w17491_
	);
	LUT2 #(
		.INIT('h2)
	) name13445 (
		_w17487_,
		_w17491_,
		_w17492_
	);
	LUT2 #(
		.INIT('h1)
	) name13446 (
		_w17485_,
		_w17492_,
		_w17493_
	);
	LUT2 #(
		.INIT('h4)
	) name13447 (
		_w17426_,
		_w17430_,
		_w17494_
	);
	LUT2 #(
		.INIT('h1)
	) name13448 (
		_w17431_,
		_w17494_,
		_w17495_
	);
	LUT2 #(
		.INIT('h2)
	) name13449 (
		_w17433_,
		_w17447_,
		_w17496_
	);
	LUT2 #(
		.INIT('h1)
	) name13450 (
		_w17448_,
		_w17496_,
		_w17497_
	);
	LUT2 #(
		.INIT('h8)
	) name13451 (
		_w17495_,
		_w17497_,
		_w17498_
	);
	LUT2 #(
		.INIT('h1)
	) name13452 (
		_w17495_,
		_w17497_,
		_w17499_
	);
	LUT2 #(
		.INIT('h1)
	) name13453 (
		_w17498_,
		_w17499_,
		_w17500_
	);
	LUT2 #(
		.INIT('h8)
	) name13454 (
		_w17493_,
		_w17500_,
		_w17501_
	);
	LUT2 #(
		.INIT('h1)
	) name13455 (
		_w17494_,
		_w17496_,
		_w17502_
	);
	LUT2 #(
		.INIT('h1)
	) name13456 (
		_w17500_,
		_w17502_,
		_w17503_
	);
	LUT2 #(
		.INIT('h1)
	) name13457 (
		_w17501_,
		_w17503_,
		_w17504_
	);
	LUT2 #(
		.INIT('h4)
	) name13458 (
		_w17478_,
		_w17504_,
		_w17505_
	);
	LUT2 #(
		.INIT('h4)
	) name13459 (
		_w17387_,
		_w17394_,
		_w17506_
	);
	LUT2 #(
		.INIT('h1)
	) name13460 (
		_w17395_,
		_w17506_,
		_w17507_
	);
	LUT2 #(
		.INIT('h8)
	) name13461 (
		_w17343_,
		_w17350_,
		_w17508_
	);
	LUT2 #(
		.INIT('h1)
	) name13462 (
		_w17351_,
		_w17508_,
		_w17509_
	);
	LUT2 #(
		.INIT('h1)
	) name13463 (
		_w15781_,
		_w17509_,
		_w17510_
	);
	LUT2 #(
		.INIT('h1)
	) name13464 (
		_w15800_,
		_w15809_,
		_w17511_
	);
	LUT2 #(
		.INIT('h1)
	) name13465 (
		_w15801_,
		_w17511_,
		_w17512_
	);
	LUT2 #(
		.INIT('h1)
	) name13466 (
		_w17371_,
		_w17380_,
		_w17513_
	);
	LUT2 #(
		.INIT('h2)
	) name13467 (
		_w17378_,
		_w17513_,
		_w17514_
	);
	LUT2 #(
		.INIT('h4)
	) name13468 (
		_w17378_,
		_w17513_,
		_w17515_
	);
	LUT2 #(
		.INIT('h1)
	) name13469 (
		_w17514_,
		_w17515_,
		_w17516_
	);
	LUT2 #(
		.INIT('h2)
	) name13470 (
		_w17512_,
		_w17516_,
		_w17517_
	);
	LUT2 #(
		.INIT('h1)
	) name13471 (
		_w17510_,
		_w17517_,
		_w17518_
	);
	LUT2 #(
		.INIT('h4)
	) name13472 (
		_w17381_,
		_w17385_,
		_w17519_
	);
	LUT2 #(
		.INIT('h1)
	) name13473 (
		_w17386_,
		_w17519_,
		_w17520_
	);
	LUT2 #(
		.INIT('h8)
	) name13474 (
		_w17351_,
		_w17355_,
		_w17521_
	);
	LUT2 #(
		.INIT('h1)
	) name13475 (
		_w17356_,
		_w17521_,
		_w17522_
	);
	LUT2 #(
		.INIT('h8)
	) name13476 (
		_w17520_,
		_w17522_,
		_w17523_
	);
	LUT2 #(
		.INIT('h1)
	) name13477 (
		_w17520_,
		_w17522_,
		_w17524_
	);
	LUT2 #(
		.INIT('h1)
	) name13478 (
		_w17523_,
		_w17524_,
		_w17525_
	);
	LUT2 #(
		.INIT('h8)
	) name13479 (
		_w17518_,
		_w17525_,
		_w17526_
	);
	LUT2 #(
		.INIT('h1)
	) name13480 (
		_w17519_,
		_w17521_,
		_w17527_
	);
	LUT2 #(
		.INIT('h1)
	) name13481 (
		_w17525_,
		_w17527_,
		_w17528_
	);
	LUT2 #(
		.INIT('h1)
	) name13482 (
		_w17526_,
		_w17528_,
		_w17529_
	);
	LUT2 #(
		.INIT('h4)
	) name13483 (
		_w17507_,
		_w17529_,
		_w17530_
	);
	LUT2 #(
		.INIT('h1)
	) name13484 (
		_w17505_,
		_w17530_,
		_w17531_
	);
	LUT2 #(
		.INIT('h2)
	) name13485 (
		_w17401_,
		_w17460_,
		_w17532_
	);
	LUT2 #(
		.INIT('h1)
	) name13486 (
		_w17461_,
		_w17532_,
		_w17533_
	);
	LUT2 #(
		.INIT('h1)
	) name13487 (
		_w17339_,
		_w17398_,
		_w17534_
	);
	LUT2 #(
		.INIT('h1)
	) name13488 (
		_w17399_,
		_w17534_,
		_w17535_
	);
	LUT2 #(
		.INIT('h8)
	) name13489 (
		_w17533_,
		_w17535_,
		_w17536_
	);
	LUT2 #(
		.INIT('h1)
	) name13490 (
		_w17533_,
		_w17535_,
		_w17537_
	);
	LUT2 #(
		.INIT('h1)
	) name13491 (
		_w17536_,
		_w17537_,
		_w17538_
	);
	LUT2 #(
		.INIT('h8)
	) name13492 (
		_w17531_,
		_w17538_,
		_w17539_
	);
	LUT2 #(
		.INIT('h1)
	) name13493 (
		_w17532_,
		_w17534_,
		_w17540_
	);
	LUT2 #(
		.INIT('h1)
	) name13494 (
		_w17538_,
		_w17540_,
		_w17541_
	);
	LUT2 #(
		.INIT('h1)
	) name13495 (
		_w17539_,
		_w17541_,
		_w17542_
	);
	LUT2 #(
		.INIT('h8)
	) name13496 (
		_w17476_,
		_w17542_,
		_w17543_
	);
	LUT2 #(
		.INIT('h1)
	) name13497 (
		_w17474_,
		_w17543_,
		_w17544_
	);
	LUT2 #(
		.INIT('h1)
	) name13498 (
		_w17322_,
		_w17330_,
		_w17545_
	);
	LUT2 #(
		.INIT('h1)
	) name13499 (
		_w16860_,
		_w16926_,
		_w17546_
	);
	LUT2 #(
		.INIT('h1)
	) name13500 (
		_w16927_,
		_w17546_,
		_w17547_
	);
	LUT2 #(
		.INIT('h2)
	) name13501 (
		_w16963_,
		_w16965_,
		_w17548_
	);
	LUT2 #(
		.INIT('h1)
	) name13502 (
		_w16966_,
		_w17548_,
		_w17549_
	);
	LUT2 #(
		.INIT('h8)
	) name13503 (
		_w17547_,
		_w17549_,
		_w17550_
	);
	LUT2 #(
		.INIT('h1)
	) name13504 (
		_w17547_,
		_w17549_,
		_w17551_
	);
	LUT2 #(
		.INIT('h1)
	) name13505 (
		_w17550_,
		_w17551_,
		_w17552_
	);
	LUT2 #(
		.INIT('h1)
	) name13506 (
		_w17545_,
		_w17552_,
		_w17553_
	);
	LUT2 #(
		.INIT('h8)
	) name13507 (
		_w17545_,
		_w17552_,
		_w17554_
	);
	LUT2 #(
		.INIT('h1)
	) name13508 (
		_w17553_,
		_w17554_,
		_w17555_
	);
	LUT2 #(
		.INIT('h1)
	) name13509 (
		_w17323_,
		_w17329_,
		_w17556_
	);
	LUT2 #(
		.INIT('h1)
	) name13510 (
		_w17334_,
		_w17556_,
		_w17557_
	);
	LUT2 #(
		.INIT('h1)
	) name13511 (
		_w17336_,
		_w17557_,
		_w17558_
	);
	LUT2 #(
		.INIT('h4)
	) name13512 (
		_w17555_,
		_w17558_,
		_w17559_
	);
	LUT2 #(
		.INIT('h1)
	) name13513 (
		_w17546_,
		_w17548_,
		_w17560_
	);
	LUT2 #(
		.INIT('h1)
	) name13514 (
		_w17552_,
		_w17560_,
		_w17561_
	);
	LUT2 #(
		.INIT('h1)
	) name13515 (
		_w17554_,
		_w17561_,
		_w17562_
	);
	LUT2 #(
		.INIT('h2)
	) name13516 (
		_w16967_,
		_w16974_,
		_w17563_
	);
	LUT2 #(
		.INIT('h1)
	) name13517 (
		_w16975_,
		_w17563_,
		_w17564_
	);
	LUT2 #(
		.INIT('h8)
	) name13518 (
		_w17562_,
		_w17564_,
		_w17565_
	);
	LUT2 #(
		.INIT('h1)
	) name13519 (
		_w17559_,
		_w17565_,
		_w17566_
	);
	LUT2 #(
		.INIT('h8)
	) name13520 (
		_w17544_,
		_w17566_,
		_w17567_
	);
	LUT2 #(
		.INIT('h8)
	) name13521 (
		_w17098_,
		_w17567_,
		_w17568_
	);
	LUT2 #(
		.INIT('h1)
	) name13522 (
		_w17531_,
		_w17538_,
		_w17569_
	);
	LUT2 #(
		.INIT('h1)
	) name13523 (
		_w17539_,
		_w17569_,
		_w17570_
	);
	LUT2 #(
		.INIT('h1)
	) name13524 (
		_w17493_,
		_w17500_,
		_w17571_
	);
	LUT2 #(
		.INIT('h1)
	) name13525 (
		_w17501_,
		_w17571_,
		_w17572_
	);
	LUT2 #(
		.INIT('h1)
	) name13526 (
		_w15852_,
		_w15874_,
		_w17573_
	);
	LUT2 #(
		.INIT('h4)
	) name13527 (
		_w17487_,
		_w17491_,
		_w17574_
	);
	LUT2 #(
		.INIT('h1)
	) name13528 (
		_w17492_,
		_w17574_,
		_w17575_
	);
	LUT2 #(
		.INIT('h4)
	) name13529 (
		_w17480_,
		_w17484_,
		_w17576_
	);
	LUT2 #(
		.INIT('h1)
	) name13530 (
		_w17485_,
		_w17576_,
		_w17577_
	);
	LUT2 #(
		.INIT('h2)
	) name13531 (
		_w17575_,
		_w17577_,
		_w17578_
	);
	LUT2 #(
		.INIT('h4)
	) name13532 (
		_w17575_,
		_w17577_,
		_w17579_
	);
	LUT2 #(
		.INIT('h1)
	) name13533 (
		_w17578_,
		_w17579_,
		_w17580_
	);
	LUT2 #(
		.INIT('h1)
	) name13534 (
		_w17573_,
		_w17580_,
		_w17581_
	);
	LUT2 #(
		.INIT('h1)
	) name13535 (
		_w17574_,
		_w17576_,
		_w17582_
	);
	LUT2 #(
		.INIT('h8)
	) name13536 (
		_w17580_,
		_w17582_,
		_w17583_
	);
	LUT2 #(
		.INIT('h1)
	) name13537 (
		_w17581_,
		_w17583_,
		_w17584_
	);
	LUT2 #(
		.INIT('h1)
	) name13538 (
		_w17572_,
		_w17584_,
		_w17585_
	);
	LUT2 #(
		.INIT('h1)
	) name13539 (
		_w17518_,
		_w17525_,
		_w17586_
	);
	LUT2 #(
		.INIT('h1)
	) name13540 (
		_w17526_,
		_w17586_,
		_w17587_
	);
	LUT2 #(
		.INIT('h2)
	) name13541 (
		_w15783_,
		_w15814_,
		_w17588_
	);
	LUT2 #(
		.INIT('h4)
	) name13542 (
		_w17512_,
		_w17516_,
		_w17589_
	);
	LUT2 #(
		.INIT('h1)
	) name13543 (
		_w17517_,
		_w17589_,
		_w17590_
	);
	LUT2 #(
		.INIT('h8)
	) name13544 (
		_w15781_,
		_w17509_,
		_w17591_
	);
	LUT2 #(
		.INIT('h1)
	) name13545 (
		_w17510_,
		_w17591_,
		_w17592_
	);
	LUT2 #(
		.INIT('h2)
	) name13546 (
		_w17590_,
		_w17592_,
		_w17593_
	);
	LUT2 #(
		.INIT('h4)
	) name13547 (
		_w17590_,
		_w17592_,
		_w17594_
	);
	LUT2 #(
		.INIT('h1)
	) name13548 (
		_w17593_,
		_w17594_,
		_w17595_
	);
	LUT2 #(
		.INIT('h1)
	) name13549 (
		_w17588_,
		_w17595_,
		_w17596_
	);
	LUT2 #(
		.INIT('h1)
	) name13550 (
		_w17589_,
		_w17591_,
		_w17597_
	);
	LUT2 #(
		.INIT('h8)
	) name13551 (
		_w17595_,
		_w17597_,
		_w17598_
	);
	LUT2 #(
		.INIT('h1)
	) name13552 (
		_w17596_,
		_w17598_,
		_w17599_
	);
	LUT2 #(
		.INIT('h1)
	) name13553 (
		_w17587_,
		_w17599_,
		_w17600_
	);
	LUT2 #(
		.INIT('h1)
	) name13554 (
		_w17585_,
		_w17600_,
		_w17601_
	);
	LUT2 #(
		.INIT('h2)
	) name13555 (
		_w17478_,
		_w17504_,
		_w17602_
	);
	LUT2 #(
		.INIT('h1)
	) name13556 (
		_w17505_,
		_w17602_,
		_w17603_
	);
	LUT2 #(
		.INIT('h2)
	) name13557 (
		_w17507_,
		_w17529_,
		_w17604_
	);
	LUT2 #(
		.INIT('h1)
	) name13558 (
		_w17530_,
		_w17604_,
		_w17605_
	);
	LUT2 #(
		.INIT('h8)
	) name13559 (
		_w17603_,
		_w17605_,
		_w17606_
	);
	LUT2 #(
		.INIT('h1)
	) name13560 (
		_w17603_,
		_w17605_,
		_w17607_
	);
	LUT2 #(
		.INIT('h1)
	) name13561 (
		_w17606_,
		_w17607_,
		_w17608_
	);
	LUT2 #(
		.INIT('h8)
	) name13562 (
		_w17601_,
		_w17608_,
		_w17609_
	);
	LUT2 #(
		.INIT('h1)
	) name13563 (
		_w17602_,
		_w17604_,
		_w17610_
	);
	LUT2 #(
		.INIT('h1)
	) name13564 (
		_w17608_,
		_w17610_,
		_w17611_
	);
	LUT2 #(
		.INIT('h1)
	) name13565 (
		_w17609_,
		_w17611_,
		_w17612_
	);
	LUT2 #(
		.INIT('h4)
	) name13566 (
		_w17570_,
		_w17612_,
		_w17613_
	);
	LUT2 #(
		.INIT('h1)
	) name13567 (
		_w17601_,
		_w17608_,
		_w17614_
	);
	LUT2 #(
		.INIT('h1)
	) name13568 (
		_w17609_,
		_w17614_,
		_w17615_
	);
	LUT2 #(
		.INIT('h8)
	) name13569 (
		_w17573_,
		_w17580_,
		_w17616_
	);
	LUT2 #(
		.INIT('h1)
	) name13570 (
		_w17581_,
		_w17616_,
		_w17617_
	);
	LUT2 #(
		.INIT('h1)
	) name13571 (
		_w15853_,
		_w15875_,
		_w17618_
	);
	LUT2 #(
		.INIT('h4)
	) name13572 (
		_w15879_,
		_w17618_,
		_w17619_
	);
	LUT2 #(
		.INIT('h1)
	) name13573 (
		_w15880_,
		_w17619_,
		_w17620_
	);
	LUT2 #(
		.INIT('h2)
	) name13574 (
		_w17617_,
		_w17620_,
		_w17621_
	);
	LUT2 #(
		.INIT('h4)
	) name13575 (
		_w15783_,
		_w15813_,
		_w17622_
	);
	LUT2 #(
		.INIT('h8)
	) name13576 (
		_w17588_,
		_w17595_,
		_w17623_
	);
	LUT2 #(
		.INIT('h1)
	) name13577 (
		_w17596_,
		_w17622_,
		_w17624_
	);
	LUT2 #(
		.INIT('h4)
	) name13578 (
		_w17623_,
		_w17624_,
		_w17625_
	);
	LUT2 #(
		.INIT('h1)
	) name13579 (
		_w17621_,
		_w17625_,
		_w17626_
	);
	LUT2 #(
		.INIT('h8)
	) name13580 (
		_w17572_,
		_w17584_,
		_w17627_
	);
	LUT2 #(
		.INIT('h1)
	) name13581 (
		_w17585_,
		_w17627_,
		_w17628_
	);
	LUT2 #(
		.INIT('h8)
	) name13582 (
		_w17587_,
		_w17599_,
		_w17629_
	);
	LUT2 #(
		.INIT('h1)
	) name13583 (
		_w17600_,
		_w17629_,
		_w17630_
	);
	LUT2 #(
		.INIT('h2)
	) name13584 (
		_w17628_,
		_w17630_,
		_w17631_
	);
	LUT2 #(
		.INIT('h4)
	) name13585 (
		_w17628_,
		_w17630_,
		_w17632_
	);
	LUT2 #(
		.INIT('h1)
	) name13586 (
		_w17631_,
		_w17632_,
		_w17633_
	);
	LUT2 #(
		.INIT('h1)
	) name13587 (
		_w17626_,
		_w17633_,
		_w17634_
	);
	LUT2 #(
		.INIT('h1)
	) name13588 (
		_w17627_,
		_w17629_,
		_w17635_
	);
	LUT2 #(
		.INIT('h8)
	) name13589 (
		_w17633_,
		_w17635_,
		_w17636_
	);
	LUT2 #(
		.INIT('h1)
	) name13590 (
		_w17634_,
		_w17636_,
		_w17637_
	);
	LUT2 #(
		.INIT('h1)
	) name13591 (
		_w17615_,
		_w17637_,
		_w17638_
	);
	LUT2 #(
		.INIT('h1)
	) name13592 (
		_w17613_,
		_w17638_,
		_w17639_
	);
	LUT2 #(
		.INIT('h8)
	) name13593 (
		_w17626_,
		_w17633_,
		_w17640_
	);
	LUT2 #(
		.INIT('h1)
	) name13594 (
		_w17634_,
		_w17640_,
		_w17641_
	);
	LUT2 #(
		.INIT('h1)
	) name13595 (
		_w15819_,
		_w15886_,
		_w17642_
	);
	LUT2 #(
		.INIT('h4)
	) name13596 (
		_w17617_,
		_w17620_,
		_w17643_
	);
	LUT2 #(
		.INIT('h1)
	) name13597 (
		_w17621_,
		_w17643_,
		_w17644_
	);
	LUT2 #(
		.INIT('h4)
	) name13598 (
		_w17595_,
		_w17622_,
		_w17645_
	);
	LUT2 #(
		.INIT('h1)
	) name13599 (
		_w17625_,
		_w17645_,
		_w17646_
	);
	LUT2 #(
		.INIT('h8)
	) name13600 (
		_w17644_,
		_w17646_,
		_w17647_
	);
	LUT2 #(
		.INIT('h1)
	) name13601 (
		_w17644_,
		_w17646_,
		_w17648_
	);
	LUT2 #(
		.INIT('h1)
	) name13602 (
		_w17647_,
		_w17648_,
		_w17649_
	);
	LUT2 #(
		.INIT('h4)
	) name13603 (
		_w17642_,
		_w17649_,
		_w17650_
	);
	LUT2 #(
		.INIT('h1)
	) name13604 (
		_w17643_,
		_w17645_,
		_w17651_
	);
	LUT2 #(
		.INIT('h4)
	) name13605 (
		_w17649_,
		_w17651_,
		_w17652_
	);
	LUT2 #(
		.INIT('h1)
	) name13606 (
		_w17650_,
		_w17652_,
		_w17653_
	);
	LUT2 #(
		.INIT('h2)
	) name13607 (
		_w17641_,
		_w17653_,
		_w17654_
	);
	LUT2 #(
		.INIT('h2)
	) name13608 (
		_w17642_,
		_w17649_,
		_w17655_
	);
	LUT2 #(
		.INIT('h1)
	) name13609 (
		_w17650_,
		_w17655_,
		_w17656_
	);
	LUT2 #(
		.INIT('h1)
	) name13610 (
		_w15820_,
		_w15887_,
		_w17657_
	);
	LUT2 #(
		.INIT('h4)
	) name13611 (
		_w15891_,
		_w17657_,
		_w17658_
	);
	LUT2 #(
		.INIT('h1)
	) name13612 (
		_w15892_,
		_w17658_,
		_w17659_
	);
	LUT2 #(
		.INIT('h2)
	) name13613 (
		_w17656_,
		_w17659_,
		_w17660_
	);
	LUT2 #(
		.INIT('h1)
	) name13614 (
		_w17654_,
		_w17660_,
		_w17661_
	);
	LUT2 #(
		.INIT('h8)
	) name13615 (
		_w17639_,
		_w17661_,
		_w17662_
	);
	LUT2 #(
		.INIT('h8)
	) name13616 (
		_w17568_,
		_w17662_,
		_w17663_
	);
	LUT2 #(
		.INIT('h4)
	) name13617 (
		_w16363_,
		_w17663_,
		_w17664_
	);
	LUT2 #(
		.INIT('h8)
	) name13618 (
		_w17615_,
		_w17637_,
		_w17665_
	);
	LUT2 #(
		.INIT('h4)
	) name13619 (
		_w17613_,
		_w17665_,
		_w17666_
	);
	LUT2 #(
		.INIT('h4)
	) name13620 (
		_w17641_,
		_w17653_,
		_w17667_
	);
	LUT2 #(
		.INIT('h4)
	) name13621 (
		_w17656_,
		_w17659_,
		_w17668_
	);
	LUT2 #(
		.INIT('h1)
	) name13622 (
		_w17667_,
		_w17668_,
		_w17669_
	);
	LUT2 #(
		.INIT('h1)
	) name13623 (
		_w17654_,
		_w17669_,
		_w17670_
	);
	LUT2 #(
		.INIT('h8)
	) name13624 (
		_w17639_,
		_w17670_,
		_w17671_
	);
	LUT2 #(
		.INIT('h2)
	) name13625 (
		_w17570_,
		_w17612_,
		_w17672_
	);
	LUT2 #(
		.INIT('h1)
	) name13626 (
		_w17666_,
		_w17672_,
		_w17673_
	);
	LUT2 #(
		.INIT('h4)
	) name13627 (
		_w17671_,
		_w17673_,
		_w17674_
	);
	LUT2 #(
		.INIT('h2)
	) name13628 (
		_w17568_,
		_w17674_,
		_w17675_
	);
	LUT2 #(
		.INIT('h1)
	) name13629 (
		_w17476_,
		_w17542_,
		_w17676_
	);
	LUT2 #(
		.INIT('h8)
	) name13630 (
		_w17337_,
		_w17473_,
		_w17677_
	);
	LUT2 #(
		.INIT('h1)
	) name13631 (
		_w17676_,
		_w17677_,
		_w17678_
	);
	LUT2 #(
		.INIT('h1)
	) name13632 (
		_w17474_,
		_w17678_,
		_w17679_
	);
	LUT2 #(
		.INIT('h8)
	) name13633 (
		_w17566_,
		_w17679_,
		_w17680_
	);
	LUT2 #(
		.INIT('h1)
	) name13634 (
		_w17562_,
		_w17564_,
		_w17681_
	);
	LUT2 #(
		.INIT('h2)
	) name13635 (
		_w17555_,
		_w17558_,
		_w17682_
	);
	LUT2 #(
		.INIT('h4)
	) name13636 (
		_w17565_,
		_w17682_,
		_w17683_
	);
	LUT2 #(
		.INIT('h1)
	) name13637 (
		_w17681_,
		_w17683_,
		_w17684_
	);
	LUT2 #(
		.INIT('h4)
	) name13638 (
		_w17680_,
		_w17684_,
		_w17685_
	);
	LUT2 #(
		.INIT('h2)
	) name13639 (
		_w17098_,
		_w17685_,
		_w17686_
	);
	LUT2 #(
		.INIT('h1)
	) name13640 (
		_w16739_,
		_w16855_,
		_w17687_
	);
	LUT2 #(
		.INIT('h8)
	) name13641 (
		_w16858_,
		_w16978_,
		_w17688_
	);
	LUT2 #(
		.INIT('h4)
	) name13642 (
		_w16856_,
		_w17688_,
		_w17689_
	);
	LUT2 #(
		.INIT('h1)
	) name13643 (
		_w17687_,
		_w17689_,
		_w17690_
	);
	LUT2 #(
		.INIT('h1)
	) name13644 (
		_w17097_,
		_w17690_,
		_w17691_
	);
	LUT2 #(
		.INIT('h4)
	) name13645 (
		_w17088_,
		_w17091_,
		_w17692_
	);
	LUT2 #(
		.INIT('h1)
	) name13646 (
		_w17095_,
		_w17692_,
		_w17693_
	);
	LUT2 #(
		.INIT('h1)
	) name13647 (
		_w17079_,
		_w17693_,
		_w17694_
	);
	LUT2 #(
		.INIT('h1)
	) name13648 (
		_w17691_,
		_w17694_,
		_w17695_
	);
	LUT2 #(
		.INIT('h4)
	) name13649 (
		_w17675_,
		_w17695_,
		_w17696_
	);
	LUT2 #(
		.INIT('h4)
	) name13650 (
		_w17686_,
		_w17696_,
		_w17697_
	);
	LUT2 #(
		.INIT('h4)
	) name13651 (
		_w17664_,
		_w17697_,
		_w17698_
	);
	LUT2 #(
		.INIT('h1)
	) name13652 (
		_w17051_,
		_w17060_,
		_w17699_
	);
	LUT2 #(
		.INIT('h2)
	) name13653 (
		_w15253_,
		_w15272_,
		_w17700_
	);
	LUT2 #(
		.INIT('h1)
	) name13654 (
		_w15273_,
		_w17700_,
		_w17701_
	);
	LUT2 #(
		.INIT('h4)
	) name13655 (
		_w15288_,
		_w15291_,
		_w17702_
	);
	LUT2 #(
		.INIT('h1)
	) name13656 (
		_w15292_,
		_w17702_,
		_w17703_
	);
	LUT2 #(
		.INIT('h2)
	) name13657 (
		_w17701_,
		_w17703_,
		_w17704_
	);
	LUT2 #(
		.INIT('h4)
	) name13658 (
		_w17701_,
		_w17703_,
		_w17705_
	);
	LUT2 #(
		.INIT('h1)
	) name13659 (
		_w17704_,
		_w17705_,
		_w17706_
	);
	LUT2 #(
		.INIT('h1)
	) name13660 (
		_w17699_,
		_w17706_,
		_w17707_
	);
	LUT2 #(
		.INIT('h8)
	) name13661 (
		_w17699_,
		_w17706_,
		_w17708_
	);
	LUT2 #(
		.INIT('h1)
	) name13662 (
		_w17707_,
		_w17708_,
		_w17709_
	);
	LUT2 #(
		.INIT('h1)
	) name13663 (
		_w17050_,
		_w17059_,
		_w17710_
	);
	LUT2 #(
		.INIT('h4)
	) name13664 (
		_w17064_,
		_w17710_,
		_w17711_
	);
	LUT2 #(
		.INIT('h1)
	) name13665 (
		_w17066_,
		_w17711_,
		_w17712_
	);
	LUT2 #(
		.INIT('h2)
	) name13666 (
		_w17709_,
		_w17712_,
		_w17713_
	);
	LUT2 #(
		.INIT('h1)
	) name13667 (
		_w14853_,
		_w17713_,
		_w17714_
	);
	LUT2 #(
		.INIT('h2)
	) name13668 (
		_w15293_,
		_w15300_,
		_w17715_
	);
	LUT2 #(
		.INIT('h1)
	) name13669 (
		_w15301_,
		_w17715_,
		_w17716_
	);
	LUT2 #(
		.INIT('h1)
	) name13670 (
		_w17700_,
		_w17702_,
		_w17717_
	);
	LUT2 #(
		.INIT('h8)
	) name13671 (
		_w17706_,
		_w17717_,
		_w17718_
	);
	LUT2 #(
		.INIT('h1)
	) name13672 (
		_w17707_,
		_w17718_,
		_w17719_
	);
	LUT2 #(
		.INIT('h4)
	) name13673 (
		_w17716_,
		_w17719_,
		_w17720_
	);
	LUT2 #(
		.INIT('h2)
	) name13674 (
		_w17716_,
		_w17719_,
		_w17721_
	);
	LUT2 #(
		.INIT('h1)
	) name13675 (
		_w17720_,
		_w17721_,
		_w17722_
	);
	LUT2 #(
		.INIT('h8)
	) name13676 (
		_w14853_,
		_w17722_,
		_w17723_
	);
	LUT2 #(
		.INIT('h1)
	) name13677 (
		_w14853_,
		_w17722_,
		_w17724_
	);
	LUT2 #(
		.INIT('h1)
	) name13678 (
		_w17723_,
		_w17724_,
		_w17725_
	);
	LUT2 #(
		.INIT('h1)
	) name13679 (
		_w17714_,
		_w17725_,
		_w17726_
	);
	LUT2 #(
		.INIT('h8)
	) name13680 (
		_w17714_,
		_w17722_,
		_w17727_
	);
	LUT2 #(
		.INIT('h1)
	) name13681 (
		_w17726_,
		_w17727_,
		_w17728_
	);
	LUT2 #(
		.INIT('h1)
	) name13682 (
		_w14853_,
		_w17071_,
		_w17729_
	);
	LUT2 #(
		.INIT('h4)
	) name13683 (
		_w17709_,
		_w17712_,
		_w17730_
	);
	LUT2 #(
		.INIT('h1)
	) name13684 (
		_w17713_,
		_w17730_,
		_w17731_
	);
	LUT2 #(
		.INIT('h8)
	) name13685 (
		_w14853_,
		_w17731_,
		_w17732_
	);
	LUT2 #(
		.INIT('h1)
	) name13686 (
		_w14853_,
		_w17731_,
		_w17733_
	);
	LUT2 #(
		.INIT('h1)
	) name13687 (
		_w17732_,
		_w17733_,
		_w17734_
	);
	LUT2 #(
		.INIT('h1)
	) name13688 (
		_w17729_,
		_w17734_,
		_w17735_
	);
	LUT2 #(
		.INIT('h8)
	) name13689 (
		_w17729_,
		_w17731_,
		_w17736_
	);
	LUT2 #(
		.INIT('h1)
	) name13690 (
		_w17735_,
		_w17736_,
		_w17737_
	);
	LUT2 #(
		.INIT('h1)
	) name13691 (
		_w17728_,
		_w17737_,
		_w17738_
	);
	LUT2 #(
		.INIT('h4)
	) name13692 (
		_w17730_,
		_w17734_,
		_w17739_
	);
	LUT2 #(
		.INIT('h1)
	) name13693 (
		_w17735_,
		_w17739_,
		_w17740_
	);
	LUT2 #(
		.INIT('h2)
	) name13694 (
		_w17728_,
		_w17740_,
		_w17741_
	);
	LUT2 #(
		.INIT('h4)
	) name13695 (
		_w17072_,
		_w17076_,
		_w17742_
	);
	LUT2 #(
		.INIT('h1)
	) name13696 (
		_w17077_,
		_w17742_,
		_w17743_
	);
	LUT2 #(
		.INIT('h4)
	) name13697 (
		_w17741_,
		_w17743_,
		_w17744_
	);
	LUT2 #(
		.INIT('h1)
	) name13698 (
		_w17738_,
		_w17744_,
		_w17745_
	);
	LUT2 #(
		.INIT('h8)
	) name13699 (
		_w15306_,
		_w15308_,
		_w17746_
	);
	LUT2 #(
		.INIT('h1)
	) name13700 (
		_w15312_,
		_w17746_,
		_w17747_
	);
	LUT2 #(
		.INIT('h4)
	) name13701 (
		_w17720_,
		_w17725_,
		_w17748_
	);
	LUT2 #(
		.INIT('h1)
	) name13702 (
		_w17726_,
		_w17748_,
		_w17749_
	);
	LUT2 #(
		.INIT('h1)
	) name13703 (
		_w14853_,
		_w17721_,
		_w17750_
	);
	LUT2 #(
		.INIT('h4)
	) name13704 (
		_w15249_,
		_w15304_,
		_w17751_
	);
	LUT2 #(
		.INIT('h1)
	) name13705 (
		_w15305_,
		_w17751_,
		_w17752_
	);
	LUT2 #(
		.INIT('h8)
	) name13706 (
		_w14853_,
		_w17752_,
		_w17753_
	);
	LUT2 #(
		.INIT('h1)
	) name13707 (
		_w14853_,
		_w17752_,
		_w17754_
	);
	LUT2 #(
		.INIT('h1)
	) name13708 (
		_w17753_,
		_w17754_,
		_w17755_
	);
	LUT2 #(
		.INIT('h1)
	) name13709 (
		_w17750_,
		_w17755_,
		_w17756_
	);
	LUT2 #(
		.INIT('h8)
	) name13710 (
		_w17750_,
		_w17752_,
		_w17757_
	);
	LUT2 #(
		.INIT('h1)
	) name13711 (
		_w17756_,
		_w17757_,
		_w17758_
	);
	LUT2 #(
		.INIT('h4)
	) name13712 (
		_w17749_,
		_w17758_,
		_w17759_
	);
	LUT2 #(
		.INIT('h1)
	) name13713 (
		_w17747_,
		_w17759_,
		_w17760_
	);
	LUT2 #(
		.INIT('h4)
	) name13714 (
		_w17751_,
		_w17755_,
		_w17761_
	);
	LUT2 #(
		.INIT('h1)
	) name13715 (
		_w17756_,
		_w17761_,
		_w17762_
	);
	LUT2 #(
		.INIT('h8)
	) name13716 (
		_w17749_,
		_w17762_,
		_w17763_
	);
	LUT2 #(
		.INIT('h1)
	) name13717 (
		_w17760_,
		_w17763_,
		_w17764_
	);
	LUT2 #(
		.INIT('h1)
	) name13718 (
		_w17745_,
		_w17764_,
		_w17765_
	);
	LUT2 #(
		.INIT('h4)
	) name13719 (
		_w17698_,
		_w17765_,
		_w17766_
	);
	LUT2 #(
		.INIT('h2)
	) name13720 (
		_w17747_,
		_w17762_,
		_w17767_
	);
	LUT2 #(
		.INIT('h2)
	) name13721 (
		_w17749_,
		_w17758_,
		_w17768_
	);
	LUT2 #(
		.INIT('h4)
	) name13722 (
		_w17767_,
		_w17768_,
		_w17769_
	);
	LUT2 #(
		.INIT('h4)
	) name13723 (
		_w17728_,
		_w17740_,
		_w17770_
	);
	LUT2 #(
		.INIT('h8)
	) name13724 (
		_w17738_,
		_w17743_,
		_w17771_
	);
	LUT2 #(
		.INIT('h1)
	) name13725 (
		_w17770_,
		_w17771_,
		_w17772_
	);
	LUT2 #(
		.INIT('h1)
	) name13726 (
		_w17764_,
		_w17772_,
		_w17773_
	);
	LUT2 #(
		.INIT('h4)
	) name13727 (
		_w17747_,
		_w17762_,
		_w17774_
	);
	LUT2 #(
		.INIT('h1)
	) name13728 (
		_w17769_,
		_w17774_,
		_w17775_
	);
	LUT2 #(
		.INIT('h4)
	) name13729 (
		_w17773_,
		_w17775_,
		_w17776_
	);
	LUT2 #(
		.INIT('h4)
	) name13730 (
		_w17766_,
		_w17776_,
		_w17777_
	);
	LUT2 #(
		.INIT('h4)
	) name13731 (
		_w15314_,
		_w17777_,
		_w17778_
	);
	LUT2 #(
		.INIT('h1)
	) name13732 (
		_w15244_,
		_w17778_,
		_w17779_
	);
	LUT2 #(
		.INIT('h4)
	) name13733 (
		_w15319_,
		_w17779_,
		_w17780_
	);
	LUT2 #(
		.INIT('h4)
	) name13734 (
		_w15246_,
		_w15316_,
		_w17781_
	);
	LUT2 #(
		.INIT('h8)
	) name13735 (
		_w15247_,
		_w15314_,
		_w17782_
	);
	LUT2 #(
		.INIT('h1)
	) name13736 (
		_w17781_,
		_w17782_,
		_w17783_
	);
	LUT2 #(
		.INIT('h4)
	) name13737 (
		_w17780_,
		_w17783_,
		_w17784_
	);
	LUT2 #(
		.INIT('h1)
	) name13738 (
		_w15183_,
		_w17784_,
		_w17785_
	);
	LUT2 #(
		.INIT('h1)
	) name13739 (
		_w15182_,
		_w17785_,
		_w17786_
	);
	LUT2 #(
		.INIT('h2)
	) name13740 (
		_w15122_,
		_w17786_,
		_w17787_
	);
	LUT2 #(
		.INIT('h4)
	) name13741 (
		_w15122_,
		_w17786_,
		_w17788_
	);
	LUT2 #(
		.INIT('h1)
	) name13742 (
		_w17787_,
		_w17788_,
		_w17789_
	);
	LUT2 #(
		.INIT('h2)
	) name13743 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17789_,
		_w17790_
	);
	LUT2 #(
		.INIT('h1)
	) name13744 (
		_w15182_,
		_w15183_,
		_w17791_
	);
	LUT2 #(
		.INIT('h8)
	) name13745 (
		_w17784_,
		_w17791_,
		_w17792_
	);
	LUT2 #(
		.INIT('h1)
	) name13746 (
		_w17784_,
		_w17791_,
		_w17793_
	);
	LUT2 #(
		.INIT('h1)
	) name13747 (
		_w17792_,
		_w17793_,
		_w17794_
	);
	LUT2 #(
		.INIT('h4)
	) name13748 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17794_,
		_w17795_
	);
	LUT2 #(
		.INIT('h1)
	) name13749 (
		_w17790_,
		_w17795_,
		_w17796_
	);
	LUT2 #(
		.INIT('h2)
	) name13750 (
		_w14752_,
		_w17796_,
		_w17797_
	);
	LUT2 #(
		.INIT('h4)
	) name13751 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w5951_,
		_w17798_
	);
	LUT2 #(
		.INIT('h8)
	) name13752 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		_w17798_,
		_w17799_
	);
	LUT2 #(
		.INIT('h1)
	) name13753 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 ,
		_w17799_,
		_w17800_
	);
	LUT2 #(
		.INIT('h4)
	) name13754 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR2_E_reg/P0001 ,
		_w17801_
	);
	LUT2 #(
		.INIT('h4)
	) name13755 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w17802_
	);
	LUT2 #(
		.INIT('h2)
	) name13756 (
		\core_c_dec_satMR_E_reg/P0001 ,
		_w4174_,
		_w17803_
	);
	LUT2 #(
		.INIT('h4)
	) name13757 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w17803_,
		_w17804_
	);
	LUT2 #(
		.INIT('h1)
	) name13758 (
		_w17802_,
		_w17804_,
		_w17805_
	);
	LUT2 #(
		.INIT('h4)
	) name13759 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w17805_,
		_w17806_
	);
	LUT2 #(
		.INIT('h4)
	) name13760 (
		_w17801_,
		_w17806_,
		_w17807_
	);
	LUT2 #(
		.INIT('h1)
	) name13761 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w17807_,
		_w17808_
	);
	LUT2 #(
		.INIT('h2)
	) name13762 (
		_w13801_,
		_w17805_,
		_w17809_
	);
	LUT2 #(
		.INIT('h1)
	) name13763 (
		_w17799_,
		_w17809_,
		_w17810_
	);
	LUT2 #(
		.INIT('h2)
	) name13764 (
		_w17808_,
		_w17810_,
		_w17811_
	);
	LUT2 #(
		.INIT('h1)
	) name13765 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8715_,
		_w17812_
	);
	LUT2 #(
		.INIT('h2)
	) name13766 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12836_,
		_w17813_
	);
	LUT2 #(
		.INIT('h1)
	) name13767 (
		_w17812_,
		_w17813_,
		_w17814_
	);
	LUT2 #(
		.INIT('h4)
	) name13768 (
		_w17809_,
		_w17814_,
		_w17815_
	);
	LUT2 #(
		.INIT('h2)
	) name13769 (
		_w17811_,
		_w17815_,
		_w17816_
	);
	LUT2 #(
		.INIT('h1)
	) name13770 (
		_w17800_,
		_w17816_,
		_w17817_
	);
	LUT2 #(
		.INIT('h1)
	) name13771 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12743_,
		_w17818_
	);
	LUT2 #(
		.INIT('h2)
	) name13772 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12771_,
		_w17819_
	);
	LUT2 #(
		.INIT('h1)
	) name13773 (
		_w17818_,
		_w17819_,
		_w17820_
	);
	LUT2 #(
		.INIT('h2)
	) name13774 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w17803_,
		_w17821_
	);
	LUT2 #(
		.INIT('h8)
	) name13775 (
		_w17820_,
		_w17821_,
		_w17822_
	);
	LUT2 #(
		.INIT('h8)
	) name13776 (
		_w17798_,
		_w17822_,
		_w17823_
	);
	LUT2 #(
		.INIT('h1)
	) name13777 (
		_w17817_,
		_w17823_,
		_w17824_
	);
	LUT2 #(
		.INIT('h1)
	) name13778 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[2]/P0001 ,
		_w17808_,
		_w17825_
	);
	LUT2 #(
		.INIT('h1)
	) name13779 (
		_w17824_,
		_w17825_,
		_w17826_
	);
	LUT2 #(
		.INIT('h8)
	) name13780 (
		_w17798_,
		_w17803_,
		_w17827_
	);
	LUT2 #(
		.INIT('h8)
	) name13781 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		_w17827_,
		_w17828_
	);
	LUT2 #(
		.INIT('h1)
	) name13782 (
		_w14752_,
		_w17828_,
		_w17829_
	);
	LUT2 #(
		.INIT('h4)
	) name13783 (
		_w17826_,
		_w17829_,
		_w17830_
	);
	LUT2 #(
		.INIT('h1)
	) name13784 (
		_w17797_,
		_w17830_,
		_w17831_
	);
	LUT2 #(
		.INIT('h1)
	) name13785 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		\core_c_dec_updSR_E_reg/P0001 ,
		_w17832_
	);
	LUT2 #(
		.INIT('h2)
	) name13786 (
		_w13804_,
		_w17832_,
		_w17833_
	);
	LUT2 #(
		.INIT('h1)
	) name13787 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7340_,
		_w17834_
	);
	LUT2 #(
		.INIT('h2)
	) name13788 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12658_,
		_w17835_
	);
	LUT2 #(
		.INIT('h1)
	) name13789 (
		_w17834_,
		_w17835_,
		_w17836_
	);
	LUT2 #(
		.INIT('h2)
	) name13790 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w17836_,
		_w17837_
	);
	LUT2 #(
		.INIT('h8)
	) name13791 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w17838_
	);
	LUT2 #(
		.INIT('h2)
	) name13792 (
		\core_c_dec_SHTop_E_reg/P0001 ,
		_w17838_,
		_w17839_
	);
	LUT2 #(
		.INIT('h4)
	) name13793 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w17840_
	);
	LUT2 #(
		.INIT('h8)
	) name13794 (
		_w7373_,
		_w9272_,
		_w17841_
	);
	LUT2 #(
		.INIT('h1)
	) name13795 (
		_w7373_,
		_w9272_,
		_w17842_
	);
	LUT2 #(
		.INIT('h1)
	) name13796 (
		_w17841_,
		_w17842_,
		_w17843_
	);
	LUT2 #(
		.INIT('h2)
	) name13797 (
		_w17840_,
		_w17843_,
		_w17844_
	);
	LUT2 #(
		.INIT('h8)
	) name13798 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w17845_
	);
	LUT2 #(
		.INIT('h1)
	) name13799 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w9272_,
		_w17846_
	);
	LUT2 #(
		.INIT('h1)
	) name13800 (
		_w17840_,
		_w17845_,
		_w17847_
	);
	LUT2 #(
		.INIT('h4)
	) name13801 (
		_w17846_,
		_w17847_,
		_w17848_
	);
	LUT2 #(
		.INIT('h1)
	) name13802 (
		_w17844_,
		_w17848_,
		_w17849_
	);
	LUT2 #(
		.INIT('h8)
	) name13803 (
		_w17839_,
		_w17849_,
		_w17850_
	);
	LUT2 #(
		.INIT('h8)
	) name13804 (
		_w8501_,
		_w17841_,
		_w17851_
	);
	LUT2 #(
		.INIT('h1)
	) name13805 (
		_w7995_,
		_w17851_,
		_w17852_
	);
	LUT2 #(
		.INIT('h8)
	) name13806 (
		_w7995_,
		_w17851_,
		_w17853_
	);
	LUT2 #(
		.INIT('h1)
	) name13807 (
		_w17852_,
		_w17853_,
		_w17854_
	);
	LUT2 #(
		.INIT('h2)
	) name13808 (
		_w17840_,
		_w17854_,
		_w17855_
	);
	LUT2 #(
		.INIT('h8)
	) name13809 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w17856_
	);
	LUT2 #(
		.INIT('h1)
	) name13810 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w7995_,
		_w17857_
	);
	LUT2 #(
		.INIT('h1)
	) name13811 (
		_w17840_,
		_w17856_,
		_w17858_
	);
	LUT2 #(
		.INIT('h4)
	) name13812 (
		_w17857_,
		_w17858_,
		_w17859_
	);
	LUT2 #(
		.INIT('h1)
	) name13813 (
		_w17855_,
		_w17859_,
		_w17860_
	);
	LUT2 #(
		.INIT('h8)
	) name13814 (
		_w17839_,
		_w17860_,
		_w17861_
	);
	LUT2 #(
		.INIT('h1)
	) name13815 (
		_w17850_,
		_w17861_,
		_w17862_
	);
	LUT2 #(
		.INIT('h8)
	) name13816 (
		_w9939_,
		_w17853_,
		_w17863_
	);
	LUT2 #(
		.INIT('h1)
	) name13817 (
		_w9939_,
		_w17853_,
		_w17864_
	);
	LUT2 #(
		.INIT('h1)
	) name13818 (
		_w17863_,
		_w17864_,
		_w17865_
	);
	LUT2 #(
		.INIT('h2)
	) name13819 (
		_w17840_,
		_w17865_,
		_w17866_
	);
	LUT2 #(
		.INIT('h8)
	) name13820 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w17867_
	);
	LUT2 #(
		.INIT('h1)
	) name13821 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w9939_,
		_w17868_
	);
	LUT2 #(
		.INIT('h1)
	) name13822 (
		_w17840_,
		_w17867_,
		_w17869_
	);
	LUT2 #(
		.INIT('h4)
	) name13823 (
		_w17868_,
		_w17869_,
		_w17870_
	);
	LUT2 #(
		.INIT('h1)
	) name13824 (
		_w17866_,
		_w17870_,
		_w17871_
	);
	LUT2 #(
		.INIT('h8)
	) name13825 (
		_w17839_,
		_w17871_,
		_w17872_
	);
	LUT2 #(
		.INIT('h1)
	) name13826 (
		_w8501_,
		_w17841_,
		_w17873_
	);
	LUT2 #(
		.INIT('h1)
	) name13827 (
		_w17851_,
		_w17873_,
		_w17874_
	);
	LUT2 #(
		.INIT('h2)
	) name13828 (
		_w17840_,
		_w17874_,
		_w17875_
	);
	LUT2 #(
		.INIT('h8)
	) name13829 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w17876_
	);
	LUT2 #(
		.INIT('h1)
	) name13830 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w8501_,
		_w17877_
	);
	LUT2 #(
		.INIT('h1)
	) name13831 (
		_w17840_,
		_w17876_,
		_w17878_
	);
	LUT2 #(
		.INIT('h4)
	) name13832 (
		_w17877_,
		_w17878_,
		_w17879_
	);
	LUT2 #(
		.INIT('h1)
	) name13833 (
		_w17875_,
		_w17879_,
		_w17880_
	);
	LUT2 #(
		.INIT('h8)
	) name13834 (
		_w17839_,
		_w17880_,
		_w17881_
	);
	LUT2 #(
		.INIT('h1)
	) name13835 (
		_w17872_,
		_w17881_,
		_w17882_
	);
	LUT2 #(
		.INIT('h8)
	) name13836 (
		_w17862_,
		_w17882_,
		_w17883_
	);
	LUT2 #(
		.INIT('h8)
	) name13837 (
		_w10789_,
		_w17863_,
		_w17884_
	);
	LUT2 #(
		.INIT('h8)
	) name13838 (
		_w11303_,
		_w17884_,
		_w17885_
	);
	LUT2 #(
		.INIT('h1)
	) name13839 (
		_w11303_,
		_w17884_,
		_w17886_
	);
	LUT2 #(
		.INIT('h1)
	) name13840 (
		_w17885_,
		_w17886_,
		_w17887_
	);
	LUT2 #(
		.INIT('h2)
	) name13841 (
		_w17840_,
		_w17887_,
		_w17888_
	);
	LUT2 #(
		.INIT('h8)
	) name13842 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w17889_
	);
	LUT2 #(
		.INIT('h1)
	) name13843 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w11303_,
		_w17890_
	);
	LUT2 #(
		.INIT('h1)
	) name13844 (
		_w17840_,
		_w17889_,
		_w17891_
	);
	LUT2 #(
		.INIT('h4)
	) name13845 (
		_w17890_,
		_w17891_,
		_w17892_
	);
	LUT2 #(
		.INIT('h1)
	) name13846 (
		_w17888_,
		_w17892_,
		_w17893_
	);
	LUT2 #(
		.INIT('h8)
	) name13847 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w17894_
	);
	LUT2 #(
		.INIT('h1)
	) name13848 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w7172_,
		_w17895_
	);
	LUT2 #(
		.INIT('h1)
	) name13849 (
		_w17840_,
		_w17894_,
		_w17896_
	);
	LUT2 #(
		.INIT('h4)
	) name13850 (
		_w17895_,
		_w17896_,
		_w17897_
	);
	LUT2 #(
		.INIT('h4)
	) name13851 (
		_w7172_,
		_w17885_,
		_w17898_
	);
	LUT2 #(
		.INIT('h2)
	) name13852 (
		_w7172_,
		_w17885_,
		_w17899_
	);
	LUT2 #(
		.INIT('h2)
	) name13853 (
		_w17840_,
		_w17898_,
		_w17900_
	);
	LUT2 #(
		.INIT('h4)
	) name13854 (
		_w17899_,
		_w17900_,
		_w17901_
	);
	LUT2 #(
		.INIT('h1)
	) name13855 (
		_w17897_,
		_w17901_,
		_w17902_
	);
	LUT2 #(
		.INIT('h1)
	) name13856 (
		_w17893_,
		_w17902_,
		_w17903_
	);
	LUT2 #(
		.INIT('h1)
	) name13857 (
		_w10789_,
		_w17863_,
		_w17904_
	);
	LUT2 #(
		.INIT('h1)
	) name13858 (
		_w17884_,
		_w17904_,
		_w17905_
	);
	LUT2 #(
		.INIT('h2)
	) name13859 (
		_w17840_,
		_w17905_,
		_w17906_
	);
	LUT2 #(
		.INIT('h8)
	) name13860 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w17907_
	);
	LUT2 #(
		.INIT('h1)
	) name13861 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w10789_,
		_w17908_
	);
	LUT2 #(
		.INIT('h1)
	) name13862 (
		_w17840_,
		_w17907_,
		_w17909_
	);
	LUT2 #(
		.INIT('h4)
	) name13863 (
		_w17908_,
		_w17909_,
		_w17910_
	);
	LUT2 #(
		.INIT('h1)
	) name13864 (
		_w17906_,
		_w17910_,
		_w17911_
	);
	LUT2 #(
		.INIT('h1)
	) name13865 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w17911_,
		_w17912_
	);
	LUT2 #(
		.INIT('h8)
	) name13866 (
		_w17903_,
		_w17912_,
		_w17913_
	);
	LUT2 #(
		.INIT('h2)
	) name13867 (
		_w17839_,
		_w17913_,
		_w17914_
	);
	LUT2 #(
		.INIT('h2)
	) name13868 (
		_w17883_,
		_w17914_,
		_w17915_
	);
	LUT2 #(
		.INIT('h2)
	) name13869 (
		_w17872_,
		_w17880_,
		_w17916_
	);
	LUT2 #(
		.INIT('h8)
	) name13870 (
		_w17862_,
		_w17916_,
		_w17917_
	);
	LUT2 #(
		.INIT('h8)
	) name13871 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w17839_,
		_w17918_
	);
	LUT2 #(
		.INIT('h4)
	) name13872 (
		_w17911_,
		_w17918_,
		_w17919_
	);
	LUT2 #(
		.INIT('h8)
	) name13873 (
		_w17903_,
		_w17919_,
		_w17920_
	);
	LUT2 #(
		.INIT('h8)
	) name13874 (
		_w17917_,
		_w17920_,
		_w17921_
	);
	LUT2 #(
		.INIT('h1)
	) name13875 (
		_w17915_,
		_w17921_,
		_w17922_
	);
	LUT2 #(
		.INIT('h4)
	) name13876 (
		_w7160_,
		_w13832_,
		_w17923_
	);
	LUT2 #(
		.INIT('h2)
	) name13877 (
		_w14444_,
		_w17923_,
		_w17924_
	);
	LUT2 #(
		.INIT('h2)
	) name13878 (
		_w17839_,
		_w17924_,
		_w17925_
	);
	LUT2 #(
		.INIT('h2)
	) name13879 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w17840_,
		_w17926_
	);
	LUT2 #(
		.INIT('h2)
	) name13880 (
		_w7373_,
		_w17926_,
		_w17927_
	);
	LUT2 #(
		.INIT('h4)
	) name13881 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w17926_,
		_w17928_
	);
	LUT2 #(
		.INIT('h1)
	) name13882 (
		_w17927_,
		_w17928_,
		_w17929_
	);
	LUT2 #(
		.INIT('h2)
	) name13883 (
		_w17925_,
		_w17929_,
		_w17930_
	);
	LUT2 #(
		.INIT('h8)
	) name13884 (
		_w17839_,
		_w17929_,
		_w17931_
	);
	LUT2 #(
		.INIT('h4)
	) name13885 (
		_w9124_,
		_w13832_,
		_w17932_
	);
	LUT2 #(
		.INIT('h2)
	) name13886 (
		_w14377_,
		_w17932_,
		_w17933_
	);
	LUT2 #(
		.INIT('h2)
	) name13887 (
		_w17931_,
		_w17933_,
		_w17934_
	);
	LUT2 #(
		.INIT('h1)
	) name13888 (
		_w17930_,
		_w17934_,
		_w17935_
	);
	LUT2 #(
		.INIT('h1)
	) name13889 (
		_w17922_,
		_w17935_,
		_w17936_
	);
	LUT2 #(
		.INIT('h4)
	) name13890 (
		_w11996_,
		_w13832_,
		_w17937_
	);
	LUT2 #(
		.INIT('h2)
	) name13891 (
		_w13831_,
		_w17937_,
		_w17938_
	);
	LUT2 #(
		.INIT('h2)
	) name13892 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w17939_
	);
	LUT2 #(
		.INIT('h4)
	) name13893 (
		_w17938_,
		_w17939_,
		_w17940_
	);
	LUT2 #(
		.INIT('h4)
	) name13894 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w17941_
	);
	LUT2 #(
		.INIT('h8)
	) name13895 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w17941_,
		_w17942_
	);
	LUT2 #(
		.INIT('h8)
	) name13896 (
		_w17840_,
		_w17942_,
		_w17943_
	);
	LUT2 #(
		.INIT('h1)
	) name13897 (
		_w17940_,
		_w17943_,
		_w17944_
	);
	LUT2 #(
		.INIT('h2)
	) name13898 (
		_w17839_,
		_w17944_,
		_w17945_
	);
	LUT2 #(
		.INIT('h8)
	) name13899 (
		_w17893_,
		_w17911_,
		_w17946_
	);
	LUT2 #(
		.INIT('h8)
	) name13900 (
		_w17839_,
		_w17902_,
		_w17947_
	);
	LUT2 #(
		.INIT('h8)
	) name13901 (
		_w17946_,
		_w17947_,
		_w17948_
	);
	LUT2 #(
		.INIT('h4)
	) name13902 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w17948_,
		_w17949_
	);
	LUT2 #(
		.INIT('h8)
	) name13903 (
		_w17871_,
		_w17881_,
		_w17950_
	);
	LUT2 #(
		.INIT('h8)
	) name13904 (
		_w17862_,
		_w17950_,
		_w17951_
	);
	LUT2 #(
		.INIT('h8)
	) name13905 (
		_w17949_,
		_w17951_,
		_w17952_
	);
	LUT2 #(
		.INIT('h2)
	) name13906 (
		_w17850_,
		_w17860_,
		_w17953_
	);
	LUT2 #(
		.INIT('h8)
	) name13907 (
		_w17882_,
		_w17953_,
		_w17954_
	);
	LUT2 #(
		.INIT('h8)
	) name13908 (
		_w17920_,
		_w17954_,
		_w17955_
	);
	LUT2 #(
		.INIT('h4)
	) name13909 (
		_w17931_,
		_w17955_,
		_w17956_
	);
	LUT2 #(
		.INIT('h8)
	) name13910 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w17948_,
		_w17957_
	);
	LUT2 #(
		.INIT('h8)
	) name13911 (
		_w17950_,
		_w17953_,
		_w17958_
	);
	LUT2 #(
		.INIT('h8)
	) name13912 (
		_w17957_,
		_w17958_,
		_w17959_
	);
	LUT2 #(
		.INIT('h8)
	) name13913 (
		_w17929_,
		_w17959_,
		_w17960_
	);
	LUT2 #(
		.INIT('h8)
	) name13914 (
		_w17839_,
		_w17960_,
		_w17961_
	);
	LUT2 #(
		.INIT('h1)
	) name13915 (
		_w17956_,
		_w17961_,
		_w17962_
	);
	LUT2 #(
		.INIT('h4)
	) name13916 (
		_w17952_,
		_w17962_,
		_w17963_
	);
	LUT2 #(
		.INIT('h2)
	) name13917 (
		_w17945_,
		_w17963_,
		_w17964_
	);
	LUT2 #(
		.INIT('h4)
	) name13918 (
		_w17929_,
		_w17945_,
		_w17965_
	);
	LUT2 #(
		.INIT('h4)
	) name13919 (
		_w17849_,
		_w17861_,
		_w17966_
	);
	LUT2 #(
		.INIT('h8)
	) name13920 (
		_w17950_,
		_w17966_,
		_w17967_
	);
	LUT2 #(
		.INIT('h8)
	) name13921 (
		_w17957_,
		_w17967_,
		_w17968_
	);
	LUT2 #(
		.INIT('h8)
	) name13922 (
		_w17965_,
		_w17968_,
		_w17969_
	);
	LUT2 #(
		.INIT('h8)
	) name13923 (
		_w17917_,
		_w17957_,
		_w17970_
	);
	LUT2 #(
		.INIT('h2)
	) name13924 (
		_w17931_,
		_w17944_,
		_w17971_
	);
	LUT2 #(
		.INIT('h8)
	) name13925 (
		_w17970_,
		_w17971_,
		_w17972_
	);
	LUT2 #(
		.INIT('h4)
	) name13926 (
		_w17871_,
		_w17881_,
		_w17973_
	);
	LUT2 #(
		.INIT('h8)
	) name13927 (
		_w17849_,
		_w17861_,
		_w17974_
	);
	LUT2 #(
		.INIT('h8)
	) name13928 (
		_w17973_,
		_w17974_,
		_w17975_
	);
	LUT2 #(
		.INIT('h8)
	) name13929 (
		_w17949_,
		_w17965_,
		_w17976_
	);
	LUT2 #(
		.INIT('h8)
	) name13930 (
		_w17975_,
		_w17976_,
		_w17977_
	);
	LUT2 #(
		.INIT('h1)
	) name13931 (
		_w17972_,
		_w17977_,
		_w17978_
	);
	LUT2 #(
		.INIT('h8)
	) name13932 (
		_w17931_,
		_w17949_,
		_w17979_
	);
	LUT2 #(
		.INIT('h8)
	) name13933 (
		_w17958_,
		_w17979_,
		_w17980_
	);
	LUT2 #(
		.INIT('h4)
	) name13934 (
		_w17931_,
		_w17959_,
		_w17981_
	);
	LUT2 #(
		.INIT('h1)
	) name13935 (
		_w17980_,
		_w17981_,
		_w17982_
	);
	LUT2 #(
		.INIT('h2)
	) name13936 (
		_w17945_,
		_w17982_,
		_w17983_
	);
	LUT2 #(
		.INIT('h2)
	) name13937 (
		_w17978_,
		_w17983_,
		_w17984_
	);
	LUT2 #(
		.INIT('h8)
	) name13938 (
		_w17966_,
		_w17973_,
		_w17985_
	);
	LUT2 #(
		.INIT('h8)
	) name13939 (
		_w17920_,
		_w17985_,
		_w17986_
	);
	LUT2 #(
		.INIT('h8)
	) name13940 (
		_w17965_,
		_w17986_,
		_w17987_
	);
	LUT2 #(
		.INIT('h2)
	) name13941 (
		_w17984_,
		_w17987_,
		_w17988_
	);
	LUT2 #(
		.INIT('h4)
	) name13942 (
		_w17931_,
		_w17949_,
		_w17989_
	);
	LUT2 #(
		.INIT('h8)
	) name13943 (
		_w17953_,
		_w17973_,
		_w17990_
	);
	LUT2 #(
		.INIT('h8)
	) name13944 (
		_w17989_,
		_w17990_,
		_w17991_
	);
	LUT2 #(
		.INIT('h8)
	) name13945 (
		_w17951_,
		_w17957_,
		_w17992_
	);
	LUT2 #(
		.INIT('h4)
	) name13946 (
		_w17931_,
		_w17992_,
		_w17993_
	);
	LUT2 #(
		.INIT('h1)
	) name13947 (
		_w17991_,
		_w17993_,
		_w17994_
	);
	LUT2 #(
		.INIT('h2)
	) name13948 (
		_w17945_,
		_w17994_,
		_w17995_
	);
	LUT2 #(
		.INIT('h8)
	) name13949 (
		_w17931_,
		_w17968_,
		_w17996_
	);
	LUT2 #(
		.INIT('h8)
	) name13950 (
		_w17979_,
		_w17985_,
		_w17997_
	);
	LUT2 #(
		.INIT('h1)
	) name13951 (
		_w17996_,
		_w17997_,
		_w17998_
	);
	LUT2 #(
		.INIT('h2)
	) name13952 (
		_w17945_,
		_w17998_,
		_w17999_
	);
	LUT2 #(
		.INIT('h8)
	) name13953 (
		_w17862_,
		_w17973_,
		_w18000_
	);
	LUT2 #(
		.INIT('h8)
	) name13954 (
		_w17920_,
		_w18000_,
		_w18001_
	);
	LUT2 #(
		.INIT('h8)
	) name13955 (
		_w17971_,
		_w18001_,
		_w18002_
	);
	LUT2 #(
		.INIT('h1)
	) name13956 (
		_w17969_,
		_w18002_,
		_w18003_
	);
	LUT2 #(
		.INIT('h4)
	) name13957 (
		_w17995_,
		_w18003_,
		_w18004_
	);
	LUT2 #(
		.INIT('h4)
	) name13958 (
		_w17999_,
		_w18004_,
		_w18005_
	);
	LUT2 #(
		.INIT('h8)
	) name13959 (
		_w17988_,
		_w18005_,
		_w18006_
	);
	LUT2 #(
		.INIT('h4)
	) name13960 (
		_w17964_,
		_w18006_,
		_w18007_
	);
	LUT2 #(
		.INIT('h2)
	) name13961 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w17893_,
		_w18008_
	);
	LUT2 #(
		.INIT('h8)
	) name13962 (
		_w17902_,
		_w17945_,
		_w18009_
	);
	LUT2 #(
		.INIT('h8)
	) name13963 (
		_w18008_,
		_w18009_,
		_w18010_
	);
	LUT2 #(
		.INIT('h4)
	) name13964 (
		_w17871_,
		_w17945_,
		_w18011_
	);
	LUT2 #(
		.INIT('h8)
	) name13965 (
		_w17957_,
		_w18011_,
		_w18012_
	);
	LUT2 #(
		.INIT('h1)
	) name13966 (
		_w17946_,
		_w18008_,
		_w18013_
	);
	LUT2 #(
		.INIT('h8)
	) name13967 (
		_w18009_,
		_w18013_,
		_w18014_
	);
	LUT2 #(
		.INIT('h1)
	) name13968 (
		_w18012_,
		_w18014_,
		_w18015_
	);
	LUT2 #(
		.INIT('h4)
	) name13969 (
		_w18010_,
		_w18015_,
		_w18016_
	);
	LUT2 #(
		.INIT('h8)
	) name13970 (
		_w17883_,
		_w17949_,
		_w18017_
	);
	LUT2 #(
		.INIT('h8)
	) name13971 (
		_w17945_,
		_w18017_,
		_w18018_
	);
	LUT2 #(
		.INIT('h2)
	) name13972 (
		_w18016_,
		_w18018_,
		_w18019_
	);
	LUT2 #(
		.INIT('h8)
	) name13973 (
		_w17916_,
		_w17953_,
		_w18020_
	);
	LUT2 #(
		.INIT('h8)
	) name13974 (
		_w17957_,
		_w18020_,
		_w18021_
	);
	LUT2 #(
		.INIT('h8)
	) name13975 (
		_w17931_,
		_w18021_,
		_w18022_
	);
	LUT2 #(
		.INIT('h4)
	) name13976 (
		_w17944_,
		_w18022_,
		_w18023_
	);
	LUT2 #(
		.INIT('h2)
	) name13977 (
		_w18019_,
		_w18023_,
		_w18024_
	);
	LUT2 #(
		.INIT('h8)
	) name13978 (
		_w17945_,
		_w17949_,
		_w18025_
	);
	LUT2 #(
		.INIT('h8)
	) name13979 (
		_w17954_,
		_w18025_,
		_w18026_
	);
	LUT2 #(
		.INIT('h8)
	) name13980 (
		_w17985_,
		_w17989_,
		_w18027_
	);
	LUT2 #(
		.INIT('h8)
	) name13981 (
		_w17916_,
		_w17966_,
		_w18028_
	);
	LUT2 #(
		.INIT('h8)
	) name13982 (
		_w17957_,
		_w18028_,
		_w18029_
	);
	LUT2 #(
		.INIT('h4)
	) name13983 (
		_w17931_,
		_w18029_,
		_w18030_
	);
	LUT2 #(
		.INIT('h1)
	) name13984 (
		_w18027_,
		_w18030_,
		_w18031_
	);
	LUT2 #(
		.INIT('h2)
	) name13985 (
		_w17945_,
		_w18031_,
		_w18032_
	);
	LUT2 #(
		.INIT('h8)
	) name13986 (
		_w17949_,
		_w17975_,
		_w18033_
	);
	LUT2 #(
		.INIT('h8)
	) name13987 (
		_w17971_,
		_w18033_,
		_w18034_
	);
	LUT2 #(
		.INIT('h8)
	) name13988 (
		_w17882_,
		_w17966_,
		_w18035_
	);
	LUT2 #(
		.INIT('h8)
	) name13989 (
		_w17949_,
		_w18035_,
		_w18036_
	);
	LUT2 #(
		.INIT('h8)
	) name13990 (
		_w17945_,
		_w18036_,
		_w18037_
	);
	LUT2 #(
		.INIT('h1)
	) name13991 (
		_w18034_,
		_w18037_,
		_w18038_
	);
	LUT2 #(
		.INIT('h8)
	) name13992 (
		_w17917_,
		_w17949_,
		_w18039_
	);
	LUT2 #(
		.INIT('h8)
	) name13993 (
		_w17971_,
		_w18039_,
		_w18040_
	);
	LUT2 #(
		.INIT('h2)
	) name13994 (
		_w18038_,
		_w18040_,
		_w18041_
	);
	LUT2 #(
		.INIT('h4)
	) name13995 (
		_w18032_,
		_w18041_,
		_w18042_
	);
	LUT2 #(
		.INIT('h8)
	) name13996 (
		_w17967_,
		_w17989_,
		_w18043_
	);
	LUT2 #(
		.INIT('h4)
	) name13997 (
		_w17931_,
		_w18021_,
		_w18044_
	);
	LUT2 #(
		.INIT('h8)
	) name13998 (
		_w17916_,
		_w17974_,
		_w18045_
	);
	LUT2 #(
		.INIT('h8)
	) name13999 (
		_w17979_,
		_w18045_,
		_w18046_
	);
	LUT2 #(
		.INIT('h1)
	) name14000 (
		_w18044_,
		_w18046_,
		_w18047_
	);
	LUT2 #(
		.INIT('h4)
	) name14001 (
		_w18043_,
		_w18047_,
		_w18048_
	);
	LUT2 #(
		.INIT('h2)
	) name14002 (
		_w17945_,
		_w18048_,
		_w18049_
	);
	LUT2 #(
		.INIT('h2)
	) name14003 (
		_w18042_,
		_w18049_,
		_w18050_
	);
	LUT2 #(
		.INIT('h8)
	) name14004 (
		_w17957_,
		_w18045_,
		_w18051_
	);
	LUT2 #(
		.INIT('h8)
	) name14005 (
		_w17965_,
		_w18051_,
		_w18052_
	);
	LUT2 #(
		.INIT('h8)
	) name14006 (
		_w17971_,
		_w18029_,
		_w18053_
	);
	LUT2 #(
		.INIT('h1)
	) name14007 (
		_w18052_,
		_w18053_,
		_w18054_
	);
	LUT2 #(
		.INIT('h8)
	) name14008 (
		_w17920_,
		_w18035_,
		_w18055_
	);
	LUT2 #(
		.INIT('h8)
	) name14009 (
		_w17920_,
		_w17990_,
		_w18056_
	);
	LUT2 #(
		.INIT('h1)
	) name14010 (
		_w18055_,
		_w18056_,
		_w18057_
	);
	LUT2 #(
		.INIT('h2)
	) name14011 (
		_w17965_,
		_w18057_,
		_w18058_
	);
	LUT2 #(
		.INIT('h2)
	) name14012 (
		_w18054_,
		_w18058_,
		_w18059_
	);
	LUT2 #(
		.INIT('h8)
	) name14013 (
		_w17965_,
		_w18001_,
		_w18060_
	);
	LUT2 #(
		.INIT('h1)
	) name14014 (
		_w18026_,
		_w18060_,
		_w18061_
	);
	LUT2 #(
		.INIT('h8)
	) name14015 (
		_w18059_,
		_w18061_,
		_w18062_
	);
	LUT2 #(
		.INIT('h8)
	) name14016 (
		_w18024_,
		_w18062_,
		_w18063_
	);
	LUT2 #(
		.INIT('h8)
	) name14017 (
		_w18050_,
		_w18063_,
		_w18064_
	);
	LUT2 #(
		.INIT('h2)
	) name14018 (
		_w17971_,
		_w18057_,
		_w18065_
	);
	LUT2 #(
		.INIT('h8)
	) name14019 (
		_w17950_,
		_w17974_,
		_w18066_
	);
	LUT2 #(
		.INIT('h8)
	) name14020 (
		_w17957_,
		_w18066_,
		_w18067_
	);
	LUT2 #(
		.INIT('h1)
	) name14021 (
		_w18039_,
		_w18067_,
		_w18068_
	);
	LUT2 #(
		.INIT('h2)
	) name14022 (
		_w17965_,
		_w18068_,
		_w18069_
	);
	LUT2 #(
		.INIT('h8)
	) name14023 (
		_w17989_,
		_w18045_,
		_w18070_
	);
	LUT2 #(
		.INIT('h8)
	) name14024 (
		_w17979_,
		_w18028_,
		_w18071_
	);
	LUT2 #(
		.INIT('h8)
	) name14025 (
		_w17949_,
		_w18020_,
		_w18072_
	);
	LUT2 #(
		.INIT('h1)
	) name14026 (
		_w18070_,
		_w18072_,
		_w18073_
	);
	LUT2 #(
		.INIT('h4)
	) name14027 (
		_w18071_,
		_w18073_,
		_w18074_
	);
	LUT2 #(
		.INIT('h2)
	) name14028 (
		_w17945_,
		_w18074_,
		_w18075_
	);
	LUT2 #(
		.INIT('h1)
	) name14029 (
		_w18069_,
		_w18075_,
		_w18076_
	);
	LUT2 #(
		.INIT('h8)
	) name14030 (
		_w17882_,
		_w17974_,
		_w18077_
	);
	LUT2 #(
		.INIT('h8)
	) name14031 (
		_w17949_,
		_w18077_,
		_w18078_
	);
	LUT2 #(
		.INIT('h1)
	) name14032 (
		_w18051_,
		_w18078_,
		_w18079_
	);
	LUT2 #(
		.INIT('h2)
	) name14033 (
		_w17931_,
		_w18079_,
		_w18080_
	);
	LUT2 #(
		.INIT('h8)
	) name14034 (
		_w17949_,
		_w18000_,
		_w18081_
	);
	LUT2 #(
		.INIT('h1)
	) name14035 (
		_w17992_,
		_w18081_,
		_w18082_
	);
	LUT2 #(
		.INIT('h2)
	) name14036 (
		_w17931_,
		_w18082_,
		_w18083_
	);
	LUT2 #(
		.INIT('h1)
	) name14037 (
		_w18080_,
		_w18083_,
		_w18084_
	);
	LUT2 #(
		.INIT('h2)
	) name14038 (
		_w17945_,
		_w18084_,
		_w18085_
	);
	LUT2 #(
		.INIT('h1)
	) name14039 (
		_w18065_,
		_w18085_,
		_w18086_
	);
	LUT2 #(
		.INIT('h8)
	) name14040 (
		_w18076_,
		_w18086_,
		_w18087_
	);
	LUT2 #(
		.INIT('h2)
	) name14041 (
		_w17839_,
		_w17938_,
		_w18088_
	);
	LUT2 #(
		.INIT('h8)
	) name14042 (
		_w17920_,
		_w17975_,
		_w18089_
	);
	LUT2 #(
		.INIT('h8)
	) name14043 (
		_w17949_,
		_w18066_,
		_w18090_
	);
	LUT2 #(
		.INIT('h1)
	) name14044 (
		_w18089_,
		_w18090_,
		_w18091_
	);
	LUT2 #(
		.INIT('h1)
	) name14045 (
		_w17931_,
		_w18091_,
		_w18092_
	);
	LUT2 #(
		.INIT('h8)
	) name14046 (
		_w18088_,
		_w18092_,
		_w18093_
	);
	LUT2 #(
		.INIT('h8)
	) name14047 (
		_w17920_,
		_w17967_,
		_w18094_
	);
	LUT2 #(
		.INIT('h4)
	) name14048 (
		_w17914_,
		_w17985_,
		_w18095_
	);
	LUT2 #(
		.INIT('h1)
	) name14049 (
		_w18094_,
		_w18095_,
		_w18096_
	);
	LUT2 #(
		.INIT('h4)
	) name14050 (
		_w9264_,
		_w13832_,
		_w18097_
	);
	LUT2 #(
		.INIT('h2)
	) name14051 (
		_w14178_,
		_w18097_,
		_w18098_
	);
	LUT2 #(
		.INIT('h2)
	) name14052 (
		_w17839_,
		_w18098_,
		_w18099_
	);
	LUT2 #(
		.INIT('h4)
	) name14053 (
		_w17929_,
		_w18099_,
		_w18100_
	);
	LUT2 #(
		.INIT('h4)
	) name14054 (
		_w7369_,
		_w13832_,
		_w18101_
	);
	LUT2 #(
		.INIT('h1)
	) name14055 (
		_w14217_,
		_w18101_,
		_w18102_
	);
	LUT2 #(
		.INIT('h2)
	) name14056 (
		_w17931_,
		_w18102_,
		_w18103_
	);
	LUT2 #(
		.INIT('h1)
	) name14057 (
		_w18100_,
		_w18103_,
		_w18104_
	);
	LUT2 #(
		.INIT('h1)
	) name14058 (
		_w18096_,
		_w18104_,
		_w18105_
	);
	LUT2 #(
		.INIT('h8)
	) name14059 (
		_w17920_,
		_w18020_,
		_w18106_
	);
	LUT2 #(
		.INIT('h4)
	) name14060 (
		_w17914_,
		_w17954_,
		_w18107_
	);
	LUT2 #(
		.INIT('h1)
	) name14061 (
		_w18106_,
		_w18107_,
		_w18108_
	);
	LUT2 #(
		.INIT('h4)
	) name14062 (
		_w8406_,
		_w13832_,
		_w18109_
	);
	LUT2 #(
		.INIT('h2)
	) name14063 (
		_w14290_,
		_w18109_,
		_w18110_
	);
	LUT2 #(
		.INIT('h2)
	) name14064 (
		_w17839_,
		_w18110_,
		_w18111_
	);
	LUT2 #(
		.INIT('h4)
	) name14065 (
		_w17929_,
		_w18111_,
		_w18112_
	);
	LUT2 #(
		.INIT('h4)
	) name14066 (
		_w7805_,
		_w13832_,
		_w18113_
	);
	LUT2 #(
		.INIT('h2)
	) name14067 (
		_w14332_,
		_w18113_,
		_w18114_
	);
	LUT2 #(
		.INIT('h2)
	) name14068 (
		_w17839_,
		_w18114_,
		_w18115_
	);
	LUT2 #(
		.INIT('h8)
	) name14069 (
		_w17929_,
		_w18115_,
		_w18116_
	);
	LUT2 #(
		.INIT('h1)
	) name14070 (
		_w18112_,
		_w18116_,
		_w18117_
	);
	LUT2 #(
		.INIT('h1)
	) name14071 (
		_w18108_,
		_w18117_,
		_w18118_
	);
	LUT2 #(
		.INIT('h4)
	) name14072 (
		_w17914_,
		_w18077_,
		_w18119_
	);
	LUT2 #(
		.INIT('h8)
	) name14073 (
		_w17920_,
		_w18045_,
		_w18120_
	);
	LUT2 #(
		.INIT('h1)
	) name14074 (
		_w18119_,
		_w18120_,
		_w18121_
	);
	LUT2 #(
		.INIT('h4)
	) name14075 (
		_w7979_,
		_w13832_,
		_w18122_
	);
	LUT2 #(
		.INIT('h2)
	) name14076 (
		_w14066_,
		_w18122_,
		_w18123_
	);
	LUT2 #(
		.INIT('h2)
	) name14077 (
		_w17839_,
		_w18123_,
		_w18124_
	);
	LUT2 #(
		.INIT('h4)
	) name14078 (
		_w17929_,
		_w18124_,
		_w18125_
	);
	LUT2 #(
		.INIT('h4)
	) name14079 (
		_w8485_,
		_w13832_,
		_w18126_
	);
	LUT2 #(
		.INIT('h2)
	) name14080 (
		_w14140_,
		_w18126_,
		_w18127_
	);
	LUT2 #(
		.INIT('h2)
	) name14081 (
		_w17931_,
		_w18127_,
		_w18128_
	);
	LUT2 #(
		.INIT('h1)
	) name14082 (
		_w18125_,
		_w18128_,
		_w18129_
	);
	LUT2 #(
		.INIT('h1)
	) name14083 (
		_w18121_,
		_w18129_,
		_w18130_
	);
	LUT2 #(
		.INIT('h4)
	) name14084 (
		_w17914_,
		_w18000_,
		_w18131_
	);
	LUT2 #(
		.INIT('h8)
	) name14085 (
		_w17920_,
		_w17951_,
		_w18132_
	);
	LUT2 #(
		.INIT('h1)
	) name14086 (
		_w18131_,
		_w18132_,
		_w18133_
	);
	LUT2 #(
		.INIT('h4)
	) name14087 (
		_w10571_,
		_w13832_,
		_w18134_
	);
	LUT2 #(
		.INIT('h2)
	) name14088 (
		_w13909_,
		_w18134_,
		_w18135_
	);
	LUT2 #(
		.INIT('h2)
	) name14089 (
		_w17931_,
		_w18135_,
		_w18136_
	);
	LUT2 #(
		.INIT('h4)
	) name14090 (
		_w18133_,
		_w18136_,
		_w18137_
	);
	LUT2 #(
		.INIT('h2)
	) name14091 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7156_,
		_w18138_
	);
	LUT2 #(
		.INIT('h8)
	) name14092 (
		_w17989_,
		_w18028_,
		_w18139_
	);
	LUT2 #(
		.INIT('h8)
	) name14093 (
		_w17945_,
		_w18139_,
		_w18140_
	);
	LUT2 #(
		.INIT('h8)
	) name14094 (
		_w17955_,
		_w17971_,
		_w18141_
	);
	LUT2 #(
		.INIT('h1)
	) name14095 (
		_w18140_,
		_w18141_,
		_w18142_
	);
	LUT2 #(
		.INIT('h8)
	) name14096 (
		_w17965_,
		_w17970_,
		_w18143_
	);
	LUT2 #(
		.INIT('h8)
	) name14097 (
		_w17971_,
		_w18067_,
		_w18144_
	);
	LUT2 #(
		.INIT('h1)
	) name14098 (
		_w18143_,
		_w18144_,
		_w18145_
	);
	LUT2 #(
		.INIT('h8)
	) name14099 (
		_w18142_,
		_w18145_,
		_w18146_
	);
	LUT2 #(
		.INIT('h8)
	) name14100 (
		_w17967_,
		_w17979_,
		_w18147_
	);
	LUT2 #(
		.INIT('h8)
	) name14101 (
		_w17931_,
		_w17986_,
		_w18148_
	);
	LUT2 #(
		.INIT('h1)
	) name14102 (
		_w18147_,
		_w18148_,
		_w18149_
	);
	LUT2 #(
		.INIT('h8)
	) name14103 (
		_w17979_,
		_w17990_,
		_w18150_
	);
	LUT2 #(
		.INIT('h8)
	) name14104 (
		_w17989_,
		_w18000_,
		_w18151_
	);
	LUT2 #(
		.INIT('h1)
	) name14105 (
		_w18150_,
		_w18151_,
		_w18152_
	);
	LUT2 #(
		.INIT('h8)
	) name14106 (
		_w17920_,
		_w18077_,
		_w18153_
	);
	LUT2 #(
		.INIT('h2)
	) name14107 (
		_w18149_,
		_w18153_,
		_w18154_
	);
	LUT2 #(
		.INIT('h8)
	) name14108 (
		_w18152_,
		_w18154_,
		_w18155_
	);
	LUT2 #(
		.INIT('h2)
	) name14109 (
		_w17945_,
		_w18155_,
		_w18156_
	);
	LUT2 #(
		.INIT('h4)
	) name14110 (
		_w17914_,
		_w18035_,
		_w18157_
	);
	LUT2 #(
		.INIT('h8)
	) name14111 (
		_w17920_,
		_w18028_,
		_w18158_
	);
	LUT2 #(
		.INIT('h1)
	) name14112 (
		_w18157_,
		_w18158_,
		_w18159_
	);
	LUT2 #(
		.INIT('h4)
	) name14113 (
		_w10793_,
		_w13832_,
		_w18160_
	);
	LUT2 #(
		.INIT('h2)
	) name14114 (
		_w14022_,
		_w18160_,
		_w18161_
	);
	LUT2 #(
		.INIT('h2)
	) name14115 (
		_w17839_,
		_w18161_,
		_w18162_
	);
	LUT2 #(
		.INIT('h4)
	) name14116 (
		_w17929_,
		_w18162_,
		_w18163_
	);
	LUT2 #(
		.INIT('h4)
	) name14117 (
		_w9943_,
		_w13832_,
		_w18164_
	);
	LUT2 #(
		.INIT('h2)
	) name14118 (
		_w14101_,
		_w18164_,
		_w18165_
	);
	LUT2 #(
		.INIT('h2)
	) name14119 (
		_w17931_,
		_w18165_,
		_w18166_
	);
	LUT2 #(
		.INIT('h1)
	) name14120 (
		_w18163_,
		_w18166_,
		_w18167_
	);
	LUT2 #(
		.INIT('h1)
	) name14121 (
		_w18159_,
		_w18167_,
		_w18168_
	);
	LUT2 #(
		.INIT('h4)
	) name14122 (
		_w10222_,
		_w13832_,
		_w18169_
	);
	LUT2 #(
		.INIT('h2)
	) name14123 (
		_w13864_,
		_w18169_,
		_w18170_
	);
	LUT2 #(
		.INIT('h2)
	) name14124 (
		_w17839_,
		_w18170_,
		_w18171_
	);
	LUT2 #(
		.INIT('h4)
	) name14125 (
		_w17929_,
		_w18171_,
		_w18172_
	);
	LUT2 #(
		.INIT('h4)
	) name14126 (
		_w18133_,
		_w18172_,
		_w18173_
	);
	LUT2 #(
		.INIT('h4)
	) name14127 (
		_w11850_,
		_w13832_,
		_w18174_
	);
	LUT2 #(
		.INIT('h2)
	) name14128 (
		_w14506_,
		_w18174_,
		_w18175_
	);
	LUT2 #(
		.INIT('h2)
	) name14129 (
		_w17931_,
		_w18091_,
		_w18176_
	);
	LUT2 #(
		.INIT('h4)
	) name14130 (
		_w18175_,
		_w18176_,
		_w18177_
	);
	LUT2 #(
		.INIT('h8)
	) name14131 (
		_w17920_,
		_w17958_,
		_w18178_
	);
	LUT2 #(
		.INIT('h4)
	) name14132 (
		_w17914_,
		_w17990_,
		_w18179_
	);
	LUT2 #(
		.INIT('h1)
	) name14133 (
		_w18178_,
		_w18179_,
		_w18180_
	);
	LUT2 #(
		.INIT('h4)
	) name14134 (
		_w11235_,
		_w13832_,
		_w18181_
	);
	LUT2 #(
		.INIT('h2)
	) name14135 (
		_w13946_,
		_w18181_,
		_w18182_
	);
	LUT2 #(
		.INIT('h2)
	) name14136 (
		_w17839_,
		_w18182_,
		_w18183_
	);
	LUT2 #(
		.INIT('h4)
	) name14137 (
		_w17929_,
		_w18183_,
		_w18184_
	);
	LUT2 #(
		.INIT('h4)
	) name14138 (
		_w11307_,
		_w13832_,
		_w18185_
	);
	LUT2 #(
		.INIT('h2)
	) name14139 (
		_w13984_,
		_w18185_,
		_w18186_
	);
	LUT2 #(
		.INIT('h2)
	) name14140 (
		_w17839_,
		_w18186_,
		_w18187_
	);
	LUT2 #(
		.INIT('h8)
	) name14141 (
		_w17929_,
		_w18187_,
		_w18188_
	);
	LUT2 #(
		.INIT('h1)
	) name14142 (
		_w18184_,
		_w18188_,
		_w18189_
	);
	LUT2 #(
		.INIT('h1)
	) name14143 (
		_w18180_,
		_w18189_,
		_w18190_
	);
	LUT2 #(
		.INIT('h8)
	) name14144 (
		_w17883_,
		_w17920_,
		_w18191_
	);
	LUT2 #(
		.INIT('h8)
	) name14145 (
		_w17945_,
		_w18191_,
		_w18192_
	);
	LUT2 #(
		.INIT('h1)
	) name14146 (
		_w17958_,
		_w18077_,
		_w18193_
	);
	LUT2 #(
		.INIT('h2)
	) name14147 (
		_w17976_,
		_w18193_,
		_w18194_
	);
	LUT2 #(
		.INIT('h1)
	) name14148 (
		_w18192_,
		_w18194_,
		_w18195_
	);
	LUT2 #(
		.INIT('h1)
	) name14149 (
		_w17936_,
		_w18138_,
		_w18196_
	);
	LUT2 #(
		.INIT('h1)
	) name14150 (
		_w18105_,
		_w18118_,
		_w18197_
	);
	LUT2 #(
		.INIT('h1)
	) name14151 (
		_w18130_,
		_w18137_,
		_w18198_
	);
	LUT2 #(
		.INIT('h1)
	) name14152 (
		_w18168_,
		_w18173_,
		_w18199_
	);
	LUT2 #(
		.INIT('h4)
	) name14153 (
		_w18190_,
		_w18195_,
		_w18200_
	);
	LUT2 #(
		.INIT('h8)
	) name14154 (
		_w18199_,
		_w18200_,
		_w18201_
	);
	LUT2 #(
		.INIT('h8)
	) name14155 (
		_w18197_,
		_w18198_,
		_w18202_
	);
	LUT2 #(
		.INIT('h4)
	) name14156 (
		_w18093_,
		_w18196_,
		_w18203_
	);
	LUT2 #(
		.INIT('h4)
	) name14157 (
		_w18177_,
		_w18203_,
		_w18204_
	);
	LUT2 #(
		.INIT('h8)
	) name14158 (
		_w18201_,
		_w18202_,
		_w18205_
	);
	LUT2 #(
		.INIT('h8)
	) name14159 (
		_w18146_,
		_w18205_,
		_w18206_
	);
	LUT2 #(
		.INIT('h4)
	) name14160 (
		_w18156_,
		_w18204_,
		_w18207_
	);
	LUT2 #(
		.INIT('h8)
	) name14161 (
		_w18206_,
		_w18207_,
		_w18208_
	);
	LUT2 #(
		.INIT('h8)
	) name14162 (
		_w18064_,
		_w18087_,
		_w18209_
	);
	LUT2 #(
		.INIT('h8)
	) name14163 (
		_w18208_,
		_w18209_,
		_w18210_
	);
	LUT2 #(
		.INIT('h8)
	) name14164 (
		_w18007_,
		_w18210_,
		_w18211_
	);
	LUT2 #(
		.INIT('h4)
	) name14165 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w18211_,
		_w18212_
	);
	LUT2 #(
		.INIT('h1)
	) name14166 (
		_w17837_,
		_w18212_,
		_w18213_
	);
	LUT2 #(
		.INIT('h2)
	) name14167 (
		_w17833_,
		_w18213_,
		_w18214_
	);
	LUT2 #(
		.INIT('h1)
	) name14168 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[13]/P0001 ,
		_w17833_,
		_w18215_
	);
	LUT2 #(
		.INIT('h1)
	) name14169 (
		_w18214_,
		_w18215_,
		_w18216_
	);
	LUT2 #(
		.INIT('h2)
	) name14170 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w4112_,
		_w18217_
	);
	LUT2 #(
		.INIT('h4)
	) name14171 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w14691_,
		_w18218_
	);
	LUT2 #(
		.INIT('h4)
	) name14172 (
		_w5950_,
		_w18218_,
		_w18219_
	);
	LUT2 #(
		.INIT('h1)
	) name14173 (
		_w18217_,
		_w18219_,
		_w18220_
	);
	LUT2 #(
		.INIT('h2)
	) name14174 (
		_w14713_,
		_w18220_,
		_w18221_
	);
	LUT2 #(
		.INIT('h2)
	) name14175 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001 ,
		_w18221_,
		_w18222_
	);
	LUT2 #(
		.INIT('h8)
	) name14176 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w18221_,
		_w18223_
	);
	LUT2 #(
		.INIT('h1)
	) name14177 (
		_w18222_,
		_w18223_,
		_w18224_
	);
	LUT2 #(
		.INIT('h8)
	) name14178 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w5944_,
		_w18225_
	);
	LUT2 #(
		.INIT('h8)
	) name14179 (
		_w13761_,
		_w18225_,
		_w18226_
	);
	LUT2 #(
		.INIT('h4)
	) name14180 (
		\memc_MMR_web_reg/NET0131 ,
		_w18226_,
		_w18227_
	);
	LUT2 #(
		.INIT('h8)
	) name14181 (
		_w7237_,
		_w7283_,
		_w18228_
	);
	LUT2 #(
		.INIT('h8)
	) name14182 (
		_w18227_,
		_w18228_,
		_w18229_
	);
	LUT2 #(
		.INIT('h8)
	) name14183 (
		_w7226_,
		_w7283_,
		_w18230_
	);
	LUT2 #(
		.INIT('h8)
	) name14184 (
		_w18227_,
		_w18230_,
		_w18231_
	);
	LUT2 #(
		.INIT('h8)
	) name14185 (
		_w12688_,
		_w18231_,
		_w18232_
	);
	LUT2 #(
		.INIT('h1)
	) name14186 (
		_w18229_,
		_w18232_,
		_w18233_
	);
	LUT2 #(
		.INIT('h8)
	) name14187 (
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w18233_,
		_w18234_
	);
	LUT2 #(
		.INIT('h8)
	) name14188 (
		_w12688_,
		_w18226_,
		_w18235_
	);
	LUT2 #(
		.INIT('h8)
	) name14189 (
		_w18230_,
		_w18235_,
		_w18236_
	);
	LUT2 #(
		.INIT('h2)
	) name14190 (
		_w18229_,
		_w18236_,
		_w18237_
	);
	LUT2 #(
		.INIT('h8)
	) name14191 (
		_w9178_,
		_w18237_,
		_w18238_
	);
	LUT2 #(
		.INIT('h1)
	) name14192 (
		_w18234_,
		_w18238_,
		_w18239_
	);
	LUT2 #(
		.INIT('h2)
	) name14193 (
		_w14708_,
		_w18220_,
		_w18240_
	);
	LUT2 #(
		.INIT('h2)
	) name14194 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001 ,
		_w18240_,
		_w18241_
	);
	LUT2 #(
		.INIT('h8)
	) name14195 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w18240_,
		_w18242_
	);
	LUT2 #(
		.INIT('h1)
	) name14196 (
		_w18241_,
		_w18242_,
		_w18243_
	);
	LUT2 #(
		.INIT('h2)
	) name14197 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001 ,
		_w18240_,
		_w18244_
	);
	LUT2 #(
		.INIT('h8)
	) name14198 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w18240_,
		_w18245_
	);
	LUT2 #(
		.INIT('h1)
	) name14199 (
		_w18244_,
		_w18245_,
		_w18246_
	);
	LUT2 #(
		.INIT('h2)
	) name14200 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001 ,
		_w18240_,
		_w18247_
	);
	LUT2 #(
		.INIT('h8)
	) name14201 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w18240_,
		_w18248_
	);
	LUT2 #(
		.INIT('h1)
	) name14202 (
		_w18247_,
		_w18248_,
		_w18249_
	);
	LUT2 #(
		.INIT('h2)
	) name14203 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][6]/P0001 ,
		_w18240_,
		_w18250_
	);
	LUT2 #(
		.INIT('h4)
	) name14204 (
		_w4174_,
		_w18240_,
		_w18251_
	);
	LUT2 #(
		.INIT('h1)
	) name14205 (
		_w18250_,
		_w18251_,
		_w18252_
	);
	LUT2 #(
		.INIT('h2)
	) name14206 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001 ,
		_w18240_,
		_w18253_
	);
	LUT2 #(
		.INIT('h8)
	) name14207 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w18240_,
		_w18254_
	);
	LUT2 #(
		.INIT('h1)
	) name14208 (
		_w18253_,
		_w18254_,
		_w18255_
	);
	LUT2 #(
		.INIT('h2)
	) name14209 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001 ,
		_w18240_,
		_w18256_
	);
	LUT2 #(
		.INIT('h8)
	) name14210 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w18240_,
		_w18257_
	);
	LUT2 #(
		.INIT('h1)
	) name14211 (
		_w18256_,
		_w18257_,
		_w18258_
	);
	LUT2 #(
		.INIT('h2)
	) name14212 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001 ,
		_w18240_,
		_w18259_
	);
	LUT2 #(
		.INIT('h8)
	) name14213 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w18240_,
		_w18260_
	);
	LUT2 #(
		.INIT('h1)
	) name14214 (
		_w18259_,
		_w18260_,
		_w18261_
	);
	LUT2 #(
		.INIT('h8)
	) name14215 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w14666_,
		_w18262_
	);
	LUT2 #(
		.INIT('h4)
	) name14216 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w18263_
	);
	LUT2 #(
		.INIT('h1)
	) name14217 (
		_w17804_,
		_w18263_,
		_w18264_
	);
	LUT2 #(
		.INIT('h4)
	) name14218 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w18264_,
		_w18265_
	);
	LUT2 #(
		.INIT('h2)
	) name14219 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w18265_,
		_w18266_
	);
	LUT2 #(
		.INIT('h2)
	) name14220 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 ,
		_w18266_,
		_w18267_
	);
	LUT2 #(
		.INIT('h8)
	) name14221 (
		_w14665_,
		_w17803_,
		_w18268_
	);
	LUT2 #(
		.INIT('h4)
	) name14222 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w18268_,
		_w18269_
	);
	LUT2 #(
		.INIT('h8)
	) name14223 (
		_w18266_,
		_w18269_,
		_w18270_
	);
	LUT2 #(
		.INIT('h8)
	) name14224 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w14665_,
		_w18271_
	);
	LUT2 #(
		.INIT('h1)
	) name14225 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[6]/P0001 ,
		_w18271_,
		_w18272_
	);
	LUT2 #(
		.INIT('h2)
	) name14226 (
		_w18266_,
		_w18268_,
		_w18273_
	);
	LUT2 #(
		.INIT('h1)
	) name14227 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w11525_,
		_w18274_
	);
	LUT2 #(
		.INIT('h2)
	) name14228 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12972_,
		_w18275_
	);
	LUT2 #(
		.INIT('h1)
	) name14229 (
		_w18274_,
		_w18275_,
		_w18276_
	);
	LUT2 #(
		.INIT('h2)
	) name14230 (
		_w18271_,
		_w18276_,
		_w18277_
	);
	LUT2 #(
		.INIT('h4)
	) name14231 (
		_w18272_,
		_w18273_,
		_w18278_
	);
	LUT2 #(
		.INIT('h4)
	) name14232 (
		_w18277_,
		_w18278_,
		_w18279_
	);
	LUT2 #(
		.INIT('h1)
	) name14233 (
		_w18267_,
		_w18270_,
		_w18280_
	);
	LUT2 #(
		.INIT('h4)
	) name14234 (
		_w18279_,
		_w18280_,
		_w18281_
	);
	LUT2 #(
		.INIT('h1)
	) name14235 (
		_w18262_,
		_w18281_,
		_w18282_
	);
	LUT2 #(
		.INIT('h4)
	) name14236 (
		_w16239_,
		_w16306_,
		_w18283_
	);
	LUT2 #(
		.INIT('h1)
	) name14237 (
		_w16307_,
		_w18283_,
		_w18284_
	);
	LUT2 #(
		.INIT('h1)
	) name14238 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w18284_,
		_w18285_
	);
	LUT2 #(
		.INIT('h1)
	) name14239 (
		_w16196_,
		_w16197_,
		_w18286_
	);
	LUT2 #(
		.INIT('h4)
	) name14240 (
		_w16308_,
		_w18286_,
		_w18287_
	);
	LUT2 #(
		.INIT('h2)
	) name14241 (
		_w16308_,
		_w18286_,
		_w18288_
	);
	LUT2 #(
		.INIT('h1)
	) name14242 (
		_w18287_,
		_w18288_,
		_w18289_
	);
	LUT2 #(
		.INIT('h2)
	) name14243 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w18289_,
		_w18290_
	);
	LUT2 #(
		.INIT('h1)
	) name14244 (
		_w18285_,
		_w18290_,
		_w18291_
	);
	LUT2 #(
		.INIT('h8)
	) name14245 (
		_w18262_,
		_w18291_,
		_w18292_
	);
	LUT2 #(
		.INIT('h1)
	) name14246 (
		_w18282_,
		_w18292_,
		_w18293_
	);
	LUT2 #(
		.INIT('h2)
	) name14247 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001 ,
		_w18240_,
		_w18294_
	);
	LUT2 #(
		.INIT('h8)
	) name14248 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w18240_,
		_w18295_
	);
	LUT2 #(
		.INIT('h1)
	) name14249 (
		_w18294_,
		_w18295_,
		_w18296_
	);
	LUT2 #(
		.INIT('h2)
	) name14250 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001 ,
		_w18240_,
		_w18297_
	);
	LUT2 #(
		.INIT('h8)
	) name14251 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w18240_,
		_w18298_
	);
	LUT2 #(
		.INIT('h1)
	) name14252 (
		_w18297_,
		_w18298_,
		_w18299_
	);
	LUT2 #(
		.INIT('h2)
	) name14253 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001 ,
		_w18240_,
		_w18300_
	);
	LUT2 #(
		.INIT('h8)
	) name14254 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w18240_,
		_w18301_
	);
	LUT2 #(
		.INIT('h1)
	) name14255 (
		_w18300_,
		_w18301_,
		_w18302_
	);
	LUT2 #(
		.INIT('h2)
	) name14256 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001 ,
		_w18240_,
		_w18303_
	);
	LUT2 #(
		.INIT('h8)
	) name14257 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w18240_,
		_w18304_
	);
	LUT2 #(
		.INIT('h1)
	) name14258 (
		_w18303_,
		_w18304_,
		_w18305_
	);
	LUT2 #(
		.INIT('h2)
	) name14259 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001 ,
		_w18240_,
		_w18306_
	);
	LUT2 #(
		.INIT('h8)
	) name14260 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w18240_,
		_w18307_
	);
	LUT2 #(
		.INIT('h1)
	) name14261 (
		_w18306_,
		_w18307_,
		_w18308_
	);
	LUT2 #(
		.INIT('h2)
	) name14262 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001 ,
		_w18240_,
		_w18309_
	);
	LUT2 #(
		.INIT('h8)
	) name14263 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w18240_,
		_w18310_
	);
	LUT2 #(
		.INIT('h1)
	) name14264 (
		_w18309_,
		_w18310_,
		_w18311_
	);
	LUT2 #(
		.INIT('h2)
	) name14265 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001 ,
		_w18240_,
		_w18312_
	);
	LUT2 #(
		.INIT('h8)
	) name14266 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w18240_,
		_w18313_
	);
	LUT2 #(
		.INIT('h1)
	) name14267 (
		_w18312_,
		_w18313_,
		_w18314_
	);
	LUT2 #(
		.INIT('h2)
	) name14268 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001 ,
		_w18240_,
		_w18315_
	);
	LUT2 #(
		.INIT('h8)
	) name14269 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w18240_,
		_w18316_
	);
	LUT2 #(
		.INIT('h1)
	) name14270 (
		_w18315_,
		_w18316_,
		_w18317_
	);
	LUT2 #(
		.INIT('h2)
	) name14271 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001 ,
		_w18240_,
		_w18318_
	);
	LUT2 #(
		.INIT('h8)
	) name14272 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w18240_,
		_w18319_
	);
	LUT2 #(
		.INIT('h1)
	) name14273 (
		_w18318_,
		_w18319_,
		_w18320_
	);
	LUT2 #(
		.INIT('h2)
	) name14274 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001 ,
		_w18240_,
		_w18321_
	);
	LUT2 #(
		.INIT('h8)
	) name14275 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w18240_,
		_w18322_
	);
	LUT2 #(
		.INIT('h1)
	) name14276 (
		_w18321_,
		_w18322_,
		_w18323_
	);
	LUT2 #(
		.INIT('h2)
	) name14277 (
		_w14752_,
		_w18291_,
		_w18324_
	);
	LUT2 #(
		.INIT('h2)
	) name14278 (
		_w13801_,
		_w17804_,
		_w18325_
	);
	LUT2 #(
		.INIT('h1)
	) name14279 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w18265_,
		_w18326_
	);
	LUT2 #(
		.INIT('h8)
	) name14280 (
		_w18263_,
		_w18325_,
		_w18327_
	);
	LUT2 #(
		.INIT('h8)
	) name14281 (
		_w18326_,
		_w18327_,
		_w18328_
	);
	LUT2 #(
		.INIT('h8)
	) name14282 (
		_w18276_,
		_w18328_,
		_w18329_
	);
	LUT2 #(
		.INIT('h2)
	) name14283 (
		_w13801_,
		_w18264_,
		_w18330_
	);
	LUT2 #(
		.INIT('h2)
	) name14284 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[6]/P0001 ,
		_w18330_,
		_w18331_
	);
	LUT2 #(
		.INIT('h4)
	) name14285 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		_w17827_,
		_w18332_
	);
	LUT2 #(
		.INIT('h8)
	) name14286 (
		_w18326_,
		_w18332_,
		_w18333_
	);
	LUT2 #(
		.INIT('h1)
	) name14287 (
		_w14752_,
		_w18333_,
		_w18334_
	);
	LUT2 #(
		.INIT('h4)
	) name14288 (
		_w18331_,
		_w18334_,
		_w18335_
	);
	LUT2 #(
		.INIT('h4)
	) name14289 (
		_w18329_,
		_w18335_,
		_w18336_
	);
	LUT2 #(
		.INIT('h1)
	) name14290 (
		_w18324_,
		_w18336_,
		_w18337_
	);
	LUT2 #(
		.INIT('h2)
	) name14291 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001 ,
		_w18240_,
		_w18338_
	);
	LUT2 #(
		.INIT('h8)
	) name14292 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w18240_,
		_w18339_
	);
	LUT2 #(
		.INIT('h1)
	) name14293 (
		_w18338_,
		_w18339_,
		_w18340_
	);
	LUT2 #(
		.INIT('h2)
	) name14294 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001 ,
		_w18240_,
		_w18341_
	);
	LUT2 #(
		.INIT('h8)
	) name14295 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w18240_,
		_w18342_
	);
	LUT2 #(
		.INIT('h1)
	) name14296 (
		_w18341_,
		_w18342_,
		_w18343_
	);
	LUT2 #(
		.INIT('h2)
	) name14297 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001 ,
		_w18240_,
		_w18344_
	);
	LUT2 #(
		.INIT('h8)
	) name14298 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w18240_,
		_w18345_
	);
	LUT2 #(
		.INIT('h1)
	) name14299 (
		_w18344_,
		_w18345_,
		_w18346_
	);
	LUT2 #(
		.INIT('h2)
	) name14300 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001 ,
		_w18240_,
		_w18347_
	);
	LUT2 #(
		.INIT('h8)
	) name14301 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w18240_,
		_w18348_
	);
	LUT2 #(
		.INIT('h1)
	) name14302 (
		_w18347_,
		_w18348_,
		_w18349_
	);
	LUT2 #(
		.INIT('h2)
	) name14303 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001 ,
		_w18240_,
		_w18350_
	);
	LUT2 #(
		.INIT('h8)
	) name14304 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w18240_,
		_w18351_
	);
	LUT2 #(
		.INIT('h1)
	) name14305 (
		_w18350_,
		_w18351_,
		_w18352_
	);
	LUT2 #(
		.INIT('h2)
	) name14306 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001 ,
		_w18240_,
		_w18353_
	);
	LUT2 #(
		.INIT('h8)
	) name14307 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w18240_,
		_w18354_
	);
	LUT2 #(
		.INIT('h1)
	) name14308 (
		_w18353_,
		_w18354_,
		_w18355_
	);
	LUT2 #(
		.INIT('h2)
	) name14309 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001 ,
		_w18240_,
		_w18356_
	);
	LUT2 #(
		.INIT('h8)
	) name14310 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w18240_,
		_w18357_
	);
	LUT2 #(
		.INIT('h1)
	) name14311 (
		_w18356_,
		_w18357_,
		_w18358_
	);
	LUT2 #(
		.INIT('h2)
	) name14312 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001 ,
		_w18240_,
		_w18359_
	);
	LUT2 #(
		.INIT('h8)
	) name14313 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w18240_,
		_w18360_
	);
	LUT2 #(
		.INIT('h1)
	) name14314 (
		_w18359_,
		_w18360_,
		_w18361_
	);
	LUT2 #(
		.INIT('h2)
	) name14315 (
		_w14702_,
		_w18220_,
		_w18362_
	);
	LUT2 #(
		.INIT('h2)
	) name14316 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001 ,
		_w18362_,
		_w18363_
	);
	LUT2 #(
		.INIT('h8)
	) name14317 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w18362_,
		_w18364_
	);
	LUT2 #(
		.INIT('h1)
	) name14318 (
		_w18363_,
		_w18364_,
		_w18365_
	);
	LUT2 #(
		.INIT('h2)
	) name14319 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001 ,
		_w18362_,
		_w18366_
	);
	LUT2 #(
		.INIT('h8)
	) name14320 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w18362_,
		_w18367_
	);
	LUT2 #(
		.INIT('h1)
	) name14321 (
		_w18366_,
		_w18367_,
		_w18368_
	);
	LUT2 #(
		.INIT('h1)
	) name14322 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w18369_
	);
	LUT2 #(
		.INIT('h4)
	) name14323 (
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w18369_,
		_w18370_
	);
	LUT2 #(
		.INIT('h4)
	) name14324 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w18370_,
		_w18371_
	);
	LUT2 #(
		.INIT('h4)
	) name14325 (
		\sport0_txctl_TX_reg[4]/P0001 ,
		_w18371_,
		_w18372_
	);
	LUT2 #(
		.INIT('h4)
	) name14326 (
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w18372_,
		_w18373_
	);
	LUT2 #(
		.INIT('h4)
	) name14327 (
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w18373_,
		_w18374_
	);
	LUT2 #(
		.INIT('h4)
	) name14328 (
		\sport0_txctl_TX_reg[7]/P0001 ,
		_w18374_,
		_w18375_
	);
	LUT2 #(
		.INIT('h4)
	) name14329 (
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w18375_,
		_w18376_
	);
	LUT2 #(
		.INIT('h2)
	) name14330 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18376_,
		_w18377_
	);
	LUT2 #(
		.INIT('h8)
	) name14331 (
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w18377_,
		_w18378_
	);
	LUT2 #(
		.INIT('h1)
	) name14332 (
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w18377_,
		_w18379_
	);
	LUT2 #(
		.INIT('h1)
	) name14333 (
		_w18378_,
		_w18379_,
		_w18380_
	);
	LUT2 #(
		.INIT('h2)
	) name14334 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18372_,
		_w18381_
	);
	LUT2 #(
		.INIT('h1)
	) name14335 (
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w18381_,
		_w18382_
	);
	LUT2 #(
		.INIT('h8)
	) name14336 (
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w18381_,
		_w18383_
	);
	LUT2 #(
		.INIT('h1)
	) name14337 (
		_w18382_,
		_w18383_,
		_w18384_
	);
	LUT2 #(
		.INIT('h4)
	) name14338 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18384_,
		_w18385_
	);
	LUT2 #(
		.INIT('h4)
	) name14339 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w18386_
	);
	LUT2 #(
		.INIT('h8)
	) name14340 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w18387_
	);
	LUT2 #(
		.INIT('h2)
	) name14341 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18369_,
		_w18388_
	);
	LUT2 #(
		.INIT('h4)
	) name14342 (
		_w18387_,
		_w18388_,
		_w18389_
	);
	LUT2 #(
		.INIT('h1)
	) name14343 (
		_w18386_,
		_w18389_,
		_w18390_
	);
	LUT2 #(
		.INIT('h1)
	) name14344 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18390_,
		_w18391_
	);
	LUT2 #(
		.INIT('h8)
	) name14345 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		_w18391_,
		_w18392_
	);
	LUT2 #(
		.INIT('h2)
	) name14346 (
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w18388_,
		_w18393_
	);
	LUT2 #(
		.INIT('h4)
	) name14347 (
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w18388_,
		_w18394_
	);
	LUT2 #(
		.INIT('h1)
	) name14348 (
		_w18393_,
		_w18394_,
		_w18395_
	);
	LUT2 #(
		.INIT('h2)
	) name14349 (
		_w18392_,
		_w18395_,
		_w18396_
	);
	LUT2 #(
		.INIT('h2)
	) name14350 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18370_,
		_w18397_
	);
	LUT2 #(
		.INIT('h2)
	) name14351 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w18397_,
		_w18398_
	);
	LUT2 #(
		.INIT('h4)
	) name14352 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w18397_,
		_w18399_
	);
	LUT2 #(
		.INIT('h1)
	) name14353 (
		_w18398_,
		_w18399_,
		_w18400_
	);
	LUT2 #(
		.INIT('h2)
	) name14354 (
		_w18396_,
		_w18400_,
		_w18401_
	);
	LUT2 #(
		.INIT('h4)
	) name14355 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_TX_reg[4]/P0001 ,
		_w18402_
	);
	LUT2 #(
		.INIT('h2)
	) name14356 (
		\sport0_txctl_TX_reg[4]/P0001 ,
		_w18371_,
		_w18403_
	);
	LUT2 #(
		.INIT('h2)
	) name14357 (
		_w18381_,
		_w18403_,
		_w18404_
	);
	LUT2 #(
		.INIT('h1)
	) name14358 (
		_w18402_,
		_w18404_,
		_w18405_
	);
	LUT2 #(
		.INIT('h2)
	) name14359 (
		_w18401_,
		_w18405_,
		_w18406_
	);
	LUT2 #(
		.INIT('h1)
	) name14360 (
		_w18385_,
		_w18406_,
		_w18407_
	);
	LUT2 #(
		.INIT('h2)
	) name14361 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18373_,
		_w18408_
	);
	LUT2 #(
		.INIT('h8)
	) name14362 (
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w18408_,
		_w18409_
	);
	LUT2 #(
		.INIT('h1)
	) name14363 (
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w18408_,
		_w18410_
	);
	LUT2 #(
		.INIT('h1)
	) name14364 (
		_w18409_,
		_w18410_,
		_w18411_
	);
	LUT2 #(
		.INIT('h4)
	) name14365 (
		_w18407_,
		_w18411_,
		_w18412_
	);
	LUT2 #(
		.INIT('h2)
	) name14366 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18374_,
		_w18413_
	);
	LUT2 #(
		.INIT('h8)
	) name14367 (
		\sport0_txctl_TX_reg[7]/P0001 ,
		_w18413_,
		_w18414_
	);
	LUT2 #(
		.INIT('h1)
	) name14368 (
		\sport0_txctl_TX_reg[7]/P0001 ,
		_w18413_,
		_w18415_
	);
	LUT2 #(
		.INIT('h1)
	) name14369 (
		_w18414_,
		_w18415_,
		_w18416_
	);
	LUT2 #(
		.INIT('h8)
	) name14370 (
		_w18412_,
		_w18416_,
		_w18417_
	);
	LUT2 #(
		.INIT('h2)
	) name14371 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18375_,
		_w18418_
	);
	LUT2 #(
		.INIT('h8)
	) name14372 (
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w18418_,
		_w18419_
	);
	LUT2 #(
		.INIT('h1)
	) name14373 (
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w18418_,
		_w18420_
	);
	LUT2 #(
		.INIT('h1)
	) name14374 (
		_w18419_,
		_w18420_,
		_w18421_
	);
	LUT2 #(
		.INIT('h8)
	) name14375 (
		_w18417_,
		_w18421_,
		_w18422_
	);
	LUT2 #(
		.INIT('h8)
	) name14376 (
		_w18380_,
		_w18422_,
		_w18423_
	);
	LUT2 #(
		.INIT('h4)
	) name14377 (
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w18376_,
		_w18424_
	);
	LUT2 #(
		.INIT('h2)
	) name14378 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18424_,
		_w18425_
	);
	LUT2 #(
		.INIT('h1)
	) name14379 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		_w18425_,
		_w18426_
	);
	LUT2 #(
		.INIT('h8)
	) name14380 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18427_
	);
	LUT2 #(
		.INIT('h4)
	) name14381 (
		_w18424_,
		_w18427_,
		_w18428_
	);
	LUT2 #(
		.INIT('h1)
	) name14382 (
		_w18426_,
		_w18428_,
		_w18429_
	);
	LUT2 #(
		.INIT('h8)
	) name14383 (
		_w18423_,
		_w18429_,
		_w18430_
	);
	LUT2 #(
		.INIT('h1)
	) name14384 (
		_w18425_,
		_w18427_,
		_w18431_
	);
	LUT2 #(
		.INIT('h2)
	) name14385 (
		\sport0_txctl_TX_reg[11]/P0001 ,
		_w18431_,
		_w18432_
	);
	LUT2 #(
		.INIT('h4)
	) name14386 (
		\sport0_txctl_TX_reg[11]/P0001 ,
		_w18431_,
		_w18433_
	);
	LUT2 #(
		.INIT('h1)
	) name14387 (
		_w18432_,
		_w18433_,
		_w18434_
	);
	LUT2 #(
		.INIT('h8)
	) name14388 (
		_w18430_,
		_w18434_,
		_w18435_
	);
	LUT2 #(
		.INIT('h1)
	) name14389 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		\sport0_txctl_TX_reg[11]/P0001 ,
		_w18436_
	);
	LUT2 #(
		.INIT('h2)
	) name14390 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18436_,
		_w18437_
	);
	LUT2 #(
		.INIT('h1)
	) name14391 (
		_w18425_,
		_w18437_,
		_w18438_
	);
	LUT2 #(
		.INIT('h2)
	) name14392 (
		\sport0_txctl_TX_reg[12]/P0001 ,
		_w18438_,
		_w18439_
	);
	LUT2 #(
		.INIT('h4)
	) name14393 (
		\sport0_txctl_TX_reg[12]/P0001 ,
		_w18438_,
		_w18440_
	);
	LUT2 #(
		.INIT('h1)
	) name14394 (
		_w18439_,
		_w18440_,
		_w18441_
	);
	LUT2 #(
		.INIT('h8)
	) name14395 (
		_w18435_,
		_w18441_,
		_w18442_
	);
	LUT2 #(
		.INIT('h1)
	) name14396 (
		_w18435_,
		_w18441_,
		_w18443_
	);
	LUT2 #(
		.INIT('h1)
	) name14397 (
		_w18442_,
		_w18443_,
		_w18444_
	);
	LUT2 #(
		.INIT('h8)
	) name14398 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18444_,
		_w18445_
	);
	LUT2 #(
		.INIT('h4)
	) name14399 (
		\sport0_txctl_TX_reg[12]/P0001 ,
		_w18436_,
		_w18446_
	);
	LUT2 #(
		.INIT('h8)
	) name14400 (
		_w18424_,
		_w18446_,
		_w18447_
	);
	LUT2 #(
		.INIT('h8)
	) name14401 (
		\sport0_txctl_TX_reg[13]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18448_
	);
	LUT2 #(
		.INIT('h4)
	) name14402 (
		_w18447_,
		_w18448_,
		_w18449_
	);
	LUT2 #(
		.INIT('h2)
	) name14403 (
		\sport0_txctl_TX_reg[14]/P0001 ,
		_w18449_,
		_w18450_
	);
	LUT2 #(
		.INIT('h2)
	) name14404 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18384_,
		_w18451_
	);
	LUT2 #(
		.INIT('h2)
	) name14405 (
		_w18442_,
		_w18451_,
		_w18452_
	);
	LUT2 #(
		.INIT('h1)
	) name14406 (
		\sport0_txctl_TX_reg[13]/P0001 ,
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w18453_
	);
	LUT2 #(
		.INIT('h1)
	) name14407 (
		\sport0_txctl_TX_reg[14]/P0001 ,
		_w18453_,
		_w18454_
	);
	LUT2 #(
		.INIT('h1)
	) name14408 (
		_w18450_,
		_w18454_,
		_w18455_
	);
	LUT2 #(
		.INIT('h4)
	) name14409 (
		_w18452_,
		_w18455_,
		_w18456_
	);
	LUT2 #(
		.INIT('h4)
	) name14410 (
		_w18445_,
		_w18456_,
		_w18457_
	);
	LUT2 #(
		.INIT('h2)
	) name14411 (
		_w18430_,
		_w18451_,
		_w18458_
	);
	LUT2 #(
		.INIT('h2)
	) name14412 (
		_w18434_,
		_w18458_,
		_w18459_
	);
	LUT2 #(
		.INIT('h4)
	) name14413 (
		_w18434_,
		_w18458_,
		_w18460_
	);
	LUT2 #(
		.INIT('h1)
	) name14414 (
		_w18459_,
		_w18460_,
		_w18461_
	);
	LUT2 #(
		.INIT('h1)
	) name14415 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18461_,
		_w18462_
	);
	LUT2 #(
		.INIT('h1)
	) name14416 (
		_w18423_,
		_w18429_,
		_w18463_
	);
	LUT2 #(
		.INIT('h1)
	) name14417 (
		_w18430_,
		_w18463_,
		_w18464_
	);
	LUT2 #(
		.INIT('h8)
	) name14418 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18464_,
		_w18465_
	);
	LUT2 #(
		.INIT('h1)
	) name14419 (
		_w18462_,
		_w18465_,
		_w18466_
	);
	LUT2 #(
		.INIT('h8)
	) name14420 (
		_w18457_,
		_w18466_,
		_w18467_
	);
	LUT2 #(
		.INIT('h2)
	) name14421 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18461_,
		_w18468_
	);
	LUT2 #(
		.INIT('h4)
	) name14422 (
		_w18444_,
		_w18456_,
		_w18469_
	);
	LUT2 #(
		.INIT('h4)
	) name14423 (
		_w18468_,
		_w18469_,
		_w18470_
	);
	LUT2 #(
		.INIT('h8)
	) name14424 (
		_w18467_,
		_w18470_,
		_w18471_
	);
	LUT2 #(
		.INIT('h4)
	) name14425 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18464_,
		_w18472_
	);
	LUT2 #(
		.INIT('h2)
	) name14426 (
		_w18422_,
		_w18451_,
		_w18473_
	);
	LUT2 #(
		.INIT('h2)
	) name14427 (
		_w18380_,
		_w18473_,
		_w18474_
	);
	LUT2 #(
		.INIT('h4)
	) name14428 (
		_w18380_,
		_w18473_,
		_w18475_
	);
	LUT2 #(
		.INIT('h1)
	) name14429 (
		_w18474_,
		_w18475_,
		_w18476_
	);
	LUT2 #(
		.INIT('h2)
	) name14430 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18476_,
		_w18477_
	);
	LUT2 #(
		.INIT('h1)
	) name14431 (
		_w18472_,
		_w18477_,
		_w18478_
	);
	LUT2 #(
		.INIT('h8)
	) name14432 (
		_w18457_,
		_w18478_,
		_w18479_
	);
	LUT2 #(
		.INIT('h8)
	) name14433 (
		_w18471_,
		_w18479_,
		_w18480_
	);
	LUT2 #(
		.INIT('h4)
	) name14434 (
		_w18467_,
		_w18470_,
		_w18481_
	);
	LUT2 #(
		.INIT('h1)
	) name14435 (
		_w18480_,
		_w18481_,
		_w18482_
	);
	LUT2 #(
		.INIT('h2)
	) name14436 (
		_w18407_,
		_w18411_,
		_w18483_
	);
	LUT2 #(
		.INIT('h1)
	) name14437 (
		_w18412_,
		_w18483_,
		_w18484_
	);
	LUT2 #(
		.INIT('h1)
	) name14438 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18484_,
		_w18485_
	);
	LUT2 #(
		.INIT('h1)
	) name14439 (
		_w18385_,
		_w18451_,
		_w18486_
	);
	LUT2 #(
		.INIT('h8)
	) name14440 (
		_w18406_,
		_w18486_,
		_w18487_
	);
	LUT2 #(
		.INIT('h1)
	) name14441 (
		_w18406_,
		_w18486_,
		_w18488_
	);
	LUT2 #(
		.INIT('h1)
	) name14442 (
		_w18487_,
		_w18488_,
		_w18489_
	);
	LUT2 #(
		.INIT('h2)
	) name14443 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18489_,
		_w18490_
	);
	LUT2 #(
		.INIT('h1)
	) name14444 (
		_w18485_,
		_w18490_,
		_w18491_
	);
	LUT2 #(
		.INIT('h8)
	) name14445 (
		_w18457_,
		_w18491_,
		_w18492_
	);
	LUT2 #(
		.INIT('h2)
	) name14446 (
		_w18412_,
		_w18451_,
		_w18493_
	);
	LUT2 #(
		.INIT('h2)
	) name14447 (
		_w18416_,
		_w18493_,
		_w18494_
	);
	LUT2 #(
		.INIT('h4)
	) name14448 (
		_w18416_,
		_w18493_,
		_w18495_
	);
	LUT2 #(
		.INIT('h1)
	) name14449 (
		_w18494_,
		_w18495_,
		_w18496_
	);
	LUT2 #(
		.INIT('h1)
	) name14450 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18496_,
		_w18497_
	);
	LUT2 #(
		.INIT('h8)
	) name14451 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18484_,
		_w18498_
	);
	LUT2 #(
		.INIT('h1)
	) name14452 (
		_w18497_,
		_w18498_,
		_w18499_
	);
	LUT2 #(
		.INIT('h8)
	) name14453 (
		_w18457_,
		_w18499_,
		_w18500_
	);
	LUT2 #(
		.INIT('h8)
	) name14454 (
		_w18492_,
		_w18500_,
		_w18501_
	);
	LUT2 #(
		.INIT('h2)
	) name14455 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18496_,
		_w18502_
	);
	LUT2 #(
		.INIT('h1)
	) name14456 (
		_w18417_,
		_w18421_,
		_w18503_
	);
	LUT2 #(
		.INIT('h1)
	) name14457 (
		_w18422_,
		_w18503_,
		_w18504_
	);
	LUT2 #(
		.INIT('h4)
	) name14458 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18504_,
		_w18505_
	);
	LUT2 #(
		.INIT('h1)
	) name14459 (
		_w18502_,
		_w18505_,
		_w18506_
	);
	LUT2 #(
		.INIT('h8)
	) name14460 (
		_w18457_,
		_w18506_,
		_w18507_
	);
	LUT2 #(
		.INIT('h4)
	) name14461 (
		_w18501_,
		_w18507_,
		_w18508_
	);
	LUT2 #(
		.INIT('h1)
	) name14462 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18476_,
		_w18509_
	);
	LUT2 #(
		.INIT('h8)
	) name14463 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18504_,
		_w18510_
	);
	LUT2 #(
		.INIT('h1)
	) name14464 (
		_w18509_,
		_w18510_,
		_w18511_
	);
	LUT2 #(
		.INIT('h8)
	) name14465 (
		_w18457_,
		_w18511_,
		_w18512_
	);
	LUT2 #(
		.INIT('h8)
	) name14466 (
		_w18479_,
		_w18512_,
		_w18513_
	);
	LUT2 #(
		.INIT('h8)
	) name14467 (
		_w18471_,
		_w18513_,
		_w18514_
	);
	LUT2 #(
		.INIT('h4)
	) name14468 (
		_w18508_,
		_w18514_,
		_w18515_
	);
	LUT2 #(
		.INIT('h1)
	) name14469 (
		_w18482_,
		_w18515_,
		_w18516_
	);
	LUT2 #(
		.INIT('h2)
	) name14470 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w18516_,
		_w18517_
	);
	LUT2 #(
		.INIT('h8)
	) name14471 (
		\core_c_dec_MTTX0_E_reg/P0001 ,
		_w5951_,
		_w18518_
	);
	LUT2 #(
		.INIT('h1)
	) name14472 (
		\auctl_T0Sack_reg/NET0131 ,
		_w18518_,
		_w18519_
	);
	LUT2 #(
		.INIT('h8)
	) name14473 (
		\sport0_txctl_TX_reg[4]/P0001 ,
		_w18519_,
		_w18520_
	);
	LUT2 #(
		.INIT('h2)
	) name14474 (
		_w10069_,
		_w18519_,
		_w18521_
	);
	LUT2 #(
		.INIT('h1)
	) name14475 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w18520_,
		_w18522_
	);
	LUT2 #(
		.INIT('h4)
	) name14476 (
		_w18521_,
		_w18522_,
		_w18523_
	);
	LUT2 #(
		.INIT('h1)
	) name14477 (
		_w18517_,
		_w18523_,
		_w18524_
	);
	LUT2 #(
		.INIT('h2)
	) name14478 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001 ,
		_w18362_,
		_w18525_
	);
	LUT2 #(
		.INIT('h8)
	) name14479 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w18362_,
		_w18526_
	);
	LUT2 #(
		.INIT('h1)
	) name14480 (
		_w18525_,
		_w18526_,
		_w18527_
	);
	LUT2 #(
		.INIT('h2)
	) name14481 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][6]/P0001 ,
		_w18362_,
		_w18528_
	);
	LUT2 #(
		.INIT('h4)
	) name14482 (
		_w4174_,
		_w18362_,
		_w18529_
	);
	LUT2 #(
		.INIT('h1)
	) name14483 (
		_w18528_,
		_w18529_,
		_w18530_
	);
	LUT2 #(
		.INIT('h2)
	) name14484 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001 ,
		_w18362_,
		_w18531_
	);
	LUT2 #(
		.INIT('h8)
	) name14485 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w18362_,
		_w18532_
	);
	LUT2 #(
		.INIT('h1)
	) name14486 (
		_w18531_,
		_w18532_,
		_w18533_
	);
	LUT2 #(
		.INIT('h2)
	) name14487 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001 ,
		_w18362_,
		_w18534_
	);
	LUT2 #(
		.INIT('h8)
	) name14488 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w18362_,
		_w18535_
	);
	LUT2 #(
		.INIT('h1)
	) name14489 (
		_w18534_,
		_w18535_,
		_w18536_
	);
	LUT2 #(
		.INIT('h2)
	) name14490 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001 ,
		_w18362_,
		_w18537_
	);
	LUT2 #(
		.INIT('h8)
	) name14491 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w18362_,
		_w18538_
	);
	LUT2 #(
		.INIT('h1)
	) name14492 (
		_w18537_,
		_w18538_,
		_w18539_
	);
	LUT2 #(
		.INIT('h2)
	) name14493 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001 ,
		_w18362_,
		_w18540_
	);
	LUT2 #(
		.INIT('h8)
	) name14494 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w18362_,
		_w18541_
	);
	LUT2 #(
		.INIT('h1)
	) name14495 (
		_w18540_,
		_w18541_,
		_w18542_
	);
	LUT2 #(
		.INIT('h2)
	) name14496 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001 ,
		_w18362_,
		_w18543_
	);
	LUT2 #(
		.INIT('h8)
	) name14497 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w18362_,
		_w18544_
	);
	LUT2 #(
		.INIT('h1)
	) name14498 (
		_w18543_,
		_w18544_,
		_w18545_
	);
	LUT2 #(
		.INIT('h2)
	) name14499 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001 ,
		_w18362_,
		_w18546_
	);
	LUT2 #(
		.INIT('h8)
	) name14500 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w18362_,
		_w18547_
	);
	LUT2 #(
		.INIT('h1)
	) name14501 (
		_w18546_,
		_w18547_,
		_w18548_
	);
	LUT2 #(
		.INIT('h2)
	) name14502 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001 ,
		_w18362_,
		_w18549_
	);
	LUT2 #(
		.INIT('h8)
	) name14503 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w18362_,
		_w18550_
	);
	LUT2 #(
		.INIT('h1)
	) name14504 (
		_w18549_,
		_w18550_,
		_w18551_
	);
	LUT2 #(
		.INIT('h2)
	) name14505 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001 ,
		_w18362_,
		_w18552_
	);
	LUT2 #(
		.INIT('h8)
	) name14506 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w18362_,
		_w18553_
	);
	LUT2 #(
		.INIT('h1)
	) name14507 (
		_w18552_,
		_w18553_,
		_w18554_
	);
	LUT2 #(
		.INIT('h2)
	) name14508 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001 ,
		_w18362_,
		_w18555_
	);
	LUT2 #(
		.INIT('h8)
	) name14509 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w18362_,
		_w18556_
	);
	LUT2 #(
		.INIT('h1)
	) name14510 (
		_w18555_,
		_w18556_,
		_w18557_
	);
	LUT2 #(
		.INIT('h2)
	) name14511 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001 ,
		_w18362_,
		_w18558_
	);
	LUT2 #(
		.INIT('h8)
	) name14512 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w18362_,
		_w18559_
	);
	LUT2 #(
		.INIT('h1)
	) name14513 (
		_w18558_,
		_w18559_,
		_w18560_
	);
	LUT2 #(
		.INIT('h2)
	) name14514 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001 ,
		_w18362_,
		_w18561_
	);
	LUT2 #(
		.INIT('h8)
	) name14515 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w18362_,
		_w18562_
	);
	LUT2 #(
		.INIT('h1)
	) name14516 (
		_w18561_,
		_w18562_,
		_w18563_
	);
	LUT2 #(
		.INIT('h2)
	) name14517 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001 ,
		_w18362_,
		_w18564_
	);
	LUT2 #(
		.INIT('h8)
	) name14518 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w18362_,
		_w18565_
	);
	LUT2 #(
		.INIT('h1)
	) name14519 (
		_w18564_,
		_w18565_,
		_w18566_
	);
	LUT2 #(
		.INIT('h2)
	) name14520 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001 ,
		_w18362_,
		_w18567_
	);
	LUT2 #(
		.INIT('h8)
	) name14521 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w18362_,
		_w18568_
	);
	LUT2 #(
		.INIT('h1)
	) name14522 (
		_w18567_,
		_w18568_,
		_w18569_
	);
	LUT2 #(
		.INIT('h2)
	) name14523 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001 ,
		_w18362_,
		_w18570_
	);
	LUT2 #(
		.INIT('h8)
	) name14524 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w18362_,
		_w18571_
	);
	LUT2 #(
		.INIT('h1)
	) name14525 (
		_w18570_,
		_w18571_,
		_w18572_
	);
	LUT2 #(
		.INIT('h2)
	) name14526 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001 ,
		_w18362_,
		_w18573_
	);
	LUT2 #(
		.INIT('h8)
	) name14527 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w18362_,
		_w18574_
	);
	LUT2 #(
		.INIT('h1)
	) name14528 (
		_w18573_,
		_w18574_,
		_w18575_
	);
	LUT2 #(
		.INIT('h2)
	) name14529 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001 ,
		_w18362_,
		_w18576_
	);
	LUT2 #(
		.INIT('h8)
	) name14530 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w18362_,
		_w18577_
	);
	LUT2 #(
		.INIT('h1)
	) name14531 (
		_w18576_,
		_w18577_,
		_w18578_
	);
	LUT2 #(
		.INIT('h2)
	) name14532 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001 ,
		_w18362_,
		_w18579_
	);
	LUT2 #(
		.INIT('h8)
	) name14533 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w18362_,
		_w18580_
	);
	LUT2 #(
		.INIT('h1)
	) name14534 (
		_w18579_,
		_w18580_,
		_w18581_
	);
	LUT2 #(
		.INIT('h2)
	) name14535 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001 ,
		_w18362_,
		_w18582_
	);
	LUT2 #(
		.INIT('h8)
	) name14536 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w18362_,
		_w18583_
	);
	LUT2 #(
		.INIT('h1)
	) name14537 (
		_w18582_,
		_w18583_,
		_w18584_
	);
	LUT2 #(
		.INIT('h2)
	) name14538 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001 ,
		_w18362_,
		_w18585_
	);
	LUT2 #(
		.INIT('h8)
	) name14539 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w18362_,
		_w18586_
	);
	LUT2 #(
		.INIT('h1)
	) name14540 (
		_w18585_,
		_w18586_,
		_w18587_
	);
	LUT2 #(
		.INIT('h2)
	) name14541 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001 ,
		_w18362_,
		_w18588_
	);
	LUT2 #(
		.INIT('h8)
	) name14542 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w18362_,
		_w18589_
	);
	LUT2 #(
		.INIT('h1)
	) name14543 (
		_w18588_,
		_w18589_,
		_w18590_
	);
	LUT2 #(
		.INIT('h2)
	) name14544 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001 ,
		_w18362_,
		_w18591_
	);
	LUT2 #(
		.INIT('h8)
	) name14545 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w18362_,
		_w18592_
	);
	LUT2 #(
		.INIT('h1)
	) name14546 (
		_w18591_,
		_w18592_,
		_w18593_
	);
	LUT2 #(
		.INIT('h2)
	) name14547 (
		_w14695_,
		_w18220_,
		_w18594_
	);
	LUT2 #(
		.INIT('h2)
	) name14548 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001 ,
		_w18594_,
		_w18595_
	);
	LUT2 #(
		.INIT('h8)
	) name14549 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w18594_,
		_w18596_
	);
	LUT2 #(
		.INIT('h1)
	) name14550 (
		_w18595_,
		_w18596_,
		_w18597_
	);
	LUT2 #(
		.INIT('h2)
	) name14551 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001 ,
		_w18594_,
		_w18598_
	);
	LUT2 #(
		.INIT('h8)
	) name14552 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w18594_,
		_w18599_
	);
	LUT2 #(
		.INIT('h1)
	) name14553 (
		_w18598_,
		_w18599_,
		_w18600_
	);
	LUT2 #(
		.INIT('h2)
	) name14554 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001 ,
		_w18594_,
		_w18601_
	);
	LUT2 #(
		.INIT('h8)
	) name14555 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w18594_,
		_w18602_
	);
	LUT2 #(
		.INIT('h1)
	) name14556 (
		_w18601_,
		_w18602_,
		_w18603_
	);
	LUT2 #(
		.INIT('h2)
	) name14557 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][6]/P0001 ,
		_w18594_,
		_w18604_
	);
	LUT2 #(
		.INIT('h4)
	) name14558 (
		_w4174_,
		_w18594_,
		_w18605_
	);
	LUT2 #(
		.INIT('h1)
	) name14559 (
		_w18604_,
		_w18605_,
		_w18606_
	);
	LUT2 #(
		.INIT('h2)
	) name14560 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001 ,
		_w18594_,
		_w18607_
	);
	LUT2 #(
		.INIT('h8)
	) name14561 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w18594_,
		_w18608_
	);
	LUT2 #(
		.INIT('h1)
	) name14562 (
		_w18607_,
		_w18608_,
		_w18609_
	);
	LUT2 #(
		.INIT('h2)
	) name14563 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001 ,
		_w18594_,
		_w18610_
	);
	LUT2 #(
		.INIT('h8)
	) name14564 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w18594_,
		_w18611_
	);
	LUT2 #(
		.INIT('h1)
	) name14565 (
		_w18610_,
		_w18611_,
		_w18612_
	);
	LUT2 #(
		.INIT('h2)
	) name14566 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001 ,
		_w18594_,
		_w18613_
	);
	LUT2 #(
		.INIT('h8)
	) name14567 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w18594_,
		_w18614_
	);
	LUT2 #(
		.INIT('h1)
	) name14568 (
		_w18613_,
		_w18614_,
		_w18615_
	);
	LUT2 #(
		.INIT('h2)
	) name14569 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001 ,
		_w18594_,
		_w18616_
	);
	LUT2 #(
		.INIT('h8)
	) name14570 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w18594_,
		_w18617_
	);
	LUT2 #(
		.INIT('h1)
	) name14571 (
		_w18616_,
		_w18617_,
		_w18618_
	);
	LUT2 #(
		.INIT('h2)
	) name14572 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001 ,
		_w18594_,
		_w18619_
	);
	LUT2 #(
		.INIT('h8)
	) name14573 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w18594_,
		_w18620_
	);
	LUT2 #(
		.INIT('h1)
	) name14574 (
		_w18619_,
		_w18620_,
		_w18621_
	);
	LUT2 #(
		.INIT('h2)
	) name14575 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001 ,
		_w18594_,
		_w18622_
	);
	LUT2 #(
		.INIT('h8)
	) name14576 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w18594_,
		_w18623_
	);
	LUT2 #(
		.INIT('h1)
	) name14577 (
		_w18622_,
		_w18623_,
		_w18624_
	);
	LUT2 #(
		.INIT('h2)
	) name14578 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001 ,
		_w18594_,
		_w18625_
	);
	LUT2 #(
		.INIT('h8)
	) name14579 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w18594_,
		_w18626_
	);
	LUT2 #(
		.INIT('h1)
	) name14580 (
		_w18625_,
		_w18626_,
		_w18627_
	);
	LUT2 #(
		.INIT('h2)
	) name14581 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001 ,
		_w18594_,
		_w18628_
	);
	LUT2 #(
		.INIT('h8)
	) name14582 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w18594_,
		_w18629_
	);
	LUT2 #(
		.INIT('h1)
	) name14583 (
		_w18628_,
		_w18629_,
		_w18630_
	);
	LUT2 #(
		.INIT('h2)
	) name14584 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001 ,
		_w18594_,
		_w18631_
	);
	LUT2 #(
		.INIT('h8)
	) name14585 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w18594_,
		_w18632_
	);
	LUT2 #(
		.INIT('h1)
	) name14586 (
		_w18631_,
		_w18632_,
		_w18633_
	);
	LUT2 #(
		.INIT('h2)
	) name14587 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001 ,
		_w18594_,
		_w18634_
	);
	LUT2 #(
		.INIT('h8)
	) name14588 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w18594_,
		_w18635_
	);
	LUT2 #(
		.INIT('h1)
	) name14589 (
		_w18634_,
		_w18635_,
		_w18636_
	);
	LUT2 #(
		.INIT('h2)
	) name14590 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001 ,
		_w18594_,
		_w18637_
	);
	LUT2 #(
		.INIT('h8)
	) name14591 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w18594_,
		_w18638_
	);
	LUT2 #(
		.INIT('h1)
	) name14592 (
		_w18637_,
		_w18638_,
		_w18639_
	);
	LUT2 #(
		.INIT('h2)
	) name14593 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001 ,
		_w18594_,
		_w18640_
	);
	LUT2 #(
		.INIT('h8)
	) name14594 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w18594_,
		_w18641_
	);
	LUT2 #(
		.INIT('h1)
	) name14595 (
		_w18640_,
		_w18641_,
		_w18642_
	);
	LUT2 #(
		.INIT('h2)
	) name14596 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001 ,
		_w18594_,
		_w18643_
	);
	LUT2 #(
		.INIT('h8)
	) name14597 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w18594_,
		_w18644_
	);
	LUT2 #(
		.INIT('h1)
	) name14598 (
		_w18643_,
		_w18644_,
		_w18645_
	);
	LUT2 #(
		.INIT('h2)
	) name14599 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001 ,
		_w18594_,
		_w18646_
	);
	LUT2 #(
		.INIT('h8)
	) name14600 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w18594_,
		_w18647_
	);
	LUT2 #(
		.INIT('h1)
	) name14601 (
		_w18646_,
		_w18647_,
		_w18648_
	);
	LUT2 #(
		.INIT('h2)
	) name14602 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001 ,
		_w18594_,
		_w18649_
	);
	LUT2 #(
		.INIT('h8)
	) name14603 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w18594_,
		_w18650_
	);
	LUT2 #(
		.INIT('h1)
	) name14604 (
		_w18649_,
		_w18650_,
		_w18651_
	);
	LUT2 #(
		.INIT('h8)
	) name14605 (
		_w7284_,
		_w18227_,
		_w18652_
	);
	LUT2 #(
		.INIT('h1)
	) name14606 (
		_w18232_,
		_w18652_,
		_w18653_
	);
	LUT2 #(
		.INIT('h8)
	) name14607 (
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w18653_,
		_w18654_
	);
	LUT2 #(
		.INIT('h4)
	) name14608 (
		_w18236_,
		_w18652_,
		_w18655_
	);
	LUT2 #(
		.INIT('h8)
	) name14609 (
		_w10289_,
		_w18655_,
		_w18656_
	);
	LUT2 #(
		.INIT('h1)
	) name14610 (
		_w18654_,
		_w18656_,
		_w18657_
	);
	LUT2 #(
		.INIT('h2)
	) name14611 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001 ,
		_w18594_,
		_w18658_
	);
	LUT2 #(
		.INIT('h8)
	) name14612 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w18594_,
		_w18659_
	);
	LUT2 #(
		.INIT('h1)
	) name14613 (
		_w18658_,
		_w18659_,
		_w18660_
	);
	LUT2 #(
		.INIT('h2)
	) name14614 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001 ,
		_w18594_,
		_w18661_
	);
	LUT2 #(
		.INIT('h8)
	) name14615 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w18594_,
		_w18662_
	);
	LUT2 #(
		.INIT('h1)
	) name14616 (
		_w18661_,
		_w18662_,
		_w18663_
	);
	LUT2 #(
		.INIT('h2)
	) name14617 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001 ,
		_w18594_,
		_w18664_
	);
	LUT2 #(
		.INIT('h8)
	) name14618 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w18594_,
		_w18665_
	);
	LUT2 #(
		.INIT('h1)
	) name14619 (
		_w18664_,
		_w18665_,
		_w18666_
	);
	LUT2 #(
		.INIT('h2)
	) name14620 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001 ,
		_w18594_,
		_w18667_
	);
	LUT2 #(
		.INIT('h8)
	) name14621 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w18594_,
		_w18668_
	);
	LUT2 #(
		.INIT('h1)
	) name14622 (
		_w18667_,
		_w18668_,
		_w18669_
	);
	LUT2 #(
		.INIT('h8)
	) name14623 (
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w18653_,
		_w18670_
	);
	LUT2 #(
		.INIT('h8)
	) name14624 (
		_w10638_,
		_w18655_,
		_w18671_
	);
	LUT2 #(
		.INIT('h1)
	) name14625 (
		_w18670_,
		_w18671_,
		_w18672_
	);
	LUT2 #(
		.INIT('h2)
	) name14626 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001 ,
		_w18594_,
		_w18673_
	);
	LUT2 #(
		.INIT('h8)
	) name14627 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w18594_,
		_w18674_
	);
	LUT2 #(
		.INIT('h1)
	) name14628 (
		_w18673_,
		_w18674_,
		_w18675_
	);
	LUT2 #(
		.INIT('h2)
	) name14629 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001 ,
		_w18594_,
		_w18676_
	);
	LUT2 #(
		.INIT('h8)
	) name14630 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w18594_,
		_w18677_
	);
	LUT2 #(
		.INIT('h1)
	) name14631 (
		_w18676_,
		_w18677_,
		_w18678_
	);
	LUT2 #(
		.INIT('h2)
	) name14632 (
		_w14694_,
		_w18220_,
		_w18679_
	);
	LUT2 #(
		.INIT('h1)
	) name14633 (
		_w5950_,
		_w14692_,
		_w18680_
	);
	LUT2 #(
		.INIT('h8)
	) name14634 (
		_w14696_,
		_w18680_,
		_w18681_
	);
	LUT2 #(
		.INIT('h8)
	) name14635 (
		_w14701_,
		_w18220_,
		_w18682_
	);
	LUT2 #(
		.INIT('h8)
	) name14636 (
		_w18681_,
		_w18682_,
		_w18683_
	);
	LUT2 #(
		.INIT('h1)
	) name14637 (
		_w18679_,
		_w18683_,
		_w18684_
	);
	LUT2 #(
		.INIT('h8)
	) name14638 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w18684_,
		_w18685_
	);
	LUT2 #(
		.INIT('h1)
	) name14639 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w18684_,
		_w18686_
	);
	LUT2 #(
		.INIT('h1)
	) name14640 (
		_w18685_,
		_w18686_,
		_w18687_
	);
	LUT2 #(
		.INIT('h1)
	) name14641 (
		_w14711_,
		_w18220_,
		_w18688_
	);
	LUT2 #(
		.INIT('h1)
	) name14642 (
		_w18681_,
		_w18688_,
		_w18689_
	);
	LUT2 #(
		.INIT('h1)
	) name14643 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		_w18689_,
		_w18690_
	);
	LUT2 #(
		.INIT('h8)
	) name14644 (
		\core_c_psq_ststk_ptr_reg[0]/NET0131 ,
		_w18689_,
		_w18691_
	);
	LUT2 #(
		.INIT('h1)
	) name14645 (
		_w18690_,
		_w18691_,
		_w18692_
	);
	LUT2 #(
		.INIT('h8)
	) name14646 (
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w18653_,
		_w18693_
	);
	LUT2 #(
		.INIT('h8)
	) name14647 (
		_w12688_,
		_w18655_,
		_w18694_
	);
	LUT2 #(
		.INIT('h1)
	) name14648 (
		_w18693_,
		_w18694_,
		_w18695_
	);
	LUT2 #(
		.INIT('h1)
	) name14649 (
		_w13806_,
		_w14551_,
		_w18696_
	);
	LUT2 #(
		.INIT('h2)
	) name14650 (
		_w13806_,
		_w14413_,
		_w18697_
	);
	LUT2 #(
		.INIT('h1)
	) name14651 (
		_w18696_,
		_w18697_,
		_w18698_
	);
	LUT2 #(
		.INIT('h2)
	) name14652 (
		_w14667_,
		_w18698_,
		_w18699_
	);
	LUT2 #(
		.INIT('h2)
	) name14653 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[13]/P0001 ,
		_w14667_,
		_w18700_
	);
	LUT2 #(
		.INIT('h1)
	) name14654 (
		_w18699_,
		_w18700_,
		_w18701_
	);
	LUT2 #(
		.INIT('h8)
	) name14655 (
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w18653_,
		_w18702_
	);
	LUT2 #(
		.INIT('h8)
	) name14656 (
		_w7340_,
		_w18655_,
		_w18703_
	);
	LUT2 #(
		.INIT('h1)
	) name14657 (
		_w18702_,
		_w18703_,
		_w18704_
	);
	LUT2 #(
		.INIT('h8)
	) name14658 (
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w18653_,
		_w18705_
	);
	LUT2 #(
		.INIT('h8)
	) name14659 (
		_w12743_,
		_w18655_,
		_w18706_
	);
	LUT2 #(
		.INIT('h1)
	) name14660 (
		_w18705_,
		_w18706_,
		_w18707_
	);
	LUT2 #(
		.INIT('h8)
	) name14661 (
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w18653_,
		_w18708_
	);
	LUT2 #(
		.INIT('h8)
	) name14662 (
		_w9178_,
		_w18655_,
		_w18709_
	);
	LUT2 #(
		.INIT('h1)
	) name14663 (
		_w18708_,
		_w18709_,
		_w18710_
	);
	LUT2 #(
		.INIT('h8)
	) name14664 (
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w18653_,
		_w18711_
	);
	LUT2 #(
		.INIT('h8)
	) name14665 (
		_w8460_,
		_w18655_,
		_w18712_
	);
	LUT2 #(
		.INIT('h1)
	) name14666 (
		_w18711_,
		_w18712_,
		_w18713_
	);
	LUT2 #(
		.INIT('h8)
	) name14667 (
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w18653_,
		_w18714_
	);
	LUT2 #(
		.INIT('h8)
	) name14668 (
		_w7859_,
		_w18655_,
		_w18715_
	);
	LUT2 #(
		.INIT('h1)
	) name14669 (
		_w18714_,
		_w18715_,
		_w18716_
	);
	LUT2 #(
		.INIT('h2)
	) name14670 (
		_w14666_,
		_w17832_,
		_w18717_
	);
	LUT2 #(
		.INIT('h2)
	) name14671 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w18276_,
		_w18718_
	);
	LUT2 #(
		.INIT('h8)
	) name14672 (
		_w17931_,
		_w18153_,
		_w18719_
	);
	LUT2 #(
		.INIT('h1)
	) name14673 (
		_w18046_,
		_w18719_,
		_w18720_
	);
	LUT2 #(
		.INIT('h2)
	) name14674 (
		_w18111_,
		_w18720_,
		_w18721_
	);
	LUT2 #(
		.INIT('h2)
	) name14675 (
		_w17931_,
		_w18161_,
		_w18722_
	);
	LUT2 #(
		.INIT('h4)
	) name14676 (
		_w17922_,
		_w18722_,
		_w18723_
	);
	LUT2 #(
		.INIT('h4)
	) name14677 (
		_w18032_,
		_w18145_,
		_w18724_
	);
	LUT2 #(
		.INIT('h8)
	) name14678 (
		_w18020_,
		_w18025_,
		_w18725_
	);
	LUT2 #(
		.INIT('h2)
	) name14679 (
		_w18724_,
		_w18725_,
		_w18726_
	);
	LUT2 #(
		.INIT('h2)
	) name14680 (
		_w18038_,
		_w18141_,
		_w18727_
	);
	LUT2 #(
		.INIT('h1)
	) name14681 (
		_w18040_,
		_w18069_,
		_w18728_
	);
	LUT2 #(
		.INIT('h8)
	) name14682 (
		_w18195_,
		_w18728_,
		_w18729_
	);
	LUT2 #(
		.INIT('h8)
	) name14683 (
		_w18727_,
		_w18729_,
		_w18730_
	);
	LUT2 #(
		.INIT('h8)
	) name14684 (
		_w18726_,
		_w18730_,
		_w18731_
	);
	LUT2 #(
		.INIT('h8)
	) name14685 (
		_w17931_,
		_w18090_,
		_w18732_
	);
	LUT2 #(
		.INIT('h4)
	) name14686 (
		_w18182_,
		_w18732_,
		_w18733_
	);
	LUT2 #(
		.INIT('h1)
	) name14687 (
		_w17991_,
		_w17997_,
		_w18734_
	);
	LUT2 #(
		.INIT('h2)
	) name14688 (
		_w17945_,
		_w18734_,
		_w18735_
	);
	LUT2 #(
		.INIT('h1)
	) name14689 (
		_w17968_,
		_w17993_,
		_w18736_
	);
	LUT2 #(
		.INIT('h2)
	) name14690 (
		_w17945_,
		_w18736_,
		_w18737_
	);
	LUT2 #(
		.INIT('h1)
	) name14691 (
		_w18735_,
		_w18737_,
		_w18738_
	);
	LUT2 #(
		.INIT('h2)
	) name14692 (
		_w18147_,
		_w18170_,
		_w18739_
	);
	LUT2 #(
		.INIT('h2)
	) name14693 (
		_w17839_,
		_w18127_,
		_w18740_
	);
	LUT2 #(
		.INIT('h4)
	) name14694 (
		_w17929_,
		_w18740_,
		_w18741_
	);
	LUT2 #(
		.INIT('h2)
	) name14695 (
		_w17931_,
		_w18098_,
		_w18742_
	);
	LUT2 #(
		.INIT('h1)
	) name14696 (
		_w18741_,
		_w18742_,
		_w18743_
	);
	LUT2 #(
		.INIT('h1)
	) name14697 (
		_w18133_,
		_w18743_,
		_w18744_
	);
	LUT2 #(
		.INIT('h2)
	) name14698 (
		_w17839_,
		_w18165_,
		_w18745_
	);
	LUT2 #(
		.INIT('h4)
	) name14699 (
		_w17929_,
		_w18745_,
		_w18746_
	);
	LUT2 #(
		.INIT('h4)
	) name14700 (
		_w18108_,
		_w18746_,
		_w18747_
	);
	LUT2 #(
		.INIT('h2)
	) name14701 (
		_w17839_,
		_w17933_,
		_w18748_
	);
	LUT2 #(
		.INIT('h4)
	) name14702 (
		_w17929_,
		_w18748_,
		_w18749_
	);
	LUT2 #(
		.INIT('h8)
	) name14703 (
		_w18153_,
		_w18749_,
		_w18750_
	);
	LUT2 #(
		.INIT('h2)
	) name14704 (
		_w17839_,
		_w18102_,
		_w18751_
	);
	LUT2 #(
		.INIT('h4)
	) name14705 (
		_w17929_,
		_w18751_,
		_w18752_
	);
	LUT2 #(
		.INIT('h8)
	) name14706 (
		_w18178_,
		_w18752_,
		_w18753_
	);
	LUT2 #(
		.INIT('h8)
	) name14707 (
		_w17929_,
		_w18183_,
		_w18754_
	);
	LUT2 #(
		.INIT('h8)
	) name14708 (
		_w18089_,
		_w18754_,
		_w18755_
	);
	LUT2 #(
		.INIT('h4)
	) name14709 (
		_w17929_,
		_w18187_,
		_w18756_
	);
	LUT2 #(
		.INIT('h8)
	) name14710 (
		_w17921_,
		_w18756_,
		_w18757_
	);
	LUT2 #(
		.INIT('h2)
	) name14711 (
		_w17839_,
		_w18135_,
		_w18758_
	);
	LUT2 #(
		.INIT('h4)
	) name14712 (
		_w17929_,
		_w18758_,
		_w18759_
	);
	LUT2 #(
		.INIT('h4)
	) name14713 (
		_w18091_,
		_w18759_,
		_w18760_
	);
	LUT2 #(
		.INIT('h4)
	) name14714 (
		_w17929_,
		_w17986_,
		_w18761_
	);
	LUT2 #(
		.INIT('h8)
	) name14715 (
		_w18115_,
		_w18761_,
		_w18762_
	);
	LUT2 #(
		.INIT('h8)
	) name14716 (
		_w17929_,
		_w18124_,
		_w18763_
	);
	LUT2 #(
		.INIT('h8)
	) name14717 (
		_w18106_,
		_w18763_,
		_w18764_
	);
	LUT2 #(
		.INIT('h2)
	) name14718 (
		_w17839_,
		_w18175_,
		_w18765_
	);
	LUT2 #(
		.INIT('h4)
	) name14719 (
		_w17929_,
		_w18765_,
		_w18766_
	);
	LUT2 #(
		.INIT('h8)
	) name14720 (
		_w18055_,
		_w18766_,
		_w18767_
	);
	LUT2 #(
		.INIT('h8)
	) name14721 (
		_w18139_,
		_w18765_,
		_w18768_
	);
	LUT2 #(
		.INIT('h8)
	) name14722 (
		_w18043_,
		_w18115_,
		_w18769_
	);
	LUT2 #(
		.INIT('h8)
	) name14723 (
		_w17959_,
		_w18112_,
		_w18770_
	);
	LUT2 #(
		.INIT('h8)
	) name14724 (
		_w17915_,
		_w18756_,
		_w18771_
	);
	LUT2 #(
		.INIT('h2)
	) name14725 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11311_,
		_w18772_
	);
	LUT2 #(
		.INIT('h8)
	) name14726 (
		_w18107_,
		_w18763_,
		_w18773_
	);
	LUT2 #(
		.INIT('h8)
	) name14727 (
		_w17929_,
		_w18055_,
		_w18774_
	);
	LUT2 #(
		.INIT('h1)
	) name14728 (
		_w18071_,
		_w18774_,
		_w18775_
	);
	LUT2 #(
		.INIT('h1)
	) name14729 (
		_w17924_,
		_w18775_,
		_w18776_
	);
	LUT2 #(
		.INIT('h4)
	) name14730 (
		_w17933_,
		_w18070_,
		_w18777_
	);
	LUT2 #(
		.INIT('h1)
	) name14731 (
		_w18776_,
		_w18777_,
		_w18778_
	);
	LUT2 #(
		.INIT('h2)
	) name14732 (
		_w17839_,
		_w18778_,
		_w18779_
	);
	LUT2 #(
		.INIT('h8)
	) name14733 (
		_w17931_,
		_w18056_,
		_w18780_
	);
	LUT2 #(
		.INIT('h1)
	) name14734 (
		_w17980_,
		_w18780_,
		_w18781_
	);
	LUT2 #(
		.INIT('h2)
	) name14735 (
		_w18088_,
		_w18781_,
		_w18782_
	);
	LUT2 #(
		.INIT('h8)
	) name14736 (
		_w17965_,
		_w18021_,
		_w18783_
	);
	LUT2 #(
		.INIT('h8)
	) name14737 (
		_w18179_,
		_w18752_,
		_w18784_
	);
	LUT2 #(
		.INIT('h8)
	) name14738 (
		_w17965_,
		_w18056_,
		_w18785_
	);
	LUT2 #(
		.INIT('h8)
	) name14739 (
		_w17945_,
		_w18150_,
		_w18786_
	);
	LUT2 #(
		.INIT('h4)
	) name14740 (
		_w17929_,
		_w18026_,
		_w18787_
	);
	LUT2 #(
		.INIT('h1)
	) name14741 (
		_w18010_,
		_w18023_,
		_w18788_
	);
	LUT2 #(
		.INIT('h4)
	) name14742 (
		_w18787_,
		_w18788_,
		_w18789_
	);
	LUT2 #(
		.INIT('h4)
	) name14743 (
		_w18786_,
		_w18789_,
		_w18790_
	);
	LUT2 #(
		.INIT('h4)
	) name14744 (
		_w18785_,
		_w18790_,
		_w18791_
	);
	LUT2 #(
		.INIT('h2)
	) name14745 (
		_w18148_,
		_w18170_,
		_w18792_
	);
	LUT2 #(
		.INIT('h8)
	) name14746 (
		_w17954_,
		_w17979_,
		_w18793_
	);
	LUT2 #(
		.INIT('h1)
	) name14747 (
		_w18151_,
		_w18793_,
		_w18794_
	);
	LUT2 #(
		.INIT('h2)
	) name14748 (
		_w17945_,
		_w18794_,
		_w18795_
	);
	LUT2 #(
		.INIT('h2)
	) name14749 (
		_w18015_,
		_w18795_,
		_w18796_
	);
	LUT2 #(
		.INIT('h4)
	) name14750 (
		_w18018_,
		_w18796_,
		_w18797_
	);
	LUT2 #(
		.INIT('h1)
	) name14751 (
		_w17964_,
		_w18085_,
		_w18798_
	);
	LUT2 #(
		.INIT('h8)
	) name14752 (
		_w18797_,
		_w18798_,
		_w18799_
	);
	LUT2 #(
		.INIT('h4)
	) name14753 (
		_w18060_,
		_w18799_,
		_w18800_
	);
	LUT2 #(
		.INIT('h1)
	) name14754 (
		_w18002_,
		_w18772_,
		_w18801_
	);
	LUT2 #(
		.INIT('h1)
	) name14755 (
		_w18750_,
		_w18753_,
		_w18802_
	);
	LUT2 #(
		.INIT('h1)
	) name14756 (
		_w18755_,
		_w18757_,
		_w18803_
	);
	LUT2 #(
		.INIT('h1)
	) name14757 (
		_w18764_,
		_w18767_,
		_w18804_
	);
	LUT2 #(
		.INIT('h8)
	) name14758 (
		_w18803_,
		_w18804_,
		_w18805_
	);
	LUT2 #(
		.INIT('h8)
	) name14759 (
		_w18801_,
		_w18802_,
		_w18806_
	);
	LUT2 #(
		.INIT('h1)
	) name14760 (
		_w18762_,
		_w18770_,
		_w18807_
	);
	LUT2 #(
		.INIT('h1)
	) name14761 (
		_w18771_,
		_w18773_,
		_w18808_
	);
	LUT2 #(
		.INIT('h1)
	) name14762 (
		_w18783_,
		_w18784_,
		_w18809_
	);
	LUT2 #(
		.INIT('h4)
	) name14763 (
		_w18792_,
		_w18809_,
		_w18810_
	);
	LUT2 #(
		.INIT('h8)
	) name14764 (
		_w18807_,
		_w18808_,
		_w18811_
	);
	LUT2 #(
		.INIT('h8)
	) name14765 (
		_w18805_,
		_w18806_,
		_w18812_
	);
	LUT2 #(
		.INIT('h8)
	) name14766 (
		_w17978_,
		_w18054_,
		_w18813_
	);
	LUT2 #(
		.INIT('h1)
	) name14767 (
		_w18723_,
		_w18733_,
		_w18814_
	);
	LUT2 #(
		.INIT('h1)
	) name14768 (
		_w18739_,
		_w18744_,
		_w18815_
	);
	LUT2 #(
		.INIT('h1)
	) name14769 (
		_w18747_,
		_w18760_,
		_w18816_
	);
	LUT2 #(
		.INIT('h1)
	) name14770 (
		_w18768_,
		_w18769_,
		_w18817_
	);
	LUT2 #(
		.INIT('h8)
	) name14771 (
		_w18816_,
		_w18817_,
		_w18818_
	);
	LUT2 #(
		.INIT('h8)
	) name14772 (
		_w18814_,
		_w18815_,
		_w18819_
	);
	LUT2 #(
		.INIT('h8)
	) name14773 (
		_w18812_,
		_w18813_,
		_w18820_
	);
	LUT2 #(
		.INIT('h8)
	) name14774 (
		_w18810_,
		_w18811_,
		_w18821_
	);
	LUT2 #(
		.INIT('h1)
	) name14775 (
		_w18721_,
		_w18782_,
		_w18822_
	);
	LUT2 #(
		.INIT('h8)
	) name14776 (
		_w18821_,
		_w18822_,
		_w18823_
	);
	LUT2 #(
		.INIT('h8)
	) name14777 (
		_w18819_,
		_w18820_,
		_w18824_
	);
	LUT2 #(
		.INIT('h8)
	) name14778 (
		_w18738_,
		_w18818_,
		_w18825_
	);
	LUT2 #(
		.INIT('h8)
	) name14779 (
		_w18824_,
		_w18825_,
		_w18826_
	);
	LUT2 #(
		.INIT('h4)
	) name14780 (
		_w18779_,
		_w18823_,
		_w18827_
	);
	LUT2 #(
		.INIT('h8)
	) name14781 (
		_w18826_,
		_w18827_,
		_w18828_
	);
	LUT2 #(
		.INIT('h8)
	) name14782 (
		_w18731_,
		_w18791_,
		_w18829_
	);
	LUT2 #(
		.INIT('h8)
	) name14783 (
		_w18828_,
		_w18829_,
		_w18830_
	);
	LUT2 #(
		.INIT('h8)
	) name14784 (
		_w18800_,
		_w18830_,
		_w18831_
	);
	LUT2 #(
		.INIT('h4)
	) name14785 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w18831_,
		_w18832_
	);
	LUT2 #(
		.INIT('h1)
	) name14786 (
		_w18718_,
		_w18832_,
		_w18833_
	);
	LUT2 #(
		.INIT('h2)
	) name14787 (
		_w18717_,
		_w18833_,
		_w18834_
	);
	LUT2 #(
		.INIT('h1)
	) name14788 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[6]/P0001 ,
		_w18717_,
		_w18835_
	);
	LUT2 #(
		.INIT('h1)
	) name14789 (
		_w18834_,
		_w18835_,
		_w18836_
	);
	LUT2 #(
		.INIT('h8)
	) name14790 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w4118_,
		_w18837_
	);
	LUT2 #(
		.INIT('h1)
	) name14791 (
		_w6023_,
		_w6108_,
		_w18838_
	);
	LUT2 #(
		.INIT('h8)
	) name14792 (
		_w6022_,
		_w6117_,
		_w18839_
	);
	LUT2 #(
		.INIT('h1)
	) name14793 (
		_w13577_,
		_w18839_,
		_w18840_
	);
	LUT2 #(
		.INIT('h4)
	) name14794 (
		_w14728_,
		_w18840_,
		_w18841_
	);
	LUT2 #(
		.INIT('h8)
	) name14795 (
		_w18838_,
		_w18841_,
		_w18842_
	);
	LUT2 #(
		.INIT('h1)
	) name14796 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w18843_
	);
	LUT2 #(
		.INIT('h1)
	) name14797 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w18844_
	);
	LUT2 #(
		.INIT('h8)
	) name14798 (
		_w18843_,
		_w18844_,
		_w18845_
	);
	LUT2 #(
		.INIT('h1)
	) name14799 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w18845_,
		_w18846_
	);
	LUT2 #(
		.INIT('h4)
	) name14800 (
		_w18842_,
		_w18846_,
		_w18847_
	);
	LUT2 #(
		.INIT('h4)
	) name14801 (
		_w4117_,
		_w18847_,
		_w18848_
	);
	LUT2 #(
		.INIT('h2)
	) name14802 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		_w6023_,
		_w18849_
	);
	LUT2 #(
		.INIT('h2)
	) name14803 (
		_w4116_,
		_w18849_,
		_w18850_
	);
	LUT2 #(
		.INIT('h8)
	) name14804 (
		_w18848_,
		_w18850_,
		_w18851_
	);
	LUT2 #(
		.INIT('h1)
	) name14805 (
		_w18837_,
		_w18851_,
		_w18852_
	);
	LUT2 #(
		.INIT('h2)
	) name14806 (
		_w13805_,
		_w18698_,
		_w18853_
	);
	LUT2 #(
		.INIT('h2)
	) name14807 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[13]/P0001 ,
		_w13805_,
		_w18854_
	);
	LUT2 #(
		.INIT('h1)
	) name14808 (
		_w18853_,
		_w18854_,
		_w18855_
	);
	LUT2 #(
		.INIT('h8)
	) name14809 (
		\sice_ICYC_reg[0]/NET0131 ,
		\sice_ICYC_reg[1]/NET0131 ,
		_w18856_
	);
	LUT2 #(
		.INIT('h8)
	) name14810 (
		\sice_ICYC_reg[2]/NET0131 ,
		_w18856_,
		_w18857_
	);
	LUT2 #(
		.INIT('h8)
	) name14811 (
		\sice_ICYC_reg[3]/NET0131 ,
		_w18857_,
		_w18858_
	);
	LUT2 #(
		.INIT('h8)
	) name14812 (
		\sice_ICYC_reg[4]/NET0131 ,
		_w18858_,
		_w18859_
	);
	LUT2 #(
		.INIT('h8)
	) name14813 (
		\sice_ICYC_reg[5]/NET0131 ,
		_w18859_,
		_w18860_
	);
	LUT2 #(
		.INIT('h8)
	) name14814 (
		\sice_ICYC_reg[6]/NET0131 ,
		_w18860_,
		_w18861_
	);
	LUT2 #(
		.INIT('h1)
	) name14815 (
		\sice_ICYC_reg[7]/NET0131 ,
		_w18861_,
		_w18862_
	);
	LUT2 #(
		.INIT('h8)
	) name14816 (
		\sice_ICYC_reg[7]/NET0131 ,
		_w18861_,
		_w18863_
	);
	LUT2 #(
		.INIT('h1)
	) name14817 (
		_w18862_,
		_w18863_,
		_w18864_
	);
	LUT2 #(
		.INIT('h8)
	) name14818 (
		\sice_IIRC_reg[0]/NET0131 ,
		\sice_IIRC_reg[1]/NET0131 ,
		_w18865_
	);
	LUT2 #(
		.INIT('h8)
	) name14819 (
		\sice_IIRC_reg[2]/NET0131 ,
		_w18865_,
		_w18866_
	);
	LUT2 #(
		.INIT('h8)
	) name14820 (
		\sice_IIRC_reg[3]/NET0131 ,
		_w18866_,
		_w18867_
	);
	LUT2 #(
		.INIT('h8)
	) name14821 (
		\sice_IIRC_reg[4]/NET0131 ,
		_w18867_,
		_w18868_
	);
	LUT2 #(
		.INIT('h8)
	) name14822 (
		\sice_IIRC_reg[5]/NET0131 ,
		_w18868_,
		_w18869_
	);
	LUT2 #(
		.INIT('h8)
	) name14823 (
		\sice_IIRC_reg[6]/NET0131 ,
		_w18869_,
		_w18870_
	);
	LUT2 #(
		.INIT('h8)
	) name14824 (
		\sice_IIRC_reg[7]/NET0131 ,
		_w18870_,
		_w18871_
	);
	LUT2 #(
		.INIT('h1)
	) name14825 (
		\sice_IIRC_reg[7]/NET0131 ,
		_w18870_,
		_w18872_
	);
	LUT2 #(
		.INIT('h1)
	) name14826 (
		_w18871_,
		_w18872_,
		_w18873_
	);
	LUT2 #(
		.INIT('h2)
	) name14827 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[3]/P0001 ,
		_w18848_,
		_w18874_
	);
	LUT2 #(
		.INIT('h2)
	) name14828 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w18843_,
		_w18875_
	);
	LUT2 #(
		.INIT('h8)
	) name14829 (
		_w18848_,
		_w18875_,
		_w18876_
	);
	LUT2 #(
		.INIT('h1)
	) name14830 (
		_w18874_,
		_w18876_,
		_w18877_
	);
	LUT2 #(
		.INIT('h2)
	) name14831 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[2]/P0001 ,
		_w18848_,
		_w18878_
	);
	LUT2 #(
		.INIT('h2)
	) name14832 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		_w18843_,
		_w18879_
	);
	LUT2 #(
		.INIT('h8)
	) name14833 (
		_w18848_,
		_w18879_,
		_w18880_
	);
	LUT2 #(
		.INIT('h1)
	) name14834 (
		_w18878_,
		_w18880_,
		_w18881_
	);
	LUT2 #(
		.INIT('h2)
	) name14835 (
		_w17833_,
		_w18833_,
		_w18882_
	);
	LUT2 #(
		.INIT('h1)
	) name14836 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[6]/P0001 ,
		_w17833_,
		_w18883_
	);
	LUT2 #(
		.INIT('h1)
	) name14837 (
		_w18882_,
		_w18883_,
		_w18884_
	);
	LUT2 #(
		.INIT('h1)
	) name14838 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		\core_c_dec_updSR_E_reg/P0001 ,
		_w18885_
	);
	LUT2 #(
		.INIT('h2)
	) name14839 (
		_w14666_,
		_w18885_,
		_w18886_
	);
	LUT2 #(
		.INIT('h2)
	) name14840 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w18276_,
		_w18887_
	);
	LUT2 #(
		.INIT('h1)
	) name14841 (
		_w17960_,
		_w18150_,
		_w18888_
	);
	LUT2 #(
		.INIT('h2)
	) name14842 (
		_w18088_,
		_w18888_,
		_w18889_
	);
	LUT2 #(
		.INIT('h2)
	) name14843 (
		_w17971_,
		_w18082_,
		_w18890_
	);
	LUT2 #(
		.INIT('h1)
	) name14844 (
		_w17995_,
		_w18890_,
		_w18891_
	);
	LUT2 #(
		.INIT('h8)
	) name14845 (
		_w18796_,
		_w18891_,
		_w18892_
	);
	LUT2 #(
		.INIT('h8)
	) name14846 (
		_w17958_,
		_w17989_,
		_w18893_
	);
	LUT2 #(
		.INIT('h4)
	) name14847 (
		_w17931_,
		_w18056_,
		_w18894_
	);
	LUT2 #(
		.INIT('h1)
	) name14848 (
		_w18893_,
		_w18894_,
		_w18895_
	);
	LUT2 #(
		.INIT('h2)
	) name14849 (
		_w18751_,
		_w18895_,
		_w18896_
	);
	LUT2 #(
		.INIT('h4)
	) name14850 (
		_w17931_,
		_w17968_,
		_w18897_
	);
	LUT2 #(
		.INIT('h1)
	) name14851 (
		_w18027_,
		_w18897_,
		_w18898_
	);
	LUT2 #(
		.INIT('h2)
	) name14852 (
		_w18115_,
		_w18898_,
		_w18899_
	);
	LUT2 #(
		.INIT('h8)
	) name14853 (
		_w17959_,
		_w17965_,
		_w18900_
	);
	LUT2 #(
		.INIT('h1)
	) name14854 (
		_w17972_,
		_w18900_,
		_w18901_
	);
	LUT2 #(
		.INIT('h1)
	) name14855 (
		_w18143_,
		_w18783_,
		_w18902_
	);
	LUT2 #(
		.INIT('h8)
	) name14856 (
		_w18901_,
		_w18902_,
		_w18903_
	);
	LUT2 #(
		.INIT('h8)
	) name14857 (
		_w18789_,
		_w18903_,
		_w18904_
	);
	LUT2 #(
		.INIT('h2)
	) name14858 (
		_w17931_,
		_w18110_,
		_w18905_
	);
	LUT2 #(
		.INIT('h4)
	) name14859 (
		_w18079_,
		_w18905_,
		_w18906_
	);
	LUT2 #(
		.INIT('h1)
	) name14860 (
		_w17952_,
		_w18001_,
		_w18907_
	);
	LUT2 #(
		.INIT('h1)
	) name14861 (
		_w18743_,
		_w18907_,
		_w18908_
	);
	LUT2 #(
		.INIT('h1)
	) name14862 (
		_w18029_,
		_w18036_,
		_w18909_
	);
	LUT2 #(
		.INIT('h2)
	) name14863 (
		_w18766_,
		_w18909_,
		_w18910_
	);
	LUT2 #(
		.INIT('h2)
	) name14864 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11315_,
		_w18911_
	);
	LUT2 #(
		.INIT('h1)
	) name14865 (
		_w17955_,
		_w18072_,
		_w18912_
	);
	LUT2 #(
		.INIT('h2)
	) name14866 (
		_w18746_,
		_w18912_,
		_w18913_
	);
	LUT2 #(
		.INIT('h1)
	) name14867 (
		_w18033_,
		_w18067_,
		_w18914_
	);
	LUT2 #(
		.INIT('h1)
	) name14868 (
		_w18754_,
		_w18759_,
		_w18915_
	);
	LUT2 #(
		.INIT('h1)
	) name14869 (
		_w18914_,
		_w18915_,
		_w18916_
	);
	LUT2 #(
		.INIT('h2)
	) name14870 (
		_w18763_,
		_w18912_,
		_w18917_
	);
	LUT2 #(
		.INIT('h1)
	) name14871 (
		_w18039_,
		_w18191_,
		_w18918_
	);
	LUT2 #(
		.INIT('h1)
	) name14872 (
		_w18722_,
		_w18756_,
		_w18919_
	);
	LUT2 #(
		.INIT('h1)
	) name14873 (
		_w18918_,
		_w18919_,
		_w18920_
	);
	LUT2 #(
		.INIT('h4)
	) name14874 (
		_w18079_,
		_w18749_,
		_w18921_
	);
	LUT2 #(
		.INIT('h2)
	) name14875 (
		_w17931_,
		_w18909_,
		_w18922_
	);
	LUT2 #(
		.INIT('h4)
	) name14876 (
		_w17924_,
		_w18922_,
		_w18923_
	);
	LUT2 #(
		.INIT('h4)
	) name14877 (
		_w17998_,
		_w18171_,
		_w18924_
	);
	LUT2 #(
		.INIT('h1)
	) name14878 (
		_w18018_,
		_w18911_,
		_w18925_
	);
	LUT2 #(
		.INIT('h4)
	) name14879 (
		_w18906_,
		_w18925_,
		_w18926_
	);
	LUT2 #(
		.INIT('h1)
	) name14880 (
		_w18908_,
		_w18910_,
		_w18927_
	);
	LUT2 #(
		.INIT('h1)
	) name14881 (
		_w18913_,
		_w18916_,
		_w18928_
	);
	LUT2 #(
		.INIT('h1)
	) name14882 (
		_w18917_,
		_w18920_,
		_w18929_
	);
	LUT2 #(
		.INIT('h4)
	) name14883 (
		_w18921_,
		_w18929_,
		_w18930_
	);
	LUT2 #(
		.INIT('h8)
	) name14884 (
		_w18927_,
		_w18928_,
		_w18931_
	);
	LUT2 #(
		.INIT('h4)
	) name14885 (
		_w18889_,
		_w18926_,
		_w18932_
	);
	LUT2 #(
		.INIT('h1)
	) name14886 (
		_w18896_,
		_w18899_,
		_w18933_
	);
	LUT2 #(
		.INIT('h1)
	) name14887 (
		_w18923_,
		_w18924_,
		_w18934_
	);
	LUT2 #(
		.INIT('h8)
	) name14888 (
		_w18933_,
		_w18934_,
		_w18935_
	);
	LUT2 #(
		.INIT('h8)
	) name14889 (
		_w18931_,
		_w18932_,
		_w18936_
	);
	LUT2 #(
		.INIT('h8)
	) name14890 (
		_w18930_,
		_w18936_,
		_w18937_
	);
	LUT2 #(
		.INIT('h8)
	) name14891 (
		_w18892_,
		_w18935_,
		_w18938_
	);
	LUT2 #(
		.INIT('h8)
	) name14892 (
		_w18904_,
		_w18938_,
		_w18939_
	);
	LUT2 #(
		.INIT('h8)
	) name14893 (
		_w18937_,
		_w18939_,
		_w18940_
	);
	LUT2 #(
		.INIT('h4)
	) name14894 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w18940_,
		_w18941_
	);
	LUT2 #(
		.INIT('h1)
	) name14895 (
		_w18887_,
		_w18941_,
		_w18942_
	);
	LUT2 #(
		.INIT('h2)
	) name14896 (
		_w18886_,
		_w18942_,
		_w18943_
	);
	LUT2 #(
		.INIT('h1)
	) name14897 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[6]/P0001 ,
		_w18886_,
		_w18944_
	);
	LUT2 #(
		.INIT('h1)
	) name14898 (
		_w18943_,
		_w18944_,
		_w18945_
	);
	LUT2 #(
		.INIT('h8)
	) name14899 (
		_w7270_,
		_w18227_,
		_w18946_
	);
	LUT2 #(
		.INIT('h2)
	) name14900 (
		\sport1_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w18946_,
		_w18947_
	);
	LUT2 #(
		.INIT('h4)
	) name14901 (
		_w12688_,
		_w18946_,
		_w18948_
	);
	LUT2 #(
		.INIT('h8)
	) name14902 (
		_w11265_,
		_w18948_,
		_w18949_
	);
	LUT2 #(
		.INIT('h1)
	) name14903 (
		_w18947_,
		_w18949_,
		_w18950_
	);
	LUT2 #(
		.INIT('h2)
	) name14904 (
		\sport1_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w18946_,
		_w18951_
	);
	LUT2 #(
		.INIT('h8)
	) name14905 (
		_w11525_,
		_w18948_,
		_w18952_
	);
	LUT2 #(
		.INIT('h1)
	) name14906 (
		_w18951_,
		_w18952_,
		_w18953_
	);
	LUT2 #(
		.INIT('h2)
	) name14907 (
		\sport1_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w18946_,
		_w18954_
	);
	LUT2 #(
		.INIT('h8)
	) name14908 (
		_w10911_,
		_w18948_,
		_w18955_
	);
	LUT2 #(
		.INIT('h1)
	) name14909 (
		_w18954_,
		_w18955_,
		_w18956_
	);
	LUT2 #(
		.INIT('h4)
	) name14910 (
		_w7340_,
		_w18946_,
		_w18957_
	);
	LUT2 #(
		.INIT('h1)
	) name14911 (
		\sport1_regs_MWORDreg_DO_reg[8]/NET0131 ,
		_w18946_,
		_w18958_
	);
	LUT2 #(
		.INIT('h1)
	) name14912 (
		_w18957_,
		_w18958_,
		_w18959_
	);
	LUT2 #(
		.INIT('h2)
	) name14913 (
		\sport1_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w18946_,
		_w18960_
	);
	LUT2 #(
		.INIT('h8)
	) name14914 (
		_w10069_,
		_w18948_,
		_w18961_
	);
	LUT2 #(
		.INIT('h1)
	) name14915 (
		_w18960_,
		_w18961_,
		_w18962_
	);
	LUT2 #(
		.INIT('h2)
	) name14916 (
		\sport1_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w18946_,
		_w18963_
	);
	LUT2 #(
		.INIT('h8)
	) name14917 (
		_w9435_,
		_w18948_,
		_w18964_
	);
	LUT2 #(
		.INIT('h1)
	) name14918 (
		_w18963_,
		_w18964_,
		_w18965_
	);
	LUT2 #(
		.INIT('h2)
	) name14919 (
		\sport1_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w18946_,
		_w18966_
	);
	LUT2 #(
		.INIT('h8)
	) name14920 (
		_w7607_,
		_w18948_,
		_w18967_
	);
	LUT2 #(
		.INIT('h1)
	) name14921 (
		_w18966_,
		_w18967_,
		_w18968_
	);
	LUT2 #(
		.INIT('h4)
	) name14922 (
		_w7340_,
		_w18231_,
		_w18969_
	);
	LUT2 #(
		.INIT('h1)
	) name14923 (
		\sport0_regs_MWORDreg_DO_reg[8]/NET0131 ,
		_w18231_,
		_w18970_
	);
	LUT2 #(
		.INIT('h1)
	) name14924 (
		_w18969_,
		_w18970_,
		_w18971_
	);
	LUT2 #(
		.INIT('h1)
	) name14925 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w9435_,
		_w18972_
	);
	LUT2 #(
		.INIT('h2)
	) name14926 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12802_,
		_w18973_
	);
	LUT2 #(
		.INIT('h1)
	) name14927 (
		_w18972_,
		_w18973_,
		_w18974_
	);
	LUT2 #(
		.INIT('h2)
	) name14928 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w18974_,
		_w18975_
	);
	LUT2 #(
		.INIT('h2)
	) name14929 (
		_w17930_,
		_w18082_,
		_w18976_
	);
	LUT2 #(
		.INIT('h1)
	) name14930 (
		_w18129_,
		_w18914_,
		_w18977_
	);
	LUT2 #(
		.INIT('h2)
	) name14931 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9276_,
		_w18978_
	);
	LUT2 #(
		.INIT('h1)
	) name14932 (
		_w18079_,
		_w18189_,
		_w18979_
	);
	LUT2 #(
		.INIT('h8)
	) name14933 (
		_w17954_,
		_w17989_,
		_w18980_
	);
	LUT2 #(
		.INIT('h1)
	) name14934 (
		_w18044_,
		_w18980_,
		_w18981_
	);
	LUT2 #(
		.INIT('h2)
	) name14935 (
		_w18088_,
		_w18981_,
		_w18982_
	);
	LUT2 #(
		.INIT('h1)
	) name14936 (
		_w18022_,
		_w18793_,
		_w18983_
	);
	LUT2 #(
		.INIT('h2)
	) name14937 (
		_w18765_,
		_w18983_,
		_w18984_
	);
	LUT2 #(
		.INIT('h1)
	) name14938 (
		_w17998_,
		_w18165_,
		_w18985_
	);
	LUT2 #(
		.INIT('h4)
	) name14939 (
		_w17933_,
		_w18083_,
		_w18986_
	);
	LUT2 #(
		.INIT('h1)
	) name14940 (
		_w17961_,
		_w18150_,
		_w18987_
	);
	LUT2 #(
		.INIT('h1)
	) name14941 (
		_w18114_,
		_w18987_,
		_w18988_
	);
	LUT2 #(
		.INIT('h2)
	) name14942 (
		_w18162_,
		_w18898_,
		_w18989_
	);
	LUT2 #(
		.INIT('h1)
	) name14943 (
		_w18104_,
		_w18918_,
		_w18990_
	);
	LUT2 #(
		.INIT('h1)
	) name14944 (
		_w18136_,
		_w18172_,
		_w18991_
	);
	LUT2 #(
		.INIT('h1)
	) name14945 (
		_w18909_,
		_w18991_,
		_w18992_
	);
	LUT2 #(
		.INIT('h8)
	) name14946 (
		_w17991_,
		_w18111_,
		_w18993_
	);
	LUT2 #(
		.INIT('h1)
	) name14947 (
		_w18143_,
		_w18978_,
		_w18994_
	);
	LUT2 #(
		.INIT('h8)
	) name14948 (
		_w18901_,
		_w18994_,
		_w18995_
	);
	LUT2 #(
		.INIT('h1)
	) name14949 (
		_w18976_,
		_w18977_,
		_w18996_
	);
	LUT2 #(
		.INIT('h1)
	) name14950 (
		_w18979_,
		_w18990_,
		_w18997_
	);
	LUT2 #(
		.INIT('h1)
	) name14951 (
		_w18992_,
		_w18993_,
		_w18998_
	);
	LUT2 #(
		.INIT('h8)
	) name14952 (
		_w18997_,
		_w18998_,
		_w18999_
	);
	LUT2 #(
		.INIT('h8)
	) name14953 (
		_w18995_,
		_w18996_,
		_w19000_
	);
	LUT2 #(
		.INIT('h2)
	) name14954 (
		_w18019_,
		_w18982_,
		_w19001_
	);
	LUT2 #(
		.INIT('h1)
	) name14955 (
		_w18984_,
		_w18985_,
		_w19002_
	);
	LUT2 #(
		.INIT('h1)
	) name14956 (
		_w18986_,
		_w18989_,
		_w19003_
	);
	LUT2 #(
		.INIT('h8)
	) name14957 (
		_w19002_,
		_w19003_,
		_w19004_
	);
	LUT2 #(
		.INIT('h8)
	) name14958 (
		_w19000_,
		_w19001_,
		_w19005_
	);
	LUT2 #(
		.INIT('h4)
	) name14959 (
		_w18988_,
		_w18999_,
		_w19006_
	);
	LUT2 #(
		.INIT('h8)
	) name14960 (
		_w19005_,
		_w19006_,
		_w19007_
	);
	LUT2 #(
		.INIT('h8)
	) name14961 (
		_w19004_,
		_w19007_,
		_w19008_
	);
	LUT2 #(
		.INIT('h4)
	) name14962 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w19008_,
		_w19009_
	);
	LUT2 #(
		.INIT('h1)
	) name14963 (
		_w18975_,
		_w19009_,
		_w19010_
	);
	LUT2 #(
		.INIT('h2)
	) name14964 (
		_w18886_,
		_w19010_,
		_w19011_
	);
	LUT2 #(
		.INIT('h1)
	) name14965 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[1]/P0001 ,
		_w18886_,
		_w19012_
	);
	LUT2 #(
		.INIT('h1)
	) name14966 (
		_w19011_,
		_w19012_,
		_w19013_
	);
	LUT2 #(
		.INIT('h2)
	) name14967 (
		\sport0_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w18231_,
		_w19014_
	);
	LUT2 #(
		.INIT('h4)
	) name14968 (
		_w12688_,
		_w18231_,
		_w19015_
	);
	LUT2 #(
		.INIT('h8)
	) name14969 (
		_w11265_,
		_w19015_,
		_w19016_
	);
	LUT2 #(
		.INIT('h1)
	) name14970 (
		_w19014_,
		_w19016_,
		_w19017_
	);
	LUT2 #(
		.INIT('h2)
	) name14971 (
		\sport0_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w18231_,
		_w19018_
	);
	LUT2 #(
		.INIT('h8)
	) name14972 (
		_w11525_,
		_w19015_,
		_w19019_
	);
	LUT2 #(
		.INIT('h1)
	) name14973 (
		_w19018_,
		_w19019_,
		_w19020_
	);
	LUT2 #(
		.INIT('h2)
	) name14974 (
		\sport0_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w18231_,
		_w19021_
	);
	LUT2 #(
		.INIT('h8)
	) name14975 (
		_w10911_,
		_w19015_,
		_w19022_
	);
	LUT2 #(
		.INIT('h1)
	) name14976 (
		_w19021_,
		_w19022_,
		_w19023_
	);
	LUT2 #(
		.INIT('h2)
	) name14977 (
		_w10069_,
		_w18236_,
		_w19024_
	);
	LUT2 #(
		.INIT('h2)
	) name14978 (
		_w18231_,
		_w19024_,
		_w19025_
	);
	LUT2 #(
		.INIT('h1)
	) name14979 (
		\sport0_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w18231_,
		_w19026_
	);
	LUT2 #(
		.INIT('h1)
	) name14980 (
		_w19025_,
		_w19026_,
		_w19027_
	);
	LUT2 #(
		.INIT('h2)
	) name14981 (
		\sport0_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w18231_,
		_w19028_
	);
	LUT2 #(
		.INIT('h8)
	) name14982 (
		_w9435_,
		_w19015_,
		_w19029_
	);
	LUT2 #(
		.INIT('h1)
	) name14983 (
		_w19028_,
		_w19029_,
		_w19030_
	);
	LUT2 #(
		.INIT('h2)
	) name14984 (
		\sport0_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w18231_,
		_w19031_
	);
	LUT2 #(
		.INIT('h8)
	) name14985 (
		_w7607_,
		_w19015_,
		_w19032_
	);
	LUT2 #(
		.INIT('h1)
	) name14986 (
		_w19031_,
		_w19032_,
		_w19033_
	);
	LUT2 #(
		.INIT('h2)
	) name14987 (
		_w13804_,
		_w18885_,
		_w19034_
	);
	LUT2 #(
		.INIT('h4)
	) name14988 (
		_w18942_,
		_w19034_,
		_w19035_
	);
	LUT2 #(
		.INIT('h1)
	) name14989 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[6]/P0001 ,
		_w19034_,
		_w19036_
	);
	LUT2 #(
		.INIT('h1)
	) name14990 (
		_w19035_,
		_w19036_,
		_w19037_
	);
	LUT2 #(
		.INIT('h8)
	) name14991 (
		\memc_Dread_E_reg/NET0131 ,
		_w5435_,
		_w19038_
	);
	LUT2 #(
		.INIT('h1)
	) name14992 (
		\memc_IOcmd_E_reg/NET0131 ,
		_w19038_,
		_w19039_
	);
	LUT2 #(
		.INIT('h1)
	) name14993 (
		PM_bdry_sel_pad,
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w19040_
	);
	LUT2 #(
		.INIT('h2)
	) name14994 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		_w19040_,
		_w19041_
	);
	LUT2 #(
		.INIT('h8)
	) name14995 (
		\core_c_dec_Double_E_reg/P0001 ,
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w19042_
	);
	LUT2 #(
		.INIT('h8)
	) name14996 (
		_w19041_,
		_w19042_,
		_w19043_
	);
	LUT2 #(
		.INIT('h2)
	) name14997 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4068_,
		_w19044_
	);
	LUT2 #(
		.INIT('h1)
	) name14998 (
		_w5697_,
		_w5712_,
		_w19045_
	);
	LUT2 #(
		.INIT('h1)
	) name14999 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w19045_,
		_w19046_
	);
	LUT2 #(
		.INIT('h1)
	) name15000 (
		_w19044_,
		_w19046_,
		_w19047_
	);
	LUT2 #(
		.INIT('h1)
	) name15001 (
		\core_c_psq_ECYC_reg/P0001 ,
		_w14733_,
		_w19048_
	);
	LUT2 #(
		.INIT('h4)
	) name15002 (
		_w19047_,
		_w19048_,
		_w19049_
	);
	LUT2 #(
		.INIT('h4)
	) name15003 (
		_w19043_,
		_w19049_,
		_w19050_
	);
	LUT2 #(
		.INIT('h4)
	) name15004 (
		_w14733_,
		_w19043_,
		_w19051_
	);
	LUT2 #(
		.INIT('h8)
	) name15005 (
		_w5560_,
		_w19051_,
		_w19052_
	);
	LUT2 #(
		.INIT('h8)
	) name15006 (
		_w5598_,
		_w19052_,
		_w19053_
	);
	LUT2 #(
		.INIT('h1)
	) name15007 (
		_w19050_,
		_w19053_,
		_w19054_
	);
	LUT2 #(
		.INIT('h1)
	) name15008 (
		_w19039_,
		_w19054_,
		_w19055_
	);
	LUT2 #(
		.INIT('h1)
	) name15009 (
		_w4117_,
		_w14733_,
		_w19056_
	);
	LUT2 #(
		.INIT('h2)
	) name15010 (
		\emc_DMDoe_reg/NET0131 ,
		_w19056_,
		_w19057_
	);
	LUT2 #(
		.INIT('h8)
	) name15011 (
		_w19054_,
		_w19057_,
		_w19058_
	);
	LUT2 #(
		.INIT('h1)
	) name15012 (
		_w19055_,
		_w19058_,
		_w19059_
	);
	LUT2 #(
		.INIT('h4)
	) name15013 (
		_w19010_,
		_w19034_,
		_w19060_
	);
	LUT2 #(
		.INIT('h1)
	) name15014 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[1]/P0001 ,
		_w19034_,
		_w19061_
	);
	LUT2 #(
		.INIT('h1)
	) name15015 (
		_w19060_,
		_w19061_,
		_w19062_
	);
	LUT2 #(
		.INIT('h1)
	) name15016 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w18946_,
		_w19063_
	);
	LUT2 #(
		.INIT('h1)
	) name15017 (
		_w18948_,
		_w19063_,
		_w19064_
	);
	LUT2 #(
		.INIT('h2)
	) name15018 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w18231_,
		_w19065_
	);
	LUT2 #(
		.INIT('h1)
	) name15019 (
		_w18232_,
		_w19065_,
		_w19066_
	);
	LUT2 #(
		.INIT('h4)
	) name15020 (
		\sport1_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w19067_
	);
	LUT2 #(
		.INIT('h4)
	) name15021 (
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w19068_
	);
	LUT2 #(
		.INIT('h4)
	) name15022 (
		\sport1_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w19069_
	);
	LUT2 #(
		.INIT('h2)
	) name15023 (
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w19070_
	);
	LUT2 #(
		.INIT('h2)
	) name15024 (
		\sport1_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w19071_
	);
	LUT2 #(
		.INIT('h2)
	) name15025 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w19072_
	);
	LUT2 #(
		.INIT('h2)
	) name15026 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w19073_
	);
	LUT2 #(
		.INIT('h4)
	) name15027 (
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w19074_
	);
	LUT2 #(
		.INIT('h4)
	) name15028 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w19075_
	);
	LUT2 #(
		.INIT('h2)
	) name15029 (
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w19076_
	);
	LUT2 #(
		.INIT('h4)
	) name15030 (
		\sport1_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w19077_
	);
	LUT2 #(
		.INIT('h2)
	) name15031 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w19078_
	);
	LUT2 #(
		.INIT('h4)
	) name15032 (
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w19079_
	);
	LUT2 #(
		.INIT('h2)
	) name15033 (
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w19080_
	);
	LUT2 #(
		.INIT('h1)
	) name15034 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w19081_
	);
	LUT2 #(
		.INIT('h8)
	) name15035 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w19082_
	);
	LUT2 #(
		.INIT('h1)
	) name15036 (
		_w19081_,
		_w19082_,
		_w19083_
	);
	LUT2 #(
		.INIT('h4)
	) name15037 (
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w19084_
	);
	LUT2 #(
		.INIT('h2)
	) name15038 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w19085_
	);
	LUT2 #(
		.INIT('h4)
	) name15039 (
		\sport1_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w19086_
	);
	LUT2 #(
		.INIT('h2)
	) name15040 (
		\sport1_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w19087_
	);
	LUT2 #(
		.INIT('h2)
	) name15041 (
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w19088_
	);
	LUT2 #(
		.INIT('h4)
	) name15042 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w19089_
	);
	LUT2 #(
		.INIT('h2)
	) name15043 (
		\sport1_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w19090_
	);
	LUT2 #(
		.INIT('h4)
	) name15044 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w19091_
	);
	LUT2 #(
		.INIT('h4)
	) name15045 (
		\sport1_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w19092_
	);
	LUT2 #(
		.INIT('h2)
	) name15046 (
		\sport1_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w19093_
	);
	LUT2 #(
		.INIT('h2)
	) name15047 (
		\sport1_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w19094_
	);
	LUT2 #(
		.INIT('h4)
	) name15048 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w19095_
	);
	LUT2 #(
		.INIT('h4)
	) name15049 (
		\sport1_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w19096_
	);
	LUT2 #(
		.INIT('h2)
	) name15050 (
		\sport1_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w19097_
	);
	LUT2 #(
		.INIT('h2)
	) name15051 (
		\sport1_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w19098_
	);
	LUT2 #(
		.INIT('h4)
	) name15052 (
		\sport1_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w19099_
	);
	LUT2 #(
		.INIT('h1)
	) name15053 (
		_w19067_,
		_w19068_,
		_w19100_
	);
	LUT2 #(
		.INIT('h1)
	) name15054 (
		_w19069_,
		_w19070_,
		_w19101_
	);
	LUT2 #(
		.INIT('h1)
	) name15055 (
		_w19071_,
		_w19072_,
		_w19102_
	);
	LUT2 #(
		.INIT('h1)
	) name15056 (
		_w19073_,
		_w19074_,
		_w19103_
	);
	LUT2 #(
		.INIT('h1)
	) name15057 (
		_w19075_,
		_w19076_,
		_w19104_
	);
	LUT2 #(
		.INIT('h1)
	) name15058 (
		_w19077_,
		_w19078_,
		_w19105_
	);
	LUT2 #(
		.INIT('h1)
	) name15059 (
		_w19079_,
		_w19080_,
		_w19106_
	);
	LUT2 #(
		.INIT('h1)
	) name15060 (
		_w19084_,
		_w19085_,
		_w19107_
	);
	LUT2 #(
		.INIT('h1)
	) name15061 (
		_w19086_,
		_w19087_,
		_w19108_
	);
	LUT2 #(
		.INIT('h1)
	) name15062 (
		_w19088_,
		_w19089_,
		_w19109_
	);
	LUT2 #(
		.INIT('h1)
	) name15063 (
		_w19090_,
		_w19091_,
		_w19110_
	);
	LUT2 #(
		.INIT('h1)
	) name15064 (
		_w19092_,
		_w19093_,
		_w19111_
	);
	LUT2 #(
		.INIT('h1)
	) name15065 (
		_w19094_,
		_w19095_,
		_w19112_
	);
	LUT2 #(
		.INIT('h1)
	) name15066 (
		_w19096_,
		_w19097_,
		_w19113_
	);
	LUT2 #(
		.INIT('h1)
	) name15067 (
		_w19098_,
		_w19099_,
		_w19114_
	);
	LUT2 #(
		.INIT('h8)
	) name15068 (
		_w19113_,
		_w19114_,
		_w19115_
	);
	LUT2 #(
		.INIT('h8)
	) name15069 (
		_w19111_,
		_w19112_,
		_w19116_
	);
	LUT2 #(
		.INIT('h8)
	) name15070 (
		_w19109_,
		_w19110_,
		_w19117_
	);
	LUT2 #(
		.INIT('h8)
	) name15071 (
		_w19107_,
		_w19108_,
		_w19118_
	);
	LUT2 #(
		.INIT('h8)
	) name15072 (
		_w19105_,
		_w19106_,
		_w19119_
	);
	LUT2 #(
		.INIT('h8)
	) name15073 (
		_w19103_,
		_w19104_,
		_w19120_
	);
	LUT2 #(
		.INIT('h8)
	) name15074 (
		_w19101_,
		_w19102_,
		_w19121_
	);
	LUT2 #(
		.INIT('h4)
	) name15075 (
		_w19083_,
		_w19100_,
		_w19122_
	);
	LUT2 #(
		.INIT('h8)
	) name15076 (
		_w19121_,
		_w19122_,
		_w19123_
	);
	LUT2 #(
		.INIT('h8)
	) name15077 (
		_w19119_,
		_w19120_,
		_w19124_
	);
	LUT2 #(
		.INIT('h8)
	) name15078 (
		_w19117_,
		_w19118_,
		_w19125_
	);
	LUT2 #(
		.INIT('h8)
	) name15079 (
		_w19115_,
		_w19116_,
		_w19126_
	);
	LUT2 #(
		.INIT('h8)
	) name15080 (
		_w19125_,
		_w19126_,
		_w19127_
	);
	LUT2 #(
		.INIT('h8)
	) name15081 (
		_w19123_,
		_w19124_,
		_w19128_
	);
	LUT2 #(
		.INIT('h8)
	) name15082 (
		_w19127_,
		_w19128_,
		_w19129_
	);
	LUT2 #(
		.INIT('h2)
	) name15083 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w19129_,
		_w19130_
	);
	LUT2 #(
		.INIT('h1)
	) name15084 (
		\sport1_cfg_SCLKi_h_reg/NET0131 ,
		_w19130_,
		_w19131_
	);
	LUT2 #(
		.INIT('h8)
	) name15085 (
		\sport1_cfg_SCLKi_h_reg/NET0131 ,
		_w19130_,
		_w19132_
	);
	LUT2 #(
		.INIT('h1)
	) name15086 (
		_w19131_,
		_w19132_,
		_w19133_
	);
	LUT2 #(
		.INIT('h4)
	) name15087 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w19134_
	);
	LUT2 #(
		.INIT('h4)
	) name15088 (
		\sport0_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w19135_
	);
	LUT2 #(
		.INIT('h4)
	) name15089 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w19136_
	);
	LUT2 #(
		.INIT('h2)
	) name15090 (
		\sport0_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w19137_
	);
	LUT2 #(
		.INIT('h2)
	) name15091 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w19138_
	);
	LUT2 #(
		.INIT('h2)
	) name15092 (
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w19139_
	);
	LUT2 #(
		.INIT('h2)
	) name15093 (
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w19140_
	);
	LUT2 #(
		.INIT('h4)
	) name15094 (
		\sport0_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w19141_
	);
	LUT2 #(
		.INIT('h4)
	) name15095 (
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w19142_
	);
	LUT2 #(
		.INIT('h2)
	) name15096 (
		\sport0_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w19143_
	);
	LUT2 #(
		.INIT('h4)
	) name15097 (
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w19144_
	);
	LUT2 #(
		.INIT('h2)
	) name15098 (
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w19145_
	);
	LUT2 #(
		.INIT('h4)
	) name15099 (
		\sport0_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w19146_
	);
	LUT2 #(
		.INIT('h2)
	) name15100 (
		\sport0_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w19147_
	);
	LUT2 #(
		.INIT('h1)
	) name15101 (
		\sport0_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w19148_
	);
	LUT2 #(
		.INIT('h8)
	) name15102 (
		\sport0_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w19149_
	);
	LUT2 #(
		.INIT('h1)
	) name15103 (
		_w19148_,
		_w19149_,
		_w19150_
	);
	LUT2 #(
		.INIT('h4)
	) name15104 (
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w19151_
	);
	LUT2 #(
		.INIT('h2)
	) name15105 (
		\sport0_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w19152_
	);
	LUT2 #(
		.INIT('h4)
	) name15106 (
		\sport0_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w19153_
	);
	LUT2 #(
		.INIT('h2)
	) name15107 (
		\sport0_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w19154_
	);
	LUT2 #(
		.INIT('h2)
	) name15108 (
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w19155_
	);
	LUT2 #(
		.INIT('h4)
	) name15109 (
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w19156_
	);
	LUT2 #(
		.INIT('h2)
	) name15110 (
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w19157_
	);
	LUT2 #(
		.INIT('h4)
	) name15111 (
		\sport0_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w19158_
	);
	LUT2 #(
		.INIT('h4)
	) name15112 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w19159_
	);
	LUT2 #(
		.INIT('h2)
	) name15113 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w19160_
	);
	LUT2 #(
		.INIT('h2)
	) name15114 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w19161_
	);
	LUT2 #(
		.INIT('h4)
	) name15115 (
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w19162_
	);
	LUT2 #(
		.INIT('h4)
	) name15116 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w19163_
	);
	LUT2 #(
		.INIT('h2)
	) name15117 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w19164_
	);
	LUT2 #(
		.INIT('h2)
	) name15118 (
		\sport0_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w19165_
	);
	LUT2 #(
		.INIT('h4)
	) name15119 (
		\sport0_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w19166_
	);
	LUT2 #(
		.INIT('h1)
	) name15120 (
		_w19134_,
		_w19135_,
		_w19167_
	);
	LUT2 #(
		.INIT('h1)
	) name15121 (
		_w19136_,
		_w19137_,
		_w19168_
	);
	LUT2 #(
		.INIT('h1)
	) name15122 (
		_w19138_,
		_w19139_,
		_w19169_
	);
	LUT2 #(
		.INIT('h1)
	) name15123 (
		_w19140_,
		_w19141_,
		_w19170_
	);
	LUT2 #(
		.INIT('h1)
	) name15124 (
		_w19142_,
		_w19143_,
		_w19171_
	);
	LUT2 #(
		.INIT('h1)
	) name15125 (
		_w19144_,
		_w19145_,
		_w19172_
	);
	LUT2 #(
		.INIT('h1)
	) name15126 (
		_w19146_,
		_w19147_,
		_w19173_
	);
	LUT2 #(
		.INIT('h1)
	) name15127 (
		_w19151_,
		_w19152_,
		_w19174_
	);
	LUT2 #(
		.INIT('h1)
	) name15128 (
		_w19153_,
		_w19154_,
		_w19175_
	);
	LUT2 #(
		.INIT('h1)
	) name15129 (
		_w19155_,
		_w19156_,
		_w19176_
	);
	LUT2 #(
		.INIT('h1)
	) name15130 (
		_w19157_,
		_w19158_,
		_w19177_
	);
	LUT2 #(
		.INIT('h1)
	) name15131 (
		_w19159_,
		_w19160_,
		_w19178_
	);
	LUT2 #(
		.INIT('h1)
	) name15132 (
		_w19161_,
		_w19162_,
		_w19179_
	);
	LUT2 #(
		.INIT('h1)
	) name15133 (
		_w19163_,
		_w19164_,
		_w19180_
	);
	LUT2 #(
		.INIT('h1)
	) name15134 (
		_w19165_,
		_w19166_,
		_w19181_
	);
	LUT2 #(
		.INIT('h8)
	) name15135 (
		_w19180_,
		_w19181_,
		_w19182_
	);
	LUT2 #(
		.INIT('h8)
	) name15136 (
		_w19178_,
		_w19179_,
		_w19183_
	);
	LUT2 #(
		.INIT('h8)
	) name15137 (
		_w19176_,
		_w19177_,
		_w19184_
	);
	LUT2 #(
		.INIT('h8)
	) name15138 (
		_w19174_,
		_w19175_,
		_w19185_
	);
	LUT2 #(
		.INIT('h8)
	) name15139 (
		_w19172_,
		_w19173_,
		_w19186_
	);
	LUT2 #(
		.INIT('h8)
	) name15140 (
		_w19170_,
		_w19171_,
		_w19187_
	);
	LUT2 #(
		.INIT('h8)
	) name15141 (
		_w19168_,
		_w19169_,
		_w19188_
	);
	LUT2 #(
		.INIT('h4)
	) name15142 (
		_w19150_,
		_w19167_,
		_w19189_
	);
	LUT2 #(
		.INIT('h8)
	) name15143 (
		_w19188_,
		_w19189_,
		_w19190_
	);
	LUT2 #(
		.INIT('h8)
	) name15144 (
		_w19186_,
		_w19187_,
		_w19191_
	);
	LUT2 #(
		.INIT('h8)
	) name15145 (
		_w19184_,
		_w19185_,
		_w19192_
	);
	LUT2 #(
		.INIT('h8)
	) name15146 (
		_w19182_,
		_w19183_,
		_w19193_
	);
	LUT2 #(
		.INIT('h8)
	) name15147 (
		_w19192_,
		_w19193_,
		_w19194_
	);
	LUT2 #(
		.INIT('h8)
	) name15148 (
		_w19190_,
		_w19191_,
		_w19195_
	);
	LUT2 #(
		.INIT('h8)
	) name15149 (
		_w19194_,
		_w19195_,
		_w19196_
	);
	LUT2 #(
		.INIT('h2)
	) name15150 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w19196_,
		_w19197_
	);
	LUT2 #(
		.INIT('h1)
	) name15151 (
		\sport0_cfg_SCLKi_h_reg/NET0131 ,
		_w19197_,
		_w19198_
	);
	LUT2 #(
		.INIT('h8)
	) name15152 (
		\sport0_cfg_SCLKi_h_reg/NET0131 ,
		_w19197_,
		_w19199_
	);
	LUT2 #(
		.INIT('h1)
	) name15153 (
		_w19198_,
		_w19199_,
		_w19200_
	);
	LUT2 #(
		.INIT('h8)
	) name15154 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w5951_,
		_w19201_
	);
	LUT2 #(
		.INIT('h1)
	) name15155 (
		_w18681_,
		_w19201_,
		_w19202_
	);
	LUT2 #(
		.INIT('h4)
	) name15156 (
		_w5950_,
		_w13803_,
		_w19203_
	);
	LUT2 #(
		.INIT('h8)
	) name15157 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		_w19203_,
		_w19204_
	);
	LUT2 #(
		.INIT('h2)
	) name15158 (
		_w19202_,
		_w19204_,
		_w19205_
	);
	LUT2 #(
		.INIT('h8)
	) name15159 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		_w13803_,
		_w19206_
	);
	LUT2 #(
		.INIT('h1)
	) name15160 (
		_w14494_,
		_w14534_,
		_w19207_
	);
	LUT2 #(
		.INIT('h1)
	) name15161 (
		_w14532_,
		_w19207_,
		_w19208_
	);
	LUT2 #(
		.INIT('h1)
	) name15162 (
		_w14491_,
		_w19208_,
		_w19209_
	);
	LUT2 #(
		.INIT('h2)
	) name15163 (
		_w14474_,
		_w14490_,
		_w19210_
	);
	LUT2 #(
		.INIT('h2)
	) name15164 (
		_w19208_,
		_w19210_,
		_w19211_
	);
	LUT2 #(
		.INIT('h1)
	) name15165 (
		_w13809_,
		_w19209_,
		_w19212_
	);
	LUT2 #(
		.INIT('h4)
	) name15166 (
		_w19211_,
		_w19212_,
		_w19213_
	);
	LUT2 #(
		.INIT('h8)
	) name15167 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w19213_,
		_w19214_
	);
	LUT2 #(
		.INIT('h1)
	) name15168 (
		_w13809_,
		_w19208_,
		_w19215_
	);
	LUT2 #(
		.INIT('h4)
	) name15169 (
		_w14406_,
		_w19210_,
		_w19216_
	);
	LUT2 #(
		.INIT('h2)
	) name15170 (
		_w14404_,
		_w19210_,
		_w19217_
	);
	LUT2 #(
		.INIT('h1)
	) name15171 (
		_w14491_,
		_w19216_,
		_w19218_
	);
	LUT2 #(
		.INIT('h4)
	) name15172 (
		_w19217_,
		_w19218_,
		_w19219_
	);
	LUT2 #(
		.INIT('h2)
	) name15173 (
		_w19215_,
		_w19219_,
		_w19220_
	);
	LUT2 #(
		.INIT('h4)
	) name15174 (
		_w19215_,
		_w19219_,
		_w19221_
	);
	LUT2 #(
		.INIT('h1)
	) name15175 (
		_w19220_,
		_w19221_,
		_w19222_
	);
	LUT2 #(
		.INIT('h8)
	) name15176 (
		_w19214_,
		_w19222_,
		_w19223_
	);
	LUT2 #(
		.INIT('h1)
	) name15177 (
		_w19214_,
		_w19222_,
		_w19224_
	);
	LUT2 #(
		.INIT('h1)
	) name15178 (
		_w19223_,
		_w19224_,
		_w19225_
	);
	LUT2 #(
		.INIT('h2)
	) name15179 (
		_w19206_,
		_w19225_,
		_w19226_
	);
	LUT2 #(
		.INIT('h8)
	) name15180 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w9435_,
		_w19227_
	);
	LUT2 #(
		.INIT('h8)
	) name15181 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][1]/P0001 ,
		_w14713_,
		_w19228_
	);
	LUT2 #(
		.INIT('h8)
	) name15182 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][1]/P0001 ,
		_w14702_,
		_w19229_
	);
	LUT2 #(
		.INIT('h8)
	) name15183 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001 ,
		_w14704_,
		_w19230_
	);
	LUT2 #(
		.INIT('h8)
	) name15184 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001 ,
		_w14706_,
		_w19231_
	);
	LUT2 #(
		.INIT('h8)
	) name15185 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][1]/P0001 ,
		_w14708_,
		_w19232_
	);
	LUT2 #(
		.INIT('h8)
	) name15186 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001 ,
		_w14699_,
		_w19233_
	);
	LUT2 #(
		.INIT('h8)
	) name15187 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001 ,
		_w14711_,
		_w19234_
	);
	LUT2 #(
		.INIT('h1)
	) name15188 (
		_w19228_,
		_w19229_,
		_w19235_
	);
	LUT2 #(
		.INIT('h1)
	) name15189 (
		_w19230_,
		_w19231_,
		_w19236_
	);
	LUT2 #(
		.INIT('h1)
	) name15190 (
		_w19232_,
		_w19233_,
		_w19237_
	);
	LUT2 #(
		.INIT('h4)
	) name15191 (
		_w19234_,
		_w19237_,
		_w19238_
	);
	LUT2 #(
		.INIT('h8)
	) name15192 (
		_w19235_,
		_w19236_,
		_w19239_
	);
	LUT2 #(
		.INIT('h8)
	) name15193 (
		_w19238_,
		_w19239_,
		_w19240_
	);
	LUT2 #(
		.INIT('h2)
	) name15194 (
		_w14697_,
		_w19240_,
		_w19241_
	);
	LUT2 #(
		.INIT('h1)
	) name15195 (
		_w19227_,
		_w19241_,
		_w19242_
	);
	LUT2 #(
		.INIT('h4)
	) name15196 (
		_w19226_,
		_w19242_,
		_w19243_
	);
	LUT2 #(
		.INIT('h8)
	) name15197 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w8715_,
		_w19244_
	);
	LUT2 #(
		.INIT('h8)
	) name15198 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w19245_
	);
	LUT2 #(
		.INIT('h1)
	) name15199 (
		_w19213_,
		_w19245_,
		_w19246_
	);
	LUT2 #(
		.INIT('h2)
	) name15200 (
		_w19206_,
		_w19246_,
		_w19247_
	);
	LUT2 #(
		.INIT('h8)
	) name15201 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][2]/P0001 ,
		_w14713_,
		_w19248_
	);
	LUT2 #(
		.INIT('h8)
	) name15202 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][2]/P0001 ,
		_w14702_,
		_w19249_
	);
	LUT2 #(
		.INIT('h8)
	) name15203 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001 ,
		_w14704_,
		_w19250_
	);
	LUT2 #(
		.INIT('h8)
	) name15204 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001 ,
		_w14706_,
		_w19251_
	);
	LUT2 #(
		.INIT('h8)
	) name15205 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][2]/P0001 ,
		_w14708_,
		_w19252_
	);
	LUT2 #(
		.INIT('h8)
	) name15206 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001 ,
		_w14699_,
		_w19253_
	);
	LUT2 #(
		.INIT('h8)
	) name15207 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001 ,
		_w14711_,
		_w19254_
	);
	LUT2 #(
		.INIT('h1)
	) name15208 (
		_w19248_,
		_w19249_,
		_w19255_
	);
	LUT2 #(
		.INIT('h1)
	) name15209 (
		_w19250_,
		_w19251_,
		_w19256_
	);
	LUT2 #(
		.INIT('h1)
	) name15210 (
		_w19252_,
		_w19253_,
		_w19257_
	);
	LUT2 #(
		.INIT('h4)
	) name15211 (
		_w19254_,
		_w19257_,
		_w19258_
	);
	LUT2 #(
		.INIT('h8)
	) name15212 (
		_w19255_,
		_w19256_,
		_w19259_
	);
	LUT2 #(
		.INIT('h8)
	) name15213 (
		_w19258_,
		_w19259_,
		_w19260_
	);
	LUT2 #(
		.INIT('h2)
	) name15214 (
		_w14697_,
		_w19260_,
		_w19261_
	);
	LUT2 #(
		.INIT('h1)
	) name15215 (
		_w19244_,
		_w19261_,
		_w19262_
	);
	LUT2 #(
		.INIT('h4)
	) name15216 (
		_w19247_,
		_w19262_,
		_w19263_
	);
	LUT2 #(
		.INIT('h1)
	) name15217 (
		_w19243_,
		_w19263_,
		_w19264_
	);
	LUT2 #(
		.INIT('h8)
	) name15218 (
		_w19243_,
		_w19263_,
		_w19265_
	);
	LUT2 #(
		.INIT('h1)
	) name15219 (
		_w19264_,
		_w19265_,
		_w19266_
	);
	LUT2 #(
		.INIT('h2)
	) name15220 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w19267_
	);
	LUT2 #(
		.INIT('h8)
	) name15221 (
		_w6091_,
		_w19267_,
		_w19268_
	);
	LUT2 #(
		.INIT('h4)
	) name15222 (
		_w19266_,
		_w19268_,
		_w19269_
	);
	LUT2 #(
		.INIT('h1)
	) name15223 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w19270_
	);
	LUT2 #(
		.INIT('h8)
	) name15224 (
		_w6091_,
		_w19270_,
		_w19271_
	);
	LUT2 #(
		.INIT('h8)
	) name15225 (
		_w19266_,
		_w19271_,
		_w19272_
	);
	LUT2 #(
		.INIT('h8)
	) name15226 (
		_w6095_,
		_w19267_,
		_w19273_
	);
	LUT2 #(
		.INIT('h4)
	) name15227 (
		_w14491_,
		_w19207_,
		_w19274_
	);
	LUT2 #(
		.INIT('h4)
	) name15228 (
		_w14467_,
		_w14532_,
		_w19275_
	);
	LUT2 #(
		.INIT('h1)
	) name15229 (
		_w19210_,
		_w19275_,
		_w19276_
	);
	LUT2 #(
		.INIT('h4)
	) name15230 (
		_w19274_,
		_w19276_,
		_w19277_
	);
	LUT2 #(
		.INIT('h1)
	) name15231 (
		_w13809_,
		_w19277_,
		_w19278_
	);
	LUT2 #(
		.INIT('h8)
	) name15232 (
		_w19206_,
		_w19278_,
		_w19279_
	);
	LUT2 #(
		.INIT('h8)
	) name15233 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001 ,
		_w14699_,
		_w19280_
	);
	LUT2 #(
		.INIT('h8)
	) name15234 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][3]/P0001 ,
		_w14702_,
		_w19281_
	);
	LUT2 #(
		.INIT('h8)
	) name15235 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001 ,
		_w14704_,
		_w19282_
	);
	LUT2 #(
		.INIT('h8)
	) name15236 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001 ,
		_w14706_,
		_w19283_
	);
	LUT2 #(
		.INIT('h8)
	) name15237 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][3]/P0001 ,
		_w14708_,
		_w19284_
	);
	LUT2 #(
		.INIT('h8)
	) name15238 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001 ,
		_w14711_,
		_w19285_
	);
	LUT2 #(
		.INIT('h8)
	) name15239 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][3]/P0001 ,
		_w14713_,
		_w19286_
	);
	LUT2 #(
		.INIT('h1)
	) name15240 (
		_w19280_,
		_w19281_,
		_w19287_
	);
	LUT2 #(
		.INIT('h1)
	) name15241 (
		_w19282_,
		_w19283_,
		_w19288_
	);
	LUT2 #(
		.INIT('h1)
	) name15242 (
		_w19284_,
		_w19285_,
		_w19289_
	);
	LUT2 #(
		.INIT('h4)
	) name15243 (
		_w19286_,
		_w19289_,
		_w19290_
	);
	LUT2 #(
		.INIT('h8)
	) name15244 (
		_w19287_,
		_w19288_,
		_w19291_
	);
	LUT2 #(
		.INIT('h8)
	) name15245 (
		_w19290_,
		_w19291_,
		_w19292_
	);
	LUT2 #(
		.INIT('h2)
	) name15246 (
		_w14697_,
		_w19292_,
		_w19293_
	);
	LUT2 #(
		.INIT('h8)
	) name15247 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w8113_,
		_w19294_
	);
	LUT2 #(
		.INIT('h1)
	) name15248 (
		_w19293_,
		_w19294_,
		_w19295_
	);
	LUT2 #(
		.INIT('h4)
	) name15249 (
		_w19279_,
		_w19295_,
		_w19296_
	);
	LUT2 #(
		.INIT('h8)
	) name15250 (
		_w19273_,
		_w19296_,
		_w19297_
	);
	LUT2 #(
		.INIT('h4)
	) name15251 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w19298_
	);
	LUT2 #(
		.INIT('h8)
	) name15252 (
		_w6091_,
		_w19298_,
		_w19299_
	);
	LUT2 #(
		.INIT('h4)
	) name15253 (
		_w19263_,
		_w19299_,
		_w19300_
	);
	LUT2 #(
		.INIT('h8)
	) name15254 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w19301_
	);
	LUT2 #(
		.INIT('h8)
	) name15255 (
		_w6091_,
		_w19301_,
		_w19302_
	);
	LUT2 #(
		.INIT('h8)
	) name15256 (
		_w19263_,
		_w19302_,
		_w19303_
	);
	LUT2 #(
		.INIT('h8)
	) name15257 (
		_w6095_,
		_w19270_,
		_w19304_
	);
	LUT2 #(
		.INIT('h4)
	) name15258 (
		_w19296_,
		_w19304_,
		_w19305_
	);
	LUT2 #(
		.INIT('h1)
	) name15259 (
		_w19297_,
		_w19305_,
		_w19306_
	);
	LUT2 #(
		.INIT('h4)
	) name15260 (
		_w19300_,
		_w19306_,
		_w19307_
	);
	LUT2 #(
		.INIT('h4)
	) name15261 (
		_w19303_,
		_w19307_,
		_w19308_
	);
	LUT2 #(
		.INIT('h4)
	) name15262 (
		_w19269_,
		_w19308_,
		_w19309_
	);
	LUT2 #(
		.INIT('h4)
	) name15263 (
		_w19272_,
		_w19309_,
		_w19310_
	);
	LUT2 #(
		.INIT('h1)
	) name15264 (
		_w19205_,
		_w19310_,
		_w19311_
	);
	LUT2 #(
		.INIT('h8)
	) name15265 (
		\core_eu_ea_alu_ea_dec_AMF_E_reg[4]/NET0131 ,
		_w19206_,
		_w19312_
	);
	LUT2 #(
		.INIT('h4)
	) name15266 (
		_w5950_,
		_w13811_,
		_w19313_
	);
	LUT2 #(
		.INIT('h8)
	) name15267 (
		_w19312_,
		_w19313_,
		_w19314_
	);
	LUT2 #(
		.INIT('h2)
	) name15268 (
		_w19202_,
		_w19314_,
		_w19315_
	);
	LUT2 #(
		.INIT('h1)
	) name15269 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w19301_,
		_w19316_
	);
	LUT2 #(
		.INIT('h2)
	) name15270 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w19298_,
		_w19317_
	);
	LUT2 #(
		.INIT('h1)
	) name15271 (
		_w19316_,
		_w19317_,
		_w19318_
	);
	LUT2 #(
		.INIT('h8)
	) name15272 (
		_w19315_,
		_w19318_,
		_w19319_
	);
	LUT2 #(
		.INIT('h8)
	) name15273 (
		_w13838_,
		_w19312_,
		_w19320_
	);
	LUT2 #(
		.INIT('h8)
	) name15274 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w10069_,
		_w19321_
	);
	LUT2 #(
		.INIT('h8)
	) name15275 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001 ,
		_w14699_,
		_w19322_
	);
	LUT2 #(
		.INIT('h8)
	) name15276 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][4]/P0001 ,
		_w14702_,
		_w19323_
	);
	LUT2 #(
		.INIT('h8)
	) name15277 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001 ,
		_w14711_,
		_w19324_
	);
	LUT2 #(
		.INIT('h8)
	) name15278 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001 ,
		_w14706_,
		_w19325_
	);
	LUT2 #(
		.INIT('h8)
	) name15279 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][4]/P0001 ,
		_w14713_,
		_w19326_
	);
	LUT2 #(
		.INIT('h8)
	) name15280 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001 ,
		_w14704_,
		_w19327_
	);
	LUT2 #(
		.INIT('h8)
	) name15281 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][4]/P0001 ,
		_w14708_,
		_w19328_
	);
	LUT2 #(
		.INIT('h1)
	) name15282 (
		_w19322_,
		_w19323_,
		_w19329_
	);
	LUT2 #(
		.INIT('h1)
	) name15283 (
		_w19324_,
		_w19325_,
		_w19330_
	);
	LUT2 #(
		.INIT('h1)
	) name15284 (
		_w19326_,
		_w19327_,
		_w19331_
	);
	LUT2 #(
		.INIT('h4)
	) name15285 (
		_w19328_,
		_w19331_,
		_w19332_
	);
	LUT2 #(
		.INIT('h8)
	) name15286 (
		_w19329_,
		_w19330_,
		_w19333_
	);
	LUT2 #(
		.INIT('h8)
	) name15287 (
		_w19332_,
		_w19333_,
		_w19334_
	);
	LUT2 #(
		.INIT('h2)
	) name15288 (
		_w14697_,
		_w19334_,
		_w19335_
	);
	LUT2 #(
		.INIT('h1)
	) name15289 (
		_w19320_,
		_w19321_,
		_w19336_
	);
	LUT2 #(
		.INIT('h4)
	) name15290 (
		_w19335_,
		_w19336_,
		_w19337_
	);
	LUT2 #(
		.INIT('h1)
	) name15291 (
		_w19298_,
		_w19337_,
		_w19338_
	);
	LUT2 #(
		.INIT('h4)
	) name15292 (
		_w19301_,
		_w19337_,
		_w19339_
	);
	LUT2 #(
		.INIT('h1)
	) name15293 (
		_w19315_,
		_w19338_,
		_w19340_
	);
	LUT2 #(
		.INIT('h4)
	) name15294 (
		_w19339_,
		_w19340_,
		_w19341_
	);
	LUT2 #(
		.INIT('h1)
	) name15295 (
		_w19319_,
		_w19341_,
		_w19342_
	);
	LUT2 #(
		.INIT('h2)
	) name15296 (
		_w6095_,
		_w19342_,
		_w19343_
	);
	LUT2 #(
		.INIT('h8)
	) name15297 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w19304_,
		_w19344_
	);
	LUT2 #(
		.INIT('h4)
	) name15298 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w19302_,
		_w19345_
	);
	LUT2 #(
		.INIT('h8)
	) name15299 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w19299_,
		_w19346_
	);
	LUT2 #(
		.INIT('h4)
	) name15300 (
		_w4137_,
		_w19268_,
		_w19347_
	);
	LUT2 #(
		.INIT('h8)
	) name15301 (
		_w4137_,
		_w19271_,
		_w19348_
	);
	LUT2 #(
		.INIT('h4)
	) name15302 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w19273_,
		_w19349_
	);
	LUT2 #(
		.INIT('h1)
	) name15303 (
		_w19344_,
		_w19345_,
		_w19350_
	);
	LUT2 #(
		.INIT('h1)
	) name15304 (
		_w19346_,
		_w19347_,
		_w19351_
	);
	LUT2 #(
		.INIT('h1)
	) name15305 (
		_w19348_,
		_w19349_,
		_w19352_
	);
	LUT2 #(
		.INIT('h8)
	) name15306 (
		_w19351_,
		_w19352_,
		_w19353_
	);
	LUT2 #(
		.INIT('h8)
	) name15307 (
		_w19350_,
		_w19353_,
		_w19354_
	);
	LUT2 #(
		.INIT('h2)
	) name15308 (
		_w19205_,
		_w19354_,
		_w19355_
	);
	LUT2 #(
		.INIT('h8)
	) name15309 (
		_w6097_,
		_w19301_,
		_w19356_
	);
	LUT2 #(
		.INIT('h1)
	) name15310 (
		_w4117_,
		_w19356_,
		_w19357_
	);
	LUT2 #(
		.INIT('h4)
	) name15311 (
		_w19355_,
		_w19357_,
		_w19358_
	);
	LUT2 #(
		.INIT('h4)
	) name15312 (
		_w19343_,
		_w19358_,
		_w19359_
	);
	LUT2 #(
		.INIT('h4)
	) name15313 (
		_w19311_,
		_w19359_,
		_w19360_
	);
	LUT2 #(
		.INIT('h4)
	) name15314 (
		\core_eu_ec_cun_condOK_CE_reg/P0001 ,
		_w4117_,
		_w19361_
	);
	LUT2 #(
		.INIT('h2)
	) name15315 (
		_w4149_,
		_w19361_,
		_w19362_
	);
	LUT2 #(
		.INIT('h4)
	) name15316 (
		_w19360_,
		_w19362_,
		_w19363_
	);
	LUT2 #(
		.INIT('h2)
	) name15317 (
		_w15314_,
		_w17777_,
		_w19364_
	);
	LUT2 #(
		.INIT('h1)
	) name15318 (
		_w17778_,
		_w19364_,
		_w19365_
	);
	LUT2 #(
		.INIT('h8)
	) name15319 (
		_w15244_,
		_w19365_,
		_w19366_
	);
	LUT2 #(
		.INIT('h1)
	) name15320 (
		_w15244_,
		_w19365_,
		_w19367_
	);
	LUT2 #(
		.INIT('h1)
	) name15321 (
		_w19366_,
		_w19367_,
		_w19368_
	);
	LUT2 #(
		.INIT('h2)
	) name15322 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19368_,
		_w19369_
	);
	LUT2 #(
		.INIT('h1)
	) name15323 (
		_w17767_,
		_w17774_,
		_w19370_
	);
	LUT2 #(
		.INIT('h1)
	) name15324 (
		_w17698_,
		_w17745_,
		_w19371_
	);
	LUT2 #(
		.INIT('h2)
	) name15325 (
		_w17772_,
		_w19371_,
		_w19372_
	);
	LUT2 #(
		.INIT('h1)
	) name15326 (
		_w17759_,
		_w19372_,
		_w19373_
	);
	LUT2 #(
		.INIT('h1)
	) name15327 (
		_w17768_,
		_w19373_,
		_w19374_
	);
	LUT2 #(
		.INIT('h2)
	) name15328 (
		_w19370_,
		_w19374_,
		_w19375_
	);
	LUT2 #(
		.INIT('h4)
	) name15329 (
		_w19370_,
		_w19374_,
		_w19376_
	);
	LUT2 #(
		.INIT('h1)
	) name15330 (
		_w19375_,
		_w19376_,
		_w19377_
	);
	LUT2 #(
		.INIT('h4)
	) name15331 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19377_,
		_w19378_
	);
	LUT2 #(
		.INIT('h1)
	) name15332 (
		_w19369_,
		_w19378_,
		_w19379_
	);
	LUT2 #(
		.INIT('h2)
	) name15333 (
		_w18262_,
		_w19379_,
		_w19380_
	);
	LUT2 #(
		.INIT('h2)
	) name15334 (
		_w14664_,
		_w17805_,
		_w19381_
	);
	LUT2 #(
		.INIT('h2)
	) name15335 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 ,
		_w19381_,
		_w19382_
	);
	LUT2 #(
		.INIT('h2)
	) name15336 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w17806_,
		_w19383_
	);
	LUT2 #(
		.INIT('h8)
	) name15337 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w18268_,
		_w19384_
	);
	LUT2 #(
		.INIT('h8)
	) name15338 (
		_w14665_,
		_w17822_,
		_w19385_
	);
	LUT2 #(
		.INIT('h1)
	) name15339 (
		_w19384_,
		_w19385_,
		_w19386_
	);
	LUT2 #(
		.INIT('h2)
	) name15340 (
		_w19383_,
		_w19386_,
		_w19387_
	);
	LUT2 #(
		.INIT('h1)
	) name15341 (
		_w19382_,
		_w19387_,
		_w19388_
	);
	LUT2 #(
		.INIT('h1)
	) name15342 (
		_w18262_,
		_w19388_,
		_w19389_
	);
	LUT2 #(
		.INIT('h2)
	) name15343 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[15]/P0001 ,
		_w19383_,
		_w19390_
	);
	LUT2 #(
		.INIT('h1)
	) name15344 (
		_w19389_,
		_w19390_,
		_w19391_
	);
	LUT2 #(
		.INIT('h4)
	) name15345 (
		_w19380_,
		_w19391_,
		_w19392_
	);
	LUT2 #(
		.INIT('h2)
	) name15346 (
		_w14752_,
		_w19379_,
		_w19393_
	);
	LUT2 #(
		.INIT('h2)
	) name15347 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 ,
		_w17809_,
		_w19394_
	);
	LUT2 #(
		.INIT('h1)
	) name15348 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w17806_,
		_w19395_
	);
	LUT2 #(
		.INIT('h1)
	) name15349 (
		_w17823_,
		_w17828_,
		_w19396_
	);
	LUT2 #(
		.INIT('h2)
	) name15350 (
		_w19395_,
		_w19396_,
		_w19397_
	);
	LUT2 #(
		.INIT('h1)
	) name15351 (
		_w19394_,
		_w19397_,
		_w19398_
	);
	LUT2 #(
		.INIT('h1)
	) name15352 (
		_w14752_,
		_w19398_,
		_w19399_
	);
	LUT2 #(
		.INIT('h2)
	) name15353 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[15]/P0001 ,
		_w19395_,
		_w19400_
	);
	LUT2 #(
		.INIT('h1)
	) name15354 (
		_w19399_,
		_w19400_,
		_w19401_
	);
	LUT2 #(
		.INIT('h4)
	) name15355 (
		_w19393_,
		_w19401_,
		_w19402_
	);
	LUT2 #(
		.INIT('h2)
	) name15356 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17794_,
		_w19403_
	);
	LUT2 #(
		.INIT('h1)
	) name15357 (
		_w15317_,
		_w17781_,
		_w19404_
	);
	LUT2 #(
		.INIT('h8)
	) name15358 (
		_w17779_,
		_w19404_,
		_w19405_
	);
	LUT2 #(
		.INIT('h1)
	) name15359 (
		_w17779_,
		_w19404_,
		_w19406_
	);
	LUT2 #(
		.INIT('h1)
	) name15360 (
		_w19405_,
		_w19406_,
		_w19407_
	);
	LUT2 #(
		.INIT('h4)
	) name15361 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19407_,
		_w19408_
	);
	LUT2 #(
		.INIT('h1)
	) name15362 (
		_w19403_,
		_w19408_,
		_w19409_
	);
	LUT2 #(
		.INIT('h1)
	) name15363 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		_w19410_
	);
	LUT2 #(
		.INIT('h8)
	) name15364 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		_w19411_
	);
	LUT2 #(
		.INIT('h1)
	) name15365 (
		_w19410_,
		_w19411_,
		_w19412_
	);
	LUT2 #(
		.INIT('h8)
	) name15366 (
		_w19197_,
		_w19412_,
		_w19413_
	);
	LUT2 #(
		.INIT('h2)
	) name15367 (
		_w17698_,
		_w17743_,
		_w19414_
	);
	LUT2 #(
		.INIT('h4)
	) name15368 (
		_w17698_,
		_w17743_,
		_w19415_
	);
	LUT2 #(
		.INIT('h1)
	) name15369 (
		_w19414_,
		_w19415_,
		_w19416_
	);
	LUT2 #(
		.INIT('h8)
	) name15370 (
		_w17737_,
		_w19416_,
		_w19417_
	);
	LUT2 #(
		.INIT('h1)
	) name15371 (
		_w17737_,
		_w19416_,
		_w19418_
	);
	LUT2 #(
		.INIT('h1)
	) name15372 (
		_w19417_,
		_w19418_,
		_w19419_
	);
	LUT2 #(
		.INIT('h2)
	) name15373 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19419_,
		_w19420_
	);
	LUT2 #(
		.INIT('h4)
	) name15374 (
		_w16363_,
		_w17662_,
		_w19421_
	);
	LUT2 #(
		.INIT('h2)
	) name15375 (
		_w17674_,
		_w19421_,
		_w19422_
	);
	LUT2 #(
		.INIT('h2)
	) name15376 (
		_w17567_,
		_w19422_,
		_w19423_
	);
	LUT2 #(
		.INIT('h2)
	) name15377 (
		_w17685_,
		_w19423_,
		_w19424_
	);
	LUT2 #(
		.INIT('h2)
	) name15378 (
		_w16980_,
		_w19424_,
		_w19425_
	);
	LUT2 #(
		.INIT('h2)
	) name15379 (
		_w17690_,
		_w19425_,
		_w19426_
	);
	LUT2 #(
		.INIT('h4)
	) name15380 (
		_w17692_,
		_w19426_,
		_w19427_
	);
	LUT2 #(
		.INIT('h1)
	) name15381 (
		_w17092_,
		_w19427_,
		_w19428_
	);
	LUT2 #(
		.INIT('h2)
	) name15382 (
		_w17079_,
		_w19428_,
		_w19429_
	);
	LUT2 #(
		.INIT('h4)
	) name15383 (
		_w17079_,
		_w19428_,
		_w19430_
	);
	LUT2 #(
		.INIT('h1)
	) name15384 (
		_w19429_,
		_w19430_,
		_w19431_
	);
	LUT2 #(
		.INIT('h8)
	) name15385 (
		_w17095_,
		_w19431_,
		_w19432_
	);
	LUT2 #(
		.INIT('h1)
	) name15386 (
		_w17095_,
		_w19431_,
		_w19433_
	);
	LUT2 #(
		.INIT('h1)
	) name15387 (
		_w19432_,
		_w19433_,
		_w19434_
	);
	LUT2 #(
		.INIT('h4)
	) name15388 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19434_,
		_w19435_
	);
	LUT2 #(
		.INIT('h1)
	) name15389 (
		_w19420_,
		_w19435_,
		_w19436_
	);
	LUT2 #(
		.INIT('h1)
	) name15390 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		_w19437_
	);
	LUT2 #(
		.INIT('h8)
	) name15391 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SCLKi_cnt_reg[1]/NET0131 ,
		_w19438_
	);
	LUT2 #(
		.INIT('h1)
	) name15392 (
		_w19437_,
		_w19438_,
		_w19439_
	);
	LUT2 #(
		.INIT('h8)
	) name15393 (
		_w19130_,
		_w19439_,
		_w19440_
	);
	LUT2 #(
		.INIT('h2)
	) name15394 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_ckr_reg_DO_reg[8]/NET0131 ,
		_w19441_
	);
	LUT2 #(
		.INIT('h4)
	) name15395 (
		\clkc_OUTcnt_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[14]/NET0131 ,
		_w19442_
	);
	LUT2 #(
		.INIT('h4)
	) name15396 (
		\clkc_OUTcnt_reg[2]/NET0131 ,
		\clkc_ckr_reg_DO_reg[10]/NET0131 ,
		_w19443_
	);
	LUT2 #(
		.INIT('h4)
	) name15397 (
		\clkc_OUTcnt_reg[3]/NET0131 ,
		\clkc_ckr_reg_DO_reg[11]/NET0131 ,
		_w19444_
	);
	LUT2 #(
		.INIT('h4)
	) name15398 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_ckr_reg_DO_reg[8]/NET0131 ,
		_w19445_
	);
	LUT2 #(
		.INIT('h2)
	) name15399 (
		\clkc_OUTcnt_reg[3]/NET0131 ,
		\clkc_ckr_reg_DO_reg[11]/NET0131 ,
		_w19446_
	);
	LUT2 #(
		.INIT('h2)
	) name15400 (
		\clkc_OUTcnt_reg[2]/NET0131 ,
		\clkc_ckr_reg_DO_reg[10]/NET0131 ,
		_w19447_
	);
	LUT2 #(
		.INIT('h4)
	) name15401 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		\clkc_ckr_reg_DO_reg[12]/NET0131 ,
		_w19448_
	);
	LUT2 #(
		.INIT('h2)
	) name15402 (
		\clkc_OUTcnt_reg[1]/NET0131 ,
		\clkc_ckr_reg_DO_reg[9]/NET0131 ,
		_w19449_
	);
	LUT2 #(
		.INIT('h2)
	) name15403 (
		\clkc_OUTcnt_reg[5]/NET0131 ,
		\clkc_ckr_reg_DO_reg[13]/NET0131 ,
		_w19450_
	);
	LUT2 #(
		.INIT('h4)
	) name15404 (
		\clkc_OUTcnt_reg[1]/NET0131 ,
		\clkc_ckr_reg_DO_reg[9]/NET0131 ,
		_w19451_
	);
	LUT2 #(
		.INIT('h4)
	) name15405 (
		\clkc_OUTcnt_reg[5]/NET0131 ,
		\clkc_ckr_reg_DO_reg[13]/NET0131 ,
		_w19452_
	);
	LUT2 #(
		.INIT('h2)
	) name15406 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		\clkc_ckr_reg_DO_reg[12]/NET0131 ,
		_w19453_
	);
	LUT2 #(
		.INIT('h2)
	) name15407 (
		\clkc_OUTcnt_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[14]/NET0131 ,
		_w19454_
	);
	LUT2 #(
		.INIT('h1)
	) name15408 (
		_w19442_,
		_w19443_,
		_w19455_
	);
	LUT2 #(
		.INIT('h1)
	) name15409 (
		_w19444_,
		_w19445_,
		_w19456_
	);
	LUT2 #(
		.INIT('h1)
	) name15410 (
		_w19446_,
		_w19447_,
		_w19457_
	);
	LUT2 #(
		.INIT('h1)
	) name15411 (
		_w19448_,
		_w19449_,
		_w19458_
	);
	LUT2 #(
		.INIT('h1)
	) name15412 (
		_w19450_,
		_w19451_,
		_w19459_
	);
	LUT2 #(
		.INIT('h1)
	) name15413 (
		_w19452_,
		_w19453_,
		_w19460_
	);
	LUT2 #(
		.INIT('h4)
	) name15414 (
		_w19454_,
		_w19460_,
		_w19461_
	);
	LUT2 #(
		.INIT('h8)
	) name15415 (
		_w19458_,
		_w19459_,
		_w19462_
	);
	LUT2 #(
		.INIT('h8)
	) name15416 (
		_w19456_,
		_w19457_,
		_w19463_
	);
	LUT2 #(
		.INIT('h8)
	) name15417 (
		_w19455_,
		_w19463_,
		_w19464_
	);
	LUT2 #(
		.INIT('h8)
	) name15418 (
		_w19461_,
		_w19462_,
		_w19465_
	);
	LUT2 #(
		.INIT('h8)
	) name15419 (
		_w19464_,
		_w19465_,
		_w19466_
	);
	LUT2 #(
		.INIT('h4)
	) name15420 (
		_w19441_,
		_w19466_,
		_w19467_
	);
	LUT2 #(
		.INIT('h8)
	) name15421 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_OUTcnt_reg[1]/NET0131 ,
		_w19468_
	);
	LUT2 #(
		.INIT('h8)
	) name15422 (
		\clkc_OUTcnt_reg[2]/NET0131 ,
		_w19468_,
		_w19469_
	);
	LUT2 #(
		.INIT('h8)
	) name15423 (
		\clkc_OUTcnt_reg[3]/NET0131 ,
		_w19469_,
		_w19470_
	);
	LUT2 #(
		.INIT('h8)
	) name15424 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		_w19470_,
		_w19471_
	);
	LUT2 #(
		.INIT('h8)
	) name15425 (
		\clkc_OUTcnt_reg[5]/NET0131 ,
		_w19471_,
		_w19472_
	);
	LUT2 #(
		.INIT('h1)
	) name15426 (
		\clkc_OUTcnt_reg[6]/NET0131 ,
		_w19472_,
		_w19473_
	);
	LUT2 #(
		.INIT('h8)
	) name15427 (
		\clkc_OUTcnt_reg[6]/NET0131 ,
		_w19472_,
		_w19474_
	);
	LUT2 #(
		.INIT('h1)
	) name15428 (
		_w19467_,
		_w19473_,
		_w19475_
	);
	LUT2 #(
		.INIT('h4)
	) name15429 (
		_w19474_,
		_w19475_,
		_w19476_
	);
	LUT2 #(
		.INIT('h2)
	) name15430 (
		\core_c_psq_INT_en_reg/NET0131 ,
		_w4094_,
		_w19477_
	);
	LUT2 #(
		.INIT('h2)
	) name15431 (
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		_w19477_,
		_w19478_
	);
	LUT2 #(
		.INIT('h8)
	) name15432 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		\core_c_psq_Iflag_reg[5]/NET0131 ,
		_w19479_
	);
	LUT2 #(
		.INIT('h4)
	) name15433 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w19479_,
		_w19480_
	);
	LUT2 #(
		.INIT('h8)
	) name15434 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		\core_c_psq_Iflag_reg[8]/NET0131 ,
		_w19481_
	);
	LUT2 #(
		.INIT('h1)
	) name15435 (
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		_w19481_,
		_w19482_
	);
	LUT2 #(
		.INIT('h1)
	) name15436 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w19482_,
		_w19483_
	);
	LUT2 #(
		.INIT('h2)
	) name15437 (
		_w19477_,
		_w19483_,
		_w19484_
	);
	LUT2 #(
		.INIT('h8)
	) name15438 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		\core_c_psq_Iflag_reg[9]/NET0131 ,
		_w19485_
	);
	LUT2 #(
		.INIT('h4)
	) name15439 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w19485_,
		_w19486_
	);
	LUT2 #(
		.INIT('h2)
	) name15440 (
		_w19484_,
		_w19486_,
		_w19487_
	);
	LUT2 #(
		.INIT('h8)
	) name15441 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		\core_c_psq_Iflag_reg[6]/NET0131 ,
		_w19488_
	);
	LUT2 #(
		.INIT('h4)
	) name15442 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w19488_,
		_w19489_
	);
	LUT2 #(
		.INIT('h8)
	) name15443 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		\core_c_psq_Iflag_reg[4]/NET0131 ,
		_w19490_
	);
	LUT2 #(
		.INIT('h4)
	) name15444 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w19490_,
		_w19491_
	);
	LUT2 #(
		.INIT('h8)
	) name15445 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		\core_c_psq_Iflag_reg[7]/NET0131 ,
		_w19492_
	);
	LUT2 #(
		.INIT('h4)
	) name15446 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w19492_,
		_w19493_
	);
	LUT2 #(
		.INIT('h1)
	) name15447 (
		_w19491_,
		_w19493_,
		_w19494_
	);
	LUT2 #(
		.INIT('h4)
	) name15448 (
		_w19489_,
		_w19494_,
		_w19495_
	);
	LUT2 #(
		.INIT('h8)
	) name15449 (
		_w19480_,
		_w19495_,
		_w19496_
	);
	LUT2 #(
		.INIT('h8)
	) name15450 (
		_w19487_,
		_w19496_,
		_w19497_
	);
	LUT2 #(
		.INIT('h1)
	) name15451 (
		_w19478_,
		_w19497_,
		_w19498_
	);
	LUT2 #(
		.INIT('h8)
	) name15452 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w14665_,
		_w19499_
	);
	LUT2 #(
		.INIT('h1)
	) name15453 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 ,
		_w19499_,
		_w19500_
	);
	LUT2 #(
		.INIT('h4)
	) name15454 (
		_w18268_,
		_w19383_,
		_w19501_
	);
	LUT2 #(
		.INIT('h1)
	) name15455 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w10289_,
		_w19502_
	);
	LUT2 #(
		.INIT('h2)
	) name15456 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w13075_,
		_w19503_
	);
	LUT2 #(
		.INIT('h1)
	) name15457 (
		_w19502_,
		_w19503_,
		_w19504_
	);
	LUT2 #(
		.INIT('h2)
	) name15458 (
		_w19499_,
		_w19504_,
		_w19505_
	);
	LUT2 #(
		.INIT('h4)
	) name15459 (
		_w19500_,
		_w19501_,
		_w19506_
	);
	LUT2 #(
		.INIT('h4)
	) name15460 (
		_w19505_,
		_w19506_,
		_w19507_
	);
	LUT2 #(
		.INIT('h8)
	) name15461 (
		_w18269_,
		_w19383_,
		_w19508_
	);
	LUT2 #(
		.INIT('h2)
	) name15462 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[9]/P0001 ,
		_w19383_,
		_w19509_
	);
	LUT2 #(
		.INIT('h1)
	) name15463 (
		_w19508_,
		_w19509_,
		_w19510_
	);
	LUT2 #(
		.INIT('h4)
	) name15464 (
		_w19507_,
		_w19510_,
		_w19511_
	);
	LUT2 #(
		.INIT('h1)
	) name15465 (
		_w18262_,
		_w19511_,
		_w19512_
	);
	LUT2 #(
		.INIT('h1)
	) name15466 (
		_w17092_,
		_w17692_,
		_w19513_
	);
	LUT2 #(
		.INIT('h8)
	) name15467 (
		_w19426_,
		_w19513_,
		_w19514_
	);
	LUT2 #(
		.INIT('h1)
	) name15468 (
		_w19426_,
		_w19513_,
		_w19515_
	);
	LUT2 #(
		.INIT('h1)
	) name15469 (
		_w19514_,
		_w19515_,
		_w19516_
	);
	LUT2 #(
		.INIT('h2)
	) name15470 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19516_,
		_w19517_
	);
	LUT2 #(
		.INIT('h1)
	) name15471 (
		_w16856_,
		_w17687_,
		_w19518_
	);
	LUT2 #(
		.INIT('h1)
	) name15472 (
		_w16979_,
		_w19424_,
		_w19519_
	);
	LUT2 #(
		.INIT('h1)
	) name15473 (
		_w17688_,
		_w19519_,
		_w19520_
	);
	LUT2 #(
		.INIT('h2)
	) name15474 (
		_w19518_,
		_w19520_,
		_w19521_
	);
	LUT2 #(
		.INIT('h4)
	) name15475 (
		_w19518_,
		_w19520_,
		_w19522_
	);
	LUT2 #(
		.INIT('h1)
	) name15476 (
		_w19521_,
		_w19522_,
		_w19523_
	);
	LUT2 #(
		.INIT('h4)
	) name15477 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19523_,
		_w19524_
	);
	LUT2 #(
		.INIT('h1)
	) name15478 (
		_w19517_,
		_w19524_,
		_w19525_
	);
	LUT2 #(
		.INIT('h2)
	) name15479 (
		_w18262_,
		_w19525_,
		_w19526_
	);
	LUT2 #(
		.INIT('h1)
	) name15480 (
		_w19512_,
		_w19526_,
		_w19527_
	);
	LUT2 #(
		.INIT('h4)
	) name15481 (
		\core_c_dec_SHTop_E_reg/P0001 ,
		_w4117_,
		_w19528_
	);
	LUT2 #(
		.INIT('h8)
	) name15482 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w6028_,
		_w19529_
	);
	LUT2 #(
		.INIT('h1)
	) name15483 (
		_w6119_,
		_w19529_,
		_w19530_
	);
	LUT2 #(
		.INIT('h4)
	) name15484 (
		_w4117_,
		_w19530_,
		_w19531_
	);
	LUT2 #(
		.INIT('h2)
	) name15485 (
		_w4116_,
		_w19528_,
		_w19532_
	);
	LUT2 #(
		.INIT('h4)
	) name15486 (
		_w19531_,
		_w19532_,
		_w19533_
	);
	LUT2 #(
		.INIT('h8)
	) name15487 (
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		_w19411_,
		_w19534_
	);
	LUT2 #(
		.INIT('h8)
	) name15488 (
		\sport0_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		_w19534_,
		_w19535_
	);
	LUT2 #(
		.INIT('h8)
	) name15489 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		_w19535_,
		_w19536_
	);
	LUT2 #(
		.INIT('h1)
	) name15490 (
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		_w19536_,
		_w19537_
	);
	LUT2 #(
		.INIT('h8)
	) name15491 (
		\sport0_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		_w19536_,
		_w19538_
	);
	LUT2 #(
		.INIT('h1)
	) name15492 (
		_w19537_,
		_w19538_,
		_w19539_
	);
	LUT2 #(
		.INIT('h8)
	) name15493 (
		_w19197_,
		_w19539_,
		_w19540_
	);
	LUT2 #(
		.INIT('h1)
	) name15494 (
		\sport0_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		_w19411_,
		_w19541_
	);
	LUT2 #(
		.INIT('h1)
	) name15495 (
		_w19534_,
		_w19541_,
		_w19542_
	);
	LUT2 #(
		.INIT('h8)
	) name15496 (
		_w19197_,
		_w19542_,
		_w19543_
	);
	LUT2 #(
		.INIT('h8)
	) name15497 (
		\sport0_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		_w19538_,
		_w19544_
	);
	LUT2 #(
		.INIT('h8)
	) name15498 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		_w19544_,
		_w19545_
	);
	LUT2 #(
		.INIT('h8)
	) name15499 (
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		_w19545_,
		_w19546_
	);
	LUT2 #(
		.INIT('h8)
	) name15500 (
		\sport0_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		_w19546_,
		_w19547_
	);
	LUT2 #(
		.INIT('h8)
	) name15501 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		_w19547_,
		_w19548_
	);
	LUT2 #(
		.INIT('h8)
	) name15502 (
		\sport0_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		_w19548_,
		_w19549_
	);
	LUT2 #(
		.INIT('h8)
	) name15503 (
		\sport0_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		_w19549_,
		_w19550_
	);
	LUT2 #(
		.INIT('h1)
	) name15504 (
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		_w19550_,
		_w19551_
	);
	LUT2 #(
		.INIT('h8)
	) name15505 (
		\sport0_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		_w19550_,
		_w19552_
	);
	LUT2 #(
		.INIT('h2)
	) name15506 (
		_w19197_,
		_w19551_,
		_w19553_
	);
	LUT2 #(
		.INIT('h4)
	) name15507 (
		_w19552_,
		_w19553_,
		_w19554_
	);
	LUT2 #(
		.INIT('h4)
	) name15508 (
		\sport0_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		_w19197_,
		_w19555_
	);
	LUT2 #(
		.INIT('h1)
	) name15509 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 ,
		_w19499_,
		_w19556_
	);
	LUT2 #(
		.INIT('h1)
	) name15510 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7607_,
		_w19557_
	);
	LUT2 #(
		.INIT('h2)
	) name15511 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12520_,
		_w19558_
	);
	LUT2 #(
		.INIT('h1)
	) name15512 (
		_w19557_,
		_w19558_,
		_w19559_
	);
	LUT2 #(
		.INIT('h2)
	) name15513 (
		_w19499_,
		_w19559_,
		_w19560_
	);
	LUT2 #(
		.INIT('h2)
	) name15514 (
		_w19501_,
		_w19556_,
		_w19561_
	);
	LUT2 #(
		.INIT('h4)
	) name15515 (
		_w19560_,
		_w19561_,
		_w19562_
	);
	LUT2 #(
		.INIT('h2)
	) name15516 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[0]/P0001 ,
		_w19383_,
		_w19563_
	);
	LUT2 #(
		.INIT('h1)
	) name15517 (
		_w19508_,
		_w19563_,
		_w19564_
	);
	LUT2 #(
		.INIT('h4)
	) name15518 (
		_w19562_,
		_w19564_,
		_w19565_
	);
	LUT2 #(
		.INIT('h1)
	) name15519 (
		_w18262_,
		_w19565_,
		_w19566_
	);
	LUT2 #(
		.INIT('h1)
	) name15520 (
		_w17660_,
		_w17668_,
		_w19567_
	);
	LUT2 #(
		.INIT('h8)
	) name15521 (
		_w16363_,
		_w19567_,
		_w19568_
	);
	LUT2 #(
		.INIT('h1)
	) name15522 (
		_w16363_,
		_w19567_,
		_w19569_
	);
	LUT2 #(
		.INIT('h1)
	) name15523 (
		_w19568_,
		_w19569_,
		_w19570_
	);
	LUT2 #(
		.INIT('h4)
	) name15524 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19570_,
		_w19571_
	);
	LUT2 #(
		.INIT('h1)
	) name15525 (
		_w17654_,
		_w17667_,
		_w19572_
	);
	LUT2 #(
		.INIT('h1)
	) name15526 (
		_w16363_,
		_w17660_,
		_w19573_
	);
	LUT2 #(
		.INIT('h1)
	) name15527 (
		_w17668_,
		_w19573_,
		_w19574_
	);
	LUT2 #(
		.INIT('h2)
	) name15528 (
		_w19572_,
		_w19574_,
		_w19575_
	);
	LUT2 #(
		.INIT('h4)
	) name15529 (
		_w19572_,
		_w19574_,
		_w19576_
	);
	LUT2 #(
		.INIT('h1)
	) name15530 (
		_w19575_,
		_w19576_,
		_w19577_
	);
	LUT2 #(
		.INIT('h2)
	) name15531 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19577_,
		_w19578_
	);
	LUT2 #(
		.INIT('h1)
	) name15532 (
		_w15775_,
		_w16353_,
		_w19579_
	);
	LUT2 #(
		.INIT('h2)
	) name15533 (
		_w16059_,
		_w16350_,
		_w19580_
	);
	LUT2 #(
		.INIT('h2)
	) name15534 (
		_w16358_,
		_w19580_,
		_w19581_
	);
	LUT2 #(
		.INIT('h4)
	) name15535 (
		_w19579_,
		_w19581_,
		_w19582_
	);
	LUT2 #(
		.INIT('h2)
	) name15536 (
		_w19579_,
		_w19581_,
		_w19583_
	);
	LUT2 #(
		.INIT('h1)
	) name15537 (
		_w19582_,
		_w19583_,
		_w19584_
	);
	LUT2 #(
		.INIT('h4)
	) name15538 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19584_,
		_w19585_
	);
	LUT2 #(
		.INIT('h1)
	) name15539 (
		_w15898_,
		_w16360_,
		_w19586_
	);
	LUT2 #(
		.INIT('h1)
	) name15540 (
		_w15775_,
		_w19581_,
		_w19587_
	);
	LUT2 #(
		.INIT('h1)
	) name15541 (
		_w16353_,
		_w19587_,
		_w19588_
	);
	LUT2 #(
		.INIT('h2)
	) name15542 (
		_w19586_,
		_w19588_,
		_w19589_
	);
	LUT2 #(
		.INIT('h4)
	) name15543 (
		_w19586_,
		_w19588_,
		_w19590_
	);
	LUT2 #(
		.INIT('h1)
	) name15544 (
		_w19589_,
		_w19590_,
		_w19591_
	);
	LUT2 #(
		.INIT('h8)
	) name15545 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19591_,
		_w19592_
	);
	LUT2 #(
		.INIT('h1)
	) name15546 (
		_w19585_,
		_w19592_,
		_w19593_
	);
	LUT2 #(
		.INIT('h2)
	) name15547 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19570_,
		_w19594_
	);
	LUT2 #(
		.INIT('h4)
	) name15548 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19591_,
		_w19595_
	);
	LUT2 #(
		.INIT('h1)
	) name15549 (
		_w19594_,
		_w19595_,
		_w19596_
	);
	LUT2 #(
		.INIT('h1)
	) name15550 (
		_w16058_,
		_w16356_,
		_w19597_
	);
	LUT2 #(
		.INIT('h2)
	) name15551 (
		_w16350_,
		_w19597_,
		_w19598_
	);
	LUT2 #(
		.INIT('h4)
	) name15552 (
		_w16350_,
		_w19597_,
		_w19599_
	);
	LUT2 #(
		.INIT('h1)
	) name15553 (
		_w19598_,
		_w19599_,
		_w19600_
	);
	LUT2 #(
		.INIT('h1)
	) name15554 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19600_,
		_w19601_
	);
	LUT2 #(
		.INIT('h1)
	) name15555 (
		_w15978_,
		_w16355_,
		_w19602_
	);
	LUT2 #(
		.INIT('h1)
	) name15556 (
		_w16058_,
		_w16350_,
		_w19603_
	);
	LUT2 #(
		.INIT('h1)
	) name15557 (
		_w16356_,
		_w19603_,
		_w19604_
	);
	LUT2 #(
		.INIT('h2)
	) name15558 (
		_w19602_,
		_w19604_,
		_w19605_
	);
	LUT2 #(
		.INIT('h4)
	) name15559 (
		_w19602_,
		_w19604_,
		_w19606_
	);
	LUT2 #(
		.INIT('h1)
	) name15560 (
		_w19605_,
		_w19606_,
		_w19607_
	);
	LUT2 #(
		.INIT('h2)
	) name15561 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19607_,
		_w19608_
	);
	LUT2 #(
		.INIT('h1)
	) name15562 (
		_w19601_,
		_w19608_,
		_w19609_
	);
	LUT2 #(
		.INIT('h2)
	) name15563 (
		_w16327_,
		_w16343_,
		_w19610_
	);
	LUT2 #(
		.INIT('h1)
	) name15564 (
		_w16347_,
		_w19610_,
		_w19611_
	);
	LUT2 #(
		.INIT('h1)
	) name15565 (
		_w16339_,
		_w16346_,
		_w19612_
	);
	LUT2 #(
		.INIT('h4)
	) name15566 (
		_w19611_,
		_w19612_,
		_w19613_
	);
	LUT2 #(
		.INIT('h2)
	) name15567 (
		_w19611_,
		_w19612_,
		_w19614_
	);
	LUT2 #(
		.INIT('h1)
	) name15568 (
		_w19613_,
		_w19614_,
		_w19615_
	);
	LUT2 #(
		.INIT('h4)
	) name15569 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19615_,
		_w19616_
	);
	LUT2 #(
		.INIT('h8)
	) name15570 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19600_,
		_w19617_
	);
	LUT2 #(
		.INIT('h1)
	) name15571 (
		_w19616_,
		_w19617_,
		_w19618_
	);
	LUT2 #(
		.INIT('h4)
	) name15572 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w18289_,
		_w19619_
	);
	LUT2 #(
		.INIT('h4)
	) name15573 (
		_w16159_,
		_w16310_,
		_w19620_
	);
	LUT2 #(
		.INIT('h1)
	) name15574 (
		_w16311_,
		_w19620_,
		_w19621_
	);
	LUT2 #(
		.INIT('h8)
	) name15575 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19621_,
		_w19622_
	);
	LUT2 #(
		.INIT('h1)
	) name15576 (
		_w19619_,
		_w19622_,
		_w19623_
	);
	LUT2 #(
		.INIT('h4)
	) name15577 (
		_w16276_,
		_w16304_,
		_w19624_
	);
	LUT2 #(
		.INIT('h1)
	) name15578 (
		_w16305_,
		_w19624_,
		_w19625_
	);
	LUT2 #(
		.INIT('h4)
	) name15579 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19625_,
		_w19626_
	);
	LUT2 #(
		.INIT('h8)
	) name15580 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w18284_,
		_w19627_
	);
	LUT2 #(
		.INIT('h1)
	) name15581 (
		_w19626_,
		_w19627_,
		_w19628_
	);
	LUT2 #(
		.INIT('h2)
	) name15582 (
		_w16312_,
		_w16326_,
		_w19629_
	);
	LUT2 #(
		.INIT('h1)
	) name15583 (
		_w16327_,
		_w19629_,
		_w19630_
	);
	LUT2 #(
		.INIT('h2)
	) name15584 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19630_,
		_w19631_
	);
	LUT2 #(
		.INIT('h1)
	) name15585 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19621_,
		_w19632_
	);
	LUT2 #(
		.INIT('h1)
	) name15586 (
		_w19631_,
		_w19632_,
		_w19633_
	);
	LUT2 #(
		.INIT('h4)
	) name15587 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19607_,
		_w19634_
	);
	LUT2 #(
		.INIT('h8)
	) name15588 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19584_,
		_w19635_
	);
	LUT2 #(
		.INIT('h1)
	) name15589 (
		_w19634_,
		_w19635_,
		_w19636_
	);
	LUT2 #(
		.INIT('h2)
	) name15590 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19615_,
		_w19637_
	);
	LUT2 #(
		.INIT('h1)
	) name15591 (
		_w16343_,
		_w16347_,
		_w19638_
	);
	LUT2 #(
		.INIT('h4)
	) name15592 (
		_w16327_,
		_w19638_,
		_w19639_
	);
	LUT2 #(
		.INIT('h2)
	) name15593 (
		_w16327_,
		_w19638_,
		_w19640_
	);
	LUT2 #(
		.INIT('h1)
	) name15594 (
		_w19639_,
		_w19640_,
		_w19641_
	);
	LUT2 #(
		.INIT('h4)
	) name15595 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19641_,
		_w19642_
	);
	LUT2 #(
		.INIT('h1)
	) name15596 (
		_w19637_,
		_w19642_,
		_w19643_
	);
	LUT2 #(
		.INIT('h2)
	) name15597 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19641_,
		_w19644_
	);
	LUT2 #(
		.INIT('h4)
	) name15598 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19630_,
		_w19645_
	);
	LUT2 #(
		.INIT('h1)
	) name15599 (
		_w19644_,
		_w19645_,
		_w19646_
	);
	LUT2 #(
		.INIT('h8)
	) name15600 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		_w19647_
	);
	LUT2 #(
		.INIT('h4)
	) name15601 (
		_w16286_,
		_w19647_,
		_w19648_
	);
	LUT2 #(
		.INIT('h2)
	) name15602 (
		_w16286_,
		_w19647_,
		_w19649_
	);
	LUT2 #(
		.INIT('h1)
	) name15603 (
		_w19648_,
		_w19649_,
		_w19650_
	);
	LUT2 #(
		.INIT('h2)
	) name15604 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19650_,
		_w19651_
	);
	LUT2 #(
		.INIT('h4)
	) name15605 (
		_w7469_,
		_w17341_,
		_w19652_
	);
	LUT2 #(
		.INIT('h1)
	) name15606 (
		_w19651_,
		_w19652_,
		_w19653_
	);
	LUT2 #(
		.INIT('h1)
	) name15607 (
		_w16301_,
		_w16303_,
		_w19654_
	);
	LUT2 #(
		.INIT('h4)
	) name15608 (
		_w16297_,
		_w19654_,
		_w19655_
	);
	LUT2 #(
		.INIT('h2)
	) name15609 (
		_w16297_,
		_w19654_,
		_w19656_
	);
	LUT2 #(
		.INIT('h1)
	) name15610 (
		_w19655_,
		_w19656_,
		_w19657_
	);
	LUT2 #(
		.INIT('h2)
	) name15611 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19657_,
		_w19658_
	);
	LUT2 #(
		.INIT('h1)
	) name15612 (
		_w16291_,
		_w16296_,
		_w19659_
	);
	LUT2 #(
		.INIT('h1)
	) name15613 (
		_w16297_,
		_w19659_,
		_w19660_
	);
	LUT2 #(
		.INIT('h4)
	) name15614 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19660_,
		_w19661_
	);
	LUT2 #(
		.INIT('h1)
	) name15615 (
		_w19658_,
		_w19661_,
		_w19662_
	);
	LUT2 #(
		.INIT('h4)
	) name15616 (
		_w16280_,
		_w16290_,
		_w19663_
	);
	LUT2 #(
		.INIT('h1)
	) name15617 (
		_w16291_,
		_w19663_,
		_w19664_
	);
	LUT2 #(
		.INIT('h2)
	) name15618 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19664_,
		_w19665_
	);
	LUT2 #(
		.INIT('h4)
	) name15619 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19650_,
		_w19666_
	);
	LUT2 #(
		.INIT('h1)
	) name15620 (
		_w19665_,
		_w19666_,
		_w19667_
	);
	LUT2 #(
		.INIT('h1)
	) name15621 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19657_,
		_w19668_
	);
	LUT2 #(
		.INIT('h8)
	) name15622 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19625_,
		_w19669_
	);
	LUT2 #(
		.INIT('h1)
	) name15623 (
		_w19668_,
		_w19669_,
		_w19670_
	);
	LUT2 #(
		.INIT('h4)
	) name15624 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19664_,
		_w19671_
	);
	LUT2 #(
		.INIT('h8)
	) name15625 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19660_,
		_w19672_
	);
	LUT2 #(
		.INIT('h1)
	) name15626 (
		_w19671_,
		_w19672_,
		_w19673_
	);
	LUT2 #(
		.INIT('h2)
	) name15627 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 ,
		\memc_usysr_DO_reg[10]/NET0131 ,
		_w19674_
	);
	LUT2 #(
		.INIT('h8)
	) name15628 (
		_w19653_,
		_w19674_,
		_w19675_
	);
	LUT2 #(
		.INIT('h4)
	) name15629 (
		_w19667_,
		_w19675_,
		_w19676_
	);
	LUT2 #(
		.INIT('h8)
	) name15630 (
		_w19673_,
		_w19676_,
		_w19677_
	);
	LUT2 #(
		.INIT('h8)
	) name15631 (
		_w19662_,
		_w19677_,
		_w19678_
	);
	LUT2 #(
		.INIT('h8)
	) name15632 (
		_w19670_,
		_w19678_,
		_w19679_
	);
	LUT2 #(
		.INIT('h8)
	) name15633 (
		_w19628_,
		_w19679_,
		_w19680_
	);
	LUT2 #(
		.INIT('h4)
	) name15634 (
		_w18291_,
		_w19680_,
		_w19681_
	);
	LUT2 #(
		.INIT('h8)
	) name15635 (
		_w19623_,
		_w19681_,
		_w19682_
	);
	LUT2 #(
		.INIT('h4)
	) name15636 (
		_w19633_,
		_w19682_,
		_w19683_
	);
	LUT2 #(
		.INIT('h8)
	) name15637 (
		_w19646_,
		_w19683_,
		_w19684_
	);
	LUT2 #(
		.INIT('h8)
	) name15638 (
		_w19618_,
		_w19684_,
		_w19685_
	);
	LUT2 #(
		.INIT('h4)
	) name15639 (
		_w19643_,
		_w19685_,
		_w19686_
	);
	LUT2 #(
		.INIT('h4)
	) name15640 (
		_w19609_,
		_w19686_,
		_w19687_
	);
	LUT2 #(
		.INIT('h8)
	) name15641 (
		_w19636_,
		_w19687_,
		_w19688_
	);
	LUT2 #(
		.INIT('h8)
	) name15642 (
		_w19593_,
		_w19688_,
		_w19689_
	);
	LUT2 #(
		.INIT('h8)
	) name15643 (
		_w19596_,
		_w19689_,
		_w19690_
	);
	LUT2 #(
		.INIT('h1)
	) name15644 (
		_w19571_,
		_w19578_,
		_w19691_
	);
	LUT2 #(
		.INIT('h4)
	) name15645 (
		_w19690_,
		_w19691_,
		_w19692_
	);
	LUT2 #(
		.INIT('h8)
	) name15646 (
		_w18262_,
		_w19692_,
		_w19693_
	);
	LUT2 #(
		.INIT('h1)
	) name15647 (
		_w19566_,
		_w19693_,
		_w19694_
	);
	LUT2 #(
		.INIT('h8)
	) name15648 (
		\core_c_dec_Post2_E_reg/P0001 ,
		_w4117_,
		_w19695_
	);
	LUT2 #(
		.INIT('h4)
	) name15649 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w19696_
	);
	LUT2 #(
		.INIT('h4)
	) name15650 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w19697_
	);
	LUT2 #(
		.INIT('h8)
	) name15651 (
		_w6027_,
		_w19697_,
		_w19698_
	);
	LUT2 #(
		.INIT('h8)
	) name15652 (
		_w19696_,
		_w19698_,
		_w19699_
	);
	LUT2 #(
		.INIT('h8)
	) name15653 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w19699_,
		_w19700_
	);
	LUT2 #(
		.INIT('h1)
	) name15654 (
		_w13574_,
		_w13577_,
		_w19701_
	);
	LUT2 #(
		.INIT('h4)
	) name15655 (
		_w6023_,
		_w19701_,
		_w19702_
	);
	LUT2 #(
		.INIT('h2)
	) name15656 (
		_w6121_,
		_w19700_,
		_w19703_
	);
	LUT2 #(
		.INIT('h8)
	) name15657 (
		_w19702_,
		_w19703_,
		_w19704_
	);
	LUT2 #(
		.INIT('h1)
	) name15658 (
		_w4117_,
		_w19704_,
		_w19705_
	);
	LUT2 #(
		.INIT('h1)
	) name15659 (
		_w19695_,
		_w19705_,
		_w19706_
	);
	LUT2 #(
		.INIT('h2)
	) name15660 (
		_w4116_,
		_w19706_,
		_w19707_
	);
	LUT2 #(
		.INIT('h2)
	) name15661 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w17820_,
		_w19708_
	);
	LUT2 #(
		.INIT('h8)
	) name15662 (
		_w18119_,
		_w18166_,
		_w19709_
	);
	LUT2 #(
		.INIT('h4)
	) name15663 (
		_w17931_,
		_w18001_,
		_w19710_
	);
	LUT2 #(
		.INIT('h1)
	) name15664 (
		_w18148_,
		_w19710_,
		_w19711_
	);
	LUT2 #(
		.INIT('h2)
	) name15665 (
		_w17945_,
		_w19711_,
		_w19712_
	);
	LUT2 #(
		.INIT('h8)
	) name15666 (
		_w18790_,
		_w18797_,
		_w19713_
	);
	LUT2 #(
		.INIT('h2)
	) name15667 (
		_w18050_,
		_w19712_,
		_w19714_
	);
	LUT2 #(
		.INIT('h8)
	) name15668 (
		_w19713_,
		_w19714_,
		_w19715_
	);
	LUT2 #(
		.INIT('h8)
	) name15669 (
		_w18076_,
		_w18145_,
		_w19716_
	);
	LUT2 #(
		.INIT('h2)
	) name15670 (
		_w17931_,
		_w18108_,
		_w19717_
	);
	LUT2 #(
		.INIT('h4)
	) name15671 (
		_w17933_,
		_w19717_,
		_w19718_
	);
	LUT2 #(
		.INIT('h4)
	) name15672 (
		_w18159_,
		_w18184_,
		_w19719_
	);
	LUT2 #(
		.INIT('h4)
	) name15673 (
		_w17929_,
		_w18088_,
		_w19720_
	);
	LUT2 #(
		.INIT('h8)
	) name15674 (
		_w17929_,
		_w18765_,
		_w19721_
	);
	LUT2 #(
		.INIT('h1)
	) name15675 (
		_w19720_,
		_w19721_,
		_w19722_
	);
	LUT2 #(
		.INIT('h1)
	) name15676 (
		_w17922_,
		_w19722_,
		_w19723_
	);
	LUT2 #(
		.INIT('h4)
	) name15677 (
		_w18121_,
		_w18163_,
		_w19724_
	);
	LUT2 #(
		.INIT('h1)
	) name15678 (
		_w18147_,
		_w18153_,
		_w19725_
	);
	LUT2 #(
		.INIT('h4)
	) name15679 (
		_w18176_,
		_w19725_,
		_w19726_
	);
	LUT2 #(
		.INIT('h8)
	) name15680 (
		_w18084_,
		_w19726_,
		_w19727_
	);
	LUT2 #(
		.INIT('h2)
	) name15681 (
		_w17945_,
		_w19727_,
		_w19728_
	);
	LUT2 #(
		.INIT('h2)
	) name15682 (
		_w17965_,
		_w18091_,
		_w19729_
	);
	LUT2 #(
		.INIT('h8)
	) name15683 (
		_w18059_,
		_w18195_,
		_w19730_
	);
	LUT2 #(
		.INIT('h8)
	) name15684 (
		_w18142_,
		_w19730_,
		_w19731_
	);
	LUT2 #(
		.INIT('h1)
	) name15685 (
		_w18117_,
		_w18133_,
		_w19732_
	);
	LUT2 #(
		.INIT('h8)
	) name15686 (
		_w17920_,
		_w18066_,
		_w19733_
	);
	LUT2 #(
		.INIT('h4)
	) name15687 (
		_w17914_,
		_w17975_,
		_w19734_
	);
	LUT2 #(
		.INIT('h1)
	) name15688 (
		_w19733_,
		_w19734_,
		_w19735_
	);
	LUT2 #(
		.INIT('h2)
	) name15689 (
		_w18100_,
		_w19735_,
		_w19736_
	);
	LUT2 #(
		.INIT('h1)
	) name15690 (
		_w18096_,
		_w18129_,
		_w19737_
	);
	LUT2 #(
		.INIT('h2)
	) name15691 (
		_w18171_,
		_w18180_,
		_w19738_
	);
	LUT2 #(
		.INIT('h8)
	) name15692 (
		_w17925_,
		_w18107_,
		_w19739_
	);
	LUT2 #(
		.INIT('h1)
	) name15693 (
		_w19738_,
		_w19739_,
		_w19740_
	);
	LUT2 #(
		.INIT('h1)
	) name15694 (
		_w17931_,
		_w19740_,
		_w19741_
	);
	LUT2 #(
		.INIT('h8)
	) name15695 (
		_w17930_,
		_w18106_,
		_w19742_
	);
	LUT2 #(
		.INIT('h2)
	) name15696 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w12000_,
		_w19743_
	);
	LUT2 #(
		.INIT('h8)
	) name15697 (
		_w18120_,
		_w18745_,
		_w19744_
	);
	LUT2 #(
		.INIT('h1)
	) name15698 (
		_w18102_,
		_w19735_,
		_w19745_
	);
	LUT2 #(
		.INIT('h4)
	) name15699 (
		_w18159_,
		_w18187_,
		_w19746_
	);
	LUT2 #(
		.INIT('h4)
	) name15700 (
		_w18180_,
		_w18758_,
		_w19747_
	);
	LUT2 #(
		.INIT('h1)
	) name15701 (
		_w19744_,
		_w19745_,
		_w19748_
	);
	LUT2 #(
		.INIT('h1)
	) name15702 (
		_w19746_,
		_w19747_,
		_w19749_
	);
	LUT2 #(
		.INIT('h8)
	) name15703 (
		_w19748_,
		_w19749_,
		_w19750_
	);
	LUT2 #(
		.INIT('h2)
	) name15704 (
		_w17931_,
		_w19750_,
		_w19751_
	);
	LUT2 #(
		.INIT('h1)
	) name15705 (
		_w19742_,
		_w19743_,
		_w19752_
	);
	LUT2 #(
		.INIT('h4)
	) name15706 (
		_w18065_,
		_w19752_,
		_w19753_
	);
	LUT2 #(
		.INIT('h4)
	) name15707 (
		_w19709_,
		_w19753_,
		_w19754_
	);
	LUT2 #(
		.INIT('h1)
	) name15708 (
		_w19719_,
		_w19723_,
		_w19755_
	);
	LUT2 #(
		.INIT('h1)
	) name15709 (
		_w19724_,
		_w19729_,
		_w19756_
	);
	LUT2 #(
		.INIT('h1)
	) name15710 (
		_w19732_,
		_w19736_,
		_w19757_
	);
	LUT2 #(
		.INIT('h4)
	) name15711 (
		_w19737_,
		_w19757_,
		_w19758_
	);
	LUT2 #(
		.INIT('h8)
	) name15712 (
		_w19755_,
		_w19756_,
		_w19759_
	);
	LUT2 #(
		.INIT('h4)
	) name15713 (
		_w19718_,
		_w19754_,
		_w19760_
	);
	LUT2 #(
		.INIT('h8)
	) name15714 (
		_w19759_,
		_w19760_,
		_w19761_
	);
	LUT2 #(
		.INIT('h4)
	) name15715 (
		_w19741_,
		_w19758_,
		_w19762_
	);
	LUT2 #(
		.INIT('h8)
	) name15716 (
		_w19761_,
		_w19762_,
		_w19763_
	);
	LUT2 #(
		.INIT('h4)
	) name15717 (
		_w19728_,
		_w19731_,
		_w19764_
	);
	LUT2 #(
		.INIT('h4)
	) name15718 (
		_w19751_,
		_w19764_,
		_w19765_
	);
	LUT2 #(
		.INIT('h8)
	) name15719 (
		_w19716_,
		_w19763_,
		_w19766_
	);
	LUT2 #(
		.INIT('h8)
	) name15720 (
		_w19765_,
		_w19766_,
		_w19767_
	);
	LUT2 #(
		.INIT('h8)
	) name15721 (
		_w18007_,
		_w19715_,
		_w19768_
	);
	LUT2 #(
		.INIT('h8)
	) name15722 (
		_w19767_,
		_w19768_,
		_w19769_
	);
	LUT2 #(
		.INIT('h4)
	) name15723 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w19769_,
		_w19770_
	);
	LUT2 #(
		.INIT('h1)
	) name15724 (
		_w19708_,
		_w19770_,
		_w19771_
	);
	LUT2 #(
		.INIT('h2)
	) name15725 (
		_w18717_,
		_w19771_,
		_w19772_
	);
	LUT2 #(
		.INIT('h1)
	) name15726 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[15]/P0001 ,
		_w18717_,
		_w19773_
	);
	LUT2 #(
		.INIT('h1)
	) name15727 (
		_w19772_,
		_w19773_,
		_w19774_
	);
	LUT2 #(
		.INIT('h8)
	) name15728 (
		_w14752_,
		_w19525_,
		_w19775_
	);
	LUT2 #(
		.INIT('h8)
	) name15729 (
		_w17802_,
		_w18325_,
		_w19776_
	);
	LUT2 #(
		.INIT('h8)
	) name15730 (
		_w19504_,
		_w19776_,
		_w19777_
	);
	LUT2 #(
		.INIT('h2)
	) name15731 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[9]/P0001 ,
		_w17809_,
		_w19778_
	);
	LUT2 #(
		.INIT('h8)
	) name15732 (
		_w18332_,
		_w19395_,
		_w19779_
	);
	LUT2 #(
		.INIT('h1)
	) name15733 (
		_w14752_,
		_w19779_,
		_w19780_
	);
	LUT2 #(
		.INIT('h4)
	) name15734 (
		_w19778_,
		_w19780_,
		_w19781_
	);
	LUT2 #(
		.INIT('h4)
	) name15735 (
		_w19777_,
		_w19781_,
		_w19782_
	);
	LUT2 #(
		.INIT('h1)
	) name15736 (
		_w19775_,
		_w19782_,
		_w19783_
	);
	LUT2 #(
		.INIT('h2)
	) name15737 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w17836_,
		_w19784_
	);
	LUT2 #(
		.INIT('h2)
	) name15738 (
		_w17931_,
		_w18918_,
		_w19785_
	);
	LUT2 #(
		.INIT('h4)
	) name15739 (
		_w17933_,
		_w19785_,
		_w19786_
	);
	LUT2 #(
		.INIT('h8)
	) name15740 (
		_w17976_,
		_w18077_,
		_w19787_
	);
	LUT2 #(
		.INIT('h1)
	) name15741 (
		_w18037_,
		_w19787_,
		_w19788_
	);
	LUT2 #(
		.INIT('h1)
	) name15742 (
		_w18032_,
		_w18085_,
		_w19789_
	);
	LUT2 #(
		.INIT('h8)
	) name15743 (
		_w19788_,
		_w19789_,
		_w19790_
	);
	LUT2 #(
		.INIT('h8)
	) name15744 (
		_w18902_,
		_w19790_,
		_w19791_
	);
	LUT2 #(
		.INIT('h8)
	) name15745 (
		_w18054_,
		_w19713_,
		_w19792_
	);
	LUT2 #(
		.INIT('h8)
	) name15746 (
		_w18738_,
		_w19792_,
		_w19793_
	);
	LUT2 #(
		.INIT('h8)
	) name15747 (
		_w19791_,
		_w19793_,
		_w19794_
	);
	LUT2 #(
		.INIT('h8)
	) name15748 (
		_w18070_,
		_w18124_,
		_w19795_
	);
	LUT2 #(
		.INIT('h1)
	) name15749 (
		_w18117_,
		_w18912_,
		_w19796_
	);
	LUT2 #(
		.INIT('h4)
	) name15750 (
		_w18914_,
		_w19720_,
		_w19797_
	);
	LUT2 #(
		.INIT('h8)
	) name15751 (
		_w17980_,
		_w18187_,
		_w19798_
	);
	LUT2 #(
		.INIT('h2)
	) name15752 (
		_w18056_,
		_w18189_,
		_w19799_
	);
	LUT2 #(
		.INIT('h4)
	) name15753 (
		_w18129_,
		_w18153_,
		_w19800_
	);
	LUT2 #(
		.INIT('h4)
	) name15754 (
		_w17929_,
		_w17952_,
		_w19801_
	);
	LUT2 #(
		.INIT('h1)
	) name15755 (
		_w19710_,
		_w19801_,
		_w19802_
	);
	LUT2 #(
		.INIT('h2)
	) name15756 (
		_w18171_,
		_w19802_,
		_w19803_
	);
	LUT2 #(
		.INIT('h1)
	) name15757 (
		_w18043_,
		_w18761_,
		_w19804_
	);
	LUT2 #(
		.INIT('h2)
	) name15758 (
		_w18099_,
		_w19804_,
		_w19805_
	);
	LUT2 #(
		.INIT('h8)
	) name15759 (
		_w18046_,
		_w18740_,
		_w19806_
	);
	LUT2 #(
		.INIT('h2)
	) name15760 (
		_w17930_,
		_w18918_,
		_w19807_
	);
	LUT2 #(
		.INIT('h2)
	) name15761 (
		_w17931_,
		_w18914_,
		_w19808_
	);
	LUT2 #(
		.INIT('h4)
	) name15762 (
		_w18175_,
		_w19808_,
		_w19809_
	);
	LUT2 #(
		.INIT('h8)
	) name15763 (
		_w18183_,
		_w18893_,
		_w19810_
	);
	LUT2 #(
		.INIT('h8)
	) name15764 (
		_w17945_,
		_w17959_,
		_w19811_
	);
	LUT2 #(
		.INIT('h1)
	) name15765 (
		_w17972_,
		_w19811_,
		_w19812_
	);
	LUT2 #(
		.INIT('h8)
	) name15766 (
		_w18147_,
		_w18751_,
		_w19813_
	);
	LUT2 #(
		.INIT('h8)
	) name15767 (
		_w17986_,
		_w18103_,
		_w19814_
	);
	LUT2 #(
		.INIT('h2)
	) name15768 (
		_w18745_,
		_w18775_,
		_w19815_
	);
	LUT2 #(
		.INIT('h2)
	) name15769 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7164_,
		_w19816_
	);
	LUT2 #(
		.INIT('h4)
	) name15770 (
		_w17931_,
		_w18055_,
		_w19817_
	);
	LUT2 #(
		.INIT('h1)
	) name15771 (
		_w18139_,
		_w19817_,
		_w19818_
	);
	LUT2 #(
		.INIT('h2)
	) name15772 (
		_w18162_,
		_w19818_,
		_w19819_
	);
	LUT2 #(
		.INIT('h2)
	) name15773 (
		_w18136_,
		_w18907_,
		_w19820_
	);
	LUT2 #(
		.INIT('h1)
	) name15774 (
		_w19799_,
		_w19816_,
		_w19821_
	);
	LUT2 #(
		.INIT('h1)
	) name15775 (
		_w19800_,
		_w19814_,
		_w19822_
	);
	LUT2 #(
		.INIT('h8)
	) name15776 (
		_w19821_,
		_w19822_,
		_w19823_
	);
	LUT2 #(
		.INIT('h4)
	) name15777 (
		_w19795_,
		_w19823_,
		_w19824_
	);
	LUT2 #(
		.INIT('h1)
	) name15778 (
		_w19796_,
		_w19797_,
		_w19825_
	);
	LUT2 #(
		.INIT('h1)
	) name15779 (
		_w19798_,
		_w19806_,
		_w19826_
	);
	LUT2 #(
		.INIT('h1)
	) name15780 (
		_w19807_,
		_w19810_,
		_w19827_
	);
	LUT2 #(
		.INIT('h2)
	) name15781 (
		_w19812_,
		_w19813_,
		_w19828_
	);
	LUT2 #(
		.INIT('h4)
	) name15782 (
		_w19820_,
		_w19828_,
		_w19829_
	);
	LUT2 #(
		.INIT('h8)
	) name15783 (
		_w19826_,
		_w19827_,
		_w19830_
	);
	LUT2 #(
		.INIT('h8)
	) name15784 (
		_w19824_,
		_w19825_,
		_w19831_
	);
	LUT2 #(
		.INIT('h1)
	) name15785 (
		_w19786_,
		_w19803_,
		_w19832_
	);
	LUT2 #(
		.INIT('h1)
	) name15786 (
		_w19805_,
		_w19809_,
		_w19833_
	);
	LUT2 #(
		.INIT('h1)
	) name15787 (
		_w19815_,
		_w19819_,
		_w19834_
	);
	LUT2 #(
		.INIT('h8)
	) name15788 (
		_w19833_,
		_w19834_,
		_w19835_
	);
	LUT2 #(
		.INIT('h8)
	) name15789 (
		_w19831_,
		_w19832_,
		_w19836_
	);
	LUT2 #(
		.INIT('h8)
	) name15790 (
		_w19829_,
		_w19830_,
		_w19837_
	);
	LUT2 #(
		.INIT('h8)
	) name15791 (
		_w19836_,
		_w19837_,
		_w19838_
	);
	LUT2 #(
		.INIT('h8)
	) name15792 (
		_w19835_,
		_w19838_,
		_w19839_
	);
	LUT2 #(
		.INIT('h8)
	) name15793 (
		_w19794_,
		_w19839_,
		_w19840_
	);
	LUT2 #(
		.INIT('h4)
	) name15794 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w19840_,
		_w19841_
	);
	LUT2 #(
		.INIT('h1)
	) name15795 (
		_w19784_,
		_w19841_,
		_w19842_
	);
	LUT2 #(
		.INIT('h2)
	) name15796 (
		_w18886_,
		_w19842_,
		_w19843_
	);
	LUT2 #(
		.INIT('h1)
	) name15797 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[13]/P0001 ,
		_w18886_,
		_w19844_
	);
	LUT2 #(
		.INIT('h1)
	) name15798 (
		_w19843_,
		_w19844_,
		_w19845_
	);
	LUT2 #(
		.INIT('h1)
	) name15799 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w7859_,
		_w19846_
	);
	LUT2 #(
		.INIT('h2)
	) name15800 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12556_,
		_w19847_
	);
	LUT2 #(
		.INIT('h1)
	) name15801 (
		_w19846_,
		_w19847_,
		_w19848_
	);
	LUT2 #(
		.INIT('h2)
	) name15802 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w19848_,
		_w19849_
	);
	LUT2 #(
		.INIT('h4)
	) name15803 (
		_w17938_,
		_w18080_,
		_w19850_
	);
	LUT2 #(
		.INIT('h2)
	) name15804 (
		_w17925_,
		_w17998_,
		_w19851_
	);
	LUT2 #(
		.INIT('h1)
	) name15805 (
		_w17959_,
		_w18030_,
		_w19852_
	);
	LUT2 #(
		.INIT('h2)
	) name15806 (
		_w17945_,
		_w19852_,
		_w19853_
	);
	LUT2 #(
		.INIT('h1)
	) name15807 (
		_w18143_,
		_w19853_,
		_w19854_
	);
	LUT2 #(
		.INIT('h8)
	) name15808 (
		_w18891_,
		_w19854_,
		_w19855_
	);
	LUT2 #(
		.INIT('h4)
	) name15809 (
		_w17931_,
		_w18153_,
		_w19856_
	);
	LUT2 #(
		.INIT('h1)
	) name15810 (
		_w18070_,
		_w19856_,
		_w19857_
	);
	LUT2 #(
		.INIT('h2)
	) name15811 (
		_w18751_,
		_w19857_,
		_w19858_
	);
	LUT2 #(
		.INIT('h2)
	) name15812 (
		_w18754_,
		_w18912_,
		_w19859_
	);
	LUT2 #(
		.INIT('h2)
	) name15813 (
		_w18124_,
		_w18781_,
		_w19860_
	);
	LUT2 #(
		.INIT('h8)
	) name15814 (
		_w18745_,
		_w18893_,
		_w19861_
	);
	LUT2 #(
		.INIT('h4)
	) name15815 (
		_w17929_,
		_w18115_,
		_w19862_
	);
	LUT2 #(
		.INIT('h2)
	) name15816 (
		_w17931_,
		_w18170_,
		_w19863_
	);
	LUT2 #(
		.INIT('h1)
	) name15817 (
		_w19862_,
		_w19863_,
		_w19864_
	);
	LUT2 #(
		.INIT('h1)
	) name15818 (
		_w18918_,
		_w19864_,
		_w19865_
	);
	LUT2 #(
		.INIT('h8)
	) name15819 (
		_w18056_,
		_w18746_,
		_w19866_
	);
	LUT2 #(
		.INIT('h2)
	) name15820 (
		_w18055_,
		_w18743_,
		_w19867_
	);
	LUT2 #(
		.INIT('h1)
	) name15821 (
		_w18907_,
		_w18919_,
		_w19868_
	);
	LUT2 #(
		.INIT('h2)
	) name15822 (
		_w18759_,
		_w18912_,
		_w19869_
	);
	LUT2 #(
		.INIT('h1)
	) name15823 (
		_w18749_,
		_w18905_,
		_w19870_
	);
	LUT2 #(
		.INIT('h1)
	) name15824 (
		_w18914_,
		_w19870_,
		_w19871_
	);
	LUT2 #(
		.INIT('h8)
	) name15825 (
		_w18071_,
		_w18099_,
		_w19872_
	);
	LUT2 #(
		.INIT('h1)
	) name15826 (
		_w17972_,
		_w18783_,
		_w19873_
	);
	LUT2 #(
		.INIT('h8)
	) name15827 (
		_w19788_,
		_w19873_,
		_w19874_
	);
	LUT2 #(
		.INIT('h2)
	) name15828 (
		_w18765_,
		_w18898_,
		_w19875_
	);
	LUT2 #(
		.INIT('h2)
	) name15829 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7801_,
		_w19876_
	);
	LUT2 #(
		.INIT('h8)
	) name15830 (
		_w18139_,
		_w18740_,
		_w19877_
	);
	LUT2 #(
		.INIT('h1)
	) name15831 (
		_w19866_,
		_w19876_,
		_w19878_
	);
	LUT2 #(
		.INIT('h4)
	) name15832 (
		_w19867_,
		_w19878_,
		_w19879_
	);
	LUT2 #(
		.INIT('h4)
	) name15833 (
		_w19859_,
		_w19879_,
		_w19880_
	);
	LUT2 #(
		.INIT('h1)
	) name15834 (
		_w19861_,
		_w19865_,
		_w19881_
	);
	LUT2 #(
		.INIT('h1)
	) name15835 (
		_w19868_,
		_w19869_,
		_w19882_
	);
	LUT2 #(
		.INIT('h1)
	) name15836 (
		_w19871_,
		_w19872_,
		_w19883_
	);
	LUT2 #(
		.INIT('h4)
	) name15837 (
		_w19877_,
		_w19883_,
		_w19884_
	);
	LUT2 #(
		.INIT('h8)
	) name15838 (
		_w19881_,
		_w19882_,
		_w19885_
	);
	LUT2 #(
		.INIT('h4)
	) name15839 (
		_w19850_,
		_w19880_,
		_w19886_
	);
	LUT2 #(
		.INIT('h1)
	) name15840 (
		_w19851_,
		_w19858_,
		_w19887_
	);
	LUT2 #(
		.INIT('h4)
	) name15841 (
		_w19860_,
		_w19874_,
		_w19888_
	);
	LUT2 #(
		.INIT('h4)
	) name15842 (
		_w19875_,
		_w19888_,
		_w19889_
	);
	LUT2 #(
		.INIT('h8)
	) name15843 (
		_w19886_,
		_w19887_,
		_w19890_
	);
	LUT2 #(
		.INIT('h8)
	) name15844 (
		_w19884_,
		_w19885_,
		_w19891_
	);
	LUT2 #(
		.INIT('h8)
	) name15845 (
		_w19890_,
		_w19891_,
		_w19892_
	);
	LUT2 #(
		.INIT('h8)
	) name15846 (
		_w19855_,
		_w19889_,
		_w19893_
	);
	LUT2 #(
		.INIT('h8)
	) name15847 (
		_w19892_,
		_w19893_,
		_w19894_
	);
	LUT2 #(
		.INIT('h8)
	) name15848 (
		_w19792_,
		_w19894_,
		_w19895_
	);
	LUT2 #(
		.INIT('h4)
	) name15849 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w19895_,
		_w19896_
	);
	LUT2 #(
		.INIT('h1)
	) name15850 (
		_w19849_,
		_w19896_,
		_w19897_
	);
	LUT2 #(
		.INIT('h2)
	) name15851 (
		_w18886_,
		_w19897_,
		_w19898_
	);
	LUT2 #(
		.INIT('h1)
	) name15852 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[10]/P0001 ,
		_w18886_,
		_w19899_
	);
	LUT2 #(
		.INIT('h1)
	) name15853 (
		_w19898_,
		_w19899_,
		_w19900_
	);
	LUT2 #(
		.INIT('h2)
	) name15854 (
		_w19034_,
		_w19842_,
		_w19901_
	);
	LUT2 #(
		.INIT('h1)
	) name15855 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[13]/P0001 ,
		_w19034_,
		_w19902_
	);
	LUT2 #(
		.INIT('h1)
	) name15856 (
		_w19901_,
		_w19902_,
		_w19903_
	);
	LUT2 #(
		.INIT('h8)
	) name15857 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w4117_,
		_w19904_
	);
	LUT2 #(
		.INIT('h1)
	) name15858 (
		_w18848_,
		_w19904_,
		_w19905_
	);
	LUT2 #(
		.INIT('h2)
	) name15859 (
		_w4116_,
		_w19905_,
		_w19906_
	);
	LUT2 #(
		.INIT('h2)
	) name15860 (
		_w19034_,
		_w19897_,
		_w19907_
	);
	LUT2 #(
		.INIT('h1)
	) name15861 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[10]/P0001 ,
		_w19034_,
		_w19908_
	);
	LUT2 #(
		.INIT('h1)
	) name15862 (
		_w19907_,
		_w19908_,
		_w19909_
	);
	LUT2 #(
		.INIT('h8)
	) name15863 (
		_w5730_,
		_w13751_,
		_w19910_
	);
	LUT2 #(
		.INIT('h8)
	) name15864 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		_w19910_,
		_w19911_
	);
	LUT2 #(
		.INIT('h2)
	) name15865 (
		\bdma_CMcnt_reg[1]/NET0131 ,
		_w19911_,
		_w19912_
	);
	LUT2 #(
		.INIT('h8)
	) name15866 (
		_w13146_,
		_w13751_,
		_w19913_
	);
	LUT2 #(
		.INIT('h1)
	) name15867 (
		_w19912_,
		_w19913_,
		_w19914_
	);
	LUT2 #(
		.INIT('h1)
	) name15868 (
		_w13752_,
		_w19914_,
		_w19915_
	);
	LUT2 #(
		.INIT('h1)
	) name15869 (
		\bdma_CMcnt_reg[0]/NET0131 ,
		_w19910_,
		_w19916_
	);
	LUT2 #(
		.INIT('h1)
	) name15870 (
		_w13752_,
		_w19911_,
		_w19917_
	);
	LUT2 #(
		.INIT('h4)
	) name15871 (
		_w19916_,
		_w19917_,
		_w19918_
	);
	LUT2 #(
		.INIT('h1)
	) name15872 (
		_w6921_,
		_w13151_,
		_w19919_
	);
	LUT2 #(
		.INIT('h1)
	) name15873 (
		\bdma_BMcyc_del_reg/P0001 ,
		_w19919_,
		_w19920_
	);
	LUT2 #(
		.INIT('h4)
	) name15874 (
		_w6917_,
		_w13747_,
		_w19921_
	);
	LUT2 #(
		.INIT('h4)
	) name15875 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w5533_,
		_w19922_
	);
	LUT2 #(
		.INIT('h8)
	) name15876 (
		_w5554_,
		_w19922_,
		_w19923_
	);
	LUT2 #(
		.INIT('h4)
	) name15877 (
		_w19921_,
		_w19923_,
		_w19924_
	);
	LUT2 #(
		.INIT('h1)
	) name15878 (
		\bdma_BSreq_reg/NET0131 ,
		_w19920_,
		_w19925_
	);
	LUT2 #(
		.INIT('h4)
	) name15879 (
		_w19924_,
		_w19925_,
		_w19926_
	);
	LUT2 #(
		.INIT('h2)
	) name15880 (
		_w17833_,
		_w19771_,
		_w19927_
	);
	LUT2 #(
		.INIT('h1)
	) name15881 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[15]/P0001 ,
		_w17833_,
		_w19928_
	);
	LUT2 #(
		.INIT('h1)
	) name15882 (
		_w19927_,
		_w19928_,
		_w19929_
	);
	LUT2 #(
		.INIT('h8)
	) name15883 (
		\sport0_txctl_TCS_reg[0]/NET0131 ,
		\sport0_txctl_TCS_reg[2]/NET0131 ,
		_w19930_
	);
	LUT2 #(
		.INIT('h4)
	) name15884 (
		\sport0_cfg_TFSg_d1_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w19931_
	);
	LUT2 #(
		.INIT('h4)
	) name15885 (
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w19931_,
		_w19932_
	);
	LUT2 #(
		.INIT('h1)
	) name15886 (
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w19933_
	);
	LUT2 #(
		.INIT('h4)
	) name15887 (
		\ITFS0_pad ,
		\T_TFS0_pad ,
		_w19934_
	);
	LUT2 #(
		.INIT('h2)
	) name15888 (
		\ITFS0_pad ,
		_w13725_,
		_w19935_
	);
	LUT2 #(
		.INIT('h1)
	) name15889 (
		_w19934_,
		_w19935_,
		_w19936_
	);
	LUT2 #(
		.INIT('h2)
	) name15890 (
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w19936_,
		_w19937_
	);
	LUT2 #(
		.INIT('h4)
	) name15891 (
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w19936_,
		_w19938_
	);
	LUT2 #(
		.INIT('h1)
	) name15892 (
		_w19937_,
		_w19938_,
		_w19939_
	);
	LUT2 #(
		.INIT('h2)
	) name15893 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_cfg_TFSgi_d_reg/NET0131 ,
		_w19940_
	);
	LUT2 #(
		.INIT('h8)
	) name15894 (
		_w19939_,
		_w19940_,
		_w19941_
	);
	LUT2 #(
		.INIT('h2)
	) name15895 (
		_w19933_,
		_w19941_,
		_w19942_
	);
	LUT2 #(
		.INIT('h2)
	) name15896 (
		\sport0_cfg_TFSg_d2_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w19943_
	);
	LUT2 #(
		.INIT('h8)
	) name15897 (
		\sport0_cfg_TFSg_d3_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w19944_
	);
	LUT2 #(
		.INIT('h2)
	) name15898 (
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w19943_,
		_w19945_
	);
	LUT2 #(
		.INIT('h4)
	) name15899 (
		_w19944_,
		_w19945_,
		_w19946_
	);
	LUT2 #(
		.INIT('h2)
	) name15900 (
		\sport0_txctl_TCS_reg[0]/NET0131 ,
		_w19932_,
		_w19947_
	);
	LUT2 #(
		.INIT('h4)
	) name15901 (
		_w19946_,
		_w19947_,
		_w19948_
	);
	LUT2 #(
		.INIT('h4)
	) name15902 (
		_w19942_,
		_w19948_,
		_w19949_
	);
	LUT2 #(
		.INIT('h1)
	) name15903 (
		\sport0_txctl_TCS_reg[2]/NET0131 ,
		_w19949_,
		_w19950_
	);
	LUT2 #(
		.INIT('h1)
	) name15904 (
		\sport0_txctl_TCS_reg[1]/NET0131 ,
		_w19930_,
		_w19951_
	);
	LUT2 #(
		.INIT('h4)
	) name15905 (
		_w19950_,
		_w19951_,
		_w19952_
	);
	LUT2 #(
		.INIT('h4)
	) name15906 (
		\sport0_txctl_TCS_reg[0]/NET0131 ,
		\sport0_txctl_TCS_reg[1]/NET0131 ,
		_w19953_
	);
	LUT2 #(
		.INIT('h4)
	) name15907 (
		\sport0_txctl_TCS_reg[2]/NET0131 ,
		_w19953_,
		_w19954_
	);
	LUT2 #(
		.INIT('h1)
	) name15908 (
		\sport0_txctl_Bcnt_reg[0]/NET0131 ,
		\sport0_txctl_Bcnt_reg[1]/NET0131 ,
		_w19955_
	);
	LUT2 #(
		.INIT('h4)
	) name15909 (
		\sport0_txctl_Bcnt_reg[2]/NET0131 ,
		_w19955_,
		_w19956_
	);
	LUT2 #(
		.INIT('h4)
	) name15910 (
		\sport0_txctl_Bcnt_reg[3]/NET0131 ,
		_w19956_,
		_w19957_
	);
	LUT2 #(
		.INIT('h4)
	) name15911 (
		\sport0_txctl_Bcnt_reg[4]/NET0131 ,
		_w19957_,
		_w19958_
	);
	LUT2 #(
		.INIT('h2)
	) name15912 (
		_w19954_,
		_w19958_,
		_w19959_
	);
	LUT2 #(
		.INIT('h1)
	) name15913 (
		_w19952_,
		_w19959_,
		_w19960_
	);
	LUT2 #(
		.INIT('h2)
	) name15914 (
		\sport0_txctl_TXSHT_reg[14]/P0001 ,
		_w19960_,
		_w19961_
	);
	LUT2 #(
		.INIT('h8)
	) name15915 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w19960_,
		_w19962_
	);
	LUT2 #(
		.INIT('h1)
	) name15916 (
		_w19961_,
		_w19962_,
		_w19963_
	);
	LUT2 #(
		.INIT('h2)
	) name15917 (
		_w14752_,
		_w19692_,
		_w19964_
	);
	LUT2 #(
		.INIT('h8)
	) name15918 (
		_w19559_,
		_w19776_,
		_w19965_
	);
	LUT2 #(
		.INIT('h2)
	) name15919 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[0]/P0001 ,
		_w17809_,
		_w19966_
	);
	LUT2 #(
		.INIT('h2)
	) name15920 (
		_w19780_,
		_w19966_,
		_w19967_
	);
	LUT2 #(
		.INIT('h4)
	) name15921 (
		_w19965_,
		_w19967_,
		_w19968_
	);
	LUT2 #(
		.INIT('h1)
	) name15922 (
		_w19964_,
		_w19968_,
		_w19969_
	);
	LUT2 #(
		.INIT('h1)
	) name15923 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w11265_,
		_w19970_
	);
	LUT2 #(
		.INIT('h2)
	) name15924 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w13006_,
		_w19971_
	);
	LUT2 #(
		.INIT('h1)
	) name15925 (
		_w19970_,
		_w19971_,
		_w19972_
	);
	LUT2 #(
		.INIT('h2)
	) name15926 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w19972_,
		_w19973_
	);
	LUT2 #(
		.INIT('h8)
	) name15927 (
		_w18125_,
		_w18132_,
		_w19974_
	);
	LUT2 #(
		.INIT('h4)
	) name15928 (
		_w18060_,
		_w18797_,
		_w19975_
	);
	LUT2 #(
		.INIT('h4)
	) name15929 (
		_w17964_,
		_w18195_,
		_w19976_
	);
	LUT2 #(
		.INIT('h8)
	) name15930 (
		_w19975_,
		_w19976_,
		_w19977_
	);
	LUT2 #(
		.INIT('h4)
	) name15931 (
		_w17931_,
		_w17986_,
		_w19978_
	);
	LUT2 #(
		.INIT('h1)
	) name15932 (
		_w18043_,
		_w19978_,
		_w19979_
	);
	LUT2 #(
		.INIT('h2)
	) name15933 (
		_w18111_,
		_w19979_,
		_w19980_
	);
	LUT2 #(
		.INIT('h2)
	) name15934 (
		_w18765_,
		_w18775_,
		_w19981_
	);
	LUT2 #(
		.INIT('h2)
	) name15935 (
		_w18128_,
		_w18133_,
		_w19982_
	);
	LUT2 #(
		.INIT('h8)
	) name15936 (
		_w18103_,
		_w18178_,
		_w19983_
	);
	LUT2 #(
		.INIT('h4)
	) name15937 (
		_w17981_,
		_w18720_,
		_w19984_
	);
	LUT2 #(
		.INIT('h2)
	) name15938 (
		_w18748_,
		_w19984_,
		_w19985_
	);
	LUT2 #(
		.INIT('h8)
	) name15939 (
		_w18103_,
		_w18179_,
		_w19986_
	);
	LUT2 #(
		.INIT('h8)
	) name15940 (
		_w18107_,
		_w18163_,
		_w19987_
	);
	LUT2 #(
		.INIT('h1)
	) name15941 (
		_w18069_,
		_w18725_,
		_w19988_
	);
	LUT2 #(
		.INIT('h2)
	) name15942 (
		_w18115_,
		_w18149_,
		_w19989_
	);
	LUT2 #(
		.INIT('h2)
	) name15943 (
		_w17925_,
		_w19857_,
		_w19990_
	);
	LUT2 #(
		.INIT('h2)
	) name15944 (
		_w17945_,
		_w18781_,
		_w19991_
	);
	LUT2 #(
		.INIT('h2)
	) name15945 (
		_w18088_,
		_w19818_,
		_w19992_
	);
	LUT2 #(
		.INIT('h1)
	) name15946 (
		_w18091_,
		_w18991_,
		_w19993_
	);
	LUT2 #(
		.INIT('h2)
	) name15947 (
		_w18100_,
		_w18180_,
		_w19994_
	);
	LUT2 #(
		.INIT('h8)
	) name15948 (
		_w18125_,
		_w18131_,
		_w19995_
	);
	LUT2 #(
		.INIT('h1)
	) name15949 (
		_w18002_,
		_w18737_,
		_w19996_
	);
	LUT2 #(
		.INIT('h8)
	) name15950 (
		_w17978_,
		_w19996_,
		_w19997_
	);
	LUT2 #(
		.INIT('h4)
	) name15951 (
		_w18108_,
		_w18166_,
		_w19998_
	);
	LUT2 #(
		.INIT('h2)
	) name15952 (
		_w18724_,
		_w18735_,
		_w19999_
	);
	LUT2 #(
		.INIT('h2)
	) name15953 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11239_,
		_w20000_
	);
	LUT2 #(
		.INIT('h8)
	) name15954 (
		_w18106_,
		_w18163_,
		_w20001_
	);
	LUT2 #(
		.INIT('h1)
	) name15955 (
		_w17922_,
		_w18189_,
		_w20002_
	);
	LUT2 #(
		.INIT('h1)
	) name15956 (
		_w19974_,
		_w20000_,
		_w20003_
	);
	LUT2 #(
		.INIT('h1)
	) name15957 (
		_w19983_,
		_w20001_,
		_w20004_
	);
	LUT2 #(
		.INIT('h8)
	) name15958 (
		_w20003_,
		_w20004_,
		_w20005_
	);
	LUT2 #(
		.INIT('h1)
	) name15959 (
		_w18040_,
		_w18783_,
		_w20006_
	);
	LUT2 #(
		.INIT('h1)
	) name15960 (
		_w19986_,
		_w19987_,
		_w20007_
	);
	LUT2 #(
		.INIT('h4)
	) name15961 (
		_w19995_,
		_w20007_,
		_w20008_
	);
	LUT2 #(
		.INIT('h8)
	) name15962 (
		_w20005_,
		_w20006_,
		_w20009_
	);
	LUT2 #(
		.INIT('h2)
	) name15963 (
		_w18054_,
		_w19982_,
		_w20010_
	);
	LUT2 #(
		.INIT('h1)
	) name15964 (
		_w19993_,
		_w19994_,
		_w20011_
	);
	LUT2 #(
		.INIT('h1)
	) name15965 (
		_w19998_,
		_w20002_,
		_w20012_
	);
	LUT2 #(
		.INIT('h8)
	) name15966 (
		_w20011_,
		_w20012_,
		_w20013_
	);
	LUT2 #(
		.INIT('h8)
	) name15967 (
		_w20009_,
		_w20010_,
		_w20014_
	);
	LUT2 #(
		.INIT('h8)
	) name15968 (
		_w18727_,
		_w20008_,
		_w20015_
	);
	LUT2 #(
		.INIT('h1)
	) name15969 (
		_w19980_,
		_w19981_,
		_w20016_
	);
	LUT2 #(
		.INIT('h2)
	) name15970 (
		_w19988_,
		_w19989_,
		_w20017_
	);
	LUT2 #(
		.INIT('h1)
	) name15971 (
		_w19990_,
		_w19991_,
		_w20018_
	);
	LUT2 #(
		.INIT('h4)
	) name15972 (
		_w19992_,
		_w20018_,
		_w20019_
	);
	LUT2 #(
		.INIT('h8)
	) name15973 (
		_w20016_,
		_w20017_,
		_w20020_
	);
	LUT2 #(
		.INIT('h8)
	) name15974 (
		_w20014_,
		_w20015_,
		_w20021_
	);
	LUT2 #(
		.INIT('h4)
	) name15975 (
		_w18085_,
		_w20013_,
		_w20022_
	);
	LUT2 #(
		.INIT('h4)
	) name15976 (
		_w19985_,
		_w20022_,
		_w20023_
	);
	LUT2 #(
		.INIT('h8)
	) name15977 (
		_w20020_,
		_w20021_,
		_w20024_
	);
	LUT2 #(
		.INIT('h8)
	) name15978 (
		_w19997_,
		_w20019_,
		_w20025_
	);
	LUT2 #(
		.INIT('h8)
	) name15979 (
		_w19999_,
		_w20025_,
		_w20026_
	);
	LUT2 #(
		.INIT('h8)
	) name15980 (
		_w20023_,
		_w20024_,
		_w20027_
	);
	LUT2 #(
		.INIT('h8)
	) name15981 (
		_w18791_,
		_w20027_,
		_w20028_
	);
	LUT2 #(
		.INIT('h8)
	) name15982 (
		_w19977_,
		_w20026_,
		_w20029_
	);
	LUT2 #(
		.INIT('h8)
	) name15983 (
		_w20028_,
		_w20029_,
		_w20030_
	);
	LUT2 #(
		.INIT('h4)
	) name15984 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w20030_,
		_w20031_
	);
	LUT2 #(
		.INIT('h1)
	) name15985 (
		_w19973_,
		_w20031_,
		_w20032_
	);
	LUT2 #(
		.INIT('h2)
	) name15986 (
		_w18717_,
		_w20032_,
		_w20033_
	);
	LUT2 #(
		.INIT('h1)
	) name15987 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[7]/P0001 ,
		_w18717_,
		_w20034_
	);
	LUT2 #(
		.INIT('h1)
	) name15988 (
		_w20033_,
		_w20034_,
		_w20035_
	);
	LUT2 #(
		.INIT('h4)
	) name15989 (
		\bdma_BSreq_reg/NET0131 ,
		_w5534_,
		_w20036_
	);
	LUT2 #(
		.INIT('h8)
	) name15990 (
		\bdma_BWcnt_reg[0]/NET0131 ,
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w20037_
	);
	LUT2 #(
		.INIT('h8)
	) name15991 (
		_w20036_,
		_w20037_,
		_w20038_
	);
	LUT2 #(
		.INIT('h8)
	) name15992 (
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w20038_,
		_w20039_
	);
	LUT2 #(
		.INIT('h8)
	) name15993 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w20039_,
		_w20040_
	);
	LUT2 #(
		.INIT('h1)
	) name15994 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w20040_,
		_w20041_
	);
	LUT2 #(
		.INIT('h8)
	) name15995 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w20040_,
		_w20042_
	);
	LUT2 #(
		.INIT('h1)
	) name15996 (
		_w20041_,
		_w20042_,
		_w20043_
	);
	LUT2 #(
		.INIT('h4)
	) name15997 (
		_w13750_,
		_w20043_,
		_w20044_
	);
	LUT2 #(
		.INIT('h1)
	) name15998 (
		_w13806_,
		_w14424_,
		_w20045_
	);
	LUT2 #(
		.INIT('h1)
	) name15999 (
		_w13809_,
		_w14321_,
		_w20046_
	);
	LUT2 #(
		.INIT('h2)
	) name16000 (
		_w14362_,
		_w14406_,
		_w20047_
	);
	LUT2 #(
		.INIT('h4)
	) name16001 (
		_w14362_,
		_w14404_,
		_w20048_
	);
	LUT2 #(
		.INIT('h1)
	) name16002 (
		_w14358_,
		_w20047_,
		_w20049_
	);
	LUT2 #(
		.INIT('h4)
	) name16003 (
		_w20048_,
		_w20049_,
		_w20050_
	);
	LUT2 #(
		.INIT('h2)
	) name16004 (
		_w20046_,
		_w20050_,
		_w20051_
	);
	LUT2 #(
		.INIT('h4)
	) name16005 (
		_w20046_,
		_w20050_,
		_w20052_
	);
	LUT2 #(
		.INIT('h1)
	) name16006 (
		_w20051_,
		_w20052_,
		_w20053_
	);
	LUT2 #(
		.INIT('h2)
	) name16007 (
		_w13806_,
		_w20053_,
		_w20054_
	);
	LUT2 #(
		.INIT('h1)
	) name16008 (
		_w20045_,
		_w20054_,
		_w20055_
	);
	LUT2 #(
		.INIT('h2)
	) name16009 (
		_w14667_,
		_w20055_,
		_w20056_
	);
	LUT2 #(
		.INIT('h2)
	) name16010 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[11]/P0001 ,
		_w14667_,
		_w20057_
	);
	LUT2 #(
		.INIT('h1)
	) name16011 (
		_w20056_,
		_w20057_,
		_w20058_
	);
	LUT2 #(
		.INIT('h2)
	) name16012 (
		_w13805_,
		_w20055_,
		_w20059_
	);
	LUT2 #(
		.INIT('h2)
	) name16013 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[11]/P0001 ,
		_w13805_,
		_w20060_
	);
	LUT2 #(
		.INIT('h1)
	) name16014 (
		_w20059_,
		_w20060_,
		_w20061_
	);
	LUT2 #(
		.INIT('h4)
	) name16015 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_RDCMD_d1_reg/P0001 ,
		_w20062_
	);
	LUT2 #(
		.INIT('h4)
	) name16016 (
		\idma_RDCMD_reg/P0001 ,
		_w20062_,
		_w20063_
	);
	LUT2 #(
		.INIT('h4)
	) name16017 (
		\idma_PCrd_1st_reg/NET0131 ,
		_w20063_,
		_w20064_
	);
	LUT2 #(
		.INIT('h2)
	) name16018 (
		\idma_IAL_reg/P0001 ,
		\idma_ISn_reg/P0001 ,
		_w20065_
	);
	LUT2 #(
		.INIT('h8)
	) name16019 (
		\idma_IADi_reg[15]/P0001 ,
		_w20065_,
		_w20066_
	);
	LUT2 #(
		.INIT('h8)
	) name16020 (
		_w7530_,
		_w18226_,
		_w20067_
	);
	LUT2 #(
		.INIT('h1)
	) name16021 (
		_w20066_,
		_w20067_,
		_w20068_
	);
	LUT2 #(
		.INIT('h4)
	) name16022 (
		\idma_IADi_reg[15]/P0001 ,
		_w20065_,
		_w20069_
	);
	LUT2 #(
		.INIT('h1)
	) name16023 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w20070_
	);
	LUT2 #(
		.INIT('h8)
	) name16024 (
		_w7261_,
		_w20070_,
		_w20071_
	);
	LUT2 #(
		.INIT('h8)
	) name16025 (
		_w13762_,
		_w20071_,
		_w20072_
	);
	LUT2 #(
		.INIT('h1)
	) name16026 (
		_w20069_,
		_w20072_,
		_w20073_
	);
	LUT2 #(
		.INIT('h8)
	) name16027 (
		_w20068_,
		_w20073_,
		_w20074_
	);
	LUT2 #(
		.INIT('h2)
	) name16028 (
		\idma_PCrd_1st_reg/NET0131 ,
		_w20063_,
		_w20075_
	);
	LUT2 #(
		.INIT('h1)
	) name16029 (
		_w20064_,
		_w20075_,
		_w20076_
	);
	LUT2 #(
		.INIT('h8)
	) name16030 (
		_w20074_,
		_w20076_,
		_w20077_
	);
	LUT2 #(
		.INIT('h1)
	) name16031 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w10069_,
		_w20078_
	);
	LUT2 #(
		.INIT('h2)
	) name16032 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12904_,
		_w20079_
	);
	LUT2 #(
		.INIT('h1)
	) name16033 (
		_w20078_,
		_w20079_,
		_w20080_
	);
	LUT2 #(
		.INIT('h2)
	) name16034 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w20080_,
		_w20081_
	);
	LUT2 #(
		.INIT('h2)
	) name16035 (
		_w18115_,
		_w19857_,
		_w20082_
	);
	LUT2 #(
		.INIT('h2)
	) name16036 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9947_,
		_w20083_
	);
	LUT2 #(
		.INIT('h1)
	) name16037 (
		_w18141_,
		_w18783_,
		_w20084_
	);
	LUT2 #(
		.INIT('h1)
	) name16038 (
		_w17977_,
		_w18900_,
		_w20085_
	);
	LUT2 #(
		.INIT('h8)
	) name16039 (
		_w20084_,
		_w20085_,
		_w20086_
	);
	LUT2 #(
		.INIT('h8)
	) name16040 (
		_w19988_,
		_w20086_,
		_w20087_
	);
	LUT2 #(
		.INIT('h2)
	) name16041 (
		_w18107_,
		_w18743_,
		_w20088_
	);
	LUT2 #(
		.INIT('h8)
	) name16042 (
		_w18153_,
		_w19863_,
		_w20089_
	);
	LUT2 #(
		.INIT('h8)
	) name16043 (
		_w18145_,
		_w19789_,
		_w20090_
	);
	LUT2 #(
		.INIT('h8)
	) name16044 (
		_w17951_,
		_w17976_,
		_w20091_
	);
	LUT2 #(
		.INIT('h8)
	) name16045 (
		_w17925_,
		_w17980_,
		_w20092_
	);
	LUT2 #(
		.INIT('h2)
	) name16046 (
		_w18147_,
		_w18182_,
		_w20093_
	);
	LUT2 #(
		.INIT('h8)
	) name16047 (
		_w18758_,
		_w18761_,
		_w20094_
	);
	LUT2 #(
		.INIT('h8)
	) name16048 (
		_w18131_,
		_w18752_,
		_w20095_
	);
	LUT2 #(
		.INIT('h1)
	) name16049 (
		_w18746_,
		_w18763_,
		_w20096_
	);
	LUT2 #(
		.INIT('h1)
	) name16050 (
		_w17922_,
		_w20096_,
		_w20097_
	);
	LUT2 #(
		.INIT('h8)
	) name16051 (
		_w18046_,
		_w18171_,
		_w20098_
	);
	LUT2 #(
		.INIT('h2)
	) name16052 (
		_w18106_,
		_w18743_,
		_w20099_
	);
	LUT2 #(
		.INIT('h8)
	) name16053 (
		_w18043_,
		_w18758_,
		_w20100_
	);
	LUT2 #(
		.INIT('h2)
	) name16054 (
		_w18111_,
		_w18775_,
		_w20101_
	);
	LUT2 #(
		.INIT('h8)
	) name16055 (
		_w18132_,
		_w18752_,
		_w20102_
	);
	LUT2 #(
		.INIT('h1)
	) name16056 (
		_w18091_,
		_w18919_,
		_w20103_
	);
	LUT2 #(
		.INIT('h2)
	) name16057 (
		_w17931_,
		_w18907_,
		_w20104_
	);
	LUT2 #(
		.INIT('h4)
	) name16058 (
		_w17938_,
		_w20104_,
		_w20105_
	);
	LUT2 #(
		.INIT('h8)
	) name16059 (
		_w18054_,
		_w18790_,
		_w20106_
	);
	LUT2 #(
		.INIT('h8)
	) name16060 (
		_w18738_,
		_w20106_,
		_w20107_
	);
	LUT2 #(
		.INIT('h2)
	) name16061 (
		_w18038_,
		_w19787_,
		_w20108_
	);
	LUT2 #(
		.INIT('h2)
	) name16062 (
		_w18748_,
		_w19818_,
		_w20109_
	);
	LUT2 #(
		.INIT('h4)
	) name16063 (
		_w17924_,
		_w18780_,
		_w20110_
	);
	LUT2 #(
		.INIT('h8)
	) name16064 (
		_w17986_,
		_w18754_,
		_w20111_
	);
	LUT2 #(
		.INIT('h2)
	) name16065 (
		_w17945_,
		_w17962_,
		_w20112_
	);
	LUT2 #(
		.INIT('h2)
	) name16066 (
		_w18765_,
		_w18895_,
		_w20113_
	);
	LUT2 #(
		.INIT('h1)
	) name16067 (
		_w18192_,
		_w20083_,
		_w20114_
	);
	LUT2 #(
		.INIT('h1)
	) name16068 (
		_w20089_,
		_w20099_,
		_w20115_
	);
	LUT2 #(
		.INIT('h1)
	) name16069 (
		_w20102_,
		_w20111_,
		_w20116_
	);
	LUT2 #(
		.INIT('h8)
	) name16070 (
		_w20115_,
		_w20116_,
		_w20117_
	);
	LUT2 #(
		.INIT('h4)
	) name16071 (
		_w17972_,
		_w20114_,
		_w20118_
	);
	LUT2 #(
		.INIT('h1)
	) name16072 (
		_w18040_,
		_w20088_,
		_w20119_
	);
	LUT2 #(
		.INIT('h1)
	) name16073 (
		_w20091_,
		_w20094_,
		_w20120_
	);
	LUT2 #(
		.INIT('h1)
	) name16074 (
		_w20095_,
		_w20110_,
		_w20121_
	);
	LUT2 #(
		.INIT('h8)
	) name16075 (
		_w20120_,
		_w20121_,
		_w20122_
	);
	LUT2 #(
		.INIT('h8)
	) name16076 (
		_w20118_,
		_w20119_,
		_w20123_
	);
	LUT2 #(
		.INIT('h4)
	) name16077 (
		_w20092_,
		_w20117_,
		_w20124_
	);
	LUT2 #(
		.INIT('h1)
	) name16078 (
		_w20093_,
		_w20097_,
		_w20125_
	);
	LUT2 #(
		.INIT('h1)
	) name16079 (
		_w20098_,
		_w20100_,
		_w20126_
	);
	LUT2 #(
		.INIT('h4)
	) name16080 (
		_w20103_,
		_w20126_,
		_w20127_
	);
	LUT2 #(
		.INIT('h8)
	) name16081 (
		_w20124_,
		_w20125_,
		_w20128_
	);
	LUT2 #(
		.INIT('h8)
	) name16082 (
		_w20122_,
		_w20123_,
		_w20129_
	);
	LUT2 #(
		.INIT('h1)
	) name16083 (
		_w20082_,
		_w20101_,
		_w20130_
	);
	LUT2 #(
		.INIT('h4)
	) name16084 (
		_w20105_,
		_w20108_,
		_w20131_
	);
	LUT2 #(
		.INIT('h1)
	) name16085 (
		_w20109_,
		_w20113_,
		_w20132_
	);
	LUT2 #(
		.INIT('h8)
	) name16086 (
		_w20131_,
		_w20132_,
		_w20133_
	);
	LUT2 #(
		.INIT('h8)
	) name16087 (
		_w20129_,
		_w20130_,
		_w20134_
	);
	LUT2 #(
		.INIT('h8)
	) name16088 (
		_w20127_,
		_w20128_,
		_w20135_
	);
	LUT2 #(
		.INIT('h2)
	) name16089 (
		_w20087_,
		_w20112_,
		_w20136_
	);
	LUT2 #(
		.INIT('h8)
	) name16090 (
		_w20135_,
		_w20136_,
		_w20137_
	);
	LUT2 #(
		.INIT('h8)
	) name16091 (
		_w20133_,
		_w20134_,
		_w20138_
	);
	LUT2 #(
		.INIT('h8)
	) name16092 (
		_w20137_,
		_w20138_,
		_w20139_
	);
	LUT2 #(
		.INIT('h8)
	) name16093 (
		_w19975_,
		_w20090_,
		_w20140_
	);
	LUT2 #(
		.INIT('h8)
	) name16094 (
		_w20139_,
		_w20140_,
		_w20141_
	);
	LUT2 #(
		.INIT('h8)
	) name16095 (
		_w20107_,
		_w20141_,
		_w20142_
	);
	LUT2 #(
		.INIT('h4)
	) name16096 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w20142_,
		_w20143_
	);
	LUT2 #(
		.INIT('h1)
	) name16097 (
		_w20081_,
		_w20143_,
		_w20144_
	);
	LUT2 #(
		.INIT('h2)
	) name16098 (
		_w18717_,
		_w20144_,
		_w20145_
	);
	LUT2 #(
		.INIT('h1)
	) name16099 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[4]/P0001 ,
		_w18717_,
		_w20146_
	);
	LUT2 #(
		.INIT('h1)
	) name16100 (
		_w20145_,
		_w20146_,
		_w20147_
	);
	LUT2 #(
		.INIT('h1)
	) name16101 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12688_,
		_w20148_
	);
	LUT2 #(
		.INIT('h2)
	) name16102 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12715_,
		_w20149_
	);
	LUT2 #(
		.INIT('h1)
	) name16103 (
		_w20148_,
		_w20149_,
		_w20150_
	);
	LUT2 #(
		.INIT('h2)
	) name16104 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w20150_,
		_w20151_
	);
	LUT2 #(
		.INIT('h4)
	) name16105 (
		_w17938_,
		_w18176_,
		_w20152_
	);
	LUT2 #(
		.INIT('h4)
	) name16106 (
		_w17922_,
		_w18766_,
		_w20153_
	);
	LUT2 #(
		.INIT('h8)
	) name16107 (
		_w18106_,
		_w18905_,
		_w20154_
	);
	LUT2 #(
		.INIT('h1)
	) name16108 (
		_w18159_,
		_w18919_,
		_w20155_
	);
	LUT2 #(
		.INIT('h4)
	) name16109 (
		_w18121_,
		_w18746_,
		_w20156_
	);
	LUT2 #(
		.INIT('h1)
	) name16110 (
		_w18096_,
		_w18743_,
		_w20157_
	);
	LUT2 #(
		.INIT('h4)
	) name16111 (
		_w18133_,
		_w19862_,
		_w20158_
	);
	LUT2 #(
		.INIT('h8)
	) name16112 (
		_w18146_,
		_w19976_,
		_w20159_
	);
	LUT2 #(
		.INIT('h1)
	) name16113 (
		_w17922_,
		_w17924_,
		_w20160_
	);
	LUT2 #(
		.INIT('h1)
	) name16114 (
		_w18121_,
		_w18123_,
		_w20161_
	);
	LUT2 #(
		.INIT('h2)
	) name16115 (
		_w18107_,
		_w18110_,
		_w20162_
	);
	LUT2 #(
		.INIT('h1)
	) name16116 (
		_w18133_,
		_w18170_,
		_w20163_
	);
	LUT2 #(
		.INIT('h1)
	) name16117 (
		_w18180_,
		_w18182_,
		_w20164_
	);
	LUT2 #(
		.INIT('h2)
	) name16118 (
		_w17931_,
		_w20162_,
		_w20165_
	);
	LUT2 #(
		.INIT('h4)
	) name16119 (
		_w20160_,
		_w20165_,
		_w20166_
	);
	LUT2 #(
		.INIT('h1)
	) name16120 (
		_w20161_,
		_w20163_,
		_w20167_
	);
	LUT2 #(
		.INIT('h4)
	) name16121 (
		_w20164_,
		_w20167_,
		_w20168_
	);
	LUT2 #(
		.INIT('h8)
	) name16122 (
		_w20166_,
		_w20168_,
		_w20169_
	);
	LUT2 #(
		.INIT('h2)
	) name16123 (
		_w18751_,
		_w19735_,
		_w20170_
	);
	LUT2 #(
		.INIT('h1)
	) name16124 (
		_w17931_,
		_w19747_,
		_w20171_
	);
	LUT2 #(
		.INIT('h4)
	) name16125 (
		_w20170_,
		_w20171_,
		_w20172_
	);
	LUT2 #(
		.INIT('h1)
	) name16126 (
		_w20169_,
		_w20172_,
		_w20173_
	);
	LUT2 #(
		.INIT('h2)
	) name16127 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11854_,
		_w20174_
	);
	LUT2 #(
		.INIT('h4)
	) name16128 (
		_w18108_,
		_w18749_,
		_w20175_
	);
	LUT2 #(
		.INIT('h4)
	) name16129 (
		_w18092_,
		_w19725_,
		_w20176_
	);
	LUT2 #(
		.INIT('h2)
	) name16130 (
		_w17945_,
		_w20176_,
		_w20177_
	);
	LUT2 #(
		.INIT('h1)
	) name16131 (
		_w20154_,
		_w20174_,
		_w20178_
	);
	LUT2 #(
		.INIT('h4)
	) name16132 (
		_w20153_,
		_w20178_,
		_w20179_
	);
	LUT2 #(
		.INIT('h1)
	) name16133 (
		_w20155_,
		_w20156_,
		_w20180_
	);
	LUT2 #(
		.INIT('h1)
	) name16134 (
		_w20157_,
		_w20158_,
		_w20181_
	);
	LUT2 #(
		.INIT('h4)
	) name16135 (
		_w20175_,
		_w20181_,
		_w20182_
	);
	LUT2 #(
		.INIT('h8)
	) name16136 (
		_w20179_,
		_w20180_,
		_w20183_
	);
	LUT2 #(
		.INIT('h2)
	) name16137 (
		_w18059_,
		_w20152_,
		_w20184_
	);
	LUT2 #(
		.INIT('h8)
	) name16138 (
		_w20183_,
		_w20184_,
		_w20185_
	);
	LUT2 #(
		.INIT('h4)
	) name16139 (
		_w20177_,
		_w20182_,
		_w20186_
	);
	LUT2 #(
		.INIT('h8)
	) name16140 (
		_w20185_,
		_w20186_,
		_w20187_
	);
	LUT2 #(
		.INIT('h8)
	) name16141 (
		_w18006_,
		_w20187_,
		_w20188_
	);
	LUT2 #(
		.INIT('h2)
	) name16142 (
		_w18087_,
		_w20173_,
		_w20189_
	);
	LUT2 #(
		.INIT('h8)
	) name16143 (
		_w20188_,
		_w20189_,
		_w20190_
	);
	LUT2 #(
		.INIT('h8)
	) name16144 (
		_w19715_,
		_w20159_,
		_w20191_
	);
	LUT2 #(
		.INIT('h8)
	) name16145 (
		_w20190_,
		_w20191_,
		_w20192_
	);
	LUT2 #(
		.INIT('h4)
	) name16146 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w20192_,
		_w20193_
	);
	LUT2 #(
		.INIT('h1)
	) name16147 (
		_w20151_,
		_w20193_,
		_w20194_
	);
	LUT2 #(
		.INIT('h2)
	) name16148 (
		_w18717_,
		_w20194_,
		_w20195_
	);
	LUT2 #(
		.INIT('h1)
	) name16149 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[14]/P0001 ,
		_w18717_,
		_w20196_
	);
	LUT2 #(
		.INIT('h1)
	) name16150 (
		_w20195_,
		_w20196_,
		_w20197_
	);
	LUT2 #(
		.INIT('h2)
	) name16151 (
		_w17833_,
		_w20032_,
		_w20198_
	);
	LUT2 #(
		.INIT('h1)
	) name16152 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[7]/P0001 ,
		_w17833_,
		_w20199_
	);
	LUT2 #(
		.INIT('h1)
	) name16153 (
		_w20198_,
		_w20199_,
		_w20200_
	);
	LUT2 #(
		.INIT('h1)
	) name16154 (
		_w5581_,
		_w5586_,
		_w20201_
	);
	LUT2 #(
		.INIT('h1)
	) name16155 (
		_w5519_,
		_w5587_,
		_w20202_
	);
	LUT2 #(
		.INIT('h4)
	) name16156 (
		_w20201_,
		_w20202_,
		_w20203_
	);
	LUT2 #(
		.INIT('h8)
	) name16157 (
		_w5605_,
		_w20203_,
		_w20204_
	);
	LUT2 #(
		.INIT('h4)
	) name16158 (
		_w5581_,
		_w13749_,
		_w20205_
	);
	LUT2 #(
		.INIT('h8)
	) name16159 (
		_w5586_,
		_w20205_,
		_w20206_
	);
	LUT2 #(
		.INIT('h4)
	) name16160 (
		_w12444_,
		_w20206_,
		_w20207_
	);
	LUT2 #(
		.INIT('h4)
	) name16161 (
		_w5586_,
		_w20205_,
		_w20208_
	);
	LUT2 #(
		.INIT('h4)
	) name16162 (
		_w5582_,
		_w20208_,
		_w20209_
	);
	LUT2 #(
		.INIT('h1)
	) name16163 (
		_w13750_,
		_w20204_,
		_w20210_
	);
	LUT2 #(
		.INIT('h4)
	) name16164 (
		_w20207_,
		_w20210_,
		_w20211_
	);
	LUT2 #(
		.INIT('h4)
	) name16165 (
		_w20209_,
		_w20211_,
		_w20212_
	);
	LUT2 #(
		.INIT('h4)
	) name16166 (
		_w5523_,
		_w5583_,
		_w20213_
	);
	LUT2 #(
		.INIT('h2)
	) name16167 (
		\emc_RWcnt_reg[0]/P0001 ,
		_w20213_,
		_w20214_
	);
	LUT2 #(
		.INIT('h8)
	) name16168 (
		\emc_RWcnt_reg[1]/P0001 ,
		_w20214_,
		_w20215_
	);
	LUT2 #(
		.INIT('h8)
	) name16169 (
		\emc_RWcnt_reg[2]/P0001 ,
		_w20215_,
		_w20216_
	);
	LUT2 #(
		.INIT('h8)
	) name16170 (
		\emc_RWcnt_reg[3]/P0001 ,
		_w20216_,
		_w20217_
	);
	LUT2 #(
		.INIT('h8)
	) name16171 (
		\emc_RWcnt_reg[4]/P0001 ,
		_w20217_,
		_w20218_
	);
	LUT2 #(
		.INIT('h1)
	) name16172 (
		\emc_RWcnt_reg[5]/P0001 ,
		_w20218_,
		_w20219_
	);
	LUT2 #(
		.INIT('h8)
	) name16173 (
		\emc_RWcnt_reg[5]/P0001 ,
		_w20218_,
		_w20220_
	);
	LUT2 #(
		.INIT('h1)
	) name16174 (
		_w20219_,
		_w20220_,
		_w20221_
	);
	LUT2 #(
		.INIT('h8)
	) name16175 (
		_w20212_,
		_w20221_,
		_w20222_
	);
	LUT2 #(
		.INIT('h1)
	) name16176 (
		\emc_RWcnt_reg[4]/P0001 ,
		_w20217_,
		_w20223_
	);
	LUT2 #(
		.INIT('h1)
	) name16177 (
		_w20218_,
		_w20223_,
		_w20224_
	);
	LUT2 #(
		.INIT('h8)
	) name16178 (
		_w20212_,
		_w20224_,
		_w20225_
	);
	LUT2 #(
		.INIT('h2)
	) name16179 (
		_w17833_,
		_w20144_,
		_w20226_
	);
	LUT2 #(
		.INIT('h1)
	) name16180 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[4]/P0001 ,
		_w17833_,
		_w20227_
	);
	LUT2 #(
		.INIT('h1)
	) name16181 (
		_w20226_,
		_w20227_,
		_w20228_
	);
	LUT2 #(
		.INIT('h2)
	) name16182 (
		_w17833_,
		_w20194_,
		_w20229_
	);
	LUT2 #(
		.INIT('h1)
	) name16183 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[14]/P0001 ,
		_w17833_,
		_w20230_
	);
	LUT2 #(
		.INIT('h1)
	) name16184 (
		_w20229_,
		_w20230_,
		_w20231_
	);
	LUT2 #(
		.INIT('h8)
	) name16185 (
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		_w19438_,
		_w20232_
	);
	LUT2 #(
		.INIT('h8)
	) name16186 (
		\sport1_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		_w20232_,
		_w20233_
	);
	LUT2 #(
		.INIT('h8)
	) name16187 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		_w20233_,
		_w20234_
	);
	LUT2 #(
		.INIT('h8)
	) name16188 (
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		_w20234_,
		_w20235_
	);
	LUT2 #(
		.INIT('h8)
	) name16189 (
		\sport1_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		_w20235_,
		_w20236_
	);
	LUT2 #(
		.INIT('h8)
	) name16190 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		_w20236_,
		_w20237_
	);
	LUT2 #(
		.INIT('h8)
	) name16191 (
		\sport1_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		_w20237_,
		_w20238_
	);
	LUT2 #(
		.INIT('h1)
	) name16192 (
		\sport1_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		_w20238_,
		_w20239_
	);
	LUT2 #(
		.INIT('h8)
	) name16193 (
		\sport1_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		_w20238_,
		_w20240_
	);
	LUT2 #(
		.INIT('h2)
	) name16194 (
		_w19130_,
		_w20239_,
		_w20241_
	);
	LUT2 #(
		.INIT('h4)
	) name16195 (
		_w20240_,
		_w20241_,
		_w20242_
	);
	LUT2 #(
		.INIT('h1)
	) name16196 (
		\sport1_cfg_SCLKi_cnt_reg[5]/NET0131 ,
		_w20234_,
		_w20243_
	);
	LUT2 #(
		.INIT('h1)
	) name16197 (
		_w20235_,
		_w20243_,
		_w20244_
	);
	LUT2 #(
		.INIT('h8)
	) name16198 (
		_w19130_,
		_w20244_,
		_w20245_
	);
	LUT2 #(
		.INIT('h1)
	) name16199 (
		\sport1_cfg_SCLKi_cnt_reg[2]/NET0131 ,
		_w19438_,
		_w20246_
	);
	LUT2 #(
		.INIT('h1)
	) name16200 (
		_w20232_,
		_w20246_,
		_w20247_
	);
	LUT2 #(
		.INIT('h8)
	) name16201 (
		_w19130_,
		_w20247_,
		_w20248_
	);
	LUT2 #(
		.INIT('h8)
	) name16202 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		_w20240_,
		_w20249_
	);
	LUT2 #(
		.INIT('h8)
	) name16203 (
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		_w20249_,
		_w20250_
	);
	LUT2 #(
		.INIT('h8)
	) name16204 (
		\sport1_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		_w20250_,
		_w20251_
	);
	LUT2 #(
		.INIT('h1)
	) name16205 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		_w20251_,
		_w20252_
	);
	LUT2 #(
		.INIT('h8)
	) name16206 (
		\sport1_cfg_SCLKi_cnt_reg[13]/NET0131 ,
		_w20251_,
		_w20253_
	);
	LUT2 #(
		.INIT('h2)
	) name16207 (
		_w19130_,
		_w20252_,
		_w20254_
	);
	LUT2 #(
		.INIT('h4)
	) name16208 (
		_w20253_,
		_w20254_,
		_w20255_
	);
	LUT2 #(
		.INIT('h4)
	) name16209 (
		\sport1_cfg_SCLKi_cnt_reg[0]/NET0131 ,
		_w19130_,
		_w20256_
	);
	LUT2 #(
		.INIT('h1)
	) name16210 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w10911_,
		_w20257_
	);
	LUT2 #(
		.INIT('h2)
	) name16211 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12938_,
		_w20258_
	);
	LUT2 #(
		.INIT('h1)
	) name16212 (
		_w20257_,
		_w20258_,
		_w20259_
	);
	LUT2 #(
		.INIT('h2)
	) name16213 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w20259_,
		_w20260_
	);
	LUT2 #(
		.INIT('h2)
	) name16214 (
		_w18765_,
		_w18888_,
		_w20261_
	);
	LUT2 #(
		.INIT('h1)
	) name16215 (
		_w18167_,
		_w18918_,
		_w20262_
	);
	LUT2 #(
		.INIT('h2)
	) name16216 (
		_w17930_,
		_w18909_,
		_w20263_
	);
	LUT2 #(
		.INIT('h2)
	) name16217 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w10801_,
		_w20264_
	);
	LUT2 #(
		.INIT('h1)
	) name16218 (
		_w18189_,
		_w18914_,
		_w20265_
	);
	LUT2 #(
		.INIT('h1)
	) name16219 (
		_w18079_,
		_w18117_,
		_w20266_
	);
	LUT2 #(
		.INIT('h4)
	) name16220 (
		_w17998_,
		_w18758_,
		_w20267_
	);
	LUT2 #(
		.INIT('h2)
	) name16221 (
		_w18171_,
		_w18898_,
		_w20268_
	);
	LUT2 #(
		.INIT('h1)
	) name16222 (
		_w18104_,
		_w18907_,
		_w20269_
	);
	LUT2 #(
		.INIT('h4)
	) name16223 (
		_w17933_,
		_w18922_,
		_w20270_
	);
	LUT2 #(
		.INIT('h8)
	) name16224 (
		_w17991_,
		_w18088_,
		_w20271_
	);
	LUT2 #(
		.INIT('h8)
	) name16225 (
		_w17965_,
		_w17992_,
		_w20272_
	);
	LUT2 #(
		.INIT('h1)
	) name16226 (
		_w18129_,
		_w18912_,
		_w20273_
	);
	LUT2 #(
		.INIT('h8)
	) name16227 (
		_w18797_,
		_w18904_,
		_w20274_
	);
	LUT2 #(
		.INIT('h1)
	) name16228 (
		_w20264_,
		_w20272_,
		_w20275_
	);
	LUT2 #(
		.INIT('h4)
	) name16229 (
		_w18890_,
		_w20275_,
		_w20276_
	);
	LUT2 #(
		.INIT('h1)
	) name16230 (
		_w20262_,
		_w20263_,
		_w20277_
	);
	LUT2 #(
		.INIT('h1)
	) name16231 (
		_w20265_,
		_w20266_,
		_w20278_
	);
	LUT2 #(
		.INIT('h1)
	) name16232 (
		_w20269_,
		_w20271_,
		_w20279_
	);
	LUT2 #(
		.INIT('h4)
	) name16233 (
		_w20273_,
		_w20279_,
		_w20280_
	);
	LUT2 #(
		.INIT('h8)
	) name16234 (
		_w20277_,
		_w20278_,
		_w20281_
	);
	LUT2 #(
		.INIT('h4)
	) name16235 (
		_w20261_,
		_w20276_,
		_w20282_
	);
	LUT2 #(
		.INIT('h1)
	) name16236 (
		_w20267_,
		_w20268_,
		_w20283_
	);
	LUT2 #(
		.INIT('h4)
	) name16237 (
		_w20270_,
		_w20283_,
		_w20284_
	);
	LUT2 #(
		.INIT('h8)
	) name16238 (
		_w20281_,
		_w20282_,
		_w20285_
	);
	LUT2 #(
		.INIT('h8)
	) name16239 (
		_w20280_,
		_w20285_,
		_w20286_
	);
	LUT2 #(
		.INIT('h8)
	) name16240 (
		_w20284_,
		_w20286_,
		_w20287_
	);
	LUT2 #(
		.INIT('h8)
	) name16241 (
		_w20274_,
		_w20287_,
		_w20288_
	);
	LUT2 #(
		.INIT('h4)
	) name16242 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w20288_,
		_w20289_
	);
	LUT2 #(
		.INIT('h1)
	) name16243 (
		_w20260_,
		_w20289_,
		_w20290_
	);
	LUT2 #(
		.INIT('h2)
	) name16244 (
		_w18886_,
		_w20290_,
		_w20291_
	);
	LUT2 #(
		.INIT('h1)
	) name16245 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[5]/P0001 ,
		_w18886_,
		_w20292_
	);
	LUT2 #(
		.INIT('h1)
	) name16246 (
		_w20291_,
		_w20292_,
		_w20293_
	);
	LUT2 #(
		.INIT('h2)
	) name16247 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w19559_,
		_w20294_
	);
	LUT2 #(
		.INIT('h2)
	) name16248 (
		_w18759_,
		_w18909_,
		_w20295_
	);
	LUT2 #(
		.INIT('h2)
	) name16249 (
		_w18745_,
		_w18898_,
		_w20296_
	);
	LUT2 #(
		.INIT('h1)
	) name16250 (
		_w18082_,
		_w19870_,
		_w20297_
	);
	LUT2 #(
		.INIT('h2)
	) name16251 (
		_w18765_,
		_w18981_,
		_w20298_
	);
	LUT2 #(
		.INIT('h1)
	) name16252 (
		_w18079_,
		_w18919_,
		_w20299_
	);
	LUT2 #(
		.INIT('h1)
	) name16253 (
		_w18743_,
		_w18914_,
		_w20300_
	);
	LUT2 #(
		.INIT('h8)
	) name16254 (
		_w17991_,
		_w18115_,
		_w20301_
	);
	LUT2 #(
		.INIT('h2)
	) name16255 (
		_w17925_,
		_w18983_,
		_w20302_
	);
	LUT2 #(
		.INIT('h2)
	) name16256 (
		_w18171_,
		_w18888_,
		_w20303_
	);
	LUT2 #(
		.INIT('h2)
	) name16257 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7381_,
		_w20304_
	);
	LUT2 #(
		.INIT('h2)
	) name16258 (
		_w18754_,
		_w18909_,
		_w20305_
	);
	LUT2 #(
		.INIT('h4)
	) name16259 (
		_w17998_,
		_w18124_,
		_w20306_
	);
	LUT2 #(
		.INIT('h2)
	) name16260 (
		_w18752_,
		_w18918_,
		_w20307_
	);
	LUT2 #(
		.INIT('h8)
	) name16261 (
		_w17929_,
		_w18088_,
		_w20308_
	);
	LUT2 #(
		.INIT('h1)
	) name16262 (
		_w17965_,
		_w20308_,
		_w20309_
	);
	LUT2 #(
		.INIT('h1)
	) name16263 (
		_w17970_,
		_w18017_,
		_w20310_
	);
	LUT2 #(
		.INIT('h1)
	) name16264 (
		_w20309_,
		_w20310_,
		_w20311_
	);
	LUT2 #(
		.INIT('h1)
	) name16265 (
		_w18900_,
		_w20304_,
		_w20312_
	);
	LUT2 #(
		.INIT('h8)
	) name16266 (
		_w18016_,
		_w20312_,
		_w20313_
	);
	LUT2 #(
		.INIT('h1)
	) name16267 (
		_w20295_,
		_w20297_,
		_w20314_
	);
	LUT2 #(
		.INIT('h1)
	) name16268 (
		_w20299_,
		_w20300_,
		_w20315_
	);
	LUT2 #(
		.INIT('h1)
	) name16269 (
		_w20301_,
		_w20305_,
		_w20316_
	);
	LUT2 #(
		.INIT('h1)
	) name16270 (
		_w20307_,
		_w20311_,
		_w20317_
	);
	LUT2 #(
		.INIT('h8)
	) name16271 (
		_w20316_,
		_w20317_,
		_w20318_
	);
	LUT2 #(
		.INIT('h8)
	) name16272 (
		_w20314_,
		_w20315_,
		_w20319_
	);
	LUT2 #(
		.INIT('h4)
	) name16273 (
		_w20296_,
		_w20313_,
		_w20320_
	);
	LUT2 #(
		.INIT('h1)
	) name16274 (
		_w20298_,
		_w20302_,
		_w20321_
	);
	LUT2 #(
		.INIT('h1)
	) name16275 (
		_w20303_,
		_w20306_,
		_w20322_
	);
	LUT2 #(
		.INIT('h8)
	) name16276 (
		_w20321_,
		_w20322_,
		_w20323_
	);
	LUT2 #(
		.INIT('h8)
	) name16277 (
		_w20319_,
		_w20320_,
		_w20324_
	);
	LUT2 #(
		.INIT('h8)
	) name16278 (
		_w20318_,
		_w20324_,
		_w20325_
	);
	LUT2 #(
		.INIT('h8)
	) name16279 (
		_w20323_,
		_w20325_,
		_w20326_
	);
	LUT2 #(
		.INIT('h4)
	) name16280 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w20326_,
		_w20327_
	);
	LUT2 #(
		.INIT('h1)
	) name16281 (
		_w20294_,
		_w20327_,
		_w20328_
	);
	LUT2 #(
		.INIT('h2)
	) name16282 (
		_w18886_,
		_w20328_,
		_w20329_
	);
	LUT2 #(
		.INIT('h1)
	) name16283 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[0]/P0001 ,
		_w18886_,
		_w20330_
	);
	LUT2 #(
		.INIT('h1)
	) name16284 (
		_w20329_,
		_w20330_,
		_w20331_
	);
	LUT2 #(
		.INIT('h2)
	) name16285 (
		_w19034_,
		_w20290_,
		_w20332_
	);
	LUT2 #(
		.INIT('h1)
	) name16286 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[5]/P0001 ,
		_w19034_,
		_w20333_
	);
	LUT2 #(
		.INIT('h1)
	) name16287 (
		_w20332_,
		_w20333_,
		_w20334_
	);
	LUT2 #(
		.INIT('h2)
	) name16288 (
		_w19034_,
		_w20328_,
		_w20335_
	);
	LUT2 #(
		.INIT('h1)
	) name16289 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[0]/P0001 ,
		_w19034_,
		_w20336_
	);
	LUT2 #(
		.INIT('h1)
	) name16290 (
		_w20335_,
		_w20336_,
		_w20337_
	);
	LUT2 #(
		.INIT('h1)
	) name16291 (
		\sport0_cfg_SCLKi_cnt_reg[9]/NET0131 ,
		_w19546_,
		_w20338_
	);
	LUT2 #(
		.INIT('h2)
	) name16292 (
		_w19197_,
		_w19547_,
		_w20339_
	);
	LUT2 #(
		.INIT('h4)
	) name16293 (
		_w20338_,
		_w20339_,
		_w20340_
	);
	LUT2 #(
		.INIT('h8)
	) name16294 (
		\emc_PMcst_reg/NET0131 ,
		_w14733_,
		_w20341_
	);
	LUT2 #(
		.INIT('h2)
	) name16295 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w4068_,
		_w20342_
	);
	LUT2 #(
		.INIT('h8)
	) name16296 (
		_w19041_,
		_w20342_,
		_w20343_
	);
	LUT2 #(
		.INIT('h8)
	) name16297 (
		\memc_Pread_E_reg/NET0131 ,
		_w20343_,
		_w20344_
	);
	LUT2 #(
		.INIT('h8)
	) name16298 (
		_w19049_,
		_w20344_,
		_w20345_
	);
	LUT2 #(
		.INIT('h8)
	) name16299 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w20343_,
		_w20346_
	);
	LUT2 #(
		.INIT('h8)
	) name16300 (
		_w19049_,
		_w20346_,
		_w20347_
	);
	LUT2 #(
		.INIT('h2)
	) name16301 (
		\emc_PMcst_reg/NET0131 ,
		_w5593_,
		_w20348_
	);
	LUT2 #(
		.INIT('h4)
	) name16302 (
		_w5604_,
		_w20348_,
		_w20349_
	);
	LUT2 #(
		.INIT('h4)
	) name16303 (
		_w19049_,
		_w20349_,
		_w20350_
	);
	LUT2 #(
		.INIT('h1)
	) name16304 (
		_w20341_,
		_w20345_,
		_w20351_
	);
	LUT2 #(
		.INIT('h1)
	) name16305 (
		_w20347_,
		_w20350_,
		_w20352_
	);
	LUT2 #(
		.INIT('h8)
	) name16306 (
		_w20351_,
		_w20352_,
		_w20353_
	);
	LUT2 #(
		.INIT('h4)
	) name16307 (
		\T_TMODE[0]_pad ,
		\tm_WR_TCR_TMP_GEN1_reg/P0001 ,
		_w20354_
	);
	LUT2 #(
		.INIT('h4)
	) name16308 (
		\tm_WR_TCR_TMP_GEN2_reg/P0001 ,
		_w20354_,
		_w20355_
	);
	LUT2 #(
		.INIT('h4)
	) name16309 (
		\T_TMODE[0]_pad ,
		\tm_WR_TSR_TMP_GEN1_reg/P0001 ,
		_w20356_
	);
	LUT2 #(
		.INIT('h4)
	) name16310 (
		\tm_WR_TSR_TMP_GEN2_reg/P0001 ,
		_w20356_,
		_w20357_
	);
	LUT2 #(
		.INIT('h1)
	) name16311 (
		\tm_TCR_TMP_reg[1]/NET0131 ,
		\tm_TCR_TMP_reg[2]/NET0131 ,
		_w20358_
	);
	LUT2 #(
		.INIT('h4)
	) name16312 (
		\tm_TCR_TMP_reg[3]/NET0131 ,
		_w20358_,
		_w20359_
	);
	LUT2 #(
		.INIT('h4)
	) name16313 (
		\tm_TCR_TMP_reg[0]/NET0131 ,
		_w20359_,
		_w20360_
	);
	LUT2 #(
		.INIT('h1)
	) name16314 (
		\tm_TCR_TMP_reg[4]/NET0131 ,
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w20361_
	);
	LUT2 #(
		.INIT('h1)
	) name16315 (
		\tm_TCR_TMP_reg[6]/NET0131 ,
		\tm_TCR_TMP_reg[7]/NET0131 ,
		_w20362_
	);
	LUT2 #(
		.INIT('h8)
	) name16316 (
		_w20361_,
		_w20362_,
		_w20363_
	);
	LUT2 #(
		.INIT('h8)
	) name16317 (
		_w20360_,
		_w20363_,
		_w20364_
	);
	LUT2 #(
		.INIT('h1)
	) name16318 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		\tm_TCR_TMP_reg[11]/NET0131 ,
		_w20365_
	);
	LUT2 #(
		.INIT('h1)
	) name16319 (
		\tm_TCR_TMP_reg[12]/NET0131 ,
		\tm_TCR_TMP_reg[13]/NET0131 ,
		_w20366_
	);
	LUT2 #(
		.INIT('h1)
	) name16320 (
		\tm_TCR_TMP_reg[14]/NET0131 ,
		\tm_TCR_TMP_reg[15]/NET0131 ,
		_w20367_
	);
	LUT2 #(
		.INIT('h1)
	) name16321 (
		\tm_TCR_TMP_reg[8]/NET0131 ,
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w20368_
	);
	LUT2 #(
		.INIT('h8)
	) name16322 (
		_w20367_,
		_w20368_,
		_w20369_
	);
	LUT2 #(
		.INIT('h8)
	) name16323 (
		_w20365_,
		_w20366_,
		_w20370_
	);
	LUT2 #(
		.INIT('h8)
	) name16324 (
		_w20369_,
		_w20370_,
		_w20371_
	);
	LUT2 #(
		.INIT('h8)
	) name16325 (
		_w20364_,
		_w20371_,
		_w20372_
	);
	LUT2 #(
		.INIT('h2)
	) name16326 (
		\tm_MSTAT5_syn_reg/NET0131 ,
		_w20355_,
		_w20373_
	);
	LUT2 #(
		.INIT('h4)
	) name16327 (
		_w20357_,
		_w20373_,
		_w20374_
	);
	LUT2 #(
		.INIT('h8)
	) name16328 (
		_w20372_,
		_w20374_,
		_w20375_
	);
	LUT2 #(
		.INIT('h8)
	) name16329 (
		\core_c_dec_updAF_E_reg/P0001 ,
		_w4118_,
		_w20376_
	);
	LUT2 #(
		.INIT('h2)
	) name16330 (
		_w5664_,
		_w18842_,
		_w20377_
	);
	LUT2 #(
		.INIT('h8)
	) name16331 (
		_w4116_,
		_w18849_,
		_w20378_
	);
	LUT2 #(
		.INIT('h8)
	) name16332 (
		_w20377_,
		_w20378_,
		_w20379_
	);
	LUT2 #(
		.INIT('h1)
	) name16333 (
		_w20376_,
		_w20379_,
		_w20380_
	);
	LUT2 #(
		.INIT('h1)
	) name16334 (
		\idma_WRcnt_reg[0]/NET0131 ,
		\idma_WRcnt_reg[1]/NET0131 ,
		_w20381_
	);
	LUT2 #(
		.INIT('h4)
	) name16335 (
		\idma_WRcnt_reg[2]/NET0131 ,
		_w20381_,
		_w20382_
	);
	LUT2 #(
		.INIT('h2)
	) name16336 (
		\idma_WRtrue_reg/NET0131 ,
		_w20382_,
		_w20383_
	);
	LUT2 #(
		.INIT('h4)
	) name16337 (
		\idma_WRCMD_d1_reg/P0001 ,
		\idma_WRCMD_reg/P0001 ,
		_w20384_
	);
	LUT2 #(
		.INIT('h1)
	) name16338 (
		_w20383_,
		_w20384_,
		_w20385_
	);
	LUT2 #(
		.INIT('h1)
	) name16339 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		_w20386_
	);
	LUT2 #(
		.INIT('h1)
	) name16340 (
		\idma_ISn_reg/P0001 ,
		\idma_IWRn_reg/P0001 ,
		_w20387_
	);
	LUT2 #(
		.INIT('h8)
	) name16341 (
		\idma_WRtrue_reg/NET0131 ,
		_w20387_,
		_w20388_
	);
	LUT2 #(
		.INIT('h2)
	) name16342 (
		\auctl_DSack_reg/NET0131 ,
		_w20386_,
		_w20389_
	);
	LUT2 #(
		.INIT('h1)
	) name16343 (
		\idma_RDcnt_reg[0]/NET0131 ,
		\idma_RDcnt_reg[1]/NET0131 ,
		_w20390_
	);
	LUT2 #(
		.INIT('h4)
	) name16344 (
		\idma_RDcnt_reg[2]/NET0131 ,
		_w20386_,
		_w20391_
	);
	LUT2 #(
		.INIT('h8)
	) name16345 (
		_w20390_,
		_w20391_,
		_w20392_
	);
	LUT2 #(
		.INIT('h1)
	) name16346 (
		_w20389_,
		_w20392_,
		_w20393_
	);
	LUT2 #(
		.INIT('h2)
	) name16347 (
		\idma_RDcyc_reg/NET0131 ,
		_w20393_,
		_w20394_
	);
	LUT2 #(
		.INIT('h1)
	) name16348 (
		_w20388_,
		_w20394_,
		_w20395_
	);
	LUT2 #(
		.INIT('h1)
	) name16349 (
		_w20386_,
		_w20395_,
		_w20396_
	);
	LUT2 #(
		.INIT('h2)
	) name16350 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[0]/P0001 ,
		_w18848_,
		_w20397_
	);
	LUT2 #(
		.INIT('h8)
	) name16351 (
		_w18843_,
		_w18848_,
		_w20398_
	);
	LUT2 #(
		.INIT('h1)
	) name16352 (
		_w20397_,
		_w20398_,
		_w20399_
	);
	LUT2 #(
		.INIT('h8)
	) name16353 (
		_w7226_,
		_w20070_,
		_w20400_
	);
	LUT2 #(
		.INIT('h8)
	) name16354 (
		_w18226_,
		_w20400_,
		_w20401_
	);
	LUT2 #(
		.INIT('h4)
	) name16355 (
		\memc_MMR_web_reg/NET0131 ,
		_w20401_,
		_w20402_
	);
	LUT2 #(
		.INIT('h4)
	) name16356 (
		_w10289_,
		_w20402_,
		_w20403_
	);
	LUT2 #(
		.INIT('h1)
	) name16357 (
		\sport0_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w20402_,
		_w20404_
	);
	LUT2 #(
		.INIT('h1)
	) name16358 (
		_w20403_,
		_w20404_,
		_w20405_
	);
	LUT2 #(
		.INIT('h1)
	) name16359 (
		\sport1_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[5]/NET0131 ,
		_w20406_
	);
	LUT2 #(
		.INIT('h4)
	) name16360 (
		\sport1_rxctl_Wcnt_reg[6]/NET0131 ,
		_w20406_,
		_w20407_
	);
	LUT2 #(
		.INIT('h4)
	) name16361 (
		\sport1_rxctl_Wcnt_reg[7]/NET0131 ,
		_w20407_,
		_w20408_
	);
	LUT2 #(
		.INIT('h2)
	) name16362 (
		\sport1_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[2]/NET0131 ,
		_w20409_
	);
	LUT2 #(
		.INIT('h1)
	) name16363 (
		\sport1_rxctl_Bcnt_reg[3]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[4]/NET0131 ,
		_w20410_
	);
	LUT2 #(
		.INIT('h8)
	) name16364 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[1]/NET0131 ,
		_w20411_
	);
	LUT2 #(
		.INIT('h4)
	) name16365 (
		\sport1_rxctl_Wcnt_reg[2]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		_w20412_
	);
	LUT2 #(
		.INIT('h8)
	) name16366 (
		_w20411_,
		_w20412_,
		_w20413_
	);
	LUT2 #(
		.INIT('h8)
	) name16367 (
		_w20409_,
		_w20410_,
		_w20414_
	);
	LUT2 #(
		.INIT('h8)
	) name16368 (
		_w20413_,
		_w20414_,
		_w20415_
	);
	LUT2 #(
		.INIT('h8)
	) name16369 (
		_w20408_,
		_w20415_,
		_w20416_
	);
	LUT2 #(
		.INIT('h4)
	) name16370 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		_w20416_,
		_w20417_
	);
	LUT2 #(
		.INIT('h2)
	) name16371 (
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w13720_,
		_w20418_
	);
	LUT2 #(
		.INIT('h1)
	) name16372 (
		\T_RD1_pad ,
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w20419_
	);
	LUT2 #(
		.INIT('h1)
	) name16373 (
		_w20418_,
		_w20419_,
		_w20420_
	);
	LUT2 #(
		.INIT('h2)
	) name16374 (
		_w20417_,
		_w20420_,
		_w20421_
	);
	LUT2 #(
		.INIT('h1)
	) name16375 (
		\sport1_rxctl_SLOT1_EXT_reg[2]/NET0131 ,
		_w20417_,
		_w20422_
	);
	LUT2 #(
		.INIT('h1)
	) name16376 (
		_w20421_,
		_w20422_,
		_w20423_
	);
	LUT2 #(
		.INIT('h8)
	) name16377 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		_w20416_,
		_w20424_
	);
	LUT2 #(
		.INIT('h4)
	) name16378 (
		_w20420_,
		_w20424_,
		_w20425_
	);
	LUT2 #(
		.INIT('h1)
	) name16379 (
		\sport1_rxctl_SLOT1_EXT_reg[3]/NET0131 ,
		_w20424_,
		_w20426_
	);
	LUT2 #(
		.INIT('h1)
	) name16380 (
		_w20425_,
		_w20426_,
		_w20427_
	);
	LUT2 #(
		.INIT('h1)
	) name16381 (
		\sport0_rxctl_Wcnt_reg[4]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[5]/NET0131 ,
		_w20428_
	);
	LUT2 #(
		.INIT('h4)
	) name16382 (
		\sport0_rxctl_Wcnt_reg[6]/NET0131 ,
		_w20428_,
		_w20429_
	);
	LUT2 #(
		.INIT('h4)
	) name16383 (
		\sport0_rxctl_Wcnt_reg[7]/NET0131 ,
		_w20429_,
		_w20430_
	);
	LUT2 #(
		.INIT('h2)
	) name16384 (
		\sport0_rxctl_Bcnt_reg[1]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[2]/NET0131 ,
		_w20431_
	);
	LUT2 #(
		.INIT('h1)
	) name16385 (
		\sport0_rxctl_Bcnt_reg[3]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[4]/NET0131 ,
		_w20432_
	);
	LUT2 #(
		.INIT('h8)
	) name16386 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[1]/NET0131 ,
		_w20433_
	);
	LUT2 #(
		.INIT('h4)
	) name16387 (
		\sport0_rxctl_Wcnt_reg[2]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		_w20434_
	);
	LUT2 #(
		.INIT('h8)
	) name16388 (
		_w20433_,
		_w20434_,
		_w20435_
	);
	LUT2 #(
		.INIT('h8)
	) name16389 (
		_w20431_,
		_w20432_,
		_w20436_
	);
	LUT2 #(
		.INIT('h8)
	) name16390 (
		_w20435_,
		_w20436_,
		_w20437_
	);
	LUT2 #(
		.INIT('h8)
	) name16391 (
		_w20430_,
		_w20437_,
		_w20438_
	);
	LUT2 #(
		.INIT('h4)
	) name16392 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		_w20438_,
		_w20439_
	);
	LUT2 #(
		.INIT('h2)
	) name16393 (
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w13671_,
		_w20440_
	);
	LUT2 #(
		.INIT('h1)
	) name16394 (
		\T_RD0_pad ,
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w20441_
	);
	LUT2 #(
		.INIT('h1)
	) name16395 (
		_w20440_,
		_w20441_,
		_w20442_
	);
	LUT2 #(
		.INIT('h2)
	) name16396 (
		_w20439_,
		_w20442_,
		_w20443_
	);
	LUT2 #(
		.INIT('h1)
	) name16397 (
		\sport0_rxctl_SLOT1_EXT_reg[2]/NET0131 ,
		_w20439_,
		_w20444_
	);
	LUT2 #(
		.INIT('h1)
	) name16398 (
		_w20443_,
		_w20444_,
		_w20445_
	);
	LUT2 #(
		.INIT('h8)
	) name16399 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		_w20438_,
		_w20446_
	);
	LUT2 #(
		.INIT('h4)
	) name16400 (
		_w20442_,
		_w20446_,
		_w20447_
	);
	LUT2 #(
		.INIT('h1)
	) name16401 (
		\sport0_rxctl_SLOT1_EXT_reg[3]/NET0131 ,
		_w20446_,
		_w20448_
	);
	LUT2 #(
		.INIT('h1)
	) name16402 (
		_w20447_,
		_w20448_,
		_w20449_
	);
	LUT2 #(
		.INIT('h4)
	) name16403 (
		_w10638_,
		_w20402_,
		_w20450_
	);
	LUT2 #(
		.INIT('h1)
	) name16404 (
		\sport0_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w20402_,
		_w20451_
	);
	LUT2 #(
		.INIT('h1)
	) name16405 (
		_w20450_,
		_w20451_,
		_w20452_
	);
	LUT2 #(
		.INIT('h4)
	) name16406 (
		IACKn_pad,
		\idma_IRDn_reg/P0001 ,
		_w20453_
	);
	LUT2 #(
		.INIT('h8)
	) name16407 (
		\idma_IWRn_reg/P0001 ,
		_w20453_,
		_w20454_
	);
	LUT2 #(
		.INIT('h2)
	) name16408 (
		_w20384_,
		_w20454_,
		_w20455_
	);
	LUT2 #(
		.INIT('h2)
	) name16409 (
		\idma_WRtrue_reg/NET0131 ,
		_w20454_,
		_w20456_
	);
	LUT2 #(
		.INIT('h4)
	) name16410 (
		\idma_WRcnt_reg[0]/NET0131 ,
		_w20456_,
		_w20457_
	);
	LUT2 #(
		.INIT('h2)
	) name16411 (
		\idma_WRcnt_reg[1]/NET0131 ,
		_w20457_,
		_w20458_
	);
	LUT2 #(
		.INIT('h8)
	) name16412 (
		_w20381_,
		_w20456_,
		_w20459_
	);
	LUT2 #(
		.INIT('h1)
	) name16413 (
		_w20455_,
		_w20459_,
		_w20460_
	);
	LUT2 #(
		.INIT('h4)
	) name16414 (
		_w20458_,
		_w20460_,
		_w20461_
	);
	LUT2 #(
		.INIT('h4)
	) name16415 (
		\memc_usysr_DO_reg[8]/NET0131 ,
		_w20455_,
		_w20462_
	);
	LUT2 #(
		.INIT('h1)
	) name16416 (
		_w20461_,
		_w20462_,
		_w20463_
	);
	LUT2 #(
		.INIT('h1)
	) name16417 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w20464_
	);
	LUT2 #(
		.INIT('h1)
	) name16418 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w20465_
	);
	LUT2 #(
		.INIT('h8)
	) name16419 (
		_w20464_,
		_w20465_,
		_w20466_
	);
	LUT2 #(
		.INIT('h2)
	) name16420 (
		_w14728_,
		_w20466_,
		_w20467_
	);
	LUT2 #(
		.INIT('h8)
	) name16421 (
		_w5664_,
		_w20467_,
		_w20468_
	);
	LUT2 #(
		.INIT('h2)
	) name16422 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[9]/P0001 ,
		_w20468_,
		_w20469_
	);
	LUT2 #(
		.INIT('h4)
	) name16423 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w20470_
	);
	LUT2 #(
		.INIT('h4)
	) name16424 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w20470_,
		_w20471_
	);
	LUT2 #(
		.INIT('h2)
	) name16425 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w20472_
	);
	LUT2 #(
		.INIT('h8)
	) name16426 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w20472_,
		_w20473_
	);
	LUT2 #(
		.INIT('h8)
	) name16427 (
		_w20471_,
		_w20473_,
		_w20474_
	);
	LUT2 #(
		.INIT('h8)
	) name16428 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w20475_
	);
	LUT2 #(
		.INIT('h4)
	) name16429 (
		_w20471_,
		_w20475_,
		_w20476_
	);
	LUT2 #(
		.INIT('h2)
	) name16430 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w20477_
	);
	LUT2 #(
		.INIT('h8)
	) name16431 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w20477_,
		_w20478_
	);
	LUT2 #(
		.INIT('h1)
	) name16432 (
		_w20474_,
		_w20478_,
		_w20479_
	);
	LUT2 #(
		.INIT('h4)
	) name16433 (
		_w20476_,
		_w20479_,
		_w20480_
	);
	LUT2 #(
		.INIT('h2)
	) name16434 (
		_w20468_,
		_w20480_,
		_w20481_
	);
	LUT2 #(
		.INIT('h1)
	) name16435 (
		_w20469_,
		_w20481_,
		_w20482_
	);
	LUT2 #(
		.INIT('h2)
	) name16436 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[8]/P0001 ,
		_w20468_,
		_w20483_
	);
	LUT2 #(
		.INIT('h8)
	) name16437 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w20464_,
		_w20484_
	);
	LUT2 #(
		.INIT('h8)
	) name16438 (
		_w20471_,
		_w20484_,
		_w20485_
	);
	LUT2 #(
		.INIT('h8)
	) name16439 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w20486_
	);
	LUT2 #(
		.INIT('h8)
	) name16440 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w20486_,
		_w20487_
	);
	LUT2 #(
		.INIT('h1)
	) name16441 (
		_w20476_,
		_w20487_,
		_w20488_
	);
	LUT2 #(
		.INIT('h4)
	) name16442 (
		_w20485_,
		_w20488_,
		_w20489_
	);
	LUT2 #(
		.INIT('h2)
	) name16443 (
		_w20468_,
		_w20489_,
		_w20490_
	);
	LUT2 #(
		.INIT('h1)
	) name16444 (
		_w20483_,
		_w20490_,
		_w20491_
	);
	LUT2 #(
		.INIT('h2)
	) name16445 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[7]/P0001 ,
		_w20468_,
		_w20492_
	);
	LUT2 #(
		.INIT('h2)
	) name16446 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w20493_
	);
	LUT2 #(
		.INIT('h8)
	) name16447 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w20493_,
		_w20494_
	);
	LUT2 #(
		.INIT('h2)
	) name16448 (
		_w20475_,
		_w20494_,
		_w20495_
	);
	LUT2 #(
		.INIT('h8)
	) name16449 (
		_w20473_,
		_w20494_,
		_w20496_
	);
	LUT2 #(
		.INIT('h1)
	) name16450 (
		_w20478_,
		_w20495_,
		_w20497_
	);
	LUT2 #(
		.INIT('h4)
	) name16451 (
		_w20496_,
		_w20497_,
		_w20498_
	);
	LUT2 #(
		.INIT('h2)
	) name16452 (
		_w20468_,
		_w20498_,
		_w20499_
	);
	LUT2 #(
		.INIT('h1)
	) name16453 (
		_w20492_,
		_w20499_,
		_w20500_
	);
	LUT2 #(
		.INIT('h2)
	) name16454 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[6]/P0001 ,
		_w20468_,
		_w20501_
	);
	LUT2 #(
		.INIT('h8)
	) name16455 (
		_w20484_,
		_w20494_,
		_w20502_
	);
	LUT2 #(
		.INIT('h1)
	) name16456 (
		_w20487_,
		_w20495_,
		_w20503_
	);
	LUT2 #(
		.INIT('h4)
	) name16457 (
		_w20502_,
		_w20503_,
		_w20504_
	);
	LUT2 #(
		.INIT('h2)
	) name16458 (
		_w20468_,
		_w20504_,
		_w20505_
	);
	LUT2 #(
		.INIT('h1)
	) name16459 (
		_w20501_,
		_w20505_,
		_w20506_
	);
	LUT2 #(
		.INIT('h2)
	) name16460 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[5]/P0001 ,
		_w20468_,
		_w20507_
	);
	LUT2 #(
		.INIT('h1)
	) name16461 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w20508_
	);
	LUT2 #(
		.INIT('h8)
	) name16462 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w20508_,
		_w20509_
	);
	LUT2 #(
		.INIT('h2)
	) name16463 (
		_w20475_,
		_w20509_,
		_w20510_
	);
	LUT2 #(
		.INIT('h8)
	) name16464 (
		_w20473_,
		_w20509_,
		_w20511_
	);
	LUT2 #(
		.INIT('h1)
	) name16465 (
		_w20478_,
		_w20510_,
		_w20512_
	);
	LUT2 #(
		.INIT('h4)
	) name16466 (
		_w20511_,
		_w20512_,
		_w20513_
	);
	LUT2 #(
		.INIT('h2)
	) name16467 (
		_w20468_,
		_w20513_,
		_w20514_
	);
	LUT2 #(
		.INIT('h1)
	) name16468 (
		_w20507_,
		_w20514_,
		_w20515_
	);
	LUT2 #(
		.INIT('h2)
	) name16469 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[4]/P0001 ,
		_w20468_,
		_w20516_
	);
	LUT2 #(
		.INIT('h8)
	) name16470 (
		_w20484_,
		_w20509_,
		_w20517_
	);
	LUT2 #(
		.INIT('h1)
	) name16471 (
		_w20487_,
		_w20510_,
		_w20518_
	);
	LUT2 #(
		.INIT('h4)
	) name16472 (
		_w20517_,
		_w20518_,
		_w20519_
	);
	LUT2 #(
		.INIT('h2)
	) name16473 (
		_w20468_,
		_w20519_,
		_w20520_
	);
	LUT2 #(
		.INIT('h1)
	) name16474 (
		_w20516_,
		_w20520_,
		_w20521_
	);
	LUT2 #(
		.INIT('h2)
	) name16475 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[3]/P0001 ,
		_w20468_,
		_w20522_
	);
	LUT2 #(
		.INIT('h1)
	) name16476 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w20523_
	);
	LUT2 #(
		.INIT('h8)
	) name16477 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w20523_,
		_w20524_
	);
	LUT2 #(
		.INIT('h2)
	) name16478 (
		_w20475_,
		_w20524_,
		_w20525_
	);
	LUT2 #(
		.INIT('h8)
	) name16479 (
		_w20473_,
		_w20524_,
		_w20526_
	);
	LUT2 #(
		.INIT('h1)
	) name16480 (
		_w20478_,
		_w20525_,
		_w20527_
	);
	LUT2 #(
		.INIT('h4)
	) name16481 (
		_w20526_,
		_w20527_,
		_w20528_
	);
	LUT2 #(
		.INIT('h2)
	) name16482 (
		_w20468_,
		_w20528_,
		_w20529_
	);
	LUT2 #(
		.INIT('h1)
	) name16483 (
		_w20522_,
		_w20529_,
		_w20530_
	);
	LUT2 #(
		.INIT('h2)
	) name16484 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[2]/P0001 ,
		_w20468_,
		_w20531_
	);
	LUT2 #(
		.INIT('h8)
	) name16485 (
		_w20484_,
		_w20524_,
		_w20532_
	);
	LUT2 #(
		.INIT('h1)
	) name16486 (
		_w20487_,
		_w20525_,
		_w20533_
	);
	LUT2 #(
		.INIT('h4)
	) name16487 (
		_w20532_,
		_w20533_,
		_w20534_
	);
	LUT2 #(
		.INIT('h2)
	) name16488 (
		_w20468_,
		_w20534_,
		_w20535_
	);
	LUT2 #(
		.INIT('h1)
	) name16489 (
		_w20531_,
		_w20535_,
		_w20536_
	);
	LUT2 #(
		.INIT('h2)
	) name16490 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[1]/P0001 ,
		_w20468_,
		_w20537_
	);
	LUT2 #(
		.INIT('h4)
	) name16491 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w20508_,
		_w20538_
	);
	LUT2 #(
		.INIT('h2)
	) name16492 (
		_w20475_,
		_w20538_,
		_w20539_
	);
	LUT2 #(
		.INIT('h8)
	) name16493 (
		_w20473_,
		_w20538_,
		_w20540_
	);
	LUT2 #(
		.INIT('h1)
	) name16494 (
		_w20478_,
		_w20539_,
		_w20541_
	);
	LUT2 #(
		.INIT('h4)
	) name16495 (
		_w20540_,
		_w20541_,
		_w20542_
	);
	LUT2 #(
		.INIT('h2)
	) name16496 (
		_w20468_,
		_w20542_,
		_w20543_
	);
	LUT2 #(
		.INIT('h1)
	) name16497 (
		_w20537_,
		_w20543_,
		_w20544_
	);
	LUT2 #(
		.INIT('h2)
	) name16498 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[11]/P0001 ,
		_w20468_,
		_w20545_
	);
	LUT2 #(
		.INIT('h8)
	) name16499 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w20470_,
		_w20546_
	);
	LUT2 #(
		.INIT('h2)
	) name16500 (
		_w20475_,
		_w20546_,
		_w20547_
	);
	LUT2 #(
		.INIT('h8)
	) name16501 (
		_w20473_,
		_w20546_,
		_w20548_
	);
	LUT2 #(
		.INIT('h1)
	) name16502 (
		_w20478_,
		_w20547_,
		_w20549_
	);
	LUT2 #(
		.INIT('h4)
	) name16503 (
		_w20548_,
		_w20549_,
		_w20550_
	);
	LUT2 #(
		.INIT('h2)
	) name16504 (
		_w20468_,
		_w20550_,
		_w20551_
	);
	LUT2 #(
		.INIT('h1)
	) name16505 (
		_w20545_,
		_w20551_,
		_w20552_
	);
	LUT2 #(
		.INIT('h2)
	) name16506 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[10]/P0001 ,
		_w20468_,
		_w20553_
	);
	LUT2 #(
		.INIT('h8)
	) name16507 (
		_w20484_,
		_w20546_,
		_w20554_
	);
	LUT2 #(
		.INIT('h1)
	) name16508 (
		_w20487_,
		_w20547_,
		_w20555_
	);
	LUT2 #(
		.INIT('h4)
	) name16509 (
		_w20554_,
		_w20555_,
		_w20556_
	);
	LUT2 #(
		.INIT('h2)
	) name16510 (
		_w20468_,
		_w20556_,
		_w20557_
	);
	LUT2 #(
		.INIT('h1)
	) name16511 (
		_w20553_,
		_w20557_,
		_w20558_
	);
	LUT2 #(
		.INIT('h2)
	) name16512 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[0]/P0001 ,
		_w20468_,
		_w20559_
	);
	LUT2 #(
		.INIT('h8)
	) name16513 (
		_w20484_,
		_w20538_,
		_w20560_
	);
	LUT2 #(
		.INIT('h1)
	) name16514 (
		_w20487_,
		_w20539_,
		_w20561_
	);
	LUT2 #(
		.INIT('h4)
	) name16515 (
		_w20560_,
		_w20561_,
		_w20562_
	);
	LUT2 #(
		.INIT('h2)
	) name16516 (
		_w20468_,
		_w20562_,
		_w20563_
	);
	LUT2 #(
		.INIT('h1)
	) name16517 (
		_w20559_,
		_w20563_,
		_w20564_
	);
	LUT2 #(
		.INIT('h4)
	) name16518 (
		_w8460_,
		_w20402_,
		_w20565_
	);
	LUT2 #(
		.INIT('h1)
	) name16519 (
		\sport0_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w20402_,
		_w20566_
	);
	LUT2 #(
		.INIT('h1)
	) name16520 (
		_w20565_,
		_w20566_,
		_w20567_
	);
	LUT2 #(
		.INIT('h4)
	) name16521 (
		_w7859_,
		_w20402_,
		_w20568_
	);
	LUT2 #(
		.INIT('h1)
	) name16522 (
		\sport0_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w20402_,
		_w20569_
	);
	LUT2 #(
		.INIT('h1)
	) name16523 (
		_w20568_,
		_w20569_,
		_w20570_
	);
	LUT2 #(
		.INIT('h1)
	) name16524 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\core_c_dec_MpopLP_Eg_reg/P0001 ,
		_w20571_
	);
	LUT2 #(
		.INIT('h4)
	) name16525 (
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		_w20571_,
		_w20572_
	);
	LUT2 #(
		.INIT('h4)
	) name16526 (
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w4849_,
		_w20573_
	);
	LUT2 #(
		.INIT('h2)
	) name16527 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		_w5950_,
		_w20574_
	);
	LUT2 #(
		.INIT('h4)
	) name16528 (
		_w20573_,
		_w20574_,
		_w20575_
	);
	LUT2 #(
		.INIT('h4)
	) name16529 (
		_w20572_,
		_w20575_,
		_w20576_
	);
	LUT2 #(
		.INIT('h1)
	) name16530 (
		\core_c_dec_MpopLP_Eg_reg/P0001 ,
		_w4842_,
		_w20577_
	);
	LUT2 #(
		.INIT('h1)
	) name16531 (
		_w5950_,
		_w20577_,
		_w20578_
	);
	LUT2 #(
		.INIT('h4)
	) name16532 (
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w20578_,
		_w20579_
	);
	LUT2 #(
		.INIT('h4)
	) name16533 (
		_w20572_,
		_w20579_,
		_w20580_
	);
	LUT2 #(
		.INIT('h1)
	) name16534 (
		_w20576_,
		_w20580_,
		_w20581_
	);
	LUT2 #(
		.INIT('h1)
	) name16535 (
		_w4847_,
		_w4851_,
		_w20582_
	);
	LUT2 #(
		.INIT('h2)
	) name16536 (
		_w20574_,
		_w20582_,
		_w20583_
	);
	LUT2 #(
		.INIT('h4)
	) name16537 (
		_w20575_,
		_w20582_,
		_w20584_
	);
	LUT2 #(
		.INIT('h1)
	) name16538 (
		_w20583_,
		_w20584_,
		_w20585_
	);
	LUT2 #(
		.INIT('h1)
	) name16539 (
		_w20581_,
		_w20585_,
		_w20586_
	);
	LUT2 #(
		.INIT('h8)
	) name16540 (
		\core_c_psq_lpstk_ptr_reg[1]/NET0131 ,
		_w20581_,
		_w20587_
	);
	LUT2 #(
		.INIT('h1)
	) name16541 (
		_w20586_,
		_w20587_,
		_w20588_
	);
	LUT2 #(
		.INIT('h2)
	) name16542 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		_w20581_,
		_w20589_
	);
	LUT2 #(
		.INIT('h4)
	) name16543 (
		\core_c_psq_lpstk_ptr_reg[0]/NET0131 ,
		_w20581_,
		_w20590_
	);
	LUT2 #(
		.INIT('h1)
	) name16544 (
		_w20589_,
		_w20590_,
		_w20591_
	);
	LUT2 #(
		.INIT('h2)
	) name16545 (
		\core_c_psq_Iact_E_reg[7]/NET0131 ,
		_w19477_,
		_w20592_
	);
	LUT2 #(
		.INIT('h8)
	) name16546 (
		_w19487_,
		_w19489_,
		_w20593_
	);
	LUT2 #(
		.INIT('h1)
	) name16547 (
		_w20592_,
		_w20593_,
		_w20594_
	);
	LUT2 #(
		.INIT('h8)
	) name16548 (
		_w4849_,
		_w20576_,
		_w20595_
	);
	LUT2 #(
		.INIT('h2)
	) name16549 (
		\core_c_psq_lpstk_ptr_reg[2]/NET0131 ,
		_w20595_,
		_w20596_
	);
	LUT2 #(
		.INIT('h2)
	) name16550 (
		_w4845_,
		_w20572_,
		_w20597_
	);
	LUT2 #(
		.INIT('h4)
	) name16551 (
		_w20575_,
		_w20597_,
		_w20598_
	);
	LUT2 #(
		.INIT('h8)
	) name16552 (
		_w20578_,
		_w20598_,
		_w20599_
	);
	LUT2 #(
		.INIT('h1)
	) name16553 (
		_w20596_,
		_w20599_,
		_w20600_
	);
	LUT2 #(
		.INIT('h2)
	) name16554 (
		_w6164_,
		_w10638_,
		_w20601_
	);
	LUT2 #(
		.INIT('h1)
	) name16555 (
		_w13347_,
		_w20601_,
		_w20602_
	);
	LUT2 #(
		.INIT('h4)
	) name16556 (
		_w6047_,
		_w20602_,
		_w20603_
	);
	LUT2 #(
		.INIT('h2)
	) name16557 (
		_w11609_,
		_w20603_,
		_w20604_
	);
	LUT2 #(
		.INIT('h2)
	) name16558 (
		_w6029_,
		_w20604_,
		_w20605_
	);
	LUT2 #(
		.INIT('h2)
	) name16559 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w20606_
	);
	LUT2 #(
		.INIT('h8)
	) name16560 (
		_w6118_,
		_w20606_,
		_w20607_
	);
	LUT2 #(
		.INIT('h8)
	) name16561 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w20607_,
		_w20608_
	);
	LUT2 #(
		.INIT('h1)
	) name16562 (
		_w4094_,
		_w20608_,
		_w20609_
	);
	LUT2 #(
		.INIT('h4)
	) name16563 (
		_w20605_,
		_w20609_,
		_w20610_
	);
	LUT2 #(
		.INIT('h4)
	) name16564 (
		\core_c_psq_Taddr_Eb_reg[8]/P0001 ,
		_w4094_,
		_w20611_
	);
	LUT2 #(
		.INIT('h1)
	) name16565 (
		_w20610_,
		_w20611_,
		_w20612_
	);
	LUT2 #(
		.INIT('h2)
	) name16566 (
		_w6164_,
		_w11265_,
		_w20613_
	);
	LUT2 #(
		.INIT('h1)
	) name16567 (
		_w13328_,
		_w20613_,
		_w20614_
	);
	LUT2 #(
		.INIT('h4)
	) name16568 (
		_w6047_,
		_w20614_,
		_w20615_
	);
	LUT2 #(
		.INIT('h2)
	) name16569 (
		_w11540_,
		_w20615_,
		_w20616_
	);
	LUT2 #(
		.INIT('h2)
	) name16570 (
		_w6029_,
		_w20616_,
		_w20617_
	);
	LUT2 #(
		.INIT('h8)
	) name16571 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w20607_,
		_w20618_
	);
	LUT2 #(
		.INIT('h1)
	) name16572 (
		_w4094_,
		_w20618_,
		_w20619_
	);
	LUT2 #(
		.INIT('h4)
	) name16573 (
		_w20617_,
		_w20619_,
		_w20620_
	);
	LUT2 #(
		.INIT('h4)
	) name16574 (
		\core_c_psq_Taddr_Eb_reg[7]/P0001 ,
		_w4094_,
		_w20621_
	);
	LUT2 #(
		.INIT('h1)
	) name16575 (
		_w20620_,
		_w20621_,
		_w20622_
	);
	LUT2 #(
		.INIT('h2)
	) name16576 (
		_w6164_,
		_w11525_,
		_w20623_
	);
	LUT2 #(
		.INIT('h1)
	) name16577 (
		_w13309_,
		_w20623_,
		_w20624_
	);
	LUT2 #(
		.INIT('h4)
	) name16578 (
		_w6047_,
		_w20624_,
		_w20625_
	);
	LUT2 #(
		.INIT('h2)
	) name16579 (
		_w10967_,
		_w20625_,
		_w20626_
	);
	LUT2 #(
		.INIT('h2)
	) name16580 (
		_w6029_,
		_w20626_,
		_w20627_
	);
	LUT2 #(
		.INIT('h8)
	) name16581 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w20607_,
		_w20628_
	);
	LUT2 #(
		.INIT('h1)
	) name16582 (
		_w4094_,
		_w20628_,
		_w20629_
	);
	LUT2 #(
		.INIT('h4)
	) name16583 (
		_w20627_,
		_w20629_,
		_w20630_
	);
	LUT2 #(
		.INIT('h4)
	) name16584 (
		\core_c_psq_Taddr_Eb_reg[6]/P0001 ,
		_w4094_,
		_w20631_
	);
	LUT2 #(
		.INIT('h1)
	) name16585 (
		_w20630_,
		_w20631_,
		_w20632_
	);
	LUT2 #(
		.INIT('h2)
	) name16586 (
		_w6164_,
		_w10911_,
		_w20633_
	);
	LUT2 #(
		.INIT('h1)
	) name16587 (
		_w13290_,
		_w20633_,
		_w20634_
	);
	LUT2 #(
		.INIT('h4)
	) name16588 (
		_w6047_,
		_w20634_,
		_w20635_
	);
	LUT2 #(
		.INIT('h2)
	) name16589 (
		_w10356_,
		_w20635_,
		_w20636_
	);
	LUT2 #(
		.INIT('h2)
	) name16590 (
		_w6029_,
		_w20636_,
		_w20637_
	);
	LUT2 #(
		.INIT('h8)
	) name16591 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w20607_,
		_w20638_
	);
	LUT2 #(
		.INIT('h1)
	) name16592 (
		_w4094_,
		_w20638_,
		_w20639_
	);
	LUT2 #(
		.INIT('h4)
	) name16593 (
		_w20637_,
		_w20639_,
		_w20640_
	);
	LUT2 #(
		.INIT('h4)
	) name16594 (
		\core_c_psq_Taddr_Eb_reg[5]/P0001 ,
		_w4094_,
		_w20641_
	);
	LUT2 #(
		.INIT('h1)
	) name16595 (
		_w20640_,
		_w20641_,
		_w20642_
	);
	LUT2 #(
		.INIT('h2)
	) name16596 (
		_w6164_,
		_w10069_,
		_w20643_
	);
	LUT2 #(
		.INIT('h1)
	) name16597 (
		_w13271_,
		_w20643_,
		_w20644_
	);
	LUT2 #(
		.INIT('h4)
	) name16598 (
		_w6047_,
		_w20644_,
		_w20645_
	);
	LUT2 #(
		.INIT('h2)
	) name16599 (
		_w9805_,
		_w20645_,
		_w20646_
	);
	LUT2 #(
		.INIT('h2)
	) name16600 (
		_w6029_,
		_w20646_,
		_w20647_
	);
	LUT2 #(
		.INIT('h8)
	) name16601 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w20607_,
		_w20648_
	);
	LUT2 #(
		.INIT('h1)
	) name16602 (
		_w4094_,
		_w20648_,
		_w20649_
	);
	LUT2 #(
		.INIT('h4)
	) name16603 (
		_w20647_,
		_w20649_,
		_w20650_
	);
	LUT2 #(
		.INIT('h4)
	) name16604 (
		\core_c_psq_Taddr_Eb_reg[4]/P0001 ,
		_w4094_,
		_w20651_
	);
	LUT2 #(
		.INIT('h1)
	) name16605 (
		_w20650_,
		_w20651_,
		_w20652_
	);
	LUT2 #(
		.INIT('h4)
	) name16606 (
		_w6047_,
		_w13262_,
		_w20653_
	);
	LUT2 #(
		.INIT('h2)
	) name16607 (
		_w9666_,
		_w20653_,
		_w20654_
	);
	LUT2 #(
		.INIT('h2)
	) name16608 (
		_w6029_,
		_w20654_,
		_w20655_
	);
	LUT2 #(
		.INIT('h8)
	) name16609 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w20607_,
		_w20656_
	);
	LUT2 #(
		.INIT('h1)
	) name16610 (
		_w4094_,
		_w20656_,
		_w20657_
	);
	LUT2 #(
		.INIT('h4)
	) name16611 (
		_w20655_,
		_w20657_,
		_w20658_
	);
	LUT2 #(
		.INIT('h4)
	) name16612 (
		\core_c_psq_Taddr_Eb_reg[3]/P0001 ,
		_w4094_,
		_w20659_
	);
	LUT2 #(
		.INIT('h1)
	) name16613 (
		_w20658_,
		_w20659_,
		_w20660_
	);
	LUT2 #(
		.INIT('h1)
	) name16614 (
		_w6164_,
		_w9625_,
		_w20661_
	);
	LUT2 #(
		.INIT('h8)
	) name16615 (
		_w6164_,
		_w8715_,
		_w20662_
	);
	LUT2 #(
		.INIT('h1)
	) name16616 (
		_w20661_,
		_w20662_,
		_w20663_
	);
	LUT2 #(
		.INIT('h1)
	) name16617 (
		_w6047_,
		_w20663_,
		_w20664_
	);
	LUT2 #(
		.INIT('h2)
	) name16618 (
		_w9600_,
		_w20664_,
		_w20665_
	);
	LUT2 #(
		.INIT('h2)
	) name16619 (
		_w6029_,
		_w20665_,
		_w20666_
	);
	LUT2 #(
		.INIT('h8)
	) name16620 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w20607_,
		_w20667_
	);
	LUT2 #(
		.INIT('h1)
	) name16621 (
		_w4094_,
		_w20667_,
		_w20668_
	);
	LUT2 #(
		.INIT('h4)
	) name16622 (
		_w20666_,
		_w20668_,
		_w20669_
	);
	LUT2 #(
		.INIT('h4)
	) name16623 (
		\core_c_psq_Taddr_Eb_reg[2]/P0001 ,
		_w4094_,
		_w20670_
	);
	LUT2 #(
		.INIT('h1)
	) name16624 (
		_w20669_,
		_w20670_,
		_w20671_
	);
	LUT2 #(
		.INIT('h1)
	) name16625 (
		_w6164_,
		_w9559_,
		_w20672_
	);
	LUT2 #(
		.INIT('h8)
	) name16626 (
		_w6164_,
		_w9435_,
		_w20673_
	);
	LUT2 #(
		.INIT('h1)
	) name16627 (
		_w20672_,
		_w20673_,
		_w20674_
	);
	LUT2 #(
		.INIT('h1)
	) name16628 (
		_w6047_,
		_w20674_,
		_w20675_
	);
	LUT2 #(
		.INIT('h2)
	) name16629 (
		_w9528_,
		_w20675_,
		_w20676_
	);
	LUT2 #(
		.INIT('h2)
	) name16630 (
		_w6029_,
		_w20676_,
		_w20677_
	);
	LUT2 #(
		.INIT('h8)
	) name16631 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w20607_,
		_w20678_
	);
	LUT2 #(
		.INIT('h1)
	) name16632 (
		_w4094_,
		_w20678_,
		_w20679_
	);
	LUT2 #(
		.INIT('h4)
	) name16633 (
		_w20677_,
		_w20679_,
		_w20680_
	);
	LUT2 #(
		.INIT('h4)
	) name16634 (
		\core_c_psq_Taddr_Eb_reg[1]/P0001 ,
		_w4094_,
		_w20681_
	);
	LUT2 #(
		.INIT('h1)
	) name16635 (
		_w20680_,
		_w20681_,
		_w20682_
	);
	LUT2 #(
		.INIT('h1)
	) name16636 (
		_w6164_,
		_w9497_,
		_w20683_
	);
	LUT2 #(
		.INIT('h8)
	) name16637 (
		_w6164_,
		_w7340_,
		_w20684_
	);
	LUT2 #(
		.INIT('h1)
	) name16638 (
		_w20683_,
		_w20684_,
		_w20685_
	);
	LUT2 #(
		.INIT('h1)
	) name16639 (
		_w6047_,
		_w20685_,
		_w20686_
	);
	LUT2 #(
		.INIT('h2)
	) name16640 (
		_w9452_,
		_w20686_,
		_w20687_
	);
	LUT2 #(
		.INIT('h2)
	) name16641 (
		_w6029_,
		_w20687_,
		_w20688_
	);
	LUT2 #(
		.INIT('h8)
	) name16642 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w20607_,
		_w20689_
	);
	LUT2 #(
		.INIT('h1)
	) name16643 (
		_w4094_,
		_w20689_,
		_w20690_
	);
	LUT2 #(
		.INIT('h4)
	) name16644 (
		_w20688_,
		_w20690_,
		_w20691_
	);
	LUT2 #(
		.INIT('h4)
	) name16645 (
		\core_c_psq_Taddr_Eb_reg[13]/P0001 ,
		_w4094_,
		_w20692_
	);
	LUT2 #(
		.INIT('h1)
	) name16646 (
		_w20691_,
		_w20692_,
		_w20693_
	);
	LUT2 #(
		.INIT('h1)
	) name16647 (
		_w6164_,
		_w8945_,
		_w20694_
	);
	LUT2 #(
		.INIT('h8)
	) name16648 (
		_w6164_,
		_w9178_,
		_w20695_
	);
	LUT2 #(
		.INIT('h1)
	) name16649 (
		_w20694_,
		_w20695_,
		_w20696_
	);
	LUT2 #(
		.INIT('h1)
	) name16650 (
		_w6047_,
		_w20696_,
		_w20697_
	);
	LUT2 #(
		.INIT('h2)
	) name16651 (
		_w8845_,
		_w20697_,
		_w20698_
	);
	LUT2 #(
		.INIT('h2)
	) name16652 (
		_w6029_,
		_w20698_,
		_w20699_
	);
	LUT2 #(
		.INIT('h8)
	) name16653 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w20607_,
		_w20700_
	);
	LUT2 #(
		.INIT('h1)
	) name16654 (
		_w4094_,
		_w20700_,
		_w20701_
	);
	LUT2 #(
		.INIT('h4)
	) name16655 (
		_w20699_,
		_w20701_,
		_w20702_
	);
	LUT2 #(
		.INIT('h4)
	) name16656 (
		\core_c_psq_Taddr_Eb_reg[12]/P0001 ,
		_w4094_,
		_w20703_
	);
	LUT2 #(
		.INIT('h1)
	) name16657 (
		_w20702_,
		_w20703_,
		_w20704_
	);
	LUT2 #(
		.INIT('h1)
	) name16658 (
		_w6164_,
		_w8813_,
		_w20705_
	);
	LUT2 #(
		.INIT('h8)
	) name16659 (
		_w6164_,
		_w8460_,
		_w20706_
	);
	LUT2 #(
		.INIT('h1)
	) name16660 (
		_w20705_,
		_w20706_,
		_w20707_
	);
	LUT2 #(
		.INIT('h1)
	) name16661 (
		_w6047_,
		_w20707_,
		_w20708_
	);
	LUT2 #(
		.INIT('h2)
	) name16662 (
		_w8723_,
		_w20708_,
		_w20709_
	);
	LUT2 #(
		.INIT('h2)
	) name16663 (
		_w6029_,
		_w20709_,
		_w20710_
	);
	LUT2 #(
		.INIT('h8)
	) name16664 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w20607_,
		_w20711_
	);
	LUT2 #(
		.INIT('h1)
	) name16665 (
		_w4094_,
		_w20711_,
		_w20712_
	);
	LUT2 #(
		.INIT('h4)
	) name16666 (
		_w20710_,
		_w20712_,
		_w20713_
	);
	LUT2 #(
		.INIT('h4)
	) name16667 (
		\core_c_psq_Taddr_Eb_reg[11]/P0001 ,
		_w4094_,
		_w20714_
	);
	LUT2 #(
		.INIT('h1)
	) name16668 (
		_w20713_,
		_w20714_,
		_w20715_
	);
	LUT2 #(
		.INIT('h2)
	) name16669 (
		_w6164_,
		_w7859_,
		_w20716_
	);
	LUT2 #(
		.INIT('h4)
	) name16670 (
		_w6164_,
		_w8211_,
		_w20717_
	);
	LUT2 #(
		.INIT('h1)
	) name16671 (
		_w20716_,
		_w20717_,
		_w20718_
	);
	LUT2 #(
		.INIT('h4)
	) name16672 (
		_w6047_,
		_w20718_,
		_w20719_
	);
	LUT2 #(
		.INIT('h2)
	) name16673 (
		_w8121_,
		_w20719_,
		_w20720_
	);
	LUT2 #(
		.INIT('h2)
	) name16674 (
		_w6029_,
		_w20720_,
		_w20721_
	);
	LUT2 #(
		.INIT('h8)
	) name16675 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w20607_,
		_w20722_
	);
	LUT2 #(
		.INIT('h1)
	) name16676 (
		_w4094_,
		_w20722_,
		_w20723_
	);
	LUT2 #(
		.INIT('h4)
	) name16677 (
		_w20721_,
		_w20723_,
		_w20724_
	);
	LUT2 #(
		.INIT('h4)
	) name16678 (
		\core_c_psq_Taddr_Eb_reg[10]/P0001 ,
		_w4094_,
		_w20725_
	);
	LUT2 #(
		.INIT('h1)
	) name16679 (
		_w20724_,
		_w20725_,
		_w20726_
	);
	LUT2 #(
		.INIT('h1)
	) name16680 (
		_w6164_,
		_w6911_,
		_w20727_
	);
	LUT2 #(
		.INIT('h8)
	) name16681 (
		_w6164_,
		_w7607_,
		_w20728_
	);
	LUT2 #(
		.INIT('h1)
	) name16682 (
		_w20727_,
		_w20728_,
		_w20729_
	);
	LUT2 #(
		.INIT('h1)
	) name16683 (
		_w6047_,
		_w20729_,
		_w20730_
	);
	LUT2 #(
		.INIT('h2)
	) name16684 (
		_w6980_,
		_w20730_,
		_w20731_
	);
	LUT2 #(
		.INIT('h2)
	) name16685 (
		_w6029_,
		_w20731_,
		_w20732_
	);
	LUT2 #(
		.INIT('h8)
	) name16686 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w20607_,
		_w20733_
	);
	LUT2 #(
		.INIT('h1)
	) name16687 (
		_w4094_,
		_w20733_,
		_w20734_
	);
	LUT2 #(
		.INIT('h4)
	) name16688 (
		_w20732_,
		_w20734_,
		_w20735_
	);
	LUT2 #(
		.INIT('h4)
	) name16689 (
		\core_c_psq_Taddr_Eb_reg[0]/P0001 ,
		_w4094_,
		_w20736_
	);
	LUT2 #(
		.INIT('h1)
	) name16690 (
		_w20735_,
		_w20736_,
		_w20737_
	);
	LUT2 #(
		.INIT('h8)
	) name16691 (
		\sice_ICYC_reg[8]/NET0131 ,
		_w18863_,
		_w20738_
	);
	LUT2 #(
		.INIT('h8)
	) name16692 (
		\sice_ICYC_reg[9]/NET0131 ,
		_w20738_,
		_w20739_
	);
	LUT2 #(
		.INIT('h8)
	) name16693 (
		\sice_ICYC_reg[10]/NET0131 ,
		_w20739_,
		_w20740_
	);
	LUT2 #(
		.INIT('h8)
	) name16694 (
		\sice_ICYC_reg[11]/NET0131 ,
		_w20740_,
		_w20741_
	);
	LUT2 #(
		.INIT('h8)
	) name16695 (
		\sice_ICYC_reg[12]/NET0131 ,
		_w20741_,
		_w20742_
	);
	LUT2 #(
		.INIT('h8)
	) name16696 (
		\sice_ICYC_reg[13]/NET0131 ,
		_w20742_,
		_w20743_
	);
	LUT2 #(
		.INIT('h8)
	) name16697 (
		\sice_ICYC_reg[14]/NET0131 ,
		_w20743_,
		_w20744_
	);
	LUT2 #(
		.INIT('h8)
	) name16698 (
		\sice_ICYC_reg[15]/NET0131 ,
		_w20744_,
		_w20745_
	);
	LUT2 #(
		.INIT('h8)
	) name16699 (
		\sice_ICYC_reg[16]/NET0131 ,
		_w20745_,
		_w20746_
	);
	LUT2 #(
		.INIT('h8)
	) name16700 (
		\sice_ICYC_reg[17]/NET0131 ,
		_w20746_,
		_w20747_
	);
	LUT2 #(
		.INIT('h8)
	) name16701 (
		\sice_ICYC_reg[18]/NET0131 ,
		_w20747_,
		_w20748_
	);
	LUT2 #(
		.INIT('h8)
	) name16702 (
		\sice_ICYC_reg[19]/NET0131 ,
		_w20748_,
		_w20749_
	);
	LUT2 #(
		.INIT('h8)
	) name16703 (
		\sice_ICYC_reg[20]/NET0131 ,
		_w20749_,
		_w20750_
	);
	LUT2 #(
		.INIT('h1)
	) name16704 (
		\sice_ICYC_reg[21]/NET0131 ,
		_w20750_,
		_w20751_
	);
	LUT2 #(
		.INIT('h8)
	) name16705 (
		\sice_ICYC_reg[21]/NET0131 ,
		_w20750_,
		_w20752_
	);
	LUT2 #(
		.INIT('h1)
	) name16706 (
		_w20751_,
		_w20752_,
		_w20753_
	);
	LUT2 #(
		.INIT('h2)
	) name16707 (
		_w6164_,
		_w10289_,
		_w20754_
	);
	LUT2 #(
		.INIT('h1)
	) name16708 (
		_w13366_,
		_w20754_,
		_w20755_
	);
	LUT2 #(
		.INIT('h4)
	) name16709 (
		_w6047_,
		_w20755_,
		_w20756_
	);
	LUT2 #(
		.INIT('h2)
	) name16710 (
		_w11668_,
		_w20756_,
		_w20757_
	);
	LUT2 #(
		.INIT('h2)
	) name16711 (
		_w6029_,
		_w20757_,
		_w20758_
	);
	LUT2 #(
		.INIT('h8)
	) name16712 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		_w20607_,
		_w20759_
	);
	LUT2 #(
		.INIT('h1)
	) name16713 (
		_w4094_,
		_w20759_,
		_w20760_
	);
	LUT2 #(
		.INIT('h4)
	) name16714 (
		_w20758_,
		_w20760_,
		_w20761_
	);
	LUT2 #(
		.INIT('h4)
	) name16715 (
		\core_c_psq_Taddr_Eb_reg[9]/P0001 ,
		_w4094_,
		_w20762_
	);
	LUT2 #(
		.INIT('h1)
	) name16716 (
		_w20761_,
		_w20762_,
		_w20763_
	);
	LUT2 #(
		.INIT('h8)
	) name16717 (
		_w13762_,
		_w20070_,
		_w20764_
	);
	LUT2 #(
		.INIT('h8)
	) name16718 (
		_w7237_,
		_w20764_,
		_w20765_
	);
	LUT2 #(
		.INIT('h1)
	) name16719 (
		\bdma_BEAD_reg[0]/NET0131 ,
		_w13147_,
		_w20766_
	);
	LUT2 #(
		.INIT('h2)
	) name16720 (
		_w13751_,
		_w20766_,
		_w20767_
	);
	LUT2 #(
		.INIT('h1)
	) name16721 (
		\bdma_BEAD_reg[1]/NET0131 ,
		_w20767_,
		_w20768_
	);
	LUT2 #(
		.INIT('h8)
	) name16722 (
		\bdma_BEAD_reg[1]/NET0131 ,
		_w20767_,
		_w20769_
	);
	LUT2 #(
		.INIT('h1)
	) name16723 (
		_w20765_,
		_w20768_,
		_w20770_
	);
	LUT2 #(
		.INIT('h4)
	) name16724 (
		_w20769_,
		_w20770_,
		_w20771_
	);
	LUT2 #(
		.INIT('h8)
	) name16725 (
		_w9435_,
		_w20765_,
		_w20772_
	);
	LUT2 #(
		.INIT('h1)
	) name16726 (
		_w20771_,
		_w20772_,
		_w20773_
	);
	LUT2 #(
		.INIT('h4)
	) name16727 (
		_w13147_,
		_w13751_,
		_w20774_
	);
	LUT2 #(
		.INIT('h2)
	) name16728 (
		\bdma_BEAD_reg[0]/NET0131 ,
		_w20774_,
		_w20775_
	);
	LUT2 #(
		.INIT('h4)
	) name16729 (
		\bdma_BEAD_reg[0]/NET0131 ,
		_w20774_,
		_w20776_
	);
	LUT2 #(
		.INIT('h1)
	) name16730 (
		_w20775_,
		_w20776_,
		_w20777_
	);
	LUT2 #(
		.INIT('h1)
	) name16731 (
		_w20765_,
		_w20777_,
		_w20778_
	);
	LUT2 #(
		.INIT('h8)
	) name16732 (
		_w7607_,
		_w20765_,
		_w20779_
	);
	LUT2 #(
		.INIT('h1)
	) name16733 (
		_w20778_,
		_w20779_,
		_w20780_
	);
	LUT2 #(
		.INIT('h2)
	) name16734 (
		\clkc_CLKOUT_reg/NET0131 ,
		_w19467_,
		_w20781_
	);
	LUT2 #(
		.INIT('h4)
	) name16735 (
		\clkc_CLKOUT_reg/NET0131 ,
		_w19467_,
		_w20782_
	);
	LUT2 #(
		.INIT('h1)
	) name16736 (
		_w20781_,
		_w20782_,
		_w20783_
	);
	LUT2 #(
		.INIT('h1)
	) name16737 (
		\sice_ICYC_reg[22]/NET0131 ,
		_w20752_,
		_w20784_
	);
	LUT2 #(
		.INIT('h8)
	) name16738 (
		\sice_ICYC_reg[22]/NET0131 ,
		_w20752_,
		_w20785_
	);
	LUT2 #(
		.INIT('h1)
	) name16739 (
		_w20784_,
		_w20785_,
		_w20786_
	);
	LUT2 #(
		.INIT('h8)
	) name16740 (
		_w7513_,
		_w18226_,
		_w20787_
	);
	LUT2 #(
		.INIT('h4)
	) name16741 (
		\memc_MMR_web_reg/NET0131 ,
		_w20787_,
		_w20788_
	);
	LUT2 #(
		.INIT('h4)
	) name16742 (
		_w11265_,
		_w20788_,
		_w20789_
	);
	LUT2 #(
		.INIT('h1)
	) name16743 (
		\tm_tsr_reg_DO_reg[7]/NET0131 ,
		_w20788_,
		_w20790_
	);
	LUT2 #(
		.INIT('h1)
	) name16744 (
		_w20789_,
		_w20790_,
		_w20791_
	);
	LUT2 #(
		.INIT('h4)
	) name16745 (
		_w11525_,
		_w20788_,
		_w20792_
	);
	LUT2 #(
		.INIT('h1)
	) name16746 (
		\tm_tsr_reg_DO_reg[6]/NET0131 ,
		_w20788_,
		_w20793_
	);
	LUT2 #(
		.INIT('h1)
	) name16747 (
		_w20792_,
		_w20793_,
		_w20794_
	);
	LUT2 #(
		.INIT('h4)
	) name16748 (
		_w10911_,
		_w20788_,
		_w20795_
	);
	LUT2 #(
		.INIT('h1)
	) name16749 (
		\tm_tsr_reg_DO_reg[5]/NET0131 ,
		_w20788_,
		_w20796_
	);
	LUT2 #(
		.INIT('h1)
	) name16750 (
		_w20795_,
		_w20796_,
		_w20797_
	);
	LUT2 #(
		.INIT('h4)
	) name16751 (
		_w8113_,
		_w20788_,
		_w20798_
	);
	LUT2 #(
		.INIT('h1)
	) name16752 (
		\tm_tsr_reg_DO_reg[3]/NET0131 ,
		_w20788_,
		_w20799_
	);
	LUT2 #(
		.INIT('h1)
	) name16753 (
		_w20798_,
		_w20799_,
		_w20800_
	);
	LUT2 #(
		.INIT('h4)
	) name16754 (
		_w8715_,
		_w20788_,
		_w20801_
	);
	LUT2 #(
		.INIT('h1)
	) name16755 (
		\tm_tsr_reg_DO_reg[2]/NET0131 ,
		_w20788_,
		_w20802_
	);
	LUT2 #(
		.INIT('h1)
	) name16756 (
		_w20801_,
		_w20802_,
		_w20803_
	);
	LUT2 #(
		.INIT('h4)
	) name16757 (
		_w10069_,
		_w20788_,
		_w20804_
	);
	LUT2 #(
		.INIT('h1)
	) name16758 (
		\tm_tsr_reg_DO_reg[4]/NET0131 ,
		_w20788_,
		_w20805_
	);
	LUT2 #(
		.INIT('h1)
	) name16759 (
		_w20804_,
		_w20805_,
		_w20806_
	);
	LUT2 #(
		.INIT('h4)
	) name16760 (
		_w9435_,
		_w20788_,
		_w20807_
	);
	LUT2 #(
		.INIT('h1)
	) name16761 (
		\tm_tsr_reg_DO_reg[1]/NET0131 ,
		_w20788_,
		_w20808_
	);
	LUT2 #(
		.INIT('h1)
	) name16762 (
		_w20807_,
		_w20808_,
		_w20809_
	);
	LUT2 #(
		.INIT('h4)
	) name16763 (
		_w7607_,
		_w20788_,
		_w20810_
	);
	LUT2 #(
		.INIT('h1)
	) name16764 (
		\tm_tsr_reg_DO_reg[0]/NET0131 ,
		_w20788_,
		_w20811_
	);
	LUT2 #(
		.INIT('h1)
	) name16765 (
		_w20810_,
		_w20811_,
		_w20812_
	);
	LUT2 #(
		.INIT('h4)
	) name16766 (
		_w12743_,
		_w20788_,
		_w20813_
	);
	LUT2 #(
		.INIT('h1)
	) name16767 (
		\tm_tsr_reg_DO_reg[8]/NET0131 ,
		_w20788_,
		_w20814_
	);
	LUT2 #(
		.INIT('h1)
	) name16768 (
		_w20813_,
		_w20814_,
		_w20815_
	);
	LUT2 #(
		.INIT('h4)
	) name16769 (
		\memc_usysr_DO_reg[7]/NET0131 ,
		_w20455_,
		_w20816_
	);
	LUT2 #(
		.INIT('h2)
	) name16770 (
		\idma_WRcnt_reg[0]/NET0131 ,
		_w20456_,
		_w20817_
	);
	LUT2 #(
		.INIT('h1)
	) name16771 (
		_w20455_,
		_w20457_,
		_w20818_
	);
	LUT2 #(
		.INIT('h4)
	) name16772 (
		_w20817_,
		_w20818_,
		_w20819_
	);
	LUT2 #(
		.INIT('h1)
	) name16773 (
		_w20816_,
		_w20819_,
		_w20820_
	);
	LUT2 #(
		.INIT('h4)
	) name16774 (
		\idma_RDCMD_d1_reg/P0001 ,
		\idma_RDCMD_reg/P0001 ,
		_w20821_
	);
	LUT2 #(
		.INIT('h1)
	) name16775 (
		\idma_DCTL_reg[14]/NET0131 ,
		_w20454_,
		_w20822_
	);
	LUT2 #(
		.INIT('h4)
	) name16776 (
		\idma_PM_1st_reg/NET0131 ,
		_w20822_,
		_w20823_
	);
	LUT2 #(
		.INIT('h8)
	) name16777 (
		_w20821_,
		_w20823_,
		_w20824_
	);
	LUT2 #(
		.INIT('h8)
	) name16778 (
		\idma_RDcyc_reg/NET0131 ,
		_w20823_,
		_w20825_
	);
	LUT2 #(
		.INIT('h4)
	) name16779 (
		\idma_RDcnt_reg[0]/NET0131 ,
		_w20825_,
		_w20826_
	);
	LUT2 #(
		.INIT('h2)
	) name16780 (
		\idma_RDcnt_reg[1]/NET0131 ,
		_w20826_,
		_w20827_
	);
	LUT2 #(
		.INIT('h8)
	) name16781 (
		_w20390_,
		_w20825_,
		_w20828_
	);
	LUT2 #(
		.INIT('h1)
	) name16782 (
		_w20824_,
		_w20828_,
		_w20829_
	);
	LUT2 #(
		.INIT('h4)
	) name16783 (
		_w20827_,
		_w20829_,
		_w20830_
	);
	LUT2 #(
		.INIT('h4)
	) name16784 (
		\memc_usysr_DO_reg[5]/NET0131 ,
		_w20824_,
		_w20831_
	);
	LUT2 #(
		.INIT('h1)
	) name16785 (
		_w20830_,
		_w20831_,
		_w20832_
	);
	LUT2 #(
		.INIT('h4)
	) name16786 (
		\memc_usysr_DO_reg[4]/NET0131 ,
		_w20824_,
		_w20833_
	);
	LUT2 #(
		.INIT('h2)
	) name16787 (
		\idma_RDcnt_reg[0]/NET0131 ,
		_w20825_,
		_w20834_
	);
	LUT2 #(
		.INIT('h1)
	) name16788 (
		_w20824_,
		_w20826_,
		_w20835_
	);
	LUT2 #(
		.INIT('h4)
	) name16789 (
		_w20834_,
		_w20835_,
		_w20836_
	);
	LUT2 #(
		.INIT('h1)
	) name16790 (
		_w20833_,
		_w20836_,
		_w20837_
	);
	LUT2 #(
		.INIT('h8)
	) name16791 (
		\core_c_dec_updAR_E_reg/P0001 ,
		_w4118_,
		_w20838_
	);
	LUT2 #(
		.INIT('h8)
	) name16792 (
		_w18850_,
		_w20377_,
		_w20839_
	);
	LUT2 #(
		.INIT('h1)
	) name16793 (
		_w20838_,
		_w20839_,
		_w20840_
	);
	LUT2 #(
		.INIT('h1)
	) name16794 (
		\sice_ICYC_reg[3]/NET0131 ,
		_w18857_,
		_w20841_
	);
	LUT2 #(
		.INIT('h1)
	) name16795 (
		_w18858_,
		_w20841_,
		_w20842_
	);
	LUT2 #(
		.INIT('h1)
	) name16796 (
		\sice_IIRC_reg[3]/NET0131 ,
		_w18866_,
		_w20843_
	);
	LUT2 #(
		.INIT('h1)
	) name16797 (
		_w18867_,
		_w20843_,
		_w20844_
	);
	LUT2 #(
		.INIT('h8)
	) name16798 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[1]/NET0131 ,
		_w20845_
	);
	LUT2 #(
		.INIT('h2)
	) name16799 (
		\clkc_oscntr_reg_DO_reg[2]/NET0131 ,
		_w20845_,
		_w20846_
	);
	LUT2 #(
		.INIT('h8)
	) name16800 (
		\clkc_oscntr_reg_DO_reg[2]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[3]/NET0131 ,
		_w20847_
	);
	LUT2 #(
		.INIT('h1)
	) name16801 (
		\clkc_oscntr_reg_DO_reg[2]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[3]/NET0131 ,
		_w20848_
	);
	LUT2 #(
		.INIT('h1)
	) name16802 (
		_w20847_,
		_w20848_,
		_w20849_
	);
	LUT2 #(
		.INIT('h1)
	) name16803 (
		_w20846_,
		_w20849_,
		_w20850_
	);
	LUT2 #(
		.INIT('h8)
	) name16804 (
		_w20846_,
		_w20849_,
		_w20851_
	);
	LUT2 #(
		.INIT('h1)
	) name16805 (
		_w20850_,
		_w20851_,
		_w20852_
	);
	LUT2 #(
		.INIT('h8)
	) name16806 (
		\sice_IIRC_reg[8]/NET0131 ,
		_w18871_,
		_w20853_
	);
	LUT2 #(
		.INIT('h8)
	) name16807 (
		\sice_IIRC_reg[9]/NET0131 ,
		_w20853_,
		_w20854_
	);
	LUT2 #(
		.INIT('h8)
	) name16808 (
		\sice_IIRC_reg[10]/NET0131 ,
		_w20854_,
		_w20855_
	);
	LUT2 #(
		.INIT('h8)
	) name16809 (
		\sice_IIRC_reg[11]/NET0131 ,
		_w20855_,
		_w20856_
	);
	LUT2 #(
		.INIT('h8)
	) name16810 (
		\sice_IIRC_reg[12]/NET0131 ,
		_w20856_,
		_w20857_
	);
	LUT2 #(
		.INIT('h8)
	) name16811 (
		\sice_IIRC_reg[13]/NET0131 ,
		_w20857_,
		_w20858_
	);
	LUT2 #(
		.INIT('h8)
	) name16812 (
		\sice_IIRC_reg[14]/NET0131 ,
		_w20858_,
		_w20859_
	);
	LUT2 #(
		.INIT('h1)
	) name16813 (
		\sice_IIRC_reg[14]/NET0131 ,
		_w20858_,
		_w20860_
	);
	LUT2 #(
		.INIT('h1)
	) name16814 (
		_w20859_,
		_w20860_,
		_w20861_
	);
	LUT2 #(
		.INIT('h1)
	) name16815 (
		\sice_ICYC_reg[14]/NET0131 ,
		_w20743_,
		_w20862_
	);
	LUT2 #(
		.INIT('h1)
	) name16816 (
		_w20744_,
		_w20862_,
		_w20863_
	);
	LUT2 #(
		.INIT('h8)
	) name16817 (
		\core_c_dec_updMF_E_reg/P0001 ,
		_w14666_,
		_w20864_
	);
	LUT2 #(
		.INIT('h2)
	) name16818 (
		\core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001 ,
		_w20864_,
		_w20865_
	);
	LUT2 #(
		.INIT('h4)
	) name16819 (
		_w19525_,
		_w20864_,
		_w20866_
	);
	LUT2 #(
		.INIT('h1)
	) name16820 (
		_w20865_,
		_w20866_,
		_w20867_
	);
	LUT2 #(
		.INIT('h2)
	) name16821 (
		\sport0_rxctl_a_sync1_reg/P0001 ,
		\sport0_rxctl_a_sync2_reg/P0001 ,
		_w20868_
	);
	LUT2 #(
		.INIT('h8)
	) name16822 (
		\core_c_dec_MTRX0_E_reg/P0001 ,
		_w5951_,
		_w20869_
	);
	LUT2 #(
		.INIT('h1)
	) name16823 (
		_w20868_,
		_w20869_,
		_w20870_
	);
	LUT2 #(
		.INIT('h4)
	) name16824 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w20870_,
		_w20871_
	);
	LUT2 #(
		.INIT('h4)
	) name16825 (
		\sport0_rxctl_RXSHT_reg[5]/P0001 ,
		_w20868_,
		_w20872_
	);
	LUT2 #(
		.INIT('h4)
	) name16826 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w20873_
	);
	LUT2 #(
		.INIT('h8)
	) name16827 (
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w20873_,
		_w20874_
	);
	LUT2 #(
		.INIT('h8)
	) name16828 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w20875_
	);
	LUT2 #(
		.INIT('h2)
	) name16829 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w20876_
	);
	LUT2 #(
		.INIT('h4)
	) name16830 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w20877_
	);
	LUT2 #(
		.INIT('h1)
	) name16831 (
		_w20876_,
		_w20877_,
		_w20878_
	);
	LUT2 #(
		.INIT('h2)
	) name16832 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20878_,
		_w20879_
	);
	LUT2 #(
		.INIT('h1)
	) name16833 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w20879_,
		_w20880_
	);
	LUT2 #(
		.INIT('h8)
	) name16834 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20879_,
		_w20881_
	);
	LUT2 #(
		.INIT('h2)
	) name16835 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w20881_,
		_w20882_
	);
	LUT2 #(
		.INIT('h8)
	) name16836 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20883_
	);
	LUT2 #(
		.INIT('h8)
	) name16837 (
		_w20878_,
		_w20883_,
		_w20884_
	);
	LUT2 #(
		.INIT('h4)
	) name16838 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20885_
	);
	LUT2 #(
		.INIT('h2)
	) name16839 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		_w20886_
	);
	LUT2 #(
		.INIT('h4)
	) name16840 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[1]/P0001 ,
		_w20887_
	);
	LUT2 #(
		.INIT('h1)
	) name16841 (
		_w20886_,
		_w20887_,
		_w20888_
	);
	LUT2 #(
		.INIT('h4)
	) name16842 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20888_,
		_w20889_
	);
	LUT2 #(
		.INIT('h1)
	) name16843 (
		_w20878_,
		_w20885_,
		_w20890_
	);
	LUT2 #(
		.INIT('h4)
	) name16844 (
		_w20889_,
		_w20890_,
		_w20891_
	);
	LUT2 #(
		.INIT('h2)
	) name16845 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20884_,
		_w20892_
	);
	LUT2 #(
		.INIT('h4)
	) name16846 (
		_w20891_,
		_w20892_,
		_w20893_
	);
	LUT2 #(
		.INIT('h2)
	) name16847 (
		_w20882_,
		_w20893_,
		_w20894_
	);
	LUT2 #(
		.INIT('h1)
	) name16848 (
		_w20878_,
		_w20888_,
		_w20895_
	);
	LUT2 #(
		.INIT('h8)
	) name16849 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20895_,
		_w20896_
	);
	LUT2 #(
		.INIT('h1)
	) name16850 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		_w20878_,
		_w20897_
	);
	LUT2 #(
		.INIT('h1)
	) name16851 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20897_,
		_w20898_
	);
	LUT2 #(
		.INIT('h2)
	) name16852 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20896_,
		_w20899_
	);
	LUT2 #(
		.INIT('h4)
	) name16853 (
		_w20898_,
		_w20899_,
		_w20900_
	);
	LUT2 #(
		.INIT('h1)
	) name16854 (
		_w20882_,
		_w20900_,
		_w20901_
	);
	LUT2 #(
		.INIT('h1)
	) name16855 (
		_w20894_,
		_w20901_,
		_w20902_
	);
	LUT2 #(
		.INIT('h2)
	) name16856 (
		_w20880_,
		_w20902_,
		_w20903_
	);
	LUT2 #(
		.INIT('h8)
	) name16857 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20878_,
		_w20904_
	);
	LUT2 #(
		.INIT('h8)
	) name16858 (
		_w20888_,
		_w20904_,
		_w20905_
	);
	LUT2 #(
		.INIT('h2)
	) name16859 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w20878_,
		_w20906_
	);
	LUT2 #(
		.INIT('h8)
	) name16860 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		_w20878_,
		_w20907_
	);
	LUT2 #(
		.INIT('h1)
	) name16861 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20906_,
		_w20908_
	);
	LUT2 #(
		.INIT('h4)
	) name16862 (
		_w20907_,
		_w20908_,
		_w20909_
	);
	LUT2 #(
		.INIT('h1)
	) name16863 (
		_w20905_,
		_w20909_,
		_w20910_
	);
	LUT2 #(
		.INIT('h2)
	) name16864 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20910_,
		_w20911_
	);
	LUT2 #(
		.INIT('h2)
	) name16865 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		_w20912_
	);
	LUT2 #(
		.INIT('h4)
	) name16866 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_rxctl_RX_reg[3]/P0001 ,
		_w20913_
	);
	LUT2 #(
		.INIT('h1)
	) name16867 (
		_w20912_,
		_w20913_,
		_w20914_
	);
	LUT2 #(
		.INIT('h2)
	) name16868 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20914_,
		_w20915_
	);
	LUT2 #(
		.INIT('h2)
	) name16869 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20878_,
		_w20916_
	);
	LUT2 #(
		.INIT('h4)
	) name16870 (
		_w20915_,
		_w20916_,
		_w20917_
	);
	LUT2 #(
		.INIT('h1)
	) name16871 (
		_w20911_,
		_w20917_,
		_w20918_
	);
	LUT2 #(
		.INIT('h2)
	) name16872 (
		_w20882_,
		_w20918_,
		_w20919_
	);
	LUT2 #(
		.INIT('h4)
	) name16873 (
		_w20882_,
		_w20893_,
		_w20920_
	);
	LUT2 #(
		.INIT('h1)
	) name16874 (
		_w20919_,
		_w20920_,
		_w20921_
	);
	LUT2 #(
		.INIT('h8)
	) name16875 (
		_w20903_,
		_w20921_,
		_w20922_
	);
	LUT2 #(
		.INIT('h1)
	) name16876 (
		_w20878_,
		_w20883_,
		_w20923_
	);
	LUT2 #(
		.INIT('h1)
	) name16877 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20923_,
		_w20924_
	);
	LUT2 #(
		.INIT('h2)
	) name16878 (
		_w20878_,
		_w20888_,
		_w20925_
	);
	LUT2 #(
		.INIT('h1)
	) name16879 (
		_w20878_,
		_w20914_,
		_w20926_
	);
	LUT2 #(
		.INIT('h8)
	) name16880 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20926_,
		_w20927_
	);
	LUT2 #(
		.INIT('h1)
	) name16881 (
		_w20925_,
		_w20927_,
		_w20928_
	);
	LUT2 #(
		.INIT('h1)
	) name16882 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20928_,
		_w20929_
	);
	LUT2 #(
		.INIT('h8)
	) name16883 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w20878_,
		_w20930_
	);
	LUT2 #(
		.INIT('h8)
	) name16884 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20930_,
		_w20931_
	);
	LUT2 #(
		.INIT('h1)
	) name16885 (
		_w20924_,
		_w20931_,
		_w20932_
	);
	LUT2 #(
		.INIT('h4)
	) name16886 (
		_w20929_,
		_w20932_,
		_w20933_
	);
	LUT2 #(
		.INIT('h2)
	) name16887 (
		_w20882_,
		_w20933_,
		_w20934_
	);
	LUT2 #(
		.INIT('h4)
	) name16888 (
		_w20882_,
		_w20918_,
		_w20935_
	);
	LUT2 #(
		.INIT('h1)
	) name16889 (
		_w20934_,
		_w20935_,
		_w20936_
	);
	LUT2 #(
		.INIT('h4)
	) name16890 (
		_w20922_,
		_w20936_,
		_w20937_
	);
	LUT2 #(
		.INIT('h1)
	) name16891 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w20881_,
		_w20938_
	);
	LUT2 #(
		.INIT('h2)
	) name16892 (
		_w20879_,
		_w20938_,
		_w20939_
	);
	LUT2 #(
		.INIT('h8)
	) name16893 (
		_w20882_,
		_w20900_,
		_w20940_
	);
	LUT2 #(
		.INIT('h2)
	) name16894 (
		_w20879_,
		_w20883_,
		_w20941_
	);
	LUT2 #(
		.INIT('h4)
	) name16895 (
		_w20882_,
		_w20941_,
		_w20942_
	);
	LUT2 #(
		.INIT('h1)
	) name16896 (
		_w20940_,
		_w20942_,
		_w20943_
	);
	LUT2 #(
		.INIT('h1)
	) name16897 (
		_w20902_,
		_w20939_,
		_w20944_
	);
	LUT2 #(
		.INIT('h8)
	) name16898 (
		_w20943_,
		_w20944_,
		_w20945_
	);
	LUT2 #(
		.INIT('h8)
	) name16899 (
		_w20921_,
		_w20945_,
		_w20946_
	);
	LUT2 #(
		.INIT('h4)
	) name16900 (
		_w20936_,
		_w20946_,
		_w20947_
	);
	LUT2 #(
		.INIT('h4)
	) name16901 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w20947_,
		_w20948_
	);
	LUT2 #(
		.INIT('h1)
	) name16902 (
		_w20937_,
		_w20948_,
		_w20949_
	);
	LUT2 #(
		.INIT('h4)
	) name16903 (
		_w20880_,
		_w20902_,
		_w20950_
	);
	LUT2 #(
		.INIT('h1)
	) name16904 (
		_w20903_,
		_w20950_,
		_w20951_
	);
	LUT2 #(
		.INIT('h8)
	) name16905 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20876_,
		_w20952_
	);
	LUT2 #(
		.INIT('h1)
	) name16906 (
		_w20938_,
		_w20952_,
		_w20953_
	);
	LUT2 #(
		.INIT('h8)
	) name16907 (
		_w20943_,
		_w20953_,
		_w20954_
	);
	LUT2 #(
		.INIT('h8)
	) name16908 (
		_w20951_,
		_w20954_,
		_w20955_
	);
	LUT2 #(
		.INIT('h8)
	) name16909 (
		_w20921_,
		_w20955_,
		_w20956_
	);
	LUT2 #(
		.INIT('h8)
	) name16910 (
		_w20949_,
		_w20956_,
		_w20957_
	);
	LUT2 #(
		.INIT('h1)
	) name16911 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w20957_,
		_w20958_
	);
	LUT2 #(
		.INIT('h1)
	) name16912 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20895_,
		_w20959_
	);
	LUT2 #(
		.INIT('h8)
	) name16913 (
		_w20878_,
		_w20914_,
		_w20960_
	);
	LUT2 #(
		.INIT('h2)
	) name16914 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20960_,
		_w20961_
	);
	LUT2 #(
		.INIT('h4)
	) name16915 (
		_w20959_,
		_w20961_,
		_w20962_
	);
	LUT2 #(
		.INIT('h1)
	) name16916 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20897_,
		_w20963_
	);
	LUT2 #(
		.INIT('h1)
	) name16917 (
		_w20930_,
		_w20963_,
		_w20964_
	);
	LUT2 #(
		.INIT('h1)
	) name16918 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20964_,
		_w20965_
	);
	LUT2 #(
		.INIT('h1)
	) name16919 (
		_w20962_,
		_w20965_,
		_w20966_
	);
	LUT2 #(
		.INIT('h8)
	) name16920 (
		_w20882_,
		_w20966_,
		_w20967_
	);
	LUT2 #(
		.INIT('h4)
	) name16921 (
		_w20882_,
		_w20933_,
		_w20968_
	);
	LUT2 #(
		.INIT('h1)
	) name16922 (
		_w20967_,
		_w20968_,
		_w20969_
	);
	LUT2 #(
		.INIT('h8)
	) name16923 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20952_,
		_w20970_
	);
	LUT2 #(
		.INIT('h1)
	) name16924 (
		_w20969_,
		_w20970_,
		_w20971_
	);
	LUT2 #(
		.INIT('h2)
	) name16925 (
		_w20947_,
		_w20971_,
		_w20972_
	);
	LUT2 #(
		.INIT('h4)
	) name16926 (
		_w20947_,
		_w20971_,
		_w20973_
	);
	LUT2 #(
		.INIT('h1)
	) name16927 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w20973_,
		_w20974_
	);
	LUT2 #(
		.INIT('h4)
	) name16928 (
		_w20972_,
		_w20974_,
		_w20975_
	);
	LUT2 #(
		.INIT('h1)
	) name16929 (
		_w20967_,
		_w20975_,
		_w20976_
	);
	LUT2 #(
		.INIT('h4)
	) name16930 (
		_w20958_,
		_w20976_,
		_w20977_
	);
	LUT2 #(
		.INIT('h2)
	) name16931 (
		_w20958_,
		_w20976_,
		_w20978_
	);
	LUT2 #(
		.INIT('h2)
	) name16932 (
		_w20875_,
		_w20977_,
		_w20979_
	);
	LUT2 #(
		.INIT('h4)
	) name16933 (
		_w20978_,
		_w20979_,
		_w20980_
	);
	LUT2 #(
		.INIT('h4)
	) name16934 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w10911_,
		_w20981_
	);
	LUT2 #(
		.INIT('h1)
	) name16935 (
		_w20868_,
		_w20874_,
		_w20982_
	);
	LUT2 #(
		.INIT('h4)
	) name16936 (
		_w20981_,
		_w20982_,
		_w20983_
	);
	LUT2 #(
		.INIT('h4)
	) name16937 (
		_w20980_,
		_w20983_,
		_w20984_
	);
	LUT2 #(
		.INIT('h1)
	) name16938 (
		_w20871_,
		_w20872_,
		_w20985_
	);
	LUT2 #(
		.INIT('h4)
	) name16939 (
		_w20984_,
		_w20985_,
		_w20986_
	);
	LUT2 #(
		.INIT('h8)
	) name16940 (
		\sport0_rxctl_RX_reg[5]/P0001 ,
		_w20871_,
		_w20987_
	);
	LUT2 #(
		.INIT('h1)
	) name16941 (
		_w20986_,
		_w20987_,
		_w20988_
	);
	LUT2 #(
		.INIT('h1)
	) name16942 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		_w19466_,
		_w20989_
	);
	LUT2 #(
		.INIT('h8)
	) name16943 (
		\core_c_dec_updMF_E_reg/P0001 ,
		_w13804_,
		_w20990_
	);
	LUT2 #(
		.INIT('h2)
	) name16944 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001 ,
		_w20990_,
		_w20991_
	);
	LUT2 #(
		.INIT('h4)
	) name16945 (
		_w19525_,
		_w20990_,
		_w20992_
	);
	LUT2 #(
		.INIT('h1)
	) name16946 (
		_w20991_,
		_w20992_,
		_w20993_
	);
	LUT2 #(
		.INIT('h2)
	) name16947 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w18974_,
		_w20994_
	);
	LUT2 #(
		.INIT('h2)
	) name16948 (
		_w18153_,
		_w18189_,
		_w20995_
	);
	LUT2 #(
		.INIT('h2)
	) name16949 (
		_w17931_,
		_w18912_,
		_w20996_
	);
	LUT2 #(
		.INIT('h4)
	) name16950 (
		_w18175_,
		_w20996_,
		_w20997_
	);
	LUT2 #(
		.INIT('h4)
	) name16951 (
		_w18069_,
		_w19873_,
		_w20998_
	);
	LUT2 #(
		.INIT('h8)
	) name16952 (
		_w20085_,
		_w20998_,
		_w20999_
	);
	LUT2 #(
		.INIT('h8)
	) name16953 (
		_w18147_,
		_w18745_,
		_w21000_
	);
	LUT2 #(
		.INIT('h1)
	) name16954 (
		_w17922_,
		_w18104_,
		_w21001_
	);
	LUT2 #(
		.INIT('h2)
	) name16955 (
		_w17930_,
		_w18907_,
		_w21002_
	);
	LUT2 #(
		.INIT('h4)
	) name16956 (
		_w18091_,
		_w18125_,
		_w21003_
	);
	LUT2 #(
		.INIT('h4)
	) name16957 (
		_w18912_,
		_w19720_,
		_w21004_
	);
	LUT2 #(
		.INIT('h8)
	) name16958 (
		_w18139_,
		_w18171_,
		_w21005_
	);
	LUT2 #(
		.INIT('h8)
	) name16959 (
		_w18043_,
		_w18162_,
		_w21006_
	);
	LUT2 #(
		.INIT('h8)
	) name16960 (
		_w18046_,
		_w18187_,
		_w21007_
	);
	LUT2 #(
		.INIT('h4)
	) name16961 (
		_w17933_,
		_w20104_,
		_w21008_
	);
	LUT2 #(
		.INIT('h2)
	) name16962 (
		_w18758_,
		_w18775_,
		_w21009_
	);
	LUT2 #(
		.INIT('h8)
	) name16963 (
		_w17945_,
		_w17960_,
		_w21010_
	);
	LUT2 #(
		.INIT('h2)
	) name16964 (
		_w18115_,
		_w18781_,
		_w21011_
	);
	LUT2 #(
		.INIT('h8)
	) name16965 (
		_w18055_,
		_w18172_,
		_w21012_
	);
	LUT2 #(
		.INIT('h8)
	) name16966 (
		_w18070_,
		_w18183_,
		_w21013_
	);
	LUT2 #(
		.INIT('h4)
	) name16967 (
		_w18127_,
		_w18732_,
		_w21014_
	);
	LUT2 #(
		.INIT('h8)
	) name16968 (
		_w18089_,
		_w18128_,
		_w21015_
	);
	LUT2 #(
		.INIT('h8)
	) name16969 (
		_w18056_,
		_w18112_,
		_w21016_
	);
	LUT2 #(
		.INIT('h8)
	) name16970 (
		_w18111_,
		_w18893_,
		_w21017_
	);
	LUT2 #(
		.INIT('h2)
	) name16971 (
		_w17986_,
		_w18167_,
		_w21018_
	);
	LUT2 #(
		.INIT('h2)
	) name16972 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9280_,
		_w21019_
	);
	LUT2 #(
		.INIT('h1)
	) name16973 (
		_w18192_,
		_w21019_,
		_w21020_
	);
	LUT2 #(
		.INIT('h1)
	) name16974 (
		_w20995_,
		_w21012_,
		_w21021_
	);
	LUT2 #(
		.INIT('h1)
	) name16975 (
		_w21015_,
		_w21016_,
		_w21022_
	);
	LUT2 #(
		.INIT('h4)
	) name16976 (
		_w21018_,
		_w21022_,
		_w21023_
	);
	LUT2 #(
		.INIT('h8)
	) name16977 (
		_w21020_,
		_w21021_,
		_w21024_
	);
	LUT2 #(
		.INIT('h4)
	) name16978 (
		_w18040_,
		_w21024_,
		_w21025_
	);
	LUT2 #(
		.INIT('h4)
	) name16979 (
		_w21000_,
		_w21023_,
		_w21026_
	);
	LUT2 #(
		.INIT('h1)
	) name16980 (
		_w21001_,
		_w21002_,
		_w21027_
	);
	LUT2 #(
		.INIT('h1)
	) name16981 (
		_w21003_,
		_w21004_,
		_w21028_
	);
	LUT2 #(
		.INIT('h1)
	) name16982 (
		_w21005_,
		_w21006_,
		_w21029_
	);
	LUT2 #(
		.INIT('h1)
	) name16983 (
		_w21007_,
		_w21010_,
		_w21030_
	);
	LUT2 #(
		.INIT('h1)
	) name16984 (
		_w21013_,
		_w21014_,
		_w21031_
	);
	LUT2 #(
		.INIT('h4)
	) name16985 (
		_w21017_,
		_w21031_,
		_w21032_
	);
	LUT2 #(
		.INIT('h8)
	) name16986 (
		_w21029_,
		_w21030_,
		_w21033_
	);
	LUT2 #(
		.INIT('h8)
	) name16987 (
		_w21027_,
		_w21028_,
		_w21034_
	);
	LUT2 #(
		.INIT('h8)
	) name16988 (
		_w21025_,
		_w21026_,
		_w21035_
	);
	LUT2 #(
		.INIT('h2)
	) name16989 (
		_w20108_,
		_w20997_,
		_w21036_
	);
	LUT2 #(
		.INIT('h1)
	) name16990 (
		_w21008_,
		_w21009_,
		_w21037_
	);
	LUT2 #(
		.INIT('h4)
	) name16991 (
		_w21011_,
		_w21037_,
		_w21038_
	);
	LUT2 #(
		.INIT('h8)
	) name16992 (
		_w21035_,
		_w21036_,
		_w21039_
	);
	LUT2 #(
		.INIT('h8)
	) name16993 (
		_w21033_,
		_w21034_,
		_w21040_
	);
	LUT2 #(
		.INIT('h8)
	) name16994 (
		_w20999_,
		_w21032_,
		_w21041_
	);
	LUT2 #(
		.INIT('h8)
	) name16995 (
		_w21040_,
		_w21041_,
		_w21042_
	);
	LUT2 #(
		.INIT('h8)
	) name16996 (
		_w21038_,
		_w21039_,
		_w21043_
	);
	LUT2 #(
		.INIT('h8)
	) name16997 (
		_w21042_,
		_w21043_,
		_w21044_
	);
	LUT2 #(
		.INIT('h8)
	) name16998 (
		_w20090_,
		_w21044_,
		_w21045_
	);
	LUT2 #(
		.INIT('h8)
	) name16999 (
		_w19793_,
		_w21045_,
		_w21046_
	);
	LUT2 #(
		.INIT('h4)
	) name17000 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w21046_,
		_w21047_
	);
	LUT2 #(
		.INIT('h1)
	) name17001 (
		_w20994_,
		_w21047_,
		_w21048_
	);
	LUT2 #(
		.INIT('h2)
	) name17002 (
		_w18717_,
		_w21048_,
		_w21049_
	);
	LUT2 #(
		.INIT('h1)
	) name17003 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[1]/P0001 ,
		_w18717_,
		_w21050_
	);
	LUT2 #(
		.INIT('h1)
	) name17004 (
		_w21049_,
		_w21050_,
		_w21051_
	);
	LUT2 #(
		.INIT('h1)
	) name17005 (
		\clkc_OUTcnt_reg[5]/NET0131 ,
		_w19471_,
		_w21052_
	);
	LUT2 #(
		.INIT('h1)
	) name17006 (
		_w19472_,
		_w21052_,
		_w21053_
	);
	LUT2 #(
		.INIT('h4)
	) name17007 (
		_w19467_,
		_w21053_,
		_w21054_
	);
	LUT2 #(
		.INIT('h2)
	) name17008 (
		_w17833_,
		_w21048_,
		_w21055_
	);
	LUT2 #(
		.INIT('h1)
	) name17009 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[1]/P0001 ,
		_w17833_,
		_w21056_
	);
	LUT2 #(
		.INIT('h1)
	) name17010 (
		_w21055_,
		_w21056_,
		_w21057_
	);
	LUT2 #(
		.INIT('h1)
	) name17011 (
		\clkc_OUTcnt_reg[2]/NET0131 ,
		_w19468_,
		_w21058_
	);
	LUT2 #(
		.INIT('h1)
	) name17012 (
		_w19469_,
		_w21058_,
		_w21059_
	);
	LUT2 #(
		.INIT('h4)
	) name17013 (
		_w19467_,
		_w21059_,
		_w21060_
	);
	LUT2 #(
		.INIT('h2)
	) name17014 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 ,
		_w18266_,
		_w21061_
	);
	LUT2 #(
		.INIT('h1)
	) name17015 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[5]/P0001 ,
		_w18271_,
		_w21062_
	);
	LUT2 #(
		.INIT('h2)
	) name17016 (
		_w18271_,
		_w20259_,
		_w21063_
	);
	LUT2 #(
		.INIT('h2)
	) name17017 (
		_w18273_,
		_w21062_,
		_w21064_
	);
	LUT2 #(
		.INIT('h4)
	) name17018 (
		_w21063_,
		_w21064_,
		_w21065_
	);
	LUT2 #(
		.INIT('h1)
	) name17019 (
		_w18270_,
		_w21061_,
		_w21066_
	);
	LUT2 #(
		.INIT('h4)
	) name17020 (
		_w21065_,
		_w21066_,
		_w21067_
	);
	LUT2 #(
		.INIT('h1)
	) name17021 (
		_w18262_,
		_w21067_,
		_w21068_
	);
	LUT2 #(
		.INIT('h2)
	) name17022 (
		_w18262_,
		_w19628_,
		_w21069_
	);
	LUT2 #(
		.INIT('h1)
	) name17023 (
		_w21068_,
		_w21069_,
		_w21070_
	);
	LUT2 #(
		.INIT('h8)
	) name17024 (
		_w14752_,
		_w19628_,
		_w21071_
	);
	LUT2 #(
		.INIT('h8)
	) name17025 (
		_w18328_,
		_w20259_,
		_w21072_
	);
	LUT2 #(
		.INIT('h2)
	) name17026 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[5]/P0001 ,
		_w18330_,
		_w21073_
	);
	LUT2 #(
		.INIT('h2)
	) name17027 (
		_w18334_,
		_w21073_,
		_w21074_
	);
	LUT2 #(
		.INIT('h4)
	) name17028 (
		_w21072_,
		_w21074_,
		_w21075_
	);
	LUT2 #(
		.INIT('h1)
	) name17029 (
		_w21071_,
		_w21075_,
		_w21076_
	);
	LUT2 #(
		.INIT('h2)
	) name17030 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w17814_,
		_w21077_
	);
	LUT2 #(
		.INIT('h8)
	) name17031 (
		_w18171_,
		_w18774_,
		_w21078_
	);
	LUT2 #(
		.INIT('h1)
	) name17032 (
		_w18034_,
		_w18192_,
		_w21079_
	);
	LUT2 #(
		.INIT('h4)
	) name17033 (
		_w18040_,
		_w21079_,
		_w21080_
	);
	LUT2 #(
		.INIT('h8)
	) name17034 (
		_w18145_,
		_w21080_,
		_w21081_
	);
	LUT2 #(
		.INIT('h4)
	) name17035 (
		_w20112_,
		_w21081_,
		_w21082_
	);
	LUT2 #(
		.INIT('h8)
	) name17036 (
		_w19790_,
		_w21082_,
		_w21083_
	);
	LUT2 #(
		.INIT('h8)
	) name17037 (
		_w19793_,
		_w21083_,
		_w21084_
	);
	LUT2 #(
		.INIT('h2)
	) name17038 (
		_w18758_,
		_w19857_,
		_w21085_
	);
	LUT2 #(
		.INIT('h8)
	) name17039 (
		_w18046_,
		_w18183_,
		_w21086_
	);
	LUT2 #(
		.INIT('h1)
	) name17040 (
		_w18091_,
		_w20096_,
		_w21087_
	);
	LUT2 #(
		.INIT('h8)
	) name17041 (
		_w18071_,
		_w18171_,
		_w21088_
	);
	LUT2 #(
		.INIT('h8)
	) name17042 (
		_w17980_,
		_w18111_,
		_w21089_
	);
	LUT2 #(
		.INIT('h1)
	) name17043 (
		_w17922_,
		_w18743_,
		_w21090_
	);
	LUT2 #(
		.INIT('h8)
	) name17044 (
		_w18147_,
		_w18162_,
		_w21091_
	);
	LUT2 #(
		.INIT('h2)
	) name17045 (
		_w18766_,
		_w18907_,
		_w21092_
	);
	LUT2 #(
		.INIT('h8)
	) name17046 (
		_w18056_,
		_w18905_,
		_w21093_
	);
	LUT2 #(
		.INIT('h2)
	) name17047 (
		_w18748_,
		_w18895_,
		_w21094_
	);
	LUT2 #(
		.INIT('h4)
	) name17048 (
		_w18912_,
		_w20308_,
		_w21095_
	);
	LUT2 #(
		.INIT('h2)
	) name17049 (
		_w18187_,
		_w19804_,
		_w21096_
	);
	LUT2 #(
		.INIT('h8)
	) name17050 (
		_w17965_,
		_w18072_,
		_w21097_
	);
	LUT2 #(
		.INIT('h2)
	) name17051 (
		_w18115_,
		_w19818_,
		_w21098_
	);
	LUT2 #(
		.INIT('h4)
	) name17052 (
		_w17924_,
		_w20104_,
		_w21099_
	);
	LUT2 #(
		.INIT('h2)
	) name17053 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w8497_,
		_w21100_
	);
	LUT2 #(
		.INIT('h8)
	) name17054 (
		_w17986_,
		_w18722_,
		_w21101_
	);
	LUT2 #(
		.INIT('h4)
	) name17055 (
		_w18108_,
		_w18752_,
		_w21102_
	);
	LUT2 #(
		.INIT('h4)
	) name17056 (
		_w18182_,
		_w18719_,
		_w21103_
	);
	LUT2 #(
		.INIT('h1)
	) name17057 (
		_w21093_,
		_w21100_,
		_w21104_
	);
	LUT2 #(
		.INIT('h4)
	) name17058 (
		_w21101_,
		_w21104_,
		_w21105_
	);
	LUT2 #(
		.INIT('h1)
	) name17059 (
		_w21078_,
		_w21097_,
		_w21106_
	);
	LUT2 #(
		.INIT('h4)
	) name17060 (
		_w21103_,
		_w21106_,
		_w21107_
	);
	LUT2 #(
		.INIT('h4)
	) name17061 (
		_w21086_,
		_w21105_,
		_w21108_
	);
	LUT2 #(
		.INIT('h1)
	) name17062 (
		_w21087_,
		_w21088_,
		_w21109_
	);
	LUT2 #(
		.INIT('h1)
	) name17063 (
		_w21089_,
		_w21090_,
		_w21110_
	);
	LUT2 #(
		.INIT('h1)
	) name17064 (
		_w21091_,
		_w21092_,
		_w21111_
	);
	LUT2 #(
		.INIT('h1)
	) name17065 (
		_w21095_,
		_w21102_,
		_w21112_
	);
	LUT2 #(
		.INIT('h8)
	) name17066 (
		_w21111_,
		_w21112_,
		_w21113_
	);
	LUT2 #(
		.INIT('h8)
	) name17067 (
		_w21109_,
		_w21110_,
		_w21114_
	);
	LUT2 #(
		.INIT('h8)
	) name17068 (
		_w21107_,
		_w21108_,
		_w21115_
	);
	LUT2 #(
		.INIT('h1)
	) name17069 (
		_w21085_,
		_w21094_,
		_w21116_
	);
	LUT2 #(
		.INIT('h1)
	) name17070 (
		_w21096_,
		_w21098_,
		_w21117_
	);
	LUT2 #(
		.INIT('h4)
	) name17071 (
		_w21099_,
		_w21117_,
		_w21118_
	);
	LUT2 #(
		.INIT('h8)
	) name17072 (
		_w21115_,
		_w21116_,
		_w21119_
	);
	LUT2 #(
		.INIT('h8)
	) name17073 (
		_w21113_,
		_w21114_,
		_w21120_
	);
	LUT2 #(
		.INIT('h8)
	) name17074 (
		_w20999_,
		_w21120_,
		_w21121_
	);
	LUT2 #(
		.INIT('h8)
	) name17075 (
		_w21118_,
		_w21119_,
		_w21122_
	);
	LUT2 #(
		.INIT('h8)
	) name17076 (
		_w21121_,
		_w21122_,
		_w21123_
	);
	LUT2 #(
		.INIT('h8)
	) name17077 (
		_w21084_,
		_w21123_,
		_w21124_
	);
	LUT2 #(
		.INIT('h4)
	) name17078 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w21124_,
		_w21125_
	);
	LUT2 #(
		.INIT('h1)
	) name17079 (
		_w21077_,
		_w21125_,
		_w21126_
	);
	LUT2 #(
		.INIT('h2)
	) name17080 (
		_w18717_,
		_w21126_,
		_w21127_
	);
	LUT2 #(
		.INIT('h1)
	) name17081 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[2]/P0001 ,
		_w18717_,
		_w21128_
	);
	LUT2 #(
		.INIT('h1)
	) name17082 (
		_w21127_,
		_w21128_,
		_w21129_
	);
	LUT2 #(
		.INIT('h2)
	) name17083 (
		_w17833_,
		_w21126_,
		_w21130_
	);
	LUT2 #(
		.INIT('h1)
	) name17084 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[2]/P0001 ,
		_w17833_,
		_w21131_
	);
	LUT2 #(
		.INIT('h1)
	) name17085 (
		_w21130_,
		_w21131_,
		_w21132_
	);
	LUT2 #(
		.INIT('h2)
	) name17086 (
		\core_c_dec_Call_Ed_reg/P0001 ,
		_w4184_,
		_w21133_
	);
	LUT2 #(
		.INIT('h1)
	) name17087 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w21134_
	);
	LUT2 #(
		.INIT('h4)
	) name17088 (
		_w21133_,
		_w21134_,
		_w21135_
	);
	LUT2 #(
		.INIT('h1)
	) name17089 (
		_w5950_,
		_w21135_,
		_w21136_
	);
	LUT2 #(
		.INIT('h1)
	) name17090 (
		_w18217_,
		_w21136_,
		_w21137_
	);
	LUT2 #(
		.INIT('h4)
	) name17091 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w4215_,
		_w21138_
	);
	LUT2 #(
		.INIT('h4)
	) name17092 (
		_w21137_,
		_w21138_,
		_w21139_
	);
	LUT2 #(
		.INIT('h1)
	) name17093 (
		\core_c_psq_SSTAT_reg[1]/NET0131 ,
		_w21139_,
		_w21140_
	);
	LUT2 #(
		.INIT('h2)
	) name17094 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w17814_,
		_w21141_
	);
	LUT2 #(
		.INIT('h2)
	) name17095 (
		_w18187_,
		_w18898_,
		_w21142_
	);
	LUT2 #(
		.INIT('h4)
	) name17096 (
		_w18082_,
		_w18766_,
		_w21143_
	);
	LUT2 #(
		.INIT('h4)
	) name17097 (
		_w18098_,
		_w19785_,
		_w21144_
	);
	LUT2 #(
		.INIT('h1)
	) name17098 (
		_w18110_,
		_w18987_,
		_w21145_
	);
	LUT2 #(
		.INIT('h1)
	) name17099 (
		_w18909_,
		_w19864_,
		_w21146_
	);
	LUT2 #(
		.INIT('h4)
	) name17100 (
		_w17998_,
		_w18162_,
		_w21147_
	);
	LUT2 #(
		.INIT('h1)
	) name17101 (
		_w18079_,
		_w18915_,
		_w21148_
	);
	LUT2 #(
		.INIT('h4)
	) name17102 (
		_w18123_,
		_w19808_,
		_w21149_
	);
	LUT2 #(
		.INIT('h8)
	) name17103 (
		_w17991_,
		_w18748_,
		_w21150_
	);
	LUT2 #(
		.INIT('h2)
	) name17104 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w8493_,
		_w21151_
	);
	LUT2 #(
		.INIT('h2)
	) name17105 (
		_w18752_,
		_w18912_,
		_w21152_
	);
	LUT2 #(
		.INIT('h4)
	) name17106 (
		_w17924_,
		_w18083_,
		_w21153_
	);
	LUT2 #(
		.INIT('h2)
	) name17107 (
		_w18088_,
		_w18983_,
		_w21154_
	);
	LUT2 #(
		.INIT('h2)
	) name17108 (
		_w18745_,
		_w18914_,
		_w21155_
	);
	LUT2 #(
		.INIT('h2)
	) name17109 (
		_w18740_,
		_w18918_,
		_w21156_
	);
	LUT2 #(
		.INIT('h1)
	) name17110 (
		_w21155_,
		_w21156_,
		_w21157_
	);
	LUT2 #(
		.INIT('h4)
	) name17111 (
		_w18026_,
		_w21157_,
		_w21158_
	);
	LUT2 #(
		.INIT('h1)
	) name17112 (
		_w17931_,
		_w21158_,
		_w21159_
	);
	LUT2 #(
		.INIT('h1)
	) name17113 (
		_w21143_,
		_w21151_,
		_w21160_
	);
	LUT2 #(
		.INIT('h1)
	) name17114 (
		_w21146_,
		_w21148_,
		_w21161_
	);
	LUT2 #(
		.INIT('h1)
	) name17115 (
		_w21150_,
		_w21152_,
		_w21162_
	);
	LUT2 #(
		.INIT('h8)
	) name17116 (
		_w21161_,
		_w21162_,
		_w21163_
	);
	LUT2 #(
		.INIT('h8)
	) name17117 (
		_w18019_,
		_w21160_,
		_w21164_
	);
	LUT2 #(
		.INIT('h2)
	) name17118 (
		_w18903_,
		_w21142_,
		_w21165_
	);
	LUT2 #(
		.INIT('h1)
	) name17119 (
		_w21144_,
		_w21147_,
		_w21166_
	);
	LUT2 #(
		.INIT('h1)
	) name17120 (
		_w21149_,
		_w21153_,
		_w21167_
	);
	LUT2 #(
		.INIT('h4)
	) name17121 (
		_w21154_,
		_w21167_,
		_w21168_
	);
	LUT2 #(
		.INIT('h8)
	) name17122 (
		_w21165_,
		_w21166_,
		_w21169_
	);
	LUT2 #(
		.INIT('h8)
	) name17123 (
		_w21163_,
		_w21164_,
		_w21170_
	);
	LUT2 #(
		.INIT('h4)
	) name17124 (
		_w21145_,
		_w21170_,
		_w21171_
	);
	LUT2 #(
		.INIT('h8)
	) name17125 (
		_w21168_,
		_w21169_,
		_w21172_
	);
	LUT2 #(
		.INIT('h4)
	) name17126 (
		_w21159_,
		_w21172_,
		_w21173_
	);
	LUT2 #(
		.INIT('h8)
	) name17127 (
		_w21171_,
		_w21173_,
		_w21174_
	);
	LUT2 #(
		.INIT('h4)
	) name17128 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w21174_,
		_w21175_
	);
	LUT2 #(
		.INIT('h1)
	) name17129 (
		_w21141_,
		_w21175_,
		_w21176_
	);
	LUT2 #(
		.INIT('h2)
	) name17130 (
		_w18886_,
		_w21176_,
		_w21177_
	);
	LUT2 #(
		.INIT('h1)
	) name17131 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[2]/P0001 ,
		_w18886_,
		_w21178_
	);
	LUT2 #(
		.INIT('h1)
	) name17132 (
		_w21177_,
		_w21178_,
		_w21179_
	);
	LUT2 #(
		.INIT('h2)
	) name17133 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w20150_,
		_w21180_
	);
	LUT2 #(
		.INIT('h2)
	) name17134 (
		_w18187_,
		_w19818_,
		_w21181_
	);
	LUT2 #(
		.INIT('h2)
	) name17135 (
		_w18001_,
		_w19864_,
		_w21182_
	);
	LUT2 #(
		.INIT('h2)
	) name17136 (
		_w18758_,
		_w18895_,
		_w21183_
	);
	LUT2 #(
		.INIT('h2)
	) name17137 (
		_w18740_,
		_w19804_,
		_w21184_
	);
	LUT2 #(
		.INIT('h2)
	) name17138 (
		_w18099_,
		_w18149_,
		_w21185_
	);
	LUT2 #(
		.INIT('h2)
	) name17139 (
		_w18905_,
		_w18912_,
		_w21186_
	);
	LUT2 #(
		.INIT('h2)
	) name17140 (
		_w18749_,
		_w18912_,
		_w21187_
	);
	LUT2 #(
		.INIT('h2)
	) name17141 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11846_,
		_w21188_
	);
	LUT2 #(
		.INIT('h8)
	) name17142 (
		_w18046_,
		_w18124_,
		_w21189_
	);
	LUT2 #(
		.INIT('h4)
	) name17143 (
		_w18914_,
		_w20308_,
		_w21190_
	);
	LUT2 #(
		.INIT('h8)
	) name17144 (
		_w18055_,
		_w18722_,
		_w21191_
	);
	LUT2 #(
		.INIT('h4)
	) name17145 (
		_w18091_,
		_w18752_,
		_w21192_
	);
	LUT2 #(
		.INIT('h8)
	) name17146 (
		_w18070_,
		_w18745_,
		_w21193_
	);
	LUT2 #(
		.INIT('h2)
	) name17147 (
		_w18153_,
		_w20096_,
		_w21194_
	);
	LUT2 #(
		.INIT('h8)
	) name17148 (
		_w17952_,
		_w19862_,
		_w21195_
	);
	LUT2 #(
		.INIT('h8)
	) name17149 (
		_w18191_,
		_w18766_,
		_w21196_
	);
	LUT2 #(
		.INIT('h8)
	) name17150 (
		_w17952_,
		_w19863_,
		_w21197_
	);
	LUT2 #(
		.INIT('h8)
	) name17151 (
		_w18039_,
		_w18766_,
		_w21198_
	);
	LUT2 #(
		.INIT('h8)
	) name17152 (
		_w17965_,
		_w18067_,
		_w21199_
	);
	LUT2 #(
		.INIT('h8)
	) name17153 (
		_w18071_,
		_w18162_,
		_w21200_
	);
	LUT2 #(
		.INIT('h2)
	) name17154 (
		_w18183_,
		_w18781_,
		_w21201_
	);
	LUT2 #(
		.INIT('h4)
	) name17155 (
		_w17924_,
		_w19785_,
		_w21202_
	);
	LUT2 #(
		.INIT('h1)
	) name17156 (
		_w21182_,
		_w21188_,
		_w21203_
	);
	LUT2 #(
		.INIT('h1)
	) name17157 (
		_w21191_,
		_w21194_,
		_w21204_
	);
	LUT2 #(
		.INIT('h4)
	) name17158 (
		_w21196_,
		_w21204_,
		_w21205_
	);
	LUT2 #(
		.INIT('h4)
	) name17159 (
		_w19811_,
		_w21203_,
		_w21206_
	);
	LUT2 #(
		.INIT('h1)
	) name17160 (
		_w21195_,
		_w21197_,
		_w21207_
	);
	LUT2 #(
		.INIT('h1)
	) name17161 (
		_w21198_,
		_w21199_,
		_w21208_
	);
	LUT2 #(
		.INIT('h8)
	) name17162 (
		_w21207_,
		_w21208_,
		_w21209_
	);
	LUT2 #(
		.INIT('h8)
	) name17163 (
		_w21205_,
		_w21206_,
		_w21210_
	);
	LUT2 #(
		.INIT('h2)
	) name17164 (
		_w17978_,
		_w21186_,
		_w21211_
	);
	LUT2 #(
		.INIT('h1)
	) name17165 (
		_w21187_,
		_w21189_,
		_w21212_
	);
	LUT2 #(
		.INIT('h1)
	) name17166 (
		_w21190_,
		_w21192_,
		_w21213_
	);
	LUT2 #(
		.INIT('h1)
	) name17167 (
		_w21193_,
		_w21200_,
		_w21214_
	);
	LUT2 #(
		.INIT('h8)
	) name17168 (
		_w21213_,
		_w21214_,
		_w21215_
	);
	LUT2 #(
		.INIT('h8)
	) name17169 (
		_w21211_,
		_w21212_,
		_w21216_
	);
	LUT2 #(
		.INIT('h8)
	) name17170 (
		_w21209_,
		_w21210_,
		_w21217_
	);
	LUT2 #(
		.INIT('h1)
	) name17171 (
		_w21181_,
		_w21183_,
		_w21218_
	);
	LUT2 #(
		.INIT('h1)
	) name17172 (
		_w21184_,
		_w21185_,
		_w21219_
	);
	LUT2 #(
		.INIT('h1)
	) name17173 (
		_w21201_,
		_w21202_,
		_w21220_
	);
	LUT2 #(
		.INIT('h8)
	) name17174 (
		_w21219_,
		_w21220_,
		_w21221_
	);
	LUT2 #(
		.INIT('h8)
	) name17175 (
		_w21217_,
		_w21218_,
		_w21222_
	);
	LUT2 #(
		.INIT('h8)
	) name17176 (
		_w21215_,
		_w21216_,
		_w21223_
	);
	LUT2 #(
		.INIT('h8)
	) name17177 (
		_w21222_,
		_w21223_,
		_w21224_
	);
	LUT2 #(
		.INIT('h8)
	) name17178 (
		_w21221_,
		_w21224_,
		_w21225_
	);
	LUT2 #(
		.INIT('h8)
	) name17179 (
		_w19794_,
		_w21225_,
		_w21226_
	);
	LUT2 #(
		.INIT('h4)
	) name17180 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w21226_,
		_w21227_
	);
	LUT2 #(
		.INIT('h1)
	) name17181 (
		_w21180_,
		_w21227_,
		_w21228_
	);
	LUT2 #(
		.INIT('h2)
	) name17182 (
		_w18886_,
		_w21228_,
		_w21229_
	);
	LUT2 #(
		.INIT('h1)
	) name17183 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[14]/P0001 ,
		_w18886_,
		_w21230_
	);
	LUT2 #(
		.INIT('h1)
	) name17184 (
		_w21229_,
		_w21230_,
		_w21231_
	);
	LUT2 #(
		.INIT('h2)
	) name17185 (
		_w19034_,
		_w21176_,
		_w21232_
	);
	LUT2 #(
		.INIT('h1)
	) name17186 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[2]/P0001 ,
		_w19034_,
		_w21233_
	);
	LUT2 #(
		.INIT('h1)
	) name17187 (
		_w21232_,
		_w21233_,
		_w21234_
	);
	LUT2 #(
		.INIT('h2)
	) name17188 (
		_w19034_,
		_w21228_,
		_w21235_
	);
	LUT2 #(
		.INIT('h1)
	) name17189 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[14]/P0001 ,
		_w19034_,
		_w21236_
	);
	LUT2 #(
		.INIT('h1)
	) name17190 (
		_w21235_,
		_w21236_,
		_w21237_
	);
	LUT2 #(
		.INIT('h8)
	) name17191 (
		\core_c_psq_PCS_reg[14]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w21238_
	);
	LUT2 #(
		.INIT('h8)
	) name17192 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		_w4068_,
		_w21239_
	);
	LUT2 #(
		.INIT('h8)
	) name17193 (
		_w4105_,
		_w21239_,
		_w21240_
	);
	LUT2 #(
		.INIT('h1)
	) name17194 (
		_w21238_,
		_w21240_,
		_w21241_
	);
	LUT2 #(
		.INIT('h8)
	) name17195 (
		_w4094_,
		_w21241_,
		_w21242_
	);
	LUT2 #(
		.INIT('h4)
	) name17196 (
		\core_c_psq_Eqend_D_reg/P0001 ,
		_w21242_,
		_w21243_
	);
	LUT2 #(
		.INIT('h1)
	) name17197 (
		_w5046_,
		_w21242_,
		_w21244_
	);
	LUT2 #(
		.INIT('h2)
	) name17198 (
		_w4116_,
		_w21243_,
		_w21245_
	);
	LUT2 #(
		.INIT('h4)
	) name17199 (
		_w21244_,
		_w21245_,
		_w21246_
	);
	LUT2 #(
		.INIT('h8)
	) name17200 (
		\core_c_dec_MpopLP_Eg_reg/P0001 ,
		_w4117_,
		_w21247_
	);
	LUT2 #(
		.INIT('h8)
	) name17201 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w21248_
	);
	LUT2 #(
		.INIT('h8)
	) name17202 (
		_w6027_,
		_w6116_,
		_w21249_
	);
	LUT2 #(
		.INIT('h8)
	) name17203 (
		_w21248_,
		_w21249_,
		_w21250_
	);
	LUT2 #(
		.INIT('h8)
	) name17204 (
		_w11742_,
		_w21250_,
		_w21251_
	);
	LUT2 #(
		.INIT('h8)
	) name17205 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w21251_,
		_w21252_
	);
	LUT2 #(
		.INIT('h1)
	) name17206 (
		_w21247_,
		_w21252_,
		_w21253_
	);
	LUT2 #(
		.INIT('h2)
	) name17207 (
		_w4116_,
		_w21253_,
		_w21254_
	);
	LUT2 #(
		.INIT('h8)
	) name17208 (
		\core_c_dec_Call_Ed_reg/P0001 ,
		_w4117_,
		_w21255_
	);
	LUT2 #(
		.INIT('h1)
	) name17209 (
		_w6029_,
		_w20607_,
		_w21256_
	);
	LUT2 #(
		.INIT('h2)
	) name17210 (
		_w11742_,
		_w21256_,
		_w21257_
	);
	LUT2 #(
		.INIT('h1)
	) name17211 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w20607_,
		_w21258_
	);
	LUT2 #(
		.INIT('h2)
	) name17212 (
		_w21257_,
		_w21258_,
		_w21259_
	);
	LUT2 #(
		.INIT('h1)
	) name17213 (
		_w21255_,
		_w21259_,
		_w21260_
	);
	LUT2 #(
		.INIT('h2)
	) name17214 (
		_w4116_,
		_w21260_,
		_w21261_
	);
	LUT2 #(
		.INIT('h8)
	) name17215 (
		\core_c_dec_ALUop_E_reg/P0001 ,
		_w4117_,
		_w21262_
	);
	LUT2 #(
		.INIT('h1)
	) name17216 (
		_w20377_,
		_w21262_,
		_w21263_
	);
	LUT2 #(
		.INIT('h2)
	) name17217 (
		_w4116_,
		_w21263_,
		_w21264_
	);
	LUT2 #(
		.INIT('h1)
	) name17218 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w20039_,
		_w21265_
	);
	LUT2 #(
		.INIT('h1)
	) name17219 (
		_w20040_,
		_w21265_,
		_w21266_
	);
	LUT2 #(
		.INIT('h4)
	) name17220 (
		_w13750_,
		_w21266_,
		_w21267_
	);
	LUT2 #(
		.INIT('h8)
	) name17221 (
		_w13762_,
		_w20400_,
		_w21268_
	);
	LUT2 #(
		.INIT('h8)
	) name17222 (
		_w11265_,
		_w21268_,
		_w21269_
	);
	LUT2 #(
		.INIT('h4)
	) name17223 (
		_w10069_,
		_w21268_,
		_w21270_
	);
	LUT2 #(
		.INIT('h1)
	) name17224 (
		_w10911_,
		_w11265_,
		_w21271_
	);
	LUT2 #(
		.INIT('h4)
	) name17225 (
		_w11525_,
		_w21271_,
		_w21272_
	);
	LUT2 #(
		.INIT('h8)
	) name17226 (
		_w21270_,
		_w21272_,
		_w21273_
	);
	LUT2 #(
		.INIT('h2)
	) name17227 (
		\bdma_BCTL_reg[7]/NET0131 ,
		_w21268_,
		_w21274_
	);
	LUT2 #(
		.INIT('h1)
	) name17228 (
		_w21269_,
		_w21274_,
		_w21275_
	);
	LUT2 #(
		.INIT('h4)
	) name17229 (
		_w21273_,
		_w21275_,
		_w21276_
	);
	LUT2 #(
		.INIT('h8)
	) name17230 (
		_w11525_,
		_w21268_,
		_w21277_
	);
	LUT2 #(
		.INIT('h2)
	) name17231 (
		\bdma_BCTL_reg[6]/NET0131 ,
		_w21268_,
		_w21278_
	);
	LUT2 #(
		.INIT('h1)
	) name17232 (
		_w21277_,
		_w21278_,
		_w21279_
	);
	LUT2 #(
		.INIT('h4)
	) name17233 (
		_w21273_,
		_w21279_,
		_w21280_
	);
	LUT2 #(
		.INIT('h8)
	) name17234 (
		_w10911_,
		_w21268_,
		_w21281_
	);
	LUT2 #(
		.INIT('h2)
	) name17235 (
		\bdma_BCTL_reg[5]/NET0131 ,
		_w21268_,
		_w21282_
	);
	LUT2 #(
		.INIT('h1)
	) name17236 (
		_w21281_,
		_w21282_,
		_w21283_
	);
	LUT2 #(
		.INIT('h4)
	) name17237 (
		_w21273_,
		_w21283_,
		_w21284_
	);
	LUT2 #(
		.INIT('h1)
	) name17238 (
		\bdma_BCTL_reg[4]/NET0131 ,
		_w21268_,
		_w21285_
	);
	LUT2 #(
		.INIT('h1)
	) name17239 (
		_w21270_,
		_w21285_,
		_w21286_
	);
	LUT2 #(
		.INIT('h1)
	) name17240 (
		_w21273_,
		_w21286_,
		_w21287_
	);
	LUT2 #(
		.INIT('h1)
	) name17241 (
		\clkc_OUTcnt_reg[0]/NET0131 ,
		\clkc_OUTcnt_reg[1]/NET0131 ,
		_w21288_
	);
	LUT2 #(
		.INIT('h1)
	) name17242 (
		_w19468_,
		_w21288_,
		_w21289_
	);
	LUT2 #(
		.INIT('h4)
	) name17243 (
		_w19467_,
		_w21289_,
		_w21290_
	);
	LUT2 #(
		.INIT('h8)
	) name17244 (
		_w7270_,
		_w13762_,
		_w21291_
	);
	LUT2 #(
		.INIT('h2)
	) name17245 (
		\pio_PIO_RES_OUT_reg[8]/P0001 ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w21292_
	);
	LUT2 #(
		.INIT('h4)
	) name17246 (
		\pio_PIO_RES_OUT_reg[8]/P0001 ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w21293_
	);
	LUT2 #(
		.INIT('h1)
	) name17247 (
		_w21292_,
		_w21293_,
		_w21294_
	);
	LUT2 #(
		.INIT('h4)
	) name17248 (
		\PIO_oe[8]_pad ,
		\pio_pmask_reg_DO_reg[8]/NET0131 ,
		_w21295_
	);
	LUT2 #(
		.INIT('h4)
	) name17249 (
		_w21294_,
		_w21295_,
		_w21296_
	);
	LUT2 #(
		.INIT('h1)
	) name17250 (
		\pio_PINT_reg[8]/NET0131 ,
		_w21296_,
		_w21297_
	);
	LUT2 #(
		.INIT('h4)
	) name17251 (
		_w21291_,
		_w21297_,
		_w21298_
	);
	LUT2 #(
		.INIT('h4)
	) name17252 (
		_w9178_,
		_w21291_,
		_w21299_
	);
	LUT2 #(
		.INIT('h1)
	) name17253 (
		_w21298_,
		_w21299_,
		_w21300_
	);
	LUT2 #(
		.INIT('h1)
	) name17254 (
		\tm_WR_TSR_KEEP_TO_TMCLK_p_reg/NET0131 ,
		\tm_WR_TSR_p_reg/P0001 ,
		_w21301_
	);
	LUT2 #(
		.INIT('h1)
	) name17255 (
		\emc_RWcnt_reg[3]/P0001 ,
		_w20216_,
		_w21302_
	);
	LUT2 #(
		.INIT('h1)
	) name17256 (
		_w20217_,
		_w21302_,
		_w21303_
	);
	LUT2 #(
		.INIT('h8)
	) name17257 (
		_w20212_,
		_w21303_,
		_w21304_
	);
	LUT2 #(
		.INIT('h1)
	) name17258 (
		\emc_RWcnt_reg[2]/P0001 ,
		_w20215_,
		_w21305_
	);
	LUT2 #(
		.INIT('h1)
	) name17259 (
		_w20216_,
		_w21305_,
		_w21306_
	);
	LUT2 #(
		.INIT('h8)
	) name17260 (
		_w20212_,
		_w21306_,
		_w21307_
	);
	LUT2 #(
		.INIT('h1)
	) name17261 (
		\emc_RWcnt_reg[1]/P0001 ,
		_w20214_,
		_w21308_
	);
	LUT2 #(
		.INIT('h1)
	) name17262 (
		_w20215_,
		_w21308_,
		_w21309_
	);
	LUT2 #(
		.INIT('h8)
	) name17263 (
		_w20212_,
		_w21309_,
		_w21310_
	);
	LUT2 #(
		.INIT('h4)
	) name17264 (
		\emc_RWcnt_reg[0]/P0001 ,
		_w20213_,
		_w21311_
	);
	LUT2 #(
		.INIT('h1)
	) name17265 (
		_w20214_,
		_w21311_,
		_w21312_
	);
	LUT2 #(
		.INIT('h8)
	) name17266 (
		_w20212_,
		_w21312_,
		_w21313_
	);
	LUT2 #(
		.INIT('h8)
	) name17267 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w19203_,
		_w21314_
	);
	LUT2 #(
		.INIT('h2)
	) name17268 (
		_w19202_,
		_w21314_,
		_w21315_
	);
	LUT2 #(
		.INIT('h1)
	) name17269 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w18519_,
		_w21316_
	);
	LUT2 #(
		.INIT('h8)
	) name17270 (
		_w10289_,
		_w21316_,
		_w21317_
	);
	LUT2 #(
		.INIT('h4)
	) name17271 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w18519_,
		_w21318_
	);
	LUT2 #(
		.INIT('h8)
	) name17272 (
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w21318_,
		_w21319_
	);
	LUT2 #(
		.INIT('h4)
	) name17273 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w21320_
	);
	LUT2 #(
		.INIT('h1)
	) name17274 (
		_w21319_,
		_w21320_,
		_w21321_
	);
	LUT2 #(
		.INIT('h4)
	) name17275 (
		_w21317_,
		_w21321_,
		_w21322_
	);
	LUT2 #(
		.INIT('h8)
	) name17276 (
		_w10638_,
		_w21316_,
		_w21323_
	);
	LUT2 #(
		.INIT('h8)
	) name17277 (
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w21318_,
		_w21324_
	);
	LUT2 #(
		.INIT('h1)
	) name17278 (
		_w21320_,
		_w21324_,
		_w21325_
	);
	LUT2 #(
		.INIT('h4)
	) name17279 (
		_w21323_,
		_w21325_,
		_w21326_
	);
	LUT2 #(
		.INIT('h8)
	) name17280 (
		_w11265_,
		_w21316_,
		_w21327_
	);
	LUT2 #(
		.INIT('h8)
	) name17281 (
		\sport0_txctl_TX_reg[7]/P0001 ,
		_w21318_,
		_w21328_
	);
	LUT2 #(
		.INIT('h1)
	) name17282 (
		_w21320_,
		_w21328_,
		_w21329_
	);
	LUT2 #(
		.INIT('h4)
	) name17283 (
		_w21327_,
		_w21329_,
		_w21330_
	);
	LUT2 #(
		.INIT('h2)
	) name17284 (
		\pio_PIO_RES_OUT_reg[9]/P0001 ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w21331_
	);
	LUT2 #(
		.INIT('h4)
	) name17285 (
		\pio_PIO_RES_OUT_reg[9]/P0001 ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w21332_
	);
	LUT2 #(
		.INIT('h1)
	) name17286 (
		_w21331_,
		_w21332_,
		_w21333_
	);
	LUT2 #(
		.INIT('h4)
	) name17287 (
		\PIO_oe[9]_pad ,
		\pio_pmask_reg_DO_reg[9]/NET0131 ,
		_w21334_
	);
	LUT2 #(
		.INIT('h4)
	) name17288 (
		_w21333_,
		_w21334_,
		_w21335_
	);
	LUT2 #(
		.INIT('h1)
	) name17289 (
		\pio_PINT_reg[9]/NET0131 ,
		_w21335_,
		_w21336_
	);
	LUT2 #(
		.INIT('h4)
	) name17290 (
		_w21291_,
		_w21336_,
		_w21337_
	);
	LUT2 #(
		.INIT('h4)
	) name17291 (
		_w7340_,
		_w21291_,
		_w21338_
	);
	LUT2 #(
		.INIT('h1)
	) name17292 (
		_w21337_,
		_w21338_,
		_w21339_
	);
	LUT2 #(
		.INIT('h8)
	) name17293 (
		\sport0_txctl_TX_reg[15]/P0001 ,
		_w21318_,
		_w21340_
	);
	LUT2 #(
		.INIT('h8)
	) name17294 (
		_w12743_,
		_w21316_,
		_w21341_
	);
	LUT2 #(
		.INIT('h1)
	) name17295 (
		_w21320_,
		_w21340_,
		_w21342_
	);
	LUT2 #(
		.INIT('h4)
	) name17296 (
		_w21341_,
		_w21342_,
		_w21343_
	);
	LUT2 #(
		.INIT('h8)
	) name17297 (
		_w7340_,
		_w21316_,
		_w21344_
	);
	LUT2 #(
		.INIT('h8)
	) name17298 (
		\sport0_txctl_TX_reg[13]/P0001 ,
		_w21318_,
		_w21345_
	);
	LUT2 #(
		.INIT('h1)
	) name17299 (
		_w21320_,
		_w21345_,
		_w21346_
	);
	LUT2 #(
		.INIT('h4)
	) name17300 (
		_w21344_,
		_w21346_,
		_w21347_
	);
	LUT2 #(
		.INIT('h8)
	) name17301 (
		_w12688_,
		_w21316_,
		_w21348_
	);
	LUT2 #(
		.INIT('h8)
	) name17302 (
		\sport0_txctl_TX_reg[14]/P0001 ,
		_w21318_,
		_w21349_
	);
	LUT2 #(
		.INIT('h1)
	) name17303 (
		_w21320_,
		_w21349_,
		_w21350_
	);
	LUT2 #(
		.INIT('h4)
	) name17304 (
		_w21348_,
		_w21350_,
		_w21351_
	);
	LUT2 #(
		.INIT('h8)
	) name17305 (
		_w9178_,
		_w21316_,
		_w21352_
	);
	LUT2 #(
		.INIT('h8)
	) name17306 (
		\sport0_txctl_TX_reg[12]/P0001 ,
		_w21318_,
		_w21353_
	);
	LUT2 #(
		.INIT('h1)
	) name17307 (
		_w21320_,
		_w21353_,
		_w21354_
	);
	LUT2 #(
		.INIT('h4)
	) name17308 (
		_w21352_,
		_w21354_,
		_w21355_
	);
	LUT2 #(
		.INIT('h8)
	) name17309 (
		_w8460_,
		_w21316_,
		_w21356_
	);
	LUT2 #(
		.INIT('h8)
	) name17310 (
		\sport0_txctl_TX_reg[11]/P0001 ,
		_w21318_,
		_w21357_
	);
	LUT2 #(
		.INIT('h1)
	) name17311 (
		_w21320_,
		_w21357_,
		_w21358_
	);
	LUT2 #(
		.INIT('h4)
	) name17312 (
		_w21356_,
		_w21358_,
		_w21359_
	);
	LUT2 #(
		.INIT('h8)
	) name17313 (
		_w7859_,
		_w21316_,
		_w21360_
	);
	LUT2 #(
		.INIT('h8)
	) name17314 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		_w21318_,
		_w21361_
	);
	LUT2 #(
		.INIT('h1)
	) name17315 (
		_w21320_,
		_w21361_,
		_w21362_
	);
	LUT2 #(
		.INIT('h4)
	) name17316 (
		_w21360_,
		_w21362_,
		_w21363_
	);
	LUT2 #(
		.INIT('h2)
	) name17317 (
		\core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001 ,
		_w20864_,
		_w21364_
	);
	LUT2 #(
		.INIT('h8)
	) name17318 (
		_w19692_,
		_w20864_,
		_w21365_
	);
	LUT2 #(
		.INIT('h1)
	) name17319 (
		_w21364_,
		_w21365_,
		_w21366_
	);
	LUT2 #(
		.INIT('h1)
	) name17320 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w20870_,
		_w21367_
	);
	LUT2 #(
		.INIT('h1)
	) name17321 (
		_w20875_,
		_w21367_,
		_w21368_
	);
	LUT2 #(
		.INIT('h8)
	) name17322 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w21369_
	);
	LUT2 #(
		.INIT('h4)
	) name17323 (
		_w21368_,
		_w21369_,
		_w21370_
	);
	LUT2 #(
		.INIT('h1)
	) name17324 (
		\sport0_rxctl_RSreq_reg/NET0131 ,
		_w21370_,
		_w21371_
	);
	LUT2 #(
		.INIT('h2)
	) name17325 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001 ,
		_w20990_,
		_w21372_
	);
	LUT2 #(
		.INIT('h8)
	) name17326 (
		_w19692_,
		_w20990_,
		_w21373_
	);
	LUT2 #(
		.INIT('h1)
	) name17327 (
		_w21372_,
		_w21373_,
		_w21374_
	);
	LUT2 #(
		.INIT('h4)
	) name17328 (
		\IRFS1_pad ,
		\T_RFS1_pad ,
		_w21375_
	);
	LUT2 #(
		.INIT('h2)
	) name17329 (
		\IRFS1_pad ,
		_w13618_,
		_w21376_
	);
	LUT2 #(
		.INIT('h1)
	) name17330 (
		_w21375_,
		_w21376_,
		_w21377_
	);
	LUT2 #(
		.INIT('h4)
	) name17331 (
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w21377_,
		_w21378_
	);
	LUT2 #(
		.INIT('h2)
	) name17332 (
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w21377_,
		_w21379_
	);
	LUT2 #(
		.INIT('h1)
	) name17333 (
		_w21378_,
		_w21379_,
		_w21380_
	);
	LUT2 #(
		.INIT('h4)
	) name17334 (
		\sport1_cfg_RFSgi_d_reg/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w21381_
	);
	LUT2 #(
		.INIT('h8)
	) name17335 (
		_w21380_,
		_w21381_,
		_w21382_
	);
	LUT2 #(
		.INIT('h4)
	) name17336 (
		\IRFS0_pad ,
		\T_RFS0_pad ,
		_w21383_
	);
	LUT2 #(
		.INIT('h2)
	) name17337 (
		\IRFS0_pad ,
		_w13613_,
		_w21384_
	);
	LUT2 #(
		.INIT('h1)
	) name17338 (
		_w21383_,
		_w21384_,
		_w21385_
	);
	LUT2 #(
		.INIT('h4)
	) name17339 (
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w21385_,
		_w21386_
	);
	LUT2 #(
		.INIT('h2)
	) name17340 (
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w21385_,
		_w21387_
	);
	LUT2 #(
		.INIT('h1)
	) name17341 (
		_w21386_,
		_w21387_,
		_w21388_
	);
	LUT2 #(
		.INIT('h4)
	) name17342 (
		\sport0_cfg_RFSgi_d_reg/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w21389_
	);
	LUT2 #(
		.INIT('h8)
	) name17343 (
		_w21388_,
		_w21389_,
		_w21390_
	);
	LUT2 #(
		.INIT('h2)
	) name17344 (
		\core_c_psq_Iact_E_reg[9]/NET0131 ,
		_w4116_,
		_w21391_
	);
	LUT2 #(
		.INIT('h1)
	) name17345 (
		\core_c_psq_IFC_reg[7]/NET0131 ,
		_w21391_,
		_w21392_
	);
	LUT2 #(
		.INIT('h2)
	) name17346 (
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		_w21392_,
		_w21393_
	);
	LUT2 #(
		.INIT('h8)
	) name17347 (
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		\core_c_psq_T_IRQ2_s1_reg/P0001 ,
		_w21394_
	);
	LUT2 #(
		.INIT('h2)
	) name17348 (
		\core_c_psq_irq2_de_OUT_reg/P0001 ,
		_w21394_,
		_w21395_
	);
	LUT2 #(
		.INIT('h1)
	) name17349 (
		\core_c_psq_IFC_reg[15]/NET0131 ,
		\core_c_psq_Iflag_reg[9]/NET0131 ,
		_w21396_
	);
	LUT2 #(
		.INIT('h2)
	) name17350 (
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		_w21396_,
		_w21397_
	);
	LUT2 #(
		.INIT('h1)
	) name17351 (
		_w21395_,
		_w21397_,
		_w21398_
	);
	LUT2 #(
		.INIT('h1)
	) name17352 (
		_w21393_,
		_w21398_,
		_w21399_
	);
	LUT2 #(
		.INIT('h4)
	) name17353 (
		\core_c_psq_ICNTL_reg_DO_reg[1]/NET0131 ,
		\core_c_psq_irq1_de_OUT_reg/P0001 ,
		_w21400_
	);
	LUT2 #(
		.INIT('h4)
	) name17354 (
		\core_c_psq_T_IRQ1_s1_reg/P0001 ,
		\core_c_psq_irq1_de_OUT_reg/P0001 ,
		_w21401_
	);
	LUT2 #(
		.INIT('h1)
	) name17355 (
		\core_c_psq_IFC_reg[10]/NET0131 ,
		_w21401_,
		_w21402_
	);
	LUT2 #(
		.INIT('h1)
	) name17356 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w21402_,
		_w21403_
	);
	LUT2 #(
		.INIT('h1)
	) name17357 (
		\core_c_psq_Iflag_reg[12]/NET0131 ,
		_w21403_,
		_w21404_
	);
	LUT2 #(
		.INIT('h2)
	) name17358 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		_w4116_,
		_w21405_
	);
	LUT2 #(
		.INIT('h1)
	) name17359 (
		\core_c_psq_IFC_reg[2]/NET0131 ,
		_w21405_,
		_w21406_
	);
	LUT2 #(
		.INIT('h2)
	) name17360 (
		\core_c_psq_ICNTL_reg_DO_reg[1]/NET0131 ,
		_w21404_,
		_w21407_
	);
	LUT2 #(
		.INIT('h8)
	) name17361 (
		_w21406_,
		_w21407_,
		_w21408_
	);
	LUT2 #(
		.INIT('h1)
	) name17362 (
		_w21400_,
		_w21408_,
		_w21409_
	);
	LUT2 #(
		.INIT('h4)
	) name17363 (
		\core_c_psq_ICNTL_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_irq0_de_OUT_reg/P0001 ,
		_w21410_
	);
	LUT2 #(
		.INIT('h4)
	) name17364 (
		\core_c_psq_T_IRQ0_s1_reg/P0001 ,
		\core_c_psq_irq0_de_OUT_reg/P0001 ,
		_w21411_
	);
	LUT2 #(
		.INIT('h1)
	) name17365 (
		\core_c_psq_IFC_reg[9]/NET0131 ,
		_w21411_,
		_w21412_
	);
	LUT2 #(
		.INIT('h1)
	) name17366 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w21412_,
		_w21413_
	);
	LUT2 #(
		.INIT('h1)
	) name17367 (
		\core_c_psq_Iflag_reg[11]/NET0131 ,
		_w21413_,
		_w21414_
	);
	LUT2 #(
		.INIT('h2)
	) name17368 (
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		_w4116_,
		_w21415_
	);
	LUT2 #(
		.INIT('h1)
	) name17369 (
		\core_c_psq_IFC_reg[1]/NET0131 ,
		_w21415_,
		_w21416_
	);
	LUT2 #(
		.INIT('h2)
	) name17370 (
		\core_c_psq_ICNTL_reg_DO_reg[0]/NET0131 ,
		_w21414_,
		_w21417_
	);
	LUT2 #(
		.INIT('h8)
	) name17371 (
		_w21416_,
		_w21417_,
		_w21418_
	);
	LUT2 #(
		.INIT('h1)
	) name17372 (
		_w21410_,
		_w21418_,
		_w21419_
	);
	LUT2 #(
		.INIT('h8)
	) name17373 (
		\core_c_dec_updSR_E_reg/P0001 ,
		_w4118_,
		_w21420_
	);
	LUT2 #(
		.INIT('h2)
	) name17374 (
		_w4116_,
		_w4117_,
		_w21421_
	);
	LUT2 #(
		.INIT('h8)
	) name17375 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w21422_
	);
	LUT2 #(
		.INIT('h1)
	) name17376 (
		_w19530_,
		_w21422_,
		_w21423_
	);
	LUT2 #(
		.INIT('h8)
	) name17377 (
		_w21421_,
		_w21423_,
		_w21424_
	);
	LUT2 #(
		.INIT('h1)
	) name17378 (
		_w21420_,
		_w21424_,
		_w21425_
	);
	LUT2 #(
		.INIT('h8)
	) name17379 (
		\core_c_dec_Nseq_Ed_reg/P0001 ,
		_w4117_,
		_w21426_
	);
	LUT2 #(
		.INIT('h8)
	) name17380 (
		_w6115_,
		_w19698_,
		_w21427_
	);
	LUT2 #(
		.INIT('h4)
	) name17381 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w21427_,
		_w21428_
	);
	LUT2 #(
		.INIT('h8)
	) name17382 (
		_w11742_,
		_w21428_,
		_w21429_
	);
	LUT2 #(
		.INIT('h1)
	) name17383 (
		_w21257_,
		_w21426_,
		_w21430_
	);
	LUT2 #(
		.INIT('h4)
	) name17384 (
		_w21429_,
		_w21430_,
		_w21431_
	);
	LUT2 #(
		.INIT('h2)
	) name17385 (
		_w4116_,
		_w21431_,
		_w21432_
	);
	LUT2 #(
		.INIT('h8)
	) name17386 (
		\core_c_dec_Nrti_Ed_reg/P0001 ,
		_w4117_,
		_w21433_
	);
	LUT2 #(
		.INIT('h4)
	) name17387 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w21429_,
		_w21434_
	);
	LUT2 #(
		.INIT('h1)
	) name17388 (
		_w21257_,
		_w21433_,
		_w21435_
	);
	LUT2 #(
		.INIT('h4)
	) name17389 (
		_w21434_,
		_w21435_,
		_w21436_
	);
	LUT2 #(
		.INIT('h2)
	) name17390 (
		_w4116_,
		_w21436_,
		_w21437_
	);
	LUT2 #(
		.INIT('h2)
	) name17391 (
		\pio_PIO_RES_OUT_reg[5]/P0001 ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w21438_
	);
	LUT2 #(
		.INIT('h4)
	) name17392 (
		\pio_PIO_RES_OUT_reg[5]/P0001 ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w21439_
	);
	LUT2 #(
		.INIT('h1)
	) name17393 (
		_w21438_,
		_w21439_,
		_w21440_
	);
	LUT2 #(
		.INIT('h4)
	) name17394 (
		\PIO_oe[5]_pad ,
		\pio_pmask_reg_DO_reg[5]/NET0131 ,
		_w21441_
	);
	LUT2 #(
		.INIT('h4)
	) name17395 (
		_w21440_,
		_w21441_,
		_w21442_
	);
	LUT2 #(
		.INIT('h1)
	) name17396 (
		\pio_PINT_reg[5]/NET0131 ,
		_w21442_,
		_w21443_
	);
	LUT2 #(
		.INIT('h4)
	) name17397 (
		_w21291_,
		_w21443_,
		_w21444_
	);
	LUT2 #(
		.INIT('h4)
	) name17398 (
		_w10911_,
		_w21291_,
		_w21445_
	);
	LUT2 #(
		.INIT('h1)
	) name17399 (
		_w21444_,
		_w21445_,
		_w21446_
	);
	LUT2 #(
		.INIT('h2)
	) name17400 (
		\pio_PIO_RES_OUT_reg[4]/P0001 ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w21447_
	);
	LUT2 #(
		.INIT('h4)
	) name17401 (
		\pio_PIO_RES_OUT_reg[4]/P0001 ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w21448_
	);
	LUT2 #(
		.INIT('h1)
	) name17402 (
		_w21447_,
		_w21448_,
		_w21449_
	);
	LUT2 #(
		.INIT('h4)
	) name17403 (
		\PIO_oe[4]_pad ,
		\pio_pmask_reg_DO_reg[4]/NET0131 ,
		_w21450_
	);
	LUT2 #(
		.INIT('h4)
	) name17404 (
		_w21449_,
		_w21450_,
		_w21451_
	);
	LUT2 #(
		.INIT('h1)
	) name17405 (
		\pio_PINT_reg[4]/NET0131 ,
		_w21451_,
		_w21452_
	);
	LUT2 #(
		.INIT('h4)
	) name17406 (
		_w21291_,
		_w21452_,
		_w21453_
	);
	LUT2 #(
		.INIT('h4)
	) name17407 (
		_w10069_,
		_w21291_,
		_w21454_
	);
	LUT2 #(
		.INIT('h1)
	) name17408 (
		_w21453_,
		_w21454_,
		_w21455_
	);
	LUT2 #(
		.INIT('h2)
	) name17409 (
		\pio_PIO_RES_OUT_reg[11]/P0001 ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w21456_
	);
	LUT2 #(
		.INIT('h4)
	) name17410 (
		\pio_PIO_RES_OUT_reg[11]/P0001 ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w21457_
	);
	LUT2 #(
		.INIT('h1)
	) name17411 (
		_w21456_,
		_w21457_,
		_w21458_
	);
	LUT2 #(
		.INIT('h4)
	) name17412 (
		\PIO_oe[11]_pad ,
		\pio_pmask_reg_DO_reg[11]/NET0131 ,
		_w21459_
	);
	LUT2 #(
		.INIT('h4)
	) name17413 (
		_w21458_,
		_w21459_,
		_w21460_
	);
	LUT2 #(
		.INIT('h1)
	) name17414 (
		\pio_PINT_reg[11]/NET0131 ,
		_w21460_,
		_w21461_
	);
	LUT2 #(
		.INIT('h4)
	) name17415 (
		_w21291_,
		_w21461_,
		_w21462_
	);
	LUT2 #(
		.INIT('h4)
	) name17416 (
		_w12743_,
		_w21291_,
		_w21463_
	);
	LUT2 #(
		.INIT('h1)
	) name17417 (
		_w21462_,
		_w21463_,
		_w21464_
	);
	LUT2 #(
		.INIT('h2)
	) name17418 (
		\pio_PIO_RES_OUT_reg[2]/P0001 ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w21465_
	);
	LUT2 #(
		.INIT('h4)
	) name17419 (
		\pio_PIO_RES_OUT_reg[2]/P0001 ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w21466_
	);
	LUT2 #(
		.INIT('h1)
	) name17420 (
		_w21465_,
		_w21466_,
		_w21467_
	);
	LUT2 #(
		.INIT('h4)
	) name17421 (
		\PIO_oe[2]_pad ,
		\pio_pmask_reg_DO_reg[2]/NET0131 ,
		_w21468_
	);
	LUT2 #(
		.INIT('h4)
	) name17422 (
		_w21467_,
		_w21468_,
		_w21469_
	);
	LUT2 #(
		.INIT('h1)
	) name17423 (
		\pio_PINT_reg[2]/NET0131 ,
		_w21469_,
		_w21470_
	);
	LUT2 #(
		.INIT('h4)
	) name17424 (
		_w21291_,
		_w21470_,
		_w21471_
	);
	LUT2 #(
		.INIT('h4)
	) name17425 (
		_w8715_,
		_w21291_,
		_w21472_
	);
	LUT2 #(
		.INIT('h1)
	) name17426 (
		_w21471_,
		_w21472_,
		_w21473_
	);
	LUT2 #(
		.INIT('h2)
	) name17427 (
		\pio_PIO_RES_OUT_reg[10]/P0001 ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w21474_
	);
	LUT2 #(
		.INIT('h4)
	) name17428 (
		\pio_PIO_RES_OUT_reg[10]/P0001 ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w21475_
	);
	LUT2 #(
		.INIT('h1)
	) name17429 (
		_w21474_,
		_w21475_,
		_w21476_
	);
	LUT2 #(
		.INIT('h4)
	) name17430 (
		\PIO_oe[10]_pad ,
		\pio_pmask_reg_DO_reg[10]/NET0131 ,
		_w21477_
	);
	LUT2 #(
		.INIT('h4)
	) name17431 (
		_w21476_,
		_w21477_,
		_w21478_
	);
	LUT2 #(
		.INIT('h1)
	) name17432 (
		\pio_PINT_reg[10]/NET0131 ,
		_w21478_,
		_w21479_
	);
	LUT2 #(
		.INIT('h4)
	) name17433 (
		_w21291_,
		_w21479_,
		_w21480_
	);
	LUT2 #(
		.INIT('h4)
	) name17434 (
		_w12688_,
		_w21291_,
		_w21481_
	);
	LUT2 #(
		.INIT('h1)
	) name17435 (
		_w21480_,
		_w21481_,
		_w21482_
	);
	LUT2 #(
		.INIT('h2)
	) name17436 (
		\pio_PIO_RES_OUT_reg[0]/P0001 ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w21483_
	);
	LUT2 #(
		.INIT('h4)
	) name17437 (
		\pio_PIO_RES_OUT_reg[0]/P0001 ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w21484_
	);
	LUT2 #(
		.INIT('h1)
	) name17438 (
		_w21483_,
		_w21484_,
		_w21485_
	);
	LUT2 #(
		.INIT('h4)
	) name17439 (
		\PIO_oe[0]_pad ,
		\pio_pmask_reg_DO_reg[0]/NET0131 ,
		_w21486_
	);
	LUT2 #(
		.INIT('h4)
	) name17440 (
		_w21485_,
		_w21486_,
		_w21487_
	);
	LUT2 #(
		.INIT('h1)
	) name17441 (
		\pio_PINT_reg[0]/NET0131 ,
		_w21487_,
		_w21488_
	);
	LUT2 #(
		.INIT('h4)
	) name17442 (
		_w21291_,
		_w21488_,
		_w21489_
	);
	LUT2 #(
		.INIT('h4)
	) name17443 (
		_w7607_,
		_w21291_,
		_w21490_
	);
	LUT2 #(
		.INIT('h1)
	) name17444 (
		_w21489_,
		_w21490_,
		_w21491_
	);
	LUT2 #(
		.INIT('h2)
	) name17445 (
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		_w19477_,
		_w21492_
	);
	LUT2 #(
		.INIT('h4)
	) name17446 (
		_w19488_,
		_w19491_,
		_w21493_
	);
	LUT2 #(
		.INIT('h4)
	) name17447 (
		_w19493_,
		_w21493_,
		_w21494_
	);
	LUT2 #(
		.INIT('h8)
	) name17448 (
		_w19487_,
		_w21494_,
		_w21495_
	);
	LUT2 #(
		.INIT('h1)
	) name17449 (
		_w21492_,
		_w21495_,
		_w21496_
	);
	LUT2 #(
		.INIT('h2)
	) name17450 (
		\pio_PIO_RES_OUT_reg[1]/P0001 ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w21497_
	);
	LUT2 #(
		.INIT('h4)
	) name17451 (
		\pio_PIO_RES_OUT_reg[1]/P0001 ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w21498_
	);
	LUT2 #(
		.INIT('h1)
	) name17452 (
		_w21497_,
		_w21498_,
		_w21499_
	);
	LUT2 #(
		.INIT('h4)
	) name17453 (
		\PIO_oe[1]_pad ,
		\pio_pmask_reg_DO_reg[1]/NET0131 ,
		_w21500_
	);
	LUT2 #(
		.INIT('h4)
	) name17454 (
		_w21499_,
		_w21500_,
		_w21501_
	);
	LUT2 #(
		.INIT('h1)
	) name17455 (
		\pio_PINT_reg[1]/NET0131 ,
		_w21501_,
		_w21502_
	);
	LUT2 #(
		.INIT('h4)
	) name17456 (
		_w21291_,
		_w21502_,
		_w21503_
	);
	LUT2 #(
		.INIT('h4)
	) name17457 (
		_w9435_,
		_w21291_,
		_w21504_
	);
	LUT2 #(
		.INIT('h1)
	) name17458 (
		_w21503_,
		_w21504_,
		_w21505_
	);
	LUT2 #(
		.INIT('h2)
	) name17459 (
		\pio_PIO_RES_OUT_reg[3]/P0001 ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w21506_
	);
	LUT2 #(
		.INIT('h4)
	) name17460 (
		\pio_PIO_RES_OUT_reg[3]/P0001 ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w21507_
	);
	LUT2 #(
		.INIT('h1)
	) name17461 (
		_w21506_,
		_w21507_,
		_w21508_
	);
	LUT2 #(
		.INIT('h4)
	) name17462 (
		\PIO_oe[3]_pad ,
		\pio_pmask_reg_DO_reg[3]/NET0131 ,
		_w21509_
	);
	LUT2 #(
		.INIT('h4)
	) name17463 (
		_w21508_,
		_w21509_,
		_w21510_
	);
	LUT2 #(
		.INIT('h1)
	) name17464 (
		\pio_PINT_reg[3]/NET0131 ,
		_w21510_,
		_w21511_
	);
	LUT2 #(
		.INIT('h4)
	) name17465 (
		_w21291_,
		_w21511_,
		_w21512_
	);
	LUT2 #(
		.INIT('h4)
	) name17466 (
		_w8113_,
		_w21291_,
		_w21513_
	);
	LUT2 #(
		.INIT('h1)
	) name17467 (
		_w21512_,
		_w21513_,
		_w21514_
	);
	LUT2 #(
		.INIT('h2)
	) name17468 (
		\pio_PIO_RES_OUT_reg[6]/P0001 ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w21515_
	);
	LUT2 #(
		.INIT('h4)
	) name17469 (
		\pio_PIO_RES_OUT_reg[6]/P0001 ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w21516_
	);
	LUT2 #(
		.INIT('h1)
	) name17470 (
		_w21515_,
		_w21516_,
		_w21517_
	);
	LUT2 #(
		.INIT('h4)
	) name17471 (
		\PIO_oe[6]_pad ,
		\pio_pmask_reg_DO_reg[6]/NET0131 ,
		_w21518_
	);
	LUT2 #(
		.INIT('h4)
	) name17472 (
		_w21517_,
		_w21518_,
		_w21519_
	);
	LUT2 #(
		.INIT('h1)
	) name17473 (
		\pio_PINT_reg[6]/NET0131 ,
		_w21519_,
		_w21520_
	);
	LUT2 #(
		.INIT('h4)
	) name17474 (
		_w21291_,
		_w21520_,
		_w21521_
	);
	LUT2 #(
		.INIT('h4)
	) name17475 (
		_w11525_,
		_w21291_,
		_w21522_
	);
	LUT2 #(
		.INIT('h1)
	) name17476 (
		_w21521_,
		_w21522_,
		_w21523_
	);
	LUT2 #(
		.INIT('h2)
	) name17477 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[15]/P0001 ,
		_w20468_,
		_w21524_
	);
	LUT2 #(
		.INIT('h8)
	) name17478 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w14728_,
		_w21525_
	);
	LUT2 #(
		.INIT('h8)
	) name17479 (
		_w5664_,
		_w21525_,
		_w21526_
	);
	LUT2 #(
		.INIT('h8)
	) name17480 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w21527_
	);
	LUT2 #(
		.INIT('h8)
	) name17481 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w21527_,
		_w21528_
	);
	LUT2 #(
		.INIT('h2)
	) name17482 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w21528_,
		_w21529_
	);
	LUT2 #(
		.INIT('h4)
	) name17483 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w21530_
	);
	LUT2 #(
		.INIT('h8)
	) name17484 (
		_w21528_,
		_w21530_,
		_w21531_
	);
	LUT2 #(
		.INIT('h1)
	) name17485 (
		_w20477_,
		_w21529_,
		_w21532_
	);
	LUT2 #(
		.INIT('h4)
	) name17486 (
		_w21531_,
		_w21532_,
		_w21533_
	);
	LUT2 #(
		.INIT('h2)
	) name17487 (
		_w21526_,
		_w21533_,
		_w21534_
	);
	LUT2 #(
		.INIT('h1)
	) name17488 (
		_w21524_,
		_w21534_,
		_w21535_
	);
	LUT2 #(
		.INIT('h2)
	) name17489 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[14]/P0001 ,
		_w20468_,
		_w21536_
	);
	LUT2 #(
		.INIT('h8)
	) name17490 (
		_w20464_,
		_w21528_,
		_w21537_
	);
	LUT2 #(
		.INIT('h1)
	) name17491 (
		_w20486_,
		_w21529_,
		_w21538_
	);
	LUT2 #(
		.INIT('h4)
	) name17492 (
		_w21537_,
		_w21538_,
		_w21539_
	);
	LUT2 #(
		.INIT('h2)
	) name17493 (
		_w21526_,
		_w21539_,
		_w21540_
	);
	LUT2 #(
		.INIT('h1)
	) name17494 (
		_w21536_,
		_w21540_,
		_w21541_
	);
	LUT2 #(
		.INIT('h2)
	) name17495 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[13]/P0001 ,
		_w20468_,
		_w21542_
	);
	LUT2 #(
		.INIT('h4)
	) name17496 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w21527_,
		_w21543_
	);
	LUT2 #(
		.INIT('h2)
	) name17497 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w21543_,
		_w21544_
	);
	LUT2 #(
		.INIT('h8)
	) name17498 (
		_w21530_,
		_w21543_,
		_w21545_
	);
	LUT2 #(
		.INIT('h1)
	) name17499 (
		_w20477_,
		_w21544_,
		_w21546_
	);
	LUT2 #(
		.INIT('h4)
	) name17500 (
		_w21545_,
		_w21546_,
		_w21547_
	);
	LUT2 #(
		.INIT('h2)
	) name17501 (
		_w21526_,
		_w21547_,
		_w21548_
	);
	LUT2 #(
		.INIT('h1)
	) name17502 (
		_w21542_,
		_w21548_,
		_w21549_
	);
	LUT2 #(
		.INIT('h2)
	) name17503 (
		\core_eu_ea_alu_ea_dec_piconst_DO_reg[12]/P0001 ,
		_w20468_,
		_w21550_
	);
	LUT2 #(
		.INIT('h8)
	) name17504 (
		_w20464_,
		_w21543_,
		_w21551_
	);
	LUT2 #(
		.INIT('h1)
	) name17505 (
		_w20486_,
		_w21544_,
		_w21552_
	);
	LUT2 #(
		.INIT('h4)
	) name17506 (
		_w21551_,
		_w21552_,
		_w21553_
	);
	LUT2 #(
		.INIT('h2)
	) name17507 (
		_w21526_,
		_w21553_,
		_w21554_
	);
	LUT2 #(
		.INIT('h1)
	) name17508 (
		_w21550_,
		_w21554_,
		_w21555_
	);
	LUT2 #(
		.INIT('h8)
	) name17509 (
		_w6027_,
		_w20606_,
		_w21556_
	);
	LUT2 #(
		.INIT('h4)
	) name17510 (
		_w4117_,
		_w21556_,
		_w21557_
	);
	LUT2 #(
		.INIT('h8)
	) name17511 (
		_w6115_,
		_w21557_,
		_w21558_
	);
	LUT2 #(
		.INIT('h4)
	) name17512 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w5615_,
		_w21559_
	);
	LUT2 #(
		.INIT('h8)
	) name17513 (
		_w19698_,
		_w21559_,
		_w21560_
	);
	LUT2 #(
		.INIT('h1)
	) name17514 (
		_w20377_,
		_w21558_,
		_w21561_
	);
	LUT2 #(
		.INIT('h4)
	) name17515 (
		_w21560_,
		_w21561_,
		_w21562_
	);
	LUT2 #(
		.INIT('h4)
	) name17516 (
		\sport0_rxctl_RXSHT_reg[4]/P0001 ,
		_w20868_,
		_w21563_
	);
	LUT2 #(
		.INIT('h8)
	) name17517 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20873_,
		_w21564_
	);
	LUT2 #(
		.INIT('h4)
	) name17518 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w10069_,
		_w21565_
	);
	LUT2 #(
		.INIT('h1)
	) name17519 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w20956_,
		_w21566_
	);
	LUT2 #(
		.INIT('h2)
	) name17520 (
		_w20949_,
		_w21566_,
		_w21567_
	);
	LUT2 #(
		.INIT('h4)
	) name17521 (
		_w20949_,
		_w21566_,
		_w21568_
	);
	LUT2 #(
		.INIT('h2)
	) name17522 (
		_w20875_,
		_w21567_,
		_w21569_
	);
	LUT2 #(
		.INIT('h4)
	) name17523 (
		_w21568_,
		_w21569_,
		_w21570_
	);
	LUT2 #(
		.INIT('h1)
	) name17524 (
		_w20868_,
		_w21564_,
		_w21571_
	);
	LUT2 #(
		.INIT('h4)
	) name17525 (
		_w21570_,
		_w21571_,
		_w21572_
	);
	LUT2 #(
		.INIT('h4)
	) name17526 (
		_w21565_,
		_w21572_,
		_w21573_
	);
	LUT2 #(
		.INIT('h1)
	) name17527 (
		_w20871_,
		_w21563_,
		_w21574_
	);
	LUT2 #(
		.INIT('h4)
	) name17528 (
		_w21573_,
		_w21574_,
		_w21575_
	);
	LUT2 #(
		.INIT('h8)
	) name17529 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20871_,
		_w21576_
	);
	LUT2 #(
		.INIT('h1)
	) name17530 (
		_w21575_,
		_w21576_,
		_w21577_
	);
	LUT2 #(
		.INIT('h2)
	) name17531 (
		_w5692_,
		_w5936_,
		_w21578_
	);
	LUT2 #(
		.INIT('h4)
	) name17532 (
		_w19705_,
		_w21578_,
		_w21579_
	);
	LUT2 #(
		.INIT('h2)
	) name17533 (
		\pio_PIO_RES_OUT_reg[7]/P0001 ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w21580_
	);
	LUT2 #(
		.INIT('h4)
	) name17534 (
		\pio_PIO_RES_OUT_reg[7]/P0001 ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w21581_
	);
	LUT2 #(
		.INIT('h1)
	) name17535 (
		_w21580_,
		_w21581_,
		_w21582_
	);
	LUT2 #(
		.INIT('h4)
	) name17536 (
		\PIO_oe[7]_pad ,
		\pio_pmask_reg_DO_reg[7]/NET0131 ,
		_w21583_
	);
	LUT2 #(
		.INIT('h4)
	) name17537 (
		_w21582_,
		_w21583_,
		_w21584_
	);
	LUT2 #(
		.INIT('h1)
	) name17538 (
		\pio_PINT_reg[7]/NET0131 ,
		_w21584_,
		_w21585_
	);
	LUT2 #(
		.INIT('h4)
	) name17539 (
		_w21291_,
		_w21585_,
		_w21586_
	);
	LUT2 #(
		.INIT('h4)
	) name17540 (
		_w11265_,
		_w21291_,
		_w21587_
	);
	LUT2 #(
		.INIT('h1)
	) name17541 (
		_w21586_,
		_w21587_,
		_w21588_
	);
	LUT2 #(
		.INIT('h4)
	) name17542 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w19699_,
		_w21589_
	);
	LUT2 #(
		.INIT('h2)
	) name17543 (
		_w6111_,
		_w21589_,
		_w21590_
	);
	LUT2 #(
		.INIT('h1)
	) name17544 (
		_w4117_,
		_w21590_,
		_w21591_
	);
	LUT2 #(
		.INIT('h2)
	) name17545 (
		_w21578_,
		_w21591_,
		_w21592_
	);
	LUT2 #(
		.INIT('h2)
	) name17546 (
		\core_c_psq_SSTAT_reg[4]/NET0131 ,
		_w18217_,
		_w21593_
	);
	LUT2 #(
		.INIT('h4)
	) name17547 (
		_w18680_,
		_w21593_,
		_w21594_
	);
	LUT2 #(
		.INIT('h1)
	) name17548 (
		_w14695_,
		_w14702_,
		_w21595_
	);
	LUT2 #(
		.INIT('h1)
	) name17549 (
		_w14693_,
		_w21595_,
		_w21596_
	);
	LUT2 #(
		.INIT('h8)
	) name17550 (
		_w18680_,
		_w21596_,
		_w21597_
	);
	LUT2 #(
		.INIT('h1)
	) name17551 (
		_w21594_,
		_w21597_,
		_w21598_
	);
	LUT2 #(
		.INIT('h2)
	) name17552 (
		\emc_PMDoe_reg/NET0131 ,
		_w19049_,
		_w21599_
	);
	LUT2 #(
		.INIT('h4)
	) name17553 (
		_w19056_,
		_w21599_,
		_w21600_
	);
	LUT2 #(
		.INIT('h1)
	) name17554 (
		_w20345_,
		_w21600_,
		_w21601_
	);
	LUT2 #(
		.INIT('h1)
	) name17555 (
		_w14698_,
		_w14710_,
		_w21602_
	);
	LUT2 #(
		.INIT('h4)
	) name17556 (
		_w18220_,
		_w21602_,
		_w21603_
	);
	LUT2 #(
		.INIT('h1)
	) name17557 (
		_w18688_,
		_w21602_,
		_w21604_
	);
	LUT2 #(
		.INIT('h1)
	) name17558 (
		_w21603_,
		_w21604_,
		_w21605_
	);
	LUT2 #(
		.INIT('h8)
	) name17559 (
		_w4851_,
		_w20576_,
		_w21606_
	);
	LUT2 #(
		.INIT('h2)
	) name17560 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][9]/P0001 ,
		_w21606_,
		_w21607_
	);
	LUT2 #(
		.INIT('h8)
	) name17561 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w21606_,
		_w21608_
	);
	LUT2 #(
		.INIT('h1)
	) name17562 (
		_w21607_,
		_w21608_,
		_w21609_
	);
	LUT2 #(
		.INIT('h2)
	) name17563 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][8]/P0001 ,
		_w21606_,
		_w21610_
	);
	LUT2 #(
		.INIT('h8)
	) name17564 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w21606_,
		_w21611_
	);
	LUT2 #(
		.INIT('h1)
	) name17565 (
		_w21610_,
		_w21611_,
		_w21612_
	);
	LUT2 #(
		.INIT('h2)
	) name17566 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][7]/P0001 ,
		_w21606_,
		_w21613_
	);
	LUT2 #(
		.INIT('h8)
	) name17567 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w21606_,
		_w21614_
	);
	LUT2 #(
		.INIT('h1)
	) name17568 (
		_w21613_,
		_w21614_,
		_w21615_
	);
	LUT2 #(
		.INIT('h2)
	) name17569 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][6]/P0001 ,
		_w21606_,
		_w21616_
	);
	LUT2 #(
		.INIT('h8)
	) name17570 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w21606_,
		_w21617_
	);
	LUT2 #(
		.INIT('h1)
	) name17571 (
		_w21616_,
		_w21617_,
		_w21618_
	);
	LUT2 #(
		.INIT('h2)
	) name17572 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][5]/P0001 ,
		_w21606_,
		_w21619_
	);
	LUT2 #(
		.INIT('h8)
	) name17573 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w21606_,
		_w21620_
	);
	LUT2 #(
		.INIT('h1)
	) name17574 (
		_w21619_,
		_w21620_,
		_w21621_
	);
	LUT2 #(
		.INIT('h2)
	) name17575 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][4]/P0001 ,
		_w21606_,
		_w21622_
	);
	LUT2 #(
		.INIT('h8)
	) name17576 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w21606_,
		_w21623_
	);
	LUT2 #(
		.INIT('h1)
	) name17577 (
		_w21622_,
		_w21623_,
		_w21624_
	);
	LUT2 #(
		.INIT('h2)
	) name17578 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][21]/P0001 ,
		_w21606_,
		_w21625_
	);
	LUT2 #(
		.INIT('h8)
	) name17579 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w21606_,
		_w21626_
	);
	LUT2 #(
		.INIT('h1)
	) name17580 (
		_w21625_,
		_w21626_,
		_w21627_
	);
	LUT2 #(
		.INIT('h2)
	) name17581 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][20]/P0001 ,
		_w21606_,
		_w21628_
	);
	LUT2 #(
		.INIT('h8)
	) name17582 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w21606_,
		_w21629_
	);
	LUT2 #(
		.INIT('h1)
	) name17583 (
		_w21628_,
		_w21629_,
		_w21630_
	);
	LUT2 #(
		.INIT('h2)
	) name17584 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][19]/P0001 ,
		_w21606_,
		_w21631_
	);
	LUT2 #(
		.INIT('h8)
	) name17585 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w21606_,
		_w21632_
	);
	LUT2 #(
		.INIT('h1)
	) name17586 (
		_w21631_,
		_w21632_,
		_w21633_
	);
	LUT2 #(
		.INIT('h2)
	) name17587 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][18]/P0001 ,
		_w21606_,
		_w21634_
	);
	LUT2 #(
		.INIT('h8)
	) name17588 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w21606_,
		_w21635_
	);
	LUT2 #(
		.INIT('h1)
	) name17589 (
		_w21634_,
		_w21635_,
		_w21636_
	);
	LUT2 #(
		.INIT('h2)
	) name17590 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][17]/P0001 ,
		_w21606_,
		_w21637_
	);
	LUT2 #(
		.INIT('h8)
	) name17591 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w21606_,
		_w21638_
	);
	LUT2 #(
		.INIT('h1)
	) name17592 (
		_w21637_,
		_w21638_,
		_w21639_
	);
	LUT2 #(
		.INIT('h2)
	) name17593 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][16]/P0001 ,
		_w21606_,
		_w21640_
	);
	LUT2 #(
		.INIT('h8)
	) name17594 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w21606_,
		_w21641_
	);
	LUT2 #(
		.INIT('h1)
	) name17595 (
		_w21640_,
		_w21641_,
		_w21642_
	);
	LUT2 #(
		.INIT('h2)
	) name17596 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][15]/P0001 ,
		_w21606_,
		_w21643_
	);
	LUT2 #(
		.INIT('h8)
	) name17597 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w21606_,
		_w21644_
	);
	LUT2 #(
		.INIT('h1)
	) name17598 (
		_w21643_,
		_w21644_,
		_w21645_
	);
	LUT2 #(
		.INIT('h2)
	) name17599 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][14]/P0001 ,
		_w21606_,
		_w21646_
	);
	LUT2 #(
		.INIT('h8)
	) name17600 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w21606_,
		_w21647_
	);
	LUT2 #(
		.INIT('h1)
	) name17601 (
		_w21646_,
		_w21647_,
		_w21648_
	);
	LUT2 #(
		.INIT('h2)
	) name17602 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][13]/P0001 ,
		_w21606_,
		_w21649_
	);
	LUT2 #(
		.INIT('h8)
	) name17603 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w21606_,
		_w21650_
	);
	LUT2 #(
		.INIT('h1)
	) name17604 (
		_w21649_,
		_w21650_,
		_w21651_
	);
	LUT2 #(
		.INIT('h2)
	) name17605 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][12]/P0001 ,
		_w21606_,
		_w21652_
	);
	LUT2 #(
		.INIT('h8)
	) name17606 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w21606_,
		_w21653_
	);
	LUT2 #(
		.INIT('h1)
	) name17607 (
		_w21652_,
		_w21653_,
		_w21654_
	);
	LUT2 #(
		.INIT('h2)
	) name17608 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][11]/P0001 ,
		_w21606_,
		_w21655_
	);
	LUT2 #(
		.INIT('h8)
	) name17609 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w21606_,
		_w21656_
	);
	LUT2 #(
		.INIT('h1)
	) name17610 (
		_w21655_,
		_w21656_,
		_w21657_
	);
	LUT2 #(
		.INIT('h2)
	) name17611 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][10]/P0001 ,
		_w21606_,
		_w21658_
	);
	LUT2 #(
		.INIT('h8)
	) name17612 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w21606_,
		_w21659_
	);
	LUT2 #(
		.INIT('h1)
	) name17613 (
		_w21658_,
		_w21659_,
		_w21660_
	);
	LUT2 #(
		.INIT('h1)
	) name17614 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8113_,
		_w21661_
	);
	LUT2 #(
		.INIT('h2)
	) name17615 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12870_,
		_w21662_
	);
	LUT2 #(
		.INIT('h1)
	) name17616 (
		_w21661_,
		_w21662_,
		_w21663_
	);
	LUT2 #(
		.INIT('h2)
	) name17617 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w21663_,
		_w21664_
	);
	LUT2 #(
		.INIT('h8)
	) name17618 (
		_w18088_,
		_w19801_,
		_w21665_
	);
	LUT2 #(
		.INIT('h2)
	) name17619 (
		_w18111_,
		_w19818_,
		_w21666_
	);
	LUT2 #(
		.INIT('h2)
	) name17620 (
		_w18171_,
		_w19857_,
		_w21667_
	);
	LUT2 #(
		.INIT('h2)
	) name17621 (
		_w18115_,
		_w18775_,
		_w21668_
	);
	LUT2 #(
		.INIT('h2)
	) name17622 (
		_w17925_,
		_w18895_,
		_w21669_
	);
	LUT2 #(
		.INIT('h2)
	) name17623 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7991_,
		_w21670_
	);
	LUT2 #(
		.INIT('h8)
	) name17624 (
		_w18046_,
		_w18758_,
		_w21671_
	);
	LUT2 #(
		.INIT('h8)
	) name17625 (
		_w18001_,
		_w19720_,
		_w21672_
	);
	LUT2 #(
		.INIT('h1)
	) name17626 (
		_w17922_,
		_w18129_,
		_w21673_
	);
	LUT2 #(
		.INIT('h8)
	) name17627 (
		_w18147_,
		_w18187_,
		_w21674_
	);
	LUT2 #(
		.INIT('h4)
	) name17628 (
		_w18175_,
		_w20104_,
		_w21675_
	);
	LUT2 #(
		.INIT('h2)
	) name17629 (
		_w17986_,
		_w18189_,
		_w21676_
	);
	LUT2 #(
		.INIT('h1)
	) name17630 (
		_w17933_,
		_w18781_,
		_w21677_
	);
	LUT2 #(
		.INIT('h1)
	) name17631 (
		_w18091_,
		_w18167_,
		_w21678_
	);
	LUT2 #(
		.INIT('h1)
	) name17632 (
		_w18104_,
		_w18108_,
		_w21679_
	);
	LUT2 #(
		.INIT('h8)
	) name17633 (
		_w18043_,
		_w18183_,
		_w21680_
	);
	LUT2 #(
		.INIT('h8)
	) name17634 (
		_w18136_,
		_w18153_,
		_w21681_
	);
	LUT2 #(
		.INIT('h1)
	) name17635 (
		_w21670_,
		_w21672_,
		_w21682_
	);
	LUT2 #(
		.INIT('h1)
	) name17636 (
		_w21676_,
		_w21681_,
		_w21683_
	);
	LUT2 #(
		.INIT('h8)
	) name17637 (
		_w21682_,
		_w21683_,
		_w21684_
	);
	LUT2 #(
		.INIT('h4)
	) name17638 (
		_w17972_,
		_w21684_,
		_w21685_
	);
	LUT2 #(
		.INIT('h1)
	) name17639 (
		_w21665_,
		_w21671_,
		_w21686_
	);
	LUT2 #(
		.INIT('h1)
	) name17640 (
		_w21673_,
		_w21674_,
		_w21687_
	);
	LUT2 #(
		.INIT('h1)
	) name17641 (
		_w21678_,
		_w21679_,
		_w21688_
	);
	LUT2 #(
		.INIT('h4)
	) name17642 (
		_w21680_,
		_w21688_,
		_w21689_
	);
	LUT2 #(
		.INIT('h8)
	) name17643 (
		_w21686_,
		_w21687_,
		_w21690_
	);
	LUT2 #(
		.INIT('h4)
	) name17644 (
		_w21666_,
		_w21685_,
		_w21691_
	);
	LUT2 #(
		.INIT('h1)
	) name17645 (
		_w21667_,
		_w21668_,
		_w21692_
	);
	LUT2 #(
		.INIT('h1)
	) name17646 (
		_w21669_,
		_w21675_,
		_w21693_
	);
	LUT2 #(
		.INIT('h4)
	) name17647 (
		_w21677_,
		_w21693_,
		_w21694_
	);
	LUT2 #(
		.INIT('h8)
	) name17648 (
		_w21691_,
		_w21692_,
		_w21695_
	);
	LUT2 #(
		.INIT('h8)
	) name17649 (
		_w21689_,
		_w21690_,
		_w21696_
	);
	LUT2 #(
		.INIT('h8)
	) name17650 (
		_w20087_,
		_w21696_,
		_w21697_
	);
	LUT2 #(
		.INIT('h8)
	) name17651 (
		_w21694_,
		_w21695_,
		_w21698_
	);
	LUT2 #(
		.INIT('h8)
	) name17652 (
		_w21697_,
		_w21698_,
		_w21699_
	);
	LUT2 #(
		.INIT('h8)
	) name17653 (
		_w21084_,
		_w21699_,
		_w21700_
	);
	LUT2 #(
		.INIT('h4)
	) name17654 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w21700_,
		_w21701_
	);
	LUT2 #(
		.INIT('h1)
	) name17655 (
		_w21664_,
		_w21701_,
		_w21702_
	);
	LUT2 #(
		.INIT('h2)
	) name17656 (
		_w18717_,
		_w21702_,
		_w21703_
	);
	LUT2 #(
		.INIT('h1)
	) name17657 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[3]/P0001 ,
		_w18717_,
		_w21704_
	);
	LUT2 #(
		.INIT('h1)
	) name17658 (
		_w21703_,
		_w21704_,
		_w21705_
	);
	LUT2 #(
		.INIT('h8)
	) name17659 (
		_w4847_,
		_w20576_,
		_w21706_
	);
	LUT2 #(
		.INIT('h2)
	) name17660 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][9]/P0001 ,
		_w21706_,
		_w21707_
	);
	LUT2 #(
		.INIT('h8)
	) name17661 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w21706_,
		_w21708_
	);
	LUT2 #(
		.INIT('h1)
	) name17662 (
		_w21707_,
		_w21708_,
		_w21709_
	);
	LUT2 #(
		.INIT('h2)
	) name17663 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][8]/P0001 ,
		_w21706_,
		_w21710_
	);
	LUT2 #(
		.INIT('h8)
	) name17664 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w21706_,
		_w21711_
	);
	LUT2 #(
		.INIT('h1)
	) name17665 (
		_w21710_,
		_w21711_,
		_w21712_
	);
	LUT2 #(
		.INIT('h2)
	) name17666 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][7]/P0001 ,
		_w21706_,
		_w21713_
	);
	LUT2 #(
		.INIT('h8)
	) name17667 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w21706_,
		_w21714_
	);
	LUT2 #(
		.INIT('h1)
	) name17668 (
		_w21713_,
		_w21714_,
		_w21715_
	);
	LUT2 #(
		.INIT('h2)
	) name17669 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][6]/P0001 ,
		_w21706_,
		_w21716_
	);
	LUT2 #(
		.INIT('h8)
	) name17670 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w21706_,
		_w21717_
	);
	LUT2 #(
		.INIT('h1)
	) name17671 (
		_w21716_,
		_w21717_,
		_w21718_
	);
	LUT2 #(
		.INIT('h2)
	) name17672 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][5]/P0001 ,
		_w21706_,
		_w21719_
	);
	LUT2 #(
		.INIT('h8)
	) name17673 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w21706_,
		_w21720_
	);
	LUT2 #(
		.INIT('h1)
	) name17674 (
		_w21719_,
		_w21720_,
		_w21721_
	);
	LUT2 #(
		.INIT('h2)
	) name17675 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][4]/P0001 ,
		_w21706_,
		_w21722_
	);
	LUT2 #(
		.INIT('h8)
	) name17676 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w21706_,
		_w21723_
	);
	LUT2 #(
		.INIT('h1)
	) name17677 (
		_w21722_,
		_w21723_,
		_w21724_
	);
	LUT2 #(
		.INIT('h2)
	) name17678 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][21]/P0001 ,
		_w21706_,
		_w21725_
	);
	LUT2 #(
		.INIT('h8)
	) name17679 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w21706_,
		_w21726_
	);
	LUT2 #(
		.INIT('h1)
	) name17680 (
		_w21725_,
		_w21726_,
		_w21727_
	);
	LUT2 #(
		.INIT('h2)
	) name17681 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][20]/P0001 ,
		_w21706_,
		_w21728_
	);
	LUT2 #(
		.INIT('h8)
	) name17682 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w21706_,
		_w21729_
	);
	LUT2 #(
		.INIT('h1)
	) name17683 (
		_w21728_,
		_w21729_,
		_w21730_
	);
	LUT2 #(
		.INIT('h2)
	) name17684 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][19]/P0001 ,
		_w21706_,
		_w21731_
	);
	LUT2 #(
		.INIT('h8)
	) name17685 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w21706_,
		_w21732_
	);
	LUT2 #(
		.INIT('h1)
	) name17686 (
		_w21731_,
		_w21732_,
		_w21733_
	);
	LUT2 #(
		.INIT('h2)
	) name17687 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][18]/P0001 ,
		_w21706_,
		_w21734_
	);
	LUT2 #(
		.INIT('h8)
	) name17688 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w21706_,
		_w21735_
	);
	LUT2 #(
		.INIT('h1)
	) name17689 (
		_w21734_,
		_w21735_,
		_w21736_
	);
	LUT2 #(
		.INIT('h2)
	) name17690 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][17]/P0001 ,
		_w21706_,
		_w21737_
	);
	LUT2 #(
		.INIT('h8)
	) name17691 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w21706_,
		_w21738_
	);
	LUT2 #(
		.INIT('h1)
	) name17692 (
		_w21737_,
		_w21738_,
		_w21739_
	);
	LUT2 #(
		.INIT('h2)
	) name17693 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][16]/P0001 ,
		_w21706_,
		_w21740_
	);
	LUT2 #(
		.INIT('h8)
	) name17694 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w21706_,
		_w21741_
	);
	LUT2 #(
		.INIT('h1)
	) name17695 (
		_w21740_,
		_w21741_,
		_w21742_
	);
	LUT2 #(
		.INIT('h2)
	) name17696 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][15]/P0001 ,
		_w21706_,
		_w21743_
	);
	LUT2 #(
		.INIT('h8)
	) name17697 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w21706_,
		_w21744_
	);
	LUT2 #(
		.INIT('h1)
	) name17698 (
		_w21743_,
		_w21744_,
		_w21745_
	);
	LUT2 #(
		.INIT('h2)
	) name17699 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][14]/P0001 ,
		_w21706_,
		_w21746_
	);
	LUT2 #(
		.INIT('h8)
	) name17700 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w21706_,
		_w21747_
	);
	LUT2 #(
		.INIT('h1)
	) name17701 (
		_w21746_,
		_w21747_,
		_w21748_
	);
	LUT2 #(
		.INIT('h2)
	) name17702 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][13]/P0001 ,
		_w21706_,
		_w21749_
	);
	LUT2 #(
		.INIT('h8)
	) name17703 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w21706_,
		_w21750_
	);
	LUT2 #(
		.INIT('h1)
	) name17704 (
		_w21749_,
		_w21750_,
		_w21751_
	);
	LUT2 #(
		.INIT('h2)
	) name17705 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][12]/P0001 ,
		_w21706_,
		_w21752_
	);
	LUT2 #(
		.INIT('h8)
	) name17706 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w21706_,
		_w21753_
	);
	LUT2 #(
		.INIT('h1)
	) name17707 (
		_w21752_,
		_w21753_,
		_w21754_
	);
	LUT2 #(
		.INIT('h2)
	) name17708 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][11]/P0001 ,
		_w21706_,
		_w21755_
	);
	LUT2 #(
		.INIT('h8)
	) name17709 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w21706_,
		_w21756_
	);
	LUT2 #(
		.INIT('h1)
	) name17710 (
		_w21755_,
		_w21756_,
		_w21757_
	);
	LUT2 #(
		.INIT('h2)
	) name17711 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][10]/P0001 ,
		_w21706_,
		_w21758_
	);
	LUT2 #(
		.INIT('h8)
	) name17712 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w21706_,
		_w21759_
	);
	LUT2 #(
		.INIT('h1)
	) name17713 (
		_w21758_,
		_w21759_,
		_w21760_
	);
	LUT2 #(
		.INIT('h8)
	) name17714 (
		_w20575_,
		_w20597_,
		_w21761_
	);
	LUT2 #(
		.INIT('h2)
	) name17715 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][9]/P0001 ,
		_w21761_,
		_w21762_
	);
	LUT2 #(
		.INIT('h8)
	) name17716 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w21761_,
		_w21763_
	);
	LUT2 #(
		.INIT('h1)
	) name17717 (
		_w21762_,
		_w21763_,
		_w21764_
	);
	LUT2 #(
		.INIT('h2)
	) name17718 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][8]/P0001 ,
		_w21761_,
		_w21765_
	);
	LUT2 #(
		.INIT('h8)
	) name17719 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w21761_,
		_w21766_
	);
	LUT2 #(
		.INIT('h1)
	) name17720 (
		_w21765_,
		_w21766_,
		_w21767_
	);
	LUT2 #(
		.INIT('h2)
	) name17721 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][7]/P0001 ,
		_w21761_,
		_w21768_
	);
	LUT2 #(
		.INIT('h8)
	) name17722 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w21761_,
		_w21769_
	);
	LUT2 #(
		.INIT('h1)
	) name17723 (
		_w21768_,
		_w21769_,
		_w21770_
	);
	LUT2 #(
		.INIT('h2)
	) name17724 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][6]/P0001 ,
		_w21761_,
		_w21771_
	);
	LUT2 #(
		.INIT('h8)
	) name17725 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w21761_,
		_w21772_
	);
	LUT2 #(
		.INIT('h1)
	) name17726 (
		_w21771_,
		_w21772_,
		_w21773_
	);
	LUT2 #(
		.INIT('h2)
	) name17727 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][5]/P0001 ,
		_w21761_,
		_w21774_
	);
	LUT2 #(
		.INIT('h8)
	) name17728 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w21761_,
		_w21775_
	);
	LUT2 #(
		.INIT('h1)
	) name17729 (
		_w21774_,
		_w21775_,
		_w21776_
	);
	LUT2 #(
		.INIT('h2)
	) name17730 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][4]/P0001 ,
		_w21761_,
		_w21777_
	);
	LUT2 #(
		.INIT('h8)
	) name17731 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w21761_,
		_w21778_
	);
	LUT2 #(
		.INIT('h1)
	) name17732 (
		_w21777_,
		_w21778_,
		_w21779_
	);
	LUT2 #(
		.INIT('h2)
	) name17733 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][21]/P0001 ,
		_w21761_,
		_w21780_
	);
	LUT2 #(
		.INIT('h8)
	) name17734 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w21761_,
		_w21781_
	);
	LUT2 #(
		.INIT('h1)
	) name17735 (
		_w21780_,
		_w21781_,
		_w21782_
	);
	LUT2 #(
		.INIT('h2)
	) name17736 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][20]/P0001 ,
		_w21761_,
		_w21783_
	);
	LUT2 #(
		.INIT('h8)
	) name17737 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w21761_,
		_w21784_
	);
	LUT2 #(
		.INIT('h1)
	) name17738 (
		_w21783_,
		_w21784_,
		_w21785_
	);
	LUT2 #(
		.INIT('h2)
	) name17739 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][19]/P0001 ,
		_w21761_,
		_w21786_
	);
	LUT2 #(
		.INIT('h8)
	) name17740 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w21761_,
		_w21787_
	);
	LUT2 #(
		.INIT('h1)
	) name17741 (
		_w21786_,
		_w21787_,
		_w21788_
	);
	LUT2 #(
		.INIT('h2)
	) name17742 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][18]/P0001 ,
		_w21761_,
		_w21789_
	);
	LUT2 #(
		.INIT('h8)
	) name17743 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w21761_,
		_w21790_
	);
	LUT2 #(
		.INIT('h1)
	) name17744 (
		_w21789_,
		_w21790_,
		_w21791_
	);
	LUT2 #(
		.INIT('h2)
	) name17745 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][17]/P0001 ,
		_w21761_,
		_w21792_
	);
	LUT2 #(
		.INIT('h8)
	) name17746 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w21761_,
		_w21793_
	);
	LUT2 #(
		.INIT('h1)
	) name17747 (
		_w21792_,
		_w21793_,
		_w21794_
	);
	LUT2 #(
		.INIT('h2)
	) name17748 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][16]/P0001 ,
		_w21761_,
		_w21795_
	);
	LUT2 #(
		.INIT('h8)
	) name17749 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w21761_,
		_w21796_
	);
	LUT2 #(
		.INIT('h1)
	) name17750 (
		_w21795_,
		_w21796_,
		_w21797_
	);
	LUT2 #(
		.INIT('h2)
	) name17751 (
		_w13806_,
		_w14649_,
		_w21798_
	);
	LUT2 #(
		.INIT('h1)
	) name17752 (
		_w13806_,
		_w20053_,
		_w21799_
	);
	LUT2 #(
		.INIT('h1)
	) name17753 (
		_w21798_,
		_w21799_,
		_w21800_
	);
	LUT2 #(
		.INIT('h2)
	) name17754 (
		_w14667_,
		_w21800_,
		_w21801_
	);
	LUT2 #(
		.INIT('h2)
	) name17755 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[10]/P0001 ,
		_w14667_,
		_w21802_
	);
	LUT2 #(
		.INIT('h1)
	) name17756 (
		_w21801_,
		_w21802_,
		_w21803_
	);
	LUT2 #(
		.INIT('h2)
	) name17757 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][15]/P0001 ,
		_w21761_,
		_w21804_
	);
	LUT2 #(
		.INIT('h8)
	) name17758 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w21761_,
		_w21805_
	);
	LUT2 #(
		.INIT('h1)
	) name17759 (
		_w21804_,
		_w21805_,
		_w21806_
	);
	LUT2 #(
		.INIT('h2)
	) name17760 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][14]/P0001 ,
		_w21761_,
		_w21807_
	);
	LUT2 #(
		.INIT('h8)
	) name17761 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w21761_,
		_w21808_
	);
	LUT2 #(
		.INIT('h1)
	) name17762 (
		_w21807_,
		_w21808_,
		_w21809_
	);
	LUT2 #(
		.INIT('h2)
	) name17763 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][12]/P0001 ,
		_w21761_,
		_w21810_
	);
	LUT2 #(
		.INIT('h8)
	) name17764 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w21761_,
		_w21811_
	);
	LUT2 #(
		.INIT('h1)
	) name17765 (
		_w21810_,
		_w21811_,
		_w21812_
	);
	LUT2 #(
		.INIT('h2)
	) name17766 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][11]/P0001 ,
		_w21761_,
		_w21813_
	);
	LUT2 #(
		.INIT('h8)
	) name17767 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w21761_,
		_w21814_
	);
	LUT2 #(
		.INIT('h1)
	) name17768 (
		_w21813_,
		_w21814_,
		_w21815_
	);
	LUT2 #(
		.INIT('h2)
	) name17769 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][10]/P0001 ,
		_w21761_,
		_w21816_
	);
	LUT2 #(
		.INIT('h8)
	) name17770 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w21761_,
		_w21817_
	);
	LUT2 #(
		.INIT('h1)
	) name17771 (
		_w21816_,
		_w21817_,
		_w21818_
	);
	LUT2 #(
		.INIT('h2)
	) name17772 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][9]/P0001 ,
		_w20595_,
		_w21819_
	);
	LUT2 #(
		.INIT('h8)
	) name17773 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w20595_,
		_w21820_
	);
	LUT2 #(
		.INIT('h1)
	) name17774 (
		_w21819_,
		_w21820_,
		_w21821_
	);
	LUT2 #(
		.INIT('h2)
	) name17775 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][8]/P0001 ,
		_w20595_,
		_w21822_
	);
	LUT2 #(
		.INIT('h8)
	) name17776 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		_w20595_,
		_w21823_
	);
	LUT2 #(
		.INIT('h1)
	) name17777 (
		_w21822_,
		_w21823_,
		_w21824_
	);
	LUT2 #(
		.INIT('h2)
	) name17778 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][6]/P0001 ,
		_w20595_,
		_w21825_
	);
	LUT2 #(
		.INIT('h8)
	) name17779 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w20595_,
		_w21826_
	);
	LUT2 #(
		.INIT('h1)
	) name17780 (
		_w21825_,
		_w21826_,
		_w21827_
	);
	LUT2 #(
		.INIT('h2)
	) name17781 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][5]/P0001 ,
		_w20595_,
		_w21828_
	);
	LUT2 #(
		.INIT('h8)
	) name17782 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w20595_,
		_w21829_
	);
	LUT2 #(
		.INIT('h1)
	) name17783 (
		_w21828_,
		_w21829_,
		_w21830_
	);
	LUT2 #(
		.INIT('h2)
	) name17784 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][4]/P0001 ,
		_w20595_,
		_w21831_
	);
	LUT2 #(
		.INIT('h8)
	) name17785 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w20595_,
		_w21832_
	);
	LUT2 #(
		.INIT('h1)
	) name17786 (
		_w21831_,
		_w21832_,
		_w21833_
	);
	LUT2 #(
		.INIT('h2)
	) name17787 (
		_w13805_,
		_w21800_,
		_w21834_
	);
	LUT2 #(
		.INIT('h2)
	) name17788 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[10]/P0001 ,
		_w13805_,
		_w21835_
	);
	LUT2 #(
		.INIT('h1)
	) name17789 (
		_w21834_,
		_w21835_,
		_w21836_
	);
	LUT2 #(
		.INIT('h2)
	) name17790 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][21]/P0001 ,
		_w20595_,
		_w21837_
	);
	LUT2 #(
		.INIT('h8)
	) name17791 (
		\core_c_dec_IRE_reg[17]/NET0131 ,
		_w20595_,
		_w21838_
	);
	LUT2 #(
		.INIT('h1)
	) name17792 (
		_w21837_,
		_w21838_,
		_w21839_
	);
	LUT2 #(
		.INIT('h2)
	) name17793 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][20]/P0001 ,
		_w20595_,
		_w21840_
	);
	LUT2 #(
		.INIT('h8)
	) name17794 (
		\core_c_dec_IRE_reg[16]/NET0131 ,
		_w20595_,
		_w21841_
	);
	LUT2 #(
		.INIT('h1)
	) name17795 (
		_w21840_,
		_w21841_,
		_w21842_
	);
	LUT2 #(
		.INIT('h2)
	) name17796 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][19]/P0001 ,
		_w20595_,
		_w21843_
	);
	LUT2 #(
		.INIT('h8)
	) name17797 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w20595_,
		_w21844_
	);
	LUT2 #(
		.INIT('h1)
	) name17798 (
		_w21843_,
		_w21844_,
		_w21845_
	);
	LUT2 #(
		.INIT('h2)
	) name17799 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][18]/P0001 ,
		_w20595_,
		_w21846_
	);
	LUT2 #(
		.INIT('h8)
	) name17800 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		_w20595_,
		_w21847_
	);
	LUT2 #(
		.INIT('h1)
	) name17801 (
		_w21846_,
		_w21847_,
		_w21848_
	);
	LUT2 #(
		.INIT('h2)
	) name17802 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][17]/P0001 ,
		_w20595_,
		_w21849_
	);
	LUT2 #(
		.INIT('h8)
	) name17803 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w20595_,
		_w21850_
	);
	LUT2 #(
		.INIT('h1)
	) name17804 (
		_w21849_,
		_w21850_,
		_w21851_
	);
	LUT2 #(
		.INIT('h2)
	) name17805 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][15]/P0001 ,
		_w20595_,
		_w21852_
	);
	LUT2 #(
		.INIT('h8)
	) name17806 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w20595_,
		_w21853_
	);
	LUT2 #(
		.INIT('h1)
	) name17807 (
		_w21852_,
		_w21853_,
		_w21854_
	);
	LUT2 #(
		.INIT('h2)
	) name17808 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][14]/P0001 ,
		_w20595_,
		_w21855_
	);
	LUT2 #(
		.INIT('h8)
	) name17809 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		_w20595_,
		_w21856_
	);
	LUT2 #(
		.INIT('h1)
	) name17810 (
		_w21855_,
		_w21856_,
		_w21857_
	);
	LUT2 #(
		.INIT('h2)
	) name17811 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][13]/P0001 ,
		_w20595_,
		_w21858_
	);
	LUT2 #(
		.INIT('h8)
	) name17812 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w20595_,
		_w21859_
	);
	LUT2 #(
		.INIT('h1)
	) name17813 (
		_w21858_,
		_w21859_,
		_w21860_
	);
	LUT2 #(
		.INIT('h2)
	) name17814 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][12]/P0001 ,
		_w20595_,
		_w21861_
	);
	LUT2 #(
		.INIT('h8)
	) name17815 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w20595_,
		_w21862_
	);
	LUT2 #(
		.INIT('h1)
	) name17816 (
		_w21861_,
		_w21862_,
		_w21863_
	);
	LUT2 #(
		.INIT('h2)
	) name17817 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][11]/P0001 ,
		_w20595_,
		_w21864_
	);
	LUT2 #(
		.INIT('h8)
	) name17818 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w20595_,
		_w21865_
	);
	LUT2 #(
		.INIT('h1)
	) name17819 (
		_w21864_,
		_w21865_,
		_w21866_
	);
	LUT2 #(
		.INIT('h2)
	) name17820 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][10]/P0001 ,
		_w20595_,
		_w21867_
	);
	LUT2 #(
		.INIT('h8)
	) name17821 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w20595_,
		_w21868_
	);
	LUT2 #(
		.INIT('h1)
	) name17822 (
		_w21867_,
		_w21868_,
		_w21869_
	);
	LUT2 #(
		.INIT('h1)
	) name17823 (
		_w13789_,
		_w13794_,
		_w21870_
	);
	LUT2 #(
		.INIT('h8)
	) name17824 (
		_w13779_,
		_w21870_,
		_w21871_
	);
	LUT2 #(
		.INIT('h1)
	) name17825 (
		_w13778_,
		_w21870_,
		_w21872_
	);
	LUT2 #(
		.INIT('h1)
	) name17826 (
		_w21871_,
		_w21872_,
		_w21873_
	);
	LUT2 #(
		.INIT('h2)
	) name17827 (
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		_w4116_,
		_w21874_
	);
	LUT2 #(
		.INIT('h2)
	) name17828 (
		\core_c_psq_T_IRQE1_reg/P0001 ,
		\core_c_psq_T_IRQE1_s1_reg/P0001 ,
		_w21875_
	);
	LUT2 #(
		.INIT('h1)
	) name17829 (
		\core_c_psq_IFC_reg[12]/NET0131 ,
		\core_c_psq_Iflag_reg[4]/NET0131 ,
		_w21876_
	);
	LUT2 #(
		.INIT('h4)
	) name17830 (
		_w21875_,
		_w21876_,
		_w21877_
	);
	LUT2 #(
		.INIT('h1)
	) name17831 (
		\core_c_psq_IFC_reg[4]/NET0131 ,
		_w21877_,
		_w21878_
	);
	LUT2 #(
		.INIT('h4)
	) name17832 (
		_w21874_,
		_w21878_,
		_w21879_
	);
	LUT2 #(
		.INIT('h2)
	) name17833 (
		_w14711_,
		_w18220_,
		_w21880_
	);
	LUT2 #(
		.INIT('h1)
	) name17834 (
		\core_c_psq_SSTAT_reg[5]/NET0131 ,
		_w21880_,
		_w21881_
	);
	LUT2 #(
		.INIT('h2)
	) name17835 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][16]/P0001 ,
		_w20595_,
		_w21882_
	);
	LUT2 #(
		.INIT('h8)
	) name17836 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w20595_,
		_w21883_
	);
	LUT2 #(
		.INIT('h1)
	) name17837 (
		_w21882_,
		_w21883_,
		_w21884_
	);
	LUT2 #(
		.INIT('h2)
	) name17838 (
		\bdma_DM_2nd_reg/NET0131 ,
		_w13753_,
		_w21885_
	);
	LUT2 #(
		.INIT('h4)
	) name17839 (
		\bdma_DM_2nd_reg/NET0131 ,
		_w13753_,
		_w21886_
	);
	LUT2 #(
		.INIT('h1)
	) name17840 (
		_w21885_,
		_w21886_,
		_w21887_
	);
	LUT2 #(
		.INIT('h2)
	) name17841 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][7]/P0001 ,
		_w20595_,
		_w21888_
	);
	LUT2 #(
		.INIT('h8)
	) name17842 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w20595_,
		_w21889_
	);
	LUT2 #(
		.INIT('h1)
	) name17843 (
		_w21888_,
		_w21889_,
		_w21890_
	);
	LUT2 #(
		.INIT('h4)
	) name17844 (
		\memc_MMR_web_reg/NET0131 ,
		_w13762_,
		_w21891_
	);
	LUT2 #(
		.INIT('h8)
	) name17845 (
		_w18230_,
		_w21891_,
		_w21892_
	);
	LUT2 #(
		.INIT('h4)
	) name17846 (
		_w7340_,
		_w21892_,
		_w21893_
	);
	LUT2 #(
		.INIT('h1)
	) name17847 (
		\pio_pmask_reg_DO_reg[9]/NET0131 ,
		_w21892_,
		_w21894_
	);
	LUT2 #(
		.INIT('h1)
	) name17848 (
		_w21893_,
		_w21894_,
		_w21895_
	);
	LUT2 #(
		.INIT('h8)
	) name17849 (
		_w18228_,
		_w21891_,
		_w21896_
	);
	LUT2 #(
		.INIT('h4)
	) name17850 (
		_w9178_,
		_w21896_,
		_w21897_
	);
	LUT2 #(
		.INIT('h1)
	) name17851 (
		\PIO_oe[8]_pad ,
		_w21896_,
		_w21898_
	);
	LUT2 #(
		.INIT('h1)
	) name17852 (
		_w21897_,
		_w21898_,
		_w21899_
	);
	LUT2 #(
		.INIT('h2)
	) name17853 (
		_w17833_,
		_w21702_,
		_w21900_
	);
	LUT2 #(
		.INIT('h1)
	) name17854 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[3]/P0001 ,
		_w17833_,
		_w21901_
	);
	LUT2 #(
		.INIT('h1)
	) name17855 (
		_w21900_,
		_w21901_,
		_w21902_
	);
	LUT2 #(
		.INIT('h2)
	) name17856 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][13]/P0001 ,
		_w21761_,
		_w21903_
	);
	LUT2 #(
		.INIT('h8)
	) name17857 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		_w21761_,
		_w21904_
	);
	LUT2 #(
		.INIT('h1)
	) name17858 (
		_w21903_,
		_w21904_,
		_w21905_
	);
	LUT2 #(
		.INIT('h8)
	) name17859 (
		_w7526_,
		_w18227_,
		_w21906_
	);
	LUT2 #(
		.INIT('h4)
	) name17860 (
		_w10289_,
		_w21906_,
		_w21907_
	);
	LUT2 #(
		.INIT('h1)
	) name17861 (
		\memc_usysr_DO_reg[9]/NET0131 ,
		_w21906_,
		_w21908_
	);
	LUT2 #(
		.INIT('h1)
	) name17862 (
		_w21907_,
		_w21908_,
		_w21909_
	);
	LUT2 #(
		.INIT('h4)
	) name17863 (
		_w10638_,
		_w21906_,
		_w21910_
	);
	LUT2 #(
		.INIT('h1)
	) name17864 (
		\memc_usysr_DO_reg[8]/NET0131 ,
		_w21906_,
		_w21911_
	);
	LUT2 #(
		.INIT('h1)
	) name17865 (
		_w21910_,
		_w21911_,
		_w21912_
	);
	LUT2 #(
		.INIT('h4)
	) name17866 (
		_w7340_,
		_w21906_,
		_w21913_
	);
	LUT2 #(
		.INIT('h1)
	) name17867 (
		\memc_usysr_DO_reg[13]/NET0131 ,
		_w21906_,
		_w21914_
	);
	LUT2 #(
		.INIT('h1)
	) name17868 (
		_w21913_,
		_w21914_,
		_w21915_
	);
	LUT2 #(
		.INIT('h4)
	) name17869 (
		_w8460_,
		_w21906_,
		_w21916_
	);
	LUT2 #(
		.INIT('h1)
	) name17870 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w21906_,
		_w21917_
	);
	LUT2 #(
		.INIT('h1)
	) name17871 (
		_w21916_,
		_w21917_,
		_w21918_
	);
	LUT2 #(
		.INIT('h4)
	) name17872 (
		_w7859_,
		_w21906_,
		_w21919_
	);
	LUT2 #(
		.INIT('h1)
	) name17873 (
		\memc_usysr_DO_reg[10]/NET0131 ,
		_w21906_,
		_w21920_
	);
	LUT2 #(
		.INIT('h1)
	) name17874 (
		_w21919_,
		_w21920_,
		_w21921_
	);
	LUT2 #(
		.INIT('h8)
	) name17875 (
		_w7232_,
		_w18227_,
		_w21922_
	);
	LUT2 #(
		.INIT('h8)
	) name17876 (
		_w20070_,
		_w21922_,
		_w21923_
	);
	LUT2 #(
		.INIT('h4)
	) name17877 (
		_w10289_,
		_w21923_,
		_w21924_
	);
	LUT2 #(
		.INIT('h1)
	) name17878 (
		\sport1_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w21923_,
		_w21925_
	);
	LUT2 #(
		.INIT('h1)
	) name17879 (
		_w21924_,
		_w21925_,
		_w21926_
	);
	LUT2 #(
		.INIT('h4)
	) name17880 (
		_w10638_,
		_w21923_,
		_w21927_
	);
	LUT2 #(
		.INIT('h1)
	) name17881 (
		\sport1_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w21923_,
		_w21928_
	);
	LUT2 #(
		.INIT('h1)
	) name17882 (
		_w21927_,
		_w21928_,
		_w21929_
	);
	LUT2 #(
		.INIT('h2)
	) name17883 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w21663_,
		_w21930_
	);
	LUT2 #(
		.INIT('h1)
	) name17884 (
		_w18117_,
		_w18909_,
		_w21931_
	);
	LUT2 #(
		.INIT('h1)
	) name17885 (
		_w18079_,
		_w18991_,
		_w21932_
	);
	LUT2 #(
		.INIT('h2)
	) name17886 (
		_w17931_,
		_w21157_,
		_w21933_
	);
	LUT2 #(
		.INIT('h1)
	) name17887 (
		_w18104_,
		_w18912_,
		_w21934_
	);
	LUT2 #(
		.INIT('h2)
	) name17888 (
		_w18083_,
		_w18175_,
		_w21935_
	);
	LUT2 #(
		.INIT('h2)
	) name17889 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7987_,
		_w21936_
	);
	LUT2 #(
		.INIT('h8)
	) name17890 (
		_w17925_,
		_w17991_,
		_w21937_
	);
	LUT2 #(
		.INIT('h2)
	) name17891 (
		_w18748_,
		_w18888_,
		_w21938_
	);
	LUT2 #(
		.INIT('h2)
	) name17892 (
		_w18125_,
		_w18918_,
		_w21939_
	);
	LUT2 #(
		.INIT('h4)
	) name17893 (
		_w18082_,
		_w19720_,
		_w21940_
	);
	LUT2 #(
		.INIT('h4)
	) name17894 (
		_w17998_,
		_w18187_,
		_w21941_
	);
	LUT2 #(
		.INIT('h2)
	) name17895 (
		_w18183_,
		_w18898_,
		_w21942_
	);
	LUT2 #(
		.INIT('h2)
	) name17896 (
		_w18163_,
		_w18914_,
		_w21943_
	);
	LUT2 #(
		.INIT('h1)
	) name17897 (
		_w18026_,
		_w21936_,
		_w21944_
	);
	LUT2 #(
		.INIT('h4)
	) name17898 (
		_w21931_,
		_w21944_,
		_w21945_
	);
	LUT2 #(
		.INIT('h1)
	) name17899 (
		_w21932_,
		_w21934_,
		_w21946_
	);
	LUT2 #(
		.INIT('h1)
	) name17900 (
		_w21937_,
		_w21939_,
		_w21947_
	);
	LUT2 #(
		.INIT('h1)
	) name17901 (
		_w21940_,
		_w21943_,
		_w21948_
	);
	LUT2 #(
		.INIT('h8)
	) name17902 (
		_w21947_,
		_w21948_,
		_w21949_
	);
	LUT2 #(
		.INIT('h8)
	) name17903 (
		_w21945_,
		_w21946_,
		_w21950_
	);
	LUT2 #(
		.INIT('h2)
	) name17904 (
		_w18903_,
		_w21935_,
		_w21951_
	);
	LUT2 #(
		.INIT('h1)
	) name17905 (
		_w21938_,
		_w21941_,
		_w21952_
	);
	LUT2 #(
		.INIT('h4)
	) name17906 (
		_w21942_,
		_w21952_,
		_w21953_
	);
	LUT2 #(
		.INIT('h8)
	) name17907 (
		_w21950_,
		_w21951_,
		_w21954_
	);
	LUT2 #(
		.INIT('h8)
	) name17908 (
		_w18024_,
		_w21949_,
		_w21955_
	);
	LUT2 #(
		.INIT('h4)
	) name17909 (
		_w21933_,
		_w21955_,
		_w21956_
	);
	LUT2 #(
		.INIT('h8)
	) name17910 (
		_w21953_,
		_w21954_,
		_w21957_
	);
	LUT2 #(
		.INIT('h8)
	) name17911 (
		_w21956_,
		_w21957_,
		_w21958_
	);
	LUT2 #(
		.INIT('h4)
	) name17912 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w21958_,
		_w21959_
	);
	LUT2 #(
		.INIT('h1)
	) name17913 (
		_w21930_,
		_w21959_,
		_w21960_
	);
	LUT2 #(
		.INIT('h2)
	) name17914 (
		_w18886_,
		_w21960_,
		_w21961_
	);
	LUT2 #(
		.INIT('h1)
	) name17915 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[3]/P0001 ,
		_w18886_,
		_w21962_
	);
	LUT2 #(
		.INIT('h1)
	) name17916 (
		_w21961_,
		_w21962_,
		_w21963_
	);
	LUT2 #(
		.INIT('h4)
	) name17917 (
		_w7340_,
		_w21923_,
		_w21964_
	);
	LUT2 #(
		.INIT('h1)
	) name17918 (
		\sport1_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w21923_,
		_w21965_
	);
	LUT2 #(
		.INIT('h1)
	) name17919 (
		_w21964_,
		_w21965_,
		_w21966_
	);
	LUT2 #(
		.INIT('h4)
	) name17920 (
		_w9178_,
		_w21923_,
		_w21967_
	);
	LUT2 #(
		.INIT('h1)
	) name17921 (
		\sport1_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w21923_,
		_w21968_
	);
	LUT2 #(
		.INIT('h1)
	) name17922 (
		_w21967_,
		_w21968_,
		_w21969_
	);
	LUT2 #(
		.INIT('h4)
	) name17923 (
		_w8460_,
		_w21923_,
		_w21970_
	);
	LUT2 #(
		.INIT('h1)
	) name17924 (
		\sport1_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w21923_,
		_w21971_
	);
	LUT2 #(
		.INIT('h1)
	) name17925 (
		_w21970_,
		_w21971_,
		_w21972_
	);
	LUT2 #(
		.INIT('h4)
	) name17926 (
		_w7859_,
		_w21923_,
		_w21973_
	);
	LUT2 #(
		.INIT('h1)
	) name17927 (
		\sport1_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w21923_,
		_w21974_
	);
	LUT2 #(
		.INIT('h1)
	) name17928 (
		_w21973_,
		_w21974_,
		_w21975_
	);
	LUT2 #(
		.INIT('h8)
	) name17929 (
		_w7526_,
		_w21891_,
		_w21976_
	);
	LUT2 #(
		.INIT('h4)
	) name17930 (
		_w10638_,
		_w21976_,
		_w21977_
	);
	LUT2 #(
		.INIT('h1)
	) name17931 (
		\sport1_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w21976_,
		_w21978_
	);
	LUT2 #(
		.INIT('h1)
	) name17932 (
		_w21977_,
		_w21978_,
		_w21979_
	);
	LUT2 #(
		.INIT('h4)
	) name17933 (
		_w10289_,
		_w21976_,
		_w21980_
	);
	LUT2 #(
		.INIT('h1)
	) name17934 (
		\sport1_regs_AUTOreg_DO_reg[9]/NET0131 ,
		_w21976_,
		_w21981_
	);
	LUT2 #(
		.INIT('h1)
	) name17935 (
		_w21980_,
		_w21981_,
		_w21982_
	);
	LUT2 #(
		.INIT('h4)
	) name17936 (
		_w8460_,
		_w21976_,
		_w21983_
	);
	LUT2 #(
		.INIT('h1)
	) name17937 (
		\sport1_regs_AUTOreg_DO_reg[11]/NET0131 ,
		_w21976_,
		_w21984_
	);
	LUT2 #(
		.INIT('h1)
	) name17938 (
		_w21983_,
		_w21984_,
		_w21985_
	);
	LUT2 #(
		.INIT('h4)
	) name17939 (
		_w7859_,
		_w21976_,
		_w21986_
	);
	LUT2 #(
		.INIT('h1)
	) name17940 (
		\sport1_regs_AUTOreg_DO_reg[10]/NET0131 ,
		_w21976_,
		_w21987_
	);
	LUT2 #(
		.INIT('h1)
	) name17941 (
		_w21986_,
		_w21987_,
		_w21988_
	);
	LUT2 #(
		.INIT('h4)
	) name17942 (
		\core_c_dec_MTAY0_E_reg/P0001 ,
		_w13799_,
		_w21989_
	);
	LUT2 #(
		.INIT('h2)
	) name17943 (
		_w14665_,
		_w21989_,
		_w21990_
	);
	LUT2 #(
		.INIT('h1)
	) name17944 (
		\core_c_dec_Double_E_reg/P0001 ,
		\core_c_dec_accPM_E_reg/P0001 ,
		_w21991_
	);
	LUT2 #(
		.INIT('h4)
	) name17945 (
		_w10289_,
		_w21991_,
		_w21992_
	);
	LUT2 #(
		.INIT('h1)
	) name17946 (
		_w13075_,
		_w21991_,
		_w21993_
	);
	LUT2 #(
		.INIT('h1)
	) name17947 (
		_w21992_,
		_w21993_,
		_w21994_
	);
	LUT2 #(
		.INIT('h1)
	) name17948 (
		_w13806_,
		_w21994_,
		_w21995_
	);
	LUT2 #(
		.INIT('h8)
	) name17949 (
		_w10453_,
		_w13806_,
		_w21996_
	);
	LUT2 #(
		.INIT('h1)
	) name17950 (
		_w21995_,
		_w21996_,
		_w21997_
	);
	LUT2 #(
		.INIT('h2)
	) name17951 (
		_w21990_,
		_w21997_,
		_w21998_
	);
	LUT2 #(
		.INIT('h1)
	) name17952 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[9]/P0001 ,
		_w21990_,
		_w21999_
	);
	LUT2 #(
		.INIT('h1)
	) name17953 (
		_w21998_,
		_w21999_,
		_w22000_
	);
	LUT2 #(
		.INIT('h2)
	) name17954 (
		_w13041_,
		_w21991_,
		_w22001_
	);
	LUT2 #(
		.INIT('h8)
	) name17955 (
		_w10638_,
		_w21991_,
		_w22002_
	);
	LUT2 #(
		.INIT('h1)
	) name17956 (
		_w22001_,
		_w22002_,
		_w22003_
	);
	LUT2 #(
		.INIT('h4)
	) name17957 (
		_w13806_,
		_w22003_,
		_w22004_
	);
	LUT2 #(
		.INIT('h8)
	) name17958 (
		_w11054_,
		_w13806_,
		_w22005_
	);
	LUT2 #(
		.INIT('h1)
	) name17959 (
		_w22004_,
		_w22005_,
		_w22006_
	);
	LUT2 #(
		.INIT('h2)
	) name17960 (
		_w21990_,
		_w22006_,
		_w22007_
	);
	LUT2 #(
		.INIT('h1)
	) name17961 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[8]/P0001 ,
		_w21990_,
		_w22008_
	);
	LUT2 #(
		.INIT('h1)
	) name17962 (
		_w22007_,
		_w22008_,
		_w22009_
	);
	LUT2 #(
		.INIT('h4)
	) name17963 (
		_w11265_,
		_w21991_,
		_w22010_
	);
	LUT2 #(
		.INIT('h1)
	) name17964 (
		_w13006_,
		_w21991_,
		_w22011_
	);
	LUT2 #(
		.INIT('h1)
	) name17965 (
		_w22010_,
		_w22011_,
		_w22012_
	);
	LUT2 #(
		.INIT('h1)
	) name17966 (
		_w13806_,
		_w22012_,
		_w22013_
	);
	LUT2 #(
		.INIT('h8)
	) name17967 (
		_w11329_,
		_w13806_,
		_w22014_
	);
	LUT2 #(
		.INIT('h1)
	) name17968 (
		_w22013_,
		_w22014_,
		_w22015_
	);
	LUT2 #(
		.INIT('h2)
	) name17969 (
		_w21990_,
		_w22015_,
		_w22016_
	);
	LUT2 #(
		.INIT('h1)
	) name17970 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[7]/P0001 ,
		_w21990_,
		_w22017_
	);
	LUT2 #(
		.INIT('h1)
	) name17971 (
		_w22016_,
		_w22017_,
		_w22018_
	);
	LUT2 #(
		.INIT('h4)
	) name17972 (
		_w11525_,
		_w21991_,
		_w22019_
	);
	LUT2 #(
		.INIT('h1)
	) name17973 (
		_w12972_,
		_w21991_,
		_w22020_
	);
	LUT2 #(
		.INIT('h1)
	) name17974 (
		_w22019_,
		_w22020_,
		_w22021_
	);
	LUT2 #(
		.INIT('h1)
	) name17975 (
		_w13806_,
		_w22021_,
		_w22022_
	);
	LUT2 #(
		.INIT('h8)
	) name17976 (
		_w10686_,
		_w13806_,
		_w22023_
	);
	LUT2 #(
		.INIT('h1)
	) name17977 (
		_w22022_,
		_w22023_,
		_w22024_
	);
	LUT2 #(
		.INIT('h2)
	) name17978 (
		_w21990_,
		_w22024_,
		_w22025_
	);
	LUT2 #(
		.INIT('h1)
	) name17979 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[6]/P0001 ,
		_w21990_,
		_w22026_
	);
	LUT2 #(
		.INIT('h1)
	) name17980 (
		_w22025_,
		_w22026_,
		_w22027_
	);
	LUT2 #(
		.INIT('h4)
	) name17981 (
		_w10911_,
		_w21991_,
		_w22028_
	);
	LUT2 #(
		.INIT('h1)
	) name17982 (
		_w12938_,
		_w21991_,
		_w22029_
	);
	LUT2 #(
		.INIT('h1)
	) name17983 (
		_w22028_,
		_w22029_,
		_w22030_
	);
	LUT2 #(
		.INIT('h1)
	) name17984 (
		_w13806_,
		_w22030_,
		_w22031_
	);
	LUT2 #(
		.INIT('h8)
	) name17985 (
		_w9904_,
		_w13806_,
		_w22032_
	);
	LUT2 #(
		.INIT('h1)
	) name17986 (
		_w22031_,
		_w22032_,
		_w22033_
	);
	LUT2 #(
		.INIT('h2)
	) name17987 (
		_w21990_,
		_w22033_,
		_w22034_
	);
	LUT2 #(
		.INIT('h1)
	) name17988 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[5]/P0001 ,
		_w21990_,
		_w22035_
	);
	LUT2 #(
		.INIT('h1)
	) name17989 (
		_w22034_,
		_w22035_,
		_w22036_
	);
	LUT2 #(
		.INIT('h4)
	) name17990 (
		_w10069_,
		_w21991_,
		_w22037_
	);
	LUT2 #(
		.INIT('h1)
	) name17991 (
		_w12904_,
		_w21991_,
		_w22038_
	);
	LUT2 #(
		.INIT('h1)
	) name17992 (
		_w22037_,
		_w22038_,
		_w22039_
	);
	LUT2 #(
		.INIT('h1)
	) name17993 (
		_w13806_,
		_w22039_,
		_w22040_
	);
	LUT2 #(
		.INIT('h8)
	) name17994 (
		_w7944_,
		_w13806_,
		_w22041_
	);
	LUT2 #(
		.INIT('h1)
	) name17995 (
		_w22040_,
		_w22041_,
		_w22042_
	);
	LUT2 #(
		.INIT('h2)
	) name17996 (
		_w21990_,
		_w22042_,
		_w22043_
	);
	LUT2 #(
		.INIT('h1)
	) name17997 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[4]/P0001 ,
		_w21990_,
		_w22044_
	);
	LUT2 #(
		.INIT('h1)
	) name17998 (
		_w22043_,
		_w22044_,
		_w22045_
	);
	LUT2 #(
		.INIT('h4)
	) name17999 (
		_w8113_,
		_w21991_,
		_w22046_
	);
	LUT2 #(
		.INIT('h1)
	) name18000 (
		_w12870_,
		_w21991_,
		_w22047_
	);
	LUT2 #(
		.INIT('h1)
	) name18001 (
		_w22046_,
		_w22047_,
		_w22048_
	);
	LUT2 #(
		.INIT('h1)
	) name18002 (
		_w13806_,
		_w22048_,
		_w22049_
	);
	LUT2 #(
		.INIT('h8)
	) name18003 (
		_w8577_,
		_w13806_,
		_w22050_
	);
	LUT2 #(
		.INIT('h1)
	) name18004 (
		_w22049_,
		_w22050_,
		_w22051_
	);
	LUT2 #(
		.INIT('h2)
	) name18005 (
		_w21990_,
		_w22051_,
		_w22052_
	);
	LUT2 #(
		.INIT('h1)
	) name18006 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[3]/P0001 ,
		_w21990_,
		_w22053_
	);
	LUT2 #(
		.INIT('h1)
	) name18007 (
		_w22052_,
		_w22053_,
		_w22054_
	);
	LUT2 #(
		.INIT('h4)
	) name18008 (
		_w8715_,
		_w21991_,
		_w22055_
	);
	LUT2 #(
		.INIT('h1)
	) name18009 (
		_w12836_,
		_w21991_,
		_w22056_
	);
	LUT2 #(
		.INIT('h1)
	) name18010 (
		_w22055_,
		_w22056_,
		_w22057_
	);
	LUT2 #(
		.INIT('h1)
	) name18011 (
		_w13806_,
		_w22057_,
		_w22058_
	);
	LUT2 #(
		.INIT('h8)
	) name18012 (
		_w9305_,
		_w13806_,
		_w22059_
	);
	LUT2 #(
		.INIT('h1)
	) name18013 (
		_w22058_,
		_w22059_,
		_w22060_
	);
	LUT2 #(
		.INIT('h2)
	) name18014 (
		_w21990_,
		_w22060_,
		_w22061_
	);
	LUT2 #(
		.INIT('h1)
	) name18015 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[2]/P0001 ,
		_w21990_,
		_w22062_
	);
	LUT2 #(
		.INIT('h1)
	) name18016 (
		_w22061_,
		_w22062_,
		_w22063_
	);
	LUT2 #(
		.INIT('h4)
	) name18017 (
		_w12743_,
		_w21991_,
		_w22064_
	);
	LUT2 #(
		.INIT('h1)
	) name18018 (
		_w12771_,
		_w21991_,
		_w22065_
	);
	LUT2 #(
		.INIT('h1)
	) name18019 (
		_w22064_,
		_w22065_,
		_w22066_
	);
	LUT2 #(
		.INIT('h1)
	) name18020 (
		_w13806_,
		_w22066_,
		_w22067_
	);
	LUT2 #(
		.INIT('h8)
	) name18021 (
		_w11829_,
		_w13806_,
		_w22068_
	);
	LUT2 #(
		.INIT('h1)
	) name18022 (
		_w22067_,
		_w22068_,
		_w22069_
	);
	LUT2 #(
		.INIT('h2)
	) name18023 (
		_w21990_,
		_w22069_,
		_w22070_
	);
	LUT2 #(
		.INIT('h1)
	) name18024 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[15]/P0001 ,
		_w21990_,
		_w22071_
	);
	LUT2 #(
		.INIT('h1)
	) name18025 (
		_w22070_,
		_w22071_,
		_w22072_
	);
	LUT2 #(
		.INIT('h4)
	) name18026 (
		_w12688_,
		_w21991_,
		_w22073_
	);
	LUT2 #(
		.INIT('h1)
	) name18027 (
		_w12715_,
		_w21991_,
		_w22074_
	);
	LUT2 #(
		.INIT('h1)
	) name18028 (
		_w22073_,
		_w22074_,
		_w22075_
	);
	LUT2 #(
		.INIT('h1)
	) name18029 (
		_w13806_,
		_w22075_,
		_w22076_
	);
	LUT2 #(
		.INIT('h8)
	) name18030 (
		_w7104_,
		_w13806_,
		_w22077_
	);
	LUT2 #(
		.INIT('h1)
	) name18031 (
		_w22076_,
		_w22077_,
		_w22078_
	);
	LUT2 #(
		.INIT('h2)
	) name18032 (
		_w21990_,
		_w22078_,
		_w22079_
	);
	LUT2 #(
		.INIT('h1)
	) name18033 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[14]/P0001 ,
		_w21990_,
		_w22080_
	);
	LUT2 #(
		.INIT('h1)
	) name18034 (
		_w22079_,
		_w22080_,
		_w22081_
	);
	LUT2 #(
		.INIT('h4)
	) name18035 (
		_w7340_,
		_w21991_,
		_w22082_
	);
	LUT2 #(
		.INIT('h1)
	) name18036 (
		_w12658_,
		_w21991_,
		_w22083_
	);
	LUT2 #(
		.INIT('h1)
	) name18037 (
		_w22082_,
		_w22083_,
		_w22084_
	);
	LUT2 #(
		.INIT('h1)
	) name18038 (
		_w13806_,
		_w22084_,
		_w22085_
	);
	LUT2 #(
		.INIT('h8)
	) name18039 (
		_w9095_,
		_w13806_,
		_w22086_
	);
	LUT2 #(
		.INIT('h1)
	) name18040 (
		_w22085_,
		_w22086_,
		_w22087_
	);
	LUT2 #(
		.INIT('h2)
	) name18041 (
		_w21990_,
		_w22087_,
		_w22088_
	);
	LUT2 #(
		.INIT('h1)
	) name18042 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[13]/P0001 ,
		_w21990_,
		_w22089_
	);
	LUT2 #(
		.INIT('h1)
	) name18043 (
		_w22088_,
		_w22089_,
		_w22090_
	);
	LUT2 #(
		.INIT('h2)
	) name18044 (
		_w12624_,
		_w21991_,
		_w22091_
	);
	LUT2 #(
		.INIT('h8)
	) name18045 (
		_w9178_,
		_w21991_,
		_w22092_
	);
	LUT2 #(
		.INIT('h1)
	) name18046 (
		_w22091_,
		_w22092_,
		_w22093_
	);
	LUT2 #(
		.INIT('h4)
	) name18047 (
		_w13806_,
		_w22093_,
		_w22094_
	);
	LUT2 #(
		.INIT('h8)
	) name18048 (
		_w8377_,
		_w13806_,
		_w22095_
	);
	LUT2 #(
		.INIT('h1)
	) name18049 (
		_w22094_,
		_w22095_,
		_w22096_
	);
	LUT2 #(
		.INIT('h2)
	) name18050 (
		_w21990_,
		_w22096_,
		_w22097_
	);
	LUT2 #(
		.INIT('h1)
	) name18051 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[12]/P0001 ,
		_w21990_,
		_w22098_
	);
	LUT2 #(
		.INIT('h1)
	) name18052 (
		_w22097_,
		_w22098_,
		_w22099_
	);
	LUT2 #(
		.INIT('h2)
	) name18053 (
		_w19034_,
		_w21960_,
		_w22100_
	);
	LUT2 #(
		.INIT('h1)
	) name18054 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[3]/P0001 ,
		_w19034_,
		_w22101_
	);
	LUT2 #(
		.INIT('h1)
	) name18055 (
		_w22100_,
		_w22101_,
		_w22102_
	);
	LUT2 #(
		.INIT('h2)
	) name18056 (
		_w12590_,
		_w21991_,
		_w22103_
	);
	LUT2 #(
		.INIT('h8)
	) name18057 (
		_w8460_,
		_w21991_,
		_w22104_
	);
	LUT2 #(
		.INIT('h1)
	) name18058 (
		_w22103_,
		_w22104_,
		_w22105_
	);
	LUT2 #(
		.INIT('h4)
	) name18059 (
		_w13806_,
		_w22105_,
		_w22106_
	);
	LUT2 #(
		.INIT('h8)
	) name18060 (
		_w7776_,
		_w13806_,
		_w22107_
	);
	LUT2 #(
		.INIT('h1)
	) name18061 (
		_w22106_,
		_w22107_,
		_w22108_
	);
	LUT2 #(
		.INIT('h2)
	) name18062 (
		_w21990_,
		_w22108_,
		_w22109_
	);
	LUT2 #(
		.INIT('h1)
	) name18063 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[11]/P0001 ,
		_w21990_,
		_w22110_
	);
	LUT2 #(
		.INIT('h1)
	) name18064 (
		_w22109_,
		_w22110_,
		_w22111_
	);
	LUT2 #(
		.INIT('h4)
	) name18065 (
		_w7859_,
		_w21991_,
		_w22112_
	);
	LUT2 #(
		.INIT('h1)
	) name18066 (
		_w12556_,
		_w21991_,
		_w22113_
	);
	LUT2 #(
		.INIT('h1)
	) name18067 (
		_w22112_,
		_w22113_,
		_w22114_
	);
	LUT2 #(
		.INIT('h1)
	) name18068 (
		_w13806_,
		_w22114_,
		_w22115_
	);
	LUT2 #(
		.INIT('h8)
	) name18069 (
		_w10183_,
		_w13806_,
		_w22116_
	);
	LUT2 #(
		.INIT('h1)
	) name18070 (
		_w22115_,
		_w22116_,
		_w22117_
	);
	LUT2 #(
		.INIT('h2)
	) name18071 (
		_w21990_,
		_w22117_,
		_w22118_
	);
	LUT2 #(
		.INIT('h1)
	) name18072 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[10]/P0001 ,
		_w21990_,
		_w22119_
	);
	LUT2 #(
		.INIT('h1)
	) name18073 (
		_w22118_,
		_w22119_,
		_w22120_
	);
	LUT2 #(
		.INIT('h4)
	) name18074 (
		_w7340_,
		_w21896_,
		_w22121_
	);
	LUT2 #(
		.INIT('h1)
	) name18075 (
		\PIO_oe[9]_pad ,
		_w21896_,
		_w22122_
	);
	LUT2 #(
		.INIT('h1)
	) name18076 (
		_w22121_,
		_w22122_,
		_w22123_
	);
	LUT2 #(
		.INIT('h8)
	) name18077 (
		_w7283_,
		_w21922_,
		_w22124_
	);
	LUT2 #(
		.INIT('h4)
	) name18078 (
		_w10289_,
		_w22124_,
		_w22125_
	);
	LUT2 #(
		.INIT('h1)
	) name18079 (
		\sport0_regs_SCLKDIVreg_DO_reg[9]/NET0131 ,
		_w22124_,
		_w22126_
	);
	LUT2 #(
		.INIT('h1)
	) name18080 (
		_w22125_,
		_w22126_,
		_w22127_
	);
	LUT2 #(
		.INIT('h4)
	) name18081 (
		_w10638_,
		_w22124_,
		_w22128_
	);
	LUT2 #(
		.INIT('h1)
	) name18082 (
		\sport0_regs_SCLKDIVreg_DO_reg[8]/NET0131 ,
		_w22124_,
		_w22129_
	);
	LUT2 #(
		.INIT('h1)
	) name18083 (
		_w22128_,
		_w22129_,
		_w22130_
	);
	LUT2 #(
		.INIT('h4)
	) name18084 (
		_w7340_,
		_w22124_,
		_w22131_
	);
	LUT2 #(
		.INIT('h1)
	) name18085 (
		\sport0_regs_SCLKDIVreg_DO_reg[13]/NET0131 ,
		_w22124_,
		_w22132_
	);
	LUT2 #(
		.INIT('h1)
	) name18086 (
		_w22131_,
		_w22132_,
		_w22133_
	);
	LUT2 #(
		.INIT('h4)
	) name18087 (
		_w9178_,
		_w22124_,
		_w22134_
	);
	LUT2 #(
		.INIT('h1)
	) name18088 (
		\sport0_regs_SCLKDIVreg_DO_reg[12]/NET0131 ,
		_w22124_,
		_w22135_
	);
	LUT2 #(
		.INIT('h1)
	) name18089 (
		_w22134_,
		_w22135_,
		_w22136_
	);
	LUT2 #(
		.INIT('h4)
	) name18090 (
		_w8460_,
		_w22124_,
		_w22137_
	);
	LUT2 #(
		.INIT('h1)
	) name18091 (
		\sport0_regs_SCLKDIVreg_DO_reg[11]/NET0131 ,
		_w22124_,
		_w22138_
	);
	LUT2 #(
		.INIT('h1)
	) name18092 (
		_w22137_,
		_w22138_,
		_w22139_
	);
	LUT2 #(
		.INIT('h4)
	) name18093 (
		_w7859_,
		_w22124_,
		_w22140_
	);
	LUT2 #(
		.INIT('h1)
	) name18094 (
		\sport0_regs_SCLKDIVreg_DO_reg[10]/NET0131 ,
		_w22124_,
		_w22141_
	);
	LUT2 #(
		.INIT('h1)
	) name18095 (
		_w22140_,
		_w22141_,
		_w22142_
	);
	LUT2 #(
		.INIT('h4)
	) name18096 (
		_w9178_,
		_w21892_,
		_w22143_
	);
	LUT2 #(
		.INIT('h1)
	) name18097 (
		\pio_pmask_reg_DO_reg[8]/NET0131 ,
		_w21892_,
		_w22144_
	);
	LUT2 #(
		.INIT('h1)
	) name18098 (
		_w22143_,
		_w22144_,
		_w22145_
	);
	LUT2 #(
		.INIT('h4)
	) name18099 (
		_w9178_,
		_w20401_,
		_w22146_
	);
	LUT2 #(
		.INIT('h1)
	) name18100 (
		\sport0_regs_AUTO_a_reg[12]/NET0131 ,
		_w20401_,
		_w22147_
	);
	LUT2 #(
		.INIT('h1)
	) name18101 (
		_w22146_,
		_w22147_,
		_w22148_
	);
	LUT2 #(
		.INIT('h4)
	) name18102 (
		_w9435_,
		_w21991_,
		_w22149_
	);
	LUT2 #(
		.INIT('h1)
	) name18103 (
		_w12802_,
		_w21991_,
		_w22150_
	);
	LUT2 #(
		.INIT('h1)
	) name18104 (
		_w22149_,
		_w22150_,
		_w22151_
	);
	LUT2 #(
		.INIT('h4)
	) name18105 (
		_w13806_,
		_w22151_,
		_w22152_
	);
	LUT2 #(
		.INIT('h4)
	) name18106 (
		_w7414_,
		_w13806_,
		_w22153_
	);
	LUT2 #(
		.INIT('h1)
	) name18107 (
		_w22152_,
		_w22153_,
		_w22154_
	);
	LUT2 #(
		.INIT('h2)
	) name18108 (
		_w21990_,
		_w22154_,
		_w22155_
	);
	LUT2 #(
		.INIT('h2)
	) name18109 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[1]/P0001 ,
		_w21990_,
		_w22156_
	);
	LUT2 #(
		.INIT('h1)
	) name18110 (
		_w22155_,
		_w22156_,
		_w22157_
	);
	LUT2 #(
		.INIT('h2)
	) name18111 (
		_w17798_,
		_w21989_,
		_w22158_
	);
	LUT2 #(
		.INIT('h4)
	) name18112 (
		_w21997_,
		_w22158_,
		_w22159_
	);
	LUT2 #(
		.INIT('h1)
	) name18113 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[9]/P0001 ,
		_w22158_,
		_w22160_
	);
	LUT2 #(
		.INIT('h1)
	) name18114 (
		_w22159_,
		_w22160_,
		_w22161_
	);
	LUT2 #(
		.INIT('h4)
	) name18115 (
		_w22006_,
		_w22158_,
		_w22162_
	);
	LUT2 #(
		.INIT('h1)
	) name18116 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[8]/P0001 ,
		_w22158_,
		_w22163_
	);
	LUT2 #(
		.INIT('h1)
	) name18117 (
		_w22162_,
		_w22163_,
		_w22164_
	);
	LUT2 #(
		.INIT('h4)
	) name18118 (
		_w22015_,
		_w22158_,
		_w22165_
	);
	LUT2 #(
		.INIT('h1)
	) name18119 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[7]/P0001 ,
		_w22158_,
		_w22166_
	);
	LUT2 #(
		.INIT('h1)
	) name18120 (
		_w22165_,
		_w22166_,
		_w22167_
	);
	LUT2 #(
		.INIT('h4)
	) name18121 (
		_w22024_,
		_w22158_,
		_w22168_
	);
	LUT2 #(
		.INIT('h1)
	) name18122 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[6]/P0001 ,
		_w22158_,
		_w22169_
	);
	LUT2 #(
		.INIT('h1)
	) name18123 (
		_w22168_,
		_w22169_,
		_w22170_
	);
	LUT2 #(
		.INIT('h4)
	) name18124 (
		_w22033_,
		_w22158_,
		_w22171_
	);
	LUT2 #(
		.INIT('h1)
	) name18125 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[5]/P0001 ,
		_w22158_,
		_w22172_
	);
	LUT2 #(
		.INIT('h1)
	) name18126 (
		_w22171_,
		_w22172_,
		_w22173_
	);
	LUT2 #(
		.INIT('h4)
	) name18127 (
		_w22042_,
		_w22158_,
		_w22174_
	);
	LUT2 #(
		.INIT('h1)
	) name18128 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[4]/P0001 ,
		_w22158_,
		_w22175_
	);
	LUT2 #(
		.INIT('h1)
	) name18129 (
		_w22174_,
		_w22175_,
		_w22176_
	);
	LUT2 #(
		.INIT('h4)
	) name18130 (
		_w22051_,
		_w22158_,
		_w22177_
	);
	LUT2 #(
		.INIT('h1)
	) name18131 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[3]/P0001 ,
		_w22158_,
		_w22178_
	);
	LUT2 #(
		.INIT('h1)
	) name18132 (
		_w22177_,
		_w22178_,
		_w22179_
	);
	LUT2 #(
		.INIT('h4)
	) name18133 (
		_w22060_,
		_w22158_,
		_w22180_
	);
	LUT2 #(
		.INIT('h1)
	) name18134 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[2]/P0001 ,
		_w22158_,
		_w22181_
	);
	LUT2 #(
		.INIT('h1)
	) name18135 (
		_w22180_,
		_w22181_,
		_w22182_
	);
	LUT2 #(
		.INIT('h4)
	) name18136 (
		_w22154_,
		_w22158_,
		_w22183_
	);
	LUT2 #(
		.INIT('h2)
	) name18137 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[1]/P0001 ,
		_w22158_,
		_w22184_
	);
	LUT2 #(
		.INIT('h1)
	) name18138 (
		_w22183_,
		_w22184_,
		_w22185_
	);
	LUT2 #(
		.INIT('h4)
	) name18139 (
		_w22069_,
		_w22158_,
		_w22186_
	);
	LUT2 #(
		.INIT('h1)
	) name18140 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[15]/P0001 ,
		_w22158_,
		_w22187_
	);
	LUT2 #(
		.INIT('h1)
	) name18141 (
		_w22186_,
		_w22187_,
		_w22188_
	);
	LUT2 #(
		.INIT('h4)
	) name18142 (
		_w22078_,
		_w22158_,
		_w22189_
	);
	LUT2 #(
		.INIT('h1)
	) name18143 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[14]/P0001 ,
		_w22158_,
		_w22190_
	);
	LUT2 #(
		.INIT('h1)
	) name18144 (
		_w22189_,
		_w22190_,
		_w22191_
	);
	LUT2 #(
		.INIT('h4)
	) name18145 (
		_w22087_,
		_w22158_,
		_w22192_
	);
	LUT2 #(
		.INIT('h1)
	) name18146 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[13]/P0001 ,
		_w22158_,
		_w22193_
	);
	LUT2 #(
		.INIT('h1)
	) name18147 (
		_w22192_,
		_w22193_,
		_w22194_
	);
	LUT2 #(
		.INIT('h4)
	) name18148 (
		_w22096_,
		_w22158_,
		_w22195_
	);
	LUT2 #(
		.INIT('h1)
	) name18149 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[12]/P0001 ,
		_w22158_,
		_w22196_
	);
	LUT2 #(
		.INIT('h1)
	) name18150 (
		_w22195_,
		_w22196_,
		_w22197_
	);
	LUT2 #(
		.INIT('h4)
	) name18151 (
		_w22108_,
		_w22158_,
		_w22198_
	);
	LUT2 #(
		.INIT('h1)
	) name18152 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[11]/P0001 ,
		_w22158_,
		_w22199_
	);
	LUT2 #(
		.INIT('h1)
	) name18153 (
		_w22198_,
		_w22199_,
		_w22200_
	);
	LUT2 #(
		.INIT('h4)
	) name18154 (
		_w22117_,
		_w22158_,
		_w22201_
	);
	LUT2 #(
		.INIT('h1)
	) name18155 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[10]/P0001 ,
		_w22158_,
		_w22202_
	);
	LUT2 #(
		.INIT('h1)
	) name18156 (
		_w22201_,
		_w22202_,
		_w22203_
	);
	LUT2 #(
		.INIT('h4)
	) name18157 (
		_w12743_,
		_w22124_,
		_w22204_
	);
	LUT2 #(
		.INIT('h1)
	) name18158 (
		\sport0_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w22124_,
		_w22205_
	);
	LUT2 #(
		.INIT('h1)
	) name18159 (
		_w22204_,
		_w22205_,
		_w22206_
	);
	LUT2 #(
		.INIT('h4)
	) name18160 (
		_w8113_,
		_w22124_,
		_w22207_
	);
	LUT2 #(
		.INIT('h1)
	) name18161 (
		\sport0_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w22124_,
		_w22208_
	);
	LUT2 #(
		.INIT('h1)
	) name18162 (
		_w22207_,
		_w22208_,
		_w22209_
	);
	LUT2 #(
		.INIT('h4)
	) name18163 (
		_w10911_,
		_w22124_,
		_w22210_
	);
	LUT2 #(
		.INIT('h1)
	) name18164 (
		\sport0_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w22124_,
		_w22211_
	);
	LUT2 #(
		.INIT('h1)
	) name18165 (
		_w22210_,
		_w22211_,
		_w22212_
	);
	LUT2 #(
		.INIT('h4)
	) name18166 (
		_w12743_,
		_w20401_,
		_w22213_
	);
	LUT2 #(
		.INIT('h1)
	) name18167 (
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w20401_,
		_w22214_
	);
	LUT2 #(
		.INIT('h1)
	) name18168 (
		_w22213_,
		_w22214_,
		_w22215_
	);
	LUT2 #(
		.INIT('h4)
	) name18169 (
		_w11265_,
		_w21892_,
		_w22216_
	);
	LUT2 #(
		.INIT('h1)
	) name18170 (
		\pio_pmask_reg_DO_reg[7]/NET0131 ,
		_w21892_,
		_w22217_
	);
	LUT2 #(
		.INIT('h1)
	) name18171 (
		_w22216_,
		_w22217_,
		_w22218_
	);
	LUT2 #(
		.INIT('h4)
	) name18172 (
		_w11525_,
		_w21892_,
		_w22219_
	);
	LUT2 #(
		.INIT('h1)
	) name18173 (
		\pio_pmask_reg_DO_reg[6]/NET0131 ,
		_w21892_,
		_w22220_
	);
	LUT2 #(
		.INIT('h1)
	) name18174 (
		_w22219_,
		_w22220_,
		_w22221_
	);
	LUT2 #(
		.INIT('h4)
	) name18175 (
		_w8113_,
		_w21892_,
		_w22222_
	);
	LUT2 #(
		.INIT('h1)
	) name18176 (
		\pio_pmask_reg_DO_reg[3]/NET0131 ,
		_w21892_,
		_w22223_
	);
	LUT2 #(
		.INIT('h1)
	) name18177 (
		_w22222_,
		_w22223_,
		_w22224_
	);
	LUT2 #(
		.INIT('h4)
	) name18178 (
		_w12743_,
		_w21892_,
		_w22225_
	);
	LUT2 #(
		.INIT('h1)
	) name18179 (
		\pio_pmask_reg_DO_reg[11]/NET0131 ,
		_w21892_,
		_w22226_
	);
	LUT2 #(
		.INIT('h1)
	) name18180 (
		_w22225_,
		_w22226_,
		_w22227_
	);
	LUT2 #(
		.INIT('h1)
	) name18181 (
		\sice_ICYC_reg[18]/NET0131 ,
		_w20747_,
		_w22228_
	);
	LUT2 #(
		.INIT('h1)
	) name18182 (
		_w20748_,
		_w22228_,
		_w22229_
	);
	LUT2 #(
		.INIT('h4)
	) name18183 (
		_w8715_,
		_w21892_,
		_w22230_
	);
	LUT2 #(
		.INIT('h1)
	) name18184 (
		\pio_pmask_reg_DO_reg[2]/NET0131 ,
		_w21892_,
		_w22231_
	);
	LUT2 #(
		.INIT('h1)
	) name18185 (
		_w22230_,
		_w22231_,
		_w22232_
	);
	LUT2 #(
		.INIT('h4)
	) name18186 (
		_w7607_,
		_w21892_,
		_w22233_
	);
	LUT2 #(
		.INIT('h1)
	) name18187 (
		\pio_pmask_reg_DO_reg[0]/NET0131 ,
		_w21892_,
		_w22234_
	);
	LUT2 #(
		.INIT('h1)
	) name18188 (
		_w22233_,
		_w22234_,
		_w22235_
	);
	LUT2 #(
		.INIT('h4)
	) name18189 (
		_w11265_,
		_w21896_,
		_w22236_
	);
	LUT2 #(
		.INIT('h1)
	) name18190 (
		\PIO_oe[7]_pad ,
		_w21896_,
		_w22237_
	);
	LUT2 #(
		.INIT('h1)
	) name18191 (
		_w22236_,
		_w22237_,
		_w22238_
	);
	LUT2 #(
		.INIT('h4)
	) name18192 (
		_w11525_,
		_w21896_,
		_w22239_
	);
	LUT2 #(
		.INIT('h1)
	) name18193 (
		\PIO_oe[6]_pad ,
		_w21896_,
		_w22240_
	);
	LUT2 #(
		.INIT('h1)
	) name18194 (
		_w22239_,
		_w22240_,
		_w22241_
	);
	LUT2 #(
		.INIT('h4)
	) name18195 (
		_w10069_,
		_w21896_,
		_w22242_
	);
	LUT2 #(
		.INIT('h1)
	) name18196 (
		\PIO_oe[4]_pad ,
		_w21896_,
		_w22243_
	);
	LUT2 #(
		.INIT('h1)
	) name18197 (
		_w22242_,
		_w22243_,
		_w22244_
	);
	LUT2 #(
		.INIT('h4)
	) name18198 (
		_w8715_,
		_w21896_,
		_w22245_
	);
	LUT2 #(
		.INIT('h1)
	) name18199 (
		\PIO_oe[2]_pad ,
		_w21896_,
		_w22246_
	);
	LUT2 #(
		.INIT('h1)
	) name18200 (
		_w22245_,
		_w22246_,
		_w22247_
	);
	LUT2 #(
		.INIT('h4)
	) name18201 (
		_w9435_,
		_w21896_,
		_w22248_
	);
	LUT2 #(
		.INIT('h1)
	) name18202 (
		\PIO_oe[1]_pad ,
		_w21896_,
		_w22249_
	);
	LUT2 #(
		.INIT('h1)
	) name18203 (
		_w22248_,
		_w22249_,
		_w22250_
	);
	LUT2 #(
		.INIT('h4)
	) name18204 (
		_w12743_,
		_w21896_,
		_w22251_
	);
	LUT2 #(
		.INIT('h1)
	) name18205 (
		\PIO_oe[11]_pad ,
		_w21896_,
		_w22252_
	);
	LUT2 #(
		.INIT('h1)
	) name18206 (
		_w22251_,
		_w22252_,
		_w22253_
	);
	LUT2 #(
		.INIT('h4)
	) name18207 (
		_w11265_,
		_w21906_,
		_w22254_
	);
	LUT2 #(
		.INIT('h1)
	) name18208 (
		\memc_usysr_DO_reg[7]/NET0131 ,
		_w21906_,
		_w22255_
	);
	LUT2 #(
		.INIT('h1)
	) name18209 (
		_w22254_,
		_w22255_,
		_w22256_
	);
	LUT2 #(
		.INIT('h4)
	) name18210 (
		_w12688_,
		_w21892_,
		_w22257_
	);
	LUT2 #(
		.INIT('h1)
	) name18211 (
		\pio_pmask_reg_DO_reg[10]/NET0131 ,
		_w21892_,
		_w22258_
	);
	LUT2 #(
		.INIT('h1)
	) name18212 (
		_w22257_,
		_w22258_,
		_w22259_
	);
	LUT2 #(
		.INIT('h4)
	) name18213 (
		_w10911_,
		_w21892_,
		_w22260_
	);
	LUT2 #(
		.INIT('h1)
	) name18214 (
		\pio_pmask_reg_DO_reg[5]/NET0131 ,
		_w21892_,
		_w22261_
	);
	LUT2 #(
		.INIT('h1)
	) name18215 (
		_w22260_,
		_w22261_,
		_w22262_
	);
	LUT2 #(
		.INIT('h4)
	) name18216 (
		_w10911_,
		_w21906_,
		_w22263_
	);
	LUT2 #(
		.INIT('h1)
	) name18217 (
		\memc_usysr_DO_reg[5]/NET0131 ,
		_w21906_,
		_w22264_
	);
	LUT2 #(
		.INIT('h1)
	) name18218 (
		_w22263_,
		_w22264_,
		_w22265_
	);
	LUT2 #(
		.INIT('h4)
	) name18219 (
		_w11525_,
		_w21906_,
		_w22266_
	);
	LUT2 #(
		.INIT('h1)
	) name18220 (
		\memc_usysr_DO_reg[6]/NET0131 ,
		_w21906_,
		_w22267_
	);
	LUT2 #(
		.INIT('h1)
	) name18221 (
		_w22266_,
		_w22267_,
		_w22268_
	);
	LUT2 #(
		.INIT('h4)
	) name18222 (
		_w10069_,
		_w21906_,
		_w22269_
	);
	LUT2 #(
		.INIT('h1)
	) name18223 (
		\memc_usysr_DO_reg[4]/NET0131 ,
		_w21906_,
		_w22270_
	);
	LUT2 #(
		.INIT('h1)
	) name18224 (
		_w22269_,
		_w22270_,
		_w22271_
	);
	LUT2 #(
		.INIT('h4)
	) name18225 (
		_w8715_,
		_w21906_,
		_w22272_
	);
	LUT2 #(
		.INIT('h1)
	) name18226 (
		\memc_usysr_DO_reg[2]/NET0131 ,
		_w21906_,
		_w22273_
	);
	LUT2 #(
		.INIT('h1)
	) name18227 (
		_w22272_,
		_w22273_,
		_w22274_
	);
	LUT2 #(
		.INIT('h4)
	) name18228 (
		_w9435_,
		_w21906_,
		_w22275_
	);
	LUT2 #(
		.INIT('h1)
	) name18229 (
		\memc_usysr_DO_reg[1]/NET0131 ,
		_w21906_,
		_w22276_
	);
	LUT2 #(
		.INIT('h1)
	) name18230 (
		_w22275_,
		_w22276_,
		_w22277_
	);
	LUT2 #(
		.INIT('h4)
	) name18231 (
		_w12743_,
		_w21906_,
		_w22278_
	);
	LUT2 #(
		.INIT('h1)
	) name18232 (
		\memc_usysr_DO_reg[15]/NET0131 ,
		_w21906_,
		_w22279_
	);
	LUT2 #(
		.INIT('h1)
	) name18233 (
		_w22278_,
		_w22279_,
		_w22280_
	);
	LUT2 #(
		.INIT('h4)
	) name18234 (
		_w12688_,
		_w21906_,
		_w22281_
	);
	LUT2 #(
		.INIT('h1)
	) name18235 (
		\memc_usysr_DO_reg[14]/NET0131 ,
		_w21906_,
		_w22282_
	);
	LUT2 #(
		.INIT('h1)
	) name18236 (
		_w22281_,
		_w22282_,
		_w22283_
	);
	LUT2 #(
		.INIT('h4)
	) name18237 (
		_w7607_,
		_w21906_,
		_w22284_
	);
	LUT2 #(
		.INIT('h1)
	) name18238 (
		\memc_usysr_DO_reg[0]/NET0131 ,
		_w21906_,
		_w22285_
	);
	LUT2 #(
		.INIT('h1)
	) name18239 (
		_w22284_,
		_w22285_,
		_w22286_
	);
	LUT2 #(
		.INIT('h8)
	) name18240 (
		\idma_RDcyc_reg/NET0131 ,
		_w20393_,
		_w22287_
	);
	LUT2 #(
		.INIT('h1)
	) name18241 (
		_w20821_,
		_w22287_,
		_w22288_
	);
	LUT2 #(
		.INIT('h8)
	) name18242 (
		_w7261_,
		_w7525_,
		_w22289_
	);
	LUT2 #(
		.INIT('h8)
	) name18243 (
		_w18226_,
		_w22289_,
		_w22290_
	);
	LUT2 #(
		.INIT('h4)
	) name18244 (
		\memc_MMR_web_reg/NET0131 ,
		_w22290_,
		_w22291_
	);
	LUT2 #(
		.INIT('h4)
	) name18245 (
		_w8460_,
		_w22291_,
		_w22292_
	);
	LUT2 #(
		.INIT('h1)
	) name18246 (
		\tm_tcr_reg_DO_reg[11]/NET0131 ,
		_w22291_,
		_w22293_
	);
	LUT2 #(
		.INIT('h1)
	) name18247 (
		_w22292_,
		_w22293_,
		_w22294_
	);
	LUT2 #(
		.INIT('h4)
	) name18248 (
		_w8113_,
		_w21896_,
		_w22295_
	);
	LUT2 #(
		.INIT('h1)
	) name18249 (
		\PIO_oe[3]_pad ,
		_w21896_,
		_w22296_
	);
	LUT2 #(
		.INIT('h1)
	) name18250 (
		_w22295_,
		_w22296_,
		_w22297_
	);
	LUT2 #(
		.INIT('h8)
	) name18251 (
		_w7513_,
		_w21891_,
		_w22298_
	);
	LUT2 #(
		.INIT('h4)
	) name18252 (
		_w11265_,
		_w22298_,
		_w22299_
	);
	LUT2 #(
		.INIT('h1)
	) name18253 (
		\emc_WSCRext_reg_DO_reg[7]/NET0131 ,
		_w22298_,
		_w22300_
	);
	LUT2 #(
		.INIT('h1)
	) name18254 (
		_w22299_,
		_w22300_,
		_w22301_
	);
	LUT2 #(
		.INIT('h4)
	) name18255 (
		_w11525_,
		_w22298_,
		_w22302_
	);
	LUT2 #(
		.INIT('h1)
	) name18256 (
		\emc_WSCRext_reg_DO_reg[6]/NET0131 ,
		_w22298_,
		_w22303_
	);
	LUT2 #(
		.INIT('h1)
	) name18257 (
		_w22302_,
		_w22303_,
		_w22304_
	);
	LUT2 #(
		.INIT('h4)
	) name18258 (
		_w10911_,
		_w22298_,
		_w22305_
	);
	LUT2 #(
		.INIT('h1)
	) name18259 (
		\emc_WSCRext_reg_DO_reg[5]/NET0131 ,
		_w22298_,
		_w22306_
	);
	LUT2 #(
		.INIT('h1)
	) name18260 (
		_w22305_,
		_w22306_,
		_w22307_
	);
	LUT2 #(
		.INIT('h4)
	) name18261 (
		_w10069_,
		_w22298_,
		_w22308_
	);
	LUT2 #(
		.INIT('h1)
	) name18262 (
		\emc_WSCRext_reg_DO_reg[4]/NET0131 ,
		_w22298_,
		_w22309_
	);
	LUT2 #(
		.INIT('h1)
	) name18263 (
		_w22308_,
		_w22309_,
		_w22310_
	);
	LUT2 #(
		.INIT('h4)
	) name18264 (
		_w8113_,
		_w22298_,
		_w22311_
	);
	LUT2 #(
		.INIT('h1)
	) name18265 (
		\emc_WSCRext_reg_DO_reg[3]/NET0131 ,
		_w22298_,
		_w22312_
	);
	LUT2 #(
		.INIT('h1)
	) name18266 (
		_w22311_,
		_w22312_,
		_w22313_
	);
	LUT2 #(
		.INIT('h4)
	) name18267 (
		_w8715_,
		_w22298_,
		_w22314_
	);
	LUT2 #(
		.INIT('h1)
	) name18268 (
		\emc_WSCRext_reg_DO_reg[2]/NET0131 ,
		_w22298_,
		_w22315_
	);
	LUT2 #(
		.INIT('h1)
	) name18269 (
		_w22314_,
		_w22315_,
		_w22316_
	);
	LUT2 #(
		.INIT('h4)
	) name18270 (
		_w9435_,
		_w22298_,
		_w22317_
	);
	LUT2 #(
		.INIT('h1)
	) name18271 (
		\emc_WSCRext_reg_DO_reg[1]/NET0131 ,
		_w22298_,
		_w22318_
	);
	LUT2 #(
		.INIT('h1)
	) name18272 (
		_w22317_,
		_w22318_,
		_w22319_
	);
	LUT2 #(
		.INIT('h4)
	) name18273 (
		_w7607_,
		_w22298_,
		_w22320_
	);
	LUT2 #(
		.INIT('h1)
	) name18274 (
		\emc_WSCRext_reg_DO_reg[0]/NET0131 ,
		_w22298_,
		_w22321_
	);
	LUT2 #(
		.INIT('h1)
	) name18275 (
		_w22320_,
		_w22321_,
		_w22322_
	);
	LUT2 #(
		.INIT('h4)
	) name18276 (
		_w11265_,
		_w21923_,
		_w22323_
	);
	LUT2 #(
		.INIT('h1)
	) name18277 (
		\sport1_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w21923_,
		_w22324_
	);
	LUT2 #(
		.INIT('h1)
	) name18278 (
		_w22323_,
		_w22324_,
		_w22325_
	);
	LUT2 #(
		.INIT('h4)
	) name18279 (
		_w11525_,
		_w21923_,
		_w22326_
	);
	LUT2 #(
		.INIT('h1)
	) name18280 (
		\sport1_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w21923_,
		_w22327_
	);
	LUT2 #(
		.INIT('h1)
	) name18281 (
		_w22326_,
		_w22327_,
		_w22328_
	);
	LUT2 #(
		.INIT('h4)
	) name18282 (
		_w10911_,
		_w21923_,
		_w22329_
	);
	LUT2 #(
		.INIT('h1)
	) name18283 (
		\sport1_regs_SCLKDIVreg_DO_reg[5]/NET0131 ,
		_w21923_,
		_w22330_
	);
	LUT2 #(
		.INIT('h1)
	) name18284 (
		_w22329_,
		_w22330_,
		_w22331_
	);
	LUT2 #(
		.INIT('h4)
	) name18285 (
		_w10069_,
		_w21923_,
		_w22332_
	);
	LUT2 #(
		.INIT('h1)
	) name18286 (
		\sport1_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w21923_,
		_w22333_
	);
	LUT2 #(
		.INIT('h1)
	) name18287 (
		_w22332_,
		_w22333_,
		_w22334_
	);
	LUT2 #(
		.INIT('h4)
	) name18288 (
		_w8113_,
		_w21923_,
		_w22335_
	);
	LUT2 #(
		.INIT('h1)
	) name18289 (
		\sport1_regs_SCLKDIVreg_DO_reg[3]/NET0131 ,
		_w21923_,
		_w22336_
	);
	LUT2 #(
		.INIT('h1)
	) name18290 (
		_w22335_,
		_w22336_,
		_w22337_
	);
	LUT2 #(
		.INIT('h4)
	) name18291 (
		_w8715_,
		_w21923_,
		_w22338_
	);
	LUT2 #(
		.INIT('h1)
	) name18292 (
		\sport1_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w21923_,
		_w22339_
	);
	LUT2 #(
		.INIT('h1)
	) name18293 (
		_w22338_,
		_w22339_,
		_w22340_
	);
	LUT2 #(
		.INIT('h4)
	) name18294 (
		_w9435_,
		_w21923_,
		_w22341_
	);
	LUT2 #(
		.INIT('h1)
	) name18295 (
		\sport1_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w21923_,
		_w22342_
	);
	LUT2 #(
		.INIT('h1)
	) name18296 (
		_w22341_,
		_w22342_,
		_w22343_
	);
	LUT2 #(
		.INIT('h4)
	) name18297 (
		_w12743_,
		_w21923_,
		_w22344_
	);
	LUT2 #(
		.INIT('h1)
	) name18298 (
		\sport1_regs_SCLKDIVreg_DO_reg[15]/NET0131 ,
		_w21923_,
		_w22345_
	);
	LUT2 #(
		.INIT('h1)
	) name18299 (
		_w22344_,
		_w22345_,
		_w22346_
	);
	LUT2 #(
		.INIT('h4)
	) name18300 (
		_w12688_,
		_w21923_,
		_w22347_
	);
	LUT2 #(
		.INIT('h1)
	) name18301 (
		\sport1_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w21923_,
		_w22348_
	);
	LUT2 #(
		.INIT('h1)
	) name18302 (
		_w22347_,
		_w22348_,
		_w22349_
	);
	LUT2 #(
		.INIT('h4)
	) name18303 (
		_w7607_,
		_w21923_,
		_w22350_
	);
	LUT2 #(
		.INIT('h1)
	) name18304 (
		\sport1_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w21923_,
		_w22351_
	);
	LUT2 #(
		.INIT('h1)
	) name18305 (
		_w22350_,
		_w22351_,
		_w22352_
	);
	LUT2 #(
		.INIT('h4)
	) name18306 (
		_w11265_,
		_w21976_,
		_w22353_
	);
	LUT2 #(
		.INIT('h1)
	) name18307 (
		\sport1_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w21976_,
		_w22354_
	);
	LUT2 #(
		.INIT('h1)
	) name18308 (
		_w22353_,
		_w22354_,
		_w22355_
	);
	LUT2 #(
		.INIT('h4)
	) name18309 (
		_w11525_,
		_w21976_,
		_w22356_
	);
	LUT2 #(
		.INIT('h1)
	) name18310 (
		\sport1_regs_AUTOreg_DO_reg[6]/NET0131 ,
		_w21976_,
		_w22357_
	);
	LUT2 #(
		.INIT('h1)
	) name18311 (
		_w22356_,
		_w22357_,
		_w22358_
	);
	LUT2 #(
		.INIT('h4)
	) name18312 (
		_w10911_,
		_w21976_,
		_w22359_
	);
	LUT2 #(
		.INIT('h1)
	) name18313 (
		\sport1_regs_AUTOreg_DO_reg[5]/NET0131 ,
		_w21976_,
		_w22360_
	);
	LUT2 #(
		.INIT('h1)
	) name18314 (
		_w22359_,
		_w22360_,
		_w22361_
	);
	LUT2 #(
		.INIT('h4)
	) name18315 (
		_w10069_,
		_w21976_,
		_w22362_
	);
	LUT2 #(
		.INIT('h1)
	) name18316 (
		\sport1_regs_AUTOreg_DO_reg[4]/NET0131 ,
		_w21976_,
		_w22363_
	);
	LUT2 #(
		.INIT('h1)
	) name18317 (
		_w22362_,
		_w22363_,
		_w22364_
	);
	LUT2 #(
		.INIT('h4)
	) name18318 (
		_w8113_,
		_w21976_,
		_w22365_
	);
	LUT2 #(
		.INIT('h1)
	) name18319 (
		\sport1_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w21976_,
		_w22366_
	);
	LUT2 #(
		.INIT('h1)
	) name18320 (
		_w22365_,
		_w22366_,
		_w22367_
	);
	LUT2 #(
		.INIT('h4)
	) name18321 (
		_w8715_,
		_w21976_,
		_w22368_
	);
	LUT2 #(
		.INIT('h1)
	) name18322 (
		\sport1_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w21976_,
		_w22369_
	);
	LUT2 #(
		.INIT('h1)
	) name18323 (
		_w22368_,
		_w22369_,
		_w22370_
	);
	LUT2 #(
		.INIT('h4)
	) name18324 (
		_w9435_,
		_w21976_,
		_w22371_
	);
	LUT2 #(
		.INIT('h1)
	) name18325 (
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w21976_,
		_w22372_
	);
	LUT2 #(
		.INIT('h1)
	) name18326 (
		_w22371_,
		_w22372_,
		_w22373_
	);
	LUT2 #(
		.INIT('h4)
	) name18327 (
		_w7607_,
		_w21976_,
		_w22374_
	);
	LUT2 #(
		.INIT('h1)
	) name18328 (
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w21976_,
		_w22375_
	);
	LUT2 #(
		.INIT('h1)
	) name18329 (
		_w22374_,
		_w22375_,
		_w22376_
	);
	LUT2 #(
		.INIT('h4)
	) name18330 (
		_w10911_,
		_w21896_,
		_w22377_
	);
	LUT2 #(
		.INIT('h1)
	) name18331 (
		\PIO_oe[5]_pad ,
		_w21896_,
		_w22378_
	);
	LUT2 #(
		.INIT('h1)
	) name18332 (
		_w22377_,
		_w22378_,
		_w22379_
	);
	LUT2 #(
		.INIT('h4)
	) name18333 (
		_w10069_,
		_w21892_,
		_w22380_
	);
	LUT2 #(
		.INIT('h1)
	) name18334 (
		\pio_pmask_reg_DO_reg[4]/NET0131 ,
		_w21892_,
		_w22381_
	);
	LUT2 #(
		.INIT('h1)
	) name18335 (
		_w22380_,
		_w22381_,
		_w22382_
	);
	LUT2 #(
		.INIT('h4)
	) name18336 (
		_w7607_,
		_w21896_,
		_w22383_
	);
	LUT2 #(
		.INIT('h1)
	) name18337 (
		\PIO_oe[0]_pad ,
		_w21896_,
		_w22384_
	);
	LUT2 #(
		.INIT('h1)
	) name18338 (
		_w22383_,
		_w22384_,
		_w22385_
	);
	LUT2 #(
		.INIT('h2)
	) name18339 (
		\sport0_regs_AUTO_a_reg[14]/NET0131 ,
		_w20401_,
		_w22386_
	);
	LUT2 #(
		.INIT('h8)
	) name18340 (
		_w18235_,
		_w20400_,
		_w22387_
	);
	LUT2 #(
		.INIT('h1)
	) name18341 (
		_w22386_,
		_w22387_,
		_w22388_
	);
	LUT2 #(
		.INIT('h4)
	) name18342 (
		_w9435_,
		_w21892_,
		_w22389_
	);
	LUT2 #(
		.INIT('h1)
	) name18343 (
		\pio_pmask_reg_DO_reg[1]/NET0131 ,
		_w21892_,
		_w22390_
	);
	LUT2 #(
		.INIT('h1)
	) name18344 (
		_w22389_,
		_w22390_,
		_w22391_
	);
	LUT2 #(
		.INIT('h4)
	) name18345 (
		_w8113_,
		_w21906_,
		_w22392_
	);
	LUT2 #(
		.INIT('h1)
	) name18346 (
		\memc_usysr_DO_reg[3]/NET0131 ,
		_w21906_,
		_w22393_
	);
	LUT2 #(
		.INIT('h1)
	) name18347 (
		_w22392_,
		_w22393_,
		_w22394_
	);
	LUT2 #(
		.INIT('h4)
	) name18348 (
		_w12688_,
		_w21896_,
		_w22395_
	);
	LUT2 #(
		.INIT('h1)
	) name18349 (
		\PIO_oe[10]_pad ,
		_w21896_,
		_w22396_
	);
	LUT2 #(
		.INIT('h1)
	) name18350 (
		_w22395_,
		_w22396_,
		_w22397_
	);
	LUT2 #(
		.INIT('h8)
	) name18351 (
		\tm_tcr_reg_DO_reg[10]/NET0131 ,
		_w20355_,
		_w22398_
	);
	LUT2 #(
		.INIT('h4)
	) name18352 (
		\T_TMODE[0]_pad ,
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w22399_
	);
	LUT2 #(
		.INIT('h8)
	) name18353 (
		_w20372_,
		_w22399_,
		_w22400_
	);
	LUT2 #(
		.INIT('h4)
	) name18354 (
		\tm_tpr_reg_DO_reg[10]/NET0131 ,
		_w22400_,
		_w22401_
	);
	LUT2 #(
		.INIT('h1)
	) name18355 (
		\tm_TSR_TMP_reg[1]/NET0131 ,
		\tm_TSR_TMP_reg[2]/NET0131 ,
		_w22402_
	);
	LUT2 #(
		.INIT('h1)
	) name18356 (
		\tm_TSR_TMP_reg[0]/NET0131 ,
		\tm_TSR_TMP_reg[3]/NET0131 ,
		_w22403_
	);
	LUT2 #(
		.INIT('h8)
	) name18357 (
		_w22402_,
		_w22403_,
		_w22404_
	);
	LUT2 #(
		.INIT('h1)
	) name18358 (
		\tm_TSR_TMP_reg[4]/NET0131 ,
		\tm_TSR_TMP_reg[5]/NET0131 ,
		_w22405_
	);
	LUT2 #(
		.INIT('h1)
	) name18359 (
		\tm_TSR_TMP_reg[6]/NET0131 ,
		\tm_TSR_TMP_reg[7]/NET0131 ,
		_w22406_
	);
	LUT2 #(
		.INIT('h8)
	) name18360 (
		_w22405_,
		_w22406_,
		_w22407_
	);
	LUT2 #(
		.INIT('h8)
	) name18361 (
		_w22404_,
		_w22407_,
		_w22408_
	);
	LUT2 #(
		.INIT('h8)
	) name18362 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w22408_,
		_w22409_
	);
	LUT2 #(
		.INIT('h1)
	) name18363 (
		\T_TMODE[0]_pad ,
		_w22409_,
		_w22410_
	);
	LUT2 #(
		.INIT('h1)
	) name18364 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w22410_,
		_w22411_
	);
	LUT2 #(
		.INIT('h1)
	) name18365 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		_w22411_,
		_w22412_
	);
	LUT2 #(
		.INIT('h1)
	) name18366 (
		\T_TMODE[0]_pad ,
		_w20364_,
		_w22413_
	);
	LUT2 #(
		.INIT('h8)
	) name18367 (
		\tm_TCR_TMP_reg[8]/NET0131 ,
		_w22413_,
		_w22414_
	);
	LUT2 #(
		.INIT('h8)
	) name18368 (
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w22414_,
		_w22415_
	);
	LUT2 #(
		.INIT('h1)
	) name18369 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		_w22415_,
		_w22416_
	);
	LUT2 #(
		.INIT('h8)
	) name18370 (
		\tm_TCR_TMP_reg[10]/NET0131 ,
		_w22415_,
		_w22417_
	);
	LUT2 #(
		.INIT('h1)
	) name18371 (
		_w22416_,
		_w22417_,
		_w22418_
	);
	LUT2 #(
		.INIT('h1)
	) name18372 (
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w22414_,
		_w22419_
	);
	LUT2 #(
		.INIT('h1)
	) name18373 (
		_w22415_,
		_w22419_,
		_w22420_
	);
	LUT2 #(
		.INIT('h1)
	) name18374 (
		\tm_TCR_TMP_reg[8]/NET0131 ,
		_w22413_,
		_w22421_
	);
	LUT2 #(
		.INIT('h1)
	) name18375 (
		_w22414_,
		_w22421_,
		_w22422_
	);
	LUT2 #(
		.INIT('h1)
	) name18376 (
		_w22420_,
		_w22422_,
		_w22423_
	);
	LUT2 #(
		.INIT('h4)
	) name18377 (
		_w22418_,
		_w22423_,
		_w22424_
	);
	LUT2 #(
		.INIT('h2)
	) name18378 (
		_w22418_,
		_w22423_,
		_w22425_
	);
	LUT2 #(
		.INIT('h2)
	) name18379 (
		_w22411_,
		_w22424_,
		_w22426_
	);
	LUT2 #(
		.INIT('h4)
	) name18380 (
		_w22425_,
		_w22426_,
		_w22427_
	);
	LUT2 #(
		.INIT('h1)
	) name18381 (
		_w22412_,
		_w22427_,
		_w22428_
	);
	LUT2 #(
		.INIT('h1)
	) name18382 (
		_w22400_,
		_w22428_,
		_w22429_
	);
	LUT2 #(
		.INIT('h1)
	) name18383 (
		_w20355_,
		_w22401_,
		_w22430_
	);
	LUT2 #(
		.INIT('h4)
	) name18384 (
		_w22429_,
		_w22430_,
		_w22431_
	);
	LUT2 #(
		.INIT('h1)
	) name18385 (
		_w22398_,
		_w22431_,
		_w22432_
	);
	LUT2 #(
		.INIT('h4)
	) name18386 (
		_w11265_,
		_w22124_,
		_w22433_
	);
	LUT2 #(
		.INIT('h1)
	) name18387 (
		\sport0_regs_SCLKDIVreg_DO_reg[7]/NET0131 ,
		_w22124_,
		_w22434_
	);
	LUT2 #(
		.INIT('h1)
	) name18388 (
		_w22433_,
		_w22434_,
		_w22435_
	);
	LUT2 #(
		.INIT('h4)
	) name18389 (
		_w11525_,
		_w22124_,
		_w22436_
	);
	LUT2 #(
		.INIT('h1)
	) name18390 (
		\sport0_regs_SCLKDIVreg_DO_reg[6]/NET0131 ,
		_w22124_,
		_w22437_
	);
	LUT2 #(
		.INIT('h1)
	) name18391 (
		_w22436_,
		_w22437_,
		_w22438_
	);
	LUT2 #(
		.INIT('h4)
	) name18392 (
		_w10069_,
		_w22124_,
		_w22439_
	);
	LUT2 #(
		.INIT('h1)
	) name18393 (
		\sport0_regs_SCLKDIVreg_DO_reg[4]/NET0131 ,
		_w22124_,
		_w22440_
	);
	LUT2 #(
		.INIT('h1)
	) name18394 (
		_w22439_,
		_w22440_,
		_w22441_
	);
	LUT2 #(
		.INIT('h4)
	) name18395 (
		_w8715_,
		_w22124_,
		_w22442_
	);
	LUT2 #(
		.INIT('h1)
	) name18396 (
		\sport0_regs_SCLKDIVreg_DO_reg[2]/NET0131 ,
		_w22124_,
		_w22443_
	);
	LUT2 #(
		.INIT('h1)
	) name18397 (
		_w22442_,
		_w22443_,
		_w22444_
	);
	LUT2 #(
		.INIT('h4)
	) name18398 (
		_w9435_,
		_w22124_,
		_w22445_
	);
	LUT2 #(
		.INIT('h1)
	) name18399 (
		\sport0_regs_SCLKDIVreg_DO_reg[1]/NET0131 ,
		_w22124_,
		_w22446_
	);
	LUT2 #(
		.INIT('h1)
	) name18400 (
		_w22445_,
		_w22446_,
		_w22447_
	);
	LUT2 #(
		.INIT('h4)
	) name18401 (
		_w12688_,
		_w22124_,
		_w22448_
	);
	LUT2 #(
		.INIT('h1)
	) name18402 (
		\sport0_regs_SCLKDIVreg_DO_reg[14]/NET0131 ,
		_w22124_,
		_w22449_
	);
	LUT2 #(
		.INIT('h1)
	) name18403 (
		_w22448_,
		_w22449_,
		_w22450_
	);
	LUT2 #(
		.INIT('h4)
	) name18404 (
		_w7607_,
		_w22124_,
		_w22451_
	);
	LUT2 #(
		.INIT('h1)
	) name18405 (
		\sport0_regs_SCLKDIVreg_DO_reg[0]/NET0131 ,
		_w22124_,
		_w22452_
	);
	LUT2 #(
		.INIT('h1)
	) name18406 (
		_w22451_,
		_w22452_,
		_w22453_
	);
	LUT2 #(
		.INIT('h2)
	) name18407 (
		\core_c_psq_Iact_E_reg[8]/NET0131 ,
		_w19477_,
		_w22454_
	);
	LUT2 #(
		.INIT('h8)
	) name18408 (
		_w19484_,
		_w19486_,
		_w22455_
	);
	LUT2 #(
		.INIT('h1)
	) name18409 (
		_w22454_,
		_w22455_,
		_w22456_
	);
	LUT2 #(
		.INIT('h8)
	) name18410 (
		_w7237_,
		_w18227_,
		_w22457_
	);
	LUT2 #(
		.INIT('h8)
	) name18411 (
		_w7269_,
		_w22457_,
		_w22458_
	);
	LUT2 #(
		.INIT('h4)
	) name18412 (
		_w10289_,
		_w22458_,
		_w22459_
	);
	LUT2 #(
		.INIT('h1)
	) name18413 (
		\clkc_ckr_reg_DO_reg[9]/NET0131 ,
		_w22458_,
		_w22460_
	);
	LUT2 #(
		.INIT('h1)
	) name18414 (
		_w22459_,
		_w22460_,
		_w22461_
	);
	LUT2 #(
		.INIT('h4)
	) name18415 (
		_w10638_,
		_w22458_,
		_w22462_
	);
	LUT2 #(
		.INIT('h1)
	) name18416 (
		\clkc_ckr_reg_DO_reg[8]/NET0131 ,
		_w22458_,
		_w22463_
	);
	LUT2 #(
		.INIT('h1)
	) name18417 (
		_w22462_,
		_w22463_,
		_w22464_
	);
	LUT2 #(
		.INIT('h4)
	) name18418 (
		_w7340_,
		_w22458_,
		_w22465_
	);
	LUT2 #(
		.INIT('h1)
	) name18419 (
		\clkc_ckr_reg_DO_reg[13]/NET0131 ,
		_w22458_,
		_w22466_
	);
	LUT2 #(
		.INIT('h1)
	) name18420 (
		_w22465_,
		_w22466_,
		_w22467_
	);
	LUT2 #(
		.INIT('h4)
	) name18421 (
		_w9178_,
		_w22458_,
		_w22468_
	);
	LUT2 #(
		.INIT('h1)
	) name18422 (
		\clkc_ckr_reg_DO_reg[12]/NET0131 ,
		_w22458_,
		_w22469_
	);
	LUT2 #(
		.INIT('h1)
	) name18423 (
		_w22468_,
		_w22469_,
		_w22470_
	);
	LUT2 #(
		.INIT('h4)
	) name18424 (
		_w7859_,
		_w22458_,
		_w22471_
	);
	LUT2 #(
		.INIT('h1)
	) name18425 (
		\clkc_ckr_reg_DO_reg[10]/NET0131 ,
		_w22458_,
		_w22472_
	);
	LUT2 #(
		.INIT('h1)
	) name18426 (
		_w22471_,
		_w22472_,
		_w22473_
	);
	LUT2 #(
		.INIT('h4)
	) name18427 (
		_w8460_,
		_w22458_,
		_w22474_
	);
	LUT2 #(
		.INIT('h1)
	) name18428 (
		\clkc_ckr_reg_DO_reg[11]/NET0131 ,
		_w22458_,
		_w22475_
	);
	LUT2 #(
		.INIT('h1)
	) name18429 (
		_w22474_,
		_w22475_,
		_w22476_
	);
	LUT2 #(
		.INIT('h8)
	) name18430 (
		_w7525_,
		_w21922_,
		_w22477_
	);
	LUT2 #(
		.INIT('h4)
	) name18431 (
		_w8460_,
		_w22477_,
		_w22478_
	);
	LUT2 #(
		.INIT('h1)
	) name18432 (
		\tm_tpr_reg_DO_reg[11]/NET0131 ,
		_w22477_,
		_w22479_
	);
	LUT2 #(
		.INIT('h1)
	) name18433 (
		_w22478_,
		_w22479_,
		_w22480_
	);
	LUT2 #(
		.INIT('h4)
	) name18434 (
		_w7859_,
		_w22477_,
		_w22481_
	);
	LUT2 #(
		.INIT('h1)
	) name18435 (
		\tm_tpr_reg_DO_reg[10]/NET0131 ,
		_w22477_,
		_w22482_
	);
	LUT2 #(
		.INIT('h1)
	) name18436 (
		_w22481_,
		_w22482_,
		_w22483_
	);
	LUT2 #(
		.INIT('h8)
	) name18437 (
		_w7525_,
		_w22457_,
		_w22484_
	);
	LUT2 #(
		.INIT('h4)
	) name18438 (
		_w10289_,
		_w22484_,
		_w22485_
	);
	LUT2 #(
		.INIT('h1)
	) name18439 (
		\emc_WSCRreg_DO_reg[9]/NET0131 ,
		_w22484_,
		_w22486_
	);
	LUT2 #(
		.INIT('h1)
	) name18440 (
		_w22485_,
		_w22486_,
		_w22487_
	);
	LUT2 #(
		.INIT('h4)
	) name18441 (
		_w10638_,
		_w22484_,
		_w22488_
	);
	LUT2 #(
		.INIT('h1)
	) name18442 (
		\emc_WSCRreg_DO_reg[8]/NET0131 ,
		_w22484_,
		_w22489_
	);
	LUT2 #(
		.INIT('h1)
	) name18443 (
		_w22488_,
		_w22489_,
		_w22490_
	);
	LUT2 #(
		.INIT('h4)
	) name18444 (
		_w7340_,
		_w22484_,
		_w22491_
	);
	LUT2 #(
		.INIT('h1)
	) name18445 (
		\emc_WSCRreg_DO_reg[13]/NET0131 ,
		_w22484_,
		_w22492_
	);
	LUT2 #(
		.INIT('h1)
	) name18446 (
		_w22491_,
		_w22492_,
		_w22493_
	);
	LUT2 #(
		.INIT('h4)
	) name18447 (
		_w9178_,
		_w22484_,
		_w22494_
	);
	LUT2 #(
		.INIT('h1)
	) name18448 (
		\emc_WSCRreg_DO_reg[12]/NET0131 ,
		_w22484_,
		_w22495_
	);
	LUT2 #(
		.INIT('h1)
	) name18449 (
		_w22494_,
		_w22495_,
		_w22496_
	);
	LUT2 #(
		.INIT('h4)
	) name18450 (
		_w8460_,
		_w22484_,
		_w22497_
	);
	LUT2 #(
		.INIT('h1)
	) name18451 (
		\emc_WSCRreg_DO_reg[11]/NET0131 ,
		_w22484_,
		_w22498_
	);
	LUT2 #(
		.INIT('h1)
	) name18452 (
		_w22497_,
		_w22498_,
		_w22499_
	);
	LUT2 #(
		.INIT('h4)
	) name18453 (
		_w7859_,
		_w22484_,
		_w22500_
	);
	LUT2 #(
		.INIT('h1)
	) name18454 (
		\emc_WSCRreg_DO_reg[10]/NET0131 ,
		_w22484_,
		_w22501_
	);
	LUT2 #(
		.INIT('h1)
	) name18455 (
		_w22500_,
		_w22501_,
		_w22502_
	);
	LUT2 #(
		.INIT('h1)
	) name18456 (
		\sice_ICYC_reg[10]/NET0131 ,
		_w20739_,
		_w22503_
	);
	LUT2 #(
		.INIT('h1)
	) name18457 (
		_w20740_,
		_w22503_,
		_w22504_
	);
	LUT2 #(
		.INIT('h1)
	) name18458 (
		\sice_IIRC_reg[10]/NET0131 ,
		_w20854_,
		_w22505_
	);
	LUT2 #(
		.INIT('h1)
	) name18459 (
		_w20855_,
		_w22505_,
		_w22506_
	);
	LUT2 #(
		.INIT('h2)
	) name18460 (
		\emc_PMDreg_reg[7]/P0001 ,
		_w14745_,
		_w22507_
	);
	LUT2 #(
		.INIT('h8)
	) name18461 (
		\T_ED[7]_pad ,
		_w14745_,
		_w22508_
	);
	LUT2 #(
		.INIT('h1)
	) name18462 (
		_w22507_,
		_w22508_,
		_w22509_
	);
	LUT2 #(
		.INIT('h2)
	) name18463 (
		\emc_PMDreg_reg[6]/P0001 ,
		_w14745_,
		_w22510_
	);
	LUT2 #(
		.INIT('h8)
	) name18464 (
		\T_ED[6]_pad ,
		_w14745_,
		_w22511_
	);
	LUT2 #(
		.INIT('h1)
	) name18465 (
		_w22510_,
		_w22511_,
		_w22512_
	);
	LUT2 #(
		.INIT('h2)
	) name18466 (
		\emc_PMDreg_reg[5]/P0001 ,
		_w14745_,
		_w22513_
	);
	LUT2 #(
		.INIT('h8)
	) name18467 (
		\T_ED[5]_pad ,
		_w14745_,
		_w22514_
	);
	LUT2 #(
		.INIT('h1)
	) name18468 (
		_w22513_,
		_w22514_,
		_w22515_
	);
	LUT2 #(
		.INIT('h2)
	) name18469 (
		\emc_PMDreg_reg[4]/P0001 ,
		_w14745_,
		_w22516_
	);
	LUT2 #(
		.INIT('h8)
	) name18470 (
		\T_ED[4]_pad ,
		_w14745_,
		_w22517_
	);
	LUT2 #(
		.INIT('h1)
	) name18471 (
		_w22516_,
		_w22517_,
		_w22518_
	);
	LUT2 #(
		.INIT('h2)
	) name18472 (
		\emc_PMDreg_reg[3]/P0001 ,
		_w14745_,
		_w22519_
	);
	LUT2 #(
		.INIT('h8)
	) name18473 (
		\T_ED[3]_pad ,
		_w14745_,
		_w22520_
	);
	LUT2 #(
		.INIT('h1)
	) name18474 (
		_w22519_,
		_w22520_,
		_w22521_
	);
	LUT2 #(
		.INIT('h2)
	) name18475 (
		\emc_PMDreg_reg[2]/P0001 ,
		_w14745_,
		_w22522_
	);
	LUT2 #(
		.INIT('h8)
	) name18476 (
		\T_ED[2]_pad ,
		_w14745_,
		_w22523_
	);
	LUT2 #(
		.INIT('h1)
	) name18477 (
		_w22522_,
		_w22523_,
		_w22524_
	);
	LUT2 #(
		.INIT('h2)
	) name18478 (
		\emc_PMDreg_reg[1]/P0001 ,
		_w14745_,
		_w22525_
	);
	LUT2 #(
		.INIT('h8)
	) name18479 (
		\T_ED[1]_pad ,
		_w14745_,
		_w22526_
	);
	LUT2 #(
		.INIT('h1)
	) name18480 (
		_w22525_,
		_w22526_,
		_w22527_
	);
	LUT2 #(
		.INIT('h2)
	) name18481 (
		\emc_PMDreg_reg[15]/P0001 ,
		_w14745_,
		_w22528_
	);
	LUT2 #(
		.INIT('h8)
	) name18482 (
		\T_ED[15]_pad ,
		_w14745_,
		_w22529_
	);
	LUT2 #(
		.INIT('h1)
	) name18483 (
		_w22528_,
		_w22529_,
		_w22530_
	);
	LUT2 #(
		.INIT('h2)
	) name18484 (
		\emc_PMDreg_reg[14]/P0001 ,
		_w14745_,
		_w22531_
	);
	LUT2 #(
		.INIT('h8)
	) name18485 (
		\T_ED[14]_pad ,
		_w14745_,
		_w22532_
	);
	LUT2 #(
		.INIT('h1)
	) name18486 (
		_w22531_,
		_w22532_,
		_w22533_
	);
	LUT2 #(
		.INIT('h2)
	) name18487 (
		\emc_PMDreg_reg[13]/P0001 ,
		_w14745_,
		_w22534_
	);
	LUT2 #(
		.INIT('h8)
	) name18488 (
		\T_ED[13]_pad ,
		_w14745_,
		_w22535_
	);
	LUT2 #(
		.INIT('h1)
	) name18489 (
		_w22534_,
		_w22535_,
		_w22536_
	);
	LUT2 #(
		.INIT('h2)
	) name18490 (
		\emc_PMDreg_reg[12]/P0001 ,
		_w14745_,
		_w22537_
	);
	LUT2 #(
		.INIT('h8)
	) name18491 (
		\T_ED[12]_pad ,
		_w14745_,
		_w22538_
	);
	LUT2 #(
		.INIT('h1)
	) name18492 (
		_w22537_,
		_w22538_,
		_w22539_
	);
	LUT2 #(
		.INIT('h2)
	) name18493 (
		\emc_PMDreg_reg[11]/P0001 ,
		_w14745_,
		_w22540_
	);
	LUT2 #(
		.INIT('h8)
	) name18494 (
		\T_ED[11]_pad ,
		_w14745_,
		_w22541_
	);
	LUT2 #(
		.INIT('h1)
	) name18495 (
		_w22540_,
		_w22541_,
		_w22542_
	);
	LUT2 #(
		.INIT('h2)
	) name18496 (
		\emc_PMDreg_reg[10]/P0001 ,
		_w14745_,
		_w22543_
	);
	LUT2 #(
		.INIT('h8)
	) name18497 (
		\T_ED[10]_pad ,
		_w14745_,
		_w22544_
	);
	LUT2 #(
		.INIT('h1)
	) name18498 (
		_w22543_,
		_w22544_,
		_w22545_
	);
	LUT2 #(
		.INIT('h2)
	) name18499 (
		\emc_PMDreg_reg[0]/P0001 ,
		_w14745_,
		_w22546_
	);
	LUT2 #(
		.INIT('h8)
	) name18500 (
		\T_ED[0]_pad ,
		_w14745_,
		_w22547_
	);
	LUT2 #(
		.INIT('h1)
	) name18501 (
		_w22546_,
		_w22547_,
		_w22548_
	);
	LUT2 #(
		.INIT('h4)
	) name18502 (
		_w11265_,
		_w22458_,
		_w22549_
	);
	LUT2 #(
		.INIT('h1)
	) name18503 (
		\clkc_ckr_reg_DO_reg[7]/NET0131 ,
		_w22458_,
		_w22550_
	);
	LUT2 #(
		.INIT('h1)
	) name18504 (
		_w22549_,
		_w22550_,
		_w22551_
	);
	LUT2 #(
		.INIT('h4)
	) name18505 (
		_w11525_,
		_w22458_,
		_w22552_
	);
	LUT2 #(
		.INIT('h1)
	) name18506 (
		\clkc_ckr_reg_DO_reg[6]/NET0131 ,
		_w22458_,
		_w22553_
	);
	LUT2 #(
		.INIT('h1)
	) name18507 (
		_w22552_,
		_w22553_,
		_w22554_
	);
	LUT2 #(
		.INIT('h4)
	) name18508 (
		_w10911_,
		_w22458_,
		_w22555_
	);
	LUT2 #(
		.INIT('h1)
	) name18509 (
		\clkc_ckr_reg_DO_reg[5]/NET0131 ,
		_w22458_,
		_w22556_
	);
	LUT2 #(
		.INIT('h1)
	) name18510 (
		_w22555_,
		_w22556_,
		_w22557_
	);
	LUT2 #(
		.INIT('h4)
	) name18511 (
		_w10069_,
		_w22458_,
		_w22558_
	);
	LUT2 #(
		.INIT('h1)
	) name18512 (
		\clkc_ckr_reg_DO_reg[4]/NET0131 ,
		_w22458_,
		_w22559_
	);
	LUT2 #(
		.INIT('h1)
	) name18513 (
		_w22558_,
		_w22559_,
		_w22560_
	);
	LUT2 #(
		.INIT('h4)
	) name18514 (
		_w8113_,
		_w22458_,
		_w22561_
	);
	LUT2 #(
		.INIT('h1)
	) name18515 (
		\clkc_ckr_reg_DO_reg[3]/NET0131 ,
		_w22458_,
		_w22562_
	);
	LUT2 #(
		.INIT('h1)
	) name18516 (
		_w22561_,
		_w22562_,
		_w22563_
	);
	LUT2 #(
		.INIT('h4)
	) name18517 (
		_w8715_,
		_w22458_,
		_w22564_
	);
	LUT2 #(
		.INIT('h1)
	) name18518 (
		\clkc_ckr_reg_DO_reg[2]/NET0131 ,
		_w22458_,
		_w22565_
	);
	LUT2 #(
		.INIT('h1)
	) name18519 (
		_w22564_,
		_w22565_,
		_w22566_
	);
	LUT2 #(
		.INIT('h4)
	) name18520 (
		_w9435_,
		_w22458_,
		_w22567_
	);
	LUT2 #(
		.INIT('h1)
	) name18521 (
		\clkc_ckr_reg_DO_reg[1]/NET0131 ,
		_w22458_,
		_w22568_
	);
	LUT2 #(
		.INIT('h1)
	) name18522 (
		_w22567_,
		_w22568_,
		_w22569_
	);
	LUT2 #(
		.INIT('h4)
	) name18523 (
		_w12743_,
		_w22458_,
		_w22570_
	);
	LUT2 #(
		.INIT('h1)
	) name18524 (
		\clkc_ckr_reg_DO_reg[15]/NET0131 ,
		_w22458_,
		_w22571_
	);
	LUT2 #(
		.INIT('h1)
	) name18525 (
		_w22570_,
		_w22571_,
		_w22572_
	);
	LUT2 #(
		.INIT('h4)
	) name18526 (
		_w12688_,
		_w22458_,
		_w22573_
	);
	LUT2 #(
		.INIT('h1)
	) name18527 (
		\clkc_ckr_reg_DO_reg[14]/NET0131 ,
		_w22458_,
		_w22574_
	);
	LUT2 #(
		.INIT('h1)
	) name18528 (
		_w22573_,
		_w22574_,
		_w22575_
	);
	LUT2 #(
		.INIT('h4)
	) name18529 (
		_w7607_,
		_w22458_,
		_w22576_
	);
	LUT2 #(
		.INIT('h1)
	) name18530 (
		\clkc_ckr_reg_DO_reg[0]/NET0131 ,
		_w22458_,
		_w22577_
	);
	LUT2 #(
		.INIT('h1)
	) name18531 (
		_w22576_,
		_w22577_,
		_w22578_
	);
	LUT2 #(
		.INIT('h1)
	) name18532 (
		\sice_ICYC_reg[17]/NET0131 ,
		_w20746_,
		_w22579_
	);
	LUT2 #(
		.INIT('h1)
	) name18533 (
		_w20747_,
		_w22579_,
		_w22580_
	);
	LUT2 #(
		.INIT('h8)
	) name18534 (
		\sice_IIRC_reg[15]/NET0131 ,
		_w20859_,
		_w22581_
	);
	LUT2 #(
		.INIT('h8)
	) name18535 (
		\sice_IIRC_reg[16]/NET0131 ,
		_w22581_,
		_w22582_
	);
	LUT2 #(
		.INIT('h1)
	) name18536 (
		\sice_IIRC_reg[17]/NET0131 ,
		_w22582_,
		_w22583_
	);
	LUT2 #(
		.INIT('h8)
	) name18537 (
		\sice_IIRC_reg[17]/NET0131 ,
		_w22582_,
		_w22584_
	);
	LUT2 #(
		.INIT('h1)
	) name18538 (
		_w22583_,
		_w22584_,
		_w22585_
	);
	LUT2 #(
		.INIT('h1)
	) name18539 (
		\sice_IIRC_reg[13]/NET0131 ,
		_w20857_,
		_w22586_
	);
	LUT2 #(
		.INIT('h1)
	) name18540 (
		_w20858_,
		_w22586_,
		_w22587_
	);
	LUT2 #(
		.INIT('h1)
	) name18541 (
		\sice_ICYC_reg[13]/NET0131 ,
		_w20742_,
		_w22588_
	);
	LUT2 #(
		.INIT('h1)
	) name18542 (
		_w20743_,
		_w22588_,
		_w22589_
	);
	LUT2 #(
		.INIT('h4)
	) name18543 (
		_w11265_,
		_w22477_,
		_w22590_
	);
	LUT2 #(
		.INIT('h1)
	) name18544 (
		\tm_tpr_reg_DO_reg[7]/NET0131 ,
		_w22477_,
		_w22591_
	);
	LUT2 #(
		.INIT('h1)
	) name18545 (
		_w22590_,
		_w22591_,
		_w22592_
	);
	LUT2 #(
		.INIT('h4)
	) name18546 (
		_w11525_,
		_w22477_,
		_w22593_
	);
	LUT2 #(
		.INIT('h1)
	) name18547 (
		\tm_tpr_reg_DO_reg[6]/NET0131 ,
		_w22477_,
		_w22594_
	);
	LUT2 #(
		.INIT('h1)
	) name18548 (
		_w22593_,
		_w22594_,
		_w22595_
	);
	LUT2 #(
		.INIT('h4)
	) name18549 (
		_w10911_,
		_w22477_,
		_w22596_
	);
	LUT2 #(
		.INIT('h1)
	) name18550 (
		\tm_tpr_reg_DO_reg[5]/NET0131 ,
		_w22477_,
		_w22597_
	);
	LUT2 #(
		.INIT('h1)
	) name18551 (
		_w22596_,
		_w22597_,
		_w22598_
	);
	LUT2 #(
		.INIT('h4)
	) name18552 (
		_w8113_,
		_w22477_,
		_w22599_
	);
	LUT2 #(
		.INIT('h1)
	) name18553 (
		\tm_tpr_reg_DO_reg[3]/NET0131 ,
		_w22477_,
		_w22600_
	);
	LUT2 #(
		.INIT('h1)
	) name18554 (
		_w22599_,
		_w22600_,
		_w22601_
	);
	LUT2 #(
		.INIT('h4)
	) name18555 (
		_w8715_,
		_w22477_,
		_w22602_
	);
	LUT2 #(
		.INIT('h1)
	) name18556 (
		\tm_tpr_reg_DO_reg[2]/NET0131 ,
		_w22477_,
		_w22603_
	);
	LUT2 #(
		.INIT('h1)
	) name18557 (
		_w22602_,
		_w22603_,
		_w22604_
	);
	LUT2 #(
		.INIT('h4)
	) name18558 (
		_w9435_,
		_w22477_,
		_w22605_
	);
	LUT2 #(
		.INIT('h1)
	) name18559 (
		\tm_tpr_reg_DO_reg[1]/NET0131 ,
		_w22477_,
		_w22606_
	);
	LUT2 #(
		.INIT('h1)
	) name18560 (
		_w22605_,
		_w22606_,
		_w22607_
	);
	LUT2 #(
		.INIT('h4)
	) name18561 (
		_w10069_,
		_w22477_,
		_w22608_
	);
	LUT2 #(
		.INIT('h1)
	) name18562 (
		\tm_tpr_reg_DO_reg[4]/NET0131 ,
		_w22477_,
		_w22609_
	);
	LUT2 #(
		.INIT('h1)
	) name18563 (
		_w22608_,
		_w22609_,
		_w22610_
	);
	LUT2 #(
		.INIT('h4)
	) name18564 (
		_w12743_,
		_w22477_,
		_w22611_
	);
	LUT2 #(
		.INIT('h1)
	) name18565 (
		\tm_tpr_reg_DO_reg[15]/NET0131 ,
		_w22477_,
		_w22612_
	);
	LUT2 #(
		.INIT('h1)
	) name18566 (
		_w22611_,
		_w22612_,
		_w22613_
	);
	LUT2 #(
		.INIT('h4)
	) name18567 (
		_w12688_,
		_w22477_,
		_w22614_
	);
	LUT2 #(
		.INIT('h1)
	) name18568 (
		\tm_tpr_reg_DO_reg[14]/NET0131 ,
		_w22477_,
		_w22615_
	);
	LUT2 #(
		.INIT('h1)
	) name18569 (
		_w22614_,
		_w22615_,
		_w22616_
	);
	LUT2 #(
		.INIT('h4)
	) name18570 (
		_w7607_,
		_w22477_,
		_w22617_
	);
	LUT2 #(
		.INIT('h1)
	) name18571 (
		\tm_tpr_reg_DO_reg[0]/NET0131 ,
		_w22477_,
		_w22618_
	);
	LUT2 #(
		.INIT('h1)
	) name18572 (
		_w22617_,
		_w22618_,
		_w22619_
	);
	LUT2 #(
		.INIT('h4)
	) name18573 (
		_w11265_,
		_w22484_,
		_w22620_
	);
	LUT2 #(
		.INIT('h1)
	) name18574 (
		\emc_WSCRreg_DO_reg[7]/NET0131 ,
		_w22484_,
		_w22621_
	);
	LUT2 #(
		.INIT('h1)
	) name18575 (
		_w22620_,
		_w22621_,
		_w22622_
	);
	LUT2 #(
		.INIT('h4)
	) name18576 (
		_w11525_,
		_w22484_,
		_w22623_
	);
	LUT2 #(
		.INIT('h1)
	) name18577 (
		\emc_WSCRreg_DO_reg[6]/NET0131 ,
		_w22484_,
		_w22624_
	);
	LUT2 #(
		.INIT('h1)
	) name18578 (
		_w22623_,
		_w22624_,
		_w22625_
	);
	LUT2 #(
		.INIT('h4)
	) name18579 (
		_w10911_,
		_w22484_,
		_w22626_
	);
	LUT2 #(
		.INIT('h1)
	) name18580 (
		\emc_WSCRreg_DO_reg[5]/NET0131 ,
		_w22484_,
		_w22627_
	);
	LUT2 #(
		.INIT('h1)
	) name18581 (
		_w22626_,
		_w22627_,
		_w22628_
	);
	LUT2 #(
		.INIT('h4)
	) name18582 (
		_w10069_,
		_w22484_,
		_w22629_
	);
	LUT2 #(
		.INIT('h1)
	) name18583 (
		\emc_WSCRreg_DO_reg[4]/NET0131 ,
		_w22484_,
		_w22630_
	);
	LUT2 #(
		.INIT('h1)
	) name18584 (
		_w22629_,
		_w22630_,
		_w22631_
	);
	LUT2 #(
		.INIT('h4)
	) name18585 (
		_w8113_,
		_w22484_,
		_w22632_
	);
	LUT2 #(
		.INIT('h1)
	) name18586 (
		\emc_WSCRreg_DO_reg[3]/NET0131 ,
		_w22484_,
		_w22633_
	);
	LUT2 #(
		.INIT('h1)
	) name18587 (
		_w22632_,
		_w22633_,
		_w22634_
	);
	LUT2 #(
		.INIT('h4)
	) name18588 (
		_w8715_,
		_w22484_,
		_w22635_
	);
	LUT2 #(
		.INIT('h1)
	) name18589 (
		\emc_WSCRreg_DO_reg[2]/NET0131 ,
		_w22484_,
		_w22636_
	);
	LUT2 #(
		.INIT('h1)
	) name18590 (
		_w22635_,
		_w22636_,
		_w22637_
	);
	LUT2 #(
		.INIT('h4)
	) name18591 (
		_w9435_,
		_w22484_,
		_w22638_
	);
	LUT2 #(
		.INIT('h1)
	) name18592 (
		\emc_WSCRreg_DO_reg[1]/NET0131 ,
		_w22484_,
		_w22639_
	);
	LUT2 #(
		.INIT('h1)
	) name18593 (
		_w22638_,
		_w22639_,
		_w22640_
	);
	LUT2 #(
		.INIT('h4)
	) name18594 (
		_w12688_,
		_w22484_,
		_w22641_
	);
	LUT2 #(
		.INIT('h1)
	) name18595 (
		\emc_WSCRreg_DO_reg[14]/NET0131 ,
		_w22484_,
		_w22642_
	);
	LUT2 #(
		.INIT('h1)
	) name18596 (
		_w22641_,
		_w22642_,
		_w22643_
	);
	LUT2 #(
		.INIT('h4)
	) name18597 (
		_w7607_,
		_w22484_,
		_w22644_
	);
	LUT2 #(
		.INIT('h1)
	) name18598 (
		\emc_WSCRreg_DO_reg[0]/NET0131 ,
		_w22484_,
		_w22645_
	);
	LUT2 #(
		.INIT('h1)
	) name18599 (
		_w22644_,
		_w22645_,
		_w22646_
	);
	LUT2 #(
		.INIT('h8)
	) name18600 (
		\sport1_txctl_TCS_reg[0]/NET0131 ,
		\sport1_txctl_TCS_reg[2]/NET0131 ,
		_w22647_
	);
	LUT2 #(
		.INIT('h4)
	) name18601 (
		\sport1_cfg_TFSg_d1_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w22648_
	);
	LUT2 #(
		.INIT('h4)
	) name18602 (
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w22648_,
		_w22649_
	);
	LUT2 #(
		.INIT('h1)
	) name18603 (
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w22650_
	);
	LUT2 #(
		.INIT('h4)
	) name18604 (
		\ITFS1_pad ,
		\T_TFS1_pad ,
		_w22651_
	);
	LUT2 #(
		.INIT('h2)
	) name18605 (
		\ITFS1_pad ,
		_w13729_,
		_w22652_
	);
	LUT2 #(
		.INIT('h1)
	) name18606 (
		_w22651_,
		_w22652_,
		_w22653_
	);
	LUT2 #(
		.INIT('h2)
	) name18607 (
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w22653_,
		_w22654_
	);
	LUT2 #(
		.INIT('h4)
	) name18608 (
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w22653_,
		_w22655_
	);
	LUT2 #(
		.INIT('h1)
	) name18609 (
		_w22654_,
		_w22655_,
		_w22656_
	);
	LUT2 #(
		.INIT('h2)
	) name18610 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_cfg_TFSgi_d_reg/NET0131 ,
		_w22657_
	);
	LUT2 #(
		.INIT('h8)
	) name18611 (
		_w22656_,
		_w22657_,
		_w22658_
	);
	LUT2 #(
		.INIT('h2)
	) name18612 (
		_w22650_,
		_w22658_,
		_w22659_
	);
	LUT2 #(
		.INIT('h2)
	) name18613 (
		\sport1_cfg_TFSg_d2_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w22660_
	);
	LUT2 #(
		.INIT('h8)
	) name18614 (
		\sport1_cfg_TFSg_d3_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w22661_
	);
	LUT2 #(
		.INIT('h2)
	) name18615 (
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w22660_,
		_w22662_
	);
	LUT2 #(
		.INIT('h4)
	) name18616 (
		_w22661_,
		_w22662_,
		_w22663_
	);
	LUT2 #(
		.INIT('h2)
	) name18617 (
		\sport1_txctl_TCS_reg[0]/NET0131 ,
		_w22649_,
		_w22664_
	);
	LUT2 #(
		.INIT('h4)
	) name18618 (
		_w22663_,
		_w22664_,
		_w22665_
	);
	LUT2 #(
		.INIT('h4)
	) name18619 (
		_w22659_,
		_w22665_,
		_w22666_
	);
	LUT2 #(
		.INIT('h1)
	) name18620 (
		\sport1_txctl_TCS_reg[2]/NET0131 ,
		_w22666_,
		_w22667_
	);
	LUT2 #(
		.INIT('h1)
	) name18621 (
		\sport1_txctl_TCS_reg[1]/NET0131 ,
		_w22647_,
		_w22668_
	);
	LUT2 #(
		.INIT('h4)
	) name18622 (
		_w22667_,
		_w22668_,
		_w22669_
	);
	LUT2 #(
		.INIT('h4)
	) name18623 (
		\sport1_txctl_TCS_reg[0]/NET0131 ,
		\sport1_txctl_TCS_reg[1]/NET0131 ,
		_w22670_
	);
	LUT2 #(
		.INIT('h4)
	) name18624 (
		\sport1_txctl_TCS_reg[2]/NET0131 ,
		_w22670_,
		_w22671_
	);
	LUT2 #(
		.INIT('h1)
	) name18625 (
		\sport1_txctl_Bcnt_reg[0]/NET0131 ,
		\sport1_txctl_Bcnt_reg[1]/NET0131 ,
		_w22672_
	);
	LUT2 #(
		.INIT('h4)
	) name18626 (
		\sport1_txctl_Bcnt_reg[2]/NET0131 ,
		_w22672_,
		_w22673_
	);
	LUT2 #(
		.INIT('h4)
	) name18627 (
		\sport1_txctl_Bcnt_reg[3]/NET0131 ,
		_w22673_,
		_w22674_
	);
	LUT2 #(
		.INIT('h4)
	) name18628 (
		\sport1_txctl_Bcnt_reg[4]/NET0131 ,
		_w22674_,
		_w22675_
	);
	LUT2 #(
		.INIT('h2)
	) name18629 (
		_w22671_,
		_w22675_,
		_w22676_
	);
	LUT2 #(
		.INIT('h1)
	) name18630 (
		_w22669_,
		_w22676_,
		_w22677_
	);
	LUT2 #(
		.INIT('h2)
	) name18631 (
		\sport1_txctl_TXSHT_reg[9]/P0001 ,
		_w22677_,
		_w22678_
	);
	LUT2 #(
		.INIT('h8)
	) name18632 (
		\sport1_txctl_TX_reg[10]/P0001 ,
		_w22677_,
		_w22679_
	);
	LUT2 #(
		.INIT('h1)
	) name18633 (
		_w22678_,
		_w22679_,
		_w22680_
	);
	LUT2 #(
		.INIT('h2)
	) name18634 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 ,
		_w18266_,
		_w22681_
	);
	LUT2 #(
		.INIT('h1)
	) name18635 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[4]/P0001 ,
		_w18271_,
		_w22682_
	);
	LUT2 #(
		.INIT('h2)
	) name18636 (
		_w18271_,
		_w20080_,
		_w22683_
	);
	LUT2 #(
		.INIT('h2)
	) name18637 (
		_w18273_,
		_w22682_,
		_w22684_
	);
	LUT2 #(
		.INIT('h4)
	) name18638 (
		_w22683_,
		_w22684_,
		_w22685_
	);
	LUT2 #(
		.INIT('h1)
	) name18639 (
		_w18270_,
		_w22681_,
		_w22686_
	);
	LUT2 #(
		.INIT('h4)
	) name18640 (
		_w22685_,
		_w22686_,
		_w22687_
	);
	LUT2 #(
		.INIT('h1)
	) name18641 (
		_w18262_,
		_w22687_,
		_w22688_
	);
	LUT2 #(
		.INIT('h2)
	) name18642 (
		_w18262_,
		_w19670_,
		_w22689_
	);
	LUT2 #(
		.INIT('h1)
	) name18643 (
		_w22688_,
		_w22689_,
		_w22690_
	);
	LUT2 #(
		.INIT('h8)
	) name18644 (
		_w14752_,
		_w19670_,
		_w22691_
	);
	LUT2 #(
		.INIT('h8)
	) name18645 (
		_w18328_,
		_w20080_,
		_w22692_
	);
	LUT2 #(
		.INIT('h2)
	) name18646 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[4]/P0001 ,
		_w18330_,
		_w22693_
	);
	LUT2 #(
		.INIT('h2)
	) name18647 (
		_w18334_,
		_w22693_,
		_w22694_
	);
	LUT2 #(
		.INIT('h4)
	) name18648 (
		_w22692_,
		_w22694_,
		_w22695_
	);
	LUT2 #(
		.INIT('h1)
	) name18649 (
		_w22691_,
		_w22695_,
		_w22696_
	);
	LUT2 #(
		.INIT('h8)
	) name18650 (
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w21318_,
		_w22697_
	);
	LUT2 #(
		.INIT('h8)
	) name18651 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w18514_,
		_w22698_
	);
	LUT2 #(
		.INIT('h8)
	) name18652 (
		_w11525_,
		_w21316_,
		_w22699_
	);
	LUT2 #(
		.INIT('h1)
	) name18653 (
		_w22697_,
		_w22699_,
		_w22700_
	);
	LUT2 #(
		.INIT('h4)
	) name18654 (
		_w22698_,
		_w22700_,
		_w22701_
	);
	LUT2 #(
		.INIT('h1)
	) name18655 (
		_w15120_,
		_w15183_,
		_w22702_
	);
	LUT2 #(
		.INIT('h4)
	) name18656 (
		_w15319_,
		_w22702_,
		_w22703_
	);
	LUT2 #(
		.INIT('h4)
	) name18657 (
		_w17777_,
		_w22703_,
		_w22704_
	);
	LUT2 #(
		.INIT('h4)
	) name18658 (
		_w15120_,
		_w15182_,
		_w22705_
	);
	LUT2 #(
		.INIT('h4)
	) name18659 (
		_w17783_,
		_w22702_,
		_w22706_
	);
	LUT2 #(
		.INIT('h1)
	) name18660 (
		_w15121_,
		_w22705_,
		_w22707_
	);
	LUT2 #(
		.INIT('h4)
	) name18661 (
		_w22706_,
		_w22707_,
		_w22708_
	);
	LUT2 #(
		.INIT('h4)
	) name18662 (
		_w22704_,
		_w22708_,
		_w22709_
	);
	LUT2 #(
		.INIT('h1)
	) name18663 (
		_w14933_,
		_w15053_,
		_w22710_
	);
	LUT2 #(
		.INIT('h4)
	) name18664 (
		_w9865_,
		_w14993_,
		_w22711_
	);
	LUT2 #(
		.INIT('h8)
	) name18665 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w15046_,
		_w22712_
	);
	LUT2 #(
		.INIT('h1)
	) name18666 (
		_w22711_,
		_w22712_,
		_w22713_
	);
	LUT2 #(
		.INIT('h1)
	) name18667 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w22713_,
		_w22714_
	);
	LUT2 #(
		.INIT('h4)
	) name18668 (
		_w14972_,
		_w22714_,
		_w22715_
	);
	LUT2 #(
		.INIT('h2)
	) name18669 (
		_w14972_,
		_w22714_,
		_w22716_
	);
	LUT2 #(
		.INIT('h1)
	) name18670 (
		_w22715_,
		_w22716_,
		_w22717_
	);
	LUT2 #(
		.INIT('h1)
	) name18671 (
		_w15051_,
		_w22717_,
		_w22718_
	);
	LUT2 #(
		.INIT('h8)
	) name18672 (
		_w15051_,
		_w22713_,
		_w22719_
	);
	LUT2 #(
		.INIT('h1)
	) name18673 (
		_w22718_,
		_w22719_,
		_w22720_
	);
	LUT2 #(
		.INIT('h2)
	) name18674 (
		_w14992_,
		_w22720_,
		_w22721_
	);
	LUT2 #(
		.INIT('h4)
	) name18675 (
		_w14992_,
		_w22720_,
		_w22722_
	);
	LUT2 #(
		.INIT('h1)
	) name18676 (
		_w22721_,
		_w22722_,
		_w22723_
	);
	LUT2 #(
		.INIT('h1)
	) name18677 (
		_w22710_,
		_w22723_,
		_w22724_
	);
	LUT2 #(
		.INIT('h8)
	) name18678 (
		_w22710_,
		_w22723_,
		_w22725_
	);
	LUT2 #(
		.INIT('h1)
	) name18679 (
		_w22724_,
		_w22725_,
		_w22726_
	);
	LUT2 #(
		.INIT('h1)
	) name18680 (
		_w14991_,
		_w15054_,
		_w22727_
	);
	LUT2 #(
		.INIT('h8)
	) name18681 (
		_w15058_,
		_w22727_,
		_w22728_
	);
	LUT2 #(
		.INIT('h1)
	) name18682 (
		_w15059_,
		_w22728_,
		_w22729_
	);
	LUT2 #(
		.INIT('h2)
	) name18683 (
		_w22726_,
		_w22729_,
		_w22730_
	);
	LUT2 #(
		.INIT('h1)
	) name18684 (
		_w14853_,
		_w22730_,
		_w22731_
	);
	LUT2 #(
		.INIT('h1)
	) name18685 (
		_w14933_,
		_w22718_,
		_w22732_
	);
	LUT2 #(
		.INIT('h4)
	) name18686 (
		_w10882_,
		_w14993_,
		_w22733_
	);
	LUT2 #(
		.INIT('h4)
	) name18687 (
		_w9865_,
		_w15044_,
		_w22734_
	);
	LUT2 #(
		.INIT('h1)
	) name18688 (
		_w22733_,
		_w22734_,
		_w22735_
	);
	LUT2 #(
		.INIT('h1)
	) name18689 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w22735_,
		_w22736_
	);
	LUT2 #(
		.INIT('h4)
	) name18690 (
		_w14972_,
		_w22736_,
		_w22737_
	);
	LUT2 #(
		.INIT('h2)
	) name18691 (
		_w14972_,
		_w22736_,
		_w22738_
	);
	LUT2 #(
		.INIT('h1)
	) name18692 (
		_w22737_,
		_w22738_,
		_w22739_
	);
	LUT2 #(
		.INIT('h1)
	) name18693 (
		_w22715_,
		_w22739_,
		_w22740_
	);
	LUT2 #(
		.INIT('h8)
	) name18694 (
		_w22715_,
		_w22735_,
		_w22741_
	);
	LUT2 #(
		.INIT('h1)
	) name18695 (
		_w22740_,
		_w22741_,
		_w22742_
	);
	LUT2 #(
		.INIT('h2)
	) name18696 (
		_w14992_,
		_w22742_,
		_w22743_
	);
	LUT2 #(
		.INIT('h4)
	) name18697 (
		_w14992_,
		_w22742_,
		_w22744_
	);
	LUT2 #(
		.INIT('h1)
	) name18698 (
		_w22743_,
		_w22744_,
		_w22745_
	);
	LUT2 #(
		.INIT('h2)
	) name18699 (
		_w22732_,
		_w22745_,
		_w22746_
	);
	LUT2 #(
		.INIT('h4)
	) name18700 (
		_w22732_,
		_w22745_,
		_w22747_
	);
	LUT2 #(
		.INIT('h1)
	) name18701 (
		_w22746_,
		_w22747_,
		_w22748_
	);
	LUT2 #(
		.INIT('h1)
	) name18702 (
		_w14991_,
		_w22719_,
		_w22749_
	);
	LUT2 #(
		.INIT('h8)
	) name18703 (
		_w22723_,
		_w22749_,
		_w22750_
	);
	LUT2 #(
		.INIT('h1)
	) name18704 (
		_w22724_,
		_w22750_,
		_w22751_
	);
	LUT2 #(
		.INIT('h1)
	) name18705 (
		_w22748_,
		_w22751_,
		_w22752_
	);
	LUT2 #(
		.INIT('h8)
	) name18706 (
		_w22748_,
		_w22751_,
		_w22753_
	);
	LUT2 #(
		.INIT('h1)
	) name18707 (
		_w22752_,
		_w22753_,
		_w22754_
	);
	LUT2 #(
		.INIT('h8)
	) name18708 (
		_w14853_,
		_w22754_,
		_w22755_
	);
	LUT2 #(
		.INIT('h1)
	) name18709 (
		_w14853_,
		_w22754_,
		_w22756_
	);
	LUT2 #(
		.INIT('h1)
	) name18710 (
		_w22755_,
		_w22756_,
		_w22757_
	);
	LUT2 #(
		.INIT('h1)
	) name18711 (
		_w22731_,
		_w22757_,
		_w22758_
	);
	LUT2 #(
		.INIT('h8)
	) name18712 (
		_w22731_,
		_w22754_,
		_w22759_
	);
	LUT2 #(
		.INIT('h1)
	) name18713 (
		_w22758_,
		_w22759_,
		_w22760_
	);
	LUT2 #(
		.INIT('h4)
	) name18714 (
		_w14853_,
		_w15065_,
		_w22761_
	);
	LUT2 #(
		.INIT('h4)
	) name18715 (
		_w22726_,
		_w22729_,
		_w22762_
	);
	LUT2 #(
		.INIT('h1)
	) name18716 (
		_w22730_,
		_w22762_,
		_w22763_
	);
	LUT2 #(
		.INIT('h8)
	) name18717 (
		_w22761_,
		_w22763_,
		_w22764_
	);
	LUT2 #(
		.INIT('h1)
	) name18718 (
		_w22761_,
		_w22763_,
		_w22765_
	);
	LUT2 #(
		.INIT('h1)
	) name18719 (
		_w22764_,
		_w22765_,
		_w22766_
	);
	LUT2 #(
		.INIT('h4)
	) name18720 (
		_w22760_,
		_w22766_,
		_w22767_
	);
	LUT2 #(
		.INIT('h2)
	) name18721 (
		_w14853_,
		_w22729_,
		_w22768_
	);
	LUT2 #(
		.INIT('h2)
	) name18722 (
		_w22765_,
		_w22768_,
		_w22769_
	);
	LUT2 #(
		.INIT('h2)
	) name18723 (
		_w22760_,
		_w22769_,
		_w22770_
	);
	LUT2 #(
		.INIT('h1)
	) name18724 (
		_w15066_,
		_w15070_,
		_w22771_
	);
	LUT2 #(
		.INIT('h1)
	) name18725 (
		_w15071_,
		_w22771_,
		_w22772_
	);
	LUT2 #(
		.INIT('h4)
	) name18726 (
		_w22770_,
		_w22772_,
		_w22773_
	);
	LUT2 #(
		.INIT('h1)
	) name18727 (
		_w22767_,
		_w22773_,
		_w22774_
	);
	LUT2 #(
		.INIT('h1)
	) name18728 (
		_w22709_,
		_w22774_,
		_w22775_
	);
	LUT2 #(
		.INIT('h4)
	) name18729 (
		_w22760_,
		_w22769_,
		_w22776_
	);
	LUT2 #(
		.INIT('h8)
	) name18730 (
		_w22767_,
		_w22772_,
		_w22777_
	);
	LUT2 #(
		.INIT('h1)
	) name18731 (
		_w22776_,
		_w22777_,
		_w22778_
	);
	LUT2 #(
		.INIT('h4)
	) name18732 (
		_w22775_,
		_w22778_,
		_w22779_
	);
	LUT2 #(
		.INIT('h1)
	) name18733 (
		_w14853_,
		_w22752_,
		_w22780_
	);
	LUT2 #(
		.INIT('h1)
	) name18734 (
		_w14933_,
		_w22740_,
		_w22781_
	);
	LUT2 #(
		.INIT('h4)
	) name18735 (
		_w11424_,
		_w14993_,
		_w22782_
	);
	LUT2 #(
		.INIT('h4)
	) name18736 (
		_w10882_,
		_w15044_,
		_w22783_
	);
	LUT2 #(
		.INIT('h1)
	) name18737 (
		_w22782_,
		_w22783_,
		_w22784_
	);
	LUT2 #(
		.INIT('h1)
	) name18738 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w22784_,
		_w22785_
	);
	LUT2 #(
		.INIT('h4)
	) name18739 (
		_w14972_,
		_w22785_,
		_w22786_
	);
	LUT2 #(
		.INIT('h2)
	) name18740 (
		_w14972_,
		_w22785_,
		_w22787_
	);
	LUT2 #(
		.INIT('h1)
	) name18741 (
		_w22786_,
		_w22787_,
		_w22788_
	);
	LUT2 #(
		.INIT('h1)
	) name18742 (
		_w22737_,
		_w22788_,
		_w22789_
	);
	LUT2 #(
		.INIT('h8)
	) name18743 (
		_w22737_,
		_w22784_,
		_w22790_
	);
	LUT2 #(
		.INIT('h1)
	) name18744 (
		_w22789_,
		_w22790_,
		_w22791_
	);
	LUT2 #(
		.INIT('h2)
	) name18745 (
		_w14992_,
		_w22791_,
		_w22792_
	);
	LUT2 #(
		.INIT('h4)
	) name18746 (
		_w14992_,
		_w22791_,
		_w22793_
	);
	LUT2 #(
		.INIT('h1)
	) name18747 (
		_w22792_,
		_w22793_,
		_w22794_
	);
	LUT2 #(
		.INIT('h2)
	) name18748 (
		_w22781_,
		_w22794_,
		_w22795_
	);
	LUT2 #(
		.INIT('h4)
	) name18749 (
		_w22781_,
		_w22794_,
		_w22796_
	);
	LUT2 #(
		.INIT('h1)
	) name18750 (
		_w22795_,
		_w22796_,
		_w22797_
	);
	LUT2 #(
		.INIT('h1)
	) name18751 (
		_w14991_,
		_w22741_,
		_w22798_
	);
	LUT2 #(
		.INIT('h2)
	) name18752 (
		_w22745_,
		_w22798_,
		_w22799_
	);
	LUT2 #(
		.INIT('h1)
	) name18753 (
		_w22746_,
		_w22799_,
		_w22800_
	);
	LUT2 #(
		.INIT('h4)
	) name18754 (
		_w22797_,
		_w22800_,
		_w22801_
	);
	LUT2 #(
		.INIT('h2)
	) name18755 (
		_w22797_,
		_w22800_,
		_w22802_
	);
	LUT2 #(
		.INIT('h1)
	) name18756 (
		_w22801_,
		_w22802_,
		_w22803_
	);
	LUT2 #(
		.INIT('h8)
	) name18757 (
		_w14853_,
		_w22803_,
		_w22804_
	);
	LUT2 #(
		.INIT('h1)
	) name18758 (
		_w14853_,
		_w22803_,
		_w22805_
	);
	LUT2 #(
		.INIT('h1)
	) name18759 (
		_w22804_,
		_w22805_,
		_w22806_
	);
	LUT2 #(
		.INIT('h1)
	) name18760 (
		_w22780_,
		_w22806_,
		_w22807_
	);
	LUT2 #(
		.INIT('h4)
	) name18761 (
		_w22802_,
		_w22806_,
		_w22808_
	);
	LUT2 #(
		.INIT('h1)
	) name18762 (
		_w22807_,
		_w22808_,
		_w22809_
	);
	LUT2 #(
		.INIT('h1)
	) name18763 (
		_w14933_,
		_w22789_,
		_w22810_
	);
	LUT2 #(
		.INIT('h4)
	) name18764 (
		_w7206_,
		_w14993_,
		_w22811_
	);
	LUT2 #(
		.INIT('h4)
	) name18765 (
		_w11424_,
		_w15044_,
		_w22812_
	);
	LUT2 #(
		.INIT('h1)
	) name18766 (
		_w22811_,
		_w22812_,
		_w22813_
	);
	LUT2 #(
		.INIT('h1)
	) name18767 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w22813_,
		_w22814_
	);
	LUT2 #(
		.INIT('h1)
	) name18768 (
		_w14972_,
		_w22814_,
		_w22815_
	);
	LUT2 #(
		.INIT('h8)
	) name18769 (
		_w14972_,
		_w22814_,
		_w22816_
	);
	LUT2 #(
		.INIT('h1)
	) name18770 (
		_w22786_,
		_w22815_,
		_w22817_
	);
	LUT2 #(
		.INIT('h4)
	) name18771 (
		_w22816_,
		_w22817_,
		_w22818_
	);
	LUT2 #(
		.INIT('h2)
	) name18772 (
		_w22786_,
		_w22814_,
		_w22819_
	);
	LUT2 #(
		.INIT('h1)
	) name18773 (
		_w22818_,
		_w22819_,
		_w22820_
	);
	LUT2 #(
		.INIT('h2)
	) name18774 (
		_w14992_,
		_w22820_,
		_w22821_
	);
	LUT2 #(
		.INIT('h4)
	) name18775 (
		_w14992_,
		_w22820_,
		_w22822_
	);
	LUT2 #(
		.INIT('h1)
	) name18776 (
		_w22821_,
		_w22822_,
		_w22823_
	);
	LUT2 #(
		.INIT('h4)
	) name18777 (
		_w22810_,
		_w22823_,
		_w22824_
	);
	LUT2 #(
		.INIT('h2)
	) name18778 (
		_w22810_,
		_w22823_,
		_w22825_
	);
	LUT2 #(
		.INIT('h1)
	) name18779 (
		_w22824_,
		_w22825_,
		_w22826_
	);
	LUT2 #(
		.INIT('h1)
	) name18780 (
		_w14991_,
		_w22790_,
		_w22827_
	);
	LUT2 #(
		.INIT('h2)
	) name18781 (
		_w22794_,
		_w22827_,
		_w22828_
	);
	LUT2 #(
		.INIT('h1)
	) name18782 (
		_w22795_,
		_w22828_,
		_w22829_
	);
	LUT2 #(
		.INIT('h4)
	) name18783 (
		_w22826_,
		_w22829_,
		_w22830_
	);
	LUT2 #(
		.INIT('h2)
	) name18784 (
		_w22826_,
		_w22829_,
		_w22831_
	);
	LUT2 #(
		.INIT('h1)
	) name18785 (
		_w22830_,
		_w22831_,
		_w22832_
	);
	LUT2 #(
		.INIT('h4)
	) name18786 (
		_w14853_,
		_w22801_,
		_w22833_
	);
	LUT2 #(
		.INIT('h4)
	) name18787 (
		_w22832_,
		_w22833_,
		_w22834_
	);
	LUT2 #(
		.INIT('h2)
	) name18788 (
		_w22832_,
		_w22833_,
		_w22835_
	);
	LUT2 #(
		.INIT('h1)
	) name18789 (
		_w22834_,
		_w22835_,
		_w22836_
	);
	LUT2 #(
		.INIT('h4)
	) name18790 (
		_w22809_,
		_w22836_,
		_w22837_
	);
	LUT2 #(
		.INIT('h4)
	) name18791 (
		_w22753_,
		_w22757_,
		_w22838_
	);
	LUT2 #(
		.INIT('h1)
	) name18792 (
		_w22758_,
		_w22838_,
		_w22839_
	);
	LUT2 #(
		.INIT('h8)
	) name18793 (
		_w22780_,
		_w22803_,
		_w22840_
	);
	LUT2 #(
		.INIT('h1)
	) name18794 (
		_w22807_,
		_w22840_,
		_w22841_
	);
	LUT2 #(
		.INIT('h4)
	) name18795 (
		_w22839_,
		_w22841_,
		_w22842_
	);
	LUT2 #(
		.INIT('h1)
	) name18796 (
		_w22837_,
		_w22842_,
		_w22843_
	);
	LUT2 #(
		.INIT('h4)
	) name18797 (
		_w22779_,
		_w22843_,
		_w22844_
	);
	LUT2 #(
		.INIT('h2)
	) name18798 (
		_w22809_,
		_w22836_,
		_w22845_
	);
	LUT2 #(
		.INIT('h2)
	) name18799 (
		_w22839_,
		_w22841_,
		_w22846_
	);
	LUT2 #(
		.INIT('h4)
	) name18800 (
		_w22837_,
		_w22846_,
		_w22847_
	);
	LUT2 #(
		.INIT('h1)
	) name18801 (
		_w22845_,
		_w22847_,
		_w22848_
	);
	LUT2 #(
		.INIT('h4)
	) name18802 (
		_w22844_,
		_w22848_,
		_w22849_
	);
	LUT2 #(
		.INIT('h4)
	) name18803 (
		_w7206_,
		_w17443_,
		_w22850_
	);
	LUT2 #(
		.INIT('h1)
	) name18804 (
		_w14991_,
		_w22819_,
		_w22851_
	);
	LUT2 #(
		.INIT('h2)
	) name18805 (
		_w22823_,
		_w22851_,
		_w22852_
	);
	LUT2 #(
		.INIT('h1)
	) name18806 (
		_w22825_,
		_w22852_,
		_w22853_
	);
	LUT2 #(
		.INIT('h2)
	) name18807 (
		_w22815_,
		_w22853_,
		_w22854_
	);
	LUT2 #(
		.INIT('h4)
	) name18808 (
		_w22815_,
		_w22853_,
		_w22855_
	);
	LUT2 #(
		.INIT('h1)
	) name18809 (
		_w22854_,
		_w22855_,
		_w22856_
	);
	LUT2 #(
		.INIT('h8)
	) name18810 (
		_w22850_,
		_w22856_,
		_w22857_
	);
	LUT2 #(
		.INIT('h1)
	) name18811 (
		_w22850_,
		_w22856_,
		_w22858_
	);
	LUT2 #(
		.INIT('h1)
	) name18812 (
		_w22857_,
		_w22858_,
		_w22859_
	);
	LUT2 #(
		.INIT('h4)
	) name18813 (
		_w22830_,
		_w22833_,
		_w22860_
	);
	LUT2 #(
		.INIT('h1)
	) name18814 (
		_w22831_,
		_w22833_,
		_w22861_
	);
	LUT2 #(
		.INIT('h1)
	) name18815 (
		_w22860_,
		_w22861_,
		_w22862_
	);
	LUT2 #(
		.INIT('h2)
	) name18816 (
		_w22859_,
		_w22862_,
		_w22863_
	);
	LUT2 #(
		.INIT('h4)
	) name18817 (
		_w22859_,
		_w22862_,
		_w22864_
	);
	LUT2 #(
		.INIT('h1)
	) name18818 (
		_w22863_,
		_w22864_,
		_w22865_
	);
	LUT2 #(
		.INIT('h1)
	) name18819 (
		_w14991_,
		_w22818_,
		_w22866_
	);
	LUT2 #(
		.INIT('h4)
	) name18820 (
		_w14992_,
		_w22818_,
		_w22867_
	);
	LUT2 #(
		.INIT('h1)
	) name18821 (
		_w22866_,
		_w22867_,
		_w22868_
	);
	LUT2 #(
		.INIT('h2)
	) name18822 (
		_w22865_,
		_w22868_,
		_w22869_
	);
	LUT2 #(
		.INIT('h4)
	) name18823 (
		_w22865_,
		_w22868_,
		_w22870_
	);
	LUT2 #(
		.INIT('h1)
	) name18824 (
		_w22869_,
		_w22870_,
		_w22871_
	);
	LUT2 #(
		.INIT('h8)
	) name18825 (
		_w22849_,
		_w22871_,
		_w22872_
	);
	LUT2 #(
		.INIT('h1)
	) name18826 (
		_w22849_,
		_w22871_,
		_w22873_
	);
	LUT2 #(
		.INIT('h1)
	) name18827 (
		_w22872_,
		_w22873_,
		_w22874_
	);
	LUT2 #(
		.INIT('h2)
	) name18828 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22874_,
		_w22875_
	);
	LUT2 #(
		.INIT('h1)
	) name18829 (
		_w22837_,
		_w22845_,
		_w22876_
	);
	LUT2 #(
		.INIT('h1)
	) name18830 (
		_w22779_,
		_w22842_,
		_w22877_
	);
	LUT2 #(
		.INIT('h1)
	) name18831 (
		_w22846_,
		_w22877_,
		_w22878_
	);
	LUT2 #(
		.INIT('h2)
	) name18832 (
		_w22876_,
		_w22878_,
		_w22879_
	);
	LUT2 #(
		.INIT('h4)
	) name18833 (
		_w22876_,
		_w22878_,
		_w22880_
	);
	LUT2 #(
		.INIT('h1)
	) name18834 (
		_w22879_,
		_w22880_,
		_w22881_
	);
	LUT2 #(
		.INIT('h4)
	) name18835 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22881_,
		_w22882_
	);
	LUT2 #(
		.INIT('h1)
	) name18836 (
		_w22875_,
		_w22882_,
		_w22883_
	);
	LUT2 #(
		.INIT('h2)
	) name18837 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w20080_,
		_w22884_
	);
	LUT2 #(
		.INIT('h1)
	) name18838 (
		_w18909_,
		_w19870_,
		_w22885_
	);
	LUT2 #(
		.INIT('h2)
	) name18839 (
		_w18752_,
		_w18907_,
		_w22886_
	);
	LUT2 #(
		.INIT('h1)
	) name18840 (
		_w18914_,
		_w18919_,
		_w22887_
	);
	LUT2 #(
		.INIT('h2)
	) name18841 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9951_,
		_w22888_
	);
	LUT2 #(
		.INIT('h2)
	) name18842 (
		_w18763_,
		_w18918_,
		_w22889_
	);
	LUT2 #(
		.INIT('h1)
	) name18843 (
		_w18079_,
		_w19864_,
		_w22890_
	);
	LUT2 #(
		.INIT('h2)
	) name18844 (
		_w18746_,
		_w18918_,
		_w22891_
	);
	LUT2 #(
		.INIT('h2)
	) name18845 (
		_w18758_,
		_w18898_,
		_w22892_
	);
	LUT2 #(
		.INIT('h1)
	) name18846 (
		_w18743_,
		_w18912_,
		_w22893_
	);
	LUT2 #(
		.INIT('h2)
	) name18847 (
		_w17925_,
		_w18888_,
		_w22894_
	);
	LUT2 #(
		.INIT('h4)
	) name18848 (
		_w17938_,
		_w18083_,
		_w22895_
	);
	LUT2 #(
		.INIT('h4)
	) name18849 (
		_w17998_,
		_w18183_,
		_w22896_
	);
	LUT2 #(
		.INIT('h8)
	) name18850 (
		_w17991_,
		_w18765_,
		_w22897_
	);
	LUT2 #(
		.INIT('h1)
	) name18851 (
		_w20272_,
		_w22888_,
		_w22898_
	);
	LUT2 #(
		.INIT('h4)
	) name18852 (
		_w22885_,
		_w22898_,
		_w22899_
	);
	LUT2 #(
		.INIT('h1)
	) name18853 (
		_w22886_,
		_w22887_,
		_w22900_
	);
	LUT2 #(
		.INIT('h1)
	) name18854 (
		_w22889_,
		_w22890_,
		_w22901_
	);
	LUT2 #(
		.INIT('h1)
	) name18855 (
		_w22891_,
		_w22893_,
		_w22902_
	);
	LUT2 #(
		.INIT('h4)
	) name18856 (
		_w22897_,
		_w22902_,
		_w22903_
	);
	LUT2 #(
		.INIT('h8)
	) name18857 (
		_w22900_,
		_w22901_,
		_w22904_
	);
	LUT2 #(
		.INIT('h4)
	) name18858 (
		_w22892_,
		_w22899_,
		_w22905_
	);
	LUT2 #(
		.INIT('h1)
	) name18859 (
		_w22894_,
		_w22895_,
		_w22906_
	);
	LUT2 #(
		.INIT('h4)
	) name18860 (
		_w22896_,
		_w22906_,
		_w22907_
	);
	LUT2 #(
		.INIT('h8)
	) name18861 (
		_w22904_,
		_w22905_,
		_w22908_
	);
	LUT2 #(
		.INIT('h8)
	) name18862 (
		_w22903_,
		_w22908_,
		_w22909_
	);
	LUT2 #(
		.INIT('h8)
	) name18863 (
		_w22907_,
		_w22909_,
		_w22910_
	);
	LUT2 #(
		.INIT('h8)
	) name18864 (
		_w20274_,
		_w22910_,
		_w22911_
	);
	LUT2 #(
		.INIT('h4)
	) name18865 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w22911_,
		_w22912_
	);
	LUT2 #(
		.INIT('h1)
	) name18866 (
		_w22884_,
		_w22912_,
		_w22913_
	);
	LUT2 #(
		.INIT('h2)
	) name18867 (
		_w18886_,
		_w22913_,
		_w22914_
	);
	LUT2 #(
		.INIT('h1)
	) name18868 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[4]/P0001 ,
		_w18886_,
		_w22915_
	);
	LUT2 #(
		.INIT('h1)
	) name18869 (
		_w22914_,
		_w22915_,
		_w22916_
	);
	LUT2 #(
		.INIT('h2)
	) name18870 (
		_w19034_,
		_w22913_,
		_w22917_
	);
	LUT2 #(
		.INIT('h1)
	) name18871 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[4]/P0001 ,
		_w19034_,
		_w22918_
	);
	LUT2 #(
		.INIT('h1)
	) name18872 (
		_w22917_,
		_w22918_,
		_w22919_
	);
	LUT2 #(
		.INIT('h8)
	) name18873 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22881_,
		_w22920_
	);
	LUT2 #(
		.INIT('h1)
	) name18874 (
		_w22842_,
		_w22846_,
		_w22921_
	);
	LUT2 #(
		.INIT('h4)
	) name18875 (
		_w22779_,
		_w22921_,
		_w22922_
	);
	LUT2 #(
		.INIT('h2)
	) name18876 (
		_w22779_,
		_w22921_,
		_w22923_
	);
	LUT2 #(
		.INIT('h1)
	) name18877 (
		_w22922_,
		_w22923_,
		_w22924_
	);
	LUT2 #(
		.INIT('h4)
	) name18878 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22924_,
		_w22925_
	);
	LUT2 #(
		.INIT('h1)
	) name18879 (
		_w22920_,
		_w22925_,
		_w22926_
	);
	LUT2 #(
		.INIT('h2)
	) name18880 (
		\core_eu_em_mac_em_reg_mrovfwe_DO_reg[0]/P0001 ,
		_w21314_,
		_w22927_
	);
	LUT2 #(
		.INIT('h4)
	) name18881 (
		_w19379_,
		_w21314_,
		_w22928_
	);
	LUT2 #(
		.INIT('h1)
	) name18882 (
		_w22927_,
		_w22928_,
		_w22929_
	);
	LUT2 #(
		.INIT('h8)
	) name18883 (
		\core_c_dec_satMR_E_reg/P0001 ,
		_w4117_,
		_w22930_
	);
	LUT2 #(
		.INIT('h8)
	) name18884 (
		_w19696_,
		_w21557_,
		_w22931_
	);
	LUT2 #(
		.INIT('h1)
	) name18885 (
		_w22930_,
		_w22931_,
		_w22932_
	);
	LUT2 #(
		.INIT('h2)
	) name18886 (
		_w4116_,
		_w22932_,
		_w22933_
	);
	LUT2 #(
		.INIT('h8)
	) name18887 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w4117_,
		_w22934_
	);
	LUT2 #(
		.INIT('h1)
	) name18888 (
		_w21558_,
		_w22934_,
		_w22935_
	);
	LUT2 #(
		.INIT('h2)
	) name18889 (
		_w4116_,
		_w22935_,
		_w22936_
	);
	LUT2 #(
		.INIT('h1)
	) name18890 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 ,
		_w19499_,
		_w22937_
	);
	LUT2 #(
		.INIT('h2)
	) name18891 (
		_w19499_,
		_w19972_,
		_w22938_
	);
	LUT2 #(
		.INIT('h2)
	) name18892 (
		_w19501_,
		_w22937_,
		_w22939_
	);
	LUT2 #(
		.INIT('h4)
	) name18893 (
		_w22938_,
		_w22939_,
		_w22940_
	);
	LUT2 #(
		.INIT('h2)
	) name18894 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[7]/P0001 ,
		_w19383_,
		_w22941_
	);
	LUT2 #(
		.INIT('h1)
	) name18895 (
		_w19508_,
		_w22941_,
		_w22942_
	);
	LUT2 #(
		.INIT('h4)
	) name18896 (
		_w22940_,
		_w22942_,
		_w22943_
	);
	LUT2 #(
		.INIT('h1)
	) name18897 (
		_w18262_,
		_w22943_,
		_w22944_
	);
	LUT2 #(
		.INIT('h1)
	) name18898 (
		_w16979_,
		_w17688_,
		_w22945_
	);
	LUT2 #(
		.INIT('h4)
	) name18899 (
		_w19424_,
		_w22945_,
		_w22946_
	);
	LUT2 #(
		.INIT('h2)
	) name18900 (
		_w19424_,
		_w22945_,
		_w22947_
	);
	LUT2 #(
		.INIT('h1)
	) name18901 (
		_w22946_,
		_w22947_,
		_w22948_
	);
	LUT2 #(
		.INIT('h2)
	) name18902 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22948_,
		_w22949_
	);
	LUT2 #(
		.INIT('h2)
	) name18903 (
		_w17544_,
		_w19422_,
		_w22950_
	);
	LUT2 #(
		.INIT('h1)
	) name18904 (
		_w17679_,
		_w22950_,
		_w22951_
	);
	LUT2 #(
		.INIT('h1)
	) name18905 (
		_w17559_,
		_w22951_,
		_w22952_
	);
	LUT2 #(
		.INIT('h1)
	) name18906 (
		_w17682_,
		_w22952_,
		_w22953_
	);
	LUT2 #(
		.INIT('h1)
	) name18907 (
		_w17565_,
		_w17681_,
		_w22954_
	);
	LUT2 #(
		.INIT('h8)
	) name18908 (
		_w22953_,
		_w22954_,
		_w22955_
	);
	LUT2 #(
		.INIT('h1)
	) name18909 (
		_w22953_,
		_w22954_,
		_w22956_
	);
	LUT2 #(
		.INIT('h1)
	) name18910 (
		_w22955_,
		_w22956_,
		_w22957_
	);
	LUT2 #(
		.INIT('h4)
	) name18911 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22957_,
		_w22958_
	);
	LUT2 #(
		.INIT('h1)
	) name18912 (
		_w22949_,
		_w22958_,
		_w22959_
	);
	LUT2 #(
		.INIT('h8)
	) name18913 (
		_w18262_,
		_w22959_,
		_w22960_
	);
	LUT2 #(
		.INIT('h1)
	) name18914 (
		_w22944_,
		_w22960_,
		_w22961_
	);
	LUT2 #(
		.INIT('h8)
	) name18915 (
		_w7340_,
		_w20401_,
		_w22962_
	);
	LUT2 #(
		.INIT('h4)
	) name18916 (
		\core_eu_ec_cun_TERM_E_reg[3]/P0001 ,
		_w4117_,
		_w22963_
	);
	LUT2 #(
		.INIT('h8)
	) name18917 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001 ,
		_w4845_,
		_w22964_
	);
	LUT2 #(
		.INIT('h8)
	) name18918 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001 ,
		_w4847_,
		_w22965_
	);
	LUT2 #(
		.INIT('h8)
	) name18919 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001 ,
		_w4851_,
		_w22966_
	);
	LUT2 #(
		.INIT('h8)
	) name18920 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001 ,
		_w4849_,
		_w22967_
	);
	LUT2 #(
		.INIT('h1)
	) name18921 (
		_w22964_,
		_w22965_,
		_w22968_
	);
	LUT2 #(
		.INIT('h1)
	) name18922 (
		_w22966_,
		_w22967_,
		_w22969_
	);
	LUT2 #(
		.INIT('h8)
	) name18923 (
		_w22968_,
		_w22969_,
		_w22970_
	);
	LUT2 #(
		.INIT('h4)
	) name18924 (
		_w4117_,
		_w22970_,
		_w22971_
	);
	LUT2 #(
		.INIT('h2)
	) name18925 (
		_w4150_,
		_w22963_,
		_w22972_
	);
	LUT2 #(
		.INIT('h4)
	) name18926 (
		_w22971_,
		_w22972_,
		_w22973_
	);
	LUT2 #(
		.INIT('h4)
	) name18927 (
		\core_eu_ec_cun_TERM_E_reg[2]/P0001 ,
		_w4117_,
		_w22974_
	);
	LUT2 #(
		.INIT('h8)
	) name18928 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001 ,
		_w4845_,
		_w22975_
	);
	LUT2 #(
		.INIT('h8)
	) name18929 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001 ,
		_w4847_,
		_w22976_
	);
	LUT2 #(
		.INIT('h8)
	) name18930 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001 ,
		_w4851_,
		_w22977_
	);
	LUT2 #(
		.INIT('h8)
	) name18931 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001 ,
		_w4849_,
		_w22978_
	);
	LUT2 #(
		.INIT('h1)
	) name18932 (
		_w22975_,
		_w22976_,
		_w22979_
	);
	LUT2 #(
		.INIT('h1)
	) name18933 (
		_w22977_,
		_w22978_,
		_w22980_
	);
	LUT2 #(
		.INIT('h8)
	) name18934 (
		_w22979_,
		_w22980_,
		_w22981_
	);
	LUT2 #(
		.INIT('h4)
	) name18935 (
		_w4117_,
		_w22981_,
		_w22982_
	);
	LUT2 #(
		.INIT('h2)
	) name18936 (
		_w4150_,
		_w22974_,
		_w22983_
	);
	LUT2 #(
		.INIT('h4)
	) name18937 (
		_w22982_,
		_w22983_,
		_w22984_
	);
	LUT2 #(
		.INIT('h1)
	) name18938 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 ,
		_w19499_,
		_w22985_
	);
	LUT2 #(
		.INIT('h2)
	) name18939 (
		_w19499_,
		_w20150_,
		_w22986_
	);
	LUT2 #(
		.INIT('h2)
	) name18940 (
		_w19501_,
		_w22985_,
		_w22987_
	);
	LUT2 #(
		.INIT('h4)
	) name18941 (
		_w22986_,
		_w22987_,
		_w22988_
	);
	LUT2 #(
		.INIT('h2)
	) name18942 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[14]/P0001 ,
		_w19383_,
		_w22989_
	);
	LUT2 #(
		.INIT('h1)
	) name18943 (
		_w19508_,
		_w22989_,
		_w22990_
	);
	LUT2 #(
		.INIT('h4)
	) name18944 (
		_w22988_,
		_w22990_,
		_w22991_
	);
	LUT2 #(
		.INIT('h1)
	) name18945 (
		_w18262_,
		_w22991_,
		_w22992_
	);
	LUT2 #(
		.INIT('h1)
	) name18946 (
		_w17759_,
		_w17768_,
		_w22993_
	);
	LUT2 #(
		.INIT('h4)
	) name18947 (
		_w19372_,
		_w22993_,
		_w22994_
	);
	LUT2 #(
		.INIT('h2)
	) name18948 (
		_w19372_,
		_w22993_,
		_w22995_
	);
	LUT2 #(
		.INIT('h1)
	) name18949 (
		_w22994_,
		_w22995_,
		_w22996_
	);
	LUT2 #(
		.INIT('h4)
	) name18950 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22996_,
		_w22997_
	);
	LUT2 #(
		.INIT('h8)
	) name18951 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19377_,
		_w22998_
	);
	LUT2 #(
		.INIT('h1)
	) name18952 (
		_w22997_,
		_w22998_,
		_w22999_
	);
	LUT2 #(
		.INIT('h2)
	) name18953 (
		_w18262_,
		_w22999_,
		_w23000_
	);
	LUT2 #(
		.INIT('h1)
	) name18954 (
		_w22992_,
		_w23000_,
		_w23001_
	);
	LUT2 #(
		.INIT('h8)
	) name18955 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		_w4117_,
		_w23002_
	);
	LUT2 #(
		.INIT('h1)
	) name18956 (
		_w21257_,
		_w23002_,
		_w23003_
	);
	LUT2 #(
		.INIT('h2)
	) name18957 (
		_w4116_,
		_w23003_,
		_w23004_
	);
	LUT2 #(
		.INIT('h8)
	) name18958 (
		\core_c_dec_imSHT_E_reg/P0001 ,
		_w4117_,
		_w23005_
	);
	LUT2 #(
		.INIT('h8)
	) name18959 (
		_w6119_,
		_w21559_,
		_w23006_
	);
	LUT2 #(
		.INIT('h1)
	) name18960 (
		_w23005_,
		_w23006_,
		_w23007_
	);
	LUT2 #(
		.INIT('h2)
	) name18961 (
		_w4116_,
		_w23007_,
		_w23008_
	);
	LUT2 #(
		.INIT('h8)
	) name18962 (
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w4117_,
		_w23009_
	);
	LUT2 #(
		.INIT('h1)
	) name18963 (
		_w21251_,
		_w23009_,
		_w23010_
	);
	LUT2 #(
		.INIT('h2)
	) name18964 (
		_w4116_,
		_w23010_,
		_w23011_
	);
	LUT2 #(
		.INIT('h2)
	) name18965 (
		_w14752_,
		_w22959_,
		_w23012_
	);
	LUT2 #(
		.INIT('h8)
	) name18966 (
		_w19776_,
		_w19972_,
		_w23013_
	);
	LUT2 #(
		.INIT('h2)
	) name18967 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[7]/P0001 ,
		_w17809_,
		_w23014_
	);
	LUT2 #(
		.INIT('h2)
	) name18968 (
		_w19780_,
		_w23014_,
		_w23015_
	);
	LUT2 #(
		.INIT('h4)
	) name18969 (
		_w23013_,
		_w23015_,
		_w23016_
	);
	LUT2 #(
		.INIT('h1)
	) name18970 (
		_w23012_,
		_w23016_,
		_w23017_
	);
	LUT2 #(
		.INIT('h1)
	) name18971 (
		\sice_GOICE_1_reg/NET0131 ,
		\sice_GOICE_2_reg/NET0131 ,
		_w23018_
	);
	LUT2 #(
		.INIT('h1)
	) name18972 (
		\sice_GOICE_s1_reg/NET0131 ,
		_w23018_,
		_w23019_
	);
	LUT2 #(
		.INIT('h8)
	) name18973 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		_w23020_
	);
	LUT2 #(
		.INIT('h4)
	) name18974 (
		\clkc_RSTtext_reg/P0001 ,
		_w23020_,
		_w23021_
	);
	LUT2 #(
		.INIT('h2)
	) name18975 (
		_w4149_,
		_w23019_,
		_w23022_
	);
	LUT2 #(
		.INIT('h8)
	) name18976 (
		_w23021_,
		_w23022_,
		_w23023_
	);
	LUT2 #(
		.INIT('h1)
	) name18977 (
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w20038_,
		_w23024_
	);
	LUT2 #(
		.INIT('h1)
	) name18978 (
		_w20039_,
		_w23024_,
		_w23025_
	);
	LUT2 #(
		.INIT('h4)
	) name18979 (
		_w13750_,
		_w23025_,
		_w23026_
	);
	LUT2 #(
		.INIT('h2)
	) name18980 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w23027_
	);
	LUT2 #(
		.INIT('h1)
	) name18981 (
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		_w23028_
	);
	LUT2 #(
		.INIT('h8)
	) name18982 (
		_w23027_,
		_w23028_,
		_w23029_
	);
	LUT2 #(
		.INIT('h2)
	) name18983 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		_w23030_
	);
	LUT2 #(
		.INIT('h8)
	) name18984 (
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w23031_
	);
	LUT2 #(
		.INIT('h8)
	) name18985 (
		_w23030_,
		_w23031_,
		_w23032_
	);
	LUT2 #(
		.INIT('h8)
	) name18986 (
		_w23029_,
		_w23032_,
		_w23033_
	);
	LUT2 #(
		.INIT('h4)
	) name18987 (
		\sice_IRST_reg/NET0131 ,
		\sice_SPC_reg[18]/P0001 ,
		_w23034_
	);
	LUT2 #(
		.INIT('h8)
	) name18988 (
		_w23033_,
		_w23034_,
		_w23035_
	);
	LUT2 #(
		.INIT('h4)
	) name18989 (
		\sice_CLR_I_reg/NET0131 ,
		\sice_SPC_reg[21]/P0001 ,
		_w23036_
	);
	LUT2 #(
		.INIT('h8)
	) name18990 (
		_w23033_,
		_w23036_,
		_w23037_
	);
	LUT2 #(
		.INIT('h4)
	) name18991 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18489_,
		_w23038_
	);
	LUT2 #(
		.INIT('h4)
	) name18992 (
		_w18401_,
		_w18405_,
		_w23039_
	);
	LUT2 #(
		.INIT('h1)
	) name18993 (
		_w18406_,
		_w23039_,
		_w23040_
	);
	LUT2 #(
		.INIT('h8)
	) name18994 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23040_,
		_w23041_
	);
	LUT2 #(
		.INIT('h1)
	) name18995 (
		_w23038_,
		_w23041_,
		_w23042_
	);
	LUT2 #(
		.INIT('h2)
	) name18996 (
		_w18457_,
		_w23042_,
		_w23043_
	);
	LUT2 #(
		.INIT('h8)
	) name18997 (
		_w18500_,
		_w18507_,
		_w23044_
	);
	LUT2 #(
		.INIT('h2)
	) name18998 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18492_,
		_w23045_
	);
	LUT2 #(
		.INIT('h8)
	) name18999 (
		_w23044_,
		_w23045_,
		_w23046_
	);
	LUT2 #(
		.INIT('h8)
	) name19000 (
		_w18514_,
		_w23046_,
		_w23047_
	);
	LUT2 #(
		.INIT('h4)
	) name19001 (
		_w23043_,
		_w23047_,
		_w23048_
	);
	LUT2 #(
		.INIT('h8)
	) name19002 (
		_w18500_,
		_w18512_,
		_w23049_
	);
	LUT2 #(
		.INIT('h1)
	) name19003 (
		_w18507_,
		_w23049_,
		_w23050_
	);
	LUT2 #(
		.INIT('h2)
	) name19004 (
		_w18480_,
		_w18512_,
		_w23051_
	);
	LUT2 #(
		.INIT('h4)
	) name19005 (
		_w18507_,
		_w18514_,
		_w23052_
	);
	LUT2 #(
		.INIT('h8)
	) name19006 (
		_w18507_,
		_w18514_,
		_w23053_
	);
	LUT2 #(
		.INIT('h4)
	) name19007 (
		_w18500_,
		_w23053_,
		_w23054_
	);
	LUT2 #(
		.INIT('h4)
	) name19008 (
		_w18396_,
		_w18400_,
		_w23055_
	);
	LUT2 #(
		.INIT('h1)
	) name19009 (
		_w18401_,
		_w23055_,
		_w23056_
	);
	LUT2 #(
		.INIT('h8)
	) name19010 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23056_,
		_w23057_
	);
	LUT2 #(
		.INIT('h4)
	) name19011 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23040_,
		_w23058_
	);
	LUT2 #(
		.INIT('h1)
	) name19012 (
		_w23057_,
		_w23058_,
		_w23059_
	);
	LUT2 #(
		.INIT('h2)
	) name19013 (
		_w18457_,
		_w23059_,
		_w23060_
	);
	LUT2 #(
		.INIT('h8)
	) name19014 (
		_w18501_,
		_w23053_,
		_w23061_
	);
	LUT2 #(
		.INIT('h4)
	) name19015 (
		_w23054_,
		_w23060_,
		_w23062_
	);
	LUT2 #(
		.INIT('h4)
	) name19016 (
		_w23061_,
		_w23062_,
		_w23063_
	);
	LUT2 #(
		.INIT('h8)
	) name19017 (
		_w18500_,
		_w23042_,
		_w23064_
	);
	LUT2 #(
		.INIT('h2)
	) name19018 (
		_w18492_,
		_w23064_,
		_w23065_
	);
	LUT2 #(
		.INIT('h8)
	) name19019 (
		_w23053_,
		_w23065_,
		_w23066_
	);
	LUT2 #(
		.INIT('h1)
	) name19020 (
		_w23063_,
		_w23066_,
		_w23067_
	);
	LUT2 #(
		.INIT('h1)
	) name19021 (
		_w23051_,
		_w23052_,
		_w23068_
	);
	LUT2 #(
		.INIT('h4)
	) name19022 (
		_w23067_,
		_w23068_,
		_w23069_
	);
	LUT2 #(
		.INIT('h1)
	) name19023 (
		_w23050_,
		_w23069_,
		_w23070_
	);
	LUT2 #(
		.INIT('h2)
	) name19024 (
		_w18479_,
		_w23070_,
		_w23071_
	);
	LUT2 #(
		.INIT('h2)
	) name19025 (
		_w18471_,
		_w23071_,
		_w23072_
	);
	LUT2 #(
		.INIT('h1)
	) name19026 (
		_w18481_,
		_w23072_,
		_w23073_
	);
	LUT2 #(
		.INIT('h2)
	) name19027 (
		_w18479_,
		_w23073_,
		_w23074_
	);
	LUT2 #(
		.INIT('h8)
	) name19028 (
		_w18512_,
		_w23072_,
		_w23075_
	);
	LUT2 #(
		.INIT('h1)
	) name19029 (
		_w23074_,
		_w23075_,
		_w23076_
	);
	LUT2 #(
		.INIT('h1)
	) name19030 (
		_w23047_,
		_w23076_,
		_w23077_
	);
	LUT2 #(
		.INIT('h2)
	) name19031 (
		_w18467_,
		_w18470_,
		_w23078_
	);
	LUT2 #(
		.INIT('h1)
	) name19032 (
		_w23048_,
		_w23078_,
		_w23079_
	);
	LUT2 #(
		.INIT('h4)
	) name19033 (
		_w23077_,
		_w23079_,
		_w23080_
	);
	LUT2 #(
		.INIT('h1)
	) name19034 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23080_,
		_w23081_
	);
	LUT2 #(
		.INIT('h8)
	) name19035 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23080_,
		_w23082_
	);
	LUT2 #(
		.INIT('h1)
	) name19036 (
		_w23081_,
		_w23082_,
		_w23083_
	);
	LUT2 #(
		.INIT('h2)
	) name19037 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w23083_,
		_w23084_
	);
	LUT2 #(
		.INIT('h4)
	) name19038 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w8113_,
		_w23085_
	);
	LUT2 #(
		.INIT('h1)
	) name19039 (
		_w23084_,
		_w23085_,
		_w23086_
	);
	LUT2 #(
		.INIT('h1)
	) name19040 (
		_w21318_,
		_w23086_,
		_w23087_
	);
	LUT2 #(
		.INIT('h8)
	) name19041 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w21318_,
		_w23088_
	);
	LUT2 #(
		.INIT('h1)
	) name19042 (
		_w23087_,
		_w23088_,
		_w23089_
	);
	LUT2 #(
		.INIT('h4)
	) name19043 (
		\sice_CLR_M_reg/NET0131 ,
		\sice_SPC_reg[22]/P0001 ,
		_w23090_
	);
	LUT2 #(
		.INIT('h8)
	) name19044 (
		_w23033_,
		_w23090_,
		_w23091_
	);
	LUT2 #(
		.INIT('h8)
	) name19045 (
		\clkc_OSCoff_set_reg/P0001 ,
		\clkc_SLEEP_reg/NET0131 ,
		_w23092_
	);
	LUT2 #(
		.INIT('h1)
	) name19046 (
		\clkc_OSCoff_reg/NET0131 ,
		_w23092_,
		_w23093_
	);
	LUT2 #(
		.INIT('h8)
	) name19047 (
		\pio_PINT_reg[3]/NET0131 ,
		\pio_pmask_reg_DO_reg[3]/NET0131 ,
		_w23094_
	);
	LUT2 #(
		.INIT('h8)
	) name19048 (
		\pio_PINT_reg[8]/NET0131 ,
		\pio_pmask_reg_DO_reg[8]/NET0131 ,
		_w23095_
	);
	LUT2 #(
		.INIT('h8)
	) name19049 (
		\pio_PINT_reg[7]/NET0131 ,
		\pio_pmask_reg_DO_reg[7]/NET0131 ,
		_w23096_
	);
	LUT2 #(
		.INIT('h8)
	) name19050 (
		\pio_PINT_reg[1]/NET0131 ,
		\pio_pmask_reg_DO_reg[1]/NET0131 ,
		_w23097_
	);
	LUT2 #(
		.INIT('h8)
	) name19051 (
		\pio_PINT_reg[6]/NET0131 ,
		\pio_pmask_reg_DO_reg[6]/NET0131 ,
		_w23098_
	);
	LUT2 #(
		.INIT('h8)
	) name19052 (
		\pio_PINT_reg[10]/NET0131 ,
		\pio_pmask_reg_DO_reg[10]/NET0131 ,
		_w23099_
	);
	LUT2 #(
		.INIT('h8)
	) name19053 (
		\pio_PINT_reg[4]/NET0131 ,
		\pio_pmask_reg_DO_reg[4]/NET0131 ,
		_w23100_
	);
	LUT2 #(
		.INIT('h8)
	) name19054 (
		\pio_PINT_reg[0]/NET0131 ,
		\pio_pmask_reg_DO_reg[0]/NET0131 ,
		_w23101_
	);
	LUT2 #(
		.INIT('h8)
	) name19055 (
		\pio_PINT_reg[5]/NET0131 ,
		\pio_pmask_reg_DO_reg[5]/NET0131 ,
		_w23102_
	);
	LUT2 #(
		.INIT('h8)
	) name19056 (
		\pio_PINT_reg[11]/NET0131 ,
		\pio_pmask_reg_DO_reg[11]/NET0131 ,
		_w23103_
	);
	LUT2 #(
		.INIT('h8)
	) name19057 (
		\pio_PINT_reg[2]/NET0131 ,
		\pio_pmask_reg_DO_reg[2]/NET0131 ,
		_w23104_
	);
	LUT2 #(
		.INIT('h8)
	) name19058 (
		\pio_PINT_reg[9]/NET0131 ,
		\pio_pmask_reg_DO_reg[9]/NET0131 ,
		_w23105_
	);
	LUT2 #(
		.INIT('h1)
	) name19059 (
		_w23094_,
		_w23095_,
		_w23106_
	);
	LUT2 #(
		.INIT('h1)
	) name19060 (
		_w23096_,
		_w23097_,
		_w23107_
	);
	LUT2 #(
		.INIT('h1)
	) name19061 (
		_w23098_,
		_w23099_,
		_w23108_
	);
	LUT2 #(
		.INIT('h1)
	) name19062 (
		_w23100_,
		_w23101_,
		_w23109_
	);
	LUT2 #(
		.INIT('h1)
	) name19063 (
		_w23102_,
		_w23103_,
		_w23110_
	);
	LUT2 #(
		.INIT('h1)
	) name19064 (
		_w23104_,
		_w23105_,
		_w23111_
	);
	LUT2 #(
		.INIT('h8)
	) name19065 (
		_w23110_,
		_w23111_,
		_w23112_
	);
	LUT2 #(
		.INIT('h8)
	) name19066 (
		_w23108_,
		_w23109_,
		_w23113_
	);
	LUT2 #(
		.INIT('h8)
	) name19067 (
		_w23106_,
		_w23107_,
		_w23114_
	);
	LUT2 #(
		.INIT('h8)
	) name19068 (
		_w23113_,
		_w23114_,
		_w23115_
	);
	LUT2 #(
		.INIT('h8)
	) name19069 (
		_w23112_,
		_w23115_,
		_w23116_
	);
	LUT2 #(
		.INIT('h2)
	) name19070 (
		_w4149_,
		_w20357_,
		_w23117_
	);
	LUT2 #(
		.INIT('h1)
	) name19071 (
		\tm_WR_TCR_KEEP_TO_TMCLK_p_reg/NET0131 ,
		\tm_WR_TCR_p_reg/P0001 ,
		_w23118_
	);
	LUT2 #(
		.INIT('h8)
	) name19072 (
		_w14752_,
		_w22999_,
		_w23119_
	);
	LUT2 #(
		.INIT('h8)
	) name19073 (
		_w19776_,
		_w20150_,
		_w23120_
	);
	LUT2 #(
		.INIT('h2)
	) name19074 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[14]/P0001 ,
		_w17809_,
		_w23121_
	);
	LUT2 #(
		.INIT('h2)
	) name19075 (
		_w19780_,
		_w23121_,
		_w23122_
	);
	LUT2 #(
		.INIT('h4)
	) name19076 (
		_w23120_,
		_w23122_,
		_w23123_
	);
	LUT2 #(
		.INIT('h1)
	) name19077 (
		_w23119_,
		_w23123_,
		_w23124_
	);
	LUT2 #(
		.INIT('h4)
	) name19078 (
		\core_eu_ec_cun_TERM_E_reg[1]/P0001 ,
		_w4117_,
		_w23125_
	);
	LUT2 #(
		.INIT('h8)
	) name19079 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001 ,
		_w4849_,
		_w23126_
	);
	LUT2 #(
		.INIT('h8)
	) name19080 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001 ,
		_w4851_,
		_w23127_
	);
	LUT2 #(
		.INIT('h8)
	) name19081 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001 ,
		_w4847_,
		_w23128_
	);
	LUT2 #(
		.INIT('h8)
	) name19082 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001 ,
		_w4845_,
		_w23129_
	);
	LUT2 #(
		.INIT('h1)
	) name19083 (
		_w23126_,
		_w23127_,
		_w23130_
	);
	LUT2 #(
		.INIT('h1)
	) name19084 (
		_w23128_,
		_w23129_,
		_w23131_
	);
	LUT2 #(
		.INIT('h8)
	) name19085 (
		_w23130_,
		_w23131_,
		_w23132_
	);
	LUT2 #(
		.INIT('h4)
	) name19086 (
		_w4117_,
		_w23132_,
		_w23133_
	);
	LUT2 #(
		.INIT('h2)
	) name19087 (
		_w4150_,
		_w23125_,
		_w23134_
	);
	LUT2 #(
		.INIT('h4)
	) name19088 (
		_w23133_,
		_w23134_,
		_w23135_
	);
	LUT2 #(
		.INIT('h4)
	) name19089 (
		\core_eu_ec_cun_TERM_E_reg[0]/P0001 ,
		_w4117_,
		_w23136_
	);
	LUT2 #(
		.INIT('h8)
	) name19090 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001 ,
		_w4845_,
		_w23137_
	);
	LUT2 #(
		.INIT('h8)
	) name19091 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001 ,
		_w4847_,
		_w23138_
	);
	LUT2 #(
		.INIT('h8)
	) name19092 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001 ,
		_w4851_,
		_w23139_
	);
	LUT2 #(
		.INIT('h8)
	) name19093 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001 ,
		_w4849_,
		_w23140_
	);
	LUT2 #(
		.INIT('h1)
	) name19094 (
		_w23137_,
		_w23138_,
		_w23141_
	);
	LUT2 #(
		.INIT('h1)
	) name19095 (
		_w23139_,
		_w23140_,
		_w23142_
	);
	LUT2 #(
		.INIT('h8)
	) name19096 (
		_w23141_,
		_w23142_,
		_w23143_
	);
	LUT2 #(
		.INIT('h4)
	) name19097 (
		_w4117_,
		_w23143_,
		_w23144_
	);
	LUT2 #(
		.INIT('h2)
	) name19098 (
		_w4150_,
		_w23136_,
		_w23145_
	);
	LUT2 #(
		.INIT('h4)
	) name19099 (
		_w23144_,
		_w23145_,
		_w23146_
	);
	LUT2 #(
		.INIT('h2)
	) name19100 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18395_,
		_w23147_
	);
	LUT2 #(
		.INIT('h4)
	) name19101 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23056_,
		_w23148_
	);
	LUT2 #(
		.INIT('h1)
	) name19102 (
		_w23147_,
		_w23148_,
		_w23149_
	);
	LUT2 #(
		.INIT('h2)
	) name19103 (
		_w18457_,
		_w23149_,
		_w23150_
	);
	LUT2 #(
		.INIT('h2)
	) name19104 (
		_w23047_,
		_w23150_,
		_w23151_
	);
	LUT2 #(
		.INIT('h8)
	) name19105 (
		_w18481_,
		_w18507_,
		_w23152_
	);
	LUT2 #(
		.INIT('h1)
	) name19106 (
		_w18479_,
		_w18500_,
		_w23153_
	);
	LUT2 #(
		.INIT('h4)
	) name19107 (
		_w18492_,
		_w23051_,
		_w23154_
	);
	LUT2 #(
		.INIT('h8)
	) name19108 (
		_w23043_,
		_w23052_,
		_w23155_
	);
	LUT2 #(
		.INIT('h2)
	) name19109 (
		_w23054_,
		_w23060_,
		_w23156_
	);
	LUT2 #(
		.INIT('h8)
	) name19110 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w18390_,
		_w23157_
	);
	LUT2 #(
		.INIT('h4)
	) name19111 (
		_w18392_,
		_w18395_,
		_w23158_
	);
	LUT2 #(
		.INIT('h1)
	) name19112 (
		_w18396_,
		_w23158_,
		_w23159_
	);
	LUT2 #(
		.INIT('h1)
	) name19113 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23159_,
		_w23160_
	);
	LUT2 #(
		.INIT('h1)
	) name19114 (
		_w23157_,
		_w23160_,
		_w23161_
	);
	LUT2 #(
		.INIT('h8)
	) name19115 (
		_w18457_,
		_w23161_,
		_w23162_
	);
	LUT2 #(
		.INIT('h1)
	) name19116 (
		_w23061_,
		_w23162_,
		_w23163_
	);
	LUT2 #(
		.INIT('h2)
	) name19117 (
		_w23061_,
		_w23150_,
		_w23164_
	);
	LUT2 #(
		.INIT('h1)
	) name19118 (
		_w23163_,
		_w23164_,
		_w23165_
	);
	LUT2 #(
		.INIT('h1)
	) name19119 (
		_w23054_,
		_w23165_,
		_w23166_
	);
	LUT2 #(
		.INIT('h1)
	) name19120 (
		_w23052_,
		_w23156_,
		_w23167_
	);
	LUT2 #(
		.INIT('h4)
	) name19121 (
		_w23166_,
		_w23167_,
		_w23168_
	);
	LUT2 #(
		.INIT('h1)
	) name19122 (
		_w23051_,
		_w23155_,
		_w23169_
	);
	LUT2 #(
		.INIT('h4)
	) name19123 (
		_w23168_,
		_w23169_,
		_w23170_
	);
	LUT2 #(
		.INIT('h2)
	) name19124 (
		_w18479_,
		_w23154_,
		_w23171_
	);
	LUT2 #(
		.INIT('h4)
	) name19125 (
		_w23170_,
		_w23171_,
		_w23172_
	);
	LUT2 #(
		.INIT('h2)
	) name19126 (
		_w18471_,
		_w23153_,
		_w23173_
	);
	LUT2 #(
		.INIT('h4)
	) name19127 (
		_w23172_,
		_w23173_,
		_w23174_
	);
	LUT2 #(
		.INIT('h1)
	) name19128 (
		_w23152_,
		_w23174_,
		_w23175_
	);
	LUT2 #(
		.INIT('h1)
	) name19129 (
		_w23047_,
		_w23175_,
		_w23176_
	);
	LUT2 #(
		.INIT('h4)
	) name19130 (
		_w18470_,
		_w18512_,
		_w23177_
	);
	LUT2 #(
		.INIT('h1)
	) name19131 (
		_w23151_,
		_w23177_,
		_w23178_
	);
	LUT2 #(
		.INIT('h4)
	) name19132 (
		_w23176_,
		_w23178_,
		_w23179_
	);
	LUT2 #(
		.INIT('h1)
	) name19133 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23179_,
		_w23180_
	);
	LUT2 #(
		.INIT('h8)
	) name19134 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w23179_,
		_w23181_
	);
	LUT2 #(
		.INIT('h1)
	) name19135 (
		_w23180_,
		_w23181_,
		_w23182_
	);
	LUT2 #(
		.INIT('h2)
	) name19136 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w23182_,
		_w23183_
	);
	LUT2 #(
		.INIT('h4)
	) name19137 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w9435_,
		_w23184_
	);
	LUT2 #(
		.INIT('h1)
	) name19138 (
		_w23183_,
		_w23184_,
		_w23185_
	);
	LUT2 #(
		.INIT('h1)
	) name19139 (
		_w21318_,
		_w23185_,
		_w23186_
	);
	LUT2 #(
		.INIT('h8)
	) name19140 (
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w21318_,
		_w23187_
	);
	LUT2 #(
		.INIT('h1)
	) name19141 (
		_w23186_,
		_w23187_,
		_w23188_
	);
	LUT2 #(
		.INIT('h4)
	) name19142 (
		\sport0_rxctl_RXSHT_reg[3]/P0001 ,
		_w20868_,
		_w23189_
	);
	LUT2 #(
		.INIT('h8)
	) name19143 (
		\sport0_rxctl_RX_reg[3]/P0001 ,
		_w20873_,
		_w23190_
	);
	LUT2 #(
		.INIT('h4)
	) name19144 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w8113_,
		_w23191_
	);
	LUT2 #(
		.INIT('h1)
	) name19145 (
		_w20903_,
		_w20921_,
		_w23192_
	);
	LUT2 #(
		.INIT('h1)
	) name19146 (
		_w20922_,
		_w23192_,
		_w23193_
	);
	LUT2 #(
		.INIT('h1)
	) name19147 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w20955_,
		_w23194_
	);
	LUT2 #(
		.INIT('h2)
	) name19148 (
		_w23193_,
		_w23194_,
		_w23195_
	);
	LUT2 #(
		.INIT('h4)
	) name19149 (
		_w23193_,
		_w23194_,
		_w23196_
	);
	LUT2 #(
		.INIT('h2)
	) name19150 (
		_w20875_,
		_w23195_,
		_w23197_
	);
	LUT2 #(
		.INIT('h4)
	) name19151 (
		_w23196_,
		_w23197_,
		_w23198_
	);
	LUT2 #(
		.INIT('h1)
	) name19152 (
		_w20868_,
		_w23190_,
		_w23199_
	);
	LUT2 #(
		.INIT('h4)
	) name19153 (
		_w23198_,
		_w23199_,
		_w23200_
	);
	LUT2 #(
		.INIT('h4)
	) name19154 (
		_w23191_,
		_w23200_,
		_w23201_
	);
	LUT2 #(
		.INIT('h1)
	) name19155 (
		_w20871_,
		_w23189_,
		_w23202_
	);
	LUT2 #(
		.INIT('h4)
	) name19156 (
		_w23201_,
		_w23202_,
		_w23203_
	);
	LUT2 #(
		.INIT('h8)
	) name19157 (
		\sport0_rxctl_RX_reg[3]/P0001 ,
		_w20871_,
		_w23204_
	);
	LUT2 #(
		.INIT('h1)
	) name19158 (
		_w23203_,
		_w23204_,
		_w23205_
	);
	LUT2 #(
		.INIT('h1)
	) name19159 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 ,
		_w19499_,
		_w23206_
	);
	LUT2 #(
		.INIT('h4)
	) name19160 (
		_w18276_,
		_w19499_,
		_w23207_
	);
	LUT2 #(
		.INIT('h2)
	) name19161 (
		_w19501_,
		_w23206_,
		_w23208_
	);
	LUT2 #(
		.INIT('h4)
	) name19162 (
		_w23207_,
		_w23208_,
		_w23209_
	);
	LUT2 #(
		.INIT('h2)
	) name19163 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[6]/P0001 ,
		_w19383_,
		_w23210_
	);
	LUT2 #(
		.INIT('h1)
	) name19164 (
		_w19508_,
		_w23210_,
		_w23211_
	);
	LUT2 #(
		.INIT('h4)
	) name19165 (
		_w23209_,
		_w23211_,
		_w23212_
	);
	LUT2 #(
		.INIT('h1)
	) name19166 (
		_w18262_,
		_w23212_,
		_w23213_
	);
	LUT2 #(
		.INIT('h2)
	) name19167 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22957_,
		_w23214_
	);
	LUT2 #(
		.INIT('h1)
	) name19168 (
		_w17559_,
		_w17682_,
		_w23215_
	);
	LUT2 #(
		.INIT('h2)
	) name19169 (
		_w22951_,
		_w23215_,
		_w23216_
	);
	LUT2 #(
		.INIT('h4)
	) name19170 (
		_w22951_,
		_w23215_,
		_w23217_
	);
	LUT2 #(
		.INIT('h1)
	) name19171 (
		_w23216_,
		_w23217_,
		_w23218_
	);
	LUT2 #(
		.INIT('h4)
	) name19172 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w23218_,
		_w23219_
	);
	LUT2 #(
		.INIT('h1)
	) name19173 (
		_w23214_,
		_w23219_,
		_w23220_
	);
	LUT2 #(
		.INIT('h2)
	) name19174 (
		_w18262_,
		_w23220_,
		_w23221_
	);
	LUT2 #(
		.INIT('h1)
	) name19175 (
		_w23213_,
		_w23221_,
		_w23222_
	);
	LUT2 #(
		.INIT('h8)
	) name19176 (
		_w14752_,
		_w23220_,
		_w23223_
	);
	LUT2 #(
		.INIT('h8)
	) name19177 (
		_w18276_,
		_w19776_,
		_w23224_
	);
	LUT2 #(
		.INIT('h2)
	) name19178 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[6]/P0001 ,
		_w17809_,
		_w23225_
	);
	LUT2 #(
		.INIT('h2)
	) name19179 (
		_w19780_,
		_w23225_,
		_w23226_
	);
	LUT2 #(
		.INIT('h4)
	) name19180 (
		_w23224_,
		_w23226_,
		_w23227_
	);
	LUT2 #(
		.INIT('h1)
	) name19181 (
		_w23223_,
		_w23227_,
		_w23228_
	);
	LUT2 #(
		.INIT('h8)
	) name19182 (
		\core_c_dec_IDLE_Eg_reg/P0001 ,
		_w4118_,
		_w23229_
	);
	LUT2 #(
		.INIT('h8)
	) name19183 (
		_w6024_,
		_w21249_,
		_w23230_
	);
	LUT2 #(
		.INIT('h8)
	) name19184 (
		_w11741_,
		_w21421_,
		_w23231_
	);
	LUT2 #(
		.INIT('h4)
	) name19185 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w23230_,
		_w23232_
	);
	LUT2 #(
		.INIT('h8)
	) name19186 (
		_w23231_,
		_w23232_,
		_w23233_
	);
	LUT2 #(
		.INIT('h1)
	) name19187 (
		_w23229_,
		_w23233_,
		_w23234_
	);
	LUT2 #(
		.INIT('h8)
	) name19188 (
		_w4117_,
		_w5696_,
		_w23235_
	);
	LUT2 #(
		.INIT('h8)
	) name19189 (
		\memc_ldSREG_E_reg/NET0131 ,
		_w23235_,
		_w23236_
	);
	LUT2 #(
		.INIT('h2)
	) name19190 (
		_w11751_,
		_w11753_,
		_w23237_
	);
	LUT2 #(
		.INIT('h2)
	) name19191 (
		_w11734_,
		_w23235_,
		_w23238_
	);
	LUT2 #(
		.INIT('h4)
	) name19192 (
		_w23237_,
		_w23238_,
		_w23239_
	);
	LUT2 #(
		.INIT('h1)
	) name19193 (
		_w23236_,
		_w23239_,
		_w23240_
	);
	LUT2 #(
		.INIT('h1)
	) name19194 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w23241_
	);
	LUT2 #(
		.INIT('h4)
	) name19195 (
		_w14697_,
		_w23241_,
		_w23242_
	);
	LUT2 #(
		.INIT('h1)
	) name19196 (
		_w5950_,
		_w23242_,
		_w23243_
	);
	LUT2 #(
		.INIT('h2)
	) name19197 (
		_w14273_,
		_w14406_,
		_w23244_
	);
	LUT2 #(
		.INIT('h4)
	) name19198 (
		_w14273_,
		_w14404_,
		_w23245_
	);
	LUT2 #(
		.INIT('h1)
	) name19199 (
		_w13972_,
		_w23244_,
		_w23246_
	);
	LUT2 #(
		.INIT('h4)
	) name19200 (
		_w23245_,
		_w23246_,
		_w23247_
	);
	LUT2 #(
		.INIT('h2)
	) name19201 (
		_w14270_,
		_w14274_,
		_w23248_
	);
	LUT2 #(
		.INIT('h1)
	) name19202 (
		_w13809_,
		_w14010_,
		_w23249_
	);
	LUT2 #(
		.INIT('h4)
	) name19203 (
		_w23248_,
		_w23249_,
		_w23250_
	);
	LUT2 #(
		.INIT('h4)
	) name19204 (
		_w23247_,
		_w23250_,
		_w23251_
	);
	LUT2 #(
		.INIT('h2)
	) name19205 (
		_w23247_,
		_w23250_,
		_w23252_
	);
	LUT2 #(
		.INIT('h1)
	) name19206 (
		_w23251_,
		_w23252_,
		_w23253_
	);
	LUT2 #(
		.INIT('h2)
	) name19207 (
		_w13806_,
		_w23253_,
		_w23254_
	);
	LUT2 #(
		.INIT('h1)
	) name19208 (
		_w13806_,
		_w14658_,
		_w23255_
	);
	LUT2 #(
		.INIT('h1)
	) name19209 (
		_w23254_,
		_w23255_,
		_w23256_
	);
	LUT2 #(
		.INIT('h2)
	) name19210 (
		_w14667_,
		_w23256_,
		_w23257_
	);
	LUT2 #(
		.INIT('h2)
	) name19211 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[8]/P0001 ,
		_w14667_,
		_w23258_
	);
	LUT2 #(
		.INIT('h1)
	) name19212 (
		_w23257_,
		_w23258_,
		_w23259_
	);
	LUT2 #(
		.INIT('h2)
	) name19213 (
		_w13805_,
		_w23256_,
		_w23260_
	);
	LUT2 #(
		.INIT('h2)
	) name19214 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[8]/P0001 ,
		_w13805_,
		_w23261_
	);
	LUT2 #(
		.INIT('h1)
	) name19215 (
		_w23260_,
		_w23261_,
		_w23262_
	);
	LUT2 #(
		.INIT('h1)
	) name19216 (
		_w22669_,
		_w22671_,
		_w23263_
	);
	LUT2 #(
		.INIT('h8)
	) name19217 (
		_w22671_,
		_w22675_,
		_w23264_
	);
	LUT2 #(
		.INIT('h1)
	) name19218 (
		_w23263_,
		_w23264_,
		_w23265_
	);
	LUT2 #(
		.INIT('h1)
	) name19219 (
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		\sport1_txctl_Wcnt_reg[1]/NET0131 ,
		_w23266_
	);
	LUT2 #(
		.INIT('h1)
	) name19220 (
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		_w23267_
	);
	LUT2 #(
		.INIT('h1)
	) name19221 (
		\sport1_txctl_Wcnt_reg[4]/NET0131 ,
		\sport1_txctl_Wcnt_reg[5]/NET0131 ,
		_w23268_
	);
	LUT2 #(
		.INIT('h1)
	) name19222 (
		\sport1_txctl_Wcnt_reg[6]/NET0131 ,
		\sport1_txctl_Wcnt_reg[7]/NET0131 ,
		_w23269_
	);
	LUT2 #(
		.INIT('h8)
	) name19223 (
		_w23268_,
		_w23269_,
		_w23270_
	);
	LUT2 #(
		.INIT('h8)
	) name19224 (
		_w23266_,
		_w23267_,
		_w23271_
	);
	LUT2 #(
		.INIT('h8)
	) name19225 (
		_w23270_,
		_w23271_,
		_w23272_
	);
	LUT2 #(
		.INIT('h1)
	) name19226 (
		_w23263_,
		_w23272_,
		_w23273_
	);
	LUT2 #(
		.INIT('h1)
	) name19227 (
		_w23265_,
		_w23273_,
		_w23274_
	);
	LUT2 #(
		.INIT('h1)
	) name19228 (
		_w19952_,
		_w19954_,
		_w23275_
	);
	LUT2 #(
		.INIT('h8)
	) name19229 (
		_w19954_,
		_w19958_,
		_w23276_
	);
	LUT2 #(
		.INIT('h1)
	) name19230 (
		_w23275_,
		_w23276_,
		_w23277_
	);
	LUT2 #(
		.INIT('h1)
	) name19231 (
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		\sport0_txctl_Wcnt_reg[1]/NET0131 ,
		_w23278_
	);
	LUT2 #(
		.INIT('h1)
	) name19232 (
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		_w23279_
	);
	LUT2 #(
		.INIT('h1)
	) name19233 (
		\sport0_txctl_Wcnt_reg[4]/NET0131 ,
		\sport0_txctl_Wcnt_reg[5]/NET0131 ,
		_w23280_
	);
	LUT2 #(
		.INIT('h1)
	) name19234 (
		\sport0_txctl_Wcnt_reg[6]/NET0131 ,
		\sport0_txctl_Wcnt_reg[7]/NET0131 ,
		_w23281_
	);
	LUT2 #(
		.INIT('h8)
	) name19235 (
		_w23280_,
		_w23281_,
		_w23282_
	);
	LUT2 #(
		.INIT('h8)
	) name19236 (
		_w23278_,
		_w23279_,
		_w23283_
	);
	LUT2 #(
		.INIT('h8)
	) name19237 (
		_w23282_,
		_w23283_,
		_w23284_
	);
	LUT2 #(
		.INIT('h1)
	) name19238 (
		_w23275_,
		_w23284_,
		_w23285_
	);
	LUT2 #(
		.INIT('h1)
	) name19239 (
		_w23277_,
		_w23285_,
		_w23286_
	);
	LUT2 #(
		.INIT('h2)
	) name19240 (
		\core_c_psq_SSTAT_reg[6]/NET0131 ,
		_w20574_,
		_w23287_
	);
	LUT2 #(
		.INIT('h1)
	) name19241 (
		_w20578_,
		_w23287_,
		_w23288_
	);
	LUT2 #(
		.INIT('h4)
	) name19242 (
		_w4845_,
		_w20579_,
		_w23289_
	);
	LUT2 #(
		.INIT('h1)
	) name19243 (
		_w23288_,
		_w23289_,
		_w23290_
	);
	LUT2 #(
		.INIT('h2)
	) name19244 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w21242_,
		_w23291_
	);
	LUT2 #(
		.INIT('h8)
	) name19245 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w21242_,
		_w23292_
	);
	LUT2 #(
		.INIT('h1)
	) name19246 (
		_w23291_,
		_w23292_,
		_w23293_
	);
	LUT2 #(
		.INIT('h2)
	) name19247 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w21242_,
		_w23294_
	);
	LUT2 #(
		.INIT('h8)
	) name19248 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w21242_,
		_w23295_
	);
	LUT2 #(
		.INIT('h1)
	) name19249 (
		_w23294_,
		_w23295_,
		_w23296_
	);
	LUT2 #(
		.INIT('h2)
	) name19250 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w21242_,
		_w23297_
	);
	LUT2 #(
		.INIT('h8)
	) name19251 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w21242_,
		_w23298_
	);
	LUT2 #(
		.INIT('h1)
	) name19252 (
		_w23297_,
		_w23298_,
		_w23299_
	);
	LUT2 #(
		.INIT('h2)
	) name19253 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w21242_,
		_w23300_
	);
	LUT2 #(
		.INIT('h8)
	) name19254 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w21242_,
		_w23301_
	);
	LUT2 #(
		.INIT('h1)
	) name19255 (
		_w23300_,
		_w23301_,
		_w23302_
	);
	LUT2 #(
		.INIT('h2)
	) name19256 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w21242_,
		_w23303_
	);
	LUT2 #(
		.INIT('h8)
	) name19257 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w21242_,
		_w23304_
	);
	LUT2 #(
		.INIT('h1)
	) name19258 (
		_w23303_,
		_w23304_,
		_w23305_
	);
	LUT2 #(
		.INIT('h2)
	) name19259 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w21242_,
		_w23306_
	);
	LUT2 #(
		.INIT('h8)
	) name19260 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w21242_,
		_w23307_
	);
	LUT2 #(
		.INIT('h1)
	) name19261 (
		_w23306_,
		_w23307_,
		_w23308_
	);
	LUT2 #(
		.INIT('h2)
	) name19262 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w21242_,
		_w23309_
	);
	LUT2 #(
		.INIT('h8)
	) name19263 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w21242_,
		_w23310_
	);
	LUT2 #(
		.INIT('h1)
	) name19264 (
		_w23309_,
		_w23310_,
		_w23311_
	);
	LUT2 #(
		.INIT('h2)
	) name19265 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w21242_,
		_w23312_
	);
	LUT2 #(
		.INIT('h8)
	) name19266 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w21242_,
		_w23313_
	);
	LUT2 #(
		.INIT('h1)
	) name19267 (
		_w23312_,
		_w23313_,
		_w23314_
	);
	LUT2 #(
		.INIT('h2)
	) name19268 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w21242_,
		_w23315_
	);
	LUT2 #(
		.INIT('h8)
	) name19269 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w21242_,
		_w23316_
	);
	LUT2 #(
		.INIT('h1)
	) name19270 (
		_w23315_,
		_w23316_,
		_w23317_
	);
	LUT2 #(
		.INIT('h2)
	) name19271 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w21242_,
		_w23318_
	);
	LUT2 #(
		.INIT('h8)
	) name19272 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w21242_,
		_w23319_
	);
	LUT2 #(
		.INIT('h1)
	) name19273 (
		_w23318_,
		_w23319_,
		_w23320_
	);
	LUT2 #(
		.INIT('h2)
	) name19274 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w21242_,
		_w23321_
	);
	LUT2 #(
		.INIT('h8)
	) name19275 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w21242_,
		_w23322_
	);
	LUT2 #(
		.INIT('h1)
	) name19276 (
		_w23321_,
		_w23322_,
		_w23323_
	);
	LUT2 #(
		.INIT('h2)
	) name19277 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w21242_,
		_w23324_
	);
	LUT2 #(
		.INIT('h8)
	) name19278 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w21242_,
		_w23325_
	);
	LUT2 #(
		.INIT('h1)
	) name19279 (
		_w23324_,
		_w23325_,
		_w23326_
	);
	LUT2 #(
		.INIT('h2)
	) name19280 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w21242_,
		_w23327_
	);
	LUT2 #(
		.INIT('h8)
	) name19281 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w21242_,
		_w23328_
	);
	LUT2 #(
		.INIT('h1)
	) name19282 (
		_w23327_,
		_w23328_,
		_w23329_
	);
	LUT2 #(
		.INIT('h2)
	) name19283 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w21242_,
		_w23330_
	);
	LUT2 #(
		.INIT('h8)
	) name19284 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w21242_,
		_w23331_
	);
	LUT2 #(
		.INIT('h1)
	) name19285 (
		_w23330_,
		_w23331_,
		_w23332_
	);
	LUT2 #(
		.INIT('h8)
	) name19286 (
		\core_c_dec_Post1_E_reg/P0001 ,
		_w4118_,
		_w23333_
	);
	LUT2 #(
		.INIT('h2)
	) name19287 (
		_w21421_,
		_w21590_,
		_w23334_
	);
	LUT2 #(
		.INIT('h1)
	) name19288 (
		_w23333_,
		_w23334_,
		_w23335_
	);
	LUT2 #(
		.INIT('h1)
	) name19289 (
		_w4117_,
		_w19702_,
		_w23336_
	);
	LUT2 #(
		.INIT('h2)
	) name19290 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		_w23336_,
		_w23337_
	);
	LUT2 #(
		.INIT('h4)
	) name19291 (
		_w20687_,
		_w23336_,
		_w23338_
	);
	LUT2 #(
		.INIT('h1)
	) name19292 (
		_w23337_,
		_w23338_,
		_w23339_
	);
	LUT2 #(
		.INIT('h2)
	) name19293 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w23336_,
		_w23340_
	);
	LUT2 #(
		.INIT('h4)
	) name19294 (
		_w20698_,
		_w23336_,
		_w23341_
	);
	LUT2 #(
		.INIT('h1)
	) name19295 (
		_w23340_,
		_w23341_,
		_w23342_
	);
	LUT2 #(
		.INIT('h1)
	) name19296 (
		_w4057_,
		_w5950_,
		_w23343_
	);
	LUT2 #(
		.INIT('h4)
	) name19297 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		_w23344_
	);
	LUT2 #(
		.INIT('h8)
	) name19298 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		_w23345_
	);
	LUT2 #(
		.INIT('h1)
	) name19299 (
		_w23344_,
		_w23345_,
		_w23346_
	);
	LUT2 #(
		.INIT('h2)
	) name19300 (
		_w23343_,
		_w23346_,
		_w23347_
	);
	LUT2 #(
		.INIT('h2)
	) name19301 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[9]/NET0131 ,
		_w23343_,
		_w23348_
	);
	LUT2 #(
		.INIT('h1)
	) name19302 (
		_w23347_,
		_w23348_,
		_w23349_
	);
	LUT2 #(
		.INIT('h4)
	) name19303 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		_w23350_
	);
	LUT2 #(
		.INIT('h8)
	) name19304 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		_w23351_
	);
	LUT2 #(
		.INIT('h1)
	) name19305 (
		_w23350_,
		_w23351_,
		_w23352_
	);
	LUT2 #(
		.INIT('h2)
	) name19306 (
		_w23343_,
		_w23352_,
		_w23353_
	);
	LUT2 #(
		.INIT('h2)
	) name19307 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[8]/NET0131 ,
		_w23343_,
		_w23354_
	);
	LUT2 #(
		.INIT('h1)
	) name19308 (
		_w23353_,
		_w23354_,
		_w23355_
	);
	LUT2 #(
		.INIT('h4)
	) name19309 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		_w23356_
	);
	LUT2 #(
		.INIT('h8)
	) name19310 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		_w23357_
	);
	LUT2 #(
		.INIT('h1)
	) name19311 (
		_w23356_,
		_w23357_,
		_w23358_
	);
	LUT2 #(
		.INIT('h2)
	) name19312 (
		_w23343_,
		_w23358_,
		_w23359_
	);
	LUT2 #(
		.INIT('h2)
	) name19313 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[7]/NET0131 ,
		_w23343_,
		_w23360_
	);
	LUT2 #(
		.INIT('h1)
	) name19314 (
		_w23359_,
		_w23360_,
		_w23361_
	);
	LUT2 #(
		.INIT('h4)
	) name19315 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		_w23362_
	);
	LUT2 #(
		.INIT('h8)
	) name19316 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		_w23363_
	);
	LUT2 #(
		.INIT('h1)
	) name19317 (
		_w23362_,
		_w23363_,
		_w23364_
	);
	LUT2 #(
		.INIT('h2)
	) name19318 (
		_w23343_,
		_w23364_,
		_w23365_
	);
	LUT2 #(
		.INIT('h2)
	) name19319 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[6]/NET0131 ,
		_w23343_,
		_w23366_
	);
	LUT2 #(
		.INIT('h1)
	) name19320 (
		_w23365_,
		_w23366_,
		_w23367_
	);
	LUT2 #(
		.INIT('h4)
	) name19321 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		_w23368_
	);
	LUT2 #(
		.INIT('h8)
	) name19322 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		_w23369_
	);
	LUT2 #(
		.INIT('h1)
	) name19323 (
		_w23368_,
		_w23369_,
		_w23370_
	);
	LUT2 #(
		.INIT('h2)
	) name19324 (
		_w23343_,
		_w23370_,
		_w23371_
	);
	LUT2 #(
		.INIT('h2)
	) name19325 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[5]/NET0131 ,
		_w23343_,
		_w23372_
	);
	LUT2 #(
		.INIT('h1)
	) name19326 (
		_w23371_,
		_w23372_,
		_w23373_
	);
	LUT2 #(
		.INIT('h4)
	) name19327 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		_w23374_
	);
	LUT2 #(
		.INIT('h8)
	) name19328 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		_w23375_
	);
	LUT2 #(
		.INIT('h1)
	) name19329 (
		_w23374_,
		_w23375_,
		_w23376_
	);
	LUT2 #(
		.INIT('h2)
	) name19330 (
		_w23343_,
		_w23376_,
		_w23377_
	);
	LUT2 #(
		.INIT('h2)
	) name19331 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[13]/NET0131 ,
		_w23343_,
		_w23378_
	);
	LUT2 #(
		.INIT('h1)
	) name19332 (
		_w23377_,
		_w23378_,
		_w23379_
	);
	LUT2 #(
		.INIT('h4)
	) name19333 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		_w23380_
	);
	LUT2 #(
		.INIT('h8)
	) name19334 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		_w23381_
	);
	LUT2 #(
		.INIT('h1)
	) name19335 (
		_w23380_,
		_w23381_,
		_w23382_
	);
	LUT2 #(
		.INIT('h2)
	) name19336 (
		_w23343_,
		_w23382_,
		_w23383_
	);
	LUT2 #(
		.INIT('h2)
	) name19337 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[12]/NET0131 ,
		_w23343_,
		_w23384_
	);
	LUT2 #(
		.INIT('h1)
	) name19338 (
		_w23383_,
		_w23384_,
		_w23385_
	);
	LUT2 #(
		.INIT('h4)
	) name19339 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w23386_
	);
	LUT2 #(
		.INIT('h8)
	) name19340 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		_w23387_
	);
	LUT2 #(
		.INIT('h1)
	) name19341 (
		_w23386_,
		_w23387_,
		_w23388_
	);
	LUT2 #(
		.INIT('h2)
	) name19342 (
		_w23343_,
		_w23388_,
		_w23389_
	);
	LUT2 #(
		.INIT('h2)
	) name19343 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[11]/NET0131 ,
		_w23343_,
		_w23390_
	);
	LUT2 #(
		.INIT('h1)
	) name19344 (
		_w23389_,
		_w23390_,
		_w23391_
	);
	LUT2 #(
		.INIT('h4)
	) name19345 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w23392_
	);
	LUT2 #(
		.INIT('h8)
	) name19346 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w23393_
	);
	LUT2 #(
		.INIT('h1)
	) name19347 (
		_w23392_,
		_w23393_,
		_w23394_
	);
	LUT2 #(
		.INIT('h2)
	) name19348 (
		_w23343_,
		_w23394_,
		_w23395_
	);
	LUT2 #(
		.INIT('h2)
	) name19349 (
		\core_dag_ilm1reg_STAC_pi_DO_reg[10]/NET0131 ,
		_w23343_,
		_w23396_
	);
	LUT2 #(
		.INIT('h1)
	) name19350 (
		_w23395_,
		_w23396_,
		_w23397_
	);
	LUT2 #(
		.INIT('h2)
	) name19351 (
		_w5429_,
		_w14733_,
		_w23398_
	);
	LUT2 #(
		.INIT('h2)
	) name19352 (
		\emc_IOcst_reg/NET0131 ,
		_w23398_,
		_w23399_
	);
	LUT2 #(
		.INIT('h4)
	) name19353 (
		_w19049_,
		_w23399_,
		_w23400_
	);
	LUT2 #(
		.INIT('h2)
	) name19354 (
		\memc_IOcmd_E_reg/NET0131 ,
		_w4068_,
		_w23401_
	);
	LUT2 #(
		.INIT('h8)
	) name19355 (
		_w19049_,
		_w23401_,
		_w23402_
	);
	LUT2 #(
		.INIT('h1)
	) name19356 (
		_w23400_,
		_w23402_,
		_w23403_
	);
	LUT2 #(
		.INIT('h2)
	) name19357 (
		\core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001 ,
		_w20864_,
		_w23404_
	);
	LUT2 #(
		.INIT('h4)
	) name19358 (
		_w19379_,
		_w20864_,
		_w23405_
	);
	LUT2 #(
		.INIT('h1)
	) name19359 (
		_w23404_,
		_w23405_,
		_w23406_
	);
	LUT2 #(
		.INIT('h8)
	) name19360 (
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		_w23407_
	);
	LUT2 #(
		.INIT('h1)
	) name19361 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w23408_
	);
	LUT2 #(
		.INIT('h8)
	) name19362 (
		_w23407_,
		_w23408_,
		_w23409_
	);
	LUT2 #(
		.INIT('h8)
	) name19363 (
		_w23032_,
		_w23409_,
		_w23410_
	);
	LUT2 #(
		.INIT('h2)
	) name19364 (
		\sice_ICYC_en_reg/NET0131 ,
		_w23410_,
		_w23411_
	);
	LUT2 #(
		.INIT('h8)
	) name19365 (
		\sice_SPC_reg[23]/P0001 ,
		_w23410_,
		_w23412_
	);
	LUT2 #(
		.INIT('h1)
	) name19366 (
		_w23411_,
		_w23412_,
		_w23413_
	);
	LUT2 #(
		.INIT('h2)
	) name19367 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001 ,
		_w20990_,
		_w23414_
	);
	LUT2 #(
		.INIT('h4)
	) name19368 (
		_w19379_,
		_w20990_,
		_w23415_
	);
	LUT2 #(
		.INIT('h1)
	) name19369 (
		_w23414_,
		_w23415_,
		_w23416_
	);
	LUT2 #(
		.INIT('h8)
	) name19370 (
		_w20845_,
		_w20847_,
		_w23417_
	);
	LUT2 #(
		.INIT('h8)
	) name19371 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		_w23417_,
		_w23418_
	);
	LUT2 #(
		.INIT('h8)
	) name19372 (
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		_w23418_,
		_w23419_
	);
	LUT2 #(
		.INIT('h8)
	) name19373 (
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		_w23419_,
		_w23420_
	);
	LUT2 #(
		.INIT('h8)
	) name19374 (
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		_w23420_,
		_w23421_
	);
	LUT2 #(
		.INIT('h8)
	) name19375 (
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		_w23421_,
		_w23422_
	);
	LUT2 #(
		.INIT('h1)
	) name19376 (
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w23422_,
		_w23423_
	);
	LUT2 #(
		.INIT('h8)
	) name19377 (
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w23422_,
		_w23424_
	);
	LUT2 #(
		.INIT('h1)
	) name19378 (
		_w23423_,
		_w23424_,
		_w23425_
	);
	LUT2 #(
		.INIT('h2)
	) name19379 (
		\core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001 ,
		_w20864_,
		_w23426_
	);
	LUT2 #(
		.INIT('h2)
	) name19380 (
		_w20864_,
		_w23220_,
		_w23427_
	);
	LUT2 #(
		.INIT('h1)
	) name19381 (
		_w23426_,
		_w23427_,
		_w23428_
	);
	LUT2 #(
		.INIT('h2)
	) name19382 (
		\sport1_rxctl_a_sync1_reg/P0001 ,
		\sport1_rxctl_a_sync2_reg/P0001 ,
		_w23429_
	);
	LUT2 #(
		.INIT('h8)
	) name19383 (
		\core_c_dec_MTRX1_E_reg/P0001 ,
		_w5951_,
		_w23430_
	);
	LUT2 #(
		.INIT('h2)
	) name19384 (
		\sport1_rxctl_RX_reg[9]/P0001 ,
		_w23430_,
		_w23431_
	);
	LUT2 #(
		.INIT('h8)
	) name19385 (
		_w10289_,
		_w23430_,
		_w23432_
	);
	LUT2 #(
		.INIT('h1)
	) name19386 (
		_w23431_,
		_w23432_,
		_w23433_
	);
	LUT2 #(
		.INIT('h1)
	) name19387 (
		_w23429_,
		_w23433_,
		_w23434_
	);
	LUT2 #(
		.INIT('h8)
	) name19388 (
		\sport1_rxctl_RXSHT_reg[9]/P0001 ,
		_w23429_,
		_w23435_
	);
	LUT2 #(
		.INIT('h1)
	) name19389 (
		_w23434_,
		_w23435_,
		_w23436_
	);
	LUT2 #(
		.INIT('h2)
	) name19390 (
		\sport1_rxctl_RX_reg[8]/P0001 ,
		_w23430_,
		_w23437_
	);
	LUT2 #(
		.INIT('h8)
	) name19391 (
		_w10638_,
		_w23430_,
		_w23438_
	);
	LUT2 #(
		.INIT('h1)
	) name19392 (
		_w23437_,
		_w23438_,
		_w23439_
	);
	LUT2 #(
		.INIT('h1)
	) name19393 (
		_w23429_,
		_w23439_,
		_w23440_
	);
	LUT2 #(
		.INIT('h8)
	) name19394 (
		\sport1_rxctl_RXSHT_reg[8]/P0001 ,
		_w23429_,
		_w23441_
	);
	LUT2 #(
		.INIT('h1)
	) name19395 (
		_w23440_,
		_w23441_,
		_w23442_
	);
	LUT2 #(
		.INIT('h2)
	) name19396 (
		\sport1_rxctl_RX_reg[7]/P0001 ,
		_w23430_,
		_w23443_
	);
	LUT2 #(
		.INIT('h8)
	) name19397 (
		_w11265_,
		_w23430_,
		_w23444_
	);
	LUT2 #(
		.INIT('h1)
	) name19398 (
		_w23443_,
		_w23444_,
		_w23445_
	);
	LUT2 #(
		.INIT('h1)
	) name19399 (
		_w23429_,
		_w23445_,
		_w23446_
	);
	LUT2 #(
		.INIT('h8)
	) name19400 (
		\sport1_rxctl_RXSHT_reg[7]/P0001 ,
		_w23429_,
		_w23447_
	);
	LUT2 #(
		.INIT('h1)
	) name19401 (
		_w23446_,
		_w23447_,
		_w23448_
	);
	LUT2 #(
		.INIT('h2)
	) name19402 (
		\sport1_rxctl_RX_reg[4]/P0001 ,
		_w23430_,
		_w23449_
	);
	LUT2 #(
		.INIT('h8)
	) name19403 (
		_w10069_,
		_w23430_,
		_w23450_
	);
	LUT2 #(
		.INIT('h1)
	) name19404 (
		_w23449_,
		_w23450_,
		_w23451_
	);
	LUT2 #(
		.INIT('h1)
	) name19405 (
		_w23429_,
		_w23451_,
		_w23452_
	);
	LUT2 #(
		.INIT('h8)
	) name19406 (
		\sport1_rxctl_RXSHT_reg[4]/P0001 ,
		_w23429_,
		_w23453_
	);
	LUT2 #(
		.INIT('h1)
	) name19407 (
		_w23452_,
		_w23453_,
		_w23454_
	);
	LUT2 #(
		.INIT('h2)
	) name19408 (
		\sport1_rxctl_RX_reg[6]/P0001 ,
		_w23430_,
		_w23455_
	);
	LUT2 #(
		.INIT('h8)
	) name19409 (
		_w11525_,
		_w23430_,
		_w23456_
	);
	LUT2 #(
		.INIT('h1)
	) name19410 (
		_w23455_,
		_w23456_,
		_w23457_
	);
	LUT2 #(
		.INIT('h1)
	) name19411 (
		_w23429_,
		_w23457_,
		_w23458_
	);
	LUT2 #(
		.INIT('h8)
	) name19412 (
		\sport1_rxctl_RXSHT_reg[6]/P0001 ,
		_w23429_,
		_w23459_
	);
	LUT2 #(
		.INIT('h1)
	) name19413 (
		_w23458_,
		_w23459_,
		_w23460_
	);
	LUT2 #(
		.INIT('h2)
	) name19414 (
		\sport1_rxctl_RX_reg[3]/P0001 ,
		_w23430_,
		_w23461_
	);
	LUT2 #(
		.INIT('h8)
	) name19415 (
		_w8113_,
		_w23430_,
		_w23462_
	);
	LUT2 #(
		.INIT('h1)
	) name19416 (
		_w23461_,
		_w23462_,
		_w23463_
	);
	LUT2 #(
		.INIT('h1)
	) name19417 (
		_w23429_,
		_w23463_,
		_w23464_
	);
	LUT2 #(
		.INIT('h8)
	) name19418 (
		\sport1_rxctl_RXSHT_reg[3]/P0001 ,
		_w23429_,
		_w23465_
	);
	LUT2 #(
		.INIT('h1)
	) name19419 (
		_w23464_,
		_w23465_,
		_w23466_
	);
	LUT2 #(
		.INIT('h2)
	) name19420 (
		\sport1_rxctl_RX_reg[5]/P0001 ,
		_w23430_,
		_w23467_
	);
	LUT2 #(
		.INIT('h8)
	) name19421 (
		_w10911_,
		_w23430_,
		_w23468_
	);
	LUT2 #(
		.INIT('h1)
	) name19422 (
		_w23467_,
		_w23468_,
		_w23469_
	);
	LUT2 #(
		.INIT('h1)
	) name19423 (
		_w23429_,
		_w23469_,
		_w23470_
	);
	LUT2 #(
		.INIT('h8)
	) name19424 (
		\sport1_rxctl_RXSHT_reg[5]/P0001 ,
		_w23429_,
		_w23471_
	);
	LUT2 #(
		.INIT('h1)
	) name19425 (
		_w23470_,
		_w23471_,
		_w23472_
	);
	LUT2 #(
		.INIT('h2)
	) name19426 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001 ,
		_w20990_,
		_w23473_
	);
	LUT2 #(
		.INIT('h2)
	) name19427 (
		_w20990_,
		_w23220_,
		_w23474_
	);
	LUT2 #(
		.INIT('h1)
	) name19428 (
		_w23473_,
		_w23474_,
		_w23475_
	);
	LUT2 #(
		.INIT('h2)
	) name19429 (
		\sport1_rxctl_RX_reg[2]/P0001 ,
		_w23430_,
		_w23476_
	);
	LUT2 #(
		.INIT('h8)
	) name19430 (
		_w8715_,
		_w23430_,
		_w23477_
	);
	LUT2 #(
		.INIT('h1)
	) name19431 (
		_w23476_,
		_w23477_,
		_w23478_
	);
	LUT2 #(
		.INIT('h1)
	) name19432 (
		_w23429_,
		_w23478_,
		_w23479_
	);
	LUT2 #(
		.INIT('h8)
	) name19433 (
		\sport1_rxctl_RXSHT_reg[2]/P0001 ,
		_w23429_,
		_w23480_
	);
	LUT2 #(
		.INIT('h1)
	) name19434 (
		_w23479_,
		_w23480_,
		_w23481_
	);
	LUT2 #(
		.INIT('h2)
	) name19435 (
		\sport1_rxctl_RX_reg[1]/P0001 ,
		_w23430_,
		_w23482_
	);
	LUT2 #(
		.INIT('h8)
	) name19436 (
		_w9435_,
		_w23430_,
		_w23483_
	);
	LUT2 #(
		.INIT('h1)
	) name19437 (
		_w23482_,
		_w23483_,
		_w23484_
	);
	LUT2 #(
		.INIT('h1)
	) name19438 (
		_w23429_,
		_w23484_,
		_w23485_
	);
	LUT2 #(
		.INIT('h8)
	) name19439 (
		\sport1_rxctl_RXSHT_reg[1]/P0001 ,
		_w23429_,
		_w23486_
	);
	LUT2 #(
		.INIT('h1)
	) name19440 (
		_w23485_,
		_w23486_,
		_w23487_
	);
	LUT2 #(
		.INIT('h2)
	) name19441 (
		\sport1_rxctl_RX_reg[15]/P0001 ,
		_w23430_,
		_w23488_
	);
	LUT2 #(
		.INIT('h8)
	) name19442 (
		_w12743_,
		_w23430_,
		_w23489_
	);
	LUT2 #(
		.INIT('h1)
	) name19443 (
		_w23488_,
		_w23489_,
		_w23490_
	);
	LUT2 #(
		.INIT('h1)
	) name19444 (
		_w23429_,
		_w23490_,
		_w23491_
	);
	LUT2 #(
		.INIT('h8)
	) name19445 (
		\sport1_rxctl_RXSHT_reg[15]/P0001 ,
		_w23429_,
		_w23492_
	);
	LUT2 #(
		.INIT('h1)
	) name19446 (
		_w23491_,
		_w23492_,
		_w23493_
	);
	LUT2 #(
		.INIT('h2)
	) name19447 (
		\sport1_rxctl_RX_reg[14]/P0001 ,
		_w23430_,
		_w23494_
	);
	LUT2 #(
		.INIT('h8)
	) name19448 (
		_w12688_,
		_w23430_,
		_w23495_
	);
	LUT2 #(
		.INIT('h1)
	) name19449 (
		_w23494_,
		_w23495_,
		_w23496_
	);
	LUT2 #(
		.INIT('h1)
	) name19450 (
		_w23429_,
		_w23496_,
		_w23497_
	);
	LUT2 #(
		.INIT('h8)
	) name19451 (
		\sport1_rxctl_RXSHT_reg[14]/P0001 ,
		_w23429_,
		_w23498_
	);
	LUT2 #(
		.INIT('h1)
	) name19452 (
		_w23497_,
		_w23498_,
		_w23499_
	);
	LUT2 #(
		.INIT('h2)
	) name19453 (
		\sport1_rxctl_RX_reg[13]/P0001 ,
		_w23430_,
		_w23500_
	);
	LUT2 #(
		.INIT('h8)
	) name19454 (
		_w7340_,
		_w23430_,
		_w23501_
	);
	LUT2 #(
		.INIT('h1)
	) name19455 (
		_w23500_,
		_w23501_,
		_w23502_
	);
	LUT2 #(
		.INIT('h1)
	) name19456 (
		_w23429_,
		_w23502_,
		_w23503_
	);
	LUT2 #(
		.INIT('h8)
	) name19457 (
		\sport1_rxctl_RXSHT_reg[13]/P0001 ,
		_w23429_,
		_w23504_
	);
	LUT2 #(
		.INIT('h1)
	) name19458 (
		_w23503_,
		_w23504_,
		_w23505_
	);
	LUT2 #(
		.INIT('h2)
	) name19459 (
		\sport1_rxctl_RX_reg[12]/P0001 ,
		_w23430_,
		_w23506_
	);
	LUT2 #(
		.INIT('h8)
	) name19460 (
		_w9178_,
		_w23430_,
		_w23507_
	);
	LUT2 #(
		.INIT('h1)
	) name19461 (
		_w23506_,
		_w23507_,
		_w23508_
	);
	LUT2 #(
		.INIT('h1)
	) name19462 (
		_w23429_,
		_w23508_,
		_w23509_
	);
	LUT2 #(
		.INIT('h8)
	) name19463 (
		\sport1_rxctl_RXSHT_reg[12]/P0001 ,
		_w23429_,
		_w23510_
	);
	LUT2 #(
		.INIT('h1)
	) name19464 (
		_w23509_,
		_w23510_,
		_w23511_
	);
	LUT2 #(
		.INIT('h2)
	) name19465 (
		\sport1_rxctl_RX_reg[11]/P0001 ,
		_w23430_,
		_w23512_
	);
	LUT2 #(
		.INIT('h8)
	) name19466 (
		_w8460_,
		_w23430_,
		_w23513_
	);
	LUT2 #(
		.INIT('h1)
	) name19467 (
		_w23512_,
		_w23513_,
		_w23514_
	);
	LUT2 #(
		.INIT('h1)
	) name19468 (
		_w23429_,
		_w23514_,
		_w23515_
	);
	LUT2 #(
		.INIT('h8)
	) name19469 (
		\sport1_rxctl_RXSHT_reg[11]/P0001 ,
		_w23429_,
		_w23516_
	);
	LUT2 #(
		.INIT('h1)
	) name19470 (
		_w23515_,
		_w23516_,
		_w23517_
	);
	LUT2 #(
		.INIT('h2)
	) name19471 (
		\sport1_rxctl_RX_reg[10]/P0001 ,
		_w23430_,
		_w23518_
	);
	LUT2 #(
		.INIT('h8)
	) name19472 (
		_w7859_,
		_w23430_,
		_w23519_
	);
	LUT2 #(
		.INIT('h1)
	) name19473 (
		_w23518_,
		_w23519_,
		_w23520_
	);
	LUT2 #(
		.INIT('h1)
	) name19474 (
		_w23429_,
		_w23520_,
		_w23521_
	);
	LUT2 #(
		.INIT('h8)
	) name19475 (
		\sport1_rxctl_RXSHT_reg[10]/P0001 ,
		_w23429_,
		_w23522_
	);
	LUT2 #(
		.INIT('h1)
	) name19476 (
		_w23521_,
		_w23522_,
		_w23523_
	);
	LUT2 #(
		.INIT('h2)
	) name19477 (
		\sport1_rxctl_RX_reg[0]/P0001 ,
		_w23430_,
		_w23524_
	);
	LUT2 #(
		.INIT('h8)
	) name19478 (
		_w7607_,
		_w23430_,
		_w23525_
	);
	LUT2 #(
		.INIT('h1)
	) name19479 (
		_w23524_,
		_w23525_,
		_w23526_
	);
	LUT2 #(
		.INIT('h1)
	) name19480 (
		_w23429_,
		_w23526_,
		_w23527_
	);
	LUT2 #(
		.INIT('h8)
	) name19481 (
		\sport1_rxctl_RXSHT_reg[0]/P0001 ,
		_w23429_,
		_w23528_
	);
	LUT2 #(
		.INIT('h1)
	) name19482 (
		_w23527_,
		_w23528_,
		_w23529_
	);
	LUT2 #(
		.INIT('h2)
	) name19483 (
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		_w4116_,
		_w23530_
	);
	LUT2 #(
		.INIT('h2)
	) name19484 (
		\core_c_psq_T_PWRDN_reg/P0001 ,
		\core_c_psq_T_PWRDN_s1_reg/P0001 ,
		_w23531_
	);
	LUT2 #(
		.INIT('h1)
	) name19485 (
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		\sport0_regs_AUTO_a_reg[13]/NET0131 ,
		_w23532_
	);
	LUT2 #(
		.INIT('h4)
	) name19486 (
		_w23531_,
		_w23532_,
		_w23533_
	);
	LUT2 #(
		.INIT('h1)
	) name19487 (
		_w23530_,
		_w23533_,
		_w23534_
	);
	LUT2 #(
		.INIT('h1)
	) name19488 (
		\sice_ICYC_reg[9]/NET0131 ,
		_w20738_,
		_w23535_
	);
	LUT2 #(
		.INIT('h1)
	) name19489 (
		_w20739_,
		_w23535_,
		_w23536_
	);
	LUT2 #(
		.INIT('h1)
	) name19490 (
		\sice_IIRC_reg[6]/NET0131 ,
		_w18869_,
		_w23537_
	);
	LUT2 #(
		.INIT('h1)
	) name19491 (
		_w18870_,
		_w23537_,
		_w23538_
	);
	LUT2 #(
		.INIT('h1)
	) name19492 (
		\sice_IIRC_reg[9]/NET0131 ,
		_w20853_,
		_w23539_
	);
	LUT2 #(
		.INIT('h1)
	) name19493 (
		_w20854_,
		_w23539_,
		_w23540_
	);
	LUT2 #(
		.INIT('h1)
	) name19494 (
		\sice_ICYC_reg[6]/NET0131 ,
		_w18860_,
		_w23541_
	);
	LUT2 #(
		.INIT('h1)
	) name19495 (
		_w18861_,
		_w23541_,
		_w23542_
	);
	LUT2 #(
		.INIT('h2)
	) name19496 (
		\emc_DMDreg_reg[7]/P0001 ,
		_w14737_,
		_w23543_
	);
	LUT2 #(
		.INIT('h8)
	) name19497 (
		\T_ED[7]_pad ,
		_w14737_,
		_w23544_
	);
	LUT2 #(
		.INIT('h1)
	) name19498 (
		_w23543_,
		_w23544_,
		_w23545_
	);
	LUT2 #(
		.INIT('h2)
	) name19499 (
		\emc_DMDreg_reg[6]/P0001 ,
		_w14737_,
		_w23546_
	);
	LUT2 #(
		.INIT('h8)
	) name19500 (
		\T_ED[6]_pad ,
		_w14737_,
		_w23547_
	);
	LUT2 #(
		.INIT('h1)
	) name19501 (
		_w23546_,
		_w23547_,
		_w23548_
	);
	LUT2 #(
		.INIT('h2)
	) name19502 (
		\emc_DMDreg_reg[5]/P0001 ,
		_w14737_,
		_w23549_
	);
	LUT2 #(
		.INIT('h8)
	) name19503 (
		\T_ED[5]_pad ,
		_w14737_,
		_w23550_
	);
	LUT2 #(
		.INIT('h1)
	) name19504 (
		_w23549_,
		_w23550_,
		_w23551_
	);
	LUT2 #(
		.INIT('h2)
	) name19505 (
		\emc_DMDreg_reg[4]/P0001 ,
		_w14737_,
		_w23552_
	);
	LUT2 #(
		.INIT('h8)
	) name19506 (
		\T_ED[4]_pad ,
		_w14737_,
		_w23553_
	);
	LUT2 #(
		.INIT('h1)
	) name19507 (
		_w23552_,
		_w23553_,
		_w23554_
	);
	LUT2 #(
		.INIT('h2)
	) name19508 (
		\emc_DMDreg_reg[3]/P0001 ,
		_w14737_,
		_w23555_
	);
	LUT2 #(
		.INIT('h8)
	) name19509 (
		\T_ED[3]_pad ,
		_w14737_,
		_w23556_
	);
	LUT2 #(
		.INIT('h1)
	) name19510 (
		_w23555_,
		_w23556_,
		_w23557_
	);
	LUT2 #(
		.INIT('h2)
	) name19511 (
		\emc_DMDreg_reg[2]/P0001 ,
		_w14737_,
		_w23558_
	);
	LUT2 #(
		.INIT('h8)
	) name19512 (
		\T_ED[2]_pad ,
		_w14737_,
		_w23559_
	);
	LUT2 #(
		.INIT('h1)
	) name19513 (
		_w23558_,
		_w23559_,
		_w23560_
	);
	LUT2 #(
		.INIT('h2)
	) name19514 (
		\emc_DMDreg_reg[1]/P0001 ,
		_w14737_,
		_w23561_
	);
	LUT2 #(
		.INIT('h8)
	) name19515 (
		\T_ED[1]_pad ,
		_w14737_,
		_w23562_
	);
	LUT2 #(
		.INIT('h1)
	) name19516 (
		_w23561_,
		_w23562_,
		_w23563_
	);
	LUT2 #(
		.INIT('h2)
	) name19517 (
		\emc_DMDreg_reg[15]/P0001 ,
		_w14737_,
		_w23564_
	);
	LUT2 #(
		.INIT('h8)
	) name19518 (
		\T_ED[15]_pad ,
		_w14737_,
		_w23565_
	);
	LUT2 #(
		.INIT('h1)
	) name19519 (
		_w23564_,
		_w23565_,
		_w23566_
	);
	LUT2 #(
		.INIT('h2)
	) name19520 (
		\emc_DMDreg_reg[14]/P0001 ,
		_w14737_,
		_w23567_
	);
	LUT2 #(
		.INIT('h8)
	) name19521 (
		\T_ED[14]_pad ,
		_w14737_,
		_w23568_
	);
	LUT2 #(
		.INIT('h1)
	) name19522 (
		_w23567_,
		_w23568_,
		_w23569_
	);
	LUT2 #(
		.INIT('h2)
	) name19523 (
		\emc_DMDreg_reg[13]/P0001 ,
		_w14737_,
		_w23570_
	);
	LUT2 #(
		.INIT('h8)
	) name19524 (
		\T_ED[13]_pad ,
		_w14737_,
		_w23571_
	);
	LUT2 #(
		.INIT('h1)
	) name19525 (
		_w23570_,
		_w23571_,
		_w23572_
	);
	LUT2 #(
		.INIT('h2)
	) name19526 (
		\emc_DMDreg_reg[12]/P0001 ,
		_w14737_,
		_w23573_
	);
	LUT2 #(
		.INIT('h8)
	) name19527 (
		\T_ED[12]_pad ,
		_w14737_,
		_w23574_
	);
	LUT2 #(
		.INIT('h1)
	) name19528 (
		_w23573_,
		_w23574_,
		_w23575_
	);
	LUT2 #(
		.INIT('h2)
	) name19529 (
		\emc_DMDreg_reg[11]/P0001 ,
		_w14737_,
		_w23576_
	);
	LUT2 #(
		.INIT('h8)
	) name19530 (
		\T_ED[11]_pad ,
		_w14737_,
		_w23577_
	);
	LUT2 #(
		.INIT('h1)
	) name19531 (
		_w23576_,
		_w23577_,
		_w23578_
	);
	LUT2 #(
		.INIT('h2)
	) name19532 (
		\emc_DMDreg_reg[10]/P0001 ,
		_w14737_,
		_w23579_
	);
	LUT2 #(
		.INIT('h8)
	) name19533 (
		\T_ED[10]_pad ,
		_w14737_,
		_w23580_
	);
	LUT2 #(
		.INIT('h1)
	) name19534 (
		_w23579_,
		_w23580_,
		_w23581_
	);
	LUT2 #(
		.INIT('h2)
	) name19535 (
		\emc_DMDreg_reg[0]/P0001 ,
		_w14737_,
		_w23582_
	);
	LUT2 #(
		.INIT('h8)
	) name19536 (
		\T_ED[0]_pad ,
		_w14737_,
		_w23583_
	);
	LUT2 #(
		.INIT('h1)
	) name19537 (
		_w23582_,
		_w23583_,
		_w23584_
	);
	LUT2 #(
		.INIT('h8)
	) name19538 (
		\core_c_dec_SHTop_E_reg/P0001 ,
		_w17838_,
		_w23585_
	);
	LUT2 #(
		.INIT('h4)
	) name19539 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w23585_,
		_w23586_
	);
	LUT2 #(
		.INIT('h8)
	) name19540 (
		_w14033_,
		_w23585_,
		_w23587_
	);
	LUT2 #(
		.INIT('h1)
	) name19541 (
		_w7172_,
		_w7373_,
		_w23588_
	);
	LUT2 #(
		.INIT('h8)
	) name19542 (
		_w7995_,
		_w8501_,
		_w23589_
	);
	LUT2 #(
		.INIT('h2)
	) name19543 (
		_w9272_,
		_w9939_,
		_w23590_
	);
	LUT2 #(
		.INIT('h1)
	) name19544 (
		_w10789_,
		_w11303_,
		_w23591_
	);
	LUT2 #(
		.INIT('h8)
	) name19545 (
		_w23590_,
		_w23591_,
		_w23592_
	);
	LUT2 #(
		.INIT('h8)
	) name19546 (
		_w23588_,
		_w23589_,
		_w23593_
	);
	LUT2 #(
		.INIT('h8)
	) name19547 (
		_w23587_,
		_w23593_,
		_w23594_
	);
	LUT2 #(
		.INIT('h8)
	) name19548 (
		_w23592_,
		_w23594_,
		_w23595_
	);
	LUT2 #(
		.INIT('h1)
	) name19549 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w23586_,
		_w23596_
	);
	LUT2 #(
		.INIT('h4)
	) name19550 (
		_w23595_,
		_w23596_,
		_w23597_
	);
	LUT2 #(
		.INIT('h2)
	) name19551 (
		_w13804_,
		_w23597_,
		_w23598_
	);
	LUT2 #(
		.INIT('h2)
	) name19552 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w19559_,
		_w23599_
	);
	LUT2 #(
		.INIT('h8)
	) name19553 (
		_w17938_,
		_w23585_,
		_w23600_
	);
	LUT2 #(
		.INIT('h4)
	) name19554 (
		_w18123_,
		_w23600_,
		_w23601_
	);
	LUT2 #(
		.INIT('h4)
	) name19555 (
		_w17938_,
		_w23585_,
		_w23602_
	);
	LUT2 #(
		.INIT('h8)
	) name19556 (
		_w18123_,
		_w23602_,
		_w23603_
	);
	LUT2 #(
		.INIT('h1)
	) name19557 (
		_w23601_,
		_w23603_,
		_w23604_
	);
	LUT2 #(
		.INIT('h4)
	) name19558 (
		_w18127_,
		_w23600_,
		_w23605_
	);
	LUT2 #(
		.INIT('h8)
	) name19559 (
		_w18127_,
		_w23602_,
		_w23606_
	);
	LUT2 #(
		.INIT('h1)
	) name19560 (
		_w23605_,
		_w23606_,
		_w23607_
	);
	LUT2 #(
		.INIT('h4)
	) name19561 (
		_w17938_,
		_w18098_,
		_w23608_
	);
	LUT2 #(
		.INIT('h1)
	) name19562 (
		_w18098_,
		_w23602_,
		_w23609_
	);
	LUT2 #(
		.INIT('h1)
	) name19563 (
		_w23608_,
		_w23609_,
		_w23610_
	);
	LUT2 #(
		.INIT('h2)
	) name19564 (
		_w17938_,
		_w18102_,
		_w23611_
	);
	LUT2 #(
		.INIT('h4)
	) name19565 (
		_w17938_,
		_w18102_,
		_w23612_
	);
	LUT2 #(
		.INIT('h1)
	) name19566 (
		_w23611_,
		_w23612_,
		_w23613_
	);
	LUT2 #(
		.INIT('h8)
	) name19567 (
		_w23585_,
		_w23610_,
		_w23614_
	);
	LUT2 #(
		.INIT('h4)
	) name19568 (
		_w23613_,
		_w23614_,
		_w23615_
	);
	LUT2 #(
		.INIT('h2)
	) name19569 (
		_w23607_,
		_w23615_,
		_w23616_
	);
	LUT2 #(
		.INIT('h2)
	) name19570 (
		_w23604_,
		_w23616_,
		_w23617_
	);
	LUT2 #(
		.INIT('h4)
	) name19571 (
		_w18165_,
		_w23600_,
		_w23618_
	);
	LUT2 #(
		.INIT('h8)
	) name19572 (
		_w18165_,
		_w23602_,
		_w23619_
	);
	LUT2 #(
		.INIT('h1)
	) name19573 (
		_w23618_,
		_w23619_,
		_w23620_
	);
	LUT2 #(
		.INIT('h4)
	) name19574 (
		_w23617_,
		_w23620_,
		_w23621_
	);
	LUT2 #(
		.INIT('h1)
	) name19575 (
		_w17938_,
		_w18161_,
		_w23622_
	);
	LUT2 #(
		.INIT('h8)
	) name19576 (
		_w17938_,
		_w18161_,
		_w23623_
	);
	LUT2 #(
		.INIT('h2)
	) name19577 (
		_w23585_,
		_w23622_,
		_w23624_
	);
	LUT2 #(
		.INIT('h4)
	) name19578 (
		_w23623_,
		_w23624_,
		_w23625_
	);
	LUT2 #(
		.INIT('h1)
	) name19579 (
		_w23621_,
		_w23625_,
		_w23626_
	);
	LUT2 #(
		.INIT('h1)
	) name19580 (
		_w17938_,
		_w18186_,
		_w23627_
	);
	LUT2 #(
		.INIT('h8)
	) name19581 (
		_w17938_,
		_w18186_,
		_w23628_
	);
	LUT2 #(
		.INIT('h2)
	) name19582 (
		_w23585_,
		_w23627_,
		_w23629_
	);
	LUT2 #(
		.INIT('h4)
	) name19583 (
		_w23628_,
		_w23629_,
		_w23630_
	);
	LUT2 #(
		.INIT('h1)
	) name19584 (
		_w23626_,
		_w23630_,
		_w23631_
	);
	LUT2 #(
		.INIT('h4)
	) name19585 (
		_w18182_,
		_w23600_,
		_w23632_
	);
	LUT2 #(
		.INIT('h8)
	) name19586 (
		_w18182_,
		_w23602_,
		_w23633_
	);
	LUT2 #(
		.INIT('h1)
	) name19587 (
		_w23632_,
		_w23633_,
		_w23634_
	);
	LUT2 #(
		.INIT('h4)
	) name19588 (
		_w23631_,
		_w23634_,
		_w23635_
	);
	LUT2 #(
		.INIT('h4)
	) name19589 (
		_w18135_,
		_w23600_,
		_w23636_
	);
	LUT2 #(
		.INIT('h8)
	) name19590 (
		_w18135_,
		_w23602_,
		_w23637_
	);
	LUT2 #(
		.INIT('h1)
	) name19591 (
		_w23636_,
		_w23637_,
		_w23638_
	);
	LUT2 #(
		.INIT('h4)
	) name19592 (
		_w23635_,
		_w23638_,
		_w23639_
	);
	LUT2 #(
		.INIT('h4)
	) name19593 (
		_w18170_,
		_w23600_,
		_w23640_
	);
	LUT2 #(
		.INIT('h8)
	) name19594 (
		_w18170_,
		_w23602_,
		_w23641_
	);
	LUT2 #(
		.INIT('h1)
	) name19595 (
		_w23640_,
		_w23641_,
		_w23642_
	);
	LUT2 #(
		.INIT('h4)
	) name19596 (
		_w23639_,
		_w23642_,
		_w23643_
	);
	LUT2 #(
		.INIT('h4)
	) name19597 (
		_w18114_,
		_w23600_,
		_w23644_
	);
	LUT2 #(
		.INIT('h8)
	) name19598 (
		_w18114_,
		_w23602_,
		_w23645_
	);
	LUT2 #(
		.INIT('h1)
	) name19599 (
		_w23644_,
		_w23645_,
		_w23646_
	);
	LUT2 #(
		.INIT('h4)
	) name19600 (
		_w23643_,
		_w23646_,
		_w23647_
	);
	LUT2 #(
		.INIT('h4)
	) name19601 (
		_w18110_,
		_w23600_,
		_w23648_
	);
	LUT2 #(
		.INIT('h8)
	) name19602 (
		_w18110_,
		_w23602_,
		_w23649_
	);
	LUT2 #(
		.INIT('h1)
	) name19603 (
		_w23648_,
		_w23649_,
		_w23650_
	);
	LUT2 #(
		.INIT('h4)
	) name19604 (
		_w23647_,
		_w23650_,
		_w23651_
	);
	LUT2 #(
		.INIT('h4)
	) name19605 (
		_w17933_,
		_w23600_,
		_w23652_
	);
	LUT2 #(
		.INIT('h8)
	) name19606 (
		_w17933_,
		_w23602_,
		_w23653_
	);
	LUT2 #(
		.INIT('h1)
	) name19607 (
		_w23652_,
		_w23653_,
		_w23654_
	);
	LUT2 #(
		.INIT('h4)
	) name19608 (
		_w23651_,
		_w23654_,
		_w23655_
	);
	LUT2 #(
		.INIT('h4)
	) name19609 (
		_w17924_,
		_w23600_,
		_w23656_
	);
	LUT2 #(
		.INIT('h8)
	) name19610 (
		_w17924_,
		_w23602_,
		_w23657_
	);
	LUT2 #(
		.INIT('h1)
	) name19611 (
		_w23656_,
		_w23657_,
		_w23658_
	);
	LUT2 #(
		.INIT('h4)
	) name19612 (
		_w23655_,
		_w23658_,
		_w23659_
	);
	LUT2 #(
		.INIT('h4)
	) name19613 (
		_w18175_,
		_w23600_,
		_w23660_
	);
	LUT2 #(
		.INIT('h8)
	) name19614 (
		_w18175_,
		_w23602_,
		_w23661_
	);
	LUT2 #(
		.INIT('h1)
	) name19615 (
		_w23660_,
		_w23661_,
		_w23662_
	);
	LUT2 #(
		.INIT('h4)
	) name19616 (
		_w23659_,
		_w23662_,
		_w23663_
	);
	LUT2 #(
		.INIT('h8)
	) name19617 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w13881_,
		_w23664_
	);
	LUT2 #(
		.INIT('h8)
	) name19618 (
		_w23585_,
		_w23664_,
		_w23665_
	);
	LUT2 #(
		.INIT('h4)
	) name19619 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w17938_,
		_w23666_
	);
	LUT2 #(
		.INIT('h8)
	) name19620 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w23602_,
		_w23667_
	);
	LUT2 #(
		.INIT('h2)
	) name19621 (
		_w23587_,
		_w23666_,
		_w23668_
	);
	LUT2 #(
		.INIT('h4)
	) name19622 (
		_w23667_,
		_w23668_,
		_w23669_
	);
	LUT2 #(
		.INIT('h1)
	) name19623 (
		_w23665_,
		_w23669_,
		_w23670_
	);
	LUT2 #(
		.INIT('h4)
	) name19624 (
		_w23663_,
		_w23670_,
		_w23671_
	);
	LUT2 #(
		.INIT('h4)
	) name19625 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w23671_,
		_w23672_
	);
	LUT2 #(
		.INIT('h1)
	) name19626 (
		_w23599_,
		_w23672_,
		_w23673_
	);
	LUT2 #(
		.INIT('h2)
	) name19627 (
		_w23598_,
		_w23673_,
		_w23674_
	);
	LUT2 #(
		.INIT('h1)
	) name19628 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[0]/P0001 ,
		_w23598_,
		_w23675_
	);
	LUT2 #(
		.INIT('h1)
	) name19629 (
		_w23674_,
		_w23675_,
		_w23676_
	);
	LUT2 #(
		.INIT('h2)
	) name19630 (
		_w14666_,
		_w23597_,
		_w23677_
	);
	LUT2 #(
		.INIT('h4)
	) name19631 (
		_w23673_,
		_w23677_,
		_w23678_
	);
	LUT2 #(
		.INIT('h1)
	) name19632 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[0]/P0001 ,
		_w23677_,
		_w23679_
	);
	LUT2 #(
		.INIT('h1)
	) name19633 (
		_w23678_,
		_w23679_,
		_w23680_
	);
	LUT2 #(
		.INIT('h4)
	) name19634 (
		_w13806_,
		_w23253_,
		_w23681_
	);
	LUT2 #(
		.INIT('h8)
	) name19635 (
		_w13806_,
		_w14623_,
		_w23682_
	);
	LUT2 #(
		.INIT('h1)
	) name19636 (
		_w23681_,
		_w23682_,
		_w23683_
	);
	LUT2 #(
		.INIT('h2)
	) name19637 (
		_w14667_,
		_w23683_,
		_w23684_
	);
	LUT2 #(
		.INIT('h1)
	) name19638 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[7]/P0001 ,
		_w14667_,
		_w23685_
	);
	LUT2 #(
		.INIT('h1)
	) name19639 (
		_w23684_,
		_w23685_,
		_w23686_
	);
	LUT2 #(
		.INIT('h2)
	) name19640 (
		_w13805_,
		_w23683_,
		_w23687_
	);
	LUT2 #(
		.INIT('h1)
	) name19641 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[7]/P0001 ,
		_w13805_,
		_w23688_
	);
	LUT2 #(
		.INIT('h1)
	) name19642 (
		_w23687_,
		_w23688_,
		_w23689_
	);
	LUT2 #(
		.INIT('h2)
	) name19643 (
		_w4149_,
		_w20355_,
		_w23690_
	);
	LUT2 #(
		.INIT('h2)
	) name19644 (
		_w12234_,
		_w23019_,
		_w23691_
	);
	LUT2 #(
		.INIT('h4)
	) name19645 (
		\core_c_dec_cdAM_E_reg/P0001 ,
		_w4117_,
		_w23692_
	);
	LUT2 #(
		.INIT('h2)
	) name19646 (
		_w4116_,
		_w14729_,
		_w23693_
	);
	LUT2 #(
		.INIT('h4)
	) name19647 (
		_w23692_,
		_w23693_,
		_w23694_
	);
	LUT2 #(
		.INIT('h8)
	) name19648 (
		\tm_tcr_reg_DO_reg[9]/NET0131 ,
		_w20355_,
		_w23695_
	);
	LUT2 #(
		.INIT('h4)
	) name19649 (
		\tm_tpr_reg_DO_reg[9]/NET0131 ,
		_w22400_,
		_w23696_
	);
	LUT2 #(
		.INIT('h2)
	) name19650 (
		_w22411_,
		_w22422_,
		_w23697_
	);
	LUT2 #(
		.INIT('h2)
	) name19651 (
		\tm_TCR_TMP_reg[9]/NET0131 ,
		_w23697_,
		_w23698_
	);
	LUT2 #(
		.INIT('h8)
	) name19652 (
		_w22411_,
		_w22423_,
		_w23699_
	);
	LUT2 #(
		.INIT('h1)
	) name19653 (
		_w22400_,
		_w23698_,
		_w23700_
	);
	LUT2 #(
		.INIT('h4)
	) name19654 (
		_w23699_,
		_w23700_,
		_w23701_
	);
	LUT2 #(
		.INIT('h1)
	) name19655 (
		_w20355_,
		_w23696_,
		_w23702_
	);
	LUT2 #(
		.INIT('h4)
	) name19656 (
		_w23701_,
		_w23702_,
		_w23703_
	);
	LUT2 #(
		.INIT('h1)
	) name19657 (
		_w23695_,
		_w23703_,
		_w23704_
	);
	LUT2 #(
		.INIT('h8)
	) name19658 (
		_w13776_,
		_w13778_,
		_w23705_
	);
	LUT2 #(
		.INIT('h1)
	) name19659 (
		\core_c_psq_SSTAT_reg[3]/NET0131 ,
		_w23705_,
		_w23706_
	);
	LUT2 #(
		.INIT('h8)
	) name19660 (
		\core_c_dec_DIVQ_E_reg/P0001 ,
		_w4117_,
		_w23707_
	);
	LUT2 #(
		.INIT('h1)
	) name19661 (
		_w21560_,
		_w23707_,
		_w23708_
	);
	LUT2 #(
		.INIT('h2)
	) name19662 (
		_w4116_,
		_w23708_,
		_w23709_
	);
	LUT2 #(
		.INIT('h8)
	) name19663 (
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w20036_,
		_w23710_
	);
	LUT2 #(
		.INIT('h1)
	) name19664 (
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w23710_,
		_w23711_
	);
	LUT2 #(
		.INIT('h1)
	) name19665 (
		_w20038_,
		_w23711_,
		_w23712_
	);
	LUT2 #(
		.INIT('h4)
	) name19666 (
		_w13750_,
		_w23712_,
		_w23713_
	);
	LUT2 #(
		.INIT('h1)
	) name19667 (
		\clkc_SlowDn_reg/NET0131 ,
		\clkc_SlowDn_s1_reg/P0001 ,
		_w23714_
	);
	LUT2 #(
		.INIT('h4)
	) name19668 (
		\clkc_SlowDn_s2_reg/P0001 ,
		_w23714_,
		_w23715_
	);
	LUT2 #(
		.INIT('h8)
	) name19669 (
		_w4071_,
		_w6929_,
		_w23716_
	);
	LUT2 #(
		.INIT('h8)
	) name19670 (
		_w4112_,
		_w23716_,
		_w23717_
	);
	LUT2 #(
		.INIT('h4)
	) name19671 (
		_w23018_,
		_w23715_,
		_w23718_
	);
	LUT2 #(
		.INIT('h8)
	) name19672 (
		_w23717_,
		_w23718_,
		_w23719_
	);
	LUT2 #(
		.INIT('h8)
	) name19673 (
		\core_c_dec_NOP_E_reg/P0001 ,
		_w4117_,
		_w23720_
	);
	LUT2 #(
		.INIT('h2)
	) name19674 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w23721_
	);
	LUT2 #(
		.INIT('h8)
	) name19675 (
		_w21249_,
		_w23721_,
		_w23722_
	);
	LUT2 #(
		.INIT('h8)
	) name19676 (
		_w5664_,
		_w23722_,
		_w23723_
	);
	LUT2 #(
		.INIT('h1)
	) name19677 (
		_w23720_,
		_w23723_,
		_w23724_
	);
	LUT2 #(
		.INIT('h2)
	) name19678 (
		_w4116_,
		_w23724_,
		_w23725_
	);
	LUT2 #(
		.INIT('h2)
	) name19679 (
		_w23264_,
		_w23272_,
		_w23726_
	);
	LUT2 #(
		.INIT('h1)
	) name19680 (
		_w23429_,
		_w23430_,
		_w23727_
	);
	LUT2 #(
		.INIT('h8)
	) name19681 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w23728_
	);
	LUT2 #(
		.INIT('h4)
	) name19682 (
		_w23727_,
		_w23728_,
		_w23729_
	);
	LUT2 #(
		.INIT('h1)
	) name19683 (
		\sport1_rxctl_RSreq_reg/NET0131 ,
		_w23729_,
		_w23730_
	);
	LUT2 #(
		.INIT('h8)
	) name19684 (
		\emc_eRDY_reg/NET0131 ,
		_w4118_,
		_w23731_
	);
	LUT2 #(
		.INIT('h4)
	) name19685 (
		\T_TMODE[1]_pad ,
		_w5581_,
		_w23732_
	);
	LUT2 #(
		.INIT('h8)
	) name19686 (
		_w5560_,
		_w23732_,
		_w23733_
	);
	LUT2 #(
		.INIT('h2)
	) name19687 (
		\T_TMODE[1]_pad ,
		_w5581_,
		_w23734_
	);
	LUT2 #(
		.INIT('h8)
	) name19688 (
		_w5605_,
		_w23734_,
		_w23735_
	);
	LUT2 #(
		.INIT('h1)
	) name19689 (
		_w23733_,
		_w23735_,
		_w23736_
	);
	LUT2 #(
		.INIT('h1)
	) name19690 (
		\emc_eRDY_reg/NET0131 ,
		_w5586_,
		_w23737_
	);
	LUT2 #(
		.INIT('h4)
	) name19691 (
		_w23736_,
		_w23737_,
		_w23738_
	);
	LUT2 #(
		.INIT('h1)
	) name19692 (
		_w23731_,
		_w23738_,
		_w23739_
	);
	LUT2 #(
		.INIT('h4)
	) name19693 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w20868_,
		_w23740_
	);
	LUT2 #(
		.INIT('h1)
	) name19694 (
		_w20875_,
		_w23740_,
		_w23741_
	);
	LUT2 #(
		.INIT('h2)
	) name19695 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w23741_,
		_w23742_
	);
	LUT2 #(
		.INIT('h8)
	) name19696 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_txctl_b_sync1_reg/P0001 ,
		_w23743_
	);
	LUT2 #(
		.INIT('h2)
	) name19697 (
		_w23276_,
		_w23284_,
		_w23744_
	);
	LUT2 #(
		.INIT('h8)
	) name19698 (
		\memc_LDaST_Eg_reg/NET0131 ,
		_w4117_,
		_w23745_
	);
	LUT2 #(
		.INIT('h2)
	) name19699 (
		_w5946_,
		_w11748_,
		_w23746_
	);
	LUT2 #(
		.INIT('h2)
	) name19700 (
		_w13130_,
		_w13580_,
		_w23747_
	);
	LUT2 #(
		.INIT('h1)
	) name19701 (
		_w23746_,
		_w23747_,
		_w23748_
	);
	LUT2 #(
		.INIT('h2)
	) name19702 (
		_w6931_,
		_w23748_,
		_w23749_
	);
	LUT2 #(
		.INIT('h8)
	) name19703 (
		_w11741_,
		_w23749_,
		_w23750_
	);
	LUT2 #(
		.INIT('h1)
	) name19704 (
		_w23745_,
		_w23750_,
		_w23751_
	);
	LUT2 #(
		.INIT('h8)
	) name19705 (
		\memc_selMIO_E_reg/P0001 ,
		_w23235_,
		_w23752_
	);
	LUT2 #(
		.INIT('h1)
	) name19706 (
		_w23238_,
		_w23752_,
		_w23753_
	);
	LUT2 #(
		.INIT('h8)
	) name19707 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		_w14665_,
		_w23754_
	);
	LUT2 #(
		.INIT('h1)
	) name19708 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w8460_,
		_w23755_
	);
	LUT2 #(
		.INIT('h2)
	) name19709 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12590_,
		_w23756_
	);
	LUT2 #(
		.INIT('h1)
	) name19710 (
		_w23755_,
		_w23756_,
		_w23757_
	);
	LUT2 #(
		.INIT('h2)
	) name19711 (
		_w23754_,
		_w23757_,
		_w23758_
	);
	LUT2 #(
		.INIT('h1)
	) name19712 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[11]/P0001 ,
		_w23754_,
		_w23759_
	);
	LUT2 #(
		.INIT('h1)
	) name19713 (
		_w23758_,
		_w23759_,
		_w23760_
	);
	LUT2 #(
		.INIT('h2)
	) name19714 (
		_w6106_,
		_w7859_,
		_w23761_
	);
	LUT2 #(
		.INIT('h4)
	) name19715 (
		_w6106_,
		_w7644_,
		_w23762_
	);
	LUT2 #(
		.INIT('h1)
	) name19716 (
		_w23761_,
		_w23762_,
		_w23763_
	);
	LUT2 #(
		.INIT('h4)
	) name19717 (
		_w6084_,
		_w23763_,
		_w23764_
	);
	LUT2 #(
		.INIT('h1)
	) name19718 (
		_w8133_,
		_w23764_,
		_w23765_
	);
	LUT2 #(
		.INIT('h8)
	) name19719 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		_w14665_,
		_w23766_
	);
	LUT2 #(
		.INIT('h4)
	) name19720 (
		_w21994_,
		_w23766_,
		_w23767_
	);
	LUT2 #(
		.INIT('h1)
	) name19721 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[9]/P0001 ,
		_w23766_,
		_w23768_
	);
	LUT2 #(
		.INIT('h1)
	) name19722 (
		_w23767_,
		_w23768_,
		_w23769_
	);
	LUT2 #(
		.INIT('h2)
	) name19723 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[8]/P0001 ,
		_w23766_,
		_w23770_
	);
	LUT2 #(
		.INIT('h4)
	) name19724 (
		_w22003_,
		_w23766_,
		_w23771_
	);
	LUT2 #(
		.INIT('h1)
	) name19725 (
		_w23770_,
		_w23771_,
		_w23772_
	);
	LUT2 #(
		.INIT('h4)
	) name19726 (
		_w22084_,
		_w23766_,
		_w23773_
	);
	LUT2 #(
		.INIT('h1)
	) name19727 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[13]/P0001 ,
		_w23766_,
		_w23774_
	);
	LUT2 #(
		.INIT('h1)
	) name19728 (
		_w23773_,
		_w23774_,
		_w23775_
	);
	LUT2 #(
		.INIT('h2)
	) name19729 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[12]/P0001 ,
		_w23766_,
		_w23776_
	);
	LUT2 #(
		.INIT('h4)
	) name19730 (
		_w22093_,
		_w23766_,
		_w23777_
	);
	LUT2 #(
		.INIT('h1)
	) name19731 (
		_w23776_,
		_w23777_,
		_w23778_
	);
	LUT2 #(
		.INIT('h2)
	) name19732 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[11]/P0001 ,
		_w23766_,
		_w23779_
	);
	LUT2 #(
		.INIT('h4)
	) name19733 (
		_w22105_,
		_w23766_,
		_w23780_
	);
	LUT2 #(
		.INIT('h1)
	) name19734 (
		_w23779_,
		_w23780_,
		_w23781_
	);
	LUT2 #(
		.INIT('h8)
	) name19735 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		_w17798_,
		_w23782_
	);
	LUT2 #(
		.INIT('h4)
	) name19736 (
		_w21994_,
		_w23782_,
		_w23783_
	);
	LUT2 #(
		.INIT('h1)
	) name19737 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[9]/P0001 ,
		_w23782_,
		_w23784_
	);
	LUT2 #(
		.INIT('h1)
	) name19738 (
		_w23783_,
		_w23784_,
		_w23785_
	);
	LUT2 #(
		.INIT('h4)
	) name19739 (
		_w22084_,
		_w23782_,
		_w23786_
	);
	LUT2 #(
		.INIT('h1)
	) name19740 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[13]/P0001 ,
		_w23782_,
		_w23787_
	);
	LUT2 #(
		.INIT('h1)
	) name19741 (
		_w23786_,
		_w23787_,
		_w23788_
	);
	LUT2 #(
		.INIT('h2)
	) name19742 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[12]/P0001 ,
		_w23782_,
		_w23789_
	);
	LUT2 #(
		.INIT('h4)
	) name19743 (
		_w22093_,
		_w23782_,
		_w23790_
	);
	LUT2 #(
		.INIT('h1)
	) name19744 (
		_w23789_,
		_w23790_,
		_w23791_
	);
	LUT2 #(
		.INIT('h2)
	) name19745 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[11]/P0001 ,
		_w23782_,
		_w23792_
	);
	LUT2 #(
		.INIT('h4)
	) name19746 (
		_w22105_,
		_w23782_,
		_w23793_
	);
	LUT2 #(
		.INIT('h1)
	) name19747 (
		_w23792_,
		_w23793_,
		_w23794_
	);
	LUT2 #(
		.INIT('h4)
	) name19748 (
		_w22114_,
		_w23782_,
		_w23795_
	);
	LUT2 #(
		.INIT('h1)
	) name19749 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[10]/P0001 ,
		_w23782_,
		_w23796_
	);
	LUT2 #(
		.INIT('h1)
	) name19750 (
		_w23795_,
		_w23796_,
		_w23797_
	);
	LUT2 #(
		.INIT('h8)
	) name19751 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		_w14665_,
		_w23798_
	);
	LUT2 #(
		.INIT('h4)
	) name19752 (
		_w21994_,
		_w23798_,
		_w23799_
	);
	LUT2 #(
		.INIT('h1)
	) name19753 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[9]/P0001 ,
		_w23798_,
		_w23800_
	);
	LUT2 #(
		.INIT('h1)
	) name19754 (
		_w23799_,
		_w23800_,
		_w23801_
	);
	LUT2 #(
		.INIT('h2)
	) name19755 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[8]/P0001 ,
		_w23798_,
		_w23802_
	);
	LUT2 #(
		.INIT('h4)
	) name19756 (
		_w22003_,
		_w23798_,
		_w23803_
	);
	LUT2 #(
		.INIT('h1)
	) name19757 (
		_w23802_,
		_w23803_,
		_w23804_
	);
	LUT2 #(
		.INIT('h2)
	) name19758 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[12]/P0001 ,
		_w23798_,
		_w23805_
	);
	LUT2 #(
		.INIT('h4)
	) name19759 (
		_w22093_,
		_w23798_,
		_w23806_
	);
	LUT2 #(
		.INIT('h1)
	) name19760 (
		_w23805_,
		_w23806_,
		_w23807_
	);
	LUT2 #(
		.INIT('h2)
	) name19761 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[11]/P0001 ,
		_w23798_,
		_w23808_
	);
	LUT2 #(
		.INIT('h4)
	) name19762 (
		_w22105_,
		_w23798_,
		_w23809_
	);
	LUT2 #(
		.INIT('h1)
	) name19763 (
		_w23808_,
		_w23809_,
		_w23810_
	);
	LUT2 #(
		.INIT('h4)
	) name19764 (
		_w22114_,
		_w23798_,
		_w23811_
	);
	LUT2 #(
		.INIT('h1)
	) name19765 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[10]/P0001 ,
		_w23798_,
		_w23812_
	);
	LUT2 #(
		.INIT('h1)
	) name19766 (
		_w23811_,
		_w23812_,
		_w23813_
	);
	LUT2 #(
		.INIT('h8)
	) name19767 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		_w17798_,
		_w23814_
	);
	LUT2 #(
		.INIT('h4)
	) name19768 (
		_w21994_,
		_w23814_,
		_w23815_
	);
	LUT2 #(
		.INIT('h1)
	) name19769 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[9]/P0001 ,
		_w23814_,
		_w23816_
	);
	LUT2 #(
		.INIT('h1)
	) name19770 (
		_w23815_,
		_w23816_,
		_w23817_
	);
	LUT2 #(
		.INIT('h2)
	) name19771 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[8]/P0001 ,
		_w23814_,
		_w23818_
	);
	LUT2 #(
		.INIT('h4)
	) name19772 (
		_w22003_,
		_w23814_,
		_w23819_
	);
	LUT2 #(
		.INIT('h1)
	) name19773 (
		_w23818_,
		_w23819_,
		_w23820_
	);
	LUT2 #(
		.INIT('h2)
	) name19774 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[12]/P0001 ,
		_w23814_,
		_w23821_
	);
	LUT2 #(
		.INIT('h4)
	) name19775 (
		_w22093_,
		_w23814_,
		_w23822_
	);
	LUT2 #(
		.INIT('h1)
	) name19776 (
		_w23821_,
		_w23822_,
		_w23823_
	);
	LUT2 #(
		.INIT('h4)
	) name19777 (
		_w22114_,
		_w23814_,
		_w23824_
	);
	LUT2 #(
		.INIT('h1)
	) name19778 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[10]/P0001 ,
		_w23814_,
		_w23825_
	);
	LUT2 #(
		.INIT('h1)
	) name19779 (
		_w23824_,
		_w23825_,
		_w23826_
	);
	LUT2 #(
		.INIT('h8)
	) name19780 (
		_w7530_,
		_w13762_,
		_w23827_
	);
	LUT2 #(
		.INIT('h4)
	) name19781 (
		_w10289_,
		_w23827_,
		_w23828_
	);
	LUT2 #(
		.INIT('h1)
	) name19782 (
		\bdma_BOVL_reg[9]/NET0131 ,
		_w23827_,
		_w23829_
	);
	LUT2 #(
		.INIT('h1)
	) name19783 (
		_w23828_,
		_w23829_,
		_w23830_
	);
	LUT2 #(
		.INIT('h4)
	) name19784 (
		_w10638_,
		_w23827_,
		_w23831_
	);
	LUT2 #(
		.INIT('h1)
	) name19785 (
		\bdma_BOVL_reg[8]/NET0131 ,
		_w23827_,
		_w23832_
	);
	LUT2 #(
		.INIT('h1)
	) name19786 (
		_w23831_,
		_w23832_,
		_w23833_
	);
	LUT2 #(
		.INIT('h4)
	) name19787 (
		_w8460_,
		_w23827_,
		_w23834_
	);
	LUT2 #(
		.INIT('h1)
	) name19788 (
		\bdma_BOVL_reg[11]/NET0131 ,
		_w23827_,
		_w23835_
	);
	LUT2 #(
		.INIT('h1)
	) name19789 (
		_w23834_,
		_w23835_,
		_w23836_
	);
	LUT2 #(
		.INIT('h4)
	) name19790 (
		_w7859_,
		_w23827_,
		_w23837_
	);
	LUT2 #(
		.INIT('h1)
	) name19791 (
		\bdma_BOVL_reg[10]/NET0131 ,
		_w23827_,
		_w23838_
	);
	LUT2 #(
		.INIT('h1)
	) name19792 (
		_w23837_,
		_w23838_,
		_w23839_
	);
	LUT2 #(
		.INIT('h4)
	) name19793 (
		_w10289_,
		_w21268_,
		_w23840_
	);
	LUT2 #(
		.INIT('h1)
	) name19794 (
		\bdma_BCTL_reg[9]/NET0131 ,
		_w21268_,
		_w23841_
	);
	LUT2 #(
		.INIT('h1)
	) name19795 (
		_w23840_,
		_w23841_,
		_w23842_
	);
	LUT2 #(
		.INIT('h4)
	) name19796 (
		_w10638_,
		_w21268_,
		_w23843_
	);
	LUT2 #(
		.INIT('h1)
	) name19797 (
		\bdma_BCTL_reg[8]/NET0131 ,
		_w21268_,
		_w23844_
	);
	LUT2 #(
		.INIT('h1)
	) name19798 (
		_w23843_,
		_w23844_,
		_w23845_
	);
	LUT2 #(
		.INIT('h4)
	) name19799 (
		_w7340_,
		_w21268_,
		_w23846_
	);
	LUT2 #(
		.INIT('h1)
	) name19800 (
		\bdma_BCTL_reg[13]/NET0131 ,
		_w21268_,
		_w23847_
	);
	LUT2 #(
		.INIT('h1)
	) name19801 (
		_w23846_,
		_w23847_,
		_w23848_
	);
	LUT2 #(
		.INIT('h4)
	) name19802 (
		_w9178_,
		_w21268_,
		_w23849_
	);
	LUT2 #(
		.INIT('h1)
	) name19803 (
		\bdma_BCTL_reg[12]/NET0131 ,
		_w21268_,
		_w23850_
	);
	LUT2 #(
		.INIT('h1)
	) name19804 (
		_w23849_,
		_w23850_,
		_w23851_
	);
	LUT2 #(
		.INIT('h4)
	) name19805 (
		_w8460_,
		_w21268_,
		_w23852_
	);
	LUT2 #(
		.INIT('h1)
	) name19806 (
		\bdma_BCTL_reg[11]/NET0131 ,
		_w21268_,
		_w23853_
	);
	LUT2 #(
		.INIT('h1)
	) name19807 (
		_w23852_,
		_w23853_,
		_w23854_
	);
	LUT2 #(
		.INIT('h4)
	) name19808 (
		_w7859_,
		_w21268_,
		_w23855_
	);
	LUT2 #(
		.INIT('h1)
	) name19809 (
		\bdma_BCTL_reg[10]/NET0131 ,
		_w21268_,
		_w23856_
	);
	LUT2 #(
		.INIT('h1)
	) name19810 (
		_w23855_,
		_w23856_,
		_w23857_
	);
	LUT2 #(
		.INIT('h1)
	) name19811 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w10638_,
		_w23858_
	);
	LUT2 #(
		.INIT('h2)
	) name19812 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w13041_,
		_w23859_
	);
	LUT2 #(
		.INIT('h1)
	) name19813 (
		_w23858_,
		_w23859_,
		_w23860_
	);
	LUT2 #(
		.INIT('h2)
	) name19814 (
		_w23754_,
		_w23860_,
		_w23861_
	);
	LUT2 #(
		.INIT('h1)
	) name19815 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[8]/P0001 ,
		_w23754_,
		_w23862_
	);
	LUT2 #(
		.INIT('h1)
	) name19816 (
		_w23861_,
		_w23862_,
		_w23863_
	);
	LUT2 #(
		.INIT('h8)
	) name19817 (
		\core_c_dec_MTTX1_E_reg/P0001 ,
		_w5951_,
		_w23864_
	);
	LUT2 #(
		.INIT('h1)
	) name19818 (
		\auctl_T1Sack_reg/NET0131 ,
		_w23864_,
		_w23865_
	);
	LUT2 #(
		.INIT('h2)
	) name19819 (
		_w10289_,
		_w23865_,
		_w23866_
	);
	LUT2 #(
		.INIT('h8)
	) name19820 (
		\sport1_txctl_TX_reg[9]/P0001 ,
		_w23865_,
		_w23867_
	);
	LUT2 #(
		.INIT('h1)
	) name19821 (
		_w23866_,
		_w23867_,
		_w23868_
	);
	LUT2 #(
		.INIT('h2)
	) name19822 (
		_w10638_,
		_w23865_,
		_w23869_
	);
	LUT2 #(
		.INIT('h8)
	) name19823 (
		\sport1_txctl_TX_reg[8]/P0001 ,
		_w23865_,
		_w23870_
	);
	LUT2 #(
		.INIT('h1)
	) name19824 (
		_w23869_,
		_w23870_,
		_w23871_
	);
	LUT2 #(
		.INIT('h2)
	) name19825 (
		_w9178_,
		_w23865_,
		_w23872_
	);
	LUT2 #(
		.INIT('h8)
	) name19826 (
		\sport1_txctl_TX_reg[12]/P0001 ,
		_w23865_,
		_w23873_
	);
	LUT2 #(
		.INIT('h1)
	) name19827 (
		_w23872_,
		_w23873_,
		_w23874_
	);
	LUT2 #(
		.INIT('h2)
	) name19828 (
		_w8460_,
		_w23865_,
		_w23875_
	);
	LUT2 #(
		.INIT('h8)
	) name19829 (
		\sport1_txctl_TX_reg[11]/P0001 ,
		_w23865_,
		_w23876_
	);
	LUT2 #(
		.INIT('h1)
	) name19830 (
		_w23875_,
		_w23876_,
		_w23877_
	);
	LUT2 #(
		.INIT('h2)
	) name19831 (
		_w7859_,
		_w23865_,
		_w23878_
	);
	LUT2 #(
		.INIT('h8)
	) name19832 (
		\sport1_txctl_TX_reg[10]/P0001 ,
		_w23865_,
		_w23879_
	);
	LUT2 #(
		.INIT('h1)
	) name19833 (
		_w23878_,
		_w23879_,
		_w23880_
	);
	LUT2 #(
		.INIT('h2)
	) name19834 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[8]/P0001 ,
		_w23782_,
		_w23881_
	);
	LUT2 #(
		.INIT('h4)
	) name19835 (
		_w22003_,
		_w23782_,
		_w23882_
	);
	LUT2 #(
		.INIT('h1)
	) name19836 (
		_w23881_,
		_w23882_,
		_w23883_
	);
	LUT2 #(
		.INIT('h2)
	) name19837 (
		_w6106_,
		_w8113_,
		_w23884_
	);
	LUT2 #(
		.INIT('h4)
	) name19838 (
		_w6106_,
		_w8224_,
		_w23885_
	);
	LUT2 #(
		.INIT('h1)
	) name19839 (
		_w23884_,
		_w23885_,
		_w23886_
	);
	LUT2 #(
		.INIT('h4)
	) name19840 (
		_w6084_,
		_w23886_,
		_w23887_
	);
	LUT2 #(
		.INIT('h1)
	) name19841 (
		_w8177_,
		_w23887_,
		_w23888_
	);
	LUT2 #(
		.INIT('h8)
	) name19842 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		_w14665_,
		_w23889_
	);
	LUT2 #(
		.INIT('h4)
	) name19843 (
		_w21994_,
		_w23889_,
		_w23890_
	);
	LUT2 #(
		.INIT('h1)
	) name19844 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[9]/P0001 ,
		_w23889_,
		_w23891_
	);
	LUT2 #(
		.INIT('h1)
	) name19845 (
		_w23890_,
		_w23891_,
		_w23892_
	);
	LUT2 #(
		.INIT('h2)
	) name19846 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[8]/P0001 ,
		_w23889_,
		_w23893_
	);
	LUT2 #(
		.INIT('h4)
	) name19847 (
		_w22003_,
		_w23889_,
		_w23894_
	);
	LUT2 #(
		.INIT('h1)
	) name19848 (
		_w23893_,
		_w23894_,
		_w23895_
	);
	LUT2 #(
		.INIT('h4)
	) name19849 (
		_w22084_,
		_w23889_,
		_w23896_
	);
	LUT2 #(
		.INIT('h1)
	) name19850 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[13]/P0001 ,
		_w23889_,
		_w23897_
	);
	LUT2 #(
		.INIT('h1)
	) name19851 (
		_w23896_,
		_w23897_,
		_w23898_
	);
	LUT2 #(
		.INIT('h2)
	) name19852 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[12]/P0001 ,
		_w23889_,
		_w23899_
	);
	LUT2 #(
		.INIT('h4)
	) name19853 (
		_w22093_,
		_w23889_,
		_w23900_
	);
	LUT2 #(
		.INIT('h1)
	) name19854 (
		_w23899_,
		_w23900_,
		_w23901_
	);
	LUT2 #(
		.INIT('h2)
	) name19855 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[11]/P0001 ,
		_w23889_,
		_w23902_
	);
	LUT2 #(
		.INIT('h4)
	) name19856 (
		_w22105_,
		_w23889_,
		_w23903_
	);
	LUT2 #(
		.INIT('h1)
	) name19857 (
		_w23902_,
		_w23903_,
		_w23904_
	);
	LUT2 #(
		.INIT('h4)
	) name19858 (
		_w22114_,
		_w23889_,
		_w23905_
	);
	LUT2 #(
		.INIT('h1)
	) name19859 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[10]/P0001 ,
		_w23889_,
		_w23906_
	);
	LUT2 #(
		.INIT('h1)
	) name19860 (
		_w23905_,
		_w23906_,
		_w23907_
	);
	LUT2 #(
		.INIT('h8)
	) name19861 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		_w14665_,
		_w23908_
	);
	LUT2 #(
		.INIT('h4)
	) name19862 (
		_w19504_,
		_w23908_,
		_w23909_
	);
	LUT2 #(
		.INIT('h1)
	) name19863 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[9]/P0001 ,
		_w23908_,
		_w23910_
	);
	LUT2 #(
		.INIT('h1)
	) name19864 (
		_w23909_,
		_w23910_,
		_w23911_
	);
	LUT2 #(
		.INIT('h4)
	) name19865 (
		_w23860_,
		_w23908_,
		_w23912_
	);
	LUT2 #(
		.INIT('h1)
	) name19866 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[8]/P0001 ,
		_w23908_,
		_w23913_
	);
	LUT2 #(
		.INIT('h1)
	) name19867 (
		_w23912_,
		_w23913_,
		_w23914_
	);
	LUT2 #(
		.INIT('h4)
	) name19868 (
		_w17836_,
		_w23908_,
		_w23915_
	);
	LUT2 #(
		.INIT('h1)
	) name19869 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[13]/P0001 ,
		_w23908_,
		_w23916_
	);
	LUT2 #(
		.INIT('h1)
	) name19870 (
		_w23915_,
		_w23916_,
		_w23917_
	);
	LUT2 #(
		.INIT('h1)
	) name19871 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w9178_,
		_w23918_
	);
	LUT2 #(
		.INIT('h2)
	) name19872 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w12624_,
		_w23919_
	);
	LUT2 #(
		.INIT('h1)
	) name19873 (
		_w23918_,
		_w23919_,
		_w23920_
	);
	LUT2 #(
		.INIT('h2)
	) name19874 (
		_w23908_,
		_w23920_,
		_w23921_
	);
	LUT2 #(
		.INIT('h1)
	) name19875 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[12]/P0001 ,
		_w23908_,
		_w23922_
	);
	LUT2 #(
		.INIT('h1)
	) name19876 (
		_w23921_,
		_w23922_,
		_w23923_
	);
	LUT2 #(
		.INIT('h4)
	) name19877 (
		_w23757_,
		_w23908_,
		_w23924_
	);
	LUT2 #(
		.INIT('h1)
	) name19878 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[11]/P0001 ,
		_w23908_,
		_w23925_
	);
	LUT2 #(
		.INIT('h1)
	) name19879 (
		_w23924_,
		_w23925_,
		_w23926_
	);
	LUT2 #(
		.INIT('h4)
	) name19880 (
		_w19848_,
		_w23908_,
		_w23927_
	);
	LUT2 #(
		.INIT('h1)
	) name19881 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[10]/P0001 ,
		_w23908_,
		_w23928_
	);
	LUT2 #(
		.INIT('h1)
	) name19882 (
		_w23927_,
		_w23928_,
		_w23929_
	);
	LUT2 #(
		.INIT('h8)
	) name19883 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		_w14665_,
		_w23930_
	);
	LUT2 #(
		.INIT('h4)
	) name19884 (
		_w19504_,
		_w23930_,
		_w23931_
	);
	LUT2 #(
		.INIT('h1)
	) name19885 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[9]/P0001 ,
		_w23930_,
		_w23932_
	);
	LUT2 #(
		.INIT('h1)
	) name19886 (
		_w23931_,
		_w23932_,
		_w23933_
	);
	LUT2 #(
		.INIT('h4)
	) name19887 (
		_w23860_,
		_w23930_,
		_w23934_
	);
	LUT2 #(
		.INIT('h1)
	) name19888 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[8]/P0001 ,
		_w23930_,
		_w23935_
	);
	LUT2 #(
		.INIT('h1)
	) name19889 (
		_w23934_,
		_w23935_,
		_w23936_
	);
	LUT2 #(
		.INIT('h4)
	) name19890 (
		_w17836_,
		_w23930_,
		_w23937_
	);
	LUT2 #(
		.INIT('h1)
	) name19891 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[13]/P0001 ,
		_w23930_,
		_w23938_
	);
	LUT2 #(
		.INIT('h1)
	) name19892 (
		_w23937_,
		_w23938_,
		_w23939_
	);
	LUT2 #(
		.INIT('h4)
	) name19893 (
		_w23920_,
		_w23930_,
		_w23940_
	);
	LUT2 #(
		.INIT('h1)
	) name19894 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[12]/P0001 ,
		_w23930_,
		_w23941_
	);
	LUT2 #(
		.INIT('h1)
	) name19895 (
		_w23940_,
		_w23941_,
		_w23942_
	);
	LUT2 #(
		.INIT('h4)
	) name19896 (
		_w23757_,
		_w23930_,
		_w23943_
	);
	LUT2 #(
		.INIT('h1)
	) name19897 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[11]/P0001 ,
		_w23930_,
		_w23944_
	);
	LUT2 #(
		.INIT('h1)
	) name19898 (
		_w23943_,
		_w23944_,
		_w23945_
	);
	LUT2 #(
		.INIT('h4)
	) name19899 (
		_w19848_,
		_w23930_,
		_w23946_
	);
	LUT2 #(
		.INIT('h1)
	) name19900 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[10]/P0001 ,
		_w23930_,
		_w23947_
	);
	LUT2 #(
		.INIT('h1)
	) name19901 (
		_w23946_,
		_w23947_,
		_w23948_
	);
	LUT2 #(
		.INIT('h2)
	) name19902 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[11]/P0001 ,
		_w23814_,
		_w23949_
	);
	LUT2 #(
		.INIT('h4)
	) name19903 (
		_w22105_,
		_w23814_,
		_w23950_
	);
	LUT2 #(
		.INIT('h1)
	) name19904 (
		_w23949_,
		_w23950_,
		_w23951_
	);
	LUT2 #(
		.INIT('h4)
	) name19905 (
		_w22084_,
		_w23814_,
		_w23952_
	);
	LUT2 #(
		.INIT('h1)
	) name19906 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[13]/P0001 ,
		_w23814_,
		_w23953_
	);
	LUT2 #(
		.INIT('h1)
	) name19907 (
		_w23952_,
		_w23953_,
		_w23954_
	);
	LUT2 #(
		.INIT('h4)
	) name19908 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIreg_E_reg[7]/P0001 ,
		_w23955_
	);
	LUT2 #(
		.INIT('h1)
	) name19909 (
		_w5999_,
		_w23955_,
		_w23956_
	);
	LUT2 #(
		.INIT('h4)
	) name19910 (
		_w5994_,
		_w23956_,
		_w23957_
	);
	LUT2 #(
		.INIT('h1)
	) name19911 (
		_w6000_,
		_w23957_,
		_w23958_
	);
	LUT2 #(
		.INIT('h2)
	) name19912 (
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w23958_,
		_w23959_
	);
	LUT2 #(
		.INIT('h4)
	) name19913 (
		_w6000_,
		_w20755_,
		_w23960_
	);
	LUT2 #(
		.INIT('h1)
	) name19914 (
		_w23959_,
		_w23960_,
		_w23961_
	);
	LUT2 #(
		.INIT('h2)
	) name19915 (
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w23958_,
		_w23962_
	);
	LUT2 #(
		.INIT('h4)
	) name19916 (
		_w6000_,
		_w20624_,
		_w23963_
	);
	LUT2 #(
		.INIT('h1)
	) name19917 (
		_w23962_,
		_w23963_,
		_w23964_
	);
	LUT2 #(
		.INIT('h2)
	) name19918 (
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w23958_,
		_w23965_
	);
	LUT2 #(
		.INIT('h4)
	) name19919 (
		_w6000_,
		_w20634_,
		_w23966_
	);
	LUT2 #(
		.INIT('h1)
	) name19920 (
		_w23965_,
		_w23966_,
		_w23967_
	);
	LUT2 #(
		.INIT('h2)
	) name19921 (
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w23958_,
		_w23968_
	);
	LUT2 #(
		.INIT('h1)
	) name19922 (
		_w6000_,
		_w20685_,
		_w23969_
	);
	LUT2 #(
		.INIT('h1)
	) name19923 (
		_w23968_,
		_w23969_,
		_w23970_
	);
	LUT2 #(
		.INIT('h2)
	) name19924 (
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w23958_,
		_w23971_
	);
	LUT2 #(
		.INIT('h1)
	) name19925 (
		_w6000_,
		_w20696_,
		_w23972_
	);
	LUT2 #(
		.INIT('h1)
	) name19926 (
		_w23971_,
		_w23972_,
		_w23973_
	);
	LUT2 #(
		.INIT('h4)
	) name19927 (
		_w6008_,
		_w20755_,
		_w23974_
	);
	LUT2 #(
		.INIT('h8)
	) name19928 (
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w6008_,
		_w23975_
	);
	LUT2 #(
		.INIT('h1)
	) name19929 (
		_w23974_,
		_w23975_,
		_w23976_
	);
	LUT2 #(
		.INIT('h4)
	) name19930 (
		_w6008_,
		_w20602_,
		_w23977_
	);
	LUT2 #(
		.INIT('h8)
	) name19931 (
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w6008_,
		_w23978_
	);
	LUT2 #(
		.INIT('h1)
	) name19932 (
		_w23977_,
		_w23978_,
		_w23979_
	);
	LUT2 #(
		.INIT('h4)
	) name19933 (
		_w6008_,
		_w20614_,
		_w23980_
	);
	LUT2 #(
		.INIT('h8)
	) name19934 (
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w6008_,
		_w23981_
	);
	LUT2 #(
		.INIT('h1)
	) name19935 (
		_w23980_,
		_w23981_,
		_w23982_
	);
	LUT2 #(
		.INIT('h4)
	) name19936 (
		_w6008_,
		_w20624_,
		_w23983_
	);
	LUT2 #(
		.INIT('h8)
	) name19937 (
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w6008_,
		_w23984_
	);
	LUT2 #(
		.INIT('h1)
	) name19938 (
		_w23983_,
		_w23984_,
		_w23985_
	);
	LUT2 #(
		.INIT('h4)
	) name19939 (
		_w6008_,
		_w20634_,
		_w23986_
	);
	LUT2 #(
		.INIT('h8)
	) name19940 (
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w6008_,
		_w23987_
	);
	LUT2 #(
		.INIT('h1)
	) name19941 (
		_w23986_,
		_w23987_,
		_w23988_
	);
	LUT2 #(
		.INIT('h1)
	) name19942 (
		_w6008_,
		_w20685_,
		_w23989_
	);
	LUT2 #(
		.INIT('h8)
	) name19943 (
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w6008_,
		_w23990_
	);
	LUT2 #(
		.INIT('h1)
	) name19944 (
		_w23989_,
		_w23990_,
		_w23991_
	);
	LUT2 #(
		.INIT('h1)
	) name19945 (
		_w6008_,
		_w20696_,
		_w23992_
	);
	LUT2 #(
		.INIT('h8)
	) name19946 (
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w6008_,
		_w23993_
	);
	LUT2 #(
		.INIT('h1)
	) name19947 (
		_w23992_,
		_w23993_,
		_w23994_
	);
	LUT2 #(
		.INIT('h1)
	) name19948 (
		_w6008_,
		_w20707_,
		_w23995_
	);
	LUT2 #(
		.INIT('h8)
	) name19949 (
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w6008_,
		_w23996_
	);
	LUT2 #(
		.INIT('h1)
	) name19950 (
		_w23995_,
		_w23996_,
		_w23997_
	);
	LUT2 #(
		.INIT('h4)
	) name19951 (
		_w6008_,
		_w20718_,
		_w23998_
	);
	LUT2 #(
		.INIT('h8)
	) name19952 (
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w6008_,
		_w23999_
	);
	LUT2 #(
		.INIT('h1)
	) name19953 (
		_w23998_,
		_w23999_,
		_w24000_
	);
	LUT2 #(
		.INIT('h4)
	) name19954 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIreg_E_reg[5]/P0001 ,
		_w24001_
	);
	LUT2 #(
		.INIT('h1)
	) name19955 (
		_w6014_,
		_w24001_,
		_w24002_
	);
	LUT2 #(
		.INIT('h4)
	) name19956 (
		_w6011_,
		_w24002_,
		_w24003_
	);
	LUT2 #(
		.INIT('h1)
	) name19957 (
		_w6015_,
		_w24003_,
		_w24004_
	);
	LUT2 #(
		.INIT('h2)
	) name19958 (
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w24004_,
		_w24005_
	);
	LUT2 #(
		.INIT('h4)
	) name19959 (
		_w6015_,
		_w20755_,
		_w24006_
	);
	LUT2 #(
		.INIT('h1)
	) name19960 (
		_w24005_,
		_w24006_,
		_w24007_
	);
	LUT2 #(
		.INIT('h2)
	) name19961 (
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		_w24004_,
		_w24008_
	);
	LUT2 #(
		.INIT('h4)
	) name19962 (
		_w6015_,
		_w20624_,
		_w24009_
	);
	LUT2 #(
		.INIT('h1)
	) name19963 (
		_w24008_,
		_w24009_,
		_w24010_
	);
	LUT2 #(
		.INIT('h2)
	) name19964 (
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		_w24004_,
		_w24011_
	);
	LUT2 #(
		.INIT('h4)
	) name19965 (
		_w6015_,
		_w20634_,
		_w24012_
	);
	LUT2 #(
		.INIT('h1)
	) name19966 (
		_w24011_,
		_w24012_,
		_w24013_
	);
	LUT2 #(
		.INIT('h2)
	) name19967 (
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		_w24004_,
		_w24014_
	);
	LUT2 #(
		.INIT('h1)
	) name19968 (
		_w6015_,
		_w20685_,
		_w24015_
	);
	LUT2 #(
		.INIT('h1)
	) name19969 (
		_w24014_,
		_w24015_,
		_w24016_
	);
	LUT2 #(
		.INIT('h2)
	) name19970 (
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		_w24004_,
		_w24017_
	);
	LUT2 #(
		.INIT('h1)
	) name19971 (
		_w6015_,
		_w20696_,
		_w24018_
	);
	LUT2 #(
		.INIT('h1)
	) name19972 (
		_w24017_,
		_w24018_,
		_w24019_
	);
	LUT2 #(
		.INIT('h4)
	) name19973 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIreg_E_reg[4]/P0001 ,
		_w24020_
	);
	LUT2 #(
		.INIT('h1)
	) name19974 (
		_w5963_,
		_w24020_,
		_w24021_
	);
	LUT2 #(
		.INIT('h4)
	) name19975 (
		_w5958_,
		_w24021_,
		_w24022_
	);
	LUT2 #(
		.INIT('h1)
	) name19976 (
		_w5964_,
		_w24022_,
		_w24023_
	);
	LUT2 #(
		.INIT('h2)
	) name19977 (
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w24023_,
		_w24024_
	);
	LUT2 #(
		.INIT('h4)
	) name19978 (
		_w5964_,
		_w20755_,
		_w24025_
	);
	LUT2 #(
		.INIT('h1)
	) name19979 (
		_w24024_,
		_w24025_,
		_w24026_
	);
	LUT2 #(
		.INIT('h2)
	) name19980 (
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		_w24023_,
		_w24027_
	);
	LUT2 #(
		.INIT('h8)
	) name19981 (
		_w20602_,
		_w24023_,
		_w24028_
	);
	LUT2 #(
		.INIT('h1)
	) name19982 (
		_w24027_,
		_w24028_,
		_w24029_
	);
	LUT2 #(
		.INIT('h2)
	) name19983 (
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w24023_,
		_w24030_
	);
	LUT2 #(
		.INIT('h8)
	) name19984 (
		_w20614_,
		_w24023_,
		_w24031_
	);
	LUT2 #(
		.INIT('h1)
	) name19985 (
		_w24030_,
		_w24031_,
		_w24032_
	);
	LUT2 #(
		.INIT('h2)
	) name19986 (
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w24023_,
		_w24033_
	);
	LUT2 #(
		.INIT('h4)
	) name19987 (
		_w5964_,
		_w20624_,
		_w24034_
	);
	LUT2 #(
		.INIT('h1)
	) name19988 (
		_w24033_,
		_w24034_,
		_w24035_
	);
	LUT2 #(
		.INIT('h2)
	) name19989 (
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w24023_,
		_w24036_
	);
	LUT2 #(
		.INIT('h4)
	) name19990 (
		_w5964_,
		_w20634_,
		_w24037_
	);
	LUT2 #(
		.INIT('h1)
	) name19991 (
		_w24036_,
		_w24037_,
		_w24038_
	);
	LUT2 #(
		.INIT('h2)
	) name19992 (
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w24023_,
		_w24039_
	);
	LUT2 #(
		.INIT('h1)
	) name19993 (
		_w5964_,
		_w20685_,
		_w24040_
	);
	LUT2 #(
		.INIT('h1)
	) name19994 (
		_w24039_,
		_w24040_,
		_w24041_
	);
	LUT2 #(
		.INIT('h2)
	) name19995 (
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w24023_,
		_w24042_
	);
	LUT2 #(
		.INIT('h1)
	) name19996 (
		_w5964_,
		_w20696_,
		_w24043_
	);
	LUT2 #(
		.INIT('h1)
	) name19997 (
		_w24042_,
		_w24043_,
		_w24044_
	);
	LUT2 #(
		.INIT('h4)
	) name19998 (
		_w20707_,
		_w24023_,
		_w24045_
	);
	LUT2 #(
		.INIT('h2)
	) name19999 (
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		_w24023_,
		_w24046_
	);
	LUT2 #(
		.INIT('h1)
	) name20000 (
		_w24045_,
		_w24046_,
		_w24047_
	);
	LUT2 #(
		.INIT('h4)
	) name20001 (
		_w20718_,
		_w24023_,
		_w24048_
	);
	LUT2 #(
		.INIT('h1)
	) name20002 (
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		_w24023_,
		_w24049_
	);
	LUT2 #(
		.INIT('h1)
	) name20003 (
		_w24048_,
		_w24049_,
		_w24050_
	);
	LUT2 #(
		.INIT('h4)
	) name20004 (
		_w19504_,
		_w23754_,
		_w24051_
	);
	LUT2 #(
		.INIT('h1)
	) name20005 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[9]/P0001 ,
		_w23754_,
		_w24052_
	);
	LUT2 #(
		.INIT('h1)
	) name20006 (
		_w24051_,
		_w24052_,
		_w24053_
	);
	LUT2 #(
		.INIT('h2)
	) name20007 (
		_w23754_,
		_w23920_,
		_w24054_
	);
	LUT2 #(
		.INIT('h1)
	) name20008 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[12]/P0001 ,
		_w23754_,
		_w24055_
	);
	LUT2 #(
		.INIT('h1)
	) name20009 (
		_w24054_,
		_w24055_,
		_w24056_
	);
	LUT2 #(
		.INIT('h4)
	) name20010 (
		_w22084_,
		_w23798_,
		_w24057_
	);
	LUT2 #(
		.INIT('h1)
	) name20011 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[13]/P0001 ,
		_w23798_,
		_w24058_
	);
	LUT2 #(
		.INIT('h1)
	) name20012 (
		_w24057_,
		_w24058_,
		_w24059_
	);
	LUT2 #(
		.INIT('h2)
	) name20013 (
		_w6106_,
		_w10638_,
		_w24060_
	);
	LUT2 #(
		.INIT('h4)
	) name20014 (
		_w6106_,
		_w10343_,
		_w24061_
	);
	LUT2 #(
		.INIT('h1)
	) name20015 (
		_w24060_,
		_w24061_,
		_w24062_
	);
	LUT2 #(
		.INIT('h4)
	) name20016 (
		_w6075_,
		_w24062_,
		_w24063_
	);
	LUT2 #(
		.INIT('h8)
	) name20017 (
		\core_dag_ilm1reg_I3_we_DO_reg[8]/NET0131 ,
		_w6075_,
		_w24064_
	);
	LUT2 #(
		.INIT('h1)
	) name20018 (
		_w24063_,
		_w24064_,
		_w24065_
	);
	LUT2 #(
		.INIT('h2)
	) name20019 (
		_w6106_,
		_w10911_,
		_w24066_
	);
	LUT2 #(
		.INIT('h4)
	) name20020 (
		_w6106_,
		_w10663_,
		_w24067_
	);
	LUT2 #(
		.INIT('h1)
	) name20021 (
		_w24066_,
		_w24067_,
		_w24068_
	);
	LUT2 #(
		.INIT('h1)
	) name20022 (
		_w6075_,
		_w24068_,
		_w24069_
	);
	LUT2 #(
		.INIT('h4)
	) name20023 (
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w6075_,
		_w24070_
	);
	LUT2 #(
		.INIT('h1)
	) name20024 (
		_w24069_,
		_w24070_,
		_w24071_
	);
	LUT2 #(
		.INIT('h2)
	) name20025 (
		_w6106_,
		_w9435_,
		_w24072_
	);
	LUT2 #(
		.INIT('h4)
	) name20026 (
		_w6106_,
		_w8926_,
		_w24073_
	);
	LUT2 #(
		.INIT('h1)
	) name20027 (
		_w24072_,
		_w24073_,
		_w24074_
	);
	LUT2 #(
		.INIT('h1)
	) name20028 (
		_w6075_,
		_w24074_,
		_w24075_
	);
	LUT2 #(
		.INIT('h4)
	) name20029 (
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w6075_,
		_w24076_
	);
	LUT2 #(
		.INIT('h1)
	) name20030 (
		_w24075_,
		_w24076_,
		_w24077_
	);
	LUT2 #(
		.INIT('h2)
	) name20031 (
		_w6106_,
		_w7340_,
		_w24078_
	);
	LUT2 #(
		.INIT('h4)
	) name20032 (
		_w6106_,
		_w6546_,
		_w24079_
	);
	LUT2 #(
		.INIT('h1)
	) name20033 (
		_w24078_,
		_w24079_,
		_w24080_
	);
	LUT2 #(
		.INIT('h4)
	) name20034 (
		_w6075_,
		_w24080_,
		_w24081_
	);
	LUT2 #(
		.INIT('h8)
	) name20035 (
		\core_dag_ilm1reg_I3_we_DO_reg[13]/NET0131 ,
		_w6075_,
		_w24082_
	);
	LUT2 #(
		.INIT('h1)
	) name20036 (
		_w24081_,
		_w24082_,
		_w24083_
	);
	LUT2 #(
		.INIT('h1)
	) name20037 (
		_w6106_,
		_w8962_,
		_w24084_
	);
	LUT2 #(
		.INIT('h8)
	) name20038 (
		_w6106_,
		_w9178_,
		_w24085_
	);
	LUT2 #(
		.INIT('h1)
	) name20039 (
		_w24084_,
		_w24085_,
		_w24086_
	);
	LUT2 #(
		.INIT('h1)
	) name20040 (
		_w6075_,
		_w24086_,
		_w24087_
	);
	LUT2 #(
		.INIT('h1)
	) name20041 (
		_w8869_,
		_w24087_,
		_w24088_
	);
	LUT2 #(
		.INIT('h1)
	) name20042 (
		_w6106_,
		_w8246_,
		_w24089_
	);
	LUT2 #(
		.INIT('h8)
	) name20043 (
		_w6106_,
		_w8460_,
		_w24090_
	);
	LUT2 #(
		.INIT('h1)
	) name20044 (
		_w24089_,
		_w24090_,
		_w24091_
	);
	LUT2 #(
		.INIT('h1)
	) name20045 (
		_w6075_,
		_w24091_,
		_w24092_
	);
	LUT2 #(
		.INIT('h1)
	) name20046 (
		_w8738_,
		_w24092_,
		_w24093_
	);
	LUT2 #(
		.INIT('h4)
	) name20047 (
		_w6075_,
		_w23763_,
		_w24094_
	);
	LUT2 #(
		.INIT('h1)
	) name20048 (
		_w8137_,
		_w24094_,
		_w24095_
	);
	LUT2 #(
		.INIT('h1)
	) name20049 (
		_w6106_,
		_w9752_,
		_w24096_
	);
	LUT2 #(
		.INIT('h8)
	) name20050 (
		_w6106_,
		_w10289_,
		_w24097_
	);
	LUT2 #(
		.INIT('h1)
	) name20051 (
		_w24096_,
		_w24097_,
		_w24098_
	);
	LUT2 #(
		.INIT('h1)
	) name20052 (
		_w6084_,
		_w24098_,
		_w24099_
	);
	LUT2 #(
		.INIT('h8)
	) name20053 (
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w6084_,
		_w24100_
	);
	LUT2 #(
		.INIT('h1)
	) name20054 (
		_w24099_,
		_w24100_,
		_w24101_
	);
	LUT2 #(
		.INIT('h4)
	) name20055 (
		_w6084_,
		_w24062_,
		_w24102_
	);
	LUT2 #(
		.INIT('h1)
	) name20056 (
		_w10398_,
		_w24102_,
		_w24103_
	);
	LUT2 #(
		.INIT('h1)
	) name20057 (
		_w6106_,
		_w10954_,
		_w24104_
	);
	LUT2 #(
		.INIT('h8)
	) name20058 (
		_w6106_,
		_w11265_,
		_w24105_
	);
	LUT2 #(
		.INIT('h1)
	) name20059 (
		_w24104_,
		_w24105_,
		_w24106_
	);
	LUT2 #(
		.INIT('h1)
	) name20060 (
		_w6084_,
		_w24106_,
		_w24107_
	);
	LUT2 #(
		.INIT('h1)
	) name20061 (
		_w11008_,
		_w24107_,
		_w24108_
	);
	LUT2 #(
		.INIT('h1)
	) name20062 (
		_w6106_,
		_w11280_,
		_w24109_
	);
	LUT2 #(
		.INIT('h8)
	) name20063 (
		_w6106_,
		_w11525_,
		_w24110_
	);
	LUT2 #(
		.INIT('h1)
	) name20064 (
		_w24109_,
		_w24110_,
		_w24111_
	);
	LUT2 #(
		.INIT('h1)
	) name20065 (
		_w6084_,
		_w24111_,
		_w24112_
	);
	LUT2 #(
		.INIT('h1)
	) name20066 (
		_w10979_,
		_w24112_,
		_w24113_
	);
	LUT2 #(
		.INIT('h4)
	) name20067 (
		_w6084_,
		_w24068_,
		_w24114_
	);
	LUT2 #(
		.INIT('h1)
	) name20068 (
		_w10371_,
		_w24114_,
		_w24115_
	);
	LUT2 #(
		.INIT('h1)
	) name20069 (
		_w6106_,
		_w10302_,
		_w24116_
	);
	LUT2 #(
		.INIT('h8)
	) name20070 (
		_w6106_,
		_w10069_,
		_w24117_
	);
	LUT2 #(
		.INIT('h1)
	) name20071 (
		_w24116_,
		_w24117_,
		_w24118_
	);
	LUT2 #(
		.INIT('h1)
	) name20072 (
		_w6084_,
		_w24118_,
		_w24119_
	);
	LUT2 #(
		.INIT('h8)
	) name20073 (
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w6084_,
		_w24120_
	);
	LUT2 #(
		.INIT('h1)
	) name20074 (
		_w24119_,
		_w24120_,
		_w24121_
	);
	LUT2 #(
		.INIT('h1)
	) name20075 (
		_w6106_,
		_w8794_,
		_w24122_
	);
	LUT2 #(
		.INIT('h8)
	) name20076 (
		_w6106_,
		_w8715_,
		_w24123_
	);
	LUT2 #(
		.INIT('h1)
	) name20077 (
		_w24122_,
		_w24123_,
		_w24124_
	);
	LUT2 #(
		.INIT('h1)
	) name20078 (
		_w6084_,
		_w24124_,
		_w24125_
	);
	LUT2 #(
		.INIT('h1)
	) name20079 (
		_w8766_,
		_w24125_,
		_w24126_
	);
	LUT2 #(
		.INIT('h1)
	) name20080 (
		_w6084_,
		_w24074_,
		_w24127_
	);
	LUT2 #(
		.INIT('h4)
	) name20081 (
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w6084_,
		_w24128_
	);
	LUT2 #(
		.INIT('h1)
	) name20082 (
		_w24127_,
		_w24128_,
		_w24129_
	);
	LUT2 #(
		.INIT('h4)
	) name20083 (
		_w6084_,
		_w24080_,
		_w24130_
	);
	LUT2 #(
		.INIT('h8)
	) name20084 (
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w6084_,
		_w24131_
	);
	LUT2 #(
		.INIT('h1)
	) name20085 (
		_w24130_,
		_w24131_,
		_w24132_
	);
	LUT2 #(
		.INIT('h1)
	) name20086 (
		_w6084_,
		_w24086_,
		_w24133_
	);
	LUT2 #(
		.INIT('h8)
	) name20087 (
		\core_dag_ilm1reg_I2_we_DO_reg[12]/NET0131 ,
		_w6084_,
		_w24134_
	);
	LUT2 #(
		.INIT('h1)
	) name20088 (
		_w24133_,
		_w24134_,
		_w24135_
	);
	LUT2 #(
		.INIT('h1)
	) name20089 (
		_w6084_,
		_w24091_,
		_w24136_
	);
	LUT2 #(
		.INIT('h1)
	) name20090 (
		_w8734_,
		_w24136_,
		_w24137_
	);
	LUT2 #(
		.INIT('h2)
	) name20091 (
		_w7340_,
		_w23865_,
		_w24138_
	);
	LUT2 #(
		.INIT('h8)
	) name20092 (
		\sport1_txctl_TX_reg[13]/P0001 ,
		_w23865_,
		_w24139_
	);
	LUT2 #(
		.INIT('h1)
	) name20093 (
		_w24138_,
		_w24139_,
		_w24140_
	);
	LUT2 #(
		.INIT('h1)
	) name20094 (
		_w6106_,
		_w7622_,
		_w24141_
	);
	LUT2 #(
		.INIT('h8)
	) name20095 (
		_w6106_,
		_w7607_,
		_w24142_
	);
	LUT2 #(
		.INIT('h1)
	) name20096 (
		_w24141_,
		_w24142_,
		_w24143_
	);
	LUT2 #(
		.INIT('h1)
	) name20097 (
		_w6084_,
		_w24143_,
		_w24144_
	);
	LUT2 #(
		.INIT('h8)
	) name20098 (
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w6084_,
		_w24145_
	);
	LUT2 #(
		.INIT('h1)
	) name20099 (
		_w24144_,
		_w24145_,
		_w24146_
	);
	LUT2 #(
		.INIT('h4)
	) name20100 (
		_w6067_,
		_w24062_,
		_w24147_
	);
	LUT2 #(
		.INIT('h1)
	) name20101 (
		_w10402_,
		_w24147_,
		_w24148_
	);
	LUT2 #(
		.INIT('h8)
	) name20102 (
		\core_dag_ilm1reg_I1_we_DO_reg[5]/NET0131 ,
		_w6067_,
		_w24149_
	);
	LUT2 #(
		.INIT('h4)
	) name20103 (
		_w6067_,
		_w24068_,
		_w24150_
	);
	LUT2 #(
		.INIT('h1)
	) name20104 (
		_w24149_,
		_w24150_,
		_w24151_
	);
	LUT2 #(
		.INIT('h4)
	) name20105 (
		_w6067_,
		_w24074_,
		_w24152_
	);
	LUT2 #(
		.INIT('h1)
	) name20106 (
		_w8891_,
		_w24152_,
		_w24153_
	);
	LUT2 #(
		.INIT('h8)
	) name20107 (
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w6067_,
		_w24154_
	);
	LUT2 #(
		.INIT('h4)
	) name20108 (
		_w6067_,
		_w24080_,
		_w24155_
	);
	LUT2 #(
		.INIT('h1)
	) name20109 (
		_w24154_,
		_w24155_,
		_w24156_
	);
	LUT2 #(
		.INIT('h4)
	) name20110 (
		_w6067_,
		_w24086_,
		_w24157_
	);
	LUT2 #(
		.INIT('h4)
	) name20111 (
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w6067_,
		_w24158_
	);
	LUT2 #(
		.INIT('h1)
	) name20112 (
		_w24157_,
		_w24158_,
		_w24159_
	);
	LUT2 #(
		.INIT('h1)
	) name20113 (
		_w6067_,
		_w24091_,
		_w24160_
	);
	LUT2 #(
		.INIT('h1)
	) name20114 (
		_w8736_,
		_w24160_,
		_w24161_
	);
	LUT2 #(
		.INIT('h4)
	) name20115 (
		_w6067_,
		_w23763_,
		_w24162_
	);
	LUT2 #(
		.INIT('h1)
	) name20116 (
		_w8135_,
		_w24162_,
		_w24163_
	);
	LUT2 #(
		.INIT('h1)
	) name20117 (
		_w6058_,
		_w24098_,
		_w24164_
	);
	LUT2 #(
		.INIT('h1)
	) name20118 (
		_w9718_,
		_w24164_,
		_w24165_
	);
	LUT2 #(
		.INIT('h8)
	) name20119 (
		\core_dag_ilm1reg_I0_we_DO_reg[8]/NET0131 ,
		_w6058_,
		_w24166_
	);
	LUT2 #(
		.INIT('h4)
	) name20120 (
		_w6058_,
		_w24062_,
		_w24167_
	);
	LUT2 #(
		.INIT('h1)
	) name20121 (
		_w24166_,
		_w24167_,
		_w24168_
	);
	LUT2 #(
		.INIT('h1)
	) name20122 (
		_w6058_,
		_w24106_,
		_w24169_
	);
	LUT2 #(
		.INIT('h8)
	) name20123 (
		\core_dag_ilm1reg_I0_we_DO_reg[7]/NET0131 ,
		_w6058_,
		_w24170_
	);
	LUT2 #(
		.INIT('h1)
	) name20124 (
		_w24169_,
		_w24170_,
		_w24171_
	);
	LUT2 #(
		.INIT('h1)
	) name20125 (
		_w6058_,
		_w24111_,
		_w24172_
	);
	LUT2 #(
		.INIT('h8)
	) name20126 (
		\core_dag_ilm1reg_I0_we_DO_reg[6]/NET0131 ,
		_w6058_,
		_w24173_
	);
	LUT2 #(
		.INIT('h1)
	) name20127 (
		_w24172_,
		_w24173_,
		_w24174_
	);
	LUT2 #(
		.INIT('h4)
	) name20128 (
		_w6058_,
		_w24068_,
		_w24175_
	);
	LUT2 #(
		.INIT('h1)
	) name20129 (
		_w10369_,
		_w24175_,
		_w24176_
	);
	LUT2 #(
		.INIT('h1)
	) name20130 (
		_w6058_,
		_w24118_,
		_w24177_
	);
	LUT2 #(
		.INIT('h1)
	) name20131 (
		_w9771_,
		_w24177_,
		_w24178_
	);
	LUT2 #(
		.INIT('h4)
	) name20132 (
		_w6058_,
		_w23886_,
		_w24179_
	);
	LUT2 #(
		.INIT('h1)
	) name20133 (
		_w8186_,
		_w24179_,
		_w24180_
	);
	LUT2 #(
		.INIT('h1)
	) name20134 (
		_w6058_,
		_w24124_,
		_w24181_
	);
	LUT2 #(
		.INIT('h8)
	) name20135 (
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w6058_,
		_w24182_
	);
	LUT2 #(
		.INIT('h1)
	) name20136 (
		_w24181_,
		_w24182_,
		_w24183_
	);
	LUT2 #(
		.INIT('h4)
	) name20137 (
		_w6058_,
		_w24074_,
		_w24184_
	);
	LUT2 #(
		.INIT('h1)
	) name20138 (
		_w8888_,
		_w24184_,
		_w24185_
	);
	LUT2 #(
		.INIT('h4)
	) name20139 (
		_w6058_,
		_w24080_,
		_w24186_
	);
	LUT2 #(
		.INIT('h1)
	) name20140 (
		_w6136_,
		_w24186_,
		_w24187_
	);
	LUT2 #(
		.INIT('h1)
	) name20141 (
		_w6058_,
		_w24086_,
		_w24188_
	);
	LUT2 #(
		.INIT('h1)
	) name20142 (
		_w8859_,
		_w24188_,
		_w24189_
	);
	LUT2 #(
		.INIT('h8)
	) name20143 (
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w6058_,
		_w24190_
	);
	LUT2 #(
		.INIT('h1)
	) name20144 (
		_w6058_,
		_w24091_,
		_w24191_
	);
	LUT2 #(
		.INIT('h1)
	) name20145 (
		_w24190_,
		_w24191_,
		_w24192_
	);
	LUT2 #(
		.INIT('h8)
	) name20146 (
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w6058_,
		_w24193_
	);
	LUT2 #(
		.INIT('h4)
	) name20147 (
		_w6058_,
		_w23763_,
		_w24194_
	);
	LUT2 #(
		.INIT('h1)
	) name20148 (
		_w24193_,
		_w24194_,
		_w24195_
	);
	LUT2 #(
		.INIT('h1)
	) name20149 (
		_w6058_,
		_w24143_,
		_w24196_
	);
	LUT2 #(
		.INIT('h1)
	) name20150 (
		_w6936_,
		_w24196_,
		_w24197_
	);
	LUT2 #(
		.INIT('h4)
	) name20151 (
		_w22114_,
		_w23766_,
		_w24198_
	);
	LUT2 #(
		.INIT('h1)
	) name20152 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[10]/P0001 ,
		_w23766_,
		_w24199_
	);
	LUT2 #(
		.INIT('h1)
	) name20153 (
		_w24198_,
		_w24199_,
		_w24200_
	);
	LUT2 #(
		.INIT('h4)
	) name20154 (
		_w17836_,
		_w23754_,
		_w24201_
	);
	LUT2 #(
		.INIT('h1)
	) name20155 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[13]/P0001 ,
		_w23754_,
		_w24202_
	);
	LUT2 #(
		.INIT('h1)
	) name20156 (
		_w24201_,
		_w24202_,
		_w24203_
	);
	LUT2 #(
		.INIT('h4)
	) name20157 (
		_w19848_,
		_w23754_,
		_w24204_
	);
	LUT2 #(
		.INIT('h1)
	) name20158 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[10]/P0001 ,
		_w23754_,
		_w24205_
	);
	LUT2 #(
		.INIT('h1)
	) name20159 (
		_w24204_,
		_w24205_,
		_w24206_
	);
	LUT2 #(
		.INIT('h2)
	) name20160 (
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w23958_,
		_w24207_
	);
	LUT2 #(
		.INIT('h4)
	) name20161 (
		_w6000_,
		_w20644_,
		_w24208_
	);
	LUT2 #(
		.INIT('h1)
	) name20162 (
		_w24207_,
		_w24208_,
		_w24209_
	);
	LUT2 #(
		.INIT('h2)
	) name20163 (
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w23958_,
		_w24210_
	);
	LUT2 #(
		.INIT('h4)
	) name20164 (
		_w6000_,
		_w13262_,
		_w24211_
	);
	LUT2 #(
		.INIT('h1)
	) name20165 (
		_w24210_,
		_w24211_,
		_w24212_
	);
	LUT2 #(
		.INIT('h2)
	) name20166 (
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w23958_,
		_w24213_
	);
	LUT2 #(
		.INIT('h1)
	) name20167 (
		_w6000_,
		_w20663_,
		_w24214_
	);
	LUT2 #(
		.INIT('h1)
	) name20168 (
		_w24213_,
		_w24214_,
		_w24215_
	);
	LUT2 #(
		.INIT('h2)
	) name20169 (
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w23958_,
		_w24216_
	);
	LUT2 #(
		.INIT('h1)
	) name20170 (
		_w6000_,
		_w20674_,
		_w24217_
	);
	LUT2 #(
		.INIT('h1)
	) name20171 (
		_w24216_,
		_w24217_,
		_w24218_
	);
	LUT2 #(
		.INIT('h2)
	) name20172 (
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w23958_,
		_w24219_
	);
	LUT2 #(
		.INIT('h1)
	) name20173 (
		_w6000_,
		_w20729_,
		_w24220_
	);
	LUT2 #(
		.INIT('h1)
	) name20174 (
		_w24219_,
		_w24220_,
		_w24221_
	);
	LUT2 #(
		.INIT('h4)
	) name20175 (
		_w6008_,
		_w20644_,
		_w24222_
	);
	LUT2 #(
		.INIT('h8)
	) name20176 (
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w6008_,
		_w24223_
	);
	LUT2 #(
		.INIT('h1)
	) name20177 (
		_w24222_,
		_w24223_,
		_w24224_
	);
	LUT2 #(
		.INIT('h4)
	) name20178 (
		_w6008_,
		_w13262_,
		_w24225_
	);
	LUT2 #(
		.INIT('h8)
	) name20179 (
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w6008_,
		_w24226_
	);
	LUT2 #(
		.INIT('h1)
	) name20180 (
		_w24225_,
		_w24226_,
		_w24227_
	);
	LUT2 #(
		.INIT('h1)
	) name20181 (
		_w6008_,
		_w20663_,
		_w24228_
	);
	LUT2 #(
		.INIT('h8)
	) name20182 (
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w6008_,
		_w24229_
	);
	LUT2 #(
		.INIT('h1)
	) name20183 (
		_w24228_,
		_w24229_,
		_w24230_
	);
	LUT2 #(
		.INIT('h1)
	) name20184 (
		_w6008_,
		_w20674_,
		_w24231_
	);
	LUT2 #(
		.INIT('h8)
	) name20185 (
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w6008_,
		_w24232_
	);
	LUT2 #(
		.INIT('h1)
	) name20186 (
		_w24231_,
		_w24232_,
		_w24233_
	);
	LUT2 #(
		.INIT('h1)
	) name20187 (
		_w6008_,
		_w20729_,
		_w24234_
	);
	LUT2 #(
		.INIT('h8)
	) name20188 (
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w6008_,
		_w24235_
	);
	LUT2 #(
		.INIT('h1)
	) name20189 (
		_w24234_,
		_w24235_,
		_w24236_
	);
	LUT2 #(
		.INIT('h2)
	) name20190 (
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		_w24004_,
		_w24237_
	);
	LUT2 #(
		.INIT('h4)
	) name20191 (
		_w6015_,
		_w20644_,
		_w24238_
	);
	LUT2 #(
		.INIT('h1)
	) name20192 (
		_w24237_,
		_w24238_,
		_w24239_
	);
	LUT2 #(
		.INIT('h2)
	) name20193 (
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		_w24004_,
		_w24240_
	);
	LUT2 #(
		.INIT('h4)
	) name20194 (
		_w6015_,
		_w13262_,
		_w24241_
	);
	LUT2 #(
		.INIT('h1)
	) name20195 (
		_w24240_,
		_w24241_,
		_w24242_
	);
	LUT2 #(
		.INIT('h2)
	) name20196 (
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		_w24004_,
		_w24243_
	);
	LUT2 #(
		.INIT('h1)
	) name20197 (
		_w6015_,
		_w20663_,
		_w24244_
	);
	LUT2 #(
		.INIT('h1)
	) name20198 (
		_w24243_,
		_w24244_,
		_w24245_
	);
	LUT2 #(
		.INIT('h2)
	) name20199 (
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		_w24004_,
		_w24246_
	);
	LUT2 #(
		.INIT('h1)
	) name20200 (
		_w6015_,
		_w20674_,
		_w24247_
	);
	LUT2 #(
		.INIT('h1)
	) name20201 (
		_w24246_,
		_w24247_,
		_w24248_
	);
	LUT2 #(
		.INIT('h2)
	) name20202 (
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		_w24004_,
		_w24249_
	);
	LUT2 #(
		.INIT('h1)
	) name20203 (
		_w6015_,
		_w20729_,
		_w24250_
	);
	LUT2 #(
		.INIT('h1)
	) name20204 (
		_w24249_,
		_w24250_,
		_w24251_
	);
	LUT2 #(
		.INIT('h2)
	) name20205 (
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w24023_,
		_w24252_
	);
	LUT2 #(
		.INIT('h4)
	) name20206 (
		_w5964_,
		_w20644_,
		_w24253_
	);
	LUT2 #(
		.INIT('h1)
	) name20207 (
		_w24252_,
		_w24253_,
		_w24254_
	);
	LUT2 #(
		.INIT('h2)
	) name20208 (
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w24023_,
		_w24255_
	);
	LUT2 #(
		.INIT('h4)
	) name20209 (
		_w5964_,
		_w13262_,
		_w24256_
	);
	LUT2 #(
		.INIT('h1)
	) name20210 (
		_w24255_,
		_w24256_,
		_w24257_
	);
	LUT2 #(
		.INIT('h2)
	) name20211 (
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w24023_,
		_w24258_
	);
	LUT2 #(
		.INIT('h1)
	) name20212 (
		_w5964_,
		_w20663_,
		_w24259_
	);
	LUT2 #(
		.INIT('h1)
	) name20213 (
		_w24258_,
		_w24259_,
		_w24260_
	);
	LUT2 #(
		.INIT('h2)
	) name20214 (
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w24023_,
		_w24261_
	);
	LUT2 #(
		.INIT('h1)
	) name20215 (
		_w5964_,
		_w20674_,
		_w24262_
	);
	LUT2 #(
		.INIT('h1)
	) name20216 (
		_w24261_,
		_w24262_,
		_w24263_
	);
	LUT2 #(
		.INIT('h2)
	) name20217 (
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w24023_,
		_w24264_
	);
	LUT2 #(
		.INIT('h1)
	) name20218 (
		_w5964_,
		_w20729_,
		_w24265_
	);
	LUT2 #(
		.INIT('h1)
	) name20219 (
		_w24264_,
		_w24265_,
		_w24266_
	);
	LUT2 #(
		.INIT('h8)
	) name20220 (
		_w23027_,
		_w23407_,
		_w24267_
	);
	LUT2 #(
		.INIT('h4)
	) name20221 (
		\sice_ICYC_clr_reg/NET0131 ,
		\sice_SPC_reg[23]/P0001 ,
		_w24268_
	);
	LUT2 #(
		.INIT('h8)
	) name20222 (
		_w23032_,
		_w24268_,
		_w24269_
	);
	LUT2 #(
		.INIT('h8)
	) name20223 (
		_w24267_,
		_w24269_,
		_w24270_
	);
	LUT2 #(
		.INIT('h2)
	) name20224 (
		\core_c_psq_Iact_E_reg[9]/NET0131 ,
		_w19477_,
		_w24271_
	);
	LUT2 #(
		.INIT('h1)
	) name20225 (
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w24272_
	);
	LUT2 #(
		.INIT('h8)
	) name20226 (
		_w19481_,
		_w24272_,
		_w24273_
	);
	LUT2 #(
		.INIT('h8)
	) name20227 (
		_w19477_,
		_w24273_,
		_w24274_
	);
	LUT2 #(
		.INIT('h1)
	) name20228 (
		_w24271_,
		_w24274_,
		_w24275_
	);
	LUT2 #(
		.INIT('h4)
	) name20229 (
		_w22021_,
		_w23782_,
		_w24276_
	);
	LUT2 #(
		.INIT('h1)
	) name20230 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[6]/P0001 ,
		_w23782_,
		_w24277_
	);
	LUT2 #(
		.INIT('h1)
	) name20231 (
		_w24276_,
		_w24277_,
		_w24278_
	);
	LUT2 #(
		.INIT('h2)
	) name20232 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][3]/P0001 ,
		_w4851_,
		_w24279_
	);
	LUT2 #(
		.INIT('h8)
	) name20233 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4851_,
		_w24280_
	);
	LUT2 #(
		.INIT('h1)
	) name20234 (
		_w24279_,
		_w24280_,
		_w24281_
	);
	LUT2 #(
		.INIT('h2)
	) name20235 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][2]/P0001 ,
		_w4851_,
		_w24282_
	);
	LUT2 #(
		.INIT('h8)
	) name20236 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4851_,
		_w24283_
	);
	LUT2 #(
		.INIT('h1)
	) name20237 (
		_w24282_,
		_w24283_,
		_w24284_
	);
	LUT2 #(
		.INIT('h2)
	) name20238 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][1]/P0001 ,
		_w4851_,
		_w24285_
	);
	LUT2 #(
		.INIT('h8)
	) name20239 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4851_,
		_w24286_
	);
	LUT2 #(
		.INIT('h1)
	) name20240 (
		_w24285_,
		_w24286_,
		_w24287_
	);
	LUT2 #(
		.INIT('h2)
	) name20241 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[3][0]/P0001 ,
		_w4851_,
		_w24288_
	);
	LUT2 #(
		.INIT('h8)
	) name20242 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4851_,
		_w24289_
	);
	LUT2 #(
		.INIT('h1)
	) name20243 (
		_w24288_,
		_w24289_,
		_w24290_
	);
	LUT2 #(
		.INIT('h2)
	) name20244 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][3]/P0001 ,
		_w4847_,
		_w24291_
	);
	LUT2 #(
		.INIT('h8)
	) name20245 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4847_,
		_w24292_
	);
	LUT2 #(
		.INIT('h1)
	) name20246 (
		_w24291_,
		_w24292_,
		_w24293_
	);
	LUT2 #(
		.INIT('h2)
	) name20247 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][1]/P0001 ,
		_w4847_,
		_w24294_
	);
	LUT2 #(
		.INIT('h8)
	) name20248 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4847_,
		_w24295_
	);
	LUT2 #(
		.INIT('h1)
	) name20249 (
		_w24294_,
		_w24295_,
		_w24296_
	);
	LUT2 #(
		.INIT('h2)
	) name20250 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][2]/P0001 ,
		_w4845_,
		_w24297_
	);
	LUT2 #(
		.INIT('h8)
	) name20251 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4845_,
		_w24298_
	);
	LUT2 #(
		.INIT('h1)
	) name20252 (
		_w24297_,
		_w24298_,
		_w24299_
	);
	LUT2 #(
		.INIT('h2)
	) name20253 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][0]/P0001 ,
		_w4845_,
		_w24300_
	);
	LUT2 #(
		.INIT('h8)
	) name20254 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4845_,
		_w24301_
	);
	LUT2 #(
		.INIT('h1)
	) name20255 (
		_w24300_,
		_w24301_,
		_w24302_
	);
	LUT2 #(
		.INIT('h2)
	) name20256 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][3]/P0001 ,
		_w4849_,
		_w24303_
	);
	LUT2 #(
		.INIT('h8)
	) name20257 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4849_,
		_w24304_
	);
	LUT2 #(
		.INIT('h1)
	) name20258 (
		_w24303_,
		_w24304_,
		_w24305_
	);
	LUT2 #(
		.INIT('h2)
	) name20259 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][2]/P0001 ,
		_w4849_,
		_w24306_
	);
	LUT2 #(
		.INIT('h8)
	) name20260 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4849_,
		_w24307_
	);
	LUT2 #(
		.INIT('h1)
	) name20261 (
		_w24306_,
		_w24307_,
		_w24308_
	);
	LUT2 #(
		.INIT('h2)
	) name20262 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][1]/P0001 ,
		_w4849_,
		_w24309_
	);
	LUT2 #(
		.INIT('h8)
	) name20263 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4849_,
		_w24310_
	);
	LUT2 #(
		.INIT('h1)
	) name20264 (
		_w24309_,
		_w24310_,
		_w24311_
	);
	LUT2 #(
		.INIT('h2)
	) name20265 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][2]/P0001 ,
		_w4847_,
		_w24312_
	);
	LUT2 #(
		.INIT('h8)
	) name20266 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w4847_,
		_w24313_
	);
	LUT2 #(
		.INIT('h1)
	) name20267 (
		_w24312_,
		_w24313_,
		_w24314_
	);
	LUT2 #(
		.INIT('h2)
	) name20268 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001 ,
		_w13794_,
		_w24315_
	);
	LUT2 #(
		.INIT('h8)
	) name20269 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w13794_,
		_w24316_
	);
	LUT2 #(
		.INIT('h1)
	) name20270 (
		_w24315_,
		_w24316_,
		_w24317_
	);
	LUT2 #(
		.INIT('h2)
	) name20271 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001 ,
		_w13794_,
		_w24318_
	);
	LUT2 #(
		.INIT('h8)
	) name20272 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w13794_,
		_w24319_
	);
	LUT2 #(
		.INIT('h1)
	) name20273 (
		_w24318_,
		_w24319_,
		_w24320_
	);
	LUT2 #(
		.INIT('h2)
	) name20274 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001 ,
		_w13794_,
		_w24321_
	);
	LUT2 #(
		.INIT('h8)
	) name20275 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w13794_,
		_w24322_
	);
	LUT2 #(
		.INIT('h1)
	) name20276 (
		_w24321_,
		_w24322_,
		_w24323_
	);
	LUT2 #(
		.INIT('h2)
	) name20277 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001 ,
		_w13794_,
		_w24324_
	);
	LUT2 #(
		.INIT('h8)
	) name20278 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w13794_,
		_w24325_
	);
	LUT2 #(
		.INIT('h1)
	) name20279 (
		_w24324_,
		_w24325_,
		_w24326_
	);
	LUT2 #(
		.INIT('h2)
	) name20280 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001 ,
		_w13794_,
		_w24327_
	);
	LUT2 #(
		.INIT('h8)
	) name20281 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w13794_,
		_w24328_
	);
	LUT2 #(
		.INIT('h1)
	) name20282 (
		_w24327_,
		_w24328_,
		_w24329_
	);
	LUT2 #(
		.INIT('h2)
	) name20283 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001 ,
		_w13794_,
		_w24330_
	);
	LUT2 #(
		.INIT('h8)
	) name20284 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w13794_,
		_w24331_
	);
	LUT2 #(
		.INIT('h1)
	) name20285 (
		_w24330_,
		_w24331_,
		_w24332_
	);
	LUT2 #(
		.INIT('h2)
	) name20286 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001 ,
		_w13794_,
		_w24333_
	);
	LUT2 #(
		.INIT('h8)
	) name20287 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w13794_,
		_w24334_
	);
	LUT2 #(
		.INIT('h1)
	) name20288 (
		_w24333_,
		_w24334_,
		_w24335_
	);
	LUT2 #(
		.INIT('h2)
	) name20289 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001 ,
		_w13794_,
		_w24336_
	);
	LUT2 #(
		.INIT('h8)
	) name20290 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w13794_,
		_w24337_
	);
	LUT2 #(
		.INIT('h1)
	) name20291 (
		_w24336_,
		_w24337_,
		_w24338_
	);
	LUT2 #(
		.INIT('h2)
	) name20292 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001 ,
		_w13794_,
		_w24339_
	);
	LUT2 #(
		.INIT('h8)
	) name20293 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w13794_,
		_w24340_
	);
	LUT2 #(
		.INIT('h1)
	) name20294 (
		_w24339_,
		_w24340_,
		_w24341_
	);
	LUT2 #(
		.INIT('h2)
	) name20295 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001 ,
		_w13794_,
		_w24342_
	);
	LUT2 #(
		.INIT('h8)
	) name20296 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w13794_,
		_w24343_
	);
	LUT2 #(
		.INIT('h1)
	) name20297 (
		_w24342_,
		_w24343_,
		_w24344_
	);
	LUT2 #(
		.INIT('h2)
	) name20298 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001 ,
		_w13794_,
		_w24345_
	);
	LUT2 #(
		.INIT('h8)
	) name20299 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		_w13794_,
		_w24346_
	);
	LUT2 #(
		.INIT('h1)
	) name20300 (
		_w24345_,
		_w24346_,
		_w24347_
	);
	LUT2 #(
		.INIT('h2)
	) name20301 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001 ,
		_w13789_,
		_w24348_
	);
	LUT2 #(
		.INIT('h8)
	) name20302 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w13789_,
		_w24349_
	);
	LUT2 #(
		.INIT('h1)
	) name20303 (
		_w24348_,
		_w24349_,
		_w24350_
	);
	LUT2 #(
		.INIT('h2)
	) name20304 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001 ,
		_w13789_,
		_w24351_
	);
	LUT2 #(
		.INIT('h8)
	) name20305 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w13789_,
		_w24352_
	);
	LUT2 #(
		.INIT('h1)
	) name20306 (
		_w24351_,
		_w24352_,
		_w24353_
	);
	LUT2 #(
		.INIT('h2)
	) name20307 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001 ,
		_w13789_,
		_w24354_
	);
	LUT2 #(
		.INIT('h8)
	) name20308 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w13789_,
		_w24355_
	);
	LUT2 #(
		.INIT('h1)
	) name20309 (
		_w24354_,
		_w24355_,
		_w24356_
	);
	LUT2 #(
		.INIT('h2)
	) name20310 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001 ,
		_w13789_,
		_w24357_
	);
	LUT2 #(
		.INIT('h8)
	) name20311 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w13789_,
		_w24358_
	);
	LUT2 #(
		.INIT('h1)
	) name20312 (
		_w24357_,
		_w24358_,
		_w24359_
	);
	LUT2 #(
		.INIT('h2)
	) name20313 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001 ,
		_w13789_,
		_w24360_
	);
	LUT2 #(
		.INIT('h8)
	) name20314 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w13789_,
		_w24361_
	);
	LUT2 #(
		.INIT('h1)
	) name20315 (
		_w24360_,
		_w24361_,
		_w24362_
	);
	LUT2 #(
		.INIT('h2)
	) name20316 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001 ,
		_w13789_,
		_w24363_
	);
	LUT2 #(
		.INIT('h8)
	) name20317 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		_w13789_,
		_w24364_
	);
	LUT2 #(
		.INIT('h1)
	) name20318 (
		_w24363_,
		_w24364_,
		_w24365_
	);
	LUT2 #(
		.INIT('h2)
	) name20319 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001 ,
		_w13784_,
		_w24366_
	);
	LUT2 #(
		.INIT('h8)
	) name20320 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w13784_,
		_w24367_
	);
	LUT2 #(
		.INIT('h1)
	) name20321 (
		_w24366_,
		_w24367_,
		_w24368_
	);
	LUT2 #(
		.INIT('h2)
	) name20322 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001 ,
		_w13784_,
		_w24369_
	);
	LUT2 #(
		.INIT('h8)
	) name20323 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w13784_,
		_w24370_
	);
	LUT2 #(
		.INIT('h1)
	) name20324 (
		_w24369_,
		_w24370_,
		_w24371_
	);
	LUT2 #(
		.INIT('h2)
	) name20325 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001 ,
		_w13784_,
		_w24372_
	);
	LUT2 #(
		.INIT('h8)
	) name20326 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w13784_,
		_w24373_
	);
	LUT2 #(
		.INIT('h1)
	) name20327 (
		_w24372_,
		_w24373_,
		_w24374_
	);
	LUT2 #(
		.INIT('h2)
	) name20328 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001 ,
		_w13784_,
		_w24375_
	);
	LUT2 #(
		.INIT('h8)
	) name20329 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w13784_,
		_w24376_
	);
	LUT2 #(
		.INIT('h1)
	) name20330 (
		_w24375_,
		_w24376_,
		_w24377_
	);
	LUT2 #(
		.INIT('h2)
	) name20331 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001 ,
		_w13784_,
		_w24378_
	);
	LUT2 #(
		.INIT('h8)
	) name20332 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w13784_,
		_w24379_
	);
	LUT2 #(
		.INIT('h1)
	) name20333 (
		_w24378_,
		_w24379_,
		_w24380_
	);
	LUT2 #(
		.INIT('h2)
	) name20334 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001 ,
		_w13784_,
		_w24381_
	);
	LUT2 #(
		.INIT('h8)
	) name20335 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w13784_,
		_w24382_
	);
	LUT2 #(
		.INIT('h1)
	) name20336 (
		_w24381_,
		_w24382_,
		_w24383_
	);
	LUT2 #(
		.INIT('h2)
	) name20337 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001 ,
		_w13784_,
		_w24384_
	);
	LUT2 #(
		.INIT('h8)
	) name20338 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w13784_,
		_w24385_
	);
	LUT2 #(
		.INIT('h1)
	) name20339 (
		_w24384_,
		_w24385_,
		_w24386_
	);
	LUT2 #(
		.INIT('h2)
	) name20340 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001 ,
		_w13784_,
		_w24387_
	);
	LUT2 #(
		.INIT('h8)
	) name20341 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w13784_,
		_w24388_
	);
	LUT2 #(
		.INIT('h1)
	) name20342 (
		_w24387_,
		_w24388_,
		_w24389_
	);
	LUT2 #(
		.INIT('h2)
	) name20343 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001 ,
		_w13784_,
		_w24390_
	);
	LUT2 #(
		.INIT('h8)
	) name20344 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w13784_,
		_w24391_
	);
	LUT2 #(
		.INIT('h1)
	) name20345 (
		_w24390_,
		_w24391_,
		_w24392_
	);
	LUT2 #(
		.INIT('h2)
	) name20346 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001 ,
		_w13775_,
		_w24393_
	);
	LUT2 #(
		.INIT('h8)
	) name20347 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w13775_,
		_w24394_
	);
	LUT2 #(
		.INIT('h1)
	) name20348 (
		_w24393_,
		_w24394_,
		_w24395_
	);
	LUT2 #(
		.INIT('h4)
	) name20349 (
		_w18276_,
		_w23754_,
		_w24396_
	);
	LUT2 #(
		.INIT('h1)
	) name20350 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[6]/P0001 ,
		_w23754_,
		_w24397_
	);
	LUT2 #(
		.INIT('h1)
	) name20351 (
		_w24396_,
		_w24397_,
		_w24398_
	);
	LUT2 #(
		.INIT('h4)
	) name20352 (
		_w22048_,
		_w23814_,
		_w24399_
	);
	LUT2 #(
		.INIT('h1)
	) name20353 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[3]/P0001 ,
		_w23814_,
		_w24400_
	);
	LUT2 #(
		.INIT('h1)
	) name20354 (
		_w24399_,
		_w24400_,
		_w24401_
	);
	LUT2 #(
		.INIT('h8)
	) name20355 (
		\core_c_dec_MTPMOVL_E_reg/P0001 ,
		_w5951_,
		_w24402_
	);
	LUT2 #(
		.INIT('h8)
	) name20356 (
		_w7607_,
		_w8113_,
		_w24403_
	);
	LUT2 #(
		.INIT('h8)
	) name20357 (
		_w8715_,
		_w9435_,
		_w24404_
	);
	LUT2 #(
		.INIT('h8)
	) name20358 (
		_w24403_,
		_w24404_,
		_w24405_
	);
	LUT2 #(
		.INIT('h2)
	) name20359 (
		_w24402_,
		_w24405_,
		_w24406_
	);
	LUT2 #(
		.INIT('h1)
	) name20360 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w24406_,
		_w24407_
	);
	LUT2 #(
		.INIT('h4)
	) name20361 (
		_w8113_,
		_w24402_,
		_w24408_
	);
	LUT2 #(
		.INIT('h1)
	) name20362 (
		_w24407_,
		_w24408_,
		_w24409_
	);
	LUT2 #(
		.INIT('h1)
	) name20363 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		_w24406_,
		_w24410_
	);
	LUT2 #(
		.INIT('h4)
	) name20364 (
		_w8715_,
		_w24402_,
		_w24411_
	);
	LUT2 #(
		.INIT('h1)
	) name20365 (
		_w24410_,
		_w24411_,
		_w24412_
	);
	LUT2 #(
		.INIT('h4)
	) name20366 (
		_w9435_,
		_w24406_,
		_w24413_
	);
	LUT2 #(
		.INIT('h1)
	) name20367 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w24406_,
		_w24414_
	);
	LUT2 #(
		.INIT('h1)
	) name20368 (
		_w24413_,
		_w24414_,
		_w24415_
	);
	LUT2 #(
		.INIT('h4)
	) name20369 (
		_w7607_,
		_w24406_,
		_w24416_
	);
	LUT2 #(
		.INIT('h1)
	) name20370 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w24406_,
		_w24417_
	);
	LUT2 #(
		.INIT('h1)
	) name20371 (
		_w24416_,
		_w24417_,
		_w24418_
	);
	LUT2 #(
		.INIT('h8)
	) name20372 (
		_w10069_,
		_w10911_,
		_w24419_
	);
	LUT2 #(
		.INIT('h8)
	) name20373 (
		_w11265_,
		_w24419_,
		_w24420_
	);
	LUT2 #(
		.INIT('h8)
	) name20374 (
		_w11525_,
		_w24420_,
		_w24421_
	);
	LUT2 #(
		.INIT('h2)
	) name20375 (
		_w24402_,
		_w24421_,
		_w24422_
	);
	LUT2 #(
		.INIT('h1)
	) name20376 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w24422_,
		_w24423_
	);
	LUT2 #(
		.INIT('h4)
	) name20377 (
		_w11265_,
		_w24402_,
		_w24424_
	);
	LUT2 #(
		.INIT('h1)
	) name20378 (
		_w24423_,
		_w24424_,
		_w24425_
	);
	LUT2 #(
		.INIT('h4)
	) name20379 (
		_w11525_,
		_w24422_,
		_w24426_
	);
	LUT2 #(
		.INIT('h1)
	) name20380 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		_w24422_,
		_w24427_
	);
	LUT2 #(
		.INIT('h1)
	) name20381 (
		_w24426_,
		_w24427_,
		_w24428_
	);
	LUT2 #(
		.INIT('h1)
	) name20382 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		_w24422_,
		_w24429_
	);
	LUT2 #(
		.INIT('h4)
	) name20383 (
		_w10911_,
		_w24402_,
		_w24430_
	);
	LUT2 #(
		.INIT('h1)
	) name20384 (
		_w24429_,
		_w24430_,
		_w24431_
	);
	LUT2 #(
		.INIT('h4)
	) name20385 (
		_w19972_,
		_w23754_,
		_w24432_
	);
	LUT2 #(
		.INIT('h1)
	) name20386 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[7]/P0001 ,
		_w23754_,
		_w24433_
	);
	LUT2 #(
		.INIT('h1)
	) name20387 (
		_w24432_,
		_w24433_,
		_w24434_
	);
	LUT2 #(
		.INIT('h2)
	) name20388 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001 ,
		_w13784_,
		_w24435_
	);
	LUT2 #(
		.INIT('h8)
	) name20389 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w13784_,
		_w24436_
	);
	LUT2 #(
		.INIT('h1)
	) name20390 (
		_w24435_,
		_w24436_,
		_w24437_
	);
	LUT2 #(
		.INIT('h2)
	) name20391 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001 ,
		_w13775_,
		_w24438_
	);
	LUT2 #(
		.INIT('h8)
	) name20392 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w13775_,
		_w24439_
	);
	LUT2 #(
		.INIT('h1)
	) name20393 (
		_w24438_,
		_w24439_,
		_w24440_
	);
	LUT2 #(
		.INIT('h8)
	) name20394 (
		_w6117_,
		_w13576_,
		_w24441_
	);
	LUT2 #(
		.INIT('h1)
	) name20395 (
		_w6107_,
		_w24441_,
		_w24442_
	);
	LUT2 #(
		.INIT('h4)
	) name20396 (
		_w4117_,
		_w24442_,
		_w24443_
	);
	LUT2 #(
		.INIT('h4)
	) name20397 (
		\core_c_dec_imm16_E_reg/P0001 ,
		_w4117_,
		_w24444_
	);
	LUT2 #(
		.INIT('h1)
	) name20398 (
		_w24443_,
		_w24444_,
		_w24445_
	);
	LUT2 #(
		.INIT('h4)
	) name20399 (
		_w10069_,
		_w24422_,
		_w24446_
	);
	LUT2 #(
		.INIT('h1)
	) name20400 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		_w24422_,
		_w24447_
	);
	LUT2 #(
		.INIT('h1)
	) name20401 (
		_w24446_,
		_w24447_,
		_w24448_
	);
	LUT2 #(
		.INIT('h2)
	) name20402 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[2][0]/P0001 ,
		_w4847_,
		_w24449_
	);
	LUT2 #(
		.INIT('h8)
	) name20403 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4847_,
		_w24450_
	);
	LUT2 #(
		.INIT('h1)
	) name20404 (
		_w24449_,
		_w24450_,
		_w24451_
	);
	LUT2 #(
		.INIT('h2)
	) name20405 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001 ,
		_w13775_,
		_w24452_
	);
	LUT2 #(
		.INIT('h8)
	) name20406 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w13775_,
		_w24453_
	);
	LUT2 #(
		.INIT('h1)
	) name20407 (
		_w24452_,
		_w24453_,
		_w24454_
	);
	LUT2 #(
		.INIT('h2)
	) name20408 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[0][0]/P0001 ,
		_w4849_,
		_w24455_
	);
	LUT2 #(
		.INIT('h8)
	) name20409 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		_w4849_,
		_w24456_
	);
	LUT2 #(
		.INIT('h1)
	) name20410 (
		_w24455_,
		_w24456_,
		_w24457_
	);
	LUT2 #(
		.INIT('h4)
	) name20411 (
		_w22012_,
		_w23766_,
		_w24458_
	);
	LUT2 #(
		.INIT('h1)
	) name20412 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[7]/P0001 ,
		_w23766_,
		_w24459_
	);
	LUT2 #(
		.INIT('h1)
	) name20413 (
		_w24458_,
		_w24459_,
		_w24460_
	);
	LUT2 #(
		.INIT('h4)
	) name20414 (
		_w22021_,
		_w23766_,
		_w24461_
	);
	LUT2 #(
		.INIT('h1)
	) name20415 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[6]/P0001 ,
		_w23766_,
		_w24462_
	);
	LUT2 #(
		.INIT('h1)
	) name20416 (
		_w24461_,
		_w24462_,
		_w24463_
	);
	LUT2 #(
		.INIT('h4)
	) name20417 (
		_w22030_,
		_w23766_,
		_w24464_
	);
	LUT2 #(
		.INIT('h1)
	) name20418 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[5]/P0001 ,
		_w23766_,
		_w24465_
	);
	LUT2 #(
		.INIT('h1)
	) name20419 (
		_w24464_,
		_w24465_,
		_w24466_
	);
	LUT2 #(
		.INIT('h4)
	) name20420 (
		_w22039_,
		_w23766_,
		_w24467_
	);
	LUT2 #(
		.INIT('h1)
	) name20421 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[4]/P0001 ,
		_w23766_,
		_w24468_
	);
	LUT2 #(
		.INIT('h1)
	) name20422 (
		_w24467_,
		_w24468_,
		_w24469_
	);
	LUT2 #(
		.INIT('h4)
	) name20423 (
		_w22048_,
		_w23766_,
		_w24470_
	);
	LUT2 #(
		.INIT('h1)
	) name20424 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[3]/P0001 ,
		_w23766_,
		_w24471_
	);
	LUT2 #(
		.INIT('h1)
	) name20425 (
		_w24470_,
		_w24471_,
		_w24472_
	);
	LUT2 #(
		.INIT('h4)
	) name20426 (
		_w22057_,
		_w23766_,
		_w24473_
	);
	LUT2 #(
		.INIT('h1)
	) name20427 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[2]/P0001 ,
		_w23766_,
		_w24474_
	);
	LUT2 #(
		.INIT('h1)
	) name20428 (
		_w24473_,
		_w24474_,
		_w24475_
	);
	LUT2 #(
		.INIT('h4)
	) name20429 (
		_w22151_,
		_w23766_,
		_w24476_
	);
	LUT2 #(
		.INIT('h1)
	) name20430 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[1]/P0001 ,
		_w23766_,
		_w24477_
	);
	LUT2 #(
		.INIT('h1)
	) name20431 (
		_w24476_,
		_w24477_,
		_w24478_
	);
	LUT2 #(
		.INIT('h4)
	) name20432 (
		_w22066_,
		_w23766_,
		_w24479_
	);
	LUT2 #(
		.INIT('h1)
	) name20433 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[15]/P0001 ,
		_w23766_,
		_w24480_
	);
	LUT2 #(
		.INIT('h1)
	) name20434 (
		_w24479_,
		_w24480_,
		_w24481_
	);
	LUT2 #(
		.INIT('h4)
	) name20435 (
		_w22075_,
		_w23766_,
		_w24482_
	);
	LUT2 #(
		.INIT('h1)
	) name20436 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[14]/P0001 ,
		_w23766_,
		_w24483_
	);
	LUT2 #(
		.INIT('h1)
	) name20437 (
		_w24482_,
		_w24483_,
		_w24484_
	);
	LUT2 #(
		.INIT('h4)
	) name20438 (
		_w22012_,
		_w23782_,
		_w24485_
	);
	LUT2 #(
		.INIT('h1)
	) name20439 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[7]/P0001 ,
		_w23782_,
		_w24486_
	);
	LUT2 #(
		.INIT('h1)
	) name20440 (
		_w24485_,
		_w24486_,
		_w24487_
	);
	LUT2 #(
		.INIT('h4)
	) name20441 (
		_w22039_,
		_w23782_,
		_w24488_
	);
	LUT2 #(
		.INIT('h1)
	) name20442 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[4]/P0001 ,
		_w23782_,
		_w24489_
	);
	LUT2 #(
		.INIT('h1)
	) name20443 (
		_w24488_,
		_w24489_,
		_w24490_
	);
	LUT2 #(
		.INIT('h4)
	) name20444 (
		_w22048_,
		_w23782_,
		_w24491_
	);
	LUT2 #(
		.INIT('h1)
	) name20445 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[3]/P0001 ,
		_w23782_,
		_w24492_
	);
	LUT2 #(
		.INIT('h1)
	) name20446 (
		_w24491_,
		_w24492_,
		_w24493_
	);
	LUT2 #(
		.INIT('h4)
	) name20447 (
		_w22151_,
		_w23782_,
		_w24494_
	);
	LUT2 #(
		.INIT('h1)
	) name20448 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[1]/P0001 ,
		_w23782_,
		_w24495_
	);
	LUT2 #(
		.INIT('h1)
	) name20449 (
		_w24494_,
		_w24495_,
		_w24496_
	);
	LUT2 #(
		.INIT('h4)
	) name20450 (
		_w22066_,
		_w23782_,
		_w24497_
	);
	LUT2 #(
		.INIT('h1)
	) name20451 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[15]/P0001 ,
		_w23782_,
		_w24498_
	);
	LUT2 #(
		.INIT('h1)
	) name20452 (
		_w24497_,
		_w24498_,
		_w24499_
	);
	LUT2 #(
		.INIT('h4)
	) name20453 (
		_w22075_,
		_w23782_,
		_w24500_
	);
	LUT2 #(
		.INIT('h1)
	) name20454 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[14]/P0001 ,
		_w23782_,
		_w24501_
	);
	LUT2 #(
		.INIT('h1)
	) name20455 (
		_w24500_,
		_w24501_,
		_w24502_
	);
	LUT2 #(
		.INIT('h4)
	) name20456 (
		_w22039_,
		_w23798_,
		_w24503_
	);
	LUT2 #(
		.INIT('h1)
	) name20457 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[4]/P0001 ,
		_w23798_,
		_w24504_
	);
	LUT2 #(
		.INIT('h1)
	) name20458 (
		_w24503_,
		_w24504_,
		_w24505_
	);
	LUT2 #(
		.INIT('h4)
	) name20459 (
		_w22021_,
		_w23798_,
		_w24506_
	);
	LUT2 #(
		.INIT('h1)
	) name20460 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[6]/P0001 ,
		_w23798_,
		_w24507_
	);
	LUT2 #(
		.INIT('h1)
	) name20461 (
		_w24506_,
		_w24507_,
		_w24508_
	);
	LUT2 #(
		.INIT('h4)
	) name20462 (
		_w22048_,
		_w23798_,
		_w24509_
	);
	LUT2 #(
		.INIT('h1)
	) name20463 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[3]/P0001 ,
		_w23798_,
		_w24510_
	);
	LUT2 #(
		.INIT('h1)
	) name20464 (
		_w24509_,
		_w24510_,
		_w24511_
	);
	LUT2 #(
		.INIT('h4)
	) name20465 (
		_w22151_,
		_w23798_,
		_w24512_
	);
	LUT2 #(
		.INIT('h1)
	) name20466 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[1]/P0001 ,
		_w23798_,
		_w24513_
	);
	LUT2 #(
		.INIT('h1)
	) name20467 (
		_w24512_,
		_w24513_,
		_w24514_
	);
	LUT2 #(
		.INIT('h4)
	) name20468 (
		_w7607_,
		_w21991_,
		_w24515_
	);
	LUT2 #(
		.INIT('h1)
	) name20469 (
		_w12520_,
		_w21991_,
		_w24516_
	);
	LUT2 #(
		.INIT('h1)
	) name20470 (
		_w24515_,
		_w24516_,
		_w24517_
	);
	LUT2 #(
		.INIT('h2)
	) name20471 (
		_w23798_,
		_w24517_,
		_w24518_
	);
	LUT2 #(
		.INIT('h1)
	) name20472 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[0]/P0001 ,
		_w23798_,
		_w24519_
	);
	LUT2 #(
		.INIT('h1)
	) name20473 (
		_w24518_,
		_w24519_,
		_w24520_
	);
	LUT2 #(
		.INIT('h4)
	) name20474 (
		_w22012_,
		_w23814_,
		_w24521_
	);
	LUT2 #(
		.INIT('h1)
	) name20475 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[7]/P0001 ,
		_w23814_,
		_w24522_
	);
	LUT2 #(
		.INIT('h1)
	) name20476 (
		_w24521_,
		_w24522_,
		_w24523_
	);
	LUT2 #(
		.INIT('h4)
	) name20477 (
		_w22030_,
		_w23814_,
		_w24524_
	);
	LUT2 #(
		.INIT('h1)
	) name20478 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[5]/P0001 ,
		_w23814_,
		_w24525_
	);
	LUT2 #(
		.INIT('h1)
	) name20479 (
		_w24524_,
		_w24525_,
		_w24526_
	);
	LUT2 #(
		.INIT('h4)
	) name20480 (
		_w22039_,
		_w23814_,
		_w24527_
	);
	LUT2 #(
		.INIT('h1)
	) name20481 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[4]/P0001 ,
		_w23814_,
		_w24528_
	);
	LUT2 #(
		.INIT('h1)
	) name20482 (
		_w24527_,
		_w24528_,
		_w24529_
	);
	LUT2 #(
		.INIT('h4)
	) name20483 (
		_w22057_,
		_w23814_,
		_w24530_
	);
	LUT2 #(
		.INIT('h1)
	) name20484 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[2]/P0001 ,
		_w23814_,
		_w24531_
	);
	LUT2 #(
		.INIT('h1)
	) name20485 (
		_w24530_,
		_w24531_,
		_w24532_
	);
	LUT2 #(
		.INIT('h2)
	) name20486 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][3]/P0001 ,
		_w4845_,
		_w24533_
	);
	LUT2 #(
		.INIT('h8)
	) name20487 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		_w4845_,
		_w24534_
	);
	LUT2 #(
		.INIT('h1)
	) name20488 (
		_w24533_,
		_w24534_,
		_w24535_
	);
	LUT2 #(
		.INIT('h4)
	) name20489 (
		_w22075_,
		_w23814_,
		_w24536_
	);
	LUT2 #(
		.INIT('h1)
	) name20490 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[14]/P0001 ,
		_w23814_,
		_w24537_
	);
	LUT2 #(
		.INIT('h1)
	) name20491 (
		_w24536_,
		_w24537_,
		_w24538_
	);
	LUT2 #(
		.INIT('h2)
	) name20492 (
		_w23814_,
		_w24517_,
		_w24539_
	);
	LUT2 #(
		.INIT('h1)
	) name20493 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[0]/P0001 ,
		_w23814_,
		_w24540_
	);
	LUT2 #(
		.INIT('h1)
	) name20494 (
		_w24539_,
		_w24540_,
		_w24541_
	);
	LUT2 #(
		.INIT('h2)
	) name20495 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001 ,
		_w13784_,
		_w24542_
	);
	LUT2 #(
		.INIT('h8)
	) name20496 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w13784_,
		_w24543_
	);
	LUT2 #(
		.INIT('h1)
	) name20497 (
		_w24542_,
		_w24543_,
		_w24544_
	);
	LUT2 #(
		.INIT('h4)
	) name20498 (
		_w11265_,
		_w23827_,
		_w24545_
	);
	LUT2 #(
		.INIT('h1)
	) name20499 (
		\bdma_BOVL_reg[7]/NET0131 ,
		_w23827_,
		_w24546_
	);
	LUT2 #(
		.INIT('h1)
	) name20500 (
		_w24545_,
		_w24546_,
		_w24547_
	);
	LUT2 #(
		.INIT('h4)
	) name20501 (
		_w11525_,
		_w23827_,
		_w24548_
	);
	LUT2 #(
		.INIT('h1)
	) name20502 (
		\bdma_BOVL_reg[6]/NET0131 ,
		_w23827_,
		_w24549_
	);
	LUT2 #(
		.INIT('h1)
	) name20503 (
		_w24548_,
		_w24549_,
		_w24550_
	);
	LUT2 #(
		.INIT('h4)
	) name20504 (
		_w10911_,
		_w23827_,
		_w24551_
	);
	LUT2 #(
		.INIT('h1)
	) name20505 (
		\bdma_BOVL_reg[5]/NET0131 ,
		_w23827_,
		_w24552_
	);
	LUT2 #(
		.INIT('h1)
	) name20506 (
		_w24551_,
		_w24552_,
		_w24553_
	);
	LUT2 #(
		.INIT('h4)
	) name20507 (
		_w10069_,
		_w23827_,
		_w24554_
	);
	LUT2 #(
		.INIT('h1)
	) name20508 (
		\bdma_BOVL_reg[4]/NET0131 ,
		_w23827_,
		_w24555_
	);
	LUT2 #(
		.INIT('h1)
	) name20509 (
		_w24554_,
		_w24555_,
		_w24556_
	);
	LUT2 #(
		.INIT('h4)
	) name20510 (
		_w8113_,
		_w23827_,
		_w24557_
	);
	LUT2 #(
		.INIT('h1)
	) name20511 (
		\bdma_BOVL_reg[3]/NET0131 ,
		_w23827_,
		_w24558_
	);
	LUT2 #(
		.INIT('h1)
	) name20512 (
		_w24557_,
		_w24558_,
		_w24559_
	);
	LUT2 #(
		.INIT('h4)
	) name20513 (
		_w8715_,
		_w23827_,
		_w24560_
	);
	LUT2 #(
		.INIT('h1)
	) name20514 (
		\bdma_BOVL_reg[2]/NET0131 ,
		_w23827_,
		_w24561_
	);
	LUT2 #(
		.INIT('h1)
	) name20515 (
		_w24560_,
		_w24561_,
		_w24562_
	);
	LUT2 #(
		.INIT('h4)
	) name20516 (
		_w9435_,
		_w23827_,
		_w24563_
	);
	LUT2 #(
		.INIT('h1)
	) name20517 (
		\bdma_BOVL_reg[1]/NET0131 ,
		_w23827_,
		_w24564_
	);
	LUT2 #(
		.INIT('h1)
	) name20518 (
		_w24563_,
		_w24564_,
		_w24565_
	);
	LUT2 #(
		.INIT('h4)
	) name20519 (
		_w7607_,
		_w23827_,
		_w24566_
	);
	LUT2 #(
		.INIT('h1)
	) name20520 (
		\bdma_BOVL_reg[0]/NET0131 ,
		_w23827_,
		_w24567_
	);
	LUT2 #(
		.INIT('h1)
	) name20521 (
		_w24566_,
		_w24567_,
		_w24568_
	);
	LUT2 #(
		.INIT('h4)
	) name20522 (
		_w8113_,
		_w21268_,
		_w24569_
	);
	LUT2 #(
		.INIT('h1)
	) name20523 (
		\bdma_BCTL_reg[3]/NET0131 ,
		_w21268_,
		_w24570_
	);
	LUT2 #(
		.INIT('h1)
	) name20524 (
		_w24569_,
		_w24570_,
		_w24571_
	);
	LUT2 #(
		.INIT('h4)
	) name20525 (
		_w8715_,
		_w21268_,
		_w24572_
	);
	LUT2 #(
		.INIT('h1)
	) name20526 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w21268_,
		_w24573_
	);
	LUT2 #(
		.INIT('h1)
	) name20527 (
		_w24572_,
		_w24573_,
		_w24574_
	);
	LUT2 #(
		.INIT('h4)
	) name20528 (
		_w9435_,
		_w21268_,
		_w24575_
	);
	LUT2 #(
		.INIT('h1)
	) name20529 (
		\bdma_BCTL_reg[1]/NET0131 ,
		_w21268_,
		_w24576_
	);
	LUT2 #(
		.INIT('h1)
	) name20530 (
		_w24575_,
		_w24576_,
		_w24577_
	);
	LUT2 #(
		.INIT('h4)
	) name20531 (
		_w12743_,
		_w21268_,
		_w24578_
	);
	LUT2 #(
		.INIT('h1)
	) name20532 (
		\bdma_BCTL_reg[15]/NET0131 ,
		_w21268_,
		_w24579_
	);
	LUT2 #(
		.INIT('h1)
	) name20533 (
		_w24578_,
		_w24579_,
		_w24580_
	);
	LUT2 #(
		.INIT('h4)
	) name20534 (
		_w12688_,
		_w21268_,
		_w24581_
	);
	LUT2 #(
		.INIT('h1)
	) name20535 (
		\bdma_BCTL_reg[14]/NET0131 ,
		_w21268_,
		_w24582_
	);
	LUT2 #(
		.INIT('h1)
	) name20536 (
		_w24581_,
		_w24582_,
		_w24583_
	);
	LUT2 #(
		.INIT('h4)
	) name20537 (
		_w7607_,
		_w21268_,
		_w24584_
	);
	LUT2 #(
		.INIT('h1)
	) name20538 (
		\bdma_BCTL_reg[0]/NET0131 ,
		_w21268_,
		_w24585_
	);
	LUT2 #(
		.INIT('h1)
	) name20539 (
		_w24584_,
		_w24585_,
		_w24586_
	);
	LUT2 #(
		.INIT('h2)
	) name20540 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001 ,
		_w13789_,
		_w24587_
	);
	LUT2 #(
		.INIT('h8)
	) name20541 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w13789_,
		_w24588_
	);
	LUT2 #(
		.INIT('h1)
	) name20542 (
		_w24587_,
		_w24588_,
		_w24589_
	);
	LUT2 #(
		.INIT('h2)
	) name20543 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001 ,
		_w13789_,
		_w24590_
	);
	LUT2 #(
		.INIT('h8)
	) name20544 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w13789_,
		_w24591_
	);
	LUT2 #(
		.INIT('h1)
	) name20545 (
		_w24590_,
		_w24591_,
		_w24592_
	);
	LUT2 #(
		.INIT('h2)
	) name20546 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001 ,
		_w13775_,
		_w24593_
	);
	LUT2 #(
		.INIT('h8)
	) name20547 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w13775_,
		_w24594_
	);
	LUT2 #(
		.INIT('h1)
	) name20548 (
		_w24593_,
		_w24594_,
		_w24595_
	);
	LUT2 #(
		.INIT('h1)
	) name20549 (
		\sice_ICYC_reg[5]/NET0131 ,
		_w18859_,
		_w24596_
	);
	LUT2 #(
		.INIT('h1)
	) name20550 (
		_w18860_,
		_w24596_,
		_w24597_
	);
	LUT2 #(
		.INIT('h2)
	) name20551 (
		\core_c_psq_lpstk_lps4x22_LPcell_reg[1][1]/P0001 ,
		_w4845_,
		_w24598_
	);
	LUT2 #(
		.INIT('h8)
	) name20552 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		_w4845_,
		_w24599_
	);
	LUT2 #(
		.INIT('h1)
	) name20553 (
		_w24598_,
		_w24599_,
		_w24600_
	);
	LUT2 #(
		.INIT('h2)
	) name20554 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001 ,
		_w13789_,
		_w24601_
	);
	LUT2 #(
		.INIT('h8)
	) name20555 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w13789_,
		_w24602_
	);
	LUT2 #(
		.INIT('h1)
	) name20556 (
		_w24601_,
		_w24602_,
		_w24603_
	);
	LUT2 #(
		.INIT('h2)
	) name20557 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001 ,
		_w13789_,
		_w24604_
	);
	LUT2 #(
		.INIT('h8)
	) name20558 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w13789_,
		_w24605_
	);
	LUT2 #(
		.INIT('h1)
	) name20559 (
		_w24604_,
		_w24605_,
		_w24606_
	);
	LUT2 #(
		.INIT('h2)
	) name20560 (
		_w23766_,
		_w24517_,
		_w24607_
	);
	LUT2 #(
		.INIT('h1)
	) name20561 (
		\core_eu_em_mac_em_reg_my1swe_DO_reg[0]/P0001 ,
		_w23766_,
		_w24608_
	);
	LUT2 #(
		.INIT('h1)
	) name20562 (
		_w24607_,
		_w24608_,
		_w24609_
	);
	LUT2 #(
		.INIT('h2)
	) name20563 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001 ,
		_w13775_,
		_w24610_
	);
	LUT2 #(
		.INIT('h8)
	) name20564 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w13775_,
		_w24611_
	);
	LUT2 #(
		.INIT('h1)
	) name20565 (
		_w24610_,
		_w24611_,
		_w24612_
	);
	LUT2 #(
		.INIT('h2)
	) name20566 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001 ,
		_w13775_,
		_w24613_
	);
	LUT2 #(
		.INIT('h8)
	) name20567 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w13775_,
		_w24614_
	);
	LUT2 #(
		.INIT('h1)
	) name20568 (
		_w24613_,
		_w24614_,
		_w24615_
	);
	LUT2 #(
		.INIT('h2)
	) name20569 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001 ,
		_w13789_,
		_w24616_
	);
	LUT2 #(
		.INIT('h8)
	) name20570 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w13789_,
		_w24617_
	);
	LUT2 #(
		.INIT('h1)
	) name20571 (
		_w24616_,
		_w24617_,
		_w24618_
	);
	LUT2 #(
		.INIT('h2)
	) name20572 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001 ,
		_w13789_,
		_w24619_
	);
	LUT2 #(
		.INIT('h8)
	) name20573 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w13789_,
		_w24620_
	);
	LUT2 #(
		.INIT('h1)
	) name20574 (
		_w24619_,
		_w24620_,
		_w24621_
	);
	LUT2 #(
		.INIT('h2)
	) name20575 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001 ,
		_w13775_,
		_w24622_
	);
	LUT2 #(
		.INIT('h8)
	) name20576 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w13775_,
		_w24623_
	);
	LUT2 #(
		.INIT('h1)
	) name20577 (
		_w24622_,
		_w24623_,
		_w24624_
	);
	LUT2 #(
		.INIT('h2)
	) name20578 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001 ,
		_w13789_,
		_w24625_
	);
	LUT2 #(
		.INIT('h8)
	) name20579 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w13789_,
		_w24626_
	);
	LUT2 #(
		.INIT('h1)
	) name20580 (
		_w24625_,
		_w24626_,
		_w24627_
	);
	LUT2 #(
		.INIT('h4)
	) name20581 (
		_w20150_,
		_w23754_,
		_w24628_
	);
	LUT2 #(
		.INIT('h1)
	) name20582 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[14]/P0001 ,
		_w23754_,
		_w24629_
	);
	LUT2 #(
		.INIT('h1)
	) name20583 (
		_w24628_,
		_w24629_,
		_w24630_
	);
	LUT2 #(
		.INIT('h4)
	) name20584 (
		_w17814_,
		_w23754_,
		_w24631_
	);
	LUT2 #(
		.INIT('h1)
	) name20585 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[2]/P0001 ,
		_w23754_,
		_w24632_
	);
	LUT2 #(
		.INIT('h1)
	) name20586 (
		_w24631_,
		_w24632_,
		_w24633_
	);
	LUT2 #(
		.INIT('h2)
	) name20587 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001 ,
		_w13775_,
		_w24634_
	);
	LUT2 #(
		.INIT('h8)
	) name20588 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w13775_,
		_w24635_
	);
	LUT2 #(
		.INIT('h1)
	) name20589 (
		_w24634_,
		_w24635_,
		_w24636_
	);
	LUT2 #(
		.INIT('h4)
	) name20590 (
		_w18974_,
		_w23754_,
		_w24637_
	);
	LUT2 #(
		.INIT('h1)
	) name20591 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[1]/P0001 ,
		_w23754_,
		_w24638_
	);
	LUT2 #(
		.INIT('h1)
	) name20592 (
		_w24637_,
		_w24638_,
		_w24639_
	);
	LUT2 #(
		.INIT('h2)
	) name20593 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001 ,
		_w13775_,
		_w24640_
	);
	LUT2 #(
		.INIT('h8)
	) name20594 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w13775_,
		_w24641_
	);
	LUT2 #(
		.INIT('h1)
	) name20595 (
		_w24640_,
		_w24641_,
		_w24642_
	);
	LUT2 #(
		.INIT('h8)
	) name20596 (
		\memc_Dwrite_E_reg/NET0131 ,
		_w4117_,
		_w24643_
	);
	LUT2 #(
		.INIT('h8)
	) name20597 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w6956_,
		_w24644_
	);
	LUT2 #(
		.INIT('h8)
	) name20598 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w6120_,
		_w24645_
	);
	LUT2 #(
		.INIT('h8)
	) name20599 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w6108_,
		_w24646_
	);
	LUT2 #(
		.INIT('h1)
	) name20600 (
		_w6107_,
		_w24644_,
		_w24647_
	);
	LUT2 #(
		.INIT('h4)
	) name20601 (
		_w24646_,
		_w24647_,
		_w24648_
	);
	LUT2 #(
		.INIT('h4)
	) name20602 (
		_w24645_,
		_w24648_,
		_w24649_
	);
	LUT2 #(
		.INIT('h2)
	) name20603 (
		_w11742_,
		_w24649_,
		_w24650_
	);
	LUT2 #(
		.INIT('h1)
	) name20604 (
		_w24643_,
		_w24650_,
		_w24651_
	);
	LUT2 #(
		.INIT('h2)
	) name20605 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001 ,
		_w13794_,
		_w24652_
	);
	LUT2 #(
		.INIT('h8)
	) name20606 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w13794_,
		_w24653_
	);
	LUT2 #(
		.INIT('h1)
	) name20607 (
		_w24652_,
		_w24653_,
		_w24654_
	);
	LUT2 #(
		.INIT('h4)
	) name20608 (
		_w21663_,
		_w23754_,
		_w24655_
	);
	LUT2 #(
		.INIT('h1)
	) name20609 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[3]/P0001 ,
		_w23754_,
		_w24656_
	);
	LUT2 #(
		.INIT('h1)
	) name20610 (
		_w24655_,
		_w24656_,
		_w24657_
	);
	LUT2 #(
		.INIT('h2)
	) name20611 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001 ,
		_w13784_,
		_w24658_
	);
	LUT2 #(
		.INIT('h8)
	) name20612 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w13784_,
		_w24659_
	);
	LUT2 #(
		.INIT('h1)
	) name20613 (
		_w24658_,
		_w24659_,
		_w24660_
	);
	LUT2 #(
		.INIT('h2)
	) name20614 (
		_w11265_,
		_w23865_,
		_w24661_
	);
	LUT2 #(
		.INIT('h8)
	) name20615 (
		\sport1_txctl_TX_reg[7]/P0001 ,
		_w23865_,
		_w24662_
	);
	LUT2 #(
		.INIT('h1)
	) name20616 (
		_w24661_,
		_w24662_,
		_w24663_
	);
	LUT2 #(
		.INIT('h2)
	) name20617 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001 ,
		_w13784_,
		_w24664_
	);
	LUT2 #(
		.INIT('h8)
	) name20618 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		_w13784_,
		_w24665_
	);
	LUT2 #(
		.INIT('h1)
	) name20619 (
		_w24664_,
		_w24665_,
		_w24666_
	);
	LUT2 #(
		.INIT('h2)
	) name20620 (
		_w11525_,
		_w23865_,
		_w24667_
	);
	LUT2 #(
		.INIT('h8)
	) name20621 (
		\sport1_txctl_TX_reg[6]/P0001 ,
		_w23865_,
		_w24668_
	);
	LUT2 #(
		.INIT('h1)
	) name20622 (
		_w24667_,
		_w24668_,
		_w24669_
	);
	LUT2 #(
		.INIT('h2)
	) name20623 (
		_w10911_,
		_w23865_,
		_w24670_
	);
	LUT2 #(
		.INIT('h8)
	) name20624 (
		\sport1_txctl_TX_reg[5]/P0001 ,
		_w23865_,
		_w24671_
	);
	LUT2 #(
		.INIT('h1)
	) name20625 (
		_w24670_,
		_w24671_,
		_w24672_
	);
	LUT2 #(
		.INIT('h2)
	) name20626 (
		_w10069_,
		_w23865_,
		_w24673_
	);
	LUT2 #(
		.INIT('h8)
	) name20627 (
		\sport1_txctl_TX_reg[4]/P0001 ,
		_w23865_,
		_w24674_
	);
	LUT2 #(
		.INIT('h1)
	) name20628 (
		_w24673_,
		_w24674_,
		_w24675_
	);
	LUT2 #(
		.INIT('h2)
	) name20629 (
		_w8113_,
		_w23865_,
		_w24676_
	);
	LUT2 #(
		.INIT('h8)
	) name20630 (
		\sport1_txctl_TX_reg[3]/P0001 ,
		_w23865_,
		_w24677_
	);
	LUT2 #(
		.INIT('h1)
	) name20631 (
		_w24676_,
		_w24677_,
		_w24678_
	);
	LUT2 #(
		.INIT('h2)
	) name20632 (
		_w8715_,
		_w23865_,
		_w24679_
	);
	LUT2 #(
		.INIT('h8)
	) name20633 (
		\sport1_txctl_TX_reg[2]/P0001 ,
		_w23865_,
		_w24680_
	);
	LUT2 #(
		.INIT('h1)
	) name20634 (
		_w24679_,
		_w24680_,
		_w24681_
	);
	LUT2 #(
		.INIT('h2)
	) name20635 (
		_w9435_,
		_w23865_,
		_w24682_
	);
	LUT2 #(
		.INIT('h8)
	) name20636 (
		\sport1_txctl_TX_reg[1]/P0001 ,
		_w23865_,
		_w24683_
	);
	LUT2 #(
		.INIT('h1)
	) name20637 (
		_w24682_,
		_w24683_,
		_w24684_
	);
	LUT2 #(
		.INIT('h2)
	) name20638 (
		_w12743_,
		_w23865_,
		_w24685_
	);
	LUT2 #(
		.INIT('h8)
	) name20639 (
		\sport1_txctl_TX_reg[15]/P0001 ,
		_w23865_,
		_w24686_
	);
	LUT2 #(
		.INIT('h1)
	) name20640 (
		_w24685_,
		_w24686_,
		_w24687_
	);
	LUT2 #(
		.INIT('h2)
	) name20641 (
		_w12688_,
		_w23865_,
		_w24688_
	);
	LUT2 #(
		.INIT('h8)
	) name20642 (
		\sport1_txctl_TX_reg[14]/P0001 ,
		_w23865_,
		_w24689_
	);
	LUT2 #(
		.INIT('h1)
	) name20643 (
		_w24688_,
		_w24689_,
		_w24690_
	);
	LUT2 #(
		.INIT('h2)
	) name20644 (
		_w7607_,
		_w23865_,
		_w24691_
	);
	LUT2 #(
		.INIT('h8)
	) name20645 (
		\sport1_txctl_TX_reg[0]/P0001 ,
		_w23865_,
		_w24692_
	);
	LUT2 #(
		.INIT('h1)
	) name20646 (
		_w24691_,
		_w24692_,
		_w24693_
	);
	LUT2 #(
		.INIT('h4)
	) name20647 (
		_w20080_,
		_w23754_,
		_w24694_
	);
	LUT2 #(
		.INIT('h1)
	) name20648 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[4]/P0001 ,
		_w23754_,
		_w24695_
	);
	LUT2 #(
		.INIT('h1)
	) name20649 (
		_w24694_,
		_w24695_,
		_w24696_
	);
	LUT2 #(
		.INIT('h2)
	) name20650 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001 ,
		_w13775_,
		_w24697_
	);
	LUT2 #(
		.INIT('h8)
	) name20651 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w13775_,
		_w24698_
	);
	LUT2 #(
		.INIT('h1)
	) name20652 (
		_w24697_,
		_w24698_,
		_w24699_
	);
	LUT2 #(
		.INIT('h2)
	) name20653 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001 ,
		_w13775_,
		_w24700_
	);
	LUT2 #(
		.INIT('h8)
	) name20654 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w13775_,
		_w24701_
	);
	LUT2 #(
		.INIT('h1)
	) name20655 (
		_w24700_,
		_w24701_,
		_w24702_
	);
	LUT2 #(
		.INIT('h4)
	) name20656 (
		_w22021_,
		_w23814_,
		_w24703_
	);
	LUT2 #(
		.INIT('h1)
	) name20657 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[6]/P0001 ,
		_w23814_,
		_w24704_
	);
	LUT2 #(
		.INIT('h1)
	) name20658 (
		_w24703_,
		_w24704_,
		_w24705_
	);
	LUT2 #(
		.INIT('h4)
	) name20659 (
		_w22030_,
		_w23798_,
		_w24706_
	);
	LUT2 #(
		.INIT('h1)
	) name20660 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[5]/P0001 ,
		_w23798_,
		_w24707_
	);
	LUT2 #(
		.INIT('h1)
	) name20661 (
		_w24706_,
		_w24707_,
		_w24708_
	);
	LUT2 #(
		.INIT('h8)
	) name20662 (
		\core_eu_ec_cun_updateMV_C_reg/P0001 ,
		_w5950_,
		_w24709_
	);
	LUT2 #(
		.INIT('h1)
	) name20663 (
		_w21314_,
		_w24709_,
		_w24710_
	);
	LUT2 #(
		.INIT('h2)
	) name20664 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22924_,
		_w24711_
	);
	LUT2 #(
		.INIT('h1)
	) name20665 (
		_w22770_,
		_w22776_,
		_w24712_
	);
	LUT2 #(
		.INIT('h1)
	) name20666 (
		_w22766_,
		_w22772_,
		_w24713_
	);
	LUT2 #(
		.INIT('h8)
	) name20667 (
		_w22766_,
		_w22772_,
		_w24714_
	);
	LUT2 #(
		.INIT('h2)
	) name20668 (
		_w22709_,
		_w24714_,
		_w24715_
	);
	LUT2 #(
		.INIT('h1)
	) name20669 (
		_w24713_,
		_w24715_,
		_w24716_
	);
	LUT2 #(
		.INIT('h2)
	) name20670 (
		_w24712_,
		_w24716_,
		_w24717_
	);
	LUT2 #(
		.INIT('h4)
	) name20671 (
		_w24712_,
		_w24716_,
		_w24718_
	);
	LUT2 #(
		.INIT('h1)
	) name20672 (
		_w24717_,
		_w24718_,
		_w24719_
	);
	LUT2 #(
		.INIT('h4)
	) name20673 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w24719_,
		_w24720_
	);
	LUT2 #(
		.INIT('h1)
	) name20674 (
		_w24711_,
		_w24720_,
		_w24721_
	);
	LUT2 #(
		.INIT('h4)
	) name20675 (
		_w22012_,
		_w23889_,
		_w24722_
	);
	LUT2 #(
		.INIT('h1)
	) name20676 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[7]/P0001 ,
		_w23889_,
		_w24723_
	);
	LUT2 #(
		.INIT('h1)
	) name20677 (
		_w24722_,
		_w24723_,
		_w24724_
	);
	LUT2 #(
		.INIT('h4)
	) name20678 (
		_w22021_,
		_w23889_,
		_w24725_
	);
	LUT2 #(
		.INIT('h1)
	) name20679 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[6]/P0001 ,
		_w23889_,
		_w24726_
	);
	LUT2 #(
		.INIT('h1)
	) name20680 (
		_w24725_,
		_w24726_,
		_w24727_
	);
	LUT2 #(
		.INIT('h4)
	) name20681 (
		_w22030_,
		_w23889_,
		_w24728_
	);
	LUT2 #(
		.INIT('h1)
	) name20682 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[5]/P0001 ,
		_w23889_,
		_w24729_
	);
	LUT2 #(
		.INIT('h1)
	) name20683 (
		_w24728_,
		_w24729_,
		_w24730_
	);
	LUT2 #(
		.INIT('h4)
	) name20684 (
		_w22039_,
		_w23889_,
		_w24731_
	);
	LUT2 #(
		.INIT('h1)
	) name20685 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[4]/P0001 ,
		_w23889_,
		_w24732_
	);
	LUT2 #(
		.INIT('h1)
	) name20686 (
		_w24731_,
		_w24732_,
		_w24733_
	);
	LUT2 #(
		.INIT('h4)
	) name20687 (
		_w22048_,
		_w23889_,
		_w24734_
	);
	LUT2 #(
		.INIT('h1)
	) name20688 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[3]/P0001 ,
		_w23889_,
		_w24735_
	);
	LUT2 #(
		.INIT('h1)
	) name20689 (
		_w24734_,
		_w24735_,
		_w24736_
	);
	LUT2 #(
		.INIT('h4)
	) name20690 (
		_w22057_,
		_w23889_,
		_w24737_
	);
	LUT2 #(
		.INIT('h1)
	) name20691 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[2]/P0001 ,
		_w23889_,
		_w24738_
	);
	LUT2 #(
		.INIT('h1)
	) name20692 (
		_w24737_,
		_w24738_,
		_w24739_
	);
	LUT2 #(
		.INIT('h4)
	) name20693 (
		_w22151_,
		_w23889_,
		_w24740_
	);
	LUT2 #(
		.INIT('h1)
	) name20694 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[1]/P0001 ,
		_w23889_,
		_w24741_
	);
	LUT2 #(
		.INIT('h1)
	) name20695 (
		_w24740_,
		_w24741_,
		_w24742_
	);
	LUT2 #(
		.INIT('h4)
	) name20696 (
		_w22066_,
		_w23889_,
		_w24743_
	);
	LUT2 #(
		.INIT('h1)
	) name20697 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[15]/P0001 ,
		_w23889_,
		_w24744_
	);
	LUT2 #(
		.INIT('h1)
	) name20698 (
		_w24743_,
		_w24744_,
		_w24745_
	);
	LUT2 #(
		.INIT('h4)
	) name20699 (
		_w22075_,
		_w23889_,
		_w24746_
	);
	LUT2 #(
		.INIT('h1)
	) name20700 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[14]/P0001 ,
		_w23889_,
		_w24747_
	);
	LUT2 #(
		.INIT('h1)
	) name20701 (
		_w24746_,
		_w24747_,
		_w24748_
	);
	LUT2 #(
		.INIT('h2)
	) name20702 (
		_w23889_,
		_w24517_,
		_w24749_
	);
	LUT2 #(
		.INIT('h1)
	) name20703 (
		\core_eu_ea_alu_ea_reg_ay1swe_DO_reg[0]/P0001 ,
		_w23889_,
		_w24750_
	);
	LUT2 #(
		.INIT('h1)
	) name20704 (
		_w24749_,
		_w24750_,
		_w24751_
	);
	LUT2 #(
		.INIT('h4)
	) name20705 (
		_w19972_,
		_w23908_,
		_w24752_
	);
	LUT2 #(
		.INIT('h1)
	) name20706 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[7]/P0001 ,
		_w23908_,
		_w24753_
	);
	LUT2 #(
		.INIT('h1)
	) name20707 (
		_w24752_,
		_w24753_,
		_w24754_
	);
	LUT2 #(
		.INIT('h4)
	) name20708 (
		_w18276_,
		_w23908_,
		_w24755_
	);
	LUT2 #(
		.INIT('h1)
	) name20709 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[6]/P0001 ,
		_w23908_,
		_w24756_
	);
	LUT2 #(
		.INIT('h1)
	) name20710 (
		_w24755_,
		_w24756_,
		_w24757_
	);
	LUT2 #(
		.INIT('h4)
	) name20711 (
		_w20259_,
		_w23908_,
		_w24758_
	);
	LUT2 #(
		.INIT('h1)
	) name20712 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[5]/P0001 ,
		_w23908_,
		_w24759_
	);
	LUT2 #(
		.INIT('h1)
	) name20713 (
		_w24758_,
		_w24759_,
		_w24760_
	);
	LUT2 #(
		.INIT('h4)
	) name20714 (
		_w20080_,
		_w23908_,
		_w24761_
	);
	LUT2 #(
		.INIT('h1)
	) name20715 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[4]/P0001 ,
		_w23908_,
		_w24762_
	);
	LUT2 #(
		.INIT('h1)
	) name20716 (
		_w24761_,
		_w24762_,
		_w24763_
	);
	LUT2 #(
		.INIT('h4)
	) name20717 (
		_w21663_,
		_w23908_,
		_w24764_
	);
	LUT2 #(
		.INIT('h1)
	) name20718 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[3]/P0001 ,
		_w23908_,
		_w24765_
	);
	LUT2 #(
		.INIT('h1)
	) name20719 (
		_w24764_,
		_w24765_,
		_w24766_
	);
	LUT2 #(
		.INIT('h4)
	) name20720 (
		_w17814_,
		_w23908_,
		_w24767_
	);
	LUT2 #(
		.INIT('h1)
	) name20721 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[2]/P0001 ,
		_w23908_,
		_w24768_
	);
	LUT2 #(
		.INIT('h1)
	) name20722 (
		_w24767_,
		_w24768_,
		_w24769_
	);
	LUT2 #(
		.INIT('h4)
	) name20723 (
		_w18974_,
		_w23908_,
		_w24770_
	);
	LUT2 #(
		.INIT('h1)
	) name20724 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[1]/P0001 ,
		_w23908_,
		_w24771_
	);
	LUT2 #(
		.INIT('h1)
	) name20725 (
		_w24770_,
		_w24771_,
		_w24772_
	);
	LUT2 #(
		.INIT('h4)
	) name20726 (
		_w17820_,
		_w23908_,
		_w24773_
	);
	LUT2 #(
		.INIT('h1)
	) name20727 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[15]/P0001 ,
		_w23908_,
		_w24774_
	);
	LUT2 #(
		.INIT('h1)
	) name20728 (
		_w24773_,
		_w24774_,
		_w24775_
	);
	LUT2 #(
		.INIT('h4)
	) name20729 (
		_w20150_,
		_w23908_,
		_w24776_
	);
	LUT2 #(
		.INIT('h1)
	) name20730 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[14]/P0001 ,
		_w23908_,
		_w24777_
	);
	LUT2 #(
		.INIT('h1)
	) name20731 (
		_w24776_,
		_w24777_,
		_w24778_
	);
	LUT2 #(
		.INIT('h4)
	) name20732 (
		_w19559_,
		_w23908_,
		_w24779_
	);
	LUT2 #(
		.INIT('h1)
	) name20733 (
		\core_eu_ea_alu_ea_reg_ax1swe_DO_reg[0]/P0001 ,
		_w23908_,
		_w24780_
	);
	LUT2 #(
		.INIT('h1)
	) name20734 (
		_w24779_,
		_w24780_,
		_w24781_
	);
	LUT2 #(
		.INIT('h4)
	) name20735 (
		_w19972_,
		_w23930_,
		_w24782_
	);
	LUT2 #(
		.INIT('h1)
	) name20736 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[7]/P0001 ,
		_w23930_,
		_w24783_
	);
	LUT2 #(
		.INIT('h1)
	) name20737 (
		_w24782_,
		_w24783_,
		_w24784_
	);
	LUT2 #(
		.INIT('h4)
	) name20738 (
		_w18276_,
		_w23930_,
		_w24785_
	);
	LUT2 #(
		.INIT('h1)
	) name20739 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[6]/P0001 ,
		_w23930_,
		_w24786_
	);
	LUT2 #(
		.INIT('h1)
	) name20740 (
		_w24785_,
		_w24786_,
		_w24787_
	);
	LUT2 #(
		.INIT('h4)
	) name20741 (
		_w20259_,
		_w23930_,
		_w24788_
	);
	LUT2 #(
		.INIT('h1)
	) name20742 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[5]/P0001 ,
		_w23930_,
		_w24789_
	);
	LUT2 #(
		.INIT('h1)
	) name20743 (
		_w24788_,
		_w24789_,
		_w24790_
	);
	LUT2 #(
		.INIT('h4)
	) name20744 (
		_w20080_,
		_w23930_,
		_w24791_
	);
	LUT2 #(
		.INIT('h1)
	) name20745 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[4]/P0001 ,
		_w23930_,
		_w24792_
	);
	LUT2 #(
		.INIT('h1)
	) name20746 (
		_w24791_,
		_w24792_,
		_w24793_
	);
	LUT2 #(
		.INIT('h4)
	) name20747 (
		_w21663_,
		_w23930_,
		_w24794_
	);
	LUT2 #(
		.INIT('h1)
	) name20748 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[3]/P0001 ,
		_w23930_,
		_w24795_
	);
	LUT2 #(
		.INIT('h1)
	) name20749 (
		_w24794_,
		_w24795_,
		_w24796_
	);
	LUT2 #(
		.INIT('h4)
	) name20750 (
		_w17814_,
		_w23930_,
		_w24797_
	);
	LUT2 #(
		.INIT('h1)
	) name20751 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[2]/P0001 ,
		_w23930_,
		_w24798_
	);
	LUT2 #(
		.INIT('h1)
	) name20752 (
		_w24797_,
		_w24798_,
		_w24799_
	);
	LUT2 #(
		.INIT('h4)
	) name20753 (
		_w18974_,
		_w23930_,
		_w24800_
	);
	LUT2 #(
		.INIT('h1)
	) name20754 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[1]/P0001 ,
		_w23930_,
		_w24801_
	);
	LUT2 #(
		.INIT('h1)
	) name20755 (
		_w24800_,
		_w24801_,
		_w24802_
	);
	LUT2 #(
		.INIT('h4)
	) name20756 (
		_w17820_,
		_w23930_,
		_w24803_
	);
	LUT2 #(
		.INIT('h1)
	) name20757 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[15]/P0001 ,
		_w23930_,
		_w24804_
	);
	LUT2 #(
		.INIT('h1)
	) name20758 (
		_w24803_,
		_w24804_,
		_w24805_
	);
	LUT2 #(
		.INIT('h4)
	) name20759 (
		_w20150_,
		_w23930_,
		_w24806_
	);
	LUT2 #(
		.INIT('h1)
	) name20760 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[14]/P0001 ,
		_w23930_,
		_w24807_
	);
	LUT2 #(
		.INIT('h1)
	) name20761 (
		_w24806_,
		_w24807_,
		_w24808_
	);
	LUT2 #(
		.INIT('h4)
	) name20762 (
		_w19559_,
		_w23930_,
		_w24809_
	);
	LUT2 #(
		.INIT('h1)
	) name20763 (
		\core_eu_ea_alu_ea_reg_ax0swe_DO_reg[0]/P0001 ,
		_w23930_,
		_w24810_
	);
	LUT2 #(
		.INIT('h1)
	) name20764 (
		_w24809_,
		_w24810_,
		_w24811_
	);
	LUT2 #(
		.INIT('h4)
	) name20765 (
		_w22066_,
		_w23798_,
		_w24812_
	);
	LUT2 #(
		.INIT('h1)
	) name20766 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[15]/P0001 ,
		_w23798_,
		_w24813_
	);
	LUT2 #(
		.INIT('h1)
	) name20767 (
		_w24812_,
		_w24813_,
		_w24814_
	);
	LUT2 #(
		.INIT('h8)
	) name20768 (
		_w19698_,
		_w21248_,
		_w24815_
	);
	LUT2 #(
		.INIT('h8)
	) name20769 (
		_w23231_,
		_w24815_,
		_w24816_
	);
	LUT2 #(
		.INIT('h8)
	) name20770 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w4118_,
		_w24817_
	);
	LUT2 #(
		.INIT('h1)
	) name20771 (
		_w24816_,
		_w24817_,
		_w24818_
	);
	LUT2 #(
		.INIT('h4)
	) name20772 (
		_w22066_,
		_w23814_,
		_w24819_
	);
	LUT2 #(
		.INIT('h1)
	) name20773 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[15]/P0001 ,
		_w23814_,
		_w24820_
	);
	LUT2 #(
		.INIT('h1)
	) name20774 (
		_w24819_,
		_w24820_,
		_w24821_
	);
	LUT2 #(
		.INIT('h2)
	) name20775 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001 ,
		_w13775_,
		_w24822_
	);
	LUT2 #(
		.INIT('h8)
	) name20776 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		_w13775_,
		_w24823_
	);
	LUT2 #(
		.INIT('h1)
	) name20777 (
		_w24822_,
		_w24823_,
		_w24824_
	);
	LUT2 #(
		.INIT('h4)
	) name20778 (
		_w22151_,
		_w23814_,
		_w24825_
	);
	LUT2 #(
		.INIT('h1)
	) name20779 (
		\core_eu_em_mac_em_reg_my0rwe_DO_reg[1]/P0001 ,
		_w23814_,
		_w24826_
	);
	LUT2 #(
		.INIT('h1)
	) name20780 (
		_w24825_,
		_w24826_,
		_w24827_
	);
	LUT2 #(
		.INIT('h2)
	) name20781 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001 ,
		_w13794_,
		_w24828_
	);
	LUT2 #(
		.INIT('h8)
	) name20782 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w13794_,
		_w24829_
	);
	LUT2 #(
		.INIT('h1)
	) name20783 (
		_w24828_,
		_w24829_,
		_w24830_
	);
	LUT2 #(
		.INIT('h4)
	) name20784 (
		_w20259_,
		_w23754_,
		_w24831_
	);
	LUT2 #(
		.INIT('h1)
	) name20785 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[5]/P0001 ,
		_w23754_,
		_w24832_
	);
	LUT2 #(
		.INIT('h1)
	) name20786 (
		_w24831_,
		_w24832_,
		_w24833_
	);
	LUT2 #(
		.INIT('h2)
	) name20787 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001 ,
		_w13775_,
		_w24834_
	);
	LUT2 #(
		.INIT('h8)
	) name20788 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w13775_,
		_w24835_
	);
	LUT2 #(
		.INIT('h1)
	) name20789 (
		_w24834_,
		_w24835_,
		_w24836_
	);
	LUT2 #(
		.INIT('h4)
	) name20790 (
		_w22075_,
		_w23798_,
		_w24837_
	);
	LUT2 #(
		.INIT('h1)
	) name20791 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[14]/P0001 ,
		_w23798_,
		_w24838_
	);
	LUT2 #(
		.INIT('h1)
	) name20792 (
		_w24837_,
		_w24838_,
		_w24839_
	);
	LUT2 #(
		.INIT('h4)
	) name20793 (
		_w22057_,
		_w23798_,
		_w24840_
	);
	LUT2 #(
		.INIT('h1)
	) name20794 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[2]/P0001 ,
		_w23798_,
		_w24841_
	);
	LUT2 #(
		.INIT('h1)
	) name20795 (
		_w24840_,
		_w24841_,
		_w24842_
	);
	LUT2 #(
		.INIT('h4)
	) name20796 (
		_w22012_,
		_w23798_,
		_w24843_
	);
	LUT2 #(
		.INIT('h1)
	) name20797 (
		\core_eu_em_mac_em_reg_my0swe_DO_reg[7]/P0001 ,
		_w23798_,
		_w24844_
	);
	LUT2 #(
		.INIT('h1)
	) name20798 (
		_w24843_,
		_w24844_,
		_w24845_
	);
	LUT2 #(
		.INIT('h2)
	) name20799 (
		_w23782_,
		_w24517_,
		_w24846_
	);
	LUT2 #(
		.INIT('h1)
	) name20800 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[0]/P0001 ,
		_w23782_,
		_w24847_
	);
	LUT2 #(
		.INIT('h1)
	) name20801 (
		_w24846_,
		_w24847_,
		_w24848_
	);
	LUT2 #(
		.INIT('h4)
	) name20802 (
		_w22057_,
		_w23782_,
		_w24849_
	);
	LUT2 #(
		.INIT('h1)
	) name20803 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[2]/P0001 ,
		_w23782_,
		_w24850_
	);
	LUT2 #(
		.INIT('h1)
	) name20804 (
		_w24849_,
		_w24850_,
		_w24851_
	);
	LUT2 #(
		.INIT('h4)
	) name20805 (
		_w17820_,
		_w23754_,
		_w24852_
	);
	LUT2 #(
		.INIT('h1)
	) name20806 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[15]/P0001 ,
		_w23754_,
		_w24853_
	);
	LUT2 #(
		.INIT('h1)
	) name20807 (
		_w24852_,
		_w24853_,
		_w24854_
	);
	LUT2 #(
		.INIT('h4)
	) name20808 (
		_w19559_,
		_w23754_,
		_w24855_
	);
	LUT2 #(
		.INIT('h1)
	) name20809 (
		\core_eu_es_sht_es_reg_siswe_DO_reg[0]/P0001 ,
		_w23754_,
		_w24856_
	);
	LUT2 #(
		.INIT('h1)
	) name20810 (
		_w24855_,
		_w24856_,
		_w24857_
	);
	LUT2 #(
		.INIT('h4)
	) name20811 (
		_w22030_,
		_w23782_,
		_w24858_
	);
	LUT2 #(
		.INIT('h1)
	) name20812 (
		\core_eu_em_mac_em_reg_my1rwe_DO_reg[5]/P0001 ,
		_w23782_,
		_w24859_
	);
	LUT2 #(
		.INIT('h1)
	) name20813 (
		_w24858_,
		_w24859_,
		_w24860_
	);
	LUT2 #(
		.INIT('h8)
	) name20814 (
		\sice_IDONE_reg/NET0131 ,
		_w5950_,
		_w24861_
	);
	LUT2 #(
		.INIT('h4)
	) name20815 (
		\core_c_dec_NOP_E_reg/P0001 ,
		_w19203_,
		_w24862_
	);
	LUT2 #(
		.INIT('h1)
	) name20816 (
		_w24861_,
		_w24862_,
		_w24863_
	);
	LUT2 #(
		.INIT('h1)
	) name20817 (
		\sice_IIRC_reg[2]/NET0131 ,
		_w18865_,
		_w24864_
	);
	LUT2 #(
		.INIT('h1)
	) name20818 (
		_w18866_,
		_w24864_,
		_w24865_
	);
	LUT2 #(
		.INIT('h4)
	) name20819 (
		\clkc_oscntr_reg_DO_reg[2]/NET0131 ,
		_w20845_,
		_w24866_
	);
	LUT2 #(
		.INIT('h1)
	) name20820 (
		_w20846_,
		_w24866_,
		_w24867_
	);
	LUT2 #(
		.INIT('h1)
	) name20821 (
		\sice_ICYC_reg[2]/NET0131 ,
		_w18856_,
		_w24868_
	);
	LUT2 #(
		.INIT('h1)
	) name20822 (
		_w18857_,
		_w24868_,
		_w24869_
	);
	LUT2 #(
		.INIT('h8)
	) name20823 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		_w17798_,
		_w24870_
	);
	LUT2 #(
		.INIT('h4)
	) name20824 (
		_w21994_,
		_w24870_,
		_w24871_
	);
	LUT2 #(
		.INIT('h1)
	) name20825 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[9]/P0001 ,
		_w24870_,
		_w24872_
	);
	LUT2 #(
		.INIT('h1)
	) name20826 (
		_w24871_,
		_w24872_,
		_w24873_
	);
	LUT2 #(
		.INIT('h2)
	) name20827 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[8]/P0001 ,
		_w24870_,
		_w24874_
	);
	LUT2 #(
		.INIT('h4)
	) name20828 (
		_w22003_,
		_w24870_,
		_w24875_
	);
	LUT2 #(
		.INIT('h1)
	) name20829 (
		_w24874_,
		_w24875_,
		_w24876_
	);
	LUT2 #(
		.INIT('h4)
	) name20830 (
		_w22012_,
		_w24870_,
		_w24877_
	);
	LUT2 #(
		.INIT('h1)
	) name20831 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[7]/P0001 ,
		_w24870_,
		_w24878_
	);
	LUT2 #(
		.INIT('h1)
	) name20832 (
		_w24877_,
		_w24878_,
		_w24879_
	);
	LUT2 #(
		.INIT('h4)
	) name20833 (
		_w22021_,
		_w24870_,
		_w24880_
	);
	LUT2 #(
		.INIT('h1)
	) name20834 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[6]/P0001 ,
		_w24870_,
		_w24881_
	);
	LUT2 #(
		.INIT('h1)
	) name20835 (
		_w24880_,
		_w24881_,
		_w24882_
	);
	LUT2 #(
		.INIT('h4)
	) name20836 (
		_w22030_,
		_w24870_,
		_w24883_
	);
	LUT2 #(
		.INIT('h1)
	) name20837 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[5]/P0001 ,
		_w24870_,
		_w24884_
	);
	LUT2 #(
		.INIT('h1)
	) name20838 (
		_w24883_,
		_w24884_,
		_w24885_
	);
	LUT2 #(
		.INIT('h4)
	) name20839 (
		_w22039_,
		_w24870_,
		_w24886_
	);
	LUT2 #(
		.INIT('h1)
	) name20840 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[4]/P0001 ,
		_w24870_,
		_w24887_
	);
	LUT2 #(
		.INIT('h1)
	) name20841 (
		_w24886_,
		_w24887_,
		_w24888_
	);
	LUT2 #(
		.INIT('h4)
	) name20842 (
		_w22048_,
		_w24870_,
		_w24889_
	);
	LUT2 #(
		.INIT('h1)
	) name20843 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[3]/P0001 ,
		_w24870_,
		_w24890_
	);
	LUT2 #(
		.INIT('h1)
	) name20844 (
		_w24889_,
		_w24890_,
		_w24891_
	);
	LUT2 #(
		.INIT('h4)
	) name20845 (
		_w22057_,
		_w24870_,
		_w24892_
	);
	LUT2 #(
		.INIT('h1)
	) name20846 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[2]/P0001 ,
		_w24870_,
		_w24893_
	);
	LUT2 #(
		.INIT('h1)
	) name20847 (
		_w24892_,
		_w24893_,
		_w24894_
	);
	LUT2 #(
		.INIT('h4)
	) name20848 (
		_w22151_,
		_w24870_,
		_w24895_
	);
	LUT2 #(
		.INIT('h1)
	) name20849 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[1]/P0001 ,
		_w24870_,
		_w24896_
	);
	LUT2 #(
		.INIT('h1)
	) name20850 (
		_w24895_,
		_w24896_,
		_w24897_
	);
	LUT2 #(
		.INIT('h4)
	) name20851 (
		_w22066_,
		_w24870_,
		_w24898_
	);
	LUT2 #(
		.INIT('h1)
	) name20852 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[15]/P0001 ,
		_w24870_,
		_w24899_
	);
	LUT2 #(
		.INIT('h1)
	) name20853 (
		_w24898_,
		_w24899_,
		_w24900_
	);
	LUT2 #(
		.INIT('h4)
	) name20854 (
		_w22075_,
		_w24870_,
		_w24901_
	);
	LUT2 #(
		.INIT('h1)
	) name20855 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[14]/P0001 ,
		_w24870_,
		_w24902_
	);
	LUT2 #(
		.INIT('h1)
	) name20856 (
		_w24901_,
		_w24902_,
		_w24903_
	);
	LUT2 #(
		.INIT('h4)
	) name20857 (
		_w22084_,
		_w24870_,
		_w24904_
	);
	LUT2 #(
		.INIT('h1)
	) name20858 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[13]/P0001 ,
		_w24870_,
		_w24905_
	);
	LUT2 #(
		.INIT('h1)
	) name20859 (
		_w24904_,
		_w24905_,
		_w24906_
	);
	LUT2 #(
		.INIT('h2)
	) name20860 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[12]/P0001 ,
		_w24870_,
		_w24907_
	);
	LUT2 #(
		.INIT('h4)
	) name20861 (
		_w22093_,
		_w24870_,
		_w24908_
	);
	LUT2 #(
		.INIT('h1)
	) name20862 (
		_w24907_,
		_w24908_,
		_w24909_
	);
	LUT2 #(
		.INIT('h2)
	) name20863 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[11]/P0001 ,
		_w24870_,
		_w24910_
	);
	LUT2 #(
		.INIT('h4)
	) name20864 (
		_w22105_,
		_w24870_,
		_w24911_
	);
	LUT2 #(
		.INIT('h1)
	) name20865 (
		_w24910_,
		_w24911_,
		_w24912_
	);
	LUT2 #(
		.INIT('h4)
	) name20866 (
		_w22114_,
		_w24870_,
		_w24913_
	);
	LUT2 #(
		.INIT('h1)
	) name20867 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[10]/P0001 ,
		_w24870_,
		_w24914_
	);
	LUT2 #(
		.INIT('h1)
	) name20868 (
		_w24913_,
		_w24914_,
		_w24915_
	);
	LUT2 #(
		.INIT('h4)
	) name20869 (
		_w24517_,
		_w24870_,
		_w24916_
	);
	LUT2 #(
		.INIT('h1)
	) name20870 (
		\core_eu_ea_alu_ea_reg_ay1rwe_DO_reg[0]/P0001 ,
		_w24870_,
		_w24917_
	);
	LUT2 #(
		.INIT('h1)
	) name20871 (
		_w24916_,
		_w24917_,
		_w24918_
	);
	LUT2 #(
		.INIT('h1)
	) name20872 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 ,
		_w19499_,
		_w24919_
	);
	LUT2 #(
		.INIT('h2)
	) name20873 (
		_w19499_,
		_w23860_,
		_w24920_
	);
	LUT2 #(
		.INIT('h2)
	) name20874 (
		_w19501_,
		_w24919_,
		_w24921_
	);
	LUT2 #(
		.INIT('h4)
	) name20875 (
		_w24920_,
		_w24921_,
		_w24922_
	);
	LUT2 #(
		.INIT('h2)
	) name20876 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[8]/P0001 ,
		_w19383_,
		_w24923_
	);
	LUT2 #(
		.INIT('h1)
	) name20877 (
		_w19508_,
		_w24923_,
		_w24924_
	);
	LUT2 #(
		.INIT('h4)
	) name20878 (
		_w24922_,
		_w24924_,
		_w24925_
	);
	LUT2 #(
		.INIT('h1)
	) name20879 (
		_w18262_,
		_w24925_,
		_w24926_
	);
	LUT2 #(
		.INIT('h4)
	) name20880 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22948_,
		_w24927_
	);
	LUT2 #(
		.INIT('h8)
	) name20881 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19523_,
		_w24928_
	);
	LUT2 #(
		.INIT('h1)
	) name20882 (
		_w24927_,
		_w24928_,
		_w24929_
	);
	LUT2 #(
		.INIT('h2)
	) name20883 (
		_w18262_,
		_w24929_,
		_w24930_
	);
	LUT2 #(
		.INIT('h1)
	) name20884 (
		_w24926_,
		_w24930_,
		_w24931_
	);
	LUT2 #(
		.INIT('h4)
	) name20885 (
		\sport0_rxctl_RXSHT_reg[2]/P0001 ,
		_w20868_,
		_w24932_
	);
	LUT2 #(
		.INIT('h8)
	) name20886 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w20873_,
		_w24933_
	);
	LUT2 #(
		.INIT('h4)
	) name20887 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w8715_,
		_w24934_
	);
	LUT2 #(
		.INIT('h1)
	) name20888 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w20954_,
		_w24935_
	);
	LUT2 #(
		.INIT('h2)
	) name20889 (
		_w20951_,
		_w24935_,
		_w24936_
	);
	LUT2 #(
		.INIT('h4)
	) name20890 (
		_w20951_,
		_w24935_,
		_w24937_
	);
	LUT2 #(
		.INIT('h2)
	) name20891 (
		_w20875_,
		_w24936_,
		_w24938_
	);
	LUT2 #(
		.INIT('h4)
	) name20892 (
		_w24937_,
		_w24938_,
		_w24939_
	);
	LUT2 #(
		.INIT('h1)
	) name20893 (
		_w20868_,
		_w24933_,
		_w24940_
	);
	LUT2 #(
		.INIT('h4)
	) name20894 (
		_w24939_,
		_w24940_,
		_w24941_
	);
	LUT2 #(
		.INIT('h4)
	) name20895 (
		_w24934_,
		_w24941_,
		_w24942_
	);
	LUT2 #(
		.INIT('h1)
	) name20896 (
		_w20871_,
		_w24932_,
		_w24943_
	);
	LUT2 #(
		.INIT('h4)
	) name20897 (
		_w24942_,
		_w24943_,
		_w24944_
	);
	LUT2 #(
		.INIT('h8)
	) name20898 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w20871_,
		_w24945_
	);
	LUT2 #(
		.INIT('h1)
	) name20899 (
		_w24944_,
		_w24945_,
		_w24946_
	);
	LUT2 #(
		.INIT('h1)
	) name20900 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 ,
		_w19499_,
		_w24947_
	);
	LUT2 #(
		.INIT('h4)
	) name20901 (
		_w17836_,
		_w19499_,
		_w24948_
	);
	LUT2 #(
		.INIT('h2)
	) name20902 (
		_w19501_,
		_w24947_,
		_w24949_
	);
	LUT2 #(
		.INIT('h4)
	) name20903 (
		_w24948_,
		_w24949_,
		_w24950_
	);
	LUT2 #(
		.INIT('h2)
	) name20904 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[13]/P0001 ,
		_w19383_,
		_w24951_
	);
	LUT2 #(
		.INIT('h1)
	) name20905 (
		_w19508_,
		_w24951_,
		_w24952_
	);
	LUT2 #(
		.INIT('h4)
	) name20906 (
		_w24950_,
		_w24952_,
		_w24953_
	);
	LUT2 #(
		.INIT('h1)
	) name20907 (
		_w18262_,
		_w24953_,
		_w24954_
	);
	LUT2 #(
		.INIT('h1)
	) name20908 (
		_w17741_,
		_w17770_,
		_w24955_
	);
	LUT2 #(
		.INIT('h1)
	) name20909 (
		_w17737_,
		_w19414_,
		_w24956_
	);
	LUT2 #(
		.INIT('h1)
	) name20910 (
		_w19415_,
		_w24956_,
		_w24957_
	);
	LUT2 #(
		.INIT('h8)
	) name20911 (
		_w24955_,
		_w24957_,
		_w24958_
	);
	LUT2 #(
		.INIT('h1)
	) name20912 (
		_w24955_,
		_w24957_,
		_w24959_
	);
	LUT2 #(
		.INIT('h1)
	) name20913 (
		_w24958_,
		_w24959_,
		_w24960_
	);
	LUT2 #(
		.INIT('h1)
	) name20914 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w24960_,
		_w24961_
	);
	LUT2 #(
		.INIT('h8)
	) name20915 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w22996_,
		_w24962_
	);
	LUT2 #(
		.INIT('h1)
	) name20916 (
		_w24961_,
		_w24962_,
		_w24963_
	);
	LUT2 #(
		.INIT('h2)
	) name20917 (
		_w18262_,
		_w24963_,
		_w24964_
	);
	LUT2 #(
		.INIT('h1)
	) name20918 (
		_w24954_,
		_w24964_,
		_w24965_
	);
	LUT2 #(
		.INIT('h1)
	) name20919 (
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		_w23418_,
		_w24966_
	);
	LUT2 #(
		.INIT('h1)
	) name20920 (
		_w23419_,
		_w24966_,
		_w24967_
	);
	LUT2 #(
		.INIT('h2)
	) name20921 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		_w24968_
	);
	LUT2 #(
		.INIT('h2)
	) name20922 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 ,
		_w18266_,
		_w24969_
	);
	LUT2 #(
		.INIT('h1)
	) name20923 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[3]/P0001 ,
		_w18271_,
		_w24970_
	);
	LUT2 #(
		.INIT('h2)
	) name20924 (
		_w18271_,
		_w21663_,
		_w24971_
	);
	LUT2 #(
		.INIT('h2)
	) name20925 (
		_w18273_,
		_w24970_,
		_w24972_
	);
	LUT2 #(
		.INIT('h4)
	) name20926 (
		_w24971_,
		_w24972_,
		_w24973_
	);
	LUT2 #(
		.INIT('h1)
	) name20927 (
		_w18270_,
		_w24969_,
		_w24974_
	);
	LUT2 #(
		.INIT('h4)
	) name20928 (
		_w24973_,
		_w24974_,
		_w24975_
	);
	LUT2 #(
		.INIT('h1)
	) name20929 (
		_w18262_,
		_w24975_,
		_w24976_
	);
	LUT2 #(
		.INIT('h2)
	) name20930 (
		_w18262_,
		_w19662_,
		_w24977_
	);
	LUT2 #(
		.INIT('h1)
	) name20931 (
		_w24976_,
		_w24977_,
		_w24978_
	);
	LUT2 #(
		.INIT('h8)
	) name20932 (
		_w14752_,
		_w19662_,
		_w24979_
	);
	LUT2 #(
		.INIT('h8)
	) name20933 (
		_w18328_,
		_w21663_,
		_w24980_
	);
	LUT2 #(
		.INIT('h2)
	) name20934 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[3]/P0001 ,
		_w18330_,
		_w24981_
	);
	LUT2 #(
		.INIT('h2)
	) name20935 (
		_w18334_,
		_w24981_,
		_w24982_
	);
	LUT2 #(
		.INIT('h4)
	) name20936 (
		_w24980_,
		_w24982_,
		_w24983_
	);
	LUT2 #(
		.INIT('h1)
	) name20937 (
		_w24979_,
		_w24983_,
		_w24984_
	);
	LUT2 #(
		.INIT('h1)
	) name20938 (
		_w13806_,
		_w14634_,
		_w24985_
	);
	LUT2 #(
		.INIT('h2)
	) name20939 (
		_w13806_,
		_w14600_,
		_w24986_
	);
	LUT2 #(
		.INIT('h1)
	) name20940 (
		_w24985_,
		_w24986_,
		_w24987_
	);
	LUT2 #(
		.INIT('h2)
	) name20941 (
		_w14667_,
		_w24987_,
		_w24988_
	);
	LUT2 #(
		.INIT('h2)
	) name20942 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[5]/P0001 ,
		_w14667_,
		_w24989_
	);
	LUT2 #(
		.INIT('h1)
	) name20943 (
		_w24988_,
		_w24989_,
		_w24990_
	);
	LUT2 #(
		.INIT('h2)
	) name20944 (
		_w13805_,
		_w24987_,
		_w24991_
	);
	LUT2 #(
		.INIT('h2)
	) name20945 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[5]/P0001 ,
		_w13805_,
		_w24992_
	);
	LUT2 #(
		.INIT('h1)
	) name20946 (
		_w24991_,
		_w24992_,
		_w24993_
	);
	LUT2 #(
		.INIT('h1)
	) name20947 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 ,
		_w19499_,
		_w24994_
	);
	LUT2 #(
		.INIT('h2)
	) name20948 (
		_w19499_,
		_w23920_,
		_w24995_
	);
	LUT2 #(
		.INIT('h2)
	) name20949 (
		_w19501_,
		_w24994_,
		_w24996_
	);
	LUT2 #(
		.INIT('h4)
	) name20950 (
		_w24995_,
		_w24996_,
		_w24997_
	);
	LUT2 #(
		.INIT('h2)
	) name20951 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[12]/P0001 ,
		_w19383_,
		_w24998_
	);
	LUT2 #(
		.INIT('h1)
	) name20952 (
		_w19508_,
		_w24998_,
		_w24999_
	);
	LUT2 #(
		.INIT('h4)
	) name20953 (
		_w24997_,
		_w24999_,
		_w25000_
	);
	LUT2 #(
		.INIT('h1)
	) name20954 (
		_w18262_,
		_w25000_,
		_w25001_
	);
	LUT2 #(
		.INIT('h8)
	) name20955 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w24960_,
		_w25002_
	);
	LUT2 #(
		.INIT('h4)
	) name20956 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19419_,
		_w25003_
	);
	LUT2 #(
		.INIT('h1)
	) name20957 (
		_w25002_,
		_w25003_,
		_w25004_
	);
	LUT2 #(
		.INIT('h8)
	) name20958 (
		_w18262_,
		_w25004_,
		_w25005_
	);
	LUT2 #(
		.INIT('h1)
	) name20959 (
		_w25001_,
		_w25005_,
		_w25006_
	);
	LUT2 #(
		.INIT('h1)
	) name20960 (
		_w6107_,
		_w6956_,
		_w25007_
	);
	LUT2 #(
		.INIT('h4)
	) name20961 (
		_w6120_,
		_w25007_,
		_w25008_
	);
	LUT2 #(
		.INIT('h8)
	) name20962 (
		_w18838_,
		_w25008_,
		_w25009_
	);
	LUT2 #(
		.INIT('h4)
	) name20963 (
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		_w25010_
	);
	LUT2 #(
		.INIT('h8)
	) name20964 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w25011_
	);
	LUT2 #(
		.INIT('h8)
	) name20965 (
		_w25010_,
		_w25011_,
		_w25012_
	);
	LUT2 #(
		.INIT('h8)
	) name20966 (
		_w23032_,
		_w25012_,
		_w25013_
	);
	LUT2 #(
		.INIT('h8)
	) name20967 (
		_w14752_,
		_w24929_,
		_w25014_
	);
	LUT2 #(
		.INIT('h8)
	) name20968 (
		_w19776_,
		_w23860_,
		_w25015_
	);
	LUT2 #(
		.INIT('h2)
	) name20969 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[8]/P0001 ,
		_w17809_,
		_w25016_
	);
	LUT2 #(
		.INIT('h2)
	) name20970 (
		_w19780_,
		_w25016_,
		_w25017_
	);
	LUT2 #(
		.INIT('h4)
	) name20971 (
		_w25015_,
		_w25017_,
		_w25018_
	);
	LUT2 #(
		.INIT('h1)
	) name20972 (
		_w25014_,
		_w25018_,
		_w25019_
	);
	LUT2 #(
		.INIT('h8)
	) name20973 (
		\core_c_dec_EXIT_E_reg/P0001 ,
		_w4118_,
		_w25020_
	);
	LUT2 #(
		.INIT('h8)
	) name20974 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w21427_,
		_w25021_
	);
	LUT2 #(
		.INIT('h8)
	) name20975 (
		_w21421_,
		_w25021_,
		_w25022_
	);
	LUT2 #(
		.INIT('h1)
	) name20976 (
		_w25020_,
		_w25022_,
		_w25023_
	);
	LUT2 #(
		.INIT('h8)
	) name20977 (
		_w13150_,
		_w19923_,
		_w25024_
	);
	LUT2 #(
		.INIT('h8)
	) name20978 (
		_w23407_,
		_w25011_,
		_w25025_
	);
	LUT2 #(
		.INIT('h8)
	) name20979 (
		_w23032_,
		_w25025_,
		_w25026_
	);
	LUT2 #(
		.INIT('h8)
	) name20980 (
		_w14752_,
		_w24963_,
		_w25027_
	);
	LUT2 #(
		.INIT('h8)
	) name20981 (
		_w17836_,
		_w19776_,
		_w25028_
	);
	LUT2 #(
		.INIT('h2)
	) name20982 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[13]/P0001 ,
		_w17809_,
		_w25029_
	);
	LUT2 #(
		.INIT('h2)
	) name20983 (
		_w19780_,
		_w25029_,
		_w25030_
	);
	LUT2 #(
		.INIT('h4)
	) name20984 (
		_w25028_,
		_w25030_,
		_w25031_
	);
	LUT2 #(
		.INIT('h1)
	) name20985 (
		_w25027_,
		_w25031_,
		_w25032_
	);
	LUT2 #(
		.INIT('h2)
	) name20986 (
		\sice_IAR_reg[1]/NET0131 ,
		\sice_IAR_reg[2]/NET0131 ,
		_w25033_
	);
	LUT2 #(
		.INIT('h8)
	) name20987 (
		_w25011_,
		_w25033_,
		_w25034_
	);
	LUT2 #(
		.INIT('h8)
	) name20988 (
		_w23032_,
		_w25034_,
		_w25035_
	);
	LUT2 #(
		.INIT('h2)
	) name20989 (
		_w14752_,
		_w25004_,
		_w25036_
	);
	LUT2 #(
		.INIT('h8)
	) name20990 (
		_w19776_,
		_w23920_,
		_w25037_
	);
	LUT2 #(
		.INIT('h2)
	) name20991 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[12]/P0001 ,
		_w17809_,
		_w25038_
	);
	LUT2 #(
		.INIT('h2)
	) name20992 (
		_w19780_,
		_w25038_,
		_w25039_
	);
	LUT2 #(
		.INIT('h4)
	) name20993 (
		_w25037_,
		_w25039_,
		_w25040_
	);
	LUT2 #(
		.INIT('h1)
	) name20994 (
		_w25036_,
		_w25040_,
		_w25041_
	);
	LUT2 #(
		.INIT('h4)
	) name20995 (
		\clkc_RSTtext_reg/P0001 ,
		_w12234_,
		_w25042_
	);
	LUT2 #(
		.INIT('h8)
	) name20996 (
		_w23020_,
		_w25042_,
		_w25043_
	);
	LUT2 #(
		.INIT('h8)
	) name20997 (
		_w20573_,
		_w20574_,
		_w25044_
	);
	LUT2 #(
		.INIT('h1)
	) name20998 (
		\core_c_psq_SSTAT_reg[7]/NET0131 ,
		_w25044_,
		_w25045_
	);
	LUT2 #(
		.INIT('h4)
	) name20999 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w4117_,
		_w25046_
	);
	LUT2 #(
		.INIT('h4)
	) name21000 (
		_w4117_,
		_w19701_,
		_w25047_
	);
	LUT2 #(
		.INIT('h2)
	) name21001 (
		_w4116_,
		_w25046_,
		_w25048_
	);
	LUT2 #(
		.INIT('h4)
	) name21002 (
		_w25047_,
		_w25048_,
		_w25049_
	);
	LUT2 #(
		.INIT('h8)
	) name21003 (
		\core_c_dec_RET_Ed_reg/P0001 ,
		_w4117_,
		_w25050_
	);
	LUT2 #(
		.INIT('h1)
	) name21004 (
		_w21429_,
		_w25050_,
		_w25051_
	);
	LUT2 #(
		.INIT('h2)
	) name21005 (
		_w4116_,
		_w25051_,
		_w25052_
	);
	LUT2 #(
		.INIT('h4)
	) name21006 (
		\sice_IAR_reg[0]/NET0131 ,
		\sice_IAR_reg[3]/NET0131 ,
		_w25053_
	);
	LUT2 #(
		.INIT('h8)
	) name21007 (
		_w25010_,
		_w25053_,
		_w25054_
	);
	LUT2 #(
		.INIT('h8)
	) name21008 (
		_w23032_,
		_w25054_,
		_w25055_
	);
	LUT2 #(
		.INIT('h2)
	) name21009 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_txctl_TCS_reg[1]/NET0131 ,
		_w25056_
	);
	LUT2 #(
		.INIT('h4)
	) name21010 (
		_w19960_,
		_w25056_,
		_w25057_
	);
	LUT2 #(
		.INIT('h8)
	) name21011 (
		\sport0_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w25057_,
		_w25058_
	);
	LUT2 #(
		.INIT('h1)
	) name21012 (
		\sport0_txctl_TSreqi_reg/NET0131 ,
		_w25058_,
		_w25059_
	);
	LUT2 #(
		.INIT('h1)
	) name21013 (
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w20036_,
		_w25060_
	);
	LUT2 #(
		.INIT('h1)
	) name21014 (
		_w23710_,
		_w25060_,
		_w25061_
	);
	LUT2 #(
		.INIT('h4)
	) name21015 (
		_w13750_,
		_w25061_,
		_w25062_
	);
	LUT2 #(
		.INIT('h2)
	) name21016 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w24719_,
		_w25063_
	);
	LUT2 #(
		.INIT('h1)
	) name21017 (
		_w24713_,
		_w24714_,
		_w25064_
	);
	LUT2 #(
		.INIT('h2)
	) name21018 (
		_w22709_,
		_w25064_,
		_w25065_
	);
	LUT2 #(
		.INIT('h4)
	) name21019 (
		_w22709_,
		_w25064_,
		_w25066_
	);
	LUT2 #(
		.INIT('h1)
	) name21020 (
		_w25065_,
		_w25066_,
		_w25067_
	);
	LUT2 #(
		.INIT('h4)
	) name21021 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w25067_,
		_w25068_
	);
	LUT2 #(
		.INIT('h1)
	) name21022 (
		_w25063_,
		_w25068_,
		_w25069_
	);
	LUT2 #(
		.INIT('h2)
	) name21023 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_txctl_TCS_reg[1]/NET0131 ,
		_w25070_
	);
	LUT2 #(
		.INIT('h4)
	) name21024 (
		_w22677_,
		_w25070_,
		_w25071_
	);
	LUT2 #(
		.INIT('h8)
	) name21025 (
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w25071_,
		_w25072_
	);
	LUT2 #(
		.INIT('h1)
	) name21026 (
		\sport1_txctl_TSreqi_reg/NET0131 ,
		_w25072_,
		_w25073_
	);
	LUT2 #(
		.INIT('h8)
	) name21027 (
		_w23028_,
		_w25011_,
		_w25074_
	);
	LUT2 #(
		.INIT('h8)
	) name21028 (
		_w23032_,
		_w25074_,
		_w25075_
	);
	LUT2 #(
		.INIT('h1)
	) name21029 (
		\bdma_BWcnt_reg[2]/NET0131 ,
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w25076_
	);
	LUT2 #(
		.INIT('h4)
	) name21030 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w25076_,
		_w25077_
	);
	LUT2 #(
		.INIT('h8)
	) name21031 (
		_w12525_,
		_w20037_,
		_w25078_
	);
	LUT2 #(
		.INIT('h8)
	) name21032 (
		_w25077_,
		_w25078_,
		_w25079_
	);
	LUT2 #(
		.INIT('h4)
	) name21033 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w19696_,
		_w25080_
	);
	LUT2 #(
		.INIT('h8)
	) name21034 (
		_w21249_,
		_w25080_,
		_w25081_
	);
	LUT2 #(
		.INIT('h8)
	) name21035 (
		_w11741_,
		_w25081_,
		_w25082_
	);
	LUT2 #(
		.INIT('h4)
	) name21036 (
		\sice_IAR_reg[1]/NET0131 ,
		_w23408_,
		_w25083_
	);
	LUT2 #(
		.INIT('h8)
	) name21037 (
		\sice_IAR_reg[2]/NET0131 ,
		_w25083_,
		_w25084_
	);
	LUT2 #(
		.INIT('h8)
	) name21038 (
		_w23032_,
		_w25084_,
		_w25085_
	);
	LUT2 #(
		.INIT('h2)
	) name21039 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19407_,
		_w25086_
	);
	LUT2 #(
		.INIT('h4)
	) name21040 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19368_,
		_w25087_
	);
	LUT2 #(
		.INIT('h1)
	) name21041 (
		_w25086_,
		_w25087_,
		_w25088_
	);
	LUT2 #(
		.INIT('h8)
	) name21042 (
		\core_c_psq_T_IRQ1p_reg/P0001 ,
		\core_c_psq_irq1_de_OUT_reg/P0001 ,
		_w25089_
	);
	LUT2 #(
		.INIT('h1)
	) name21043 (
		\core_c_psq_T_IRQ1p_reg/P0001 ,
		\core_c_psq_irq1_de_OUT_reg/P0001 ,
		_w25090_
	);
	LUT2 #(
		.INIT('h2)
	) name21044 (
		\core_c_psq_irq1_de_IN_syn_reg/P0001 ,
		_w25090_,
		_w25091_
	);
	LUT2 #(
		.INIT('h1)
	) name21045 (
		_w25089_,
		_w25091_,
		_w25092_
	);
	LUT2 #(
		.INIT('h8)
	) name21046 (
		\core_c_psq_T_IRQ0p_reg/P0001 ,
		\core_c_psq_irq0_de_OUT_reg/P0001 ,
		_w25093_
	);
	LUT2 #(
		.INIT('h1)
	) name21047 (
		\core_c_psq_T_IRQ0p_reg/P0001 ,
		\core_c_psq_irq0_de_OUT_reg/P0001 ,
		_w25094_
	);
	LUT2 #(
		.INIT('h2)
	) name21048 (
		\core_c_psq_irq0_de_IN_syn_reg/P0001 ,
		_w25094_,
		_w25095_
	);
	LUT2 #(
		.INIT('h1)
	) name21049 (
		_w25093_,
		_w25095_,
		_w25096_
	);
	LUT2 #(
		.INIT('h2)
	) name21050 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		_w5950_,
		_w25097_
	);
	LUT2 #(
		.INIT('h8)
	) name21051 (
		_w8460_,
		_w25097_,
		_w25098_
	);
	LUT2 #(
		.INIT('h2)
	) name21052 (
		\core_c_psq_IFC_reg[10]/NET0131 ,
		\core_c_psq_IFC_reg[11]/NET0131 ,
		_w25099_
	);
	LUT2 #(
		.INIT('h4)
	) name21053 (
		_w25097_,
		_w25099_,
		_w25100_
	);
	LUT2 #(
		.INIT('h1)
	) name21054 (
		_w25098_,
		_w25100_,
		_w25101_
	);
	LUT2 #(
		.INIT('h8)
	) name21055 (
		\core_c_psq_T_IRQ2p_reg/P0001 ,
		\core_c_psq_irq2_de_OUT_reg/P0001 ,
		_w25102_
	);
	LUT2 #(
		.INIT('h1)
	) name21056 (
		\core_c_psq_T_IRQ2p_reg/P0001 ,
		\core_c_psq_irq2_de_OUT_reg/P0001 ,
		_w25103_
	);
	LUT2 #(
		.INIT('h2)
	) name21057 (
		\core_c_psq_irq2_de_IN_syn_reg/P0001 ,
		_w25103_,
		_w25104_
	);
	LUT2 #(
		.INIT('h1)
	) name21058 (
		_w25102_,
		_w25104_,
		_w25105_
	);
	LUT2 #(
		.INIT('h8)
	) name21059 (
		_w10289_,
		_w25097_,
		_w25106_
	);
	LUT2 #(
		.INIT('h2)
	) name21060 (
		\core_c_psq_IFC_reg[8]/NET0131 ,
		\core_c_psq_IFC_reg[9]/NET0131 ,
		_w25107_
	);
	LUT2 #(
		.INIT('h4)
	) name21061 (
		_w25097_,
		_w25107_,
		_w25108_
	);
	LUT2 #(
		.INIT('h1)
	) name21062 (
		_w25106_,
		_w25108_,
		_w25109_
	);
	LUT2 #(
		.INIT('h8)
	) name21063 (
		\core_c_psq_T_IRQL1p_reg/P0001 ,
		\core_c_psq_irql1_de_OUT_reg/P0001 ,
		_w25110_
	);
	LUT2 #(
		.INIT('h1)
	) name21064 (
		\core_c_psq_T_IRQL1p_reg/P0001 ,
		\core_c_psq_irql1_de_OUT_reg/P0001 ,
		_w25111_
	);
	LUT2 #(
		.INIT('h2)
	) name21065 (
		\core_c_psq_irql1_de_IN_syn_reg/P0001 ,
		_w25111_,
		_w25112_
	);
	LUT2 #(
		.INIT('h1)
	) name21066 (
		_w25110_,
		_w25112_,
		_w25113_
	);
	LUT2 #(
		.INIT('h8)
	) name21067 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		_w17798_,
		_w25114_
	);
	LUT2 #(
		.INIT('h4)
	) name21068 (
		_w17836_,
		_w25114_,
		_w25115_
	);
	LUT2 #(
		.INIT('h1)
	) name21069 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[13]/P0001 ,
		_w25114_,
		_w25116_
	);
	LUT2 #(
		.INIT('h1)
	) name21070 (
		_w25115_,
		_w25116_,
		_w25117_
	);
	LUT2 #(
		.INIT('h8)
	) name21071 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		_w17798_,
		_w25118_
	);
	LUT2 #(
		.INIT('h4)
	) name21072 (
		_w19848_,
		_w25118_,
		_w25119_
	);
	LUT2 #(
		.INIT('h1)
	) name21073 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[10]/P0001 ,
		_w25118_,
		_w25120_
	);
	LUT2 #(
		.INIT('h1)
	) name21074 (
		_w25119_,
		_w25120_,
		_w25121_
	);
	LUT2 #(
		.INIT('h4)
	) name21075 (
		_w23920_,
		_w25118_,
		_w25122_
	);
	LUT2 #(
		.INIT('h1)
	) name21076 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[12]/P0001 ,
		_w25118_,
		_w25123_
	);
	LUT2 #(
		.INIT('h1)
	) name21077 (
		_w25122_,
		_w25123_,
		_w25124_
	);
	LUT2 #(
		.INIT('h8)
	) name21078 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		_w14665_,
		_w25125_
	);
	LUT2 #(
		.INIT('h4)
	) name21079 (
		_w23920_,
		_w25125_,
		_w25126_
	);
	LUT2 #(
		.INIT('h1)
	) name21080 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[12]/P0001 ,
		_w25125_,
		_w25127_
	);
	LUT2 #(
		.INIT('h1)
	) name21081 (
		_w25126_,
		_w25127_,
		_w25128_
	);
	LUT2 #(
		.INIT('h4)
	) name21082 (
		_w23920_,
		_w25114_,
		_w25129_
	);
	LUT2 #(
		.INIT('h1)
	) name21083 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[12]/P0001 ,
		_w25114_,
		_w25130_
	);
	LUT2 #(
		.INIT('h1)
	) name21084 (
		_w25129_,
		_w25130_,
		_w25131_
	);
	LUT2 #(
		.INIT('h8)
	) name21085 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		_w14665_,
		_w25132_
	);
	LUT2 #(
		.INIT('h4)
	) name21086 (
		_w19504_,
		_w25132_,
		_w25133_
	);
	LUT2 #(
		.INIT('h1)
	) name21087 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[9]/P0001 ,
		_w25132_,
		_w25134_
	);
	LUT2 #(
		.INIT('h1)
	) name21088 (
		_w25133_,
		_w25134_,
		_w25135_
	);
	LUT2 #(
		.INIT('h4)
	) name21089 (
		_w17836_,
		_w25132_,
		_w25136_
	);
	LUT2 #(
		.INIT('h1)
	) name21090 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[13]/P0001 ,
		_w25132_,
		_w25137_
	);
	LUT2 #(
		.INIT('h1)
	) name21091 (
		_w25136_,
		_w25137_,
		_w25138_
	);
	LUT2 #(
		.INIT('h4)
	) name21092 (
		_w23920_,
		_w25132_,
		_w25139_
	);
	LUT2 #(
		.INIT('h1)
	) name21093 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[12]/P0001 ,
		_w25132_,
		_w25140_
	);
	LUT2 #(
		.INIT('h1)
	) name21094 (
		_w25139_,
		_w25140_,
		_w25141_
	);
	LUT2 #(
		.INIT('h4)
	) name21095 (
		_w19848_,
		_w25132_,
		_w25142_
	);
	LUT2 #(
		.INIT('h1)
	) name21096 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[10]/P0001 ,
		_w25132_,
		_w25143_
	);
	LUT2 #(
		.INIT('h1)
	) name21097 (
		_w25142_,
		_w25143_,
		_w25144_
	);
	LUT2 #(
		.INIT('h4)
	) name21098 (
		_w23860_,
		_w25114_,
		_w25145_
	);
	LUT2 #(
		.INIT('h1)
	) name21099 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[8]/P0001 ,
		_w25114_,
		_w25146_
	);
	LUT2 #(
		.INIT('h1)
	) name21100 (
		_w25145_,
		_w25146_,
		_w25147_
	);
	LUT2 #(
		.INIT('h4)
	) name21101 (
		_w23860_,
		_w25125_,
		_w25148_
	);
	LUT2 #(
		.INIT('h1)
	) name21102 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[8]/P0001 ,
		_w25125_,
		_w25149_
	);
	LUT2 #(
		.INIT('h1)
	) name21103 (
		_w25148_,
		_w25149_,
		_w25150_
	);
	LUT2 #(
		.INIT('h4)
	) name21104 (
		_w17836_,
		_w25125_,
		_w25151_
	);
	LUT2 #(
		.INIT('h1)
	) name21105 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[13]/P0001 ,
		_w25125_,
		_w25152_
	);
	LUT2 #(
		.INIT('h1)
	) name21106 (
		_w25151_,
		_w25152_,
		_w25153_
	);
	LUT2 #(
		.INIT('h4)
	) name21107 (
		_w23757_,
		_w25125_,
		_w25154_
	);
	LUT2 #(
		.INIT('h1)
	) name21108 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[11]/P0001 ,
		_w25125_,
		_w25155_
	);
	LUT2 #(
		.INIT('h1)
	) name21109 (
		_w25154_,
		_w25155_,
		_w25156_
	);
	LUT2 #(
		.INIT('h4)
	) name21110 (
		_w23860_,
		_w25118_,
		_w25157_
	);
	LUT2 #(
		.INIT('h1)
	) name21111 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[8]/P0001 ,
		_w25118_,
		_w25158_
	);
	LUT2 #(
		.INIT('h1)
	) name21112 (
		_w25157_,
		_w25158_,
		_w25159_
	);
	LUT2 #(
		.INIT('h4)
	) name21113 (
		_w17836_,
		_w25118_,
		_w25160_
	);
	LUT2 #(
		.INIT('h1)
	) name21114 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[13]/P0001 ,
		_w25118_,
		_w25161_
	);
	LUT2 #(
		.INIT('h1)
	) name21115 (
		_w25160_,
		_w25161_,
		_w25162_
	);
	LUT2 #(
		.INIT('h4)
	) name21116 (
		_w19504_,
		_w25118_,
		_w25163_
	);
	LUT2 #(
		.INIT('h1)
	) name21117 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[9]/P0001 ,
		_w25118_,
		_w25164_
	);
	LUT2 #(
		.INIT('h1)
	) name21118 (
		_w25163_,
		_w25164_,
		_w25165_
	);
	LUT2 #(
		.INIT('h4)
	) name21119 (
		_w23757_,
		_w25118_,
		_w25166_
	);
	LUT2 #(
		.INIT('h1)
	) name21120 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[11]/P0001 ,
		_w25118_,
		_w25167_
	);
	LUT2 #(
		.INIT('h1)
	) name21121 (
		_w25166_,
		_w25167_,
		_w25168_
	);
	LUT2 #(
		.INIT('h4)
	) name21122 (
		_w23757_,
		_w25132_,
		_w25169_
	);
	LUT2 #(
		.INIT('h1)
	) name21123 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[11]/P0001 ,
		_w25132_,
		_w25170_
	);
	LUT2 #(
		.INIT('h1)
	) name21124 (
		_w25169_,
		_w25170_,
		_w25171_
	);
	LUT2 #(
		.INIT('h4)
	) name21125 (
		_w19848_,
		_w25125_,
		_w25172_
	);
	LUT2 #(
		.INIT('h1)
	) name21126 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[10]/P0001 ,
		_w25125_,
		_w25173_
	);
	LUT2 #(
		.INIT('h1)
	) name21127 (
		_w25172_,
		_w25173_,
		_w25174_
	);
	LUT2 #(
		.INIT('h4)
	) name21128 (
		_w19504_,
		_w25125_,
		_w25175_
	);
	LUT2 #(
		.INIT('h1)
	) name21129 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[9]/P0001 ,
		_w25125_,
		_w25176_
	);
	LUT2 #(
		.INIT('h1)
	) name21130 (
		_w25175_,
		_w25176_,
		_w25177_
	);
	LUT2 #(
		.INIT('h4)
	) name21131 (
		_w23860_,
		_w25132_,
		_w25178_
	);
	LUT2 #(
		.INIT('h1)
	) name21132 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[8]/P0001 ,
		_w25132_,
		_w25179_
	);
	LUT2 #(
		.INIT('h1)
	) name21133 (
		_w25178_,
		_w25179_,
		_w25180_
	);
	LUT2 #(
		.INIT('h4)
	) name21134 (
		_w23757_,
		_w25114_,
		_w25181_
	);
	LUT2 #(
		.INIT('h1)
	) name21135 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[11]/P0001 ,
		_w25114_,
		_w25182_
	);
	LUT2 #(
		.INIT('h1)
	) name21136 (
		_w25181_,
		_w25182_,
		_w25183_
	);
	LUT2 #(
		.INIT('h4)
	) name21137 (
		_w19848_,
		_w25114_,
		_w25184_
	);
	LUT2 #(
		.INIT('h1)
	) name21138 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[10]/P0001 ,
		_w25114_,
		_w25185_
	);
	LUT2 #(
		.INIT('h1)
	) name21139 (
		_w25184_,
		_w25185_,
		_w25186_
	);
	LUT2 #(
		.INIT('h4)
	) name21140 (
		_w19504_,
		_w25114_,
		_w25187_
	);
	LUT2 #(
		.INIT('h1)
	) name21141 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[9]/P0001 ,
		_w25114_,
		_w25188_
	);
	LUT2 #(
		.INIT('h1)
	) name21142 (
		_w25187_,
		_w25188_,
		_w25189_
	);
	LUT2 #(
		.INIT('h2)
	) name21143 (
		_w4099_,
		_w5950_,
		_w25190_
	);
	LUT2 #(
		.INIT('h2)
	) name21144 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12918_,
		_w25191_
	);
	LUT2 #(
		.INIT('h1)
	) name21145 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w10905_,
		_w25192_
	);
	LUT2 #(
		.INIT('h1)
	) name21146 (
		_w25191_,
		_w25192_,
		_w25193_
	);
	LUT2 #(
		.INIT('h2)
	) name21147 (
		_w25190_,
		_w25193_,
		_w25194_
	);
	LUT2 #(
		.INIT('h2)
	) name21148 (
		\regout_STD_C_reg[5]/P0001 ,
		_w25190_,
		_w25195_
	);
	LUT2 #(
		.INIT('h1)
	) name21149 (
		_w25194_,
		_w25195_,
		_w25196_
	);
	LUT2 #(
		.INIT('h4)
	) name21150 (
		_w17814_,
		_w25132_,
		_w25197_
	);
	LUT2 #(
		.INIT('h1)
	) name21151 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[2]/P0001 ,
		_w25132_,
		_w25198_
	);
	LUT2 #(
		.INIT('h1)
	) name21152 (
		_w25197_,
		_w25198_,
		_w25199_
	);
	LUT2 #(
		.INIT('h4)
	) name21153 (
		\core_c_psq_PCS_reg[10]/NET0131 ,
		_w4094_,
		_w25200_
	);
	LUT2 #(
		.INIT('h1)
	) name21154 (
		T_BRn_pad,
		_w25200_,
		_w25201_
	);
	LUT2 #(
		.INIT('h8)
	) name21155 (
		\core_c_psq_MREQ_reg/NET0131 ,
		_w5679_,
		_w25202_
	);
	LUT2 #(
		.INIT('h8)
	) name21156 (
		_w4112_,
		_w25202_,
		_w25203_
	);
	LUT2 #(
		.INIT('h8)
	) name21157 (
		_w25200_,
		_w25203_,
		_w25204_
	);
	LUT2 #(
		.INIT('h1)
	) name21158 (
		_w25201_,
		_w25204_,
		_w25205_
	);
	LUT2 #(
		.INIT('h8)
	) name21159 (
		\core_c_dec_IRE_reg[6]/NET0131 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w25206_
	);
	LUT2 #(
		.INIT('h4)
	) name21160 (
		_w5950_,
		_w25206_,
		_w25207_
	);
	LUT2 #(
		.INIT('h2)
	) name21161 (
		\core_c_psq_INT_en_reg/NET0131 ,
		_w25207_,
		_w25208_
	);
	LUT2 #(
		.INIT('h8)
	) name21162 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		_w25207_,
		_w25209_
	);
	LUT2 #(
		.INIT('h1)
	) name21163 (
		_w25208_,
		_w25209_,
		_w25210_
	);
	LUT2 #(
		.INIT('h2)
	) name21164 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12751_,
		_w25211_
	);
	LUT2 #(
		.INIT('h1)
	) name21165 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12095_,
		_w25212_
	);
	LUT2 #(
		.INIT('h1)
	) name21166 (
		_w25211_,
		_w25212_,
		_w25213_
	);
	LUT2 #(
		.INIT('h2)
	) name21167 (
		_w25190_,
		_w25213_,
		_w25214_
	);
	LUT2 #(
		.INIT('h2)
	) name21168 (
		\regout_STD_C_reg[15]/P0001 ,
		_w25190_,
		_w25215_
	);
	LUT2 #(
		.INIT('h1)
	) name21169 (
		_w25214_,
		_w25215_,
		_w25216_
	);
	LUT2 #(
		.INIT('h8)
	) name21170 (
		_w10638_,
		_w25097_,
		_w25217_
	);
	LUT2 #(
		.INIT('h4)
	) name21171 (
		\core_c_psq_IFC_reg[8]/NET0131 ,
		\core_c_psq_IFC_reg[9]/NET0131 ,
		_w25218_
	);
	LUT2 #(
		.INIT('h4)
	) name21172 (
		_w25097_,
		_w25218_,
		_w25219_
	);
	LUT2 #(
		.INIT('h1)
	) name21173 (
		_w25217_,
		_w25219_,
		_w25220_
	);
	LUT2 #(
		.INIT('h8)
	) name21174 (
		_w11265_,
		_w25097_,
		_w25221_
	);
	LUT2 #(
		.INIT('h2)
	) name21175 (
		\core_c_psq_IFC_reg[6]/NET0131 ,
		\core_c_psq_IFC_reg[7]/NET0131 ,
		_w25222_
	);
	LUT2 #(
		.INIT('h4)
	) name21176 (
		_w25097_,
		_w25222_,
		_w25223_
	);
	LUT2 #(
		.INIT('h1)
	) name21177 (
		_w25221_,
		_w25223_,
		_w25224_
	);
	LUT2 #(
		.INIT('h8)
	) name21178 (
		\core_c_dec_MTDMOVL_E_reg/P0001 ,
		_w5951_,
		_w25225_
	);
	LUT2 #(
		.INIT('h4)
	) name21179 (
		_w8113_,
		_w25225_,
		_w25226_
	);
	LUT2 #(
		.INIT('h1)
	) name21180 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		_w25225_,
		_w25227_
	);
	LUT2 #(
		.INIT('h1)
	) name21181 (
		_w25226_,
		_w25227_,
		_w25228_
	);
	LUT2 #(
		.INIT('h4)
	) name21182 (
		_w8715_,
		_w25225_,
		_w25229_
	);
	LUT2 #(
		.INIT('h1)
	) name21183 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		_w25225_,
		_w25230_
	);
	LUT2 #(
		.INIT('h1)
	) name21184 (
		_w25229_,
		_w25230_,
		_w25231_
	);
	LUT2 #(
		.INIT('h4)
	) name21185 (
		_w9435_,
		_w25225_,
		_w25232_
	);
	LUT2 #(
		.INIT('h1)
	) name21186 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		_w25225_,
		_w25233_
	);
	LUT2 #(
		.INIT('h1)
	) name21187 (
		_w25232_,
		_w25233_,
		_w25234_
	);
	LUT2 #(
		.INIT('h4)
	) name21188 (
		_w7607_,
		_w25225_,
		_w25235_
	);
	LUT2 #(
		.INIT('h1)
	) name21189 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		_w25225_,
		_w25236_
	);
	LUT2 #(
		.INIT('h1)
	) name21190 (
		_w25235_,
		_w25236_,
		_w25237_
	);
	LUT2 #(
		.INIT('h2)
	) name21191 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12638_,
		_w25238_
	);
	LUT2 #(
		.INIT('h1)
	) name21192 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7334_,
		_w25239_
	);
	LUT2 #(
		.INIT('h1)
	) name21193 (
		_w25238_,
		_w25239_,
		_w25240_
	);
	LUT2 #(
		.INIT('h2)
	) name21194 (
		_w25190_,
		_w25240_,
		_w25241_
	);
	LUT2 #(
		.INIT('h2)
	) name21195 (
		\regout_STD_C_reg[13]/P0001 ,
		_w25190_,
		_w25242_
	);
	LUT2 #(
		.INIT('h1)
	) name21196 (
		_w25241_,
		_w25242_,
		_w25243_
	);
	LUT2 #(
		.INIT('h8)
	) name21197 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w14727_,
		_w25244_
	);
	LUT2 #(
		.INIT('h4)
	) name21198 (
		_w4117_,
		_w25244_,
		_w25245_
	);
	LUT2 #(
		.INIT('h8)
	) name21199 (
		\core_c_dec_imm14_E_reg/P0001 ,
		_w4117_,
		_w25246_
	);
	LUT2 #(
		.INIT('h1)
	) name21200 (
		_w25245_,
		_w25246_,
		_w25247_
	);
	LUT2 #(
		.INIT('h8)
	) name21201 (
		\core_c_dec_DU_Eg_reg/P0001 ,
		_w4118_,
		_w25248_
	);
	LUT2 #(
		.INIT('h8)
	) name21202 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w6118_,
		_w25249_
	);
	LUT2 #(
		.INIT('h8)
	) name21203 (
		_w23231_,
		_w25249_,
		_w25250_
	);
	LUT2 #(
		.INIT('h1)
	) name21204 (
		_w25248_,
		_w25250_,
		_w25251_
	);
	LUT2 #(
		.INIT('h4)
	) name21205 (
		_w20259_,
		_w25114_,
		_w25252_
	);
	LUT2 #(
		.INIT('h1)
	) name21206 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[5]/P0001 ,
		_w25114_,
		_w25253_
	);
	LUT2 #(
		.INIT('h1)
	) name21207 (
		_w25252_,
		_w25253_,
		_w25254_
	);
	LUT2 #(
		.INIT('h4)
	) name21208 (
		_w20259_,
		_w25118_,
		_w25255_
	);
	LUT2 #(
		.INIT('h1)
	) name21209 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[5]/P0001 ,
		_w25118_,
		_w25256_
	);
	LUT2 #(
		.INIT('h1)
	) name21210 (
		_w25255_,
		_w25256_,
		_w25257_
	);
	LUT2 #(
		.INIT('h4)
	) name21211 (
		_w20150_,
		_w25125_,
		_w25258_
	);
	LUT2 #(
		.INIT('h1)
	) name21212 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[14]/P0001 ,
		_w25125_,
		_w25259_
	);
	LUT2 #(
		.INIT('h1)
	) name21213 (
		_w25258_,
		_w25259_,
		_w25260_
	);
	LUT2 #(
		.INIT('h4)
	) name21214 (
		_w19972_,
		_w25132_,
		_w25261_
	);
	LUT2 #(
		.INIT('h1)
	) name21215 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[7]/P0001 ,
		_w25132_,
		_w25262_
	);
	LUT2 #(
		.INIT('h1)
	) name21216 (
		_w25261_,
		_w25262_,
		_w25263_
	);
	LUT2 #(
		.INIT('h4)
	) name21217 (
		_w20259_,
		_w25132_,
		_w25264_
	);
	LUT2 #(
		.INIT('h1)
	) name21218 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[5]/P0001 ,
		_w25132_,
		_w25265_
	);
	LUT2 #(
		.INIT('h1)
	) name21219 (
		_w25264_,
		_w25265_,
		_w25266_
	);
	LUT2 #(
		.INIT('h4)
	) name21220 (
		_w21663_,
		_w25132_,
		_w25267_
	);
	LUT2 #(
		.INIT('h1)
	) name21221 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[3]/P0001 ,
		_w25132_,
		_w25268_
	);
	LUT2 #(
		.INIT('h1)
	) name21222 (
		_w25267_,
		_w25268_,
		_w25269_
	);
	LUT2 #(
		.INIT('h4)
	) name21223 (
		_w18974_,
		_w25132_,
		_w25270_
	);
	LUT2 #(
		.INIT('h1)
	) name21224 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[1]/P0001 ,
		_w25132_,
		_w25271_
	);
	LUT2 #(
		.INIT('h1)
	) name21225 (
		_w25270_,
		_w25271_,
		_w25272_
	);
	LUT2 #(
		.INIT('h4)
	) name21226 (
		_w18276_,
		_w25114_,
		_w25273_
	);
	LUT2 #(
		.INIT('h1)
	) name21227 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[6]/P0001 ,
		_w25114_,
		_w25274_
	);
	LUT2 #(
		.INIT('h1)
	) name21228 (
		_w25273_,
		_w25274_,
		_w25275_
	);
	LUT2 #(
		.INIT('h4)
	) name21229 (
		_w21663_,
		_w25114_,
		_w25276_
	);
	LUT2 #(
		.INIT('h1)
	) name21230 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[3]/P0001 ,
		_w25114_,
		_w25277_
	);
	LUT2 #(
		.INIT('h1)
	) name21231 (
		_w25276_,
		_w25277_,
		_w25278_
	);
	LUT2 #(
		.INIT('h4)
	) name21232 (
		_w17814_,
		_w25114_,
		_w25279_
	);
	LUT2 #(
		.INIT('h1)
	) name21233 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[2]/P0001 ,
		_w25114_,
		_w25280_
	);
	LUT2 #(
		.INIT('h1)
	) name21234 (
		_w25279_,
		_w25280_,
		_w25281_
	);
	LUT2 #(
		.INIT('h4)
	) name21235 (
		_w17820_,
		_w25114_,
		_w25282_
	);
	LUT2 #(
		.INIT('h1)
	) name21236 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[15]/P0001 ,
		_w25114_,
		_w25283_
	);
	LUT2 #(
		.INIT('h1)
	) name21237 (
		_w25282_,
		_w25283_,
		_w25284_
	);
	LUT2 #(
		.INIT('h4)
	) name21238 (
		_w19559_,
		_w25114_,
		_w25285_
	);
	LUT2 #(
		.INIT('h1)
	) name21239 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[0]/P0001 ,
		_w25114_,
		_w25286_
	);
	LUT2 #(
		.INIT('h1)
	) name21240 (
		_w25285_,
		_w25286_,
		_w25287_
	);
	LUT2 #(
		.INIT('h4)
	) name21241 (
		_w19972_,
		_w25125_,
		_w25288_
	);
	LUT2 #(
		.INIT('h1)
	) name21242 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[7]/P0001 ,
		_w25125_,
		_w25289_
	);
	LUT2 #(
		.INIT('h1)
	) name21243 (
		_w25288_,
		_w25289_,
		_w25290_
	);
	LUT2 #(
		.INIT('h4)
	) name21244 (
		_w18276_,
		_w25125_,
		_w25291_
	);
	LUT2 #(
		.INIT('h1)
	) name21245 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[6]/P0001 ,
		_w25125_,
		_w25292_
	);
	LUT2 #(
		.INIT('h1)
	) name21246 (
		_w25291_,
		_w25292_,
		_w25293_
	);
	LUT2 #(
		.INIT('h4)
	) name21247 (
		_w21663_,
		_w25125_,
		_w25294_
	);
	LUT2 #(
		.INIT('h1)
	) name21248 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[3]/P0001 ,
		_w25125_,
		_w25295_
	);
	LUT2 #(
		.INIT('h1)
	) name21249 (
		_w25294_,
		_w25295_,
		_w25296_
	);
	LUT2 #(
		.INIT('h4)
	) name21250 (
		_w17814_,
		_w25125_,
		_w25297_
	);
	LUT2 #(
		.INIT('h1)
	) name21251 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[2]/P0001 ,
		_w25125_,
		_w25298_
	);
	LUT2 #(
		.INIT('h1)
	) name21252 (
		_w25297_,
		_w25298_,
		_w25299_
	);
	LUT2 #(
		.INIT('h4)
	) name21253 (
		_w18276_,
		_w25118_,
		_w25300_
	);
	LUT2 #(
		.INIT('h1)
	) name21254 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[6]/P0001 ,
		_w25118_,
		_w25301_
	);
	LUT2 #(
		.INIT('h1)
	) name21255 (
		_w25300_,
		_w25301_,
		_w25302_
	);
	LUT2 #(
		.INIT('h4)
	) name21256 (
		_w21663_,
		_w25118_,
		_w25303_
	);
	LUT2 #(
		.INIT('h1)
	) name21257 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[3]/P0001 ,
		_w25118_,
		_w25304_
	);
	LUT2 #(
		.INIT('h1)
	) name21258 (
		_w25303_,
		_w25304_,
		_w25305_
	);
	LUT2 #(
		.INIT('h4)
	) name21259 (
		_w17814_,
		_w25118_,
		_w25306_
	);
	LUT2 #(
		.INIT('h1)
	) name21260 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[2]/P0001 ,
		_w25118_,
		_w25307_
	);
	LUT2 #(
		.INIT('h1)
	) name21261 (
		_w25306_,
		_w25307_,
		_w25308_
	);
	LUT2 #(
		.INIT('h4)
	) name21262 (
		_w20150_,
		_w25118_,
		_w25309_
	);
	LUT2 #(
		.INIT('h1)
	) name21263 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[14]/P0001 ,
		_w25118_,
		_w25310_
	);
	LUT2 #(
		.INIT('h1)
	) name21264 (
		_w25309_,
		_w25310_,
		_w25311_
	);
	LUT2 #(
		.INIT('h4)
	) name21265 (
		_w19559_,
		_w25118_,
		_w25312_
	);
	LUT2 #(
		.INIT('h1)
	) name21266 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[0]/P0001 ,
		_w25118_,
		_w25313_
	);
	LUT2 #(
		.INIT('h1)
	) name21267 (
		_w25312_,
		_w25313_,
		_w25314_
	);
	LUT2 #(
		.INIT('h8)
	) name21268 (
		\core_c_dec_RTI_Ed_reg/P0001 ,
		_w4118_,
		_w25315_
	);
	LUT2 #(
		.INIT('h8)
	) name21269 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w4116_,
		_w25316_
	);
	LUT2 #(
		.INIT('h8)
	) name21270 (
		_w21429_,
		_w25316_,
		_w25317_
	);
	LUT2 #(
		.INIT('h1)
	) name21271 (
		_w25315_,
		_w25317_,
		_w25318_
	);
	LUT2 #(
		.INIT('h2)
	) name21272 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w13055_,
		_w25319_
	);
	LUT2 #(
		.INIT('h1)
	) name21273 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w10283_,
		_w25320_
	);
	LUT2 #(
		.INIT('h1)
	) name21274 (
		_w25319_,
		_w25320_,
		_w25321_
	);
	LUT2 #(
		.INIT('h2)
	) name21275 (
		_w25190_,
		_w25321_,
		_w25322_
	);
	LUT2 #(
		.INIT('h2)
	) name21276 (
		\regout_STD_C_reg[9]/P0001 ,
		_w25190_,
		_w25323_
	);
	LUT2 #(
		.INIT('h1)
	) name21277 (
		_w25322_,
		_w25323_,
		_w25324_
	);
	LUT2 #(
		.INIT('h2)
	) name21278 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12850_,
		_w25325_
	);
	LUT2 #(
		.INIT('h1)
	) name21279 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8107_,
		_w25326_
	);
	LUT2 #(
		.INIT('h1)
	) name21280 (
		_w25325_,
		_w25326_,
		_w25327_
	);
	LUT2 #(
		.INIT('h2)
	) name21281 (
		_w25190_,
		_w25327_,
		_w25328_
	);
	LUT2 #(
		.INIT('h2)
	) name21282 (
		\regout_STD_C_reg[3]/P0001 ,
		_w25190_,
		_w25329_
	);
	LUT2 #(
		.INIT('h1)
	) name21283 (
		_w25328_,
		_w25329_,
		_w25330_
	);
	LUT2 #(
		.INIT('h2)
	) name21284 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12570_,
		_w25331_
	);
	LUT2 #(
		.INIT('h1)
	) name21285 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8454_,
		_w25332_
	);
	LUT2 #(
		.INIT('h1)
	) name21286 (
		_w25331_,
		_w25332_,
		_w25333_
	);
	LUT2 #(
		.INIT('h2)
	) name21287 (
		_w25190_,
		_w25333_,
		_w25334_
	);
	LUT2 #(
		.INIT('h2)
	) name21288 (
		\regout_STD_C_reg[11]/P0001 ,
		_w25190_,
		_w25335_
	);
	LUT2 #(
		.INIT('h1)
	) name21289 (
		_w25334_,
		_w25335_,
		_w25336_
	);
	LUT2 #(
		.INIT('h4)
	) name21290 (
		_w18974_,
		_w25125_,
		_w25337_
	);
	LUT2 #(
		.INIT('h1)
	) name21291 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[1]/P0001 ,
		_w25125_,
		_w25338_
	);
	LUT2 #(
		.INIT('h1)
	) name21292 (
		_w25337_,
		_w25338_,
		_w25339_
	);
	LUT2 #(
		.INIT('h8)
	) name21293 (
		_w7859_,
		_w25097_,
		_w25340_
	);
	LUT2 #(
		.INIT('h4)
	) name21294 (
		\core_c_psq_IFC_reg[10]/NET0131 ,
		\core_c_psq_IFC_reg[11]/NET0131 ,
		_w25341_
	);
	LUT2 #(
		.INIT('h4)
	) name21295 (
		_w25097_,
		_w25341_,
		_w25342_
	);
	LUT2 #(
		.INIT('h1)
	) name21296 (
		_w25340_,
		_w25342_,
		_w25343_
	);
	LUT2 #(
		.INIT('h4)
	) name21297 (
		_w20150_,
		_w25114_,
		_w25344_
	);
	LUT2 #(
		.INIT('h1)
	) name21298 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[14]/P0001 ,
		_w25114_,
		_w25345_
	);
	LUT2 #(
		.INIT('h1)
	) name21299 (
		_w25344_,
		_w25345_,
		_w25346_
	);
	LUT2 #(
		.INIT('h4)
	) name21300 (
		_w20080_,
		_w25132_,
		_w25347_
	);
	LUT2 #(
		.INIT('h1)
	) name21301 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[4]/P0001 ,
		_w25132_,
		_w25348_
	);
	LUT2 #(
		.INIT('h1)
	) name21302 (
		_w25347_,
		_w25348_,
		_w25349_
	);
	LUT2 #(
		.INIT('h4)
	) name21303 (
		_w19559_,
		_w25125_,
		_w25350_
	);
	LUT2 #(
		.INIT('h1)
	) name21304 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[0]/P0001 ,
		_w25125_,
		_w25351_
	);
	LUT2 #(
		.INIT('h1)
	) name21305 (
		_w25350_,
		_w25351_,
		_w25352_
	);
	LUT2 #(
		.INIT('h8)
	) name21306 (
		_w8113_,
		_w25097_,
		_w25353_
	);
	LUT2 #(
		.INIT('h2)
	) name21307 (
		\core_c_psq_IFC_reg[2]/NET0131 ,
		\core_c_psq_IFC_reg[3]/NET0131 ,
		_w25354_
	);
	LUT2 #(
		.INIT('h4)
	) name21308 (
		_w25097_,
		_w25354_,
		_w25355_
	);
	LUT2 #(
		.INIT('h1)
	) name21309 (
		_w25353_,
		_w25355_,
		_w25356_
	);
	LUT2 #(
		.INIT('h8)
	) name21310 (
		_w10911_,
		_w25097_,
		_w25357_
	);
	LUT2 #(
		.INIT('h2)
	) name21311 (
		\core_c_psq_IFC_reg[4]/NET0131 ,
		\core_c_psq_IFC_reg[5]/NET0131 ,
		_w25358_
	);
	LUT2 #(
		.INIT('h4)
	) name21312 (
		_w25097_,
		_w25358_,
		_w25359_
	);
	LUT2 #(
		.INIT('h1)
	) name21313 (
		_w25357_,
		_w25359_,
		_w25360_
	);
	LUT2 #(
		.INIT('h4)
	) name21314 (
		_w17820_,
		_w25125_,
		_w25361_
	);
	LUT2 #(
		.INIT('h1)
	) name21315 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[15]/P0001 ,
		_w25125_,
		_w25362_
	);
	LUT2 #(
		.INIT('h1)
	) name21316 (
		_w25361_,
		_w25362_,
		_w25363_
	);
	LUT2 #(
		.INIT('h2)
	) name21317 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12695_,
		_w25364_
	);
	LUT2 #(
		.INIT('h1)
	) name21318 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w11953_,
		_w25365_
	);
	LUT2 #(
		.INIT('h1)
	) name21319 (
		_w25364_,
		_w25365_,
		_w25366_
	);
	LUT2 #(
		.INIT('h2)
	) name21320 (
		_w25190_,
		_w25366_,
		_w25367_
	);
	LUT2 #(
		.INIT('h2)
	) name21321 (
		\regout_STD_C_reg[14]/P0001 ,
		_w25190_,
		_w25368_
	);
	LUT2 #(
		.INIT('h1)
	) name21322 (
		_w25367_,
		_w25368_,
		_w25369_
	);
	LUT2 #(
		.INIT('h4)
	) name21323 (
		_w17820_,
		_w25118_,
		_w25370_
	);
	LUT2 #(
		.INIT('h1)
	) name21324 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[15]/P0001 ,
		_w25118_,
		_w25371_
	);
	LUT2 #(
		.INIT('h1)
	) name21325 (
		_w25370_,
		_w25371_,
		_w25372_
	);
	LUT2 #(
		.INIT('h2)
	) name21326 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12782_,
		_w25373_
	);
	LUT2 #(
		.INIT('h1)
	) name21327 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w9429_,
		_w25374_
	);
	LUT2 #(
		.INIT('h1)
	) name21328 (
		_w25373_,
		_w25374_,
		_w25375_
	);
	LUT2 #(
		.INIT('h2)
	) name21329 (
		_w25190_,
		_w25375_,
		_w25376_
	);
	LUT2 #(
		.INIT('h2)
	) name21330 (
		\regout_STD_C_reg[1]/P0001 ,
		_w25190_,
		_w25377_
	);
	LUT2 #(
		.INIT('h1)
	) name21331 (
		_w25376_,
		_w25377_,
		_w25378_
	);
	LUT2 #(
		.INIT('h4)
	) name21332 (
		_w19972_,
		_w25118_,
		_w25379_
	);
	LUT2 #(
		.INIT('h1)
	) name21333 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[7]/P0001 ,
		_w25118_,
		_w25380_
	);
	LUT2 #(
		.INIT('h1)
	) name21334 (
		_w25379_,
		_w25380_,
		_w25381_
	);
	LUT2 #(
		.INIT('h4)
	) name21335 (
		_w20080_,
		_w25125_,
		_w25382_
	);
	LUT2 #(
		.INIT('h1)
	) name21336 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[4]/P0001 ,
		_w25125_,
		_w25383_
	);
	LUT2 #(
		.INIT('h1)
	) name21337 (
		_w25382_,
		_w25383_,
		_w25384_
	);
	LUT2 #(
		.INIT('h4)
	) name21338 (
		_w18974_,
		_w25114_,
		_w25385_
	);
	LUT2 #(
		.INIT('h1)
	) name21339 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[1]/P0001 ,
		_w25114_,
		_w25386_
	);
	LUT2 #(
		.INIT('h1)
	) name21340 (
		_w25385_,
		_w25386_,
		_w25387_
	);
	LUT2 #(
		.INIT('h2)
	) name21341 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w13021_,
		_w25388_
	);
	LUT2 #(
		.INIT('h1)
	) name21342 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w10632_,
		_w25389_
	);
	LUT2 #(
		.INIT('h1)
	) name21343 (
		_w25388_,
		_w25389_,
		_w25390_
	);
	LUT2 #(
		.INIT('h2)
	) name21344 (
		_w25190_,
		_w25390_,
		_w25391_
	);
	LUT2 #(
		.INIT('h2)
	) name21345 (
		\regout_STD_C_reg[8]/P0001 ,
		_w25190_,
		_w25392_
	);
	LUT2 #(
		.INIT('h1)
	) name21346 (
		_w25391_,
		_w25392_,
		_w25393_
	);
	LUT2 #(
		.INIT('h2)
	) name21347 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12884_,
		_w25394_
	);
	LUT2 #(
		.INIT('h1)
	) name21348 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w10063_,
		_w25395_
	);
	LUT2 #(
		.INIT('h1)
	) name21349 (
		_w25394_,
		_w25395_,
		_w25396_
	);
	LUT2 #(
		.INIT('h2)
	) name21350 (
		_w25190_,
		_w25396_,
		_w25397_
	);
	LUT2 #(
		.INIT('h2)
	) name21351 (
		\regout_STD_C_reg[4]/P0001 ,
		_w25190_,
		_w25398_
	);
	LUT2 #(
		.INIT('h1)
	) name21352 (
		_w25397_,
		_w25398_,
		_w25399_
	);
	LUT2 #(
		.INIT('h4)
	) name21353 (
		_w18276_,
		_w25132_,
		_w25400_
	);
	LUT2 #(
		.INIT('h1)
	) name21354 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[6]/P0001 ,
		_w25132_,
		_w25401_
	);
	LUT2 #(
		.INIT('h1)
	) name21355 (
		_w25400_,
		_w25401_,
		_w25402_
	);
	LUT2 #(
		.INIT('h4)
	) name21356 (
		_w20150_,
		_w25132_,
		_w25403_
	);
	LUT2 #(
		.INIT('h1)
	) name21357 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[14]/P0001 ,
		_w25132_,
		_w25404_
	);
	LUT2 #(
		.INIT('h1)
	) name21358 (
		_w25403_,
		_w25404_,
		_w25405_
	);
	LUT2 #(
		.INIT('h2)
	) name21359 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12473_,
		_w25406_
	);
	LUT2 #(
		.INIT('h1)
	) name21360 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7601_,
		_w25407_
	);
	LUT2 #(
		.INIT('h1)
	) name21361 (
		_w25406_,
		_w25407_,
		_w25408_
	);
	LUT2 #(
		.INIT('h2)
	) name21362 (
		_w25190_,
		_w25408_,
		_w25409_
	);
	LUT2 #(
		.INIT('h2)
	) name21363 (
		\regout_STD_C_reg[0]/P0001 ,
		_w25190_,
		_w25410_
	);
	LUT2 #(
		.INIT('h1)
	) name21364 (
		_w25409_,
		_w25410_,
		_w25411_
	);
	LUT2 #(
		.INIT('h2)
	) name21365 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12986_,
		_w25412_
	);
	LUT2 #(
		.INIT('h1)
	) name21366 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w11259_,
		_w25413_
	);
	LUT2 #(
		.INIT('h1)
	) name21367 (
		_w25412_,
		_w25413_,
		_w25414_
	);
	LUT2 #(
		.INIT('h2)
	) name21368 (
		_w25190_,
		_w25414_,
		_w25415_
	);
	LUT2 #(
		.INIT('h2)
	) name21369 (
		\regout_STD_C_reg[7]/P0001 ,
		_w25190_,
		_w25416_
	);
	LUT2 #(
		.INIT('h1)
	) name21370 (
		_w25415_,
		_w25416_,
		_w25417_
	);
	LUT2 #(
		.INIT('h8)
	) name21371 (
		_w9435_,
		_w25097_,
		_w25418_
	);
	LUT2 #(
		.INIT('h2)
	) name21372 (
		\core_c_psq_IFC_reg[0]/NET0131 ,
		\core_c_psq_IFC_reg[1]/NET0131 ,
		_w25419_
	);
	LUT2 #(
		.INIT('h4)
	) name21373 (
		_w25097_,
		_w25419_,
		_w25420_
	);
	LUT2 #(
		.INIT('h1)
	) name21374 (
		_w25418_,
		_w25420_,
		_w25421_
	);
	LUT2 #(
		.INIT('h2)
	) name21375 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12604_,
		_w25422_
	);
	LUT2 #(
		.INIT('h1)
	) name21376 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w9172_,
		_w25423_
	);
	LUT2 #(
		.INIT('h1)
	) name21377 (
		_w25422_,
		_w25423_,
		_w25424_
	);
	LUT2 #(
		.INIT('h2)
	) name21378 (
		_w25190_,
		_w25424_,
		_w25425_
	);
	LUT2 #(
		.INIT('h2)
	) name21379 (
		\regout_STD_C_reg[12]/P0001 ,
		_w25190_,
		_w25426_
	);
	LUT2 #(
		.INIT('h1)
	) name21380 (
		_w25425_,
		_w25426_,
		_w25427_
	);
	LUT2 #(
		.INIT('h2)
	) name21381 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12816_,
		_w25428_
	);
	LUT2 #(
		.INIT('h1)
	) name21382 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w8709_,
		_w25429_
	);
	LUT2 #(
		.INIT('h1)
	) name21383 (
		_w25428_,
		_w25429_,
		_w25430_
	);
	LUT2 #(
		.INIT('h2)
	) name21384 (
		_w25190_,
		_w25430_,
		_w25431_
	);
	LUT2 #(
		.INIT('h2)
	) name21385 (
		\regout_STD_C_reg[2]/P0001 ,
		_w25190_,
		_w25432_
	);
	LUT2 #(
		.INIT('h1)
	) name21386 (
		_w25431_,
		_w25432_,
		_w25433_
	);
	LUT2 #(
		.INIT('h4)
	) name21387 (
		_w19559_,
		_w25132_,
		_w25434_
	);
	LUT2 #(
		.INIT('h1)
	) name21388 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[0]/P0001 ,
		_w25132_,
		_w25435_
	);
	LUT2 #(
		.INIT('h1)
	) name21389 (
		_w25434_,
		_w25435_,
		_w25436_
	);
	LUT2 #(
		.INIT('h2)
	) name21390 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12536_,
		_w25437_
	);
	LUT2 #(
		.INIT('h1)
	) name21391 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w7853_,
		_w25438_
	);
	LUT2 #(
		.INIT('h1)
	) name21392 (
		_w25437_,
		_w25438_,
		_w25439_
	);
	LUT2 #(
		.INIT('h2)
	) name21393 (
		_w25190_,
		_w25439_,
		_w25440_
	);
	LUT2 #(
		.INIT('h2)
	) name21394 (
		\regout_STD_C_reg[10]/P0001 ,
		_w25190_,
		_w25441_
	);
	LUT2 #(
		.INIT('h1)
	) name21395 (
		_w25440_,
		_w25441_,
		_w25442_
	);
	LUT2 #(
		.INIT('h4)
	) name21396 (
		_w20080_,
		_w25118_,
		_w25443_
	);
	LUT2 #(
		.INIT('h1)
	) name21397 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[4]/P0001 ,
		_w25118_,
		_w25444_
	);
	LUT2 #(
		.INIT('h1)
	) name21398 (
		_w25443_,
		_w25444_,
		_w25445_
	);
	LUT2 #(
		.INIT('h2)
	) name21399 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w12968_,
		_w25446_
	);
	LUT2 #(
		.INIT('h1)
	) name21400 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w11519_,
		_w25447_
	);
	LUT2 #(
		.INIT('h1)
	) name21401 (
		_w25446_,
		_w25447_,
		_w25448_
	);
	LUT2 #(
		.INIT('h2)
	) name21402 (
		_w25190_,
		_w25448_,
		_w25449_
	);
	LUT2 #(
		.INIT('h2)
	) name21403 (
		\regout_STD_C_reg[6]/P0001 ,
		_w25190_,
		_w25450_
	);
	LUT2 #(
		.INIT('h1)
	) name21404 (
		_w25449_,
		_w25450_,
		_w25451_
	);
	LUT2 #(
		.INIT('h4)
	) name21405 (
		_w20080_,
		_w25114_,
		_w25452_
	);
	LUT2 #(
		.INIT('h1)
	) name21406 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[4]/P0001 ,
		_w25114_,
		_w25453_
	);
	LUT2 #(
		.INIT('h1)
	) name21407 (
		_w25452_,
		_w25453_,
		_w25454_
	);
	LUT2 #(
		.INIT('h4)
	) name21408 (
		_w19972_,
		_w25114_,
		_w25455_
	);
	LUT2 #(
		.INIT('h1)
	) name21409 (
		\core_eu_em_mac_em_reg_mx1rwe_DO_reg[7]/P0001 ,
		_w25114_,
		_w25456_
	);
	LUT2 #(
		.INIT('h1)
	) name21410 (
		_w25455_,
		_w25456_,
		_w25457_
	);
	LUT2 #(
		.INIT('h4)
	) name21411 (
		_w20259_,
		_w25125_,
		_w25458_
	);
	LUT2 #(
		.INIT('h1)
	) name21412 (
		\core_eu_em_mac_em_reg_mx0swe_DO_reg[5]/P0001 ,
		_w25125_,
		_w25459_
	);
	LUT2 #(
		.INIT('h1)
	) name21413 (
		_w25458_,
		_w25459_,
		_w25460_
	);
	LUT2 #(
		.INIT('h4)
	) name21414 (
		_w17820_,
		_w25132_,
		_w25461_
	);
	LUT2 #(
		.INIT('h1)
	) name21415 (
		\core_eu_em_mac_em_reg_mx1swe_DO_reg[15]/P0001 ,
		_w25132_,
		_w25462_
	);
	LUT2 #(
		.INIT('h1)
	) name21416 (
		_w25461_,
		_w25462_,
		_w25463_
	);
	LUT2 #(
		.INIT('h4)
	) name21417 (
		_w18974_,
		_w25118_,
		_w25464_
	);
	LUT2 #(
		.INIT('h1)
	) name21418 (
		\core_eu_em_mac_em_reg_mx0rwe_DO_reg[1]/P0001 ,
		_w25118_,
		_w25465_
	);
	LUT2 #(
		.INIT('h1)
	) name21419 (
		_w25464_,
		_w25465_,
		_w25466_
	);
	LUT2 #(
		.INIT('h8)
	) name21420 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w4117_,
		_w25467_
	);
	LUT2 #(
		.INIT('h8)
	) name21421 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w13574_,
		_w25468_
	);
	LUT2 #(
		.INIT('h8)
	) name21422 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w13577_,
		_w25469_
	);
	LUT2 #(
		.INIT('h1)
	) name21423 (
		_w25468_,
		_w25469_,
		_w25470_
	);
	LUT2 #(
		.INIT('h2)
	) name21424 (
		_w11742_,
		_w25470_,
		_w25471_
	);
	LUT2 #(
		.INIT('h1)
	) name21425 (
		_w25467_,
		_w25471_,
		_w25472_
	);
	LUT2 #(
		.INIT('h8)
	) name21426 (
		_w11525_,
		_w25097_,
		_w25473_
	);
	LUT2 #(
		.INIT('h4)
	) name21427 (
		\core_c_psq_IFC_reg[6]/NET0131 ,
		\core_c_psq_IFC_reg[7]/NET0131 ,
		_w25474_
	);
	LUT2 #(
		.INIT('h4)
	) name21428 (
		_w25097_,
		_w25474_,
		_w25475_
	);
	LUT2 #(
		.INIT('h1)
	) name21429 (
		_w25473_,
		_w25475_,
		_w25476_
	);
	LUT2 #(
		.INIT('h8)
	) name21430 (
		_w10069_,
		_w25097_,
		_w25477_
	);
	LUT2 #(
		.INIT('h4)
	) name21431 (
		\core_c_psq_IFC_reg[4]/NET0131 ,
		\core_c_psq_IFC_reg[5]/NET0131 ,
		_w25478_
	);
	LUT2 #(
		.INIT('h4)
	) name21432 (
		_w25097_,
		_w25478_,
		_w25479_
	);
	LUT2 #(
		.INIT('h1)
	) name21433 (
		_w25477_,
		_w25479_,
		_w25480_
	);
	LUT2 #(
		.INIT('h8)
	) name21434 (
		_w8715_,
		_w25097_,
		_w25481_
	);
	LUT2 #(
		.INIT('h4)
	) name21435 (
		\core_c_psq_IFC_reg[2]/NET0131 ,
		\core_c_psq_IFC_reg[3]/NET0131 ,
		_w25482_
	);
	LUT2 #(
		.INIT('h4)
	) name21436 (
		_w25097_,
		_w25482_,
		_w25483_
	);
	LUT2 #(
		.INIT('h1)
	) name21437 (
		_w25481_,
		_w25483_,
		_w25484_
	);
	LUT2 #(
		.INIT('h8)
	) name21438 (
		_w7607_,
		_w25097_,
		_w25485_
	);
	LUT2 #(
		.INIT('h4)
	) name21439 (
		\core_c_psq_IFC_reg[0]/NET0131 ,
		\core_c_psq_IFC_reg[1]/NET0131 ,
		_w25486_
	);
	LUT2 #(
		.INIT('h4)
	) name21440 (
		_w25097_,
		_w25486_,
		_w25487_
	);
	LUT2 #(
		.INIT('h1)
	) name21441 (
		_w25485_,
		_w25487_,
		_w25488_
	);
	LUT2 #(
		.INIT('h2)
	) name21442 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w22408_,
		_w25489_
	);
	LUT2 #(
		.INIT('h1)
	) name21443 (
		\T_TMODE[0]_pad ,
		_w25489_,
		_w25490_
	);
	LUT2 #(
		.INIT('h1)
	) name21444 (
		_w20357_,
		_w25490_,
		_w25491_
	);
	LUT2 #(
		.INIT('h1)
	) name21445 (
		\T_TMODE[0]_pad ,
		_w22404_,
		_w25492_
	);
	LUT2 #(
		.INIT('h1)
	) name21446 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w25492_,
		_w25493_
	);
	LUT2 #(
		.INIT('h4)
	) name21447 (
		\tm_TSR_TMP_reg[4]/NET0131 ,
		_w25493_,
		_w25494_
	);
	LUT2 #(
		.INIT('h4)
	) name21448 (
		\tm_TSR_TMP_reg[5]/NET0131 ,
		_w25494_,
		_w25495_
	);
	LUT2 #(
		.INIT('h4)
	) name21449 (
		\tm_TSR_TMP_reg[6]/NET0131 ,
		_w25495_,
		_w25496_
	);
	LUT2 #(
		.INIT('h2)
	) name21450 (
		\tm_TSR_TMP_reg[7]/NET0131 ,
		_w25496_,
		_w25497_
	);
	LUT2 #(
		.INIT('h4)
	) name21451 (
		\tm_TSR_TMP_reg[7]/NET0131 ,
		_w25496_,
		_w25498_
	);
	LUT2 #(
		.INIT('h1)
	) name21452 (
		_w25497_,
		_w25498_,
		_w25499_
	);
	LUT2 #(
		.INIT('h2)
	) name21453 (
		_w25491_,
		_w25499_,
		_w25500_
	);
	LUT2 #(
		.INIT('h2)
	) name21454 (
		\tm_tsr_reg_DO_reg[7]/NET0131 ,
		_w25491_,
		_w25501_
	);
	LUT2 #(
		.INIT('h1)
	) name21455 (
		_w25500_,
		_w25501_,
		_w25502_
	);
	LUT2 #(
		.INIT('h8)
	) name21456 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		_w17798_,
		_w25503_
	);
	LUT2 #(
		.INIT('h4)
	) name21457 (
		_w19504_,
		_w25503_,
		_w25504_
	);
	LUT2 #(
		.INIT('h1)
	) name21458 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[9]/P0001 ,
		_w25503_,
		_w25505_
	);
	LUT2 #(
		.INIT('h1)
	) name21459 (
		_w25504_,
		_w25505_,
		_w25506_
	);
	LUT2 #(
		.INIT('h4)
	) name21460 (
		_w17836_,
		_w25503_,
		_w25507_
	);
	LUT2 #(
		.INIT('h1)
	) name21461 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[13]/P0001 ,
		_w25503_,
		_w25508_
	);
	LUT2 #(
		.INIT('h1)
	) name21462 (
		_w25507_,
		_w25508_,
		_w25509_
	);
	LUT2 #(
		.INIT('h4)
	) name21463 (
		_w23860_,
		_w25503_,
		_w25510_
	);
	LUT2 #(
		.INIT('h1)
	) name21464 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[8]/P0001 ,
		_w25503_,
		_w25511_
	);
	LUT2 #(
		.INIT('h1)
	) name21465 (
		_w25510_,
		_w25511_,
		_w25512_
	);
	LUT2 #(
		.INIT('h4)
	) name21466 (
		_w18276_,
		_w25503_,
		_w25513_
	);
	LUT2 #(
		.INIT('h1)
	) name21467 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[6]/P0001 ,
		_w25503_,
		_w25514_
	);
	LUT2 #(
		.INIT('h1)
	) name21468 (
		_w25513_,
		_w25514_,
		_w25515_
	);
	LUT2 #(
		.INIT('h4)
	) name21469 (
		_w17814_,
		_w25503_,
		_w25516_
	);
	LUT2 #(
		.INIT('h1)
	) name21470 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[2]/P0001 ,
		_w25503_,
		_w25517_
	);
	LUT2 #(
		.INIT('h1)
	) name21471 (
		_w25516_,
		_w25517_,
		_w25518_
	);
	LUT2 #(
		.INIT('h4)
	) name21472 (
		_w23757_,
		_w25503_,
		_w25519_
	);
	LUT2 #(
		.INIT('h1)
	) name21473 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[11]/P0001 ,
		_w25503_,
		_w25520_
	);
	LUT2 #(
		.INIT('h1)
	) name21474 (
		_w25519_,
		_w25520_,
		_w25521_
	);
	LUT2 #(
		.INIT('h4)
	) name21475 (
		_w19559_,
		_w25503_,
		_w25522_
	);
	LUT2 #(
		.INIT('h1)
	) name21476 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[0]/P0001 ,
		_w25503_,
		_w25523_
	);
	LUT2 #(
		.INIT('h1)
	) name21477 (
		_w25522_,
		_w25523_,
		_w25524_
	);
	LUT2 #(
		.INIT('h4)
	) name21478 (
		_w20259_,
		_w25503_,
		_w25525_
	);
	LUT2 #(
		.INIT('h1)
	) name21479 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[5]/P0001 ,
		_w25503_,
		_w25526_
	);
	LUT2 #(
		.INIT('h1)
	) name21480 (
		_w25525_,
		_w25526_,
		_w25527_
	);
	LUT2 #(
		.INIT('h8)
	) name21481 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		_w17798_,
		_w25528_
	);
	LUT2 #(
		.INIT('h4)
	) name21482 (
		_w23860_,
		_w25528_,
		_w25529_
	);
	LUT2 #(
		.INIT('h1)
	) name21483 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[8]/P0001 ,
		_w25528_,
		_w25530_
	);
	LUT2 #(
		.INIT('h1)
	) name21484 (
		_w25529_,
		_w25530_,
		_w25531_
	);
	LUT2 #(
		.INIT('h4)
	) name21485 (
		_w17820_,
		_w25503_,
		_w25532_
	);
	LUT2 #(
		.INIT('h1)
	) name21486 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[15]/P0001 ,
		_w25503_,
		_w25533_
	);
	LUT2 #(
		.INIT('h1)
	) name21487 (
		_w25532_,
		_w25533_,
		_w25534_
	);
	LUT2 #(
		.INIT('h8)
	) name21488 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		_w17798_,
		_w25535_
	);
	LUT2 #(
		.INIT('h4)
	) name21489 (
		_w19504_,
		_w25535_,
		_w25536_
	);
	LUT2 #(
		.INIT('h1)
	) name21490 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[9]/P0001 ,
		_w25535_,
		_w25537_
	);
	LUT2 #(
		.INIT('h1)
	) name21491 (
		_w25536_,
		_w25537_,
		_w25538_
	);
	LUT2 #(
		.INIT('h4)
	) name21492 (
		_w23860_,
		_w25535_,
		_w25539_
	);
	LUT2 #(
		.INIT('h1)
	) name21493 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[8]/P0001 ,
		_w25535_,
		_w25540_
	);
	LUT2 #(
		.INIT('h1)
	) name21494 (
		_w25539_,
		_w25540_,
		_w25541_
	);
	LUT2 #(
		.INIT('h4)
	) name21495 (
		_w19972_,
		_w25535_,
		_w25542_
	);
	LUT2 #(
		.INIT('h1)
	) name21496 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[7]/P0001 ,
		_w25535_,
		_w25543_
	);
	LUT2 #(
		.INIT('h1)
	) name21497 (
		_w25542_,
		_w25543_,
		_w25544_
	);
	LUT2 #(
		.INIT('h4)
	) name21498 (
		_w18276_,
		_w25535_,
		_w25545_
	);
	LUT2 #(
		.INIT('h1)
	) name21499 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[6]/P0001 ,
		_w25535_,
		_w25546_
	);
	LUT2 #(
		.INIT('h1)
	) name21500 (
		_w25545_,
		_w25546_,
		_w25547_
	);
	LUT2 #(
		.INIT('h4)
	) name21501 (
		_w20259_,
		_w25535_,
		_w25548_
	);
	LUT2 #(
		.INIT('h1)
	) name21502 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[5]/P0001 ,
		_w25535_,
		_w25549_
	);
	LUT2 #(
		.INIT('h1)
	) name21503 (
		_w25548_,
		_w25549_,
		_w25550_
	);
	LUT2 #(
		.INIT('h4)
	) name21504 (
		_w20080_,
		_w25535_,
		_w25551_
	);
	LUT2 #(
		.INIT('h1)
	) name21505 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[4]/P0001 ,
		_w25535_,
		_w25552_
	);
	LUT2 #(
		.INIT('h1)
	) name21506 (
		_w25551_,
		_w25552_,
		_w25553_
	);
	LUT2 #(
		.INIT('h4)
	) name21507 (
		_w21663_,
		_w25535_,
		_w25554_
	);
	LUT2 #(
		.INIT('h1)
	) name21508 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[3]/P0001 ,
		_w25535_,
		_w25555_
	);
	LUT2 #(
		.INIT('h1)
	) name21509 (
		_w25554_,
		_w25555_,
		_w25556_
	);
	LUT2 #(
		.INIT('h4)
	) name21510 (
		_w17814_,
		_w25535_,
		_w25557_
	);
	LUT2 #(
		.INIT('h1)
	) name21511 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[2]/P0001 ,
		_w25535_,
		_w25558_
	);
	LUT2 #(
		.INIT('h1)
	) name21512 (
		_w25557_,
		_w25558_,
		_w25559_
	);
	LUT2 #(
		.INIT('h4)
	) name21513 (
		_w18974_,
		_w25535_,
		_w25560_
	);
	LUT2 #(
		.INIT('h1)
	) name21514 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[1]/P0001 ,
		_w25535_,
		_w25561_
	);
	LUT2 #(
		.INIT('h1)
	) name21515 (
		_w25560_,
		_w25561_,
		_w25562_
	);
	LUT2 #(
		.INIT('h4)
	) name21516 (
		_w17820_,
		_w25535_,
		_w25563_
	);
	LUT2 #(
		.INIT('h1)
	) name21517 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[15]/P0001 ,
		_w25535_,
		_w25564_
	);
	LUT2 #(
		.INIT('h1)
	) name21518 (
		_w25563_,
		_w25564_,
		_w25565_
	);
	LUT2 #(
		.INIT('h4)
	) name21519 (
		_w20150_,
		_w25535_,
		_w25566_
	);
	LUT2 #(
		.INIT('h1)
	) name21520 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[14]/P0001 ,
		_w25535_,
		_w25567_
	);
	LUT2 #(
		.INIT('h1)
	) name21521 (
		_w25566_,
		_w25567_,
		_w25568_
	);
	LUT2 #(
		.INIT('h4)
	) name21522 (
		_w17836_,
		_w25535_,
		_w25569_
	);
	LUT2 #(
		.INIT('h1)
	) name21523 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[13]/P0001 ,
		_w25535_,
		_w25570_
	);
	LUT2 #(
		.INIT('h1)
	) name21524 (
		_w25569_,
		_w25570_,
		_w25571_
	);
	LUT2 #(
		.INIT('h4)
	) name21525 (
		_w23920_,
		_w25535_,
		_w25572_
	);
	LUT2 #(
		.INIT('h1)
	) name21526 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[12]/P0001 ,
		_w25535_,
		_w25573_
	);
	LUT2 #(
		.INIT('h1)
	) name21527 (
		_w25572_,
		_w25573_,
		_w25574_
	);
	LUT2 #(
		.INIT('h4)
	) name21528 (
		_w23757_,
		_w25535_,
		_w25575_
	);
	LUT2 #(
		.INIT('h1)
	) name21529 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[11]/P0001 ,
		_w25535_,
		_w25576_
	);
	LUT2 #(
		.INIT('h1)
	) name21530 (
		_w25575_,
		_w25576_,
		_w25577_
	);
	LUT2 #(
		.INIT('h4)
	) name21531 (
		_w19848_,
		_w25535_,
		_w25578_
	);
	LUT2 #(
		.INIT('h1)
	) name21532 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[10]/P0001 ,
		_w25535_,
		_w25579_
	);
	LUT2 #(
		.INIT('h1)
	) name21533 (
		_w25578_,
		_w25579_,
		_w25580_
	);
	LUT2 #(
		.INIT('h4)
	) name21534 (
		_w19559_,
		_w25535_,
		_w25581_
	);
	LUT2 #(
		.INIT('h1)
	) name21535 (
		\core_eu_ea_alu_ea_reg_ax1rwe_DO_reg[0]/P0001 ,
		_w25535_,
		_w25582_
	);
	LUT2 #(
		.INIT('h1)
	) name21536 (
		_w25581_,
		_w25582_,
		_w25583_
	);
	LUT2 #(
		.INIT('h4)
	) name21537 (
		_w19504_,
		_w25528_,
		_w25584_
	);
	LUT2 #(
		.INIT('h1)
	) name21538 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[9]/P0001 ,
		_w25528_,
		_w25585_
	);
	LUT2 #(
		.INIT('h1)
	) name21539 (
		_w25584_,
		_w25585_,
		_w25586_
	);
	LUT2 #(
		.INIT('h4)
	) name21540 (
		_w19972_,
		_w25528_,
		_w25587_
	);
	LUT2 #(
		.INIT('h1)
	) name21541 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[7]/P0001 ,
		_w25528_,
		_w25588_
	);
	LUT2 #(
		.INIT('h1)
	) name21542 (
		_w25587_,
		_w25588_,
		_w25589_
	);
	LUT2 #(
		.INIT('h4)
	) name21543 (
		_w18276_,
		_w25528_,
		_w25590_
	);
	LUT2 #(
		.INIT('h1)
	) name21544 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[6]/P0001 ,
		_w25528_,
		_w25591_
	);
	LUT2 #(
		.INIT('h1)
	) name21545 (
		_w25590_,
		_w25591_,
		_w25592_
	);
	LUT2 #(
		.INIT('h4)
	) name21546 (
		_w20259_,
		_w25528_,
		_w25593_
	);
	LUT2 #(
		.INIT('h1)
	) name21547 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[5]/P0001 ,
		_w25528_,
		_w25594_
	);
	LUT2 #(
		.INIT('h1)
	) name21548 (
		_w25593_,
		_w25594_,
		_w25595_
	);
	LUT2 #(
		.INIT('h4)
	) name21549 (
		_w20080_,
		_w25528_,
		_w25596_
	);
	LUT2 #(
		.INIT('h1)
	) name21550 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[4]/P0001 ,
		_w25528_,
		_w25597_
	);
	LUT2 #(
		.INIT('h1)
	) name21551 (
		_w25596_,
		_w25597_,
		_w25598_
	);
	LUT2 #(
		.INIT('h4)
	) name21552 (
		_w21663_,
		_w25528_,
		_w25599_
	);
	LUT2 #(
		.INIT('h1)
	) name21553 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[3]/P0001 ,
		_w25528_,
		_w25600_
	);
	LUT2 #(
		.INIT('h1)
	) name21554 (
		_w25599_,
		_w25600_,
		_w25601_
	);
	LUT2 #(
		.INIT('h4)
	) name21555 (
		_w17814_,
		_w25528_,
		_w25602_
	);
	LUT2 #(
		.INIT('h1)
	) name21556 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[2]/P0001 ,
		_w25528_,
		_w25603_
	);
	LUT2 #(
		.INIT('h1)
	) name21557 (
		_w25602_,
		_w25603_,
		_w25604_
	);
	LUT2 #(
		.INIT('h4)
	) name21558 (
		_w18974_,
		_w25528_,
		_w25605_
	);
	LUT2 #(
		.INIT('h1)
	) name21559 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[1]/P0001 ,
		_w25528_,
		_w25606_
	);
	LUT2 #(
		.INIT('h1)
	) name21560 (
		_w25605_,
		_w25606_,
		_w25607_
	);
	LUT2 #(
		.INIT('h4)
	) name21561 (
		_w17836_,
		_w25528_,
		_w25608_
	);
	LUT2 #(
		.INIT('h1)
	) name21562 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[13]/P0001 ,
		_w25528_,
		_w25609_
	);
	LUT2 #(
		.INIT('h1)
	) name21563 (
		_w25608_,
		_w25609_,
		_w25610_
	);
	LUT2 #(
		.INIT('h4)
	) name21564 (
		_w23920_,
		_w25528_,
		_w25611_
	);
	LUT2 #(
		.INIT('h1)
	) name21565 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[12]/P0001 ,
		_w25528_,
		_w25612_
	);
	LUT2 #(
		.INIT('h1)
	) name21566 (
		_w25611_,
		_w25612_,
		_w25613_
	);
	LUT2 #(
		.INIT('h4)
	) name21567 (
		_w23757_,
		_w25528_,
		_w25614_
	);
	LUT2 #(
		.INIT('h1)
	) name21568 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[11]/P0001 ,
		_w25528_,
		_w25615_
	);
	LUT2 #(
		.INIT('h1)
	) name21569 (
		_w25614_,
		_w25615_,
		_w25616_
	);
	LUT2 #(
		.INIT('h4)
	) name21570 (
		_w19848_,
		_w25528_,
		_w25617_
	);
	LUT2 #(
		.INIT('h1)
	) name21571 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[10]/P0001 ,
		_w25528_,
		_w25618_
	);
	LUT2 #(
		.INIT('h1)
	) name21572 (
		_w25617_,
		_w25618_,
		_w25619_
	);
	LUT2 #(
		.INIT('h4)
	) name21573 (
		_w19559_,
		_w25528_,
		_w25620_
	);
	LUT2 #(
		.INIT('h1)
	) name21574 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[0]/P0001 ,
		_w25528_,
		_w25621_
	);
	LUT2 #(
		.INIT('h1)
	) name21575 (
		_w25620_,
		_w25621_,
		_w25622_
	);
	LUT2 #(
		.INIT('h4)
	) name21576 (
		_w19972_,
		_w25503_,
		_w25623_
	);
	LUT2 #(
		.INIT('h1)
	) name21577 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[7]/P0001 ,
		_w25503_,
		_w25624_
	);
	LUT2 #(
		.INIT('h1)
	) name21578 (
		_w25623_,
		_w25624_,
		_w25625_
	);
	LUT2 #(
		.INIT('h4)
	) name21579 (
		_w20080_,
		_w25503_,
		_w25626_
	);
	LUT2 #(
		.INIT('h1)
	) name21580 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[4]/P0001 ,
		_w25503_,
		_w25627_
	);
	LUT2 #(
		.INIT('h1)
	) name21581 (
		_w25626_,
		_w25627_,
		_w25628_
	);
	LUT2 #(
		.INIT('h4)
	) name21582 (
		_w21663_,
		_w25503_,
		_w25629_
	);
	LUT2 #(
		.INIT('h1)
	) name21583 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[3]/P0001 ,
		_w25503_,
		_w25630_
	);
	LUT2 #(
		.INIT('h1)
	) name21584 (
		_w25629_,
		_w25630_,
		_w25631_
	);
	LUT2 #(
		.INIT('h4)
	) name21585 (
		_w18974_,
		_w25503_,
		_w25632_
	);
	LUT2 #(
		.INIT('h1)
	) name21586 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[1]/P0001 ,
		_w25503_,
		_w25633_
	);
	LUT2 #(
		.INIT('h1)
	) name21587 (
		_w25632_,
		_w25633_,
		_w25634_
	);
	LUT2 #(
		.INIT('h4)
	) name21588 (
		_w20150_,
		_w25503_,
		_w25635_
	);
	LUT2 #(
		.INIT('h1)
	) name21589 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[14]/P0001 ,
		_w25503_,
		_w25636_
	);
	LUT2 #(
		.INIT('h1)
	) name21590 (
		_w25635_,
		_w25636_,
		_w25637_
	);
	LUT2 #(
		.INIT('h4)
	) name21591 (
		_w23920_,
		_w25503_,
		_w25638_
	);
	LUT2 #(
		.INIT('h1)
	) name21592 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[12]/P0001 ,
		_w25503_,
		_w25639_
	);
	LUT2 #(
		.INIT('h1)
	) name21593 (
		_w25638_,
		_w25639_,
		_w25640_
	);
	LUT2 #(
		.INIT('h4)
	) name21594 (
		_w19848_,
		_w25503_,
		_w25641_
	);
	LUT2 #(
		.INIT('h1)
	) name21595 (
		\core_eu_es_sht_es_reg_sirwe_DO_reg[10]/P0001 ,
		_w25503_,
		_w25642_
	);
	LUT2 #(
		.INIT('h1)
	) name21596 (
		_w25641_,
		_w25642_,
		_w25643_
	);
	LUT2 #(
		.INIT('h4)
	) name21597 (
		_w20150_,
		_w25528_,
		_w25644_
	);
	LUT2 #(
		.INIT('h1)
	) name21598 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[14]/P0001 ,
		_w25528_,
		_w25645_
	);
	LUT2 #(
		.INIT('h1)
	) name21599 (
		_w25644_,
		_w25645_,
		_w25646_
	);
	LUT2 #(
		.INIT('h4)
	) name21600 (
		_w17820_,
		_w25528_,
		_w25647_
	);
	LUT2 #(
		.INIT('h1)
	) name21601 (
		\core_eu_ea_alu_ea_reg_ax0rwe_DO_reg[15]/P0001 ,
		_w25528_,
		_w25648_
	);
	LUT2 #(
		.INIT('h1)
	) name21602 (
		_w25647_,
		_w25648_,
		_w25649_
	);
	LUT2 #(
		.INIT('h8)
	) name21603 (
		\PIO_oe[8]_pad ,
		\PIO_oe[9]_pad ,
		_w25650_
	);
	LUT2 #(
		.INIT('h8)
	) name21604 (
		\memc_MMR_web_reg/NET0131 ,
		_w25650_,
		_w25651_
	);
	LUT2 #(
		.INIT('h2)
	) name21605 (
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w25651_,
		_w25652_
	);
	LUT2 #(
		.INIT('h8)
	) name21606 (
		\pio_PIO_RES_OUT_reg[9]/P0001 ,
		_w25651_,
		_w25653_
	);
	LUT2 #(
		.INIT('h1)
	) name21607 (
		_w25652_,
		_w25653_,
		_w25654_
	);
	LUT2 #(
		.INIT('h8)
	) name21608 (
		\PIO_oe[0]_pad ,
		\PIO_oe[1]_pad ,
		_w25655_
	);
	LUT2 #(
		.INIT('h8)
	) name21609 (
		\memc_MMR_web_reg/NET0131 ,
		_w25655_,
		_w25656_
	);
	LUT2 #(
		.INIT('h2)
	) name21610 (
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w25656_,
		_w25657_
	);
	LUT2 #(
		.INIT('h8)
	) name21611 (
		\pio_PIO_RES_OUT_reg[1]/P0001 ,
		_w25656_,
		_w25658_
	);
	LUT2 #(
		.INIT('h1)
	) name21612 (
		_w25657_,
		_w25658_,
		_w25659_
	);
	LUT2 #(
		.INIT('h8)
	) name21613 (
		\PIO_oe[10]_pad ,
		\PIO_oe[11]_pad ,
		_w25660_
	);
	LUT2 #(
		.INIT('h8)
	) name21614 (
		\memc_MMR_web_reg/NET0131 ,
		_w25660_,
		_w25661_
	);
	LUT2 #(
		.INIT('h2)
	) name21615 (
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w25661_,
		_w25662_
	);
	LUT2 #(
		.INIT('h8)
	) name21616 (
		\pio_PIO_RES_OUT_reg[11]/P0001 ,
		_w25661_,
		_w25663_
	);
	LUT2 #(
		.INIT('h1)
	) name21617 (
		_w25662_,
		_w25663_,
		_w25664_
	);
	LUT2 #(
		.INIT('h8)
	) name21618 (
		\PIO_oe[2]_pad ,
		\PIO_oe[3]_pad ,
		_w25665_
	);
	LUT2 #(
		.INIT('h8)
	) name21619 (
		\memc_MMR_web_reg/NET0131 ,
		_w25665_,
		_w25666_
	);
	LUT2 #(
		.INIT('h2)
	) name21620 (
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w25666_,
		_w25667_
	);
	LUT2 #(
		.INIT('h8)
	) name21621 (
		\pio_PIO_RES_OUT_reg[3]/P0001 ,
		_w25666_,
		_w25668_
	);
	LUT2 #(
		.INIT('h1)
	) name21622 (
		_w25667_,
		_w25668_,
		_w25669_
	);
	LUT2 #(
		.INIT('h8)
	) name21623 (
		\PIO_oe[6]_pad ,
		\PIO_oe[7]_pad ,
		_w25670_
	);
	LUT2 #(
		.INIT('h8)
	) name21624 (
		\memc_MMR_web_reg/NET0131 ,
		_w25670_,
		_w25671_
	);
	LUT2 #(
		.INIT('h2)
	) name21625 (
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w25671_,
		_w25672_
	);
	LUT2 #(
		.INIT('h8)
	) name21626 (
		\pio_PIO_RES_OUT_reg[7]/P0001 ,
		_w25671_,
		_w25673_
	);
	LUT2 #(
		.INIT('h1)
	) name21627 (
		_w25672_,
		_w25673_,
		_w25674_
	);
	LUT2 #(
		.INIT('h2)
	) name21628 (
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w25651_,
		_w25675_
	);
	LUT2 #(
		.INIT('h8)
	) name21629 (
		\pio_PIO_RES_OUT_reg[8]/P0001 ,
		_w25651_,
		_w25676_
	);
	LUT2 #(
		.INIT('h1)
	) name21630 (
		_w25675_,
		_w25676_,
		_w25677_
	);
	LUT2 #(
		.INIT('h8)
	) name21631 (
		\PIO_oe[4]_pad ,
		\PIO_oe[5]_pad ,
		_w25678_
	);
	LUT2 #(
		.INIT('h8)
	) name21632 (
		\memc_MMR_web_reg/NET0131 ,
		_w25678_,
		_w25679_
	);
	LUT2 #(
		.INIT('h2)
	) name21633 (
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w25679_,
		_w25680_
	);
	LUT2 #(
		.INIT('h8)
	) name21634 (
		\pio_PIO_RES_OUT_reg[5]/P0001 ,
		_w25679_,
		_w25681_
	);
	LUT2 #(
		.INIT('h1)
	) name21635 (
		_w25680_,
		_w25681_,
		_w25682_
	);
	LUT2 #(
		.INIT('h2)
	) name21636 (
		PWDACK_pad,
		\clkc_SLEEP_reg/NET0131 ,
		_w25683_
	);
	LUT2 #(
		.INIT('h8)
	) name21637 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w25683_,
		_w25684_
	);
	LUT2 #(
		.INIT('h2)
	) name21638 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		_w25684_,
		_w25685_
	);
	LUT2 #(
		.INIT('h4)
	) name21639 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		_w25684_,
		_w25686_
	);
	LUT2 #(
		.INIT('h1)
	) name21640 (
		_w25685_,
		_w25686_,
		_w25687_
	);
	LUT2 #(
		.INIT('h2)
	) name21641 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w6023_,
		_w25688_
	);
	LUT2 #(
		.INIT('h8)
	) name21642 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w6023_,
		_w25689_
	);
	LUT2 #(
		.INIT('h1)
	) name21643 (
		_w25688_,
		_w25689_,
		_w25690_
	);
	LUT2 #(
		.INIT('h1)
	) name21644 (
		_w4117_,
		_w25690_,
		_w25691_
	);
	LUT2 #(
		.INIT('h8)
	) name21645 (
		\core_dag_ilm2reg_M_E_reg[1]/NET0131 ,
		_w4117_,
		_w25692_
	);
	LUT2 #(
		.INIT('h1)
	) name21646 (
		_w25691_,
		_w25692_,
		_w25693_
	);
	LUT2 #(
		.INIT('h2)
	) name21647 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w6023_,
		_w25694_
	);
	LUT2 #(
		.INIT('h8)
	) name21648 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w6023_,
		_w25695_
	);
	LUT2 #(
		.INIT('h1)
	) name21649 (
		_w25694_,
		_w25695_,
		_w25696_
	);
	LUT2 #(
		.INIT('h1)
	) name21650 (
		_w4117_,
		_w25696_,
		_w25697_
	);
	LUT2 #(
		.INIT('h8)
	) name21651 (
		\core_dag_ilm2reg_M_E_reg[0]/NET0131 ,
		_w4117_,
		_w25698_
	);
	LUT2 #(
		.INIT('h1)
	) name21652 (
		_w25697_,
		_w25698_,
		_w25699_
	);
	LUT2 #(
		.INIT('h4)
	) name21653 (
		_w13585_,
		_w13593_,
		_w25700_
	);
	LUT2 #(
		.INIT('h2)
	) name21654 (
		_w13563_,
		_w13585_,
		_w25701_
	);
	LUT2 #(
		.INIT('h4)
	) name21655 (
		_w13585_,
		_w13590_,
		_w25702_
	);
	LUT2 #(
		.INIT('h4)
	) name21656 (
		_w13585_,
		_w13600_,
		_w25703_
	);
	LUT2 #(
		.INIT('h8)
	) name21657 (
		\tm_tcr_reg_DO_reg[8]/NET0131 ,
		_w20355_,
		_w25704_
	);
	LUT2 #(
		.INIT('h4)
	) name21658 (
		\tm_tpr_reg_DO_reg[8]/NET0131 ,
		_w22400_,
		_w25705_
	);
	LUT2 #(
		.INIT('h2)
	) name21659 (
		\tm_TCR_TMP_reg[8]/NET0131 ,
		_w22411_,
		_w25706_
	);
	LUT2 #(
		.INIT('h1)
	) name21660 (
		_w22400_,
		_w25706_,
		_w25707_
	);
	LUT2 #(
		.INIT('h4)
	) name21661 (
		_w23697_,
		_w25707_,
		_w25708_
	);
	LUT2 #(
		.INIT('h1)
	) name21662 (
		_w20355_,
		_w25705_,
		_w25709_
	);
	LUT2 #(
		.INIT('h4)
	) name21663 (
		_w25708_,
		_w25709_,
		_w25710_
	);
	LUT2 #(
		.INIT('h1)
	) name21664 (
		_w25704_,
		_w25710_,
		_w25711_
	);
	LUT2 #(
		.INIT('h4)
	) name21665 (
		_w11758_,
		_w12232_,
		_w25712_
	);
	LUT2 #(
		.INIT('h4)
	) name21666 (
		_w11758_,
		_w12230_,
		_w25713_
	);
	LUT2 #(
		.INIT('h4)
	) name21667 (
		_w11758_,
		_w12228_,
		_w25714_
	);
	LUT2 #(
		.INIT('h4)
	) name21668 (
		_w11758_,
		_w12225_,
		_w25715_
	);
	LUT2 #(
		.INIT('h4)
	) name21669 (
		_w11758_,
		_w12221_,
		_w25716_
	);
	LUT2 #(
		.INIT('h4)
	) name21670 (
		_w11758_,
		_w12219_,
		_w25717_
	);
	LUT2 #(
		.INIT('h4)
	) name21671 (
		_w11758_,
		_w12216_,
		_w25718_
	);
	LUT2 #(
		.INIT('h4)
	) name21672 (
		_w11758_,
		_w12213_,
		_w25719_
	);
	LUT2 #(
		.INIT('h2)
	) name21673 (
		_w11735_,
		_w11758_,
		_w25720_
	);
	LUT2 #(
		.INIT('h4)
	) name21674 (
		_w13585_,
		_w13607_,
		_w25721_
	);
	LUT2 #(
		.INIT('h4)
	) name21675 (
		_w13585_,
		_w13595_,
		_w25722_
	);
	LUT2 #(
		.INIT('h4)
	) name21676 (
		_w13585_,
		_w13603_,
		_w25723_
	);
	LUT2 #(
		.INIT('h4)
	) name21677 (
		_w13585_,
		_w13605_,
		_w25724_
	);
	LUT2 #(
		.INIT('h4)
	) name21678 (
		_w4117_,
		_w6023_,
		_w25725_
	);
	LUT2 #(
		.INIT('h8)
	) name21679 (
		\core_c_dec_Double_E_reg/P0001 ,
		_w4117_,
		_w25726_
	);
	LUT2 #(
		.INIT('h1)
	) name21680 (
		_w25725_,
		_w25726_,
		_w25727_
	);
	LUT2 #(
		.INIT('h2)
	) name21681 (
		_w4116_,
		_w25727_,
		_w25728_
	);
	LUT2 #(
		.INIT('h1)
	) name21682 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w4117_,
		_w25729_
	);
	LUT2 #(
		.INIT('h4)
	) name21683 (
		\core_eu_ec_cun_COND_E_reg[0]/P0001 ,
		_w4117_,
		_w25730_
	);
	LUT2 #(
		.INIT('h2)
	) name21684 (
		_w4150_,
		_w25729_,
		_w25731_
	);
	LUT2 #(
		.INIT('h4)
	) name21685 (
		_w25730_,
		_w25731_,
		_w25732_
	);
	LUT2 #(
		.INIT('h8)
	) name21686 (
		\core_eu_ec_cun_COND_E_reg[1]/P0001 ,
		_w4117_,
		_w25733_
	);
	LUT2 #(
		.INIT('h2)
	) name21687 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w4117_,
		_w25734_
	);
	LUT2 #(
		.INIT('h1)
	) name21688 (
		_w25733_,
		_w25734_,
		_w25735_
	);
	LUT2 #(
		.INIT('h2)
	) name21689 (
		_w4150_,
		_w25735_,
		_w25736_
	);
	LUT2 #(
		.INIT('h4)
	) name21690 (
		\clkc_Awake_reg/NET0131 ,
		_w25042_,
		_w25737_
	);
	LUT2 #(
		.INIT('h8)
	) name21691 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w23429_,
		_w25738_
	);
	LUT2 #(
		.INIT('h1)
	) name21692 (
		_w11739_,
		_w11749_,
		_w25739_
	);
	LUT2 #(
		.INIT('h1)
	) name21693 (
		_w13581_,
		_w13583_,
		_w25740_
	);
	LUT2 #(
		.INIT('h4)
	) name21694 (
		_w22981_,
		_w23132_,
		_w25741_
	);
	LUT2 #(
		.INIT('h2)
	) name21695 (
		_w22970_,
		_w23143_,
		_w25742_
	);
	LUT2 #(
		.INIT('h8)
	) name21696 (
		_w25741_,
		_w25742_,
		_w25743_
	);
	LUT2 #(
		.INIT('h8)
	) name21697 (
		_w19266_,
		_w25743_,
		_w25744_
	);
	LUT2 #(
		.INIT('h8)
	) name21698 (
		_w22970_,
		_w23143_,
		_w25745_
	);
	LUT2 #(
		.INIT('h8)
	) name21699 (
		_w25741_,
		_w25745_,
		_w25746_
	);
	LUT2 #(
		.INIT('h4)
	) name21700 (
		_w19266_,
		_w25746_,
		_w25747_
	);
	LUT2 #(
		.INIT('h8)
	) name21701 (
		_w22981_,
		_w23132_,
		_w25748_
	);
	LUT2 #(
		.INIT('h4)
	) name21702 (
		_w22970_,
		_w23143_,
		_w25749_
	);
	LUT2 #(
		.INIT('h8)
	) name21703 (
		_w25748_,
		_w25749_,
		_w25750_
	);
	LUT2 #(
		.INIT('h8)
	) name21704 (
		_w19296_,
		_w25750_,
		_w25751_
	);
	LUT2 #(
		.INIT('h1)
	) name21705 (
		_w22981_,
		_w23132_,
		_w25752_
	);
	LUT2 #(
		.INIT('h8)
	) name21706 (
		_w25745_,
		_w25752_,
		_w25753_
	);
	LUT2 #(
		.INIT('h8)
	) name21707 (
		_w19263_,
		_w25753_,
		_w25754_
	);
	LUT2 #(
		.INIT('h8)
	) name21708 (
		_w25742_,
		_w25752_,
		_w25755_
	);
	LUT2 #(
		.INIT('h4)
	) name21709 (
		_w19263_,
		_w25755_,
		_w25756_
	);
	LUT2 #(
		.INIT('h1)
	) name21710 (
		_w22970_,
		_w23143_,
		_w25757_
	);
	LUT2 #(
		.INIT('h8)
	) name21711 (
		_w25748_,
		_w25757_,
		_w25758_
	);
	LUT2 #(
		.INIT('h4)
	) name21712 (
		_w19296_,
		_w25758_,
		_w25759_
	);
	LUT2 #(
		.INIT('h1)
	) name21713 (
		_w25751_,
		_w25759_,
		_w25760_
	);
	LUT2 #(
		.INIT('h4)
	) name21714 (
		_w25754_,
		_w25760_,
		_w25761_
	);
	LUT2 #(
		.INIT('h4)
	) name21715 (
		_w25756_,
		_w25761_,
		_w25762_
	);
	LUT2 #(
		.INIT('h4)
	) name21716 (
		_w25744_,
		_w25762_,
		_w25763_
	);
	LUT2 #(
		.INIT('h4)
	) name21717 (
		_w25747_,
		_w25763_,
		_w25764_
	);
	LUT2 #(
		.INIT('h1)
	) name21718 (
		_w19205_,
		_w25764_,
		_w25765_
	);
	LUT2 #(
		.INIT('h8)
	) name21719 (
		_w4137_,
		_w25743_,
		_w25766_
	);
	LUT2 #(
		.INIT('h2)
	) name21720 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w25755_,
		_w25767_
	);
	LUT2 #(
		.INIT('h1)
	) name21721 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w25753_,
		_w25768_
	);
	LUT2 #(
		.INIT('h1)
	) name21722 (
		_w25767_,
		_w25768_,
		_w25769_
	);
	LUT2 #(
		.INIT('h4)
	) name21723 (
		_w4137_,
		_w25746_,
		_w25770_
	);
	LUT2 #(
		.INIT('h4)
	) name21724 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w25750_,
		_w25771_
	);
	LUT2 #(
		.INIT('h8)
	) name21725 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w25758_,
		_w25772_
	);
	LUT2 #(
		.INIT('h1)
	) name21726 (
		_w25766_,
		_w25770_,
		_w25773_
	);
	LUT2 #(
		.INIT('h1)
	) name21727 (
		_w25771_,
		_w25772_,
		_w25774_
	);
	LUT2 #(
		.INIT('h8)
	) name21728 (
		_w25773_,
		_w25774_,
		_w25775_
	);
	LUT2 #(
		.INIT('h4)
	) name21729 (
		_w25769_,
		_w25775_,
		_w25776_
	);
	LUT2 #(
		.INIT('h2)
	) name21730 (
		_w19205_,
		_w25776_,
		_w25777_
	);
	LUT2 #(
		.INIT('h1)
	) name21731 (
		_w19315_,
		_w19337_,
		_w25778_
	);
	LUT2 #(
		.INIT('h8)
	) name21732 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w19315_,
		_w25779_
	);
	LUT2 #(
		.INIT('h1)
	) name21733 (
		_w25778_,
		_w25779_,
		_w25780_
	);
	LUT2 #(
		.INIT('h2)
	) name21734 (
		_w23143_,
		_w25780_,
		_w25781_
	);
	LUT2 #(
		.INIT('h4)
	) name21735 (
		_w23143_,
		_w25780_,
		_w25782_
	);
	LUT2 #(
		.INIT('h4)
	) name21736 (
		_w22970_,
		_w22981_,
		_w25783_
	);
	LUT2 #(
		.INIT('h4)
	) name21737 (
		_w23132_,
		_w25783_,
		_w25784_
	);
	LUT2 #(
		.INIT('h4)
	) name21738 (
		_w25781_,
		_w25784_,
		_w25785_
	);
	LUT2 #(
		.INIT('h4)
	) name21739 (
		_w25782_,
		_w25785_,
		_w25786_
	);
	LUT2 #(
		.INIT('h1)
	) name21740 (
		_w4117_,
		_w25777_,
		_w25787_
	);
	LUT2 #(
		.INIT('h4)
	) name21741 (
		_w25786_,
		_w25787_,
		_w25788_
	);
	LUT2 #(
		.INIT('h4)
	) name21742 (
		_w25765_,
		_w25788_,
		_w25789_
	);
	LUT2 #(
		.INIT('h4)
	) name21743 (
		\core_eu_ec_cun_termOK_CE_reg/P0001 ,
		_w4117_,
		_w25790_
	);
	LUT2 #(
		.INIT('h2)
	) name21744 (
		_w4149_,
		_w25790_,
		_w25791_
	);
	LUT2 #(
		.INIT('h4)
	) name21745 (
		_w25789_,
		_w25791_,
		_w25792_
	);
	LUT2 #(
		.INIT('h1)
	) name21746 (
		\T_PIOin[3]_pad ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w25793_
	);
	LUT2 #(
		.INIT('h8)
	) name21747 (
		\T_PIOin[3]_pad ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w25794_
	);
	LUT2 #(
		.INIT('h1)
	) name21748 (
		\pio_PIO_IN_P_reg[3]/P0001 ,
		_w25794_,
		_w25795_
	);
	LUT2 #(
		.INIT('h1)
	) name21749 (
		_w25793_,
		_w25795_,
		_w25796_
	);
	LUT2 #(
		.INIT('h1)
	) name21750 (
		\T_PIOin[1]_pad ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w25797_
	);
	LUT2 #(
		.INIT('h8)
	) name21751 (
		\T_PIOin[1]_pad ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w25798_
	);
	LUT2 #(
		.INIT('h1)
	) name21752 (
		\pio_PIO_IN_P_reg[1]/P0001 ,
		_w25798_,
		_w25799_
	);
	LUT2 #(
		.INIT('h1)
	) name21753 (
		_w25797_,
		_w25799_,
		_w25800_
	);
	LUT2 #(
		.INIT('h1)
	) name21754 (
		\T_PIOin[10]_pad ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w25801_
	);
	LUT2 #(
		.INIT('h8)
	) name21755 (
		\T_PIOin[10]_pad ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w25802_
	);
	LUT2 #(
		.INIT('h1)
	) name21756 (
		\pio_PIO_IN_P_reg[10]/P0001 ,
		_w25802_,
		_w25803_
	);
	LUT2 #(
		.INIT('h1)
	) name21757 (
		_w25801_,
		_w25803_,
		_w25804_
	);
	LUT2 #(
		.INIT('h1)
	) name21758 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w5950_,
		_w25805_
	);
	LUT2 #(
		.INIT('h4)
	) name21759 (
		\core_c_dec_Long_Cg_reg/P0001 ,
		_w5950_,
		_w25806_
	);
	LUT2 #(
		.INIT('h2)
	) name21760 (
		_w4116_,
		_w25805_,
		_w25807_
	);
	LUT2 #(
		.INIT('h4)
	) name21761 (
		_w25806_,
		_w25807_,
		_w25808_
	);
	LUT2 #(
		.INIT('h4)
	) name21762 (
		\auctl_T0Sack_reg/NET0131 ,
		_w4050_,
		_w25809_
	);
	LUT2 #(
		.INIT('h4)
	) name21763 (
		_w4097_,
		_w25809_,
		_w25810_
	);
	LUT2 #(
		.INIT('h4)
	) name21764 (
		\auctl_R1Sack_reg/NET0131 ,
		_w11772_,
		_w25811_
	);
	LUT2 #(
		.INIT('h1)
	) name21765 (
		\T_PIOin[8]_pad ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w25812_
	);
	LUT2 #(
		.INIT('h8)
	) name21766 (
		\T_PIOin[8]_pad ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w25813_
	);
	LUT2 #(
		.INIT('h1)
	) name21767 (
		\pio_PIO_IN_P_reg[8]/P0001 ,
		_w25813_,
		_w25814_
	);
	LUT2 #(
		.INIT('h1)
	) name21768 (
		_w25812_,
		_w25814_,
		_w25815_
	);
	LUT2 #(
		.INIT('h1)
	) name21769 (
		\T_PIOin[5]_pad ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w25816_
	);
	LUT2 #(
		.INIT('h8)
	) name21770 (
		\T_PIOin[5]_pad ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w25817_
	);
	LUT2 #(
		.INIT('h1)
	) name21771 (
		\pio_PIO_IN_P_reg[5]/P0001 ,
		_w25817_,
		_w25818_
	);
	LUT2 #(
		.INIT('h1)
	) name21772 (
		_w25816_,
		_w25818_,
		_w25819_
	);
	LUT2 #(
		.INIT('h1)
	) name21773 (
		\T_PIOin[6]_pad ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w25820_
	);
	LUT2 #(
		.INIT('h8)
	) name21774 (
		\T_PIOin[6]_pad ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w25821_
	);
	LUT2 #(
		.INIT('h1)
	) name21775 (
		\pio_PIO_IN_P_reg[6]/P0001 ,
		_w25821_,
		_w25822_
	);
	LUT2 #(
		.INIT('h1)
	) name21776 (
		_w25820_,
		_w25822_,
		_w25823_
	);
	LUT2 #(
		.INIT('h1)
	) name21777 (
		\T_PIOin[11]_pad ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w25824_
	);
	LUT2 #(
		.INIT('h8)
	) name21778 (
		\T_PIOin[11]_pad ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w25825_
	);
	LUT2 #(
		.INIT('h1)
	) name21779 (
		\pio_PIO_IN_P_reg[11]/P0001 ,
		_w25825_,
		_w25826_
	);
	LUT2 #(
		.INIT('h1)
	) name21780 (
		_w25824_,
		_w25826_,
		_w25827_
	);
	LUT2 #(
		.INIT('h4)
	) name21781 (
		\auctl_R0Sack_reg/NET0131 ,
		_w11774_,
		_w25828_
	);
	LUT2 #(
		.INIT('h4)
	) name21782 (
		\auctl_T1Sack_reg/NET0131 ,
		_w5968_,
		_w25829_
	);
	LUT2 #(
		.INIT('h4)
	) name21783 (
		_w4097_,
		_w25829_,
		_w25830_
	);
	LUT2 #(
		.INIT('h8)
	) name21784 (
		\tm_tcr_reg_DO_reg[15]/NET0131 ,
		_w20355_,
		_w25831_
	);
	LUT2 #(
		.INIT('h4)
	) name21785 (
		\tm_tpr_reg_DO_reg[15]/NET0131 ,
		_w22400_,
		_w25832_
	);
	LUT2 #(
		.INIT('h1)
	) name21786 (
		\tm_TCR_TMP_reg[11]/NET0131 ,
		_w22417_,
		_w25833_
	);
	LUT2 #(
		.INIT('h8)
	) name21787 (
		_w22424_,
		_w25833_,
		_w25834_
	);
	LUT2 #(
		.INIT('h8)
	) name21788 (
		\tm_TCR_TMP_reg[11]/NET0131 ,
		_w22417_,
		_w25835_
	);
	LUT2 #(
		.INIT('h4)
	) name21789 (
		_w22423_,
		_w25835_,
		_w25836_
	);
	LUT2 #(
		.INIT('h1)
	) name21790 (
		\T_TMODE[0]_pad ,
		_w25836_,
		_w25837_
	);
	LUT2 #(
		.INIT('h4)
	) name21791 (
		_w25834_,
		_w25837_,
		_w25838_
	);
	LUT2 #(
		.INIT('h2)
	) name21792 (
		_w22411_,
		_w25838_,
		_w25839_
	);
	LUT2 #(
		.INIT('h4)
	) name21793 (
		\tm_TCR_TMP_reg[12]/NET0131 ,
		_w25839_,
		_w25840_
	);
	LUT2 #(
		.INIT('h4)
	) name21794 (
		\tm_TCR_TMP_reg[13]/NET0131 ,
		_w25840_,
		_w25841_
	);
	LUT2 #(
		.INIT('h4)
	) name21795 (
		\tm_TCR_TMP_reg[14]/NET0131 ,
		_w25841_,
		_w25842_
	);
	LUT2 #(
		.INIT('h1)
	) name21796 (
		\tm_TCR_TMP_reg[15]/NET0131 ,
		_w25842_,
		_w25843_
	);
	LUT2 #(
		.INIT('h8)
	) name21797 (
		\tm_TCR_TMP_reg[15]/NET0131 ,
		_w25842_,
		_w25844_
	);
	LUT2 #(
		.INIT('h1)
	) name21798 (
		_w25843_,
		_w25844_,
		_w25845_
	);
	LUT2 #(
		.INIT('h1)
	) name21799 (
		_w22400_,
		_w25845_,
		_w25846_
	);
	LUT2 #(
		.INIT('h1)
	) name21800 (
		_w20355_,
		_w25832_,
		_w25847_
	);
	LUT2 #(
		.INIT('h4)
	) name21801 (
		_w25846_,
		_w25847_,
		_w25848_
	);
	LUT2 #(
		.INIT('h1)
	) name21802 (
		_w25831_,
		_w25848_,
		_w25849_
	);
	LUT2 #(
		.INIT('h4)
	) name21803 (
		\T_TMODE[1]_pad ,
		\core_c_dec_PPclr_reg/P0001 ,
		_w25850_
	);
	LUT2 #(
		.INIT('h8)
	) name21804 (
		\core_eu_ec_cun_COND_E_reg[2]/P0001 ,
		_w4117_,
		_w25851_
	);
	LUT2 #(
		.INIT('h2)
	) name21805 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w4117_,
		_w25852_
	);
	LUT2 #(
		.INIT('h1)
	) name21806 (
		_w25851_,
		_w25852_,
		_w25853_
	);
	LUT2 #(
		.INIT('h2)
	) name21807 (
		_w4150_,
		_w25853_,
		_w25854_
	);
	LUT2 #(
		.INIT('h1)
	) name21808 (
		\T_PIOin[4]_pad ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w25855_
	);
	LUT2 #(
		.INIT('h8)
	) name21809 (
		\T_PIOin[4]_pad ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w25856_
	);
	LUT2 #(
		.INIT('h1)
	) name21810 (
		\pio_PIO_IN_P_reg[4]/P0001 ,
		_w25856_,
		_w25857_
	);
	LUT2 #(
		.INIT('h1)
	) name21811 (
		_w25855_,
		_w25857_,
		_w25858_
	);
	LUT2 #(
		.INIT('h1)
	) name21812 (
		\T_PIOin[7]_pad ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w25859_
	);
	LUT2 #(
		.INIT('h8)
	) name21813 (
		\T_PIOin[7]_pad ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w25860_
	);
	LUT2 #(
		.INIT('h1)
	) name21814 (
		\pio_PIO_IN_P_reg[7]/P0001 ,
		_w25860_,
		_w25861_
	);
	LUT2 #(
		.INIT('h1)
	) name21815 (
		_w25859_,
		_w25861_,
		_w25862_
	);
	LUT2 #(
		.INIT('h8)
	) name21816 (
		\core_eu_ec_cun_COND_E_reg[3]/P0001 ,
		_w4117_,
		_w25863_
	);
	LUT2 #(
		.INIT('h2)
	) name21817 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w4117_,
		_w25864_
	);
	LUT2 #(
		.INIT('h1)
	) name21818 (
		_w25863_,
		_w25864_,
		_w25865_
	);
	LUT2 #(
		.INIT('h2)
	) name21819 (
		_w4150_,
		_w25865_,
		_w25866_
	);
	LUT2 #(
		.INIT('h1)
	) name21820 (
		\T_PIOin[9]_pad ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w25867_
	);
	LUT2 #(
		.INIT('h8)
	) name21821 (
		\T_PIOin[9]_pad ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w25868_
	);
	LUT2 #(
		.INIT('h1)
	) name21822 (
		\pio_PIO_IN_P_reg[9]/P0001 ,
		_w25868_,
		_w25869_
	);
	LUT2 #(
		.INIT('h1)
	) name21823 (
		_w25867_,
		_w25869_,
		_w25870_
	);
	LUT2 #(
		.INIT('h8)
	) name21824 (
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w21318_,
		_w25871_
	);
	LUT2 #(
		.INIT('h8)
	) name21825 (
		_w8715_,
		_w21316_,
		_w25872_
	);
	LUT2 #(
		.INIT('h4)
	) name21826 (
		_w18470_,
		_w18479_,
		_w25873_
	);
	LUT2 #(
		.INIT('h2)
	) name21827 (
		_w18470_,
		_w23047_,
		_w25874_
	);
	LUT2 #(
		.INIT('h4)
	) name21828 (
		_w18467_,
		_w18512_,
		_w25875_
	);
	LUT2 #(
		.INIT('h2)
	) name21829 (
		_w18471_,
		_w18479_,
		_w25876_
	);
	LUT2 #(
		.INIT('h8)
	) name21830 (
		_w18507_,
		_w25876_,
		_w25877_
	);
	LUT2 #(
		.INIT('h4)
	) name21831 (
		_w18500_,
		_w23051_,
		_w25878_
	);
	LUT2 #(
		.INIT('h1)
	) name21832 (
		_w18481_,
		_w25876_,
		_w25879_
	);
	LUT2 #(
		.INIT('h4)
	) name21833 (
		_w18492_,
		_w23052_,
		_w25880_
	);
	LUT2 #(
		.INIT('h8)
	) name21834 (
		_w23043_,
		_w23054_,
		_w25881_
	);
	LUT2 #(
		.INIT('h1)
	) name21835 (
		_w23061_,
		_w23150_,
		_w25882_
	);
	LUT2 #(
		.INIT('h4)
	) name21836 (
		_w23060_,
		_w23061_,
		_w25883_
	);
	LUT2 #(
		.INIT('h1)
	) name21837 (
		_w23054_,
		_w25882_,
		_w25884_
	);
	LUT2 #(
		.INIT('h4)
	) name21838 (
		_w25883_,
		_w25884_,
		_w25885_
	);
	LUT2 #(
		.INIT('h1)
	) name21839 (
		_w23052_,
		_w25881_,
		_w25886_
	);
	LUT2 #(
		.INIT('h4)
	) name21840 (
		_w25885_,
		_w25886_,
		_w25887_
	);
	LUT2 #(
		.INIT('h1)
	) name21841 (
		_w23051_,
		_w25880_,
		_w25888_
	);
	LUT2 #(
		.INIT('h4)
	) name21842 (
		_w25887_,
		_w25888_,
		_w25889_
	);
	LUT2 #(
		.INIT('h4)
	) name21843 (
		_w25878_,
		_w25879_,
		_w25890_
	);
	LUT2 #(
		.INIT('h4)
	) name21844 (
		_w25889_,
		_w25890_,
		_w25891_
	);
	LUT2 #(
		.INIT('h1)
	) name21845 (
		_w25875_,
		_w25877_,
		_w25892_
	);
	LUT2 #(
		.INIT('h4)
	) name21846 (
		_w25891_,
		_w25892_,
		_w25893_
	);
	LUT2 #(
		.INIT('h2)
	) name21847 (
		_w25874_,
		_w25893_,
		_w25894_
	);
	LUT2 #(
		.INIT('h2)
	) name21848 (
		_w23047_,
		_w23060_,
		_w25895_
	);
	LUT2 #(
		.INIT('h1)
	) name21849 (
		_w25873_,
		_w25895_,
		_w25896_
	);
	LUT2 #(
		.INIT('h4)
	) name21850 (
		_w25894_,
		_w25896_,
		_w25897_
	);
	LUT2 #(
		.INIT('h2)
	) name21851 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w25897_,
		_w25898_
	);
	LUT2 #(
		.INIT('h1)
	) name21852 (
		_w25871_,
		_w25872_,
		_w25899_
	);
	LUT2 #(
		.INIT('h4)
	) name21853 (
		_w25898_,
		_w25899_,
		_w25900_
	);
	LUT2 #(
		.INIT('h1)
	) name21854 (
		\T_PIOin[2]_pad ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w25901_
	);
	LUT2 #(
		.INIT('h8)
	) name21855 (
		\T_PIOin[2]_pad ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w25902_
	);
	LUT2 #(
		.INIT('h1)
	) name21856 (
		\pio_PIO_IN_P_reg[2]/P0001 ,
		_w25902_,
		_w25903_
	);
	LUT2 #(
		.INIT('h1)
	) name21857 (
		_w25901_,
		_w25903_,
		_w25904_
	);
	LUT2 #(
		.INIT('h8)
	) name21858 (
		\T_TMODE[1]_pad ,
		_w20206_,
		_w25905_
	);
	LUT2 #(
		.INIT('h8)
	) name21859 (
		\T_TMODE[1]_pad ,
		_w5518_,
		_w25906_
	);
	LUT2 #(
		.INIT('h8)
	) name21860 (
		_w5592_,
		_w25906_,
		_w25907_
	);
	LUT2 #(
		.INIT('h2)
	) name21861 (
		\emc_ECMcs_reg/NET0131 ,
		_w25907_,
		_w25908_
	);
	LUT2 #(
		.INIT('h1)
	) name21862 (
		_w25905_,
		_w25908_,
		_w25909_
	);
	LUT2 #(
		.INIT('h1)
	) name21863 (
		\T_PIOin[0]_pad ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w25910_
	);
	LUT2 #(
		.INIT('h8)
	) name21864 (
		\T_PIOin[0]_pad ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w25911_
	);
	LUT2 #(
		.INIT('h1)
	) name21865 (
		\pio_PIO_IN_P_reg[0]/P0001 ,
		_w25911_,
		_w25912_
	);
	LUT2 #(
		.INIT('h1)
	) name21866 (
		_w25910_,
		_w25912_,
		_w25913_
	);
	LUT2 #(
		.INIT('h8)
	) name21867 (
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		_w4094_,
		_w25914_
	);
	LUT2 #(
		.INIT('h2)
	) name21868 (
		\core_c_psq_Eqend_D_reg/P0001 ,
		_w4094_,
		_w25915_
	);
	LUT2 #(
		.INIT('h8)
	) name21869 (
		_w11741_,
		_w25915_,
		_w25916_
	);
	LUT2 #(
		.INIT('h1)
	) name21870 (
		_w25914_,
		_w25916_,
		_w25917_
	);
	LUT2 #(
		.INIT('h2)
	) name21871 (
		_w4116_,
		_w25917_,
		_w25918_
	);
	LUT2 #(
		.INIT('h8)
	) name21872 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		_w21318_,
		_w25919_
	);
	LUT2 #(
		.INIT('h4)
	) name21873 (
		_w18470_,
		_w18507_,
		_w25920_
	);
	LUT2 #(
		.INIT('h2)
	) name21874 (
		_w23047_,
		_w23162_,
		_w25921_
	);
	LUT2 #(
		.INIT('h4)
	) name21875 (
		_w18467_,
		_w18500_,
		_w25922_
	);
	LUT2 #(
		.INIT('h4)
	) name21876 (
		_w18492_,
		_w25876_,
		_w25923_
	);
	LUT2 #(
		.INIT('h8)
	) name21877 (
		_w23042_,
		_w23051_,
		_w25924_
	);
	LUT2 #(
		.INIT('h2)
	) name21878 (
		_w23052_,
		_w23059_,
		_w25925_
	);
	LUT2 #(
		.INIT('h8)
	) name21879 (
		_w23061_,
		_w23161_,
		_w25926_
	);
	LUT2 #(
		.INIT('h1)
	) name21880 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		_w18391_,
		_w25927_
	);
	LUT2 #(
		.INIT('h1)
	) name21881 (
		_w18392_,
		_w25927_,
		_w25928_
	);
	LUT2 #(
		.INIT('h4)
	) name21882 (
		_w23061_,
		_w25928_,
		_w25929_
	);
	LUT2 #(
		.INIT('h1)
	) name21883 (
		_w23054_,
		_w25926_,
		_w25930_
	);
	LUT2 #(
		.INIT('h4)
	) name21884 (
		_w25929_,
		_w25930_,
		_w25931_
	);
	LUT2 #(
		.INIT('h8)
	) name21885 (
		_w23054_,
		_w23149_,
		_w25932_
	);
	LUT2 #(
		.INIT('h1)
	) name21886 (
		_w23052_,
		_w25932_,
		_w25933_
	);
	LUT2 #(
		.INIT('h4)
	) name21887 (
		_w25931_,
		_w25933_,
		_w25934_
	);
	LUT2 #(
		.INIT('h1)
	) name21888 (
		_w23051_,
		_w25925_,
		_w25935_
	);
	LUT2 #(
		.INIT('h4)
	) name21889 (
		_w25934_,
		_w25935_,
		_w25936_
	);
	LUT2 #(
		.INIT('h2)
	) name21890 (
		_w18457_,
		_w25924_,
		_w25937_
	);
	LUT2 #(
		.INIT('h4)
	) name21891 (
		_w25936_,
		_w25937_,
		_w25938_
	);
	LUT2 #(
		.INIT('h2)
	) name21892 (
		_w25879_,
		_w25938_,
		_w25939_
	);
	LUT2 #(
		.INIT('h1)
	) name21893 (
		_w25922_,
		_w25923_,
		_w25940_
	);
	LUT2 #(
		.INIT('h4)
	) name21894 (
		_w25939_,
		_w25940_,
		_w25941_
	);
	LUT2 #(
		.INIT('h2)
	) name21895 (
		_w25874_,
		_w25941_,
		_w25942_
	);
	LUT2 #(
		.INIT('h1)
	) name21896 (
		_w25920_,
		_w25921_,
		_w25943_
	);
	LUT2 #(
		.INIT('h4)
	) name21897 (
		_w25942_,
		_w25943_,
		_w25944_
	);
	LUT2 #(
		.INIT('h2)
	) name21898 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w25944_,
		_w25945_
	);
	LUT2 #(
		.INIT('h8)
	) name21899 (
		_w7607_,
		_w21316_,
		_w25946_
	);
	LUT2 #(
		.INIT('h1)
	) name21900 (
		_w25919_,
		_w25946_,
		_w25947_
	);
	LUT2 #(
		.INIT('h4)
	) name21901 (
		_w25945_,
		_w25947_,
		_w25948_
	);
	LUT2 #(
		.INIT('h2)
	) name21902 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w25949_
	);
	LUT2 #(
		.INIT('h8)
	) name21903 (
		_w4115_,
		_w25949_,
		_w25950_
	);
	LUT2 #(
		.INIT('h2)
	) name21904 (
		PWDACK_pad,
		\clkc_Awake_reg/NET0131 ,
		_w25951_
	);
	LUT2 #(
		.INIT('h8)
	) name21905 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w25951_,
		_w25952_
	);
	LUT2 #(
		.INIT('h1)
	) name21906 (
		_w25950_,
		_w25952_,
		_w25953_
	);
	LUT2 #(
		.INIT('h8)
	) name21907 (
		\core_c_dec_MTLreg_E_reg[4]/P0001 ,
		_w5951_,
		_w25954_
	);
	LUT2 #(
		.INIT('h8)
	) name21908 (
		\core_c_dec_MTLreg_E_reg[5]/P0001 ,
		_w5951_,
		_w25955_
	);
	LUT2 #(
		.INIT('h8)
	) name21909 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w4117_,
		_w25956_
	);
	LUT2 #(
		.INIT('h4)
	) name21910 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w5888_,
		_w25957_
	);
	LUT2 #(
		.INIT('h1)
	) name21911 (
		_w25956_,
		_w25957_,
		_w25958_
	);
	LUT2 #(
		.INIT('h8)
	) name21912 (
		\core_c_dec_MTLreg_E_reg[7]/P0001 ,
		_w5951_,
		_w25959_
	);
	LUT2 #(
		.INIT('h4)
	) name21913 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w11736_,
		_w25960_
	);
	LUT2 #(
		.INIT('h1)
	) name21914 (
		_w13760_,
		_w25960_,
		_w25961_
	);
	LUT2 #(
		.INIT('h8)
	) name21915 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w25962_
	);
	LUT2 #(
		.INIT('h4)
	) name21916 (
		\sport1_txctl_SP_EN_D1_reg/P0001 ,
		_w25962_,
		_w25963_
	);
	LUT2 #(
		.INIT('h1)
	) name21917 (
		\sport1_txctl_TSreqi_reg/NET0131 ,
		_w25963_,
		_w25964_
	);
	LUT2 #(
		.INIT('h8)
	) name21918 (
		\core_c_dec_MTLreg_E_reg[6]/P0001 ,
		_w5951_,
		_w25965_
	);
	LUT2 #(
		.INIT('h8)
	) name21919 (
		\memc_usysr_DO_reg[12]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w25966_
	);
	LUT2 #(
		.INIT('h4)
	) name21920 (
		\sport0_txctl_SP_EN_D1_reg/P0001 ,
		_w25966_,
		_w25967_
	);
	LUT2 #(
		.INIT('h1)
	) name21921 (
		\sport0_txctl_TSreqi_reg/NET0131 ,
		_w25967_,
		_w25968_
	);
	LUT2 #(
		.INIT('h4)
	) name21922 (
		IACKn_pad,
		\sice_RCS_reg[0]/NET0131 ,
		_w25969_
	);
	LUT2 #(
		.INIT('h4)
	) name21923 (
		\sice_RCS_reg[1]/NET0131 ,
		_w25969_,
		_w25970_
	);
	LUT2 #(
		.INIT('h4)
	) name21924 (
		\sice_RCS_reg[0]/NET0131 ,
		\sice_RCS_reg[1]/NET0131 ,
		_w25971_
	);
	LUT2 #(
		.INIT('h1)
	) name21925 (
		_w25970_,
		_w25971_,
		_w25972_
	);
	LUT2 #(
		.INIT('h8)
	) name21926 (
		\core_c_dec_MTLreg_E_reg[2]/P0001 ,
		_w5951_,
		_w25973_
	);
	LUT2 #(
		.INIT('h8)
	) name21927 (
		\core_c_dec_MTLreg_E_reg[1]/P0001 ,
		_w5951_,
		_w25974_
	);
	LUT2 #(
		.INIT('h8)
	) name21928 (
		\core_c_dec_MTLreg_E_reg[0]/P0001 ,
		_w5951_,
		_w25975_
	);
	LUT2 #(
		.INIT('h8)
	) name21929 (
		\core_c_dec_MTLreg_E_reg[3]/P0001 ,
		_w5951_,
		_w25976_
	);
	LUT2 #(
		.INIT('h2)
	) name21930 (
		\core_c_psq_Iact_E_reg[10]/NET0131 ,
		_w19477_,
		_w25977_
	);
	LUT2 #(
		.INIT('h2)
	) name21931 (
		\core_c_psq_Iflag_reg[10]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w25978_
	);
	LUT2 #(
		.INIT('h8)
	) name21932 (
		_w19477_,
		_w25978_,
		_w25979_
	);
	LUT2 #(
		.INIT('h1)
	) name21933 (
		_w25977_,
		_w25979_,
		_w25980_
	);
	LUT2 #(
		.INIT('h8)
	) name21934 (
		\clkc_SLEEP_reg/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w25981_
	);
	LUT2 #(
		.INIT('h1)
	) name21935 (
		_w25950_,
		_w25981_,
		_w25982_
	);
	LUT2 #(
		.INIT('h1)
	) name21936 (
		_w13806_,
		_w14610_,
		_w25983_
	);
	LUT2 #(
		.INIT('h2)
	) name21937 (
		_w13806_,
		_w14586_,
		_w25984_
	);
	LUT2 #(
		.INIT('h1)
	) name21938 (
		_w25983_,
		_w25984_,
		_w25985_
	);
	LUT2 #(
		.INIT('h2)
	) name21939 (
		_w14667_,
		_w25985_,
		_w25986_
	);
	LUT2 #(
		.INIT('h2)
	) name21940 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[3]/P0001 ,
		_w14667_,
		_w25987_
	);
	LUT2 #(
		.INIT('h1)
	) name21941 (
		_w25986_,
		_w25987_,
		_w25988_
	);
	LUT2 #(
		.INIT('h2)
	) name21942 (
		\core_c_dec_MTICNTL_Eg_reg/P0001 ,
		_w5950_,
		_w25989_
	);
	LUT2 #(
		.INIT('h4)
	) name21943 (
		_w10069_,
		_w25989_,
		_w25990_
	);
	LUT2 #(
		.INIT('h1)
	) name21944 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w25989_,
		_w25991_
	);
	LUT2 #(
		.INIT('h1)
	) name21945 (
		_w25990_,
		_w25991_,
		_w25992_
	);
	LUT2 #(
		.INIT('h4)
	) name21946 (
		_w8715_,
		_w25989_,
		_w25993_
	);
	LUT2 #(
		.INIT('h1)
	) name21947 (
		\core_c_psq_ICNTL_reg_DO_reg[2]/NET0131 ,
		_w25989_,
		_w25994_
	);
	LUT2 #(
		.INIT('h1)
	) name21948 (
		_w25993_,
		_w25994_,
		_w25995_
	);
	LUT2 #(
		.INIT('h2)
	) name21949 (
		_w13805_,
		_w25985_,
		_w25996_
	);
	LUT2 #(
		.INIT('h2)
	) name21950 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[3]/P0001 ,
		_w13805_,
		_w25997_
	);
	LUT2 #(
		.INIT('h1)
	) name21951 (
		_w25996_,
		_w25997_,
		_w25998_
	);
	LUT2 #(
		.INIT('h8)
	) name21952 (
		\memc_STI_Cg_reg/NET0131 ,
		_w5950_,
		_w25999_
	);
	LUT2 #(
		.INIT('h1)
	) name21953 (
		_w5946_,
		_w13130_,
		_w26000_
	);
	LUT2 #(
		.INIT('h2)
	) name21954 (
		_w5951_,
		_w26000_,
		_w26001_
	);
	LUT2 #(
		.INIT('h1)
	) name21955 (
		_w25999_,
		_w26001_,
		_w26002_
	);
	LUT2 #(
		.INIT('h1)
	) name21956 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 ,
		_w19499_,
		_w26003_
	);
	LUT2 #(
		.INIT('h2)
	) name21957 (
		_w19499_,
		_w20259_,
		_w26004_
	);
	LUT2 #(
		.INIT('h2)
	) name21958 (
		_w19501_,
		_w26003_,
		_w26005_
	);
	LUT2 #(
		.INIT('h4)
	) name21959 (
		_w26004_,
		_w26005_,
		_w26006_
	);
	LUT2 #(
		.INIT('h2)
	) name21960 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[5]/P0001 ,
		_w19383_,
		_w26007_
	);
	LUT2 #(
		.INIT('h1)
	) name21961 (
		_w19508_,
		_w26007_,
		_w26008_
	);
	LUT2 #(
		.INIT('h4)
	) name21962 (
		_w26006_,
		_w26008_,
		_w26009_
	);
	LUT2 #(
		.INIT('h1)
	) name21963 (
		_w18262_,
		_w26009_,
		_w26010_
	);
	LUT2 #(
		.INIT('h1)
	) name21964 (
		_w17543_,
		_w19422_,
		_w26011_
	);
	LUT2 #(
		.INIT('h1)
	) name21965 (
		_w17676_,
		_w26011_,
		_w26012_
	);
	LUT2 #(
		.INIT('h1)
	) name21966 (
		_w17474_,
		_w17677_,
		_w26013_
	);
	LUT2 #(
		.INIT('h4)
	) name21967 (
		_w26012_,
		_w26013_,
		_w26014_
	);
	LUT2 #(
		.INIT('h2)
	) name21968 (
		_w26012_,
		_w26013_,
		_w26015_
	);
	LUT2 #(
		.INIT('h1)
	) name21969 (
		_w26014_,
		_w26015_,
		_w26016_
	);
	LUT2 #(
		.INIT('h4)
	) name21970 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w26016_,
		_w26017_
	);
	LUT2 #(
		.INIT('h8)
	) name21971 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w23218_,
		_w26018_
	);
	LUT2 #(
		.INIT('h1)
	) name21972 (
		_w26017_,
		_w26018_,
		_w26019_
	);
	LUT2 #(
		.INIT('h2)
	) name21973 (
		_w18262_,
		_w26019_,
		_w26020_
	);
	LUT2 #(
		.INIT('h1)
	) name21974 (
		_w26010_,
		_w26020_,
		_w26021_
	);
	LUT2 #(
		.INIT('h2)
	) name21975 (
		\tm_TSR_TMP_reg[6]/NET0131 ,
		_w25495_,
		_w26022_
	);
	LUT2 #(
		.INIT('h1)
	) name21976 (
		_w25496_,
		_w26022_,
		_w26023_
	);
	LUT2 #(
		.INIT('h2)
	) name21977 (
		_w25491_,
		_w26023_,
		_w26024_
	);
	LUT2 #(
		.INIT('h2)
	) name21978 (
		\tm_tsr_reg_DO_reg[6]/NET0131 ,
		_w25491_,
		_w26025_
	);
	LUT2 #(
		.INIT('h1)
	) name21979 (
		_w26024_,
		_w26025_,
		_w26026_
	);
	LUT2 #(
		.INIT('h2)
	) name21980 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w5950_,
		_w26027_
	);
	LUT2 #(
		.INIT('h4)
	) name21981 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w13565_,
		_w26028_
	);
	LUT2 #(
		.INIT('h1)
	) name21982 (
		_w26027_,
		_w26028_,
		_w26029_
	);
	LUT2 #(
		.INIT('h2)
	) name21983 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		\core_c_psq_TRAP_R_L_reg/NET0131 ,
		_w26030_
	);
	LUT2 #(
		.INIT('h8)
	) name21984 (
		\clkc_STBY_reg/NET0131 ,
		_w26030_,
		_w26031_
	);
	LUT2 #(
		.INIT('h1)
	) name21985 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w26032_
	);
	LUT2 #(
		.INIT('h8)
	) name21986 (
		_w4115_,
		_w26032_,
		_w26033_
	);
	LUT2 #(
		.INIT('h1)
	) name21987 (
		_w26031_,
		_w26033_,
		_w26034_
	);
	LUT2 #(
		.INIT('h8)
	) name21988 (
		_w14752_,
		_w26019_,
		_w26035_
	);
	LUT2 #(
		.INIT('h8)
	) name21989 (
		_w19776_,
		_w20259_,
		_w26036_
	);
	LUT2 #(
		.INIT('h2)
	) name21990 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[5]/P0001 ,
		_w17809_,
		_w26037_
	);
	LUT2 #(
		.INIT('h2)
	) name21991 (
		_w19780_,
		_w26037_,
		_w26038_
	);
	LUT2 #(
		.INIT('h4)
	) name21992 (
		_w26036_,
		_w26038_,
		_w26039_
	);
	LUT2 #(
		.INIT('h1)
	) name21993 (
		_w26035_,
		_w26039_,
		_w26040_
	);
	LUT2 #(
		.INIT('h1)
	) name21994 (
		\sice_IIRC_reg[0]/NET0131 ,
		\sice_IIRC_reg[1]/NET0131 ,
		_w26041_
	);
	LUT2 #(
		.INIT('h1)
	) name21995 (
		_w18865_,
		_w26041_,
		_w26042_
	);
	LUT2 #(
		.INIT('h1)
	) name21996 (
		\sice_ICYC_reg[0]/NET0131 ,
		\sice_ICYC_reg[1]/NET0131 ,
		_w26043_
	);
	LUT2 #(
		.INIT('h1)
	) name21997 (
		_w18856_,
		_w26043_,
		_w26044_
	);
	LUT2 #(
		.INIT('h1)
	) name21998 (
		\clkc_oscntr_reg_DO_reg[0]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[1]/NET0131 ,
		_w26045_
	);
	LUT2 #(
		.INIT('h1)
	) name21999 (
		_w20845_,
		_w26045_,
		_w26046_
	);
	LUT2 #(
		.INIT('h2)
	) name22000 (
		\core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001 ,
		_w20864_,
		_w26047_
	);
	LUT2 #(
		.INIT('h2)
	) name22001 (
		_w20864_,
		_w26019_,
		_w26048_
	);
	LUT2 #(
		.INIT('h1)
	) name22002 (
		_w26047_,
		_w26048_,
		_w26049_
	);
	LUT2 #(
		.INIT('h8)
	) name22003 (
		_w12743_,
		_w25097_,
		_w26050_
	);
	LUT2 #(
		.INIT('h8)
	) name22004 (
		_w19045_,
		_w25202_,
		_w26051_
	);
	LUT2 #(
		.INIT('h8)
	) name22005 (
		_w5524_,
		_w5575_,
		_w26052_
	);
	LUT2 #(
		.INIT('h8)
	) name22006 (
		_w12688_,
		_w25097_,
		_w26053_
	);
	LUT2 #(
		.INIT('h1)
	) name22007 (
		\clkc_SIDLE_s2_reg/NET0131 ,
		\clkc_STBY_reg/NET0131 ,
		_w26054_
	);
	LUT2 #(
		.INIT('h2)
	) name22008 (
		_w12241_,
		_w26054_,
		_w26055_
	);
	LUT2 #(
		.INIT('h2)
	) name22009 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001 ,
		_w20990_,
		_w26056_
	);
	LUT2 #(
		.INIT('h2)
	) name22010 (
		_w20990_,
		_w26019_,
		_w26057_
	);
	LUT2 #(
		.INIT('h1)
	) name22011 (
		_w26056_,
		_w26057_,
		_w26058_
	);
	LUT2 #(
		.INIT('h8)
	) name22012 (
		\core_c_dec_MTMreg_E_reg[6]/P0001 ,
		_w5951_,
		_w26059_
	);
	LUT2 #(
		.INIT('h8)
	) name22013 (
		\core_c_dec_MTMreg_E_reg[5]/P0001 ,
		_w5951_,
		_w26060_
	);
	LUT2 #(
		.INIT('h4)
	) name22014 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4098_,
		_w26061_
	);
	LUT2 #(
		.INIT('h4)
	) name22015 (
		\auctl_DSack_reg/NET0131 ,
		_w5068_,
		_w26062_
	);
	LUT2 #(
		.INIT('h4)
	) name22016 (
		_w26061_,
		_w26062_,
		_w26063_
	);
	LUT2 #(
		.INIT('h4)
	) name22017 (
		T_IMS_pad,
		\sice_ICS_reg[1]/NET0131 ,
		_w26064_
	);
	LUT2 #(
		.INIT('h4)
	) name22018 (
		\sice_ICS_reg[2]/NET0131 ,
		_w26064_,
		_w26065_
	);
	LUT2 #(
		.INIT('h8)
	) name22019 (
		_w7340_,
		_w25097_,
		_w26066_
	);
	LUT2 #(
		.INIT('h4)
	) name22020 (
		\auctl_BSack_reg/NET0131 ,
		_w5644_,
		_w26067_
	);
	LUT2 #(
		.INIT('h1)
	) name22021 (
		\auctl_DSack_reg/NET0131 ,
		\auctl_RST_reg/P0001 ,
		_w26068_
	);
	LUT2 #(
		.INIT('h8)
	) name22022 (
		\clkc_DSPoff_reg/NET0131 ,
		\clkc_SLEEP_reg/NET0131 ,
		_w26069_
	);
	LUT2 #(
		.INIT('h8)
	) name22023 (
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w26069_,
		_w26070_
	);
	LUT2 #(
		.INIT('h8)
	) name22024 (
		_w9178_,
		_w25097_,
		_w26071_
	);
	LUT2 #(
		.INIT('h8)
	) name22025 (
		\core_eu_ec_cun_mven_FFout_reg/NET0131 ,
		_w12245_,
		_w26072_
	);
	LUT2 #(
		.INIT('h2)
	) name22026 (
		_w4149_,
		_w26072_,
		_w26073_
	);
	LUT2 #(
		.INIT('h8)
	) name22027 (
		\core_c_dec_MTMreg_E_reg[7]/P0001 ,
		_w5951_,
		_w26074_
	);
	LUT2 #(
		.INIT('h8)
	) name22028 (
		\core_c_dec_MTMreg_E_reg[4]/P0001 ,
		_w5951_,
		_w26075_
	);
	LUT2 #(
		.INIT('h8)
	) name22029 (
		\core_c_dec_MTMreg_E_reg[1]/P0001 ,
		_w5951_,
		_w26076_
	);
	LUT2 #(
		.INIT('h8)
	) name22030 (
		\core_c_dec_MTMreg_E_reg[3]/P0001 ,
		_w5951_,
		_w26077_
	);
	LUT2 #(
		.INIT('h1)
	) name22031 (
		\auctl_BSack_reg/NET0131 ,
		\auctl_RST_reg/P0001 ,
		_w26078_
	);
	LUT2 #(
		.INIT('h8)
	) name22032 (
		\core_c_dec_MTMreg_E_reg[2]/P0001 ,
		_w5951_,
		_w26079_
	);
	LUT2 #(
		.INIT('h8)
	) name22033 (
		\core_c_dec_MTMreg_E_reg[0]/P0001 ,
		_w5951_,
		_w26080_
	);
	LUT2 #(
		.INIT('h1)
	) name22034 (
		\core_c_psq_PCS2or3_reg/NET0131 ,
		\core_c_psq_PCS_reg[4]/NET0131 ,
		_w26081_
	);
	LUT2 #(
		.INIT('h2)
	) name22035 (
		\auctl_STEAL_reg/NET0131 ,
		_w26081_,
		_w26082_
	);
	LUT2 #(
		.INIT('h4)
	) name22036 (
		\clkc_SIDLE_s1_reg/NET0131 ,
		\clkc_SIDLE_s2_reg/NET0131 ,
		_w26083_
	);
	LUT2 #(
		.INIT('h2)
	) name22037 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w26083_,
		_w26084_
	);
	LUT2 #(
		.INIT('h2)
	) name22038 (
		\bdma_RST_pin_reg/P0001 ,
		_w13733_,
		_w26085_
	);
	LUT2 #(
		.INIT('h8)
	) name22039 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w4117_,
		_w26086_
	);
	LUT2 #(
		.INIT('h1)
	) name22040 (
		_w25864_,
		_w26086_,
		_w26087_
	);
	LUT2 #(
		.INIT('h2)
	) name22041 (
		T_BMODE_pad,
		T_MMAP_pad,
		_w26088_
	);
	LUT2 #(
		.INIT('h2)
	) name22042 (
		\bdma_RST_pin_reg/P0001 ,
		_w26088_,
		_w26089_
	);
	LUT2 #(
		.INIT('h8)
	) name22043 (
		\bdma_RST_pin_reg/P0001 ,
		_w26088_,
		_w26090_
	);
	LUT2 #(
		.INIT('h8)
	) name22044 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w4117_,
		_w26091_
	);
	LUT2 #(
		.INIT('h1)
	) name22045 (
		_w25852_,
		_w26091_,
		_w26092_
	);
	LUT2 #(
		.INIT('h1)
	) name22046 (
		\bdma_BDMAmode_reg/NET0131 ,
		_w4116_,
		_w26093_
	);
	LUT2 #(
		.INIT('h2)
	) name22047 (
		_w4149_,
		_w26093_,
		_w26094_
	);
	LUT2 #(
		.INIT('h4)
	) name22048 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w4117_,
		_w26095_
	);
	LUT2 #(
		.INIT('h1)
	) name22049 (
		_w11742_,
		_w26095_,
		_w26096_
	);
	LUT2 #(
		.INIT('h4)
	) name22050 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		_w26097_
	);
	LUT2 #(
		.INIT('h8)
	) name22051 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		_w26098_
	);
	LUT2 #(
		.INIT('h1)
	) name22052 (
		_w26097_,
		_w26098_,
		_w26099_
	);
	LUT2 #(
		.INIT('h2)
	) name22053 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w4117_,
		_w26100_
	);
	LUT2 #(
		.INIT('h8)
	) name22054 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w4117_,
		_w26101_
	);
	LUT2 #(
		.INIT('h1)
	) name22055 (
		_w26100_,
		_w26101_,
		_w26102_
	);
	LUT2 #(
		.INIT('h8)
	) name22056 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w4117_,
		_w26103_
	);
	LUT2 #(
		.INIT('h1)
	) name22057 (
		_w25734_,
		_w26103_,
		_w26104_
	);
	LUT2 #(
		.INIT('h4)
	) name22058 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w26105_
	);
	LUT2 #(
		.INIT('h8)
	) name22059 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		_w26106_
	);
	LUT2 #(
		.INIT('h1)
	) name22060 (
		_w26105_,
		_w26106_,
		_w26107_
	);
	LUT2 #(
		.INIT('h4)
	) name22061 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w26108_
	);
	LUT2 #(
		.INIT('h8)
	) name22062 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		_w26109_
	);
	LUT2 #(
		.INIT('h1)
	) name22063 (
		_w26108_,
		_w26109_,
		_w26110_
	);
	LUT2 #(
		.INIT('h4)
	) name22064 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		_w26111_
	);
	LUT2 #(
		.INIT('h8)
	) name22065 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		_w26112_
	);
	LUT2 #(
		.INIT('h1)
	) name22066 (
		_w26111_,
		_w26112_,
		_w26113_
	);
	LUT2 #(
		.INIT('h4)
	) name22067 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w26114_
	);
	LUT2 #(
		.INIT('h8)
	) name22068 (
		\core_c_dec_accPM_E_reg/P0001 ,
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		_w26115_
	);
	LUT2 #(
		.INIT('h1)
	) name22069 (
		_w26114_,
		_w26115_,
		_w26116_
	);
	LUT2 #(
		.INIT('h1)
	) name22070 (
		\tm_tsr_reg_DO_reg[8]/NET0131 ,
		_w12245_,
		_w26117_
	);
	LUT2 #(
		.INIT('h2)
	) name22071 (
		\tm_tsr_reg_DO_reg[8]/NET0131 ,
		_w12241_,
		_w26118_
	);
	LUT2 #(
		.INIT('h1)
	) name22072 (
		_w26117_,
		_w26118_,
		_w26119_
	);
	LUT2 #(
		.INIT('h4)
	) name22073 (
		\clkc_DSPoff_reg/NET0131 ,
		\clkc_SLEEP_reg/NET0131 ,
		_w26120_
	);
	LUT2 #(
		.INIT('h4)
	) name22074 (
		\clkc_Cnt4096_reg/NET0131 ,
		\clkc_DSPoff_reg/NET0131 ,
		_w26121_
	);
	LUT2 #(
		.INIT('h1)
	) name22075 (
		_w26120_,
		_w26121_,
		_w26122_
	);
	LUT2 #(
		.INIT('h2)
	) name22076 (
		\sport1_txctl_TXSHT_reg[13]/P0001 ,
		_w22677_,
		_w26123_
	);
	LUT2 #(
		.INIT('h8)
	) name22077 (
		\sport1_txctl_TX_reg[14]/P0001 ,
		_w22677_,
		_w26124_
	);
	LUT2 #(
		.INIT('h1)
	) name22078 (
		_w26123_,
		_w26124_,
		_w26125_
	);
	LUT2 #(
		.INIT('h8)
	) name22079 (
		_w4094_,
		_w4116_,
		_w26126_
	);
	LUT2 #(
		.INIT('h1)
	) name22080 (
		_w5635_,
		_w26126_,
		_w26127_
	);
	LUT2 #(
		.INIT('h8)
	) name22081 (
		\core_c_psq_IFA_reg[12]/P0001 ,
		_w26126_,
		_w26128_
	);
	LUT2 #(
		.INIT('h1)
	) name22082 (
		_w26127_,
		_w26128_,
		_w26129_
	);
	LUT2 #(
		.INIT('h1)
	) name22083 (
		_w5419_,
		_w26126_,
		_w26130_
	);
	LUT2 #(
		.INIT('h8)
	) name22084 (
		\core_c_psq_IFA_reg[9]/P0001 ,
		_w26126_,
		_w26131_
	);
	LUT2 #(
		.INIT('h1)
	) name22085 (
		_w26130_,
		_w26131_,
		_w26132_
	);
	LUT2 #(
		.INIT('h1)
	) name22086 (
		_w5338_,
		_w26126_,
		_w26133_
	);
	LUT2 #(
		.INIT('h8)
	) name22087 (
		\core_c_psq_IFA_reg[6]/P0001 ,
		_w26126_,
		_w26134_
	);
	LUT2 #(
		.INIT('h1)
	) name22088 (
		_w26133_,
		_w26134_,
		_w26135_
	);
	LUT2 #(
		.INIT('h1)
	) name22089 (
		_w5311_,
		_w26126_,
		_w26136_
	);
	LUT2 #(
		.INIT('h8)
	) name22090 (
		\core_c_psq_IFA_reg[5]/P0001 ,
		_w26126_,
		_w26137_
	);
	LUT2 #(
		.INIT('h1)
	) name22091 (
		_w26136_,
		_w26137_,
		_w26138_
	);
	LUT2 #(
		.INIT('h1)
	) name22092 (
		_w5208_,
		_w26126_,
		_w26139_
	);
	LUT2 #(
		.INIT('h8)
	) name22093 (
		\core_c_psq_IFA_reg[2]/P0001 ,
		_w26126_,
		_w26140_
	);
	LUT2 #(
		.INIT('h1)
	) name22094 (
		_w26139_,
		_w26140_,
		_w26141_
	);
	LUT2 #(
		.INIT('h1)
	) name22095 (
		_w5169_,
		_w26126_,
		_w26142_
	);
	LUT2 #(
		.INIT('h8)
	) name22096 (
		\core_c_psq_IFA_reg[1]/P0001 ,
		_w26126_,
		_w26143_
	);
	LUT2 #(
		.INIT('h1)
	) name22097 (
		_w26142_,
		_w26143_,
		_w26144_
	);
	LUT2 #(
		.INIT('h1)
	) name22098 (
		_w5142_,
		_w26126_,
		_w26145_
	);
	LUT2 #(
		.INIT('h8)
	) name22099 (
		\core_c_psq_IFA_reg[11]/P0001 ,
		_w26126_,
		_w26146_
	);
	LUT2 #(
		.INIT('h1)
	) name22100 (
		_w26145_,
		_w26146_,
		_w26147_
	);
	LUT2 #(
		.INIT('h1)
	) name22101 (
		_w5064_,
		_w26126_,
		_w26148_
	);
	LUT2 #(
		.INIT('h8)
	) name22102 (
		\core_c_psq_IFA_reg[0]/P0001 ,
		_w26126_,
		_w26149_
	);
	LUT2 #(
		.INIT('h1)
	) name22103 (
		_w26148_,
		_w26149_,
		_w26150_
	);
	LUT2 #(
		.INIT('h2)
	) name22104 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		_w4094_,
		_w26151_
	);
	LUT2 #(
		.INIT('h8)
	) name22105 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		_w4094_,
		_w26152_
	);
	LUT2 #(
		.INIT('h1)
	) name22106 (
		_w26151_,
		_w26152_,
		_w26153_
	);
	LUT2 #(
		.INIT('h2)
	) name22107 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		_w4094_,
		_w26154_
	);
	LUT2 #(
		.INIT('h8)
	) name22108 (
		\core_c_psq_EXA_reg[6]/P0001 ,
		_w4094_,
		_w26155_
	);
	LUT2 #(
		.INIT('h1)
	) name22109 (
		_w26154_,
		_w26155_,
		_w26156_
	);
	LUT2 #(
		.INIT('h2)
	) name22110 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		_w4094_,
		_w26157_
	);
	LUT2 #(
		.INIT('h8)
	) name22111 (
		\core_c_psq_EXA_reg[3]/P0001 ,
		_w4094_,
		_w26158_
	);
	LUT2 #(
		.INIT('h1)
	) name22112 (
		_w26157_,
		_w26158_,
		_w26159_
	);
	LUT2 #(
		.INIT('h2)
	) name22113 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		_w4094_,
		_w26160_
	);
	LUT2 #(
		.INIT('h8)
	) name22114 (
		\core_c_psq_EXA_reg[2]/P0001 ,
		_w4094_,
		_w26161_
	);
	LUT2 #(
		.INIT('h1)
	) name22115 (
		_w26160_,
		_w26161_,
		_w26162_
	);
	LUT2 #(
		.INIT('h2)
	) name22116 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		_w4094_,
		_w26163_
	);
	LUT2 #(
		.INIT('h8)
	) name22117 (
		\core_c_psq_EXA_reg[13]/P0001 ,
		_w4094_,
		_w26164_
	);
	LUT2 #(
		.INIT('h1)
	) name22118 (
		_w26163_,
		_w26164_,
		_w26165_
	);
	LUT2 #(
		.INIT('h2)
	) name22119 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		_w4094_,
		_w26166_
	);
	LUT2 #(
		.INIT('h8)
	) name22120 (
		\core_c_psq_EXA_reg[12]/P0001 ,
		_w4094_,
		_w26167_
	);
	LUT2 #(
		.INIT('h1)
	) name22121 (
		_w26166_,
		_w26167_,
		_w26168_
	);
	LUT2 #(
		.INIT('h8)
	) name22122 (
		\core_c_dec_accCM_E_reg/NET0131 ,
		_w4117_,
		_w26169_
	);
	LUT2 #(
		.INIT('h1)
	) name22123 (
		_w5888_,
		_w26169_,
		_w26170_
	);
	LUT2 #(
		.INIT('h1)
	) name22124 (
		_w5245_,
		_w26126_,
		_w26171_
	);
	LUT2 #(
		.INIT('h8)
	) name22125 (
		\core_c_psq_IFA_reg[3]/P0001 ,
		_w26126_,
		_w26172_
	);
	LUT2 #(
		.INIT('h1)
	) name22126 (
		_w26171_,
		_w26172_,
		_w26173_
	);
	LUT2 #(
		.INIT('h2)
	) name22127 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		_w4094_,
		_w26174_
	);
	LUT2 #(
		.INIT('h8)
	) name22128 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		_w4094_,
		_w26175_
	);
	LUT2 #(
		.INIT('h1)
	) name22129 (
		_w26174_,
		_w26175_,
		_w26176_
	);
	LUT2 #(
		.INIT('h2)
	) name22130 (
		_w4829_,
		_w5950_,
		_w26177_
	);
	LUT2 #(
		.INIT('h8)
	) name22131 (
		\core_c_dec_Prderr_Cg_reg/NET0131 ,
		_w5950_,
		_w26178_
	);
	LUT2 #(
		.INIT('h1)
	) name22132 (
		_w26177_,
		_w26178_,
		_w26179_
	);
	LUT2 #(
		.INIT('h2)
	) name22133 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		_w4094_,
		_w26180_
	);
	LUT2 #(
		.INIT('h8)
	) name22134 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		_w4094_,
		_w26181_
	);
	LUT2 #(
		.INIT('h1)
	) name22135 (
		_w26180_,
		_w26181_,
		_w26182_
	);
	LUT2 #(
		.INIT('h2)
	) name22136 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		_w4117_,
		_w26183_
	);
	LUT2 #(
		.INIT('h8)
	) name22137 (
		\core_c_dec_IRE_reg[18]/NET0131 ,
		_w4117_,
		_w26184_
	);
	LUT2 #(
		.INIT('h1)
	) name22138 (
		_w26183_,
		_w26184_,
		_w26185_
	);
	LUT2 #(
		.INIT('h2)
	) name22139 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w4117_,
		_w26186_
	);
	LUT2 #(
		.INIT('h8)
	) name22140 (
		\core_c_dec_IRE_reg[19]/NET0131 ,
		_w4117_,
		_w26187_
	);
	LUT2 #(
		.INIT('h1)
	) name22141 (
		_w26186_,
		_w26187_,
		_w26188_
	);
	LUT2 #(
		.INIT('h1)
	) name22142 (
		_w5365_,
		_w26126_,
		_w26189_
	);
	LUT2 #(
		.INIT('h8)
	) name22143 (
		\core_c_psq_IFA_reg[7]/P0001 ,
		_w26126_,
		_w26190_
	);
	LUT2 #(
		.INIT('h1)
	) name22144 (
		_w26189_,
		_w26190_,
		_w26191_
	);
	LUT2 #(
		.INIT('h2)
	) name22145 (
		\sport1_txctl_TXSHT_reg[14]/P0001 ,
		_w22677_,
		_w26192_
	);
	LUT2 #(
		.INIT('h8)
	) name22146 (
		\sport1_txctl_TX_reg[15]/P0001 ,
		_w22677_,
		_w26193_
	);
	LUT2 #(
		.INIT('h1)
	) name22147 (
		_w26192_,
		_w26193_,
		_w26194_
	);
	LUT2 #(
		.INIT('h1)
	) name22148 (
		_w4117_,
		_w6033_,
		_w26195_
	);
	LUT2 #(
		.INIT('h8)
	) name22149 (
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w4117_,
		_w26196_
	);
	LUT2 #(
		.INIT('h1)
	) name22150 (
		_w26195_,
		_w26196_,
		_w26197_
	);
	LUT2 #(
		.INIT('h1)
	) name22151 (
		_w4117_,
		_w6036_,
		_w26198_
	);
	LUT2 #(
		.INIT('h8)
	) name22152 (
		\core_dag_ilm2reg_IL_E_reg[0]/P0001 ,
		_w4117_,
		_w26199_
	);
	LUT2 #(
		.INIT('h1)
	) name22153 (
		_w26198_,
		_w26199_,
		_w26200_
	);
	LUT2 #(
		.INIT('h2)
	) name22154 (
		_w4099_,
		_w5981_,
		_w26201_
	);
	LUT2 #(
		.INIT('h2)
	) name22155 (
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w4099_,
		_w26202_
	);
	LUT2 #(
		.INIT('h1)
	) name22156 (
		_w26201_,
		_w26202_,
		_w26203_
	);
	LUT2 #(
		.INIT('h2)
	) name22157 (
		_w4099_,
		_w5974_,
		_w26204_
	);
	LUT2 #(
		.INIT('h2)
	) name22158 (
		\core_dag_ilm1reg_STEALI_E_reg[1]/P0001 ,
		_w4099_,
		_w26205_
	);
	LUT2 #(
		.INIT('h1)
	) name22159 (
		_w26204_,
		_w26205_,
		_w26206_
	);
	LUT2 #(
		.INIT('h2)
	) name22160 (
		_w4099_,
		_w5989_,
		_w26207_
	);
	LUT2 #(
		.INIT('h2)
	) name22161 (
		\core_dag_ilm1reg_STEALI_E_reg[0]/P0001 ,
		_w4099_,
		_w26208_
	);
	LUT2 #(
		.INIT('h1)
	) name22162 (
		_w26207_,
		_w26208_,
		_w26209_
	);
	LUT2 #(
		.INIT('h2)
	) name22163 (
		\sport1_txctl_TXSHT_reg[12]/P0001 ,
		_w22677_,
		_w26210_
	);
	LUT2 #(
		.INIT('h8)
	) name22164 (
		\sport1_txctl_TX_reg[13]/P0001 ,
		_w22677_,
		_w26211_
	);
	LUT2 #(
		.INIT('h1)
	) name22165 (
		_w26210_,
		_w26211_,
		_w26212_
	);
	LUT2 #(
		.INIT('h2)
	) name22166 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		_w4094_,
		_w26213_
	);
	LUT2 #(
		.INIT('h8)
	) name22167 (
		\core_c_psq_EXA_reg[1]/P0001 ,
		_w4094_,
		_w26214_
	);
	LUT2 #(
		.INIT('h1)
	) name22168 (
		_w26213_,
		_w26214_,
		_w26215_
	);
	LUT2 #(
		.INIT('h2)
	) name22169 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		_w4094_,
		_w26216_
	);
	LUT2 #(
		.INIT('h8)
	) name22170 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		_w4094_,
		_w26217_
	);
	LUT2 #(
		.INIT('h1)
	) name22171 (
		_w26216_,
		_w26217_,
		_w26218_
	);
	LUT2 #(
		.INIT('h2)
	) name22172 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		_w4094_,
		_w26219_
	);
	LUT2 #(
		.INIT('h8)
	) name22173 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		_w4094_,
		_w26220_
	);
	LUT2 #(
		.INIT('h1)
	) name22174 (
		_w26219_,
		_w26220_,
		_w26221_
	);
	LUT2 #(
		.INIT('h2)
	) name22175 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		_w4094_,
		_w26222_
	);
	LUT2 #(
		.INIT('h8)
	) name22176 (
		\core_c_psq_EXA_reg[5]/P0001 ,
		_w4094_,
		_w26223_
	);
	LUT2 #(
		.INIT('h1)
	) name22177 (
		_w26222_,
		_w26223_,
		_w26224_
	);
	LUT2 #(
		.INIT('h2)
	) name22178 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		_w4094_,
		_w26225_
	);
	LUT2 #(
		.INIT('h8)
	) name22179 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		_w4094_,
		_w26226_
	);
	LUT2 #(
		.INIT('h1)
	) name22180 (
		_w26225_,
		_w26226_,
		_w26227_
	);
	LUT2 #(
		.INIT('h2)
	) name22181 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		_w4094_,
		_w26228_
	);
	LUT2 #(
		.INIT('h8)
	) name22182 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		_w4094_,
		_w26229_
	);
	LUT2 #(
		.INIT('h1)
	) name22183 (
		_w26228_,
		_w26229_,
		_w26230_
	);
	LUT2 #(
		.INIT('h1)
	) name22184 (
		_w5113_,
		_w26126_,
		_w26231_
	);
	LUT2 #(
		.INIT('h8)
	) name22185 (
		\core_c_psq_IFA_reg[10]/P0001 ,
		_w26126_,
		_w26232_
	);
	LUT2 #(
		.INIT('h1)
	) name22186 (
		_w26231_,
		_w26232_,
		_w26233_
	);
	LUT2 #(
		.INIT('h1)
	) name22187 (
		_w5660_,
		_w26126_,
		_w26234_
	);
	LUT2 #(
		.INIT('h8)
	) name22188 (
		\core_c_psq_IFA_reg[13]/P0001 ,
		_w26126_,
		_w26235_
	);
	LUT2 #(
		.INIT('h1)
	) name22189 (
		_w26234_,
		_w26235_,
		_w26236_
	);
	LUT2 #(
		.INIT('h1)
	) name22190 (
		_w5279_,
		_w26126_,
		_w26237_
	);
	LUT2 #(
		.INIT('h8)
	) name22191 (
		\core_c_psq_IFA_reg[4]/P0001 ,
		_w26126_,
		_w26238_
	);
	LUT2 #(
		.INIT('h1)
	) name22192 (
		_w26237_,
		_w26238_,
		_w26239_
	);
	LUT2 #(
		.INIT('h1)
	) name22193 (
		_w5392_,
		_w26126_,
		_w26240_
	);
	LUT2 #(
		.INIT('h8)
	) name22194 (
		\core_c_psq_IFA_reg[8]/P0001 ,
		_w26126_,
		_w26241_
	);
	LUT2 #(
		.INIT('h1)
	) name22195 (
		_w26240_,
		_w26241_,
		_w26242_
	);
	LUT2 #(
		.INIT('h4)
	) name22196 (
		\sport0_rxctl_RXSHT_reg[1]/P0001 ,
		_w20868_,
		_w26243_
	);
	LUT2 #(
		.INIT('h8)
	) name22197 (
		\sport0_rxctl_RX_reg[1]/P0001 ,
		_w20873_,
		_w26244_
	);
	LUT2 #(
		.INIT('h4)
	) name22198 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w9435_,
		_w26245_
	);
	LUT2 #(
		.INIT('h1)
	) name22199 (
		_w20938_,
		_w20943_,
		_w26246_
	);
	LUT2 #(
		.INIT('h1)
	) name22200 (
		_w20880_,
		_w26246_,
		_w26247_
	);
	LUT2 #(
		.INIT('h1)
	) name22201 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w20953_,
		_w26248_
	);
	LUT2 #(
		.INIT('h2)
	) name22202 (
		_w26247_,
		_w26248_,
		_w26249_
	);
	LUT2 #(
		.INIT('h4)
	) name22203 (
		_w26247_,
		_w26248_,
		_w26250_
	);
	LUT2 #(
		.INIT('h2)
	) name22204 (
		_w20875_,
		_w26249_,
		_w26251_
	);
	LUT2 #(
		.INIT('h4)
	) name22205 (
		_w26250_,
		_w26251_,
		_w26252_
	);
	LUT2 #(
		.INIT('h1)
	) name22206 (
		_w20868_,
		_w26244_,
		_w26253_
	);
	LUT2 #(
		.INIT('h4)
	) name22207 (
		_w26252_,
		_w26253_,
		_w26254_
	);
	LUT2 #(
		.INIT('h4)
	) name22208 (
		_w26245_,
		_w26254_,
		_w26255_
	);
	LUT2 #(
		.INIT('h1)
	) name22209 (
		_w20871_,
		_w26243_,
		_w26256_
	);
	LUT2 #(
		.INIT('h4)
	) name22210 (
		_w26255_,
		_w26256_,
		_w26257_
	);
	LUT2 #(
		.INIT('h8)
	) name22211 (
		\sport0_rxctl_RX_reg[1]/P0001 ,
		_w20871_,
		_w26258_
	);
	LUT2 #(
		.INIT('h1)
	) name22212 (
		_w26257_,
		_w26258_,
		_w26259_
	);
	LUT2 #(
		.INIT('h2)
	) name22213 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w18974_,
		_w26260_
	);
	LUT2 #(
		.INIT('h4)
	) name22214 (
		_w23630_,
		_w23634_,
		_w26261_
	);
	LUT2 #(
		.INIT('h2)
	) name22215 (
		_w23620_,
		_w23625_,
		_w26262_
	);
	LUT2 #(
		.INIT('h8)
	) name22216 (
		_w23604_,
		_w23607_,
		_w26263_
	);
	LUT2 #(
		.INIT('h8)
	) name22217 (
		_w23610_,
		_w23613_,
		_w26264_
	);
	LUT2 #(
		.INIT('h8)
	) name22218 (
		_w23585_,
		_w26263_,
		_w26265_
	);
	LUT2 #(
		.INIT('h4)
	) name22219 (
		_w26264_,
		_w26265_,
		_w26266_
	);
	LUT2 #(
		.INIT('h2)
	) name22220 (
		_w26262_,
		_w26266_,
		_w26267_
	);
	LUT2 #(
		.INIT('h2)
	) name22221 (
		_w26261_,
		_w26267_,
		_w26268_
	);
	LUT2 #(
		.INIT('h8)
	) name22222 (
		_w23638_,
		_w23642_,
		_w26269_
	);
	LUT2 #(
		.INIT('h4)
	) name22223 (
		_w26268_,
		_w26269_,
		_w26270_
	);
	LUT2 #(
		.INIT('h8)
	) name22224 (
		_w23646_,
		_w23650_,
		_w26271_
	);
	LUT2 #(
		.INIT('h4)
	) name22225 (
		_w26270_,
		_w26271_,
		_w26272_
	);
	LUT2 #(
		.INIT('h8)
	) name22226 (
		_w23654_,
		_w23658_,
		_w26273_
	);
	LUT2 #(
		.INIT('h4)
	) name22227 (
		_w26272_,
		_w26273_,
		_w26274_
	);
	LUT2 #(
		.INIT('h8)
	) name22228 (
		_w23662_,
		_w23670_,
		_w26275_
	);
	LUT2 #(
		.INIT('h4)
	) name22229 (
		_w26274_,
		_w26275_,
		_w26276_
	);
	LUT2 #(
		.INIT('h1)
	) name22230 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w26276_,
		_w26277_
	);
	LUT2 #(
		.INIT('h1)
	) name22231 (
		_w26260_,
		_w26277_,
		_w26278_
	);
	LUT2 #(
		.INIT('h2)
	) name22232 (
		_w23677_,
		_w26278_,
		_w26279_
	);
	LUT2 #(
		.INIT('h1)
	) name22233 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[1]/P0001 ,
		_w23677_,
		_w26280_
	);
	LUT2 #(
		.INIT('h1)
	) name22234 (
		_w26279_,
		_w26280_,
		_w26281_
	);
	LUT2 #(
		.INIT('h2)
	) name22235 (
		_w23598_,
		_w26278_,
		_w26282_
	);
	LUT2 #(
		.INIT('h1)
	) name22236 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[1]/P0001 ,
		_w23598_,
		_w26283_
	);
	LUT2 #(
		.INIT('h1)
	) name22237 (
		_w26282_,
		_w26283_,
		_w26284_
	);
	LUT2 #(
		.INIT('h4)
	) name22238 (
		\clkc_CTR_cnt_reg[0]/NET0131 ,
		\clkc_CTR_cnt_reg[1]/NET0131 ,
		_w26285_
	);
	LUT2 #(
		.INIT('h1)
	) name22239 (
		_w24968_,
		_w26285_,
		_w26286_
	);
	LUT2 #(
		.INIT('h1)
	) name22240 (
		\auctl_R0Sack_reg/NET0131 ,
		\auctl_RST_reg/P0001 ,
		_w26287_
	);
	LUT2 #(
		.INIT('h1)
	) name22241 (
		\auctl_RST_reg/P0001 ,
		\auctl_T0Sack_reg/NET0131 ,
		_w26288_
	);
	LUT2 #(
		.INIT('h1)
	) name22242 (
		\auctl_R1Sack_reg/NET0131 ,
		\auctl_RST_reg/P0001 ,
		_w26289_
	);
	LUT2 #(
		.INIT('h8)
	) name22243 (
		\sice_ICYC_en_syn_reg/P0001 ,
		_w12245_,
		_w26290_
	);
	LUT2 #(
		.INIT('h1)
	) name22244 (
		\auctl_RST_reg/P0001 ,
		\auctl_T1Sack_reg/NET0131 ,
		_w26291_
	);
	LUT2 #(
		.INIT('h8)
	) name22245 (
		_w4116_,
		_w4149_,
		_w26292_
	);
	LUT2 #(
		.INIT('h8)
	) name22246 (
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		_w26293_
	);
	LUT2 #(
		.INIT('h1)
	) name22247 (
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[1]/NET0131 ,
		_w26294_
	);
	LUT2 #(
		.INIT('h2)
	) name22248 (
		T_IMS_pad,
		_w26293_,
		_w26295_
	);
	LUT2 #(
		.INIT('h4)
	) name22249 (
		_w26294_,
		_w26295_,
		_w26296_
	);
	LUT2 #(
		.INIT('h2)
	) name22250 (
		\sice_ICS_reg[2]/NET0131 ,
		_w26296_,
		_w26297_
	);
	LUT2 #(
		.INIT('h2)
	) name22251 (
		\sice_ICS_reg[0]/NET0131 ,
		\sice_ICS_reg[2]/NET0131 ,
		_w26298_
	);
	LUT2 #(
		.INIT('h1)
	) name22252 (
		_w23030_,
		_w26064_,
		_w26299_
	);
	LUT2 #(
		.INIT('h8)
	) name22253 (
		_w26298_,
		_w26299_,
		_w26300_
	);
	LUT2 #(
		.INIT('h1)
	) name22254 (
		_w26297_,
		_w26300_,
		_w26301_
	);
	LUT2 #(
		.INIT('h2)
	) name22255 (
		_w12234_,
		_w26301_,
		_w26302_
	);
	LUT2 #(
		.INIT('h1)
	) name22256 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 ,
		_w19499_,
		_w26303_
	);
	LUT2 #(
		.INIT('h2)
	) name22257 (
		_w19499_,
		_w20080_,
		_w26304_
	);
	LUT2 #(
		.INIT('h2)
	) name22258 (
		_w19501_,
		_w26303_,
		_w26305_
	);
	LUT2 #(
		.INIT('h4)
	) name22259 (
		_w26304_,
		_w26305_,
		_w26306_
	);
	LUT2 #(
		.INIT('h2)
	) name22260 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[4]/P0001 ,
		_w19383_,
		_w26307_
	);
	LUT2 #(
		.INIT('h1)
	) name22261 (
		_w19508_,
		_w26307_,
		_w26308_
	);
	LUT2 #(
		.INIT('h4)
	) name22262 (
		_w26306_,
		_w26308_,
		_w26309_
	);
	LUT2 #(
		.INIT('h1)
	) name22263 (
		_w18262_,
		_w26309_,
		_w26310_
	);
	LUT2 #(
		.INIT('h8)
	) name22264 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w26016_,
		_w26311_
	);
	LUT2 #(
		.INIT('h1)
	) name22265 (
		_w17543_,
		_w17676_,
		_w26312_
	);
	LUT2 #(
		.INIT('h2)
	) name22266 (
		_w19422_,
		_w26312_,
		_w26313_
	);
	LUT2 #(
		.INIT('h4)
	) name22267 (
		_w19422_,
		_w26312_,
		_w26314_
	);
	LUT2 #(
		.INIT('h1)
	) name22268 (
		_w26313_,
		_w26314_,
		_w26315_
	);
	LUT2 #(
		.INIT('h4)
	) name22269 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w26315_,
		_w26316_
	);
	LUT2 #(
		.INIT('h1)
	) name22270 (
		_w26311_,
		_w26316_,
		_w26317_
	);
	LUT2 #(
		.INIT('h2)
	) name22271 (
		_w18262_,
		_w26317_,
		_w26318_
	);
	LUT2 #(
		.INIT('h1)
	) name22272 (
		_w26310_,
		_w26318_,
		_w26319_
	);
	LUT2 #(
		.INIT('h4)
	) name22273 (
		\clkc_ckr_reg_DO_reg[15]/NET0131 ,
		_w12245_,
		_w26320_
	);
	LUT2 #(
		.INIT('h8)
	) name22274 (
		_w14752_,
		_w26317_,
		_w26321_
	);
	LUT2 #(
		.INIT('h8)
	) name22275 (
		_w19776_,
		_w20080_,
		_w26322_
	);
	LUT2 #(
		.INIT('h2)
	) name22276 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[4]/P0001 ,
		_w17809_,
		_w26323_
	);
	LUT2 #(
		.INIT('h2)
	) name22277 (
		_w19780_,
		_w26323_,
		_w26324_
	);
	LUT2 #(
		.INIT('h4)
	) name22278 (
		_w26322_,
		_w26324_,
		_w26325_
	);
	LUT2 #(
		.INIT('h1)
	) name22279 (
		_w26321_,
		_w26325_,
		_w26326_
	);
	LUT2 #(
		.INIT('h1)
	) name22280 (
		T_ISn_pad,
		T_IWRn_pad,
		_w26327_
	);
	LUT2 #(
		.INIT('h4)
	) name22281 (
		\sice_ICS_reg[2]/NET0131 ,
		_w26294_,
		_w26328_
	);
	LUT2 #(
		.INIT('h2)
	) name22282 (
		T_IMS_pad,
		_w23031_,
		_w26329_
	);
	LUT2 #(
		.INIT('h1)
	) name22283 (
		\sice_ICS_reg[1]/NET0131 ,
		_w26329_,
		_w26330_
	);
	LUT2 #(
		.INIT('h8)
	) name22284 (
		\sice_ICS_reg[1]/NET0131 ,
		_w26329_,
		_w26331_
	);
	LUT2 #(
		.INIT('h1)
	) name22285 (
		_w26328_,
		_w26330_,
		_w26332_
	);
	LUT2 #(
		.INIT('h4)
	) name22286 (
		_w26331_,
		_w26332_,
		_w26333_
	);
	LUT2 #(
		.INIT('h8)
	) name22287 (
		_w12234_,
		_w26333_,
		_w26334_
	);
	LUT2 #(
		.INIT('h4)
	) name22288 (
		\sice_ICS_reg[1]/NET0131 ,
		_w26298_,
		_w26335_
	);
	LUT2 #(
		.INIT('h1)
	) name22289 (
		T_IMS_pad,
		_w26335_,
		_w26336_
	);
	LUT2 #(
		.INIT('h8)
	) name22290 (
		_w12234_,
		_w26336_,
		_w26337_
	);
	LUT2 #(
		.INIT('h4)
	) name22291 (
		\sice_ICYC_clr_reg/NET0131 ,
		_w4149_,
		_w26338_
	);
	LUT2 #(
		.INIT('h4)
	) name22292 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w26339_
	);
	LUT2 #(
		.INIT('h4)
	) name22293 (
		_w18264_,
		_w26339_,
		_w26340_
	);
	LUT2 #(
		.INIT('h4)
	) name22294 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w26341_
	);
	LUT2 #(
		.INIT('h4)
	) name22295 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w26342_
	);
	LUT2 #(
		.INIT('h8)
	) name22296 (
		_w26341_,
		_w26342_,
		_w26343_
	);
	LUT2 #(
		.INIT('h1)
	) name22297 (
		_w26340_,
		_w26343_,
		_w26344_
	);
	LUT2 #(
		.INIT('h2)
	) name22298 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w26344_,
		_w26345_
	);
	LUT2 #(
		.INIT('h2)
	) name22299 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w26346_
	);
	LUT2 #(
		.INIT('h8)
	) name22300 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w17801_,
		_w26347_
	);
	LUT2 #(
		.INIT('h2)
	) name22301 (
		_w17805_,
		_w26347_,
		_w26348_
	);
	LUT2 #(
		.INIT('h2)
	) name22302 (
		_w26346_,
		_w26348_,
		_w26349_
	);
	LUT2 #(
		.INIT('h2)
	) name22303 (
		\core_c_dec_updAR_E_reg/P0001 ,
		_w13802_,
		_w26350_
	);
	LUT2 #(
		.INIT('h1)
	) name22304 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w26350_,
		_w26351_
	);
	LUT2 #(
		.INIT('h1)
	) name22305 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w26352_
	);
	LUT2 #(
		.INIT('h8)
	) name22306 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w26352_,
		_w26353_
	);
	LUT2 #(
		.INIT('h4)
	) name22307 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w26353_,
		_w26354_
	);
	LUT2 #(
		.INIT('h4)
	) name22308 (
		_w26351_,
		_w26354_,
		_w26355_
	);
	LUT2 #(
		.INIT('h8)
	) name22309 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w26356_
	);
	LUT2 #(
		.INIT('h8)
	) name22310 (
		\core_c_dec_updSR_E_reg/P0001 ,
		_w13803_,
		_w26357_
	);
	LUT2 #(
		.INIT('h8)
	) name22311 (
		_w18846_,
		_w21525_,
		_w26358_
	);
	LUT2 #(
		.INIT('h2)
	) name22312 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w26358_,
		_w26359_
	);
	LUT2 #(
		.INIT('h2)
	) name22313 (
		_w26356_,
		_w26359_,
		_w26360_
	);
	LUT2 #(
		.INIT('h8)
	) name22314 (
		_w26357_,
		_w26360_,
		_w26361_
	);
	LUT2 #(
		.INIT('h4)
	) name22315 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w26362_
	);
	LUT2 #(
		.INIT('h1)
	) name22316 (
		_w26357_,
		_w26362_,
		_w26363_
	);
	LUT2 #(
		.INIT('h8)
	) name22317 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w26356_,
		_w26364_
	);
	LUT2 #(
		.INIT('h4)
	) name22318 (
		_w26363_,
		_w26364_,
		_w26365_
	);
	LUT2 #(
		.INIT('h1)
	) name22319 (
		_w26345_,
		_w26349_,
		_w26366_
	);
	LUT2 #(
		.INIT('h4)
	) name22320 (
		_w26355_,
		_w26366_,
		_w26367_
	);
	LUT2 #(
		.INIT('h4)
	) name22321 (
		_w26361_,
		_w26367_,
		_w26368_
	);
	LUT2 #(
		.INIT('h4)
	) name22322 (
		_w26365_,
		_w26368_,
		_w26369_
	);
	LUT2 #(
		.INIT('h2)
	) name22323 (
		_w18847_,
		_w26369_,
		_w26370_
	);
	LUT2 #(
		.INIT('h8)
	) name22324 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w26339_,
		_w26371_
	);
	LUT2 #(
		.INIT('h8)
	) name22325 (
		_w18263_,
		_w26371_,
		_w26372_
	);
	LUT2 #(
		.INIT('h1)
	) name22326 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w26373_
	);
	LUT2 #(
		.INIT('h8)
	) name22327 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w26341_,
		_w26374_
	);
	LUT2 #(
		.INIT('h8)
	) name22328 (
		_w26373_,
		_w26374_,
		_w26375_
	);
	LUT2 #(
		.INIT('h1)
	) name22329 (
		_w26372_,
		_w26375_,
		_w26376_
	);
	LUT2 #(
		.INIT('h2)
	) name22330 (
		_w26370_,
		_w26376_,
		_w26377_
	);
	LUT2 #(
		.INIT('h4)
	) name22331 (
		_w5689_,
		_w26377_,
		_w26378_
	);
	LUT2 #(
		.INIT('h4)
	) name22332 (
		_w5689_,
		_w26346_,
		_w26379_
	);
	LUT2 #(
		.INIT('h8)
	) name22333 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w26379_,
		_w26380_
	);
	LUT2 #(
		.INIT('h8)
	) name22334 (
		_w17802_,
		_w26380_,
		_w26381_
	);
	LUT2 #(
		.INIT('h8)
	) name22335 (
		_w26370_,
		_w26381_,
		_w26382_
	);
	LUT2 #(
		.INIT('h1)
	) name22336 (
		_w26378_,
		_w26382_,
		_w26383_
	);
	LUT2 #(
		.INIT('h8)
	) name22337 (
		_w26346_,
		_w26347_,
		_w26384_
	);
	LUT2 #(
		.INIT('h8)
	) name22338 (
		_w18847_,
		_w26384_,
		_w26385_
	);
	LUT2 #(
		.INIT('h8)
	) name22339 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w26385_,
		_w26386_
	);
	LUT2 #(
		.INIT('h4)
	) name22340 (
		_w5689_,
		_w26386_,
		_w26387_
	);
	LUT2 #(
		.INIT('h2)
	) name22341 (
		_w26383_,
		_w26387_,
		_w26388_
	);
	LUT2 #(
		.INIT('h8)
	) name22342 (
		_w26383_,
		_w26387_,
		_w26389_
	);
	LUT2 #(
		.INIT('h1)
	) name22343 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w5689_,
		_w26390_
	);
	LUT2 #(
		.INIT('h8)
	) name22344 (
		_w26385_,
		_w26390_,
		_w26391_
	);
	LUT2 #(
		.INIT('h1)
	) name22345 (
		_w26386_,
		_w26391_,
		_w26392_
	);
	LUT2 #(
		.INIT('h8)
	) name22346 (
		_w26382_,
		_w26392_,
		_w26393_
	);
	LUT2 #(
		.INIT('h1)
	) name22347 (
		_w26389_,
		_w26393_,
		_w26394_
	);
	LUT2 #(
		.INIT('h4)
	) name22348 (
		_w26378_,
		_w26394_,
		_w26395_
	);
	LUT2 #(
		.INIT('h4)
	) name22349 (
		_w26388_,
		_w26395_,
		_w26396_
	);
	LUT2 #(
		.INIT('h2)
	) name22350 (
		\sport0_txctl_TXSHT_reg[12]/P0001 ,
		_w19960_,
		_w26397_
	);
	LUT2 #(
		.INIT('h8)
	) name22351 (
		\sport0_txctl_TX_reg[13]/P0001 ,
		_w19960_,
		_w26398_
	);
	LUT2 #(
		.INIT('h1)
	) name22352 (
		_w26397_,
		_w26398_,
		_w26399_
	);
	LUT2 #(
		.INIT('h1)
	) name22353 (
		\core_c_psq_PCS_reg[0]/NET0131 ,
		\core_c_psq_PCS_reg[15]/NET0131 ,
		_w26400_
	);
	LUT2 #(
		.INIT('h4)
	) name22354 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		\sice_GOICE_syn_reg/P0001 ,
		_w26401_
	);
	LUT2 #(
		.INIT('h8)
	) name22355 (
		_w26400_,
		_w26401_,
		_w26402_
	);
	LUT2 #(
		.INIT('h8)
	) name22356 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		\sice_ITR_reg[0]/NET0131 ,
		_w26403_
	);
	LUT2 #(
		.INIT('h8)
	) name22357 (
		_w23230_,
		_w26403_,
		_w26404_
	);
	LUT2 #(
		.INIT('h1)
	) name22358 (
		\sice_DBR1_reg[11]/P0001 ,
		\sice_DMR1_reg[11]/NET0131 ,
		_w26405_
	);
	LUT2 #(
		.INIT('h8)
	) name22359 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		_w26405_,
		_w26406_
	);
	LUT2 #(
		.INIT('h1)
	) name22360 (
		\sice_DBR1_reg[10]/P0001 ,
		\sice_DMR1_reg[10]/NET0131 ,
		_w26407_
	);
	LUT2 #(
		.INIT('h8)
	) name22361 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w26407_,
		_w26408_
	);
	LUT2 #(
		.INIT('h2)
	) name22362 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[16]/P0001 ,
		_w26409_
	);
	LUT2 #(
		.INIT('h4)
	) name22363 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[16]/P0001 ,
		_w26410_
	);
	LUT2 #(
		.INIT('h1)
	) name22364 (
		_w26409_,
		_w26410_,
		_w26411_
	);
	LUT2 #(
		.INIT('h1)
	) name22365 (
		\sice_DMR1_reg[16]/NET0131 ,
		_w26411_,
		_w26412_
	);
	LUT2 #(
		.INIT('h1)
	) name22366 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[1]/P0001 ,
		_w26413_
	);
	LUT2 #(
		.INIT('h8)
	) name22367 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[1]/P0001 ,
		_w26414_
	);
	LUT2 #(
		.INIT('h1)
	) name22368 (
		\sice_DMR1_reg[1]/NET0131 ,
		_w26413_,
		_w26415_
	);
	LUT2 #(
		.INIT('h4)
	) name22369 (
		_w26414_,
		_w26415_,
		_w26416_
	);
	LUT2 #(
		.INIT('h1)
	) name22370 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[3]/P0001 ,
		_w26417_
	);
	LUT2 #(
		.INIT('h8)
	) name22371 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[3]/P0001 ,
		_w26418_
	);
	LUT2 #(
		.INIT('h1)
	) name22372 (
		\sice_DMR1_reg[3]/NET0131 ,
		_w26417_,
		_w26419_
	);
	LUT2 #(
		.INIT('h4)
	) name22373 (
		_w26418_,
		_w26419_,
		_w26420_
	);
	LUT2 #(
		.INIT('h1)
	) name22374 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[15]/P0001 ,
		_w26421_
	);
	LUT2 #(
		.INIT('h8)
	) name22375 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[15]/P0001 ,
		_w26422_
	);
	LUT2 #(
		.INIT('h1)
	) name22376 (
		\sice_DMR1_reg[15]/NET0131 ,
		_w26421_,
		_w26423_
	);
	LUT2 #(
		.INIT('h4)
	) name22377 (
		_w26422_,
		_w26423_,
		_w26424_
	);
	LUT2 #(
		.INIT('h1)
	) name22378 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[17]/P0001 ,
		_w26425_
	);
	LUT2 #(
		.INIT('h8)
	) name22379 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[17]/P0001 ,
		_w26426_
	);
	LUT2 #(
		.INIT('h1)
	) name22380 (
		_w26425_,
		_w26426_,
		_w26427_
	);
	LUT2 #(
		.INIT('h1)
	) name22381 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[2]/P0001 ,
		_w26428_
	);
	LUT2 #(
		.INIT('h8)
	) name22382 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[2]/P0001 ,
		_w26429_
	);
	LUT2 #(
		.INIT('h1)
	) name22383 (
		\sice_DMR1_reg[2]/NET0131 ,
		_w26428_,
		_w26430_
	);
	LUT2 #(
		.INIT('h4)
	) name22384 (
		_w26429_,
		_w26430_,
		_w26431_
	);
	LUT2 #(
		.INIT('h2)
	) name22385 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[14]/P0001 ,
		_w26432_
	);
	LUT2 #(
		.INIT('h4)
	) name22386 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[14]/P0001 ,
		_w26433_
	);
	LUT2 #(
		.INIT('h1)
	) name22387 (
		_w26432_,
		_w26433_,
		_w26434_
	);
	LUT2 #(
		.INIT('h1)
	) name22388 (
		\sice_DMR1_reg[14]/NET0131 ,
		_w26434_,
		_w26435_
	);
	LUT2 #(
		.INIT('h1)
	) name22389 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR1_reg[4]/P0001 ,
		_w26436_
	);
	LUT2 #(
		.INIT('h8)
	) name22390 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR1_reg[4]/P0001 ,
		_w26437_
	);
	LUT2 #(
		.INIT('h1)
	) name22391 (
		\sice_DMR1_reg[4]/NET0131 ,
		_w26436_,
		_w26438_
	);
	LUT2 #(
		.INIT('h4)
	) name22392 (
		_w26437_,
		_w26438_,
		_w26439_
	);
	LUT2 #(
		.INIT('h1)
	) name22393 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR1_reg[13]/P0001 ,
		_w26440_
	);
	LUT2 #(
		.INIT('h8)
	) name22394 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR1_reg[13]/P0001 ,
		_w26441_
	);
	LUT2 #(
		.INIT('h1)
	) name22395 (
		\sice_DMR1_reg[13]/NET0131 ,
		_w26440_,
		_w26442_
	);
	LUT2 #(
		.INIT('h4)
	) name22396 (
		_w26441_,
		_w26442_,
		_w26443_
	);
	LUT2 #(
		.INIT('h2)
	) name22397 (
		\sice_DBR1_reg[10]/P0001 ,
		\sice_DMR1_reg[10]/NET0131 ,
		_w26444_
	);
	LUT2 #(
		.INIT('h4)
	) name22398 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w26444_,
		_w26445_
	);
	LUT2 #(
		.INIT('h2)
	) name22399 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR1_reg[5]/P0001 ,
		_w26446_
	);
	LUT2 #(
		.INIT('h4)
	) name22400 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR1_reg[5]/P0001 ,
		_w26447_
	);
	LUT2 #(
		.INIT('h1)
	) name22401 (
		_w26446_,
		_w26447_,
		_w26448_
	);
	LUT2 #(
		.INIT('h1)
	) name22402 (
		\sice_DMR1_reg[5]/NET0131 ,
		_w26448_,
		_w26449_
	);
	LUT2 #(
		.INIT('h1)
	) name22403 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR1_reg[12]/P0001 ,
		_w26450_
	);
	LUT2 #(
		.INIT('h8)
	) name22404 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR1_reg[12]/P0001 ,
		_w26451_
	);
	LUT2 #(
		.INIT('h1)
	) name22405 (
		\sice_DMR1_reg[12]/NET0131 ,
		_w26450_,
		_w26452_
	);
	LUT2 #(
		.INIT('h4)
	) name22406 (
		_w26451_,
		_w26452_,
		_w26453_
	);
	LUT2 #(
		.INIT('h2)
	) name22407 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR1_reg[8]/P0001 ,
		_w26454_
	);
	LUT2 #(
		.INIT('h4)
	) name22408 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR1_reg[8]/P0001 ,
		_w26455_
	);
	LUT2 #(
		.INIT('h1)
	) name22409 (
		_w26454_,
		_w26455_,
		_w26456_
	);
	LUT2 #(
		.INIT('h1)
	) name22410 (
		\sice_DMR1_reg[8]/NET0131 ,
		_w26456_,
		_w26457_
	);
	LUT2 #(
		.INIT('h1)
	) name22411 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[0]/P0001 ,
		_w26458_
	);
	LUT2 #(
		.INIT('h8)
	) name22412 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[0]/P0001 ,
		_w26459_
	);
	LUT2 #(
		.INIT('h1)
	) name22413 (
		\sice_DMR1_reg[0]/NET0131 ,
		_w26458_,
		_w26460_
	);
	LUT2 #(
		.INIT('h4)
	) name22414 (
		_w26459_,
		_w26460_,
		_w26461_
	);
	LUT2 #(
		.INIT('h1)
	) name22415 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR1_reg[6]/P0001 ,
		_w26462_
	);
	LUT2 #(
		.INIT('h8)
	) name22416 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR1_reg[6]/P0001 ,
		_w26463_
	);
	LUT2 #(
		.INIT('h1)
	) name22417 (
		\sice_DMR1_reg[6]/NET0131 ,
		_w26462_,
		_w26464_
	);
	LUT2 #(
		.INIT('h4)
	) name22418 (
		_w26463_,
		_w26464_,
		_w26465_
	);
	LUT2 #(
		.INIT('h2)
	) name22419 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR1_reg[9]/P0001 ,
		_w26466_
	);
	LUT2 #(
		.INIT('h4)
	) name22420 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR1_reg[9]/P0001 ,
		_w26467_
	);
	LUT2 #(
		.INIT('h1)
	) name22421 (
		_w26466_,
		_w26467_,
		_w26468_
	);
	LUT2 #(
		.INIT('h1)
	) name22422 (
		\sice_DMR1_reg[9]/NET0131 ,
		_w26468_,
		_w26469_
	);
	LUT2 #(
		.INIT('h2)
	) name22423 (
		\sice_DBR1_reg[11]/P0001 ,
		\sice_DMR1_reg[11]/NET0131 ,
		_w26470_
	);
	LUT2 #(
		.INIT('h4)
	) name22424 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		_w26470_,
		_w26471_
	);
	LUT2 #(
		.INIT('h1)
	) name22425 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR1_reg[7]/P0001 ,
		_w26472_
	);
	LUT2 #(
		.INIT('h8)
	) name22426 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR1_reg[7]/P0001 ,
		_w26473_
	);
	LUT2 #(
		.INIT('h1)
	) name22427 (
		\sice_DMR1_reg[7]/NET0131 ,
		_w26472_,
		_w26474_
	);
	LUT2 #(
		.INIT('h4)
	) name22428 (
		_w26473_,
		_w26474_,
		_w26475_
	);
	LUT2 #(
		.INIT('h4)
	) name22429 (
		\sice_DBR1_reg[18]/P0001 ,
		\sice_DMR1_reg[17]/NET0131 ,
		_w26476_
	);
	LUT2 #(
		.INIT('h4)
	) name22430 (
		_w26406_,
		_w26476_,
		_w26477_
	);
	LUT2 #(
		.INIT('h1)
	) name22431 (
		_w26408_,
		_w26427_,
		_w26478_
	);
	LUT2 #(
		.INIT('h1)
	) name22432 (
		_w26445_,
		_w26471_,
		_w26479_
	);
	LUT2 #(
		.INIT('h8)
	) name22433 (
		_w26478_,
		_w26479_,
		_w26480_
	);
	LUT2 #(
		.INIT('h4)
	) name22434 (
		_w26412_,
		_w26477_,
		_w26481_
	);
	LUT2 #(
		.INIT('h1)
	) name22435 (
		_w26416_,
		_w26420_,
		_w26482_
	);
	LUT2 #(
		.INIT('h1)
	) name22436 (
		_w26424_,
		_w26431_,
		_w26483_
	);
	LUT2 #(
		.INIT('h1)
	) name22437 (
		_w26435_,
		_w26439_,
		_w26484_
	);
	LUT2 #(
		.INIT('h1)
	) name22438 (
		_w26443_,
		_w26449_,
		_w26485_
	);
	LUT2 #(
		.INIT('h1)
	) name22439 (
		_w26453_,
		_w26457_,
		_w26486_
	);
	LUT2 #(
		.INIT('h1)
	) name22440 (
		_w26461_,
		_w26465_,
		_w26487_
	);
	LUT2 #(
		.INIT('h1)
	) name22441 (
		_w26469_,
		_w26475_,
		_w26488_
	);
	LUT2 #(
		.INIT('h8)
	) name22442 (
		_w26487_,
		_w26488_,
		_w26489_
	);
	LUT2 #(
		.INIT('h8)
	) name22443 (
		_w26485_,
		_w26486_,
		_w26490_
	);
	LUT2 #(
		.INIT('h8)
	) name22444 (
		_w26483_,
		_w26484_,
		_w26491_
	);
	LUT2 #(
		.INIT('h8)
	) name22445 (
		_w26481_,
		_w26482_,
		_w26492_
	);
	LUT2 #(
		.INIT('h8)
	) name22446 (
		_w26480_,
		_w26492_,
		_w26493_
	);
	LUT2 #(
		.INIT('h8)
	) name22447 (
		_w26490_,
		_w26491_,
		_w26494_
	);
	LUT2 #(
		.INIT('h8)
	) name22448 (
		_w26489_,
		_w26494_,
		_w26495_
	);
	LUT2 #(
		.INIT('h8)
	) name22449 (
		_w26493_,
		_w26495_,
		_w26496_
	);
	LUT2 #(
		.INIT('h1)
	) name22450 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR2_reg[9]/P0001 ,
		_w26497_
	);
	LUT2 #(
		.INIT('h8)
	) name22451 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR2_reg[9]/P0001 ,
		_w26498_
	);
	LUT2 #(
		.INIT('h1)
	) name22452 (
		\sice_DMR2_reg[9]/NET0131 ,
		_w26497_,
		_w26499_
	);
	LUT2 #(
		.INIT('h4)
	) name22453 (
		_w26498_,
		_w26499_,
		_w26500_
	);
	LUT2 #(
		.INIT('h1)
	) name22454 (
		\sice_DBR2_reg[5]/P0001 ,
		\sice_DMR2_reg[5]/NET0131 ,
		_w26501_
	);
	LUT2 #(
		.INIT('h8)
	) name22455 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		_w26501_,
		_w26502_
	);
	LUT2 #(
		.INIT('h1)
	) name22456 (
		\sice_DBR2_reg[10]/P0001 ,
		\sice_DMR2_reg[10]/NET0131 ,
		_w26503_
	);
	LUT2 #(
		.INIT('h8)
	) name22457 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w26503_,
		_w26504_
	);
	LUT2 #(
		.INIT('h2)
	) name22458 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR2_reg[11]/P0001 ,
		_w26505_
	);
	LUT2 #(
		.INIT('h4)
	) name22459 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR2_reg[11]/P0001 ,
		_w26506_
	);
	LUT2 #(
		.INIT('h1)
	) name22460 (
		_w26505_,
		_w26506_,
		_w26507_
	);
	LUT2 #(
		.INIT('h1)
	) name22461 (
		\sice_DMR2_reg[11]/NET0131 ,
		_w26507_,
		_w26508_
	);
	LUT2 #(
		.INIT('h2)
	) name22462 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR2_reg[4]/P0001 ,
		_w26509_
	);
	LUT2 #(
		.INIT('h4)
	) name22463 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR2_reg[4]/P0001 ,
		_w26510_
	);
	LUT2 #(
		.INIT('h1)
	) name22464 (
		_w26509_,
		_w26510_,
		_w26511_
	);
	LUT2 #(
		.INIT('h1)
	) name22465 (
		\sice_DMR2_reg[4]/NET0131 ,
		_w26511_,
		_w26512_
	);
	LUT2 #(
		.INIT('h1)
	) name22466 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[14]/P0001 ,
		_w26513_
	);
	LUT2 #(
		.INIT('h8)
	) name22467 (
		\core_c_psq_PMOVL_regh_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[14]/P0001 ,
		_w26514_
	);
	LUT2 #(
		.INIT('h1)
	) name22468 (
		\sice_DMR2_reg[14]/NET0131 ,
		_w26513_,
		_w26515_
	);
	LUT2 #(
		.INIT('h4)
	) name22469 (
		_w26514_,
		_w26515_,
		_w26516_
	);
	LUT2 #(
		.INIT('h2)
	) name22470 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR2_reg[8]/P0001 ,
		_w26517_
	);
	LUT2 #(
		.INIT('h4)
	) name22471 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR2_reg[8]/P0001 ,
		_w26518_
	);
	LUT2 #(
		.INIT('h1)
	) name22472 (
		_w26517_,
		_w26518_,
		_w26519_
	);
	LUT2 #(
		.INIT('h1)
	) name22473 (
		\sice_DMR2_reg[8]/NET0131 ,
		_w26519_,
		_w26520_
	);
	LUT2 #(
		.INIT('h1)
	) name22474 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[15]/P0001 ,
		_w26521_
	);
	LUT2 #(
		.INIT('h8)
	) name22475 (
		\core_c_psq_PMOVL_regh_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[15]/P0001 ,
		_w26522_
	);
	LUT2 #(
		.INIT('h1)
	) name22476 (
		\sice_DMR2_reg[15]/NET0131 ,
		_w26521_,
		_w26523_
	);
	LUT2 #(
		.INIT('h4)
	) name22477 (
		_w26522_,
		_w26523_,
		_w26524_
	);
	LUT2 #(
		.INIT('h1)
	) name22478 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR2_reg[6]/P0001 ,
		_w26525_
	);
	LUT2 #(
		.INIT('h8)
	) name22479 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR2_reg[6]/P0001 ,
		_w26526_
	);
	LUT2 #(
		.INIT('h1)
	) name22480 (
		\sice_DMR2_reg[6]/NET0131 ,
		_w26525_,
		_w26527_
	);
	LUT2 #(
		.INIT('h4)
	) name22481 (
		_w26526_,
		_w26527_,
		_w26528_
	);
	LUT2 #(
		.INIT('h2)
	) name22482 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[3]/P0001 ,
		_w26529_
	);
	LUT2 #(
		.INIT('h4)
	) name22483 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[3]/P0001 ,
		_w26530_
	);
	LUT2 #(
		.INIT('h1)
	) name22484 (
		_w26529_,
		_w26530_,
		_w26531_
	);
	LUT2 #(
		.INIT('h1)
	) name22485 (
		\sice_DMR2_reg[3]/NET0131 ,
		_w26531_,
		_w26532_
	);
	LUT2 #(
		.INIT('h1)
	) name22486 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR2_reg[12]/P0001 ,
		_w26533_
	);
	LUT2 #(
		.INIT('h8)
	) name22487 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR2_reg[12]/P0001 ,
		_w26534_
	);
	LUT2 #(
		.INIT('h1)
	) name22488 (
		\sice_DMR2_reg[12]/NET0131 ,
		_w26533_,
		_w26535_
	);
	LUT2 #(
		.INIT('h4)
	) name22489 (
		_w26534_,
		_w26535_,
		_w26536_
	);
	LUT2 #(
		.INIT('h1)
	) name22490 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[1]/P0001 ,
		_w26537_
	);
	LUT2 #(
		.INIT('h8)
	) name22491 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[1]/P0001 ,
		_w26538_
	);
	LUT2 #(
		.INIT('h1)
	) name22492 (
		\sice_DMR2_reg[1]/NET0131 ,
		_w26537_,
		_w26539_
	);
	LUT2 #(
		.INIT('h4)
	) name22493 (
		_w26538_,
		_w26539_,
		_w26540_
	);
	LUT2 #(
		.INIT('h1)
	) name22494 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[16]/P0001 ,
		_w26541_
	);
	LUT2 #(
		.INIT('h8)
	) name22495 (
		\core_c_psq_PMOVL_regh_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[16]/P0001 ,
		_w26542_
	);
	LUT2 #(
		.INIT('h1)
	) name22496 (
		\sice_DMR2_reg[16]/NET0131 ,
		_w26541_,
		_w26543_
	);
	LUT2 #(
		.INIT('h4)
	) name22497 (
		_w26542_,
		_w26543_,
		_w26544_
	);
	LUT2 #(
		.INIT('h2)
	) name22498 (
		\sice_DBR2_reg[10]/P0001 ,
		\sice_DMR2_reg[10]/NET0131 ,
		_w26545_
	);
	LUT2 #(
		.INIT('h4)
	) name22499 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[10]/NET0131 ,
		_w26545_,
		_w26546_
	);
	LUT2 #(
		.INIT('h2)
	) name22500 (
		\sice_DBR2_reg[5]/P0001 ,
		\sice_DMR2_reg[5]/NET0131 ,
		_w26547_
	);
	LUT2 #(
		.INIT('h4)
	) name22501 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[5]/NET0131 ,
		_w26547_,
		_w26548_
	);
	LUT2 #(
		.INIT('h2)
	) name22502 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR2_reg[7]/P0001 ,
		_w26549_
	);
	LUT2 #(
		.INIT('h4)
	) name22503 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR2_reg[7]/P0001 ,
		_w26550_
	);
	LUT2 #(
		.INIT('h1)
	) name22504 (
		_w26549_,
		_w26550_,
		_w26551_
	);
	LUT2 #(
		.INIT('h1)
	) name22505 (
		\sice_DMR2_reg[7]/NET0131 ,
		_w26551_,
		_w26552_
	);
	LUT2 #(
		.INIT('h2)
	) name22506 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[2]/P0001 ,
		_w26553_
	);
	LUT2 #(
		.INIT('h4)
	) name22507 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[2]/P0001 ,
		_w26554_
	);
	LUT2 #(
		.INIT('h1)
	) name22508 (
		_w26553_,
		_w26554_,
		_w26555_
	);
	LUT2 #(
		.INIT('h1)
	) name22509 (
		\sice_DMR2_reg[2]/NET0131 ,
		_w26555_,
		_w26556_
	);
	LUT2 #(
		.INIT('h1)
	) name22510 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[0]/P0001 ,
		_w26557_
	);
	LUT2 #(
		.INIT('h8)
	) name22511 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[0]/P0001 ,
		_w26558_
	);
	LUT2 #(
		.INIT('h1)
	) name22512 (
		\sice_DMR2_reg[0]/NET0131 ,
		_w26557_,
		_w26559_
	);
	LUT2 #(
		.INIT('h4)
	) name22513 (
		_w26558_,
		_w26559_,
		_w26560_
	);
	LUT2 #(
		.INIT('h1)
	) name22514 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR2_reg[13]/P0001 ,
		_w26561_
	);
	LUT2 #(
		.INIT('h8)
	) name22515 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR2_reg[13]/P0001 ,
		_w26562_
	);
	LUT2 #(
		.INIT('h1)
	) name22516 (
		\sice_DMR2_reg[13]/NET0131 ,
		_w26561_,
		_w26563_
	);
	LUT2 #(
		.INIT('h4)
	) name22517 (
		_w26562_,
		_w26563_,
		_w26564_
	);
	LUT2 #(
		.INIT('h2)
	) name22518 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[17]/P0001 ,
		_w26565_
	);
	LUT2 #(
		.INIT('h4)
	) name22519 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[17]/P0001 ,
		_w26566_
	);
	LUT2 #(
		.INIT('h4)
	) name22520 (
		\sice_DBR2_reg[18]/P0001 ,
		\sice_DMR2_reg[17]/NET0131 ,
		_w26567_
	);
	LUT2 #(
		.INIT('h4)
	) name22521 (
		_w26565_,
		_w26567_,
		_w26568_
	);
	LUT2 #(
		.INIT('h4)
	) name22522 (
		_w26566_,
		_w26568_,
		_w26569_
	);
	LUT2 #(
		.INIT('h1)
	) name22523 (
		_w26502_,
		_w26504_,
		_w26570_
	);
	LUT2 #(
		.INIT('h1)
	) name22524 (
		_w26546_,
		_w26548_,
		_w26571_
	);
	LUT2 #(
		.INIT('h8)
	) name22525 (
		_w26570_,
		_w26571_,
		_w26572_
	);
	LUT2 #(
		.INIT('h4)
	) name22526 (
		_w26500_,
		_w26569_,
		_w26573_
	);
	LUT2 #(
		.INIT('h1)
	) name22527 (
		_w26508_,
		_w26512_,
		_w26574_
	);
	LUT2 #(
		.INIT('h1)
	) name22528 (
		_w26516_,
		_w26520_,
		_w26575_
	);
	LUT2 #(
		.INIT('h1)
	) name22529 (
		_w26524_,
		_w26528_,
		_w26576_
	);
	LUT2 #(
		.INIT('h1)
	) name22530 (
		_w26532_,
		_w26536_,
		_w26577_
	);
	LUT2 #(
		.INIT('h1)
	) name22531 (
		_w26540_,
		_w26544_,
		_w26578_
	);
	LUT2 #(
		.INIT('h1)
	) name22532 (
		_w26552_,
		_w26556_,
		_w26579_
	);
	LUT2 #(
		.INIT('h1)
	) name22533 (
		_w26560_,
		_w26564_,
		_w26580_
	);
	LUT2 #(
		.INIT('h8)
	) name22534 (
		_w26579_,
		_w26580_,
		_w26581_
	);
	LUT2 #(
		.INIT('h8)
	) name22535 (
		_w26577_,
		_w26578_,
		_w26582_
	);
	LUT2 #(
		.INIT('h8)
	) name22536 (
		_w26575_,
		_w26576_,
		_w26583_
	);
	LUT2 #(
		.INIT('h8)
	) name22537 (
		_w26573_,
		_w26574_,
		_w26584_
	);
	LUT2 #(
		.INIT('h8)
	) name22538 (
		_w26572_,
		_w26584_,
		_w26585_
	);
	LUT2 #(
		.INIT('h8)
	) name22539 (
		_w26582_,
		_w26583_,
		_w26586_
	);
	LUT2 #(
		.INIT('h8)
	) name22540 (
		_w26581_,
		_w26586_,
		_w26587_
	);
	LUT2 #(
		.INIT('h8)
	) name22541 (
		_w26585_,
		_w26587_,
		_w26588_
	);
	LUT2 #(
		.INIT('h1)
	) name22542 (
		_w26496_,
		_w26588_,
		_w26589_
	);
	LUT2 #(
		.INIT('h4)
	) name22543 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\memc_accPM_E_reg/NET0131 ,
		_w26590_
	);
	LUT2 #(
		.INIT('h4)
	) name22544 (
		_w26589_,
		_w26590_,
		_w26591_
	);
	LUT2 #(
		.INIT('h4)
	) name22545 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w26545_,
		_w26592_
	);
	LUT2 #(
		.INIT('h4)
	) name22546 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		_w26547_,
		_w26593_
	);
	LUT2 #(
		.INIT('h2)
	) name22547 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[3]/P0001 ,
		_w26594_
	);
	LUT2 #(
		.INIT('h4)
	) name22548 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[3]/P0001 ,
		_w26595_
	);
	LUT2 #(
		.INIT('h1)
	) name22549 (
		_w26594_,
		_w26595_,
		_w26596_
	);
	LUT2 #(
		.INIT('h1)
	) name22550 (
		\sice_DMR2_reg[3]/NET0131 ,
		_w26596_,
		_w26597_
	);
	LUT2 #(
		.INIT('h1)
	) name22551 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[1]/P0001 ,
		_w26598_
	);
	LUT2 #(
		.INIT('h8)
	) name22552 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[1]/P0001 ,
		_w26599_
	);
	LUT2 #(
		.INIT('h1)
	) name22553 (
		\sice_DMR2_reg[1]/NET0131 ,
		_w26598_,
		_w26600_
	);
	LUT2 #(
		.INIT('h4)
	) name22554 (
		_w26599_,
		_w26600_,
		_w26601_
	);
	LUT2 #(
		.INIT('h2)
	) name22555 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR2_reg[11]/P0001 ,
		_w26602_
	);
	LUT2 #(
		.INIT('h4)
	) name22556 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		\sice_DBR2_reg[11]/P0001 ,
		_w26603_
	);
	LUT2 #(
		.INIT('h1)
	) name22557 (
		_w26602_,
		_w26603_,
		_w26604_
	);
	LUT2 #(
		.INIT('h1)
	) name22558 (
		\sice_DMR2_reg[11]/NET0131 ,
		_w26604_,
		_w26605_
	);
	LUT2 #(
		.INIT('h1)
	) name22559 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR2_reg[12]/P0001 ,
		_w26606_
	);
	LUT2 #(
		.INIT('h8)
	) name22560 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR2_reg[12]/P0001 ,
		_w26607_
	);
	LUT2 #(
		.INIT('h1)
	) name22561 (
		\sice_DMR2_reg[12]/NET0131 ,
		_w26606_,
		_w26608_
	);
	LUT2 #(
		.INIT('h4)
	) name22562 (
		_w26607_,
		_w26608_,
		_w26609_
	);
	LUT2 #(
		.INIT('h1)
	) name22563 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR2_reg[6]/P0001 ,
		_w26610_
	);
	LUT2 #(
		.INIT('h8)
	) name22564 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR2_reg[6]/P0001 ,
		_w26611_
	);
	LUT2 #(
		.INIT('h1)
	) name22565 (
		\sice_DMR2_reg[6]/NET0131 ,
		_w26610_,
		_w26612_
	);
	LUT2 #(
		.INIT('h4)
	) name22566 (
		_w26611_,
		_w26612_,
		_w26613_
	);
	LUT2 #(
		.INIT('h1)
	) name22567 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR2_reg[8]/P0001 ,
		_w26614_
	);
	LUT2 #(
		.INIT('h8)
	) name22568 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR2_reg[8]/P0001 ,
		_w26615_
	);
	LUT2 #(
		.INIT('h1)
	) name22569 (
		\sice_DMR2_reg[8]/NET0131 ,
		_w26614_,
		_w26616_
	);
	LUT2 #(
		.INIT('h4)
	) name22570 (
		_w26615_,
		_w26616_,
		_w26617_
	);
	LUT2 #(
		.INIT('h2)
	) name22571 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[16]/P0001 ,
		_w26618_
	);
	LUT2 #(
		.INIT('h4)
	) name22572 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[16]/P0001 ,
		_w26619_
	);
	LUT2 #(
		.INIT('h1)
	) name22573 (
		_w26618_,
		_w26619_,
		_w26620_
	);
	LUT2 #(
		.INIT('h1)
	) name22574 (
		\sice_DMR2_reg[16]/NET0131 ,
		_w26620_,
		_w26621_
	);
	LUT2 #(
		.INIT('h1)
	) name22575 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR2_reg[9]/P0001 ,
		_w26622_
	);
	LUT2 #(
		.INIT('h8)
	) name22576 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR2_reg[9]/P0001 ,
		_w26623_
	);
	LUT2 #(
		.INIT('h1)
	) name22577 (
		\sice_DMR2_reg[9]/NET0131 ,
		_w26622_,
		_w26624_
	);
	LUT2 #(
		.INIT('h4)
	) name22578 (
		_w26623_,
		_w26624_,
		_w26625_
	);
	LUT2 #(
		.INIT('h1)
	) name22579 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[0]/P0001 ,
		_w26626_
	);
	LUT2 #(
		.INIT('h8)
	) name22580 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[0]/P0001 ,
		_w26627_
	);
	LUT2 #(
		.INIT('h1)
	) name22581 (
		\sice_DMR2_reg[0]/NET0131 ,
		_w26626_,
		_w26628_
	);
	LUT2 #(
		.INIT('h4)
	) name22582 (
		_w26627_,
		_w26628_,
		_w26629_
	);
	LUT2 #(
		.INIT('h4)
	) name22583 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[17]/P0001 ,
		_w26630_
	);
	LUT2 #(
		.INIT('h4)
	) name22584 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\memc_accDM_E_reg/NET0131 ,
		_w26631_
	);
	LUT2 #(
		.INIT('h2)
	) name22585 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\sice_DBR2_reg[17]/P0001 ,
		_w26632_
	);
	LUT2 #(
		.INIT('h1)
	) name22586 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[15]/P0001 ,
		_w26633_
	);
	LUT2 #(
		.INIT('h8)
	) name22587 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		\sice_DBR2_reg[15]/P0001 ,
		_w26634_
	);
	LUT2 #(
		.INIT('h1)
	) name22588 (
		\sice_DMR2_reg[15]/NET0131 ,
		_w26633_,
		_w26635_
	);
	LUT2 #(
		.INIT('h4)
	) name22589 (
		_w26634_,
		_w26635_,
		_w26636_
	);
	LUT2 #(
		.INIT('h2)
	) name22590 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[14]/P0001 ,
		_w26637_
	);
	LUT2 #(
		.INIT('h4)
	) name22591 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		\sice_DBR2_reg[14]/P0001 ,
		_w26638_
	);
	LUT2 #(
		.INIT('h1)
	) name22592 (
		_w26637_,
		_w26638_,
		_w26639_
	);
	LUT2 #(
		.INIT('h1)
	) name22593 (
		\sice_DMR2_reg[14]/NET0131 ,
		_w26639_,
		_w26640_
	);
	LUT2 #(
		.INIT('h1)
	) name22594 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR2_reg[13]/P0001 ,
		_w26641_
	);
	LUT2 #(
		.INIT('h8)
	) name22595 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR2_reg[13]/P0001 ,
		_w26642_
	);
	LUT2 #(
		.INIT('h1)
	) name22596 (
		\sice_DMR2_reg[13]/NET0131 ,
		_w26641_,
		_w26643_
	);
	LUT2 #(
		.INIT('h4)
	) name22597 (
		_w26642_,
		_w26643_,
		_w26644_
	);
	LUT2 #(
		.INIT('h8)
	) name22598 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w26503_,
		_w26645_
	);
	LUT2 #(
		.INIT('h8)
	) name22599 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		_w26501_,
		_w26646_
	);
	LUT2 #(
		.INIT('h2)
	) name22600 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR2_reg[7]/P0001 ,
		_w26647_
	);
	LUT2 #(
		.INIT('h4)
	) name22601 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR2_reg[7]/P0001 ,
		_w26648_
	);
	LUT2 #(
		.INIT('h1)
	) name22602 (
		_w26647_,
		_w26648_,
		_w26649_
	);
	LUT2 #(
		.INIT('h1)
	) name22603 (
		\sice_DMR2_reg[7]/NET0131 ,
		_w26649_,
		_w26650_
	);
	LUT2 #(
		.INIT('h1)
	) name22604 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[2]/P0001 ,
		_w26651_
	);
	LUT2 #(
		.INIT('h8)
	) name22605 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR2_reg[2]/P0001 ,
		_w26652_
	);
	LUT2 #(
		.INIT('h1)
	) name22606 (
		\sice_DMR2_reg[2]/NET0131 ,
		_w26651_,
		_w26653_
	);
	LUT2 #(
		.INIT('h4)
	) name22607 (
		_w26652_,
		_w26653_,
		_w26654_
	);
	LUT2 #(
		.INIT('h1)
	) name22608 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR2_reg[4]/P0001 ,
		_w26655_
	);
	LUT2 #(
		.INIT('h8)
	) name22609 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR2_reg[4]/P0001 ,
		_w26656_
	);
	LUT2 #(
		.INIT('h1)
	) name22610 (
		\sice_DMR2_reg[4]/NET0131 ,
		_w26655_,
		_w26657_
	);
	LUT2 #(
		.INIT('h4)
	) name22611 (
		_w26656_,
		_w26657_,
		_w26658_
	);
	LUT2 #(
		.INIT('h8)
	) name22612 (
		\sice_DBR2_reg[18]/P0001 ,
		\sice_DMR2_reg[17]/NET0131 ,
		_w26659_
	);
	LUT2 #(
		.INIT('h4)
	) name22613 (
		_w26630_,
		_w26659_,
		_w26660_
	);
	LUT2 #(
		.INIT('h2)
	) name22614 (
		_w26631_,
		_w26632_,
		_w26661_
	);
	LUT2 #(
		.INIT('h8)
	) name22615 (
		_w26660_,
		_w26661_,
		_w26662_
	);
	LUT2 #(
		.INIT('h1)
	) name22616 (
		_w26592_,
		_w26593_,
		_w26663_
	);
	LUT2 #(
		.INIT('h1)
	) name22617 (
		_w26645_,
		_w26646_,
		_w26664_
	);
	LUT2 #(
		.INIT('h8)
	) name22618 (
		_w26663_,
		_w26664_,
		_w26665_
	);
	LUT2 #(
		.INIT('h4)
	) name22619 (
		_w26597_,
		_w26662_,
		_w26666_
	);
	LUT2 #(
		.INIT('h1)
	) name22620 (
		_w26601_,
		_w26605_,
		_w26667_
	);
	LUT2 #(
		.INIT('h1)
	) name22621 (
		_w26609_,
		_w26613_,
		_w26668_
	);
	LUT2 #(
		.INIT('h1)
	) name22622 (
		_w26617_,
		_w26621_,
		_w26669_
	);
	LUT2 #(
		.INIT('h1)
	) name22623 (
		_w26625_,
		_w26629_,
		_w26670_
	);
	LUT2 #(
		.INIT('h1)
	) name22624 (
		_w26636_,
		_w26640_,
		_w26671_
	);
	LUT2 #(
		.INIT('h1)
	) name22625 (
		_w26644_,
		_w26650_,
		_w26672_
	);
	LUT2 #(
		.INIT('h1)
	) name22626 (
		_w26654_,
		_w26658_,
		_w26673_
	);
	LUT2 #(
		.INIT('h8)
	) name22627 (
		_w26672_,
		_w26673_,
		_w26674_
	);
	LUT2 #(
		.INIT('h8)
	) name22628 (
		_w26670_,
		_w26671_,
		_w26675_
	);
	LUT2 #(
		.INIT('h8)
	) name22629 (
		_w26668_,
		_w26669_,
		_w26676_
	);
	LUT2 #(
		.INIT('h8)
	) name22630 (
		_w26666_,
		_w26667_,
		_w26677_
	);
	LUT2 #(
		.INIT('h8)
	) name22631 (
		_w26665_,
		_w26677_,
		_w26678_
	);
	LUT2 #(
		.INIT('h8)
	) name22632 (
		_w26675_,
		_w26676_,
		_w26679_
	);
	LUT2 #(
		.INIT('h8)
	) name22633 (
		_w26674_,
		_w26679_,
		_w26680_
	);
	LUT2 #(
		.INIT('h8)
	) name22634 (
		_w26678_,
		_w26680_,
		_w26681_
	);
	LUT2 #(
		.INIT('h8)
	) name22635 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w26407_,
		_w26682_
	);
	LUT2 #(
		.INIT('h4)
	) name22636 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w26444_,
		_w26683_
	);
	LUT2 #(
		.INIT('h2)
	) name22637 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[2]/P0001 ,
		_w26684_
	);
	LUT2 #(
		.INIT('h4)
	) name22638 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[2]/P0001 ,
		_w26685_
	);
	LUT2 #(
		.INIT('h1)
	) name22639 (
		_w26684_,
		_w26685_,
		_w26686_
	);
	LUT2 #(
		.INIT('h1)
	) name22640 (
		\sice_DMR1_reg[2]/NET0131 ,
		_w26686_,
		_w26687_
	);
	LUT2 #(
		.INIT('h1)
	) name22641 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[16]/P0001 ,
		_w26688_
	);
	LUT2 #(
		.INIT('h8)
	) name22642 (
		\core_c_psq_DMOVL_reg_DO_reg[2]/NET0131 ,
		\sice_DBR1_reg[16]/P0001 ,
		_w26689_
	);
	LUT2 #(
		.INIT('h1)
	) name22643 (
		\sice_DMR1_reg[16]/NET0131 ,
		_w26688_,
		_w26690_
	);
	LUT2 #(
		.INIT('h4)
	) name22644 (
		_w26689_,
		_w26690_,
		_w26691_
	);
	LUT2 #(
		.INIT('h1)
	) name22645 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR1_reg[5]/P0001 ,
		_w26692_
	);
	LUT2 #(
		.INIT('h8)
	) name22646 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		\sice_DBR1_reg[5]/P0001 ,
		_w26693_
	);
	LUT2 #(
		.INIT('h1)
	) name22647 (
		\sice_DMR1_reg[5]/NET0131 ,
		_w26692_,
		_w26694_
	);
	LUT2 #(
		.INIT('h4)
	) name22648 (
		_w26693_,
		_w26694_,
		_w26695_
	);
	LUT2 #(
		.INIT('h1)
	) name22649 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR1_reg[7]/P0001 ,
		_w26696_
	);
	LUT2 #(
		.INIT('h8)
	) name22650 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		\sice_DBR1_reg[7]/P0001 ,
		_w26697_
	);
	LUT2 #(
		.INIT('h1)
	) name22651 (
		\sice_DMR1_reg[7]/NET0131 ,
		_w26696_,
		_w26698_
	);
	LUT2 #(
		.INIT('h4)
	) name22652 (
		_w26697_,
		_w26698_,
		_w26699_
	);
	LUT2 #(
		.INIT('h1)
	) name22653 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR1_reg[12]/P0001 ,
		_w26700_
	);
	LUT2 #(
		.INIT('h8)
	) name22654 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		\sice_DBR1_reg[12]/P0001 ,
		_w26701_
	);
	LUT2 #(
		.INIT('h1)
	) name22655 (
		\sice_DMR1_reg[12]/NET0131 ,
		_w26700_,
		_w26702_
	);
	LUT2 #(
		.INIT('h4)
	) name22656 (
		_w26701_,
		_w26702_,
		_w26703_
	);
	LUT2 #(
		.INIT('h4)
	) name22657 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w26470_,
		_w26704_
	);
	LUT2 #(
		.INIT('h2)
	) name22658 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[1]/P0001 ,
		_w26705_
	);
	LUT2 #(
		.INIT('h4)
	) name22659 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[1]/P0001 ,
		_w26706_
	);
	LUT2 #(
		.INIT('h1)
	) name22660 (
		_w26705_,
		_w26706_,
		_w26707_
	);
	LUT2 #(
		.INIT('h1)
	) name22661 (
		\sice_DMR1_reg[1]/NET0131 ,
		_w26707_,
		_w26708_
	);
	LUT2 #(
		.INIT('h1)
	) name22662 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR1_reg[9]/P0001 ,
		_w26709_
	);
	LUT2 #(
		.INIT('h8)
	) name22663 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		\sice_DBR1_reg[9]/P0001 ,
		_w26710_
	);
	LUT2 #(
		.INIT('h1)
	) name22664 (
		\sice_DMR1_reg[9]/NET0131 ,
		_w26709_,
		_w26711_
	);
	LUT2 #(
		.INIT('h4)
	) name22665 (
		_w26710_,
		_w26711_,
		_w26712_
	);
	LUT2 #(
		.INIT('h1)
	) name22666 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR1_reg[13]/P0001 ,
		_w26713_
	);
	LUT2 #(
		.INIT('h8)
	) name22667 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		\sice_DBR1_reg[13]/P0001 ,
		_w26714_
	);
	LUT2 #(
		.INIT('h1)
	) name22668 (
		\sice_DMR1_reg[13]/NET0131 ,
		_w26713_,
		_w26715_
	);
	LUT2 #(
		.INIT('h4)
	) name22669 (
		_w26714_,
		_w26715_,
		_w26716_
	);
	LUT2 #(
		.INIT('h1)
	) name22670 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[17]/P0001 ,
		_w26717_
	);
	LUT2 #(
		.INIT('h8)
	) name22671 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[17]/P0001 ,
		_w26718_
	);
	LUT2 #(
		.INIT('h1)
	) name22672 (
		_w26717_,
		_w26718_,
		_w26719_
	);
	LUT2 #(
		.INIT('h2)
	) name22673 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[15]/P0001 ,
		_w26720_
	);
	LUT2 #(
		.INIT('h4)
	) name22674 (
		\core_c_psq_DMOVL_reg_DO_reg[1]/NET0131 ,
		\sice_DBR1_reg[15]/P0001 ,
		_w26721_
	);
	LUT2 #(
		.INIT('h1)
	) name22675 (
		_w26720_,
		_w26721_,
		_w26722_
	);
	LUT2 #(
		.INIT('h1)
	) name22676 (
		\sice_DMR1_reg[15]/NET0131 ,
		_w26722_,
		_w26723_
	);
	LUT2 #(
		.INIT('h1)
	) name22677 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[14]/P0001 ,
		_w26724_
	);
	LUT2 #(
		.INIT('h8)
	) name22678 (
		\core_c_psq_DMOVL_reg_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[14]/P0001 ,
		_w26725_
	);
	LUT2 #(
		.INIT('h1)
	) name22679 (
		\sice_DMR1_reg[14]/NET0131 ,
		_w26724_,
		_w26726_
	);
	LUT2 #(
		.INIT('h4)
	) name22680 (
		_w26725_,
		_w26726_,
		_w26727_
	);
	LUT2 #(
		.INIT('h2)
	) name22681 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[3]/P0001 ,
		_w26728_
	);
	LUT2 #(
		.INIT('h4)
	) name22682 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		\sice_DBR1_reg[3]/P0001 ,
		_w26729_
	);
	LUT2 #(
		.INIT('h1)
	) name22683 (
		_w26728_,
		_w26729_,
		_w26730_
	);
	LUT2 #(
		.INIT('h1)
	) name22684 (
		\sice_DMR1_reg[3]/NET0131 ,
		_w26730_,
		_w26731_
	);
	LUT2 #(
		.INIT('h1)
	) name22685 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR1_reg[8]/P0001 ,
		_w26732_
	);
	LUT2 #(
		.INIT('h8)
	) name22686 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		\sice_DBR1_reg[8]/P0001 ,
		_w26733_
	);
	LUT2 #(
		.INIT('h1)
	) name22687 (
		\sice_DMR1_reg[8]/NET0131 ,
		_w26732_,
		_w26734_
	);
	LUT2 #(
		.INIT('h4)
	) name22688 (
		_w26733_,
		_w26734_,
		_w26735_
	);
	LUT2 #(
		.INIT('h1)
	) name22689 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR1_reg[4]/P0001 ,
		_w26736_
	);
	LUT2 #(
		.INIT('h8)
	) name22690 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		\sice_DBR1_reg[4]/P0001 ,
		_w26737_
	);
	LUT2 #(
		.INIT('h1)
	) name22691 (
		\sice_DMR1_reg[4]/NET0131 ,
		_w26736_,
		_w26738_
	);
	LUT2 #(
		.INIT('h4)
	) name22692 (
		_w26737_,
		_w26738_,
		_w26739_
	);
	LUT2 #(
		.INIT('h2)
	) name22693 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR1_reg[6]/P0001 ,
		_w26740_
	);
	LUT2 #(
		.INIT('h4)
	) name22694 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		\sice_DBR1_reg[6]/P0001 ,
		_w26741_
	);
	LUT2 #(
		.INIT('h1)
	) name22695 (
		_w26740_,
		_w26741_,
		_w26742_
	);
	LUT2 #(
		.INIT('h1)
	) name22696 (
		\sice_DMR1_reg[6]/NET0131 ,
		_w26742_,
		_w26743_
	);
	LUT2 #(
		.INIT('h8)
	) name22697 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w26405_,
		_w26744_
	);
	LUT2 #(
		.INIT('h1)
	) name22698 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[0]/P0001 ,
		_w26745_
	);
	LUT2 #(
		.INIT('h8)
	) name22699 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		\sice_DBR1_reg[0]/P0001 ,
		_w26746_
	);
	LUT2 #(
		.INIT('h1)
	) name22700 (
		\sice_DMR1_reg[0]/NET0131 ,
		_w26745_,
		_w26747_
	);
	LUT2 #(
		.INIT('h4)
	) name22701 (
		_w26746_,
		_w26747_,
		_w26748_
	);
	LUT2 #(
		.INIT('h8)
	) name22702 (
		\sice_DBR1_reg[18]/P0001 ,
		\sice_DMR1_reg[17]/NET0131 ,
		_w26749_
	);
	LUT2 #(
		.INIT('h8)
	) name22703 (
		_w26631_,
		_w26749_,
		_w26750_
	);
	LUT2 #(
		.INIT('h4)
	) name22704 (
		_w26682_,
		_w26750_,
		_w26751_
	);
	LUT2 #(
		.INIT('h1)
	) name22705 (
		_w26683_,
		_w26704_,
		_w26752_
	);
	LUT2 #(
		.INIT('h1)
	) name22706 (
		_w26719_,
		_w26744_,
		_w26753_
	);
	LUT2 #(
		.INIT('h8)
	) name22707 (
		_w26752_,
		_w26753_,
		_w26754_
	);
	LUT2 #(
		.INIT('h4)
	) name22708 (
		_w26687_,
		_w26751_,
		_w26755_
	);
	LUT2 #(
		.INIT('h1)
	) name22709 (
		_w26691_,
		_w26695_,
		_w26756_
	);
	LUT2 #(
		.INIT('h1)
	) name22710 (
		_w26699_,
		_w26703_,
		_w26757_
	);
	LUT2 #(
		.INIT('h1)
	) name22711 (
		_w26708_,
		_w26712_,
		_w26758_
	);
	LUT2 #(
		.INIT('h1)
	) name22712 (
		_w26716_,
		_w26723_,
		_w26759_
	);
	LUT2 #(
		.INIT('h1)
	) name22713 (
		_w26727_,
		_w26731_,
		_w26760_
	);
	LUT2 #(
		.INIT('h1)
	) name22714 (
		_w26735_,
		_w26739_,
		_w26761_
	);
	LUT2 #(
		.INIT('h1)
	) name22715 (
		_w26743_,
		_w26748_,
		_w26762_
	);
	LUT2 #(
		.INIT('h8)
	) name22716 (
		_w26761_,
		_w26762_,
		_w26763_
	);
	LUT2 #(
		.INIT('h8)
	) name22717 (
		_w26759_,
		_w26760_,
		_w26764_
	);
	LUT2 #(
		.INIT('h8)
	) name22718 (
		_w26757_,
		_w26758_,
		_w26765_
	);
	LUT2 #(
		.INIT('h8)
	) name22719 (
		_w26755_,
		_w26756_,
		_w26766_
	);
	LUT2 #(
		.INIT('h8)
	) name22720 (
		_w26754_,
		_w26766_,
		_w26767_
	);
	LUT2 #(
		.INIT('h8)
	) name22721 (
		_w26764_,
		_w26765_,
		_w26768_
	);
	LUT2 #(
		.INIT('h8)
	) name22722 (
		_w26763_,
		_w26768_,
		_w26769_
	);
	LUT2 #(
		.INIT('h8)
	) name22723 (
		_w26767_,
		_w26769_,
		_w26770_
	);
	LUT2 #(
		.INIT('h1)
	) name22724 (
		_w26681_,
		_w26770_,
		_w26771_
	);
	LUT2 #(
		.INIT('h4)
	) name22725 (
		_w26591_,
		_w26771_,
		_w26772_
	);
	LUT2 #(
		.INIT('h2)
	) name22726 (
		\sice_ITR_reg[2]/NET0131 ,
		_w26772_,
		_w26773_
	);
	LUT2 #(
		.INIT('h2)
	) name22727 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\sice_IBR1_reg[16]/P0001 ,
		_w26774_
	);
	LUT2 #(
		.INIT('h4)
	) name22728 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\sice_IBR1_reg[16]/P0001 ,
		_w26775_
	);
	LUT2 #(
		.INIT('h1)
	) name22729 (
		_w26774_,
		_w26775_,
		_w26776_
	);
	LUT2 #(
		.INIT('h1)
	) name22730 (
		\sice_IMR1_reg[16]/NET0131 ,
		_w26776_,
		_w26777_
	);
	LUT2 #(
		.INIT('h2)
	) name22731 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		\sice_IBR1_reg[13]/P0001 ,
		_w26778_
	);
	LUT2 #(
		.INIT('h4)
	) name22732 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		\sice_IBR1_reg[13]/P0001 ,
		_w26779_
	);
	LUT2 #(
		.INIT('h1)
	) name22733 (
		_w26778_,
		_w26779_,
		_w26780_
	);
	LUT2 #(
		.INIT('h1)
	) name22734 (
		\sice_IMR1_reg[13]/NET0131 ,
		_w26780_,
		_w26781_
	);
	LUT2 #(
		.INIT('h1)
	) name22735 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		\sice_IBR1_reg[6]/P0001 ,
		_w26782_
	);
	LUT2 #(
		.INIT('h8)
	) name22736 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		\sice_IBR1_reg[6]/P0001 ,
		_w26783_
	);
	LUT2 #(
		.INIT('h1)
	) name22737 (
		\sice_IMR1_reg[6]/NET0131 ,
		_w26782_,
		_w26784_
	);
	LUT2 #(
		.INIT('h4)
	) name22738 (
		_w26783_,
		_w26784_,
		_w26785_
	);
	LUT2 #(
		.INIT('h2)
	) name22739 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		\sice_IBR1_reg[12]/P0001 ,
		_w26786_
	);
	LUT2 #(
		.INIT('h4)
	) name22740 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		\sice_IBR1_reg[12]/P0001 ,
		_w26787_
	);
	LUT2 #(
		.INIT('h1)
	) name22741 (
		_w26786_,
		_w26787_,
		_w26788_
	);
	LUT2 #(
		.INIT('h1)
	) name22742 (
		\sice_IMR1_reg[12]/NET0131 ,
		_w26788_,
		_w26789_
	);
	LUT2 #(
		.INIT('h1)
	) name22743 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		\sice_IBR1_reg[8]/P0001 ,
		_w26790_
	);
	LUT2 #(
		.INIT('h8)
	) name22744 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		\sice_IBR1_reg[8]/P0001 ,
		_w26791_
	);
	LUT2 #(
		.INIT('h1)
	) name22745 (
		\sice_IMR1_reg[8]/NET0131 ,
		_w26790_,
		_w26792_
	);
	LUT2 #(
		.INIT('h4)
	) name22746 (
		_w26791_,
		_w26792_,
		_w26793_
	);
	LUT2 #(
		.INIT('h1)
	) name22747 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		\sice_IBR1_reg[5]/P0001 ,
		_w26794_
	);
	LUT2 #(
		.INIT('h8)
	) name22748 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		\sice_IBR1_reg[5]/P0001 ,
		_w26795_
	);
	LUT2 #(
		.INIT('h1)
	) name22749 (
		\sice_IMR1_reg[5]/NET0131 ,
		_w26794_,
		_w26796_
	);
	LUT2 #(
		.INIT('h4)
	) name22750 (
		_w26795_,
		_w26796_,
		_w26797_
	);
	LUT2 #(
		.INIT('h2)
	) name22751 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		\sice_IBR1_reg[10]/P0001 ,
		_w26798_
	);
	LUT2 #(
		.INIT('h4)
	) name22752 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		\sice_IBR1_reg[10]/P0001 ,
		_w26799_
	);
	LUT2 #(
		.INIT('h1)
	) name22753 (
		_w26798_,
		_w26799_,
		_w26800_
	);
	LUT2 #(
		.INIT('h1)
	) name22754 (
		\sice_IMR1_reg[10]/NET0131 ,
		_w26800_,
		_w26801_
	);
	LUT2 #(
		.INIT('h1)
	) name22755 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\sice_IBR1_reg[15]/P0001 ,
		_w26802_
	);
	LUT2 #(
		.INIT('h8)
	) name22756 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\sice_IBR1_reg[15]/P0001 ,
		_w26803_
	);
	LUT2 #(
		.INIT('h1)
	) name22757 (
		\sice_IMR1_reg[15]/NET0131 ,
		_w26802_,
		_w26804_
	);
	LUT2 #(
		.INIT('h4)
	) name22758 (
		_w26803_,
		_w26804_,
		_w26805_
	);
	LUT2 #(
		.INIT('h2)
	) name22759 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		\sice_IBR1_reg[7]/P0001 ,
		_w26806_
	);
	LUT2 #(
		.INIT('h4)
	) name22760 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		\sice_IBR1_reg[7]/P0001 ,
		_w26807_
	);
	LUT2 #(
		.INIT('h1)
	) name22761 (
		_w26806_,
		_w26807_,
		_w26808_
	);
	LUT2 #(
		.INIT('h1)
	) name22762 (
		\sice_IMR1_reg[7]/NET0131 ,
		_w26808_,
		_w26809_
	);
	LUT2 #(
		.INIT('h1)
	) name22763 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		\sice_IBR1_reg[1]/P0001 ,
		_w26810_
	);
	LUT2 #(
		.INIT('h8)
	) name22764 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		\sice_IBR1_reg[1]/P0001 ,
		_w26811_
	);
	LUT2 #(
		.INIT('h1)
	) name22765 (
		\sice_IMR1_reg[1]/NET0131 ,
		_w26810_,
		_w26812_
	);
	LUT2 #(
		.INIT('h4)
	) name22766 (
		_w26811_,
		_w26812_,
		_w26813_
	);
	LUT2 #(
		.INIT('h1)
	) name22767 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		\sice_IBR1_reg[4]/P0001 ,
		_w26814_
	);
	LUT2 #(
		.INIT('h8)
	) name22768 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		\sice_IBR1_reg[4]/P0001 ,
		_w26815_
	);
	LUT2 #(
		.INIT('h1)
	) name22769 (
		\sice_IMR1_reg[4]/NET0131 ,
		_w26814_,
		_w26816_
	);
	LUT2 #(
		.INIT('h4)
	) name22770 (
		_w26815_,
		_w26816_,
		_w26817_
	);
	LUT2 #(
		.INIT('h1)
	) name22771 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		\sice_IBR1_reg[11]/P0001 ,
		_w26818_
	);
	LUT2 #(
		.INIT('h8)
	) name22772 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		\sice_IBR1_reg[11]/P0001 ,
		_w26819_
	);
	LUT2 #(
		.INIT('h1)
	) name22773 (
		\sice_IMR1_reg[11]/NET0131 ,
		_w26818_,
		_w26820_
	);
	LUT2 #(
		.INIT('h4)
	) name22774 (
		_w26819_,
		_w26820_,
		_w26821_
	);
	LUT2 #(
		.INIT('h2)
	) name22775 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\sice_IBR1_reg[14]/P0001 ,
		_w26822_
	);
	LUT2 #(
		.INIT('h4)
	) name22776 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\sice_IBR1_reg[14]/P0001 ,
		_w26823_
	);
	LUT2 #(
		.INIT('h1)
	) name22777 (
		_w26822_,
		_w26823_,
		_w26824_
	);
	LUT2 #(
		.INIT('h1)
	) name22778 (
		\sice_IMR1_reg[14]/NET0131 ,
		_w26824_,
		_w26825_
	);
	LUT2 #(
		.INIT('h2)
	) name22779 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		\sice_IBR1_reg[3]/P0001 ,
		_w26826_
	);
	LUT2 #(
		.INIT('h4)
	) name22780 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		\sice_IBR1_reg[3]/P0001 ,
		_w26827_
	);
	LUT2 #(
		.INIT('h1)
	) name22781 (
		_w26826_,
		_w26827_,
		_w26828_
	);
	LUT2 #(
		.INIT('h1)
	) name22782 (
		\sice_IMR1_reg[3]/NET0131 ,
		_w26828_,
		_w26829_
	);
	LUT2 #(
		.INIT('h1)
	) name22783 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		\sice_IBR1_reg[0]/P0001 ,
		_w26830_
	);
	LUT2 #(
		.INIT('h8)
	) name22784 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		\sice_IBR1_reg[0]/P0001 ,
		_w26831_
	);
	LUT2 #(
		.INIT('h1)
	) name22785 (
		\sice_IMR1_reg[0]/NET0131 ,
		_w26830_,
		_w26832_
	);
	LUT2 #(
		.INIT('h4)
	) name22786 (
		_w26831_,
		_w26832_,
		_w26833_
	);
	LUT2 #(
		.INIT('h2)
	) name22787 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		\sice_IBR1_reg[9]/P0001 ,
		_w26834_
	);
	LUT2 #(
		.INIT('h4)
	) name22788 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		\sice_IBR1_reg[9]/P0001 ,
		_w26835_
	);
	LUT2 #(
		.INIT('h1)
	) name22789 (
		_w26834_,
		_w26835_,
		_w26836_
	);
	LUT2 #(
		.INIT('h1)
	) name22790 (
		\sice_IMR1_reg[9]/NET0131 ,
		_w26836_,
		_w26837_
	);
	LUT2 #(
		.INIT('h1)
	) name22791 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		\sice_IBR1_reg[2]/P0001 ,
		_w26838_
	);
	LUT2 #(
		.INIT('h8)
	) name22792 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		\sice_IBR1_reg[2]/P0001 ,
		_w26839_
	);
	LUT2 #(
		.INIT('h1)
	) name22793 (
		\sice_IMR1_reg[2]/NET0131 ,
		_w26838_,
		_w26840_
	);
	LUT2 #(
		.INIT('h4)
	) name22794 (
		_w26839_,
		_w26840_,
		_w26841_
	);
	LUT2 #(
		.INIT('h2)
	) name22795 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\sice_IBR1_reg[17]/P0001 ,
		_w26842_
	);
	LUT2 #(
		.INIT('h4)
	) name22796 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\sice_IBR1_reg[17]/P0001 ,
		_w26843_
	);
	LUT2 #(
		.INIT('h8)
	) name22797 (
		\sice_IMR1_reg[17]/NET0131 ,
		\sice_ITR_reg[1]/NET0131 ,
		_w26844_
	);
	LUT2 #(
		.INIT('h4)
	) name22798 (
		_w26842_,
		_w26844_,
		_w26845_
	);
	LUT2 #(
		.INIT('h4)
	) name22799 (
		_w26843_,
		_w26845_,
		_w26846_
	);
	LUT2 #(
		.INIT('h4)
	) name22800 (
		_w26777_,
		_w26846_,
		_w26847_
	);
	LUT2 #(
		.INIT('h1)
	) name22801 (
		_w26781_,
		_w26785_,
		_w26848_
	);
	LUT2 #(
		.INIT('h1)
	) name22802 (
		_w26789_,
		_w26793_,
		_w26849_
	);
	LUT2 #(
		.INIT('h1)
	) name22803 (
		_w26797_,
		_w26801_,
		_w26850_
	);
	LUT2 #(
		.INIT('h1)
	) name22804 (
		_w26805_,
		_w26809_,
		_w26851_
	);
	LUT2 #(
		.INIT('h1)
	) name22805 (
		_w26813_,
		_w26817_,
		_w26852_
	);
	LUT2 #(
		.INIT('h1)
	) name22806 (
		_w26821_,
		_w26825_,
		_w26853_
	);
	LUT2 #(
		.INIT('h1)
	) name22807 (
		_w26829_,
		_w26833_,
		_w26854_
	);
	LUT2 #(
		.INIT('h1)
	) name22808 (
		_w26837_,
		_w26841_,
		_w26855_
	);
	LUT2 #(
		.INIT('h8)
	) name22809 (
		_w26854_,
		_w26855_,
		_w26856_
	);
	LUT2 #(
		.INIT('h8)
	) name22810 (
		_w26852_,
		_w26853_,
		_w26857_
	);
	LUT2 #(
		.INIT('h8)
	) name22811 (
		_w26850_,
		_w26851_,
		_w26858_
	);
	LUT2 #(
		.INIT('h8)
	) name22812 (
		_w26848_,
		_w26849_,
		_w26859_
	);
	LUT2 #(
		.INIT('h8)
	) name22813 (
		_w26847_,
		_w26859_,
		_w26860_
	);
	LUT2 #(
		.INIT('h8)
	) name22814 (
		_w26857_,
		_w26858_,
		_w26861_
	);
	LUT2 #(
		.INIT('h8)
	) name22815 (
		_w26856_,
		_w26861_,
		_w26862_
	);
	LUT2 #(
		.INIT('h8)
	) name22816 (
		_w26860_,
		_w26862_,
		_w26863_
	);
	LUT2 #(
		.INIT('h2)
	) name22817 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		\sice_IBR2_reg[6]/P0001 ,
		_w26864_
	);
	LUT2 #(
		.INIT('h4)
	) name22818 (
		\core_c_psq_DRA_reg[6]/P0001 ,
		\sice_IBR2_reg[6]/P0001 ,
		_w26865_
	);
	LUT2 #(
		.INIT('h1)
	) name22819 (
		_w26864_,
		_w26865_,
		_w26866_
	);
	LUT2 #(
		.INIT('h1)
	) name22820 (
		\sice_IMR2_reg[6]/NET0131 ,
		_w26866_,
		_w26867_
	);
	LUT2 #(
		.INIT('h1)
	) name22821 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		\sice_IBR2_reg[12]/P0001 ,
		_w26868_
	);
	LUT2 #(
		.INIT('h8)
	) name22822 (
		\core_c_psq_DRA_reg[12]/P0001 ,
		\sice_IBR2_reg[12]/P0001 ,
		_w26869_
	);
	LUT2 #(
		.INIT('h1)
	) name22823 (
		\sice_IMR2_reg[12]/NET0131 ,
		_w26868_,
		_w26870_
	);
	LUT2 #(
		.INIT('h4)
	) name22824 (
		_w26869_,
		_w26870_,
		_w26871_
	);
	LUT2 #(
		.INIT('h2)
	) name22825 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		\sice_IBR2_reg[9]/P0001 ,
		_w26872_
	);
	LUT2 #(
		.INIT('h4)
	) name22826 (
		\core_c_psq_DRA_reg[9]/P0001 ,
		\sice_IBR2_reg[9]/P0001 ,
		_w26873_
	);
	LUT2 #(
		.INIT('h1)
	) name22827 (
		_w26872_,
		_w26873_,
		_w26874_
	);
	LUT2 #(
		.INIT('h1)
	) name22828 (
		\sice_IMR2_reg[9]/NET0131 ,
		_w26874_,
		_w26875_
	);
	LUT2 #(
		.INIT('h1)
	) name22829 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		\sice_IBR2_reg[4]/P0001 ,
		_w26876_
	);
	LUT2 #(
		.INIT('h8)
	) name22830 (
		\core_c_psq_DRA_reg[4]/P0001 ,
		\sice_IBR2_reg[4]/P0001 ,
		_w26877_
	);
	LUT2 #(
		.INIT('h1)
	) name22831 (
		\sice_IMR2_reg[4]/NET0131 ,
		_w26876_,
		_w26878_
	);
	LUT2 #(
		.INIT('h4)
	) name22832 (
		_w26877_,
		_w26878_,
		_w26879_
	);
	LUT2 #(
		.INIT('h1)
	) name22833 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\sice_IBR2_reg[16]/P0001 ,
		_w26880_
	);
	LUT2 #(
		.INIT('h8)
	) name22834 (
		\core_c_psq_PMOVL_regl_DO_reg[2]/NET0131 ,
		\sice_IBR2_reg[16]/P0001 ,
		_w26881_
	);
	LUT2 #(
		.INIT('h1)
	) name22835 (
		\sice_IMR2_reg[16]/NET0131 ,
		_w26880_,
		_w26882_
	);
	LUT2 #(
		.INIT('h4)
	) name22836 (
		_w26881_,
		_w26882_,
		_w26883_
	);
	LUT2 #(
		.INIT('h2)
	) name22837 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		\sice_IBR2_reg[1]/P0001 ,
		_w26884_
	);
	LUT2 #(
		.INIT('h4)
	) name22838 (
		\core_c_psq_DRA_reg[1]/P0001 ,
		\sice_IBR2_reg[1]/P0001 ,
		_w26885_
	);
	LUT2 #(
		.INIT('h1)
	) name22839 (
		_w26884_,
		_w26885_,
		_w26886_
	);
	LUT2 #(
		.INIT('h1)
	) name22840 (
		\sice_IMR2_reg[1]/NET0131 ,
		_w26886_,
		_w26887_
	);
	LUT2 #(
		.INIT('h2)
	) name22841 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		\sice_IBR2_reg[2]/P0001 ,
		_w26888_
	);
	LUT2 #(
		.INIT('h4)
	) name22842 (
		\core_c_psq_DRA_reg[2]/P0001 ,
		\sice_IBR2_reg[2]/P0001 ,
		_w26889_
	);
	LUT2 #(
		.INIT('h1)
	) name22843 (
		_w26888_,
		_w26889_,
		_w26890_
	);
	LUT2 #(
		.INIT('h1)
	) name22844 (
		\sice_IMR2_reg[2]/NET0131 ,
		_w26890_,
		_w26891_
	);
	LUT2 #(
		.INIT('h2)
	) name22845 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		\sice_IBR2_reg[0]/P0001 ,
		_w26892_
	);
	LUT2 #(
		.INIT('h4)
	) name22846 (
		\core_c_psq_DRA_reg[0]/P0001 ,
		\sice_IBR2_reg[0]/P0001 ,
		_w26893_
	);
	LUT2 #(
		.INIT('h1)
	) name22847 (
		_w26892_,
		_w26893_,
		_w26894_
	);
	LUT2 #(
		.INIT('h1)
	) name22848 (
		\sice_IMR2_reg[0]/NET0131 ,
		_w26894_,
		_w26895_
	);
	LUT2 #(
		.INIT('h1)
	) name22849 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		\sice_IBR2_reg[8]/P0001 ,
		_w26896_
	);
	LUT2 #(
		.INIT('h8)
	) name22850 (
		\core_c_psq_DRA_reg[8]/P0001 ,
		\sice_IBR2_reg[8]/P0001 ,
		_w26897_
	);
	LUT2 #(
		.INIT('h1)
	) name22851 (
		\sice_IMR2_reg[8]/NET0131 ,
		_w26896_,
		_w26898_
	);
	LUT2 #(
		.INIT('h4)
	) name22852 (
		_w26897_,
		_w26898_,
		_w26899_
	);
	LUT2 #(
		.INIT('h2)
	) name22853 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		\sice_IBR2_reg[13]/P0001 ,
		_w26900_
	);
	LUT2 #(
		.INIT('h4)
	) name22854 (
		\core_c_psq_DRA_reg[13]/P0001 ,
		\sice_IBR2_reg[13]/P0001 ,
		_w26901_
	);
	LUT2 #(
		.INIT('h1)
	) name22855 (
		_w26900_,
		_w26901_,
		_w26902_
	);
	LUT2 #(
		.INIT('h1)
	) name22856 (
		\sice_IMR2_reg[13]/NET0131 ,
		_w26902_,
		_w26903_
	);
	LUT2 #(
		.INIT('h1)
	) name22857 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		\sice_IBR2_reg[5]/P0001 ,
		_w26904_
	);
	LUT2 #(
		.INIT('h8)
	) name22858 (
		\core_c_psq_DRA_reg[5]/P0001 ,
		\sice_IBR2_reg[5]/P0001 ,
		_w26905_
	);
	LUT2 #(
		.INIT('h1)
	) name22859 (
		\sice_IMR2_reg[5]/NET0131 ,
		_w26904_,
		_w26906_
	);
	LUT2 #(
		.INIT('h4)
	) name22860 (
		_w26905_,
		_w26906_,
		_w26907_
	);
	LUT2 #(
		.INIT('h1)
	) name22861 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\sice_IBR2_reg[14]/P0001 ,
		_w26908_
	);
	LUT2 #(
		.INIT('h8)
	) name22862 (
		\core_c_psq_PMOVL_regl_DO_reg[0]/NET0131 ,
		\sice_IBR2_reg[14]/P0001 ,
		_w26909_
	);
	LUT2 #(
		.INIT('h1)
	) name22863 (
		\sice_IMR2_reg[14]/NET0131 ,
		_w26908_,
		_w26910_
	);
	LUT2 #(
		.INIT('h4)
	) name22864 (
		_w26909_,
		_w26910_,
		_w26911_
	);
	LUT2 #(
		.INIT('h2)
	) name22865 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		\sice_IBR2_reg[7]/P0001 ,
		_w26912_
	);
	LUT2 #(
		.INIT('h4)
	) name22866 (
		\core_c_psq_DRA_reg[7]/P0001 ,
		\sice_IBR2_reg[7]/P0001 ,
		_w26913_
	);
	LUT2 #(
		.INIT('h1)
	) name22867 (
		_w26912_,
		_w26913_,
		_w26914_
	);
	LUT2 #(
		.INIT('h1)
	) name22868 (
		\sice_IMR2_reg[7]/NET0131 ,
		_w26914_,
		_w26915_
	);
	LUT2 #(
		.INIT('h2)
	) name22869 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		\sice_IBR2_reg[11]/P0001 ,
		_w26916_
	);
	LUT2 #(
		.INIT('h4)
	) name22870 (
		\core_c_psq_DRA_reg[11]/P0001 ,
		\sice_IBR2_reg[11]/P0001 ,
		_w26917_
	);
	LUT2 #(
		.INIT('h1)
	) name22871 (
		_w26916_,
		_w26917_,
		_w26918_
	);
	LUT2 #(
		.INIT('h1)
	) name22872 (
		\sice_IMR2_reg[11]/NET0131 ,
		_w26918_,
		_w26919_
	);
	LUT2 #(
		.INIT('h1)
	) name22873 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		\sice_IBR2_reg[3]/P0001 ,
		_w26920_
	);
	LUT2 #(
		.INIT('h8)
	) name22874 (
		\core_c_psq_DRA_reg[3]/P0001 ,
		\sice_IBR2_reg[3]/P0001 ,
		_w26921_
	);
	LUT2 #(
		.INIT('h1)
	) name22875 (
		\sice_IMR2_reg[3]/NET0131 ,
		_w26920_,
		_w26922_
	);
	LUT2 #(
		.INIT('h4)
	) name22876 (
		_w26921_,
		_w26922_,
		_w26923_
	);
	LUT2 #(
		.INIT('h2)
	) name22877 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\sice_IBR2_reg[15]/P0001 ,
		_w26924_
	);
	LUT2 #(
		.INIT('h4)
	) name22878 (
		\core_c_psq_PMOVL_regl_DO_reg[1]/NET0131 ,
		\sice_IBR2_reg[15]/P0001 ,
		_w26925_
	);
	LUT2 #(
		.INIT('h1)
	) name22879 (
		_w26924_,
		_w26925_,
		_w26926_
	);
	LUT2 #(
		.INIT('h1)
	) name22880 (
		\sice_IMR2_reg[15]/NET0131 ,
		_w26926_,
		_w26927_
	);
	LUT2 #(
		.INIT('h1)
	) name22881 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		\sice_IBR2_reg[10]/P0001 ,
		_w26928_
	);
	LUT2 #(
		.INIT('h8)
	) name22882 (
		\core_c_psq_DRA_reg[10]/P0001 ,
		\sice_IBR2_reg[10]/P0001 ,
		_w26929_
	);
	LUT2 #(
		.INIT('h1)
	) name22883 (
		\sice_IMR2_reg[10]/NET0131 ,
		_w26928_,
		_w26930_
	);
	LUT2 #(
		.INIT('h4)
	) name22884 (
		_w26929_,
		_w26930_,
		_w26931_
	);
	LUT2 #(
		.INIT('h2)
	) name22885 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\sice_IBR2_reg[17]/P0001 ,
		_w26932_
	);
	LUT2 #(
		.INIT('h4)
	) name22886 (
		\core_c_psq_PMOVL_regl_DO_reg[3]/NET0131 ,
		\sice_IBR2_reg[17]/P0001 ,
		_w26933_
	);
	LUT2 #(
		.INIT('h8)
	) name22887 (
		\sice_IMR2_reg[17]/NET0131 ,
		\sice_ITR_reg[1]/NET0131 ,
		_w26934_
	);
	LUT2 #(
		.INIT('h4)
	) name22888 (
		_w26932_,
		_w26934_,
		_w26935_
	);
	LUT2 #(
		.INIT('h4)
	) name22889 (
		_w26933_,
		_w26935_,
		_w26936_
	);
	LUT2 #(
		.INIT('h4)
	) name22890 (
		_w26867_,
		_w26936_,
		_w26937_
	);
	LUT2 #(
		.INIT('h1)
	) name22891 (
		_w26871_,
		_w26875_,
		_w26938_
	);
	LUT2 #(
		.INIT('h1)
	) name22892 (
		_w26879_,
		_w26883_,
		_w26939_
	);
	LUT2 #(
		.INIT('h1)
	) name22893 (
		_w26887_,
		_w26891_,
		_w26940_
	);
	LUT2 #(
		.INIT('h1)
	) name22894 (
		_w26895_,
		_w26899_,
		_w26941_
	);
	LUT2 #(
		.INIT('h1)
	) name22895 (
		_w26903_,
		_w26907_,
		_w26942_
	);
	LUT2 #(
		.INIT('h1)
	) name22896 (
		_w26911_,
		_w26915_,
		_w26943_
	);
	LUT2 #(
		.INIT('h1)
	) name22897 (
		_w26919_,
		_w26923_,
		_w26944_
	);
	LUT2 #(
		.INIT('h1)
	) name22898 (
		_w26927_,
		_w26931_,
		_w26945_
	);
	LUT2 #(
		.INIT('h8)
	) name22899 (
		_w26944_,
		_w26945_,
		_w26946_
	);
	LUT2 #(
		.INIT('h8)
	) name22900 (
		_w26942_,
		_w26943_,
		_w26947_
	);
	LUT2 #(
		.INIT('h8)
	) name22901 (
		_w26940_,
		_w26941_,
		_w26948_
	);
	LUT2 #(
		.INIT('h8)
	) name22902 (
		_w26938_,
		_w26939_,
		_w26949_
	);
	LUT2 #(
		.INIT('h8)
	) name22903 (
		_w26937_,
		_w26949_,
		_w26950_
	);
	LUT2 #(
		.INIT('h8)
	) name22904 (
		_w26947_,
		_w26948_,
		_w26951_
	);
	LUT2 #(
		.INIT('h8)
	) name22905 (
		_w26946_,
		_w26951_,
		_w26952_
	);
	LUT2 #(
		.INIT('h8)
	) name22906 (
		_w26950_,
		_w26952_,
		_w26953_
	);
	LUT2 #(
		.INIT('h1)
	) name22907 (
		_w26402_,
		_w26404_,
		_w26954_
	);
	LUT2 #(
		.INIT('h4)
	) name22908 (
		_w26863_,
		_w26954_,
		_w26955_
	);
	LUT2 #(
		.INIT('h4)
	) name22909 (
		_w26953_,
		_w26955_,
		_w26956_
	);
	LUT2 #(
		.INIT('h4)
	) name22910 (
		_w26773_,
		_w26956_,
		_w26957_
	);
	LUT2 #(
		.INIT('h1)
	) name22911 (
		_w4093_,
		_w26957_,
		_w26958_
	);
	LUT2 #(
		.INIT('h8)
	) name22912 (
		_w11741_,
		_w26958_,
		_w26959_
	);
	LUT2 #(
		.INIT('h1)
	) name22913 (
		\sice_HALT_E_reg/P0001 ,
		_w26959_,
		_w26960_
	);
	LUT2 #(
		.INIT('h8)
	) name22914 (
		_w12234_,
		_w23717_,
		_w26961_
	);
	LUT2 #(
		.INIT('h4)
	) name22915 (
		_w26960_,
		_w26961_,
		_w26962_
	);
	LUT2 #(
		.INIT('h8)
	) name22916 (
		_w26377_,
		_w26390_,
		_w26963_
	);
	LUT2 #(
		.INIT('h2)
	) name22917 (
		_w26388_,
		_w26391_,
		_w26964_
	);
	LUT2 #(
		.INIT('h1)
	) name22918 (
		_w26389_,
		_w26963_,
		_w26965_
	);
	LUT2 #(
		.INIT('h4)
	) name22919 (
		_w26964_,
		_w26965_,
		_w26966_
	);
	LUT2 #(
		.INIT('h2)
	) name22920 (
		\sice_UpdDR_sd1_reg/P0001 ,
		\sice_UpdDR_sd2_reg/P0001 ,
		_w26967_
	);
	LUT2 #(
		.INIT('h8)
	) name22921 (
		_w23408_,
		_w25033_,
		_w26968_
	);
	LUT2 #(
		.INIT('h8)
	) name22922 (
		_w26967_,
		_w26968_,
		_w26969_
	);
	LUT2 #(
		.INIT('h4)
	) name22923 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTIDR_E_reg/P0001 ,
		_w26970_
	);
	LUT2 #(
		.INIT('h1)
	) name22924 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w26970_,
		_w26971_
	);
	LUT2 #(
		.INIT('h1)
	) name22925 (
		_w5950_,
		_w26971_,
		_w26972_
	);
	LUT2 #(
		.INIT('h1)
	) name22926 (
		_w26969_,
		_w26972_,
		_w26973_
	);
	LUT2 #(
		.INIT('h8)
	) name22927 (
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w26973_,
		_w26974_
	);
	LUT2 #(
		.INIT('h8)
	) name22928 (
		_w12743_,
		_w26970_,
		_w26975_
	);
	LUT2 #(
		.INIT('h8)
	) name22929 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[15]/P0001 ,
		_w26976_
	);
	LUT2 #(
		.INIT('h1)
	) name22930 (
		\idma_CMo_oe3_reg/P0001 ,
		\idma_CMo_oe4_reg/P0001 ,
		_w26977_
	);
	LUT2 #(
		.INIT('h4)
	) name22931 (
		\idma_CMo_oe5_reg/P0001 ,
		_w26977_,
		_w26978_
	);
	LUT2 #(
		.INIT('h4)
	) name22932 (
		\idma_CMo_oe6_reg/P0001 ,
		_w26978_,
		_w26979_
	);
	LUT2 #(
		.INIT('h1)
	) name22933 (
		\idma_CM_oe_reg/P0001 ,
		\idma_CMo_oe0_reg/P0001 ,
		_w26980_
	);
	LUT2 #(
		.INIT('h4)
	) name22934 (
		\idma_CMo_oe7_reg/P0001 ,
		_w26980_,
		_w26981_
	);
	LUT2 #(
		.INIT('h8)
	) name22935 (
		_w26979_,
		_w26981_,
		_w26982_
	);
	LUT2 #(
		.INIT('h2)
	) name22936 (
		\idma_CMo_oe1_reg/P0001 ,
		\idma_CMo_oe2_reg/P0001 ,
		_w26983_
	);
	LUT2 #(
		.INIT('h8)
	) name22937 (
		_w26982_,
		_w26983_,
		_w26984_
	);
	LUT2 #(
		.INIT('h8)
	) name22938 (
		\CM_rd1[15]_pad ,
		_w26984_,
		_w26985_
	);
	LUT2 #(
		.INIT('h1)
	) name22939 (
		\idma_CMo_oe1_reg/P0001 ,
		\idma_CMo_oe2_reg/P0001 ,
		_w26986_
	);
	LUT2 #(
		.INIT('h8)
	) name22940 (
		_w26981_,
		_w26986_,
		_w26987_
	);
	LUT2 #(
		.INIT('h8)
	) name22941 (
		\idma_CMo_oe6_reg/P0001 ,
		_w26978_,
		_w26988_
	);
	LUT2 #(
		.INIT('h8)
	) name22942 (
		_w26987_,
		_w26988_,
		_w26989_
	);
	LUT2 #(
		.INIT('h8)
	) name22943 (
		\CM_rd6[15]_pad ,
		_w26989_,
		_w26990_
	);
	LUT2 #(
		.INIT('h8)
	) name22944 (
		_w26979_,
		_w26986_,
		_w26991_
	);
	LUT2 #(
		.INIT('h4)
	) name22945 (
		\idma_CM_oe_reg/P0001 ,
		\idma_CMo_oe0_reg/P0001 ,
		_w26992_
	);
	LUT2 #(
		.INIT('h4)
	) name22946 (
		\idma_CMo_oe7_reg/P0001 ,
		_w26992_,
		_w26993_
	);
	LUT2 #(
		.INIT('h8)
	) name22947 (
		_w26991_,
		_w26993_,
		_w26994_
	);
	LUT2 #(
		.INIT('h8)
	) name22948 (
		\CM_rd0[15]_pad ,
		_w26994_,
		_w26995_
	);
	LUT2 #(
		.INIT('h8)
	) name22949 (
		\idma_CMo_oe7_reg/P0001 ,
		_w26980_,
		_w26996_
	);
	LUT2 #(
		.INIT('h8)
	) name22950 (
		_w26991_,
		_w26996_,
		_w26997_
	);
	LUT2 #(
		.INIT('h8)
	) name22951 (
		\CM_rd7[15]_pad ,
		_w26997_,
		_w26998_
	);
	LUT2 #(
		.INIT('h4)
	) name22952 (
		\idma_CMo_oe1_reg/P0001 ,
		\idma_CMo_oe2_reg/P0001 ,
		_w26999_
	);
	LUT2 #(
		.INIT('h8)
	) name22953 (
		_w26982_,
		_w26999_,
		_w27000_
	);
	LUT2 #(
		.INIT('h8)
	) name22954 (
		\CM_rd2[15]_pad ,
		_w27000_,
		_w27001_
	);
	LUT2 #(
		.INIT('h4)
	) name22955 (
		\idma_CMo_oe6_reg/P0001 ,
		_w26987_,
		_w27002_
	);
	LUT2 #(
		.INIT('h8)
	) name22956 (
		\idma_CMo_oe5_reg/P0001 ,
		_w26977_,
		_w27003_
	);
	LUT2 #(
		.INIT('h8)
	) name22957 (
		_w27002_,
		_w27003_,
		_w27004_
	);
	LUT2 #(
		.INIT('h8)
	) name22958 (
		\CM_rd5[15]_pad ,
		_w27004_,
		_w27005_
	);
	LUT2 #(
		.INIT('h4)
	) name22959 (
		\idma_CMo_oe5_reg/P0001 ,
		_w27002_,
		_w27006_
	);
	LUT2 #(
		.INIT('h4)
	) name22960 (
		\idma_CMo_oe3_reg/P0001 ,
		\idma_CMo_oe4_reg/P0001 ,
		_w27007_
	);
	LUT2 #(
		.INIT('h8)
	) name22961 (
		_w27006_,
		_w27007_,
		_w27008_
	);
	LUT2 #(
		.INIT('h8)
	) name22962 (
		\CM_rd4[15]_pad ,
		_w27008_,
		_w27009_
	);
	LUT2 #(
		.INIT('h2)
	) name22963 (
		\idma_CMo_oe3_reg/P0001 ,
		\idma_CMo_oe4_reg/P0001 ,
		_w27010_
	);
	LUT2 #(
		.INIT('h8)
	) name22964 (
		_w27006_,
		_w27010_,
		_w27011_
	);
	LUT2 #(
		.INIT('h1)
	) name22965 (
		_w26984_,
		_w26989_,
		_w27012_
	);
	LUT2 #(
		.INIT('h1)
	) name22966 (
		_w26994_,
		_w26997_,
		_w27013_
	);
	LUT2 #(
		.INIT('h1)
	) name22967 (
		_w27000_,
		_w27004_,
		_w27014_
	);
	LUT2 #(
		.INIT('h8)
	) name22968 (
		_w27013_,
		_w27014_,
		_w27015_
	);
	LUT2 #(
		.INIT('h4)
	) name22969 (
		_w27008_,
		_w27012_,
		_w27016_
	);
	LUT2 #(
		.INIT('h4)
	) name22970 (
		_w27011_,
		_w27016_,
		_w27017_
	);
	LUT2 #(
		.INIT('h8)
	) name22971 (
		_w27015_,
		_w27017_,
		_w27018_
	);
	LUT2 #(
		.INIT('h8)
	) name22972 (
		\CM_rdm[15]_pad ,
		_w27018_,
		_w27019_
	);
	LUT2 #(
		.INIT('h8)
	) name22973 (
		\CM_rd3[15]_pad ,
		_w27011_,
		_w27020_
	);
	LUT2 #(
		.INIT('h1)
	) name22974 (
		_w26985_,
		_w26990_,
		_w27021_
	);
	LUT2 #(
		.INIT('h1)
	) name22975 (
		_w26995_,
		_w26998_,
		_w27022_
	);
	LUT2 #(
		.INIT('h1)
	) name22976 (
		_w27001_,
		_w27005_,
		_w27023_
	);
	LUT2 #(
		.INIT('h8)
	) name22977 (
		_w27022_,
		_w27023_,
		_w27024_
	);
	LUT2 #(
		.INIT('h4)
	) name22978 (
		_w27009_,
		_w27021_,
		_w27025_
	);
	LUT2 #(
		.INIT('h4)
	) name22979 (
		_w27020_,
		_w27025_,
		_w27026_
	);
	LUT2 #(
		.INIT('h8)
	) name22980 (
		_w27024_,
		_w27026_,
		_w27027_
	);
	LUT2 #(
		.INIT('h4)
	) name22981 (
		_w27019_,
		_w27027_,
		_w27028_
	);
	LUT2 #(
		.INIT('h1)
	) name22982 (
		\T_TMODE[1]_pad ,
		_w27028_,
		_w27029_
	);
	LUT2 #(
		.INIT('h1)
	) name22983 (
		_w26976_,
		_w27029_,
		_w27030_
	);
	LUT2 #(
		.INIT('h2)
	) name22984 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27030_,
		_w27031_
	);
	LUT2 #(
		.INIT('h1)
	) name22985 (
		_w26975_,
		_w27031_,
		_w27032_
	);
	LUT2 #(
		.INIT('h1)
	) name22986 (
		_w26973_,
		_w27032_,
		_w27033_
	);
	LUT2 #(
		.INIT('h8)
	) name22987 (
		\sice_SPC_reg[15]/P0001 ,
		_w26969_,
		_w27034_
	);
	LUT2 #(
		.INIT('h1)
	) name22988 (
		_w26974_,
		_w27034_,
		_w27035_
	);
	LUT2 #(
		.INIT('h4)
	) name22989 (
		_w27033_,
		_w27035_,
		_w27036_
	);
	LUT2 #(
		.INIT('h1)
	) name22990 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 ,
		_w19499_,
		_w27037_
	);
	LUT2 #(
		.INIT('h4)
	) name22991 (
		_w18974_,
		_w19499_,
		_w27038_
	);
	LUT2 #(
		.INIT('h2)
	) name22992 (
		_w19501_,
		_w27037_,
		_w27039_
	);
	LUT2 #(
		.INIT('h4)
	) name22993 (
		_w27038_,
		_w27039_,
		_w27040_
	);
	LUT2 #(
		.INIT('h2)
	) name22994 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[1]/P0001 ,
		_w19383_,
		_w27041_
	);
	LUT2 #(
		.INIT('h1)
	) name22995 (
		_w19508_,
		_w27041_,
		_w27042_
	);
	LUT2 #(
		.INIT('h4)
	) name22996 (
		_w27040_,
		_w27042_,
		_w27043_
	);
	LUT2 #(
		.INIT('h1)
	) name22997 (
		_w18262_,
		_w27043_,
		_w27044_
	);
	LUT2 #(
		.INIT('h4)
	) name22998 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19577_,
		_w27045_
	);
	LUT2 #(
		.INIT('h1)
	) name22999 (
		_w17638_,
		_w17665_,
		_w27046_
	);
	LUT2 #(
		.INIT('h4)
	) name23000 (
		_w16363_,
		_w17661_,
		_w27047_
	);
	LUT2 #(
		.INIT('h1)
	) name23001 (
		_w17670_,
		_w27047_,
		_w27048_
	);
	LUT2 #(
		.INIT('h4)
	) name23002 (
		_w27046_,
		_w27048_,
		_w27049_
	);
	LUT2 #(
		.INIT('h2)
	) name23003 (
		_w27046_,
		_w27048_,
		_w27050_
	);
	LUT2 #(
		.INIT('h1)
	) name23004 (
		_w27049_,
		_w27050_,
		_w27051_
	);
	LUT2 #(
		.INIT('h8)
	) name23005 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w27051_,
		_w27052_
	);
	LUT2 #(
		.INIT('h1)
	) name23006 (
		_w27045_,
		_w27052_,
		_w27053_
	);
	LUT2 #(
		.INIT('h2)
	) name23007 (
		_w18262_,
		_w27053_,
		_w27054_
	);
	LUT2 #(
		.INIT('h1)
	) name23008 (
		_w27044_,
		_w27054_,
		_w27055_
	);
	LUT2 #(
		.INIT('h8)
	) name23009 (
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w26973_,
		_w27056_
	);
	LUT2 #(
		.INIT('h8)
	) name23010 (
		_w12688_,
		_w26970_,
		_w27057_
	);
	LUT2 #(
		.INIT('h8)
	) name23011 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[14]/P0001 ,
		_w27058_
	);
	LUT2 #(
		.INIT('h8)
	) name23012 (
		\CM_rd1[14]_pad ,
		_w26984_,
		_w27059_
	);
	LUT2 #(
		.INIT('h8)
	) name23013 (
		\CM_rd6[14]_pad ,
		_w26989_,
		_w27060_
	);
	LUT2 #(
		.INIT('h8)
	) name23014 (
		\CM_rd0[14]_pad ,
		_w26994_,
		_w27061_
	);
	LUT2 #(
		.INIT('h8)
	) name23015 (
		\CM_rd7[14]_pad ,
		_w26997_,
		_w27062_
	);
	LUT2 #(
		.INIT('h8)
	) name23016 (
		\CM_rd2[14]_pad ,
		_w27000_,
		_w27063_
	);
	LUT2 #(
		.INIT('h8)
	) name23017 (
		\CM_rd5[14]_pad ,
		_w27004_,
		_w27064_
	);
	LUT2 #(
		.INIT('h8)
	) name23018 (
		\CM_rd4[14]_pad ,
		_w27008_,
		_w27065_
	);
	LUT2 #(
		.INIT('h8)
	) name23019 (
		\CM_rdm[14]_pad ,
		_w27018_,
		_w27066_
	);
	LUT2 #(
		.INIT('h8)
	) name23020 (
		\CM_rd3[14]_pad ,
		_w27011_,
		_w27067_
	);
	LUT2 #(
		.INIT('h1)
	) name23021 (
		_w27059_,
		_w27060_,
		_w27068_
	);
	LUT2 #(
		.INIT('h1)
	) name23022 (
		_w27061_,
		_w27062_,
		_w27069_
	);
	LUT2 #(
		.INIT('h1)
	) name23023 (
		_w27063_,
		_w27064_,
		_w27070_
	);
	LUT2 #(
		.INIT('h8)
	) name23024 (
		_w27069_,
		_w27070_,
		_w27071_
	);
	LUT2 #(
		.INIT('h4)
	) name23025 (
		_w27065_,
		_w27068_,
		_w27072_
	);
	LUT2 #(
		.INIT('h4)
	) name23026 (
		_w27067_,
		_w27072_,
		_w27073_
	);
	LUT2 #(
		.INIT('h8)
	) name23027 (
		_w27071_,
		_w27073_,
		_w27074_
	);
	LUT2 #(
		.INIT('h4)
	) name23028 (
		_w27066_,
		_w27074_,
		_w27075_
	);
	LUT2 #(
		.INIT('h1)
	) name23029 (
		\T_TMODE[1]_pad ,
		_w27075_,
		_w27076_
	);
	LUT2 #(
		.INIT('h1)
	) name23030 (
		_w27058_,
		_w27076_,
		_w27077_
	);
	LUT2 #(
		.INIT('h2)
	) name23031 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27077_,
		_w27078_
	);
	LUT2 #(
		.INIT('h1)
	) name23032 (
		_w27057_,
		_w27078_,
		_w27079_
	);
	LUT2 #(
		.INIT('h1)
	) name23033 (
		_w26973_,
		_w27079_,
		_w27080_
	);
	LUT2 #(
		.INIT('h8)
	) name23034 (
		\sice_SPC_reg[14]/P0001 ,
		_w26969_,
		_w27081_
	);
	LUT2 #(
		.INIT('h1)
	) name23035 (
		_w27056_,
		_w27081_,
		_w27082_
	);
	LUT2 #(
		.INIT('h4)
	) name23036 (
		_w27080_,
		_w27082_,
		_w27083_
	);
	LUT2 #(
		.INIT('h8)
	) name23037 (
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w26973_,
		_w27084_
	);
	LUT2 #(
		.INIT('h8)
	) name23038 (
		_w11265_,
		_w26970_,
		_w27085_
	);
	LUT2 #(
		.INIT('h8)
	) name23039 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[7]/P0001 ,
		_w27086_
	);
	LUT2 #(
		.INIT('h8)
	) name23040 (
		\CM_rd1[7]_pad ,
		_w26984_,
		_w27087_
	);
	LUT2 #(
		.INIT('h8)
	) name23041 (
		\CM_rd6[7]_pad ,
		_w26989_,
		_w27088_
	);
	LUT2 #(
		.INIT('h8)
	) name23042 (
		\CM_rd0[7]_pad ,
		_w26994_,
		_w27089_
	);
	LUT2 #(
		.INIT('h8)
	) name23043 (
		\CM_rd7[7]_pad ,
		_w26997_,
		_w27090_
	);
	LUT2 #(
		.INIT('h8)
	) name23044 (
		\CM_rd2[7]_pad ,
		_w27000_,
		_w27091_
	);
	LUT2 #(
		.INIT('h8)
	) name23045 (
		\CM_rd5[7]_pad ,
		_w27004_,
		_w27092_
	);
	LUT2 #(
		.INIT('h8)
	) name23046 (
		\CM_rd4[7]_pad ,
		_w27008_,
		_w27093_
	);
	LUT2 #(
		.INIT('h8)
	) name23047 (
		\CM_rdm[7]_pad ,
		_w27018_,
		_w27094_
	);
	LUT2 #(
		.INIT('h8)
	) name23048 (
		\CM_rd3[7]_pad ,
		_w27011_,
		_w27095_
	);
	LUT2 #(
		.INIT('h1)
	) name23049 (
		_w27087_,
		_w27088_,
		_w27096_
	);
	LUT2 #(
		.INIT('h1)
	) name23050 (
		_w27089_,
		_w27090_,
		_w27097_
	);
	LUT2 #(
		.INIT('h1)
	) name23051 (
		_w27091_,
		_w27092_,
		_w27098_
	);
	LUT2 #(
		.INIT('h8)
	) name23052 (
		_w27097_,
		_w27098_,
		_w27099_
	);
	LUT2 #(
		.INIT('h4)
	) name23053 (
		_w27093_,
		_w27096_,
		_w27100_
	);
	LUT2 #(
		.INIT('h4)
	) name23054 (
		_w27095_,
		_w27100_,
		_w27101_
	);
	LUT2 #(
		.INIT('h8)
	) name23055 (
		_w27099_,
		_w27101_,
		_w27102_
	);
	LUT2 #(
		.INIT('h4)
	) name23056 (
		_w27094_,
		_w27102_,
		_w27103_
	);
	LUT2 #(
		.INIT('h1)
	) name23057 (
		\T_TMODE[1]_pad ,
		_w27103_,
		_w27104_
	);
	LUT2 #(
		.INIT('h1)
	) name23058 (
		_w27086_,
		_w27104_,
		_w27105_
	);
	LUT2 #(
		.INIT('h2)
	) name23059 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27105_,
		_w27106_
	);
	LUT2 #(
		.INIT('h1)
	) name23060 (
		_w27085_,
		_w27106_,
		_w27107_
	);
	LUT2 #(
		.INIT('h1)
	) name23061 (
		_w26973_,
		_w27107_,
		_w27108_
	);
	LUT2 #(
		.INIT('h8)
	) name23062 (
		\sice_SPC_reg[7]/P0001 ,
		_w26969_,
		_w27109_
	);
	LUT2 #(
		.INIT('h1)
	) name23063 (
		_w27084_,
		_w27109_,
		_w27110_
	);
	LUT2 #(
		.INIT('h4)
	) name23064 (
		_w27108_,
		_w27110_,
		_w27111_
	);
	LUT2 #(
		.INIT('h8)
	) name23065 (
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w26973_,
		_w27112_
	);
	LUT2 #(
		.INIT('h8)
	) name23066 (
		_w11525_,
		_w26970_,
		_w27113_
	);
	LUT2 #(
		.INIT('h8)
	) name23067 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[6]/P0001 ,
		_w27114_
	);
	LUT2 #(
		.INIT('h8)
	) name23068 (
		\CM_rd1[6]_pad ,
		_w26984_,
		_w27115_
	);
	LUT2 #(
		.INIT('h8)
	) name23069 (
		\CM_rd6[6]_pad ,
		_w26989_,
		_w27116_
	);
	LUT2 #(
		.INIT('h8)
	) name23070 (
		\CM_rd0[6]_pad ,
		_w26994_,
		_w27117_
	);
	LUT2 #(
		.INIT('h8)
	) name23071 (
		\CM_rd7[6]_pad ,
		_w26997_,
		_w27118_
	);
	LUT2 #(
		.INIT('h8)
	) name23072 (
		\CM_rd2[6]_pad ,
		_w27000_,
		_w27119_
	);
	LUT2 #(
		.INIT('h8)
	) name23073 (
		\CM_rd5[6]_pad ,
		_w27004_,
		_w27120_
	);
	LUT2 #(
		.INIT('h8)
	) name23074 (
		\CM_rd4[6]_pad ,
		_w27008_,
		_w27121_
	);
	LUT2 #(
		.INIT('h8)
	) name23075 (
		\CM_rdm[6]_pad ,
		_w27018_,
		_w27122_
	);
	LUT2 #(
		.INIT('h8)
	) name23076 (
		\CM_rd3[6]_pad ,
		_w27011_,
		_w27123_
	);
	LUT2 #(
		.INIT('h1)
	) name23077 (
		_w27115_,
		_w27116_,
		_w27124_
	);
	LUT2 #(
		.INIT('h1)
	) name23078 (
		_w27117_,
		_w27118_,
		_w27125_
	);
	LUT2 #(
		.INIT('h1)
	) name23079 (
		_w27119_,
		_w27120_,
		_w27126_
	);
	LUT2 #(
		.INIT('h8)
	) name23080 (
		_w27125_,
		_w27126_,
		_w27127_
	);
	LUT2 #(
		.INIT('h4)
	) name23081 (
		_w27121_,
		_w27124_,
		_w27128_
	);
	LUT2 #(
		.INIT('h4)
	) name23082 (
		_w27123_,
		_w27128_,
		_w27129_
	);
	LUT2 #(
		.INIT('h8)
	) name23083 (
		_w27127_,
		_w27129_,
		_w27130_
	);
	LUT2 #(
		.INIT('h4)
	) name23084 (
		_w27122_,
		_w27130_,
		_w27131_
	);
	LUT2 #(
		.INIT('h1)
	) name23085 (
		\T_TMODE[1]_pad ,
		_w27131_,
		_w27132_
	);
	LUT2 #(
		.INIT('h1)
	) name23086 (
		_w27114_,
		_w27132_,
		_w27133_
	);
	LUT2 #(
		.INIT('h2)
	) name23087 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27133_,
		_w27134_
	);
	LUT2 #(
		.INIT('h1)
	) name23088 (
		_w27113_,
		_w27134_,
		_w27135_
	);
	LUT2 #(
		.INIT('h1)
	) name23089 (
		_w26973_,
		_w27135_,
		_w27136_
	);
	LUT2 #(
		.INIT('h8)
	) name23090 (
		\sice_SPC_reg[6]/P0001 ,
		_w26969_,
		_w27137_
	);
	LUT2 #(
		.INIT('h1)
	) name23091 (
		_w27112_,
		_w27137_,
		_w27138_
	);
	LUT2 #(
		.INIT('h4)
	) name23092 (
		_w27136_,
		_w27138_,
		_w27139_
	);
	LUT2 #(
		.INIT('h8)
	) name23093 (
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w26973_,
		_w27140_
	);
	LUT2 #(
		.INIT('h8)
	) name23094 (
		_w10911_,
		_w26970_,
		_w27141_
	);
	LUT2 #(
		.INIT('h8)
	) name23095 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[5]/P0001 ,
		_w27142_
	);
	LUT2 #(
		.INIT('h8)
	) name23096 (
		\CM_rd1[5]_pad ,
		_w26984_,
		_w27143_
	);
	LUT2 #(
		.INIT('h8)
	) name23097 (
		\CM_rd6[5]_pad ,
		_w26989_,
		_w27144_
	);
	LUT2 #(
		.INIT('h8)
	) name23098 (
		\CM_rd0[5]_pad ,
		_w26994_,
		_w27145_
	);
	LUT2 #(
		.INIT('h8)
	) name23099 (
		\CM_rd7[5]_pad ,
		_w26997_,
		_w27146_
	);
	LUT2 #(
		.INIT('h8)
	) name23100 (
		\CM_rd2[5]_pad ,
		_w27000_,
		_w27147_
	);
	LUT2 #(
		.INIT('h8)
	) name23101 (
		\CM_rd5[5]_pad ,
		_w27004_,
		_w27148_
	);
	LUT2 #(
		.INIT('h8)
	) name23102 (
		\CM_rd4[5]_pad ,
		_w27008_,
		_w27149_
	);
	LUT2 #(
		.INIT('h8)
	) name23103 (
		\CM_rdm[5]_pad ,
		_w27018_,
		_w27150_
	);
	LUT2 #(
		.INIT('h8)
	) name23104 (
		\CM_rd3[5]_pad ,
		_w27011_,
		_w27151_
	);
	LUT2 #(
		.INIT('h1)
	) name23105 (
		_w27143_,
		_w27144_,
		_w27152_
	);
	LUT2 #(
		.INIT('h1)
	) name23106 (
		_w27145_,
		_w27146_,
		_w27153_
	);
	LUT2 #(
		.INIT('h1)
	) name23107 (
		_w27147_,
		_w27148_,
		_w27154_
	);
	LUT2 #(
		.INIT('h8)
	) name23108 (
		_w27153_,
		_w27154_,
		_w27155_
	);
	LUT2 #(
		.INIT('h4)
	) name23109 (
		_w27149_,
		_w27152_,
		_w27156_
	);
	LUT2 #(
		.INIT('h4)
	) name23110 (
		_w27151_,
		_w27156_,
		_w27157_
	);
	LUT2 #(
		.INIT('h8)
	) name23111 (
		_w27155_,
		_w27157_,
		_w27158_
	);
	LUT2 #(
		.INIT('h4)
	) name23112 (
		_w27150_,
		_w27158_,
		_w27159_
	);
	LUT2 #(
		.INIT('h1)
	) name23113 (
		\T_TMODE[1]_pad ,
		_w27159_,
		_w27160_
	);
	LUT2 #(
		.INIT('h1)
	) name23114 (
		_w27142_,
		_w27160_,
		_w27161_
	);
	LUT2 #(
		.INIT('h2)
	) name23115 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27161_,
		_w27162_
	);
	LUT2 #(
		.INIT('h1)
	) name23116 (
		_w27141_,
		_w27162_,
		_w27163_
	);
	LUT2 #(
		.INIT('h1)
	) name23117 (
		_w26973_,
		_w27163_,
		_w27164_
	);
	LUT2 #(
		.INIT('h8)
	) name23118 (
		\sice_SPC_reg[5]/P0001 ,
		_w26969_,
		_w27165_
	);
	LUT2 #(
		.INIT('h1)
	) name23119 (
		_w27140_,
		_w27165_,
		_w27166_
	);
	LUT2 #(
		.INIT('h4)
	) name23120 (
		_w27164_,
		_w27166_,
		_w27167_
	);
	LUT2 #(
		.INIT('h8)
	) name23121 (
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w26973_,
		_w27168_
	);
	LUT2 #(
		.INIT('h8)
	) name23122 (
		_w10069_,
		_w26970_,
		_w27169_
	);
	LUT2 #(
		.INIT('h8)
	) name23123 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[4]/P0001 ,
		_w27170_
	);
	LUT2 #(
		.INIT('h8)
	) name23124 (
		\CM_rd1[4]_pad ,
		_w26984_,
		_w27171_
	);
	LUT2 #(
		.INIT('h8)
	) name23125 (
		\CM_rd6[4]_pad ,
		_w26989_,
		_w27172_
	);
	LUT2 #(
		.INIT('h8)
	) name23126 (
		\CM_rd0[4]_pad ,
		_w26994_,
		_w27173_
	);
	LUT2 #(
		.INIT('h8)
	) name23127 (
		\CM_rd7[4]_pad ,
		_w26997_,
		_w27174_
	);
	LUT2 #(
		.INIT('h8)
	) name23128 (
		\CM_rd2[4]_pad ,
		_w27000_,
		_w27175_
	);
	LUT2 #(
		.INIT('h8)
	) name23129 (
		\CM_rd5[4]_pad ,
		_w27004_,
		_w27176_
	);
	LUT2 #(
		.INIT('h8)
	) name23130 (
		\CM_rd4[4]_pad ,
		_w27008_,
		_w27177_
	);
	LUT2 #(
		.INIT('h8)
	) name23131 (
		\CM_rdm[4]_pad ,
		_w27018_,
		_w27178_
	);
	LUT2 #(
		.INIT('h8)
	) name23132 (
		\CM_rd3[4]_pad ,
		_w27011_,
		_w27179_
	);
	LUT2 #(
		.INIT('h1)
	) name23133 (
		_w27171_,
		_w27172_,
		_w27180_
	);
	LUT2 #(
		.INIT('h1)
	) name23134 (
		_w27173_,
		_w27174_,
		_w27181_
	);
	LUT2 #(
		.INIT('h1)
	) name23135 (
		_w27175_,
		_w27176_,
		_w27182_
	);
	LUT2 #(
		.INIT('h8)
	) name23136 (
		_w27181_,
		_w27182_,
		_w27183_
	);
	LUT2 #(
		.INIT('h4)
	) name23137 (
		_w27177_,
		_w27180_,
		_w27184_
	);
	LUT2 #(
		.INIT('h4)
	) name23138 (
		_w27179_,
		_w27184_,
		_w27185_
	);
	LUT2 #(
		.INIT('h8)
	) name23139 (
		_w27183_,
		_w27185_,
		_w27186_
	);
	LUT2 #(
		.INIT('h4)
	) name23140 (
		_w27178_,
		_w27186_,
		_w27187_
	);
	LUT2 #(
		.INIT('h1)
	) name23141 (
		\T_TMODE[1]_pad ,
		_w27187_,
		_w27188_
	);
	LUT2 #(
		.INIT('h1)
	) name23142 (
		_w27170_,
		_w27188_,
		_w27189_
	);
	LUT2 #(
		.INIT('h2)
	) name23143 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27189_,
		_w27190_
	);
	LUT2 #(
		.INIT('h1)
	) name23144 (
		_w27169_,
		_w27190_,
		_w27191_
	);
	LUT2 #(
		.INIT('h1)
	) name23145 (
		_w26973_,
		_w27191_,
		_w27192_
	);
	LUT2 #(
		.INIT('h8)
	) name23146 (
		\sice_SPC_reg[4]/P0001 ,
		_w26969_,
		_w27193_
	);
	LUT2 #(
		.INIT('h1)
	) name23147 (
		_w27168_,
		_w27193_,
		_w27194_
	);
	LUT2 #(
		.INIT('h4)
	) name23148 (
		_w27192_,
		_w27194_,
		_w27195_
	);
	LUT2 #(
		.INIT('h8)
	) name23149 (
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w26973_,
		_w27196_
	);
	LUT2 #(
		.INIT('h8)
	) name23150 (
		_w8113_,
		_w26970_,
		_w27197_
	);
	LUT2 #(
		.INIT('h8)
	) name23151 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[3]/P0001 ,
		_w27198_
	);
	LUT2 #(
		.INIT('h8)
	) name23152 (
		\CM_rd1[3]_pad ,
		_w26984_,
		_w27199_
	);
	LUT2 #(
		.INIT('h8)
	) name23153 (
		\CM_rd6[3]_pad ,
		_w26989_,
		_w27200_
	);
	LUT2 #(
		.INIT('h8)
	) name23154 (
		\CM_rd0[3]_pad ,
		_w26994_,
		_w27201_
	);
	LUT2 #(
		.INIT('h8)
	) name23155 (
		\CM_rd7[3]_pad ,
		_w26997_,
		_w27202_
	);
	LUT2 #(
		.INIT('h8)
	) name23156 (
		\CM_rd2[3]_pad ,
		_w27000_,
		_w27203_
	);
	LUT2 #(
		.INIT('h8)
	) name23157 (
		\CM_rd5[3]_pad ,
		_w27004_,
		_w27204_
	);
	LUT2 #(
		.INIT('h8)
	) name23158 (
		\CM_rd4[3]_pad ,
		_w27008_,
		_w27205_
	);
	LUT2 #(
		.INIT('h8)
	) name23159 (
		\CM_rdm[3]_pad ,
		_w27018_,
		_w27206_
	);
	LUT2 #(
		.INIT('h8)
	) name23160 (
		\CM_rd3[3]_pad ,
		_w27011_,
		_w27207_
	);
	LUT2 #(
		.INIT('h1)
	) name23161 (
		_w27199_,
		_w27200_,
		_w27208_
	);
	LUT2 #(
		.INIT('h1)
	) name23162 (
		_w27201_,
		_w27202_,
		_w27209_
	);
	LUT2 #(
		.INIT('h1)
	) name23163 (
		_w27203_,
		_w27204_,
		_w27210_
	);
	LUT2 #(
		.INIT('h8)
	) name23164 (
		_w27209_,
		_w27210_,
		_w27211_
	);
	LUT2 #(
		.INIT('h4)
	) name23165 (
		_w27205_,
		_w27208_,
		_w27212_
	);
	LUT2 #(
		.INIT('h4)
	) name23166 (
		_w27207_,
		_w27212_,
		_w27213_
	);
	LUT2 #(
		.INIT('h8)
	) name23167 (
		_w27211_,
		_w27213_,
		_w27214_
	);
	LUT2 #(
		.INIT('h4)
	) name23168 (
		_w27206_,
		_w27214_,
		_w27215_
	);
	LUT2 #(
		.INIT('h1)
	) name23169 (
		\T_TMODE[1]_pad ,
		_w27215_,
		_w27216_
	);
	LUT2 #(
		.INIT('h1)
	) name23170 (
		_w27198_,
		_w27216_,
		_w27217_
	);
	LUT2 #(
		.INIT('h2)
	) name23171 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27217_,
		_w27218_
	);
	LUT2 #(
		.INIT('h1)
	) name23172 (
		_w27197_,
		_w27218_,
		_w27219_
	);
	LUT2 #(
		.INIT('h1)
	) name23173 (
		_w26973_,
		_w27219_,
		_w27220_
	);
	LUT2 #(
		.INIT('h8)
	) name23174 (
		\sice_SPC_reg[3]/P0001 ,
		_w26969_,
		_w27221_
	);
	LUT2 #(
		.INIT('h1)
	) name23175 (
		_w27196_,
		_w27221_,
		_w27222_
	);
	LUT2 #(
		.INIT('h4)
	) name23176 (
		_w27220_,
		_w27222_,
		_w27223_
	);
	LUT2 #(
		.INIT('h8)
	) name23177 (
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w26973_,
		_w27224_
	);
	LUT2 #(
		.INIT('h8)
	) name23178 (
		_w8715_,
		_w26970_,
		_w27225_
	);
	LUT2 #(
		.INIT('h8)
	) name23179 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[2]/P0001 ,
		_w27226_
	);
	LUT2 #(
		.INIT('h8)
	) name23180 (
		\CM_rd1[2]_pad ,
		_w26984_,
		_w27227_
	);
	LUT2 #(
		.INIT('h8)
	) name23181 (
		\CM_rd6[2]_pad ,
		_w26989_,
		_w27228_
	);
	LUT2 #(
		.INIT('h8)
	) name23182 (
		\CM_rd0[2]_pad ,
		_w26994_,
		_w27229_
	);
	LUT2 #(
		.INIT('h8)
	) name23183 (
		\CM_rd7[2]_pad ,
		_w26997_,
		_w27230_
	);
	LUT2 #(
		.INIT('h8)
	) name23184 (
		\CM_rd2[2]_pad ,
		_w27000_,
		_w27231_
	);
	LUT2 #(
		.INIT('h8)
	) name23185 (
		\CM_rd5[2]_pad ,
		_w27004_,
		_w27232_
	);
	LUT2 #(
		.INIT('h8)
	) name23186 (
		\CM_rd4[2]_pad ,
		_w27008_,
		_w27233_
	);
	LUT2 #(
		.INIT('h8)
	) name23187 (
		\CM_rdm[2]_pad ,
		_w27018_,
		_w27234_
	);
	LUT2 #(
		.INIT('h8)
	) name23188 (
		\CM_rd3[2]_pad ,
		_w27011_,
		_w27235_
	);
	LUT2 #(
		.INIT('h1)
	) name23189 (
		_w27227_,
		_w27228_,
		_w27236_
	);
	LUT2 #(
		.INIT('h1)
	) name23190 (
		_w27229_,
		_w27230_,
		_w27237_
	);
	LUT2 #(
		.INIT('h1)
	) name23191 (
		_w27231_,
		_w27232_,
		_w27238_
	);
	LUT2 #(
		.INIT('h8)
	) name23192 (
		_w27237_,
		_w27238_,
		_w27239_
	);
	LUT2 #(
		.INIT('h4)
	) name23193 (
		_w27233_,
		_w27236_,
		_w27240_
	);
	LUT2 #(
		.INIT('h4)
	) name23194 (
		_w27235_,
		_w27240_,
		_w27241_
	);
	LUT2 #(
		.INIT('h8)
	) name23195 (
		_w27239_,
		_w27241_,
		_w27242_
	);
	LUT2 #(
		.INIT('h4)
	) name23196 (
		_w27234_,
		_w27242_,
		_w27243_
	);
	LUT2 #(
		.INIT('h1)
	) name23197 (
		\T_TMODE[1]_pad ,
		_w27243_,
		_w27244_
	);
	LUT2 #(
		.INIT('h1)
	) name23198 (
		_w27226_,
		_w27244_,
		_w27245_
	);
	LUT2 #(
		.INIT('h2)
	) name23199 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27245_,
		_w27246_
	);
	LUT2 #(
		.INIT('h1)
	) name23200 (
		_w27225_,
		_w27246_,
		_w27247_
	);
	LUT2 #(
		.INIT('h1)
	) name23201 (
		_w26973_,
		_w27247_,
		_w27248_
	);
	LUT2 #(
		.INIT('h8)
	) name23202 (
		\sice_SPC_reg[2]/P0001 ,
		_w26969_,
		_w27249_
	);
	LUT2 #(
		.INIT('h1)
	) name23203 (
		_w27224_,
		_w27249_,
		_w27250_
	);
	LUT2 #(
		.INIT('h4)
	) name23204 (
		_w27248_,
		_w27250_,
		_w27251_
	);
	LUT2 #(
		.INIT('h8)
	) name23205 (
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w26973_,
		_w27252_
	);
	LUT2 #(
		.INIT('h8)
	) name23206 (
		_w9435_,
		_w26970_,
		_w27253_
	);
	LUT2 #(
		.INIT('h8)
	) name23207 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[1]/P0001 ,
		_w27254_
	);
	LUT2 #(
		.INIT('h8)
	) name23208 (
		\CM_rd1[1]_pad ,
		_w26984_,
		_w27255_
	);
	LUT2 #(
		.INIT('h8)
	) name23209 (
		\CM_rd6[1]_pad ,
		_w26989_,
		_w27256_
	);
	LUT2 #(
		.INIT('h8)
	) name23210 (
		\CM_rd0[1]_pad ,
		_w26994_,
		_w27257_
	);
	LUT2 #(
		.INIT('h8)
	) name23211 (
		\CM_rd7[1]_pad ,
		_w26997_,
		_w27258_
	);
	LUT2 #(
		.INIT('h8)
	) name23212 (
		\CM_rd2[1]_pad ,
		_w27000_,
		_w27259_
	);
	LUT2 #(
		.INIT('h8)
	) name23213 (
		\CM_rd5[1]_pad ,
		_w27004_,
		_w27260_
	);
	LUT2 #(
		.INIT('h8)
	) name23214 (
		\CM_rd4[1]_pad ,
		_w27008_,
		_w27261_
	);
	LUT2 #(
		.INIT('h8)
	) name23215 (
		\CM_rdm[1]_pad ,
		_w27018_,
		_w27262_
	);
	LUT2 #(
		.INIT('h8)
	) name23216 (
		\CM_rd3[1]_pad ,
		_w27011_,
		_w27263_
	);
	LUT2 #(
		.INIT('h1)
	) name23217 (
		_w27255_,
		_w27256_,
		_w27264_
	);
	LUT2 #(
		.INIT('h1)
	) name23218 (
		_w27257_,
		_w27258_,
		_w27265_
	);
	LUT2 #(
		.INIT('h1)
	) name23219 (
		_w27259_,
		_w27260_,
		_w27266_
	);
	LUT2 #(
		.INIT('h8)
	) name23220 (
		_w27265_,
		_w27266_,
		_w27267_
	);
	LUT2 #(
		.INIT('h4)
	) name23221 (
		_w27261_,
		_w27264_,
		_w27268_
	);
	LUT2 #(
		.INIT('h4)
	) name23222 (
		_w27263_,
		_w27268_,
		_w27269_
	);
	LUT2 #(
		.INIT('h8)
	) name23223 (
		_w27267_,
		_w27269_,
		_w27270_
	);
	LUT2 #(
		.INIT('h4)
	) name23224 (
		_w27262_,
		_w27270_,
		_w27271_
	);
	LUT2 #(
		.INIT('h1)
	) name23225 (
		\T_TMODE[1]_pad ,
		_w27271_,
		_w27272_
	);
	LUT2 #(
		.INIT('h1)
	) name23226 (
		_w27254_,
		_w27272_,
		_w27273_
	);
	LUT2 #(
		.INIT('h2)
	) name23227 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27273_,
		_w27274_
	);
	LUT2 #(
		.INIT('h1)
	) name23228 (
		_w27253_,
		_w27274_,
		_w27275_
	);
	LUT2 #(
		.INIT('h1)
	) name23229 (
		_w26973_,
		_w27275_,
		_w27276_
	);
	LUT2 #(
		.INIT('h8)
	) name23230 (
		\sice_SPC_reg[1]/P0001 ,
		_w26969_,
		_w27277_
	);
	LUT2 #(
		.INIT('h1)
	) name23231 (
		_w27252_,
		_w27277_,
		_w27278_
	);
	LUT2 #(
		.INIT('h4)
	) name23232 (
		_w27276_,
		_w27278_,
		_w27279_
	);
	LUT2 #(
		.INIT('h8)
	) name23233 (
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w26973_,
		_w27280_
	);
	LUT2 #(
		.INIT('h8)
	) name23234 (
		_w7607_,
		_w26970_,
		_w27281_
	);
	LUT2 #(
		.INIT('h8)
	) name23235 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[0]/P0001 ,
		_w27282_
	);
	LUT2 #(
		.INIT('h8)
	) name23236 (
		\CM_rd1[0]_pad ,
		_w26984_,
		_w27283_
	);
	LUT2 #(
		.INIT('h8)
	) name23237 (
		\CM_rd6[0]_pad ,
		_w26989_,
		_w27284_
	);
	LUT2 #(
		.INIT('h8)
	) name23238 (
		\CM_rd0[0]_pad ,
		_w26994_,
		_w27285_
	);
	LUT2 #(
		.INIT('h8)
	) name23239 (
		\CM_rd7[0]_pad ,
		_w26997_,
		_w27286_
	);
	LUT2 #(
		.INIT('h8)
	) name23240 (
		\CM_rd2[0]_pad ,
		_w27000_,
		_w27287_
	);
	LUT2 #(
		.INIT('h8)
	) name23241 (
		\CM_rd5[0]_pad ,
		_w27004_,
		_w27288_
	);
	LUT2 #(
		.INIT('h8)
	) name23242 (
		\CM_rd4[0]_pad ,
		_w27008_,
		_w27289_
	);
	LUT2 #(
		.INIT('h8)
	) name23243 (
		\CM_rdm[0]_pad ,
		_w27018_,
		_w27290_
	);
	LUT2 #(
		.INIT('h8)
	) name23244 (
		\CM_rd3[0]_pad ,
		_w27011_,
		_w27291_
	);
	LUT2 #(
		.INIT('h1)
	) name23245 (
		_w27283_,
		_w27284_,
		_w27292_
	);
	LUT2 #(
		.INIT('h1)
	) name23246 (
		_w27285_,
		_w27286_,
		_w27293_
	);
	LUT2 #(
		.INIT('h1)
	) name23247 (
		_w27287_,
		_w27288_,
		_w27294_
	);
	LUT2 #(
		.INIT('h8)
	) name23248 (
		_w27293_,
		_w27294_,
		_w27295_
	);
	LUT2 #(
		.INIT('h4)
	) name23249 (
		_w27289_,
		_w27292_,
		_w27296_
	);
	LUT2 #(
		.INIT('h4)
	) name23250 (
		_w27291_,
		_w27296_,
		_w27297_
	);
	LUT2 #(
		.INIT('h8)
	) name23251 (
		_w27295_,
		_w27297_,
		_w27298_
	);
	LUT2 #(
		.INIT('h4)
	) name23252 (
		_w27290_,
		_w27298_,
		_w27299_
	);
	LUT2 #(
		.INIT('h1)
	) name23253 (
		\T_TMODE[1]_pad ,
		_w27299_,
		_w27300_
	);
	LUT2 #(
		.INIT('h1)
	) name23254 (
		_w27282_,
		_w27300_,
		_w27301_
	);
	LUT2 #(
		.INIT('h2)
	) name23255 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27301_,
		_w27302_
	);
	LUT2 #(
		.INIT('h1)
	) name23256 (
		_w27281_,
		_w27302_,
		_w27303_
	);
	LUT2 #(
		.INIT('h1)
	) name23257 (
		_w26973_,
		_w27303_,
		_w27304_
	);
	LUT2 #(
		.INIT('h8)
	) name23258 (
		\sice_SPC_reg[0]/P0001 ,
		_w26969_,
		_w27305_
	);
	LUT2 #(
		.INIT('h1)
	) name23259 (
		_w27280_,
		_w27305_,
		_w27306_
	);
	LUT2 #(
		.INIT('h4)
	) name23260 (
		_w27304_,
		_w27306_,
		_w27307_
	);
	LUT2 #(
		.INIT('h8)
	) name23261 (
		_w14752_,
		_w27053_,
		_w27308_
	);
	LUT2 #(
		.INIT('h8)
	) name23262 (
		_w18974_,
		_w19776_,
		_w27309_
	);
	LUT2 #(
		.INIT('h2)
	) name23263 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[1]/P0001 ,
		_w17809_,
		_w27310_
	);
	LUT2 #(
		.INIT('h2)
	) name23264 (
		_w19780_,
		_w27310_,
		_w27311_
	);
	LUT2 #(
		.INIT('h4)
	) name23265 (
		_w27309_,
		_w27311_,
		_w27312_
	);
	LUT2 #(
		.INIT('h1)
	) name23266 (
		_w27308_,
		_w27312_,
		_w27313_
	);
	LUT2 #(
		.INIT('h8)
	) name23267 (
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w26973_,
		_w27314_
	);
	LUT2 #(
		.INIT('h8)
	) name23268 (
		_w7340_,
		_w26970_,
		_w27315_
	);
	LUT2 #(
		.INIT('h8)
	) name23269 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[13]/P0001 ,
		_w27316_
	);
	LUT2 #(
		.INIT('h8)
	) name23270 (
		\CM_rd1[13]_pad ,
		_w26984_,
		_w27317_
	);
	LUT2 #(
		.INIT('h8)
	) name23271 (
		\CM_rd6[13]_pad ,
		_w26989_,
		_w27318_
	);
	LUT2 #(
		.INIT('h8)
	) name23272 (
		\CM_rd0[13]_pad ,
		_w26994_,
		_w27319_
	);
	LUT2 #(
		.INIT('h8)
	) name23273 (
		\CM_rd7[13]_pad ,
		_w26997_,
		_w27320_
	);
	LUT2 #(
		.INIT('h8)
	) name23274 (
		\CM_rd2[13]_pad ,
		_w27000_,
		_w27321_
	);
	LUT2 #(
		.INIT('h8)
	) name23275 (
		\CM_rd5[13]_pad ,
		_w27004_,
		_w27322_
	);
	LUT2 #(
		.INIT('h8)
	) name23276 (
		\CM_rd4[13]_pad ,
		_w27008_,
		_w27323_
	);
	LUT2 #(
		.INIT('h8)
	) name23277 (
		\CM_rdm[13]_pad ,
		_w27018_,
		_w27324_
	);
	LUT2 #(
		.INIT('h8)
	) name23278 (
		\CM_rd3[13]_pad ,
		_w27011_,
		_w27325_
	);
	LUT2 #(
		.INIT('h1)
	) name23279 (
		_w27317_,
		_w27318_,
		_w27326_
	);
	LUT2 #(
		.INIT('h1)
	) name23280 (
		_w27319_,
		_w27320_,
		_w27327_
	);
	LUT2 #(
		.INIT('h1)
	) name23281 (
		_w27321_,
		_w27322_,
		_w27328_
	);
	LUT2 #(
		.INIT('h8)
	) name23282 (
		_w27327_,
		_w27328_,
		_w27329_
	);
	LUT2 #(
		.INIT('h4)
	) name23283 (
		_w27323_,
		_w27326_,
		_w27330_
	);
	LUT2 #(
		.INIT('h4)
	) name23284 (
		_w27325_,
		_w27330_,
		_w27331_
	);
	LUT2 #(
		.INIT('h8)
	) name23285 (
		_w27329_,
		_w27331_,
		_w27332_
	);
	LUT2 #(
		.INIT('h4)
	) name23286 (
		_w27324_,
		_w27332_,
		_w27333_
	);
	LUT2 #(
		.INIT('h1)
	) name23287 (
		\T_TMODE[1]_pad ,
		_w27333_,
		_w27334_
	);
	LUT2 #(
		.INIT('h1)
	) name23288 (
		_w27316_,
		_w27334_,
		_w27335_
	);
	LUT2 #(
		.INIT('h2)
	) name23289 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27335_,
		_w27336_
	);
	LUT2 #(
		.INIT('h1)
	) name23290 (
		_w27315_,
		_w27336_,
		_w27337_
	);
	LUT2 #(
		.INIT('h1)
	) name23291 (
		_w26973_,
		_w27337_,
		_w27338_
	);
	LUT2 #(
		.INIT('h8)
	) name23292 (
		\sice_SPC_reg[13]/P0001 ,
		_w26969_,
		_w27339_
	);
	LUT2 #(
		.INIT('h1)
	) name23293 (
		_w27314_,
		_w27339_,
		_w27340_
	);
	LUT2 #(
		.INIT('h4)
	) name23294 (
		_w27338_,
		_w27340_,
		_w27341_
	);
	LUT2 #(
		.INIT('h8)
	) name23295 (
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w26973_,
		_w27342_
	);
	LUT2 #(
		.INIT('h8)
	) name23296 (
		_w9178_,
		_w26970_,
		_w27343_
	);
	LUT2 #(
		.INIT('h8)
	) name23297 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[12]/P0001 ,
		_w27344_
	);
	LUT2 #(
		.INIT('h8)
	) name23298 (
		\CM_rd1[12]_pad ,
		_w26984_,
		_w27345_
	);
	LUT2 #(
		.INIT('h8)
	) name23299 (
		\CM_rd6[12]_pad ,
		_w26989_,
		_w27346_
	);
	LUT2 #(
		.INIT('h8)
	) name23300 (
		\CM_rd0[12]_pad ,
		_w26994_,
		_w27347_
	);
	LUT2 #(
		.INIT('h8)
	) name23301 (
		\CM_rd7[12]_pad ,
		_w26997_,
		_w27348_
	);
	LUT2 #(
		.INIT('h8)
	) name23302 (
		\CM_rd2[12]_pad ,
		_w27000_,
		_w27349_
	);
	LUT2 #(
		.INIT('h8)
	) name23303 (
		\CM_rd5[12]_pad ,
		_w27004_,
		_w27350_
	);
	LUT2 #(
		.INIT('h8)
	) name23304 (
		\CM_rd4[12]_pad ,
		_w27008_,
		_w27351_
	);
	LUT2 #(
		.INIT('h8)
	) name23305 (
		\CM_rdm[12]_pad ,
		_w27018_,
		_w27352_
	);
	LUT2 #(
		.INIT('h8)
	) name23306 (
		\CM_rd3[12]_pad ,
		_w27011_,
		_w27353_
	);
	LUT2 #(
		.INIT('h1)
	) name23307 (
		_w27345_,
		_w27346_,
		_w27354_
	);
	LUT2 #(
		.INIT('h1)
	) name23308 (
		_w27347_,
		_w27348_,
		_w27355_
	);
	LUT2 #(
		.INIT('h1)
	) name23309 (
		_w27349_,
		_w27350_,
		_w27356_
	);
	LUT2 #(
		.INIT('h8)
	) name23310 (
		_w27355_,
		_w27356_,
		_w27357_
	);
	LUT2 #(
		.INIT('h4)
	) name23311 (
		_w27351_,
		_w27354_,
		_w27358_
	);
	LUT2 #(
		.INIT('h4)
	) name23312 (
		_w27353_,
		_w27358_,
		_w27359_
	);
	LUT2 #(
		.INIT('h8)
	) name23313 (
		_w27357_,
		_w27359_,
		_w27360_
	);
	LUT2 #(
		.INIT('h4)
	) name23314 (
		_w27352_,
		_w27360_,
		_w27361_
	);
	LUT2 #(
		.INIT('h1)
	) name23315 (
		\T_TMODE[1]_pad ,
		_w27361_,
		_w27362_
	);
	LUT2 #(
		.INIT('h1)
	) name23316 (
		_w27344_,
		_w27362_,
		_w27363_
	);
	LUT2 #(
		.INIT('h2)
	) name23317 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27363_,
		_w27364_
	);
	LUT2 #(
		.INIT('h1)
	) name23318 (
		_w27343_,
		_w27364_,
		_w27365_
	);
	LUT2 #(
		.INIT('h1)
	) name23319 (
		_w26973_,
		_w27365_,
		_w27366_
	);
	LUT2 #(
		.INIT('h8)
	) name23320 (
		\sice_SPC_reg[12]/P0001 ,
		_w26969_,
		_w27367_
	);
	LUT2 #(
		.INIT('h1)
	) name23321 (
		_w27342_,
		_w27367_,
		_w27368_
	);
	LUT2 #(
		.INIT('h4)
	) name23322 (
		_w27366_,
		_w27368_,
		_w27369_
	);
	LUT2 #(
		.INIT('h8)
	) name23323 (
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w26973_,
		_w27370_
	);
	LUT2 #(
		.INIT('h8)
	) name23324 (
		_w10638_,
		_w26970_,
		_w27371_
	);
	LUT2 #(
		.INIT('h8)
	) name23325 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[8]/P0001 ,
		_w27372_
	);
	LUT2 #(
		.INIT('h8)
	) name23326 (
		\CM_rd1[8]_pad ,
		_w26984_,
		_w27373_
	);
	LUT2 #(
		.INIT('h8)
	) name23327 (
		\CM_rd6[8]_pad ,
		_w26989_,
		_w27374_
	);
	LUT2 #(
		.INIT('h8)
	) name23328 (
		\CM_rd0[8]_pad ,
		_w26994_,
		_w27375_
	);
	LUT2 #(
		.INIT('h8)
	) name23329 (
		\CM_rd7[8]_pad ,
		_w26997_,
		_w27376_
	);
	LUT2 #(
		.INIT('h8)
	) name23330 (
		\CM_rd2[8]_pad ,
		_w27000_,
		_w27377_
	);
	LUT2 #(
		.INIT('h8)
	) name23331 (
		\CM_rd5[8]_pad ,
		_w27004_,
		_w27378_
	);
	LUT2 #(
		.INIT('h8)
	) name23332 (
		\CM_rd4[8]_pad ,
		_w27008_,
		_w27379_
	);
	LUT2 #(
		.INIT('h8)
	) name23333 (
		\CM_rdm[8]_pad ,
		_w27018_,
		_w27380_
	);
	LUT2 #(
		.INIT('h8)
	) name23334 (
		\CM_rd3[8]_pad ,
		_w27011_,
		_w27381_
	);
	LUT2 #(
		.INIT('h1)
	) name23335 (
		_w27373_,
		_w27374_,
		_w27382_
	);
	LUT2 #(
		.INIT('h1)
	) name23336 (
		_w27375_,
		_w27376_,
		_w27383_
	);
	LUT2 #(
		.INIT('h1)
	) name23337 (
		_w27377_,
		_w27378_,
		_w27384_
	);
	LUT2 #(
		.INIT('h8)
	) name23338 (
		_w27383_,
		_w27384_,
		_w27385_
	);
	LUT2 #(
		.INIT('h4)
	) name23339 (
		_w27379_,
		_w27382_,
		_w27386_
	);
	LUT2 #(
		.INIT('h4)
	) name23340 (
		_w27381_,
		_w27386_,
		_w27387_
	);
	LUT2 #(
		.INIT('h8)
	) name23341 (
		_w27385_,
		_w27387_,
		_w27388_
	);
	LUT2 #(
		.INIT('h4)
	) name23342 (
		_w27380_,
		_w27388_,
		_w27389_
	);
	LUT2 #(
		.INIT('h1)
	) name23343 (
		\T_TMODE[1]_pad ,
		_w27389_,
		_w27390_
	);
	LUT2 #(
		.INIT('h1)
	) name23344 (
		_w27372_,
		_w27390_,
		_w27391_
	);
	LUT2 #(
		.INIT('h2)
	) name23345 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27391_,
		_w27392_
	);
	LUT2 #(
		.INIT('h1)
	) name23346 (
		_w27371_,
		_w27392_,
		_w27393_
	);
	LUT2 #(
		.INIT('h1)
	) name23347 (
		_w26973_,
		_w27393_,
		_w27394_
	);
	LUT2 #(
		.INIT('h8)
	) name23348 (
		\sice_SPC_reg[8]/P0001 ,
		_w26969_,
		_w27395_
	);
	LUT2 #(
		.INIT('h1)
	) name23349 (
		_w27370_,
		_w27395_,
		_w27396_
	);
	LUT2 #(
		.INIT('h4)
	) name23350 (
		_w27394_,
		_w27396_,
		_w27397_
	);
	LUT2 #(
		.INIT('h8)
	) name23351 (
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w26973_,
		_w27398_
	);
	LUT2 #(
		.INIT('h8)
	) name23352 (
		_w10289_,
		_w26970_,
		_w27399_
	);
	LUT2 #(
		.INIT('h8)
	) name23353 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[9]/P0001 ,
		_w27400_
	);
	LUT2 #(
		.INIT('h8)
	) name23354 (
		\CM_rd1[9]_pad ,
		_w26984_,
		_w27401_
	);
	LUT2 #(
		.INIT('h8)
	) name23355 (
		\CM_rd6[9]_pad ,
		_w26989_,
		_w27402_
	);
	LUT2 #(
		.INIT('h8)
	) name23356 (
		\CM_rd0[9]_pad ,
		_w26994_,
		_w27403_
	);
	LUT2 #(
		.INIT('h8)
	) name23357 (
		\CM_rd7[9]_pad ,
		_w26997_,
		_w27404_
	);
	LUT2 #(
		.INIT('h8)
	) name23358 (
		\CM_rd2[9]_pad ,
		_w27000_,
		_w27405_
	);
	LUT2 #(
		.INIT('h8)
	) name23359 (
		\CM_rd5[9]_pad ,
		_w27004_,
		_w27406_
	);
	LUT2 #(
		.INIT('h8)
	) name23360 (
		\CM_rd4[9]_pad ,
		_w27008_,
		_w27407_
	);
	LUT2 #(
		.INIT('h8)
	) name23361 (
		\CM_rdm[9]_pad ,
		_w27018_,
		_w27408_
	);
	LUT2 #(
		.INIT('h8)
	) name23362 (
		\CM_rd3[9]_pad ,
		_w27011_,
		_w27409_
	);
	LUT2 #(
		.INIT('h1)
	) name23363 (
		_w27401_,
		_w27402_,
		_w27410_
	);
	LUT2 #(
		.INIT('h1)
	) name23364 (
		_w27403_,
		_w27404_,
		_w27411_
	);
	LUT2 #(
		.INIT('h1)
	) name23365 (
		_w27405_,
		_w27406_,
		_w27412_
	);
	LUT2 #(
		.INIT('h8)
	) name23366 (
		_w27411_,
		_w27412_,
		_w27413_
	);
	LUT2 #(
		.INIT('h4)
	) name23367 (
		_w27407_,
		_w27410_,
		_w27414_
	);
	LUT2 #(
		.INIT('h4)
	) name23368 (
		_w27409_,
		_w27414_,
		_w27415_
	);
	LUT2 #(
		.INIT('h8)
	) name23369 (
		_w27413_,
		_w27415_,
		_w27416_
	);
	LUT2 #(
		.INIT('h4)
	) name23370 (
		_w27408_,
		_w27416_,
		_w27417_
	);
	LUT2 #(
		.INIT('h1)
	) name23371 (
		\T_TMODE[1]_pad ,
		_w27417_,
		_w27418_
	);
	LUT2 #(
		.INIT('h1)
	) name23372 (
		_w27400_,
		_w27418_,
		_w27419_
	);
	LUT2 #(
		.INIT('h2)
	) name23373 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27419_,
		_w27420_
	);
	LUT2 #(
		.INIT('h1)
	) name23374 (
		_w27399_,
		_w27420_,
		_w27421_
	);
	LUT2 #(
		.INIT('h1)
	) name23375 (
		_w26973_,
		_w27421_,
		_w27422_
	);
	LUT2 #(
		.INIT('h8)
	) name23376 (
		\sice_SPC_reg[9]/P0001 ,
		_w26969_,
		_w27423_
	);
	LUT2 #(
		.INIT('h1)
	) name23377 (
		_w27398_,
		_w27423_,
		_w27424_
	);
	LUT2 #(
		.INIT('h4)
	) name23378 (
		_w27422_,
		_w27424_,
		_w27425_
	);
	LUT2 #(
		.INIT('h8)
	) name23379 (
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w26973_,
		_w27426_
	);
	LUT2 #(
		.INIT('h8)
	) name23380 (
		_w8460_,
		_w26970_,
		_w27427_
	);
	LUT2 #(
		.INIT('h8)
	) name23381 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[11]/P0001 ,
		_w27428_
	);
	LUT2 #(
		.INIT('h8)
	) name23382 (
		\CM_rd1[11]_pad ,
		_w26984_,
		_w27429_
	);
	LUT2 #(
		.INIT('h8)
	) name23383 (
		\CM_rd6[11]_pad ,
		_w26989_,
		_w27430_
	);
	LUT2 #(
		.INIT('h8)
	) name23384 (
		\CM_rd0[11]_pad ,
		_w26994_,
		_w27431_
	);
	LUT2 #(
		.INIT('h8)
	) name23385 (
		\CM_rd7[11]_pad ,
		_w26997_,
		_w27432_
	);
	LUT2 #(
		.INIT('h8)
	) name23386 (
		\CM_rd2[11]_pad ,
		_w27000_,
		_w27433_
	);
	LUT2 #(
		.INIT('h8)
	) name23387 (
		\CM_rd5[11]_pad ,
		_w27004_,
		_w27434_
	);
	LUT2 #(
		.INIT('h8)
	) name23388 (
		\CM_rd4[11]_pad ,
		_w27008_,
		_w27435_
	);
	LUT2 #(
		.INIT('h8)
	) name23389 (
		\CM_rdm[11]_pad ,
		_w27018_,
		_w27436_
	);
	LUT2 #(
		.INIT('h8)
	) name23390 (
		\CM_rd3[11]_pad ,
		_w27011_,
		_w27437_
	);
	LUT2 #(
		.INIT('h1)
	) name23391 (
		_w27429_,
		_w27430_,
		_w27438_
	);
	LUT2 #(
		.INIT('h1)
	) name23392 (
		_w27431_,
		_w27432_,
		_w27439_
	);
	LUT2 #(
		.INIT('h1)
	) name23393 (
		_w27433_,
		_w27434_,
		_w27440_
	);
	LUT2 #(
		.INIT('h8)
	) name23394 (
		_w27439_,
		_w27440_,
		_w27441_
	);
	LUT2 #(
		.INIT('h4)
	) name23395 (
		_w27435_,
		_w27438_,
		_w27442_
	);
	LUT2 #(
		.INIT('h4)
	) name23396 (
		_w27437_,
		_w27442_,
		_w27443_
	);
	LUT2 #(
		.INIT('h8)
	) name23397 (
		_w27441_,
		_w27443_,
		_w27444_
	);
	LUT2 #(
		.INIT('h4)
	) name23398 (
		_w27436_,
		_w27444_,
		_w27445_
	);
	LUT2 #(
		.INIT('h1)
	) name23399 (
		\T_TMODE[1]_pad ,
		_w27445_,
		_w27446_
	);
	LUT2 #(
		.INIT('h1)
	) name23400 (
		_w27428_,
		_w27446_,
		_w27447_
	);
	LUT2 #(
		.INIT('h2)
	) name23401 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27447_,
		_w27448_
	);
	LUT2 #(
		.INIT('h1)
	) name23402 (
		_w27427_,
		_w27448_,
		_w27449_
	);
	LUT2 #(
		.INIT('h1)
	) name23403 (
		_w26973_,
		_w27449_,
		_w27450_
	);
	LUT2 #(
		.INIT('h8)
	) name23404 (
		\sice_SPC_reg[11]/P0001 ,
		_w26969_,
		_w27451_
	);
	LUT2 #(
		.INIT('h1)
	) name23405 (
		_w27426_,
		_w27451_,
		_w27452_
	);
	LUT2 #(
		.INIT('h4)
	) name23406 (
		_w27450_,
		_w27452_,
		_w27453_
	);
	LUT2 #(
		.INIT('h8)
	) name23407 (
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w26973_,
		_w27454_
	);
	LUT2 #(
		.INIT('h8)
	) name23408 (
		_w7859_,
		_w26970_,
		_w27455_
	);
	LUT2 #(
		.INIT('h8)
	) name23409 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[10]/P0001 ,
		_w27456_
	);
	LUT2 #(
		.INIT('h8)
	) name23410 (
		\CM_rd1[10]_pad ,
		_w26984_,
		_w27457_
	);
	LUT2 #(
		.INIT('h8)
	) name23411 (
		\CM_rd6[10]_pad ,
		_w26989_,
		_w27458_
	);
	LUT2 #(
		.INIT('h8)
	) name23412 (
		\CM_rd0[10]_pad ,
		_w26994_,
		_w27459_
	);
	LUT2 #(
		.INIT('h8)
	) name23413 (
		\CM_rd7[10]_pad ,
		_w26997_,
		_w27460_
	);
	LUT2 #(
		.INIT('h8)
	) name23414 (
		\CM_rd2[10]_pad ,
		_w27000_,
		_w27461_
	);
	LUT2 #(
		.INIT('h8)
	) name23415 (
		\CM_rd5[10]_pad ,
		_w27004_,
		_w27462_
	);
	LUT2 #(
		.INIT('h8)
	) name23416 (
		\CM_rd4[10]_pad ,
		_w27008_,
		_w27463_
	);
	LUT2 #(
		.INIT('h8)
	) name23417 (
		\CM_rdm[10]_pad ,
		_w27018_,
		_w27464_
	);
	LUT2 #(
		.INIT('h8)
	) name23418 (
		\CM_rd3[10]_pad ,
		_w27011_,
		_w27465_
	);
	LUT2 #(
		.INIT('h1)
	) name23419 (
		_w27457_,
		_w27458_,
		_w27466_
	);
	LUT2 #(
		.INIT('h1)
	) name23420 (
		_w27459_,
		_w27460_,
		_w27467_
	);
	LUT2 #(
		.INIT('h1)
	) name23421 (
		_w27461_,
		_w27462_,
		_w27468_
	);
	LUT2 #(
		.INIT('h8)
	) name23422 (
		_w27467_,
		_w27468_,
		_w27469_
	);
	LUT2 #(
		.INIT('h4)
	) name23423 (
		_w27463_,
		_w27466_,
		_w27470_
	);
	LUT2 #(
		.INIT('h4)
	) name23424 (
		_w27465_,
		_w27470_,
		_w27471_
	);
	LUT2 #(
		.INIT('h8)
	) name23425 (
		_w27469_,
		_w27471_,
		_w27472_
	);
	LUT2 #(
		.INIT('h4)
	) name23426 (
		_w27464_,
		_w27472_,
		_w27473_
	);
	LUT2 #(
		.INIT('h1)
	) name23427 (
		\T_TMODE[1]_pad ,
		_w27473_,
		_w27474_
	);
	LUT2 #(
		.INIT('h1)
	) name23428 (
		_w27456_,
		_w27474_,
		_w27475_
	);
	LUT2 #(
		.INIT('h2)
	) name23429 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w27475_,
		_w27476_
	);
	LUT2 #(
		.INIT('h1)
	) name23430 (
		_w27455_,
		_w27476_,
		_w27477_
	);
	LUT2 #(
		.INIT('h1)
	) name23431 (
		_w26973_,
		_w27477_,
		_w27478_
	);
	LUT2 #(
		.INIT('h8)
	) name23432 (
		\sice_SPC_reg[10]/P0001 ,
		_w26969_,
		_w27479_
	);
	LUT2 #(
		.INIT('h1)
	) name23433 (
		_w27454_,
		_w27479_,
		_w27480_
	);
	LUT2 #(
		.INIT('h4)
	) name23434 (
		_w27478_,
		_w27480_,
		_w27481_
	);
	LUT2 #(
		.INIT('h2)
	) name23435 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w17814_,
		_w27482_
	);
	LUT2 #(
		.INIT('h8)
	) name23436 (
		_w26262_,
		_w26263_,
		_w27483_
	);
	LUT2 #(
		.INIT('h8)
	) name23437 (
		_w26261_,
		_w26269_,
		_w27484_
	);
	LUT2 #(
		.INIT('h4)
	) name23438 (
		_w27483_,
		_w27484_,
		_w27485_
	);
	LUT2 #(
		.INIT('h8)
	) name23439 (
		_w26271_,
		_w26273_,
		_w27486_
	);
	LUT2 #(
		.INIT('h4)
	) name23440 (
		_w27485_,
		_w27486_,
		_w27487_
	);
	LUT2 #(
		.INIT('h2)
	) name23441 (
		_w26275_,
		_w27487_,
		_w27488_
	);
	LUT2 #(
		.INIT('h1)
	) name23442 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w27488_,
		_w27489_
	);
	LUT2 #(
		.INIT('h1)
	) name23443 (
		_w27482_,
		_w27489_,
		_w27490_
	);
	LUT2 #(
		.INIT('h2)
	) name23444 (
		_w23677_,
		_w27490_,
		_w27491_
	);
	LUT2 #(
		.INIT('h1)
	) name23445 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[2]/P0001 ,
		_w23677_,
		_w27492_
	);
	LUT2 #(
		.INIT('h1)
	) name23446 (
		_w27491_,
		_w27492_,
		_w27493_
	);
	LUT2 #(
		.INIT('h2)
	) name23447 (
		_w23598_,
		_w27490_,
		_w27494_
	);
	LUT2 #(
		.INIT('h1)
	) name23448 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[2]/P0001 ,
		_w23598_,
		_w27495_
	);
	LUT2 #(
		.INIT('h1)
	) name23449 (
		_w27494_,
		_w27495_,
		_w27496_
	);
	LUT2 #(
		.INIT('h4)
	) name23450 (
		_w13006_,
		_w13570_,
		_w27497_
	);
	LUT2 #(
		.INIT('h2)
	) name23451 (
		_w13569_,
		_w27028_,
		_w27498_
	);
	LUT2 #(
		.INIT('h4)
	) name23452 (
		_w5882_,
		_w13569_,
		_w27499_
	);
	LUT2 #(
		.INIT('h2)
	) name23453 (
		\idma_IADi_reg[7]/P0001 ,
		_w27499_,
		_w27500_
	);
	LUT2 #(
		.INIT('h1)
	) name23454 (
		_w13570_,
		_w27500_,
		_w27501_
	);
	LUT2 #(
		.INIT('h4)
	) name23455 (
		_w27498_,
		_w27501_,
		_w27502_
	);
	LUT2 #(
		.INIT('h1)
	) name23456 (
		_w11752_,
		_w27497_,
		_w27503_
	);
	LUT2 #(
		.INIT('h4)
	) name23457 (
		_w27502_,
		_w27503_,
		_w27504_
	);
	LUT2 #(
		.INIT('h8)
	) name23458 (
		_w11265_,
		_w11752_,
		_w27505_
	);
	LUT2 #(
		.INIT('h1)
	) name23459 (
		_w27504_,
		_w27505_,
		_w27506_
	);
	LUT2 #(
		.INIT('h4)
	) name23460 (
		_w12972_,
		_w13570_,
		_w27507_
	);
	LUT2 #(
		.INIT('h2)
	) name23461 (
		_w13569_,
		_w27075_,
		_w27508_
	);
	LUT2 #(
		.INIT('h2)
	) name23462 (
		\idma_IADi_reg[6]/P0001 ,
		_w27499_,
		_w27509_
	);
	LUT2 #(
		.INIT('h1)
	) name23463 (
		_w13570_,
		_w27509_,
		_w27510_
	);
	LUT2 #(
		.INIT('h4)
	) name23464 (
		_w27508_,
		_w27510_,
		_w27511_
	);
	LUT2 #(
		.INIT('h1)
	) name23465 (
		_w11752_,
		_w27511_,
		_w27512_
	);
	LUT2 #(
		.INIT('h4)
	) name23466 (
		_w27507_,
		_w27512_,
		_w27513_
	);
	LUT2 #(
		.INIT('h8)
	) name23467 (
		_w11525_,
		_w11752_,
		_w27514_
	);
	LUT2 #(
		.INIT('h1)
	) name23468 (
		_w27513_,
		_w27514_,
		_w27515_
	);
	LUT2 #(
		.INIT('h4)
	) name23469 (
		_w12938_,
		_w13570_,
		_w27516_
	);
	LUT2 #(
		.INIT('h2)
	) name23470 (
		_w13569_,
		_w27333_,
		_w27517_
	);
	LUT2 #(
		.INIT('h2)
	) name23471 (
		\idma_IADi_reg[5]/P0001 ,
		_w27499_,
		_w27518_
	);
	LUT2 #(
		.INIT('h1)
	) name23472 (
		_w13570_,
		_w27518_,
		_w27519_
	);
	LUT2 #(
		.INIT('h4)
	) name23473 (
		_w27517_,
		_w27519_,
		_w27520_
	);
	LUT2 #(
		.INIT('h1)
	) name23474 (
		_w11752_,
		_w27516_,
		_w27521_
	);
	LUT2 #(
		.INIT('h4)
	) name23475 (
		_w27520_,
		_w27521_,
		_w27522_
	);
	LUT2 #(
		.INIT('h8)
	) name23476 (
		_w10911_,
		_w11752_,
		_w27523_
	);
	LUT2 #(
		.INIT('h1)
	) name23477 (
		_w27522_,
		_w27523_,
		_w27524_
	);
	LUT2 #(
		.INIT('h4)
	) name23478 (
		_w12904_,
		_w13570_,
		_w27525_
	);
	LUT2 #(
		.INIT('h2)
	) name23479 (
		_w13569_,
		_w27361_,
		_w27526_
	);
	LUT2 #(
		.INIT('h2)
	) name23480 (
		\idma_IADi_reg[4]/P0001 ,
		_w27499_,
		_w27527_
	);
	LUT2 #(
		.INIT('h1)
	) name23481 (
		_w13570_,
		_w27527_,
		_w27528_
	);
	LUT2 #(
		.INIT('h4)
	) name23482 (
		_w27526_,
		_w27528_,
		_w27529_
	);
	LUT2 #(
		.INIT('h1)
	) name23483 (
		_w11752_,
		_w27525_,
		_w27530_
	);
	LUT2 #(
		.INIT('h4)
	) name23484 (
		_w27529_,
		_w27530_,
		_w27531_
	);
	LUT2 #(
		.INIT('h8)
	) name23485 (
		_w10069_,
		_w11752_,
		_w27532_
	);
	LUT2 #(
		.INIT('h1)
	) name23486 (
		_w27531_,
		_w27532_,
		_w27533_
	);
	LUT2 #(
		.INIT('h4)
	) name23487 (
		_w12870_,
		_w13570_,
		_w27534_
	);
	LUT2 #(
		.INIT('h2)
	) name23488 (
		_w13569_,
		_w27445_,
		_w27535_
	);
	LUT2 #(
		.INIT('h2)
	) name23489 (
		\idma_IADi_reg[3]/P0001 ,
		_w27499_,
		_w27536_
	);
	LUT2 #(
		.INIT('h1)
	) name23490 (
		_w13570_,
		_w27536_,
		_w27537_
	);
	LUT2 #(
		.INIT('h4)
	) name23491 (
		_w27535_,
		_w27537_,
		_w27538_
	);
	LUT2 #(
		.INIT('h1)
	) name23492 (
		_w11752_,
		_w27534_,
		_w27539_
	);
	LUT2 #(
		.INIT('h4)
	) name23493 (
		_w27538_,
		_w27539_,
		_w27540_
	);
	LUT2 #(
		.INIT('h8)
	) name23494 (
		_w8113_,
		_w11752_,
		_w27541_
	);
	LUT2 #(
		.INIT('h1)
	) name23495 (
		_w27540_,
		_w27541_,
		_w27542_
	);
	LUT2 #(
		.INIT('h4)
	) name23496 (
		_w12836_,
		_w13570_,
		_w27543_
	);
	LUT2 #(
		.INIT('h2)
	) name23497 (
		_w13569_,
		_w27473_,
		_w27544_
	);
	LUT2 #(
		.INIT('h2)
	) name23498 (
		\idma_IADi_reg[2]/P0001 ,
		_w27499_,
		_w27545_
	);
	LUT2 #(
		.INIT('h1)
	) name23499 (
		_w13570_,
		_w27545_,
		_w27546_
	);
	LUT2 #(
		.INIT('h4)
	) name23500 (
		_w27544_,
		_w27546_,
		_w27547_
	);
	LUT2 #(
		.INIT('h1)
	) name23501 (
		_w11752_,
		_w27543_,
		_w27548_
	);
	LUT2 #(
		.INIT('h4)
	) name23502 (
		_w27547_,
		_w27548_,
		_w27549_
	);
	LUT2 #(
		.INIT('h8)
	) name23503 (
		_w8715_,
		_w11752_,
		_w27550_
	);
	LUT2 #(
		.INIT('h1)
	) name23504 (
		_w27549_,
		_w27550_,
		_w27551_
	);
	LUT2 #(
		.INIT('h4)
	) name23505 (
		_w12802_,
		_w13570_,
		_w27552_
	);
	LUT2 #(
		.INIT('h2)
	) name23506 (
		_w13569_,
		_w27417_,
		_w27553_
	);
	LUT2 #(
		.INIT('h2)
	) name23507 (
		\idma_IADi_reg[1]/P0001 ,
		_w27499_,
		_w27554_
	);
	LUT2 #(
		.INIT('h1)
	) name23508 (
		_w13570_,
		_w27554_,
		_w27555_
	);
	LUT2 #(
		.INIT('h4)
	) name23509 (
		_w27553_,
		_w27555_,
		_w27556_
	);
	LUT2 #(
		.INIT('h1)
	) name23510 (
		_w11752_,
		_w27552_,
		_w27557_
	);
	LUT2 #(
		.INIT('h4)
	) name23511 (
		_w27556_,
		_w27557_,
		_w27558_
	);
	LUT2 #(
		.INIT('h8)
	) name23512 (
		_w9435_,
		_w11752_,
		_w27559_
	);
	LUT2 #(
		.INIT('h1)
	) name23513 (
		_w27558_,
		_w27559_,
		_w27560_
	);
	LUT2 #(
		.INIT('h8)
	) name23514 (
		\CM_rd1[23]_pad ,
		_w26984_,
		_w27561_
	);
	LUT2 #(
		.INIT('h8)
	) name23515 (
		\CM_rd6[23]_pad ,
		_w26989_,
		_w27562_
	);
	LUT2 #(
		.INIT('h8)
	) name23516 (
		\CM_rd0[23]_pad ,
		_w26994_,
		_w27563_
	);
	LUT2 #(
		.INIT('h8)
	) name23517 (
		\CM_rd7[23]_pad ,
		_w26997_,
		_w27564_
	);
	LUT2 #(
		.INIT('h8)
	) name23518 (
		\CM_rd2[23]_pad ,
		_w27000_,
		_w27565_
	);
	LUT2 #(
		.INIT('h8)
	) name23519 (
		\CM_rd5[23]_pad ,
		_w27004_,
		_w27566_
	);
	LUT2 #(
		.INIT('h8)
	) name23520 (
		\CM_rd4[23]_pad ,
		_w27008_,
		_w27567_
	);
	LUT2 #(
		.INIT('h8)
	) name23521 (
		\CM_rdm[23]_pad ,
		_w27018_,
		_w27568_
	);
	LUT2 #(
		.INIT('h8)
	) name23522 (
		\CM_rd3[23]_pad ,
		_w27011_,
		_w27569_
	);
	LUT2 #(
		.INIT('h1)
	) name23523 (
		_w27561_,
		_w27562_,
		_w27570_
	);
	LUT2 #(
		.INIT('h1)
	) name23524 (
		_w27563_,
		_w27564_,
		_w27571_
	);
	LUT2 #(
		.INIT('h1)
	) name23525 (
		_w27565_,
		_w27566_,
		_w27572_
	);
	LUT2 #(
		.INIT('h8)
	) name23526 (
		_w27571_,
		_w27572_,
		_w27573_
	);
	LUT2 #(
		.INIT('h4)
	) name23527 (
		_w27567_,
		_w27570_,
		_w27574_
	);
	LUT2 #(
		.INIT('h4)
	) name23528 (
		_w27569_,
		_w27574_,
		_w27575_
	);
	LUT2 #(
		.INIT('h8)
	) name23529 (
		_w27573_,
		_w27575_,
		_w27576_
	);
	LUT2 #(
		.INIT('h4)
	) name23530 (
		_w27568_,
		_w27576_,
		_w27577_
	);
	LUT2 #(
		.INIT('h2)
	) name23531 (
		_w27499_,
		_w27577_,
		_w27578_
	);
	LUT2 #(
		.INIT('h2)
	) name23532 (
		\idma_IADi_reg[15]/P0001 ,
		_w27499_,
		_w27579_
	);
	LUT2 #(
		.INIT('h1)
	) name23533 (
		_w27578_,
		_w27579_,
		_w27580_
	);
	LUT2 #(
		.INIT('h1)
	) name23534 (
		_w13570_,
		_w27580_,
		_w27581_
	);
	LUT2 #(
		.INIT('h8)
	) name23535 (
		_w12771_,
		_w13570_,
		_w27582_
	);
	LUT2 #(
		.INIT('h1)
	) name23536 (
		_w27581_,
		_w27582_,
		_w27583_
	);
	LUT2 #(
		.INIT('h1)
	) name23537 (
		_w11752_,
		_w27583_,
		_w27584_
	);
	LUT2 #(
		.INIT('h8)
	) name23538 (
		_w11752_,
		_w12743_,
		_w27585_
	);
	LUT2 #(
		.INIT('h1)
	) name23539 (
		_w27584_,
		_w27585_,
		_w27586_
	);
	LUT2 #(
		.INIT('h8)
	) name23540 (
		\CM_rd1[22]_pad ,
		_w26984_,
		_w27587_
	);
	LUT2 #(
		.INIT('h8)
	) name23541 (
		\CM_rd6[22]_pad ,
		_w26989_,
		_w27588_
	);
	LUT2 #(
		.INIT('h8)
	) name23542 (
		\CM_rd0[22]_pad ,
		_w26994_,
		_w27589_
	);
	LUT2 #(
		.INIT('h8)
	) name23543 (
		\CM_rd7[22]_pad ,
		_w26997_,
		_w27590_
	);
	LUT2 #(
		.INIT('h8)
	) name23544 (
		\CM_rd2[22]_pad ,
		_w27000_,
		_w27591_
	);
	LUT2 #(
		.INIT('h8)
	) name23545 (
		\CM_rd5[22]_pad ,
		_w27004_,
		_w27592_
	);
	LUT2 #(
		.INIT('h8)
	) name23546 (
		\CM_rd4[22]_pad ,
		_w27008_,
		_w27593_
	);
	LUT2 #(
		.INIT('h8)
	) name23547 (
		\CM_rdm[22]_pad ,
		_w27018_,
		_w27594_
	);
	LUT2 #(
		.INIT('h8)
	) name23548 (
		\CM_rd3[22]_pad ,
		_w27011_,
		_w27595_
	);
	LUT2 #(
		.INIT('h1)
	) name23549 (
		_w27587_,
		_w27588_,
		_w27596_
	);
	LUT2 #(
		.INIT('h1)
	) name23550 (
		_w27589_,
		_w27590_,
		_w27597_
	);
	LUT2 #(
		.INIT('h1)
	) name23551 (
		_w27591_,
		_w27592_,
		_w27598_
	);
	LUT2 #(
		.INIT('h8)
	) name23552 (
		_w27597_,
		_w27598_,
		_w27599_
	);
	LUT2 #(
		.INIT('h4)
	) name23553 (
		_w27593_,
		_w27596_,
		_w27600_
	);
	LUT2 #(
		.INIT('h4)
	) name23554 (
		_w27595_,
		_w27600_,
		_w27601_
	);
	LUT2 #(
		.INIT('h8)
	) name23555 (
		_w27599_,
		_w27601_,
		_w27602_
	);
	LUT2 #(
		.INIT('h4)
	) name23556 (
		_w27594_,
		_w27602_,
		_w27603_
	);
	LUT2 #(
		.INIT('h2)
	) name23557 (
		_w27499_,
		_w27603_,
		_w27604_
	);
	LUT2 #(
		.INIT('h2)
	) name23558 (
		\idma_IADi_reg[14]/P0001 ,
		_w27499_,
		_w27605_
	);
	LUT2 #(
		.INIT('h1)
	) name23559 (
		_w27604_,
		_w27605_,
		_w27606_
	);
	LUT2 #(
		.INIT('h1)
	) name23560 (
		_w13570_,
		_w27606_,
		_w27607_
	);
	LUT2 #(
		.INIT('h8)
	) name23561 (
		_w12715_,
		_w13570_,
		_w27608_
	);
	LUT2 #(
		.INIT('h1)
	) name23562 (
		_w27607_,
		_w27608_,
		_w27609_
	);
	LUT2 #(
		.INIT('h1)
	) name23563 (
		_w11752_,
		_w27609_,
		_w27610_
	);
	LUT2 #(
		.INIT('h8)
	) name23564 (
		_w11752_,
		_w12688_,
		_w27611_
	);
	LUT2 #(
		.INIT('h1)
	) name23565 (
		_w27610_,
		_w27611_,
		_w27612_
	);
	LUT2 #(
		.INIT('h4)
	) name23566 (
		_w12520_,
		_w13570_,
		_w27613_
	);
	LUT2 #(
		.INIT('h2)
	) name23567 (
		_w13569_,
		_w27389_,
		_w27614_
	);
	LUT2 #(
		.INIT('h2)
	) name23568 (
		\idma_IADi_reg[0]/P0001 ,
		_w27499_,
		_w27615_
	);
	LUT2 #(
		.INIT('h1)
	) name23569 (
		_w13570_,
		_w27615_,
		_w27616_
	);
	LUT2 #(
		.INIT('h4)
	) name23570 (
		_w27614_,
		_w27616_,
		_w27617_
	);
	LUT2 #(
		.INIT('h1)
	) name23571 (
		_w11752_,
		_w27613_,
		_w27618_
	);
	LUT2 #(
		.INIT('h4)
	) name23572 (
		_w27617_,
		_w27618_,
		_w27619_
	);
	LUT2 #(
		.INIT('h8)
	) name23573 (
		_w7607_,
		_w11752_,
		_w27620_
	);
	LUT2 #(
		.INIT('h1)
	) name23574 (
		_w27619_,
		_w27620_,
		_w27621_
	);
	LUT2 #(
		.INIT('h2)
	) name23575 (
		\tm_TSR_TMP_reg[5]/NET0131 ,
		_w25494_,
		_w27622_
	);
	LUT2 #(
		.INIT('h1)
	) name23576 (
		_w25495_,
		_w27622_,
		_w27623_
	);
	LUT2 #(
		.INIT('h2)
	) name23577 (
		_w25491_,
		_w27623_,
		_w27624_
	);
	LUT2 #(
		.INIT('h2)
	) name23578 (
		\tm_tsr_reg_DO_reg[5]/NET0131 ,
		_w25491_,
		_w27625_
	);
	LUT2 #(
		.INIT('h1)
	) name23579 (
		_w27624_,
		_w27625_,
		_w27626_
	);
	LUT2 #(
		.INIT('h8)
	) name23580 (
		\CM_rd1[17]_pad ,
		_w26984_,
		_w27627_
	);
	LUT2 #(
		.INIT('h8)
	) name23581 (
		\CM_rd6[17]_pad ,
		_w26989_,
		_w27628_
	);
	LUT2 #(
		.INIT('h8)
	) name23582 (
		\CM_rd0[17]_pad ,
		_w26994_,
		_w27629_
	);
	LUT2 #(
		.INIT('h8)
	) name23583 (
		\CM_rd7[17]_pad ,
		_w26997_,
		_w27630_
	);
	LUT2 #(
		.INIT('h8)
	) name23584 (
		\CM_rd2[17]_pad ,
		_w27000_,
		_w27631_
	);
	LUT2 #(
		.INIT('h8)
	) name23585 (
		\CM_rd5[17]_pad ,
		_w27004_,
		_w27632_
	);
	LUT2 #(
		.INIT('h8)
	) name23586 (
		\CM_rd4[17]_pad ,
		_w27008_,
		_w27633_
	);
	LUT2 #(
		.INIT('h8)
	) name23587 (
		\CM_rdm[17]_pad ,
		_w27018_,
		_w27634_
	);
	LUT2 #(
		.INIT('h8)
	) name23588 (
		\CM_rd3[17]_pad ,
		_w27011_,
		_w27635_
	);
	LUT2 #(
		.INIT('h1)
	) name23589 (
		_w27627_,
		_w27628_,
		_w27636_
	);
	LUT2 #(
		.INIT('h1)
	) name23590 (
		_w27629_,
		_w27630_,
		_w27637_
	);
	LUT2 #(
		.INIT('h1)
	) name23591 (
		_w27631_,
		_w27632_,
		_w27638_
	);
	LUT2 #(
		.INIT('h8)
	) name23592 (
		_w27637_,
		_w27638_,
		_w27639_
	);
	LUT2 #(
		.INIT('h4)
	) name23593 (
		_w27633_,
		_w27636_,
		_w27640_
	);
	LUT2 #(
		.INIT('h4)
	) name23594 (
		_w27635_,
		_w27640_,
		_w27641_
	);
	LUT2 #(
		.INIT('h8)
	) name23595 (
		_w27639_,
		_w27641_,
		_w27642_
	);
	LUT2 #(
		.INIT('h4)
	) name23596 (
		_w27634_,
		_w27642_,
		_w27643_
	);
	LUT2 #(
		.INIT('h2)
	) name23597 (
		_w27499_,
		_w27643_,
		_w27644_
	);
	LUT2 #(
		.INIT('h2)
	) name23598 (
		\idma_IADi_reg[9]/P0001 ,
		_w27499_,
		_w27645_
	);
	LUT2 #(
		.INIT('h1)
	) name23599 (
		_w27644_,
		_w27645_,
		_w27646_
	);
	LUT2 #(
		.INIT('h1)
	) name23600 (
		_w13570_,
		_w27646_,
		_w27647_
	);
	LUT2 #(
		.INIT('h8)
	) name23601 (
		_w13075_,
		_w13570_,
		_w27648_
	);
	LUT2 #(
		.INIT('h1)
	) name23602 (
		_w27647_,
		_w27648_,
		_w27649_
	);
	LUT2 #(
		.INIT('h1)
	) name23603 (
		_w11752_,
		_w27649_,
		_w27650_
	);
	LUT2 #(
		.INIT('h8)
	) name23604 (
		_w10289_,
		_w11752_,
		_w27651_
	);
	LUT2 #(
		.INIT('h1)
	) name23605 (
		_w27650_,
		_w27651_,
		_w27652_
	);
	LUT2 #(
		.INIT('h8)
	) name23606 (
		\CM_rd1[16]_pad ,
		_w26984_,
		_w27653_
	);
	LUT2 #(
		.INIT('h8)
	) name23607 (
		\CM_rd6[16]_pad ,
		_w26989_,
		_w27654_
	);
	LUT2 #(
		.INIT('h8)
	) name23608 (
		\CM_rd0[16]_pad ,
		_w26994_,
		_w27655_
	);
	LUT2 #(
		.INIT('h8)
	) name23609 (
		\CM_rd7[16]_pad ,
		_w26997_,
		_w27656_
	);
	LUT2 #(
		.INIT('h8)
	) name23610 (
		\CM_rd2[16]_pad ,
		_w27000_,
		_w27657_
	);
	LUT2 #(
		.INIT('h8)
	) name23611 (
		\CM_rd5[16]_pad ,
		_w27004_,
		_w27658_
	);
	LUT2 #(
		.INIT('h8)
	) name23612 (
		\CM_rd4[16]_pad ,
		_w27008_,
		_w27659_
	);
	LUT2 #(
		.INIT('h8)
	) name23613 (
		\CM_rdm[16]_pad ,
		_w27018_,
		_w27660_
	);
	LUT2 #(
		.INIT('h8)
	) name23614 (
		\CM_rd3[16]_pad ,
		_w27011_,
		_w27661_
	);
	LUT2 #(
		.INIT('h1)
	) name23615 (
		_w27653_,
		_w27654_,
		_w27662_
	);
	LUT2 #(
		.INIT('h1)
	) name23616 (
		_w27655_,
		_w27656_,
		_w27663_
	);
	LUT2 #(
		.INIT('h1)
	) name23617 (
		_w27657_,
		_w27658_,
		_w27664_
	);
	LUT2 #(
		.INIT('h8)
	) name23618 (
		_w27663_,
		_w27664_,
		_w27665_
	);
	LUT2 #(
		.INIT('h4)
	) name23619 (
		_w27659_,
		_w27662_,
		_w27666_
	);
	LUT2 #(
		.INIT('h4)
	) name23620 (
		_w27661_,
		_w27666_,
		_w27667_
	);
	LUT2 #(
		.INIT('h8)
	) name23621 (
		_w27665_,
		_w27667_,
		_w27668_
	);
	LUT2 #(
		.INIT('h4)
	) name23622 (
		_w27660_,
		_w27668_,
		_w27669_
	);
	LUT2 #(
		.INIT('h2)
	) name23623 (
		_w27499_,
		_w27669_,
		_w27670_
	);
	LUT2 #(
		.INIT('h2)
	) name23624 (
		\idma_IADi_reg[8]/P0001 ,
		_w27499_,
		_w27671_
	);
	LUT2 #(
		.INIT('h1)
	) name23625 (
		_w27670_,
		_w27671_,
		_w27672_
	);
	LUT2 #(
		.INIT('h1)
	) name23626 (
		_w13570_,
		_w27672_,
		_w27673_
	);
	LUT2 #(
		.INIT('h8)
	) name23627 (
		_w13041_,
		_w13570_,
		_w27674_
	);
	LUT2 #(
		.INIT('h1)
	) name23628 (
		_w27673_,
		_w27674_,
		_w27675_
	);
	LUT2 #(
		.INIT('h1)
	) name23629 (
		_w11752_,
		_w27675_,
		_w27676_
	);
	LUT2 #(
		.INIT('h8)
	) name23630 (
		_w10638_,
		_w11752_,
		_w27677_
	);
	LUT2 #(
		.INIT('h1)
	) name23631 (
		_w27676_,
		_w27677_,
		_w27678_
	);
	LUT2 #(
		.INIT('h8)
	) name23632 (
		\CM_rd1[21]_pad ,
		_w26984_,
		_w27679_
	);
	LUT2 #(
		.INIT('h8)
	) name23633 (
		\CM_rd6[21]_pad ,
		_w26989_,
		_w27680_
	);
	LUT2 #(
		.INIT('h8)
	) name23634 (
		\CM_rd0[21]_pad ,
		_w26994_,
		_w27681_
	);
	LUT2 #(
		.INIT('h8)
	) name23635 (
		\CM_rd7[21]_pad ,
		_w26997_,
		_w27682_
	);
	LUT2 #(
		.INIT('h8)
	) name23636 (
		\CM_rd2[21]_pad ,
		_w27000_,
		_w27683_
	);
	LUT2 #(
		.INIT('h8)
	) name23637 (
		\CM_rd5[21]_pad ,
		_w27004_,
		_w27684_
	);
	LUT2 #(
		.INIT('h8)
	) name23638 (
		\CM_rd4[21]_pad ,
		_w27008_,
		_w27685_
	);
	LUT2 #(
		.INIT('h8)
	) name23639 (
		\CM_rdm[21]_pad ,
		_w27018_,
		_w27686_
	);
	LUT2 #(
		.INIT('h8)
	) name23640 (
		\CM_rd3[21]_pad ,
		_w27011_,
		_w27687_
	);
	LUT2 #(
		.INIT('h1)
	) name23641 (
		_w27679_,
		_w27680_,
		_w27688_
	);
	LUT2 #(
		.INIT('h1)
	) name23642 (
		_w27681_,
		_w27682_,
		_w27689_
	);
	LUT2 #(
		.INIT('h1)
	) name23643 (
		_w27683_,
		_w27684_,
		_w27690_
	);
	LUT2 #(
		.INIT('h8)
	) name23644 (
		_w27689_,
		_w27690_,
		_w27691_
	);
	LUT2 #(
		.INIT('h4)
	) name23645 (
		_w27685_,
		_w27688_,
		_w27692_
	);
	LUT2 #(
		.INIT('h4)
	) name23646 (
		_w27687_,
		_w27692_,
		_w27693_
	);
	LUT2 #(
		.INIT('h8)
	) name23647 (
		_w27691_,
		_w27693_,
		_w27694_
	);
	LUT2 #(
		.INIT('h4)
	) name23648 (
		_w27686_,
		_w27694_,
		_w27695_
	);
	LUT2 #(
		.INIT('h2)
	) name23649 (
		_w27499_,
		_w27695_,
		_w27696_
	);
	LUT2 #(
		.INIT('h2)
	) name23650 (
		\idma_IADi_reg[13]/P0001 ,
		_w27499_,
		_w27697_
	);
	LUT2 #(
		.INIT('h1)
	) name23651 (
		_w27696_,
		_w27697_,
		_w27698_
	);
	LUT2 #(
		.INIT('h1)
	) name23652 (
		_w13570_,
		_w27698_,
		_w27699_
	);
	LUT2 #(
		.INIT('h8)
	) name23653 (
		_w12658_,
		_w13570_,
		_w27700_
	);
	LUT2 #(
		.INIT('h1)
	) name23654 (
		_w27699_,
		_w27700_,
		_w27701_
	);
	LUT2 #(
		.INIT('h1)
	) name23655 (
		_w11752_,
		_w27701_,
		_w27702_
	);
	LUT2 #(
		.INIT('h8)
	) name23656 (
		_w7340_,
		_w11752_,
		_w27703_
	);
	LUT2 #(
		.INIT('h1)
	) name23657 (
		_w27702_,
		_w27703_,
		_w27704_
	);
	LUT2 #(
		.INIT('h8)
	) name23658 (
		\CM_rd1[20]_pad ,
		_w26984_,
		_w27705_
	);
	LUT2 #(
		.INIT('h8)
	) name23659 (
		\CM_rd6[20]_pad ,
		_w26989_,
		_w27706_
	);
	LUT2 #(
		.INIT('h8)
	) name23660 (
		\CM_rd0[20]_pad ,
		_w26994_,
		_w27707_
	);
	LUT2 #(
		.INIT('h8)
	) name23661 (
		\CM_rd7[20]_pad ,
		_w26997_,
		_w27708_
	);
	LUT2 #(
		.INIT('h8)
	) name23662 (
		\CM_rd2[20]_pad ,
		_w27000_,
		_w27709_
	);
	LUT2 #(
		.INIT('h8)
	) name23663 (
		\CM_rd5[20]_pad ,
		_w27004_,
		_w27710_
	);
	LUT2 #(
		.INIT('h8)
	) name23664 (
		\CM_rd4[20]_pad ,
		_w27008_,
		_w27711_
	);
	LUT2 #(
		.INIT('h8)
	) name23665 (
		\CM_rdm[20]_pad ,
		_w27018_,
		_w27712_
	);
	LUT2 #(
		.INIT('h8)
	) name23666 (
		\CM_rd3[20]_pad ,
		_w27011_,
		_w27713_
	);
	LUT2 #(
		.INIT('h1)
	) name23667 (
		_w27705_,
		_w27706_,
		_w27714_
	);
	LUT2 #(
		.INIT('h1)
	) name23668 (
		_w27707_,
		_w27708_,
		_w27715_
	);
	LUT2 #(
		.INIT('h1)
	) name23669 (
		_w27709_,
		_w27710_,
		_w27716_
	);
	LUT2 #(
		.INIT('h8)
	) name23670 (
		_w27715_,
		_w27716_,
		_w27717_
	);
	LUT2 #(
		.INIT('h4)
	) name23671 (
		_w27711_,
		_w27714_,
		_w27718_
	);
	LUT2 #(
		.INIT('h4)
	) name23672 (
		_w27713_,
		_w27718_,
		_w27719_
	);
	LUT2 #(
		.INIT('h8)
	) name23673 (
		_w27717_,
		_w27719_,
		_w27720_
	);
	LUT2 #(
		.INIT('h4)
	) name23674 (
		_w27712_,
		_w27720_,
		_w27721_
	);
	LUT2 #(
		.INIT('h2)
	) name23675 (
		_w27499_,
		_w27721_,
		_w27722_
	);
	LUT2 #(
		.INIT('h2)
	) name23676 (
		\idma_IADi_reg[12]/P0001 ,
		_w27499_,
		_w27723_
	);
	LUT2 #(
		.INIT('h1)
	) name23677 (
		_w27722_,
		_w27723_,
		_w27724_
	);
	LUT2 #(
		.INIT('h1)
	) name23678 (
		_w13570_,
		_w27724_,
		_w27725_
	);
	LUT2 #(
		.INIT('h8)
	) name23679 (
		_w12624_,
		_w13570_,
		_w27726_
	);
	LUT2 #(
		.INIT('h1)
	) name23680 (
		_w27725_,
		_w27726_,
		_w27727_
	);
	LUT2 #(
		.INIT('h1)
	) name23681 (
		_w11752_,
		_w27727_,
		_w27728_
	);
	LUT2 #(
		.INIT('h8)
	) name23682 (
		_w9178_,
		_w11752_,
		_w27729_
	);
	LUT2 #(
		.INIT('h1)
	) name23683 (
		_w27728_,
		_w27729_,
		_w27730_
	);
	LUT2 #(
		.INIT('h8)
	) name23684 (
		\CM_rd1[19]_pad ,
		_w26984_,
		_w27731_
	);
	LUT2 #(
		.INIT('h8)
	) name23685 (
		\CM_rd6[19]_pad ,
		_w26989_,
		_w27732_
	);
	LUT2 #(
		.INIT('h8)
	) name23686 (
		\CM_rd0[19]_pad ,
		_w26994_,
		_w27733_
	);
	LUT2 #(
		.INIT('h8)
	) name23687 (
		\CM_rd7[19]_pad ,
		_w26997_,
		_w27734_
	);
	LUT2 #(
		.INIT('h8)
	) name23688 (
		\CM_rd2[19]_pad ,
		_w27000_,
		_w27735_
	);
	LUT2 #(
		.INIT('h8)
	) name23689 (
		\CM_rd5[19]_pad ,
		_w27004_,
		_w27736_
	);
	LUT2 #(
		.INIT('h8)
	) name23690 (
		\CM_rd4[19]_pad ,
		_w27008_,
		_w27737_
	);
	LUT2 #(
		.INIT('h8)
	) name23691 (
		\CM_rdm[19]_pad ,
		_w27018_,
		_w27738_
	);
	LUT2 #(
		.INIT('h8)
	) name23692 (
		\CM_rd3[19]_pad ,
		_w27011_,
		_w27739_
	);
	LUT2 #(
		.INIT('h1)
	) name23693 (
		_w27731_,
		_w27732_,
		_w27740_
	);
	LUT2 #(
		.INIT('h1)
	) name23694 (
		_w27733_,
		_w27734_,
		_w27741_
	);
	LUT2 #(
		.INIT('h1)
	) name23695 (
		_w27735_,
		_w27736_,
		_w27742_
	);
	LUT2 #(
		.INIT('h8)
	) name23696 (
		_w27741_,
		_w27742_,
		_w27743_
	);
	LUT2 #(
		.INIT('h4)
	) name23697 (
		_w27737_,
		_w27740_,
		_w27744_
	);
	LUT2 #(
		.INIT('h4)
	) name23698 (
		_w27739_,
		_w27744_,
		_w27745_
	);
	LUT2 #(
		.INIT('h8)
	) name23699 (
		_w27743_,
		_w27745_,
		_w27746_
	);
	LUT2 #(
		.INIT('h4)
	) name23700 (
		_w27738_,
		_w27746_,
		_w27747_
	);
	LUT2 #(
		.INIT('h2)
	) name23701 (
		_w27499_,
		_w27747_,
		_w27748_
	);
	LUT2 #(
		.INIT('h2)
	) name23702 (
		\idma_IADi_reg[11]/P0001 ,
		_w27499_,
		_w27749_
	);
	LUT2 #(
		.INIT('h1)
	) name23703 (
		_w27748_,
		_w27749_,
		_w27750_
	);
	LUT2 #(
		.INIT('h1)
	) name23704 (
		_w13570_,
		_w27750_,
		_w27751_
	);
	LUT2 #(
		.INIT('h8)
	) name23705 (
		_w12590_,
		_w13570_,
		_w27752_
	);
	LUT2 #(
		.INIT('h1)
	) name23706 (
		_w27751_,
		_w27752_,
		_w27753_
	);
	LUT2 #(
		.INIT('h1)
	) name23707 (
		_w11752_,
		_w27753_,
		_w27754_
	);
	LUT2 #(
		.INIT('h8)
	) name23708 (
		_w8460_,
		_w11752_,
		_w27755_
	);
	LUT2 #(
		.INIT('h1)
	) name23709 (
		_w27754_,
		_w27755_,
		_w27756_
	);
	LUT2 #(
		.INIT('h8)
	) name23710 (
		\CM_rd1[18]_pad ,
		_w26984_,
		_w27757_
	);
	LUT2 #(
		.INIT('h8)
	) name23711 (
		\CM_rd6[18]_pad ,
		_w26989_,
		_w27758_
	);
	LUT2 #(
		.INIT('h8)
	) name23712 (
		\CM_rd0[18]_pad ,
		_w26994_,
		_w27759_
	);
	LUT2 #(
		.INIT('h8)
	) name23713 (
		\CM_rd7[18]_pad ,
		_w26997_,
		_w27760_
	);
	LUT2 #(
		.INIT('h8)
	) name23714 (
		\CM_rd2[18]_pad ,
		_w27000_,
		_w27761_
	);
	LUT2 #(
		.INIT('h8)
	) name23715 (
		\CM_rd5[18]_pad ,
		_w27004_,
		_w27762_
	);
	LUT2 #(
		.INIT('h8)
	) name23716 (
		\CM_rd4[18]_pad ,
		_w27008_,
		_w27763_
	);
	LUT2 #(
		.INIT('h8)
	) name23717 (
		\CM_rdm[18]_pad ,
		_w27018_,
		_w27764_
	);
	LUT2 #(
		.INIT('h8)
	) name23718 (
		\CM_rd3[18]_pad ,
		_w27011_,
		_w27765_
	);
	LUT2 #(
		.INIT('h1)
	) name23719 (
		_w27757_,
		_w27758_,
		_w27766_
	);
	LUT2 #(
		.INIT('h1)
	) name23720 (
		_w27759_,
		_w27760_,
		_w27767_
	);
	LUT2 #(
		.INIT('h1)
	) name23721 (
		_w27761_,
		_w27762_,
		_w27768_
	);
	LUT2 #(
		.INIT('h8)
	) name23722 (
		_w27767_,
		_w27768_,
		_w27769_
	);
	LUT2 #(
		.INIT('h4)
	) name23723 (
		_w27763_,
		_w27766_,
		_w27770_
	);
	LUT2 #(
		.INIT('h4)
	) name23724 (
		_w27765_,
		_w27770_,
		_w27771_
	);
	LUT2 #(
		.INIT('h8)
	) name23725 (
		_w27769_,
		_w27771_,
		_w27772_
	);
	LUT2 #(
		.INIT('h4)
	) name23726 (
		_w27764_,
		_w27772_,
		_w27773_
	);
	LUT2 #(
		.INIT('h2)
	) name23727 (
		_w27499_,
		_w27773_,
		_w27774_
	);
	LUT2 #(
		.INIT('h2)
	) name23728 (
		\idma_IADi_reg[10]/P0001 ,
		_w27499_,
		_w27775_
	);
	LUT2 #(
		.INIT('h1)
	) name23729 (
		_w27774_,
		_w27775_,
		_w27776_
	);
	LUT2 #(
		.INIT('h1)
	) name23730 (
		_w13570_,
		_w27776_,
		_w27777_
	);
	LUT2 #(
		.INIT('h8)
	) name23731 (
		_w12556_,
		_w13570_,
		_w27778_
	);
	LUT2 #(
		.INIT('h1)
	) name23732 (
		_w27777_,
		_w27778_,
		_w27779_
	);
	LUT2 #(
		.INIT('h1)
	) name23733 (
		_w11752_,
		_w27779_,
		_w27780_
	);
	LUT2 #(
		.INIT('h8)
	) name23734 (
		_w7859_,
		_w11752_,
		_w27781_
	);
	LUT2 #(
		.INIT('h1)
	) name23735 (
		_w27780_,
		_w27781_,
		_w27782_
	);
	LUT2 #(
		.INIT('h1)
	) name23736 (
		_w6931_,
		_w6988_,
		_w27783_
	);
	LUT2 #(
		.INIT('h1)
	) name23737 (
		_w13567_,
		_w27783_,
		_w27784_
	);
	LUT2 #(
		.INIT('h2)
	) name23738 (
		_w13564_,
		_w27784_,
		_w27785_
	);
	LUT2 #(
		.INIT('h2)
	) name23739 (
		_w13597_,
		_w27785_,
		_w27786_
	);
	LUT2 #(
		.INIT('h1)
	) name23740 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 ,
		_w19499_,
		_w27787_
	);
	LUT2 #(
		.INIT('h4)
	) name23741 (
		_w17814_,
		_w19499_,
		_w27788_
	);
	LUT2 #(
		.INIT('h2)
	) name23742 (
		_w19501_,
		_w27787_,
		_w27789_
	);
	LUT2 #(
		.INIT('h4)
	) name23743 (
		_w27788_,
		_w27789_,
		_w27790_
	);
	LUT2 #(
		.INIT('h2)
	) name23744 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[2]/P0001 ,
		_w19383_,
		_w27791_
	);
	LUT2 #(
		.INIT('h1)
	) name23745 (
		_w19508_,
		_w27791_,
		_w27792_
	);
	LUT2 #(
		.INIT('h4)
	) name23746 (
		_w27790_,
		_w27792_,
		_w27793_
	);
	LUT2 #(
		.INIT('h1)
	) name23747 (
		_w18262_,
		_w27793_,
		_w27794_
	);
	LUT2 #(
		.INIT('h1)
	) name23748 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w27051_,
		_w27795_
	);
	LUT2 #(
		.INIT('h1)
	) name23749 (
		_w17613_,
		_w17672_,
		_w27796_
	);
	LUT2 #(
		.INIT('h1)
	) name23750 (
		_w17638_,
		_w27048_,
		_w27797_
	);
	LUT2 #(
		.INIT('h1)
	) name23751 (
		_w17665_,
		_w27797_,
		_w27798_
	);
	LUT2 #(
		.INIT('h2)
	) name23752 (
		_w27796_,
		_w27798_,
		_w27799_
	);
	LUT2 #(
		.INIT('h4)
	) name23753 (
		_w27796_,
		_w27798_,
		_w27800_
	);
	LUT2 #(
		.INIT('h1)
	) name23754 (
		_w27799_,
		_w27800_,
		_w27801_
	);
	LUT2 #(
		.INIT('h2)
	) name23755 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w27801_,
		_w27802_
	);
	LUT2 #(
		.INIT('h1)
	) name23756 (
		_w27795_,
		_w27802_,
		_w27803_
	);
	LUT2 #(
		.INIT('h8)
	) name23757 (
		_w18262_,
		_w27803_,
		_w27804_
	);
	LUT2 #(
		.INIT('h1)
	) name23758 (
		_w27794_,
		_w27804_,
		_w27805_
	);
	LUT2 #(
		.INIT('h1)
	) name23759 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 ,
		_w19499_,
		_w27806_
	);
	LUT2 #(
		.INIT('h2)
	) name23760 (
		_w19499_,
		_w21663_,
		_w27807_
	);
	LUT2 #(
		.INIT('h2)
	) name23761 (
		_w19501_,
		_w27806_,
		_w27808_
	);
	LUT2 #(
		.INIT('h4)
	) name23762 (
		_w27807_,
		_w27808_,
		_w27809_
	);
	LUT2 #(
		.INIT('h2)
	) name23763 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[3]/P0001 ,
		_w19383_,
		_w27810_
	);
	LUT2 #(
		.INIT('h1)
	) name23764 (
		_w19508_,
		_w27810_,
		_w27811_
	);
	LUT2 #(
		.INIT('h4)
	) name23765 (
		_w27809_,
		_w27811_,
		_w27812_
	);
	LUT2 #(
		.INIT('h1)
	) name23766 (
		_w18262_,
		_w27812_,
		_w27813_
	);
	LUT2 #(
		.INIT('h4)
	) name23767 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w27801_,
		_w27814_
	);
	LUT2 #(
		.INIT('h8)
	) name23768 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w26315_,
		_w27815_
	);
	LUT2 #(
		.INIT('h1)
	) name23769 (
		_w27814_,
		_w27815_,
		_w27816_
	);
	LUT2 #(
		.INIT('h2)
	) name23770 (
		_w18262_,
		_w27816_,
		_w27817_
	);
	LUT2 #(
		.INIT('h1)
	) name23771 (
		_w27813_,
		_w27817_,
		_w27818_
	);
	LUT2 #(
		.INIT('h8)
	) name23772 (
		_w14752_,
		_w27816_,
		_w27819_
	);
	LUT2 #(
		.INIT('h8)
	) name23773 (
		_w19776_,
		_w21663_,
		_w27820_
	);
	LUT2 #(
		.INIT('h2)
	) name23774 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[3]/P0001 ,
		_w17809_,
		_w27821_
	);
	LUT2 #(
		.INIT('h2)
	) name23775 (
		_w19780_,
		_w27821_,
		_w27822_
	);
	LUT2 #(
		.INIT('h4)
	) name23776 (
		_w27820_,
		_w27822_,
		_w27823_
	);
	LUT2 #(
		.INIT('h1)
	) name23777 (
		_w27819_,
		_w27823_,
		_w27824_
	);
	LUT2 #(
		.INIT('h2)
	) name23778 (
		_w14752_,
		_w27803_,
		_w27825_
	);
	LUT2 #(
		.INIT('h8)
	) name23779 (
		_w17814_,
		_w19776_,
		_w27826_
	);
	LUT2 #(
		.INIT('h2)
	) name23780 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[2]/P0001 ,
		_w17809_,
		_w27827_
	);
	LUT2 #(
		.INIT('h2)
	) name23781 (
		_w19780_,
		_w27827_,
		_w27828_
	);
	LUT2 #(
		.INIT('h4)
	) name23782 (
		_w27826_,
		_w27828_,
		_w27829_
	);
	LUT2 #(
		.INIT('h1)
	) name23783 (
		_w27825_,
		_w27829_,
		_w27830_
	);
	LUT2 #(
		.INIT('h2)
	) name23784 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 ,
		_w18266_,
		_w27831_
	);
	LUT2 #(
		.INIT('h1)
	) name23785 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[14]/P0001 ,
		_w18271_,
		_w27832_
	);
	LUT2 #(
		.INIT('h2)
	) name23786 (
		_w18271_,
		_w20150_,
		_w27833_
	);
	LUT2 #(
		.INIT('h2)
	) name23787 (
		_w18273_,
		_w27832_,
		_w27834_
	);
	LUT2 #(
		.INIT('h4)
	) name23788 (
		_w27833_,
		_w27834_,
		_w27835_
	);
	LUT2 #(
		.INIT('h1)
	) name23789 (
		_w18270_,
		_w27831_,
		_w27836_
	);
	LUT2 #(
		.INIT('h4)
	) name23790 (
		_w27835_,
		_w27836_,
		_w27837_
	);
	LUT2 #(
		.INIT('h1)
	) name23791 (
		_w18262_,
		_w27837_,
		_w27838_
	);
	LUT2 #(
		.INIT('h2)
	) name23792 (
		_w18262_,
		_w19593_,
		_w27839_
	);
	LUT2 #(
		.INIT('h1)
	) name23793 (
		_w27838_,
		_w27839_,
		_w27840_
	);
	LUT2 #(
		.INIT('h8)
	) name23794 (
		_w14752_,
		_w19593_,
		_w27841_
	);
	LUT2 #(
		.INIT('h8)
	) name23795 (
		_w18328_,
		_w20150_,
		_w27842_
	);
	LUT2 #(
		.INIT('h2)
	) name23796 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[14]/P0001 ,
		_w18330_,
		_w27843_
	);
	LUT2 #(
		.INIT('h2)
	) name23797 (
		_w18334_,
		_w27843_,
		_w27844_
	);
	LUT2 #(
		.INIT('h4)
	) name23798 (
		_w27842_,
		_w27844_,
		_w27845_
	);
	LUT2 #(
		.INIT('h1)
	) name23799 (
		_w27841_,
		_w27845_,
		_w27846_
	);
	LUT2 #(
		.INIT('h2)
	) name23800 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 ,
		_w18266_,
		_w27847_
	);
	LUT2 #(
		.INIT('h1)
	) name23801 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[2]/P0001 ,
		_w18271_,
		_w27848_
	);
	LUT2 #(
		.INIT('h4)
	) name23802 (
		_w17814_,
		_w18271_,
		_w27849_
	);
	LUT2 #(
		.INIT('h2)
	) name23803 (
		_w18273_,
		_w27848_,
		_w27850_
	);
	LUT2 #(
		.INIT('h4)
	) name23804 (
		_w27849_,
		_w27850_,
		_w27851_
	);
	LUT2 #(
		.INIT('h1)
	) name23805 (
		_w18270_,
		_w27847_,
		_w27852_
	);
	LUT2 #(
		.INIT('h4)
	) name23806 (
		_w27851_,
		_w27852_,
		_w27853_
	);
	LUT2 #(
		.INIT('h1)
	) name23807 (
		_w18262_,
		_w27853_,
		_w27854_
	);
	LUT2 #(
		.INIT('h2)
	) name23808 (
		_w18262_,
		_w19673_,
		_w27855_
	);
	LUT2 #(
		.INIT('h1)
	) name23809 (
		_w27854_,
		_w27855_,
		_w27856_
	);
	LUT2 #(
		.INIT('h8)
	) name23810 (
		_w14752_,
		_w19673_,
		_w27857_
	);
	LUT2 #(
		.INIT('h8)
	) name23811 (
		_w17814_,
		_w18328_,
		_w27858_
	);
	LUT2 #(
		.INIT('h2)
	) name23812 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[2]/P0001 ,
		_w18330_,
		_w27859_
	);
	LUT2 #(
		.INIT('h2)
	) name23813 (
		_w18334_,
		_w27859_,
		_w27860_
	);
	LUT2 #(
		.INIT('h4)
	) name23814 (
		_w27858_,
		_w27860_,
		_w27861_
	);
	LUT2 #(
		.INIT('h1)
	) name23815 (
		_w27857_,
		_w27861_,
		_w27862_
	);
	LUT2 #(
		.INIT('h2)
	) name23816 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 ,
		_w18266_,
		_w27863_
	);
	LUT2 #(
		.INIT('h1)
	) name23817 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[15]/P0001 ,
		_w18271_,
		_w27864_
	);
	LUT2 #(
		.INIT('h4)
	) name23818 (
		_w17820_,
		_w18271_,
		_w27865_
	);
	LUT2 #(
		.INIT('h2)
	) name23819 (
		_w18273_,
		_w27864_,
		_w27866_
	);
	LUT2 #(
		.INIT('h4)
	) name23820 (
		_w27865_,
		_w27866_,
		_w27867_
	);
	LUT2 #(
		.INIT('h1)
	) name23821 (
		_w18270_,
		_w27863_,
		_w27868_
	);
	LUT2 #(
		.INIT('h4)
	) name23822 (
		_w27867_,
		_w27868_,
		_w27869_
	);
	LUT2 #(
		.INIT('h1)
	) name23823 (
		_w18262_,
		_w27869_,
		_w27870_
	);
	LUT2 #(
		.INIT('h2)
	) name23824 (
		_w18262_,
		_w19596_,
		_w27871_
	);
	LUT2 #(
		.INIT('h1)
	) name23825 (
		_w27870_,
		_w27871_,
		_w27872_
	);
	LUT2 #(
		.INIT('h4)
	) name23826 (
		_w13806_,
		_w14564_,
		_w27873_
	);
	LUT2 #(
		.INIT('h8)
	) name23827 (
		_w11975_,
		_w13806_,
		_w27874_
	);
	LUT2 #(
		.INIT('h1)
	) name23828 (
		_w27873_,
		_w27874_,
		_w27875_
	);
	LUT2 #(
		.INIT('h2)
	) name23829 (
		_w14667_,
		_w27875_,
		_w27876_
	);
	LUT2 #(
		.INIT('h1)
	) name23830 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[0]/P0001 ,
		_w14667_,
		_w27877_
	);
	LUT2 #(
		.INIT('h1)
	) name23831 (
		_w27876_,
		_w27877_,
		_w27878_
	);
	LUT2 #(
		.INIT('h2)
	) name23832 (
		_w13805_,
		_w27875_,
		_w27879_
	);
	LUT2 #(
		.INIT('h1)
	) name23833 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[0]/P0001 ,
		_w13805_,
		_w27880_
	);
	LUT2 #(
		.INIT('h1)
	) name23834 (
		_w27879_,
		_w27880_,
		_w27881_
	);
	LUT2 #(
		.INIT('h8)
	) name23835 (
		_w14752_,
		_w19596_,
		_w27882_
	);
	LUT2 #(
		.INIT('h8)
	) name23836 (
		_w17820_,
		_w18328_,
		_w27883_
	);
	LUT2 #(
		.INIT('h2)
	) name23837 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[15]/P0001 ,
		_w18330_,
		_w27884_
	);
	LUT2 #(
		.INIT('h2)
	) name23838 (
		_w18334_,
		_w27884_,
		_w27885_
	);
	LUT2 #(
		.INIT('h4)
	) name23839 (
		_w27883_,
		_w27885_,
		_w27886_
	);
	LUT2 #(
		.INIT('h1)
	) name23840 (
		_w27882_,
		_w27886_,
		_w27887_
	);
	LUT2 #(
		.INIT('h8)
	) name23841 (
		\tm_tcr_reg_DO_reg[7]/NET0131 ,
		_w20355_,
		_w27888_
	);
	LUT2 #(
		.INIT('h4)
	) name23842 (
		\tm_tpr_reg_DO_reg[7]/NET0131 ,
		_w22400_,
		_w27889_
	);
	LUT2 #(
		.INIT('h1)
	) name23843 (
		\T_TMODE[0]_pad ,
		_w20360_,
		_w27890_
	);
	LUT2 #(
		.INIT('h2)
	) name23844 (
		_w20363_,
		_w27890_,
		_w27891_
	);
	LUT2 #(
		.INIT('h8)
	) name23845 (
		_w22411_,
		_w27891_,
		_w27892_
	);
	LUT2 #(
		.INIT('h1)
	) name23846 (
		\tm_TCR_TMP_reg[4]/NET0131 ,
		_w27890_,
		_w27893_
	);
	LUT2 #(
		.INIT('h4)
	) name23847 (
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w27893_,
		_w27894_
	);
	LUT2 #(
		.INIT('h8)
	) name23848 (
		_w22411_,
		_w27894_,
		_w27895_
	);
	LUT2 #(
		.INIT('h4)
	) name23849 (
		\tm_TCR_TMP_reg[6]/NET0131 ,
		_w27895_,
		_w27896_
	);
	LUT2 #(
		.INIT('h2)
	) name23850 (
		\tm_TCR_TMP_reg[7]/NET0131 ,
		_w27896_,
		_w27897_
	);
	LUT2 #(
		.INIT('h1)
	) name23851 (
		_w22400_,
		_w27892_,
		_w27898_
	);
	LUT2 #(
		.INIT('h4)
	) name23852 (
		_w27897_,
		_w27898_,
		_w27899_
	);
	LUT2 #(
		.INIT('h1)
	) name23853 (
		_w20355_,
		_w27889_,
		_w27900_
	);
	LUT2 #(
		.INIT('h4)
	) name23854 (
		_w27899_,
		_w27900_,
		_w27901_
	);
	LUT2 #(
		.INIT('h1)
	) name23855 (
		_w27888_,
		_w27901_,
		_w27902_
	);
	LUT2 #(
		.INIT('h8)
	) name23856 (
		_w23407_,
		_w25053_,
		_w27903_
	);
	LUT2 #(
		.INIT('h8)
	) name23857 (
		_w23032_,
		_w27903_,
		_w27904_
	);
	LUT2 #(
		.INIT('h8)
	) name23858 (
		_w25749_,
		_w25752_,
		_w27905_
	);
	LUT2 #(
		.INIT('h8)
	) name23859 (
		_w4186_,
		_w27905_,
		_w27906_
	);
	LUT2 #(
		.INIT('h8)
	) name23860 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w27907_
	);
	LUT2 #(
		.INIT('h1)
	) name23861 (
		\core_c_dec_MTCNTR_Eg_reg/P0001 ,
		\core_c_dec_MTOWRCNTR_Eg_reg/P0001 ,
		_w27908_
	);
	LUT2 #(
		.INIT('h2)
	) name23862 (
		\core_c_dec_BR_Ed_reg/P0001 ,
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w27909_
	);
	LUT2 #(
		.INIT('h8)
	) name23863 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w27909_,
		_w27910_
	);
	LUT2 #(
		.INIT('h8)
	) name23864 (
		_w6071_,
		_w27910_,
		_w27911_
	);
	LUT2 #(
		.INIT('h4)
	) name23865 (
		_w27907_,
		_w27908_,
		_w27912_
	);
	LUT2 #(
		.INIT('h4)
	) name23866 (
		_w27911_,
		_w27912_,
		_w27913_
	);
	LUT2 #(
		.INIT('h4)
	) name23867 (
		_w27906_,
		_w27913_,
		_w27914_
	);
	LUT2 #(
		.INIT('h1)
	) name23868 (
		_w5950_,
		_w27914_,
		_w27915_
	);
	LUT2 #(
		.INIT('h2)
	) name23869 (
		\core_c_psq_CE_reg/NET0131 ,
		_w27915_,
		_w27916_
	);
	LUT2 #(
		.INIT('h8)
	) name23870 (
		\core_c_psq_CE_reg/NET0131 ,
		_w27911_,
		_w27917_
	);
	LUT2 #(
		.INIT('h8)
	) name23871 (
		_w4842_,
		_w27905_,
		_w27918_
	);
	LUT2 #(
		.INIT('h1)
	) name23872 (
		_w27907_,
		_w27917_,
		_w27919_
	);
	LUT2 #(
		.INIT('h4)
	) name23873 (
		_w27918_,
		_w27919_,
		_w27920_
	);
	LUT2 #(
		.INIT('h1)
	) name23874 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w27920_,
		_w27921_
	);
	LUT2 #(
		.INIT('h1)
	) name23875 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w27922_
	);
	LUT2 #(
		.INIT('h4)
	) name23876 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w27922_,
		_w27923_
	);
	LUT2 #(
		.INIT('h4)
	) name23877 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w27923_,
		_w27924_
	);
	LUT2 #(
		.INIT('h4)
	) name23878 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w27924_,
		_w27925_
	);
	LUT2 #(
		.INIT('h4)
	) name23879 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w27925_,
		_w27926_
	);
	LUT2 #(
		.INIT('h4)
	) name23880 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w27926_,
		_w27927_
	);
	LUT2 #(
		.INIT('h4)
	) name23881 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w27927_,
		_w27928_
	);
	LUT2 #(
		.INIT('h4)
	) name23882 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w27928_,
		_w27929_
	);
	LUT2 #(
		.INIT('h4)
	) name23883 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w27929_,
		_w27930_
	);
	LUT2 #(
		.INIT('h4)
	) name23884 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w27930_,
		_w27931_
	);
	LUT2 #(
		.INIT('h4)
	) name23885 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w27931_,
		_w27932_
	);
	LUT2 #(
		.INIT('h4)
	) name23886 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w27932_,
		_w27933_
	);
	LUT2 #(
		.INIT('h2)
	) name23887 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w27932_,
		_w27934_
	);
	LUT2 #(
		.INIT('h1)
	) name23888 (
		_w27933_,
		_w27934_,
		_w27935_
	);
	LUT2 #(
		.INIT('h1)
	) name23889 (
		_w27921_,
		_w27935_,
		_w27936_
	);
	LUT2 #(
		.INIT('h8)
	) name23890 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][12]/P0001 ,
		_w13775_,
		_w27937_
	);
	LUT2 #(
		.INIT('h8)
	) name23891 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][12]/P0001 ,
		_w13789_,
		_w27938_
	);
	LUT2 #(
		.INIT('h8)
	) name23892 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][12]/P0001 ,
		_w13794_,
		_w27939_
	);
	LUT2 #(
		.INIT('h8)
	) name23893 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][12]/P0001 ,
		_w13784_,
		_w27940_
	);
	LUT2 #(
		.INIT('h1)
	) name23894 (
		_w27937_,
		_w27938_,
		_w27941_
	);
	LUT2 #(
		.INIT('h1)
	) name23895 (
		_w27939_,
		_w27940_,
		_w27942_
	);
	LUT2 #(
		.INIT('h8)
	) name23896 (
		_w27941_,
		_w27942_,
		_w27943_
	);
	LUT2 #(
		.INIT('h2)
	) name23897 (
		_w27921_,
		_w27943_,
		_w27944_
	);
	LUT2 #(
		.INIT('h1)
	) name23898 (
		_w27936_,
		_w27944_,
		_w27945_
	);
	LUT2 #(
		.INIT('h2)
	) name23899 (
		_w27908_,
		_w27945_,
		_w27946_
	);
	LUT2 #(
		.INIT('h2)
	) name23900 (
		_w9178_,
		_w27908_,
		_w27947_
	);
	LUT2 #(
		.INIT('h1)
	) name23901 (
		_w27946_,
		_w27947_,
		_w27948_
	);
	LUT2 #(
		.INIT('h2)
	) name23902 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w27930_,
		_w27949_
	);
	LUT2 #(
		.INIT('h1)
	) name23903 (
		_w27931_,
		_w27949_,
		_w27950_
	);
	LUT2 #(
		.INIT('h1)
	) name23904 (
		_w27921_,
		_w27950_,
		_w27951_
	);
	LUT2 #(
		.INIT('h8)
	) name23905 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][10]/P0001 ,
		_w13775_,
		_w27952_
	);
	LUT2 #(
		.INIT('h8)
	) name23906 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][10]/P0001 ,
		_w13784_,
		_w27953_
	);
	LUT2 #(
		.INIT('h8)
	) name23907 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][10]/P0001 ,
		_w13789_,
		_w27954_
	);
	LUT2 #(
		.INIT('h8)
	) name23908 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][10]/P0001 ,
		_w13794_,
		_w27955_
	);
	LUT2 #(
		.INIT('h1)
	) name23909 (
		_w27952_,
		_w27953_,
		_w27956_
	);
	LUT2 #(
		.INIT('h1)
	) name23910 (
		_w27954_,
		_w27955_,
		_w27957_
	);
	LUT2 #(
		.INIT('h8)
	) name23911 (
		_w27956_,
		_w27957_,
		_w27958_
	);
	LUT2 #(
		.INIT('h2)
	) name23912 (
		_w27921_,
		_w27958_,
		_w27959_
	);
	LUT2 #(
		.INIT('h1)
	) name23913 (
		_w27951_,
		_w27959_,
		_w27960_
	);
	LUT2 #(
		.INIT('h2)
	) name23914 (
		_w27908_,
		_w27960_,
		_w27961_
	);
	LUT2 #(
		.INIT('h2)
	) name23915 (
		_w7859_,
		_w27908_,
		_w27962_
	);
	LUT2 #(
		.INIT('h1)
	) name23916 (
		_w27961_,
		_w27962_,
		_w27963_
	);
	LUT2 #(
		.INIT('h2)
	) name23917 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w27928_,
		_w27964_
	);
	LUT2 #(
		.INIT('h1)
	) name23918 (
		_w27929_,
		_w27964_,
		_w27965_
	);
	LUT2 #(
		.INIT('h1)
	) name23919 (
		_w27921_,
		_w27965_,
		_w27966_
	);
	LUT2 #(
		.INIT('h8)
	) name23920 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][8]/P0001 ,
		_w13775_,
		_w27967_
	);
	LUT2 #(
		.INIT('h8)
	) name23921 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][8]/P0001 ,
		_w13794_,
		_w27968_
	);
	LUT2 #(
		.INIT('h8)
	) name23922 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][8]/P0001 ,
		_w13789_,
		_w27969_
	);
	LUT2 #(
		.INIT('h8)
	) name23923 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][8]/P0001 ,
		_w13784_,
		_w27970_
	);
	LUT2 #(
		.INIT('h1)
	) name23924 (
		_w27967_,
		_w27968_,
		_w27971_
	);
	LUT2 #(
		.INIT('h1)
	) name23925 (
		_w27969_,
		_w27970_,
		_w27972_
	);
	LUT2 #(
		.INIT('h8)
	) name23926 (
		_w27971_,
		_w27972_,
		_w27973_
	);
	LUT2 #(
		.INIT('h2)
	) name23927 (
		_w27921_,
		_w27973_,
		_w27974_
	);
	LUT2 #(
		.INIT('h1)
	) name23928 (
		_w27966_,
		_w27974_,
		_w27975_
	);
	LUT2 #(
		.INIT('h2)
	) name23929 (
		_w27908_,
		_w27975_,
		_w27976_
	);
	LUT2 #(
		.INIT('h2)
	) name23930 (
		_w10638_,
		_w27908_,
		_w27977_
	);
	LUT2 #(
		.INIT('h1)
	) name23931 (
		_w27976_,
		_w27977_,
		_w27978_
	);
	LUT2 #(
		.INIT('h2)
	) name23932 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w27924_,
		_w27979_
	);
	LUT2 #(
		.INIT('h1)
	) name23933 (
		_w27925_,
		_w27979_,
		_w27980_
	);
	LUT2 #(
		.INIT('h1)
	) name23934 (
		_w27921_,
		_w27980_,
		_w27981_
	);
	LUT2 #(
		.INIT('h8)
	) name23935 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][4]/P0001 ,
		_w13794_,
		_w27982_
	);
	LUT2 #(
		.INIT('h8)
	) name23936 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][4]/P0001 ,
		_w13789_,
		_w27983_
	);
	LUT2 #(
		.INIT('h8)
	) name23937 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][4]/P0001 ,
		_w13775_,
		_w27984_
	);
	LUT2 #(
		.INIT('h8)
	) name23938 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][4]/P0001 ,
		_w13784_,
		_w27985_
	);
	LUT2 #(
		.INIT('h1)
	) name23939 (
		_w27982_,
		_w27983_,
		_w27986_
	);
	LUT2 #(
		.INIT('h1)
	) name23940 (
		_w27984_,
		_w27985_,
		_w27987_
	);
	LUT2 #(
		.INIT('h8)
	) name23941 (
		_w27986_,
		_w27987_,
		_w27988_
	);
	LUT2 #(
		.INIT('h2)
	) name23942 (
		_w27921_,
		_w27988_,
		_w27989_
	);
	LUT2 #(
		.INIT('h1)
	) name23943 (
		_w27981_,
		_w27989_,
		_w27990_
	);
	LUT2 #(
		.INIT('h2)
	) name23944 (
		_w27908_,
		_w27990_,
		_w27991_
	);
	LUT2 #(
		.INIT('h2)
	) name23945 (
		_w10069_,
		_w27908_,
		_w27992_
	);
	LUT2 #(
		.INIT('h1)
	) name23946 (
		_w27991_,
		_w27992_,
		_w27993_
	);
	LUT2 #(
		.INIT('h2)
	) name23947 (
		_w9435_,
		_w27908_,
		_w27994_
	);
	LUT2 #(
		.INIT('h8)
	) name23948 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][1]/P0001 ,
		_w13784_,
		_w27995_
	);
	LUT2 #(
		.INIT('h8)
	) name23949 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][1]/P0001 ,
		_w13775_,
		_w27996_
	);
	LUT2 #(
		.INIT('h8)
	) name23950 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][1]/P0001 ,
		_w13794_,
		_w27997_
	);
	LUT2 #(
		.INIT('h8)
	) name23951 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][1]/P0001 ,
		_w13789_,
		_w27998_
	);
	LUT2 #(
		.INIT('h1)
	) name23952 (
		_w27995_,
		_w27996_,
		_w27999_
	);
	LUT2 #(
		.INIT('h1)
	) name23953 (
		_w27997_,
		_w27998_,
		_w28000_
	);
	LUT2 #(
		.INIT('h8)
	) name23954 (
		_w27999_,
		_w28000_,
		_w28001_
	);
	LUT2 #(
		.INIT('h8)
	) name23955 (
		_w27921_,
		_w28001_,
		_w28002_
	);
	LUT2 #(
		.INIT('h8)
	) name23956 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w28003_
	);
	LUT2 #(
		.INIT('h1)
	) name23957 (
		_w27922_,
		_w28003_,
		_w28004_
	);
	LUT2 #(
		.INIT('h4)
	) name23958 (
		_w27921_,
		_w28004_,
		_w28005_
	);
	LUT2 #(
		.INIT('h2)
	) name23959 (
		_w27908_,
		_w28002_,
		_w28006_
	);
	LUT2 #(
		.INIT('h4)
	) name23960 (
		_w28005_,
		_w28006_,
		_w28007_
	);
	LUT2 #(
		.INIT('h1)
	) name23961 (
		_w27994_,
		_w28007_,
		_w28008_
	);
	LUT2 #(
		.INIT('h2)
	) name23962 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w27929_,
		_w28009_
	);
	LUT2 #(
		.INIT('h1)
	) name23963 (
		_w27930_,
		_w28009_,
		_w28010_
	);
	LUT2 #(
		.INIT('h1)
	) name23964 (
		_w27921_,
		_w28010_,
		_w28011_
	);
	LUT2 #(
		.INIT('h8)
	) name23965 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][9]/P0001 ,
		_w13775_,
		_w28012_
	);
	LUT2 #(
		.INIT('h8)
	) name23966 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][9]/P0001 ,
		_w13794_,
		_w28013_
	);
	LUT2 #(
		.INIT('h8)
	) name23967 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][9]/P0001 ,
		_w13789_,
		_w28014_
	);
	LUT2 #(
		.INIT('h8)
	) name23968 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][9]/P0001 ,
		_w13784_,
		_w28015_
	);
	LUT2 #(
		.INIT('h1)
	) name23969 (
		_w28012_,
		_w28013_,
		_w28016_
	);
	LUT2 #(
		.INIT('h1)
	) name23970 (
		_w28014_,
		_w28015_,
		_w28017_
	);
	LUT2 #(
		.INIT('h8)
	) name23971 (
		_w28016_,
		_w28017_,
		_w28018_
	);
	LUT2 #(
		.INIT('h2)
	) name23972 (
		_w27921_,
		_w28018_,
		_w28019_
	);
	LUT2 #(
		.INIT('h1)
	) name23973 (
		_w28011_,
		_w28019_,
		_w28020_
	);
	LUT2 #(
		.INIT('h2)
	) name23974 (
		_w27908_,
		_w28020_,
		_w28021_
	);
	LUT2 #(
		.INIT('h2)
	) name23975 (
		_w10289_,
		_w27908_,
		_w28022_
	);
	LUT2 #(
		.INIT('h1)
	) name23976 (
		_w28021_,
		_w28022_,
		_w28023_
	);
	LUT2 #(
		.INIT('h2)
	) name23977 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w27923_,
		_w28024_
	);
	LUT2 #(
		.INIT('h1)
	) name23978 (
		_w27924_,
		_w28024_,
		_w28025_
	);
	LUT2 #(
		.INIT('h1)
	) name23979 (
		_w27921_,
		_w28025_,
		_w28026_
	);
	LUT2 #(
		.INIT('h8)
	) name23980 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][3]/P0001 ,
		_w13794_,
		_w28027_
	);
	LUT2 #(
		.INIT('h8)
	) name23981 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][3]/P0001 ,
		_w13789_,
		_w28028_
	);
	LUT2 #(
		.INIT('h8)
	) name23982 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][3]/P0001 ,
		_w13775_,
		_w28029_
	);
	LUT2 #(
		.INIT('h8)
	) name23983 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][3]/P0001 ,
		_w13784_,
		_w28030_
	);
	LUT2 #(
		.INIT('h1)
	) name23984 (
		_w28027_,
		_w28028_,
		_w28031_
	);
	LUT2 #(
		.INIT('h1)
	) name23985 (
		_w28029_,
		_w28030_,
		_w28032_
	);
	LUT2 #(
		.INIT('h8)
	) name23986 (
		_w28031_,
		_w28032_,
		_w28033_
	);
	LUT2 #(
		.INIT('h2)
	) name23987 (
		_w27921_,
		_w28033_,
		_w28034_
	);
	LUT2 #(
		.INIT('h1)
	) name23988 (
		_w28026_,
		_w28034_,
		_w28035_
	);
	LUT2 #(
		.INIT('h2)
	) name23989 (
		_w27908_,
		_w28035_,
		_w28036_
	);
	LUT2 #(
		.INIT('h2)
	) name23990 (
		_w8113_,
		_w27908_,
		_w28037_
	);
	LUT2 #(
		.INIT('h1)
	) name23991 (
		_w28036_,
		_w28037_,
		_w28038_
	);
	LUT2 #(
		.INIT('h2)
	) name23992 (
		_w7340_,
		_w27908_,
		_w28039_
	);
	LUT2 #(
		.INIT('h2)
	) name23993 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w27933_,
		_w28040_
	);
	LUT2 #(
		.INIT('h4)
	) name23994 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w27933_,
		_w28041_
	);
	LUT2 #(
		.INIT('h1)
	) name23995 (
		_w28040_,
		_w28041_,
		_w28042_
	);
	LUT2 #(
		.INIT('h4)
	) name23996 (
		_w27921_,
		_w28042_,
		_w28043_
	);
	LUT2 #(
		.INIT('h8)
	) name23997 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][13]/P0001 ,
		_w13784_,
		_w28044_
	);
	LUT2 #(
		.INIT('h8)
	) name23998 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][13]/P0001 ,
		_w13775_,
		_w28045_
	);
	LUT2 #(
		.INIT('h8)
	) name23999 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][13]/P0001 ,
		_w13794_,
		_w28046_
	);
	LUT2 #(
		.INIT('h8)
	) name24000 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][13]/P0001 ,
		_w13789_,
		_w28047_
	);
	LUT2 #(
		.INIT('h1)
	) name24001 (
		_w28044_,
		_w28045_,
		_w28048_
	);
	LUT2 #(
		.INIT('h1)
	) name24002 (
		_w28046_,
		_w28047_,
		_w28049_
	);
	LUT2 #(
		.INIT('h8)
	) name24003 (
		_w28048_,
		_w28049_,
		_w28050_
	);
	LUT2 #(
		.INIT('h8)
	) name24004 (
		_w27921_,
		_w28050_,
		_w28051_
	);
	LUT2 #(
		.INIT('h2)
	) name24005 (
		_w27908_,
		_w28043_,
		_w28052_
	);
	LUT2 #(
		.INIT('h4)
	) name24006 (
		_w28051_,
		_w28052_,
		_w28053_
	);
	LUT2 #(
		.INIT('h1)
	) name24007 (
		_w28039_,
		_w28053_,
		_w28054_
	);
	LUT2 #(
		.INIT('h2)
	) name24008 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w27922_,
		_w28055_
	);
	LUT2 #(
		.INIT('h1)
	) name24009 (
		_w27923_,
		_w28055_,
		_w28056_
	);
	LUT2 #(
		.INIT('h1)
	) name24010 (
		_w27921_,
		_w28056_,
		_w28057_
	);
	LUT2 #(
		.INIT('h8)
	) name24011 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][2]/P0001 ,
		_w13794_,
		_w28058_
	);
	LUT2 #(
		.INIT('h8)
	) name24012 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][2]/P0001 ,
		_w13789_,
		_w28059_
	);
	LUT2 #(
		.INIT('h8)
	) name24013 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][2]/P0001 ,
		_w13775_,
		_w28060_
	);
	LUT2 #(
		.INIT('h8)
	) name24014 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][2]/P0001 ,
		_w13784_,
		_w28061_
	);
	LUT2 #(
		.INIT('h1)
	) name24015 (
		_w28058_,
		_w28059_,
		_w28062_
	);
	LUT2 #(
		.INIT('h1)
	) name24016 (
		_w28060_,
		_w28061_,
		_w28063_
	);
	LUT2 #(
		.INIT('h8)
	) name24017 (
		_w28062_,
		_w28063_,
		_w28064_
	);
	LUT2 #(
		.INIT('h2)
	) name24018 (
		_w27921_,
		_w28064_,
		_w28065_
	);
	LUT2 #(
		.INIT('h1)
	) name24019 (
		_w28057_,
		_w28065_,
		_w28066_
	);
	LUT2 #(
		.INIT('h2)
	) name24020 (
		_w27908_,
		_w28066_,
		_w28067_
	);
	LUT2 #(
		.INIT('h2)
	) name24021 (
		_w8715_,
		_w27908_,
		_w28068_
	);
	LUT2 #(
		.INIT('h1)
	) name24022 (
		_w28067_,
		_w28068_,
		_w28069_
	);
	LUT2 #(
		.INIT('h1)
	) name24023 (
		_w7607_,
		_w27908_,
		_w28070_
	);
	LUT2 #(
		.INIT('h1)
	) name24024 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		_w27921_,
		_w28071_
	);
	LUT2 #(
		.INIT('h8)
	) name24025 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][0]/P0001 ,
		_w13784_,
		_w28072_
	);
	LUT2 #(
		.INIT('h8)
	) name24026 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][0]/P0001 ,
		_w13794_,
		_w28073_
	);
	LUT2 #(
		.INIT('h8)
	) name24027 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][0]/P0001 ,
		_w13789_,
		_w28074_
	);
	LUT2 #(
		.INIT('h8)
	) name24028 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][0]/P0001 ,
		_w13775_,
		_w28075_
	);
	LUT2 #(
		.INIT('h1)
	) name24029 (
		_w28072_,
		_w28073_,
		_w28076_
	);
	LUT2 #(
		.INIT('h1)
	) name24030 (
		_w28074_,
		_w28075_,
		_w28077_
	);
	LUT2 #(
		.INIT('h8)
	) name24031 (
		_w28076_,
		_w28077_,
		_w28078_
	);
	LUT2 #(
		.INIT('h2)
	) name24032 (
		_w27921_,
		_w28078_,
		_w28079_
	);
	LUT2 #(
		.INIT('h2)
	) name24033 (
		_w27908_,
		_w28071_,
		_w28080_
	);
	LUT2 #(
		.INIT('h4)
	) name24034 (
		_w28079_,
		_w28080_,
		_w28081_
	);
	LUT2 #(
		.INIT('h2)
	) name24035 (
		_w27915_,
		_w28070_,
		_w28082_
	);
	LUT2 #(
		.INIT('h4)
	) name24036 (
		_w28081_,
		_w28082_,
		_w28083_
	);
	LUT2 #(
		.INIT('h2)
	) name24037 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w27927_,
		_w28084_
	);
	LUT2 #(
		.INIT('h1)
	) name24038 (
		_w27928_,
		_w28084_,
		_w28085_
	);
	LUT2 #(
		.INIT('h1)
	) name24039 (
		_w27921_,
		_w28085_,
		_w28086_
	);
	LUT2 #(
		.INIT('h8)
	) name24040 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][7]/P0001 ,
		_w13794_,
		_w28087_
	);
	LUT2 #(
		.INIT('h8)
	) name24041 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][7]/P0001 ,
		_w13789_,
		_w28088_
	);
	LUT2 #(
		.INIT('h8)
	) name24042 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][7]/P0001 ,
		_w13784_,
		_w28089_
	);
	LUT2 #(
		.INIT('h8)
	) name24043 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][7]/P0001 ,
		_w13775_,
		_w28090_
	);
	LUT2 #(
		.INIT('h1)
	) name24044 (
		_w28087_,
		_w28088_,
		_w28091_
	);
	LUT2 #(
		.INIT('h1)
	) name24045 (
		_w28089_,
		_w28090_,
		_w28092_
	);
	LUT2 #(
		.INIT('h8)
	) name24046 (
		_w28091_,
		_w28092_,
		_w28093_
	);
	LUT2 #(
		.INIT('h2)
	) name24047 (
		_w27921_,
		_w28093_,
		_w28094_
	);
	LUT2 #(
		.INIT('h1)
	) name24048 (
		_w28086_,
		_w28094_,
		_w28095_
	);
	LUT2 #(
		.INIT('h2)
	) name24049 (
		_w27908_,
		_w28095_,
		_w28096_
	);
	LUT2 #(
		.INIT('h2)
	) name24050 (
		_w11265_,
		_w27908_,
		_w28097_
	);
	LUT2 #(
		.INIT('h1)
	) name24051 (
		_w28096_,
		_w28097_,
		_w28098_
	);
	LUT2 #(
		.INIT('h2)
	) name24052 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w27926_,
		_w28099_
	);
	LUT2 #(
		.INIT('h1)
	) name24053 (
		_w27927_,
		_w28099_,
		_w28100_
	);
	LUT2 #(
		.INIT('h1)
	) name24054 (
		_w27921_,
		_w28100_,
		_w28101_
	);
	LUT2 #(
		.INIT('h8)
	) name24055 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][6]/P0001 ,
		_w13775_,
		_w28102_
	);
	LUT2 #(
		.INIT('h8)
	) name24056 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][6]/P0001 ,
		_w13784_,
		_w28103_
	);
	LUT2 #(
		.INIT('h8)
	) name24057 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][6]/P0001 ,
		_w13789_,
		_w28104_
	);
	LUT2 #(
		.INIT('h8)
	) name24058 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][6]/P0001 ,
		_w13794_,
		_w28105_
	);
	LUT2 #(
		.INIT('h1)
	) name24059 (
		_w28102_,
		_w28103_,
		_w28106_
	);
	LUT2 #(
		.INIT('h1)
	) name24060 (
		_w28104_,
		_w28105_,
		_w28107_
	);
	LUT2 #(
		.INIT('h8)
	) name24061 (
		_w28106_,
		_w28107_,
		_w28108_
	);
	LUT2 #(
		.INIT('h2)
	) name24062 (
		_w27921_,
		_w28108_,
		_w28109_
	);
	LUT2 #(
		.INIT('h1)
	) name24063 (
		_w28101_,
		_w28109_,
		_w28110_
	);
	LUT2 #(
		.INIT('h2)
	) name24064 (
		_w27908_,
		_w28110_,
		_w28111_
	);
	LUT2 #(
		.INIT('h2)
	) name24065 (
		_w11525_,
		_w27908_,
		_w28112_
	);
	LUT2 #(
		.INIT('h1)
	) name24066 (
		_w28111_,
		_w28112_,
		_w28113_
	);
	LUT2 #(
		.INIT('h2)
	) name24067 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w27925_,
		_w28114_
	);
	LUT2 #(
		.INIT('h1)
	) name24068 (
		_w27926_,
		_w28114_,
		_w28115_
	);
	LUT2 #(
		.INIT('h1)
	) name24069 (
		_w27921_,
		_w28115_,
		_w28116_
	);
	LUT2 #(
		.INIT('h8)
	) name24070 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001 ,
		_w13775_,
		_w28117_
	);
	LUT2 #(
		.INIT('h8)
	) name24071 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001 ,
		_w13784_,
		_w28118_
	);
	LUT2 #(
		.INIT('h8)
	) name24072 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001 ,
		_w13794_,
		_w28119_
	);
	LUT2 #(
		.INIT('h8)
	) name24073 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001 ,
		_w13789_,
		_w28120_
	);
	LUT2 #(
		.INIT('h1)
	) name24074 (
		_w28117_,
		_w28118_,
		_w28121_
	);
	LUT2 #(
		.INIT('h1)
	) name24075 (
		_w28119_,
		_w28120_,
		_w28122_
	);
	LUT2 #(
		.INIT('h8)
	) name24076 (
		_w28121_,
		_w28122_,
		_w28123_
	);
	LUT2 #(
		.INIT('h2)
	) name24077 (
		_w27921_,
		_w28123_,
		_w28124_
	);
	LUT2 #(
		.INIT('h1)
	) name24078 (
		_w28116_,
		_w28124_,
		_w28125_
	);
	LUT2 #(
		.INIT('h2)
	) name24079 (
		_w27908_,
		_w28125_,
		_w28126_
	);
	LUT2 #(
		.INIT('h2)
	) name24080 (
		_w10911_,
		_w27908_,
		_w28127_
	);
	LUT2 #(
		.INIT('h1)
	) name24081 (
		_w28126_,
		_w28127_,
		_w28128_
	);
	LUT2 #(
		.INIT('h2)
	) name24082 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w27931_,
		_w28129_
	);
	LUT2 #(
		.INIT('h1)
	) name24083 (
		_w27932_,
		_w28129_,
		_w28130_
	);
	LUT2 #(
		.INIT('h1)
	) name24084 (
		_w27921_,
		_w28130_,
		_w28131_
	);
	LUT2 #(
		.INIT('h8)
	) name24085 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][11]/P0001 ,
		_w13775_,
		_w28132_
	);
	LUT2 #(
		.INIT('h8)
	) name24086 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][11]/P0001 ,
		_w13784_,
		_w28133_
	);
	LUT2 #(
		.INIT('h8)
	) name24087 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][11]/P0001 ,
		_w13789_,
		_w28134_
	);
	LUT2 #(
		.INIT('h8)
	) name24088 (
		\core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][11]/P0001 ,
		_w13794_,
		_w28135_
	);
	LUT2 #(
		.INIT('h1)
	) name24089 (
		_w28132_,
		_w28133_,
		_w28136_
	);
	LUT2 #(
		.INIT('h1)
	) name24090 (
		_w28134_,
		_w28135_,
		_w28137_
	);
	LUT2 #(
		.INIT('h8)
	) name24091 (
		_w28136_,
		_w28137_,
		_w28138_
	);
	LUT2 #(
		.INIT('h2)
	) name24092 (
		_w27921_,
		_w28138_,
		_w28139_
	);
	LUT2 #(
		.INIT('h1)
	) name24093 (
		_w28131_,
		_w28139_,
		_w28140_
	);
	LUT2 #(
		.INIT('h2)
	) name24094 (
		_w27908_,
		_w28140_,
		_w28141_
	);
	LUT2 #(
		.INIT('h2)
	) name24095 (
		_w8460_,
		_w27908_,
		_w28142_
	);
	LUT2 #(
		.INIT('h1)
	) name24096 (
		_w28141_,
		_w28142_,
		_w28143_
	);
	LUT2 #(
		.INIT('h8)
	) name24097 (
		_w27948_,
		_w27963_,
		_w28144_
	);
	LUT2 #(
		.INIT('h8)
	) name24098 (
		_w27978_,
		_w27993_,
		_w28145_
	);
	LUT2 #(
		.INIT('h8)
	) name24099 (
		_w28008_,
		_w28023_,
		_w28146_
	);
	LUT2 #(
		.INIT('h8)
	) name24100 (
		_w28038_,
		_w28054_,
		_w28147_
	);
	LUT2 #(
		.INIT('h8)
	) name24101 (
		_w28069_,
		_w28083_,
		_w28148_
	);
	LUT2 #(
		.INIT('h8)
	) name24102 (
		_w28098_,
		_w28113_,
		_w28149_
	);
	LUT2 #(
		.INIT('h8)
	) name24103 (
		_w28128_,
		_w28143_,
		_w28150_
	);
	LUT2 #(
		.INIT('h8)
	) name24104 (
		_w28149_,
		_w28150_,
		_w28151_
	);
	LUT2 #(
		.INIT('h8)
	) name24105 (
		_w28147_,
		_w28148_,
		_w28152_
	);
	LUT2 #(
		.INIT('h8)
	) name24106 (
		_w28145_,
		_w28146_,
		_w28153_
	);
	LUT2 #(
		.INIT('h8)
	) name24107 (
		_w28144_,
		_w28153_,
		_w28154_
	);
	LUT2 #(
		.INIT('h8)
	) name24108 (
		_w28151_,
		_w28152_,
		_w28155_
	);
	LUT2 #(
		.INIT('h8)
	) name24109 (
		_w28154_,
		_w28155_,
		_w28156_
	);
	LUT2 #(
		.INIT('h1)
	) name24110 (
		_w27916_,
		_w28156_,
		_w28157_
	);
	LUT2 #(
		.INIT('h4)
	) name24111 (
		_w27103_,
		_w27499_,
		_w28158_
	);
	LUT2 #(
		.INIT('h1)
	) name24112 (
		_w27500_,
		_w28158_,
		_w28159_
	);
	LUT2 #(
		.INIT('h2)
	) name24113 (
		\idma_PM_1st_reg/NET0131 ,
		_w20394_,
		_w28160_
	);
	LUT2 #(
		.INIT('h1)
	) name24114 (
		\idma_PM_1st_reg/NET0131 ,
		_w20388_,
		_w28161_
	);
	LUT2 #(
		.INIT('h2)
	) name24115 (
		_w20822_,
		_w28161_,
		_w28162_
	);
	LUT2 #(
		.INIT('h4)
	) name24116 (
		_w28160_,
		_w28162_,
		_w28163_
	);
	LUT2 #(
		.INIT('h4)
	) name24117 (
		_w13570_,
		_w28163_,
		_w28164_
	);
	LUT2 #(
		.INIT('h4)
	) name24118 (
		_w28159_,
		_w28164_,
		_w28165_
	);
	LUT2 #(
		.INIT('h2)
	) name24119 (
		\idma_DTMP_L_reg[7]/P0001 ,
		_w28163_,
		_w28166_
	);
	LUT2 #(
		.INIT('h1)
	) name24120 (
		_w28165_,
		_w28166_,
		_w28167_
	);
	LUT2 #(
		.INIT('h4)
	) name24121 (
		_w27187_,
		_w27499_,
		_w28168_
	);
	LUT2 #(
		.INIT('h1)
	) name24122 (
		_w27527_,
		_w28168_,
		_w28169_
	);
	LUT2 #(
		.INIT('h2)
	) name24123 (
		_w28164_,
		_w28169_,
		_w28170_
	);
	LUT2 #(
		.INIT('h2)
	) name24124 (
		\idma_DTMP_L_reg[4]/P0001 ,
		_w28163_,
		_w28171_
	);
	LUT2 #(
		.INIT('h1)
	) name24125 (
		_w28170_,
		_w28171_,
		_w28172_
	);
	LUT2 #(
		.INIT('h4)
	) name24126 (
		_w27215_,
		_w27499_,
		_w28173_
	);
	LUT2 #(
		.INIT('h1)
	) name24127 (
		_w27536_,
		_w28173_,
		_w28174_
	);
	LUT2 #(
		.INIT('h2)
	) name24128 (
		_w28164_,
		_w28174_,
		_w28175_
	);
	LUT2 #(
		.INIT('h2)
	) name24129 (
		\idma_DTMP_L_reg[3]/P0001 ,
		_w28163_,
		_w28176_
	);
	LUT2 #(
		.INIT('h1)
	) name24130 (
		_w28175_,
		_w28176_,
		_w28177_
	);
	LUT2 #(
		.INIT('h4)
	) name24131 (
		_w27131_,
		_w27499_,
		_w28178_
	);
	LUT2 #(
		.INIT('h1)
	) name24132 (
		_w27509_,
		_w28178_,
		_w28179_
	);
	LUT2 #(
		.INIT('h2)
	) name24133 (
		_w28164_,
		_w28179_,
		_w28180_
	);
	LUT2 #(
		.INIT('h2)
	) name24134 (
		\idma_DTMP_L_reg[6]/P0001 ,
		_w28163_,
		_w28181_
	);
	LUT2 #(
		.INIT('h1)
	) name24135 (
		_w28180_,
		_w28181_,
		_w28182_
	);
	LUT2 #(
		.INIT('h4)
	) name24136 (
		_w27243_,
		_w27499_,
		_w28183_
	);
	LUT2 #(
		.INIT('h1)
	) name24137 (
		_w27545_,
		_w28183_,
		_w28184_
	);
	LUT2 #(
		.INIT('h2)
	) name24138 (
		_w28164_,
		_w28184_,
		_w28185_
	);
	LUT2 #(
		.INIT('h2)
	) name24139 (
		\idma_DTMP_L_reg[2]/P0001 ,
		_w28163_,
		_w28186_
	);
	LUT2 #(
		.INIT('h1)
	) name24140 (
		_w28185_,
		_w28186_,
		_w28187_
	);
	LUT2 #(
		.INIT('h4)
	) name24141 (
		_w27159_,
		_w27499_,
		_w28188_
	);
	LUT2 #(
		.INIT('h1)
	) name24142 (
		_w27518_,
		_w28188_,
		_w28189_
	);
	LUT2 #(
		.INIT('h2)
	) name24143 (
		_w28164_,
		_w28189_,
		_w28190_
	);
	LUT2 #(
		.INIT('h2)
	) name24144 (
		\idma_DTMP_L_reg[5]/P0001 ,
		_w28163_,
		_w28191_
	);
	LUT2 #(
		.INIT('h1)
	) name24145 (
		_w28190_,
		_w28191_,
		_w28192_
	);
	LUT2 #(
		.INIT('h4)
	) name24146 (
		_w27271_,
		_w27499_,
		_w28193_
	);
	LUT2 #(
		.INIT('h1)
	) name24147 (
		_w27554_,
		_w28193_,
		_w28194_
	);
	LUT2 #(
		.INIT('h2)
	) name24148 (
		_w28164_,
		_w28194_,
		_w28195_
	);
	LUT2 #(
		.INIT('h2)
	) name24149 (
		\idma_DTMP_L_reg[1]/P0001 ,
		_w28163_,
		_w28196_
	);
	LUT2 #(
		.INIT('h1)
	) name24150 (
		_w28195_,
		_w28196_,
		_w28197_
	);
	LUT2 #(
		.INIT('h4)
	) name24151 (
		_w27299_,
		_w27499_,
		_w28198_
	);
	LUT2 #(
		.INIT('h1)
	) name24152 (
		_w27615_,
		_w28198_,
		_w28199_
	);
	LUT2 #(
		.INIT('h2)
	) name24153 (
		_w28164_,
		_w28199_,
		_w28200_
	);
	LUT2 #(
		.INIT('h2)
	) name24154 (
		\idma_DTMP_L_reg[0]/P0001 ,
		_w28163_,
		_w28201_
	);
	LUT2 #(
		.INIT('h1)
	) name24155 (
		_w28200_,
		_w28201_,
		_w28202_
	);
	LUT2 #(
		.INIT('h8)
	) name24156 (
		_w23027_,
		_w25033_,
		_w28203_
	);
	LUT2 #(
		.INIT('h8)
	) name24157 (
		_w26967_,
		_w28203_,
		_w28204_
	);
	LUT2 #(
		.INIT('h1)
	) name24158 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w28204_,
		_w28205_
	);
	LUT2 #(
		.INIT('h4)
	) name24159 (
		\sice_SPC_reg[9]/P0001 ,
		_w28204_,
		_w28206_
	);
	LUT2 #(
		.INIT('h1)
	) name24160 (
		_w28205_,
		_w28206_,
		_w28207_
	);
	LUT2 #(
		.INIT('h2)
	) name24161 (
		_w21242_,
		_w28207_,
		_w28208_
	);
	LUT2 #(
		.INIT('h4)
	) name24162 (
		_w21242_,
		_w27419_,
		_w28209_
	);
	LUT2 #(
		.INIT('h1)
	) name24163 (
		_w28208_,
		_w28209_,
		_w28210_
	);
	LUT2 #(
		.INIT('h1)
	) name24164 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w28204_,
		_w28211_
	);
	LUT2 #(
		.INIT('h4)
	) name24165 (
		\sice_SPC_reg[8]/P0001 ,
		_w28204_,
		_w28212_
	);
	LUT2 #(
		.INIT('h1)
	) name24166 (
		_w28211_,
		_w28212_,
		_w28213_
	);
	LUT2 #(
		.INIT('h2)
	) name24167 (
		_w21242_,
		_w28213_,
		_w28214_
	);
	LUT2 #(
		.INIT('h4)
	) name24168 (
		_w21242_,
		_w27391_,
		_w28215_
	);
	LUT2 #(
		.INIT('h1)
	) name24169 (
		_w28214_,
		_w28215_,
		_w28216_
	);
	LUT2 #(
		.INIT('h1)
	) name24170 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w28204_,
		_w28217_
	);
	LUT2 #(
		.INIT('h4)
	) name24171 (
		\sice_SPC_reg[7]/P0001 ,
		_w28204_,
		_w28218_
	);
	LUT2 #(
		.INIT('h1)
	) name24172 (
		_w28217_,
		_w28218_,
		_w28219_
	);
	LUT2 #(
		.INIT('h2)
	) name24173 (
		_w21242_,
		_w28219_,
		_w28220_
	);
	LUT2 #(
		.INIT('h4)
	) name24174 (
		_w21242_,
		_w27105_,
		_w28221_
	);
	LUT2 #(
		.INIT('h1)
	) name24175 (
		_w28220_,
		_w28221_,
		_w28222_
	);
	LUT2 #(
		.INIT('h1)
	) name24176 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w28204_,
		_w28223_
	);
	LUT2 #(
		.INIT('h4)
	) name24177 (
		\sice_SPC_reg[6]/P0001 ,
		_w28204_,
		_w28224_
	);
	LUT2 #(
		.INIT('h1)
	) name24178 (
		_w28223_,
		_w28224_,
		_w28225_
	);
	LUT2 #(
		.INIT('h2)
	) name24179 (
		_w21242_,
		_w28225_,
		_w28226_
	);
	LUT2 #(
		.INIT('h4)
	) name24180 (
		_w21242_,
		_w27133_,
		_w28227_
	);
	LUT2 #(
		.INIT('h1)
	) name24181 (
		_w28226_,
		_w28227_,
		_w28228_
	);
	LUT2 #(
		.INIT('h1)
	) name24182 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w28204_,
		_w28229_
	);
	LUT2 #(
		.INIT('h4)
	) name24183 (
		\sice_SPC_reg[5]/P0001 ,
		_w28204_,
		_w28230_
	);
	LUT2 #(
		.INIT('h1)
	) name24184 (
		_w28229_,
		_w28230_,
		_w28231_
	);
	LUT2 #(
		.INIT('h2)
	) name24185 (
		_w21242_,
		_w28231_,
		_w28232_
	);
	LUT2 #(
		.INIT('h4)
	) name24186 (
		_w21242_,
		_w27161_,
		_w28233_
	);
	LUT2 #(
		.INIT('h1)
	) name24187 (
		_w28232_,
		_w28233_,
		_w28234_
	);
	LUT2 #(
		.INIT('h1)
	) name24188 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w28204_,
		_w28235_
	);
	LUT2 #(
		.INIT('h4)
	) name24189 (
		\sice_SPC_reg[4]/P0001 ,
		_w28204_,
		_w28236_
	);
	LUT2 #(
		.INIT('h1)
	) name24190 (
		_w28235_,
		_w28236_,
		_w28237_
	);
	LUT2 #(
		.INIT('h2)
	) name24191 (
		_w21242_,
		_w28237_,
		_w28238_
	);
	LUT2 #(
		.INIT('h4)
	) name24192 (
		_w21242_,
		_w27189_,
		_w28239_
	);
	LUT2 #(
		.INIT('h1)
	) name24193 (
		_w28238_,
		_w28239_,
		_w28240_
	);
	LUT2 #(
		.INIT('h1)
	) name24194 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w28204_,
		_w28241_
	);
	LUT2 #(
		.INIT('h4)
	) name24195 (
		\sice_SPC_reg[3]/P0001 ,
		_w28204_,
		_w28242_
	);
	LUT2 #(
		.INIT('h1)
	) name24196 (
		_w28241_,
		_w28242_,
		_w28243_
	);
	LUT2 #(
		.INIT('h2)
	) name24197 (
		_w21242_,
		_w28243_,
		_w28244_
	);
	LUT2 #(
		.INIT('h4)
	) name24198 (
		_w21242_,
		_w27217_,
		_w28245_
	);
	LUT2 #(
		.INIT('h1)
	) name24199 (
		_w28244_,
		_w28245_,
		_w28246_
	);
	LUT2 #(
		.INIT('h1)
	) name24200 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w28204_,
		_w28247_
	);
	LUT2 #(
		.INIT('h4)
	) name24201 (
		\sice_SPC_reg[2]/P0001 ,
		_w28204_,
		_w28248_
	);
	LUT2 #(
		.INIT('h1)
	) name24202 (
		_w28247_,
		_w28248_,
		_w28249_
	);
	LUT2 #(
		.INIT('h2)
	) name24203 (
		_w21242_,
		_w28249_,
		_w28250_
	);
	LUT2 #(
		.INIT('h4)
	) name24204 (
		_w21242_,
		_w27245_,
		_w28251_
	);
	LUT2 #(
		.INIT('h1)
	) name24205 (
		_w28250_,
		_w28251_,
		_w28252_
	);
	LUT2 #(
		.INIT('h1)
	) name24206 (
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w28204_,
		_w28253_
	);
	LUT2 #(
		.INIT('h4)
	) name24207 (
		\sice_SPC_reg[23]/P0001 ,
		_w28204_,
		_w28254_
	);
	LUT2 #(
		.INIT('h1)
	) name24208 (
		_w28253_,
		_w28254_,
		_w28255_
	);
	LUT2 #(
		.INIT('h2)
	) name24209 (
		_w21242_,
		_w28255_,
		_w28256_
	);
	LUT2 #(
		.INIT('h8)
	) name24210 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[23]/P0001 ,
		_w28257_
	);
	LUT2 #(
		.INIT('h1)
	) name24211 (
		\T_TMODE[1]_pad ,
		_w27577_,
		_w28258_
	);
	LUT2 #(
		.INIT('h1)
	) name24212 (
		_w28257_,
		_w28258_,
		_w28259_
	);
	LUT2 #(
		.INIT('h4)
	) name24213 (
		_w21242_,
		_w28259_,
		_w28260_
	);
	LUT2 #(
		.INIT('h1)
	) name24214 (
		_w28256_,
		_w28260_,
		_w28261_
	);
	LUT2 #(
		.INIT('h1)
	) name24215 (
		\core_c_dec_IR_reg[22]/NET0131 ,
		_w28204_,
		_w28262_
	);
	LUT2 #(
		.INIT('h4)
	) name24216 (
		\sice_SPC_reg[22]/P0001 ,
		_w28204_,
		_w28263_
	);
	LUT2 #(
		.INIT('h1)
	) name24217 (
		_w28262_,
		_w28263_,
		_w28264_
	);
	LUT2 #(
		.INIT('h2)
	) name24218 (
		_w21242_,
		_w28264_,
		_w28265_
	);
	LUT2 #(
		.INIT('h8)
	) name24219 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[22]/P0001 ,
		_w28266_
	);
	LUT2 #(
		.INIT('h1)
	) name24220 (
		\T_TMODE[1]_pad ,
		_w27603_,
		_w28267_
	);
	LUT2 #(
		.INIT('h1)
	) name24221 (
		_w28266_,
		_w28267_,
		_w28268_
	);
	LUT2 #(
		.INIT('h4)
	) name24222 (
		_w21242_,
		_w28268_,
		_w28269_
	);
	LUT2 #(
		.INIT('h1)
	) name24223 (
		_w28265_,
		_w28269_,
		_w28270_
	);
	LUT2 #(
		.INIT('h1)
	) name24224 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		_w28204_,
		_w28271_
	);
	LUT2 #(
		.INIT('h4)
	) name24225 (
		\sice_SPC_reg[21]/P0001 ,
		_w28204_,
		_w28272_
	);
	LUT2 #(
		.INIT('h1)
	) name24226 (
		_w28271_,
		_w28272_,
		_w28273_
	);
	LUT2 #(
		.INIT('h2)
	) name24227 (
		_w21242_,
		_w28273_,
		_w28274_
	);
	LUT2 #(
		.INIT('h8)
	) name24228 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[21]/P0001 ,
		_w28275_
	);
	LUT2 #(
		.INIT('h1)
	) name24229 (
		\T_TMODE[1]_pad ,
		_w27695_,
		_w28276_
	);
	LUT2 #(
		.INIT('h1)
	) name24230 (
		_w28275_,
		_w28276_,
		_w28277_
	);
	LUT2 #(
		.INIT('h4)
	) name24231 (
		_w21242_,
		_w28277_,
		_w28278_
	);
	LUT2 #(
		.INIT('h1)
	) name24232 (
		_w28274_,
		_w28278_,
		_w28279_
	);
	LUT2 #(
		.INIT('h1)
	) name24233 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w28204_,
		_w28280_
	);
	LUT2 #(
		.INIT('h4)
	) name24234 (
		\sice_SPC_reg[20]/P0001 ,
		_w28204_,
		_w28281_
	);
	LUT2 #(
		.INIT('h1)
	) name24235 (
		_w28280_,
		_w28281_,
		_w28282_
	);
	LUT2 #(
		.INIT('h2)
	) name24236 (
		_w21242_,
		_w28282_,
		_w28283_
	);
	LUT2 #(
		.INIT('h8)
	) name24237 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[20]/P0001 ,
		_w28284_
	);
	LUT2 #(
		.INIT('h1)
	) name24238 (
		\T_TMODE[1]_pad ,
		_w27721_,
		_w28285_
	);
	LUT2 #(
		.INIT('h1)
	) name24239 (
		_w28284_,
		_w28285_,
		_w28286_
	);
	LUT2 #(
		.INIT('h4)
	) name24240 (
		_w21242_,
		_w28286_,
		_w28287_
	);
	LUT2 #(
		.INIT('h1)
	) name24241 (
		_w28283_,
		_w28287_,
		_w28288_
	);
	LUT2 #(
		.INIT('h1)
	) name24242 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w28204_,
		_w28289_
	);
	LUT2 #(
		.INIT('h4)
	) name24243 (
		\sice_SPC_reg[19]/P0001 ,
		_w28204_,
		_w28290_
	);
	LUT2 #(
		.INIT('h1)
	) name24244 (
		_w28289_,
		_w28290_,
		_w28291_
	);
	LUT2 #(
		.INIT('h2)
	) name24245 (
		_w21242_,
		_w28291_,
		_w28292_
	);
	LUT2 #(
		.INIT('h8)
	) name24246 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[19]/P0001 ,
		_w28293_
	);
	LUT2 #(
		.INIT('h1)
	) name24247 (
		\T_TMODE[1]_pad ,
		_w27747_,
		_w28294_
	);
	LUT2 #(
		.INIT('h1)
	) name24248 (
		_w28293_,
		_w28294_,
		_w28295_
	);
	LUT2 #(
		.INIT('h4)
	) name24249 (
		_w21242_,
		_w28295_,
		_w28296_
	);
	LUT2 #(
		.INIT('h1)
	) name24250 (
		_w28292_,
		_w28296_,
		_w28297_
	);
	LUT2 #(
		.INIT('h1)
	) name24251 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		_w28204_,
		_w28298_
	);
	LUT2 #(
		.INIT('h4)
	) name24252 (
		\sice_SPC_reg[18]/P0001 ,
		_w28204_,
		_w28299_
	);
	LUT2 #(
		.INIT('h1)
	) name24253 (
		_w28298_,
		_w28299_,
		_w28300_
	);
	LUT2 #(
		.INIT('h2)
	) name24254 (
		_w21242_,
		_w28300_,
		_w28301_
	);
	LUT2 #(
		.INIT('h8)
	) name24255 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[18]/P0001 ,
		_w28302_
	);
	LUT2 #(
		.INIT('h1)
	) name24256 (
		\T_TMODE[1]_pad ,
		_w27773_,
		_w28303_
	);
	LUT2 #(
		.INIT('h1)
	) name24257 (
		_w28302_,
		_w28303_,
		_w28304_
	);
	LUT2 #(
		.INIT('h4)
	) name24258 (
		_w21242_,
		_w28304_,
		_w28305_
	);
	LUT2 #(
		.INIT('h1)
	) name24259 (
		_w28301_,
		_w28305_,
		_w28306_
	);
	LUT2 #(
		.INIT('h1)
	) name24260 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w28204_,
		_w28307_
	);
	LUT2 #(
		.INIT('h4)
	) name24261 (
		\sice_SPC_reg[17]/P0001 ,
		_w28204_,
		_w28308_
	);
	LUT2 #(
		.INIT('h1)
	) name24262 (
		_w28307_,
		_w28308_,
		_w28309_
	);
	LUT2 #(
		.INIT('h2)
	) name24263 (
		_w21242_,
		_w28309_,
		_w28310_
	);
	LUT2 #(
		.INIT('h8)
	) name24264 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[17]/P0001 ,
		_w28311_
	);
	LUT2 #(
		.INIT('h1)
	) name24265 (
		\T_TMODE[1]_pad ,
		_w27643_,
		_w28312_
	);
	LUT2 #(
		.INIT('h1)
	) name24266 (
		_w28311_,
		_w28312_,
		_w28313_
	);
	LUT2 #(
		.INIT('h4)
	) name24267 (
		_w21242_,
		_w28313_,
		_w28314_
	);
	LUT2 #(
		.INIT('h1)
	) name24268 (
		_w28310_,
		_w28314_,
		_w28315_
	);
	LUT2 #(
		.INIT('h1)
	) name24269 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w28204_,
		_w28316_
	);
	LUT2 #(
		.INIT('h4)
	) name24270 (
		\sice_SPC_reg[16]/P0001 ,
		_w28204_,
		_w28317_
	);
	LUT2 #(
		.INIT('h1)
	) name24271 (
		_w28316_,
		_w28317_,
		_w28318_
	);
	LUT2 #(
		.INIT('h2)
	) name24272 (
		_w21242_,
		_w28318_,
		_w28319_
	);
	LUT2 #(
		.INIT('h8)
	) name24273 (
		\T_TMODE[1]_pad ,
		\emc_ECMDreg_reg[16]/P0001 ,
		_w28320_
	);
	LUT2 #(
		.INIT('h1)
	) name24274 (
		\T_TMODE[1]_pad ,
		_w27669_,
		_w28321_
	);
	LUT2 #(
		.INIT('h1)
	) name24275 (
		_w28320_,
		_w28321_,
		_w28322_
	);
	LUT2 #(
		.INIT('h4)
	) name24276 (
		_w21242_,
		_w28322_,
		_w28323_
	);
	LUT2 #(
		.INIT('h1)
	) name24277 (
		_w28319_,
		_w28323_,
		_w28324_
	);
	LUT2 #(
		.INIT('h1)
	) name24278 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w28204_,
		_w28325_
	);
	LUT2 #(
		.INIT('h4)
	) name24279 (
		\sice_SPC_reg[15]/P0001 ,
		_w28204_,
		_w28326_
	);
	LUT2 #(
		.INIT('h1)
	) name24280 (
		_w28325_,
		_w28326_,
		_w28327_
	);
	LUT2 #(
		.INIT('h2)
	) name24281 (
		_w21242_,
		_w28327_,
		_w28328_
	);
	LUT2 #(
		.INIT('h4)
	) name24282 (
		_w21242_,
		_w27030_,
		_w28329_
	);
	LUT2 #(
		.INIT('h1)
	) name24283 (
		_w28328_,
		_w28329_,
		_w28330_
	);
	LUT2 #(
		.INIT('h1)
	) name24284 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w28204_,
		_w28331_
	);
	LUT2 #(
		.INIT('h4)
	) name24285 (
		\sice_SPC_reg[14]/P0001 ,
		_w28204_,
		_w28332_
	);
	LUT2 #(
		.INIT('h1)
	) name24286 (
		_w28331_,
		_w28332_,
		_w28333_
	);
	LUT2 #(
		.INIT('h2)
	) name24287 (
		_w21242_,
		_w28333_,
		_w28334_
	);
	LUT2 #(
		.INIT('h4)
	) name24288 (
		_w21242_,
		_w27077_,
		_w28335_
	);
	LUT2 #(
		.INIT('h1)
	) name24289 (
		_w28334_,
		_w28335_,
		_w28336_
	);
	LUT2 #(
		.INIT('h1)
	) name24290 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		_w28204_,
		_w28337_
	);
	LUT2 #(
		.INIT('h4)
	) name24291 (
		\sice_SPC_reg[13]/P0001 ,
		_w28204_,
		_w28338_
	);
	LUT2 #(
		.INIT('h1)
	) name24292 (
		_w28337_,
		_w28338_,
		_w28339_
	);
	LUT2 #(
		.INIT('h2)
	) name24293 (
		_w21242_,
		_w28339_,
		_w28340_
	);
	LUT2 #(
		.INIT('h4)
	) name24294 (
		_w21242_,
		_w27335_,
		_w28341_
	);
	LUT2 #(
		.INIT('h1)
	) name24295 (
		_w28340_,
		_w28341_,
		_w28342_
	);
	LUT2 #(
		.INIT('h1)
	) name24296 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w28204_,
		_w28343_
	);
	LUT2 #(
		.INIT('h4)
	) name24297 (
		\sice_SPC_reg[12]/P0001 ,
		_w28204_,
		_w28344_
	);
	LUT2 #(
		.INIT('h1)
	) name24298 (
		_w28343_,
		_w28344_,
		_w28345_
	);
	LUT2 #(
		.INIT('h2)
	) name24299 (
		_w21242_,
		_w28345_,
		_w28346_
	);
	LUT2 #(
		.INIT('h4)
	) name24300 (
		_w21242_,
		_w27363_,
		_w28347_
	);
	LUT2 #(
		.INIT('h1)
	) name24301 (
		_w28346_,
		_w28347_,
		_w28348_
	);
	LUT2 #(
		.INIT('h1)
	) name24302 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w28204_,
		_w28349_
	);
	LUT2 #(
		.INIT('h4)
	) name24303 (
		\sice_SPC_reg[11]/P0001 ,
		_w28204_,
		_w28350_
	);
	LUT2 #(
		.INIT('h1)
	) name24304 (
		_w28349_,
		_w28350_,
		_w28351_
	);
	LUT2 #(
		.INIT('h2)
	) name24305 (
		_w21242_,
		_w28351_,
		_w28352_
	);
	LUT2 #(
		.INIT('h4)
	) name24306 (
		_w21242_,
		_w27447_,
		_w28353_
	);
	LUT2 #(
		.INIT('h1)
	) name24307 (
		_w28352_,
		_w28353_,
		_w28354_
	);
	LUT2 #(
		.INIT('h1)
	) name24308 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w28204_,
		_w28355_
	);
	LUT2 #(
		.INIT('h4)
	) name24309 (
		\sice_SPC_reg[10]/P0001 ,
		_w28204_,
		_w28356_
	);
	LUT2 #(
		.INIT('h1)
	) name24310 (
		_w28355_,
		_w28356_,
		_w28357_
	);
	LUT2 #(
		.INIT('h2)
	) name24311 (
		_w21242_,
		_w28357_,
		_w28358_
	);
	LUT2 #(
		.INIT('h4)
	) name24312 (
		_w21242_,
		_w27475_,
		_w28359_
	);
	LUT2 #(
		.INIT('h1)
	) name24313 (
		_w28358_,
		_w28359_,
		_w28360_
	);
	LUT2 #(
		.INIT('h8)
	) name24314 (
		\sice_SPC_reg[21]/P0001 ,
		_w26969_,
		_w28361_
	);
	LUT2 #(
		.INIT('h2)
	) name24315 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w28277_,
		_w28362_
	);
	LUT2 #(
		.INIT('h1)
	) name24316 (
		_w28361_,
		_w28362_,
		_w28363_
	);
	LUT2 #(
		.INIT('h8)
	) name24317 (
		\sice_SPC_reg[20]/P0001 ,
		_w26969_,
		_w28364_
	);
	LUT2 #(
		.INIT('h2)
	) name24318 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w28286_,
		_w28365_
	);
	LUT2 #(
		.INIT('h1)
	) name24319 (
		_w28364_,
		_w28365_,
		_w28366_
	);
	LUT2 #(
		.INIT('h8)
	) name24320 (
		\sice_SPC_reg[19]/P0001 ,
		_w26969_,
		_w28367_
	);
	LUT2 #(
		.INIT('h2)
	) name24321 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w28295_,
		_w28368_
	);
	LUT2 #(
		.INIT('h1)
	) name24322 (
		_w28367_,
		_w28368_,
		_w28369_
	);
	LUT2 #(
		.INIT('h8)
	) name24323 (
		\sice_SPC_reg[18]/P0001 ,
		_w26969_,
		_w28370_
	);
	LUT2 #(
		.INIT('h2)
	) name24324 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w28304_,
		_w28371_
	);
	LUT2 #(
		.INIT('h1)
	) name24325 (
		_w28370_,
		_w28371_,
		_w28372_
	);
	LUT2 #(
		.INIT('h8)
	) name24326 (
		\sice_SPC_reg[17]/P0001 ,
		_w26969_,
		_w28373_
	);
	LUT2 #(
		.INIT('h2)
	) name24327 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w28313_,
		_w28374_
	);
	LUT2 #(
		.INIT('h1)
	) name24328 (
		_w28373_,
		_w28374_,
		_w28375_
	);
	LUT2 #(
		.INIT('h8)
	) name24329 (
		\sice_SPC_reg[16]/P0001 ,
		_w26969_,
		_w28376_
	);
	LUT2 #(
		.INIT('h2)
	) name24330 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w28322_,
		_w28377_
	);
	LUT2 #(
		.INIT('h1)
	) name24331 (
		_w28376_,
		_w28377_,
		_w28378_
	);
	LUT2 #(
		.INIT('h8)
	) name24332 (
		\sice_SPC_reg[23]/P0001 ,
		_w26969_,
		_w28379_
	);
	LUT2 #(
		.INIT('h2)
	) name24333 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w28259_,
		_w28380_
	);
	LUT2 #(
		.INIT('h1)
	) name24334 (
		_w28379_,
		_w28380_,
		_w28381_
	);
	LUT2 #(
		.INIT('h8)
	) name24335 (
		\sice_SPC_reg[22]/P0001 ,
		_w26969_,
		_w28382_
	);
	LUT2 #(
		.INIT('h2)
	) name24336 (
		\core_c_dec_rdCM_E_reg/NET0131 ,
		_w28268_,
		_w28383_
	);
	LUT2 #(
		.INIT('h1)
	) name24337 (
		_w28382_,
		_w28383_,
		_w28384_
	);
	LUT2 #(
		.INIT('h4)
	) name24338 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[8]/P0001 ,
		_w28385_
	);
	LUT2 #(
		.INIT('h8)
	) name24339 (
		_w6921_,
		_w10638_,
		_w28386_
	);
	LUT2 #(
		.INIT('h8)
	) name24340 (
		_w12520_,
		_w13152_,
		_w28387_
	);
	LUT2 #(
		.INIT('h4)
	) name24341 (
		_w5727_,
		_w13151_,
		_w28388_
	);
	LUT2 #(
		.INIT('h4)
	) name24342 (
		_w27389_,
		_w28388_,
		_w28389_
	);
	LUT2 #(
		.INIT('h1)
	) name24343 (
		_w28387_,
		_w28389_,
		_w28390_
	);
	LUT2 #(
		.INIT('h4)
	) name24344 (
		_w28386_,
		_w28390_,
		_w28391_
	);
	LUT2 #(
		.INIT('h2)
	) name24345 (
		\auctl_BSack_reg/NET0131 ,
		_w28391_,
		_w28392_
	);
	LUT2 #(
		.INIT('h1)
	) name24346 (
		_w28385_,
		_w28392_,
		_w28393_
	);
	LUT2 #(
		.INIT('h4)
	) name24347 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[9]/P0001 ,
		_w28394_
	);
	LUT2 #(
		.INIT('h8)
	) name24348 (
		_w6921_,
		_w10289_,
		_w28395_
	);
	LUT2 #(
		.INIT('h8)
	) name24349 (
		_w12802_,
		_w13152_,
		_w28396_
	);
	LUT2 #(
		.INIT('h4)
	) name24350 (
		_w27417_,
		_w28388_,
		_w28397_
	);
	LUT2 #(
		.INIT('h1)
	) name24351 (
		_w28396_,
		_w28397_,
		_w28398_
	);
	LUT2 #(
		.INIT('h4)
	) name24352 (
		_w28395_,
		_w28398_,
		_w28399_
	);
	LUT2 #(
		.INIT('h2)
	) name24353 (
		\auctl_BSack_reg/NET0131 ,
		_w28399_,
		_w28400_
	);
	LUT2 #(
		.INIT('h1)
	) name24354 (
		_w28394_,
		_w28400_,
		_w28401_
	);
	LUT2 #(
		.INIT('h4)
	) name24355 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[15]/P0001 ,
		_w28402_
	);
	LUT2 #(
		.INIT('h8)
	) name24356 (
		_w6921_,
		_w12743_,
		_w28403_
	);
	LUT2 #(
		.INIT('h8)
	) name24357 (
		_w13006_,
		_w13152_,
		_w28404_
	);
	LUT2 #(
		.INIT('h4)
	) name24358 (
		_w27028_,
		_w28388_,
		_w28405_
	);
	LUT2 #(
		.INIT('h1)
	) name24359 (
		_w28404_,
		_w28405_,
		_w28406_
	);
	LUT2 #(
		.INIT('h4)
	) name24360 (
		_w28403_,
		_w28406_,
		_w28407_
	);
	LUT2 #(
		.INIT('h2)
	) name24361 (
		\auctl_BSack_reg/NET0131 ,
		_w28407_,
		_w28408_
	);
	LUT2 #(
		.INIT('h1)
	) name24362 (
		_w28402_,
		_w28408_,
		_w28409_
	);
	LUT2 #(
		.INIT('h4)
	) name24363 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[14]/P0001 ,
		_w28410_
	);
	LUT2 #(
		.INIT('h8)
	) name24364 (
		_w6921_,
		_w12688_,
		_w28411_
	);
	LUT2 #(
		.INIT('h4)
	) name24365 (
		_w27075_,
		_w28388_,
		_w28412_
	);
	LUT2 #(
		.INIT('h8)
	) name24366 (
		_w12972_,
		_w13152_,
		_w28413_
	);
	LUT2 #(
		.INIT('h1)
	) name24367 (
		_w28411_,
		_w28412_,
		_w28414_
	);
	LUT2 #(
		.INIT('h4)
	) name24368 (
		_w28413_,
		_w28414_,
		_w28415_
	);
	LUT2 #(
		.INIT('h2)
	) name24369 (
		\auctl_BSack_reg/NET0131 ,
		_w28415_,
		_w28416_
	);
	LUT2 #(
		.INIT('h1)
	) name24370 (
		_w28410_,
		_w28416_,
		_w28417_
	);
	LUT2 #(
		.INIT('h4)
	) name24371 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[13]/P0001 ,
		_w28418_
	);
	LUT2 #(
		.INIT('h8)
	) name24372 (
		_w6921_,
		_w7340_,
		_w28419_
	);
	LUT2 #(
		.INIT('h8)
	) name24373 (
		_w12938_,
		_w13152_,
		_w28420_
	);
	LUT2 #(
		.INIT('h4)
	) name24374 (
		_w27333_,
		_w28388_,
		_w28421_
	);
	LUT2 #(
		.INIT('h1)
	) name24375 (
		_w28420_,
		_w28421_,
		_w28422_
	);
	LUT2 #(
		.INIT('h4)
	) name24376 (
		_w28419_,
		_w28422_,
		_w28423_
	);
	LUT2 #(
		.INIT('h2)
	) name24377 (
		\auctl_BSack_reg/NET0131 ,
		_w28423_,
		_w28424_
	);
	LUT2 #(
		.INIT('h1)
	) name24378 (
		_w28418_,
		_w28424_,
		_w28425_
	);
	LUT2 #(
		.INIT('h4)
	) name24379 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[12]/P0001 ,
		_w28426_
	);
	LUT2 #(
		.INIT('h8)
	) name24380 (
		_w6921_,
		_w9178_,
		_w28427_
	);
	LUT2 #(
		.INIT('h8)
	) name24381 (
		_w12904_,
		_w13152_,
		_w28428_
	);
	LUT2 #(
		.INIT('h4)
	) name24382 (
		_w27361_,
		_w28388_,
		_w28429_
	);
	LUT2 #(
		.INIT('h1)
	) name24383 (
		_w28428_,
		_w28429_,
		_w28430_
	);
	LUT2 #(
		.INIT('h4)
	) name24384 (
		_w28427_,
		_w28430_,
		_w28431_
	);
	LUT2 #(
		.INIT('h2)
	) name24385 (
		\auctl_BSack_reg/NET0131 ,
		_w28431_,
		_w28432_
	);
	LUT2 #(
		.INIT('h1)
	) name24386 (
		_w28426_,
		_w28432_,
		_w28433_
	);
	LUT2 #(
		.INIT('h4)
	) name24387 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[11]/P0001 ,
		_w28434_
	);
	LUT2 #(
		.INIT('h8)
	) name24388 (
		_w6921_,
		_w8460_,
		_w28435_
	);
	LUT2 #(
		.INIT('h8)
	) name24389 (
		_w12870_,
		_w13152_,
		_w28436_
	);
	LUT2 #(
		.INIT('h4)
	) name24390 (
		_w27445_,
		_w28388_,
		_w28437_
	);
	LUT2 #(
		.INIT('h1)
	) name24391 (
		_w28436_,
		_w28437_,
		_w28438_
	);
	LUT2 #(
		.INIT('h4)
	) name24392 (
		_w28435_,
		_w28438_,
		_w28439_
	);
	LUT2 #(
		.INIT('h2)
	) name24393 (
		\auctl_BSack_reg/NET0131 ,
		_w28439_,
		_w28440_
	);
	LUT2 #(
		.INIT('h1)
	) name24394 (
		_w28434_,
		_w28440_,
		_w28441_
	);
	LUT2 #(
		.INIT('h4)
	) name24395 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[10]/P0001 ,
		_w28442_
	);
	LUT2 #(
		.INIT('h8)
	) name24396 (
		_w6921_,
		_w7859_,
		_w28443_
	);
	LUT2 #(
		.INIT('h8)
	) name24397 (
		_w12836_,
		_w13152_,
		_w28444_
	);
	LUT2 #(
		.INIT('h4)
	) name24398 (
		_w27473_,
		_w28388_,
		_w28445_
	);
	LUT2 #(
		.INIT('h1)
	) name24399 (
		_w28444_,
		_w28445_,
		_w28446_
	);
	LUT2 #(
		.INIT('h4)
	) name24400 (
		_w28443_,
		_w28446_,
		_w28447_
	);
	LUT2 #(
		.INIT('h2)
	) name24401 (
		\auctl_BSack_reg/NET0131 ,
		_w28447_,
		_w28448_
	);
	LUT2 #(
		.INIT('h1)
	) name24402 (
		_w28442_,
		_w28448_,
		_w28449_
	);
	LUT2 #(
		.INIT('h1)
	) name24403 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w28204_,
		_w28450_
	);
	LUT2 #(
		.INIT('h4)
	) name24404 (
		\sice_SPC_reg[1]/P0001 ,
		_w28204_,
		_w28451_
	);
	LUT2 #(
		.INIT('h1)
	) name24405 (
		_w28450_,
		_w28451_,
		_w28452_
	);
	LUT2 #(
		.INIT('h2)
	) name24406 (
		_w21242_,
		_w28452_,
		_w28453_
	);
	LUT2 #(
		.INIT('h4)
	) name24407 (
		_w21242_,
		_w27273_,
		_w28454_
	);
	LUT2 #(
		.INIT('h1)
	) name24408 (
		_w28453_,
		_w28454_,
		_w28455_
	);
	LUT2 #(
		.INIT('h1)
	) name24409 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w28204_,
		_w28456_
	);
	LUT2 #(
		.INIT('h4)
	) name24410 (
		\sice_SPC_reg[0]/P0001 ,
		_w28204_,
		_w28457_
	);
	LUT2 #(
		.INIT('h1)
	) name24411 (
		_w28456_,
		_w28457_,
		_w28458_
	);
	LUT2 #(
		.INIT('h2)
	) name24412 (
		_w21242_,
		_w28458_,
		_w28459_
	);
	LUT2 #(
		.INIT('h4)
	) name24413 (
		_w21242_,
		_w27301_,
		_w28460_
	);
	LUT2 #(
		.INIT('h1)
	) name24414 (
		_w28459_,
		_w28460_,
		_w28461_
	);
	LUT2 #(
		.INIT('h4)
	) name24415 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[7]/P0001 ,
		_w28462_
	);
	LUT2 #(
		.INIT('h8)
	) name24416 (
		_w6921_,
		_w11265_,
		_w28463_
	);
	LUT2 #(
		.INIT('h4)
	) name24417 (
		_w27103_,
		_w28388_,
		_w28464_
	);
	LUT2 #(
		.INIT('h1)
	) name24418 (
		_w28463_,
		_w28464_,
		_w28465_
	);
	LUT2 #(
		.INIT('h2)
	) name24419 (
		\auctl_BSack_reg/NET0131 ,
		_w28465_,
		_w28466_
	);
	LUT2 #(
		.INIT('h1)
	) name24420 (
		_w28462_,
		_w28466_,
		_w28467_
	);
	LUT2 #(
		.INIT('h4)
	) name24421 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[6]/P0001 ,
		_w28468_
	);
	LUT2 #(
		.INIT('h8)
	) name24422 (
		_w6921_,
		_w11525_,
		_w28469_
	);
	LUT2 #(
		.INIT('h4)
	) name24423 (
		_w27131_,
		_w28388_,
		_w28470_
	);
	LUT2 #(
		.INIT('h1)
	) name24424 (
		_w28469_,
		_w28470_,
		_w28471_
	);
	LUT2 #(
		.INIT('h2)
	) name24425 (
		\auctl_BSack_reg/NET0131 ,
		_w28471_,
		_w28472_
	);
	LUT2 #(
		.INIT('h1)
	) name24426 (
		_w28468_,
		_w28472_,
		_w28473_
	);
	LUT2 #(
		.INIT('h4)
	) name24427 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[5]/P0001 ,
		_w28474_
	);
	LUT2 #(
		.INIT('h8)
	) name24428 (
		_w6921_,
		_w10911_,
		_w28475_
	);
	LUT2 #(
		.INIT('h4)
	) name24429 (
		_w27159_,
		_w28388_,
		_w28476_
	);
	LUT2 #(
		.INIT('h1)
	) name24430 (
		_w28475_,
		_w28476_,
		_w28477_
	);
	LUT2 #(
		.INIT('h2)
	) name24431 (
		\auctl_BSack_reg/NET0131 ,
		_w28477_,
		_w28478_
	);
	LUT2 #(
		.INIT('h1)
	) name24432 (
		_w28474_,
		_w28478_,
		_w28479_
	);
	LUT2 #(
		.INIT('h4)
	) name24433 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[4]/P0001 ,
		_w28480_
	);
	LUT2 #(
		.INIT('h8)
	) name24434 (
		_w6921_,
		_w10069_,
		_w28481_
	);
	LUT2 #(
		.INIT('h4)
	) name24435 (
		_w27187_,
		_w28388_,
		_w28482_
	);
	LUT2 #(
		.INIT('h1)
	) name24436 (
		_w28481_,
		_w28482_,
		_w28483_
	);
	LUT2 #(
		.INIT('h2)
	) name24437 (
		\auctl_BSack_reg/NET0131 ,
		_w28483_,
		_w28484_
	);
	LUT2 #(
		.INIT('h1)
	) name24438 (
		_w28480_,
		_w28484_,
		_w28485_
	);
	LUT2 #(
		.INIT('h4)
	) name24439 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[3]/P0001 ,
		_w28486_
	);
	LUT2 #(
		.INIT('h8)
	) name24440 (
		_w6921_,
		_w8113_,
		_w28487_
	);
	LUT2 #(
		.INIT('h4)
	) name24441 (
		_w27215_,
		_w28388_,
		_w28488_
	);
	LUT2 #(
		.INIT('h1)
	) name24442 (
		_w28487_,
		_w28488_,
		_w28489_
	);
	LUT2 #(
		.INIT('h2)
	) name24443 (
		\auctl_BSack_reg/NET0131 ,
		_w28489_,
		_w28490_
	);
	LUT2 #(
		.INIT('h1)
	) name24444 (
		_w28486_,
		_w28490_,
		_w28491_
	);
	LUT2 #(
		.INIT('h4)
	) name24445 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[2]/P0001 ,
		_w28492_
	);
	LUT2 #(
		.INIT('h8)
	) name24446 (
		_w6921_,
		_w8715_,
		_w28493_
	);
	LUT2 #(
		.INIT('h4)
	) name24447 (
		_w27243_,
		_w28388_,
		_w28494_
	);
	LUT2 #(
		.INIT('h1)
	) name24448 (
		_w28493_,
		_w28494_,
		_w28495_
	);
	LUT2 #(
		.INIT('h2)
	) name24449 (
		\auctl_BSack_reg/NET0131 ,
		_w28495_,
		_w28496_
	);
	LUT2 #(
		.INIT('h1)
	) name24450 (
		_w28492_,
		_w28496_,
		_w28497_
	);
	LUT2 #(
		.INIT('h4)
	) name24451 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[23]/P0001 ,
		_w28498_
	);
	LUT2 #(
		.INIT('h8)
	) name24452 (
		_w12771_,
		_w13152_,
		_w28499_
	);
	LUT2 #(
		.INIT('h4)
	) name24453 (
		_w27577_,
		_w28388_,
		_w28500_
	);
	LUT2 #(
		.INIT('h1)
	) name24454 (
		_w28499_,
		_w28500_,
		_w28501_
	);
	LUT2 #(
		.INIT('h2)
	) name24455 (
		\auctl_BSack_reg/NET0131 ,
		_w28501_,
		_w28502_
	);
	LUT2 #(
		.INIT('h1)
	) name24456 (
		_w28498_,
		_w28502_,
		_w28503_
	);
	LUT2 #(
		.INIT('h4)
	) name24457 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[22]/P0001 ,
		_w28504_
	);
	LUT2 #(
		.INIT('h8)
	) name24458 (
		_w12715_,
		_w13152_,
		_w28505_
	);
	LUT2 #(
		.INIT('h4)
	) name24459 (
		_w27603_,
		_w28388_,
		_w28506_
	);
	LUT2 #(
		.INIT('h1)
	) name24460 (
		_w28505_,
		_w28506_,
		_w28507_
	);
	LUT2 #(
		.INIT('h2)
	) name24461 (
		\auctl_BSack_reg/NET0131 ,
		_w28507_,
		_w28508_
	);
	LUT2 #(
		.INIT('h1)
	) name24462 (
		_w28504_,
		_w28508_,
		_w28509_
	);
	LUT2 #(
		.INIT('h4)
	) name24463 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[21]/P0001 ,
		_w28510_
	);
	LUT2 #(
		.INIT('h8)
	) name24464 (
		_w12658_,
		_w13152_,
		_w28511_
	);
	LUT2 #(
		.INIT('h4)
	) name24465 (
		_w27695_,
		_w28388_,
		_w28512_
	);
	LUT2 #(
		.INIT('h1)
	) name24466 (
		_w28511_,
		_w28512_,
		_w28513_
	);
	LUT2 #(
		.INIT('h2)
	) name24467 (
		\auctl_BSack_reg/NET0131 ,
		_w28513_,
		_w28514_
	);
	LUT2 #(
		.INIT('h1)
	) name24468 (
		_w28510_,
		_w28514_,
		_w28515_
	);
	LUT2 #(
		.INIT('h4)
	) name24469 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[20]/P0001 ,
		_w28516_
	);
	LUT2 #(
		.INIT('h8)
	) name24470 (
		_w12624_,
		_w13152_,
		_w28517_
	);
	LUT2 #(
		.INIT('h4)
	) name24471 (
		_w27721_,
		_w28388_,
		_w28518_
	);
	LUT2 #(
		.INIT('h1)
	) name24472 (
		_w28517_,
		_w28518_,
		_w28519_
	);
	LUT2 #(
		.INIT('h2)
	) name24473 (
		\auctl_BSack_reg/NET0131 ,
		_w28519_,
		_w28520_
	);
	LUT2 #(
		.INIT('h1)
	) name24474 (
		_w28516_,
		_w28520_,
		_w28521_
	);
	LUT2 #(
		.INIT('h4)
	) name24475 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[1]/P0001 ,
		_w28522_
	);
	LUT2 #(
		.INIT('h8)
	) name24476 (
		_w6921_,
		_w9435_,
		_w28523_
	);
	LUT2 #(
		.INIT('h4)
	) name24477 (
		_w27271_,
		_w28388_,
		_w28524_
	);
	LUT2 #(
		.INIT('h1)
	) name24478 (
		_w28523_,
		_w28524_,
		_w28525_
	);
	LUT2 #(
		.INIT('h2)
	) name24479 (
		\auctl_BSack_reg/NET0131 ,
		_w28525_,
		_w28526_
	);
	LUT2 #(
		.INIT('h1)
	) name24480 (
		_w28522_,
		_w28526_,
		_w28527_
	);
	LUT2 #(
		.INIT('h8)
	) name24481 (
		_w18262_,
		_w19409_,
		_w28528_
	);
	LUT2 #(
		.INIT('h1)
	) name24482 (
		_w18262_,
		_w19384_,
		_w28529_
	);
	LUT2 #(
		.INIT('h8)
	) name24483 (
		_w14664_,
		_w17801_,
		_w28530_
	);
	LUT2 #(
		.INIT('h1)
	) name24484 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 ,
		_w28530_,
		_w28531_
	);
	LUT2 #(
		.INIT('h2)
	) name24485 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w17807_,
		_w28532_
	);
	LUT2 #(
		.INIT('h1)
	) name24486 (
		_w19381_,
		_w28530_,
		_w28533_
	);
	LUT2 #(
		.INIT('h2)
	) name24487 (
		_w28532_,
		_w28533_,
		_w28534_
	);
	LUT2 #(
		.INIT('h2)
	) name24488 (
		_w18974_,
		_w19381_,
		_w28535_
	);
	LUT2 #(
		.INIT('h2)
	) name24489 (
		_w28534_,
		_w28535_,
		_w28536_
	);
	LUT2 #(
		.INIT('h1)
	) name24490 (
		_w28531_,
		_w28536_,
		_w28537_
	);
	LUT2 #(
		.INIT('h1)
	) name24491 (
		_w19385_,
		_w28537_,
		_w28538_
	);
	LUT2 #(
		.INIT('h1)
	) name24492 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[1]/P0001 ,
		_w28532_,
		_w28539_
	);
	LUT2 #(
		.INIT('h1)
	) name24493 (
		_w28538_,
		_w28539_,
		_w28540_
	);
	LUT2 #(
		.INIT('h2)
	) name24494 (
		_w28529_,
		_w28540_,
		_w28541_
	);
	LUT2 #(
		.INIT('h1)
	) name24495 (
		_w28528_,
		_w28541_,
		_w28542_
	);
	LUT2 #(
		.INIT('h1)
	) name24496 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w18847_,
		_w28543_
	);
	LUT2 #(
		.INIT('h2)
	) name24497 (
		_w4117_,
		_w5689_,
		_w28544_
	);
	LUT2 #(
		.INIT('h1)
	) name24498 (
		_w28543_,
		_w28544_,
		_w28545_
	);
	LUT2 #(
		.INIT('h2)
	) name24499 (
		_w5689_,
		_w13832_,
		_w28546_
	);
	LUT2 #(
		.INIT('h1)
	) name24500 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w28547_
	);
	LUT2 #(
		.INIT('h1)
	) name24501 (
		_w5689_,
		_w28547_,
		_w28548_
	);
	LUT2 #(
		.INIT('h1)
	) name24502 (
		_w28546_,
		_w28548_,
		_w28549_
	);
	LUT2 #(
		.INIT('h2)
	) name24503 (
		_w28545_,
		_w28549_,
		_w28550_
	);
	LUT2 #(
		.INIT('h8)
	) name24504 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w5689_,
		_w28551_
	);
	LUT2 #(
		.INIT('h8)
	) name24505 (
		_w13823_,
		_w28551_,
		_w28552_
	);
	LUT2 #(
		.INIT('h4)
	) name24506 (
		_w5689_,
		_w26356_,
		_w28553_
	);
	LUT2 #(
		.INIT('h4)
	) name24507 (
		_w26370_,
		_w28553_,
		_w28554_
	);
	LUT2 #(
		.INIT('h8)
	) name24508 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w28554_,
		_w28555_
	);
	LUT2 #(
		.INIT('h1)
	) name24509 (
		_w28552_,
		_w28555_,
		_w28556_
	);
	LUT2 #(
		.INIT('h1)
	) name24510 (
		_w8497_,
		_w28556_,
		_w28557_
	);
	LUT2 #(
		.INIT('h4)
	) name24511 (
		_w5689_,
		_w26353_,
		_w28558_
	);
	LUT2 #(
		.INIT('h8)
	) name24512 (
		_w26370_,
		_w28558_,
		_w28559_
	);
	LUT2 #(
		.INIT('h8)
	) name24513 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w17814_,
		_w28560_
	);
	LUT2 #(
		.INIT('h1)
	) name24514 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w19214_,
		_w28561_
	);
	LUT2 #(
		.INIT('h4)
	) name24515 (
		_w14586_,
		_w28561_,
		_w28562_
	);
	LUT2 #(
		.INIT('h1)
	) name24516 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w19278_,
		_w28563_
	);
	LUT2 #(
		.INIT('h8)
	) name24517 (
		_w19214_,
		_w28563_,
		_w28564_
	);
	LUT2 #(
		.INIT('h1)
	) name24518 (
		_w28560_,
		_w28564_,
		_w28565_
	);
	LUT2 #(
		.INIT('h4)
	) name24519 (
		_w28562_,
		_w28565_,
		_w28566_
	);
	LUT2 #(
		.INIT('h2)
	) name24520 (
		_w28559_,
		_w28566_,
		_w28567_
	);
	LUT2 #(
		.INIT('h8)
	) name24521 (
		\core_eu_em_mac_em_reg_s2_reg/P0000_reg_syn_2 ,
		_w26395_,
		_w28568_
	);
	LUT2 #(
		.INIT('h1)
	) name24522 (
		_w26388_,
		_w28568_,
		_w28569_
	);
	LUT2 #(
		.INIT('h4)
	) name24523 (
		_w26396_,
		_w26966_,
		_w28570_
	);
	LUT2 #(
		.INIT('h4)
	) name24524 (
		\core_eu_em_mac_em_reg_s0_reg/P0000_reg_syn_2 ,
		_w26396_,
		_w28571_
	);
	LUT2 #(
		.INIT('h1)
	) name24525 (
		_w28570_,
		_w28571_,
		_w28572_
	);
	LUT2 #(
		.INIT('h8)
	) name24526 (
		\core_eu_em_mac_em_reg_s1_reg/P0000_reg_syn_2 ,
		_w26396_,
		_w28573_
	);
	LUT2 #(
		.INIT('h2)
	) name24527 (
		_w26394_,
		_w28573_,
		_w28574_
	);
	LUT2 #(
		.INIT('h1)
	) name24528 (
		_w28572_,
		_w28574_,
		_w28575_
	);
	LUT2 #(
		.INIT('h8)
	) name24529 (
		_w17820_,
		_w28575_,
		_w28576_
	);
	LUT2 #(
		.INIT('h8)
	) name24530 (
		_w28572_,
		_w28574_,
		_w28577_
	);
	LUT2 #(
		.INIT('h1)
	) name24531 (
		_w12836_,
		_w28577_,
		_w28578_
	);
	LUT2 #(
		.INIT('h4)
	) name24532 (
		_w8715_,
		_w28577_,
		_w28579_
	);
	LUT2 #(
		.INIT('h1)
	) name24533 (
		_w28575_,
		_w28578_,
		_w28580_
	);
	LUT2 #(
		.INIT('h4)
	) name24534 (
		_w28579_,
		_w28580_,
		_w28581_
	);
	LUT2 #(
		.INIT('h1)
	) name24535 (
		_w28576_,
		_w28581_,
		_w28582_
	);
	LUT2 #(
		.INIT('h2)
	) name24536 (
		_w28569_,
		_w28582_,
		_w28583_
	);
	LUT2 #(
		.INIT('h4)
	) name24537 (
		_w28569_,
		_w28574_,
		_w28584_
	);
	LUT2 #(
		.INIT('h1)
	) name24538 (
		_w8715_,
		_w28572_,
		_w28585_
	);
	LUT2 #(
		.INIT('h4)
	) name24539 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w26379_,
		_w28586_
	);
	LUT2 #(
		.INIT('h4)
	) name24540 (
		_w26370_,
		_w28586_,
		_w28587_
	);
	LUT2 #(
		.INIT('h8)
	) name24541 (
		_w5689_,
		_w13821_,
		_w28588_
	);
	LUT2 #(
		.INIT('h1)
	) name24542 (
		_w28587_,
		_w28588_,
		_w28589_
	);
	LUT2 #(
		.INIT('h1)
	) name24543 (
		_w8558_,
		_w28589_,
		_w28590_
	);
	LUT2 #(
		.INIT('h8)
	) name24544 (
		_w5689_,
		_w13819_,
		_w28591_
	);
	LUT2 #(
		.INIT('h4)
	) name24545 (
		_w5689_,
		_w26371_,
		_w28592_
	);
	LUT2 #(
		.INIT('h4)
	) name24546 (
		_w26370_,
		_w28592_,
		_w28593_
	);
	LUT2 #(
		.INIT('h1)
	) name24547 (
		_w28591_,
		_w28593_,
		_w28594_
	);
	LUT2 #(
		.INIT('h1)
	) name24548 (
		_w8554_,
		_w28594_,
		_w28595_
	);
	LUT2 #(
		.INIT('h4)
	) name24549 (
		_w26370_,
		_w26380_,
		_w28596_
	);
	LUT2 #(
		.INIT('h8)
	) name24550 (
		_w5689_,
		_w13813_,
		_w28597_
	);
	LUT2 #(
		.INIT('h1)
	) name24551 (
		_w28596_,
		_w28597_,
		_w28598_
	);
	LUT2 #(
		.INIT('h1)
	) name24552 (
		_w8534_,
		_w28598_,
		_w28599_
	);
	LUT2 #(
		.INIT('h8)
	) name24553 (
		_w17804_,
		_w26370_,
		_w28600_
	);
	LUT2 #(
		.INIT('h8)
	) name24554 (
		_w7206_,
		_w28600_,
		_w28601_
	);
	LUT2 #(
		.INIT('h1)
	) name24555 (
		_w28586_,
		_w28592_,
		_w28602_
	);
	LUT2 #(
		.INIT('h2)
	) name24556 (
		_w28601_,
		_w28602_,
		_w28603_
	);
	LUT2 #(
		.INIT('h4)
	) name24557 (
		_w7206_,
		_w26379_,
		_w28604_
	);
	LUT2 #(
		.INIT('h8)
	) name24558 (
		_w28600_,
		_w28604_,
		_w28605_
	);
	LUT2 #(
		.INIT('h8)
	) name24559 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w28605_,
		_w28606_
	);
	LUT2 #(
		.INIT('h1)
	) name24560 (
		_w28603_,
		_w28606_,
		_w28607_
	);
	LUT2 #(
		.INIT('h1)
	) name24561 (
		_w28590_,
		_w28595_,
		_w28608_
	);
	LUT2 #(
		.INIT('h4)
	) name24562 (
		_w28599_,
		_w28608_,
		_w28609_
	);
	LUT2 #(
		.INIT('h8)
	) name24563 (
		_w28607_,
		_w28609_,
		_w28610_
	);
	LUT2 #(
		.INIT('h8)
	) name24564 (
		_w28572_,
		_w28610_,
		_w28611_
	);
	LUT2 #(
		.INIT('h2)
	) name24565 (
		_w28584_,
		_w28585_,
		_w28612_
	);
	LUT2 #(
		.INIT('h4)
	) name24566 (
		_w28611_,
		_w28612_,
		_w28613_
	);
	LUT2 #(
		.INIT('h1)
	) name24567 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w28614_
	);
	LUT2 #(
		.INIT('h2)
	) name24568 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w28615_
	);
	LUT2 #(
		.INIT('h1)
	) name24569 (
		_w28614_,
		_w28615_,
		_w28616_
	);
	LUT2 #(
		.INIT('h8)
	) name24570 (
		_w26370_,
		_w28616_,
		_w28617_
	);
	LUT2 #(
		.INIT('h8)
	) name24571 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w28553_,
		_w28618_
	);
	LUT2 #(
		.INIT('h8)
	) name24572 (
		_w28617_,
		_w28618_,
		_w28619_
	);
	LUT2 #(
		.INIT('h8)
	) name24573 (
		_w12836_,
		_w28619_,
		_w28620_
	);
	LUT2 #(
		.INIT('h4)
	) name24574 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w28554_,
		_w28621_
	);
	LUT2 #(
		.INIT('h4)
	) name24575 (
		\core_c_dec_IRE_reg[8]/NET0131 ,
		_w13823_,
		_w28622_
	);
	LUT2 #(
		.INIT('h8)
	) name24576 (
		_w5689_,
		_w28622_,
		_w28623_
	);
	LUT2 #(
		.INIT('h1)
	) name24577 (
		_w28621_,
		_w28623_,
		_w28624_
	);
	LUT2 #(
		.INIT('h1)
	) name24578 (
		_w8493_,
		_w28624_,
		_w28625_
	);
	LUT2 #(
		.INIT('h8)
	) name24579 (
		_w26370_,
		_w28553_,
		_w28626_
	);
	LUT2 #(
		.INIT('h8)
	) name24580 (
		_w28615_,
		_w28626_,
		_w28627_
	);
	LUT2 #(
		.INIT('h4)
	) name24581 (
		_w21124_,
		_w28627_,
		_w28628_
	);
	LUT2 #(
		.INIT('h4)
	) name24582 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w28553_,
		_w28629_
	);
	LUT2 #(
		.INIT('h8)
	) name24583 (
		_w28617_,
		_w28629_,
		_w28630_
	);
	LUT2 #(
		.INIT('h8)
	) name24584 (
		_w8715_,
		_w28630_,
		_w28631_
	);
	LUT2 #(
		.INIT('h8)
	) name24585 (
		_w5689_,
		_w13816_,
		_w28632_
	);
	LUT2 #(
		.INIT('h4)
	) name24586 (
		_w26370_,
		_w28558_,
		_w28633_
	);
	LUT2 #(
		.INIT('h1)
	) name24587 (
		_w28632_,
		_w28633_,
		_w28634_
	);
	LUT2 #(
		.INIT('h1)
	) name24588 (
		_w8585_,
		_w28634_,
		_w28635_
	);
	LUT2 #(
		.INIT('h8)
	) name24589 (
		_w28614_,
		_w28626_,
		_w28636_
	);
	LUT2 #(
		.INIT('h4)
	) name24590 (
		_w21174_,
		_w28636_,
		_w28637_
	);
	LUT2 #(
		.INIT('h1)
	) name24591 (
		_w28620_,
		_w28631_,
		_w28638_
	);
	LUT2 #(
		.INIT('h4)
	) name24592 (
		_w28635_,
		_w28638_,
		_w28639_
	);
	LUT2 #(
		.INIT('h1)
	) name24593 (
		_w28557_,
		_w28625_,
		_w28640_
	);
	LUT2 #(
		.INIT('h4)
	) name24594 (
		_w28637_,
		_w28640_,
		_w28641_
	);
	LUT2 #(
		.INIT('h8)
	) name24595 (
		_w28639_,
		_w28641_,
		_w28642_
	);
	LUT2 #(
		.INIT('h4)
	) name24596 (
		_w28628_,
		_w28642_,
		_w28643_
	);
	LUT2 #(
		.INIT('h4)
	) name24597 (
		_w28613_,
		_w28643_,
		_w28644_
	);
	LUT2 #(
		.INIT('h4)
	) name24598 (
		_w28583_,
		_w28644_,
		_w28645_
	);
	LUT2 #(
		.INIT('h4)
	) name24599 (
		_w28567_,
		_w28645_,
		_w28646_
	);
	LUT2 #(
		.INIT('h2)
	) name24600 (
		_w28550_,
		_w28646_,
		_w28647_
	);
	LUT2 #(
		.INIT('h8)
	) name24601 (
		\core_c_dec_MACop_E_reg/P0001 ,
		_w5689_,
		_w28648_
	);
	LUT2 #(
		.INIT('h1)
	) name24602 (
		_w18848_,
		_w28648_,
		_w28649_
	);
	LUT2 #(
		.INIT('h4)
	) name24603 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[2]/P0001 ,
		_w28649_,
		_w28650_
	);
	LUT2 #(
		.INIT('h2)
	) name24604 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w5689_,
		_w28651_
	);
	LUT2 #(
		.INIT('h1)
	) name24605 (
		_w28551_,
		_w28651_,
		_w28652_
	);
	LUT2 #(
		.INIT('h8)
	) name24606 (
		_w8550_,
		_w28652_,
		_w28653_
	);
	LUT2 #(
		.INIT('h2)
	) name24607 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTMX1_E_reg/P0001 ,
		_w28654_
	);
	LUT2 #(
		.INIT('h4)
	) name24608 (
		_w5689_,
		_w18847_,
		_w28655_
	);
	LUT2 #(
		.INIT('h1)
	) name24609 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		\core_c_dec_MTMX0_E_reg/P0001 ,
		_w28656_
	);
	LUT2 #(
		.INIT('h4)
	) name24610 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w28547_,
		_w28657_
	);
	LUT2 #(
		.INIT('h1)
	) name24611 (
		_w28654_,
		_w28656_,
		_w28658_
	);
	LUT2 #(
		.INIT('h8)
	) name24612 (
		_w28657_,
		_w28658_,
		_w28659_
	);
	LUT2 #(
		.INIT('h8)
	) name24613 (
		_w28655_,
		_w28659_,
		_w28660_
	);
	LUT2 #(
		.INIT('h2)
	) name24614 (
		_w8538_,
		_w28652_,
		_w28661_
	);
	LUT2 #(
		.INIT('h1)
	) name24615 (
		_w28653_,
		_w28660_,
		_w28662_
	);
	LUT2 #(
		.INIT('h4)
	) name24616 (
		_w28661_,
		_w28662_,
		_w28663_
	);
	LUT2 #(
		.INIT('h8)
	) name24617 (
		_w17814_,
		_w28660_,
		_w28664_
	);
	LUT2 #(
		.INIT('h1)
	) name24618 (
		_w28649_,
		_w28663_,
		_w28665_
	);
	LUT2 #(
		.INIT('h4)
	) name24619 (
		_w28664_,
		_w28665_,
		_w28666_
	);
	LUT2 #(
		.INIT('h1)
	) name24620 (
		_w28550_,
		_w28650_,
		_w28667_
	);
	LUT2 #(
		.INIT('h4)
	) name24621 (
		_w28666_,
		_w28667_,
		_w28668_
	);
	LUT2 #(
		.INIT('h1)
	) name24622 (
		_w28647_,
		_w28668_,
		_w28669_
	);
	LUT2 #(
		.INIT('h4)
	) name24623 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[19]/P0001 ,
		_w28670_
	);
	LUT2 #(
		.INIT('h8)
	) name24624 (
		_w12590_,
		_w13152_,
		_w28671_
	);
	LUT2 #(
		.INIT('h4)
	) name24625 (
		_w27747_,
		_w28388_,
		_w28672_
	);
	LUT2 #(
		.INIT('h1)
	) name24626 (
		_w28671_,
		_w28672_,
		_w28673_
	);
	LUT2 #(
		.INIT('h2)
	) name24627 (
		\auctl_BSack_reg/NET0131 ,
		_w28673_,
		_w28674_
	);
	LUT2 #(
		.INIT('h1)
	) name24628 (
		_w28670_,
		_w28674_,
		_w28675_
	);
	LUT2 #(
		.INIT('h4)
	) name24629 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[18]/P0001 ,
		_w28676_
	);
	LUT2 #(
		.INIT('h8)
	) name24630 (
		_w12556_,
		_w13152_,
		_w28677_
	);
	LUT2 #(
		.INIT('h4)
	) name24631 (
		_w27773_,
		_w28388_,
		_w28678_
	);
	LUT2 #(
		.INIT('h1)
	) name24632 (
		_w28677_,
		_w28678_,
		_w28679_
	);
	LUT2 #(
		.INIT('h2)
	) name24633 (
		\auctl_BSack_reg/NET0131 ,
		_w28679_,
		_w28680_
	);
	LUT2 #(
		.INIT('h1)
	) name24634 (
		_w28676_,
		_w28680_,
		_w28681_
	);
	LUT2 #(
		.INIT('h4)
	) name24635 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[17]/P0001 ,
		_w28682_
	);
	LUT2 #(
		.INIT('h8)
	) name24636 (
		_w13075_,
		_w13152_,
		_w28683_
	);
	LUT2 #(
		.INIT('h4)
	) name24637 (
		_w27643_,
		_w28388_,
		_w28684_
	);
	LUT2 #(
		.INIT('h1)
	) name24638 (
		_w28683_,
		_w28684_,
		_w28685_
	);
	LUT2 #(
		.INIT('h2)
	) name24639 (
		\auctl_BSack_reg/NET0131 ,
		_w28685_,
		_w28686_
	);
	LUT2 #(
		.INIT('h1)
	) name24640 (
		_w28682_,
		_w28686_,
		_w28687_
	);
	LUT2 #(
		.INIT('h4)
	) name24641 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[16]/P0001 ,
		_w28688_
	);
	LUT2 #(
		.INIT('h8)
	) name24642 (
		_w13041_,
		_w13152_,
		_w28689_
	);
	LUT2 #(
		.INIT('h4)
	) name24643 (
		_w27669_,
		_w28388_,
		_w28690_
	);
	LUT2 #(
		.INIT('h1)
	) name24644 (
		_w28689_,
		_w28690_,
		_w28691_
	);
	LUT2 #(
		.INIT('h2)
	) name24645 (
		\auctl_BSack_reg/NET0131 ,
		_w28691_,
		_w28692_
	);
	LUT2 #(
		.INIT('h1)
	) name24646 (
		_w28688_,
		_w28692_,
		_w28693_
	);
	LUT2 #(
		.INIT('h4)
	) name24647 (
		\auctl_BSack_reg/NET0131 ,
		\bdma_BWdataBUF_h_reg[0]/P0001 ,
		_w28694_
	);
	LUT2 #(
		.INIT('h8)
	) name24648 (
		_w6921_,
		_w7607_,
		_w28695_
	);
	LUT2 #(
		.INIT('h4)
	) name24649 (
		_w27299_,
		_w28388_,
		_w28696_
	);
	LUT2 #(
		.INIT('h1)
	) name24650 (
		_w28695_,
		_w28696_,
		_w28697_
	);
	LUT2 #(
		.INIT('h2)
	) name24651 (
		\auctl_BSack_reg/NET0131 ,
		_w28697_,
		_w28698_
	);
	LUT2 #(
		.INIT('h1)
	) name24652 (
		_w28694_,
		_w28698_,
		_w28699_
	);
	LUT2 #(
		.INIT('h2)
	) name24653 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w5689_,
		_w28700_
	);
	LUT2 #(
		.INIT('h8)
	) name24654 (
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w5689_,
		_w28701_
	);
	LUT2 #(
		.INIT('h1)
	) name24655 (
		_w28700_,
		_w28701_,
		_w28702_
	);
	LUT2 #(
		.INIT('h2)
	) name24656 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w5689_,
		_w28703_
	);
	LUT2 #(
		.INIT('h8)
	) name24657 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w5689_,
		_w28704_
	);
	LUT2 #(
		.INIT('h1)
	) name24658 (
		_w28703_,
		_w28704_,
		_w28705_
	);
	LUT2 #(
		.INIT('h1)
	) name24659 (
		_w28702_,
		_w28705_,
		_w28706_
	);
	LUT2 #(
		.INIT('h1)
	) name24660 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_MTMY0_E_reg/P0001 ,
		_w28707_
	);
	LUT2 #(
		.INIT('h2)
	) name24661 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		\core_c_dec_MTMY1_E_reg/P0001 ,
		_w28708_
	);
	LUT2 #(
		.INIT('h1)
	) name24662 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w28709_
	);
	LUT2 #(
		.INIT('h4)
	) name24663 (
		_w28707_,
		_w28709_,
		_w28710_
	);
	LUT2 #(
		.INIT('h4)
	) name24664 (
		_w28708_,
		_w28710_,
		_w28711_
	);
	LUT2 #(
		.INIT('h4)
	) name24665 (
		_w26358_,
		_w28711_,
		_w28712_
	);
	LUT2 #(
		.INIT('h8)
	) name24666 (
		_w28655_,
		_w28712_,
		_w28713_
	);
	LUT2 #(
		.INIT('h1)
	) name24667 (
		_w28706_,
		_w28713_,
		_w28714_
	);
	LUT2 #(
		.INIT('h1)
	) name24668 (
		_w5689_,
		_w21525_,
		_w28715_
	);
	LUT2 #(
		.INIT('h4)
	) name24669 (
		\core_eu_em_mac_em_reg_Sq_E_reg/P0001 ,
		_w5689_,
		_w28716_
	);
	LUT2 #(
		.INIT('h1)
	) name24670 (
		_w28715_,
		_w28716_,
		_w28717_
	);
	LUT2 #(
		.INIT('h8)
	) name24671 (
		_w28714_,
		_w28717_,
		_w28718_
	);
	LUT2 #(
		.INIT('h8)
	) name24672 (
		_w28550_,
		_w28718_,
		_w28719_
	);
	LUT2 #(
		.INIT('h4)
	) name24673 (
		_w28544_,
		_w28718_,
		_w28720_
	);
	LUT2 #(
		.INIT('h8)
	) name24674 (
		_w28660_,
		_w28720_,
		_w28721_
	);
	LUT2 #(
		.INIT('h4)
	) name24675 (
		_w4117_,
		_w28713_,
		_w28722_
	);
	LUT2 #(
		.INIT('h4)
	) name24676 (
		\core_c_dec_Double_E_reg/P0001 ,
		_w28722_,
		_w28723_
	);
	LUT2 #(
		.INIT('h1)
	) name24677 (
		_w28721_,
		_w28723_,
		_w28724_
	);
	LUT2 #(
		.INIT('h1)
	) name24678 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w28724_,
		_w28725_
	);
	LUT2 #(
		.INIT('h8)
	) name24679 (
		\core_c_dec_accPM_E_reg/P0001 ,
		_w28721_,
		_w28726_
	);
	LUT2 #(
		.INIT('h4)
	) name24680 (
		_w21991_,
		_w28722_,
		_w28727_
	);
	LUT2 #(
		.INIT('h1)
	) name24681 (
		_w28726_,
		_w28727_,
		_w28728_
	);
	LUT2 #(
		.INIT('h1)
	) name24682 (
		_w28725_,
		_w28728_,
		_w28729_
	);
	LUT2 #(
		.INIT('h8)
	) name24683 (
		_w12836_,
		_w28729_,
		_w28730_
	);
	LUT2 #(
		.INIT('h8)
	) name24684 (
		_w8715_,
		_w28725_,
		_w28731_
	);
	LUT2 #(
		.INIT('h8)
	) name24685 (
		_w8546_,
		_w28705_,
		_w28732_
	);
	LUT2 #(
		.INIT('h1)
	) name24686 (
		_w28544_,
		_w28717_,
		_w28733_
	);
	LUT2 #(
		.INIT('h8)
	) name24687 (
		_w28714_,
		_w28733_,
		_w28734_
	);
	LUT2 #(
		.INIT('h8)
	) name24688 (
		_w28702_,
		_w28734_,
		_w28735_
	);
	LUT2 #(
		.INIT('h2)
	) name24689 (
		_w8542_,
		_w28705_,
		_w28736_
	);
	LUT2 #(
		.INIT('h1)
	) name24690 (
		_w28732_,
		_w28736_,
		_w28737_
	);
	LUT2 #(
		.INIT('h8)
	) name24691 (
		_w28735_,
		_w28737_,
		_w28738_
	);
	LUT2 #(
		.INIT('h8)
	) name24692 (
		_w28549_,
		_w28720_,
		_w28739_
	);
	LUT2 #(
		.INIT('h8)
	) name24693 (
		_w28663_,
		_w28739_,
		_w28740_
	);
	LUT2 #(
		.INIT('h4)
	) name24694 (
		_w28702_,
		_w28734_,
		_w28741_
	);
	LUT2 #(
		.INIT('h1)
	) name24695 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[2]/P0001 ,
		_w28742_
	);
	LUT2 #(
		.INIT('h2)
	) name24696 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[2]/P0001 ,
		_w28743_
	);
	LUT2 #(
		.INIT('h1)
	) name24697 (
		_w28742_,
		_w28743_,
		_w28744_
	);
	LUT2 #(
		.INIT('h8)
	) name24698 (
		_w28741_,
		_w28744_,
		_w28745_
	);
	LUT2 #(
		.INIT('h1)
	) name24699 (
		_w28738_,
		_w28740_,
		_w28746_
	);
	LUT2 #(
		.INIT('h4)
	) name24700 (
		_w28745_,
		_w28746_,
		_w28747_
	);
	LUT2 #(
		.INIT('h4)
	) name24701 (
		_w28730_,
		_w28747_,
		_w28748_
	);
	LUT2 #(
		.INIT('h4)
	) name24702 (
		_w28731_,
		_w28748_,
		_w28749_
	);
	LUT2 #(
		.INIT('h1)
	) name24703 (
		_w28543_,
		_w28749_,
		_w28750_
	);
	LUT2 #(
		.INIT('h2)
	) name24704 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[2]/P0001 ,
		_w28545_,
		_w28751_
	);
	LUT2 #(
		.INIT('h1)
	) name24705 (
		_w28750_,
		_w28751_,
		_w28752_
	);
	LUT2 #(
		.INIT('h1)
	) name24706 (
		_w28719_,
		_w28752_,
		_w28753_
	);
	LUT2 #(
		.INIT('h4)
	) name24707 (
		_w28646_,
		_w28719_,
		_w28754_
	);
	LUT2 #(
		.INIT('h1)
	) name24708 (
		_w28753_,
		_w28754_,
		_w28755_
	);
	LUT2 #(
		.INIT('h8)
	) name24709 (
		\tm_tcr_reg_DO_reg[14]/NET0131 ,
		_w20355_,
		_w28756_
	);
	LUT2 #(
		.INIT('h4)
	) name24710 (
		\tm_tpr_reg_DO_reg[14]/NET0131 ,
		_w22400_,
		_w28757_
	);
	LUT2 #(
		.INIT('h2)
	) name24711 (
		\tm_TCR_TMP_reg[14]/NET0131 ,
		_w25841_,
		_w28758_
	);
	LUT2 #(
		.INIT('h1)
	) name24712 (
		_w22400_,
		_w25842_,
		_w28759_
	);
	LUT2 #(
		.INIT('h4)
	) name24713 (
		_w28758_,
		_w28759_,
		_w28760_
	);
	LUT2 #(
		.INIT('h1)
	) name24714 (
		_w20355_,
		_w28757_,
		_w28761_
	);
	LUT2 #(
		.INIT('h4)
	) name24715 (
		_w28760_,
		_w28761_,
		_w28762_
	);
	LUT2 #(
		.INIT('h1)
	) name24716 (
		_w28756_,
		_w28762_,
		_w28763_
	);
	LUT2 #(
		.INIT('h8)
	) name24717 (
		_w14752_,
		_w19409_,
		_w28764_
	);
	LUT2 #(
		.INIT('h1)
	) name24718 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 ,
		_w17799_,
		_w28765_
	);
	LUT2 #(
		.INIT('h4)
	) name24719 (
		_w17809_,
		_w18974_,
		_w28766_
	);
	LUT2 #(
		.INIT('h2)
	) name24720 (
		_w17811_,
		_w28766_,
		_w28767_
	);
	LUT2 #(
		.INIT('h1)
	) name24721 (
		_w28765_,
		_w28767_,
		_w28768_
	);
	LUT2 #(
		.INIT('h1)
	) name24722 (
		_w17823_,
		_w28768_,
		_w28769_
	);
	LUT2 #(
		.INIT('h1)
	) name24723 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[1]/P0001 ,
		_w17808_,
		_w28770_
	);
	LUT2 #(
		.INIT('h1)
	) name24724 (
		_w28769_,
		_w28770_,
		_w28771_
	);
	LUT2 #(
		.INIT('h2)
	) name24725 (
		_w17829_,
		_w28771_,
		_w28772_
	);
	LUT2 #(
		.INIT('h1)
	) name24726 (
		_w28764_,
		_w28772_,
		_w28773_
	);
	LUT2 #(
		.INIT('h4)
	) name24727 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[0]/P0001 ,
		_w28774_
	);
	LUT2 #(
		.INIT('h2)
	) name24728 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w20953_,
		_w28775_
	);
	LUT2 #(
		.INIT('h2)
	) name24729 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w28774_,
		_w28776_
	);
	LUT2 #(
		.INIT('h4)
	) name24730 (
		_w28775_,
		_w28776_,
		_w28777_
	);
	LUT2 #(
		.INIT('h8)
	) name24731 (
		_w7607_,
		_w20869_,
		_w28778_
	);
	LUT2 #(
		.INIT('h2)
	) name24732 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		_w20869_,
		_w28779_
	);
	LUT2 #(
		.INIT('h1)
	) name24733 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w28779_,
		_w28780_
	);
	LUT2 #(
		.INIT('h4)
	) name24734 (
		_w28778_,
		_w28780_,
		_w28781_
	);
	LUT2 #(
		.INIT('h1)
	) name24735 (
		_w28777_,
		_w28781_,
		_w28782_
	);
	LUT2 #(
		.INIT('h1)
	) name24736 (
		_w20868_,
		_w28782_,
		_w28783_
	);
	LUT2 #(
		.INIT('h4)
	) name24737 (
		\sport0_rxctl_RXSHT_reg[0]/P0001 ,
		_w20868_,
		_w28784_
	);
	LUT2 #(
		.INIT('h1)
	) name24738 (
		_w28783_,
		_w28784_,
		_w28785_
	);
	LUT2 #(
		.INIT('h4)
	) name24739 (
		\sport1_cfg_SP_ENg_D1_reg/P0001 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w28786_
	);
	LUT2 #(
		.INIT('h8)
	) name24740 (
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w28786_,
		_w28787_
	);
	LUT2 #(
		.INIT('h1)
	) name24741 (
		\IRFS1_pad ,
		\ITFS1_pad ,
		_w28788_
	);
	LUT2 #(
		.INIT('h2)
	) name24742 (
		\sport1_cfg_FSi_cnt_reg[8]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w28789_
	);
	LUT2 #(
		.INIT('h4)
	) name24743 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w28790_
	);
	LUT2 #(
		.INIT('h4)
	) name24744 (
		\sport1_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w28791_
	);
	LUT2 #(
		.INIT('h2)
	) name24745 (
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w28792_
	);
	LUT2 #(
		.INIT('h2)
	) name24746 (
		\sport1_cfg_FSi_cnt_reg[5]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w28793_
	);
	LUT2 #(
		.INIT('h4)
	) name24747 (
		\sport1_cfg_FSi_cnt_reg[8]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w28794_
	);
	LUT2 #(
		.INIT('h4)
	) name24748 (
		\sport1_cfg_FSi_cnt_reg[5]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w28795_
	);
	LUT2 #(
		.INIT('h4)
	) name24749 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w28796_
	);
	LUT2 #(
		.INIT('h4)
	) name24750 (
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w28797_
	);
	LUT2 #(
		.INIT('h4)
	) name24751 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w28798_
	);
	LUT2 #(
		.INIT('h2)
	) name24752 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w28799_
	);
	LUT2 #(
		.INIT('h4)
	) name24753 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w28800_
	);
	LUT2 #(
		.INIT('h4)
	) name24754 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w28801_
	);
	LUT2 #(
		.INIT('h4)
	) name24755 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w28802_
	);
	LUT2 #(
		.INIT('h2)
	) name24756 (
		\sport1_cfg_FSi_cnt_reg[15]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w28803_
	);
	LUT2 #(
		.INIT('h2)
	) name24757 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w28804_
	);
	LUT2 #(
		.INIT('h2)
	) name24758 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w28805_
	);
	LUT2 #(
		.INIT('h2)
	) name24759 (
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w28806_
	);
	LUT2 #(
		.INIT('h2)
	) name24760 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w28807_
	);
	LUT2 #(
		.INIT('h2)
	) name24761 (
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w28808_
	);
	LUT2 #(
		.INIT('h2)
	) name24762 (
		\sport1_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w28809_
	);
	LUT2 #(
		.INIT('h2)
	) name24763 (
		\sport1_cfg_FSi_cnt_reg[14]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w28810_
	);
	LUT2 #(
		.INIT('h4)
	) name24764 (
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w28811_
	);
	LUT2 #(
		.INIT('h2)
	) name24765 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w28812_
	);
	LUT2 #(
		.INIT('h4)
	) name24766 (
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w28813_
	);
	LUT2 #(
		.INIT('h4)
	) name24767 (
		\sport1_cfg_FSi_cnt_reg[14]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w28814_
	);
	LUT2 #(
		.INIT('h4)
	) name24768 (
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w28815_
	);
	LUT2 #(
		.INIT('h2)
	) name24769 (
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w28816_
	);
	LUT2 #(
		.INIT('h2)
	) name24770 (
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w28817_
	);
	LUT2 #(
		.INIT('h4)
	) name24771 (
		\sport1_cfg_FSi_cnt_reg[15]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w28818_
	);
	LUT2 #(
		.INIT('h2)
	) name24772 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w28819_
	);
	LUT2 #(
		.INIT('h4)
	) name24773 (
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w28820_
	);
	LUT2 #(
		.INIT('h1)
	) name24774 (
		_w28789_,
		_w28790_,
		_w28821_
	);
	LUT2 #(
		.INIT('h1)
	) name24775 (
		_w28791_,
		_w28792_,
		_w28822_
	);
	LUT2 #(
		.INIT('h1)
	) name24776 (
		_w28793_,
		_w28794_,
		_w28823_
	);
	LUT2 #(
		.INIT('h1)
	) name24777 (
		_w28795_,
		_w28796_,
		_w28824_
	);
	LUT2 #(
		.INIT('h1)
	) name24778 (
		_w28797_,
		_w28798_,
		_w28825_
	);
	LUT2 #(
		.INIT('h1)
	) name24779 (
		_w28799_,
		_w28800_,
		_w28826_
	);
	LUT2 #(
		.INIT('h1)
	) name24780 (
		_w28801_,
		_w28802_,
		_w28827_
	);
	LUT2 #(
		.INIT('h1)
	) name24781 (
		_w28803_,
		_w28804_,
		_w28828_
	);
	LUT2 #(
		.INIT('h1)
	) name24782 (
		_w28805_,
		_w28806_,
		_w28829_
	);
	LUT2 #(
		.INIT('h1)
	) name24783 (
		_w28807_,
		_w28808_,
		_w28830_
	);
	LUT2 #(
		.INIT('h1)
	) name24784 (
		_w28809_,
		_w28810_,
		_w28831_
	);
	LUT2 #(
		.INIT('h1)
	) name24785 (
		_w28811_,
		_w28812_,
		_w28832_
	);
	LUT2 #(
		.INIT('h1)
	) name24786 (
		_w28813_,
		_w28814_,
		_w28833_
	);
	LUT2 #(
		.INIT('h1)
	) name24787 (
		_w28815_,
		_w28816_,
		_w28834_
	);
	LUT2 #(
		.INIT('h1)
	) name24788 (
		_w28817_,
		_w28818_,
		_w28835_
	);
	LUT2 #(
		.INIT('h1)
	) name24789 (
		_w28819_,
		_w28820_,
		_w28836_
	);
	LUT2 #(
		.INIT('h8)
	) name24790 (
		_w28835_,
		_w28836_,
		_w28837_
	);
	LUT2 #(
		.INIT('h8)
	) name24791 (
		_w28833_,
		_w28834_,
		_w28838_
	);
	LUT2 #(
		.INIT('h8)
	) name24792 (
		_w28831_,
		_w28832_,
		_w28839_
	);
	LUT2 #(
		.INIT('h8)
	) name24793 (
		_w28829_,
		_w28830_,
		_w28840_
	);
	LUT2 #(
		.INIT('h8)
	) name24794 (
		_w28827_,
		_w28828_,
		_w28841_
	);
	LUT2 #(
		.INIT('h8)
	) name24795 (
		_w28825_,
		_w28826_,
		_w28842_
	);
	LUT2 #(
		.INIT('h8)
	) name24796 (
		_w28823_,
		_w28824_,
		_w28843_
	);
	LUT2 #(
		.INIT('h8)
	) name24797 (
		_w28821_,
		_w28822_,
		_w28844_
	);
	LUT2 #(
		.INIT('h8)
	) name24798 (
		_w28843_,
		_w28844_,
		_w28845_
	);
	LUT2 #(
		.INIT('h8)
	) name24799 (
		_w28841_,
		_w28842_,
		_w28846_
	);
	LUT2 #(
		.INIT('h8)
	) name24800 (
		_w28839_,
		_w28840_,
		_w28847_
	);
	LUT2 #(
		.INIT('h8)
	) name24801 (
		_w28837_,
		_w28838_,
		_w28848_
	);
	LUT2 #(
		.INIT('h8)
	) name24802 (
		_w28847_,
		_w28848_,
		_w28849_
	);
	LUT2 #(
		.INIT('h8)
	) name24803 (
		_w28845_,
		_w28846_,
		_w28850_
	);
	LUT2 #(
		.INIT('h8)
	) name24804 (
		_w28849_,
		_w28850_,
		_w28851_
	);
	LUT2 #(
		.INIT('h1)
	) name24805 (
		_w28788_,
		_w28851_,
		_w28852_
	);
	LUT2 #(
		.INIT('h8)
	) name24806 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w28853_
	);
	LUT2 #(
		.INIT('h4)
	) name24807 (
		_w28852_,
		_w28853_,
		_w28854_
	);
	LUT2 #(
		.INIT('h1)
	) name24808 (
		_w28786_,
		_w28854_,
		_w28855_
	);
	LUT2 #(
		.INIT('h8)
	) name24809 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w28856_
	);
	LUT2 #(
		.INIT('h8)
	) name24810 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		_w28856_,
		_w28857_
	);
	LUT2 #(
		.INIT('h8)
	) name24811 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		_w28857_,
		_w28858_
	);
	LUT2 #(
		.INIT('h8)
	) name24812 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		_w28858_,
		_w28859_
	);
	LUT2 #(
		.INIT('h8)
	) name24813 (
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		_w28859_,
		_w28860_
	);
	LUT2 #(
		.INIT('h8)
	) name24814 (
		\sport1_cfg_FSi_cnt_reg[5]/NET0131 ,
		_w28860_,
		_w28861_
	);
	LUT2 #(
		.INIT('h8)
	) name24815 (
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		_w28861_,
		_w28862_
	);
	LUT2 #(
		.INIT('h8)
	) name24816 (
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		_w28862_,
		_w28863_
	);
	LUT2 #(
		.INIT('h8)
	) name24817 (
		\sport1_cfg_FSi_cnt_reg[8]/NET0131 ,
		_w28863_,
		_w28864_
	);
	LUT2 #(
		.INIT('h8)
	) name24818 (
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w28864_,
		_w28865_
	);
	LUT2 #(
		.INIT('h8)
	) name24819 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		_w28865_,
		_w28866_
	);
	LUT2 #(
		.INIT('h8)
	) name24820 (
		\sport1_cfg_FSi_cnt_reg[11]/NET0131 ,
		_w28866_,
		_w28867_
	);
	LUT2 #(
		.INIT('h8)
	) name24821 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		_w28867_,
		_w28868_
	);
	LUT2 #(
		.INIT('h8)
	) name24822 (
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		_w28868_,
		_w28869_
	);
	LUT2 #(
		.INIT('h8)
	) name24823 (
		\sport1_cfg_FSi_cnt_reg[14]/NET0131 ,
		_w28869_,
		_w28870_
	);
	LUT2 #(
		.INIT('h1)
	) name24824 (
		\sport1_cfg_FSi_cnt_reg[15]/NET0131 ,
		_w28870_,
		_w28871_
	);
	LUT2 #(
		.INIT('h8)
	) name24825 (
		\sport1_cfg_FSi_cnt_reg[15]/NET0131 ,
		_w28870_,
		_w28872_
	);
	LUT2 #(
		.INIT('h2)
	) name24826 (
		_w28855_,
		_w28871_,
		_w28873_
	);
	LUT2 #(
		.INIT('h4)
	) name24827 (
		_w28872_,
		_w28873_,
		_w28874_
	);
	LUT2 #(
		.INIT('h1)
	) name24828 (
		_w28787_,
		_w28874_,
		_w28875_
	);
	LUT2 #(
		.INIT('h4)
	) name24829 (
		\sport0_cfg_SP_ENg_D1_reg/P0001 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w28876_
	);
	LUT2 #(
		.INIT('h8)
	) name24830 (
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w28876_,
		_w28877_
	);
	LUT2 #(
		.INIT('h1)
	) name24831 (
		\IRFS0_pad ,
		\ITFS0_pad ,
		_w28878_
	);
	LUT2 #(
		.INIT('h2)
	) name24832 (
		\sport0_cfg_FSi_cnt_reg[8]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w28879_
	);
	LUT2 #(
		.INIT('h4)
	) name24833 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w28880_
	);
	LUT2 #(
		.INIT('h4)
	) name24834 (
		\sport0_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w28881_
	);
	LUT2 #(
		.INIT('h2)
	) name24835 (
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w28882_
	);
	LUT2 #(
		.INIT('h2)
	) name24836 (
		\sport0_cfg_FSi_cnt_reg[5]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w28883_
	);
	LUT2 #(
		.INIT('h4)
	) name24837 (
		\sport0_cfg_FSi_cnt_reg[8]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w28884_
	);
	LUT2 #(
		.INIT('h4)
	) name24838 (
		\sport0_cfg_FSi_cnt_reg[5]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w28885_
	);
	LUT2 #(
		.INIT('h4)
	) name24839 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w28886_
	);
	LUT2 #(
		.INIT('h4)
	) name24840 (
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w28887_
	);
	LUT2 #(
		.INIT('h4)
	) name24841 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w28888_
	);
	LUT2 #(
		.INIT('h2)
	) name24842 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w28889_
	);
	LUT2 #(
		.INIT('h4)
	) name24843 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w28890_
	);
	LUT2 #(
		.INIT('h4)
	) name24844 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w28891_
	);
	LUT2 #(
		.INIT('h4)
	) name24845 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w28892_
	);
	LUT2 #(
		.INIT('h2)
	) name24846 (
		\sport0_cfg_FSi_cnt_reg[15]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w28893_
	);
	LUT2 #(
		.INIT('h2)
	) name24847 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w28894_
	);
	LUT2 #(
		.INIT('h2)
	) name24848 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w28895_
	);
	LUT2 #(
		.INIT('h2)
	) name24849 (
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w28896_
	);
	LUT2 #(
		.INIT('h2)
	) name24850 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w28897_
	);
	LUT2 #(
		.INIT('h2)
	) name24851 (
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w28898_
	);
	LUT2 #(
		.INIT('h2)
	) name24852 (
		\sport0_cfg_FSi_cnt_reg[11]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w28899_
	);
	LUT2 #(
		.INIT('h2)
	) name24853 (
		\sport0_cfg_FSi_cnt_reg[14]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w28900_
	);
	LUT2 #(
		.INIT('h4)
	) name24854 (
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w28901_
	);
	LUT2 #(
		.INIT('h2)
	) name24855 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w28902_
	);
	LUT2 #(
		.INIT('h4)
	) name24856 (
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w28903_
	);
	LUT2 #(
		.INIT('h4)
	) name24857 (
		\sport0_cfg_FSi_cnt_reg[14]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w28904_
	);
	LUT2 #(
		.INIT('h4)
	) name24858 (
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w28905_
	);
	LUT2 #(
		.INIT('h2)
	) name24859 (
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w28906_
	);
	LUT2 #(
		.INIT('h2)
	) name24860 (
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w28907_
	);
	LUT2 #(
		.INIT('h4)
	) name24861 (
		\sport0_cfg_FSi_cnt_reg[15]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w28908_
	);
	LUT2 #(
		.INIT('h2)
	) name24862 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w28909_
	);
	LUT2 #(
		.INIT('h4)
	) name24863 (
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w28910_
	);
	LUT2 #(
		.INIT('h1)
	) name24864 (
		_w28879_,
		_w28880_,
		_w28911_
	);
	LUT2 #(
		.INIT('h1)
	) name24865 (
		_w28881_,
		_w28882_,
		_w28912_
	);
	LUT2 #(
		.INIT('h1)
	) name24866 (
		_w28883_,
		_w28884_,
		_w28913_
	);
	LUT2 #(
		.INIT('h1)
	) name24867 (
		_w28885_,
		_w28886_,
		_w28914_
	);
	LUT2 #(
		.INIT('h1)
	) name24868 (
		_w28887_,
		_w28888_,
		_w28915_
	);
	LUT2 #(
		.INIT('h1)
	) name24869 (
		_w28889_,
		_w28890_,
		_w28916_
	);
	LUT2 #(
		.INIT('h1)
	) name24870 (
		_w28891_,
		_w28892_,
		_w28917_
	);
	LUT2 #(
		.INIT('h1)
	) name24871 (
		_w28893_,
		_w28894_,
		_w28918_
	);
	LUT2 #(
		.INIT('h1)
	) name24872 (
		_w28895_,
		_w28896_,
		_w28919_
	);
	LUT2 #(
		.INIT('h1)
	) name24873 (
		_w28897_,
		_w28898_,
		_w28920_
	);
	LUT2 #(
		.INIT('h1)
	) name24874 (
		_w28899_,
		_w28900_,
		_w28921_
	);
	LUT2 #(
		.INIT('h1)
	) name24875 (
		_w28901_,
		_w28902_,
		_w28922_
	);
	LUT2 #(
		.INIT('h1)
	) name24876 (
		_w28903_,
		_w28904_,
		_w28923_
	);
	LUT2 #(
		.INIT('h1)
	) name24877 (
		_w28905_,
		_w28906_,
		_w28924_
	);
	LUT2 #(
		.INIT('h1)
	) name24878 (
		_w28907_,
		_w28908_,
		_w28925_
	);
	LUT2 #(
		.INIT('h1)
	) name24879 (
		_w28909_,
		_w28910_,
		_w28926_
	);
	LUT2 #(
		.INIT('h8)
	) name24880 (
		_w28925_,
		_w28926_,
		_w28927_
	);
	LUT2 #(
		.INIT('h8)
	) name24881 (
		_w28923_,
		_w28924_,
		_w28928_
	);
	LUT2 #(
		.INIT('h8)
	) name24882 (
		_w28921_,
		_w28922_,
		_w28929_
	);
	LUT2 #(
		.INIT('h8)
	) name24883 (
		_w28919_,
		_w28920_,
		_w28930_
	);
	LUT2 #(
		.INIT('h8)
	) name24884 (
		_w28917_,
		_w28918_,
		_w28931_
	);
	LUT2 #(
		.INIT('h8)
	) name24885 (
		_w28915_,
		_w28916_,
		_w28932_
	);
	LUT2 #(
		.INIT('h8)
	) name24886 (
		_w28913_,
		_w28914_,
		_w28933_
	);
	LUT2 #(
		.INIT('h8)
	) name24887 (
		_w28911_,
		_w28912_,
		_w28934_
	);
	LUT2 #(
		.INIT('h8)
	) name24888 (
		_w28933_,
		_w28934_,
		_w28935_
	);
	LUT2 #(
		.INIT('h8)
	) name24889 (
		_w28931_,
		_w28932_,
		_w28936_
	);
	LUT2 #(
		.INIT('h8)
	) name24890 (
		_w28929_,
		_w28930_,
		_w28937_
	);
	LUT2 #(
		.INIT('h8)
	) name24891 (
		_w28927_,
		_w28928_,
		_w28938_
	);
	LUT2 #(
		.INIT('h8)
	) name24892 (
		_w28937_,
		_w28938_,
		_w28939_
	);
	LUT2 #(
		.INIT('h8)
	) name24893 (
		_w28935_,
		_w28936_,
		_w28940_
	);
	LUT2 #(
		.INIT('h8)
	) name24894 (
		_w28939_,
		_w28940_,
		_w28941_
	);
	LUT2 #(
		.INIT('h1)
	) name24895 (
		_w28878_,
		_w28941_,
		_w28942_
	);
	LUT2 #(
		.INIT('h8)
	) name24896 (
		\memc_usysr_DO_reg[12]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w28943_
	);
	LUT2 #(
		.INIT('h4)
	) name24897 (
		_w28942_,
		_w28943_,
		_w28944_
	);
	LUT2 #(
		.INIT('h1)
	) name24898 (
		_w28876_,
		_w28944_,
		_w28945_
	);
	LUT2 #(
		.INIT('h8)
	) name24899 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w28946_
	);
	LUT2 #(
		.INIT('h8)
	) name24900 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		_w28946_,
		_w28947_
	);
	LUT2 #(
		.INIT('h8)
	) name24901 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		_w28947_,
		_w28948_
	);
	LUT2 #(
		.INIT('h8)
	) name24902 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		_w28948_,
		_w28949_
	);
	LUT2 #(
		.INIT('h8)
	) name24903 (
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		_w28949_,
		_w28950_
	);
	LUT2 #(
		.INIT('h8)
	) name24904 (
		\sport0_cfg_FSi_cnt_reg[5]/NET0131 ,
		_w28950_,
		_w28951_
	);
	LUT2 #(
		.INIT('h8)
	) name24905 (
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		_w28951_,
		_w28952_
	);
	LUT2 #(
		.INIT('h8)
	) name24906 (
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		_w28952_,
		_w28953_
	);
	LUT2 #(
		.INIT('h8)
	) name24907 (
		\sport0_cfg_FSi_cnt_reg[8]/NET0131 ,
		_w28953_,
		_w28954_
	);
	LUT2 #(
		.INIT('h8)
	) name24908 (
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w28954_,
		_w28955_
	);
	LUT2 #(
		.INIT('h8)
	) name24909 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		_w28955_,
		_w28956_
	);
	LUT2 #(
		.INIT('h8)
	) name24910 (
		\sport0_cfg_FSi_cnt_reg[11]/NET0131 ,
		_w28956_,
		_w28957_
	);
	LUT2 #(
		.INIT('h8)
	) name24911 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		_w28957_,
		_w28958_
	);
	LUT2 #(
		.INIT('h8)
	) name24912 (
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		_w28958_,
		_w28959_
	);
	LUT2 #(
		.INIT('h8)
	) name24913 (
		\sport0_cfg_FSi_cnt_reg[14]/NET0131 ,
		_w28959_,
		_w28960_
	);
	LUT2 #(
		.INIT('h1)
	) name24914 (
		\sport0_cfg_FSi_cnt_reg[15]/NET0131 ,
		_w28960_,
		_w28961_
	);
	LUT2 #(
		.INIT('h8)
	) name24915 (
		\sport0_cfg_FSi_cnt_reg[15]/NET0131 ,
		_w28960_,
		_w28962_
	);
	LUT2 #(
		.INIT('h2)
	) name24916 (
		_w28945_,
		_w28961_,
		_w28963_
	);
	LUT2 #(
		.INIT('h4)
	) name24917 (
		_w28962_,
		_w28963_,
		_w28964_
	);
	LUT2 #(
		.INIT('h1)
	) name24918 (
		_w28877_,
		_w28964_,
		_w28965_
	);
	LUT2 #(
		.INIT('h2)
	) name24919 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 ,
		_w18266_,
		_w28966_
	);
	LUT2 #(
		.INIT('h1)
	) name24920 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[13]/P0001 ,
		_w18271_,
		_w28967_
	);
	LUT2 #(
		.INIT('h4)
	) name24921 (
		_w17836_,
		_w18271_,
		_w28968_
	);
	LUT2 #(
		.INIT('h2)
	) name24922 (
		_w18273_,
		_w28967_,
		_w28969_
	);
	LUT2 #(
		.INIT('h4)
	) name24923 (
		_w28968_,
		_w28969_,
		_w28970_
	);
	LUT2 #(
		.INIT('h1)
	) name24924 (
		_w18270_,
		_w28966_,
		_w28971_
	);
	LUT2 #(
		.INIT('h4)
	) name24925 (
		_w28970_,
		_w28971_,
		_w28972_
	);
	LUT2 #(
		.INIT('h1)
	) name24926 (
		_w18262_,
		_w28972_,
		_w28973_
	);
	LUT2 #(
		.INIT('h2)
	) name24927 (
		_w18262_,
		_w19636_,
		_w28974_
	);
	LUT2 #(
		.INIT('h1)
	) name24928 (
		_w28973_,
		_w28974_,
		_w28975_
	);
	LUT2 #(
		.INIT('h8)
	) name24929 (
		_w14752_,
		_w19636_,
		_w28976_
	);
	LUT2 #(
		.INIT('h8)
	) name24930 (
		_w17836_,
		_w18328_,
		_w28977_
	);
	LUT2 #(
		.INIT('h2)
	) name24931 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[13]/P0001 ,
		_w18330_,
		_w28978_
	);
	LUT2 #(
		.INIT('h2)
	) name24932 (
		_w18334_,
		_w28978_,
		_w28979_
	);
	LUT2 #(
		.INIT('h4)
	) name24933 (
		_w28977_,
		_w28979_,
		_w28980_
	);
	LUT2 #(
		.INIT('h1)
	) name24934 (
		_w28976_,
		_w28980_,
		_w28981_
	);
	LUT2 #(
		.INIT('h4)
	) name24935 (
		_w26301_,
		_w26333_,
		_w28982_
	);
	LUT2 #(
		.INIT('h2)
	) name24936 (
		\sport1_txctl_TXSHT_reg[11]/P0001 ,
		_w22677_,
		_w28983_
	);
	LUT2 #(
		.INIT('h8)
	) name24937 (
		\sport1_txctl_TX_reg[12]/P0001 ,
		_w22677_,
		_w28984_
	);
	LUT2 #(
		.INIT('h1)
	) name24938 (
		_w28983_,
		_w28984_,
		_w28985_
	);
	LUT2 #(
		.INIT('h1)
	) name24939 (
		_w11311_,
		_w28556_,
		_w28986_
	);
	LUT2 #(
		.INIT('h8)
	) name24940 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w18276_,
		_w28987_
	);
	LUT2 #(
		.INIT('h4)
	) name24941 (
		_w14623_,
		_w28561_,
		_w28988_
	);
	LUT2 #(
		.INIT('h1)
	) name24942 (
		_w28564_,
		_w28987_,
		_w28989_
	);
	LUT2 #(
		.INIT('h4)
	) name24943 (
		_w28988_,
		_w28989_,
		_w28990_
	);
	LUT2 #(
		.INIT('h2)
	) name24944 (
		_w28559_,
		_w28990_,
		_w28991_
	);
	LUT2 #(
		.INIT('h2)
	) name24945 (
		_w28572_,
		_w28574_,
		_w28992_
	);
	LUT2 #(
		.INIT('h8)
	) name24946 (
		_w12972_,
		_w28992_,
		_w28993_
	);
	LUT2 #(
		.INIT('h1)
	) name24947 (
		_w28576_,
		_w28993_,
		_w28994_
	);
	LUT2 #(
		.INIT('h2)
	) name24948 (
		_w28569_,
		_w28994_,
		_w28995_
	);
	LUT2 #(
		.INIT('h1)
	) name24949 (
		_w12972_,
		_w28572_,
		_w28996_
	);
	LUT2 #(
		.INIT('h8)
	) name24950 (
		_w28569_,
		_w28574_,
		_w28997_
	);
	LUT2 #(
		.INIT('h4)
	) name24951 (
		_w11525_,
		_w28572_,
		_w28998_
	);
	LUT2 #(
		.INIT('h4)
	) name24952 (
		_w28996_,
		_w28997_,
		_w28999_
	);
	LUT2 #(
		.INIT('h4)
	) name24953 (
		_w28998_,
		_w28999_,
		_w29000_
	);
	LUT2 #(
		.INIT('h1)
	) name24954 (
		_w11341_,
		_w28634_,
		_w29001_
	);
	LUT2 #(
		.INIT('h4)
	) name24955 (
		_w18940_,
		_w28636_,
		_w29002_
	);
	LUT2 #(
		.INIT('h8)
	) name24956 (
		_w11525_,
		_w28630_,
		_w29003_
	);
	LUT2 #(
		.INIT('h1)
	) name24957 (
		_w11315_,
		_w28624_,
		_w29004_
	);
	LUT2 #(
		.INIT('h8)
	) name24958 (
		_w12972_,
		_w28619_,
		_w29005_
	);
	LUT2 #(
		.INIT('h4)
	) name24959 (
		_w18831_,
		_w28627_,
		_w29006_
	);
	LUT2 #(
		.INIT('h1)
	) name24960 (
		_w11525_,
		_w28572_,
		_w29007_
	);
	LUT2 #(
		.INIT('h1)
	) name24961 (
		_w11444_,
		_w28594_,
		_w29008_
	);
	LUT2 #(
		.INIT('h1)
	) name24962 (
		_w11448_,
		_w28589_,
		_w29009_
	);
	LUT2 #(
		.INIT('h1)
	) name24963 (
		_w11424_,
		_w28598_,
		_w29010_
	);
	LUT2 #(
		.INIT('h1)
	) name24964 (
		_w29008_,
		_w29009_,
		_w29011_
	);
	LUT2 #(
		.INIT('h4)
	) name24965 (
		_w29010_,
		_w29011_,
		_w29012_
	);
	LUT2 #(
		.INIT('h8)
	) name24966 (
		_w28607_,
		_w29012_,
		_w29013_
	);
	LUT2 #(
		.INIT('h8)
	) name24967 (
		_w28572_,
		_w29013_,
		_w29014_
	);
	LUT2 #(
		.INIT('h2)
	) name24968 (
		_w28584_,
		_w29007_,
		_w29015_
	);
	LUT2 #(
		.INIT('h4)
	) name24969 (
		_w29014_,
		_w29015_,
		_w29016_
	);
	LUT2 #(
		.INIT('h1)
	) name24970 (
		_w29001_,
		_w29003_,
		_w29017_
	);
	LUT2 #(
		.INIT('h4)
	) name24971 (
		_w29005_,
		_w29017_,
		_w29018_
	);
	LUT2 #(
		.INIT('h1)
	) name24972 (
		_w28986_,
		_w29002_,
		_w29019_
	);
	LUT2 #(
		.INIT('h4)
	) name24973 (
		_w29004_,
		_w29019_,
		_w29020_
	);
	LUT2 #(
		.INIT('h4)
	) name24974 (
		_w29006_,
		_w29018_,
		_w29021_
	);
	LUT2 #(
		.INIT('h8)
	) name24975 (
		_w29020_,
		_w29021_,
		_w29022_
	);
	LUT2 #(
		.INIT('h4)
	) name24976 (
		_w29000_,
		_w29022_,
		_w29023_
	);
	LUT2 #(
		.INIT('h4)
	) name24977 (
		_w29016_,
		_w29023_,
		_w29024_
	);
	LUT2 #(
		.INIT('h4)
	) name24978 (
		_w28995_,
		_w29024_,
		_w29025_
	);
	LUT2 #(
		.INIT('h4)
	) name24979 (
		_w28991_,
		_w29025_,
		_w29026_
	);
	LUT2 #(
		.INIT('h2)
	) name24980 (
		_w28550_,
		_w29026_,
		_w29027_
	);
	LUT2 #(
		.INIT('h4)
	) name24981 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[6]/P0001 ,
		_w28649_,
		_w29028_
	);
	LUT2 #(
		.INIT('h8)
	) name24982 (
		_w11440_,
		_w28652_,
		_w29029_
	);
	LUT2 #(
		.INIT('h2)
	) name24983 (
		_w11428_,
		_w28652_,
		_w29030_
	);
	LUT2 #(
		.INIT('h1)
	) name24984 (
		_w28660_,
		_w29029_,
		_w29031_
	);
	LUT2 #(
		.INIT('h4)
	) name24985 (
		_w29030_,
		_w29031_,
		_w29032_
	);
	LUT2 #(
		.INIT('h8)
	) name24986 (
		_w18276_,
		_w28660_,
		_w29033_
	);
	LUT2 #(
		.INIT('h1)
	) name24987 (
		_w28649_,
		_w29032_,
		_w29034_
	);
	LUT2 #(
		.INIT('h4)
	) name24988 (
		_w29033_,
		_w29034_,
		_w29035_
	);
	LUT2 #(
		.INIT('h1)
	) name24989 (
		_w28550_,
		_w29028_,
		_w29036_
	);
	LUT2 #(
		.INIT('h4)
	) name24990 (
		_w29035_,
		_w29036_,
		_w29037_
	);
	LUT2 #(
		.INIT('h1)
	) name24991 (
		_w29027_,
		_w29037_,
		_w29038_
	);
	LUT2 #(
		.INIT('h4)
	) name24992 (
		_w14634_,
		_w28561_,
		_w29039_
	);
	LUT2 #(
		.INIT('h8)
	) name24993 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w20259_,
		_w29040_
	);
	LUT2 #(
		.INIT('h1)
	) name24994 (
		_w28564_,
		_w29040_,
		_w29041_
	);
	LUT2 #(
		.INIT('h4)
	) name24995 (
		_w29039_,
		_w29041_,
		_w29042_
	);
	LUT2 #(
		.INIT('h2)
	) name24996 (
		_w28559_,
		_w29042_,
		_w29043_
	);
	LUT2 #(
		.INIT('h1)
	) name24997 (
		_w10801_,
		_w28624_,
		_w29044_
	);
	LUT2 #(
		.INIT('h1)
	) name24998 (
		_w10694_,
		_w28634_,
		_w29045_
	);
	LUT2 #(
		.INIT('h2)
	) name24999 (
		_w18088_,
		_w18895_,
		_w29046_
	);
	LUT2 #(
		.INIT('h4)
	) name25000 (
		_w18002_,
		_w20107_,
		_w29047_
	);
	LUT2 #(
		.INIT('h2)
	) name25001 (
		_w17925_,
		_w19818_,
		_w29048_
	);
	LUT2 #(
		.INIT('h1)
	) name25002 (
		_w18069_,
		_w19787_,
		_w29049_
	);
	LUT2 #(
		.INIT('h1)
	) name25003 (
		_w18091_,
		_w18189_,
		_w29050_
	);
	LUT2 #(
		.INIT('h4)
	) name25004 (
		_w18114_,
		_w18719_,
		_w29051_
	);
	LUT2 #(
		.INIT('h8)
	) name25005 (
		_w17978_,
		_w20084_,
		_w29052_
	);
	LUT2 #(
		.INIT('h2)
	) name25006 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w10797_,
		_w29053_
	);
	LUT2 #(
		.INIT('h8)
	) name25007 (
		_w17934_,
		_w18055_,
		_w29054_
	);
	LUT2 #(
		.INIT('h2)
	) name25008 (
		_w18111_,
		_w19857_,
		_w29055_
	);
	LUT2 #(
		.INIT('h1)
	) name25009 (
		_w18104_,
		_w18133_,
		_w29056_
	);
	LUT2 #(
		.INIT('h1)
	) name25010 (
		_w17922_,
		_w18167_,
		_w29057_
	);
	LUT2 #(
		.INIT('h1)
	) name25011 (
		_w18108_,
		_w18129_,
		_w29058_
	);
	LUT2 #(
		.INIT('h8)
	) name25012 (
		_w18071_,
		_w18748_,
		_w29059_
	);
	LUT2 #(
		.INIT('h2)
	) name25013 (
		_w18765_,
		_w18781_,
		_w29060_
	);
	LUT2 #(
		.INIT('h2)
	) name25014 (
		_w18171_,
		_w19979_,
		_w29061_
	);
	LUT2 #(
		.INIT('h1)
	) name25015 (
		_w18135_,
		_w18149_,
		_w29062_
	);
	LUT2 #(
		.INIT('h1)
	) name25016 (
		_w17981_,
		_w18046_,
		_w29063_
	);
	LUT2 #(
		.INIT('h2)
	) name25017 (
		_w18115_,
		_w29063_,
		_w29064_
	);
	LUT2 #(
		.INIT('h1)
	) name25018 (
		_w18192_,
		_w29053_,
		_w29065_
	);
	LUT2 #(
		.INIT('h4)
	) name25019 (
		_w29054_,
		_w29065_,
		_w29066_
	);
	LUT2 #(
		.INIT('h4)
	) name25020 (
		_w29051_,
		_w29066_,
		_w29067_
	);
	LUT2 #(
		.INIT('h1)
	) name25021 (
		_w29050_,
		_w29056_,
		_w29068_
	);
	LUT2 #(
		.INIT('h1)
	) name25022 (
		_w29057_,
		_w29058_,
		_w29069_
	);
	LUT2 #(
		.INIT('h4)
	) name25023 (
		_w29059_,
		_w29069_,
		_w29070_
	);
	LUT2 #(
		.INIT('h8)
	) name25024 (
		_w29067_,
		_w29068_,
		_w29071_
	);
	LUT2 #(
		.INIT('h2)
	) name25025 (
		_w18041_,
		_w29046_,
		_w29072_
	);
	LUT2 #(
		.INIT('h4)
	) name25026 (
		_w29048_,
		_w29049_,
		_w29073_
	);
	LUT2 #(
		.INIT('h2)
	) name25027 (
		_w29052_,
		_w29055_,
		_w29074_
	);
	LUT2 #(
		.INIT('h1)
	) name25028 (
		_w29060_,
		_w29061_,
		_w29075_
	);
	LUT2 #(
		.INIT('h1)
	) name25029 (
		_w29062_,
		_w29064_,
		_w29076_
	);
	LUT2 #(
		.INIT('h8)
	) name25030 (
		_w29075_,
		_w29076_,
		_w29077_
	);
	LUT2 #(
		.INIT('h8)
	) name25031 (
		_w29073_,
		_w29074_,
		_w29078_
	);
	LUT2 #(
		.INIT('h8)
	) name25032 (
		_w29071_,
		_w29072_,
		_w29079_
	);
	LUT2 #(
		.INIT('h8)
	) name25033 (
		_w29070_,
		_w29079_,
		_w29080_
	);
	LUT2 #(
		.INIT('h8)
	) name25034 (
		_w29077_,
		_w29078_,
		_w29081_
	);
	LUT2 #(
		.INIT('h8)
	) name25035 (
		_w18726_,
		_w29081_,
		_w29082_
	);
	LUT2 #(
		.INIT('h8)
	) name25036 (
		_w29080_,
		_w29082_,
		_w29083_
	);
	LUT2 #(
		.INIT('h8)
	) name25037 (
		_w18800_,
		_w29083_,
		_w29084_
	);
	LUT2 #(
		.INIT('h8)
	) name25038 (
		_w29047_,
		_w29084_,
		_w29085_
	);
	LUT2 #(
		.INIT('h2)
	) name25039 (
		_w28627_,
		_w29085_,
		_w29086_
	);
	LUT2 #(
		.INIT('h1)
	) name25040 (
		_w10797_,
		_w28556_,
		_w29087_
	);
	LUT2 #(
		.INIT('h4)
	) name25041 (
		_w20288_,
		_w28636_,
		_w29088_
	);
	LUT2 #(
		.INIT('h1)
	) name25042 (
		_w12938_,
		_w28577_,
		_w29089_
	);
	LUT2 #(
		.INIT('h4)
	) name25043 (
		_w10911_,
		_w28577_,
		_w29090_
	);
	LUT2 #(
		.INIT('h1)
	) name25044 (
		_w28575_,
		_w29089_,
		_w29091_
	);
	LUT2 #(
		.INIT('h4)
	) name25045 (
		_w29090_,
		_w29091_,
		_w29092_
	);
	LUT2 #(
		.INIT('h1)
	) name25046 (
		_w28576_,
		_w29092_,
		_w29093_
	);
	LUT2 #(
		.INIT('h2)
	) name25047 (
		_w28569_,
		_w29093_,
		_w29094_
	);
	LUT2 #(
		.INIT('h8)
	) name25048 (
		_w10911_,
		_w28630_,
		_w29095_
	);
	LUT2 #(
		.INIT('h8)
	) name25049 (
		_w12938_,
		_w28619_,
		_w29096_
	);
	LUT2 #(
		.INIT('h1)
	) name25050 (
		_w10911_,
		_w28572_,
		_w29097_
	);
	LUT2 #(
		.INIT('h1)
	) name25051 (
		_w10882_,
		_w28598_,
		_w29098_
	);
	LUT2 #(
		.INIT('h1)
	) name25052 (
		_w10858_,
		_w28589_,
		_w29099_
	);
	LUT2 #(
		.INIT('h1)
	) name25053 (
		_w10878_,
		_w28594_,
		_w29100_
	);
	LUT2 #(
		.INIT('h1)
	) name25054 (
		_w29098_,
		_w29099_,
		_w29101_
	);
	LUT2 #(
		.INIT('h4)
	) name25055 (
		_w29100_,
		_w29101_,
		_w29102_
	);
	LUT2 #(
		.INIT('h8)
	) name25056 (
		_w28607_,
		_w29102_,
		_w29103_
	);
	LUT2 #(
		.INIT('h8)
	) name25057 (
		_w28572_,
		_w29103_,
		_w29104_
	);
	LUT2 #(
		.INIT('h2)
	) name25058 (
		_w28584_,
		_w29097_,
		_w29105_
	);
	LUT2 #(
		.INIT('h4)
	) name25059 (
		_w29104_,
		_w29105_,
		_w29106_
	);
	LUT2 #(
		.INIT('h1)
	) name25060 (
		_w29045_,
		_w29095_,
		_w29107_
	);
	LUT2 #(
		.INIT('h4)
	) name25061 (
		_w29096_,
		_w29107_,
		_w29108_
	);
	LUT2 #(
		.INIT('h1)
	) name25062 (
		_w29044_,
		_w29087_,
		_w29109_
	);
	LUT2 #(
		.INIT('h4)
	) name25063 (
		_w29088_,
		_w29109_,
		_w29110_
	);
	LUT2 #(
		.INIT('h8)
	) name25064 (
		_w29108_,
		_w29110_,
		_w29111_
	);
	LUT2 #(
		.INIT('h4)
	) name25065 (
		_w29086_,
		_w29111_,
		_w29112_
	);
	LUT2 #(
		.INIT('h4)
	) name25066 (
		_w29106_,
		_w29112_,
		_w29113_
	);
	LUT2 #(
		.INIT('h4)
	) name25067 (
		_w29094_,
		_w29113_,
		_w29114_
	);
	LUT2 #(
		.INIT('h4)
	) name25068 (
		_w29043_,
		_w29114_,
		_w29115_
	);
	LUT2 #(
		.INIT('h2)
	) name25069 (
		_w28550_,
		_w29115_,
		_w29116_
	);
	LUT2 #(
		.INIT('h4)
	) name25070 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[5]/P0001 ,
		_w28649_,
		_w29117_
	);
	LUT2 #(
		.INIT('h8)
	) name25071 (
		_w10874_,
		_w28652_,
		_w29118_
	);
	LUT2 #(
		.INIT('h2)
	) name25072 (
		_w10866_,
		_w28652_,
		_w29119_
	);
	LUT2 #(
		.INIT('h1)
	) name25073 (
		_w28660_,
		_w29118_,
		_w29120_
	);
	LUT2 #(
		.INIT('h4)
	) name25074 (
		_w29119_,
		_w29120_,
		_w29121_
	);
	LUT2 #(
		.INIT('h8)
	) name25075 (
		_w20259_,
		_w28660_,
		_w29122_
	);
	LUT2 #(
		.INIT('h1)
	) name25076 (
		_w28649_,
		_w29121_,
		_w29123_
	);
	LUT2 #(
		.INIT('h4)
	) name25077 (
		_w29122_,
		_w29123_,
		_w29124_
	);
	LUT2 #(
		.INIT('h1)
	) name25078 (
		_w28550_,
		_w29117_,
		_w29125_
	);
	LUT2 #(
		.INIT('h4)
	) name25079 (
		_w29124_,
		_w29125_,
		_w29126_
	);
	LUT2 #(
		.INIT('h1)
	) name25080 (
		_w29116_,
		_w29126_,
		_w29127_
	);
	LUT2 #(
		.INIT('h4)
	) name25081 (
		_w20142_,
		_w28627_,
		_w29128_
	);
	LUT2 #(
		.INIT('h8)
	) name25082 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w20080_,
		_w29129_
	);
	LUT2 #(
		.INIT('h4)
	) name25083 (
		_w14600_,
		_w28561_,
		_w29130_
	);
	LUT2 #(
		.INIT('h1)
	) name25084 (
		_w28564_,
		_w29129_,
		_w29131_
	);
	LUT2 #(
		.INIT('h4)
	) name25085 (
		_w29130_,
		_w29131_,
		_w29132_
	);
	LUT2 #(
		.INIT('h2)
	) name25086 (
		_w28559_,
		_w29132_,
		_w29133_
	);
	LUT2 #(
		.INIT('h8)
	) name25087 (
		_w12904_,
		_w28992_,
		_w29134_
	);
	LUT2 #(
		.INIT('h1)
	) name25088 (
		_w28576_,
		_w29134_,
		_w29135_
	);
	LUT2 #(
		.INIT('h2)
	) name25089 (
		_w28569_,
		_w29135_,
		_w29136_
	);
	LUT2 #(
		.INIT('h1)
	) name25090 (
		_w12904_,
		_w28572_,
		_w29137_
	);
	LUT2 #(
		.INIT('h4)
	) name25091 (
		_w10069_,
		_w28572_,
		_w29138_
	);
	LUT2 #(
		.INIT('h2)
	) name25092 (
		_w28997_,
		_w29137_,
		_w29139_
	);
	LUT2 #(
		.INIT('h4)
	) name25093 (
		_w29138_,
		_w29139_,
		_w29140_
	);
	LUT2 #(
		.INIT('h1)
	) name25094 (
		_w9947_,
		_w28556_,
		_w29141_
	);
	LUT2 #(
		.INIT('h1)
	) name25095 (
		_w9912_,
		_w28634_,
		_w29142_
	);
	LUT2 #(
		.INIT('h4)
	) name25096 (
		_w22911_,
		_w28636_,
		_w29143_
	);
	LUT2 #(
		.INIT('h8)
	) name25097 (
		_w10069_,
		_w28630_,
		_w29144_
	);
	LUT2 #(
		.INIT('h8)
	) name25098 (
		_w12904_,
		_w28619_,
		_w29145_
	);
	LUT2 #(
		.INIT('h1)
	) name25099 (
		_w9951_,
		_w28624_,
		_w29146_
	);
	LUT2 #(
		.INIT('h1)
	) name25100 (
		_w10069_,
		_w28572_,
		_w29147_
	);
	LUT2 #(
		.INIT('h1)
	) name25101 (
		_w9845_,
		_w28589_,
		_w29148_
	);
	LUT2 #(
		.INIT('h1)
	) name25102 (
		_w9869_,
		_w28594_,
		_w29149_
	);
	LUT2 #(
		.INIT('h1)
	) name25103 (
		_w9865_,
		_w28598_,
		_w29150_
	);
	LUT2 #(
		.INIT('h1)
	) name25104 (
		_w29148_,
		_w29149_,
		_w29151_
	);
	LUT2 #(
		.INIT('h4)
	) name25105 (
		_w29150_,
		_w29151_,
		_w29152_
	);
	LUT2 #(
		.INIT('h8)
	) name25106 (
		_w28607_,
		_w29152_,
		_w29153_
	);
	LUT2 #(
		.INIT('h8)
	) name25107 (
		_w28572_,
		_w29153_,
		_w29154_
	);
	LUT2 #(
		.INIT('h2)
	) name25108 (
		_w28584_,
		_w29147_,
		_w29155_
	);
	LUT2 #(
		.INIT('h4)
	) name25109 (
		_w29154_,
		_w29155_,
		_w29156_
	);
	LUT2 #(
		.INIT('h1)
	) name25110 (
		_w29142_,
		_w29144_,
		_w29157_
	);
	LUT2 #(
		.INIT('h4)
	) name25111 (
		_w29145_,
		_w29157_,
		_w29158_
	);
	LUT2 #(
		.INIT('h1)
	) name25112 (
		_w29141_,
		_w29143_,
		_w29159_
	);
	LUT2 #(
		.INIT('h4)
	) name25113 (
		_w29146_,
		_w29159_,
		_w29160_
	);
	LUT2 #(
		.INIT('h4)
	) name25114 (
		_w29128_,
		_w29158_,
		_w29161_
	);
	LUT2 #(
		.INIT('h8)
	) name25115 (
		_w29160_,
		_w29161_,
		_w29162_
	);
	LUT2 #(
		.INIT('h4)
	) name25116 (
		_w29140_,
		_w29162_,
		_w29163_
	);
	LUT2 #(
		.INIT('h4)
	) name25117 (
		_w29156_,
		_w29163_,
		_w29164_
	);
	LUT2 #(
		.INIT('h4)
	) name25118 (
		_w29136_,
		_w29164_,
		_w29165_
	);
	LUT2 #(
		.INIT('h4)
	) name25119 (
		_w29133_,
		_w29165_,
		_w29166_
	);
	LUT2 #(
		.INIT('h2)
	) name25120 (
		_w28550_,
		_w29166_,
		_w29167_
	);
	LUT2 #(
		.INIT('h4)
	) name25121 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[4]/P0001 ,
		_w28649_,
		_w29168_
	);
	LUT2 #(
		.INIT('h8)
	) name25122 (
		_w9861_,
		_w28652_,
		_w29169_
	);
	LUT2 #(
		.INIT('h2)
	) name25123 (
		_w9849_,
		_w28652_,
		_w29170_
	);
	LUT2 #(
		.INIT('h1)
	) name25124 (
		_w28660_,
		_w29169_,
		_w29171_
	);
	LUT2 #(
		.INIT('h4)
	) name25125 (
		_w29170_,
		_w29171_,
		_w29172_
	);
	LUT2 #(
		.INIT('h8)
	) name25126 (
		_w20080_,
		_w28660_,
		_w29173_
	);
	LUT2 #(
		.INIT('h1)
	) name25127 (
		_w28649_,
		_w29172_,
		_w29174_
	);
	LUT2 #(
		.INIT('h4)
	) name25128 (
		_w29173_,
		_w29174_,
		_w29175_
	);
	LUT2 #(
		.INIT('h1)
	) name25129 (
		_w28550_,
		_w29168_,
		_w29176_
	);
	LUT2 #(
		.INIT('h4)
	) name25130 (
		_w29175_,
		_w29176_,
		_w29177_
	);
	LUT2 #(
		.INIT('h1)
	) name25131 (
		_w29167_,
		_w29177_,
		_w29178_
	);
	LUT2 #(
		.INIT('h1)
	) name25132 (
		_w9280_,
		_w28556_,
		_w29179_
	);
	LUT2 #(
		.INIT('h8)
	) name25133 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w18974_,
		_w29180_
	);
	LUT2 #(
		.INIT('h8)
	) name25134 (
		_w14573_,
		_w28561_,
		_w29181_
	);
	LUT2 #(
		.INIT('h1)
	) name25135 (
		_w28564_,
		_w29180_,
		_w29182_
	);
	LUT2 #(
		.INIT('h4)
	) name25136 (
		_w29181_,
		_w29182_,
		_w29183_
	);
	LUT2 #(
		.INIT('h2)
	) name25137 (
		_w28559_,
		_w29183_,
		_w29184_
	);
	LUT2 #(
		.INIT('h1)
	) name25138 (
		_w12802_,
		_w28577_,
		_w29185_
	);
	LUT2 #(
		.INIT('h4)
	) name25139 (
		_w9435_,
		_w28577_,
		_w29186_
	);
	LUT2 #(
		.INIT('h1)
	) name25140 (
		_w28575_,
		_w29185_,
		_w29187_
	);
	LUT2 #(
		.INIT('h4)
	) name25141 (
		_w29186_,
		_w29187_,
		_w29188_
	);
	LUT2 #(
		.INIT('h1)
	) name25142 (
		_w28576_,
		_w29188_,
		_w29189_
	);
	LUT2 #(
		.INIT('h2)
	) name25143 (
		_w28569_,
		_w29189_,
		_w29190_
	);
	LUT2 #(
		.INIT('h1)
	) name25144 (
		_w9276_,
		_w28624_,
		_w29191_
	);
	LUT2 #(
		.INIT('h4)
	) name25145 (
		_w21046_,
		_w28627_,
		_w29192_
	);
	LUT2 #(
		.INIT('h1)
	) name25146 (
		_w9297_,
		_w28634_,
		_w29193_
	);
	LUT2 #(
		.INIT('h8)
	) name25147 (
		_w12802_,
		_w28619_,
		_w29194_
	);
	LUT2 #(
		.INIT('h8)
	) name25148 (
		_w9435_,
		_w28630_,
		_w29195_
	);
	LUT2 #(
		.INIT('h4)
	) name25149 (
		_w19008_,
		_w28636_,
		_w29196_
	);
	LUT2 #(
		.INIT('h1)
	) name25150 (
		_w9435_,
		_w28572_,
		_w29197_
	);
	LUT2 #(
		.INIT('h1)
	) name25151 (
		_w9225_,
		_w28594_,
		_w29198_
	);
	LUT2 #(
		.INIT('h1)
	) name25152 (
		_w9229_,
		_w28598_,
		_w29199_
	);
	LUT2 #(
		.INIT('h1)
	) name25153 (
		_w9205_,
		_w28589_,
		_w29200_
	);
	LUT2 #(
		.INIT('h1)
	) name25154 (
		_w29198_,
		_w29199_,
		_w29201_
	);
	LUT2 #(
		.INIT('h4)
	) name25155 (
		_w29200_,
		_w29201_,
		_w29202_
	);
	LUT2 #(
		.INIT('h8)
	) name25156 (
		_w28607_,
		_w29202_,
		_w29203_
	);
	LUT2 #(
		.INIT('h8)
	) name25157 (
		_w28572_,
		_w29203_,
		_w29204_
	);
	LUT2 #(
		.INIT('h2)
	) name25158 (
		_w28584_,
		_w29197_,
		_w29205_
	);
	LUT2 #(
		.INIT('h4)
	) name25159 (
		_w29204_,
		_w29205_,
		_w29206_
	);
	LUT2 #(
		.INIT('h1)
	) name25160 (
		_w29193_,
		_w29194_,
		_w29207_
	);
	LUT2 #(
		.INIT('h1)
	) name25161 (
		_w29195_,
		_w29196_,
		_w29208_
	);
	LUT2 #(
		.INIT('h8)
	) name25162 (
		_w29207_,
		_w29208_,
		_w29209_
	);
	LUT2 #(
		.INIT('h1)
	) name25163 (
		_w29179_,
		_w29191_,
		_w29210_
	);
	LUT2 #(
		.INIT('h8)
	) name25164 (
		_w29209_,
		_w29210_,
		_w29211_
	);
	LUT2 #(
		.INIT('h4)
	) name25165 (
		_w29192_,
		_w29211_,
		_w29212_
	);
	LUT2 #(
		.INIT('h4)
	) name25166 (
		_w29206_,
		_w29212_,
		_w29213_
	);
	LUT2 #(
		.INIT('h4)
	) name25167 (
		_w29190_,
		_w29213_,
		_w29214_
	);
	LUT2 #(
		.INIT('h4)
	) name25168 (
		_w29184_,
		_w29214_,
		_w29215_
	);
	LUT2 #(
		.INIT('h2)
	) name25169 (
		_w28550_,
		_w29215_,
		_w29216_
	);
	LUT2 #(
		.INIT('h4)
	) name25170 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[1]/P0001 ,
		_w28649_,
		_w29217_
	);
	LUT2 #(
		.INIT('h8)
	) name25171 (
		_w9221_,
		_w28652_,
		_w29218_
	);
	LUT2 #(
		.INIT('h2)
	) name25172 (
		_w9213_,
		_w28652_,
		_w29219_
	);
	LUT2 #(
		.INIT('h1)
	) name25173 (
		_w28660_,
		_w29218_,
		_w29220_
	);
	LUT2 #(
		.INIT('h4)
	) name25174 (
		_w29219_,
		_w29220_,
		_w29221_
	);
	LUT2 #(
		.INIT('h8)
	) name25175 (
		_w18974_,
		_w28660_,
		_w29222_
	);
	LUT2 #(
		.INIT('h1)
	) name25176 (
		_w28649_,
		_w29221_,
		_w29223_
	);
	LUT2 #(
		.INIT('h4)
	) name25177 (
		_w29222_,
		_w29223_,
		_w29224_
	);
	LUT2 #(
		.INIT('h1)
	) name25178 (
		_w28550_,
		_w29217_,
		_w29225_
	);
	LUT2 #(
		.INIT('h4)
	) name25179 (
		_w29224_,
		_w29225_,
		_w29226_
	);
	LUT2 #(
		.INIT('h1)
	) name25180 (
		_w29216_,
		_w29226_,
		_w29227_
	);
	LUT2 #(
		.INIT('h8)
	) name25181 (
		\sport0_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		_w19552_,
		_w29228_
	);
	LUT2 #(
		.INIT('h1)
	) name25182 (
		\sport0_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		_w29228_,
		_w29229_
	);
	LUT2 #(
		.INIT('h8)
	) name25183 (
		\sport0_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		_w29228_,
		_w29230_
	);
	LUT2 #(
		.INIT('h2)
	) name25184 (
		_w19197_,
		_w29229_,
		_w29231_
	);
	LUT2 #(
		.INIT('h4)
	) name25185 (
		_w29230_,
		_w29231_,
		_w29232_
	);
	LUT2 #(
		.INIT('h4)
	) name25186 (
		_w18127_,
		_w18148_,
		_w29233_
	);
	LUT2 #(
		.INIT('h2)
	) name25187 (
		_w18039_,
		_w19722_,
		_w29234_
	);
	LUT2 #(
		.INIT('h4)
	) name25188 (
		_w18114_,
		_w20104_,
		_w29235_
	);
	LUT2 #(
		.INIT('h2)
	) name25189 (
		_w17980_,
		_w18135_,
		_w29236_
	);
	LUT2 #(
		.INIT('h8)
	) name25190 (
		_w18171_,
		_w18893_,
		_w29237_
	);
	LUT2 #(
		.INIT('h2)
	) name25191 (
		_w18124_,
		_w19804_,
		_w29238_
	);
	LUT2 #(
		.INIT('h1)
	) name25192 (
		_w18783_,
		_w21010_,
		_w29239_
	);
	LUT2 #(
		.INIT('h8)
	) name25193 (
		_w18139_,
		_w18183_,
		_w29240_
	);
	LUT2 #(
		.INIT('h4)
	) name25194 (
		_w17935_,
		_w18072_,
		_w29241_
	);
	LUT2 #(
		.INIT('h8)
	) name25195 (
		_w17971_,
		_w18051_,
		_w29242_
	);
	LUT2 #(
		.INIT('h8)
	) name25196 (
		_w18046_,
		_w18745_,
		_w29243_
	);
	LUT2 #(
		.INIT('h1)
	) name25197 (
		_w18091_,
		_w18104_,
		_w29244_
	);
	LUT2 #(
		.INIT('h8)
	) name25198 (
		_w18071_,
		_w18187_,
		_w29245_
	);
	LUT2 #(
		.INIT('h2)
	) name25199 (
		_w18112_,
		_w18907_,
		_w29246_
	);
	LUT2 #(
		.INIT('h4)
	) name25200 (
		_w18127_,
		_w18147_,
		_w29247_
	);
	LUT2 #(
		.INIT('h8)
	) name25201 (
		_w17979_,
		_w18077_,
		_w29248_
	);
	LUT2 #(
		.INIT('h1)
	) name25202 (
		_w17981_,
		_w29248_,
		_w29249_
	);
	LUT2 #(
		.INIT('h4)
	) name25203 (
		_w18083_,
		_w29249_,
		_w29250_
	);
	LUT2 #(
		.INIT('h2)
	) name25204 (
		_w17945_,
		_w29250_,
		_w29251_
	);
	LUT2 #(
		.INIT('h2)
	) name25205 (
		_w17978_,
		_w29251_,
		_w29252_
	);
	LUT2 #(
		.INIT('h2)
	) name25206 (
		_w18055_,
		_w18189_,
		_w29253_
	);
	LUT2 #(
		.INIT('h2)
	) name25207 (
		_w18056_,
		_w18991_,
		_w29254_
	);
	LUT2 #(
		.INIT('h2)
	) name25208 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11992_,
		_w29255_
	);
	LUT2 #(
		.INIT('h2)
	) name25209 (
		_w18191_,
		_w19722_,
		_w29256_
	);
	LUT2 #(
		.INIT('h8)
	) name25210 (
		_w18153_,
		_w18166_,
		_w29257_
	);
	LUT2 #(
		.INIT('h4)
	) name25211 (
		_w17935_,
		_w17955_,
		_w29258_
	);
	LUT2 #(
		.INIT('h2)
	) name25212 (
		_w18162_,
		_w19857_,
		_w29259_
	);
	LUT2 #(
		.INIT('h1)
	) name25213 (
		_w29253_,
		_w29255_,
		_w29260_
	);
	LUT2 #(
		.INIT('h1)
	) name25214 (
		_w29254_,
		_w29256_,
		_w29261_
	);
	LUT2 #(
		.INIT('h1)
	) name25215 (
		_w29257_,
		_w29258_,
		_w29262_
	);
	LUT2 #(
		.INIT('h8)
	) name25216 (
		_w29261_,
		_w29262_,
		_w29263_
	);
	LUT2 #(
		.INIT('h4)
	) name25217 (
		_w21199_,
		_w29260_,
		_w29264_
	);
	LUT2 #(
		.INIT('h1)
	) name25218 (
		_w29233_,
		_w29234_,
		_w29265_
	);
	LUT2 #(
		.INIT('h1)
	) name25219 (
		_w29241_,
		_w29242_,
		_w29266_
	);
	LUT2 #(
		.INIT('h8)
	) name25220 (
		_w29265_,
		_w29266_,
		_w29267_
	);
	LUT2 #(
		.INIT('h8)
	) name25221 (
		_w29263_,
		_w29264_,
		_w29268_
	);
	LUT2 #(
		.INIT('h1)
	) name25222 (
		_w29236_,
		_w29237_,
		_w29269_
	);
	LUT2 #(
		.INIT('h1)
	) name25223 (
		_w29240_,
		_w29243_,
		_w29270_
	);
	LUT2 #(
		.INIT('h1)
	) name25224 (
		_w29244_,
		_w29245_,
		_w29271_
	);
	LUT2 #(
		.INIT('h1)
	) name25225 (
		_w29246_,
		_w29247_,
		_w29272_
	);
	LUT2 #(
		.INIT('h8)
	) name25226 (
		_w29271_,
		_w29272_,
		_w29273_
	);
	LUT2 #(
		.INIT('h8)
	) name25227 (
		_w29269_,
		_w29270_,
		_w29274_
	);
	LUT2 #(
		.INIT('h8)
	) name25228 (
		_w29267_,
		_w29268_,
		_w29275_
	);
	LUT2 #(
		.INIT('h2)
	) name25229 (
		_w20108_,
		_w29235_,
		_w29276_
	);
	LUT2 #(
		.INIT('h4)
	) name25230 (
		_w29238_,
		_w29239_,
		_w29277_
	);
	LUT2 #(
		.INIT('h4)
	) name25231 (
		_w29259_,
		_w29277_,
		_w29278_
	);
	LUT2 #(
		.INIT('h8)
	) name25232 (
		_w29275_,
		_w29276_,
		_w29279_
	);
	LUT2 #(
		.INIT('h8)
	) name25233 (
		_w29273_,
		_w29274_,
		_w29280_
	);
	LUT2 #(
		.INIT('h8)
	) name25234 (
		_w18724_,
		_w29280_,
		_w29281_
	);
	LUT2 #(
		.INIT('h8)
	) name25235 (
		_w29278_,
		_w29279_,
		_w29282_
	);
	LUT2 #(
		.INIT('h8)
	) name25236 (
		_w29252_,
		_w29282_,
		_w29283_
	);
	LUT2 #(
		.INIT('h8)
	) name25237 (
		_w29281_,
		_w29283_,
		_w29284_
	);
	LUT2 #(
		.INIT('h8)
	) name25238 (
		_w19793_,
		_w29284_,
		_w29285_
	);
	LUT2 #(
		.INIT('h2)
	) name25239 (
		_w28636_,
		_w29285_,
		_w29286_
	);
	LUT2 #(
		.INIT('h8)
	) name25240 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w17820_,
		_w29287_
	);
	LUT2 #(
		.INIT('h8)
	) name25241 (
		_w19214_,
		_w19278_,
		_w29288_
	);
	LUT2 #(
		.INIT('h1)
	) name25242 (
		_w19224_,
		_w29288_,
		_w29289_
	);
	LUT2 #(
		.INIT('h1)
	) name25243 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w29289_,
		_w29290_
	);
	LUT2 #(
		.INIT('h1)
	) name25244 (
		_w29287_,
		_w29290_,
		_w29291_
	);
	LUT2 #(
		.INIT('h2)
	) name25245 (
		_w28559_,
		_w29291_,
		_w29292_
	);
	LUT2 #(
		.INIT('h1)
	) name25246 (
		_w12028_,
		_w28589_,
		_w29293_
	);
	LUT2 #(
		.INIT('h8)
	) name25247 (
		_w28592_,
		_w28601_,
		_w29294_
	);
	LUT2 #(
		.INIT('h1)
	) name25248 (
		_w7206_,
		_w28598_,
		_w29295_
	);
	LUT2 #(
		.INIT('h1)
	) name25249 (
		_w12024_,
		_w28594_,
		_w29296_
	);
	LUT2 #(
		.INIT('h1)
	) name25250 (
		_w28605_,
		_w29293_,
		_w29297_
	);
	LUT2 #(
		.INIT('h1)
	) name25251 (
		_w29294_,
		_w29295_,
		_w29298_
	);
	LUT2 #(
		.INIT('h4)
	) name25252 (
		_w29296_,
		_w29298_,
		_w29299_
	);
	LUT2 #(
		.INIT('h8)
	) name25253 (
		_w29297_,
		_w29299_,
		_w29300_
	);
	LUT2 #(
		.INIT('h2)
	) name25254 (
		_w28577_,
		_w29300_,
		_w29301_
	);
	LUT2 #(
		.INIT('h2)
	) name25255 (
		_w11265_,
		_w28572_,
		_w29302_
	);
	LUT2 #(
		.INIT('h8)
	) name25256 (
		_w28574_,
		_w29302_,
		_w29303_
	);
	LUT2 #(
		.INIT('h1)
	) name25257 (
		_w29301_,
		_w29303_,
		_w29304_
	);
	LUT2 #(
		.INIT('h1)
	) name25258 (
		_w28569_,
		_w29304_,
		_w29305_
	);
	LUT2 #(
		.INIT('h8)
	) name25259 (
		_w13006_,
		_w28992_,
		_w29306_
	);
	LUT2 #(
		.INIT('h1)
	) name25260 (
		_w28576_,
		_w29306_,
		_w29307_
	);
	LUT2 #(
		.INIT('h2)
	) name25261 (
		_w28569_,
		_w29307_,
		_w29308_
	);
	LUT2 #(
		.INIT('h1)
	) name25262 (
		_w12771_,
		_w28572_,
		_w29309_
	);
	LUT2 #(
		.INIT('h4)
	) name25263 (
		_w12743_,
		_w28572_,
		_w29310_
	);
	LUT2 #(
		.INIT('h2)
	) name25264 (
		_w28997_,
		_w29309_,
		_w29311_
	);
	LUT2 #(
		.INIT('h4)
	) name25265 (
		_w29310_,
		_w29311_,
		_w29312_
	);
	LUT2 #(
		.INIT('h8)
	) name25266 (
		_w12771_,
		_w28619_,
		_w29313_
	);
	LUT2 #(
		.INIT('h1)
	) name25267 (
		_w12000_,
		_w28556_,
		_w29314_
	);
	LUT2 #(
		.INIT('h1)
	) name25268 (
		_w11992_,
		_w28624_,
		_w29315_
	);
	LUT2 #(
		.INIT('h1)
	) name25269 (
		_w11983_,
		_w28634_,
		_w29316_
	);
	LUT2 #(
		.INIT('h8)
	) name25270 (
		_w12743_,
		_w28630_,
		_w29317_
	);
	LUT2 #(
		.INIT('h4)
	) name25271 (
		_w19769_,
		_w28627_,
		_w29318_
	);
	LUT2 #(
		.INIT('h1)
	) name25272 (
		_w29313_,
		_w29316_,
		_w29319_
	);
	LUT2 #(
		.INIT('h4)
	) name25273 (
		_w29317_,
		_w29319_,
		_w29320_
	);
	LUT2 #(
		.INIT('h1)
	) name25274 (
		_w29314_,
		_w29315_,
		_w29321_
	);
	LUT2 #(
		.INIT('h8)
	) name25275 (
		_w29320_,
		_w29321_,
		_w29322_
	);
	LUT2 #(
		.INIT('h1)
	) name25276 (
		_w29286_,
		_w29318_,
		_w29323_
	);
	LUT2 #(
		.INIT('h8)
	) name25277 (
		_w29322_,
		_w29323_,
		_w29324_
	);
	LUT2 #(
		.INIT('h4)
	) name25278 (
		_w29312_,
		_w29324_,
		_w29325_
	);
	LUT2 #(
		.INIT('h4)
	) name25279 (
		_w29305_,
		_w29325_,
		_w29326_
	);
	LUT2 #(
		.INIT('h4)
	) name25280 (
		_w29308_,
		_w29326_,
		_w29327_
	);
	LUT2 #(
		.INIT('h4)
	) name25281 (
		_w29292_,
		_w29327_,
		_w29328_
	);
	LUT2 #(
		.INIT('h2)
	) name25282 (
		_w28550_,
		_w29328_,
		_w29329_
	);
	LUT2 #(
		.INIT('h4)
	) name25283 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[15]/P0001 ,
		_w28649_,
		_w29330_
	);
	LUT2 #(
		.INIT('h8)
	) name25284 (
		_w12016_,
		_w28652_,
		_w29331_
	);
	LUT2 #(
		.INIT('h2)
	) name25285 (
		_w12020_,
		_w28652_,
		_w29332_
	);
	LUT2 #(
		.INIT('h1)
	) name25286 (
		_w28660_,
		_w29331_,
		_w29333_
	);
	LUT2 #(
		.INIT('h4)
	) name25287 (
		_w29332_,
		_w29333_,
		_w29334_
	);
	LUT2 #(
		.INIT('h8)
	) name25288 (
		_w17820_,
		_w28660_,
		_w29335_
	);
	LUT2 #(
		.INIT('h1)
	) name25289 (
		_w28649_,
		_w29334_,
		_w29336_
	);
	LUT2 #(
		.INIT('h4)
	) name25290 (
		_w29335_,
		_w29336_,
		_w29337_
	);
	LUT2 #(
		.INIT('h1)
	) name25291 (
		_w28550_,
		_w29330_,
		_w29338_
	);
	LUT2 #(
		.INIT('h4)
	) name25292 (
		_w29337_,
		_w29338_,
		_w29339_
	);
	LUT2 #(
		.INIT('h1)
	) name25293 (
		_w29329_,
		_w29339_,
		_w29340_
	);
	LUT2 #(
		.INIT('h2)
	) name25294 (
		\sport0_txctl_TXSHT_reg[11]/P0001 ,
		_w19960_,
		_w29341_
	);
	LUT2 #(
		.INIT('h8)
	) name25295 (
		\sport0_txctl_TX_reg[12]/P0001 ,
		_w19960_,
		_w29342_
	);
	LUT2 #(
		.INIT('h1)
	) name25296 (
		_w29341_,
		_w29342_,
		_w29343_
	);
	LUT2 #(
		.INIT('h8)
	) name25297 (
		_w12802_,
		_w28729_,
		_w29344_
	);
	LUT2 #(
		.INIT('h8)
	) name25298 (
		_w9435_,
		_w28725_,
		_w29345_
	);
	LUT2 #(
		.INIT('h8)
	) name25299 (
		_w9209_,
		_w28705_,
		_w29346_
	);
	LUT2 #(
		.INIT('h2)
	) name25300 (
		_w9217_,
		_w28705_,
		_w29347_
	);
	LUT2 #(
		.INIT('h1)
	) name25301 (
		_w29346_,
		_w29347_,
		_w29348_
	);
	LUT2 #(
		.INIT('h8)
	) name25302 (
		_w28735_,
		_w29348_,
		_w29349_
	);
	LUT2 #(
		.INIT('h8)
	) name25303 (
		_w28739_,
		_w29221_,
		_w29350_
	);
	LUT2 #(
		.INIT('h1)
	) name25304 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[1]/P0001 ,
		_w29351_
	);
	LUT2 #(
		.INIT('h2)
	) name25305 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[1]/P0001 ,
		_w29352_
	);
	LUT2 #(
		.INIT('h1)
	) name25306 (
		_w29351_,
		_w29352_,
		_w29353_
	);
	LUT2 #(
		.INIT('h8)
	) name25307 (
		_w28741_,
		_w29353_,
		_w29354_
	);
	LUT2 #(
		.INIT('h1)
	) name25308 (
		_w29349_,
		_w29350_,
		_w29355_
	);
	LUT2 #(
		.INIT('h4)
	) name25309 (
		_w29354_,
		_w29355_,
		_w29356_
	);
	LUT2 #(
		.INIT('h4)
	) name25310 (
		_w29344_,
		_w29356_,
		_w29357_
	);
	LUT2 #(
		.INIT('h4)
	) name25311 (
		_w29345_,
		_w29357_,
		_w29358_
	);
	LUT2 #(
		.INIT('h1)
	) name25312 (
		_w28543_,
		_w29358_,
		_w29359_
	);
	LUT2 #(
		.INIT('h2)
	) name25313 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[1]/P0001 ,
		_w28545_,
		_w29360_
	);
	LUT2 #(
		.INIT('h1)
	) name25314 (
		_w29359_,
		_w29360_,
		_w29361_
	);
	LUT2 #(
		.INIT('h1)
	) name25315 (
		_w28719_,
		_w29361_,
		_w29362_
	);
	LUT2 #(
		.INIT('h2)
	) name25316 (
		_w28719_,
		_w29215_,
		_w29363_
	);
	LUT2 #(
		.INIT('h1)
	) name25317 (
		_w29362_,
		_w29363_,
		_w29364_
	);
	LUT2 #(
		.INIT('h8)
	) name25318 (
		_w12904_,
		_w28729_,
		_w29365_
	);
	LUT2 #(
		.INIT('h8)
	) name25319 (
		_w10069_,
		_w28725_,
		_w29366_
	);
	LUT2 #(
		.INIT('h8)
	) name25320 (
		_w9853_,
		_w28705_,
		_w29367_
	);
	LUT2 #(
		.INIT('h2)
	) name25321 (
		_w9857_,
		_w28705_,
		_w29368_
	);
	LUT2 #(
		.INIT('h1)
	) name25322 (
		_w29367_,
		_w29368_,
		_w29369_
	);
	LUT2 #(
		.INIT('h8)
	) name25323 (
		_w28735_,
		_w29369_,
		_w29370_
	);
	LUT2 #(
		.INIT('h8)
	) name25324 (
		_w28739_,
		_w29172_,
		_w29371_
	);
	LUT2 #(
		.INIT('h1)
	) name25325 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[4]/P0001 ,
		_w29372_
	);
	LUT2 #(
		.INIT('h2)
	) name25326 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[4]/P0001 ,
		_w29373_
	);
	LUT2 #(
		.INIT('h1)
	) name25327 (
		_w29372_,
		_w29373_,
		_w29374_
	);
	LUT2 #(
		.INIT('h8)
	) name25328 (
		_w28741_,
		_w29374_,
		_w29375_
	);
	LUT2 #(
		.INIT('h1)
	) name25329 (
		_w29370_,
		_w29371_,
		_w29376_
	);
	LUT2 #(
		.INIT('h4)
	) name25330 (
		_w29375_,
		_w29376_,
		_w29377_
	);
	LUT2 #(
		.INIT('h4)
	) name25331 (
		_w29365_,
		_w29377_,
		_w29378_
	);
	LUT2 #(
		.INIT('h4)
	) name25332 (
		_w29366_,
		_w29378_,
		_w29379_
	);
	LUT2 #(
		.INIT('h1)
	) name25333 (
		_w28543_,
		_w29379_,
		_w29380_
	);
	LUT2 #(
		.INIT('h2)
	) name25334 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[4]/P0001 ,
		_w28545_,
		_w29381_
	);
	LUT2 #(
		.INIT('h1)
	) name25335 (
		_w29380_,
		_w29381_,
		_w29382_
	);
	LUT2 #(
		.INIT('h1)
	) name25336 (
		_w28719_,
		_w29382_,
		_w29383_
	);
	LUT2 #(
		.INIT('h2)
	) name25337 (
		_w28719_,
		_w29166_,
		_w29384_
	);
	LUT2 #(
		.INIT('h1)
	) name25338 (
		_w29383_,
		_w29384_,
		_w29385_
	);
	LUT2 #(
		.INIT('h8)
	) name25339 (
		_w12972_,
		_w28729_,
		_w29386_
	);
	LUT2 #(
		.INIT('h8)
	) name25340 (
		_w11525_,
		_w28725_,
		_w29387_
	);
	LUT2 #(
		.INIT('h8)
	) name25341 (
		_w11436_,
		_w28705_,
		_w29388_
	);
	LUT2 #(
		.INIT('h2)
	) name25342 (
		_w11432_,
		_w28705_,
		_w29389_
	);
	LUT2 #(
		.INIT('h1)
	) name25343 (
		_w29388_,
		_w29389_,
		_w29390_
	);
	LUT2 #(
		.INIT('h8)
	) name25344 (
		_w28735_,
		_w29390_,
		_w29391_
	);
	LUT2 #(
		.INIT('h8)
	) name25345 (
		_w28739_,
		_w29032_,
		_w29392_
	);
	LUT2 #(
		.INIT('h1)
	) name25346 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[6]/P0001 ,
		_w29393_
	);
	LUT2 #(
		.INIT('h2)
	) name25347 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[6]/P0001 ,
		_w29394_
	);
	LUT2 #(
		.INIT('h1)
	) name25348 (
		_w29393_,
		_w29394_,
		_w29395_
	);
	LUT2 #(
		.INIT('h8)
	) name25349 (
		_w28741_,
		_w29395_,
		_w29396_
	);
	LUT2 #(
		.INIT('h1)
	) name25350 (
		_w29391_,
		_w29392_,
		_w29397_
	);
	LUT2 #(
		.INIT('h4)
	) name25351 (
		_w29396_,
		_w29397_,
		_w29398_
	);
	LUT2 #(
		.INIT('h4)
	) name25352 (
		_w29386_,
		_w29398_,
		_w29399_
	);
	LUT2 #(
		.INIT('h4)
	) name25353 (
		_w29387_,
		_w29399_,
		_w29400_
	);
	LUT2 #(
		.INIT('h1)
	) name25354 (
		_w28543_,
		_w29400_,
		_w29401_
	);
	LUT2 #(
		.INIT('h2)
	) name25355 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[6]/P0001 ,
		_w28545_,
		_w29402_
	);
	LUT2 #(
		.INIT('h1)
	) name25356 (
		_w29401_,
		_w29402_,
		_w29403_
	);
	LUT2 #(
		.INIT('h1)
	) name25357 (
		_w28719_,
		_w29403_,
		_w29404_
	);
	LUT2 #(
		.INIT('h2)
	) name25358 (
		_w28719_,
		_w29026_,
		_w29405_
	);
	LUT2 #(
		.INIT('h1)
	) name25359 (
		_w29404_,
		_w29405_,
		_w29406_
	);
	LUT2 #(
		.INIT('h8)
	) name25360 (
		\sport1_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		_w20253_,
		_w29407_
	);
	LUT2 #(
		.INIT('h1)
	) name25361 (
		\sport1_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		_w29407_,
		_w29408_
	);
	LUT2 #(
		.INIT('h8)
	) name25362 (
		\sport1_cfg_SCLKi_cnt_reg[15]/NET0131 ,
		_w29407_,
		_w29409_
	);
	LUT2 #(
		.INIT('h2)
	) name25363 (
		_w19130_,
		_w29408_,
		_w29410_
	);
	LUT2 #(
		.INIT('h4)
	) name25364 (
		_w29409_,
		_w29410_,
		_w29411_
	);
	LUT2 #(
		.INIT('h8)
	) name25365 (
		_w12938_,
		_w28729_,
		_w29412_
	);
	LUT2 #(
		.INIT('h8)
	) name25366 (
		_w10911_,
		_w28725_,
		_w29413_
	);
	LUT2 #(
		.INIT('h8)
	) name25367 (
		_w10862_,
		_w28705_,
		_w29414_
	);
	LUT2 #(
		.INIT('h2)
	) name25368 (
		_w10870_,
		_w28705_,
		_w29415_
	);
	LUT2 #(
		.INIT('h1)
	) name25369 (
		_w29414_,
		_w29415_,
		_w29416_
	);
	LUT2 #(
		.INIT('h8)
	) name25370 (
		_w28735_,
		_w29416_,
		_w29417_
	);
	LUT2 #(
		.INIT('h8)
	) name25371 (
		_w28739_,
		_w29121_,
		_w29418_
	);
	LUT2 #(
		.INIT('h1)
	) name25372 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[5]/P0001 ,
		_w29419_
	);
	LUT2 #(
		.INIT('h2)
	) name25373 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[5]/P0001 ,
		_w29420_
	);
	LUT2 #(
		.INIT('h1)
	) name25374 (
		_w29419_,
		_w29420_,
		_w29421_
	);
	LUT2 #(
		.INIT('h8)
	) name25375 (
		_w28741_,
		_w29421_,
		_w29422_
	);
	LUT2 #(
		.INIT('h1)
	) name25376 (
		_w29417_,
		_w29418_,
		_w29423_
	);
	LUT2 #(
		.INIT('h4)
	) name25377 (
		_w29422_,
		_w29423_,
		_w29424_
	);
	LUT2 #(
		.INIT('h4)
	) name25378 (
		_w29412_,
		_w29424_,
		_w29425_
	);
	LUT2 #(
		.INIT('h4)
	) name25379 (
		_w29413_,
		_w29425_,
		_w29426_
	);
	LUT2 #(
		.INIT('h1)
	) name25380 (
		_w28543_,
		_w29426_,
		_w29427_
	);
	LUT2 #(
		.INIT('h2)
	) name25381 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[5]/P0001 ,
		_w28545_,
		_w29428_
	);
	LUT2 #(
		.INIT('h1)
	) name25382 (
		_w29427_,
		_w29428_,
		_w29429_
	);
	LUT2 #(
		.INIT('h1)
	) name25383 (
		_w28719_,
		_w29429_,
		_w29430_
	);
	LUT2 #(
		.INIT('h2)
	) name25384 (
		_w28719_,
		_w29115_,
		_w29431_
	);
	LUT2 #(
		.INIT('h1)
	) name25385 (
		_w29430_,
		_w29431_,
		_w29432_
	);
	LUT2 #(
		.INIT('h8)
	) name25386 (
		_w12771_,
		_w28729_,
		_w29433_
	);
	LUT2 #(
		.INIT('h8)
	) name25387 (
		_w12743_,
		_w28725_,
		_w29434_
	);
	LUT2 #(
		.INIT('h8)
	) name25388 (
		_w12008_,
		_w28705_,
		_w29435_
	);
	LUT2 #(
		.INIT('h2)
	) name25389 (
		_w12012_,
		_w28705_,
		_w29436_
	);
	LUT2 #(
		.INIT('h1)
	) name25390 (
		_w29435_,
		_w29436_,
		_w29437_
	);
	LUT2 #(
		.INIT('h8)
	) name25391 (
		_w28735_,
		_w29437_,
		_w29438_
	);
	LUT2 #(
		.INIT('h8)
	) name25392 (
		_w28739_,
		_w29334_,
		_w29439_
	);
	LUT2 #(
		.INIT('h1)
	) name25393 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[15]/P0001 ,
		_w29440_
	);
	LUT2 #(
		.INIT('h2)
	) name25394 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[15]/P0001 ,
		_w29441_
	);
	LUT2 #(
		.INIT('h1)
	) name25395 (
		_w29440_,
		_w29441_,
		_w29442_
	);
	LUT2 #(
		.INIT('h8)
	) name25396 (
		_w28741_,
		_w29442_,
		_w29443_
	);
	LUT2 #(
		.INIT('h1)
	) name25397 (
		_w29438_,
		_w29439_,
		_w29444_
	);
	LUT2 #(
		.INIT('h4)
	) name25398 (
		_w29443_,
		_w29444_,
		_w29445_
	);
	LUT2 #(
		.INIT('h4)
	) name25399 (
		_w29434_,
		_w29445_,
		_w29446_
	);
	LUT2 #(
		.INIT('h4)
	) name25400 (
		_w29433_,
		_w29446_,
		_w29447_
	);
	LUT2 #(
		.INIT('h1)
	) name25401 (
		_w28543_,
		_w29447_,
		_w29448_
	);
	LUT2 #(
		.INIT('h2)
	) name25402 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[15]/P0001 ,
		_w28545_,
		_w29449_
	);
	LUT2 #(
		.INIT('h1)
	) name25403 (
		_w29448_,
		_w29449_,
		_w29450_
	);
	LUT2 #(
		.INIT('h1)
	) name25404 (
		_w28719_,
		_w29450_,
		_w29451_
	);
	LUT2 #(
		.INIT('h2)
	) name25405 (
		_w28719_,
		_w29328_,
		_w29452_
	);
	LUT2 #(
		.INIT('h1)
	) name25406 (
		_w29451_,
		_w29452_,
		_w29453_
	);
	LUT2 #(
		.INIT('h2)
	) name25407 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[7]/P0001 ,
		_w23598_,
		_w29454_
	);
	LUT2 #(
		.INIT('h8)
	) name25408 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w19972_,
		_w29455_
	);
	LUT2 #(
		.INIT('h1)
	) name25409 (
		_w23587_,
		_w23662_,
		_w29456_
	);
	LUT2 #(
		.INIT('h1)
	) name25410 (
		_w23665_,
		_w29456_,
		_w29457_
	);
	LUT2 #(
		.INIT('h4)
	) name25411 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w29457_,
		_w29458_
	);
	LUT2 #(
		.INIT('h1)
	) name25412 (
		_w29455_,
		_w29458_,
		_w29459_
	);
	LUT2 #(
		.INIT('h2)
	) name25413 (
		_w23598_,
		_w29459_,
		_w29460_
	);
	LUT2 #(
		.INIT('h1)
	) name25414 (
		_w29454_,
		_w29460_,
		_w29461_
	);
	LUT2 #(
		.INIT('h2)
	) name25415 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[6]/P0001 ,
		_w23598_,
		_w29462_
	);
	LUT2 #(
		.INIT('h8)
	) name25416 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w18276_,
		_w29463_
	);
	LUT2 #(
		.INIT('h1)
	) name25417 (
		_w29458_,
		_w29463_,
		_w29464_
	);
	LUT2 #(
		.INIT('h2)
	) name25418 (
		_w23598_,
		_w29464_,
		_w29465_
	);
	LUT2 #(
		.INIT('h1)
	) name25419 (
		_w29462_,
		_w29465_,
		_w29466_
	);
	LUT2 #(
		.INIT('h2)
	) name25420 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 ,
		_w18266_,
		_w29467_
	);
	LUT2 #(
		.INIT('h1)
	) name25421 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[12]/P0001 ,
		_w18271_,
		_w29468_
	);
	LUT2 #(
		.INIT('h2)
	) name25422 (
		_w18271_,
		_w23920_,
		_w29469_
	);
	LUT2 #(
		.INIT('h2)
	) name25423 (
		_w18273_,
		_w29468_,
		_w29470_
	);
	LUT2 #(
		.INIT('h4)
	) name25424 (
		_w29469_,
		_w29470_,
		_w29471_
	);
	LUT2 #(
		.INIT('h1)
	) name25425 (
		_w18270_,
		_w29467_,
		_w29472_
	);
	LUT2 #(
		.INIT('h4)
	) name25426 (
		_w29471_,
		_w29472_,
		_w29473_
	);
	LUT2 #(
		.INIT('h1)
	) name25427 (
		_w18262_,
		_w29473_,
		_w29474_
	);
	LUT2 #(
		.INIT('h8)
	) name25428 (
		_w18262_,
		_w19609_,
		_w29475_
	);
	LUT2 #(
		.INIT('h1)
	) name25429 (
		_w29474_,
		_w29475_,
		_w29476_
	);
	LUT2 #(
		.INIT('h2)
	) name25430 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w20080_,
		_w29477_
	);
	LUT2 #(
		.INIT('h8)
	) name25431 (
		_w23587_,
		_w23662_,
		_w29478_
	);
	LUT2 #(
		.INIT('h2)
	) name25432 (
		_w29457_,
		_w29478_,
		_w29479_
	);
	LUT2 #(
		.INIT('h1)
	) name25433 (
		_w23669_,
		_w29479_,
		_w29480_
	);
	LUT2 #(
		.INIT('h4)
	) name25434 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w29480_,
		_w29481_
	);
	LUT2 #(
		.INIT('h1)
	) name25435 (
		_w29477_,
		_w29481_,
		_w29482_
	);
	LUT2 #(
		.INIT('h2)
	) name25436 (
		_w23598_,
		_w29482_,
		_w29483_
	);
	LUT2 #(
		.INIT('h1)
	) name25437 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[4]/P0001 ,
		_w23598_,
		_w29484_
	);
	LUT2 #(
		.INIT('h1)
	) name25438 (
		_w29483_,
		_w29484_,
		_w29485_
	);
	LUT2 #(
		.INIT('h2)
	) name25439 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[5]/P0001 ,
		_w23598_,
		_w29486_
	);
	LUT2 #(
		.INIT('h8)
	) name25440 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w20259_,
		_w29487_
	);
	LUT2 #(
		.INIT('h1)
	) name25441 (
		_w29458_,
		_w29487_,
		_w29488_
	);
	LUT2 #(
		.INIT('h2)
	) name25442 (
		_w23598_,
		_w29488_,
		_w29489_
	);
	LUT2 #(
		.INIT('h1)
	) name25443 (
		_w29486_,
		_w29489_,
		_w29490_
	);
	LUT2 #(
		.INIT('h2)
	) name25444 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w21663_,
		_w29491_
	);
	LUT2 #(
		.INIT('h8)
	) name25445 (
		_w27484_,
		_w27486_,
		_w29492_
	);
	LUT2 #(
		.INIT('h2)
	) name25446 (
		_w26275_,
		_w29492_,
		_w29493_
	);
	LUT2 #(
		.INIT('h1)
	) name25447 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w29493_,
		_w29494_
	);
	LUT2 #(
		.INIT('h1)
	) name25448 (
		_w29491_,
		_w29494_,
		_w29495_
	);
	LUT2 #(
		.INIT('h2)
	) name25449 (
		_w23598_,
		_w29495_,
		_w29496_
	);
	LUT2 #(
		.INIT('h1)
	) name25450 (
		\core_eu_es_sht_es_reg_serwe_DO_reg[3]/P0001 ,
		_w23598_,
		_w29497_
	);
	LUT2 #(
		.INIT('h1)
	) name25451 (
		_w29496_,
		_w29497_,
		_w29498_
	);
	LUT2 #(
		.INIT('h2)
	) name25452 (
		_w14752_,
		_w19609_,
		_w29499_
	);
	LUT2 #(
		.INIT('h8)
	) name25453 (
		_w18328_,
		_w23920_,
		_w29500_
	);
	LUT2 #(
		.INIT('h2)
	) name25454 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[12]/P0001 ,
		_w18330_,
		_w29501_
	);
	LUT2 #(
		.INIT('h2)
	) name25455 (
		_w18334_,
		_w29501_,
		_w29502_
	);
	LUT2 #(
		.INIT('h4)
	) name25456 (
		_w29500_,
		_w29502_,
		_w29503_
	);
	LUT2 #(
		.INIT('h1)
	) name25457 (
		_w29499_,
		_w29503_,
		_w29504_
	);
	LUT2 #(
		.INIT('h2)
	) name25458 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[6]/P0001 ,
		_w23677_,
		_w29505_
	);
	LUT2 #(
		.INIT('h2)
	) name25459 (
		_w23677_,
		_w29464_,
		_w29506_
	);
	LUT2 #(
		.INIT('h1)
	) name25460 (
		_w29505_,
		_w29506_,
		_w29507_
	);
	LUT2 #(
		.INIT('h2)
	) name25461 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[7]/P0001 ,
		_w23677_,
		_w29508_
	);
	LUT2 #(
		.INIT('h2)
	) name25462 (
		_w23677_,
		_w29459_,
		_w29509_
	);
	LUT2 #(
		.INIT('h1)
	) name25463 (
		_w29508_,
		_w29509_,
		_w29510_
	);
	LUT2 #(
		.INIT('h2)
	) name25464 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[5]/P0001 ,
		_w23677_,
		_w29511_
	);
	LUT2 #(
		.INIT('h2)
	) name25465 (
		_w23677_,
		_w29488_,
		_w29512_
	);
	LUT2 #(
		.INIT('h1)
	) name25466 (
		_w29511_,
		_w29512_,
		_w29513_
	);
	LUT2 #(
		.INIT('h2)
	) name25467 (
		_w23677_,
		_w29482_,
		_w29514_
	);
	LUT2 #(
		.INIT('h1)
	) name25468 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[4]/P0001 ,
		_w23677_,
		_w29515_
	);
	LUT2 #(
		.INIT('h1)
	) name25469 (
		_w29514_,
		_w29515_,
		_w29516_
	);
	LUT2 #(
		.INIT('h2)
	) name25470 (
		_w23677_,
		_w29495_,
		_w29517_
	);
	LUT2 #(
		.INIT('h1)
	) name25471 (
		\core_eu_es_sht_es_reg_seswe_DO_reg[3]/P0001 ,
		_w23677_,
		_w29518_
	);
	LUT2 #(
		.INIT('h1)
	) name25472 (
		_w29517_,
		_w29518_,
		_w29519_
	);
	LUT2 #(
		.INIT('h1)
	) name25473 (
		_w18167_,
		_w18907_,
		_w29520_
	);
	LUT2 #(
		.INIT('h8)
	) name25474 (
		_w19855_,
		_w19873_,
		_w29521_
	);
	LUT2 #(
		.INIT('h8)
	) name25475 (
		_w19713_,
		_w29521_,
		_w29522_
	);
	LUT2 #(
		.INIT('h1)
	) name25476 (
		_w18189_,
		_w18912_,
		_w29523_
	);
	LUT2 #(
		.INIT('h2)
	) name25477 (
		_w18112_,
		_w18914_,
		_w29524_
	);
	LUT2 #(
		.INIT('h2)
	) name25478 (
		_w18751_,
		_w18775_,
		_w29525_
	);
	LUT2 #(
		.INIT('h4)
	) name25479 (
		_w17998_,
		_w18748_,
		_w29526_
	);
	LUT2 #(
		.INIT('h4)
	) name25480 (
		_w18079_,
		_w19720_,
		_w29527_
	);
	LUT2 #(
		.INIT('h2)
	) name25481 (
		_w18172_,
		_w18918_,
		_w29528_
	);
	LUT2 #(
		.INIT('h2)
	) name25482 (
		_w18740_,
		_w18781_,
		_w29529_
	);
	LUT2 #(
		.INIT('h2)
	) name25483 (
		_w17925_,
		_w18898_,
		_w29530_
	);
	LUT2 #(
		.INIT('h2)
	) name25484 (
		_w18099_,
		_w19818_,
		_w29531_
	);
	LUT2 #(
		.INIT('h2)
	) name25485 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w10218_,
		_w29532_
	);
	LUT2 #(
		.INIT('h4)
	) name25486 (
		_w18079_,
		_w18765_,
		_w29533_
	);
	LUT2 #(
		.INIT('h2)
	) name25487 (
		_w18758_,
		_w18918_,
		_w29534_
	);
	LUT2 #(
		.INIT('h2)
	) name25488 (
		_w18115_,
		_w18914_,
		_w29535_
	);
	LUT2 #(
		.INIT('h1)
	) name25489 (
		_w29534_,
		_w29535_,
		_w29536_
	);
	LUT2 #(
		.INIT('h2)
	) name25490 (
		_w17839_,
		_w29536_,
		_w29537_
	);
	LUT2 #(
		.INIT('h1)
	) name25491 (
		_w29533_,
		_w29537_,
		_w29538_
	);
	LUT2 #(
		.INIT('h2)
	) name25492 (
		_w17929_,
		_w29538_,
		_w29539_
	);
	LUT2 #(
		.INIT('h2)
	) name25493 (
		_w18124_,
		_w18895_,
		_w29540_
	);
	LUT2 #(
		.INIT('h1)
	) name25494 (
		_w18037_,
		_w29532_,
		_w29541_
	);
	LUT2 #(
		.INIT('h4)
	) name25495 (
		_w18053_,
		_w29541_,
		_w29542_
	);
	LUT2 #(
		.INIT('h1)
	) name25496 (
		_w29520_,
		_w29523_,
		_w29543_
	);
	LUT2 #(
		.INIT('h1)
	) name25497 (
		_w29524_,
		_w29527_,
		_w29544_
	);
	LUT2 #(
		.INIT('h4)
	) name25498 (
		_w29528_,
		_w29544_,
		_w29545_
	);
	LUT2 #(
		.INIT('h8)
	) name25499 (
		_w29542_,
		_w29543_,
		_w29546_
	);
	LUT2 #(
		.INIT('h1)
	) name25500 (
		_w29525_,
		_w29526_,
		_w29547_
	);
	LUT2 #(
		.INIT('h1)
	) name25501 (
		_w29529_,
		_w29530_,
		_w29548_
	);
	LUT2 #(
		.INIT('h1)
	) name25502 (
		_w29531_,
		_w29540_,
		_w29549_
	);
	LUT2 #(
		.INIT('h8)
	) name25503 (
		_w29548_,
		_w29549_,
		_w29550_
	);
	LUT2 #(
		.INIT('h8)
	) name25504 (
		_w29546_,
		_w29547_,
		_w29551_
	);
	LUT2 #(
		.INIT('h8)
	) name25505 (
		_w29545_,
		_w29551_,
		_w29552_
	);
	LUT2 #(
		.INIT('h8)
	) name25506 (
		_w29550_,
		_w29552_,
		_w29553_
	);
	LUT2 #(
		.INIT('h4)
	) name25507 (
		_w29539_,
		_w29553_,
		_w29554_
	);
	LUT2 #(
		.INIT('h8)
	) name25508 (
		_w29522_,
		_w29554_,
		_w29555_
	);
	LUT2 #(
		.INIT('h2)
	) name25509 (
		_w28636_,
		_w29555_,
		_w29556_
	);
	LUT2 #(
		.INIT('h8)
	) name25510 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w19504_,
		_w29557_
	);
	LUT2 #(
		.INIT('h4)
	) name25511 (
		_w14649_,
		_w28561_,
		_w29558_
	);
	LUT2 #(
		.INIT('h1)
	) name25512 (
		_w28564_,
		_w29557_,
		_w29559_
	);
	LUT2 #(
		.INIT('h4)
	) name25513 (
		_w29558_,
		_w29559_,
		_w29560_
	);
	LUT2 #(
		.INIT('h2)
	) name25514 (
		_w28559_,
		_w29560_,
		_w29561_
	);
	LUT2 #(
		.INIT('h2)
	) name25515 (
		_w28607_,
		_w29295_,
		_w29562_
	);
	LUT2 #(
		.INIT('h1)
	) name25516 (
		_w10096_,
		_w28589_,
		_w29563_
	);
	LUT2 #(
		.INIT('h1)
	) name25517 (
		_w10112_,
		_w28594_,
		_w29564_
	);
	LUT2 #(
		.INIT('h1)
	) name25518 (
		_w29563_,
		_w29564_,
		_w29565_
	);
	LUT2 #(
		.INIT('h8)
	) name25519 (
		_w29562_,
		_w29565_,
		_w29566_
	);
	LUT2 #(
		.INIT('h2)
	) name25520 (
		_w28577_,
		_w29566_,
		_w29567_
	);
	LUT2 #(
		.INIT('h1)
	) name25521 (
		_w29303_,
		_w29567_,
		_w29568_
	);
	LUT2 #(
		.INIT('h1)
	) name25522 (
		_w28569_,
		_w29568_,
		_w29569_
	);
	LUT2 #(
		.INIT('h1)
	) name25523 (
		_w10191_,
		_w28634_,
		_w29570_
	);
	LUT2 #(
		.INIT('h8)
	) name25524 (
		_w13075_,
		_w28619_,
		_w29571_
	);
	LUT2 #(
		.INIT('h8)
	) name25525 (
		_w10289_,
		_w28630_,
		_w29572_
	);
	LUT2 #(
		.INIT('h1)
	) name25526 (
		_w10218_,
		_w28624_,
		_w29573_
	);
	LUT2 #(
		.INIT('h1)
	) name25527 (
		_w10226_,
		_w28556_,
		_w29574_
	);
	LUT2 #(
		.INIT('h4)
	) name25528 (
		_w18091_,
		_w18112_,
		_w29575_
	);
	LUT2 #(
		.INIT('h8)
	) name25529 (
		_w18147_,
		_w18748_,
		_w29576_
	);
	LUT2 #(
		.INIT('h4)
	) name25530 (
		_w17922_,
		_w18136_,
		_w29577_
	);
	LUT2 #(
		.INIT('h1)
	) name25531 (
		_w18104_,
		_w18159_,
		_w29578_
	);
	LUT2 #(
		.INIT('h1)
	) name25532 (
		_w18065_,
		_w18735_,
		_w29579_
	);
	LUT2 #(
		.INIT('h2)
	) name25533 (
		_w17925_,
		_w19979_,
		_w29580_
	);
	LUT2 #(
		.INIT('h2)
	) name25534 (
		_w18107_,
		_w18189_,
		_w29581_
	);
	LUT2 #(
		.INIT('h8)
	) name25535 (
		_w18070_,
		_w18088_,
		_w29582_
	);
	LUT2 #(
		.INIT('h2)
	) name25536 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w10226_,
		_w29583_
	);
	LUT2 #(
		.INIT('h2)
	) name25537 (
		_w18106_,
		_w18189_,
		_w29584_
	);
	LUT2 #(
		.INIT('h2)
	) name25538 (
		_w18132_,
		_w18167_,
		_w29585_
	);
	LUT2 #(
		.INIT('h8)
	) name25539 (
		_w17921_,
		_w18172_,
		_w29586_
	);
	LUT2 #(
		.INIT('h8)
	) name25540 (
		_w18089_,
		_w18116_,
		_w29587_
	);
	LUT2 #(
		.INIT('h4)
	) name25541 (
		_w18114_,
		_w18732_,
		_w29588_
	);
	LUT2 #(
		.INIT('h1)
	) name25542 (
		_w17980_,
		_w18071_,
		_w29589_
	);
	LUT2 #(
		.INIT('h2)
	) name25543 (
		_w17945_,
		_w29589_,
		_w29590_
	);
	LUT2 #(
		.INIT('h4)
	) name25544 (
		_w18129_,
		_w18178_,
		_w29591_
	);
	LUT2 #(
		.INIT('h2)
	) name25545 (
		_w18153_,
		_w19722_,
		_w29592_
	);
	LUT2 #(
		.INIT('h8)
	) name25546 (
		_w17934_,
		_w17986_,
		_w29593_
	);
	LUT2 #(
		.INIT('h4)
	) name25547 (
		_w18129_,
		_w18179_,
		_w29594_
	);
	LUT2 #(
		.INIT('h2)
	) name25548 (
		_w18131_,
		_w18167_,
		_w29595_
	);
	LUT2 #(
		.INIT('h8)
	) name25549 (
		_w17915_,
		_w18172_,
		_w29596_
	);
	LUT2 #(
		.INIT('h2)
	) name25550 (
		_w18765_,
		_w29063_,
		_w29597_
	);
	LUT2 #(
		.INIT('h1)
	) name25551 (
		_w29583_,
		_w29584_,
		_w29598_
	);
	LUT2 #(
		.INIT('h1)
	) name25552 (
		_w29585_,
		_w29586_,
		_w29599_
	);
	LUT2 #(
		.INIT('h1)
	) name25553 (
		_w29587_,
		_w29591_,
		_w29600_
	);
	LUT2 #(
		.INIT('h1)
	) name25554 (
		_w29592_,
		_w29593_,
		_w29601_
	);
	LUT2 #(
		.INIT('h8)
	) name25555 (
		_w29600_,
		_w29601_,
		_w29602_
	);
	LUT2 #(
		.INIT('h8)
	) name25556 (
		_w29598_,
		_w29599_,
		_w29603_
	);
	LUT2 #(
		.INIT('h1)
	) name25557 (
		_w18058_,
		_w18783_,
		_w29604_
	);
	LUT2 #(
		.INIT('h1)
	) name25558 (
		_w29581_,
		_w29594_,
		_w29605_
	);
	LUT2 #(
		.INIT('h1)
	) name25559 (
		_w29595_,
		_w29596_,
		_w29606_
	);
	LUT2 #(
		.INIT('h8)
	) name25560 (
		_w29605_,
		_w29606_,
		_w29607_
	);
	LUT2 #(
		.INIT('h8)
	) name25561 (
		_w29603_,
		_w29604_,
		_w29608_
	);
	LUT2 #(
		.INIT('h8)
	) name25562 (
		_w17978_,
		_w29602_,
		_w29609_
	);
	LUT2 #(
		.INIT('h1)
	) name25563 (
		_w18140_,
		_w29575_,
		_w29610_
	);
	LUT2 #(
		.INIT('h1)
	) name25564 (
		_w29576_,
		_w29577_,
		_w29611_
	);
	LUT2 #(
		.INIT('h1)
	) name25565 (
		_w29578_,
		_w29582_,
		_w29612_
	);
	LUT2 #(
		.INIT('h4)
	) name25566 (
		_w29588_,
		_w29612_,
		_w29613_
	);
	LUT2 #(
		.INIT('h8)
	) name25567 (
		_w29610_,
		_w29611_,
		_w29614_
	);
	LUT2 #(
		.INIT('h8)
	) name25568 (
		_w29608_,
		_w29609_,
		_w29615_
	);
	LUT2 #(
		.INIT('h4)
	) name25569 (
		_w29580_,
		_w29607_,
		_w29616_
	);
	LUT2 #(
		.INIT('h1)
	) name25570 (
		_w29590_,
		_w29597_,
		_w29617_
	);
	LUT2 #(
		.INIT('h8)
	) name25571 (
		_w29616_,
		_w29617_,
		_w29618_
	);
	LUT2 #(
		.INIT('h8)
	) name25572 (
		_w29614_,
		_w29615_,
		_w29619_
	);
	LUT2 #(
		.INIT('h8)
	) name25573 (
		_w19996_,
		_w29613_,
		_w29620_
	);
	LUT2 #(
		.INIT('h8)
	) name25574 (
		_w29579_,
		_w29620_,
		_w29621_
	);
	LUT2 #(
		.INIT('h8)
	) name25575 (
		_w29618_,
		_w29619_,
		_w29622_
	);
	LUT2 #(
		.INIT('h8)
	) name25576 (
		_w29621_,
		_w29622_,
		_w29623_
	);
	LUT2 #(
		.INIT('h8)
	) name25577 (
		_w18731_,
		_w20106_,
		_w29624_
	);
	LUT2 #(
		.INIT('h8)
	) name25578 (
		_w29623_,
		_w29624_,
		_w29625_
	);
	LUT2 #(
		.INIT('h8)
	) name25579 (
		_w18800_,
		_w29625_,
		_w29626_
	);
	LUT2 #(
		.INIT('h2)
	) name25580 (
		_w28627_,
		_w29626_,
		_w29627_
	);
	LUT2 #(
		.INIT('h4)
	) name25581 (
		_w10289_,
		_w28572_,
		_w29628_
	);
	LUT2 #(
		.INIT('h1)
	) name25582 (
		_w13075_,
		_w28572_,
		_w29629_
	);
	LUT2 #(
		.INIT('h2)
	) name25583 (
		_w28997_,
		_w29628_,
		_w29630_
	);
	LUT2 #(
		.INIT('h4)
	) name25584 (
		_w29629_,
		_w29630_,
		_w29631_
	);
	LUT2 #(
		.INIT('h1)
	) name25585 (
		_w29570_,
		_w29571_,
		_w29632_
	);
	LUT2 #(
		.INIT('h4)
	) name25586 (
		_w29572_,
		_w29632_,
		_w29633_
	);
	LUT2 #(
		.INIT('h1)
	) name25587 (
		_w29573_,
		_w29574_,
		_w29634_
	);
	LUT2 #(
		.INIT('h8)
	) name25588 (
		_w29633_,
		_w29634_,
		_w29635_
	);
	LUT2 #(
		.INIT('h1)
	) name25589 (
		_w29556_,
		_w29627_,
		_w29636_
	);
	LUT2 #(
		.INIT('h8)
	) name25590 (
		_w29635_,
		_w29636_,
		_w29637_
	);
	LUT2 #(
		.INIT('h4)
	) name25591 (
		_w29631_,
		_w29637_,
		_w29638_
	);
	LUT2 #(
		.INIT('h4)
	) name25592 (
		_w29308_,
		_w29638_,
		_w29639_
	);
	LUT2 #(
		.INIT('h4)
	) name25593 (
		_w29569_,
		_w29639_,
		_w29640_
	);
	LUT2 #(
		.INIT('h4)
	) name25594 (
		_w29561_,
		_w29640_,
		_w29641_
	);
	LUT2 #(
		.INIT('h2)
	) name25595 (
		_w28719_,
		_w29641_,
		_w29642_
	);
	LUT2 #(
		.INIT('h4)
	) name25596 (
		_w28543_,
		_w28725_,
		_w29643_
	);
	LUT2 #(
		.INIT('h4)
	) name25597 (
		_w10289_,
		_w29643_,
		_w29644_
	);
	LUT2 #(
		.INIT('h2)
	) name25598 (
		_w13075_,
		_w28728_,
		_w29645_
	);
	LUT2 #(
		.INIT('h1)
	) name25599 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[9]/P0001 ,
		_w29646_
	);
	LUT2 #(
		.INIT('h2)
	) name25600 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[9]/P0001 ,
		_w29647_
	);
	LUT2 #(
		.INIT('h1)
	) name25601 (
		_w29646_,
		_w29647_,
		_w29648_
	);
	LUT2 #(
		.INIT('h8)
	) name25602 (
		_w28741_,
		_w29648_,
		_w29649_
	);
	LUT2 #(
		.INIT('h8)
	) name25603 (
		_w10116_,
		_w28652_,
		_w29650_
	);
	LUT2 #(
		.INIT('h2)
	) name25604 (
		_w10100_,
		_w28652_,
		_w29651_
	);
	LUT2 #(
		.INIT('h1)
	) name25605 (
		_w28660_,
		_w29650_,
		_w29652_
	);
	LUT2 #(
		.INIT('h4)
	) name25606 (
		_w29651_,
		_w29652_,
		_w29653_
	);
	LUT2 #(
		.INIT('h8)
	) name25607 (
		_w28739_,
		_w29653_,
		_w29654_
	);
	LUT2 #(
		.INIT('h8)
	) name25608 (
		_w10104_,
		_w28705_,
		_w29655_
	);
	LUT2 #(
		.INIT('h2)
	) name25609 (
		_w10108_,
		_w28705_,
		_w29656_
	);
	LUT2 #(
		.INIT('h1)
	) name25610 (
		_w29655_,
		_w29656_,
		_w29657_
	);
	LUT2 #(
		.INIT('h8)
	) name25611 (
		_w28735_,
		_w29657_,
		_w29658_
	);
	LUT2 #(
		.INIT('h2)
	) name25612 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w28545_,
		_w29659_
	);
	LUT2 #(
		.INIT('h1)
	) name25613 (
		_w29649_,
		_w29659_,
		_w29660_
	);
	LUT2 #(
		.INIT('h1)
	) name25614 (
		_w29654_,
		_w29658_,
		_w29661_
	);
	LUT2 #(
		.INIT('h8)
	) name25615 (
		_w29660_,
		_w29661_,
		_w29662_
	);
	LUT2 #(
		.INIT('h4)
	) name25616 (
		_w28725_,
		_w29662_,
		_w29663_
	);
	LUT2 #(
		.INIT('h4)
	) name25617 (
		_w29645_,
		_w29663_,
		_w29664_
	);
	LUT2 #(
		.INIT('h4)
	) name25618 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[9]/P0001 ,
		_w28543_,
		_w29665_
	);
	LUT2 #(
		.INIT('h1)
	) name25619 (
		_w28719_,
		_w29665_,
		_w29666_
	);
	LUT2 #(
		.INIT('h4)
	) name25620 (
		_w29644_,
		_w29666_,
		_w29667_
	);
	LUT2 #(
		.INIT('h4)
	) name25621 (
		_w29664_,
		_w29667_,
		_w29668_
	);
	LUT2 #(
		.INIT('h1)
	) name25622 (
		_w29642_,
		_w29668_,
		_w29669_
	);
	LUT2 #(
		.INIT('h4)
	) name25623 (
		_w18211_,
		_w28627_,
		_w29670_
	);
	LUT2 #(
		.INIT('h8)
	) name25624 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w17836_,
		_w29671_
	);
	LUT2 #(
		.INIT('h4)
	) name25625 (
		_w14551_,
		_w28561_,
		_w29672_
	);
	LUT2 #(
		.INIT('h1)
	) name25626 (
		_w28564_,
		_w29671_,
		_w29673_
	);
	LUT2 #(
		.INIT('h4)
	) name25627 (
		_w29672_,
		_w29673_,
		_w29674_
	);
	LUT2 #(
		.INIT('h2)
	) name25628 (
		_w28559_,
		_w29674_,
		_w29675_
	);
	LUT2 #(
		.INIT('h1)
	) name25629 (
		_w7202_,
		_w28589_,
		_w29676_
	);
	LUT2 #(
		.INIT('h1)
	) name25630 (
		_w7182_,
		_w28594_,
		_w29677_
	);
	LUT2 #(
		.INIT('h1)
	) name25631 (
		_w29676_,
		_w29677_,
		_w29678_
	);
	LUT2 #(
		.INIT('h8)
	) name25632 (
		_w29562_,
		_w29678_,
		_w29679_
	);
	LUT2 #(
		.INIT('h2)
	) name25633 (
		_w28577_,
		_w29679_,
		_w29680_
	);
	LUT2 #(
		.INIT('h1)
	) name25634 (
		_w29303_,
		_w29680_,
		_w29681_
	);
	LUT2 #(
		.INIT('h1)
	) name25635 (
		_w28569_,
		_w29681_,
		_w29682_
	);
	LUT2 #(
		.INIT('h1)
	) name25636 (
		_w12658_,
		_w28572_,
		_w29683_
	);
	LUT2 #(
		.INIT('h4)
	) name25637 (
		_w7340_,
		_w28572_,
		_w29684_
	);
	LUT2 #(
		.INIT('h2)
	) name25638 (
		_w28997_,
		_w29683_,
		_w29685_
	);
	LUT2 #(
		.INIT('h4)
	) name25639 (
		_w29684_,
		_w29685_,
		_w29686_
	);
	LUT2 #(
		.INIT('h8)
	) name25640 (
		_w12658_,
		_w28619_,
		_w29687_
	);
	LUT2 #(
		.INIT('h1)
	) name25641 (
		_w7112_,
		_w28634_,
		_w29688_
	);
	LUT2 #(
		.INIT('h8)
	) name25642 (
		_w7340_,
		_w28630_,
		_w29689_
	);
	LUT2 #(
		.INIT('h1)
	) name25643 (
		_w7164_,
		_w28624_,
		_w29690_
	);
	LUT2 #(
		.INIT('h1)
	) name25644 (
		_w7156_,
		_w28556_,
		_w29691_
	);
	LUT2 #(
		.INIT('h4)
	) name25645 (
		_w19840_,
		_w28636_,
		_w29692_
	);
	LUT2 #(
		.INIT('h1)
	) name25646 (
		_w29687_,
		_w29688_,
		_w29693_
	);
	LUT2 #(
		.INIT('h4)
	) name25647 (
		_w29689_,
		_w29693_,
		_w29694_
	);
	LUT2 #(
		.INIT('h1)
	) name25648 (
		_w29690_,
		_w29691_,
		_w29695_
	);
	LUT2 #(
		.INIT('h8)
	) name25649 (
		_w29694_,
		_w29695_,
		_w29696_
	);
	LUT2 #(
		.INIT('h4)
	) name25650 (
		_w29670_,
		_w29696_,
		_w29697_
	);
	LUT2 #(
		.INIT('h4)
	) name25651 (
		_w29692_,
		_w29697_,
		_w29698_
	);
	LUT2 #(
		.INIT('h4)
	) name25652 (
		_w29686_,
		_w29698_,
		_w29699_
	);
	LUT2 #(
		.INIT('h4)
	) name25653 (
		_w29308_,
		_w29699_,
		_w29700_
	);
	LUT2 #(
		.INIT('h4)
	) name25654 (
		_w29682_,
		_w29700_,
		_w29701_
	);
	LUT2 #(
		.INIT('h4)
	) name25655 (
		_w29675_,
		_w29701_,
		_w29702_
	);
	LUT2 #(
		.INIT('h2)
	) name25656 (
		_w28719_,
		_w29702_,
		_w29703_
	);
	LUT2 #(
		.INIT('h4)
	) name25657 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w28543_,
		_w29704_
	);
	LUT2 #(
		.INIT('h8)
	) name25658 (
		_w12658_,
		_w28729_,
		_w29705_
	);
	LUT2 #(
		.INIT('h8)
	) name25659 (
		_w7340_,
		_w28725_,
		_w29706_
	);
	LUT2 #(
		.INIT('h2)
	) name25660 (
		_w28725_,
		_w28727_,
		_w29707_
	);
	LUT2 #(
		.INIT('h8)
	) name25661 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[13]/P0001 ,
		_w28544_,
		_w29708_
	);
	LUT2 #(
		.INIT('h8)
	) name25662 (
		_w7194_,
		_w28652_,
		_w29709_
	);
	LUT2 #(
		.INIT('h2)
	) name25663 (
		_w7186_,
		_w28652_,
		_w29710_
	);
	LUT2 #(
		.INIT('h1)
	) name25664 (
		_w28660_,
		_w29709_,
		_w29711_
	);
	LUT2 #(
		.INIT('h4)
	) name25665 (
		_w29710_,
		_w29711_,
		_w29712_
	);
	LUT2 #(
		.INIT('h8)
	) name25666 (
		_w28739_,
		_w29712_,
		_w29713_
	);
	LUT2 #(
		.INIT('h8)
	) name25667 (
		_w7198_,
		_w28705_,
		_w29714_
	);
	LUT2 #(
		.INIT('h2)
	) name25668 (
		_w7190_,
		_w28705_,
		_w29715_
	);
	LUT2 #(
		.INIT('h1)
	) name25669 (
		_w29714_,
		_w29715_,
		_w29716_
	);
	LUT2 #(
		.INIT('h8)
	) name25670 (
		_w28735_,
		_w29716_,
		_w29717_
	);
	LUT2 #(
		.INIT('h1)
	) name25671 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[13]/P0001 ,
		_w29718_
	);
	LUT2 #(
		.INIT('h2)
	) name25672 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[13]/P0001 ,
		_w29719_
	);
	LUT2 #(
		.INIT('h1)
	) name25673 (
		_w29718_,
		_w29719_,
		_w29720_
	);
	LUT2 #(
		.INIT('h8)
	) name25674 (
		_w28741_,
		_w29720_,
		_w29721_
	);
	LUT2 #(
		.INIT('h1)
	) name25675 (
		_w29708_,
		_w29713_,
		_w29722_
	);
	LUT2 #(
		.INIT('h1)
	) name25676 (
		_w29717_,
		_w29721_,
		_w29723_
	);
	LUT2 #(
		.INIT('h8)
	) name25677 (
		_w29722_,
		_w29723_,
		_w29724_
	);
	LUT2 #(
		.INIT('h1)
	) name25678 (
		_w29707_,
		_w29724_,
		_w29725_
	);
	LUT2 #(
		.INIT('h1)
	) name25679 (
		_w28543_,
		_w29705_,
		_w29726_
	);
	LUT2 #(
		.INIT('h4)
	) name25680 (
		_w29725_,
		_w29726_,
		_w29727_
	);
	LUT2 #(
		.INIT('h4)
	) name25681 (
		_w29706_,
		_w29727_,
		_w29728_
	);
	LUT2 #(
		.INIT('h1)
	) name25682 (
		_w28719_,
		_w29704_,
		_w29729_
	);
	LUT2 #(
		.INIT('h4)
	) name25683 (
		_w29728_,
		_w29729_,
		_w29730_
	);
	LUT2 #(
		.INIT('h1)
	) name25684 (
		_w29703_,
		_w29730_,
		_w29731_
	);
	LUT2 #(
		.INIT('h1)
	) name25685 (
		_w8402_,
		_w28624_,
		_w29732_
	);
	LUT2 #(
		.INIT('h8)
	) name25686 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w23757_,
		_w29733_
	);
	LUT2 #(
		.INIT('h4)
	) name25687 (
		_w14424_,
		_w28561_,
		_w29734_
	);
	LUT2 #(
		.INIT('h1)
	) name25688 (
		_w28564_,
		_w29733_,
		_w29735_
	);
	LUT2 #(
		.INIT('h4)
	) name25689 (
		_w29734_,
		_w29735_,
		_w29736_
	);
	LUT2 #(
		.INIT('h2)
	) name25690 (
		_w28559_,
		_w29736_,
		_w29737_
	);
	LUT2 #(
		.INIT('h1)
	) name25691 (
		_w8354_,
		_w28594_,
		_w29738_
	);
	LUT2 #(
		.INIT('h1)
	) name25692 (
		_w8358_,
		_w28589_,
		_w29739_
	);
	LUT2 #(
		.INIT('h1)
	) name25693 (
		_w29738_,
		_w29739_,
		_w29740_
	);
	LUT2 #(
		.INIT('h8)
	) name25694 (
		_w29562_,
		_w29740_,
		_w29741_
	);
	LUT2 #(
		.INIT('h2)
	) name25695 (
		_w28577_,
		_w29741_,
		_w29742_
	);
	LUT2 #(
		.INIT('h1)
	) name25696 (
		_w29303_,
		_w29742_,
		_w29743_
	);
	LUT2 #(
		.INIT('h1)
	) name25697 (
		_w28569_,
		_w29743_,
		_w29744_
	);
	LUT2 #(
		.INIT('h1)
	) name25698 (
		_w8410_,
		_w28556_,
		_w29745_
	);
	LUT2 #(
		.INIT('h8)
	) name25699 (
		_w12590_,
		_w28619_,
		_w29746_
	);
	LUT2 #(
		.INIT('h2)
	) name25700 (
		_w18745_,
		_w18781_,
		_w29747_
	);
	LUT2 #(
		.INIT('h4)
	) name25701 (
		_w17995_,
		_w19792_,
		_w29748_
	);
	LUT2 #(
		.INIT('h1)
	) name25702 (
		_w18102_,
		_w18720_,
		_w29749_
	);
	LUT2 #(
		.INIT('h2)
	) name25703 (
		_w18088_,
		_w18898_,
		_w29750_
	);
	LUT2 #(
		.INIT('h2)
	) name25704 (
		_w18124_,
		_w19818_,
		_w29751_
	);
	LUT2 #(
		.INIT('h2)
	) name25705 (
		_w18099_,
		_w19857_,
		_w29752_
	);
	LUT2 #(
		.INIT('h2)
	) name25706 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w8402_,
		_w29753_
	);
	LUT2 #(
		.INIT('h2)
	) name25707 (
		_w18162_,
		_w18895_,
		_w29754_
	);
	LUT2 #(
		.INIT('h1)
	) name25708 (
		_w18189_,
		_w18907_,
		_w29755_
	);
	LUT2 #(
		.INIT('h1)
	) name25709 (
		_w17935_,
		_w18914_,
		_w29756_
	);
	LUT2 #(
		.INIT('h1)
	) name25710 (
		_w18912_,
		_w18991_,
		_w29757_
	);
	LUT2 #(
		.INIT('h1)
	) name25711 (
		_w18117_,
		_w18918_,
		_w29758_
	);
	LUT2 #(
		.INIT('h2)
	) name25712 (
		_w18740_,
		_w18775_,
		_w29759_
	);
	LUT2 #(
		.INIT('h4)
	) name25713 (
		_w17998_,
		_w18765_,
		_w29760_
	);
	LUT2 #(
		.INIT('h1)
	) name25714 (
		_w29753_,
		_w29755_,
		_w29761_
	);
	LUT2 #(
		.INIT('h1)
	) name25715 (
		_w29756_,
		_w29757_,
		_w29762_
	);
	LUT2 #(
		.INIT('h4)
	) name25716 (
		_w29758_,
		_w29762_,
		_w29763_
	);
	LUT2 #(
		.INIT('h8)
	) name25717 (
		_w19874_,
		_w29761_,
		_w29764_
	);
	LUT2 #(
		.INIT('h1)
	) name25718 (
		_w29747_,
		_w29749_,
		_w29765_
	);
	LUT2 #(
		.INIT('h1)
	) name25719 (
		_w29750_,
		_w29751_,
		_w29766_
	);
	LUT2 #(
		.INIT('h1)
	) name25720 (
		_w29752_,
		_w29754_,
		_w29767_
	);
	LUT2 #(
		.INIT('h1)
	) name25721 (
		_w29759_,
		_w29760_,
		_w29768_
	);
	LUT2 #(
		.INIT('h8)
	) name25722 (
		_w29767_,
		_w29768_,
		_w29769_
	);
	LUT2 #(
		.INIT('h8)
	) name25723 (
		_w29765_,
		_w29766_,
		_w29770_
	);
	LUT2 #(
		.INIT('h8)
	) name25724 (
		_w29763_,
		_w29764_,
		_w29771_
	);
	LUT2 #(
		.INIT('h4)
	) name25725 (
		_w18085_,
		_w19854_,
		_w29772_
	);
	LUT2 #(
		.INIT('h8)
	) name25726 (
		_w29771_,
		_w29772_,
		_w29773_
	);
	LUT2 #(
		.INIT('h8)
	) name25727 (
		_w29769_,
		_w29770_,
		_w29774_
	);
	LUT2 #(
		.INIT('h8)
	) name25728 (
		_w29773_,
		_w29774_,
		_w29775_
	);
	LUT2 #(
		.INIT('h8)
	) name25729 (
		_w29748_,
		_w29775_,
		_w29776_
	);
	LUT2 #(
		.INIT('h2)
	) name25730 (
		_w28636_,
		_w29776_,
		_w29777_
	);
	LUT2 #(
		.INIT('h8)
	) name25731 (
		_w8460_,
		_w28630_,
		_w29778_
	);
	LUT2 #(
		.INIT('h1)
	) name25732 (
		_w8385_,
		_w28634_,
		_w29779_
	);
	LUT2 #(
		.INIT('h2)
	) name25733 (
		_w17921_,
		_w18117_,
		_w29780_
	);
	LUT2 #(
		.INIT('h2)
	) name25734 (
		_w18100_,
		_w18121_,
		_w29781_
	);
	LUT2 #(
		.INIT('h8)
	) name25735 (
		_w18162_,
		_w18179_,
		_w29782_
	);
	LUT2 #(
		.INIT('h8)
	) name25736 (
		_w18124_,
		_w18157_,
		_w29783_
	);
	LUT2 #(
		.INIT('h8)
	) name25737 (
		_w18107_,
		_w18171_,
		_w29784_
	);
	LUT2 #(
		.INIT('h8)
	) name25738 (
		_w17915_,
		_w18111_,
		_w29785_
	);
	LUT2 #(
		.INIT('h1)
	) name25739 (
		_w29782_,
		_w29783_,
		_w29786_
	);
	LUT2 #(
		.INIT('h1)
	) name25740 (
		_w29784_,
		_w29785_,
		_w29787_
	);
	LUT2 #(
		.INIT('h8)
	) name25741 (
		_w29786_,
		_w29787_,
		_w29788_
	);
	LUT2 #(
		.INIT('h1)
	) name25742 (
		_w17931_,
		_w29788_,
		_w29789_
	);
	LUT2 #(
		.INIT('h4)
	) name25743 (
		_w18133_,
		_w18184_,
		_w29790_
	);
	LUT2 #(
		.INIT('h1)
	) name25744 (
		_w17935_,
		_w18091_,
		_w29791_
	);
	LUT2 #(
		.INIT('h2)
	) name25745 (
		_w18147_,
		_w18175_,
		_w29792_
	);
	LUT2 #(
		.INIT('h8)
	) name25746 (
		_w17945_,
		_w18153_,
		_w29793_
	);
	LUT2 #(
		.INIT('h2)
	) name25747 (
		_w19996_,
		_w29793_,
		_w29794_
	);
	LUT2 #(
		.INIT('h8)
	) name25748 (
		_w18076_,
		_w29794_,
		_w29795_
	);
	LUT2 #(
		.INIT('h2)
	) name25749 (
		_w17945_,
		_w18047_,
		_w29796_
	);
	LUT2 #(
		.INIT('h8)
	) name25750 (
		_w18131_,
		_w18188_,
		_w29797_
	);
	LUT2 #(
		.INIT('h8)
	) name25751 (
		_w18790_,
		_w19731_,
		_w29798_
	);
	LUT2 #(
		.INIT('h2)
	) name25752 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w8410_,
		_w29799_
	);
	LUT2 #(
		.INIT('h4)
	) name25753 (
		_w18129_,
		_w18158_,
		_w29800_
	);
	LUT2 #(
		.INIT('h8)
	) name25754 (
		_w18128_,
		_w18157_,
		_w29801_
	);
	LUT2 #(
		.INIT('h4)
	) name25755 (
		_w18167_,
		_w18178_,
		_w29802_
	);
	LUT2 #(
		.INIT('h8)
	) name25756 (
		_w18103_,
		_w18120_,
		_w29803_
	);
	LUT2 #(
		.INIT('h8)
	) name25757 (
		_w18103_,
		_w18119_,
		_w29804_
	);
	LUT2 #(
		.INIT('h2)
	) name25758 (
		_w18088_,
		_w19979_,
		_w29805_
	);
	LUT2 #(
		.INIT('h8)
	) name25759 (
		_w18132_,
		_w18188_,
		_w29806_
	);
	LUT2 #(
		.INIT('h4)
	) name25760 (
		_w18108_,
		_w18136_,
		_w29807_
	);
	LUT2 #(
		.INIT('h2)
	) name25761 (
		_w18148_,
		_w18175_,
		_w29808_
	);
	LUT2 #(
		.INIT('h8)
	) name25762 (
		_w17915_,
		_w18116_,
		_w29809_
	);
	LUT2 #(
		.INIT('h8)
	) name25763 (
		_w18166_,
		_w18179_,
		_w29810_
	);
	LUT2 #(
		.INIT('h8)
	) name25764 (
		_w18106_,
		_w18172_,
		_w29811_
	);
	LUT2 #(
		.INIT('h1)
	) name25765 (
		_w18060_,
		_w29799_,
		_w29812_
	);
	LUT2 #(
		.INIT('h1)
	) name25766 (
		_w29780_,
		_w29800_,
		_w29813_
	);
	LUT2 #(
		.INIT('h1)
	) name25767 (
		_w29802_,
		_w29803_,
		_w29814_
	);
	LUT2 #(
		.INIT('h1)
	) name25768 (
		_w29806_,
		_w29811_,
		_w29815_
	);
	LUT2 #(
		.INIT('h8)
	) name25769 (
		_w29814_,
		_w29815_,
		_w29816_
	);
	LUT2 #(
		.INIT('h8)
	) name25770 (
		_w29812_,
		_w29813_,
		_w29817_
	);
	LUT2 #(
		.INIT('h1)
	) name25771 (
		_w18065_,
		_w29797_,
		_w29818_
	);
	LUT2 #(
		.INIT('h1)
	) name25772 (
		_w29801_,
		_w29804_,
		_w29819_
	);
	LUT2 #(
		.INIT('h1)
	) name25773 (
		_w29808_,
		_w29809_,
		_w29820_
	);
	LUT2 #(
		.INIT('h4)
	) name25774 (
		_w29810_,
		_w29820_,
		_w29821_
	);
	LUT2 #(
		.INIT('h8)
	) name25775 (
		_w29818_,
		_w29819_,
		_w29822_
	);
	LUT2 #(
		.INIT('h8)
	) name25776 (
		_w29816_,
		_w29817_,
		_w29823_
	);
	LUT2 #(
		.INIT('h1)
	) name25777 (
		_w29781_,
		_w29790_,
		_w29824_
	);
	LUT2 #(
		.INIT('h1)
	) name25778 (
		_w29791_,
		_w29792_,
		_w29825_
	);
	LUT2 #(
		.INIT('h4)
	) name25779 (
		_w29807_,
		_w29825_,
		_w29826_
	);
	LUT2 #(
		.INIT('h8)
	) name25780 (
		_w29823_,
		_w29824_,
		_w29827_
	);
	LUT2 #(
		.INIT('h8)
	) name25781 (
		_w29821_,
		_w29822_,
		_w29828_
	);
	LUT2 #(
		.INIT('h2)
	) name25782 (
		_w18041_,
		_w29796_,
		_w29829_
	);
	LUT2 #(
		.INIT('h4)
	) name25783 (
		_w29805_,
		_w29829_,
		_w29830_
	);
	LUT2 #(
		.INIT('h8)
	) name25784 (
		_w29827_,
		_w29828_,
		_w29831_
	);
	LUT2 #(
		.INIT('h8)
	) name25785 (
		_w17984_,
		_w29826_,
		_w29832_
	);
	LUT2 #(
		.INIT('h4)
	) name25786 (
		_w29789_,
		_w29832_,
		_w29833_
	);
	LUT2 #(
		.INIT('h8)
	) name25787 (
		_w29830_,
		_w29831_,
		_w29834_
	);
	LUT2 #(
		.INIT('h8)
	) name25788 (
		_w19999_,
		_w29834_,
		_w29835_
	);
	LUT2 #(
		.INIT('h8)
	) name25789 (
		_w29795_,
		_w29833_,
		_w29836_
	);
	LUT2 #(
		.INIT('h8)
	) name25790 (
		_w29798_,
		_w29836_,
		_w29837_
	);
	LUT2 #(
		.INIT('h8)
	) name25791 (
		_w18799_,
		_w29835_,
		_w29838_
	);
	LUT2 #(
		.INIT('h8)
	) name25792 (
		_w29837_,
		_w29838_,
		_w29839_
	);
	LUT2 #(
		.INIT('h2)
	) name25793 (
		_w28627_,
		_w29839_,
		_w29840_
	);
	LUT2 #(
		.INIT('h1)
	) name25794 (
		_w12590_,
		_w28572_,
		_w29841_
	);
	LUT2 #(
		.INIT('h4)
	) name25795 (
		_w8460_,
		_w28572_,
		_w29842_
	);
	LUT2 #(
		.INIT('h2)
	) name25796 (
		_w28997_,
		_w29841_,
		_w29843_
	);
	LUT2 #(
		.INIT('h4)
	) name25797 (
		_w29842_,
		_w29843_,
		_w29844_
	);
	LUT2 #(
		.INIT('h1)
	) name25798 (
		_w29746_,
		_w29778_,
		_w29845_
	);
	LUT2 #(
		.INIT('h4)
	) name25799 (
		_w29779_,
		_w29845_,
		_w29846_
	);
	LUT2 #(
		.INIT('h1)
	) name25800 (
		_w29732_,
		_w29745_,
		_w29847_
	);
	LUT2 #(
		.INIT('h8)
	) name25801 (
		_w29846_,
		_w29847_,
		_w29848_
	);
	LUT2 #(
		.INIT('h1)
	) name25802 (
		_w29777_,
		_w29840_,
		_w29849_
	);
	LUT2 #(
		.INIT('h8)
	) name25803 (
		_w29848_,
		_w29849_,
		_w29850_
	);
	LUT2 #(
		.INIT('h4)
	) name25804 (
		_w29844_,
		_w29850_,
		_w29851_
	);
	LUT2 #(
		.INIT('h4)
	) name25805 (
		_w29308_,
		_w29851_,
		_w29852_
	);
	LUT2 #(
		.INIT('h4)
	) name25806 (
		_w29744_,
		_w29852_,
		_w29853_
	);
	LUT2 #(
		.INIT('h4)
	) name25807 (
		_w29737_,
		_w29853_,
		_w29854_
	);
	LUT2 #(
		.INIT('h2)
	) name25808 (
		_w28719_,
		_w29854_,
		_w29855_
	);
	LUT2 #(
		.INIT('h4)
	) name25809 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		_w28543_,
		_w29856_
	);
	LUT2 #(
		.INIT('h8)
	) name25810 (
		_w12590_,
		_w28729_,
		_w29857_
	);
	LUT2 #(
		.INIT('h8)
	) name25811 (
		_w8460_,
		_w28725_,
		_w29858_
	);
	LUT2 #(
		.INIT('h8)
	) name25812 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[11]/P0001 ,
		_w28544_,
		_w29859_
	);
	LUT2 #(
		.INIT('h8)
	) name25813 (
		_w8346_,
		_w28652_,
		_w29860_
	);
	LUT2 #(
		.INIT('h2)
	) name25814 (
		_w8350_,
		_w28652_,
		_w29861_
	);
	LUT2 #(
		.INIT('h1)
	) name25815 (
		_w28660_,
		_w29860_,
		_w29862_
	);
	LUT2 #(
		.INIT('h4)
	) name25816 (
		_w29861_,
		_w29862_,
		_w29863_
	);
	LUT2 #(
		.INIT('h8)
	) name25817 (
		_w28739_,
		_w29863_,
		_w29864_
	);
	LUT2 #(
		.INIT('h8)
	) name25818 (
		_w8338_,
		_w28705_,
		_w29865_
	);
	LUT2 #(
		.INIT('h2)
	) name25819 (
		_w8342_,
		_w28705_,
		_w29866_
	);
	LUT2 #(
		.INIT('h1)
	) name25820 (
		_w29865_,
		_w29866_,
		_w29867_
	);
	LUT2 #(
		.INIT('h8)
	) name25821 (
		_w28735_,
		_w29867_,
		_w29868_
	);
	LUT2 #(
		.INIT('h1)
	) name25822 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[11]/P0001 ,
		_w29869_
	);
	LUT2 #(
		.INIT('h2)
	) name25823 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[11]/P0001 ,
		_w29870_
	);
	LUT2 #(
		.INIT('h1)
	) name25824 (
		_w29869_,
		_w29870_,
		_w29871_
	);
	LUT2 #(
		.INIT('h8)
	) name25825 (
		_w28741_,
		_w29871_,
		_w29872_
	);
	LUT2 #(
		.INIT('h1)
	) name25826 (
		_w29859_,
		_w29864_,
		_w29873_
	);
	LUT2 #(
		.INIT('h1)
	) name25827 (
		_w29868_,
		_w29872_,
		_w29874_
	);
	LUT2 #(
		.INIT('h8)
	) name25828 (
		_w29873_,
		_w29874_,
		_w29875_
	);
	LUT2 #(
		.INIT('h1)
	) name25829 (
		_w29707_,
		_w29875_,
		_w29876_
	);
	LUT2 #(
		.INIT('h1)
	) name25830 (
		_w28543_,
		_w29857_,
		_w29877_
	);
	LUT2 #(
		.INIT('h4)
	) name25831 (
		_w29876_,
		_w29877_,
		_w29878_
	);
	LUT2 #(
		.INIT('h4)
	) name25832 (
		_w29858_,
		_w29878_,
		_w29879_
	);
	LUT2 #(
		.INIT('h1)
	) name25833 (
		_w28719_,
		_w29856_,
		_w29880_
	);
	LUT2 #(
		.INIT('h4)
	) name25834 (
		_w29879_,
		_w29880_,
		_w29881_
	);
	LUT2 #(
		.INIT('h1)
	) name25835 (
		_w29855_,
		_w29881_,
		_w29882_
	);
	LUT2 #(
		.INIT('h1)
	) name25836 (
		_w7784_,
		_w28634_,
		_w29883_
	);
	LUT2 #(
		.INIT('h8)
	) name25837 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w19848_,
		_w29884_
	);
	LUT2 #(
		.INIT('h4)
	) name25838 (
		_w20053_,
		_w28561_,
		_w29885_
	);
	LUT2 #(
		.INIT('h1)
	) name25839 (
		_w28564_,
		_w29884_,
		_w29886_
	);
	LUT2 #(
		.INIT('h4)
	) name25840 (
		_w29885_,
		_w29886_,
		_w29887_
	);
	LUT2 #(
		.INIT('h2)
	) name25841 (
		_w28559_,
		_w29887_,
		_w29888_
	);
	LUT2 #(
		.INIT('h1)
	) name25842 (
		_w7753_,
		_w28594_,
		_w29889_
	);
	LUT2 #(
		.INIT('h1)
	) name25843 (
		_w7737_,
		_w28589_,
		_w29890_
	);
	LUT2 #(
		.INIT('h1)
	) name25844 (
		_w29889_,
		_w29890_,
		_w29891_
	);
	LUT2 #(
		.INIT('h8)
	) name25845 (
		_w29562_,
		_w29891_,
		_w29892_
	);
	LUT2 #(
		.INIT('h2)
	) name25846 (
		_w28577_,
		_w29892_,
		_w29893_
	);
	LUT2 #(
		.INIT('h1)
	) name25847 (
		_w29303_,
		_w29893_,
		_w29894_
	);
	LUT2 #(
		.INIT('h1)
	) name25848 (
		_w28569_,
		_w29894_,
		_w29895_
	);
	LUT2 #(
		.INIT('h8)
	) name25849 (
		_w7859_,
		_w28630_,
		_w29896_
	);
	LUT2 #(
		.INIT('h4)
	) name25850 (
		_w19895_,
		_w28636_,
		_w29897_
	);
	LUT2 #(
		.INIT('h1)
	) name25851 (
		_w18133_,
		_w18919_,
		_w29898_
	);
	LUT2 #(
		.INIT('h1)
	) name25852 (
		_w18123_,
		_w18180_,
		_w29899_
	);
	LUT2 #(
		.INIT('h8)
	) name25853 (
		_w18099_,
		_w18157_,
		_w29900_
	);
	LUT2 #(
		.INIT('h8)
	) name25854 (
		_w18090_,
		_w18111_,
		_w29901_
	);
	LUT2 #(
		.INIT('h1)
	) name25855 (
		_w29900_,
		_w29901_,
		_w29902_
	);
	LUT2 #(
		.INIT('h4)
	) name25856 (
		_w29899_,
		_w29902_,
		_w29903_
	);
	LUT2 #(
		.INIT('h2)
	) name25857 (
		_w17931_,
		_w29903_,
		_w29904_
	);
	LUT2 #(
		.INIT('h4)
	) name25858 (
		_w18159_,
		_w18741_,
		_w29905_
	);
	LUT2 #(
		.INIT('h4)
	) name25859 (
		_w18091_,
		_w18749_,
		_w29906_
	);
	LUT2 #(
		.INIT('h4)
	) name25860 (
		_w18180_,
		_w18746_,
		_w29907_
	);
	LUT2 #(
		.INIT('h1)
	) name25861 (
		_w17922_,
		_w19864_,
		_w29908_
	);
	LUT2 #(
		.INIT('h4)
	) name25862 (
		_w18121_,
		_w18752_,
		_w29909_
	);
	LUT2 #(
		.INIT('h1)
	) name25863 (
		_w17980_,
		_w19856_,
		_w29910_
	);
	LUT2 #(
		.INIT('h2)
	) name25864 (
		_w17945_,
		_w29910_,
		_w29911_
	);
	LUT2 #(
		.INIT('h1)
	) name25865 (
		_w17981_,
		_w18719_,
		_w29912_
	);
	LUT2 #(
		.INIT('h2)
	) name25866 (
		_w17839_,
		_w29912_,
		_w29913_
	);
	LUT2 #(
		.INIT('h1)
	) name25867 (
		_w18046_,
		_w29913_,
		_w29914_
	);
	LUT2 #(
		.INIT('h1)
	) name25868 (
		_w17938_,
		_w29914_,
		_w29915_
	);
	LUT2 #(
		.INIT('h1)
	) name25869 (
		_w17924_,
		_w18149_,
		_w29916_
	);
	LUT2 #(
		.INIT('h8)
	) name25870 (
		_w18089_,
		_w18905_,
		_w29917_
	);
	LUT2 #(
		.INIT('h2)
	) name25871 (
		_w18765_,
		_w19979_,
		_w29918_
	);
	LUT2 #(
		.INIT('h2)
	) name25872 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7809_,
		_w29919_
	);
	LUT2 #(
		.INIT('h8)
	) name25873 (
		_w18158_,
		_w18742_,
		_w29920_
	);
	LUT2 #(
		.INIT('h1)
	) name25874 (
		_w18108_,
		_w18915_,
		_w29921_
	);
	LUT2 #(
		.INIT('h1)
	) name25875 (
		_w29917_,
		_w29919_,
		_w29922_
	);
	LUT2 #(
		.INIT('h4)
	) name25876 (
		_w29920_,
		_w29922_,
		_w29923_
	);
	LUT2 #(
		.INIT('h4)
	) name25877 (
		_w18783_,
		_w29923_,
		_w29924_
	);
	LUT2 #(
		.INIT('h1)
	) name25878 (
		_w29898_,
		_w29905_,
		_w29925_
	);
	LUT2 #(
		.INIT('h1)
	) name25879 (
		_w29906_,
		_w29907_,
		_w29926_
	);
	LUT2 #(
		.INIT('h1)
	) name25880 (
		_w29908_,
		_w29909_,
		_w29927_
	);
	LUT2 #(
		.INIT('h4)
	) name25881 (
		_w29921_,
		_w29927_,
		_w29928_
	);
	LUT2 #(
		.INIT('h8)
	) name25882 (
		_w29925_,
		_w29926_,
		_w29929_
	);
	LUT2 #(
		.INIT('h4)
	) name25883 (
		_w29911_,
		_w29924_,
		_w29930_
	);
	LUT2 #(
		.INIT('h1)
	) name25884 (
		_w29916_,
		_w29918_,
		_w29931_
	);
	LUT2 #(
		.INIT('h8)
	) name25885 (
		_w29930_,
		_w29931_,
		_w29932_
	);
	LUT2 #(
		.INIT('h8)
	) name25886 (
		_w29928_,
		_w29929_,
		_w29933_
	);
	LUT2 #(
		.INIT('h8)
	) name25887 (
		_w18042_,
		_w29579_,
		_w29934_
	);
	LUT2 #(
		.INIT('h4)
	) name25888 (
		_w29904_,
		_w29934_,
		_w29935_
	);
	LUT2 #(
		.INIT('h8)
	) name25889 (
		_w29932_,
		_w29933_,
		_w29936_
	);
	LUT2 #(
		.INIT('h2)
	) name25890 (
		_w19997_,
		_w29915_,
		_w29937_
	);
	LUT2 #(
		.INIT('h8)
	) name25891 (
		_w29936_,
		_w29937_,
		_w29938_
	);
	LUT2 #(
		.INIT('h8)
	) name25892 (
		_w19716_,
		_w29935_,
		_w29939_
	);
	LUT2 #(
		.INIT('h8)
	) name25893 (
		_w29798_,
		_w29939_,
		_w29940_
	);
	LUT2 #(
		.INIT('h8)
	) name25894 (
		_w29938_,
		_w29940_,
		_w29941_
	);
	LUT2 #(
		.INIT('h8)
	) name25895 (
		_w18800_,
		_w29941_,
		_w29942_
	);
	LUT2 #(
		.INIT('h2)
	) name25896 (
		_w28627_,
		_w29942_,
		_w29943_
	);
	LUT2 #(
		.INIT('h1)
	) name25897 (
		_w7801_,
		_w28624_,
		_w29944_
	);
	LUT2 #(
		.INIT('h1)
	) name25898 (
		_w7809_,
		_w28556_,
		_w29945_
	);
	LUT2 #(
		.INIT('h8)
	) name25899 (
		_w12556_,
		_w28619_,
		_w29946_
	);
	LUT2 #(
		.INIT('h1)
	) name25900 (
		_w12556_,
		_w28572_,
		_w29947_
	);
	LUT2 #(
		.INIT('h4)
	) name25901 (
		_w7859_,
		_w28572_,
		_w29948_
	);
	LUT2 #(
		.INIT('h2)
	) name25902 (
		_w28997_,
		_w29947_,
		_w29949_
	);
	LUT2 #(
		.INIT('h4)
	) name25903 (
		_w29948_,
		_w29949_,
		_w29950_
	);
	LUT2 #(
		.INIT('h1)
	) name25904 (
		_w29883_,
		_w29896_,
		_w29951_
	);
	LUT2 #(
		.INIT('h4)
	) name25905 (
		_w29946_,
		_w29951_,
		_w29952_
	);
	LUT2 #(
		.INIT('h1)
	) name25906 (
		_w29897_,
		_w29944_,
		_w29953_
	);
	LUT2 #(
		.INIT('h4)
	) name25907 (
		_w29945_,
		_w29953_,
		_w29954_
	);
	LUT2 #(
		.INIT('h8)
	) name25908 (
		_w29952_,
		_w29954_,
		_w29955_
	);
	LUT2 #(
		.INIT('h4)
	) name25909 (
		_w29943_,
		_w29955_,
		_w29956_
	);
	LUT2 #(
		.INIT('h4)
	) name25910 (
		_w29950_,
		_w29956_,
		_w29957_
	);
	LUT2 #(
		.INIT('h4)
	) name25911 (
		_w29308_,
		_w29957_,
		_w29958_
	);
	LUT2 #(
		.INIT('h4)
	) name25912 (
		_w29895_,
		_w29958_,
		_w29959_
	);
	LUT2 #(
		.INIT('h4)
	) name25913 (
		_w29888_,
		_w29959_,
		_w29960_
	);
	LUT2 #(
		.INIT('h2)
	) name25914 (
		_w28719_,
		_w29960_,
		_w29961_
	);
	LUT2 #(
		.INIT('h4)
	) name25915 (
		_w7859_,
		_w29643_,
		_w29962_
	);
	LUT2 #(
		.INIT('h2)
	) name25916 (
		_w12556_,
		_w28728_,
		_w29963_
	);
	LUT2 #(
		.INIT('h1)
	) name25917 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001 ,
		_w29964_
	);
	LUT2 #(
		.INIT('h2)
	) name25918 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001 ,
		_w29965_
	);
	LUT2 #(
		.INIT('h1)
	) name25919 (
		_w29964_,
		_w29965_,
		_w29966_
	);
	LUT2 #(
		.INIT('h8)
	) name25920 (
		_w28741_,
		_w29966_,
		_w29967_
	);
	LUT2 #(
		.INIT('h8)
	) name25921 (
		_w7757_,
		_w28652_,
		_w29968_
	);
	LUT2 #(
		.INIT('h2)
	) name25922 (
		_w7741_,
		_w28652_,
		_w29969_
	);
	LUT2 #(
		.INIT('h1)
	) name25923 (
		_w28660_,
		_w29968_,
		_w29970_
	);
	LUT2 #(
		.INIT('h4)
	) name25924 (
		_w29969_,
		_w29970_,
		_w29971_
	);
	LUT2 #(
		.INIT('h8)
	) name25925 (
		_w28739_,
		_w29971_,
		_w29972_
	);
	LUT2 #(
		.INIT('h8)
	) name25926 (
		_w7745_,
		_w28705_,
		_w29973_
	);
	LUT2 #(
		.INIT('h2)
	) name25927 (
		_w7749_,
		_w28705_,
		_w29974_
	);
	LUT2 #(
		.INIT('h1)
	) name25928 (
		_w29973_,
		_w29974_,
		_w29975_
	);
	LUT2 #(
		.INIT('h8)
	) name25929 (
		_w28735_,
		_w29975_,
		_w29976_
	);
	LUT2 #(
		.INIT('h2)
	) name25930 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		_w28545_,
		_w29977_
	);
	LUT2 #(
		.INIT('h1)
	) name25931 (
		_w29967_,
		_w29977_,
		_w29978_
	);
	LUT2 #(
		.INIT('h1)
	) name25932 (
		_w29972_,
		_w29976_,
		_w29979_
	);
	LUT2 #(
		.INIT('h8)
	) name25933 (
		_w29978_,
		_w29979_,
		_w29980_
	);
	LUT2 #(
		.INIT('h4)
	) name25934 (
		_w28725_,
		_w29980_,
		_w29981_
	);
	LUT2 #(
		.INIT('h4)
	) name25935 (
		_w29963_,
		_w29981_,
		_w29982_
	);
	LUT2 #(
		.INIT('h4)
	) name25936 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[10]/P0001 ,
		_w28543_,
		_w29983_
	);
	LUT2 #(
		.INIT('h1)
	) name25937 (
		_w28719_,
		_w29983_,
		_w29984_
	);
	LUT2 #(
		.INIT('h4)
	) name25938 (
		_w29962_,
		_w29984_,
		_w29985_
	);
	LUT2 #(
		.INIT('h4)
	) name25939 (
		_w29982_,
		_w29985_,
		_w29986_
	);
	LUT2 #(
		.INIT('h1)
	) name25940 (
		_w29961_,
		_w29986_,
		_w29987_
	);
	LUT2 #(
		.INIT('h8)
	) name25941 (
		_w19504_,
		_w28660_,
		_w29988_
	);
	LUT2 #(
		.INIT('h1)
	) name25942 (
		_w29653_,
		_w29988_,
		_w29989_
	);
	LUT2 #(
		.INIT('h1)
	) name25943 (
		_w28649_,
		_w29989_,
		_w29990_
	);
	LUT2 #(
		.INIT('h8)
	) name25944 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[9]/P0001 ,
		_w28649_,
		_w29991_
	);
	LUT2 #(
		.INIT('h1)
	) name25945 (
		_w29990_,
		_w29991_,
		_w29992_
	);
	LUT2 #(
		.INIT('h1)
	) name25946 (
		_w28550_,
		_w29992_,
		_w29993_
	);
	LUT2 #(
		.INIT('h2)
	) name25947 (
		_w28550_,
		_w29641_,
		_w29994_
	);
	LUT2 #(
		.INIT('h1)
	) name25948 (
		_w29993_,
		_w29994_,
		_w29995_
	);
	LUT2 #(
		.INIT('h8)
	) name25949 (
		_w17836_,
		_w28660_,
		_w29996_
	);
	LUT2 #(
		.INIT('h1)
	) name25950 (
		_w29712_,
		_w29996_,
		_w29997_
	);
	LUT2 #(
		.INIT('h1)
	) name25951 (
		_w28649_,
		_w29997_,
		_w29998_
	);
	LUT2 #(
		.INIT('h8)
	) name25952 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[13]/P0001 ,
		_w28649_,
		_w29999_
	);
	LUT2 #(
		.INIT('h1)
	) name25953 (
		_w29998_,
		_w29999_,
		_w30000_
	);
	LUT2 #(
		.INIT('h1)
	) name25954 (
		_w28550_,
		_w30000_,
		_w30001_
	);
	LUT2 #(
		.INIT('h2)
	) name25955 (
		_w28550_,
		_w29702_,
		_w30002_
	);
	LUT2 #(
		.INIT('h1)
	) name25956 (
		_w30001_,
		_w30002_,
		_w30003_
	);
	LUT2 #(
		.INIT('h8)
	) name25957 (
		_w23757_,
		_w28660_,
		_w30004_
	);
	LUT2 #(
		.INIT('h1)
	) name25958 (
		_w29863_,
		_w30004_,
		_w30005_
	);
	LUT2 #(
		.INIT('h1)
	) name25959 (
		_w28649_,
		_w30005_,
		_w30006_
	);
	LUT2 #(
		.INIT('h8)
	) name25960 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[11]/P0001 ,
		_w28649_,
		_w30007_
	);
	LUT2 #(
		.INIT('h1)
	) name25961 (
		_w30006_,
		_w30007_,
		_w30008_
	);
	LUT2 #(
		.INIT('h1)
	) name25962 (
		_w28550_,
		_w30008_,
		_w30009_
	);
	LUT2 #(
		.INIT('h2)
	) name25963 (
		_w28550_,
		_w29854_,
		_w30010_
	);
	LUT2 #(
		.INIT('h1)
	) name25964 (
		_w30009_,
		_w30010_,
		_w30011_
	);
	LUT2 #(
		.INIT('h8)
	) name25965 (
		_w19848_,
		_w28660_,
		_w30012_
	);
	LUT2 #(
		.INIT('h1)
	) name25966 (
		_w29971_,
		_w30012_,
		_w30013_
	);
	LUT2 #(
		.INIT('h1)
	) name25967 (
		_w28649_,
		_w30013_,
		_w30014_
	);
	LUT2 #(
		.INIT('h8)
	) name25968 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[10]/P0001 ,
		_w28649_,
		_w30015_
	);
	LUT2 #(
		.INIT('h1)
	) name25969 (
		_w30014_,
		_w30015_,
		_w30016_
	);
	LUT2 #(
		.INIT('h1)
	) name25970 (
		_w28550_,
		_w30016_,
		_w30017_
	);
	LUT2 #(
		.INIT('h2)
	) name25971 (
		_w28550_,
		_w29960_,
		_w30018_
	);
	LUT2 #(
		.INIT('h1)
	) name25972 (
		_w30017_,
		_w30018_,
		_w30019_
	);
	LUT2 #(
		.INIT('h8)
	) name25973 (
		_w12624_,
		_w28729_,
		_w30020_
	);
	LUT2 #(
		.INIT('h8)
	) name25974 (
		_w9178_,
		_w28725_,
		_w30021_
	);
	LUT2 #(
		.INIT('h8)
	) name25975 (
		_w9064_,
		_w28705_,
		_w30022_
	);
	LUT2 #(
		.INIT('h2)
	) name25976 (
		_w9068_,
		_w28705_,
		_w30023_
	);
	LUT2 #(
		.INIT('h1)
	) name25977 (
		_w30022_,
		_w30023_,
		_w30024_
	);
	LUT2 #(
		.INIT('h8)
	) name25978 (
		_w28735_,
		_w30024_,
		_w30025_
	);
	LUT2 #(
		.INIT('h8)
	) name25979 (
		_w9076_,
		_w28652_,
		_w30026_
	);
	LUT2 #(
		.INIT('h2)
	) name25980 (
		_w9060_,
		_w28652_,
		_w30027_
	);
	LUT2 #(
		.INIT('h1)
	) name25981 (
		_w28660_,
		_w30026_,
		_w30028_
	);
	LUT2 #(
		.INIT('h4)
	) name25982 (
		_w30027_,
		_w30028_,
		_w30029_
	);
	LUT2 #(
		.INIT('h8)
	) name25983 (
		_w28739_,
		_w30029_,
		_w30030_
	);
	LUT2 #(
		.INIT('h1)
	) name25984 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[12]/P0001 ,
		_w30031_
	);
	LUT2 #(
		.INIT('h2)
	) name25985 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[12]/P0001 ,
		_w30032_
	);
	LUT2 #(
		.INIT('h1)
	) name25986 (
		_w30031_,
		_w30032_,
		_w30033_
	);
	LUT2 #(
		.INIT('h8)
	) name25987 (
		_w28741_,
		_w30033_,
		_w30034_
	);
	LUT2 #(
		.INIT('h1)
	) name25988 (
		_w30025_,
		_w30030_,
		_w30035_
	);
	LUT2 #(
		.INIT('h4)
	) name25989 (
		_w30034_,
		_w30035_,
		_w30036_
	);
	LUT2 #(
		.INIT('h4)
	) name25990 (
		_w30020_,
		_w30036_,
		_w30037_
	);
	LUT2 #(
		.INIT('h4)
	) name25991 (
		_w30021_,
		_w30037_,
		_w30038_
	);
	LUT2 #(
		.INIT('h1)
	) name25992 (
		_w28543_,
		_w30038_,
		_w30039_
	);
	LUT2 #(
		.INIT('h2)
	) name25993 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[12]/P0001 ,
		_w28545_,
		_w30040_
	);
	LUT2 #(
		.INIT('h1)
	) name25994 (
		_w28719_,
		_w30040_,
		_w30041_
	);
	LUT2 #(
		.INIT('h4)
	) name25995 (
		_w30039_,
		_w30041_,
		_w30042_
	);
	LUT2 #(
		.INIT('h8)
	) name25996 (
		_w18191_,
		_w18905_,
		_w30043_
	);
	LUT2 #(
		.INIT('h2)
	) name25997 (
		_w18766_,
		_w18914_,
		_w30044_
	);
	LUT2 #(
		.INIT('h4)
	) name25998 (
		_w18912_,
		_w19862_,
		_w30045_
	);
	LUT2 #(
		.INIT('h2)
	) name25999 (
		_w18759_,
		_w18907_,
		_w30046_
	);
	LUT2 #(
		.INIT('h8)
	) name26000 (
		_w18139_,
		_w18745_,
		_w30047_
	);
	LUT2 #(
		.INIT('h8)
	) name26001 (
		_w18071_,
		_w18124_,
		_w30048_
	);
	LUT2 #(
		.INIT('h8)
	) name26002 (
		_w18187_,
		_w18893_,
		_w30049_
	);
	LUT2 #(
		.INIT('h8)
	) name26003 (
		_w18070_,
		_w18740_,
		_w30050_
	);
	LUT2 #(
		.INIT('h8)
	) name26004 (
		_w18043_,
		_w18751_,
		_w30051_
	);
	LUT2 #(
		.INIT('h4)
	) name26005 (
		_w17924_,
		_w19808_,
		_w30052_
	);
	LUT2 #(
		.INIT('h2)
	) name26006 (
		_w18099_,
		_w18720_,
		_w30053_
	);
	LUT2 #(
		.INIT('h2)
	) name26007 (
		_w18055_,
		_w20096_,
		_w30054_
	);
	LUT2 #(
		.INIT('h4)
	) name26008 (
		_w17998_,
		_w18088_,
		_w30055_
	);
	LUT2 #(
		.INIT('h2)
	) name26009 (
		_w18162_,
		_w18781_,
		_w30056_
	);
	LUT2 #(
		.INIT('h8)
	) name26010 (
		_w17986_,
		_w18752_,
		_w30057_
	);
	LUT2 #(
		.INIT('h2)
	) name26011 (
		_w18039_,
		_w19870_,
		_w30058_
	);
	LUT2 #(
		.INIT('h2)
	) name26012 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9120_,
		_w30059_
	);
	LUT2 #(
		.INIT('h8)
	) name26013 (
		_w18191_,
		_w18749_,
		_w30060_
	);
	LUT2 #(
		.INIT('h4)
	) name26014 (
		_w18170_,
		_w20996_,
		_w30061_
	);
	LUT2 #(
		.INIT('h4)
	) name26015 (
		_w18182_,
		_w20104_,
		_w30062_
	);
	LUT2 #(
		.INIT('h8)
	) name26016 (
		_w18056_,
		_w18756_,
		_w30063_
	);
	LUT2 #(
		.INIT('h8)
	) name26017 (
		_w18153_,
		_w18741_,
		_w30064_
	);
	LUT2 #(
		.INIT('h1)
	) name26018 (
		_w30043_,
		_w30059_,
		_w30065_
	);
	LUT2 #(
		.INIT('h1)
	) name26019 (
		_w30054_,
		_w30057_,
		_w30066_
	);
	LUT2 #(
		.INIT('h1)
	) name26020 (
		_w30060_,
		_w30063_,
		_w30067_
	);
	LUT2 #(
		.INIT('h4)
	) name26021 (
		_w30064_,
		_w30067_,
		_w30068_
	);
	LUT2 #(
		.INIT('h8)
	) name26022 (
		_w30065_,
		_w30066_,
		_w30069_
	);
	LUT2 #(
		.INIT('h1)
	) name26023 (
		_w17969_,
		_w30058_,
		_w30070_
	);
	LUT2 #(
		.INIT('h8)
	) name26024 (
		_w30069_,
		_w30070_,
		_w30071_
	);
	LUT2 #(
		.INIT('h8)
	) name26025 (
		_w19812_,
		_w30068_,
		_w30072_
	);
	LUT2 #(
		.INIT('h1)
	) name26026 (
		_w30044_,
		_w30045_,
		_w30073_
	);
	LUT2 #(
		.INIT('h1)
	) name26027 (
		_w30046_,
		_w30047_,
		_w30074_
	);
	LUT2 #(
		.INIT('h1)
	) name26028 (
		_w30048_,
		_w30049_,
		_w30075_
	);
	LUT2 #(
		.INIT('h1)
	) name26029 (
		_w30050_,
		_w30051_,
		_w30076_
	);
	LUT2 #(
		.INIT('h8)
	) name26030 (
		_w30075_,
		_w30076_,
		_w30077_
	);
	LUT2 #(
		.INIT('h8)
	) name26031 (
		_w30073_,
		_w30074_,
		_w30078_
	);
	LUT2 #(
		.INIT('h8)
	) name26032 (
		_w30071_,
		_w30072_,
		_w30079_
	);
	LUT2 #(
		.INIT('h1)
	) name26033 (
		_w30052_,
		_w30053_,
		_w30080_
	);
	LUT2 #(
		.INIT('h1)
	) name26034 (
		_w30055_,
		_w30056_,
		_w30081_
	);
	LUT2 #(
		.INIT('h1)
	) name26035 (
		_w30061_,
		_w30062_,
		_w30082_
	);
	LUT2 #(
		.INIT('h8)
	) name26036 (
		_w30081_,
		_w30082_,
		_w30083_
	);
	LUT2 #(
		.INIT('h8)
	) name26037 (
		_w30079_,
		_w30080_,
		_w30084_
	);
	LUT2 #(
		.INIT('h8)
	) name26038 (
		_w30077_,
		_w30078_,
		_w30085_
	);
	LUT2 #(
		.INIT('h8)
	) name26039 (
		_w30084_,
		_w30085_,
		_w30086_
	);
	LUT2 #(
		.INIT('h8)
	) name26040 (
		_w30083_,
		_w30086_,
		_w30087_
	);
	LUT2 #(
		.INIT('h8)
	) name26041 (
		_w19791_,
		_w30087_,
		_w30088_
	);
	LUT2 #(
		.INIT('h8)
	) name26042 (
		_w29748_,
		_w30088_,
		_w30089_
	);
	LUT2 #(
		.INIT('h2)
	) name26043 (
		_w28636_,
		_w30089_,
		_w30090_
	);
	LUT2 #(
		.INIT('h8)
	) name26044 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w23920_,
		_w30091_
	);
	LUT2 #(
		.INIT('h4)
	) name26045 (
		_w14413_,
		_w28561_,
		_w30092_
	);
	LUT2 #(
		.INIT('h1)
	) name26046 (
		_w28564_,
		_w30091_,
		_w30093_
	);
	LUT2 #(
		.INIT('h4)
	) name26047 (
		_w30092_,
		_w30093_,
		_w30094_
	);
	LUT2 #(
		.INIT('h2)
	) name26048 (
		_w28559_,
		_w30094_,
		_w30095_
	);
	LUT2 #(
		.INIT('h1)
	) name26049 (
		_w9072_,
		_w28594_,
		_w30096_
	);
	LUT2 #(
		.INIT('h1)
	) name26050 (
		_w9056_,
		_w28589_,
		_w30097_
	);
	LUT2 #(
		.INIT('h1)
	) name26051 (
		_w30096_,
		_w30097_,
		_w30098_
	);
	LUT2 #(
		.INIT('h8)
	) name26052 (
		_w29562_,
		_w30098_,
		_w30099_
	);
	LUT2 #(
		.INIT('h2)
	) name26053 (
		_w28577_,
		_w30099_,
		_w30100_
	);
	LUT2 #(
		.INIT('h1)
	) name26054 (
		_w29303_,
		_w30100_,
		_w30101_
	);
	LUT2 #(
		.INIT('h1)
	) name26055 (
		_w28569_,
		_w30101_,
		_w30102_
	);
	LUT2 #(
		.INIT('h1)
	) name26056 (
		_w12624_,
		_w28572_,
		_w30103_
	);
	LUT2 #(
		.INIT('h4)
	) name26057 (
		_w9178_,
		_w28572_,
		_w30104_
	);
	LUT2 #(
		.INIT('h2)
	) name26058 (
		_w28997_,
		_w30103_,
		_w30105_
	);
	LUT2 #(
		.INIT('h4)
	) name26059 (
		_w30104_,
		_w30105_,
		_w30106_
	);
	LUT2 #(
		.INIT('h1)
	) name26060 (
		_w9103_,
		_w28634_,
		_w30107_
	);
	LUT2 #(
		.INIT('h8)
	) name26061 (
		_w12624_,
		_w28619_,
		_w30108_
	);
	LUT2 #(
		.INIT('h8)
	) name26062 (
		_w9178_,
		_w28630_,
		_w30109_
	);
	LUT2 #(
		.INIT('h1)
	) name26063 (
		_w9120_,
		_w28624_,
		_w30110_
	);
	LUT2 #(
		.INIT('h1)
	) name26064 (
		_w9128_,
		_w28556_,
		_w30111_
	);
	LUT2 #(
		.INIT('h4)
	) name26065 (
		_w18170_,
		_w19717_,
		_w30112_
	);
	LUT2 #(
		.INIT('h2)
	) name26066 (
		_w17945_,
		_w18152_,
		_w30113_
	);
	LUT2 #(
		.INIT('h1)
	) name26067 (
		_w18133_,
		_w18915_,
		_w30114_
	);
	LUT2 #(
		.INIT('h1)
	) name26068 (
		_w18180_,
		_w18919_,
		_w30115_
	);
	LUT2 #(
		.INIT('h1)
	) name26069 (
		_w17938_,
		_w18149_,
		_w30116_
	);
	LUT2 #(
		.INIT('h1)
	) name26070 (
		_w17922_,
		_w19870_,
		_w30117_
	);
	LUT2 #(
		.INIT('h4)
	) name26071 (
		_w18096_,
		_w18752_,
		_w30118_
	);
	LUT2 #(
		.INIT('h4)
	) name26072 (
		_w18108_,
		_w19862_,
		_w30119_
	);
	LUT2 #(
		.INIT('h1)
	) name26073 (
		_w18159_,
		_w20096_,
		_w30120_
	);
	LUT2 #(
		.INIT('h2)
	) name26074 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w9128_,
		_w30121_
	);
	LUT2 #(
		.INIT('h4)
	) name26075 (
		_w18091_,
		_w18766_,
		_w30122_
	);
	LUT2 #(
		.INIT('h1)
	) name26076 (
		_w18121_,
		_w18743_,
		_w30123_
	);
	LUT2 #(
		.INIT('h4)
	) name26077 (
		_w17924_,
		_w18176_,
		_w30124_
	);
	LUT2 #(
		.INIT('h1)
	) name26078 (
		_w30114_,
		_w30121_,
		_w30125_
	);
	LUT2 #(
		.INIT('h1)
	) name26079 (
		_w30115_,
		_w30117_,
		_w30126_
	);
	LUT2 #(
		.INIT('h1)
	) name26080 (
		_w30118_,
		_w30119_,
		_w30127_
	);
	LUT2 #(
		.INIT('h1)
	) name26081 (
		_w30120_,
		_w30122_,
		_w30128_
	);
	LUT2 #(
		.INIT('h4)
	) name26082 (
		_w30123_,
		_w30128_,
		_w30129_
	);
	LUT2 #(
		.INIT('h8)
	) name26083 (
		_w30126_,
		_w30127_,
		_w30130_
	);
	LUT2 #(
		.INIT('h4)
	) name26084 (
		_w30112_,
		_w30125_,
		_w30131_
	);
	LUT2 #(
		.INIT('h1)
	) name26085 (
		_w30113_,
		_w30116_,
		_w30132_
	);
	LUT2 #(
		.INIT('h4)
	) name26086 (
		_w30124_,
		_w30132_,
		_w30133_
	);
	LUT2 #(
		.INIT('h8)
	) name26087 (
		_w30130_,
		_w30131_,
		_w30134_
	);
	LUT2 #(
		.INIT('h4)
	) name26088 (
		_w18085_,
		_w30129_,
		_w30135_
	);
	LUT2 #(
		.INIT('h8)
	) name26089 (
		_w29579_,
		_w30135_,
		_w30136_
	);
	LUT2 #(
		.INIT('h8)
	) name26090 (
		_w30133_,
		_w30134_,
		_w30137_
	);
	LUT2 #(
		.INIT('h8)
	) name26091 (
		_w17988_,
		_w30137_,
		_w30138_
	);
	LUT2 #(
		.INIT('h8)
	) name26092 (
		_w18064_,
		_w30136_,
		_w30139_
	);
	LUT2 #(
		.INIT('h8)
	) name26093 (
		_w29795_,
		_w30139_,
		_w30140_
	);
	LUT2 #(
		.INIT('h8)
	) name26094 (
		_w20159_,
		_w30138_,
		_w30141_
	);
	LUT2 #(
		.INIT('h8)
	) name26095 (
		_w30140_,
		_w30141_,
		_w30142_
	);
	LUT2 #(
		.INIT('h2)
	) name26096 (
		_w28627_,
		_w30142_,
		_w30143_
	);
	LUT2 #(
		.INIT('h1)
	) name26097 (
		_w30107_,
		_w30108_,
		_w30144_
	);
	LUT2 #(
		.INIT('h4)
	) name26098 (
		_w30109_,
		_w30144_,
		_w30145_
	);
	LUT2 #(
		.INIT('h1)
	) name26099 (
		_w30110_,
		_w30111_,
		_w30146_
	);
	LUT2 #(
		.INIT('h8)
	) name26100 (
		_w30145_,
		_w30146_,
		_w30147_
	);
	LUT2 #(
		.INIT('h1)
	) name26101 (
		_w30090_,
		_w30143_,
		_w30148_
	);
	LUT2 #(
		.INIT('h8)
	) name26102 (
		_w30147_,
		_w30148_,
		_w30149_
	);
	LUT2 #(
		.INIT('h4)
	) name26103 (
		_w30106_,
		_w30149_,
		_w30150_
	);
	LUT2 #(
		.INIT('h4)
	) name26104 (
		_w29308_,
		_w30150_,
		_w30151_
	);
	LUT2 #(
		.INIT('h4)
	) name26105 (
		_w30102_,
		_w30151_,
		_w30152_
	);
	LUT2 #(
		.INIT('h4)
	) name26106 (
		_w30095_,
		_w30152_,
		_w30153_
	);
	LUT2 #(
		.INIT('h8)
	) name26107 (
		_w28719_,
		_w30153_,
		_w30154_
	);
	LUT2 #(
		.INIT('h1)
	) name26108 (
		_w30042_,
		_w30154_,
		_w30155_
	);
	LUT2 #(
		.INIT('h8)
	) name26109 (
		_w23920_,
		_w28660_,
		_w30156_
	);
	LUT2 #(
		.INIT('h1)
	) name26110 (
		_w30029_,
		_w30156_,
		_w30157_
	);
	LUT2 #(
		.INIT('h1)
	) name26111 (
		_w28649_,
		_w30157_,
		_w30158_
	);
	LUT2 #(
		.INIT('h8)
	) name26112 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[12]/P0001 ,
		_w28649_,
		_w30159_
	);
	LUT2 #(
		.INIT('h1)
	) name26113 (
		_w30158_,
		_w30159_,
		_w30160_
	);
	LUT2 #(
		.INIT('h1)
	) name26114 (
		_w28550_,
		_w30160_,
		_w30161_
	);
	LUT2 #(
		.INIT('h2)
	) name26115 (
		_w28550_,
		_w30153_,
		_w30162_
	);
	LUT2 #(
		.INIT('h1)
	) name26116 (
		_w30161_,
		_w30162_,
		_w30163_
	);
	LUT2 #(
		.INIT('h8)
	) name26117 (
		_w13006_,
		_w28729_,
		_w30164_
	);
	LUT2 #(
		.INIT('h8)
	) name26118 (
		_w11265_,
		_w28725_,
		_w30165_
	);
	LUT2 #(
		.INIT('h8)
	) name26119 (
		_w11176_,
		_w28705_,
		_w30166_
	);
	LUT2 #(
		.INIT('h2)
	) name26120 (
		_w11180_,
		_w28705_,
		_w30167_
	);
	LUT2 #(
		.INIT('h1)
	) name26121 (
		_w30166_,
		_w30167_,
		_w30168_
	);
	LUT2 #(
		.INIT('h8)
	) name26122 (
		_w28735_,
		_w30168_,
		_w30169_
	);
	LUT2 #(
		.INIT('h8)
	) name26123 (
		_w11184_,
		_w28652_,
		_w30170_
	);
	LUT2 #(
		.INIT('h2)
	) name26124 (
		_w11188_,
		_w28652_,
		_w30171_
	);
	LUT2 #(
		.INIT('h1)
	) name26125 (
		_w28660_,
		_w30170_,
		_w30172_
	);
	LUT2 #(
		.INIT('h4)
	) name26126 (
		_w30171_,
		_w30172_,
		_w30173_
	);
	LUT2 #(
		.INIT('h8)
	) name26127 (
		_w28739_,
		_w30173_,
		_w30174_
	);
	LUT2 #(
		.INIT('h1)
	) name26128 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[7]/P0001 ,
		_w30175_
	);
	LUT2 #(
		.INIT('h2)
	) name26129 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[7]/P0001 ,
		_w30176_
	);
	LUT2 #(
		.INIT('h1)
	) name26130 (
		_w30175_,
		_w30176_,
		_w30177_
	);
	LUT2 #(
		.INIT('h8)
	) name26131 (
		_w28741_,
		_w30177_,
		_w30178_
	);
	LUT2 #(
		.INIT('h1)
	) name26132 (
		_w30169_,
		_w30174_,
		_w30179_
	);
	LUT2 #(
		.INIT('h4)
	) name26133 (
		_w30178_,
		_w30179_,
		_w30180_
	);
	LUT2 #(
		.INIT('h4)
	) name26134 (
		_w30164_,
		_w30180_,
		_w30181_
	);
	LUT2 #(
		.INIT('h4)
	) name26135 (
		_w30165_,
		_w30181_,
		_w30182_
	);
	LUT2 #(
		.INIT('h1)
	) name26136 (
		_w28543_,
		_w30182_,
		_w30183_
	);
	LUT2 #(
		.INIT('h2)
	) name26137 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[7]/P0001 ,
		_w28545_,
		_w30184_
	);
	LUT2 #(
		.INIT('h1)
	) name26138 (
		_w28719_,
		_w30184_,
		_w30185_
	);
	LUT2 #(
		.INIT('h4)
	) name26139 (
		_w30183_,
		_w30185_,
		_w30186_
	);
	LUT2 #(
		.INIT('h4)
	) name26140 (
		_w20030_,
		_w28627_,
		_w30187_
	);
	LUT2 #(
		.INIT('h8)
	) name26141 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w19972_,
		_w30188_
	);
	LUT2 #(
		.INIT('h4)
	) name26142 (
		_w23253_,
		_w28561_,
		_w30189_
	);
	LUT2 #(
		.INIT('h1)
	) name26143 (
		_w28564_,
		_w30188_,
		_w30190_
	);
	LUT2 #(
		.INIT('h4)
	) name26144 (
		_w30189_,
		_w30190_,
		_w30191_
	);
	LUT2 #(
		.INIT('h2)
	) name26145 (
		_w28559_,
		_w30191_,
		_w30192_
	);
	LUT2 #(
		.INIT('h1)
	) name26146 (
		_w11192_,
		_w28594_,
		_w30193_
	);
	LUT2 #(
		.INIT('h1)
	) name26147 (
		_w11196_,
		_w28589_,
		_w30194_
	);
	LUT2 #(
		.INIT('h1)
	) name26148 (
		_w30193_,
		_w30194_,
		_w30195_
	);
	LUT2 #(
		.INIT('h8)
	) name26149 (
		_w29562_,
		_w30195_,
		_w30196_
	);
	LUT2 #(
		.INIT('h2)
	) name26150 (
		_w28577_,
		_w30196_,
		_w30197_
	);
	LUT2 #(
		.INIT('h1)
	) name26151 (
		_w29303_,
		_w30197_,
		_w30198_
	);
	LUT2 #(
		.INIT('h1)
	) name26152 (
		_w28569_,
		_w30198_,
		_w30199_
	);
	LUT2 #(
		.INIT('h4)
	) name26153 (
		_w11265_,
		_w28572_,
		_w30200_
	);
	LUT2 #(
		.INIT('h1)
	) name26154 (
		_w13006_,
		_w28572_,
		_w30201_
	);
	LUT2 #(
		.INIT('h2)
	) name26155 (
		_w28997_,
		_w30200_,
		_w30202_
	);
	LUT2 #(
		.INIT('h4)
	) name26156 (
		_w30201_,
		_w30202_,
		_w30203_
	);
	LUT2 #(
		.INIT('h1)
	) name26157 (
		_w11231_,
		_w28624_,
		_w30204_
	);
	LUT2 #(
		.INIT('h8)
	) name26158 (
		_w11265_,
		_w28630_,
		_w30205_
	);
	LUT2 #(
		.INIT('h2)
	) name26159 (
		_w18111_,
		_w18898_,
		_w30206_
	);
	LUT2 #(
		.INIT('h4)
	) name26160 (
		_w18165_,
		_w20996_,
		_w30207_
	);
	LUT2 #(
		.INIT('h1)
	) name26161 (
		_w18914_,
		_w18991_,
		_w30208_
	);
	LUT2 #(
		.INIT('h1)
	) name26162 (
		_w17935_,
		_w18079_,
		_w30209_
	);
	LUT2 #(
		.INIT('h8)
	) name26163 (
		_w18039_,
		_w18188_,
		_w30210_
	);
	LUT2 #(
		.INIT('h4)
	) name26164 (
		_w18175_,
		_w18922_,
		_w30211_
	);
	LUT2 #(
		.INIT('h2)
	) name26165 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w11231_,
		_w30212_
	);
	LUT2 #(
		.INIT('h8)
	) name26166 (
		_w18124_,
		_w19801_,
		_w30213_
	);
	LUT2 #(
		.INIT('h8)
	) name26167 (
		_w18001_,
		_w18125_,
		_w30214_
	);
	LUT2 #(
		.INIT('h8)
	) name26168 (
		_w18188_,
		_w18191_,
		_w30215_
	);
	LUT2 #(
		.INIT('h2)
	) name26169 (
		_w18099_,
		_w18895_,
		_w30216_
	);
	LUT2 #(
		.INIT('h4)
	) name26170 (
		_w17998_,
		_w18115_,
		_w30217_
	);
	LUT2 #(
		.INIT('h8)
	) name26171 (
		_w18056_,
		_w18103_,
		_w30218_
	);
	LUT2 #(
		.INIT('h2)
	) name26172 (
		_w18128_,
		_w18907_,
		_w30219_
	);
	LUT2 #(
		.INIT('h2)
	) name26173 (
		_w18163_,
		_w18912_,
		_w30220_
	);
	LUT2 #(
		.INIT('h2)
	) name26174 (
		_w18184_,
		_w18918_,
		_w30221_
	);
	LUT2 #(
		.INIT('h8)
	) name26175 (
		_w17980_,
		_w18751_,
		_w30222_
	);
	LUT2 #(
		.INIT('h4)
	) name26176 (
		_w18909_,
		_w19720_,
		_w30223_
	);
	LUT2 #(
		.INIT('h1)
	) name26177 (
		_w30212_,
		_w30214_,
		_w30224_
	);
	LUT2 #(
		.INIT('h1)
	) name26178 (
		_w30215_,
		_w30218_,
		_w30225_
	);
	LUT2 #(
		.INIT('h8)
	) name26179 (
		_w30224_,
		_w30225_,
		_w30226_
	);
	LUT2 #(
		.INIT('h1)
	) name26180 (
		_w18018_,
		_w30210_,
		_w30227_
	);
	LUT2 #(
		.INIT('h8)
	) name26181 (
		_w30226_,
		_w30227_,
		_w30228_
	);
	LUT2 #(
		.INIT('h8)
	) name26182 (
		_w18902_,
		_w19812_,
		_w30229_
	);
	LUT2 #(
		.INIT('h1)
	) name26183 (
		_w30208_,
		_w30209_,
		_w30230_
	);
	LUT2 #(
		.INIT('h1)
	) name26184 (
		_w30213_,
		_w30219_,
		_w30231_
	);
	LUT2 #(
		.INIT('h1)
	) name26185 (
		_w30220_,
		_w30221_,
		_w30232_
	);
	LUT2 #(
		.INIT('h1)
	) name26186 (
		_w30222_,
		_w30223_,
		_w30233_
	);
	LUT2 #(
		.INIT('h8)
	) name26187 (
		_w30232_,
		_w30233_,
		_w30234_
	);
	LUT2 #(
		.INIT('h8)
	) name26188 (
		_w30230_,
		_w30231_,
		_w30235_
	);
	LUT2 #(
		.INIT('h8)
	) name26189 (
		_w30228_,
		_w30229_,
		_w30236_
	);
	LUT2 #(
		.INIT('h1)
	) name26190 (
		_w30206_,
		_w30207_,
		_w30237_
	);
	LUT2 #(
		.INIT('h1)
	) name26191 (
		_w30211_,
		_w30216_,
		_w30238_
	);
	LUT2 #(
		.INIT('h4)
	) name26192 (
		_w30217_,
		_w30238_,
		_w30239_
	);
	LUT2 #(
		.INIT('h8)
	) name26193 (
		_w30236_,
		_w30237_,
		_w30240_
	);
	LUT2 #(
		.INIT('h8)
	) name26194 (
		_w30234_,
		_w30235_,
		_w30241_
	);
	LUT2 #(
		.INIT('h8)
	) name26195 (
		_w30240_,
		_w30241_,
		_w30242_
	);
	LUT2 #(
		.INIT('h8)
	) name26196 (
		_w18790_,
		_w30239_,
		_w30243_
	);
	LUT2 #(
		.INIT('h8)
	) name26197 (
		_w18892_,
		_w30243_,
		_w30244_
	);
	LUT2 #(
		.INIT('h8)
	) name26198 (
		_w30242_,
		_w30244_,
		_w30245_
	);
	LUT2 #(
		.INIT('h2)
	) name26199 (
		_w28636_,
		_w30245_,
		_w30246_
	);
	LUT2 #(
		.INIT('h8)
	) name26200 (
		_w13006_,
		_w28619_,
		_w30247_
	);
	LUT2 #(
		.INIT('h1)
	) name26201 (
		_w11062_,
		_w28634_,
		_w30248_
	);
	LUT2 #(
		.INIT('h1)
	) name26202 (
		_w11239_,
		_w28556_,
		_w30249_
	);
	LUT2 #(
		.INIT('h1)
	) name26203 (
		_w30205_,
		_w30247_,
		_w30250_
	);
	LUT2 #(
		.INIT('h4)
	) name26204 (
		_w30248_,
		_w30250_,
		_w30251_
	);
	LUT2 #(
		.INIT('h1)
	) name26205 (
		_w30204_,
		_w30246_,
		_w30252_
	);
	LUT2 #(
		.INIT('h4)
	) name26206 (
		_w30249_,
		_w30252_,
		_w30253_
	);
	LUT2 #(
		.INIT('h4)
	) name26207 (
		_w30187_,
		_w30251_,
		_w30254_
	);
	LUT2 #(
		.INIT('h8)
	) name26208 (
		_w30253_,
		_w30254_,
		_w30255_
	);
	LUT2 #(
		.INIT('h4)
	) name26209 (
		_w30203_,
		_w30255_,
		_w30256_
	);
	LUT2 #(
		.INIT('h4)
	) name26210 (
		_w29308_,
		_w30256_,
		_w30257_
	);
	LUT2 #(
		.INIT('h4)
	) name26211 (
		_w30199_,
		_w30257_,
		_w30258_
	);
	LUT2 #(
		.INIT('h4)
	) name26212 (
		_w30192_,
		_w30258_,
		_w30259_
	);
	LUT2 #(
		.INIT('h8)
	) name26213 (
		_w28719_,
		_w30259_,
		_w30260_
	);
	LUT2 #(
		.INIT('h1)
	) name26214 (
		_w30186_,
		_w30260_,
		_w30261_
	);
	LUT2 #(
		.INIT('h8)
	) name26215 (
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w28786_,
		_w30262_
	);
	LUT2 #(
		.INIT('h1)
	) name26216 (
		\sport1_cfg_FSi_cnt_reg[14]/NET0131 ,
		_w28869_,
		_w30263_
	);
	LUT2 #(
		.INIT('h2)
	) name26217 (
		_w28855_,
		_w28870_,
		_w30264_
	);
	LUT2 #(
		.INIT('h4)
	) name26218 (
		_w30263_,
		_w30264_,
		_w30265_
	);
	LUT2 #(
		.INIT('h1)
	) name26219 (
		_w30262_,
		_w30265_,
		_w30266_
	);
	LUT2 #(
		.INIT('h8)
	) name26220 (
		_w12715_,
		_w28729_,
		_w30267_
	);
	LUT2 #(
		.INIT('h8)
	) name26221 (
		_w12688_,
		_w28725_,
		_w30268_
	);
	LUT2 #(
		.INIT('h8)
	) name26222 (
		_w11862_,
		_w28705_,
		_w30269_
	);
	LUT2 #(
		.INIT('h2)
	) name26223 (
		_w11866_,
		_w28705_,
		_w30270_
	);
	LUT2 #(
		.INIT('h1)
	) name26224 (
		_w30269_,
		_w30270_,
		_w30271_
	);
	LUT2 #(
		.INIT('h8)
	) name26225 (
		_w28735_,
		_w30271_,
		_w30272_
	);
	LUT2 #(
		.INIT('h8)
	) name26226 (
		_w11870_,
		_w28652_,
		_w30273_
	);
	LUT2 #(
		.INIT('h2)
	) name26227 (
		_w11874_,
		_w28652_,
		_w30274_
	);
	LUT2 #(
		.INIT('h1)
	) name26228 (
		_w28660_,
		_w30273_,
		_w30275_
	);
	LUT2 #(
		.INIT('h4)
	) name26229 (
		_w30274_,
		_w30275_,
		_w30276_
	);
	LUT2 #(
		.INIT('h8)
	) name26230 (
		_w28739_,
		_w30276_,
		_w30277_
	);
	LUT2 #(
		.INIT('h1)
	) name26231 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[14]/P0001 ,
		_w30278_
	);
	LUT2 #(
		.INIT('h2)
	) name26232 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[14]/P0001 ,
		_w30279_
	);
	LUT2 #(
		.INIT('h1)
	) name26233 (
		_w30278_,
		_w30279_,
		_w30280_
	);
	LUT2 #(
		.INIT('h8)
	) name26234 (
		_w28741_,
		_w30280_,
		_w30281_
	);
	LUT2 #(
		.INIT('h1)
	) name26235 (
		_w30272_,
		_w30277_,
		_w30282_
	);
	LUT2 #(
		.INIT('h4)
	) name26236 (
		_w30281_,
		_w30282_,
		_w30283_
	);
	LUT2 #(
		.INIT('h4)
	) name26237 (
		_w30268_,
		_w30283_,
		_w30284_
	);
	LUT2 #(
		.INIT('h4)
	) name26238 (
		_w30267_,
		_w30284_,
		_w30285_
	);
	LUT2 #(
		.INIT('h1)
	) name26239 (
		_w28543_,
		_w30285_,
		_w30286_
	);
	LUT2 #(
		.INIT('h2)
	) name26240 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[14]/P0001 ,
		_w28545_,
		_w30287_
	);
	LUT2 #(
		.INIT('h1)
	) name26241 (
		_w28719_,
		_w30287_,
		_w30288_
	);
	LUT2 #(
		.INIT('h4)
	) name26242 (
		_w30286_,
		_w30288_,
		_w30289_
	);
	LUT2 #(
		.INIT('h4)
	) name26243 (
		_w20192_,
		_w28627_,
		_w30290_
	);
	LUT2 #(
		.INIT('h8)
	) name26244 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w20150_,
		_w30291_
	);
	LUT2 #(
		.INIT('h8)
	) name26245 (
		_w14540_,
		_w28561_,
		_w30292_
	);
	LUT2 #(
		.INIT('h1)
	) name26246 (
		_w28564_,
		_w30291_,
		_w30293_
	);
	LUT2 #(
		.INIT('h4)
	) name26247 (
		_w30292_,
		_w30293_,
		_w30294_
	);
	LUT2 #(
		.INIT('h2)
	) name26248 (
		_w28559_,
		_w30294_,
		_w30295_
	);
	LUT2 #(
		.INIT('h1)
	) name26249 (
		_w11878_,
		_w28594_,
		_w30296_
	);
	LUT2 #(
		.INIT('h1)
	) name26250 (
		_w11882_,
		_w28589_,
		_w30297_
	);
	LUT2 #(
		.INIT('h1)
	) name26251 (
		_w30296_,
		_w30297_,
		_w30298_
	);
	LUT2 #(
		.INIT('h8)
	) name26252 (
		_w29562_,
		_w30298_,
		_w30299_
	);
	LUT2 #(
		.INIT('h2)
	) name26253 (
		_w28577_,
		_w30299_,
		_w30300_
	);
	LUT2 #(
		.INIT('h1)
	) name26254 (
		_w29303_,
		_w30300_,
		_w30301_
	);
	LUT2 #(
		.INIT('h1)
	) name26255 (
		_w28569_,
		_w30301_,
		_w30302_
	);
	LUT2 #(
		.INIT('h1)
	) name26256 (
		_w11837_,
		_w28634_,
		_w30303_
	);
	LUT2 #(
		.INIT('h8)
	) name26257 (
		_w12688_,
		_w28630_,
		_w30304_
	);
	LUT2 #(
		.INIT('h8)
	) name26258 (
		_w12715_,
		_w28619_,
		_w30305_
	);
	LUT2 #(
		.INIT('h1)
	) name26259 (
		_w11854_,
		_w28556_,
		_w30306_
	);
	LUT2 #(
		.INIT('h1)
	) name26260 (
		_w11846_,
		_w28624_,
		_w30307_
	);
	LUT2 #(
		.INIT('h4)
	) name26261 (
		_w21226_,
		_w28636_,
		_w30308_
	);
	LUT2 #(
		.INIT('h1)
	) name26262 (
		_w12715_,
		_w28572_,
		_w30309_
	);
	LUT2 #(
		.INIT('h4)
	) name26263 (
		_w12688_,
		_w28572_,
		_w30310_
	);
	LUT2 #(
		.INIT('h2)
	) name26264 (
		_w28997_,
		_w30309_,
		_w30311_
	);
	LUT2 #(
		.INIT('h4)
	) name26265 (
		_w30310_,
		_w30311_,
		_w30312_
	);
	LUT2 #(
		.INIT('h1)
	) name26266 (
		_w30303_,
		_w30304_,
		_w30313_
	);
	LUT2 #(
		.INIT('h4)
	) name26267 (
		_w30305_,
		_w30313_,
		_w30314_
	);
	LUT2 #(
		.INIT('h1)
	) name26268 (
		_w30306_,
		_w30307_,
		_w30315_
	);
	LUT2 #(
		.INIT('h8)
	) name26269 (
		_w30314_,
		_w30315_,
		_w30316_
	);
	LUT2 #(
		.INIT('h4)
	) name26270 (
		_w30290_,
		_w30316_,
		_w30317_
	);
	LUT2 #(
		.INIT('h4)
	) name26271 (
		_w30308_,
		_w30317_,
		_w30318_
	);
	LUT2 #(
		.INIT('h4)
	) name26272 (
		_w30312_,
		_w30318_,
		_w30319_
	);
	LUT2 #(
		.INIT('h4)
	) name26273 (
		_w29308_,
		_w30319_,
		_w30320_
	);
	LUT2 #(
		.INIT('h4)
	) name26274 (
		_w30302_,
		_w30320_,
		_w30321_
	);
	LUT2 #(
		.INIT('h4)
	) name26275 (
		_w30295_,
		_w30321_,
		_w30322_
	);
	LUT2 #(
		.INIT('h8)
	) name26276 (
		_w28719_,
		_w30322_,
		_w30323_
	);
	LUT2 #(
		.INIT('h1)
	) name26277 (
		_w30289_,
		_w30323_,
		_w30324_
	);
	LUT2 #(
		.INIT('h8)
	) name26278 (
		\sport0_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w28876_,
		_w30325_
	);
	LUT2 #(
		.INIT('h1)
	) name26279 (
		\sport0_cfg_FSi_cnt_reg[14]/NET0131 ,
		_w28959_,
		_w30326_
	);
	LUT2 #(
		.INIT('h2)
	) name26280 (
		_w28945_,
		_w28960_,
		_w30327_
	);
	LUT2 #(
		.INIT('h4)
	) name26281 (
		_w30326_,
		_w30327_,
		_w30328_
	);
	LUT2 #(
		.INIT('h1)
	) name26282 (
		_w30325_,
		_w30328_,
		_w30329_
	);
	LUT2 #(
		.INIT('h8)
	) name26283 (
		_w19972_,
		_w28660_,
		_w30330_
	);
	LUT2 #(
		.INIT('h1)
	) name26284 (
		_w30173_,
		_w30330_,
		_w30331_
	);
	LUT2 #(
		.INIT('h1)
	) name26285 (
		_w28649_,
		_w30331_,
		_w30332_
	);
	LUT2 #(
		.INIT('h8)
	) name26286 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[7]/P0001 ,
		_w28649_,
		_w30333_
	);
	LUT2 #(
		.INIT('h1)
	) name26287 (
		_w30332_,
		_w30333_,
		_w30334_
	);
	LUT2 #(
		.INIT('h1)
	) name26288 (
		_w28550_,
		_w30334_,
		_w30335_
	);
	LUT2 #(
		.INIT('h2)
	) name26289 (
		_w28550_,
		_w30259_,
		_w30336_
	);
	LUT2 #(
		.INIT('h1)
	) name26290 (
		_w30335_,
		_w30336_,
		_w30337_
	);
	LUT2 #(
		.INIT('h8)
	) name26291 (
		_w20150_,
		_w28660_,
		_w30338_
	);
	LUT2 #(
		.INIT('h1)
	) name26292 (
		_w30276_,
		_w30338_,
		_w30339_
	);
	LUT2 #(
		.INIT('h1)
	) name26293 (
		_w28649_,
		_w30339_,
		_w30340_
	);
	LUT2 #(
		.INIT('h8)
	) name26294 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[14]/P0001 ,
		_w28649_,
		_w30341_
	);
	LUT2 #(
		.INIT('h1)
	) name26295 (
		_w30340_,
		_w30341_,
		_w30342_
	);
	LUT2 #(
		.INIT('h1)
	) name26296 (
		_w28550_,
		_w30342_,
		_w30343_
	);
	LUT2 #(
		.INIT('h2)
	) name26297 (
		_w28550_,
		_w30322_,
		_w30344_
	);
	LUT2 #(
		.INIT('h1)
	) name26298 (
		_w30343_,
		_w30344_,
		_w30345_
	);
	LUT2 #(
		.INIT('h4)
	) name26299 (
		_w18161_,
		_w19717_,
		_w30346_
	);
	LUT2 #(
		.INIT('h4)
	) name26300 (
		_w18170_,
		_w18732_,
		_w30347_
	);
	LUT2 #(
		.INIT('h8)
	) name26301 (
		_w18748_,
		_w18761_,
		_w30348_
	);
	LUT2 #(
		.INIT('h8)
	) name26302 (
		_w18089_,
		_w19863_,
		_w30349_
	);
	LUT2 #(
		.INIT('h2)
	) name26303 (
		_w17925_,
		_w29063_,
		_w30350_
	);
	LUT2 #(
		.INIT('h2)
	) name26304 (
		_w18088_,
		_w18775_,
		_w30351_
	);
	LUT2 #(
		.INIT('h4)
	) name26305 (
		_w17924_,
		_w18719_,
		_w30352_
	);
	LUT2 #(
		.INIT('h1)
	) name26306 (
		_w18180_,
		_w18743_,
		_w30353_
	);
	LUT2 #(
		.INIT('h4)
	) name26307 (
		_w18159_,
		_w18752_,
		_w30354_
	);
	LUT2 #(
		.INIT('h4)
	) name26308 (
		_w18091_,
		_w19862_,
		_w30355_
	);
	LUT2 #(
		.INIT('h4)
	) name26309 (
		_w18108_,
		_w18756_,
		_w30356_
	);
	LUT2 #(
		.INIT('h8)
	) name26310 (
		_w17986_,
		_w18905_,
		_w30357_
	);
	LUT2 #(
		.INIT('h2)
	) name26311 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w10575_,
		_w30358_
	);
	LUT2 #(
		.INIT('h1)
	) name26312 (
		_w18133_,
		_w20096_,
		_w30359_
	);
	LUT2 #(
		.INIT('h8)
	) name26313 (
		_w18043_,
		_w18748_,
		_w30360_
	);
	LUT2 #(
		.INIT('h8)
	) name26314 (
		_w18070_,
		_w18765_,
		_w30361_
	);
	LUT2 #(
		.INIT('h4)
	) name26315 (
		_w18110_,
		_w18147_,
		_w30362_
	);
	LUT2 #(
		.INIT('h1)
	) name26316 (
		_w17922_,
		_w18915_,
		_w30363_
	);
	LUT2 #(
		.INIT('h8)
	) name26317 (
		_w18153_,
		_w18766_,
		_w30364_
	);
	LUT2 #(
		.INIT('h1)
	) name26318 (
		_w30349_,
		_w30358_,
		_w30365_
	);
	LUT2 #(
		.INIT('h1)
	) name26319 (
		_w30357_,
		_w30364_,
		_w30366_
	);
	LUT2 #(
		.INIT('h8)
	) name26320 (
		_w30365_,
		_w30366_,
		_w30367_
	);
	LUT2 #(
		.INIT('h1)
	) name26321 (
		_w18058_,
		_w30348_,
		_w30368_
	);
	LUT2 #(
		.INIT('h4)
	) name26322 (
		_w30352_,
		_w30368_,
		_w30369_
	);
	LUT2 #(
		.INIT('h4)
	) name26323 (
		_w18069_,
		_w30367_,
		_w30370_
	);
	LUT2 #(
		.INIT('h1)
	) name26324 (
		_w18140_,
		_w30347_,
		_w30371_
	);
	LUT2 #(
		.INIT('h1)
	) name26325 (
		_w30353_,
		_w30354_,
		_w30372_
	);
	LUT2 #(
		.INIT('h1)
	) name26326 (
		_w30355_,
		_w30356_,
		_w30373_
	);
	LUT2 #(
		.INIT('h1)
	) name26327 (
		_w30359_,
		_w30360_,
		_w30374_
	);
	LUT2 #(
		.INIT('h1)
	) name26328 (
		_w30361_,
		_w30362_,
		_w30375_
	);
	LUT2 #(
		.INIT('h4)
	) name26329 (
		_w30363_,
		_w30375_,
		_w30376_
	);
	LUT2 #(
		.INIT('h8)
	) name26330 (
		_w30373_,
		_w30374_,
		_w30377_
	);
	LUT2 #(
		.INIT('h8)
	) name26331 (
		_w30371_,
		_w30372_,
		_w30378_
	);
	LUT2 #(
		.INIT('h8)
	) name26332 (
		_w30369_,
		_w30370_,
		_w30379_
	);
	LUT2 #(
		.INIT('h2)
	) name26333 (
		_w18041_,
		_w19991_,
		_w30380_
	);
	LUT2 #(
		.INIT('h2)
	) name26334 (
		_w29052_,
		_w30346_,
		_w30381_
	);
	LUT2 #(
		.INIT('h1)
	) name26335 (
		_w30350_,
		_w30351_,
		_w30382_
	);
	LUT2 #(
		.INIT('h8)
	) name26336 (
		_w30381_,
		_w30382_,
		_w30383_
	);
	LUT2 #(
		.INIT('h8)
	) name26337 (
		_w30379_,
		_w30380_,
		_w30384_
	);
	LUT2 #(
		.INIT('h8)
	) name26338 (
		_w30377_,
		_w30378_,
		_w30385_
	);
	LUT2 #(
		.INIT('h4)
	) name26339 (
		_w18085_,
		_w30376_,
		_w30386_
	);
	LUT2 #(
		.INIT('h8)
	) name26340 (
		_w30385_,
		_w30386_,
		_w30387_
	);
	LUT2 #(
		.INIT('h8)
	) name26341 (
		_w30383_,
		_w30384_,
		_w30388_
	);
	LUT2 #(
		.INIT('h8)
	) name26342 (
		_w18726_,
		_w30388_,
		_w30389_
	);
	LUT2 #(
		.INIT('h8)
	) name26343 (
		_w30387_,
		_w30389_,
		_w30390_
	);
	LUT2 #(
		.INIT('h8)
	) name26344 (
		_w19977_,
		_w30390_,
		_w30391_
	);
	LUT2 #(
		.INIT('h8)
	) name26345 (
		_w29047_,
		_w30391_,
		_w30392_
	);
	LUT2 #(
		.INIT('h2)
	) name26346 (
		_w28627_,
		_w30392_,
		_w30393_
	);
	LUT2 #(
		.INIT('h8)
	) name26347 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w23860_,
		_w30394_
	);
	LUT2 #(
		.INIT('h4)
	) name26348 (
		_w14658_,
		_w28561_,
		_w30395_
	);
	LUT2 #(
		.INIT('h1)
	) name26349 (
		_w28564_,
		_w30394_,
		_w30396_
	);
	LUT2 #(
		.INIT('h4)
	) name26350 (
		_w30395_,
		_w30396_,
		_w30397_
	);
	LUT2 #(
		.INIT('h2)
	) name26351 (
		_w28559_,
		_w30397_,
		_w30398_
	);
	LUT2 #(
		.INIT('h1)
	) name26352 (
		_w10534_,
		_w28594_,
		_w30399_
	);
	LUT2 #(
		.INIT('h1)
	) name26353 (
		_w10538_,
		_w28589_,
		_w30400_
	);
	LUT2 #(
		.INIT('h1)
	) name26354 (
		_w30399_,
		_w30400_,
		_w30401_
	);
	LUT2 #(
		.INIT('h8)
	) name26355 (
		_w29562_,
		_w30401_,
		_w30402_
	);
	LUT2 #(
		.INIT('h2)
	) name26356 (
		_w28577_,
		_w30402_,
		_w30403_
	);
	LUT2 #(
		.INIT('h1)
	) name26357 (
		_w29303_,
		_w30403_,
		_w30404_
	);
	LUT2 #(
		.INIT('h1)
	) name26358 (
		_w28569_,
		_w30404_,
		_w30405_
	);
	LUT2 #(
		.INIT('h1)
	) name26359 (
		_w13041_,
		_w28572_,
		_w30406_
	);
	LUT2 #(
		.INIT('h4)
	) name26360 (
		_w10638_,
		_w28572_,
		_w30407_
	);
	LUT2 #(
		.INIT('h2)
	) name26361 (
		_w28997_,
		_w30406_,
		_w30408_
	);
	LUT2 #(
		.INIT('h4)
	) name26362 (
		_w30407_,
		_w30408_,
		_w30409_
	);
	LUT2 #(
		.INIT('h8)
	) name26363 (
		_w17952_,
		_w18746_,
		_w30410_
	);
	LUT2 #(
		.INIT('h2)
	) name26364 (
		_w18748_,
		_w18898_,
		_w30411_
	);
	LUT2 #(
		.INIT('h2)
	) name26365 (
		_w18740_,
		_w18895_,
		_w30412_
	);
	LUT2 #(
		.INIT('h1)
	) name26366 (
		_w18098_,
		_w18781_,
		_w30413_
	);
	LUT2 #(
		.INIT('h2)
	) name26367 (
		_w18751_,
		_w19818_,
		_w30414_
	);
	LUT2 #(
		.INIT('h4)
	) name26368 (
		_w18170_,
		_w19808_,
		_w30415_
	);
	LUT2 #(
		.INIT('h4)
	) name26369 (
		_w18182_,
		_w19785_,
		_w30416_
	);
	LUT2 #(
		.INIT('h1)
	) name26370 (
		_w18912_,
		_w18919_,
		_w30417_
	);
	LUT2 #(
		.INIT('h4)
	) name26371 (
		_w17938_,
		_w18922_,
		_w30418_
	);
	LUT2 #(
		.INIT('h4)
	) name26372 (
		_w17998_,
		_w18111_,
		_w30419_
	);
	LUT2 #(
		.INIT('h2)
	) name26373 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w10567_,
		_w30420_
	);
	LUT2 #(
		.INIT('h8)
	) name26374 (
		_w18001_,
		_w18745_,
		_w30421_
	);
	LUT2 #(
		.INIT('h1)
	) name26375 (
		_w18037_,
		_w30421_,
		_w30422_
	);
	LUT2 #(
		.INIT('h4)
	) name26376 (
		_w29533_,
		_w30422_,
		_w30423_
	);
	LUT2 #(
		.INIT('h8)
	) name26377 (
		_w29536_,
		_w30423_,
		_w30424_
	);
	LUT2 #(
		.INIT('h1)
	) name26378 (
		_w17931_,
		_w30424_,
		_w30425_
	);
	LUT2 #(
		.INIT('h4)
	) name26379 (
		_w17924_,
		_w18080_,
		_w30426_
	);
	LUT2 #(
		.INIT('h2)
	) name26380 (
		_w18763_,
		_w18907_,
		_w30427_
	);
	LUT2 #(
		.INIT('h1)
	) name26381 (
		_w30410_,
		_w30420_,
		_w30428_
	);
	LUT2 #(
		.INIT('h4)
	) name26382 (
		_w30417_,
		_w30428_,
		_w30429_
	);
	LUT2 #(
		.INIT('h4)
	) name26383 (
		_w30427_,
		_w30429_,
		_w30430_
	);
	LUT2 #(
		.INIT('h1)
	) name26384 (
		_w30411_,
		_w30412_,
		_w30431_
	);
	LUT2 #(
		.INIT('h1)
	) name26385 (
		_w30413_,
		_w30414_,
		_w30432_
	);
	LUT2 #(
		.INIT('h1)
	) name26386 (
		_w30415_,
		_w30416_,
		_w30433_
	);
	LUT2 #(
		.INIT('h1)
	) name26387 (
		_w30418_,
		_w30419_,
		_w30434_
	);
	LUT2 #(
		.INIT('h4)
	) name26388 (
		_w30426_,
		_w30434_,
		_w30435_
	);
	LUT2 #(
		.INIT('h8)
	) name26389 (
		_w30432_,
		_w30433_,
		_w30436_
	);
	LUT2 #(
		.INIT('h8)
	) name26390 (
		_w30430_,
		_w30431_,
		_w30437_
	);
	LUT2 #(
		.INIT('h8)
	) name26391 (
		_w30436_,
		_w30437_,
		_w30438_
	);
	LUT2 #(
		.INIT('h4)
	) name26392 (
		_w30425_,
		_w30435_,
		_w30439_
	);
	LUT2 #(
		.INIT('h8)
	) name26393 (
		_w30438_,
		_w30439_,
		_w30440_
	);
	LUT2 #(
		.INIT('h8)
	) name26394 (
		_w29522_,
		_w30440_,
		_w30441_
	);
	LUT2 #(
		.INIT('h2)
	) name26395 (
		_w28636_,
		_w30441_,
		_w30442_
	);
	LUT2 #(
		.INIT('h8)
	) name26396 (
		_w10638_,
		_w28630_,
		_w30443_
	);
	LUT2 #(
		.INIT('h8)
	) name26397 (
		_w13041_,
		_w28619_,
		_w30444_
	);
	LUT2 #(
		.INIT('h1)
	) name26398 (
		_w10461_,
		_w28634_,
		_w30445_
	);
	LUT2 #(
		.INIT('h1)
	) name26399 (
		_w10575_,
		_w28556_,
		_w30446_
	);
	LUT2 #(
		.INIT('h1)
	) name26400 (
		_w10567_,
		_w28624_,
		_w30447_
	);
	LUT2 #(
		.INIT('h1)
	) name26401 (
		_w30443_,
		_w30444_,
		_w30448_
	);
	LUT2 #(
		.INIT('h4)
	) name26402 (
		_w30445_,
		_w30448_,
		_w30449_
	);
	LUT2 #(
		.INIT('h1)
	) name26403 (
		_w30442_,
		_w30446_,
		_w30450_
	);
	LUT2 #(
		.INIT('h4)
	) name26404 (
		_w30447_,
		_w30450_,
		_w30451_
	);
	LUT2 #(
		.INIT('h8)
	) name26405 (
		_w30449_,
		_w30451_,
		_w30452_
	);
	LUT2 #(
		.INIT('h4)
	) name26406 (
		_w30393_,
		_w30452_,
		_w30453_
	);
	LUT2 #(
		.INIT('h4)
	) name26407 (
		_w30409_,
		_w30453_,
		_w30454_
	);
	LUT2 #(
		.INIT('h4)
	) name26408 (
		_w29308_,
		_w30454_,
		_w30455_
	);
	LUT2 #(
		.INIT('h4)
	) name26409 (
		_w30405_,
		_w30455_,
		_w30456_
	);
	LUT2 #(
		.INIT('h4)
	) name26410 (
		_w30398_,
		_w30456_,
		_w30457_
	);
	LUT2 #(
		.INIT('h2)
	) name26411 (
		_w28719_,
		_w30457_,
		_w30458_
	);
	LUT2 #(
		.INIT('h4)
	) name26412 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		_w28543_,
		_w30459_
	);
	LUT2 #(
		.INIT('h8)
	) name26413 (
		_w13041_,
		_w28729_,
		_w30460_
	);
	LUT2 #(
		.INIT('h8)
	) name26414 (
		_w10638_,
		_w28725_,
		_w30461_
	);
	LUT2 #(
		.INIT('h8)
	) name26415 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[8]/P0001 ,
		_w28544_,
		_w30462_
	);
	LUT2 #(
		.INIT('h8)
	) name26416 (
		_w10526_,
		_w28652_,
		_w30463_
	);
	LUT2 #(
		.INIT('h2)
	) name26417 (
		_w10530_,
		_w28652_,
		_w30464_
	);
	LUT2 #(
		.INIT('h1)
	) name26418 (
		_w28660_,
		_w30463_,
		_w30465_
	);
	LUT2 #(
		.INIT('h4)
	) name26419 (
		_w30464_,
		_w30465_,
		_w30466_
	);
	LUT2 #(
		.INIT('h8)
	) name26420 (
		_w28739_,
		_w30466_,
		_w30467_
	);
	LUT2 #(
		.INIT('h8)
	) name26421 (
		_w10518_,
		_w28705_,
		_w30468_
	);
	LUT2 #(
		.INIT('h2)
	) name26422 (
		_w10522_,
		_w28705_,
		_w30469_
	);
	LUT2 #(
		.INIT('h1)
	) name26423 (
		_w30468_,
		_w30469_,
		_w30470_
	);
	LUT2 #(
		.INIT('h8)
	) name26424 (
		_w28735_,
		_w30470_,
		_w30471_
	);
	LUT2 #(
		.INIT('h1)
	) name26425 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[8]/P0001 ,
		_w30472_
	);
	LUT2 #(
		.INIT('h2)
	) name26426 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[8]/P0001 ,
		_w30473_
	);
	LUT2 #(
		.INIT('h1)
	) name26427 (
		_w30472_,
		_w30473_,
		_w30474_
	);
	LUT2 #(
		.INIT('h8)
	) name26428 (
		_w28741_,
		_w30474_,
		_w30475_
	);
	LUT2 #(
		.INIT('h1)
	) name26429 (
		_w30462_,
		_w30467_,
		_w30476_
	);
	LUT2 #(
		.INIT('h1)
	) name26430 (
		_w30471_,
		_w30475_,
		_w30477_
	);
	LUT2 #(
		.INIT('h8)
	) name26431 (
		_w30476_,
		_w30477_,
		_w30478_
	);
	LUT2 #(
		.INIT('h1)
	) name26432 (
		_w29707_,
		_w30478_,
		_w30479_
	);
	LUT2 #(
		.INIT('h1)
	) name26433 (
		_w28543_,
		_w30460_,
		_w30480_
	);
	LUT2 #(
		.INIT('h4)
	) name26434 (
		_w30479_,
		_w30480_,
		_w30481_
	);
	LUT2 #(
		.INIT('h4)
	) name26435 (
		_w30461_,
		_w30481_,
		_w30482_
	);
	LUT2 #(
		.INIT('h1)
	) name26436 (
		_w28719_,
		_w30459_,
		_w30483_
	);
	LUT2 #(
		.INIT('h4)
	) name26437 (
		_w30482_,
		_w30483_,
		_w30484_
	);
	LUT2 #(
		.INIT('h1)
	) name26438 (
		_w30458_,
		_w30484_,
		_w30485_
	);
	LUT2 #(
		.INIT('h8)
	) name26439 (
		_w23860_,
		_w28660_,
		_w30486_
	);
	LUT2 #(
		.INIT('h1)
	) name26440 (
		_w30466_,
		_w30486_,
		_w30487_
	);
	LUT2 #(
		.INIT('h1)
	) name26441 (
		_w28649_,
		_w30487_,
		_w30488_
	);
	LUT2 #(
		.INIT('h8)
	) name26442 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[8]/P0001 ,
		_w28649_,
		_w30489_
	);
	LUT2 #(
		.INIT('h1)
	) name26443 (
		_w30488_,
		_w30489_,
		_w30490_
	);
	LUT2 #(
		.INIT('h1)
	) name26444 (
		_w28550_,
		_w30490_,
		_w30491_
	);
	LUT2 #(
		.INIT('h2)
	) name26445 (
		_w28550_,
		_w30457_,
		_w30492_
	);
	LUT2 #(
		.INIT('h1)
	) name26446 (
		_w30491_,
		_w30492_,
		_w30493_
	);
	LUT2 #(
		.INIT('h4)
	) name26447 (
		_w14610_,
		_w28561_,
		_w30494_
	);
	LUT2 #(
		.INIT('h8)
	) name26448 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w21663_,
		_w30495_
	);
	LUT2 #(
		.INIT('h1)
	) name26449 (
		_w28564_,
		_w30495_,
		_w30496_
	);
	LUT2 #(
		.INIT('h4)
	) name26450 (
		_w30494_,
		_w30496_,
		_w30497_
	);
	LUT2 #(
		.INIT('h2)
	) name26451 (
		_w28559_,
		_w30497_,
		_w30498_
	);
	LUT2 #(
		.INIT('h4)
	) name26452 (
		_w21958_,
		_w28636_,
		_w30499_
	);
	LUT2 #(
		.INIT('h8)
	) name26453 (
		_w8113_,
		_w28630_,
		_w30500_
	);
	LUT2 #(
		.INIT('h4)
	) name26454 (
		_w21700_,
		_w28627_,
		_w30501_
	);
	LUT2 #(
		.INIT('h1)
	) name26455 (
		_w7987_,
		_w28624_,
		_w30502_
	);
	LUT2 #(
		.INIT('h1)
	) name26456 (
		_w7991_,
		_w28556_,
		_w30503_
	);
	LUT2 #(
		.INIT('h1)
	) name26457 (
		_w12870_,
		_w28577_,
		_w30504_
	);
	LUT2 #(
		.INIT('h4)
	) name26458 (
		_w8113_,
		_w28577_,
		_w30505_
	);
	LUT2 #(
		.INIT('h1)
	) name26459 (
		_w28575_,
		_w30504_,
		_w30506_
	);
	LUT2 #(
		.INIT('h4)
	) name26460 (
		_w30505_,
		_w30506_,
		_w30507_
	);
	LUT2 #(
		.INIT('h1)
	) name26461 (
		_w28576_,
		_w30507_,
		_w30508_
	);
	LUT2 #(
		.INIT('h2)
	) name26462 (
		_w28569_,
		_w30508_,
		_w30509_
	);
	LUT2 #(
		.INIT('h1)
	) name26463 (
		_w7952_,
		_w28634_,
		_w30510_
	);
	LUT2 #(
		.INIT('h8)
	) name26464 (
		_w12870_,
		_w28619_,
		_w30511_
	);
	LUT2 #(
		.INIT('h1)
	) name26465 (
		_w8113_,
		_w28572_,
		_w30512_
	);
	LUT2 #(
		.INIT('h1)
	) name26466 (
		_w7905_,
		_w28598_,
		_w30513_
	);
	LUT2 #(
		.INIT('h1)
	) name26467 (
		_w7909_,
		_w28594_,
		_w30514_
	);
	LUT2 #(
		.INIT('h1)
	) name26468 (
		_w7885_,
		_w28589_,
		_w30515_
	);
	LUT2 #(
		.INIT('h1)
	) name26469 (
		_w30513_,
		_w30514_,
		_w30516_
	);
	LUT2 #(
		.INIT('h4)
	) name26470 (
		_w30515_,
		_w30516_,
		_w30517_
	);
	LUT2 #(
		.INIT('h8)
	) name26471 (
		_w28607_,
		_w30517_,
		_w30518_
	);
	LUT2 #(
		.INIT('h8)
	) name26472 (
		_w28572_,
		_w30518_,
		_w30519_
	);
	LUT2 #(
		.INIT('h2)
	) name26473 (
		_w28584_,
		_w30512_,
		_w30520_
	);
	LUT2 #(
		.INIT('h4)
	) name26474 (
		_w30519_,
		_w30520_,
		_w30521_
	);
	LUT2 #(
		.INIT('h1)
	) name26475 (
		_w30499_,
		_w30500_,
		_w30522_
	);
	LUT2 #(
		.INIT('h1)
	) name26476 (
		_w30510_,
		_w30511_,
		_w30523_
	);
	LUT2 #(
		.INIT('h8)
	) name26477 (
		_w30522_,
		_w30523_,
		_w30524_
	);
	LUT2 #(
		.INIT('h1)
	) name26478 (
		_w30502_,
		_w30503_,
		_w30525_
	);
	LUT2 #(
		.INIT('h8)
	) name26479 (
		_w30524_,
		_w30525_,
		_w30526_
	);
	LUT2 #(
		.INIT('h4)
	) name26480 (
		_w30501_,
		_w30526_,
		_w30527_
	);
	LUT2 #(
		.INIT('h4)
	) name26481 (
		_w30521_,
		_w30527_,
		_w30528_
	);
	LUT2 #(
		.INIT('h4)
	) name26482 (
		_w30509_,
		_w30528_,
		_w30529_
	);
	LUT2 #(
		.INIT('h4)
	) name26483 (
		_w30498_,
		_w30529_,
		_w30530_
	);
	LUT2 #(
		.INIT('h2)
	) name26484 (
		_w28550_,
		_w30530_,
		_w30531_
	);
	LUT2 #(
		.INIT('h4)
	) name26485 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[3]/P0001 ,
		_w28649_,
		_w30532_
	);
	LUT2 #(
		.INIT('h8)
	) name26486 (
		_w7889_,
		_w28652_,
		_w30533_
	);
	LUT2 #(
		.INIT('h2)
	) name26487 (
		_w7901_,
		_w28652_,
		_w30534_
	);
	LUT2 #(
		.INIT('h1)
	) name26488 (
		_w28660_,
		_w30533_,
		_w30535_
	);
	LUT2 #(
		.INIT('h4)
	) name26489 (
		_w30534_,
		_w30535_,
		_w30536_
	);
	LUT2 #(
		.INIT('h8)
	) name26490 (
		_w21663_,
		_w28660_,
		_w30537_
	);
	LUT2 #(
		.INIT('h1)
	) name26491 (
		_w28649_,
		_w30536_,
		_w30538_
	);
	LUT2 #(
		.INIT('h4)
	) name26492 (
		_w30537_,
		_w30538_,
		_w30539_
	);
	LUT2 #(
		.INIT('h1)
	) name26493 (
		_w28550_,
		_w30532_,
		_w30540_
	);
	LUT2 #(
		.INIT('h4)
	) name26494 (
		_w30539_,
		_w30540_,
		_w30541_
	);
	LUT2 #(
		.INIT('h1)
	) name26495 (
		_w30531_,
		_w30541_,
		_w30542_
	);
	LUT2 #(
		.INIT('h8)
	) name26496 (
		_w7607_,
		_w28630_,
		_w30543_
	);
	LUT2 #(
		.INIT('h8)
	) name26497 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w19559_,
		_w30544_
	);
	LUT2 #(
		.INIT('h4)
	) name26498 (
		_w14564_,
		_w28561_,
		_w30545_
	);
	LUT2 #(
		.INIT('h1)
	) name26499 (
		_w28564_,
		_w30544_,
		_w30546_
	);
	LUT2 #(
		.INIT('h4)
	) name26500 (
		_w30545_,
		_w30546_,
		_w30547_
	);
	LUT2 #(
		.INIT('h2)
	) name26501 (
		_w28559_,
		_w30547_,
		_w30548_
	);
	LUT2 #(
		.INIT('h4)
	) name26502 (
		_w7607_,
		_w28577_,
		_w30549_
	);
	LUT2 #(
		.INIT('h1)
	) name26503 (
		_w12520_,
		_w28577_,
		_w30550_
	);
	LUT2 #(
		.INIT('h1)
	) name26504 (
		_w28575_,
		_w30549_,
		_w30551_
	);
	LUT2 #(
		.INIT('h4)
	) name26505 (
		_w30550_,
		_w30551_,
		_w30552_
	);
	LUT2 #(
		.INIT('h1)
	) name26506 (
		_w28576_,
		_w30552_,
		_w30553_
	);
	LUT2 #(
		.INIT('h2)
	) name26507 (
		_w28569_,
		_w30553_,
		_w30554_
	);
	LUT2 #(
		.INIT('h1)
	) name26508 (
		_w7377_,
		_w28556_,
		_w30555_
	);
	LUT2 #(
		.INIT('h1)
	) name26509 (
		_w7381_,
		_w28624_,
		_w30556_
	);
	LUT2 #(
		.INIT('h1)
	) name26510 (
		_w7422_,
		_w28634_,
		_w30557_
	);
	LUT2 #(
		.INIT('h8)
	) name26511 (
		_w18056_,
		_w19862_,
		_w30558_
	);
	LUT2 #(
		.INIT('h8)
	) name26512 (
		_w18071_,
		_w18183_,
		_w30559_
	);
	LUT2 #(
		.INIT('h2)
	) name26513 (
		_w18905_,
		_w18907_,
		_w30560_
	);
	LUT2 #(
		.INIT('h8)
	) name26514 (
		_w18115_,
		_w18893_,
		_w30561_
	);
	LUT2 #(
		.INIT('h8)
	) name26515 (
		_w18070_,
		_w18187_,
		_w30562_
	);
	LUT2 #(
		.INIT('h8)
	) name26516 (
		_w18139_,
		_w18758_,
		_w30563_
	);
	LUT2 #(
		.INIT('h2)
	) name26517 (
		_w18171_,
		_w18781_,
		_w30564_
	);
	LUT2 #(
		.INIT('h4)
	) name26518 (
		_w17924_,
		_w20996_,
		_w30565_
	);
	LUT2 #(
		.INIT('h2)
	) name26519 (
		_w18745_,
		_w19804_,
		_w30566_
	);
	LUT2 #(
		.INIT('h2)
	) name26520 (
		_w18153_,
		_w18919_,
		_w30567_
	);
	LUT2 #(
		.INIT('h1)
	) name26521 (
		_w18091_,
		_w18743_,
		_w30568_
	);
	LUT2 #(
		.INIT('h8)
	) name26522 (
		_w18001_,
		_w18749_,
		_w30569_
	);
	LUT2 #(
		.INIT('h8)
	) name26523 (
		_w18046_,
		_w18162_,
		_w30570_
	);
	LUT2 #(
		.INIT('h8)
	) name26524 (
		_w18124_,
		_w18147_,
		_w30571_
	);
	LUT2 #(
		.INIT('h8)
	) name26525 (
		_w17952_,
		_w18749_,
		_w30572_
	);
	LUT2 #(
		.INIT('h4)
	) name26526 (
		_w18918_,
		_w20308_,
		_w30573_
	);
	LUT2 #(
		.INIT('h8)
	) name26527 (
		_w17915_,
		_w18751_,
		_w30574_
	);
	LUT2 #(
		.INIT('h1)
	) name26528 (
		_w18192_,
		_w30574_,
		_w30575_
	);
	LUT2 #(
		.INIT('h1)
	) name26529 (
		_w17929_,
		_w30575_,
		_w30576_
	);
	LUT2 #(
		.INIT('h2)
	) name26530 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		_w7377_,
		_w30577_
	);
	LUT2 #(
		.INIT('h4)
	) name26531 (
		_w18123_,
		_w18148_,
		_w30578_
	);
	LUT2 #(
		.INIT('h2)
	) name26532 (
		_w18766_,
		_w18912_,
		_w30579_
	);
	LUT2 #(
		.INIT('h8)
	) name26533 (
		_w18055_,
		_w18754_,
		_w30580_
	);
	LUT2 #(
		.INIT('h8)
	) name26534 (
		_w18055_,
		_w18759_,
		_w30581_
	);
	LUT2 #(
		.INIT('h8)
	) name26535 (
		_w17921_,
		_w18752_,
		_w30582_
	);
	LUT2 #(
		.INIT('h1)
	) name26536 (
		_w30558_,
		_w30577_,
		_w30583_
	);
	LUT2 #(
		.INIT('h1)
	) name26537 (
		_w30567_,
		_w30569_,
		_w30584_
	);
	LUT2 #(
		.INIT('h1)
	) name26538 (
		_w30580_,
		_w30581_,
		_w30585_
	);
	LUT2 #(
		.INIT('h4)
	) name26539 (
		_w30582_,
		_w30585_,
		_w30586_
	);
	LUT2 #(
		.INIT('h8)
	) name26540 (
		_w30583_,
		_w30584_,
		_w30587_
	);
	LUT2 #(
		.INIT('h1)
	) name26541 (
		_w18018_,
		_w29242_,
		_w30588_
	);
	LUT2 #(
		.INIT('h1)
	) name26542 (
		_w30572_,
		_w30578_,
		_w30589_
	);
	LUT2 #(
		.INIT('h8)
	) name26543 (
		_w30588_,
		_w30589_,
		_w30590_
	);
	LUT2 #(
		.INIT('h8)
	) name26544 (
		_w30586_,
		_w30587_,
		_w30591_
	);
	LUT2 #(
		.INIT('h2)
	) name26545 (
		_w18038_,
		_w30559_,
		_w30592_
	);
	LUT2 #(
		.INIT('h1)
	) name26546 (
		_w30560_,
		_w30561_,
		_w30593_
	);
	LUT2 #(
		.INIT('h1)
	) name26547 (
		_w30562_,
		_w30563_,
		_w30594_
	);
	LUT2 #(
		.INIT('h1)
	) name26548 (
		_w30568_,
		_w30570_,
		_w30595_
	);
	LUT2 #(
		.INIT('h1)
	) name26549 (
		_w30571_,
		_w30573_,
		_w30596_
	);
	LUT2 #(
		.INIT('h4)
	) name26550 (
		_w30579_,
		_w30596_,
		_w30597_
	);
	LUT2 #(
		.INIT('h8)
	) name26551 (
		_w30594_,
		_w30595_,
		_w30598_
	);
	LUT2 #(
		.INIT('h8)
	) name26552 (
		_w30592_,
		_w30593_,
		_w30599_
	);
	LUT2 #(
		.INIT('h8)
	) name26553 (
		_w30590_,
		_w30591_,
		_w30600_
	);
	LUT2 #(
		.INIT('h8)
	) name26554 (
		_w29049_,
		_w29239_,
		_w30601_
	);
	LUT2 #(
		.INIT('h1)
	) name26555 (
		_w30564_,
		_w30565_,
		_w30602_
	);
	LUT2 #(
		.INIT('h1)
	) name26556 (
		_w30566_,
		_w30576_,
		_w30603_
	);
	LUT2 #(
		.INIT('h8)
	) name26557 (
		_w30602_,
		_w30603_,
		_w30604_
	);
	LUT2 #(
		.INIT('h8)
	) name26558 (
		_w30600_,
		_w30601_,
		_w30605_
	);
	LUT2 #(
		.INIT('h8)
	) name26559 (
		_w30598_,
		_w30599_,
		_w30606_
	);
	LUT2 #(
		.INIT('h8)
	) name26560 (
		_w18724_,
		_w30597_,
		_w30607_
	);
	LUT2 #(
		.INIT('h8)
	) name26561 (
		_w18796_,
		_w30607_,
		_w30608_
	);
	LUT2 #(
		.INIT('h8)
	) name26562 (
		_w30605_,
		_w30606_,
		_w30609_
	);
	LUT2 #(
		.INIT('h8)
	) name26563 (
		_w29252_,
		_w30604_,
		_w30610_
	);
	LUT2 #(
		.INIT('h8)
	) name26564 (
		_w30609_,
		_w30610_,
		_w30611_
	);
	LUT2 #(
		.INIT('h8)
	) name26565 (
		_w30608_,
		_w30611_,
		_w30612_
	);
	LUT2 #(
		.INIT('h8)
	) name26566 (
		_w20107_,
		_w30612_,
		_w30613_
	);
	LUT2 #(
		.INIT('h2)
	) name26567 (
		_w28627_,
		_w30613_,
		_w30614_
	);
	LUT2 #(
		.INIT('h8)
	) name26568 (
		_w12520_,
		_w28619_,
		_w30615_
	);
	LUT2 #(
		.INIT('h4)
	) name26569 (
		_w20326_,
		_w28636_,
		_w30616_
	);
	LUT2 #(
		.INIT('h1)
	) name26570 (
		_w7607_,
		_w28572_,
		_w30617_
	);
	LUT2 #(
		.INIT('h1)
	) name26571 (
		_w7473_,
		_w28598_,
		_w30618_
	);
	LUT2 #(
		.INIT('h1)
	) name26572 (
		_w7469_,
		_w28594_,
		_w30619_
	);
	LUT2 #(
		.INIT('h1)
	) name26573 (
		_w7449_,
		_w28589_,
		_w30620_
	);
	LUT2 #(
		.INIT('h1)
	) name26574 (
		_w30618_,
		_w30619_,
		_w30621_
	);
	LUT2 #(
		.INIT('h4)
	) name26575 (
		_w30620_,
		_w30621_,
		_w30622_
	);
	LUT2 #(
		.INIT('h8)
	) name26576 (
		_w28607_,
		_w30622_,
		_w30623_
	);
	LUT2 #(
		.INIT('h8)
	) name26577 (
		_w28572_,
		_w30623_,
		_w30624_
	);
	LUT2 #(
		.INIT('h2)
	) name26578 (
		_w28584_,
		_w30617_,
		_w30625_
	);
	LUT2 #(
		.INIT('h4)
	) name26579 (
		_w30624_,
		_w30625_,
		_w30626_
	);
	LUT2 #(
		.INIT('h1)
	) name26580 (
		_w30543_,
		_w30557_,
		_w30627_
	);
	LUT2 #(
		.INIT('h1)
	) name26581 (
		_w30615_,
		_w30616_,
		_w30628_
	);
	LUT2 #(
		.INIT('h8)
	) name26582 (
		_w30627_,
		_w30628_,
		_w30629_
	);
	LUT2 #(
		.INIT('h1)
	) name26583 (
		_w30555_,
		_w30556_,
		_w30630_
	);
	LUT2 #(
		.INIT('h8)
	) name26584 (
		_w30629_,
		_w30630_,
		_w30631_
	);
	LUT2 #(
		.INIT('h4)
	) name26585 (
		_w30614_,
		_w30631_,
		_w30632_
	);
	LUT2 #(
		.INIT('h4)
	) name26586 (
		_w30626_,
		_w30632_,
		_w30633_
	);
	LUT2 #(
		.INIT('h4)
	) name26587 (
		_w30554_,
		_w30633_,
		_w30634_
	);
	LUT2 #(
		.INIT('h4)
	) name26588 (
		_w30548_,
		_w30634_,
		_w30635_
	);
	LUT2 #(
		.INIT('h2)
	) name26589 (
		_w28550_,
		_w30635_,
		_w30636_
	);
	LUT2 #(
		.INIT('h4)
	) name26590 (
		\core_eu_em_mac_em_reg_mxopwe_DO_reg[0]/P0001 ,
		_w28649_,
		_w30637_
	);
	LUT2 #(
		.INIT('h8)
	) name26591 (
		_w7465_,
		_w28652_,
		_w30638_
	);
	LUT2 #(
		.INIT('h2)
	) name26592 (
		_w7457_,
		_w28652_,
		_w30639_
	);
	LUT2 #(
		.INIT('h1)
	) name26593 (
		_w28660_,
		_w30638_,
		_w30640_
	);
	LUT2 #(
		.INIT('h4)
	) name26594 (
		_w30639_,
		_w30640_,
		_w30641_
	);
	LUT2 #(
		.INIT('h8)
	) name26595 (
		_w19559_,
		_w28660_,
		_w30642_
	);
	LUT2 #(
		.INIT('h1)
	) name26596 (
		_w28649_,
		_w30641_,
		_w30643_
	);
	LUT2 #(
		.INIT('h4)
	) name26597 (
		_w30642_,
		_w30643_,
		_w30644_
	);
	LUT2 #(
		.INIT('h1)
	) name26598 (
		_w28550_,
		_w30637_,
		_w30645_
	);
	LUT2 #(
		.INIT('h4)
	) name26599 (
		_w30644_,
		_w30645_,
		_w30646_
	);
	LUT2 #(
		.INIT('h1)
	) name26600 (
		_w30636_,
		_w30646_,
		_w30647_
	);
	LUT2 #(
		.INIT('h8)
	) name26601 (
		_w12520_,
		_w28729_,
		_w30648_
	);
	LUT2 #(
		.INIT('h8)
	) name26602 (
		_w7607_,
		_w28725_,
		_w30649_
	);
	LUT2 #(
		.INIT('h8)
	) name26603 (
		_w7453_,
		_w28705_,
		_w30650_
	);
	LUT2 #(
		.INIT('h2)
	) name26604 (
		_w7461_,
		_w28705_,
		_w30651_
	);
	LUT2 #(
		.INIT('h1)
	) name26605 (
		_w30650_,
		_w30651_,
		_w30652_
	);
	LUT2 #(
		.INIT('h8)
	) name26606 (
		_w28735_,
		_w30652_,
		_w30653_
	);
	LUT2 #(
		.INIT('h8)
	) name26607 (
		_w28739_,
		_w30641_,
		_w30654_
	);
	LUT2 #(
		.INIT('h1)
	) name26608 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[0]/P0001 ,
		_w30655_
	);
	LUT2 #(
		.INIT('h2)
	) name26609 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[0]/P0001 ,
		_w30656_
	);
	LUT2 #(
		.INIT('h1)
	) name26610 (
		_w30655_,
		_w30656_,
		_w30657_
	);
	LUT2 #(
		.INIT('h8)
	) name26611 (
		_w28741_,
		_w30657_,
		_w30658_
	);
	LUT2 #(
		.INIT('h1)
	) name26612 (
		_w30653_,
		_w30654_,
		_w30659_
	);
	LUT2 #(
		.INIT('h4)
	) name26613 (
		_w30658_,
		_w30659_,
		_w30660_
	);
	LUT2 #(
		.INIT('h4)
	) name26614 (
		_w30648_,
		_w30660_,
		_w30661_
	);
	LUT2 #(
		.INIT('h4)
	) name26615 (
		_w30649_,
		_w30661_,
		_w30662_
	);
	LUT2 #(
		.INIT('h1)
	) name26616 (
		_w28543_,
		_w30662_,
		_w30663_
	);
	LUT2 #(
		.INIT('h2)
	) name26617 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[0]/P0001 ,
		_w28545_,
		_w30664_
	);
	LUT2 #(
		.INIT('h1)
	) name26618 (
		_w30663_,
		_w30664_,
		_w30665_
	);
	LUT2 #(
		.INIT('h1)
	) name26619 (
		_w28719_,
		_w30665_,
		_w30666_
	);
	LUT2 #(
		.INIT('h2)
	) name26620 (
		_w28719_,
		_w30635_,
		_w30667_
	);
	LUT2 #(
		.INIT('h1)
	) name26621 (
		_w30666_,
		_w30667_,
		_w30668_
	);
	LUT2 #(
		.INIT('h8)
	) name26622 (
		_w12870_,
		_w28729_,
		_w30669_
	);
	LUT2 #(
		.INIT('h8)
	) name26623 (
		_w8113_,
		_w28725_,
		_w30670_
	);
	LUT2 #(
		.INIT('h8)
	) name26624 (
		_w7897_,
		_w28705_,
		_w30671_
	);
	LUT2 #(
		.INIT('h2)
	) name26625 (
		_w7893_,
		_w28705_,
		_w30672_
	);
	LUT2 #(
		.INIT('h1)
	) name26626 (
		_w30671_,
		_w30672_,
		_w30673_
	);
	LUT2 #(
		.INIT('h8)
	) name26627 (
		_w28735_,
		_w30673_,
		_w30674_
	);
	LUT2 #(
		.INIT('h8)
	) name26628 (
		_w28739_,
		_w30536_,
		_w30675_
	);
	LUT2 #(
		.INIT('h1)
	) name26629 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[3]/P0001 ,
		_w30676_
	);
	LUT2 #(
		.INIT('h2)
	) name26630 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		\core_eu_em_mac_em_reg_mfswe_DO_reg[3]/P0001 ,
		_w30677_
	);
	LUT2 #(
		.INIT('h1)
	) name26631 (
		_w30676_,
		_w30677_,
		_w30678_
	);
	LUT2 #(
		.INIT('h8)
	) name26632 (
		_w28741_,
		_w30678_,
		_w30679_
	);
	LUT2 #(
		.INIT('h1)
	) name26633 (
		_w30674_,
		_w30675_,
		_w30680_
	);
	LUT2 #(
		.INIT('h4)
	) name26634 (
		_w30679_,
		_w30680_,
		_w30681_
	);
	LUT2 #(
		.INIT('h4)
	) name26635 (
		_w30669_,
		_w30681_,
		_w30682_
	);
	LUT2 #(
		.INIT('h4)
	) name26636 (
		_w30670_,
		_w30682_,
		_w30683_
	);
	LUT2 #(
		.INIT('h1)
	) name26637 (
		_w28543_,
		_w30683_,
		_w30684_
	);
	LUT2 #(
		.INIT('h2)
	) name26638 (
		\core_eu_em_mac_em_reg_myopwe_DO_reg[3]/P0001 ,
		_w28545_,
		_w30685_
	);
	LUT2 #(
		.INIT('h1)
	) name26639 (
		_w30684_,
		_w30685_,
		_w30686_
	);
	LUT2 #(
		.INIT('h1)
	) name26640 (
		_w28719_,
		_w30686_,
		_w30687_
	);
	LUT2 #(
		.INIT('h2)
	) name26641 (
		_w28719_,
		_w30530_,
		_w30688_
	);
	LUT2 #(
		.INIT('h1)
	) name26642 (
		_w30687_,
		_w30688_,
		_w30689_
	);
	LUT2 #(
		.INIT('h8)
	) name26643 (
		_w17805_,
		_w28530_,
		_w30690_
	);
	LUT2 #(
		.INIT('h8)
	) name26644 (
		_w19972_,
		_w30690_,
		_w30691_
	);
	LUT2 #(
		.INIT('h1)
	) name26645 (
		_w19385_,
		_w30691_,
		_w30692_
	);
	LUT2 #(
		.INIT('h2)
	) name26646 (
		_w28532_,
		_w30692_,
		_w30693_
	);
	LUT2 #(
		.INIT('h4)
	) name26647 (
		_w18268_,
		_w28534_,
		_w30694_
	);
	LUT2 #(
		.INIT('h2)
	) name26648 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[7]/P0001 ,
		_w30694_,
		_w30695_
	);
	LUT2 #(
		.INIT('h1)
	) name26649 (
		_w30693_,
		_w30695_,
		_w30696_
	);
	LUT2 #(
		.INIT('h1)
	) name26650 (
		_w18262_,
		_w30696_,
		_w30697_
	);
	LUT2 #(
		.INIT('h2)
	) name26651 (
		_w18262_,
		_w22883_,
		_w30698_
	);
	LUT2 #(
		.INIT('h1)
	) name26652 (
		_w30697_,
		_w30698_,
		_w30699_
	);
	LUT2 #(
		.INIT('h8)
	) name26653 (
		\tm_tcr_reg_DO_reg[1]/NET0131 ,
		_w20355_,
		_w30700_
	);
	LUT2 #(
		.INIT('h4)
	) name26654 (
		\tm_tpr_reg_DO_reg[1]/NET0131 ,
		_w22400_,
		_w30701_
	);
	LUT2 #(
		.INIT('h4)
	) name26655 (
		\tm_TCR_TMP_reg[0]/NET0131 ,
		_w22411_,
		_w30702_
	);
	LUT2 #(
		.INIT('h2)
	) name26656 (
		\tm_TCR_TMP_reg[1]/NET0131 ,
		_w30702_,
		_w30703_
	);
	LUT2 #(
		.INIT('h4)
	) name26657 (
		\tm_TCR_TMP_reg[1]/NET0131 ,
		_w30702_,
		_w30704_
	);
	LUT2 #(
		.INIT('h1)
	) name26658 (
		_w22400_,
		_w30703_,
		_w30705_
	);
	LUT2 #(
		.INIT('h4)
	) name26659 (
		_w30704_,
		_w30705_,
		_w30706_
	);
	LUT2 #(
		.INIT('h1)
	) name26660 (
		_w20355_,
		_w30701_,
		_w30707_
	);
	LUT2 #(
		.INIT('h4)
	) name26661 (
		_w30706_,
		_w30707_,
		_w30708_
	);
	LUT2 #(
		.INIT('h1)
	) name26662 (
		_w30700_,
		_w30708_,
		_w30709_
	);
	LUT2 #(
		.INIT('h8)
	) name26663 (
		\tm_tcr_reg_DO_reg[2]/NET0131 ,
		_w20355_,
		_w30710_
	);
	LUT2 #(
		.INIT('h4)
	) name26664 (
		\tm_tpr_reg_DO_reg[2]/NET0131 ,
		_w22400_,
		_w30711_
	);
	LUT2 #(
		.INIT('h4)
	) name26665 (
		\tm_TCR_TMP_reg[2]/NET0131 ,
		_w30704_,
		_w30712_
	);
	LUT2 #(
		.INIT('h2)
	) name26666 (
		\tm_TCR_TMP_reg[2]/NET0131 ,
		_w30704_,
		_w30713_
	);
	LUT2 #(
		.INIT('h1)
	) name26667 (
		_w22400_,
		_w30712_,
		_w30714_
	);
	LUT2 #(
		.INIT('h4)
	) name26668 (
		_w30713_,
		_w30714_,
		_w30715_
	);
	LUT2 #(
		.INIT('h1)
	) name26669 (
		_w20355_,
		_w30711_,
		_w30716_
	);
	LUT2 #(
		.INIT('h4)
	) name26670 (
		_w30715_,
		_w30716_,
		_w30717_
	);
	LUT2 #(
		.INIT('h1)
	) name26671 (
		_w30710_,
		_w30717_,
		_w30718_
	);
	LUT2 #(
		.INIT('h4)
	) name26672 (
		\tm_tpr_reg_DO_reg[6]/NET0131 ,
		_w22400_,
		_w30719_
	);
	LUT2 #(
		.INIT('h2)
	) name26673 (
		\tm_TCR_TMP_reg[6]/NET0131 ,
		_w27895_,
		_w30720_
	);
	LUT2 #(
		.INIT('h1)
	) name26674 (
		_w22400_,
		_w27896_,
		_w30721_
	);
	LUT2 #(
		.INIT('h4)
	) name26675 (
		_w30720_,
		_w30721_,
		_w30722_
	);
	LUT2 #(
		.INIT('h1)
	) name26676 (
		_w30719_,
		_w30722_,
		_w30723_
	);
	LUT2 #(
		.INIT('h1)
	) name26677 (
		_w20355_,
		_w30723_,
		_w30724_
	);
	LUT2 #(
		.INIT('h4)
	) name26678 (
		\tm_tcr_reg_DO_reg[6]/NET0131 ,
		_w20355_,
		_w30725_
	);
	LUT2 #(
		.INIT('h1)
	) name26679 (
		_w30724_,
		_w30725_,
		_w30726_
	);
	LUT2 #(
		.INIT('h8)
	) name26680 (
		\tm_tcr_reg_DO_reg[5]/NET0131 ,
		_w20355_,
		_w30727_
	);
	LUT2 #(
		.INIT('h4)
	) name26681 (
		\tm_tpr_reg_DO_reg[5]/NET0131 ,
		_w22400_,
		_w30728_
	);
	LUT2 #(
		.INIT('h8)
	) name26682 (
		\tm_TCR_TMP_reg[4]/NET0131 ,
		_w27890_,
		_w30729_
	);
	LUT2 #(
		.INIT('h8)
	) name26683 (
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w30729_,
		_w30730_
	);
	LUT2 #(
		.INIT('h1)
	) name26684 (
		_w27894_,
		_w30730_,
		_w30731_
	);
	LUT2 #(
		.INIT('h2)
	) name26685 (
		_w22411_,
		_w30731_,
		_w30732_
	);
	LUT2 #(
		.INIT('h1)
	) name26686 (
		_w27893_,
		_w30729_,
		_w30733_
	);
	LUT2 #(
		.INIT('h2)
	) name26687 (
		_w22411_,
		_w30733_,
		_w30734_
	);
	LUT2 #(
		.INIT('h2)
	) name26688 (
		\tm_TCR_TMP_reg[5]/NET0131 ,
		_w30734_,
		_w30735_
	);
	LUT2 #(
		.INIT('h1)
	) name26689 (
		_w22400_,
		_w30732_,
		_w30736_
	);
	LUT2 #(
		.INIT('h4)
	) name26690 (
		_w30735_,
		_w30736_,
		_w30737_
	);
	LUT2 #(
		.INIT('h1)
	) name26691 (
		_w20355_,
		_w30728_,
		_w30738_
	);
	LUT2 #(
		.INIT('h4)
	) name26692 (
		_w30737_,
		_w30738_,
		_w30739_
	);
	LUT2 #(
		.INIT('h1)
	) name26693 (
		_w30727_,
		_w30739_,
		_w30740_
	);
	LUT2 #(
		.INIT('h4)
	) name26694 (
		\sport1_cfg_RFSg_d1_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w30741_
	);
	LUT2 #(
		.INIT('h4)
	) name26695 (
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w30741_,
		_w30742_
	);
	LUT2 #(
		.INIT('h4)
	) name26696 (
		_w21382_,
		_w22650_,
		_w30743_
	);
	LUT2 #(
		.INIT('h2)
	) name26697 (
		\sport1_cfg_RFSg_d2_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w30744_
	);
	LUT2 #(
		.INIT('h8)
	) name26698 (
		\sport1_cfg_RFSg_d3_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w30745_
	);
	LUT2 #(
		.INIT('h2)
	) name26699 (
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w30744_,
		_w30746_
	);
	LUT2 #(
		.INIT('h4)
	) name26700 (
		_w30745_,
		_w30746_,
		_w30747_
	);
	LUT2 #(
		.INIT('h1)
	) name26701 (
		_w30742_,
		_w30747_,
		_w30748_
	);
	LUT2 #(
		.INIT('h4)
	) name26702 (
		_w30743_,
		_w30748_,
		_w30749_
	);
	LUT2 #(
		.INIT('h2)
	) name26703 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		_w30749_,
		_w30750_
	);
	LUT2 #(
		.INIT('h1)
	) name26704 (
		\sport1_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[1]/NET0131 ,
		_w30751_
	);
	LUT2 #(
		.INIT('h4)
	) name26705 (
		\sport1_rxctl_LMcnt_reg[2]/NET0131 ,
		_w30751_,
		_w30752_
	);
	LUT2 #(
		.INIT('h4)
	) name26706 (
		\sport1_rxctl_LMcnt_reg[3]/NET0131 ,
		_w30752_,
		_w30753_
	);
	LUT2 #(
		.INIT('h4)
	) name26707 (
		\sport1_rxctl_LMcnt_reg[4]/NET0131 ,
		_w30753_,
		_w30754_
	);
	LUT2 #(
		.INIT('h1)
	) name26708 (
		_w30750_,
		_w30754_,
		_w30755_
	);
	LUT2 #(
		.INIT('h2)
	) name26709 (
		\sport1_rxctl_RXSHT_reg[15]/P0001 ,
		_w30755_,
		_w30756_
	);
	LUT2 #(
		.INIT('h4)
	) name26710 (
		\sport1_rxctl_sht2nd_reg/P0001 ,
		_w30755_,
		_w30757_
	);
	LUT2 #(
		.INIT('h8)
	) name26711 (
		\sport1_rxctl_RXSHT_reg[14]/P0001 ,
		_w30757_,
		_w30758_
	);
	LUT2 #(
		.INIT('h1)
	) name26712 (
		\sport1_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w30759_
	);
	LUT2 #(
		.INIT('h8)
	) name26713 (
		\sport1_rxctl_RXSHT_reg[0]/P0001 ,
		_w30755_,
		_w30760_
	);
	LUT2 #(
		.INIT('h2)
	) name26714 (
		\sport1_rxctl_sht2nd_reg/P0001 ,
		_w30759_,
		_w30761_
	);
	LUT2 #(
		.INIT('h8)
	) name26715 (
		_w30760_,
		_w30761_,
		_w30762_
	);
	LUT2 #(
		.INIT('h1)
	) name26716 (
		_w30756_,
		_w30758_,
		_w30763_
	);
	LUT2 #(
		.INIT('h4)
	) name26717 (
		_w30762_,
		_w30763_,
		_w30764_
	);
	LUT2 #(
		.INIT('h4)
	) name26718 (
		\sport0_cfg_RFSg_d1_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w30765_
	);
	LUT2 #(
		.INIT('h4)
	) name26719 (
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w30765_,
		_w30766_
	);
	LUT2 #(
		.INIT('h2)
	) name26720 (
		_w19933_,
		_w21390_,
		_w30767_
	);
	LUT2 #(
		.INIT('h2)
	) name26721 (
		\sport0_cfg_RFSg_d2_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w30768_
	);
	LUT2 #(
		.INIT('h8)
	) name26722 (
		\sport0_cfg_RFSg_d3_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w30769_
	);
	LUT2 #(
		.INIT('h2)
	) name26723 (
		\sport0_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w30768_,
		_w30770_
	);
	LUT2 #(
		.INIT('h4)
	) name26724 (
		_w30769_,
		_w30770_,
		_w30771_
	);
	LUT2 #(
		.INIT('h1)
	) name26725 (
		_w30766_,
		_w30771_,
		_w30772_
	);
	LUT2 #(
		.INIT('h4)
	) name26726 (
		_w30767_,
		_w30772_,
		_w30773_
	);
	LUT2 #(
		.INIT('h2)
	) name26727 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		_w30773_,
		_w30774_
	);
	LUT2 #(
		.INIT('h1)
	) name26728 (
		\sport0_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[1]/NET0131 ,
		_w30775_
	);
	LUT2 #(
		.INIT('h4)
	) name26729 (
		\sport0_rxctl_LMcnt_reg[2]/NET0131 ,
		_w30775_,
		_w30776_
	);
	LUT2 #(
		.INIT('h4)
	) name26730 (
		\sport0_rxctl_LMcnt_reg[3]/NET0131 ,
		_w30776_,
		_w30777_
	);
	LUT2 #(
		.INIT('h4)
	) name26731 (
		\sport0_rxctl_LMcnt_reg[4]/NET0131 ,
		_w30777_,
		_w30778_
	);
	LUT2 #(
		.INIT('h1)
	) name26732 (
		_w30774_,
		_w30778_,
		_w30779_
	);
	LUT2 #(
		.INIT('h2)
	) name26733 (
		\sport0_rxctl_RXSHT_reg[10]/P0001 ,
		_w30779_,
		_w30780_
	);
	LUT2 #(
		.INIT('h4)
	) name26734 (
		\sport0_rxctl_sht2nd_reg/P0001 ,
		_w30779_,
		_w30781_
	);
	LUT2 #(
		.INIT('h8)
	) name26735 (
		\sport0_rxctl_RXSHT_reg[9]/P0001 ,
		_w30781_,
		_w30782_
	);
	LUT2 #(
		.INIT('h1)
	) name26736 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w30783_
	);
	LUT2 #(
		.INIT('h8)
	) name26737 (
		\sport0_rxctl_RXSHT_reg[0]/P0001 ,
		_w30779_,
		_w30784_
	);
	LUT2 #(
		.INIT('h2)
	) name26738 (
		\sport0_rxctl_sht2nd_reg/P0001 ,
		_w30783_,
		_w30785_
	);
	LUT2 #(
		.INIT('h8)
	) name26739 (
		_w30784_,
		_w30785_,
		_w30786_
	);
	LUT2 #(
		.INIT('h1)
	) name26740 (
		_w30780_,
		_w30782_,
		_w30787_
	);
	LUT2 #(
		.INIT('h4)
	) name26741 (
		_w30786_,
		_w30787_,
		_w30788_
	);
	LUT2 #(
		.INIT('h2)
	) name26742 (
		\sport1_rxctl_RXSHT_reg[10]/P0001 ,
		_w30755_,
		_w30789_
	);
	LUT2 #(
		.INIT('h8)
	) name26743 (
		\sport1_rxctl_RXSHT_reg[9]/P0001 ,
		_w30757_,
		_w30790_
	);
	LUT2 #(
		.INIT('h1)
	) name26744 (
		_w30762_,
		_w30789_,
		_w30791_
	);
	LUT2 #(
		.INIT('h4)
	) name26745 (
		_w30790_,
		_w30791_,
		_w30792_
	);
	LUT2 #(
		.INIT('h2)
	) name26746 (
		\sport1_rxctl_RXSHT_reg[11]/P0001 ,
		_w30755_,
		_w30793_
	);
	LUT2 #(
		.INIT('h8)
	) name26747 (
		\sport1_rxctl_RXSHT_reg[10]/P0001 ,
		_w30757_,
		_w30794_
	);
	LUT2 #(
		.INIT('h1)
	) name26748 (
		_w30762_,
		_w30793_,
		_w30795_
	);
	LUT2 #(
		.INIT('h4)
	) name26749 (
		_w30794_,
		_w30795_,
		_w30796_
	);
	LUT2 #(
		.INIT('h8)
	) name26750 (
		_w18262_,
		_w22926_,
		_w30797_
	);
	LUT2 #(
		.INIT('h2)
	) name26751 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[6]/P0001 ,
		_w28534_,
		_w30798_
	);
	LUT2 #(
		.INIT('h8)
	) name26752 (
		_w18276_,
		_w30690_,
		_w30799_
	);
	LUT2 #(
		.INIT('h1)
	) name26753 (
		_w19385_,
		_w30799_,
		_w30800_
	);
	LUT2 #(
		.INIT('h2)
	) name26754 (
		_w28532_,
		_w30800_,
		_w30801_
	);
	LUT2 #(
		.INIT('h2)
	) name26755 (
		_w28529_,
		_w30798_,
		_w30802_
	);
	LUT2 #(
		.INIT('h4)
	) name26756 (
		_w30801_,
		_w30802_,
		_w30803_
	);
	LUT2 #(
		.INIT('h1)
	) name26757 (
		_w30797_,
		_w30803_,
		_w30804_
	);
	LUT2 #(
		.INIT('h2)
	) name26758 (
		\sport1_rxctl_RXSHT_reg[12]/P0001 ,
		_w30755_,
		_w30805_
	);
	LUT2 #(
		.INIT('h8)
	) name26759 (
		\sport1_rxctl_RXSHT_reg[11]/P0001 ,
		_w30757_,
		_w30806_
	);
	LUT2 #(
		.INIT('h1)
	) name26760 (
		_w30762_,
		_w30805_,
		_w30807_
	);
	LUT2 #(
		.INIT('h4)
	) name26761 (
		_w30806_,
		_w30807_,
		_w30808_
	);
	LUT2 #(
		.INIT('h2)
	) name26762 (
		\sport1_rxctl_RXSHT_reg[13]/P0001 ,
		_w30755_,
		_w30809_
	);
	LUT2 #(
		.INIT('h8)
	) name26763 (
		\sport1_rxctl_RXSHT_reg[12]/P0001 ,
		_w30757_,
		_w30810_
	);
	LUT2 #(
		.INIT('h1)
	) name26764 (
		_w30762_,
		_w30809_,
		_w30811_
	);
	LUT2 #(
		.INIT('h4)
	) name26765 (
		_w30810_,
		_w30811_,
		_w30812_
	);
	LUT2 #(
		.INIT('h2)
	) name26766 (
		\sport1_rxctl_RXSHT_reg[14]/P0001 ,
		_w30755_,
		_w30813_
	);
	LUT2 #(
		.INIT('h8)
	) name26767 (
		\sport1_rxctl_RXSHT_reg[13]/P0001 ,
		_w30757_,
		_w30814_
	);
	LUT2 #(
		.INIT('h1)
	) name26768 (
		_w30762_,
		_w30813_,
		_w30815_
	);
	LUT2 #(
		.INIT('h4)
	) name26769 (
		_w30814_,
		_w30815_,
		_w30816_
	);
	LUT2 #(
		.INIT('h2)
	) name26770 (
		\sport1_rxctl_RXSHT_reg[2]/P0001 ,
		_w30755_,
		_w30817_
	);
	LUT2 #(
		.INIT('h8)
	) name26771 (
		\sport1_rxctl_RXSHT_reg[1]/P0001 ,
		_w30757_,
		_w30818_
	);
	LUT2 #(
		.INIT('h1)
	) name26772 (
		_w30762_,
		_w30817_,
		_w30819_
	);
	LUT2 #(
		.INIT('h4)
	) name26773 (
		_w30818_,
		_w30819_,
		_w30820_
	);
	LUT2 #(
		.INIT('h2)
	) name26774 (
		\sport1_rxctl_RXSHT_reg[3]/P0001 ,
		_w30755_,
		_w30821_
	);
	LUT2 #(
		.INIT('h8)
	) name26775 (
		\sport1_rxctl_RXSHT_reg[2]/P0001 ,
		_w30757_,
		_w30822_
	);
	LUT2 #(
		.INIT('h1)
	) name26776 (
		_w30762_,
		_w30821_,
		_w30823_
	);
	LUT2 #(
		.INIT('h4)
	) name26777 (
		_w30822_,
		_w30823_,
		_w30824_
	);
	LUT2 #(
		.INIT('h2)
	) name26778 (
		\sport1_rxctl_RXSHT_reg[4]/P0001 ,
		_w30755_,
		_w30825_
	);
	LUT2 #(
		.INIT('h8)
	) name26779 (
		\sport1_rxctl_RXSHT_reg[3]/P0001 ,
		_w30757_,
		_w30826_
	);
	LUT2 #(
		.INIT('h1)
	) name26780 (
		_w30762_,
		_w30825_,
		_w30827_
	);
	LUT2 #(
		.INIT('h4)
	) name26781 (
		_w30826_,
		_w30827_,
		_w30828_
	);
	LUT2 #(
		.INIT('h2)
	) name26782 (
		\sport1_rxctl_RXSHT_reg[5]/P0001 ,
		_w30755_,
		_w30829_
	);
	LUT2 #(
		.INIT('h8)
	) name26783 (
		\sport1_rxctl_RXSHT_reg[4]/P0001 ,
		_w30757_,
		_w30830_
	);
	LUT2 #(
		.INIT('h1)
	) name26784 (
		_w30762_,
		_w30829_,
		_w30831_
	);
	LUT2 #(
		.INIT('h4)
	) name26785 (
		_w30830_,
		_w30831_,
		_w30832_
	);
	LUT2 #(
		.INIT('h2)
	) name26786 (
		\sport1_rxctl_RXSHT_reg[6]/P0001 ,
		_w30755_,
		_w30833_
	);
	LUT2 #(
		.INIT('h8)
	) name26787 (
		\sport1_rxctl_RXSHT_reg[5]/P0001 ,
		_w30757_,
		_w30834_
	);
	LUT2 #(
		.INIT('h1)
	) name26788 (
		_w30762_,
		_w30833_,
		_w30835_
	);
	LUT2 #(
		.INIT('h4)
	) name26789 (
		_w30834_,
		_w30835_,
		_w30836_
	);
	LUT2 #(
		.INIT('h2)
	) name26790 (
		\sport1_rxctl_RXSHT_reg[8]/P0001 ,
		_w30755_,
		_w30837_
	);
	LUT2 #(
		.INIT('h8)
	) name26791 (
		\sport1_rxctl_RXSHT_reg[7]/P0001 ,
		_w30757_,
		_w30838_
	);
	LUT2 #(
		.INIT('h1)
	) name26792 (
		_w30762_,
		_w30837_,
		_w30839_
	);
	LUT2 #(
		.INIT('h4)
	) name26793 (
		_w30838_,
		_w30839_,
		_w30840_
	);
	LUT2 #(
		.INIT('h2)
	) name26794 (
		\sport1_rxctl_RXSHT_reg[9]/P0001 ,
		_w30755_,
		_w30841_
	);
	LUT2 #(
		.INIT('h8)
	) name26795 (
		\sport1_rxctl_RXSHT_reg[8]/P0001 ,
		_w30757_,
		_w30842_
	);
	LUT2 #(
		.INIT('h1)
	) name26796 (
		_w30762_,
		_w30841_,
		_w30843_
	);
	LUT2 #(
		.INIT('h4)
	) name26797 (
		_w30842_,
		_w30843_,
		_w30844_
	);
	LUT2 #(
		.INIT('h2)
	) name26798 (
		\sport0_rxctl_RXSHT_reg[11]/P0001 ,
		_w30779_,
		_w30845_
	);
	LUT2 #(
		.INIT('h8)
	) name26799 (
		\sport0_rxctl_RXSHT_reg[10]/P0001 ,
		_w30781_,
		_w30846_
	);
	LUT2 #(
		.INIT('h1)
	) name26800 (
		_w30786_,
		_w30845_,
		_w30847_
	);
	LUT2 #(
		.INIT('h4)
	) name26801 (
		_w30846_,
		_w30847_,
		_w30848_
	);
	LUT2 #(
		.INIT('h2)
	) name26802 (
		\sport0_rxctl_RXSHT_reg[14]/P0001 ,
		_w30779_,
		_w30849_
	);
	LUT2 #(
		.INIT('h8)
	) name26803 (
		\sport0_rxctl_RXSHT_reg[13]/P0001 ,
		_w30781_,
		_w30850_
	);
	LUT2 #(
		.INIT('h1)
	) name26804 (
		_w30786_,
		_w30849_,
		_w30851_
	);
	LUT2 #(
		.INIT('h4)
	) name26805 (
		_w30850_,
		_w30851_,
		_w30852_
	);
	LUT2 #(
		.INIT('h2)
	) name26806 (
		\sport0_rxctl_RXSHT_reg[15]/P0001 ,
		_w30779_,
		_w30853_
	);
	LUT2 #(
		.INIT('h8)
	) name26807 (
		\sport0_rxctl_RXSHT_reg[14]/P0001 ,
		_w30781_,
		_w30854_
	);
	LUT2 #(
		.INIT('h1)
	) name26808 (
		_w30786_,
		_w30853_,
		_w30855_
	);
	LUT2 #(
		.INIT('h4)
	) name26809 (
		_w30854_,
		_w30855_,
		_w30856_
	);
	LUT2 #(
		.INIT('h2)
	) name26810 (
		\sport0_rxctl_RXSHT_reg[2]/P0001 ,
		_w30779_,
		_w30857_
	);
	LUT2 #(
		.INIT('h8)
	) name26811 (
		\sport0_rxctl_RXSHT_reg[1]/P0001 ,
		_w30781_,
		_w30858_
	);
	LUT2 #(
		.INIT('h1)
	) name26812 (
		_w30786_,
		_w30857_,
		_w30859_
	);
	LUT2 #(
		.INIT('h4)
	) name26813 (
		_w30858_,
		_w30859_,
		_w30860_
	);
	LUT2 #(
		.INIT('h2)
	) name26814 (
		\sport0_rxctl_RXSHT_reg[3]/P0001 ,
		_w30779_,
		_w30861_
	);
	LUT2 #(
		.INIT('h8)
	) name26815 (
		\sport0_rxctl_RXSHT_reg[2]/P0001 ,
		_w30781_,
		_w30862_
	);
	LUT2 #(
		.INIT('h1)
	) name26816 (
		_w30786_,
		_w30861_,
		_w30863_
	);
	LUT2 #(
		.INIT('h4)
	) name26817 (
		_w30862_,
		_w30863_,
		_w30864_
	);
	LUT2 #(
		.INIT('h2)
	) name26818 (
		\sport0_rxctl_RXSHT_reg[4]/P0001 ,
		_w30779_,
		_w30865_
	);
	LUT2 #(
		.INIT('h8)
	) name26819 (
		\sport0_rxctl_RXSHT_reg[3]/P0001 ,
		_w30781_,
		_w30866_
	);
	LUT2 #(
		.INIT('h1)
	) name26820 (
		_w30786_,
		_w30865_,
		_w30867_
	);
	LUT2 #(
		.INIT('h4)
	) name26821 (
		_w30866_,
		_w30867_,
		_w30868_
	);
	LUT2 #(
		.INIT('h2)
	) name26822 (
		\sport0_rxctl_RXSHT_reg[5]/P0001 ,
		_w30779_,
		_w30869_
	);
	LUT2 #(
		.INIT('h8)
	) name26823 (
		\sport0_rxctl_RXSHT_reg[4]/P0001 ,
		_w30781_,
		_w30870_
	);
	LUT2 #(
		.INIT('h1)
	) name26824 (
		_w30786_,
		_w30869_,
		_w30871_
	);
	LUT2 #(
		.INIT('h4)
	) name26825 (
		_w30870_,
		_w30871_,
		_w30872_
	);
	LUT2 #(
		.INIT('h2)
	) name26826 (
		\sport0_rxctl_RXSHT_reg[6]/P0001 ,
		_w30779_,
		_w30873_
	);
	LUT2 #(
		.INIT('h8)
	) name26827 (
		\sport0_rxctl_RXSHT_reg[5]/P0001 ,
		_w30781_,
		_w30874_
	);
	LUT2 #(
		.INIT('h1)
	) name26828 (
		_w30786_,
		_w30873_,
		_w30875_
	);
	LUT2 #(
		.INIT('h4)
	) name26829 (
		_w30874_,
		_w30875_,
		_w30876_
	);
	LUT2 #(
		.INIT('h2)
	) name26830 (
		\sport0_rxctl_RXSHT_reg[7]/P0001 ,
		_w30779_,
		_w30877_
	);
	LUT2 #(
		.INIT('h8)
	) name26831 (
		\sport0_rxctl_RXSHT_reg[6]/P0001 ,
		_w30781_,
		_w30878_
	);
	LUT2 #(
		.INIT('h1)
	) name26832 (
		_w30786_,
		_w30877_,
		_w30879_
	);
	LUT2 #(
		.INIT('h4)
	) name26833 (
		_w30878_,
		_w30879_,
		_w30880_
	);
	LUT2 #(
		.INIT('h2)
	) name26834 (
		\sport0_rxctl_RXSHT_reg[8]/P0001 ,
		_w30779_,
		_w30881_
	);
	LUT2 #(
		.INIT('h8)
	) name26835 (
		\sport0_rxctl_RXSHT_reg[7]/P0001 ,
		_w30781_,
		_w30882_
	);
	LUT2 #(
		.INIT('h1)
	) name26836 (
		_w30786_,
		_w30881_,
		_w30883_
	);
	LUT2 #(
		.INIT('h4)
	) name26837 (
		_w30882_,
		_w30883_,
		_w30884_
	);
	LUT2 #(
		.INIT('h2)
	) name26838 (
		\sport0_rxctl_RXSHT_reg[9]/P0001 ,
		_w30779_,
		_w30885_
	);
	LUT2 #(
		.INIT('h8)
	) name26839 (
		\sport0_rxctl_RXSHT_reg[8]/P0001 ,
		_w30781_,
		_w30886_
	);
	LUT2 #(
		.INIT('h1)
	) name26840 (
		_w30786_,
		_w30885_,
		_w30887_
	);
	LUT2 #(
		.INIT('h4)
	) name26841 (
		_w30886_,
		_w30887_,
		_w30888_
	);
	LUT2 #(
		.INIT('h2)
	) name26842 (
		\sport1_rxctl_RXSHT_reg[7]/P0001 ,
		_w30755_,
		_w30889_
	);
	LUT2 #(
		.INIT('h8)
	) name26843 (
		\sport1_rxctl_RXSHT_reg[6]/P0001 ,
		_w30757_,
		_w30890_
	);
	LUT2 #(
		.INIT('h1)
	) name26844 (
		_w30762_,
		_w30889_,
		_w30891_
	);
	LUT2 #(
		.INIT('h4)
	) name26845 (
		_w30890_,
		_w30891_,
		_w30892_
	);
	LUT2 #(
		.INIT('h2)
	) name26846 (
		\sport0_rxctl_RXSHT_reg[13]/P0001 ,
		_w30779_,
		_w30893_
	);
	LUT2 #(
		.INIT('h8)
	) name26847 (
		\sport0_rxctl_RXSHT_reg[12]/P0001 ,
		_w30781_,
		_w30894_
	);
	LUT2 #(
		.INIT('h1)
	) name26848 (
		_w30786_,
		_w30893_,
		_w30895_
	);
	LUT2 #(
		.INIT('h4)
	) name26849 (
		_w30894_,
		_w30895_,
		_w30896_
	);
	LUT2 #(
		.INIT('h2)
	) name26850 (
		\sport0_rxctl_RXSHT_reg[12]/P0001 ,
		_w30779_,
		_w30897_
	);
	LUT2 #(
		.INIT('h8)
	) name26851 (
		\sport0_rxctl_RXSHT_reg[11]/P0001 ,
		_w30781_,
		_w30898_
	);
	LUT2 #(
		.INIT('h1)
	) name26852 (
		_w30786_,
		_w30897_,
		_w30899_
	);
	LUT2 #(
		.INIT('h4)
	) name26853 (
		_w30898_,
		_w30899_,
		_w30900_
	);
	LUT2 #(
		.INIT('h4)
	) name26854 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w19205_,
		_w30901_
	);
	LUT2 #(
		.INIT('h4)
	) name26855 (
		_w19205_,
		_w19243_,
		_w30902_
	);
	LUT2 #(
		.INIT('h2)
	) name26856 (
		_w4150_,
		_w30901_,
		_w30903_
	);
	LUT2 #(
		.INIT('h4)
	) name26857 (
		_w30902_,
		_w30903_,
		_w30904_
	);
	LUT2 #(
		.INIT('h8)
	) name26858 (
		_w17799_,
		_w17805_,
		_w30905_
	);
	LUT2 #(
		.INIT('h8)
	) name26859 (
		_w19972_,
		_w30905_,
		_w30906_
	);
	LUT2 #(
		.INIT('h1)
	) name26860 (
		_w17823_,
		_w30906_,
		_w30907_
	);
	LUT2 #(
		.INIT('h2)
	) name26861 (
		_w17808_,
		_w30907_,
		_w30908_
	);
	LUT2 #(
		.INIT('h2)
	) name26862 (
		_w17811_,
		_w17827_,
		_w30909_
	);
	LUT2 #(
		.INIT('h2)
	) name26863 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[7]/P0001 ,
		_w30909_,
		_w30910_
	);
	LUT2 #(
		.INIT('h1)
	) name26864 (
		_w30908_,
		_w30910_,
		_w30911_
	);
	LUT2 #(
		.INIT('h1)
	) name26865 (
		_w14752_,
		_w30911_,
		_w30912_
	);
	LUT2 #(
		.INIT('h2)
	) name26866 (
		_w14752_,
		_w22883_,
		_w30913_
	);
	LUT2 #(
		.INIT('h1)
	) name26867 (
		_w30912_,
		_w30913_,
		_w30914_
	);
	LUT2 #(
		.INIT('h8)
	) name26868 (
		\tm_tcr_reg_DO_reg[13]/NET0131 ,
		_w20355_,
		_w30915_
	);
	LUT2 #(
		.INIT('h4)
	) name26869 (
		\tm_tpr_reg_DO_reg[13]/NET0131 ,
		_w22400_,
		_w30916_
	);
	LUT2 #(
		.INIT('h2)
	) name26870 (
		\tm_TCR_TMP_reg[13]/NET0131 ,
		_w25840_,
		_w30917_
	);
	LUT2 #(
		.INIT('h1)
	) name26871 (
		_w22400_,
		_w25841_,
		_w30918_
	);
	LUT2 #(
		.INIT('h4)
	) name26872 (
		_w30917_,
		_w30918_,
		_w30919_
	);
	LUT2 #(
		.INIT('h1)
	) name26873 (
		_w20355_,
		_w30916_,
		_w30920_
	);
	LUT2 #(
		.INIT('h4)
	) name26874 (
		_w30919_,
		_w30920_,
		_w30921_
	);
	LUT2 #(
		.INIT('h1)
	) name26875 (
		_w30915_,
		_w30921_,
		_w30922_
	);
	LUT2 #(
		.INIT('h8)
	) name26876 (
		_w14752_,
		_w22926_,
		_w30923_
	);
	LUT2 #(
		.INIT('h1)
	) name26877 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 ,
		_w17799_,
		_w30924_
	);
	LUT2 #(
		.INIT('h4)
	) name26878 (
		_w17809_,
		_w18276_,
		_w30925_
	);
	LUT2 #(
		.INIT('h2)
	) name26879 (
		_w17811_,
		_w30925_,
		_w30926_
	);
	LUT2 #(
		.INIT('h1)
	) name26880 (
		_w30924_,
		_w30926_,
		_w30927_
	);
	LUT2 #(
		.INIT('h1)
	) name26881 (
		_w17823_,
		_w30927_,
		_w30928_
	);
	LUT2 #(
		.INIT('h1)
	) name26882 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[6]/P0001 ,
		_w17808_,
		_w30929_
	);
	LUT2 #(
		.INIT('h1)
	) name26883 (
		_w30928_,
		_w30929_,
		_w30930_
	);
	LUT2 #(
		.INIT('h2)
	) name26884 (
		_w17829_,
		_w30930_,
		_w30931_
	);
	LUT2 #(
		.INIT('h1)
	) name26885 (
		_w30923_,
		_w30931_,
		_w30932_
	);
	LUT2 #(
		.INIT('h8)
	) name26886 (
		\core_c_dec_pMFMAC_Ei_reg/NET0131 ,
		_w4117_,
		_w30933_
	);
	LUT2 #(
		.INIT('h1)
	) name26887 (
		_w4117_,
		_w19701_,
		_w30934_
	);
	LUT2 #(
		.INIT('h8)
	) name26888 (
		_w6028_,
		_w19696_,
		_w30935_
	);
	LUT2 #(
		.INIT('h1)
	) name26889 (
		_w24644_,
		_w30935_,
		_w30936_
	);
	LUT2 #(
		.INIT('h8)
	) name26890 (
		_w6028_,
		_w21248_,
		_w30937_
	);
	LUT2 #(
		.INIT('h4)
	) name26891 (
		_w6024_,
		_w6119_,
		_w30938_
	);
	LUT2 #(
		.INIT('h8)
	) name26892 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w30938_,
		_w30939_
	);
	LUT2 #(
		.INIT('h1)
	) name26893 (
		_w18839_,
		_w25469_,
		_w30940_
	);
	LUT2 #(
		.INIT('h4)
	) name26894 (
		_w24646_,
		_w30940_,
		_w30941_
	);
	LUT2 #(
		.INIT('h4)
	) name26895 (
		_w30937_,
		_w30941_,
		_w30942_
	);
	LUT2 #(
		.INIT('h2)
	) name26896 (
		_w30936_,
		_w30939_,
		_w30943_
	);
	LUT2 #(
		.INIT('h8)
	) name26897 (
		_w30942_,
		_w30943_,
		_w30944_
	);
	LUT2 #(
		.INIT('h8)
	) name26898 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w6028_,
		_w30945_
	);
	LUT2 #(
		.INIT('h1)
	) name26899 (
		_w6956_,
		_w18839_,
		_w30946_
	);
	LUT2 #(
		.INIT('h4)
	) name26900 (
		_w25081_,
		_w30946_,
		_w30947_
	);
	LUT2 #(
		.INIT('h4)
	) name26901 (
		_w30945_,
		_w30947_,
		_w30948_
	);
	LUT2 #(
		.INIT('h2)
	) name26902 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w30948_,
		_w30949_
	);
	LUT2 #(
		.INIT('h8)
	) name26903 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w30948_,
		_w30950_
	);
	LUT2 #(
		.INIT('h1)
	) name26904 (
		_w30949_,
		_w30950_,
		_w30951_
	);
	LUT2 #(
		.INIT('h1)
	) name26905 (
		_w30944_,
		_w30951_,
		_w30952_
	);
	LUT2 #(
		.INIT('h4)
	) name26906 (
		_w6116_,
		_w6956_,
		_w30953_
	);
	LUT2 #(
		.INIT('h4)
	) name26907 (
		_w26373_,
		_w30935_,
		_w30954_
	);
	LUT2 #(
		.INIT('h1)
	) name26908 (
		_w30953_,
		_w30954_,
		_w30955_
	);
	LUT2 #(
		.INIT('h2)
	) name26909 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w30948_,
		_w30956_
	);
	LUT2 #(
		.INIT('h8)
	) name26910 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w30948_,
		_w30957_
	);
	LUT2 #(
		.INIT('h1)
	) name26911 (
		_w30956_,
		_w30957_,
		_w30958_
	);
	LUT2 #(
		.INIT('h2)
	) name26912 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w30948_,
		_w30959_
	);
	LUT2 #(
		.INIT('h8)
	) name26913 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w30948_,
		_w30960_
	);
	LUT2 #(
		.INIT('h1)
	) name26914 (
		_w30959_,
		_w30960_,
		_w30961_
	);
	LUT2 #(
		.INIT('h2)
	) name26915 (
		_w30958_,
		_w30961_,
		_w30962_
	);
	LUT2 #(
		.INIT('h8)
	) name26916 (
		_w30955_,
		_w30962_,
		_w30963_
	);
	LUT2 #(
		.INIT('h2)
	) name26917 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w30948_,
		_w30964_
	);
	LUT2 #(
		.INIT('h8)
	) name26918 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w30948_,
		_w30965_
	);
	LUT2 #(
		.INIT('h1)
	) name26919 (
		_w30964_,
		_w30965_,
		_w30966_
	);
	LUT2 #(
		.INIT('h2)
	) name26920 (
		_w30963_,
		_w30966_,
		_w30967_
	);
	LUT2 #(
		.INIT('h8)
	) name26921 (
		_w30952_,
		_w30967_,
		_w30968_
	);
	LUT2 #(
		.INIT('h1)
	) name26922 (
		_w30958_,
		_w30961_,
		_w30969_
	);
	LUT2 #(
		.INIT('h8)
	) name26923 (
		_w30952_,
		_w30955_,
		_w30970_
	);
	LUT2 #(
		.INIT('h8)
	) name26924 (
		_w30966_,
		_w30970_,
		_w30971_
	);
	LUT2 #(
		.INIT('h8)
	) name26925 (
		_w30969_,
		_w30971_,
		_w30972_
	);
	LUT2 #(
		.INIT('h4)
	) name26926 (
		_w30944_,
		_w30951_,
		_w30973_
	);
	LUT2 #(
		.INIT('h8)
	) name26927 (
		_w30955_,
		_w30973_,
		_w30974_
	);
	LUT2 #(
		.INIT('h8)
	) name26928 (
		_w30966_,
		_w30974_,
		_w30975_
	);
	LUT2 #(
		.INIT('h8)
	) name26929 (
		_w30969_,
		_w30975_,
		_w30976_
	);
	LUT2 #(
		.INIT('h4)
	) name26930 (
		_w30958_,
		_w30961_,
		_w30977_
	);
	LUT2 #(
		.INIT('h4)
	) name26931 (
		_w30966_,
		_w30977_,
		_w30978_
	);
	LUT2 #(
		.INIT('h8)
	) name26932 (
		_w30970_,
		_w30978_,
		_w30979_
	);
	LUT2 #(
		.INIT('h4)
	) name26933 (
		_w30944_,
		_w30966_,
		_w30980_
	);
	LUT2 #(
		.INIT('h8)
	) name26934 (
		_w30963_,
		_w30980_,
		_w30981_
	);
	LUT2 #(
		.INIT('h8)
	) name26935 (
		_w30974_,
		_w30978_,
		_w30982_
	);
	LUT2 #(
		.INIT('h1)
	) name26936 (
		_w30979_,
		_w30981_,
		_w30983_
	);
	LUT2 #(
		.INIT('h4)
	) name26937 (
		_w30982_,
		_w30983_,
		_w30984_
	);
	LUT2 #(
		.INIT('h1)
	) name26938 (
		_w30968_,
		_w30972_,
		_w30985_
	);
	LUT2 #(
		.INIT('h4)
	) name26939 (
		_w30976_,
		_w30985_,
		_w30986_
	);
	LUT2 #(
		.INIT('h8)
	) name26940 (
		_w30984_,
		_w30986_,
		_w30987_
	);
	LUT2 #(
		.INIT('h2)
	) name26941 (
		_w30934_,
		_w30987_,
		_w30988_
	);
	LUT2 #(
		.INIT('h1)
	) name26942 (
		_w30933_,
		_w30988_,
		_w30989_
	);
	LUT2 #(
		.INIT('h8)
	) name26943 (
		\core_c_dec_MFMAC_Ei_reg/NET0131 ,
		_w4117_,
		_w30990_
	);
	LUT2 #(
		.INIT('h2)
	) name26944 (
		_w25047_,
		_w30987_,
		_w30991_
	);
	LUT2 #(
		.INIT('h1)
	) name26945 (
		_w30990_,
		_w30991_,
		_w30992_
	);
	LUT2 #(
		.INIT('h8)
	) name26946 (
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w28786_,
		_w30993_
	);
	LUT2 #(
		.INIT('h1)
	) name26947 (
		\sport1_cfg_FSi_cnt_reg[11]/NET0131 ,
		_w28866_,
		_w30994_
	);
	LUT2 #(
		.INIT('h2)
	) name26948 (
		_w28855_,
		_w28867_,
		_w30995_
	);
	LUT2 #(
		.INIT('h4)
	) name26949 (
		_w30994_,
		_w30995_,
		_w30996_
	);
	LUT2 #(
		.INIT('h1)
	) name26950 (
		_w30993_,
		_w30996_,
		_w30997_
	);
	LUT2 #(
		.INIT('h8)
	) name26951 (
		\sport0_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w28876_,
		_w30998_
	);
	LUT2 #(
		.INIT('h1)
	) name26952 (
		\sport0_cfg_FSi_cnt_reg[11]/NET0131 ,
		_w28956_,
		_w30999_
	);
	LUT2 #(
		.INIT('h2)
	) name26953 (
		_w28945_,
		_w28957_,
		_w31000_
	);
	LUT2 #(
		.INIT('h4)
	) name26954 (
		_w30999_,
		_w31000_,
		_w31001_
	);
	LUT2 #(
		.INIT('h1)
	) name26955 (
		_w30998_,
		_w31001_,
		_w31002_
	);
	LUT2 #(
		.INIT('h8)
	) name26956 (
		\tm_tcr_reg_DO_reg[0]/NET0131 ,
		_w20355_,
		_w31003_
	);
	LUT2 #(
		.INIT('h4)
	) name26957 (
		\tm_tpr_reg_DO_reg[0]/NET0131 ,
		_w22400_,
		_w31004_
	);
	LUT2 #(
		.INIT('h2)
	) name26958 (
		\tm_TCR_TMP_reg[0]/NET0131 ,
		_w22411_,
		_w31005_
	);
	LUT2 #(
		.INIT('h1)
	) name26959 (
		_w22400_,
		_w30702_,
		_w31006_
	);
	LUT2 #(
		.INIT('h4)
	) name26960 (
		_w31005_,
		_w31006_,
		_w31007_
	);
	LUT2 #(
		.INIT('h1)
	) name26961 (
		_w20355_,
		_w31004_,
		_w31008_
	);
	LUT2 #(
		.INIT('h4)
	) name26962 (
		_w31007_,
		_w31008_,
		_w31009_
	);
	LUT2 #(
		.INIT('h1)
	) name26963 (
		_w31003_,
		_w31009_,
		_w31010_
	);
	LUT2 #(
		.INIT('h8)
	) name26964 (
		\tm_tcr_reg_DO_reg[3]/NET0131 ,
		_w20355_,
		_w31011_
	);
	LUT2 #(
		.INIT('h4)
	) name26965 (
		\tm_tpr_reg_DO_reg[3]/NET0131 ,
		_w22400_,
		_w31012_
	);
	LUT2 #(
		.INIT('h8)
	) name26966 (
		_w20359_,
		_w30702_,
		_w31013_
	);
	LUT2 #(
		.INIT('h2)
	) name26967 (
		\tm_TCR_TMP_reg[3]/NET0131 ,
		_w30712_,
		_w31014_
	);
	LUT2 #(
		.INIT('h1)
	) name26968 (
		_w22400_,
		_w31013_,
		_w31015_
	);
	LUT2 #(
		.INIT('h4)
	) name26969 (
		_w31014_,
		_w31015_,
		_w31016_
	);
	LUT2 #(
		.INIT('h1)
	) name26970 (
		_w20355_,
		_w31012_,
		_w31017_
	);
	LUT2 #(
		.INIT('h4)
	) name26971 (
		_w31016_,
		_w31017_,
		_w31018_
	);
	LUT2 #(
		.INIT('h1)
	) name26972 (
		_w31011_,
		_w31018_,
		_w31019_
	);
	LUT2 #(
		.INIT('h8)
	) name26973 (
		\tm_tcr_reg_DO_reg[4]/NET0131 ,
		_w20355_,
		_w31020_
	);
	LUT2 #(
		.INIT('h4)
	) name26974 (
		\tm_tpr_reg_DO_reg[4]/NET0131 ,
		_w22400_,
		_w31021_
	);
	LUT2 #(
		.INIT('h2)
	) name26975 (
		\tm_TCR_TMP_reg[4]/NET0131 ,
		_w22411_,
		_w31022_
	);
	LUT2 #(
		.INIT('h1)
	) name26976 (
		_w22400_,
		_w30734_,
		_w31023_
	);
	LUT2 #(
		.INIT('h4)
	) name26977 (
		_w31022_,
		_w31023_,
		_w31024_
	);
	LUT2 #(
		.INIT('h1)
	) name26978 (
		_w20355_,
		_w31021_,
		_w31025_
	);
	LUT2 #(
		.INIT('h4)
	) name26979 (
		_w31024_,
		_w31025_,
		_w31026_
	);
	LUT2 #(
		.INIT('h1)
	) name26980 (
		_w31020_,
		_w31026_,
		_w31027_
	);
	LUT2 #(
		.INIT('h8)
	) name26981 (
		\sport0_rxctl_RX_reg[12]/P0001 ,
		_w20871_,
		_w31028_
	);
	LUT2 #(
		.INIT('h1)
	) name26982 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		\sport0_rxctl_RX_reg[12]/P0001 ,
		_w31029_
	);
	LUT2 #(
		.INIT('h8)
	) name26983 (
		_w20957_,
		_w20976_,
		_w31030_
	);
	LUT2 #(
		.INIT('h4)
	) name26984 (
		_w20966_,
		_w20974_,
		_w31031_
	);
	LUT2 #(
		.INIT('h1)
	) name26985 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20914_,
		_w31032_
	);
	LUT2 #(
		.INIT('h2)
	) name26986 (
		_w20878_,
		_w31032_,
		_w31033_
	);
	LUT2 #(
		.INIT('h2)
	) name26987 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w31033_,
		_w31034_
	);
	LUT2 #(
		.INIT('h4)
	) name26988 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20884_,
		_w31035_
	);
	LUT2 #(
		.INIT('h1)
	) name26989 (
		_w20891_,
		_w31035_,
		_w31036_
	);
	LUT2 #(
		.INIT('h4)
	) name26990 (
		_w31034_,
		_w31036_,
		_w31037_
	);
	LUT2 #(
		.INIT('h8)
	) name26991 (
		_w20882_,
		_w31037_,
		_w31038_
	);
	LUT2 #(
		.INIT('h4)
	) name26992 (
		_w20882_,
		_w20966_,
		_w31039_
	);
	LUT2 #(
		.INIT('h4)
	) name26993 (
		_w20974_,
		_w31039_,
		_w31040_
	);
	LUT2 #(
		.INIT('h1)
	) name26994 (
		_w31031_,
		_w31038_,
		_w31041_
	);
	LUT2 #(
		.INIT('h4)
	) name26995 (
		_w31040_,
		_w31041_,
		_w31042_
	);
	LUT2 #(
		.INIT('h8)
	) name26996 (
		_w31030_,
		_w31042_,
		_w31043_
	);
	LUT2 #(
		.INIT('h1)
	) name26997 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w31043_,
		_w31044_
	);
	LUT2 #(
		.INIT('h4)
	) name26998 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20878_,
		_w31045_
	);
	LUT2 #(
		.INIT('h4)
	) name26999 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w31045_,
		_w31046_
	);
	LUT2 #(
		.INIT('h4)
	) name27000 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w31046_,
		_w31047_
	);
	LUT2 #(
		.INIT('h4)
	) name27001 (
		_w31044_,
		_w31047_,
		_w31048_
	);
	LUT2 #(
		.INIT('h1)
	) name27002 (
		_w31043_,
		_w31046_,
		_w31049_
	);
	LUT2 #(
		.INIT('h1)
	) name27003 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w31049_,
		_w31050_
	);
	LUT2 #(
		.INIT('h1)
	) name27004 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w31050_,
		_w31051_
	);
	LUT2 #(
		.INIT('h2)
	) name27005 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w31048_,
		_w31052_
	);
	LUT2 #(
		.INIT('h4)
	) name27006 (
		_w31051_,
		_w31052_,
		_w31053_
	);
	LUT2 #(
		.INIT('h2)
	) name27007 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w31029_,
		_w31054_
	);
	LUT2 #(
		.INIT('h4)
	) name27008 (
		_w31053_,
		_w31054_,
		_w31055_
	);
	LUT2 #(
		.INIT('h4)
	) name27009 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w20869_,
		_w31056_
	);
	LUT2 #(
		.INIT('h8)
	) name27010 (
		_w9178_,
		_w31056_,
		_w31057_
	);
	LUT2 #(
		.INIT('h1)
	) name27011 (
		_w31055_,
		_w31057_,
		_w31058_
	);
	LUT2 #(
		.INIT('h1)
	) name27012 (
		_w20868_,
		_w31058_,
		_w31059_
	);
	LUT2 #(
		.INIT('h8)
	) name27013 (
		\sport0_rxctl_RXSHT_reg[12]/P0001 ,
		_w20868_,
		_w31060_
	);
	LUT2 #(
		.INIT('h1)
	) name27014 (
		_w31028_,
		_w31060_,
		_w31061_
	);
	LUT2 #(
		.INIT('h4)
	) name27015 (
		_w31059_,
		_w31061_,
		_w31062_
	);
	LUT2 #(
		.INIT('h1)
	) name27016 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		\core_c_dec_updAR_E_reg/P0001 ,
		_w31063_
	);
	LUT2 #(
		.INIT('h2)
	) name27017 (
		_w14666_,
		_w31063_,
		_w31064_
	);
	LUT2 #(
		.INIT('h4)
	) name27018 (
		_w29291_,
		_w31064_,
		_w31065_
	);
	LUT2 #(
		.INIT('h2)
	) name27019 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[15]/P0001 ,
		_w31064_,
		_w31066_
	);
	LUT2 #(
		.INIT('h1)
	) name27020 (
		_w31065_,
		_w31066_,
		_w31067_
	);
	LUT2 #(
		.INIT('h4)
	) name27021 (
		\core_c_dec_MTMY1_E_reg/P0001 ,
		_w4117_,
		_w31068_
	);
	LUT2 #(
		.INIT('h1)
	) name27022 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		\core_c_dec_IR_reg[21]/NET0131 ,
		_w31069_
	);
	LUT2 #(
		.INIT('h2)
	) name27023 (
		\core_c_dec_IR_reg[22]/NET0131 ,
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w31070_
	);
	LUT2 #(
		.INIT('h4)
	) name27024 (
		_w31069_,
		_w31070_,
		_w31071_
	);
	LUT2 #(
		.INIT('h1)
	) name27025 (
		_w25244_,
		_w31071_,
		_w31072_
	);
	LUT2 #(
		.INIT('h4)
	) name27026 (
		_w25081_,
		_w31072_,
		_w31073_
	);
	LUT2 #(
		.INIT('h2)
	) name27027 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w31073_,
		_w31074_
	);
	LUT2 #(
		.INIT('h8)
	) name27028 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w31073_,
		_w31075_
	);
	LUT2 #(
		.INIT('h1)
	) name27029 (
		_w31074_,
		_w31075_,
		_w31076_
	);
	LUT2 #(
		.INIT('h2)
	) name27030 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w31073_,
		_w31077_
	);
	LUT2 #(
		.INIT('h8)
	) name27031 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w31073_,
		_w31078_
	);
	LUT2 #(
		.INIT('h1)
	) name27032 (
		_w31077_,
		_w31078_,
		_w31079_
	);
	LUT2 #(
		.INIT('h1)
	) name27033 (
		_w31076_,
		_w31079_,
		_w31080_
	);
	LUT2 #(
		.INIT('h1)
	) name27034 (
		_w25081_,
		_w30938_,
		_w31081_
	);
	LUT2 #(
		.INIT('h1)
	) name27035 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w31081_,
		_w31082_
	);
	LUT2 #(
		.INIT('h1)
	) name27036 (
		_w11745_,
		_w25244_,
		_w31083_
	);
	LUT2 #(
		.INIT('h1)
	) name27037 (
		_w18839_,
		_w24441_,
		_w31084_
	);
	LUT2 #(
		.INIT('h4)
	) name27038 (
		_w13578_,
		_w31084_,
		_w31085_
	);
	LUT2 #(
		.INIT('h4)
	) name27039 (
		_w11744_,
		_w31085_,
		_w31086_
	);
	LUT2 #(
		.INIT('h4)
	) name27040 (
		_w30945_,
		_w31083_,
		_w31087_
	);
	LUT2 #(
		.INIT('h8)
	) name27041 (
		_w31086_,
		_w31087_,
		_w31088_
	);
	LUT2 #(
		.INIT('h4)
	) name27042 (
		_w31082_,
		_w31088_,
		_w31089_
	);
	LUT2 #(
		.INIT('h8)
	) name27043 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w30935_,
		_w31090_
	);
	LUT2 #(
		.INIT('h8)
	) name27044 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w30935_,
		_w31091_
	);
	LUT2 #(
		.INIT('h1)
	) name27045 (
		_w25244_,
		_w30953_,
		_w31092_
	);
	LUT2 #(
		.INIT('h4)
	) name27046 (
		_w31090_,
		_w31092_,
		_w31093_
	);
	LUT2 #(
		.INIT('h4)
	) name27047 (
		_w31091_,
		_w31093_,
		_w31094_
	);
	LUT2 #(
		.INIT('h4)
	) name27048 (
		_w31089_,
		_w31094_,
		_w31095_
	);
	LUT2 #(
		.INIT('h2)
	) name27049 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w31073_,
		_w31096_
	);
	LUT2 #(
		.INIT('h8)
	) name27050 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w31073_,
		_w31097_
	);
	LUT2 #(
		.INIT('h1)
	) name27051 (
		_w31096_,
		_w31097_,
		_w31098_
	);
	LUT2 #(
		.INIT('h2)
	) name27052 (
		_w31095_,
		_w31098_,
		_w31099_
	);
	LUT2 #(
		.INIT('h2)
	) name27053 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w31073_,
		_w31100_
	);
	LUT2 #(
		.INIT('h8)
	) name27054 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w31073_,
		_w31101_
	);
	LUT2 #(
		.INIT('h1)
	) name27055 (
		_w31100_,
		_w31101_,
		_w31102_
	);
	LUT2 #(
		.INIT('h8)
	) name27056 (
		_w31099_,
		_w31102_,
		_w31103_
	);
	LUT2 #(
		.INIT('h8)
	) name27057 (
		_w31080_,
		_w31103_,
		_w31104_
	);
	LUT2 #(
		.INIT('h8)
	) name27058 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w6023_,
		_w31105_
	);
	LUT2 #(
		.INIT('h1)
	) name27059 (
		_w4117_,
		_w31105_,
		_w31106_
	);
	LUT2 #(
		.INIT('h4)
	) name27060 (
		_w31104_,
		_w31106_,
		_w31107_
	);
	LUT2 #(
		.INIT('h2)
	) name27061 (
		_w4116_,
		_w31068_,
		_w31108_
	);
	LUT2 #(
		.INIT('h4)
	) name27062 (
		_w31107_,
		_w31108_,
		_w31109_
	);
	LUT2 #(
		.INIT('h4)
	) name27063 (
		\core_c_dec_MTMY0_E_reg/P0001 ,
		_w4117_,
		_w31110_
	);
	LUT2 #(
		.INIT('h8)
	) name27064 (
		_w31095_,
		_w31098_,
		_w31111_
	);
	LUT2 #(
		.INIT('h8)
	) name27065 (
		_w31102_,
		_w31111_,
		_w31112_
	);
	LUT2 #(
		.INIT('h8)
	) name27066 (
		_w31080_,
		_w31112_,
		_w31113_
	);
	LUT2 #(
		.INIT('h4)
	) name27067 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w6023_,
		_w31114_
	);
	LUT2 #(
		.INIT('h1)
	) name27068 (
		_w4117_,
		_w31114_,
		_w31115_
	);
	LUT2 #(
		.INIT('h4)
	) name27069 (
		_w31113_,
		_w31115_,
		_w31116_
	);
	LUT2 #(
		.INIT('h2)
	) name27070 (
		_w4116_,
		_w31110_,
		_w31117_
	);
	LUT2 #(
		.INIT('h4)
	) name27071 (
		_w31116_,
		_w31117_,
		_w31118_
	);
	LUT2 #(
		.INIT('h8)
	) name27072 (
		\core_c_dec_MTAY1_E_reg/P0001 ,
		_w4117_,
		_w31119_
	);
	LUT2 #(
		.INIT('h4)
	) name27073 (
		_w4117_,
		_w31099_,
		_w31120_
	);
	LUT2 #(
		.INIT('h8)
	) name27074 (
		_w31076_,
		_w31102_,
		_w31121_
	);
	LUT2 #(
		.INIT('h4)
	) name27075 (
		_w31079_,
		_w31121_,
		_w31122_
	);
	LUT2 #(
		.INIT('h8)
	) name27076 (
		_w31120_,
		_w31122_,
		_w31123_
	);
	LUT2 #(
		.INIT('h1)
	) name27077 (
		_w31119_,
		_w31123_,
		_w31124_
	);
	LUT2 #(
		.INIT('h2)
	) name27078 (
		_w4116_,
		_w31124_,
		_w31125_
	);
	LUT2 #(
		.INIT('h8)
	) name27079 (
		\core_c_dec_MTAY0_E_reg/P0001 ,
		_w4117_,
		_w31126_
	);
	LUT2 #(
		.INIT('h4)
	) name27080 (
		_w4117_,
		_w31111_,
		_w31127_
	);
	LUT2 #(
		.INIT('h8)
	) name27081 (
		_w31122_,
		_w31127_,
		_w31128_
	);
	LUT2 #(
		.INIT('h1)
	) name27082 (
		_w31126_,
		_w31128_,
		_w31129_
	);
	LUT2 #(
		.INIT('h2)
	) name27083 (
		_w4116_,
		_w31129_,
		_w31130_
	);
	LUT2 #(
		.INIT('h1)
	) name27084 (
		\sport0_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		_w19548_,
		_w31131_
	);
	LUT2 #(
		.INIT('h2)
	) name27085 (
		_w19197_,
		_w19549_,
		_w31132_
	);
	LUT2 #(
		.INIT('h4)
	) name27086 (
		_w31131_,
		_w31132_,
		_w31133_
	);
	LUT2 #(
		.INIT('h2)
	) name27087 (
		_w13804_,
		_w31063_,
		_w31134_
	);
	LUT2 #(
		.INIT('h4)
	) name27088 (
		_w29291_,
		_w31134_,
		_w31135_
	);
	LUT2 #(
		.INIT('h2)
	) name27089 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[15]/P0001 ,
		_w31134_,
		_w31136_
	);
	LUT2 #(
		.INIT('h1)
	) name27090 (
		_w31135_,
		_w31136_,
		_w31137_
	);
	LUT2 #(
		.INIT('h2)
	) name27091 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 ,
		_w18266_,
		_w31138_
	);
	LUT2 #(
		.INIT('h1)
	) name27092 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[11]/P0001 ,
		_w18271_,
		_w31139_
	);
	LUT2 #(
		.INIT('h2)
	) name27093 (
		_w18271_,
		_w23757_,
		_w31140_
	);
	LUT2 #(
		.INIT('h2)
	) name27094 (
		_w18273_,
		_w31139_,
		_w31141_
	);
	LUT2 #(
		.INIT('h4)
	) name27095 (
		_w31140_,
		_w31141_,
		_w31142_
	);
	LUT2 #(
		.INIT('h1)
	) name27096 (
		_w18270_,
		_w31138_,
		_w31143_
	);
	LUT2 #(
		.INIT('h4)
	) name27097 (
		_w31142_,
		_w31143_,
		_w31144_
	);
	LUT2 #(
		.INIT('h1)
	) name27098 (
		_w18262_,
		_w31144_,
		_w31145_
	);
	LUT2 #(
		.INIT('h2)
	) name27099 (
		_w18262_,
		_w19618_,
		_w31146_
	);
	LUT2 #(
		.INIT('h1)
	) name27100 (
		_w31145_,
		_w31146_,
		_w31147_
	);
	LUT2 #(
		.INIT('h8)
	) name27101 (
		_w14752_,
		_w19618_,
		_w31148_
	);
	LUT2 #(
		.INIT('h8)
	) name27102 (
		_w18328_,
		_w23757_,
		_w31149_
	);
	LUT2 #(
		.INIT('h2)
	) name27103 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[11]/P0001 ,
		_w18330_,
		_w31150_
	);
	LUT2 #(
		.INIT('h2)
	) name27104 (
		_w18334_,
		_w31150_,
		_w31151_
	);
	LUT2 #(
		.INIT('h4)
	) name27105 (
		_w31149_,
		_w31151_,
		_w31152_
	);
	LUT2 #(
		.INIT('h1)
	) name27106 (
		_w31148_,
		_w31152_,
		_w31153_
	);
	LUT2 #(
		.INIT('h1)
	) name27107 (
		\sice_RCS_reg[1]/NET0131 ,
		\sice_RST_req_reg/NET0131 ,
		_w31154_
	);
	LUT2 #(
		.INIT('h1)
	) name27108 (
		\sice_RCS_reg[0]/NET0131 ,
		_w31154_,
		_w31155_
	);
	LUT2 #(
		.INIT('h8)
	) name27109 (
		IACKn_pad,
		\sice_RCS_reg[0]/NET0131 ,
		_w31156_
	);
	LUT2 #(
		.INIT('h4)
	) name27110 (
		\sice_RCS_reg[1]/NET0131 ,
		_w31156_,
		_w31157_
	);
	LUT2 #(
		.INIT('h1)
	) name27111 (
		_w31155_,
		_w31157_,
		_w31158_
	);
	LUT2 #(
		.INIT('h1)
	) name27112 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 ,
		_w19499_,
		_w31159_
	);
	LUT2 #(
		.INIT('h2)
	) name27113 (
		_w19499_,
		_w23757_,
		_w31160_
	);
	LUT2 #(
		.INIT('h2)
	) name27114 (
		_w19501_,
		_w31159_,
		_w31161_
	);
	LUT2 #(
		.INIT('h4)
	) name27115 (
		_w31160_,
		_w31161_,
		_w31162_
	);
	LUT2 #(
		.INIT('h2)
	) name27116 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[11]/P0001 ,
		_w19383_,
		_w31163_
	);
	LUT2 #(
		.INIT('h1)
	) name27117 (
		_w19508_,
		_w31163_,
		_w31164_
	);
	LUT2 #(
		.INIT('h4)
	) name27118 (
		_w31162_,
		_w31164_,
		_w31165_
	);
	LUT2 #(
		.INIT('h1)
	) name27119 (
		_w18262_,
		_w31165_,
		_w31166_
	);
	LUT2 #(
		.INIT('h2)
	) name27120 (
		_w18262_,
		_w19436_,
		_w31167_
	);
	LUT2 #(
		.INIT('h1)
	) name27121 (
		_w31166_,
		_w31167_,
		_w31168_
	);
	LUT2 #(
		.INIT('h2)
	) name27122 (
		\core_eu_ea_alu_ea_reg_ay0swe_DO_reg[0]/P0001 ,
		_w21990_,
		_w31169_
	);
	LUT2 #(
		.INIT('h1)
	) name27123 (
		_w13806_,
		_w24517_,
		_w31170_
	);
	LUT2 #(
		.INIT('h2)
	) name27124 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w14486_,
		_w31171_
	);
	LUT2 #(
		.INIT('h4)
	) name27125 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w19222_,
		_w31172_
	);
	LUT2 #(
		.INIT('h1)
	) name27126 (
		_w31171_,
		_w31172_,
		_w31173_
	);
	LUT2 #(
		.INIT('h2)
	) name27127 (
		_w13837_,
		_w31173_,
		_w31174_
	);
	LUT2 #(
		.INIT('h4)
	) name27128 (
		_w13837_,
		_w31173_,
		_w31175_
	);
	LUT2 #(
		.INIT('h1)
	) name27129 (
		_w31174_,
		_w31175_,
		_w31176_
	);
	LUT2 #(
		.INIT('h8)
	) name27130 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w31176_,
		_w31177_
	);
	LUT2 #(
		.INIT('h1)
	) name27131 (
		\core_c_dec_DIVS_E_reg/P0001 ,
		_w31176_,
		_w31178_
	);
	LUT2 #(
		.INIT('h2)
	) name27132 (
		_w13806_,
		_w31177_,
		_w31179_
	);
	LUT2 #(
		.INIT('h4)
	) name27133 (
		_w31178_,
		_w31179_,
		_w31180_
	);
	LUT2 #(
		.INIT('h1)
	) name27134 (
		_w31170_,
		_w31180_,
		_w31181_
	);
	LUT2 #(
		.INIT('h8)
	) name27135 (
		_w21990_,
		_w31181_,
		_w31182_
	);
	LUT2 #(
		.INIT('h1)
	) name27136 (
		_w31169_,
		_w31182_,
		_w31183_
	);
	LUT2 #(
		.INIT('h2)
	) name27137 (
		\core_eu_ea_alu_ea_reg_ay0rwe_DO_reg[0]/P0001 ,
		_w22158_,
		_w31184_
	);
	LUT2 #(
		.INIT('h8)
	) name27138 (
		_w22158_,
		_w31181_,
		_w31185_
	);
	LUT2 #(
		.INIT('h1)
	) name27139 (
		_w31184_,
		_w31185_,
		_w31186_
	);
	LUT2 #(
		.INIT('h1)
	) name27140 (
		\sport1_cfg_SCLKi_cnt_reg[11]/NET0131 ,
		_w20249_,
		_w31187_
	);
	LUT2 #(
		.INIT('h2)
	) name27141 (
		_w19130_,
		_w20250_,
		_w31188_
	);
	LUT2 #(
		.INIT('h4)
	) name27142 (
		_w31187_,
		_w31188_,
		_w31189_
	);
	LUT2 #(
		.INIT('h4)
	) name27143 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w19205_,
		_w31190_
	);
	LUT2 #(
		.INIT('h8)
	) name27144 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][0]/P0001 ,
		_w14713_,
		_w31191_
	);
	LUT2 #(
		.INIT('h8)
	) name27145 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][0]/P0001 ,
		_w14702_,
		_w31192_
	);
	LUT2 #(
		.INIT('h8)
	) name27146 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][0]/P0001 ,
		_w14708_,
		_w31193_
	);
	LUT2 #(
		.INIT('h8)
	) name27147 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001 ,
		_w14706_,
		_w31194_
	);
	LUT2 #(
		.INIT('h8)
	) name27148 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][0]/P0001 ,
		_w14704_,
		_w31195_
	);
	LUT2 #(
		.INIT('h8)
	) name27149 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001 ,
		_w14711_,
		_w31196_
	);
	LUT2 #(
		.INIT('h8)
	) name27150 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001 ,
		_w14699_,
		_w31197_
	);
	LUT2 #(
		.INIT('h1)
	) name27151 (
		_w31191_,
		_w31192_,
		_w31198_
	);
	LUT2 #(
		.INIT('h1)
	) name27152 (
		_w31193_,
		_w31194_,
		_w31199_
	);
	LUT2 #(
		.INIT('h1)
	) name27153 (
		_w31195_,
		_w31196_,
		_w31200_
	);
	LUT2 #(
		.INIT('h4)
	) name27154 (
		_w31197_,
		_w31200_,
		_w31201_
	);
	LUT2 #(
		.INIT('h8)
	) name27155 (
		_w31198_,
		_w31199_,
		_w31202_
	);
	LUT2 #(
		.INIT('h8)
	) name27156 (
		_w31201_,
		_w31202_,
		_w31203_
	);
	LUT2 #(
		.INIT('h2)
	) name27157 (
		_w14697_,
		_w31203_,
		_w31204_
	);
	LUT2 #(
		.INIT('h8)
	) name27158 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w7607_,
		_w31205_
	);
	LUT2 #(
		.INIT('h8)
	) name27159 (
		_w14564_,
		_w19206_,
		_w31206_
	);
	LUT2 #(
		.INIT('h4)
	) name27160 (
		_w14573_,
		_w31206_,
		_w31207_
	);
	LUT2 #(
		.INIT('h8)
	) name27161 (
		_w14586_,
		_w31207_,
		_w31208_
	);
	LUT2 #(
		.INIT('h8)
	) name27162 (
		_w14610_,
		_w31208_,
		_w31209_
	);
	LUT2 #(
		.INIT('h8)
	) name27163 (
		_w14600_,
		_w31209_,
		_w31210_
	);
	LUT2 #(
		.INIT('h8)
	) name27164 (
		_w14634_,
		_w31210_,
		_w31211_
	);
	LUT2 #(
		.INIT('h8)
	) name27165 (
		_w14623_,
		_w31211_,
		_w31212_
	);
	LUT2 #(
		.INIT('h8)
	) name27166 (
		_w23253_,
		_w31212_,
		_w31213_
	);
	LUT2 #(
		.INIT('h8)
	) name27167 (
		_w14658_,
		_w31213_,
		_w31214_
	);
	LUT2 #(
		.INIT('h8)
	) name27168 (
		_w14649_,
		_w31214_,
		_w31215_
	);
	LUT2 #(
		.INIT('h8)
	) name27169 (
		_w20053_,
		_w31215_,
		_w31216_
	);
	LUT2 #(
		.INIT('h8)
	) name27170 (
		_w14424_,
		_w31216_,
		_w31217_
	);
	LUT2 #(
		.INIT('h8)
	) name27171 (
		_w14413_,
		_w31217_,
		_w31218_
	);
	LUT2 #(
		.INIT('h8)
	) name27172 (
		_w14551_,
		_w31218_,
		_w31219_
	);
	LUT2 #(
		.INIT('h4)
	) name27173 (
		_w14540_,
		_w31219_,
		_w31220_
	);
	LUT2 #(
		.INIT('h8)
	) name27174 (
		_w19222_,
		_w31220_,
		_w31221_
	);
	LUT2 #(
		.INIT('h1)
	) name27175 (
		_w31204_,
		_w31205_,
		_w31222_
	);
	LUT2 #(
		.INIT('h4)
	) name27176 (
		_w19205_,
		_w31222_,
		_w31223_
	);
	LUT2 #(
		.INIT('h4)
	) name27177 (
		_w31221_,
		_w31223_,
		_w31224_
	);
	LUT2 #(
		.INIT('h2)
	) name27178 (
		_w4150_,
		_w31190_,
		_w31225_
	);
	LUT2 #(
		.INIT('h4)
	) name27179 (
		_w31224_,
		_w31225_,
		_w31226_
	);
	LUT2 #(
		.INIT('h8)
	) name27180 (
		_w14752_,
		_w19436_,
		_w31227_
	);
	LUT2 #(
		.INIT('h8)
	) name27181 (
		_w19776_,
		_w23757_,
		_w31228_
	);
	LUT2 #(
		.INIT('h2)
	) name27182 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[11]/P0001 ,
		_w17809_,
		_w31229_
	);
	LUT2 #(
		.INIT('h2)
	) name27183 (
		_w19780_,
		_w31229_,
		_w31230_
	);
	LUT2 #(
		.INIT('h4)
	) name27184 (
		_w31228_,
		_w31230_,
		_w31231_
	);
	LUT2 #(
		.INIT('h1)
	) name27185 (
		_w31227_,
		_w31231_,
		_w31232_
	);
	LUT2 #(
		.INIT('h4)
	) name27186 (
		_w5950_,
		_w13806_,
		_w31233_
	);
	LUT2 #(
		.INIT('h2)
	) name27187 (
		_w19202_,
		_w31233_,
		_w31234_
	);
	LUT2 #(
		.INIT('h4)
	) name27188 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w31234_,
		_w31235_
	);
	LUT2 #(
		.INIT('h8)
	) name27189 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w10911_,
		_w31236_
	);
	LUT2 #(
		.INIT('h8)
	) name27190 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][5]/P0001 ,
		_w14713_,
		_w31237_
	);
	LUT2 #(
		.INIT('h8)
	) name27191 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][5]/P0001 ,
		_w14702_,
		_w31238_
	);
	LUT2 #(
		.INIT('h8)
	) name27192 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001 ,
		_w14706_,
		_w31239_
	);
	LUT2 #(
		.INIT('h8)
	) name27193 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][5]/P0001 ,
		_w14708_,
		_w31240_
	);
	LUT2 #(
		.INIT('h8)
	) name27194 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001 ,
		_w14704_,
		_w31241_
	);
	LUT2 #(
		.INIT('h8)
	) name27195 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001 ,
		_w14699_,
		_w31242_
	);
	LUT2 #(
		.INIT('h8)
	) name27196 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001 ,
		_w14711_,
		_w31243_
	);
	LUT2 #(
		.INIT('h1)
	) name27197 (
		_w31237_,
		_w31238_,
		_w31244_
	);
	LUT2 #(
		.INIT('h1)
	) name27198 (
		_w31239_,
		_w31240_,
		_w31245_
	);
	LUT2 #(
		.INIT('h1)
	) name27199 (
		_w31241_,
		_w31242_,
		_w31246_
	);
	LUT2 #(
		.INIT('h4)
	) name27200 (
		_w31243_,
		_w31246_,
		_w31247_
	);
	LUT2 #(
		.INIT('h8)
	) name27201 (
		_w31244_,
		_w31245_,
		_w31248_
	);
	LUT2 #(
		.INIT('h8)
	) name27202 (
		_w31247_,
		_w31248_,
		_w31249_
	);
	LUT2 #(
		.INIT('h2)
	) name27203 (
		_w14697_,
		_w31249_,
		_w31250_
	);
	LUT2 #(
		.INIT('h8)
	) name27204 (
		_w13806_,
		_w31176_,
		_w31251_
	);
	LUT2 #(
		.INIT('h1)
	) name27205 (
		_w31236_,
		_w31250_,
		_w31252_
	);
	LUT2 #(
		.INIT('h4)
	) name27206 (
		_w31234_,
		_w31252_,
		_w31253_
	);
	LUT2 #(
		.INIT('h4)
	) name27207 (
		_w31251_,
		_w31253_,
		_w31254_
	);
	LUT2 #(
		.INIT('h2)
	) name27208 (
		_w4150_,
		_w31235_,
		_w31255_
	);
	LUT2 #(
		.INIT('h4)
	) name27209 (
		_w31254_,
		_w31255_,
		_w31256_
	);
	LUT2 #(
		.INIT('h8)
	) name27210 (
		\core_c_dec_pMFALU_Ei_reg/NET0131 ,
		_w4117_,
		_w31257_
	);
	LUT2 #(
		.INIT('h8)
	) name27211 (
		_w30955_,
		_w30961_,
		_w31258_
	);
	LUT2 #(
		.INIT('h8)
	) name27212 (
		_w30980_,
		_w31258_,
		_w31259_
	);
	LUT2 #(
		.INIT('h8)
	) name27213 (
		_w30967_,
		_w30973_,
		_w31260_
	);
	LUT2 #(
		.INIT('h8)
	) name27214 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w30935_,
		_w31261_
	);
	LUT2 #(
		.INIT('h2)
	) name27215 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		_w30935_,
		_w31262_
	);
	LUT2 #(
		.INIT('h1)
	) name27216 (
		_w31261_,
		_w31262_,
		_w31263_
	);
	LUT2 #(
		.INIT('h1)
	) name27217 (
		_w30936_,
		_w31263_,
		_w31264_
	);
	LUT2 #(
		.INIT('h1)
	) name27218 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w31265_
	);
	LUT2 #(
		.INIT('h8)
	) name27219 (
		_w31264_,
		_w31265_,
		_w31266_
	);
	LUT2 #(
		.INIT('h8)
	) name27220 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w30935_,
		_w31267_
	);
	LUT2 #(
		.INIT('h2)
	) name27221 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w30935_,
		_w31268_
	);
	LUT2 #(
		.INIT('h1)
	) name27222 (
		_w31267_,
		_w31268_,
		_w31269_
	);
	LUT2 #(
		.INIT('h1)
	) name27223 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w31269_,
		_w31270_
	);
	LUT2 #(
		.INIT('h4)
	) name27224 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w31270_,
		_w31271_
	);
	LUT2 #(
		.INIT('h8)
	) name27225 (
		_w31266_,
		_w31271_,
		_w31272_
	);
	LUT2 #(
		.INIT('h1)
	) name27226 (
		_w31259_,
		_w31272_,
		_w31273_
	);
	LUT2 #(
		.INIT('h4)
	) name27227 (
		_w31260_,
		_w31273_,
		_w31274_
	);
	LUT2 #(
		.INIT('h2)
	) name27228 (
		_w30934_,
		_w31274_,
		_w31275_
	);
	LUT2 #(
		.INIT('h1)
	) name27229 (
		_w31257_,
		_w31275_,
		_w31276_
	);
	LUT2 #(
		.INIT('h8)
	) name27230 (
		\core_c_dec_MFALU_Ei_reg/NET0131 ,
		_w4117_,
		_w31277_
	);
	LUT2 #(
		.INIT('h2)
	) name27231 (
		_w25047_,
		_w31274_,
		_w31278_
	);
	LUT2 #(
		.INIT('h1)
	) name27232 (
		_w31277_,
		_w31278_,
		_w31279_
	);
	LUT2 #(
		.INIT('h2)
	) name27233 (
		\sport1_txctl_TXSHT_reg[6]/P0001 ,
		_w22677_,
		_w31280_
	);
	LUT2 #(
		.INIT('h8)
	) name27234 (
		\sport1_txctl_TX_reg[7]/P0001 ,
		_w22677_,
		_w31281_
	);
	LUT2 #(
		.INIT('h1)
	) name27235 (
		_w31280_,
		_w31281_,
		_w31282_
	);
	LUT2 #(
		.INIT('h8)
	) name27236 (
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w28786_,
		_w31283_
	);
	LUT2 #(
		.INIT('h1)
	) name27237 (
		\sport1_cfg_FSi_cnt_reg[10]/NET0131 ,
		_w28865_,
		_w31284_
	);
	LUT2 #(
		.INIT('h2)
	) name27238 (
		_w28855_,
		_w28866_,
		_w31285_
	);
	LUT2 #(
		.INIT('h4)
	) name27239 (
		_w31284_,
		_w31285_,
		_w31286_
	);
	LUT2 #(
		.INIT('h1)
	) name27240 (
		_w31283_,
		_w31286_,
		_w31287_
	);
	LUT2 #(
		.INIT('h8)
	) name27241 (
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w28786_,
		_w31288_
	);
	LUT2 #(
		.INIT('h1)
	) name27242 (
		\sport1_cfg_FSi_cnt_reg[12]/NET0131 ,
		_w28867_,
		_w31289_
	);
	LUT2 #(
		.INIT('h2)
	) name27243 (
		_w28855_,
		_w28868_,
		_w31290_
	);
	LUT2 #(
		.INIT('h4)
	) name27244 (
		_w31289_,
		_w31290_,
		_w31291_
	);
	LUT2 #(
		.INIT('h1)
	) name27245 (
		_w31288_,
		_w31291_,
		_w31292_
	);
	LUT2 #(
		.INIT('h8)
	) name27246 (
		\sport0_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w28876_,
		_w31293_
	);
	LUT2 #(
		.INIT('h1)
	) name27247 (
		\sport0_cfg_FSi_cnt_reg[10]/NET0131 ,
		_w28955_,
		_w31294_
	);
	LUT2 #(
		.INIT('h2)
	) name27248 (
		_w28945_,
		_w28956_,
		_w31295_
	);
	LUT2 #(
		.INIT('h4)
	) name27249 (
		_w31294_,
		_w31295_,
		_w31296_
	);
	LUT2 #(
		.INIT('h1)
	) name27250 (
		_w31293_,
		_w31296_,
		_w31297_
	);
	LUT2 #(
		.INIT('h2)
	) name27251 (
		\sport0_txctl_TXSHT_reg[6]/P0001 ,
		_w19960_,
		_w31298_
	);
	LUT2 #(
		.INIT('h8)
	) name27252 (
		\sport0_txctl_TX_reg[7]/P0001 ,
		_w19960_,
		_w31299_
	);
	LUT2 #(
		.INIT('h1)
	) name27253 (
		_w31298_,
		_w31299_,
		_w31300_
	);
	LUT2 #(
		.INIT('h8)
	) name27254 (
		\sport0_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w28876_,
		_w31301_
	);
	LUT2 #(
		.INIT('h1)
	) name27255 (
		\sport0_cfg_FSi_cnt_reg[12]/NET0131 ,
		_w28957_,
		_w31302_
	);
	LUT2 #(
		.INIT('h2)
	) name27256 (
		_w28945_,
		_w28958_,
		_w31303_
	);
	LUT2 #(
		.INIT('h4)
	) name27257 (
		_w31302_,
		_w31303_,
		_w31304_
	);
	LUT2 #(
		.INIT('h1)
	) name27258 (
		_w31301_,
		_w31304_,
		_w31305_
	);
	LUT2 #(
		.INIT('h2)
	) name27259 (
		\core_dag_ilm2reg_M_E_reg[1]/NET0131 ,
		_w5692_,
		_w31306_
	);
	LUT2 #(
		.INIT('h2)
	) name27260 (
		_w4055_,
		_w25690_,
		_w31307_
	);
	LUT2 #(
		.INIT('h8)
	) name27261 (
		\sport0_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w5970_,
		_w31308_
	);
	LUT2 #(
		.INIT('h8)
	) name27262 (
		\sport1_regs_AUTOreg_DO_reg[3]/NET0131 ,
		_w5966_,
		_w31309_
	);
	LUT2 #(
		.INIT('h8)
	) name27263 (
		\sport1_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w5968_,
		_w31310_
	);
	LUT2 #(
		.INIT('h8)
	) name27264 (
		\sport0_regs_AUTOreg_DO_reg[8]/NET0131 ,
		_w4050_,
		_w31311_
	);
	LUT2 #(
		.INIT('h1)
	) name27265 (
		_w31308_,
		_w31311_,
		_w31312_
	);
	LUT2 #(
		.INIT('h4)
	) name27266 (
		_w31310_,
		_w31312_,
		_w31313_
	);
	LUT2 #(
		.INIT('h4)
	) name27267 (
		_w31309_,
		_w31313_,
		_w31314_
	);
	LUT2 #(
		.INIT('h4)
	) name27268 (
		_w31307_,
		_w31314_,
		_w31315_
	);
	LUT2 #(
		.INIT('h2)
	) name27269 (
		_w5692_,
		_w31315_,
		_w31316_
	);
	LUT2 #(
		.INIT('h1)
	) name27270 (
		_w31306_,
		_w31316_,
		_w31317_
	);
	LUT2 #(
		.INIT('h2)
	) name27271 (
		\core_dag_ilm2reg_M_E_reg[0]/NET0131 ,
		_w5692_,
		_w31318_
	);
	LUT2 #(
		.INIT('h2)
	) name27272 (
		_w4055_,
		_w25696_,
		_w31319_
	);
	LUT2 #(
		.INIT('h8)
	) name27273 (
		\sport0_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w4050_,
		_w31320_
	);
	LUT2 #(
		.INIT('h8)
	) name27274 (
		\sport1_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w5966_,
		_w31321_
	);
	LUT2 #(
		.INIT('h8)
	) name27275 (
		\sport1_regs_AUTOreg_DO_reg[7]/NET0131 ,
		_w5968_,
		_w31322_
	);
	LUT2 #(
		.INIT('h8)
	) name27276 (
		\sport0_regs_AUTOreg_DO_reg[2]/NET0131 ,
		_w5970_,
		_w31323_
	);
	LUT2 #(
		.INIT('h1)
	) name27277 (
		_w31320_,
		_w31323_,
		_w31324_
	);
	LUT2 #(
		.INIT('h4)
	) name27278 (
		_w31322_,
		_w31324_,
		_w31325_
	);
	LUT2 #(
		.INIT('h4)
	) name27279 (
		_w31321_,
		_w31325_,
		_w31326_
	);
	LUT2 #(
		.INIT('h4)
	) name27280 (
		_w31319_,
		_w31326_,
		_w31327_
	);
	LUT2 #(
		.INIT('h2)
	) name27281 (
		_w5692_,
		_w31327_,
		_w31328_
	);
	LUT2 #(
		.INIT('h1)
	) name27282 (
		_w31318_,
		_w31328_,
		_w31329_
	);
	LUT2 #(
		.INIT('h4)
	) name27283 (
		_w31317_,
		_w31329_,
		_w31330_
	);
	LUT2 #(
		.INIT('h4)
	) name27284 (
		_w26059_,
		_w31330_,
		_w31331_
	);
	LUT2 #(
		.INIT('h1)
	) name27285 (
		_w26060_,
		_w31329_,
		_w31332_
	);
	LUT2 #(
		.INIT('h4)
	) name27286 (
		_w26075_,
		_w31329_,
		_w31333_
	);
	LUT2 #(
		.INIT('h1)
	) name27287 (
		_w31332_,
		_w31333_,
		_w31334_
	);
	LUT2 #(
		.INIT('h2)
	) name27288 (
		_w31317_,
		_w31334_,
		_w31335_
	);
	LUT2 #(
		.INIT('h1)
	) name27289 (
		_w31317_,
		_w31329_,
		_w31336_
	);
	LUT2 #(
		.INIT('h4)
	) name27290 (
		_w26074_,
		_w31336_,
		_w31337_
	);
	LUT2 #(
		.INIT('h1)
	) name27291 (
		_w31331_,
		_w31337_,
		_w31338_
	);
	LUT2 #(
		.INIT('h4)
	) name27292 (
		_w31335_,
		_w31338_,
		_w31339_
	);
	LUT2 #(
		.INIT('h8)
	) name27293 (
		_w10289_,
		_w31339_,
		_w31340_
	);
	LUT2 #(
		.INIT('h8)
	) name27294 (
		_w31317_,
		_w31332_,
		_w31341_
	);
	LUT2 #(
		.INIT('h8)
	) name27295 (
		\core_dag_ilm2reg_M5_we_DO_reg[9]/NET0131 ,
		_w31341_,
		_w31342_
	);
	LUT2 #(
		.INIT('h8)
	) name27296 (
		\core_dag_ilm2reg_M7_we_DO_reg[9]/NET0131 ,
		_w31337_,
		_w31343_
	);
	LUT2 #(
		.INIT('h8)
	) name27297 (
		_w31317_,
		_w31333_,
		_w31344_
	);
	LUT2 #(
		.INIT('h8)
	) name27298 (
		\core_dag_ilm2reg_M4_we_DO_reg[9]/NET0131 ,
		_w31344_,
		_w31345_
	);
	LUT2 #(
		.INIT('h8)
	) name27299 (
		\core_dag_ilm2reg_M6_we_DO_reg[9]/NET0131 ,
		_w31331_,
		_w31346_
	);
	LUT2 #(
		.INIT('h1)
	) name27300 (
		_w31343_,
		_w31346_,
		_w31347_
	);
	LUT2 #(
		.INIT('h4)
	) name27301 (
		_w21579_,
		_w31347_,
		_w31348_
	);
	LUT2 #(
		.INIT('h1)
	) name27302 (
		_w31342_,
		_w31345_,
		_w31349_
	);
	LUT2 #(
		.INIT('h8)
	) name27303 (
		_w31348_,
		_w31349_,
		_w31350_
	);
	LUT2 #(
		.INIT('h4)
	) name27304 (
		_w31340_,
		_w31350_,
		_w31351_
	);
	LUT2 #(
		.INIT('h4)
	) name27305 (
		\core_dag_ilm2reg_M_reg[9]/NET0131 ,
		_w21579_,
		_w31352_
	);
	LUT2 #(
		.INIT('h1)
	) name27306 (
		_w31351_,
		_w31352_,
		_w31353_
	);
	LUT2 #(
		.INIT('h8)
	) name27307 (
		_w9178_,
		_w31339_,
		_w31354_
	);
	LUT2 #(
		.INIT('h8)
	) name27308 (
		\core_dag_ilm2reg_M5_we_DO_reg[12]/NET0131 ,
		_w31341_,
		_w31355_
	);
	LUT2 #(
		.INIT('h8)
	) name27309 (
		\core_dag_ilm2reg_M7_we_DO_reg[12]/NET0131 ,
		_w31337_,
		_w31356_
	);
	LUT2 #(
		.INIT('h8)
	) name27310 (
		\core_dag_ilm2reg_M4_we_DO_reg[12]/NET0131 ,
		_w31344_,
		_w31357_
	);
	LUT2 #(
		.INIT('h8)
	) name27311 (
		\core_dag_ilm2reg_M6_we_DO_reg[12]/NET0131 ,
		_w31331_,
		_w31358_
	);
	LUT2 #(
		.INIT('h1)
	) name27312 (
		_w31356_,
		_w31358_,
		_w31359_
	);
	LUT2 #(
		.INIT('h4)
	) name27313 (
		_w21579_,
		_w31359_,
		_w31360_
	);
	LUT2 #(
		.INIT('h1)
	) name27314 (
		_w31355_,
		_w31357_,
		_w31361_
	);
	LUT2 #(
		.INIT('h8)
	) name27315 (
		_w31360_,
		_w31361_,
		_w31362_
	);
	LUT2 #(
		.INIT('h4)
	) name27316 (
		_w31354_,
		_w31362_,
		_w31363_
	);
	LUT2 #(
		.INIT('h4)
	) name27317 (
		\core_dag_ilm2reg_M_reg[12]/NET0131 ,
		_w21579_,
		_w31364_
	);
	LUT2 #(
		.INIT('h1)
	) name27318 (
		_w31363_,
		_w31364_,
		_w31365_
	);
	LUT2 #(
		.INIT('h8)
	) name27319 (
		_w8460_,
		_w31339_,
		_w31366_
	);
	LUT2 #(
		.INIT('h8)
	) name27320 (
		\core_dag_ilm2reg_M5_we_DO_reg[11]/NET0131 ,
		_w31341_,
		_w31367_
	);
	LUT2 #(
		.INIT('h8)
	) name27321 (
		\core_dag_ilm2reg_M7_we_DO_reg[11]/NET0131 ,
		_w31337_,
		_w31368_
	);
	LUT2 #(
		.INIT('h8)
	) name27322 (
		\core_dag_ilm2reg_M4_we_DO_reg[11]/NET0131 ,
		_w31344_,
		_w31369_
	);
	LUT2 #(
		.INIT('h8)
	) name27323 (
		\core_dag_ilm2reg_M6_we_DO_reg[11]/NET0131 ,
		_w31331_,
		_w31370_
	);
	LUT2 #(
		.INIT('h1)
	) name27324 (
		_w31368_,
		_w31370_,
		_w31371_
	);
	LUT2 #(
		.INIT('h4)
	) name27325 (
		_w21579_,
		_w31371_,
		_w31372_
	);
	LUT2 #(
		.INIT('h1)
	) name27326 (
		_w31367_,
		_w31369_,
		_w31373_
	);
	LUT2 #(
		.INIT('h8)
	) name27327 (
		_w31372_,
		_w31373_,
		_w31374_
	);
	LUT2 #(
		.INIT('h4)
	) name27328 (
		_w31366_,
		_w31374_,
		_w31375_
	);
	LUT2 #(
		.INIT('h4)
	) name27329 (
		\core_dag_ilm2reg_M_reg[11]/NET0131 ,
		_w21579_,
		_w31376_
	);
	LUT2 #(
		.INIT('h1)
	) name27330 (
		_w31375_,
		_w31376_,
		_w31377_
	);
	LUT2 #(
		.INIT('h8)
	) name27331 (
		_w7859_,
		_w31339_,
		_w31378_
	);
	LUT2 #(
		.INIT('h8)
	) name27332 (
		\core_dag_ilm2reg_M5_we_DO_reg[10]/NET0131 ,
		_w31341_,
		_w31379_
	);
	LUT2 #(
		.INIT('h8)
	) name27333 (
		\core_dag_ilm2reg_M7_we_DO_reg[10]/NET0131 ,
		_w31337_,
		_w31380_
	);
	LUT2 #(
		.INIT('h8)
	) name27334 (
		\core_dag_ilm2reg_M4_we_DO_reg[10]/NET0131 ,
		_w31344_,
		_w31381_
	);
	LUT2 #(
		.INIT('h8)
	) name27335 (
		\core_dag_ilm2reg_M6_we_DO_reg[10]/NET0131 ,
		_w31331_,
		_w31382_
	);
	LUT2 #(
		.INIT('h1)
	) name27336 (
		_w31380_,
		_w31382_,
		_w31383_
	);
	LUT2 #(
		.INIT('h4)
	) name27337 (
		_w21579_,
		_w31383_,
		_w31384_
	);
	LUT2 #(
		.INIT('h1)
	) name27338 (
		_w31379_,
		_w31381_,
		_w31385_
	);
	LUT2 #(
		.INIT('h8)
	) name27339 (
		_w31384_,
		_w31385_,
		_w31386_
	);
	LUT2 #(
		.INIT('h4)
	) name27340 (
		_w31378_,
		_w31386_,
		_w31387_
	);
	LUT2 #(
		.INIT('h4)
	) name27341 (
		\core_dag_ilm2reg_M_reg[10]/NET0131 ,
		_w21579_,
		_w31388_
	);
	LUT2 #(
		.INIT('h1)
	) name27342 (
		_w31387_,
		_w31388_,
		_w31389_
	);
	LUT2 #(
		.INIT('h2)
	) name27343 (
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w5692_,
		_w31390_
	);
	LUT2 #(
		.INIT('h8)
	) name27344 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w4055_,
		_w31391_
	);
	LUT2 #(
		.INIT('h2)
	) name27345 (
		_w31314_,
		_w31391_,
		_w31392_
	);
	LUT2 #(
		.INIT('h2)
	) name27346 (
		_w5692_,
		_w31392_,
		_w31393_
	);
	LUT2 #(
		.INIT('h1)
	) name27347 (
		_w31390_,
		_w31393_,
		_w31394_
	);
	LUT2 #(
		.INIT('h2)
	) name27348 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		_w5692_,
		_w31395_
	);
	LUT2 #(
		.INIT('h8)
	) name27349 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w4055_,
		_w31396_
	);
	LUT2 #(
		.INIT('h2)
	) name27350 (
		_w31326_,
		_w31396_,
		_w31397_
	);
	LUT2 #(
		.INIT('h2)
	) name27351 (
		_w5692_,
		_w31397_,
		_w31398_
	);
	LUT2 #(
		.INIT('h1)
	) name27352 (
		_w31395_,
		_w31398_,
		_w31399_
	);
	LUT2 #(
		.INIT('h4)
	) name27353 (
		_w31394_,
		_w31399_,
		_w31400_
	);
	LUT2 #(
		.INIT('h4)
	) name27354 (
		_w26079_,
		_w31400_,
		_w31401_
	);
	LUT2 #(
		.INIT('h4)
	) name27355 (
		_w26080_,
		_w31399_,
		_w31402_
	);
	LUT2 #(
		.INIT('h1)
	) name27356 (
		_w26076_,
		_w31399_,
		_w31403_
	);
	LUT2 #(
		.INIT('h1)
	) name27357 (
		_w31402_,
		_w31403_,
		_w31404_
	);
	LUT2 #(
		.INIT('h2)
	) name27358 (
		_w31394_,
		_w31404_,
		_w31405_
	);
	LUT2 #(
		.INIT('h1)
	) name27359 (
		_w31394_,
		_w31399_,
		_w31406_
	);
	LUT2 #(
		.INIT('h4)
	) name27360 (
		_w26077_,
		_w31406_,
		_w31407_
	);
	LUT2 #(
		.INIT('h1)
	) name27361 (
		_w31401_,
		_w31407_,
		_w31408_
	);
	LUT2 #(
		.INIT('h4)
	) name27362 (
		_w31405_,
		_w31408_,
		_w31409_
	);
	LUT2 #(
		.INIT('h8)
	) name27363 (
		_w10289_,
		_w31409_,
		_w31410_
	);
	LUT2 #(
		.INIT('h8)
	) name27364 (
		_w31394_,
		_w31402_,
		_w31411_
	);
	LUT2 #(
		.INIT('h8)
	) name27365 (
		\core_dag_ilm1reg_M0_we_DO_reg[9]/NET0131 ,
		_w31411_,
		_w31412_
	);
	LUT2 #(
		.INIT('h8)
	) name27366 (
		\core_dag_ilm1reg_M3_we_DO_reg[9]/NET0131 ,
		_w31407_,
		_w31413_
	);
	LUT2 #(
		.INIT('h8)
	) name27367 (
		_w31394_,
		_w31403_,
		_w31414_
	);
	LUT2 #(
		.INIT('h8)
	) name27368 (
		\core_dag_ilm1reg_M1_we_DO_reg[9]/NET0131 ,
		_w31414_,
		_w31415_
	);
	LUT2 #(
		.INIT('h8)
	) name27369 (
		\core_dag_ilm1reg_M2_we_DO_reg[9]/NET0131 ,
		_w31401_,
		_w31416_
	);
	LUT2 #(
		.INIT('h1)
	) name27370 (
		_w31413_,
		_w31416_,
		_w31417_
	);
	LUT2 #(
		.INIT('h4)
	) name27371 (
		_w21592_,
		_w31417_,
		_w31418_
	);
	LUT2 #(
		.INIT('h1)
	) name27372 (
		_w31412_,
		_w31415_,
		_w31419_
	);
	LUT2 #(
		.INIT('h8)
	) name27373 (
		_w31418_,
		_w31419_,
		_w31420_
	);
	LUT2 #(
		.INIT('h4)
	) name27374 (
		_w31410_,
		_w31420_,
		_w31421_
	);
	LUT2 #(
		.INIT('h4)
	) name27375 (
		\core_dag_ilm1reg_M_reg[9]/NET0131 ,
		_w21592_,
		_w31422_
	);
	LUT2 #(
		.INIT('h1)
	) name27376 (
		_w31421_,
		_w31422_,
		_w31423_
	);
	LUT2 #(
		.INIT('h8)
	) name27377 (
		_w10638_,
		_w31409_,
		_w31424_
	);
	LUT2 #(
		.INIT('h8)
	) name27378 (
		\core_dag_ilm1reg_M0_we_DO_reg[8]/NET0131 ,
		_w31411_,
		_w31425_
	);
	LUT2 #(
		.INIT('h8)
	) name27379 (
		\core_dag_ilm1reg_M3_we_DO_reg[8]/NET0131 ,
		_w31407_,
		_w31426_
	);
	LUT2 #(
		.INIT('h8)
	) name27380 (
		\core_dag_ilm1reg_M1_we_DO_reg[8]/NET0131 ,
		_w31414_,
		_w31427_
	);
	LUT2 #(
		.INIT('h8)
	) name27381 (
		\core_dag_ilm1reg_M2_we_DO_reg[8]/NET0131 ,
		_w31401_,
		_w31428_
	);
	LUT2 #(
		.INIT('h1)
	) name27382 (
		_w31426_,
		_w31428_,
		_w31429_
	);
	LUT2 #(
		.INIT('h4)
	) name27383 (
		_w21592_,
		_w31429_,
		_w31430_
	);
	LUT2 #(
		.INIT('h1)
	) name27384 (
		_w31425_,
		_w31427_,
		_w31431_
	);
	LUT2 #(
		.INIT('h8)
	) name27385 (
		_w31430_,
		_w31431_,
		_w31432_
	);
	LUT2 #(
		.INIT('h4)
	) name27386 (
		_w31424_,
		_w31432_,
		_w31433_
	);
	LUT2 #(
		.INIT('h4)
	) name27387 (
		\core_dag_ilm1reg_M_reg[8]/NET0131 ,
		_w21592_,
		_w31434_
	);
	LUT2 #(
		.INIT('h1)
	) name27388 (
		_w31433_,
		_w31434_,
		_w31435_
	);
	LUT2 #(
		.INIT('h8)
	) name27389 (
		_w7340_,
		_w31409_,
		_w31436_
	);
	LUT2 #(
		.INIT('h8)
	) name27390 (
		\core_dag_ilm1reg_M0_we_DO_reg[13]/NET0131 ,
		_w31411_,
		_w31437_
	);
	LUT2 #(
		.INIT('h8)
	) name27391 (
		\core_dag_ilm1reg_M3_we_DO_reg[13]/NET0131 ,
		_w31407_,
		_w31438_
	);
	LUT2 #(
		.INIT('h8)
	) name27392 (
		\core_dag_ilm1reg_M1_we_DO_reg[13]/NET0131 ,
		_w31414_,
		_w31439_
	);
	LUT2 #(
		.INIT('h8)
	) name27393 (
		\core_dag_ilm1reg_M2_we_DO_reg[13]/NET0131 ,
		_w31401_,
		_w31440_
	);
	LUT2 #(
		.INIT('h1)
	) name27394 (
		_w31438_,
		_w31440_,
		_w31441_
	);
	LUT2 #(
		.INIT('h4)
	) name27395 (
		_w21592_,
		_w31441_,
		_w31442_
	);
	LUT2 #(
		.INIT('h1)
	) name27396 (
		_w31437_,
		_w31439_,
		_w31443_
	);
	LUT2 #(
		.INIT('h8)
	) name27397 (
		_w31442_,
		_w31443_,
		_w31444_
	);
	LUT2 #(
		.INIT('h4)
	) name27398 (
		_w31436_,
		_w31444_,
		_w31445_
	);
	LUT2 #(
		.INIT('h4)
	) name27399 (
		\core_dag_ilm1reg_M_reg[13]/NET0131 ,
		_w21592_,
		_w31446_
	);
	LUT2 #(
		.INIT('h1)
	) name27400 (
		_w31445_,
		_w31446_,
		_w31447_
	);
	LUT2 #(
		.INIT('h8)
	) name27401 (
		_w8460_,
		_w31409_,
		_w31448_
	);
	LUT2 #(
		.INIT('h8)
	) name27402 (
		\core_dag_ilm1reg_M0_we_DO_reg[11]/NET0131 ,
		_w31411_,
		_w31449_
	);
	LUT2 #(
		.INIT('h8)
	) name27403 (
		\core_dag_ilm1reg_M3_we_DO_reg[11]/NET0131 ,
		_w31407_,
		_w31450_
	);
	LUT2 #(
		.INIT('h8)
	) name27404 (
		\core_dag_ilm1reg_M1_we_DO_reg[11]/NET0131 ,
		_w31414_,
		_w31451_
	);
	LUT2 #(
		.INIT('h8)
	) name27405 (
		\core_dag_ilm1reg_M2_we_DO_reg[11]/NET0131 ,
		_w31401_,
		_w31452_
	);
	LUT2 #(
		.INIT('h1)
	) name27406 (
		_w31450_,
		_w31452_,
		_w31453_
	);
	LUT2 #(
		.INIT('h4)
	) name27407 (
		_w21592_,
		_w31453_,
		_w31454_
	);
	LUT2 #(
		.INIT('h1)
	) name27408 (
		_w31449_,
		_w31451_,
		_w31455_
	);
	LUT2 #(
		.INIT('h8)
	) name27409 (
		_w31454_,
		_w31455_,
		_w31456_
	);
	LUT2 #(
		.INIT('h4)
	) name27410 (
		_w31448_,
		_w31456_,
		_w31457_
	);
	LUT2 #(
		.INIT('h4)
	) name27411 (
		\core_dag_ilm1reg_M_reg[11]/NET0131 ,
		_w21592_,
		_w31458_
	);
	LUT2 #(
		.INIT('h1)
	) name27412 (
		_w31457_,
		_w31458_,
		_w31459_
	);
	LUT2 #(
		.INIT('h8)
	) name27413 (
		_w7859_,
		_w31409_,
		_w31460_
	);
	LUT2 #(
		.INIT('h8)
	) name27414 (
		\core_dag_ilm1reg_M0_we_DO_reg[10]/NET0131 ,
		_w31411_,
		_w31461_
	);
	LUT2 #(
		.INIT('h8)
	) name27415 (
		\core_dag_ilm1reg_M3_we_DO_reg[10]/NET0131 ,
		_w31407_,
		_w31462_
	);
	LUT2 #(
		.INIT('h8)
	) name27416 (
		\core_dag_ilm1reg_M1_we_DO_reg[10]/NET0131 ,
		_w31414_,
		_w31463_
	);
	LUT2 #(
		.INIT('h8)
	) name27417 (
		\core_dag_ilm1reg_M2_we_DO_reg[10]/NET0131 ,
		_w31401_,
		_w31464_
	);
	LUT2 #(
		.INIT('h1)
	) name27418 (
		_w31462_,
		_w31464_,
		_w31465_
	);
	LUT2 #(
		.INIT('h4)
	) name27419 (
		_w21592_,
		_w31465_,
		_w31466_
	);
	LUT2 #(
		.INIT('h1)
	) name27420 (
		_w31461_,
		_w31463_,
		_w31467_
	);
	LUT2 #(
		.INIT('h8)
	) name27421 (
		_w31466_,
		_w31467_,
		_w31468_
	);
	LUT2 #(
		.INIT('h4)
	) name27422 (
		_w31460_,
		_w31468_,
		_w31469_
	);
	LUT2 #(
		.INIT('h4)
	) name27423 (
		\core_dag_ilm1reg_M_reg[10]/NET0131 ,
		_w21592_,
		_w31470_
	);
	LUT2 #(
		.INIT('h1)
	) name27424 (
		_w31469_,
		_w31470_,
		_w31471_
	);
	LUT2 #(
		.INIT('h1)
	) name27425 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 ,
		_w19499_,
		_w31472_
	);
	LUT2 #(
		.INIT('h2)
	) name27426 (
		_w19499_,
		_w19848_,
		_w31473_
	);
	LUT2 #(
		.INIT('h2)
	) name27427 (
		_w19501_,
		_w31472_,
		_w31474_
	);
	LUT2 #(
		.INIT('h4)
	) name27428 (
		_w31473_,
		_w31474_,
		_w31475_
	);
	LUT2 #(
		.INIT('h2)
	) name27429 (
		\core_eu_em_mac_em_reg_mr1swe_DO_reg[10]/P0001 ,
		_w19383_,
		_w31476_
	);
	LUT2 #(
		.INIT('h1)
	) name27430 (
		_w19508_,
		_w31476_,
		_w31477_
	);
	LUT2 #(
		.INIT('h4)
	) name27431 (
		_w31475_,
		_w31477_,
		_w31478_
	);
	LUT2 #(
		.INIT('h1)
	) name27432 (
		_w18262_,
		_w31478_,
		_w31479_
	);
	LUT2 #(
		.INIT('h1)
	) name27433 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19516_,
		_w31480_
	);
	LUT2 #(
		.INIT('h8)
	) name27434 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w19434_,
		_w31481_
	);
	LUT2 #(
		.INIT('h1)
	) name27435 (
		_w31480_,
		_w31481_,
		_w31482_
	);
	LUT2 #(
		.INIT('h2)
	) name27436 (
		_w18262_,
		_w31482_,
		_w31483_
	);
	LUT2 #(
		.INIT('h1)
	) name27437 (
		_w31479_,
		_w31483_,
		_w31484_
	);
	LUT2 #(
		.INIT('h8)
	) name27438 (
		_w14752_,
		_w31482_,
		_w31485_
	);
	LUT2 #(
		.INIT('h8)
	) name27439 (
		_w19776_,
		_w19848_,
		_w31486_
	);
	LUT2 #(
		.INIT('h2)
	) name27440 (
		\core_eu_em_mac_em_reg_mr1rwe_DO_reg[10]/P0001 ,
		_w17809_,
		_w31487_
	);
	LUT2 #(
		.INIT('h2)
	) name27441 (
		_w19780_,
		_w31487_,
		_w31488_
	);
	LUT2 #(
		.INIT('h4)
	) name27442 (
		_w31486_,
		_w31488_,
		_w31489_
	);
	LUT2 #(
		.INIT('h1)
	) name27443 (
		_w31485_,
		_w31489_,
		_w31490_
	);
	LUT2 #(
		.INIT('h4)
	) name27444 (
		\clkc_STDcnt_reg[8]/NET0131 ,
		\clkc_ckr_reg_DO_reg[5]/NET0131 ,
		_w31491_
	);
	LUT2 #(
		.INIT('h1)
	) name27445 (
		\clkc_STDcnt_reg[9]/NET0131 ,
		\clkc_ckr_reg_DO_reg[6]/NET0131 ,
		_w31492_
	);
	LUT2 #(
		.INIT('h8)
	) name27446 (
		\clkc_STDcnt_reg[9]/NET0131 ,
		\clkc_ckr_reg_DO_reg[6]/NET0131 ,
		_w31493_
	);
	LUT2 #(
		.INIT('h1)
	) name27447 (
		_w31492_,
		_w31493_,
		_w31494_
	);
	LUT2 #(
		.INIT('h2)
	) name27448 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		\clkc_ckr_reg_DO_reg[4]/NET0131 ,
		_w31495_
	);
	LUT2 #(
		.INIT('h4)
	) name27449 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		\clkc_ckr_reg_DO_reg[4]/NET0131 ,
		_w31496_
	);
	LUT2 #(
		.INIT('h1)
	) name27450 (
		\clkc_STDcnt_reg[10]/NET0131 ,
		\clkc_ckr_reg_DO_reg[7]/NET0131 ,
		_w31497_
	);
	LUT2 #(
		.INIT('h8)
	) name27451 (
		\clkc_STDcnt_reg[10]/NET0131 ,
		\clkc_ckr_reg_DO_reg[7]/NET0131 ,
		_w31498_
	);
	LUT2 #(
		.INIT('h1)
	) name27452 (
		_w31497_,
		_w31498_,
		_w31499_
	);
	LUT2 #(
		.INIT('h4)
	) name27453 (
		\clkc_STDcnt_reg[5]/NET0131 ,
		\clkc_ckr_reg_DO_reg[2]/NET0131 ,
		_w31500_
	);
	LUT2 #(
		.INIT('h2)
	) name27454 (
		\clkc_STDcnt_reg[5]/NET0131 ,
		\clkc_ckr_reg_DO_reg[2]/NET0131 ,
		_w31501_
	);
	LUT2 #(
		.INIT('h2)
	) name27455 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		\clkc_ckr_reg_DO_reg[1]/NET0131 ,
		_w31502_
	);
	LUT2 #(
		.INIT('h4)
	) name27456 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		\clkc_ckr_reg_DO_reg[1]/NET0131 ,
		_w31503_
	);
	LUT2 #(
		.INIT('h4)
	) name27457 (
		\clkc_STDcnt_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[3]/NET0131 ,
		_w31504_
	);
	LUT2 #(
		.INIT('h2)
	) name27458 (
		\clkc_STDcnt_reg[3]/NET0131 ,
		\clkc_ckr_reg_DO_reg[0]/NET0131 ,
		_w31505_
	);
	LUT2 #(
		.INIT('h2)
	) name27459 (
		\clkc_STDcnt_reg[6]/NET0131 ,
		\clkc_ckr_reg_DO_reg[3]/NET0131 ,
		_w31506_
	);
	LUT2 #(
		.INIT('h4)
	) name27460 (
		\clkc_STDcnt_reg[3]/NET0131 ,
		\clkc_ckr_reg_DO_reg[0]/NET0131 ,
		_w31507_
	);
	LUT2 #(
		.INIT('h2)
	) name27461 (
		\clkc_STDcnt_reg[8]/NET0131 ,
		\clkc_ckr_reg_DO_reg[5]/NET0131 ,
		_w31508_
	);
	LUT2 #(
		.INIT('h1)
	) name27462 (
		_w31491_,
		_w31495_,
		_w31509_
	);
	LUT2 #(
		.INIT('h1)
	) name27463 (
		_w31496_,
		_w31500_,
		_w31510_
	);
	LUT2 #(
		.INIT('h1)
	) name27464 (
		_w31501_,
		_w31502_,
		_w31511_
	);
	LUT2 #(
		.INIT('h1)
	) name27465 (
		_w31503_,
		_w31504_,
		_w31512_
	);
	LUT2 #(
		.INIT('h1)
	) name27466 (
		_w31505_,
		_w31506_,
		_w31513_
	);
	LUT2 #(
		.INIT('h1)
	) name27467 (
		_w31507_,
		_w31508_,
		_w31514_
	);
	LUT2 #(
		.INIT('h8)
	) name27468 (
		_w31513_,
		_w31514_,
		_w31515_
	);
	LUT2 #(
		.INIT('h8)
	) name27469 (
		_w31511_,
		_w31512_,
		_w31516_
	);
	LUT2 #(
		.INIT('h8)
	) name27470 (
		_w31509_,
		_w31510_,
		_w31517_
	);
	LUT2 #(
		.INIT('h1)
	) name27471 (
		_w31494_,
		_w31499_,
		_w31518_
	);
	LUT2 #(
		.INIT('h8)
	) name27472 (
		_w31517_,
		_w31518_,
		_w31519_
	);
	LUT2 #(
		.INIT('h8)
	) name27473 (
		_w31515_,
		_w31516_,
		_w31520_
	);
	LUT2 #(
		.INIT('h8)
	) name27474 (
		_w31519_,
		_w31520_,
		_w31521_
	);
	LUT2 #(
		.INIT('h8)
	) name27475 (
		\clkc_STDcnt_reg[0]/NET0131 ,
		\clkc_STDcnt_reg[1]/NET0131 ,
		_w31522_
	);
	LUT2 #(
		.INIT('h8)
	) name27476 (
		\clkc_STDcnt_reg[2]/NET0131 ,
		_w31522_,
		_w31523_
	);
	LUT2 #(
		.INIT('h8)
	) name27477 (
		\clkc_STDcnt_reg[3]/NET0131 ,
		_w31523_,
		_w31524_
	);
	LUT2 #(
		.INIT('h8)
	) name27478 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		_w31524_,
		_w31525_
	);
	LUT2 #(
		.INIT('h8)
	) name27479 (
		\clkc_STDcnt_reg[5]/NET0131 ,
		_w31525_,
		_w31526_
	);
	LUT2 #(
		.INIT('h8)
	) name27480 (
		\clkc_STDcnt_reg[6]/NET0131 ,
		_w31526_,
		_w31527_
	);
	LUT2 #(
		.INIT('h8)
	) name27481 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		_w31527_,
		_w31528_
	);
	LUT2 #(
		.INIT('h8)
	) name27482 (
		\clkc_STDcnt_reg[8]/NET0131 ,
		_w31528_,
		_w31529_
	);
	LUT2 #(
		.INIT('h8)
	) name27483 (
		\clkc_STDcnt_reg[9]/NET0131 ,
		_w31529_,
		_w31530_
	);
	LUT2 #(
		.INIT('h1)
	) name27484 (
		\clkc_STDcnt_reg[10]/NET0131 ,
		_w31530_,
		_w31531_
	);
	LUT2 #(
		.INIT('h8)
	) name27485 (
		\clkc_STDcnt_reg[10]/NET0131 ,
		_w31530_,
		_w31532_
	);
	LUT2 #(
		.INIT('h1)
	) name27486 (
		_w31521_,
		_w31531_,
		_w31533_
	);
	LUT2 #(
		.INIT('h4)
	) name27487 (
		_w31532_,
		_w31533_,
		_w31534_
	);
	LUT2 #(
		.INIT('h2)
	) name27488 (
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		_w4116_,
		_w31535_
	);
	LUT2 #(
		.INIT('h4)
	) name27489 (
		\sport0_regs_AUTOreg_DO_reg[1]/NET0131 ,
		\sport0_txctl_c_sync1_reg/P0001 ,
		_w31536_
	);
	LUT2 #(
		.INIT('h4)
	) name27490 (
		\sport0_txctl_c_sync2_reg/P0001 ,
		_w31536_,
		_w31537_
	);
	LUT2 #(
		.INIT('h8)
	) name27491 (
		\core_dag_modulo1_T0wrap_reg/P0001 ,
		\sport0_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w31538_
	);
	LUT2 #(
		.INIT('h1)
	) name27492 (
		\core_c_psq_IFC_reg[14]/NET0131 ,
		\core_c_psq_Iflag_reg[6]/NET0131 ,
		_w31539_
	);
	LUT2 #(
		.INIT('h4)
	) name27493 (
		_w31538_,
		_w31539_,
		_w31540_
	);
	LUT2 #(
		.INIT('h4)
	) name27494 (
		_w31537_,
		_w31540_,
		_w31541_
	);
	LUT2 #(
		.INIT('h1)
	) name27495 (
		\core_c_psq_IFC_reg[6]/NET0131 ,
		_w31541_,
		_w31542_
	);
	LUT2 #(
		.INIT('h4)
	) name27496 (
		_w31535_,
		_w31542_,
		_w31543_
	);
	LUT2 #(
		.INIT('h4)
	) name27497 (
		\core_c_dec_MTMX1_E_reg/P0001 ,
		_w4117_,
		_w31544_
	);
	LUT2 #(
		.INIT('h4)
	) name27498 (
		_w31076_,
		_w31079_,
		_w31545_
	);
	LUT2 #(
		.INIT('h8)
	) name27499 (
		_w31103_,
		_w31545_,
		_w31546_
	);
	LUT2 #(
		.INIT('h8)
	) name27500 (
		_w6023_,
		_w6025_,
		_w31547_
	);
	LUT2 #(
		.INIT('h1)
	) name27501 (
		_w4117_,
		_w31547_,
		_w31548_
	);
	LUT2 #(
		.INIT('h4)
	) name27502 (
		_w31546_,
		_w31548_,
		_w31549_
	);
	LUT2 #(
		.INIT('h2)
	) name27503 (
		_w4116_,
		_w31544_,
		_w31550_
	);
	LUT2 #(
		.INIT('h4)
	) name27504 (
		_w31549_,
		_w31550_,
		_w31551_
	);
	LUT2 #(
		.INIT('h4)
	) name27505 (
		\core_c_dec_MTMX0_E_reg/P0001 ,
		_w4117_,
		_w31552_
	);
	LUT2 #(
		.INIT('h8)
	) name27506 (
		_w31112_,
		_w31545_,
		_w31553_
	);
	LUT2 #(
		.INIT('h8)
	) name27507 (
		_w6023_,
		_w19697_,
		_w31554_
	);
	LUT2 #(
		.INIT('h1)
	) name27508 (
		_w4117_,
		_w31554_,
		_w31555_
	);
	LUT2 #(
		.INIT('h4)
	) name27509 (
		_w31553_,
		_w31555_,
		_w31556_
	);
	LUT2 #(
		.INIT('h2)
	) name27510 (
		_w4116_,
		_w31552_,
		_w31557_
	);
	LUT2 #(
		.INIT('h4)
	) name27511 (
		_w31556_,
		_w31557_,
		_w31558_
	);
	LUT2 #(
		.INIT('h4)
	) name27512 (
		\core_c_dec_MTAX1_E_reg/P0001 ,
		_w4117_,
		_w31559_
	);
	LUT2 #(
		.INIT('h8)
	) name27513 (
		_w6023_,
		_w20606_,
		_w31560_
	);
	LUT2 #(
		.INIT('h2)
	) name27514 (
		_w31079_,
		_w31089_,
		_w31561_
	);
	LUT2 #(
		.INIT('h8)
	) name27515 (
		_w31094_,
		_w31121_,
		_w31562_
	);
	LUT2 #(
		.INIT('h4)
	) name27516 (
		_w31098_,
		_w31561_,
		_w31563_
	);
	LUT2 #(
		.INIT('h8)
	) name27517 (
		_w31562_,
		_w31563_,
		_w31564_
	);
	LUT2 #(
		.INIT('h1)
	) name27518 (
		_w4117_,
		_w31560_,
		_w31565_
	);
	LUT2 #(
		.INIT('h4)
	) name27519 (
		_w31564_,
		_w31565_,
		_w31566_
	);
	LUT2 #(
		.INIT('h2)
	) name27520 (
		_w4116_,
		_w31559_,
		_w31567_
	);
	LUT2 #(
		.INIT('h4)
	) name27521 (
		_w31566_,
		_w31567_,
		_w31568_
	);
	LUT2 #(
		.INIT('h1)
	) name27522 (
		\sport0_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		_w19552_,
		_w31569_
	);
	LUT2 #(
		.INIT('h2)
	) name27523 (
		_w19197_,
		_w29228_,
		_w31570_
	);
	LUT2 #(
		.INIT('h4)
	) name27524 (
		_w31569_,
		_w31570_,
		_w31571_
	);
	LUT2 #(
		.INIT('h4)
	) name27525 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w17789_,
		_w31572_
	);
	LUT2 #(
		.INIT('h8)
	) name27526 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w25067_,
		_w31573_
	);
	LUT2 #(
		.INIT('h1)
	) name27527 (
		_w31572_,
		_w31573_,
		_w31574_
	);
	LUT2 #(
		.INIT('h1)
	) name27528 (
		\sport1_cfg_SCLKi_cnt_reg[14]/NET0131 ,
		_w20253_,
		_w31575_
	);
	LUT2 #(
		.INIT('h2)
	) name27529 (
		_w19130_,
		_w29407_,
		_w31576_
	);
	LUT2 #(
		.INIT('h4)
	) name27530 (
		_w31575_,
		_w31576_,
		_w31577_
	);
	LUT2 #(
		.INIT('h8)
	) name27531 (
		_w6116_,
		_w25725_,
		_w31578_
	);
	LUT2 #(
		.INIT('h8)
	) name27532 (
		\core_c_dec_MTAX0_E_reg/P0001 ,
		_w4117_,
		_w31579_
	);
	LUT2 #(
		.INIT('h8)
	) name27533 (
		_w31098_,
		_w31561_,
		_w31580_
	);
	LUT2 #(
		.INIT('h4)
	) name27534 (
		_w4117_,
		_w31580_,
		_w31581_
	);
	LUT2 #(
		.INIT('h8)
	) name27535 (
		_w31562_,
		_w31581_,
		_w31582_
	);
	LUT2 #(
		.INIT('h1)
	) name27536 (
		_w31578_,
		_w31579_,
		_w31583_
	);
	LUT2 #(
		.INIT('h4)
	) name27537 (
		_w31582_,
		_w31583_,
		_w31584_
	);
	LUT2 #(
		.INIT('h2)
	) name27538 (
		_w4116_,
		_w31584_,
		_w31585_
	);
	LUT2 #(
		.INIT('h1)
	) name27539 (
		\sport1_cfg_FSi_reg/NET0131 ,
		_w28854_,
		_w31586_
	);
	LUT2 #(
		.INIT('h8)
	) name27540 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		_w31587_
	);
	LUT2 #(
		.INIT('h8)
	) name27541 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		_w31588_
	);
	LUT2 #(
		.INIT('h4)
	) name27542 (
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w31589_
	);
	LUT2 #(
		.INIT('h8)
	) name27543 (
		_w31588_,
		_w31589_,
		_w31590_
	);
	LUT2 #(
		.INIT('h8)
	) name27544 (
		_w31587_,
		_w31590_,
		_w31591_
	);
	LUT2 #(
		.INIT('h4)
	) name27545 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w31592_
	);
	LUT2 #(
		.INIT('h2)
	) name27546 (
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w31593_
	);
	LUT2 #(
		.INIT('h2)
	) name27547 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w31594_
	);
	LUT2 #(
		.INIT('h4)
	) name27548 (
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w31595_
	);
	LUT2 #(
		.INIT('h2)
	) name27549 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w31596_
	);
	LUT2 #(
		.INIT('h4)
	) name27550 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w31597_
	);
	LUT2 #(
		.INIT('h4)
	) name27551 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w31598_
	);
	LUT2 #(
		.INIT('h2)
	) name27552 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w31599_
	);
	LUT2 #(
		.INIT('h2)
	) name27553 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w31600_
	);
	LUT2 #(
		.INIT('h4)
	) name27554 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w31601_
	);
	LUT2 #(
		.INIT('h1)
	) name27555 (
		_w31592_,
		_w31593_,
		_w31602_
	);
	LUT2 #(
		.INIT('h1)
	) name27556 (
		_w31594_,
		_w31595_,
		_w31603_
	);
	LUT2 #(
		.INIT('h1)
	) name27557 (
		_w31596_,
		_w31597_,
		_w31604_
	);
	LUT2 #(
		.INIT('h1)
	) name27558 (
		_w31598_,
		_w31599_,
		_w31605_
	);
	LUT2 #(
		.INIT('h1)
	) name27559 (
		_w31600_,
		_w31601_,
		_w31606_
	);
	LUT2 #(
		.INIT('h8)
	) name27560 (
		_w31605_,
		_w31606_,
		_w31607_
	);
	LUT2 #(
		.INIT('h8)
	) name27561 (
		_w31603_,
		_w31604_,
		_w31608_
	);
	LUT2 #(
		.INIT('h8)
	) name27562 (
		_w31602_,
		_w31608_,
		_w31609_
	);
	LUT2 #(
		.INIT('h8)
	) name27563 (
		_w31607_,
		_w31609_,
		_w31610_
	);
	LUT2 #(
		.INIT('h8)
	) name27564 (
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		\sport1_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w31611_
	);
	LUT2 #(
		.INIT('h4)
	) name27565 (
		_w31591_,
		_w31611_,
		_w31612_
	);
	LUT2 #(
		.INIT('h4)
	) name27566 (
		_w31610_,
		_w31612_,
		_w31613_
	);
	LUT2 #(
		.INIT('h2)
	) name27567 (
		\sport1_cfg_FSi_reg/NET0131 ,
		_w31613_,
		_w31614_
	);
	LUT2 #(
		.INIT('h1)
	) name27568 (
		_w31586_,
		_w31614_,
		_w31615_
	);
	LUT2 #(
		.INIT('h1)
	) name27569 (
		\sport0_cfg_FSi_reg/NET0131 ,
		_w28944_,
		_w31616_
	);
	LUT2 #(
		.INIT('h8)
	) name27570 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		_w31617_
	);
	LUT2 #(
		.INIT('h8)
	) name27571 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		_w31618_
	);
	LUT2 #(
		.INIT('h4)
	) name27572 (
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w31619_
	);
	LUT2 #(
		.INIT('h8)
	) name27573 (
		_w31618_,
		_w31619_,
		_w31620_
	);
	LUT2 #(
		.INIT('h8)
	) name27574 (
		_w31617_,
		_w31620_,
		_w31621_
	);
	LUT2 #(
		.INIT('h4)
	) name27575 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w31622_
	);
	LUT2 #(
		.INIT('h2)
	) name27576 (
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w31623_
	);
	LUT2 #(
		.INIT('h2)
	) name27577 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w31624_
	);
	LUT2 #(
		.INIT('h4)
	) name27578 (
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w31625_
	);
	LUT2 #(
		.INIT('h2)
	) name27579 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w31626_
	);
	LUT2 #(
		.INIT('h4)
	) name27580 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w31627_
	);
	LUT2 #(
		.INIT('h4)
	) name27581 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w31628_
	);
	LUT2 #(
		.INIT('h2)
	) name27582 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w31629_
	);
	LUT2 #(
		.INIT('h2)
	) name27583 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w31630_
	);
	LUT2 #(
		.INIT('h4)
	) name27584 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w31631_
	);
	LUT2 #(
		.INIT('h1)
	) name27585 (
		_w31622_,
		_w31623_,
		_w31632_
	);
	LUT2 #(
		.INIT('h1)
	) name27586 (
		_w31624_,
		_w31625_,
		_w31633_
	);
	LUT2 #(
		.INIT('h1)
	) name27587 (
		_w31626_,
		_w31627_,
		_w31634_
	);
	LUT2 #(
		.INIT('h1)
	) name27588 (
		_w31628_,
		_w31629_,
		_w31635_
	);
	LUT2 #(
		.INIT('h1)
	) name27589 (
		_w31630_,
		_w31631_,
		_w31636_
	);
	LUT2 #(
		.INIT('h8)
	) name27590 (
		_w31635_,
		_w31636_,
		_w31637_
	);
	LUT2 #(
		.INIT('h8)
	) name27591 (
		_w31633_,
		_w31634_,
		_w31638_
	);
	LUT2 #(
		.INIT('h8)
	) name27592 (
		_w31632_,
		_w31638_,
		_w31639_
	);
	LUT2 #(
		.INIT('h8)
	) name27593 (
		_w31637_,
		_w31639_,
		_w31640_
	);
	LUT2 #(
		.INIT('h8)
	) name27594 (
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		\sport0_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w31641_
	);
	LUT2 #(
		.INIT('h4)
	) name27595 (
		_w31621_,
		_w31641_,
		_w31642_
	);
	LUT2 #(
		.INIT('h4)
	) name27596 (
		_w31640_,
		_w31642_,
		_w31643_
	);
	LUT2 #(
		.INIT('h2)
	) name27597 (
		\sport0_cfg_FSi_reg/NET0131 ,
		_w31643_,
		_w31644_
	);
	LUT2 #(
		.INIT('h1)
	) name27598 (
		_w31616_,
		_w31644_,
		_w31645_
	);
	LUT2 #(
		.INIT('h8)
	) name27599 (
		\core_c_dec_pMFSHT_Ei_reg/NET0131 ,
		_w4117_,
		_w31646_
	);
	LUT2 #(
		.INIT('h4)
	) name27600 (
		_w30966_,
		_w30969_,
		_w31647_
	);
	LUT2 #(
		.INIT('h8)
	) name27601 (
		_w30970_,
		_w31647_,
		_w31648_
	);
	LUT2 #(
		.INIT('h8)
	) name27602 (
		_w30974_,
		_w31647_,
		_w31649_
	);
	LUT2 #(
		.INIT('h8)
	) name27603 (
		_w30958_,
		_w30961_,
		_w31650_
	);
	LUT2 #(
		.INIT('h4)
	) name27604 (
		_w30966_,
		_w31650_,
		_w31651_
	);
	LUT2 #(
		.INIT('h8)
	) name27605 (
		_w30970_,
		_w31651_,
		_w31652_
	);
	LUT2 #(
		.INIT('h8)
	) name27606 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w31653_
	);
	LUT2 #(
		.INIT('h8)
	) name27607 (
		_w31264_,
		_w31653_,
		_w31654_
	);
	LUT2 #(
		.INIT('h8)
	) name27608 (
		_w31271_,
		_w31654_,
		_w31655_
	);
	LUT2 #(
		.INIT('h8)
	) name27609 (
		_w30974_,
		_w31651_,
		_w31656_
	);
	LUT2 #(
		.INIT('h1)
	) name27610 (
		_w31648_,
		_w31655_,
		_w31657_
	);
	LUT2 #(
		.INIT('h1)
	) name27611 (
		_w31649_,
		_w31652_,
		_w31658_
	);
	LUT2 #(
		.INIT('h4)
	) name27612 (
		_w31656_,
		_w31658_,
		_w31659_
	);
	LUT2 #(
		.INIT('h8)
	) name27613 (
		_w31657_,
		_w31659_,
		_w31660_
	);
	LUT2 #(
		.INIT('h2)
	) name27614 (
		_w30934_,
		_w31660_,
		_w31661_
	);
	LUT2 #(
		.INIT('h1)
	) name27615 (
		_w31646_,
		_w31661_,
		_w31662_
	);
	LUT2 #(
		.INIT('h8)
	) name27616 (
		\core_c_dec_MFSHT_Ei_reg/NET0131 ,
		_w4117_,
		_w31663_
	);
	LUT2 #(
		.INIT('h2)
	) name27617 (
		_w25047_,
		_w31660_,
		_w31664_
	);
	LUT2 #(
		.INIT('h1)
	) name27618 (
		_w31663_,
		_w31664_,
		_w31665_
	);
	LUT2 #(
		.INIT('h2)
	) name27619 (
		\tm_tsr_reg_DO_reg[4]/NET0131 ,
		_w25491_,
		_w31666_
	);
	LUT2 #(
		.INIT('h2)
	) name27620 (
		\tm_TSR_TMP_reg[4]/NET0131 ,
		_w25493_,
		_w31667_
	);
	LUT2 #(
		.INIT('h1)
	) name27621 (
		_w25494_,
		_w31667_,
		_w31668_
	);
	LUT2 #(
		.INIT('h2)
	) name27622 (
		_w25491_,
		_w31668_,
		_w31669_
	);
	LUT2 #(
		.INIT('h1)
	) name27623 (
		_w31666_,
		_w31669_,
		_w31670_
	);
	LUT2 #(
		.INIT('h8)
	) name27624 (
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w28876_,
		_w31671_
	);
	LUT2 #(
		.INIT('h1)
	) name27625 (
		\sport0_cfg_FSi_cnt_reg[7]/NET0131 ,
		_w28952_,
		_w31672_
	);
	LUT2 #(
		.INIT('h1)
	) name27626 (
		_w28953_,
		_w31672_,
		_w31673_
	);
	LUT2 #(
		.INIT('h8)
	) name27627 (
		_w28945_,
		_w31673_,
		_w31674_
	);
	LUT2 #(
		.INIT('h1)
	) name27628 (
		_w31671_,
		_w31674_,
		_w31675_
	);
	LUT2 #(
		.INIT('h8)
	) name27629 (
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w28786_,
		_w31676_
	);
	LUT2 #(
		.INIT('h1)
	) name27630 (
		\sport1_cfg_FSi_cnt_reg[7]/NET0131 ,
		_w28862_,
		_w31677_
	);
	LUT2 #(
		.INIT('h1)
	) name27631 (
		_w28863_,
		_w31677_,
		_w31678_
	);
	LUT2 #(
		.INIT('h8)
	) name27632 (
		_w28855_,
		_w31678_,
		_w31679_
	);
	LUT2 #(
		.INIT('h1)
	) name27633 (
		_w31676_,
		_w31679_,
		_w31680_
	);
	LUT2 #(
		.INIT('h8)
	) name27634 (
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w28786_,
		_w31681_
	);
	LUT2 #(
		.INIT('h1)
	) name27635 (
		\sport1_cfg_FSi_cnt_reg[8]/NET0131 ,
		_w28863_,
		_w31682_
	);
	LUT2 #(
		.INIT('h2)
	) name27636 (
		_w28855_,
		_w28864_,
		_w31683_
	);
	LUT2 #(
		.INIT('h4)
	) name27637 (
		_w31682_,
		_w31683_,
		_w31684_
	);
	LUT2 #(
		.INIT('h1)
	) name27638 (
		_w31681_,
		_w31684_,
		_w31685_
	);
	LUT2 #(
		.INIT('h8)
	) name27639 (
		\sport0_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w28876_,
		_w31686_
	);
	LUT2 #(
		.INIT('h1)
	) name27640 (
		\sport0_cfg_FSi_cnt_reg[8]/NET0131 ,
		_w28953_,
		_w31687_
	);
	LUT2 #(
		.INIT('h2)
	) name27641 (
		_w28945_,
		_w28954_,
		_w31688_
	);
	LUT2 #(
		.INIT('h4)
	) name27642 (
		_w31687_,
		_w31688_,
		_w31689_
	);
	LUT2 #(
		.INIT('h1)
	) name27643 (
		_w31686_,
		_w31689_,
		_w31690_
	);
	LUT2 #(
		.INIT('h1)
	) name27644 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[1]/NET0131 ,
		_w31691_
	);
	LUT2 #(
		.INIT('h4)
	) name27645 (
		\sport1_rxctl_Bcnt_reg[2]/NET0131 ,
		_w31691_,
		_w31692_
	);
	LUT2 #(
		.INIT('h4)
	) name27646 (
		\sport1_rxctl_Bcnt_reg[3]/NET0131 ,
		_w31692_,
		_w31693_
	);
	LUT2 #(
		.INIT('h2)
	) name27647 (
		\sport1_rxctl_Bcnt_reg[3]/NET0131 ,
		_w31692_,
		_w31694_
	);
	LUT2 #(
		.INIT('h1)
	) name27648 (
		_w31693_,
		_w31694_,
		_w31695_
	);
	LUT2 #(
		.INIT('h1)
	) name27649 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RCS_reg[2]/NET0131 ,
		_w31696_
	);
	LUT2 #(
		.INIT('h8)
	) name27650 (
		\sport1_rxctl_RCS_reg[1]/NET0131 ,
		_w31696_,
		_w31697_
	);
	LUT2 #(
		.INIT('h8)
	) name27651 (
		\sport1_rxctl_RCS_reg[0]/NET0131 ,
		\sport1_rxctl_RCS_reg[2]/NET0131 ,
		_w31698_
	);
	LUT2 #(
		.INIT('h1)
	) name27652 (
		\sport1_rxctl_RCS_reg[1]/NET0131 ,
		_w31696_,
		_w31699_
	);
	LUT2 #(
		.INIT('h4)
	) name27653 (
		_w31698_,
		_w31699_,
		_w31700_
	);
	LUT2 #(
		.INIT('h4)
	) name27654 (
		_w30750_,
		_w31700_,
		_w31701_
	);
	LUT2 #(
		.INIT('h1)
	) name27655 (
		_w31697_,
		_w31701_,
		_w31702_
	);
	LUT2 #(
		.INIT('h4)
	) name27656 (
		\sport1_rxctl_Bcnt_reg[4]/NET0131 ,
		_w31693_,
		_w31703_
	);
	LUT2 #(
		.INIT('h4)
	) name27657 (
		_w31701_,
		_w31703_,
		_w31704_
	);
	LUT2 #(
		.INIT('h1)
	) name27658 (
		_w31702_,
		_w31704_,
		_w31705_
	);
	LUT2 #(
		.INIT('h4)
	) name27659 (
		_w31695_,
		_w31705_,
		_w31706_
	);
	LUT2 #(
		.INIT('h2)
	) name27660 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w31705_,
		_w31707_
	);
	LUT2 #(
		.INIT('h1)
	) name27661 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w31706_,
		_w31708_
	);
	LUT2 #(
		.INIT('h4)
	) name27662 (
		_w31707_,
		_w31708_,
		_w31709_
	);
	LUT2 #(
		.INIT('h2)
	) name27663 (
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w31705_,
		_w31710_
	);
	LUT2 #(
		.INIT('h2)
	) name27664 (
		\sport1_rxctl_Bcnt_reg[2]/NET0131 ,
		_w31691_,
		_w31711_
	);
	LUT2 #(
		.INIT('h1)
	) name27665 (
		_w31692_,
		_w31711_,
		_w31712_
	);
	LUT2 #(
		.INIT('h2)
	) name27666 (
		_w31705_,
		_w31712_,
		_w31713_
	);
	LUT2 #(
		.INIT('h1)
	) name27667 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w31710_,
		_w31714_
	);
	LUT2 #(
		.INIT('h4)
	) name27668 (
		_w31713_,
		_w31714_,
		_w31715_
	);
	LUT2 #(
		.INIT('h2)
	) name27669 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w31705_,
		_w31716_
	);
	LUT2 #(
		.INIT('h8)
	) name27670 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Bcnt_reg[1]/NET0131 ,
		_w31717_
	);
	LUT2 #(
		.INIT('h1)
	) name27671 (
		_w31691_,
		_w31717_,
		_w31718_
	);
	LUT2 #(
		.INIT('h2)
	) name27672 (
		_w31705_,
		_w31718_,
		_w31719_
	);
	LUT2 #(
		.INIT('h1)
	) name27673 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w31716_,
		_w31720_
	);
	LUT2 #(
		.INIT('h4)
	) name27674 (
		_w31719_,
		_w31720_,
		_w31721_
	);
	LUT2 #(
		.INIT('h4)
	) name27675 (
		\sport1_rxctl_Bcnt_reg[0]/NET0131 ,
		_w31705_,
		_w31722_
	);
	LUT2 #(
		.INIT('h2)
	) name27676 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w31705_,
		_w31723_
	);
	LUT2 #(
		.INIT('h1)
	) name27677 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w31722_,
		_w31724_
	);
	LUT2 #(
		.INIT('h4)
	) name27678 (
		_w31723_,
		_w31724_,
		_w31725_
	);
	LUT2 #(
		.INIT('h8)
	) name27679 (
		_w11525_,
		_w31339_,
		_w31726_
	);
	LUT2 #(
		.INIT('h8)
	) name27680 (
		\core_dag_ilm2reg_M5_we_DO_reg[6]/NET0131 ,
		_w31341_,
		_w31727_
	);
	LUT2 #(
		.INIT('h8)
	) name27681 (
		\core_dag_ilm2reg_M6_we_DO_reg[6]/NET0131 ,
		_w31331_,
		_w31728_
	);
	LUT2 #(
		.INIT('h8)
	) name27682 (
		\core_dag_ilm2reg_M4_we_DO_reg[6]/NET0131 ,
		_w31344_,
		_w31729_
	);
	LUT2 #(
		.INIT('h8)
	) name27683 (
		\core_dag_ilm2reg_M7_we_DO_reg[6]/NET0131 ,
		_w31337_,
		_w31730_
	);
	LUT2 #(
		.INIT('h1)
	) name27684 (
		_w31728_,
		_w31730_,
		_w31731_
	);
	LUT2 #(
		.INIT('h4)
	) name27685 (
		_w31727_,
		_w31731_,
		_w31732_
	);
	LUT2 #(
		.INIT('h4)
	) name27686 (
		_w31729_,
		_w31732_,
		_w31733_
	);
	LUT2 #(
		.INIT('h4)
	) name27687 (
		_w31726_,
		_w31733_,
		_w31734_
	);
	LUT2 #(
		.INIT('h8)
	) name27688 (
		_w10911_,
		_w31339_,
		_w31735_
	);
	LUT2 #(
		.INIT('h8)
	) name27689 (
		\core_dag_ilm2reg_M5_we_DO_reg[5]/NET0131 ,
		_w31341_,
		_w31736_
	);
	LUT2 #(
		.INIT('h8)
	) name27690 (
		\core_dag_ilm2reg_M6_we_DO_reg[5]/NET0131 ,
		_w31331_,
		_w31737_
	);
	LUT2 #(
		.INIT('h8)
	) name27691 (
		\core_dag_ilm2reg_M4_we_DO_reg[5]/NET0131 ,
		_w31344_,
		_w31738_
	);
	LUT2 #(
		.INIT('h8)
	) name27692 (
		\core_dag_ilm2reg_M7_we_DO_reg[5]/NET0131 ,
		_w31337_,
		_w31739_
	);
	LUT2 #(
		.INIT('h1)
	) name27693 (
		_w31737_,
		_w31739_,
		_w31740_
	);
	LUT2 #(
		.INIT('h4)
	) name27694 (
		_w31736_,
		_w31740_,
		_w31741_
	);
	LUT2 #(
		.INIT('h4)
	) name27695 (
		_w31738_,
		_w31741_,
		_w31742_
	);
	LUT2 #(
		.INIT('h4)
	) name27696 (
		_w31735_,
		_w31742_,
		_w31743_
	);
	LUT2 #(
		.INIT('h8)
	) name27697 (
		_w10069_,
		_w31339_,
		_w31744_
	);
	LUT2 #(
		.INIT('h8)
	) name27698 (
		\core_dag_ilm2reg_M4_we_DO_reg[4]/NET0131 ,
		_w31344_,
		_w31745_
	);
	LUT2 #(
		.INIT('h8)
	) name27699 (
		\core_dag_ilm2reg_M7_we_DO_reg[4]/NET0131 ,
		_w31337_,
		_w31746_
	);
	LUT2 #(
		.INIT('h8)
	) name27700 (
		\core_dag_ilm2reg_M5_we_DO_reg[4]/NET0131 ,
		_w31341_,
		_w31747_
	);
	LUT2 #(
		.INIT('h8)
	) name27701 (
		\core_dag_ilm2reg_M6_we_DO_reg[4]/NET0131 ,
		_w31331_,
		_w31748_
	);
	LUT2 #(
		.INIT('h1)
	) name27702 (
		_w31746_,
		_w31748_,
		_w31749_
	);
	LUT2 #(
		.INIT('h4)
	) name27703 (
		_w31745_,
		_w31749_,
		_w31750_
	);
	LUT2 #(
		.INIT('h4)
	) name27704 (
		_w31747_,
		_w31750_,
		_w31751_
	);
	LUT2 #(
		.INIT('h4)
	) name27705 (
		_w31744_,
		_w31751_,
		_w31752_
	);
	LUT2 #(
		.INIT('h8)
	) name27706 (
		_w8113_,
		_w31339_,
		_w31753_
	);
	LUT2 #(
		.INIT('h8)
	) name27707 (
		\core_dag_ilm2reg_M4_we_DO_reg[3]/NET0131 ,
		_w31344_,
		_w31754_
	);
	LUT2 #(
		.INIT('h8)
	) name27708 (
		\core_dag_ilm2reg_M7_we_DO_reg[3]/NET0131 ,
		_w31337_,
		_w31755_
	);
	LUT2 #(
		.INIT('h8)
	) name27709 (
		\core_dag_ilm2reg_M5_we_DO_reg[3]/NET0131 ,
		_w31341_,
		_w31756_
	);
	LUT2 #(
		.INIT('h8)
	) name27710 (
		\core_dag_ilm2reg_M6_we_DO_reg[3]/NET0131 ,
		_w31331_,
		_w31757_
	);
	LUT2 #(
		.INIT('h1)
	) name27711 (
		_w31755_,
		_w31757_,
		_w31758_
	);
	LUT2 #(
		.INIT('h4)
	) name27712 (
		_w31754_,
		_w31758_,
		_w31759_
	);
	LUT2 #(
		.INIT('h4)
	) name27713 (
		_w31756_,
		_w31759_,
		_w31760_
	);
	LUT2 #(
		.INIT('h4)
	) name27714 (
		_w31753_,
		_w31760_,
		_w31761_
	);
	LUT2 #(
		.INIT('h8)
	) name27715 (
		_w8715_,
		_w31339_,
		_w31762_
	);
	LUT2 #(
		.INIT('h8)
	) name27716 (
		\core_dag_ilm2reg_M4_we_DO_reg[2]/NET0131 ,
		_w31344_,
		_w31763_
	);
	LUT2 #(
		.INIT('h8)
	) name27717 (
		\core_dag_ilm2reg_M7_we_DO_reg[2]/NET0131 ,
		_w31337_,
		_w31764_
	);
	LUT2 #(
		.INIT('h8)
	) name27718 (
		\core_dag_ilm2reg_M5_we_DO_reg[2]/NET0131 ,
		_w31341_,
		_w31765_
	);
	LUT2 #(
		.INIT('h8)
	) name27719 (
		\core_dag_ilm2reg_M6_we_DO_reg[2]/NET0131 ,
		_w31331_,
		_w31766_
	);
	LUT2 #(
		.INIT('h1)
	) name27720 (
		_w31764_,
		_w31766_,
		_w31767_
	);
	LUT2 #(
		.INIT('h4)
	) name27721 (
		_w31763_,
		_w31767_,
		_w31768_
	);
	LUT2 #(
		.INIT('h4)
	) name27722 (
		_w31765_,
		_w31768_,
		_w31769_
	);
	LUT2 #(
		.INIT('h4)
	) name27723 (
		_w31762_,
		_w31769_,
		_w31770_
	);
	LUT2 #(
		.INIT('h8)
	) name27724 (
		_w9435_,
		_w31339_,
		_w31771_
	);
	LUT2 #(
		.INIT('h8)
	) name27725 (
		\core_dag_ilm2reg_M4_we_DO_reg[1]/NET0131 ,
		_w31344_,
		_w31772_
	);
	LUT2 #(
		.INIT('h8)
	) name27726 (
		\core_dag_ilm2reg_M7_we_DO_reg[1]/NET0131 ,
		_w31337_,
		_w31773_
	);
	LUT2 #(
		.INIT('h8)
	) name27727 (
		\core_dag_ilm2reg_M5_we_DO_reg[1]/NET0131 ,
		_w31341_,
		_w31774_
	);
	LUT2 #(
		.INIT('h8)
	) name27728 (
		\core_dag_ilm2reg_M6_we_DO_reg[1]/NET0131 ,
		_w31331_,
		_w31775_
	);
	LUT2 #(
		.INIT('h1)
	) name27729 (
		_w31773_,
		_w31775_,
		_w31776_
	);
	LUT2 #(
		.INIT('h4)
	) name27730 (
		_w31772_,
		_w31776_,
		_w31777_
	);
	LUT2 #(
		.INIT('h4)
	) name27731 (
		_w31774_,
		_w31777_,
		_w31778_
	);
	LUT2 #(
		.INIT('h4)
	) name27732 (
		_w31771_,
		_w31778_,
		_w31779_
	);
	LUT2 #(
		.INIT('h8)
	) name27733 (
		_w8715_,
		_w31409_,
		_w31780_
	);
	LUT2 #(
		.INIT('h8)
	) name27734 (
		\core_dag_ilm1reg_M0_we_DO_reg[2]/NET0131 ,
		_w31411_,
		_w31781_
	);
	LUT2 #(
		.INIT('h8)
	) name27735 (
		\core_dag_ilm1reg_M2_we_DO_reg[2]/NET0131 ,
		_w31401_,
		_w31782_
	);
	LUT2 #(
		.INIT('h8)
	) name27736 (
		\core_dag_ilm1reg_M1_we_DO_reg[2]/NET0131 ,
		_w31414_,
		_w31783_
	);
	LUT2 #(
		.INIT('h8)
	) name27737 (
		\core_dag_ilm1reg_M3_we_DO_reg[2]/NET0131 ,
		_w31407_,
		_w31784_
	);
	LUT2 #(
		.INIT('h1)
	) name27738 (
		_w31782_,
		_w31784_,
		_w31785_
	);
	LUT2 #(
		.INIT('h4)
	) name27739 (
		_w31781_,
		_w31785_,
		_w31786_
	);
	LUT2 #(
		.INIT('h4)
	) name27740 (
		_w31783_,
		_w31786_,
		_w31787_
	);
	LUT2 #(
		.INIT('h4)
	) name27741 (
		_w31780_,
		_w31787_,
		_w31788_
	);
	LUT2 #(
		.INIT('h8)
	) name27742 (
		_w9435_,
		_w31409_,
		_w31789_
	);
	LUT2 #(
		.INIT('h8)
	) name27743 (
		\core_dag_ilm1reg_M0_we_DO_reg[1]/NET0131 ,
		_w31411_,
		_w31790_
	);
	LUT2 #(
		.INIT('h8)
	) name27744 (
		\core_dag_ilm1reg_M2_we_DO_reg[1]/NET0131 ,
		_w31401_,
		_w31791_
	);
	LUT2 #(
		.INIT('h8)
	) name27745 (
		\core_dag_ilm1reg_M1_we_DO_reg[1]/NET0131 ,
		_w31414_,
		_w31792_
	);
	LUT2 #(
		.INIT('h8)
	) name27746 (
		\core_dag_ilm1reg_M3_we_DO_reg[1]/NET0131 ,
		_w31407_,
		_w31793_
	);
	LUT2 #(
		.INIT('h1)
	) name27747 (
		_w31791_,
		_w31793_,
		_w31794_
	);
	LUT2 #(
		.INIT('h4)
	) name27748 (
		_w31790_,
		_w31794_,
		_w31795_
	);
	LUT2 #(
		.INIT('h4)
	) name27749 (
		_w31792_,
		_w31795_,
		_w31796_
	);
	LUT2 #(
		.INIT('h4)
	) name27750 (
		_w31789_,
		_w31796_,
		_w31797_
	);
	LUT2 #(
		.INIT('h8)
	) name27751 (
		_w7607_,
		_w31409_,
		_w31798_
	);
	LUT2 #(
		.INIT('h8)
	) name27752 (
		\core_dag_ilm1reg_M0_we_DO_reg[0]/NET0131 ,
		_w31411_,
		_w31799_
	);
	LUT2 #(
		.INIT('h8)
	) name27753 (
		\core_dag_ilm1reg_M2_we_DO_reg[0]/NET0131 ,
		_w31401_,
		_w31800_
	);
	LUT2 #(
		.INIT('h8)
	) name27754 (
		\core_dag_ilm1reg_M1_we_DO_reg[0]/NET0131 ,
		_w31414_,
		_w31801_
	);
	LUT2 #(
		.INIT('h8)
	) name27755 (
		\core_dag_ilm1reg_M3_we_DO_reg[0]/NET0131 ,
		_w31407_,
		_w31802_
	);
	LUT2 #(
		.INIT('h1)
	) name27756 (
		_w31800_,
		_w31802_,
		_w31803_
	);
	LUT2 #(
		.INIT('h4)
	) name27757 (
		_w31799_,
		_w31803_,
		_w31804_
	);
	LUT2 #(
		.INIT('h4)
	) name27758 (
		_w31801_,
		_w31804_,
		_w31805_
	);
	LUT2 #(
		.INIT('h4)
	) name27759 (
		_w31798_,
		_w31805_,
		_w31806_
	);
	LUT2 #(
		.INIT('h8)
	) name27760 (
		_w11525_,
		_w31409_,
		_w31807_
	);
	LUT2 #(
		.INIT('h8)
	) name27761 (
		\core_dag_ilm1reg_M1_we_DO_reg[6]/NET0131 ,
		_w31414_,
		_w31808_
	);
	LUT2 #(
		.INIT('h8)
	) name27762 (
		\core_dag_ilm1reg_M3_we_DO_reg[6]/NET0131 ,
		_w31407_,
		_w31809_
	);
	LUT2 #(
		.INIT('h8)
	) name27763 (
		\core_dag_ilm1reg_M0_we_DO_reg[6]/NET0131 ,
		_w31411_,
		_w31810_
	);
	LUT2 #(
		.INIT('h8)
	) name27764 (
		\core_dag_ilm1reg_M2_we_DO_reg[6]/NET0131 ,
		_w31401_,
		_w31811_
	);
	LUT2 #(
		.INIT('h1)
	) name27765 (
		_w31809_,
		_w31811_,
		_w31812_
	);
	LUT2 #(
		.INIT('h4)
	) name27766 (
		_w31808_,
		_w31812_,
		_w31813_
	);
	LUT2 #(
		.INIT('h4)
	) name27767 (
		_w31810_,
		_w31813_,
		_w31814_
	);
	LUT2 #(
		.INIT('h4)
	) name27768 (
		_w31807_,
		_w31814_,
		_w31815_
	);
	LUT2 #(
		.INIT('h8)
	) name27769 (
		_w10911_,
		_w31409_,
		_w31816_
	);
	LUT2 #(
		.INIT('h8)
	) name27770 (
		\core_dag_ilm1reg_M1_we_DO_reg[5]/NET0131 ,
		_w31414_,
		_w31817_
	);
	LUT2 #(
		.INIT('h8)
	) name27771 (
		\core_dag_ilm1reg_M3_we_DO_reg[5]/NET0131 ,
		_w31407_,
		_w31818_
	);
	LUT2 #(
		.INIT('h8)
	) name27772 (
		\core_dag_ilm1reg_M0_we_DO_reg[5]/NET0131 ,
		_w31411_,
		_w31819_
	);
	LUT2 #(
		.INIT('h8)
	) name27773 (
		\core_dag_ilm1reg_M2_we_DO_reg[5]/NET0131 ,
		_w31401_,
		_w31820_
	);
	LUT2 #(
		.INIT('h1)
	) name27774 (
		_w31818_,
		_w31820_,
		_w31821_
	);
	LUT2 #(
		.INIT('h4)
	) name27775 (
		_w31817_,
		_w31821_,
		_w31822_
	);
	LUT2 #(
		.INIT('h4)
	) name27776 (
		_w31819_,
		_w31822_,
		_w31823_
	);
	LUT2 #(
		.INIT('h4)
	) name27777 (
		_w31816_,
		_w31823_,
		_w31824_
	);
	LUT2 #(
		.INIT('h8)
	) name27778 (
		_w10069_,
		_w31409_,
		_w31825_
	);
	LUT2 #(
		.INIT('h8)
	) name27779 (
		\core_dag_ilm1reg_M1_we_DO_reg[4]/NET0131 ,
		_w31414_,
		_w31826_
	);
	LUT2 #(
		.INIT('h8)
	) name27780 (
		\core_dag_ilm1reg_M3_we_DO_reg[4]/NET0131 ,
		_w31407_,
		_w31827_
	);
	LUT2 #(
		.INIT('h8)
	) name27781 (
		\core_dag_ilm1reg_M0_we_DO_reg[4]/NET0131 ,
		_w31411_,
		_w31828_
	);
	LUT2 #(
		.INIT('h8)
	) name27782 (
		\core_dag_ilm1reg_M2_we_DO_reg[4]/NET0131 ,
		_w31401_,
		_w31829_
	);
	LUT2 #(
		.INIT('h1)
	) name27783 (
		_w31827_,
		_w31829_,
		_w31830_
	);
	LUT2 #(
		.INIT('h4)
	) name27784 (
		_w31826_,
		_w31830_,
		_w31831_
	);
	LUT2 #(
		.INIT('h4)
	) name27785 (
		_w31828_,
		_w31831_,
		_w31832_
	);
	LUT2 #(
		.INIT('h4)
	) name27786 (
		_w31825_,
		_w31832_,
		_w31833_
	);
	LUT2 #(
		.INIT('h1)
	) name27787 (
		\sport0_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		_w19544_,
		_w31834_
	);
	LUT2 #(
		.INIT('h2)
	) name27788 (
		_w19197_,
		_w19545_,
		_w31835_
	);
	LUT2 #(
		.INIT('h4)
	) name27789 (
		_w31834_,
		_w31835_,
		_w31836_
	);
	LUT2 #(
		.INIT('h2)
	) name27790 (
		\core_eu_em_mac_em_reg_mfswe_DO_reg[10]/P0001 ,
		_w20864_,
		_w31837_
	);
	LUT2 #(
		.INIT('h2)
	) name27791 (
		_w20864_,
		_w31482_,
		_w31838_
	);
	LUT2 #(
		.INIT('h1)
	) name27792 (
		_w31837_,
		_w31838_,
		_w31839_
	);
	LUT2 #(
		.INIT('h8)
	) name27793 (
		\core_c_dec_MACdep_Eg_reg/P0001 ,
		_w4117_,
		_w31840_
	);
	LUT2 #(
		.INIT('h1)
	) name27794 (
		_w26346_,
		_w26371_,
		_w31841_
	);
	LUT2 #(
		.INIT('h2)
	) name27795 (
		\core_c_dec_updMR_E_reg/P0001 ,
		_w31841_,
		_w31842_
	);
	LUT2 #(
		.INIT('h8)
	) name27796 (
		\core_c_dec_updMF_E_reg/P0001 ,
		_w20470_,
		_w31843_
	);
	LUT2 #(
		.INIT('h4)
	) name27797 (
		_w26358_,
		_w31843_,
		_w31844_
	);
	LUT2 #(
		.INIT('h1)
	) name27798 (
		_w31842_,
		_w31844_,
		_w31845_
	);
	LUT2 #(
		.INIT('h2)
	) name27799 (
		_w18848_,
		_w31845_,
		_w31846_
	);
	LUT2 #(
		.INIT('h8)
	) name27800 (
		_w13803_,
		_w31846_,
		_w31847_
	);
	LUT2 #(
		.INIT('h1)
	) name27801 (
		_w31840_,
		_w31847_,
		_w31848_
	);
	LUT2 #(
		.INIT('h2)
	) name27802 (
		_w4116_,
		_w31848_,
		_w31849_
	);
	LUT2 #(
		.INIT('h1)
	) name27803 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w31705_,
		_w31850_
	);
	LUT2 #(
		.INIT('h2)
	) name27804 (
		\sport1_rxctl_Bcnt_reg[4]/NET0131 ,
		_w31693_,
		_w31851_
	);
	LUT2 #(
		.INIT('h1)
	) name27805 (
		_w31703_,
		_w31851_,
		_w31852_
	);
	LUT2 #(
		.INIT('h8)
	) name27806 (
		_w31705_,
		_w31852_,
		_w31853_
	);
	LUT2 #(
		.INIT('h1)
	) name27807 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w31850_,
		_w31854_
	);
	LUT2 #(
		.INIT('h4)
	) name27808 (
		_w31853_,
		_w31854_,
		_w31855_
	);
	LUT2 #(
		.INIT('h1)
	) name27809 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RCS_reg[2]/NET0131 ,
		_w31856_
	);
	LUT2 #(
		.INIT('h8)
	) name27810 (
		\sport0_rxctl_RCS_reg[1]/NET0131 ,
		_w31856_,
		_w31857_
	);
	LUT2 #(
		.INIT('h8)
	) name27811 (
		\sport0_rxctl_RCS_reg[0]/NET0131 ,
		\sport0_rxctl_RCS_reg[2]/NET0131 ,
		_w31858_
	);
	LUT2 #(
		.INIT('h1)
	) name27812 (
		\sport0_rxctl_RCS_reg[1]/NET0131 ,
		_w31856_,
		_w31859_
	);
	LUT2 #(
		.INIT('h4)
	) name27813 (
		_w31858_,
		_w31859_,
		_w31860_
	);
	LUT2 #(
		.INIT('h4)
	) name27814 (
		_w30774_,
		_w31860_,
		_w31861_
	);
	LUT2 #(
		.INIT('h1)
	) name27815 (
		_w31857_,
		_w31861_,
		_w31862_
	);
	LUT2 #(
		.INIT('h1)
	) name27816 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[1]/NET0131 ,
		_w31863_
	);
	LUT2 #(
		.INIT('h4)
	) name27817 (
		\sport0_rxctl_Bcnt_reg[2]/NET0131 ,
		_w31863_,
		_w31864_
	);
	LUT2 #(
		.INIT('h4)
	) name27818 (
		\sport0_rxctl_Bcnt_reg[3]/NET0131 ,
		_w31864_,
		_w31865_
	);
	LUT2 #(
		.INIT('h4)
	) name27819 (
		\sport0_rxctl_Bcnt_reg[4]/NET0131 ,
		_w31865_,
		_w31866_
	);
	LUT2 #(
		.INIT('h4)
	) name27820 (
		_w31861_,
		_w31866_,
		_w31867_
	);
	LUT2 #(
		.INIT('h1)
	) name27821 (
		_w31862_,
		_w31867_,
		_w31868_
	);
	LUT2 #(
		.INIT('h1)
	) name27822 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w31868_,
		_w31869_
	);
	LUT2 #(
		.INIT('h2)
	) name27823 (
		\sport0_rxctl_Bcnt_reg[4]/NET0131 ,
		_w31865_,
		_w31870_
	);
	LUT2 #(
		.INIT('h1)
	) name27824 (
		_w31866_,
		_w31870_,
		_w31871_
	);
	LUT2 #(
		.INIT('h8)
	) name27825 (
		_w31868_,
		_w31871_,
		_w31872_
	);
	LUT2 #(
		.INIT('h1)
	) name27826 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w31869_,
		_w31873_
	);
	LUT2 #(
		.INIT('h4)
	) name27827 (
		_w31872_,
		_w31873_,
		_w31874_
	);
	LUT2 #(
		.INIT('h2)
	) name27828 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w31868_,
		_w31875_
	);
	LUT2 #(
		.INIT('h2)
	) name27829 (
		\sport0_rxctl_Bcnt_reg[3]/NET0131 ,
		_w31864_,
		_w31876_
	);
	LUT2 #(
		.INIT('h1)
	) name27830 (
		_w31865_,
		_w31876_,
		_w31877_
	);
	LUT2 #(
		.INIT('h2)
	) name27831 (
		_w31868_,
		_w31877_,
		_w31878_
	);
	LUT2 #(
		.INIT('h1)
	) name27832 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w31875_,
		_w31879_
	);
	LUT2 #(
		.INIT('h4)
	) name27833 (
		_w31878_,
		_w31879_,
		_w31880_
	);
	LUT2 #(
		.INIT('h2)
	) name27834 (
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w31868_,
		_w31881_
	);
	LUT2 #(
		.INIT('h2)
	) name27835 (
		\sport0_rxctl_Bcnt_reg[2]/NET0131 ,
		_w31863_,
		_w31882_
	);
	LUT2 #(
		.INIT('h1)
	) name27836 (
		_w31864_,
		_w31882_,
		_w31883_
	);
	LUT2 #(
		.INIT('h2)
	) name27837 (
		_w31868_,
		_w31883_,
		_w31884_
	);
	LUT2 #(
		.INIT('h1)
	) name27838 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w31881_,
		_w31885_
	);
	LUT2 #(
		.INIT('h4)
	) name27839 (
		_w31884_,
		_w31885_,
		_w31886_
	);
	LUT2 #(
		.INIT('h2)
	) name27840 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w31868_,
		_w31887_
	);
	LUT2 #(
		.INIT('h8)
	) name27841 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Bcnt_reg[1]/NET0131 ,
		_w31888_
	);
	LUT2 #(
		.INIT('h1)
	) name27842 (
		_w31863_,
		_w31888_,
		_w31889_
	);
	LUT2 #(
		.INIT('h2)
	) name27843 (
		_w31868_,
		_w31889_,
		_w31890_
	);
	LUT2 #(
		.INIT('h1)
	) name27844 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w31887_,
		_w31891_
	);
	LUT2 #(
		.INIT('h4)
	) name27845 (
		_w31890_,
		_w31891_,
		_w31892_
	);
	LUT2 #(
		.INIT('h4)
	) name27846 (
		\sport0_rxctl_Bcnt_reg[0]/NET0131 ,
		_w31868_,
		_w31893_
	);
	LUT2 #(
		.INIT('h2)
	) name27847 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w31868_,
		_w31894_
	);
	LUT2 #(
		.INIT('h1)
	) name27848 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w31893_,
		_w31895_
	);
	LUT2 #(
		.INIT('h4)
	) name27849 (
		_w31894_,
		_w31895_,
		_w31896_
	);
	LUT2 #(
		.INIT('h1)
	) name27850 (
		\sport1_cfg_SCLKi_cnt_reg[7]/NET0131 ,
		_w20236_,
		_w31897_
	);
	LUT2 #(
		.INIT('h2)
	) name27851 (
		_w19130_,
		_w20237_,
		_w31898_
	);
	LUT2 #(
		.INIT('h4)
	) name27852 (
		_w31897_,
		_w31898_,
		_w31899_
	);
	LUT2 #(
		.INIT('h2)
	) name27853 (
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		_w4116_,
		_w31900_
	);
	LUT2 #(
		.INIT('h4)
	) name27854 (
		\sport0_regs_AUTOreg_DO_reg[0]/NET0131 ,
		\sport0_rxctl_ISRa_reg/P0001 ,
		_w31901_
	);
	LUT2 #(
		.INIT('h8)
	) name27855 (
		\core_dag_modulo1_R0wrap_reg/P0001 ,
		\sport0_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w31902_
	);
	LUT2 #(
		.INIT('h1)
	) name27856 (
		\core_c_psq_IFC_reg[13]/NET0131 ,
		\core_c_psq_Iflag_reg[5]/NET0131 ,
		_w31903_
	);
	LUT2 #(
		.INIT('h4)
	) name27857 (
		_w31901_,
		_w31903_,
		_w31904_
	);
	LUT2 #(
		.INIT('h4)
	) name27858 (
		_w31902_,
		_w31904_,
		_w31905_
	);
	LUT2 #(
		.INIT('h1)
	) name27859 (
		\core_c_psq_IFC_reg[5]/NET0131 ,
		_w31905_,
		_w31906_
	);
	LUT2 #(
		.INIT('h4)
	) name27860 (
		_w31900_,
		_w31906_,
		_w31907_
	);
	LUT2 #(
		.INIT('h8)
	) name27861 (
		\sport0_regs_AUTO_a_reg[14]/NET0131 ,
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w31908_
	);
	LUT2 #(
		.INIT('h2)
	) name27862 (
		\clkc_Cnt128_reg/NET0131 ,
		_w31908_,
		_w31909_
	);
	LUT2 #(
		.INIT('h4)
	) name27863 (
		\clkc_oscntr_reg_DO_reg[10]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		_w31910_
	);
	LUT2 #(
		.INIT('h1)
	) name27864 (
		\clkc_oscntr_reg_DO_reg[10]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[11]/NET0131 ,
		_w31911_
	);
	LUT2 #(
		.INIT('h1)
	) name27865 (
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		_w31912_
	);
	LUT2 #(
		.INIT('h8)
	) name27866 (
		_w31911_,
		_w31912_,
		_w31913_
	);
	LUT2 #(
		.INIT('h2)
	) name27867 (
		\T_TMODE[0]_pad ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		_w31914_
	);
	LUT2 #(
		.INIT('h8)
	) name27868 (
		_w31913_,
		_w31914_,
		_w31915_
	);
	LUT2 #(
		.INIT('h4)
	) name27869 (
		\T_TMODE[0]_pad ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		_w31916_
	);
	LUT2 #(
		.INIT('h8)
	) name27870 (
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		_w31916_,
		_w31917_
	);
	LUT2 #(
		.INIT('h8)
	) name27871 (
		\clkc_oscntr_reg_DO_reg[11]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		_w31918_
	);
	LUT2 #(
		.INIT('h8)
	) name27872 (
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w31918_,
		_w31919_
	);
	LUT2 #(
		.INIT('h8)
	) name27873 (
		_w31917_,
		_w31919_,
		_w31920_
	);
	LUT2 #(
		.INIT('h1)
	) name27874 (
		_w31915_,
		_w31920_,
		_w31921_
	);
	LUT2 #(
		.INIT('h4)
	) name27875 (
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w31922_
	);
	LUT2 #(
		.INIT('h2)
	) name27876 (
		_w31908_,
		_w31910_,
		_w31923_
	);
	LUT2 #(
		.INIT('h4)
	) name27877 (
		_w31922_,
		_w31923_,
		_w31924_
	);
	LUT2 #(
		.INIT('h8)
	) name27878 (
		_w23418_,
		_w31924_,
		_w31925_
	);
	LUT2 #(
		.INIT('h4)
	) name27879 (
		_w31921_,
		_w31925_,
		_w31926_
	);
	LUT2 #(
		.INIT('h1)
	) name27880 (
		\clkc_Cnt4096_reg/NET0131 ,
		_w31909_,
		_w31927_
	);
	LUT2 #(
		.INIT('h4)
	) name27881 (
		_w31926_,
		_w31927_,
		_w31928_
	);
	LUT2 #(
		.INIT('h1)
	) name27882 (
		\clkc_Awake_reg/NET0131 ,
		_w31928_,
		_w31929_
	);
	LUT2 #(
		.INIT('h2)
	) name27883 (
		_w27915_,
		_w28054_,
		_w31930_
	);
	LUT2 #(
		.INIT('h2)
	) name27884 (
		\core_c_psq_CNTR_reg_DO_reg[13]/NET0131 ,
		_w27915_,
		_w31931_
	);
	LUT2 #(
		.INIT('h1)
	) name27885 (
		_w31930_,
		_w31931_,
		_w31932_
	);
	LUT2 #(
		.INIT('h2)
	) name27886 (
		\tm_tsr_reg_DO_reg[0]/NET0131 ,
		_w25491_,
		_w31933_
	);
	LUT2 #(
		.INIT('h8)
	) name27887 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TSR_TMP_reg[0]/NET0131 ,
		_w31934_
	);
	LUT2 #(
		.INIT('h1)
	) name27888 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		\tm_TSR_TMP_reg[0]/NET0131 ,
		_w31935_
	);
	LUT2 #(
		.INIT('h1)
	) name27889 (
		_w31934_,
		_w31935_,
		_w31936_
	);
	LUT2 #(
		.INIT('h2)
	) name27890 (
		_w25491_,
		_w31936_,
		_w31937_
	);
	LUT2 #(
		.INIT('h1)
	) name27891 (
		_w31933_,
		_w31937_,
		_w31938_
	);
	LUT2 #(
		.INIT('h2)
	) name27892 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 ,
		_w18266_,
		_w31939_
	);
	LUT2 #(
		.INIT('h1)
	) name27893 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[1]/P0001 ,
		_w18271_,
		_w31940_
	);
	LUT2 #(
		.INIT('h2)
	) name27894 (
		_w18271_,
		_w18974_,
		_w31941_
	);
	LUT2 #(
		.INIT('h2)
	) name27895 (
		_w18273_,
		_w31940_,
		_w31942_
	);
	LUT2 #(
		.INIT('h4)
	) name27896 (
		_w31941_,
		_w31942_,
		_w31943_
	);
	LUT2 #(
		.INIT('h1)
	) name27897 (
		_w18270_,
		_w31939_,
		_w31944_
	);
	LUT2 #(
		.INIT('h4)
	) name27898 (
		_w31943_,
		_w31944_,
		_w31945_
	);
	LUT2 #(
		.INIT('h1)
	) name27899 (
		_w18262_,
		_w31945_,
		_w31946_
	);
	LUT2 #(
		.INIT('h8)
	) name27900 (
		_w18262_,
		_w19667_,
		_w31947_
	);
	LUT2 #(
		.INIT('h1)
	) name27901 (
		_w31946_,
		_w31947_,
		_w31948_
	);
	LUT2 #(
		.INIT('h2)
	) name27902 (
		_w14752_,
		_w19667_,
		_w31949_
	);
	LUT2 #(
		.INIT('h8)
	) name27903 (
		_w18328_,
		_w18974_,
		_w31950_
	);
	LUT2 #(
		.INIT('h2)
	) name27904 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[1]/P0001 ,
		_w18330_,
		_w31951_
	);
	LUT2 #(
		.INIT('h2)
	) name27905 (
		_w18334_,
		_w31951_,
		_w31952_
	);
	LUT2 #(
		.INIT('h4)
	) name27906 (
		_w31950_,
		_w31952_,
		_w31953_
	);
	LUT2 #(
		.INIT('h1)
	) name27907 (
		_w31949_,
		_w31953_,
		_w31954_
	);
	LUT2 #(
		.INIT('h2)
	) name27908 (
		\core_eu_em_mac_em_reg_mfrwe_DO_reg[10]/P0001 ,
		_w20990_,
		_w31955_
	);
	LUT2 #(
		.INIT('h2)
	) name27909 (
		_w20990_,
		_w31482_,
		_w31956_
	);
	LUT2 #(
		.INIT('h1)
	) name27910 (
		_w31955_,
		_w31956_,
		_w31957_
	);
	LUT2 #(
		.INIT('h4)
	) name27911 (
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		\sport1_rxctl_ISRa_reg/P0001 ,
		_w31958_
	);
	LUT2 #(
		.INIT('h8)
	) name27912 (
		\core_dag_modulo1_R1wrap_reg/P0001 ,
		\sport1_regs_AUTOreg_DO_reg[0]/NET0131 ,
		_w31959_
	);
	LUT2 #(
		.INIT('h1)
	) name27913 (
		\core_c_psq_IFC_reg[9]/NET0131 ,
		_w31958_,
		_w31960_
	);
	LUT2 #(
		.INIT('h4)
	) name27914 (
		_w31959_,
		_w31960_,
		_w31961_
	);
	LUT2 #(
		.INIT('h2)
	) name27915 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w31961_,
		_w31962_
	);
	LUT2 #(
		.INIT('h1)
	) name27916 (
		\core_c_psq_Iflag_reg[1]/NET0131 ,
		_w31962_,
		_w31963_
	);
	LUT2 #(
		.INIT('h2)
	) name27917 (
		_w21416_,
		_w31963_,
		_w31964_
	);
	LUT2 #(
		.INIT('h4)
	) name27918 (
		\core_c_dec_MFDAG1_Ei_reg/NET0131 ,
		_w4117_,
		_w31965_
	);
	LUT2 #(
		.INIT('h4)
	) name27919 (
		_w30936_,
		_w31269_,
		_w31966_
	);
	LUT2 #(
		.INIT('h4)
	) name27920 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w31966_,
		_w31967_
	);
	LUT2 #(
		.INIT('h2)
	) name27921 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w31263_,
		_w31968_
	);
	LUT2 #(
		.INIT('h8)
	) name27922 (
		_w19270_,
		_w31968_,
		_w31969_
	);
	LUT2 #(
		.INIT('h8)
	) name27923 (
		_w31967_,
		_w31969_,
		_w31970_
	);
	LUT2 #(
		.INIT('h1)
	) name27924 (
		_w4117_,
		_w31970_,
		_w31971_
	);
	LUT2 #(
		.INIT('h1)
	) name27925 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w31263_,
		_w31972_
	);
	LUT2 #(
		.INIT('h8)
	) name27926 (
		_w31966_,
		_w31972_,
		_w31973_
	);
	LUT2 #(
		.INIT('h8)
	) name27927 (
		_w19298_,
		_w31968_,
		_w31974_
	);
	LUT2 #(
		.INIT('h8)
	) name27928 (
		_w31967_,
		_w31974_,
		_w31975_
	);
	LUT2 #(
		.INIT('h8)
	) name27929 (
		_w19267_,
		_w31968_,
		_w31976_
	);
	LUT2 #(
		.INIT('h8)
	) name27930 (
		_w31967_,
		_w31976_,
		_w31977_
	);
	LUT2 #(
		.INIT('h1)
	) name27931 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w31269_,
		_w31978_
	);
	LUT2 #(
		.INIT('h8)
	) name27932 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w31978_,
		_w31979_
	);
	LUT2 #(
		.INIT('h8)
	) name27933 (
		_w31654_,
		_w31979_,
		_w31980_
	);
	LUT2 #(
		.INIT('h8)
	) name27934 (
		_w19301_,
		_w31968_,
		_w31981_
	);
	LUT2 #(
		.INIT('h8)
	) name27935 (
		_w31967_,
		_w31981_,
		_w31982_
	);
	LUT2 #(
		.INIT('h1)
	) name27936 (
		_w31973_,
		_w31975_,
		_w31983_
	);
	LUT2 #(
		.INIT('h1)
	) name27937 (
		_w31977_,
		_w31980_,
		_w31984_
	);
	LUT2 #(
		.INIT('h4)
	) name27938 (
		_w31982_,
		_w31984_,
		_w31985_
	);
	LUT2 #(
		.INIT('h8)
	) name27939 (
		_w31971_,
		_w31983_,
		_w31986_
	);
	LUT2 #(
		.INIT('h8)
	) name27940 (
		_w31985_,
		_w31986_,
		_w31987_
	);
	LUT2 #(
		.INIT('h1)
	) name27941 (
		_w31965_,
		_w31987_,
		_w31988_
	);
	LUT2 #(
		.INIT('h8)
	) name27942 (
		\core_c_dec_Long_Eg_reg/P0001 ,
		_w4118_,
		_w31989_
	);
	LUT2 #(
		.INIT('h2)
	) name27943 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w30935_,
		_w31990_
	);
	LUT2 #(
		.INIT('h8)
	) name27944 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w30935_,
		_w31991_
	);
	LUT2 #(
		.INIT('h1)
	) name27945 (
		_w31990_,
		_w31991_,
		_w31992_
	);
	LUT2 #(
		.INIT('h2)
	) name27946 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w30935_,
		_w31993_
	);
	LUT2 #(
		.INIT('h8)
	) name27947 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w30935_,
		_w31994_
	);
	LUT2 #(
		.INIT('h1)
	) name27948 (
		_w31993_,
		_w31994_,
		_w31995_
	);
	LUT2 #(
		.INIT('h2)
	) name27949 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w30935_,
		_w31996_
	);
	LUT2 #(
		.INIT('h8)
	) name27950 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w30935_,
		_w31997_
	);
	LUT2 #(
		.INIT('h1)
	) name27951 (
		_w31996_,
		_w31997_,
		_w31998_
	);
	LUT2 #(
		.INIT('h1)
	) name27952 (
		_w31995_,
		_w31998_,
		_w31999_
	);
	LUT2 #(
		.INIT('h1)
	) name27953 (
		_w31090_,
		_w31262_,
		_w32000_
	);
	LUT2 #(
		.INIT('h4)
	) name27954 (
		_w30935_,
		_w31083_,
		_w32001_
	);
	LUT2 #(
		.INIT('h1)
	) name27955 (
		_w32000_,
		_w32001_,
		_w32002_
	);
	LUT2 #(
		.INIT('h1)
	) name27956 (
		_w31091_,
		_w31268_,
		_w32003_
	);
	LUT2 #(
		.INIT('h2)
	) name27957 (
		_w32002_,
		_w32003_,
		_w32004_
	);
	LUT2 #(
		.INIT('h2)
	) name27958 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w30935_,
		_w32005_
	);
	LUT2 #(
		.INIT('h8)
	) name27959 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w30935_,
		_w32006_
	);
	LUT2 #(
		.INIT('h1)
	) name27960 (
		_w32005_,
		_w32006_,
		_w32007_
	);
	LUT2 #(
		.INIT('h2)
	) name27961 (
		_w32004_,
		_w32007_,
		_w32008_
	);
	LUT2 #(
		.INIT('h4)
	) name27962 (
		_w31992_,
		_w31999_,
		_w32009_
	);
	LUT2 #(
		.INIT('h8)
	) name27963 (
		_w32008_,
		_w32009_,
		_w32010_
	);
	LUT2 #(
		.INIT('h1)
	) name27964 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w32011_
	);
	LUT2 #(
		.INIT('h4)
	) name27965 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w32011_,
		_w32012_
	);
	LUT2 #(
		.INIT('h2)
	) name27966 (
		_w24815_,
		_w32012_,
		_w32013_
	);
	LUT2 #(
		.INIT('h8)
	) name27967 (
		_w31995_,
		_w31998_,
		_w32014_
	);
	LUT2 #(
		.INIT('h8)
	) name27968 (
		_w32007_,
		_w32014_,
		_w32015_
	);
	LUT2 #(
		.INIT('h8)
	) name27969 (
		_w31992_,
		_w32004_,
		_w32016_
	);
	LUT2 #(
		.INIT('h8)
	) name27970 (
		_w32015_,
		_w32016_,
		_w32017_
	);
	LUT2 #(
		.INIT('h4)
	) name27971 (
		_w31992_,
		_w32002_,
		_w32018_
	);
	LUT2 #(
		.INIT('h8)
	) name27972 (
		_w32003_,
		_w32018_,
		_w32019_
	);
	LUT2 #(
		.INIT('h8)
	) name27973 (
		_w31999_,
		_w32019_,
		_w32020_
	);
	LUT2 #(
		.INIT('h8)
	) name27974 (
		_w31992_,
		_w31995_,
		_w32021_
	);
	LUT2 #(
		.INIT('h8)
	) name27975 (
		_w32008_,
		_w32021_,
		_w32022_
	);
	LUT2 #(
		.INIT('h2)
	) name27976 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w31269_,
		_w32023_
	);
	LUT2 #(
		.INIT('h8)
	) name27977 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w32023_,
		_w32024_
	);
	LUT2 #(
		.INIT('h8)
	) name27978 (
		_w31654_,
		_w32024_,
		_w32025_
	);
	LUT2 #(
		.INIT('h1)
	) name27979 (
		_w21250_,
		_w25249_,
		_w32026_
	);
	LUT2 #(
		.INIT('h4)
	) name27980 (
		_w32013_,
		_w32026_,
		_w32027_
	);
	LUT2 #(
		.INIT('h4)
	) name27981 (
		_w32025_,
		_w32027_,
		_w32028_
	);
	LUT2 #(
		.INIT('h4)
	) name27982 (
		_w32010_,
		_w32028_,
		_w32029_
	);
	LUT2 #(
		.INIT('h1)
	) name27983 (
		_w32017_,
		_w32020_,
		_w32030_
	);
	LUT2 #(
		.INIT('h4)
	) name27984 (
		_w32022_,
		_w32030_,
		_w32031_
	);
	LUT2 #(
		.INIT('h8)
	) name27985 (
		_w32029_,
		_w32031_,
		_w32032_
	);
	LUT2 #(
		.INIT('h2)
	) name27986 (
		_w23231_,
		_w32032_,
		_w32033_
	);
	LUT2 #(
		.INIT('h1)
	) name27987 (
		_w31989_,
		_w32033_,
		_w32034_
	);
	LUT2 #(
		.INIT('h8)
	) name27988 (
		\sice_ICYC_reg[23]/NET0131 ,
		_w20785_,
		_w32035_
	);
	LUT2 #(
		.INIT('h1)
	) name27989 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w32035_,
		_w32036_
	);
	LUT2 #(
		.INIT('h1)
	) name27990 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		_w4093_,
		_w32037_
	);
	LUT2 #(
		.INIT('h8)
	) name27991 (
		_w32036_,
		_w32037_,
		_w32038_
	);
	LUT2 #(
		.INIT('h8)
	) name27992 (
		_w22584_,
		_w32038_,
		_w32039_
	);
	LUT2 #(
		.INIT('h8)
	) name27993 (
		\sice_IIRC_reg[18]/NET0131 ,
		_w32039_,
		_w32040_
	);
	LUT2 #(
		.INIT('h8)
	) name27994 (
		\sice_IIRC_reg[19]/NET0131 ,
		_w32040_,
		_w32041_
	);
	LUT2 #(
		.INIT('h8)
	) name27995 (
		\sice_IIRC_reg[20]/NET0131 ,
		_w32041_,
		_w32042_
	);
	LUT2 #(
		.INIT('h1)
	) name27996 (
		\sice_IIRC_reg[20]/NET0131 ,
		_w32041_,
		_w32043_
	);
	LUT2 #(
		.INIT('h1)
	) name27997 (
		_w32042_,
		_w32043_,
		_w32044_
	);
	LUT2 #(
		.INIT('h2)
	) name27998 (
		_w6111_,
		_w6164_,
		_w32045_
	);
	LUT2 #(
		.INIT('h4)
	) name27999 (
		_w6121_,
		_w32045_,
		_w32046_
	);
	LUT2 #(
		.INIT('h4)
	) name28000 (
		_w6047_,
		_w32046_,
		_w32047_
	);
	LUT2 #(
		.INIT('h1)
	) name28001 (
		_w6112_,
		_w32047_,
		_w32048_
	);
	LUT2 #(
		.INIT('h8)
	) name28002 (
		_w6546_,
		_w32048_,
		_w32049_
	);
	LUT2 #(
		.INIT('h4)
	) name28003 (
		_w6101_,
		_w6121_,
		_w32050_
	);
	LUT2 #(
		.INIT('h1)
	) name28004 (
		_w6111_,
		_w32050_,
		_w32051_
	);
	LUT2 #(
		.INIT('h4)
	) name28005 (
		_w6047_,
		_w6165_,
		_w32052_
	);
	LUT2 #(
		.INIT('h2)
	) name28006 (
		_w6111_,
		_w32052_,
		_w32053_
	);
	LUT2 #(
		.INIT('h1)
	) name28007 (
		_w32051_,
		_w32053_,
		_w32054_
	);
	LUT2 #(
		.INIT('h2)
	) name28008 (
		_w7622_,
		_w32048_,
		_w32055_
	);
	LUT2 #(
		.INIT('h4)
	) name28009 (
		_w32049_,
		_w32054_,
		_w32056_
	);
	LUT2 #(
		.INIT('h4)
	) name28010 (
		_w32055_,
		_w32056_,
		_w32057_
	);
	LUT2 #(
		.INIT('h2)
	) name28011 (
		_w6047_,
		_w6121_,
		_w32058_
	);
	LUT2 #(
		.INIT('h4)
	) name28012 (
		_w9452_,
		_w32058_,
		_w32059_
	);
	LUT2 #(
		.INIT('h4)
	) name28013 (
		_w9445_,
		_w32048_,
		_w32060_
	);
	LUT2 #(
		.INIT('h4)
	) name28014 (
		_w32059_,
		_w32060_,
		_w32061_
	);
	LUT2 #(
		.INIT('h2)
	) name28015 (
		_w9497_,
		_w32048_,
		_w32062_
	);
	LUT2 #(
		.INIT('h1)
	) name28016 (
		_w32054_,
		_w32061_,
		_w32063_
	);
	LUT2 #(
		.INIT('h4)
	) name28017 (
		_w32062_,
		_w32063_,
		_w32064_
	);
	LUT2 #(
		.INIT('h1)
	) name28018 (
		_w32057_,
		_w32064_,
		_w32065_
	);
	LUT2 #(
		.INIT('h1)
	) name28019 (
		_w6106_,
		_w6111_,
		_w32066_
	);
	LUT2 #(
		.INIT('h4)
	) name28020 (
		_w6101_,
		_w32066_,
		_w32067_
	);
	LUT2 #(
		.INIT('h1)
	) name28021 (
		_w32053_,
		_w32067_,
		_w32068_
	);
	LUT2 #(
		.INIT('h1)
	) name28022 (
		_w32065_,
		_w32068_,
		_w32069_
	);
	LUT2 #(
		.INIT('h1)
	) name28023 (
		_w7607_,
		_w32048_,
		_w32070_
	);
	LUT2 #(
		.INIT('h4)
	) name28024 (
		_w7340_,
		_w32048_,
		_w32071_
	);
	LUT2 #(
		.INIT('h2)
	) name28025 (
		_w32054_,
		_w32070_,
		_w32072_
	);
	LUT2 #(
		.INIT('h4)
	) name28026 (
		_w32071_,
		_w32072_,
		_w32073_
	);
	LUT2 #(
		.INIT('h8)
	) name28027 (
		_w6158_,
		_w32048_,
		_w32074_
	);
	LUT2 #(
		.INIT('h2)
	) name28028 (
		_w6951_,
		_w32048_,
		_w32075_
	);
	LUT2 #(
		.INIT('h1)
	) name28029 (
		_w32054_,
		_w32074_,
		_w32076_
	);
	LUT2 #(
		.INIT('h4)
	) name28030 (
		_w32075_,
		_w32076_,
		_w32077_
	);
	LUT2 #(
		.INIT('h1)
	) name28031 (
		_w32073_,
		_w32077_,
		_w32078_
	);
	LUT2 #(
		.INIT('h2)
	) name28032 (
		_w32068_,
		_w32078_,
		_w32079_
	);
	LUT2 #(
		.INIT('h1)
	) name28033 (
		_w32069_,
		_w32079_,
		_w32080_
	);
	LUT2 #(
		.INIT('h2)
	) name28034 (
		\core_c_psq_DMOVL_reg_DO_reg[3]/NET0131 ,
		_w25009_,
		_w32081_
	);
	LUT2 #(
		.INIT('h8)
	) name28035 (
		_w32080_,
		_w32081_,
		_w32082_
	);
	LUT2 #(
		.INIT('h4)
	) name28036 (
		PM_bdry_sel_pad,
		_w20698_,
		_w32083_
	);
	LUT2 #(
		.INIT('h2)
	) name28037 (
		\core_c_psq_PMOVL_regh_DO_reg[3]/NET0131 ,
		_w19702_,
		_w32084_
	);
	LUT2 #(
		.INIT('h4)
	) name28038 (
		_w20687_,
		_w32084_,
		_w32085_
	);
	LUT2 #(
		.INIT('h4)
	) name28039 (
		_w32083_,
		_w32085_,
		_w32086_
	);
	LUT2 #(
		.INIT('h1)
	) name28040 (
		_w25081_,
		_w32086_,
		_w32087_
	);
	LUT2 #(
		.INIT('h4)
	) name28041 (
		_w32082_,
		_w32087_,
		_w32088_
	);
	LUT2 #(
		.INIT('h2)
	) name28042 (
		_w11741_,
		_w32088_,
		_w32089_
	);
	LUT2 #(
		.INIT('h1)
	) name28043 (
		\T_TMODE[1]_pad ,
		_w4117_,
		_w32090_
	);
	LUT2 #(
		.INIT('h4)
	) name28044 (
		_w32089_,
		_w32090_,
		_w32091_
	);
	LUT2 #(
		.INIT('h8)
	) name28045 (
		_w4068_,
		_w4117_,
		_w32092_
	);
	LUT2 #(
		.INIT('h1)
	) name28046 (
		_w32091_,
		_w32092_,
		_w32093_
	);
	LUT2 #(
		.INIT('h8)
	) name28047 (
		_w10638_,
		_w31339_,
		_w32094_
	);
	LUT2 #(
		.INIT('h8)
	) name28048 (
		\core_dag_ilm2reg_M5_we_DO_reg[8]/NET0131 ,
		_w31341_,
		_w32095_
	);
	LUT2 #(
		.INIT('h8)
	) name28049 (
		\core_dag_ilm2reg_M6_we_DO_reg[8]/NET0131 ,
		_w31331_,
		_w32096_
	);
	LUT2 #(
		.INIT('h8)
	) name28050 (
		\core_dag_ilm2reg_M4_we_DO_reg[8]/NET0131 ,
		_w31344_,
		_w32097_
	);
	LUT2 #(
		.INIT('h8)
	) name28051 (
		\core_dag_ilm2reg_M7_we_DO_reg[8]/NET0131 ,
		_w31337_,
		_w32098_
	);
	LUT2 #(
		.INIT('h1)
	) name28052 (
		_w32096_,
		_w32098_,
		_w32099_
	);
	LUT2 #(
		.INIT('h4)
	) name28053 (
		_w21579_,
		_w32099_,
		_w32100_
	);
	LUT2 #(
		.INIT('h1)
	) name28054 (
		_w32095_,
		_w32097_,
		_w32101_
	);
	LUT2 #(
		.INIT('h8)
	) name28055 (
		_w32100_,
		_w32101_,
		_w32102_
	);
	LUT2 #(
		.INIT('h4)
	) name28056 (
		_w32094_,
		_w32102_,
		_w32103_
	);
	LUT2 #(
		.INIT('h4)
	) name28057 (
		\core_dag_ilm2reg_M_reg[8]/NET0131 ,
		_w21579_,
		_w32104_
	);
	LUT2 #(
		.INIT('h1)
	) name28058 (
		_w32103_,
		_w32104_,
		_w32105_
	);
	LUT2 #(
		.INIT('h8)
	) name28059 (
		_w7340_,
		_w31339_,
		_w32106_
	);
	LUT2 #(
		.INIT('h8)
	) name28060 (
		\core_dag_ilm2reg_M4_we_DO_reg[13]/NET0131 ,
		_w31344_,
		_w32107_
	);
	LUT2 #(
		.INIT('h8)
	) name28061 (
		\core_dag_ilm2reg_M7_we_DO_reg[13]/NET0131 ,
		_w31337_,
		_w32108_
	);
	LUT2 #(
		.INIT('h8)
	) name28062 (
		\core_dag_ilm2reg_M5_we_DO_reg[13]/NET0131 ,
		_w31341_,
		_w32109_
	);
	LUT2 #(
		.INIT('h8)
	) name28063 (
		\core_dag_ilm2reg_M6_we_DO_reg[13]/NET0131 ,
		_w31331_,
		_w32110_
	);
	LUT2 #(
		.INIT('h1)
	) name28064 (
		_w32108_,
		_w32110_,
		_w32111_
	);
	LUT2 #(
		.INIT('h4)
	) name28065 (
		_w21579_,
		_w32111_,
		_w32112_
	);
	LUT2 #(
		.INIT('h1)
	) name28066 (
		_w32107_,
		_w32109_,
		_w32113_
	);
	LUT2 #(
		.INIT('h8)
	) name28067 (
		_w32112_,
		_w32113_,
		_w32114_
	);
	LUT2 #(
		.INIT('h4)
	) name28068 (
		_w32106_,
		_w32114_,
		_w32115_
	);
	LUT2 #(
		.INIT('h4)
	) name28069 (
		\core_dag_ilm2reg_M_reg[13]/NET0131 ,
		_w21579_,
		_w32116_
	);
	LUT2 #(
		.INIT('h1)
	) name28070 (
		_w32115_,
		_w32116_,
		_w32117_
	);
	LUT2 #(
		.INIT('h8)
	) name28071 (
		_w9178_,
		_w31409_,
		_w32118_
	);
	LUT2 #(
		.INIT('h8)
	) name28072 (
		\core_dag_ilm1reg_M1_we_DO_reg[12]/NET0131 ,
		_w31414_,
		_w32119_
	);
	LUT2 #(
		.INIT('h8)
	) name28073 (
		\core_dag_ilm1reg_M3_we_DO_reg[12]/NET0131 ,
		_w31407_,
		_w32120_
	);
	LUT2 #(
		.INIT('h8)
	) name28074 (
		\core_dag_ilm1reg_M0_we_DO_reg[12]/NET0131 ,
		_w31411_,
		_w32121_
	);
	LUT2 #(
		.INIT('h8)
	) name28075 (
		\core_dag_ilm1reg_M2_we_DO_reg[12]/NET0131 ,
		_w31401_,
		_w32122_
	);
	LUT2 #(
		.INIT('h1)
	) name28076 (
		_w32120_,
		_w32122_,
		_w32123_
	);
	LUT2 #(
		.INIT('h4)
	) name28077 (
		_w21592_,
		_w32123_,
		_w32124_
	);
	LUT2 #(
		.INIT('h1)
	) name28078 (
		_w32119_,
		_w32121_,
		_w32125_
	);
	LUT2 #(
		.INIT('h8)
	) name28079 (
		_w32124_,
		_w32125_,
		_w32126_
	);
	LUT2 #(
		.INIT('h4)
	) name28080 (
		_w32118_,
		_w32126_,
		_w32127_
	);
	LUT2 #(
		.INIT('h4)
	) name28081 (
		\core_dag_ilm1reg_M_reg[12]/NET0131 ,
		_w21592_,
		_w32128_
	);
	LUT2 #(
		.INIT('h1)
	) name28082 (
		_w32127_,
		_w32128_,
		_w32129_
	);
	LUT2 #(
		.INIT('h8)
	) name28083 (
		_w11265_,
		_w31339_,
		_w32130_
	);
	LUT2 #(
		.INIT('h8)
	) name28084 (
		\core_dag_ilm2reg_M4_we_DO_reg[7]/NET0131 ,
		_w31344_,
		_w32131_
	);
	LUT2 #(
		.INIT('h8)
	) name28085 (
		\core_dag_ilm2reg_M7_we_DO_reg[7]/NET0131 ,
		_w31337_,
		_w32132_
	);
	LUT2 #(
		.INIT('h8)
	) name28086 (
		\core_dag_ilm2reg_M5_we_DO_reg[7]/NET0131 ,
		_w31341_,
		_w32133_
	);
	LUT2 #(
		.INIT('h8)
	) name28087 (
		\core_dag_ilm2reg_M6_we_DO_reg[7]/NET0131 ,
		_w31331_,
		_w32134_
	);
	LUT2 #(
		.INIT('h1)
	) name28088 (
		_w32132_,
		_w32134_,
		_w32135_
	);
	LUT2 #(
		.INIT('h4)
	) name28089 (
		_w21579_,
		_w32135_,
		_w32136_
	);
	LUT2 #(
		.INIT('h1)
	) name28090 (
		_w32131_,
		_w32133_,
		_w32137_
	);
	LUT2 #(
		.INIT('h8)
	) name28091 (
		_w32136_,
		_w32137_,
		_w32138_
	);
	LUT2 #(
		.INIT('h4)
	) name28092 (
		_w32130_,
		_w32138_,
		_w32139_
	);
	LUT2 #(
		.INIT('h4)
	) name28093 (
		\core_dag_ilm2reg_M_reg[7]/NET0131 ,
		_w21579_,
		_w32140_
	);
	LUT2 #(
		.INIT('h1)
	) name28094 (
		_w32139_,
		_w32140_,
		_w32141_
	);
	LUT2 #(
		.INIT('h8)
	) name28095 (
		_w7607_,
		_w31339_,
		_w32142_
	);
	LUT2 #(
		.INIT('h8)
	) name28096 (
		\core_dag_ilm2reg_M4_we_DO_reg[0]/NET0131 ,
		_w31344_,
		_w32143_
	);
	LUT2 #(
		.INIT('h8)
	) name28097 (
		\core_dag_ilm2reg_M7_we_DO_reg[0]/NET0131 ,
		_w31337_,
		_w32144_
	);
	LUT2 #(
		.INIT('h8)
	) name28098 (
		\core_dag_ilm2reg_M5_we_DO_reg[0]/NET0131 ,
		_w31341_,
		_w32145_
	);
	LUT2 #(
		.INIT('h8)
	) name28099 (
		\core_dag_ilm2reg_M6_we_DO_reg[0]/NET0131 ,
		_w31331_,
		_w32146_
	);
	LUT2 #(
		.INIT('h1)
	) name28100 (
		_w32144_,
		_w32146_,
		_w32147_
	);
	LUT2 #(
		.INIT('h4)
	) name28101 (
		_w21579_,
		_w32147_,
		_w32148_
	);
	LUT2 #(
		.INIT('h1)
	) name28102 (
		_w32143_,
		_w32145_,
		_w32149_
	);
	LUT2 #(
		.INIT('h8)
	) name28103 (
		_w32148_,
		_w32149_,
		_w32150_
	);
	LUT2 #(
		.INIT('h4)
	) name28104 (
		_w32142_,
		_w32150_,
		_w32151_
	);
	LUT2 #(
		.INIT('h4)
	) name28105 (
		\core_dag_ilm2reg_M_reg[0]/NET0131 ,
		_w21579_,
		_w32152_
	);
	LUT2 #(
		.INIT('h1)
	) name28106 (
		_w32151_,
		_w32152_,
		_w32153_
	);
	LUT2 #(
		.INIT('h8)
	) name28107 (
		_w11265_,
		_w31409_,
		_w32154_
	);
	LUT2 #(
		.INIT('h8)
	) name28108 (
		\core_dag_ilm1reg_M1_we_DO_reg[7]/NET0131 ,
		_w31414_,
		_w32155_
	);
	LUT2 #(
		.INIT('h8)
	) name28109 (
		\core_dag_ilm1reg_M3_we_DO_reg[7]/NET0131 ,
		_w31407_,
		_w32156_
	);
	LUT2 #(
		.INIT('h8)
	) name28110 (
		\core_dag_ilm1reg_M0_we_DO_reg[7]/NET0131 ,
		_w31411_,
		_w32157_
	);
	LUT2 #(
		.INIT('h8)
	) name28111 (
		\core_dag_ilm1reg_M2_we_DO_reg[7]/NET0131 ,
		_w31401_,
		_w32158_
	);
	LUT2 #(
		.INIT('h1)
	) name28112 (
		_w32156_,
		_w32158_,
		_w32159_
	);
	LUT2 #(
		.INIT('h4)
	) name28113 (
		_w21592_,
		_w32159_,
		_w32160_
	);
	LUT2 #(
		.INIT('h1)
	) name28114 (
		_w32155_,
		_w32157_,
		_w32161_
	);
	LUT2 #(
		.INIT('h8)
	) name28115 (
		_w32160_,
		_w32161_,
		_w32162_
	);
	LUT2 #(
		.INIT('h4)
	) name28116 (
		_w32154_,
		_w32162_,
		_w32163_
	);
	LUT2 #(
		.INIT('h4)
	) name28117 (
		\core_dag_ilm1reg_M_reg[7]/NET0131 ,
		_w21592_,
		_w32164_
	);
	LUT2 #(
		.INIT('h1)
	) name28118 (
		_w32163_,
		_w32164_,
		_w32165_
	);
	LUT2 #(
		.INIT('h8)
	) name28119 (
		_w8113_,
		_w31409_,
		_w32166_
	);
	LUT2 #(
		.INIT('h8)
	) name28120 (
		\core_dag_ilm1reg_M0_we_DO_reg[3]/NET0131 ,
		_w31411_,
		_w32167_
	);
	LUT2 #(
		.INIT('h8)
	) name28121 (
		\core_dag_ilm1reg_M2_we_DO_reg[3]/NET0131 ,
		_w31401_,
		_w32168_
	);
	LUT2 #(
		.INIT('h8)
	) name28122 (
		\core_dag_ilm1reg_M1_we_DO_reg[3]/NET0131 ,
		_w31414_,
		_w32169_
	);
	LUT2 #(
		.INIT('h8)
	) name28123 (
		\core_dag_ilm1reg_M3_we_DO_reg[3]/NET0131 ,
		_w31407_,
		_w32170_
	);
	LUT2 #(
		.INIT('h1)
	) name28124 (
		_w32168_,
		_w32170_,
		_w32171_
	);
	LUT2 #(
		.INIT('h4)
	) name28125 (
		_w21592_,
		_w32171_,
		_w32172_
	);
	LUT2 #(
		.INIT('h1)
	) name28126 (
		_w32167_,
		_w32169_,
		_w32173_
	);
	LUT2 #(
		.INIT('h8)
	) name28127 (
		_w32172_,
		_w32173_,
		_w32174_
	);
	LUT2 #(
		.INIT('h4)
	) name28128 (
		_w32166_,
		_w32174_,
		_w32175_
	);
	LUT2 #(
		.INIT('h4)
	) name28129 (
		\core_dag_ilm1reg_M_reg[3]/NET0131 ,
		_w21592_,
		_w32176_
	);
	LUT2 #(
		.INIT('h1)
	) name28130 (
		_w32175_,
		_w32176_,
		_w32177_
	);
	LUT2 #(
		.INIT('h8)
	) name28131 (
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w28786_,
		_w32178_
	);
	LUT2 #(
		.INIT('h1)
	) name28132 (
		\sport1_cfg_FSi_cnt_reg[4]/NET0131 ,
		_w28859_,
		_w32179_
	);
	LUT2 #(
		.INIT('h1)
	) name28133 (
		_w28860_,
		_w32179_,
		_w32180_
	);
	LUT2 #(
		.INIT('h8)
	) name28134 (
		_w28855_,
		_w32180_,
		_w32181_
	);
	LUT2 #(
		.INIT('h1)
	) name28135 (
		_w32178_,
		_w32181_,
		_w32182_
	);
	LUT2 #(
		.INIT('h8)
	) name28136 (
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w28876_,
		_w32183_
	);
	LUT2 #(
		.INIT('h1)
	) name28137 (
		\sport0_cfg_FSi_cnt_reg[4]/NET0131 ,
		_w28949_,
		_w32184_
	);
	LUT2 #(
		.INIT('h1)
	) name28138 (
		_w28950_,
		_w32184_,
		_w32185_
	);
	LUT2 #(
		.INIT('h8)
	) name28139 (
		_w28945_,
		_w32185_,
		_w32186_
	);
	LUT2 #(
		.INIT('h1)
	) name28140 (
		_w32183_,
		_w32186_,
		_w32187_
	);
	LUT2 #(
		.INIT('h8)
	) name28141 (
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w28786_,
		_w32188_
	);
	LUT2 #(
		.INIT('h1)
	) name28142 (
		\sport1_cfg_FSi_cnt_reg[6]/NET0131 ,
		_w28861_,
		_w32189_
	);
	LUT2 #(
		.INIT('h1)
	) name28143 (
		_w28862_,
		_w32189_,
		_w32190_
	);
	LUT2 #(
		.INIT('h8)
	) name28144 (
		_w28855_,
		_w32190_,
		_w32191_
	);
	LUT2 #(
		.INIT('h1)
	) name28145 (
		_w32188_,
		_w32191_,
		_w32192_
	);
	LUT2 #(
		.INIT('h8)
	) name28146 (
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w28876_,
		_w32193_
	);
	LUT2 #(
		.INIT('h1)
	) name28147 (
		\sport0_cfg_FSi_cnt_reg[6]/NET0131 ,
		_w28951_,
		_w32194_
	);
	LUT2 #(
		.INIT('h1)
	) name28148 (
		_w28952_,
		_w32194_,
		_w32195_
	);
	LUT2 #(
		.INIT('h8)
	) name28149 (
		_w28945_,
		_w32195_,
		_w32196_
	);
	LUT2 #(
		.INIT('h1)
	) name28150 (
		_w32193_,
		_w32196_,
		_w32197_
	);
	LUT2 #(
		.INIT('h2)
	) name28151 (
		\tm_tsr_reg_DO_reg[1]/NET0131 ,
		_w25491_,
		_w32198_
	);
	LUT2 #(
		.INIT('h4)
	) name28152 (
		\tm_TSR_TMP_reg[1]/NET0131 ,
		_w31935_,
		_w32199_
	);
	LUT2 #(
		.INIT('h2)
	) name28153 (
		\tm_TSR_TMP_reg[1]/NET0131 ,
		_w31935_,
		_w32200_
	);
	LUT2 #(
		.INIT('h1)
	) name28154 (
		_w32199_,
		_w32200_,
		_w32201_
	);
	LUT2 #(
		.INIT('h2)
	) name28155 (
		_w25491_,
		_w32201_,
		_w32202_
	);
	LUT2 #(
		.INIT('h1)
	) name28156 (
		_w32198_,
		_w32202_,
		_w32203_
	);
	LUT2 #(
		.INIT('h2)
	) name28157 (
		\tm_tsr_reg_DO_reg[2]/NET0131 ,
		_w25491_,
		_w32204_
	);
	LUT2 #(
		.INIT('h2)
	) name28158 (
		\tm_TSR_TMP_reg[2]/NET0131 ,
		_w32199_,
		_w32205_
	);
	LUT2 #(
		.INIT('h8)
	) name28159 (
		_w22402_,
		_w31935_,
		_w32206_
	);
	LUT2 #(
		.INIT('h1)
	) name28160 (
		_w32205_,
		_w32206_,
		_w32207_
	);
	LUT2 #(
		.INIT('h2)
	) name28161 (
		_w25491_,
		_w32207_,
		_w32208_
	);
	LUT2 #(
		.INIT('h1)
	) name28162 (
		_w32204_,
		_w32208_,
		_w32209_
	);
	LUT2 #(
		.INIT('h2)
	) name28163 (
		\tm_TSR_TMP_reg[3]/NET0131 ,
		_w32206_,
		_w32210_
	);
	LUT2 #(
		.INIT('h4)
	) name28164 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w22404_,
		_w32211_
	);
	LUT2 #(
		.INIT('h1)
	) name28165 (
		_w32210_,
		_w32211_,
		_w32212_
	);
	LUT2 #(
		.INIT('h2)
	) name28166 (
		_w25491_,
		_w32212_,
		_w32213_
	);
	LUT2 #(
		.INIT('h2)
	) name28167 (
		\tm_tsr_reg_DO_reg[3]/NET0131 ,
		_w25491_,
		_w32214_
	);
	LUT2 #(
		.INIT('h1)
	) name28168 (
		_w32213_,
		_w32214_,
		_w32215_
	);
	LUT2 #(
		.INIT('h4)
	) name28169 (
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		\sport1_txctl_c_sync1_reg/P0001 ,
		_w32216_
	);
	LUT2 #(
		.INIT('h4)
	) name28170 (
		\sport1_txctl_c_sync2_reg/P0001 ,
		_w32216_,
		_w32217_
	);
	LUT2 #(
		.INIT('h8)
	) name28171 (
		\core_dag_modulo1_T1wrap_reg/P0001 ,
		\sport1_regs_AUTOreg_DO_reg[1]/NET0131 ,
		_w32218_
	);
	LUT2 #(
		.INIT('h1)
	) name28172 (
		\core_c_psq_IFC_reg[10]/NET0131 ,
		_w32218_,
		_w32219_
	);
	LUT2 #(
		.INIT('h4)
	) name28173 (
		_w32217_,
		_w32219_,
		_w32220_
	);
	LUT2 #(
		.INIT('h2)
	) name28174 (
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w32220_,
		_w32221_
	);
	LUT2 #(
		.INIT('h1)
	) name28175 (
		\core_c_psq_Iflag_reg[2]/NET0131 ,
		_w32221_,
		_w32222_
	);
	LUT2 #(
		.INIT('h2)
	) name28176 (
		_w21406_,
		_w32222_,
		_w32223_
	);
	LUT2 #(
		.INIT('h8)
	) name28177 (
		_w19203_,
		_w23586_,
		_w32224_
	);
	LUT2 #(
		.INIT('h2)
	) name28178 (
		_w19202_,
		_w32224_,
		_w32225_
	);
	LUT2 #(
		.INIT('h4)
	) name28179 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w32225_,
		_w32226_
	);
	LUT2 #(
		.INIT('h8)
	) name28180 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w11265_,
		_w32227_
	);
	LUT2 #(
		.INIT('h8)
	) name28181 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][7]/P0001 ,
		_w14708_,
		_w32228_
	);
	LUT2 #(
		.INIT('h8)
	) name28182 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001 ,
		_w14699_,
		_w32229_
	);
	LUT2 #(
		.INIT('h8)
	) name28183 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001 ,
		_w14711_,
		_w32230_
	);
	LUT2 #(
		.INIT('h8)
	) name28184 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001 ,
		_w14704_,
		_w32231_
	);
	LUT2 #(
		.INIT('h8)
	) name28185 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001 ,
		_w14706_,
		_w32232_
	);
	LUT2 #(
		.INIT('h8)
	) name28186 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][7]/P0001 ,
		_w14702_,
		_w32233_
	);
	LUT2 #(
		.INIT('h8)
	) name28187 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][7]/P0001 ,
		_w14713_,
		_w32234_
	);
	LUT2 #(
		.INIT('h1)
	) name28188 (
		_w32228_,
		_w32229_,
		_w32235_
	);
	LUT2 #(
		.INIT('h1)
	) name28189 (
		_w32230_,
		_w32231_,
		_w32236_
	);
	LUT2 #(
		.INIT('h1)
	) name28190 (
		_w32232_,
		_w32233_,
		_w32237_
	);
	LUT2 #(
		.INIT('h4)
	) name28191 (
		_w32234_,
		_w32237_,
		_w32238_
	);
	LUT2 #(
		.INIT('h8)
	) name28192 (
		_w32235_,
		_w32236_,
		_w32239_
	);
	LUT2 #(
		.INIT('h8)
	) name28193 (
		_w32238_,
		_w32239_,
		_w32240_
	);
	LUT2 #(
		.INIT('h2)
	) name28194 (
		_w14697_,
		_w32240_,
		_w32241_
	);
	LUT2 #(
		.INIT('h4)
	) name28195 (
		_w17938_,
		_w23664_,
		_w32242_
	);
	LUT2 #(
		.INIT('h2)
	) name28196 (
		_w17938_,
		_w23664_,
		_w32243_
	);
	LUT2 #(
		.INIT('h2)
	) name28197 (
		_w23586_,
		_w32242_,
		_w32244_
	);
	LUT2 #(
		.INIT('h4)
	) name28198 (
		_w32243_,
		_w32244_,
		_w32245_
	);
	LUT2 #(
		.INIT('h8)
	) name28199 (
		_w13803_,
		_w32245_,
		_w32246_
	);
	LUT2 #(
		.INIT('h1)
	) name28200 (
		_w32227_,
		_w32246_,
		_w32247_
	);
	LUT2 #(
		.INIT('h4)
	) name28201 (
		_w32241_,
		_w32247_,
		_w32248_
	);
	LUT2 #(
		.INIT('h4)
	) name28202 (
		_w32225_,
		_w32248_,
		_w32249_
	);
	LUT2 #(
		.INIT('h2)
	) name28203 (
		_w4150_,
		_w32226_,
		_w32250_
	);
	LUT2 #(
		.INIT('h4)
	) name28204 (
		_w32249_,
		_w32250_,
		_w32251_
	);
	LUT2 #(
		.INIT('h4)
	) name28205 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w19205_,
		_w32252_
	);
	LUT2 #(
		.INIT('h4)
	) name28206 (
		_w19205_,
		_w19263_,
		_w32253_
	);
	LUT2 #(
		.INIT('h2)
	) name28207 (
		_w4150_,
		_w32252_,
		_w32254_
	);
	LUT2 #(
		.INIT('h4)
	) name28208 (
		_w32253_,
		_w32254_,
		_w32255_
	);
	LUT2 #(
		.INIT('h1)
	) name28209 (
		\sport0_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		_w19549_,
		_w32256_
	);
	LUT2 #(
		.INIT('h2)
	) name28210 (
		_w19197_,
		_w19550_,
		_w32257_
	);
	LUT2 #(
		.INIT('h4)
	) name28211 (
		_w32256_,
		_w32257_,
		_w32258_
	);
	LUT2 #(
		.INIT('h1)
	) name28212 (
		\sport0_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		_w19547_,
		_w32259_
	);
	LUT2 #(
		.INIT('h2)
	) name28213 (
		_w19197_,
		_w19548_,
		_w32260_
	);
	LUT2 #(
		.INIT('h4)
	) name28214 (
		_w32259_,
		_w32260_,
		_w32261_
	);
	LUT2 #(
		.INIT('h2)
	) name28215 (
		\sport1_rxctl_LMcnt_reg[2]/NET0131 ,
		_w30751_,
		_w32262_
	);
	LUT2 #(
		.INIT('h1)
	) name28216 (
		_w30752_,
		_w32262_,
		_w32263_
	);
	LUT2 #(
		.INIT('h4)
	) name28217 (
		_w30754_,
		_w31705_,
		_w32264_
	);
	LUT2 #(
		.INIT('h4)
	) name28218 (
		_w32263_,
		_w32264_,
		_w32265_
	);
	LUT2 #(
		.INIT('h8)
	) name28219 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w4117_,
		_w32266_
	);
	LUT2 #(
		.INIT('h2)
	) name28220 (
		_w31080_,
		_w31102_,
		_w32267_
	);
	LUT2 #(
		.INIT('h8)
	) name28221 (
		_w31120_,
		_w32267_,
		_w32268_
	);
	LUT2 #(
		.INIT('h1)
	) name28222 (
		_w32266_,
		_w32268_,
		_w32269_
	);
	LUT2 #(
		.INIT('h2)
	) name28223 (
		_w4116_,
		_w32269_,
		_w32270_
	);
	LUT2 #(
		.INIT('h8)
	) name28224 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w4117_,
		_w32271_
	);
	LUT2 #(
		.INIT('h8)
	) name28225 (
		_w31127_,
		_w32267_,
		_w32272_
	);
	LUT2 #(
		.INIT('h1)
	) name28226 (
		_w32271_,
		_w32272_,
		_w32273_
	);
	LUT2 #(
		.INIT('h2)
	) name28227 (
		_w4116_,
		_w32273_,
		_w32274_
	);
	LUT2 #(
		.INIT('h8)
	) name28228 (
		\core_c_dec_MTSI_E_reg/P0001 ,
		_w4117_,
		_w32275_
	);
	LUT2 #(
		.INIT('h2)
	) name28229 (
		_w31076_,
		_w31102_,
		_w32276_
	);
	LUT2 #(
		.INIT('h8)
	) name28230 (
		_w31079_,
		_w32276_,
		_w32277_
	);
	LUT2 #(
		.INIT('h8)
	) name28231 (
		_w31127_,
		_w32277_,
		_w32278_
	);
	LUT2 #(
		.INIT('h1)
	) name28232 (
		_w32275_,
		_w32278_,
		_w32279_
	);
	LUT2 #(
		.INIT('h2)
	) name28233 (
		_w4116_,
		_w32279_,
		_w32280_
	);
	LUT2 #(
		.INIT('h8)
	) name28234 (
		\core_c_dec_MTSE_E_reg/P0001 ,
		_w4117_,
		_w32281_
	);
	LUT2 #(
		.INIT('h8)
	) name28235 (
		_w31120_,
		_w32277_,
		_w32282_
	);
	LUT2 #(
		.INIT('h1)
	) name28236 (
		_w32281_,
		_w32282_,
		_w32283_
	);
	LUT2 #(
		.INIT('h2)
	) name28237 (
		_w4116_,
		_w32283_,
		_w32284_
	);
	LUT2 #(
		.INIT('h8)
	) name28238 (
		\core_c_dec_MTMR2_E_reg/P0001 ,
		_w4117_,
		_w32285_
	);
	LUT2 #(
		.INIT('h4)
	) name28239 (
		_w31079_,
		_w32276_,
		_w32286_
	);
	LUT2 #(
		.INIT('h8)
	) name28240 (
		_w31120_,
		_w32286_,
		_w32287_
	);
	LUT2 #(
		.INIT('h1)
	) name28241 (
		_w32285_,
		_w32287_,
		_w32288_
	);
	LUT2 #(
		.INIT('h2)
	) name28242 (
		_w4116_,
		_w32288_,
		_w32289_
	);
	LUT2 #(
		.INIT('h8)
	) name28243 (
		\core_c_dec_MTMR1_E_reg/P0001 ,
		_w4117_,
		_w32290_
	);
	LUT2 #(
		.INIT('h8)
	) name28244 (
		_w31127_,
		_w32286_,
		_w32291_
	);
	LUT2 #(
		.INIT('h1)
	) name28245 (
		_w32290_,
		_w32291_,
		_w32292_
	);
	LUT2 #(
		.INIT('h2)
	) name28246 (
		_w4116_,
		_w32292_,
		_w32293_
	);
	LUT2 #(
		.INIT('h8)
	) name28247 (
		\core_c_dec_MTMR0_E_reg/P0001 ,
		_w4117_,
		_w32294_
	);
	LUT2 #(
		.INIT('h4)
	) name28248 (
		_w31102_,
		_w31545_,
		_w32295_
	);
	LUT2 #(
		.INIT('h8)
	) name28249 (
		_w31120_,
		_w32295_,
		_w32296_
	);
	LUT2 #(
		.INIT('h1)
	) name28250 (
		_w32294_,
		_w32296_,
		_w32297_
	);
	LUT2 #(
		.INIT('h2)
	) name28251 (
		_w4116_,
		_w32297_,
		_w32298_
	);
	LUT2 #(
		.INIT('h8)
	) name28252 (
		\core_c_dec_MTAR_E_reg/P0001 ,
		_w4117_,
		_w32299_
	);
	LUT2 #(
		.INIT('h8)
	) name28253 (
		_w31127_,
		_w32295_,
		_w32300_
	);
	LUT2 #(
		.INIT('h1)
	) name28254 (
		_w32299_,
		_w32300_,
		_w32301_
	);
	LUT2 #(
		.INIT('h2)
	) name28255 (
		_w4116_,
		_w32301_,
		_w32302_
	);
	LUT2 #(
		.INIT('h2)
	) name28256 (
		\sport1_rxctl_LMcnt_reg[3]/NET0131 ,
		_w30752_,
		_w32303_
	);
	LUT2 #(
		.INIT('h1)
	) name28257 (
		_w30753_,
		_w32303_,
		_w32304_
	);
	LUT2 #(
		.INIT('h2)
	) name28258 (
		_w32264_,
		_w32304_,
		_w32305_
	);
	LUT2 #(
		.INIT('h8)
	) name28259 (
		\sport1_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport1_rxctl_LMcnt_reg[1]/NET0131 ,
		_w32306_
	);
	LUT2 #(
		.INIT('h1)
	) name28260 (
		_w30751_,
		_w32306_,
		_w32307_
	);
	LUT2 #(
		.INIT('h2)
	) name28261 (
		_w32264_,
		_w32307_,
		_w32308_
	);
	LUT2 #(
		.INIT('h4)
	) name28262 (
		_w30778_,
		_w31868_,
		_w32309_
	);
	LUT2 #(
		.INIT('h2)
	) name28263 (
		\sport0_rxctl_LMcnt_reg[3]/NET0131 ,
		_w30776_,
		_w32310_
	);
	LUT2 #(
		.INIT('h1)
	) name28264 (
		_w30777_,
		_w32310_,
		_w32311_
	);
	LUT2 #(
		.INIT('h2)
	) name28265 (
		_w32309_,
		_w32311_,
		_w32312_
	);
	LUT2 #(
		.INIT('h2)
	) name28266 (
		\sport0_rxctl_LMcnt_reg[2]/NET0131 ,
		_w30775_,
		_w32313_
	);
	LUT2 #(
		.INIT('h1)
	) name28267 (
		_w30776_,
		_w32313_,
		_w32314_
	);
	LUT2 #(
		.INIT('h2)
	) name28268 (
		_w32309_,
		_w32314_,
		_w32315_
	);
	LUT2 #(
		.INIT('h8)
	) name28269 (
		\sport0_rxctl_LMcnt_reg[0]/NET0131 ,
		\sport0_rxctl_LMcnt_reg[1]/NET0131 ,
		_w32316_
	);
	LUT2 #(
		.INIT('h1)
	) name28270 (
		_w30775_,
		_w32316_,
		_w32317_
	);
	LUT2 #(
		.INIT('h2)
	) name28271 (
		_w32309_,
		_w32317_,
		_w32318_
	);
	LUT2 #(
		.INIT('h4)
	) name28272 (
		\sport0_rxctl_LMcnt_reg[0]/NET0131 ,
		_w32309_,
		_w32319_
	);
	LUT2 #(
		.INIT('h8)
	) name28273 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		_w31917_,
		_w32320_
	);
	LUT2 #(
		.INIT('h1)
	) name28274 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[5]/NET0131 ,
		_w32321_
	);
	LUT2 #(
		.INIT('h2)
	) name28275 (
		\T_TMODE[0]_pad ,
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		_w32322_
	);
	LUT2 #(
		.INIT('h8)
	) name28276 (
		_w32321_,
		_w32322_,
		_w32323_
	);
	LUT2 #(
		.INIT('h1)
	) name28277 (
		_w32320_,
		_w32323_,
		_w32324_
	);
	LUT2 #(
		.INIT('h2)
	) name28278 (
		_w23417_,
		_w32324_,
		_w32325_
	);
	LUT2 #(
		.INIT('h2)
	) name28279 (
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w32325_,
		_w32326_
	);
	LUT2 #(
		.INIT('h1)
	) name28280 (
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		\clkc_oscntr_reg_DO_reg[9]/NET0131 ,
		_w32327_
	);
	LUT2 #(
		.INIT('h4)
	) name28281 (
		\sport0_regs_AUTO_a_reg[15]/NET0131 ,
		_w32327_,
		_w32328_
	);
	LUT2 #(
		.INIT('h8)
	) name28282 (
		_w20848_,
		_w26045_,
		_w32329_
	);
	LUT2 #(
		.INIT('h8)
	) name28283 (
		_w32321_,
		_w32329_,
		_w32330_
	);
	LUT2 #(
		.INIT('h8)
	) name28284 (
		_w31913_,
		_w32328_,
		_w32331_
	);
	LUT2 #(
		.INIT('h8)
	) name28285 (
		_w32330_,
		_w32331_,
		_w32332_
	);
	LUT2 #(
		.INIT('h1)
	) name28286 (
		_w32326_,
		_w32332_,
		_w32333_
	);
	LUT2 #(
		.INIT('h1)
	) name28287 (
		\clkc_Cnt128_reg/NET0131 ,
		_w32333_,
		_w32334_
	);
	LUT2 #(
		.INIT('h1)
	) name28288 (
		\clkc_Awake_reg/NET0131 ,
		_w32334_,
		_w32335_
	);
	LUT2 #(
		.INIT('h1)
	) name28289 (
		\sport1_cfg_SCLKi_cnt_reg[12]/NET0131 ,
		_w20250_,
		_w32336_
	);
	LUT2 #(
		.INIT('h2)
	) name28290 (
		_w19130_,
		_w20251_,
		_w32337_
	);
	LUT2 #(
		.INIT('h4)
	) name28291 (
		_w32336_,
		_w32337_,
		_w32338_
	);
	LUT2 #(
		.INIT('h1)
	) name28292 (
		\sport1_cfg_SCLKi_cnt_reg[10]/NET0131 ,
		_w20240_,
		_w32339_
	);
	LUT2 #(
		.INIT('h2)
	) name28293 (
		_w19130_,
		_w20249_,
		_w32340_
	);
	LUT2 #(
		.INIT('h4)
	) name28294 (
		_w32339_,
		_w32340_,
		_w32341_
	);
	LUT2 #(
		.INIT('h4)
	) name28295 (
		\sport1_rxctl_LMcnt_reg[0]/NET0131 ,
		_w32264_,
		_w32342_
	);
	LUT2 #(
		.INIT('h2)
	) name28296 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w19504_,
		_w32343_
	);
	LUT2 #(
		.INIT('h4)
	) name28297 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w29626_,
		_w32344_
	);
	LUT2 #(
		.INIT('h1)
	) name28298 (
		_w32343_,
		_w32344_,
		_w32345_
	);
	LUT2 #(
		.INIT('h2)
	) name28299 (
		_w18717_,
		_w32345_,
		_w32346_
	);
	LUT2 #(
		.INIT('h1)
	) name28300 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[9]/P0001 ,
		_w18717_,
		_w32347_
	);
	LUT2 #(
		.INIT('h1)
	) name28301 (
		_w32346_,
		_w32347_,
		_w32348_
	);
	LUT2 #(
		.INIT('h2)
	) name28302 (
		\core_c_psq_Iact_E_reg[3]/NET0131 ,
		_w4116_,
		_w32349_
	);
	LUT2 #(
		.INIT('h2)
	) name28303 (
		\core_c_psq_T_IRQE0_reg/P0001 ,
		\core_c_psq_T_IRQE0_s1_reg/P0001 ,
		_w32350_
	);
	LUT2 #(
		.INIT('h8)
	) name28304 (
		_w4064_,
		_w13757_,
		_w32351_
	);
	LUT2 #(
		.INIT('h1)
	) name28305 (
		\core_c_psq_IFC_reg[11]/NET0131 ,
		\core_c_psq_Iflag_reg[3]/NET0131 ,
		_w32352_
	);
	LUT2 #(
		.INIT('h4)
	) name28306 (
		_w32350_,
		_w32352_,
		_w32353_
	);
	LUT2 #(
		.INIT('h4)
	) name28307 (
		_w32351_,
		_w32353_,
		_w32354_
	);
	LUT2 #(
		.INIT('h1)
	) name28308 (
		\core_c_psq_IFC_reg[3]/NET0131 ,
		_w32349_,
		_w32355_
	);
	LUT2 #(
		.INIT('h4)
	) name28309 (
		_w32354_,
		_w32355_,
		_w32356_
	);
	LUT2 #(
		.INIT('h2)
	) name28310 (
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		_w4116_,
		_w32357_
	);
	LUT2 #(
		.INIT('h1)
	) name28311 (
		\T_TMODE[0]_pad ,
		\tm_TINT_GEN1_reg/NET0131 ,
		_w32358_
	);
	LUT2 #(
		.INIT('h8)
	) name28312 (
		\tm_TINT_GEN2_reg/NET0131 ,
		_w32358_,
		_w32359_
	);
	LUT2 #(
		.INIT('h1)
	) name28313 (
		\core_c_psq_IFC_reg[8]/NET0131 ,
		\core_c_psq_Iflag_reg[0]/NET0131 ,
		_w32360_
	);
	LUT2 #(
		.INIT('h4)
	) name28314 (
		_w32359_,
		_w32360_,
		_w32361_
	);
	LUT2 #(
		.INIT('h1)
	) name28315 (
		\core_c_psq_IFC_reg[0]/NET0131 ,
		_w32361_,
		_w32362_
	);
	LUT2 #(
		.INIT('h4)
	) name28316 (
		_w32357_,
		_w32362_,
		_w32363_
	);
	LUT2 #(
		.INIT('h1)
	) name28317 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w4112_,
		_w32364_
	);
	LUT2 #(
		.INIT('h1)
	) name28318 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w14697_,
		_w32365_
	);
	LUT2 #(
		.INIT('h1)
	) name28319 (
		_w5950_,
		_w32365_,
		_w32366_
	);
	LUT2 #(
		.INIT('h4)
	) name28320 (
		_w32364_,
		_w32366_,
		_w32367_
	);
	LUT2 #(
		.INIT('h2)
	) name28321 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w8113_,
		_w32368_
	);
	LUT2 #(
		.INIT('h8)
	) name28322 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][18]/P0001 ,
		_w14708_,
		_w32369_
	);
	LUT2 #(
		.INIT('h8)
	) name28323 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][18]/P0001 ,
		_w14713_,
		_w32370_
	);
	LUT2 #(
		.INIT('h8)
	) name28324 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001 ,
		_w14711_,
		_w32371_
	);
	LUT2 #(
		.INIT('h8)
	) name28325 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001 ,
		_w14699_,
		_w32372_
	);
	LUT2 #(
		.INIT('h8)
	) name28326 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001 ,
		_w14704_,
		_w32373_
	);
	LUT2 #(
		.INIT('h8)
	) name28327 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][18]/P0001 ,
		_w14702_,
		_w32374_
	);
	LUT2 #(
		.INIT('h8)
	) name28328 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001 ,
		_w14706_,
		_w32375_
	);
	LUT2 #(
		.INIT('h1)
	) name28329 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w32369_,
		_w32376_
	);
	LUT2 #(
		.INIT('h1)
	) name28330 (
		_w32370_,
		_w32371_,
		_w32377_
	);
	LUT2 #(
		.INIT('h1)
	) name28331 (
		_w32372_,
		_w32373_,
		_w32378_
	);
	LUT2 #(
		.INIT('h1)
	) name28332 (
		_w32374_,
		_w32375_,
		_w32379_
	);
	LUT2 #(
		.INIT('h8)
	) name28333 (
		_w32378_,
		_w32379_,
		_w32380_
	);
	LUT2 #(
		.INIT('h8)
	) name28334 (
		_w32376_,
		_w32377_,
		_w32381_
	);
	LUT2 #(
		.INIT('h8)
	) name28335 (
		_w32380_,
		_w32381_,
		_w32382_
	);
	LUT2 #(
		.INIT('h1)
	) name28336 (
		_w32368_,
		_w32382_,
		_w32383_
	);
	LUT2 #(
		.INIT('h8)
	) name28337 (
		_w32367_,
		_w32383_,
		_w32384_
	);
	LUT2 #(
		.INIT('h4)
	) name28338 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		_w5299_,
		_w32385_
	);
	LUT2 #(
		.INIT('h2)
	) name28339 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w32385_,
		_w32386_
	);
	LUT2 #(
		.INIT('h2)
	) name28340 (
		_w32364_,
		_w32386_,
		_w32387_
	);
	LUT2 #(
		.INIT('h2)
	) name28341 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w32387_,
		_w32388_
	);
	LUT2 #(
		.INIT('h4)
	) name28342 (
		_w32367_,
		_w32388_,
		_w32389_
	);
	LUT2 #(
		.INIT('h1)
	) name28343 (
		_w32384_,
		_w32389_,
		_w32390_
	);
	LUT2 #(
		.INIT('h2)
	) name28344 (
		_w17833_,
		_w32345_,
		_w32391_
	);
	LUT2 #(
		.INIT('h1)
	) name28345 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[9]/P0001 ,
		_w17833_,
		_w32392_
	);
	LUT2 #(
		.INIT('h1)
	) name28346 (
		_w32391_,
		_w32392_,
		_w32393_
	);
	LUT2 #(
		.INIT('h4)
	) name28347 (
		\sport0_rxctl_RXSHT_reg[14]/P0001 ,
		_w20868_,
		_w32394_
	);
	LUT2 #(
		.INIT('h8)
	) name28348 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w32395_
	);
	LUT2 #(
		.INIT('h8)
	) name28349 (
		_w20913_,
		_w32395_,
		_w32396_
	);
	LUT2 #(
		.INIT('h4)
	) name28350 (
		_w20888_,
		_w32396_,
		_w32397_
	);
	LUT2 #(
		.INIT('h8)
	) name28351 (
		_w20881_,
		_w32397_,
		_w32398_
	);
	LUT2 #(
		.INIT('h4)
	) name28352 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w20875_,
		_w32399_
	);
	LUT2 #(
		.INIT('h4)
	) name28353 (
		_w32398_,
		_w32399_,
		_w32400_
	);
	LUT2 #(
		.INIT('h4)
	) name28354 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w12688_,
		_w32401_
	);
	LUT2 #(
		.INIT('h8)
	) name28355 (
		\sport0_rxctl_RX_reg[14]/P0001 ,
		_w20873_,
		_w32402_
	);
	LUT2 #(
		.INIT('h1)
	) name28356 (
		_w20868_,
		_w32402_,
		_w32403_
	);
	LUT2 #(
		.INIT('h4)
	) name28357 (
		_w32400_,
		_w32403_,
		_w32404_
	);
	LUT2 #(
		.INIT('h4)
	) name28358 (
		_w32401_,
		_w32404_,
		_w32405_
	);
	LUT2 #(
		.INIT('h1)
	) name28359 (
		_w20871_,
		_w32394_,
		_w32406_
	);
	LUT2 #(
		.INIT('h4)
	) name28360 (
		_w32405_,
		_w32406_,
		_w32407_
	);
	LUT2 #(
		.INIT('h8)
	) name28361 (
		\sport0_rxctl_RX_reg[14]/P0001 ,
		_w20871_,
		_w32408_
	);
	LUT2 #(
		.INIT('h1)
	) name28362 (
		_w32407_,
		_w32408_,
		_w32409_
	);
	LUT2 #(
		.INIT('h4)
	) name28363 (
		\sport0_rxctl_RXSHT_reg[15]/P0001 ,
		_w20868_,
		_w32410_
	);
	LUT2 #(
		.INIT('h4)
	) name28364 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w12743_,
		_w32411_
	);
	LUT2 #(
		.INIT('h8)
	) name28365 (
		\sport0_rxctl_RX_reg[15]/P0001 ,
		_w20873_,
		_w32412_
	);
	LUT2 #(
		.INIT('h1)
	) name28366 (
		_w20868_,
		_w32412_,
		_w32413_
	);
	LUT2 #(
		.INIT('h4)
	) name28367 (
		_w32400_,
		_w32413_,
		_w32414_
	);
	LUT2 #(
		.INIT('h4)
	) name28368 (
		_w32411_,
		_w32414_,
		_w32415_
	);
	LUT2 #(
		.INIT('h1)
	) name28369 (
		_w20871_,
		_w32410_,
		_w32416_
	);
	LUT2 #(
		.INIT('h4)
	) name28370 (
		_w32415_,
		_w32416_,
		_w32417_
	);
	LUT2 #(
		.INIT('h8)
	) name28371 (
		\sport0_rxctl_RX_reg[15]/P0001 ,
		_w20871_,
		_w32418_
	);
	LUT2 #(
		.INIT('h1)
	) name28372 (
		_w32417_,
		_w32418_,
		_w32419_
	);
	LUT2 #(
		.INIT('h4)
	) name28373 (
		_w29560_,
		_w31064_,
		_w32420_
	);
	LUT2 #(
		.INIT('h2)
	) name28374 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[9]/P0001 ,
		_w31064_,
		_w32421_
	);
	LUT2 #(
		.INIT('h1)
	) name28375 (
		_w32420_,
		_w32421_,
		_w32422_
	);
	LUT2 #(
		.INIT('h2)
	) name28376 (
		_w27915_,
		_w28023_,
		_w32423_
	);
	LUT2 #(
		.INIT('h2)
	) name28377 (
		\core_c_psq_CNTR_reg_DO_reg[9]/NET0131 ,
		_w27915_,
		_w32424_
	);
	LUT2 #(
		.INIT('h1)
	) name28378 (
		_w32423_,
		_w32424_,
		_w32425_
	);
	LUT2 #(
		.INIT('h2)
	) name28379 (
		_w27915_,
		_w27978_,
		_w32426_
	);
	LUT2 #(
		.INIT('h2)
	) name28380 (
		\core_c_psq_CNTR_reg_DO_reg[8]/NET0131 ,
		_w27915_,
		_w32427_
	);
	LUT2 #(
		.INIT('h1)
	) name28381 (
		_w32426_,
		_w32427_,
		_w32428_
	);
	LUT2 #(
		.INIT('h2)
	) name28382 (
		_w27915_,
		_w27993_,
		_w32429_
	);
	LUT2 #(
		.INIT('h2)
	) name28383 (
		\core_c_psq_CNTR_reg_DO_reg[4]/NET0131 ,
		_w27915_,
		_w32430_
	);
	LUT2 #(
		.INIT('h1)
	) name28384 (
		_w32429_,
		_w32430_,
		_w32431_
	);
	LUT2 #(
		.INIT('h2)
	) name28385 (
		_w27915_,
		_w28038_,
		_w32432_
	);
	LUT2 #(
		.INIT('h2)
	) name28386 (
		\core_c_psq_CNTR_reg_DO_reg[3]/NET0131 ,
		_w27915_,
		_w32433_
	);
	LUT2 #(
		.INIT('h1)
	) name28387 (
		_w32432_,
		_w32433_,
		_w32434_
	);
	LUT2 #(
		.INIT('h4)
	) name28388 (
		_w30397_,
		_w31064_,
		_w32435_
	);
	LUT2 #(
		.INIT('h2)
	) name28389 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[8]/P0001 ,
		_w31064_,
		_w32436_
	);
	LUT2 #(
		.INIT('h1)
	) name28390 (
		_w32435_,
		_w32436_,
		_w32437_
	);
	LUT2 #(
		.INIT('h2)
	) name28391 (
		_w27915_,
		_w28069_,
		_w32438_
	);
	LUT2 #(
		.INIT('h2)
	) name28392 (
		\core_c_psq_CNTR_reg_DO_reg[2]/NET0131 ,
		_w27915_,
		_w32439_
	);
	LUT2 #(
		.INIT('h1)
	) name28393 (
		_w32438_,
		_w32439_,
		_w32440_
	);
	LUT2 #(
		.INIT('h2)
	) name28394 (
		_w27915_,
		_w27948_,
		_w32441_
	);
	LUT2 #(
		.INIT('h2)
	) name28395 (
		\core_c_psq_CNTR_reg_DO_reg[12]/NET0131 ,
		_w27915_,
		_w32442_
	);
	LUT2 #(
		.INIT('h1)
	) name28396 (
		_w32441_,
		_w32442_,
		_w32443_
	);
	LUT2 #(
		.INIT('h2)
	) name28397 (
		_w27915_,
		_w28143_,
		_w32444_
	);
	LUT2 #(
		.INIT('h2)
	) name28398 (
		\core_c_psq_CNTR_reg_DO_reg[11]/NET0131 ,
		_w27915_,
		_w32445_
	);
	LUT2 #(
		.INIT('h1)
	) name28399 (
		_w32444_,
		_w32445_,
		_w32446_
	);
	LUT2 #(
		.INIT('h2)
	) name28400 (
		_w27915_,
		_w27963_,
		_w32447_
	);
	LUT2 #(
		.INIT('h2)
	) name28401 (
		\core_c_psq_CNTR_reg_DO_reg[10]/NET0131 ,
		_w27915_,
		_w32448_
	);
	LUT2 #(
		.INIT('h1)
	) name28402 (
		_w32447_,
		_w32448_,
		_w32449_
	);
	LUT2 #(
		.INIT('h4)
	) name28403 (
		_w30191_,
		_w31064_,
		_w32450_
	);
	LUT2 #(
		.INIT('h2)
	) name28404 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[7]/P0001 ,
		_w31064_,
		_w32451_
	);
	LUT2 #(
		.INIT('h1)
	) name28405 (
		_w32450_,
		_w32451_,
		_w32452_
	);
	LUT2 #(
		.INIT('h1)
	) name28406 (
		IACKn_pad,
		\idma_IAL_reg/P0001 ,
		_w32453_
	);
	LUT2 #(
		.INIT('h8)
	) name28407 (
		\memc_MMR_web_reg/NET0131 ,
		_w32453_,
		_w32454_
	);
	LUT2 #(
		.INIT('h1)
	) name28408 (
		_w20073_,
		_w32454_,
		_w32455_
	);
	LUT2 #(
		.INIT('h1)
	) name28409 (
		\idma_IAL_reg/P0001 ,
		_w10638_,
		_w32456_
	);
	LUT2 #(
		.INIT('h4)
	) name28410 (
		\idma_IADi_reg[8]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32457_
	);
	LUT2 #(
		.INIT('h1)
	) name28411 (
		_w32456_,
		_w32457_,
		_w32458_
	);
	LUT2 #(
		.INIT('h8)
	) name28412 (
		_w32455_,
		_w32458_,
		_w32459_
	);
	LUT2 #(
		.INIT('h4)
	) name28413 (
		\idma_DCTL_reg[14]/NET0131 ,
		\idma_PM_1st_reg/NET0131 ,
		_w32460_
	);
	LUT2 #(
		.INIT('h2)
	) name28414 (
		\auctl_DSack_reg/NET0131 ,
		_w32460_,
		_w32461_
	);
	LUT2 #(
		.INIT('h8)
	) name28415 (
		_w20382_,
		_w32460_,
		_w32462_
	);
	LUT2 #(
		.INIT('h1)
	) name28416 (
		_w32461_,
		_w32462_,
		_w32463_
	);
	LUT2 #(
		.INIT('h2)
	) name28417 (
		\idma_WRcyc_reg/NET0131 ,
		_w32463_,
		_w32464_
	);
	LUT2 #(
		.INIT('h1)
	) name28418 (
		_w20394_,
		_w32464_,
		_w32465_
	);
	LUT2 #(
		.INIT('h1)
	) name28419 (
		_w32454_,
		_w32460_,
		_w32466_
	);
	LUT2 #(
		.INIT('h4)
	) name28420 (
		_w32465_,
		_w32466_,
		_w32467_
	);
	LUT2 #(
		.INIT('h8)
	) name28421 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w32467_,
		_w32468_
	);
	LUT2 #(
		.INIT('h8)
	) name28422 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w32468_,
		_w32469_
	);
	LUT2 #(
		.INIT('h8)
	) name28423 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w32469_,
		_w32470_
	);
	LUT2 #(
		.INIT('h8)
	) name28424 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w32470_,
		_w32471_
	);
	LUT2 #(
		.INIT('h8)
	) name28425 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w32471_,
		_w32472_
	);
	LUT2 #(
		.INIT('h8)
	) name28426 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w32472_,
		_w32473_
	);
	LUT2 #(
		.INIT('h8)
	) name28427 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w32473_,
		_w32474_
	);
	LUT2 #(
		.INIT('h8)
	) name28428 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w32474_,
		_w32475_
	);
	LUT2 #(
		.INIT('h1)
	) name28429 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w32475_,
		_w32476_
	);
	LUT2 #(
		.INIT('h8)
	) name28430 (
		\idma_DCTL_reg[8]/NET0131 ,
		_w32475_,
		_w32477_
	);
	LUT2 #(
		.INIT('h1)
	) name28431 (
		_w32455_,
		_w32476_,
		_w32478_
	);
	LUT2 #(
		.INIT('h4)
	) name28432 (
		_w32477_,
		_w32478_,
		_w32479_
	);
	LUT2 #(
		.INIT('h1)
	) name28433 (
		_w32459_,
		_w32479_,
		_w32480_
	);
	LUT2 #(
		.INIT('h1)
	) name28434 (
		\idma_IAL_reg/P0001 ,
		_w10289_,
		_w32481_
	);
	LUT2 #(
		.INIT('h4)
	) name28435 (
		\idma_IADi_reg[9]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32482_
	);
	LUT2 #(
		.INIT('h1)
	) name28436 (
		_w32481_,
		_w32482_,
		_w32483_
	);
	LUT2 #(
		.INIT('h8)
	) name28437 (
		_w32455_,
		_w32483_,
		_w32484_
	);
	LUT2 #(
		.INIT('h1)
	) name28438 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w32477_,
		_w32485_
	);
	LUT2 #(
		.INIT('h8)
	) name28439 (
		\idma_DCTL_reg[9]/NET0131 ,
		_w32477_,
		_w32486_
	);
	LUT2 #(
		.INIT('h1)
	) name28440 (
		_w32455_,
		_w32485_,
		_w32487_
	);
	LUT2 #(
		.INIT('h4)
	) name28441 (
		_w32486_,
		_w32487_,
		_w32488_
	);
	LUT2 #(
		.INIT('h1)
	) name28442 (
		_w32484_,
		_w32488_,
		_w32489_
	);
	LUT2 #(
		.INIT('h4)
	) name28443 (
		\idma_IADi_reg[13]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32490_
	);
	LUT2 #(
		.INIT('h1)
	) name28444 (
		\idma_IAL_reg/P0001 ,
		_w7340_,
		_w32491_
	);
	LUT2 #(
		.INIT('h2)
	) name28445 (
		_w32455_,
		_w32490_,
		_w32492_
	);
	LUT2 #(
		.INIT('h4)
	) name28446 (
		_w32491_,
		_w32492_,
		_w32493_
	);
	LUT2 #(
		.INIT('h8)
	) name28447 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w32486_,
		_w32494_
	);
	LUT2 #(
		.INIT('h8)
	) name28448 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w32494_,
		_w32495_
	);
	LUT2 #(
		.INIT('h8)
	) name28449 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w32495_,
		_w32496_
	);
	LUT2 #(
		.INIT('h1)
	) name28450 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w32496_,
		_w32497_
	);
	LUT2 #(
		.INIT('h8)
	) name28451 (
		\idma_DCTL_reg[13]/NET0131 ,
		_w32496_,
		_w32498_
	);
	LUT2 #(
		.INIT('h1)
	) name28452 (
		_w32455_,
		_w32497_,
		_w32499_
	);
	LUT2 #(
		.INIT('h4)
	) name28453 (
		_w32498_,
		_w32499_,
		_w32500_
	);
	LUT2 #(
		.INIT('h1)
	) name28454 (
		_w32493_,
		_w32500_,
		_w32501_
	);
	LUT2 #(
		.INIT('h1)
	) name28455 (
		\idma_DCTL_reg[12]/NET0131 ,
		_w32495_,
		_w32502_
	);
	LUT2 #(
		.INIT('h1)
	) name28456 (
		_w32496_,
		_w32502_,
		_w32503_
	);
	LUT2 #(
		.INIT('h1)
	) name28457 (
		_w32455_,
		_w32503_,
		_w32504_
	);
	LUT2 #(
		.INIT('h4)
	) name28458 (
		\idma_IAL_reg/P0001 ,
		_w9178_,
		_w32505_
	);
	LUT2 #(
		.INIT('h8)
	) name28459 (
		\idma_IADi_reg[12]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32506_
	);
	LUT2 #(
		.INIT('h2)
	) name28460 (
		_w32455_,
		_w32506_,
		_w32507_
	);
	LUT2 #(
		.INIT('h4)
	) name28461 (
		_w32505_,
		_w32507_,
		_w32508_
	);
	LUT2 #(
		.INIT('h1)
	) name28462 (
		_w32504_,
		_w32508_,
		_w32509_
	);
	LUT2 #(
		.INIT('h1)
	) name28463 (
		\idma_IAL_reg/P0001 ,
		_w8460_,
		_w32510_
	);
	LUT2 #(
		.INIT('h4)
	) name28464 (
		\idma_IADi_reg[11]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32511_
	);
	LUT2 #(
		.INIT('h1)
	) name28465 (
		_w32510_,
		_w32511_,
		_w32512_
	);
	LUT2 #(
		.INIT('h8)
	) name28466 (
		_w32455_,
		_w32512_,
		_w32513_
	);
	LUT2 #(
		.INIT('h1)
	) name28467 (
		\idma_DCTL_reg[11]/NET0131 ,
		_w32494_,
		_w32514_
	);
	LUT2 #(
		.INIT('h1)
	) name28468 (
		_w32455_,
		_w32495_,
		_w32515_
	);
	LUT2 #(
		.INIT('h4)
	) name28469 (
		_w32514_,
		_w32515_,
		_w32516_
	);
	LUT2 #(
		.INIT('h1)
	) name28470 (
		_w32513_,
		_w32516_,
		_w32517_
	);
	LUT2 #(
		.INIT('h1)
	) name28471 (
		\idma_IAL_reg/P0001 ,
		_w7859_,
		_w32518_
	);
	LUT2 #(
		.INIT('h4)
	) name28472 (
		\idma_IADi_reg[10]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32519_
	);
	LUT2 #(
		.INIT('h1)
	) name28473 (
		_w32518_,
		_w32519_,
		_w32520_
	);
	LUT2 #(
		.INIT('h8)
	) name28474 (
		_w32455_,
		_w32520_,
		_w32521_
	);
	LUT2 #(
		.INIT('h1)
	) name28475 (
		\idma_DCTL_reg[10]/NET0131 ,
		_w32486_,
		_w32522_
	);
	LUT2 #(
		.INIT('h1)
	) name28476 (
		_w32455_,
		_w32494_,
		_w32523_
	);
	LUT2 #(
		.INIT('h4)
	) name28477 (
		_w32522_,
		_w32523_,
		_w32524_
	);
	LUT2 #(
		.INIT('h1)
	) name28478 (
		_w32521_,
		_w32524_,
		_w32525_
	);
	LUT2 #(
		.INIT('h4)
	) name28479 (
		_w28990_,
		_w31064_,
		_w32526_
	);
	LUT2 #(
		.INIT('h2)
	) name28480 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[6]/P0001 ,
		_w31064_,
		_w32527_
	);
	LUT2 #(
		.INIT('h1)
	) name28481 (
		_w32526_,
		_w32527_,
		_w32528_
	);
	LUT2 #(
		.INIT('h4)
	) name28482 (
		\sport0_rxctl_RXSHT_reg[13]/P0001 ,
		_w20868_,
		_w32529_
	);
	LUT2 #(
		.INIT('h4)
	) name28483 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w7340_,
		_w32530_
	);
	LUT2 #(
		.INIT('h8)
	) name28484 (
		\sport0_rxctl_RX_reg[13]/P0001 ,
		_w20873_,
		_w32531_
	);
	LUT2 #(
		.INIT('h1)
	) name28485 (
		_w20868_,
		_w32531_,
		_w32532_
	);
	LUT2 #(
		.INIT('h4)
	) name28486 (
		_w32400_,
		_w32532_,
		_w32533_
	);
	LUT2 #(
		.INIT('h4)
	) name28487 (
		_w32530_,
		_w32533_,
		_w32534_
	);
	LUT2 #(
		.INIT('h1)
	) name28488 (
		_w20871_,
		_w32529_,
		_w32535_
	);
	LUT2 #(
		.INIT('h4)
	) name28489 (
		_w32534_,
		_w32535_,
		_w32536_
	);
	LUT2 #(
		.INIT('h8)
	) name28490 (
		\sport0_rxctl_RX_reg[13]/P0001 ,
		_w20871_,
		_w32537_
	);
	LUT2 #(
		.INIT('h1)
	) name28491 (
		_w32536_,
		_w32537_,
		_w32538_
	);
	LUT2 #(
		.INIT('h1)
	) name28492 (
		\idma_IAL_reg/P0001 ,
		_w11265_,
		_w32539_
	);
	LUT2 #(
		.INIT('h4)
	) name28493 (
		\idma_IADi_reg[7]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32540_
	);
	LUT2 #(
		.INIT('h1)
	) name28494 (
		_w32539_,
		_w32540_,
		_w32541_
	);
	LUT2 #(
		.INIT('h8)
	) name28495 (
		_w32455_,
		_w32541_,
		_w32542_
	);
	LUT2 #(
		.INIT('h1)
	) name28496 (
		\idma_DCTL_reg[7]/NET0131 ,
		_w32474_,
		_w32543_
	);
	LUT2 #(
		.INIT('h1)
	) name28497 (
		_w32455_,
		_w32475_,
		_w32544_
	);
	LUT2 #(
		.INIT('h4)
	) name28498 (
		_w32543_,
		_w32544_,
		_w32545_
	);
	LUT2 #(
		.INIT('h1)
	) name28499 (
		_w32542_,
		_w32545_,
		_w32546_
	);
	LUT2 #(
		.INIT('h1)
	) name28500 (
		\idma_IAL_reg/P0001 ,
		_w10911_,
		_w32547_
	);
	LUT2 #(
		.INIT('h4)
	) name28501 (
		\idma_IADi_reg[5]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32548_
	);
	LUT2 #(
		.INIT('h1)
	) name28502 (
		_w32547_,
		_w32548_,
		_w32549_
	);
	LUT2 #(
		.INIT('h8)
	) name28503 (
		_w32455_,
		_w32549_,
		_w32550_
	);
	LUT2 #(
		.INIT('h1)
	) name28504 (
		\idma_DCTL_reg[5]/NET0131 ,
		_w32472_,
		_w32551_
	);
	LUT2 #(
		.INIT('h1)
	) name28505 (
		_w32473_,
		_w32551_,
		_w32552_
	);
	LUT2 #(
		.INIT('h4)
	) name28506 (
		_w32455_,
		_w32552_,
		_w32553_
	);
	LUT2 #(
		.INIT('h1)
	) name28507 (
		_w32550_,
		_w32553_,
		_w32554_
	);
	LUT2 #(
		.INIT('h1)
	) name28508 (
		\idma_IAL_reg/P0001 ,
		_w11525_,
		_w32555_
	);
	LUT2 #(
		.INIT('h4)
	) name28509 (
		\idma_IADi_reg[6]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32556_
	);
	LUT2 #(
		.INIT('h1)
	) name28510 (
		_w32555_,
		_w32556_,
		_w32557_
	);
	LUT2 #(
		.INIT('h8)
	) name28511 (
		_w32455_,
		_w32557_,
		_w32558_
	);
	LUT2 #(
		.INIT('h1)
	) name28512 (
		\idma_DCTL_reg[6]/NET0131 ,
		_w32473_,
		_w32559_
	);
	LUT2 #(
		.INIT('h1)
	) name28513 (
		_w32455_,
		_w32474_,
		_w32560_
	);
	LUT2 #(
		.INIT('h4)
	) name28514 (
		_w32559_,
		_w32560_,
		_w32561_
	);
	LUT2 #(
		.INIT('h1)
	) name28515 (
		_w32558_,
		_w32561_,
		_w32562_
	);
	LUT2 #(
		.INIT('h1)
	) name28516 (
		\idma_IAL_reg/P0001 ,
		_w10069_,
		_w32563_
	);
	LUT2 #(
		.INIT('h4)
	) name28517 (
		\idma_IADi_reg[4]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32564_
	);
	LUT2 #(
		.INIT('h1)
	) name28518 (
		_w32563_,
		_w32564_,
		_w32565_
	);
	LUT2 #(
		.INIT('h8)
	) name28519 (
		_w32455_,
		_w32565_,
		_w32566_
	);
	LUT2 #(
		.INIT('h1)
	) name28520 (
		\idma_DCTL_reg[4]/NET0131 ,
		_w32471_,
		_w32567_
	);
	LUT2 #(
		.INIT('h1)
	) name28521 (
		_w32472_,
		_w32567_,
		_w32568_
	);
	LUT2 #(
		.INIT('h4)
	) name28522 (
		_w32455_,
		_w32568_,
		_w32569_
	);
	LUT2 #(
		.INIT('h1)
	) name28523 (
		_w32566_,
		_w32569_,
		_w32570_
	);
	LUT2 #(
		.INIT('h1)
	) name28524 (
		\idma_IAL_reg/P0001 ,
		_w8113_,
		_w32571_
	);
	LUT2 #(
		.INIT('h4)
	) name28525 (
		\idma_IADi_reg[3]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32572_
	);
	LUT2 #(
		.INIT('h1)
	) name28526 (
		_w32571_,
		_w32572_,
		_w32573_
	);
	LUT2 #(
		.INIT('h8)
	) name28527 (
		_w32455_,
		_w32573_,
		_w32574_
	);
	LUT2 #(
		.INIT('h1)
	) name28528 (
		\idma_DCTL_reg[3]/NET0131 ,
		_w32470_,
		_w32575_
	);
	LUT2 #(
		.INIT('h1)
	) name28529 (
		_w32471_,
		_w32575_,
		_w32576_
	);
	LUT2 #(
		.INIT('h4)
	) name28530 (
		_w32455_,
		_w32576_,
		_w32577_
	);
	LUT2 #(
		.INIT('h1)
	) name28531 (
		_w32574_,
		_w32577_,
		_w32578_
	);
	LUT2 #(
		.INIT('h1)
	) name28532 (
		\idma_IAL_reg/P0001 ,
		_w8715_,
		_w32579_
	);
	LUT2 #(
		.INIT('h4)
	) name28533 (
		\idma_IADi_reg[2]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32580_
	);
	LUT2 #(
		.INIT('h1)
	) name28534 (
		_w32579_,
		_w32580_,
		_w32581_
	);
	LUT2 #(
		.INIT('h8)
	) name28535 (
		_w32455_,
		_w32581_,
		_w32582_
	);
	LUT2 #(
		.INIT('h1)
	) name28536 (
		\idma_DCTL_reg[2]/NET0131 ,
		_w32469_,
		_w32583_
	);
	LUT2 #(
		.INIT('h1)
	) name28537 (
		_w32470_,
		_w32583_,
		_w32584_
	);
	LUT2 #(
		.INIT('h4)
	) name28538 (
		_w32455_,
		_w32584_,
		_w32585_
	);
	LUT2 #(
		.INIT('h1)
	) name28539 (
		_w32582_,
		_w32585_,
		_w32586_
	);
	LUT2 #(
		.INIT('h1)
	) name28540 (
		\idma_IAL_reg/P0001 ,
		_w7607_,
		_w32587_
	);
	LUT2 #(
		.INIT('h4)
	) name28541 (
		\idma_IADi_reg[0]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32588_
	);
	LUT2 #(
		.INIT('h1)
	) name28542 (
		_w32587_,
		_w32588_,
		_w32589_
	);
	LUT2 #(
		.INIT('h8)
	) name28543 (
		_w32455_,
		_w32589_,
		_w32590_
	);
	LUT2 #(
		.INIT('h1)
	) name28544 (
		\idma_DCTL_reg[0]/NET0131 ,
		_w32467_,
		_w32591_
	);
	LUT2 #(
		.INIT('h1)
	) name28545 (
		_w32468_,
		_w32591_,
		_w32592_
	);
	LUT2 #(
		.INIT('h4)
	) name28546 (
		_w32455_,
		_w32592_,
		_w32593_
	);
	LUT2 #(
		.INIT('h1)
	) name28547 (
		_w32590_,
		_w32593_,
		_w32594_
	);
	LUT2 #(
		.INIT('h4)
	) name28548 (
		_w29042_,
		_w31064_,
		_w32595_
	);
	LUT2 #(
		.INIT('h2)
	) name28549 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[5]/P0001 ,
		_w31064_,
		_w32596_
	);
	LUT2 #(
		.INIT('h1)
	) name28550 (
		_w32595_,
		_w32596_,
		_w32597_
	);
	LUT2 #(
		.INIT('h2)
	) name28551 (
		_w27915_,
		_w28098_,
		_w32598_
	);
	LUT2 #(
		.INIT('h2)
	) name28552 (
		\core_c_psq_CNTR_reg_DO_reg[7]/NET0131 ,
		_w27915_,
		_w32599_
	);
	LUT2 #(
		.INIT('h1)
	) name28553 (
		_w32598_,
		_w32599_,
		_w32600_
	);
	LUT2 #(
		.INIT('h2)
	) name28554 (
		_w27915_,
		_w28113_,
		_w32601_
	);
	LUT2 #(
		.INIT('h2)
	) name28555 (
		\core_c_psq_CNTR_reg_DO_reg[6]/NET0131 ,
		_w27915_,
		_w32602_
	);
	LUT2 #(
		.INIT('h1)
	) name28556 (
		_w32601_,
		_w32602_,
		_w32603_
	);
	LUT2 #(
		.INIT('h2)
	) name28557 (
		\core_c_psq_CNTR_reg_DO_reg[0]/NET0131 ,
		_w27915_,
		_w32604_
	);
	LUT2 #(
		.INIT('h1)
	) name28558 (
		_w28083_,
		_w32604_,
		_w32605_
	);
	LUT2 #(
		.INIT('h8)
	) name28559 (
		_w31697_,
		_w31703_,
		_w32606_
	);
	LUT2 #(
		.INIT('h1)
	) name28560 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[1]/NET0131 ,
		_w32607_
	);
	LUT2 #(
		.INIT('h1)
	) name28561 (
		\sport1_rxctl_Wcnt_reg[2]/NET0131 ,
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		_w32608_
	);
	LUT2 #(
		.INIT('h8)
	) name28562 (
		_w32607_,
		_w32608_,
		_w32609_
	);
	LUT2 #(
		.INIT('h8)
	) name28563 (
		_w20408_,
		_w32609_,
		_w32610_
	);
	LUT2 #(
		.INIT('h8)
	) name28564 (
		_w32606_,
		_w32610_,
		_w32611_
	);
	LUT2 #(
		.INIT('h1)
	) name28565 (
		_w31702_,
		_w32611_,
		_w32612_
	);
	LUT2 #(
		.INIT('h2)
	) name28566 (
		_w32606_,
		_w32610_,
		_w32613_
	);
	LUT2 #(
		.INIT('h8)
	) name28567 (
		_w32607_,
		_w32613_,
		_w32614_
	);
	LUT2 #(
		.INIT('h4)
	) name28568 (
		\sport1_rxctl_Wcnt_reg[2]/NET0131 ,
		_w32614_,
		_w32615_
	);
	LUT2 #(
		.INIT('h4)
	) name28569 (
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		_w32615_,
		_w32616_
	);
	LUT2 #(
		.INIT('h2)
	) name28570 (
		\sport1_rxctl_Wcnt_reg[4]/NET0131 ,
		_w32616_,
		_w32617_
	);
	LUT2 #(
		.INIT('h4)
	) name28571 (
		\sport1_rxctl_Wcnt_reg[4]/NET0131 ,
		_w32616_,
		_w32618_
	);
	LUT2 #(
		.INIT('h1)
	) name28572 (
		_w32617_,
		_w32618_,
		_w32619_
	);
	LUT2 #(
		.INIT('h2)
	) name28573 (
		_w32612_,
		_w32619_,
		_w32620_
	);
	LUT2 #(
		.INIT('h2)
	) name28574 (
		\sport1_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w32612_,
		_w32621_
	);
	LUT2 #(
		.INIT('h1)
	) name28575 (
		_w32620_,
		_w32621_,
		_w32622_
	);
	LUT2 #(
		.INIT('h2)
	) name28576 (
		_w27915_,
		_w28128_,
		_w32623_
	);
	LUT2 #(
		.INIT('h2)
	) name28577 (
		\core_c_psq_CNTR_reg_DO_reg[5]/NET0131 ,
		_w27915_,
		_w32624_
	);
	LUT2 #(
		.INIT('h1)
	) name28578 (
		_w32623_,
		_w32624_,
		_w32625_
	);
	LUT2 #(
		.INIT('h2)
	) name28579 (
		_w27915_,
		_w28008_,
		_w32626_
	);
	LUT2 #(
		.INIT('h2)
	) name28580 (
		\core_c_psq_CNTR_reg_DO_reg[1]/NET0131 ,
		_w27915_,
		_w32627_
	);
	LUT2 #(
		.INIT('h1)
	) name28581 (
		_w32626_,
		_w32627_,
		_w32628_
	);
	LUT2 #(
		.INIT('h4)
	) name28582 (
		_w29132_,
		_w31064_,
		_w32629_
	);
	LUT2 #(
		.INIT('h2)
	) name28583 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[4]/P0001 ,
		_w31064_,
		_w32630_
	);
	LUT2 #(
		.INIT('h1)
	) name28584 (
		_w32629_,
		_w32630_,
		_w32631_
	);
	LUT2 #(
		.INIT('h8)
	) name28585 (
		\core_c_dec_MFMY1_E_reg/P0001 ,
		_w4117_,
		_w32632_
	);
	LUT2 #(
		.INIT('h4)
	) name28586 (
		_w4117_,
		_w30972_,
		_w32633_
	);
	LUT2 #(
		.INIT('h1)
	) name28587 (
		_w32632_,
		_w32633_,
		_w32634_
	);
	LUT2 #(
		.INIT('h8)
	) name28588 (
		\core_c_dec_MFMY0_E_reg/P0001 ,
		_w4117_,
		_w32635_
	);
	LUT2 #(
		.INIT('h4)
	) name28589 (
		_w4117_,
		_w30976_,
		_w32636_
	);
	LUT2 #(
		.INIT('h1)
	) name28590 (
		_w32635_,
		_w32636_,
		_w32637_
	);
	LUT2 #(
		.INIT('h8)
	) name28591 (
		\core_c_dec_MFMX0_E_reg/P0001 ,
		_w4117_,
		_w32638_
	);
	LUT2 #(
		.INIT('h4)
	) name28592 (
		_w4117_,
		_w30975_,
		_w32639_
	);
	LUT2 #(
		.INIT('h8)
	) name28593 (
		_w30962_,
		_w32639_,
		_w32640_
	);
	LUT2 #(
		.INIT('h1)
	) name28594 (
		_w32638_,
		_w32640_,
		_w32641_
	);
	LUT2 #(
		.INIT('h8)
	) name28595 (
		\core_c_dec_MFAY1_E_reg/P0001 ,
		_w4117_,
		_w32642_
	);
	LUT2 #(
		.INIT('h4)
	) name28596 (
		_w4117_,
		_w30971_,
		_w32643_
	);
	LUT2 #(
		.INIT('h8)
	) name28597 (
		_w30977_,
		_w32643_,
		_w32644_
	);
	LUT2 #(
		.INIT('h1)
	) name28598 (
		_w32642_,
		_w32644_,
		_w32645_
	);
	LUT2 #(
		.INIT('h8)
	) name28599 (
		\core_c_dec_MFAY0_E_reg/P0001 ,
		_w4117_,
		_w32646_
	);
	LUT2 #(
		.INIT('h8)
	) name28600 (
		_w30977_,
		_w32639_,
		_w32647_
	);
	LUT2 #(
		.INIT('h1)
	) name28601 (
		_w32646_,
		_w32647_,
		_w32648_
	);
	LUT2 #(
		.INIT('h4)
	) name28602 (
		_w30497_,
		_w31064_,
		_w32649_
	);
	LUT2 #(
		.INIT('h2)
	) name28603 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[3]/P0001 ,
		_w31064_,
		_w32650_
	);
	LUT2 #(
		.INIT('h1)
	) name28604 (
		_w32649_,
		_w32650_,
		_w32651_
	);
	LUT2 #(
		.INIT('h8)
	) name28605 (
		_w31857_,
		_w31866_,
		_w32652_
	);
	LUT2 #(
		.INIT('h1)
	) name28606 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[1]/NET0131 ,
		_w32653_
	);
	LUT2 #(
		.INIT('h1)
	) name28607 (
		\sport0_rxctl_Wcnt_reg[2]/NET0131 ,
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		_w32654_
	);
	LUT2 #(
		.INIT('h8)
	) name28608 (
		_w32653_,
		_w32654_,
		_w32655_
	);
	LUT2 #(
		.INIT('h8)
	) name28609 (
		_w20430_,
		_w32655_,
		_w32656_
	);
	LUT2 #(
		.INIT('h8)
	) name28610 (
		_w32652_,
		_w32656_,
		_w32657_
	);
	LUT2 #(
		.INIT('h1)
	) name28611 (
		_w31862_,
		_w32657_,
		_w32658_
	);
	LUT2 #(
		.INIT('h2)
	) name28612 (
		_w32652_,
		_w32656_,
		_w32659_
	);
	LUT2 #(
		.INIT('h8)
	) name28613 (
		_w32653_,
		_w32659_,
		_w32660_
	);
	LUT2 #(
		.INIT('h4)
	) name28614 (
		\sport0_rxctl_Wcnt_reg[2]/NET0131 ,
		_w32660_,
		_w32661_
	);
	LUT2 #(
		.INIT('h4)
	) name28615 (
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		_w32661_,
		_w32662_
	);
	LUT2 #(
		.INIT('h2)
	) name28616 (
		\sport0_rxctl_Wcnt_reg[4]/NET0131 ,
		_w32662_,
		_w32663_
	);
	LUT2 #(
		.INIT('h4)
	) name28617 (
		\sport0_rxctl_Wcnt_reg[4]/NET0131 ,
		_w32662_,
		_w32664_
	);
	LUT2 #(
		.INIT('h1)
	) name28618 (
		_w32663_,
		_w32664_,
		_w32665_
	);
	LUT2 #(
		.INIT('h2)
	) name28619 (
		_w32658_,
		_w32665_,
		_w32666_
	);
	LUT2 #(
		.INIT('h2)
	) name28620 (
		\sport0_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w32658_,
		_w32667_
	);
	LUT2 #(
		.INIT('h1)
	) name28621 (
		_w32666_,
		_w32667_,
		_w32668_
	);
	LUT2 #(
		.INIT('h4)
	) name28622 (
		_w28566_,
		_w31064_,
		_w32669_
	);
	LUT2 #(
		.INIT('h2)
	) name28623 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[2]/P0001 ,
		_w31064_,
		_w32670_
	);
	LUT2 #(
		.INIT('h1)
	) name28624 (
		_w32669_,
		_w32670_,
		_w32671_
	);
	LUT2 #(
		.INIT('h4)
	) name28625 (
		_w29183_,
		_w31064_,
		_w32672_
	);
	LUT2 #(
		.INIT('h2)
	) name28626 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[1]/P0001 ,
		_w31064_,
		_w32673_
	);
	LUT2 #(
		.INIT('h1)
	) name28627 (
		_w32672_,
		_w32673_,
		_w32674_
	);
	LUT2 #(
		.INIT('h1)
	) name28628 (
		\idma_IAL_reg/P0001 ,
		_w9435_,
		_w32675_
	);
	LUT2 #(
		.INIT('h4)
	) name28629 (
		\idma_IADi_reg[1]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w32676_
	);
	LUT2 #(
		.INIT('h1)
	) name28630 (
		_w32675_,
		_w32676_,
		_w32677_
	);
	LUT2 #(
		.INIT('h8)
	) name28631 (
		_w32455_,
		_w32677_,
		_w32678_
	);
	LUT2 #(
		.INIT('h1)
	) name28632 (
		\idma_DCTL_reg[1]/NET0131 ,
		_w32468_,
		_w32679_
	);
	LUT2 #(
		.INIT('h1)
	) name28633 (
		_w32469_,
		_w32679_,
		_w32680_
	);
	LUT2 #(
		.INIT('h4)
	) name28634 (
		_w32455_,
		_w32680_,
		_w32681_
	);
	LUT2 #(
		.INIT('h1)
	) name28635 (
		_w32678_,
		_w32681_,
		_w32682_
	);
	LUT2 #(
		.INIT('h4)
	) name28636 (
		_w30294_,
		_w31064_,
		_w32683_
	);
	LUT2 #(
		.INIT('h2)
	) name28637 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[14]/P0001 ,
		_w31064_,
		_w32684_
	);
	LUT2 #(
		.INIT('h1)
	) name28638 (
		_w32683_,
		_w32684_,
		_w32685_
	);
	LUT2 #(
		.INIT('h4)
	) name28639 (
		_w29674_,
		_w31064_,
		_w32686_
	);
	LUT2 #(
		.INIT('h2)
	) name28640 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[13]/P0001 ,
		_w31064_,
		_w32687_
	);
	LUT2 #(
		.INIT('h1)
	) name28641 (
		_w32686_,
		_w32687_,
		_w32688_
	);
	LUT2 #(
		.INIT('h4)
	) name28642 (
		_w30094_,
		_w31064_,
		_w32689_
	);
	LUT2 #(
		.INIT('h2)
	) name28643 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[12]/P0001 ,
		_w31064_,
		_w32690_
	);
	LUT2 #(
		.INIT('h1)
	) name28644 (
		_w32689_,
		_w32690_,
		_w32691_
	);
	LUT2 #(
		.INIT('h4)
	) name28645 (
		_w29736_,
		_w31064_,
		_w32692_
	);
	LUT2 #(
		.INIT('h2)
	) name28646 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[11]/P0001 ,
		_w31064_,
		_w32693_
	);
	LUT2 #(
		.INIT('h1)
	) name28647 (
		_w32692_,
		_w32693_,
		_w32694_
	);
	LUT2 #(
		.INIT('h4)
	) name28648 (
		_w29887_,
		_w31064_,
		_w32695_
	);
	LUT2 #(
		.INIT('h2)
	) name28649 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[10]/P0001 ,
		_w31064_,
		_w32696_
	);
	LUT2 #(
		.INIT('h1)
	) name28650 (
		_w32695_,
		_w32696_,
		_w32697_
	);
	LUT2 #(
		.INIT('h4)
	) name28651 (
		_w30547_,
		_w31064_,
		_w32698_
	);
	LUT2 #(
		.INIT('h2)
	) name28652 (
		\core_eu_ea_alu_ea_reg_arswe_DO_reg[0]/P0001 ,
		_w31064_,
		_w32699_
	);
	LUT2 #(
		.INIT('h1)
	) name28653 (
		_w32698_,
		_w32699_,
		_w32700_
	);
	LUT2 #(
		.INIT('h4)
	) name28654 (
		_w29560_,
		_w31134_,
		_w32701_
	);
	LUT2 #(
		.INIT('h2)
	) name28655 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[9]/P0001 ,
		_w31134_,
		_w32702_
	);
	LUT2 #(
		.INIT('h1)
	) name28656 (
		_w32701_,
		_w32702_,
		_w32703_
	);
	LUT2 #(
		.INIT('h4)
	) name28657 (
		_w30397_,
		_w31134_,
		_w32704_
	);
	LUT2 #(
		.INIT('h2)
	) name28658 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[8]/P0001 ,
		_w31134_,
		_w32705_
	);
	LUT2 #(
		.INIT('h1)
	) name28659 (
		_w32704_,
		_w32705_,
		_w32706_
	);
	LUT2 #(
		.INIT('h4)
	) name28660 (
		_w30191_,
		_w31134_,
		_w32707_
	);
	LUT2 #(
		.INIT('h2)
	) name28661 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[7]/P0001 ,
		_w31134_,
		_w32708_
	);
	LUT2 #(
		.INIT('h1)
	) name28662 (
		_w32707_,
		_w32708_,
		_w32709_
	);
	LUT2 #(
		.INIT('h4)
	) name28663 (
		_w28990_,
		_w31134_,
		_w32710_
	);
	LUT2 #(
		.INIT('h2)
	) name28664 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[6]/P0001 ,
		_w31134_,
		_w32711_
	);
	LUT2 #(
		.INIT('h1)
	) name28665 (
		_w32710_,
		_w32711_,
		_w32712_
	);
	LUT2 #(
		.INIT('h4)
	) name28666 (
		_w29132_,
		_w31134_,
		_w32713_
	);
	LUT2 #(
		.INIT('h2)
	) name28667 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[4]/P0001 ,
		_w31134_,
		_w32714_
	);
	LUT2 #(
		.INIT('h1)
	) name28668 (
		_w32713_,
		_w32714_,
		_w32715_
	);
	LUT2 #(
		.INIT('h4)
	) name28669 (
		_w30497_,
		_w31134_,
		_w32716_
	);
	LUT2 #(
		.INIT('h2)
	) name28670 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[3]/P0001 ,
		_w31134_,
		_w32717_
	);
	LUT2 #(
		.INIT('h1)
	) name28671 (
		_w32716_,
		_w32717_,
		_w32718_
	);
	LUT2 #(
		.INIT('h4)
	) name28672 (
		_w29042_,
		_w31134_,
		_w32719_
	);
	LUT2 #(
		.INIT('h2)
	) name28673 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[5]/P0001 ,
		_w31134_,
		_w32720_
	);
	LUT2 #(
		.INIT('h1)
	) name28674 (
		_w32719_,
		_w32720_,
		_w32721_
	);
	LUT2 #(
		.INIT('h1)
	) name28675 (
		\clkc_STDcnt_reg[8]/NET0131 ,
		_w31528_,
		_w32722_
	);
	LUT2 #(
		.INIT('h1)
	) name28676 (
		_w31521_,
		_w31529_,
		_w32723_
	);
	LUT2 #(
		.INIT('h4)
	) name28677 (
		_w32722_,
		_w32723_,
		_w32724_
	);
	LUT2 #(
		.INIT('h1)
	) name28678 (
		\clkc_STDcnt_reg[6]/NET0131 ,
		_w31526_,
		_w32725_
	);
	LUT2 #(
		.INIT('h1)
	) name28679 (
		_w31521_,
		_w31527_,
		_w32726_
	);
	LUT2 #(
		.INIT('h4)
	) name28680 (
		_w32725_,
		_w32726_,
		_w32727_
	);
	LUT2 #(
		.INIT('h1)
	) name28681 (
		\sport0_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		_w19545_,
		_w32728_
	);
	LUT2 #(
		.INIT('h2)
	) name28682 (
		_w19197_,
		_w19546_,
		_w32729_
	);
	LUT2 #(
		.INIT('h4)
	) name28683 (
		_w32728_,
		_w32729_,
		_w32730_
	);
	LUT2 #(
		.INIT('h4)
	) name28684 (
		_w28566_,
		_w31134_,
		_w32731_
	);
	LUT2 #(
		.INIT('h2)
	) name28685 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[2]/P0001 ,
		_w31134_,
		_w32732_
	);
	LUT2 #(
		.INIT('h1)
	) name28686 (
		_w32731_,
		_w32732_,
		_w32733_
	);
	LUT2 #(
		.INIT('h1)
	) name28687 (
		\sport1_cfg_SCLKi_cnt_reg[8]/NET0131 ,
		_w20237_,
		_w32734_
	);
	LUT2 #(
		.INIT('h2)
	) name28688 (
		_w19130_,
		_w20238_,
		_w32735_
	);
	LUT2 #(
		.INIT('h4)
	) name28689 (
		_w32734_,
		_w32735_,
		_w32736_
	);
	LUT2 #(
		.INIT('h4)
	) name28690 (
		_w29183_,
		_w31134_,
		_w32737_
	);
	LUT2 #(
		.INIT('h2)
	) name28691 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[1]/P0001 ,
		_w31134_,
		_w32738_
	);
	LUT2 #(
		.INIT('h1)
	) name28692 (
		_w32737_,
		_w32738_,
		_w32739_
	);
	LUT2 #(
		.INIT('h4)
	) name28693 (
		_w30294_,
		_w31134_,
		_w32740_
	);
	LUT2 #(
		.INIT('h2)
	) name28694 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[14]/P0001 ,
		_w31134_,
		_w32741_
	);
	LUT2 #(
		.INIT('h1)
	) name28695 (
		_w32740_,
		_w32741_,
		_w32742_
	);
	LUT2 #(
		.INIT('h4)
	) name28696 (
		_w29674_,
		_w31134_,
		_w32743_
	);
	LUT2 #(
		.INIT('h2)
	) name28697 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[13]/P0001 ,
		_w31134_,
		_w32744_
	);
	LUT2 #(
		.INIT('h1)
	) name28698 (
		_w32743_,
		_w32744_,
		_w32745_
	);
	LUT2 #(
		.INIT('h4)
	) name28699 (
		_w30094_,
		_w31134_,
		_w32746_
	);
	LUT2 #(
		.INIT('h2)
	) name28700 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[12]/P0001 ,
		_w31134_,
		_w32747_
	);
	LUT2 #(
		.INIT('h1)
	) name28701 (
		_w32746_,
		_w32747_,
		_w32748_
	);
	LUT2 #(
		.INIT('h4)
	) name28702 (
		_w29736_,
		_w31134_,
		_w32749_
	);
	LUT2 #(
		.INIT('h2)
	) name28703 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[11]/P0001 ,
		_w31134_,
		_w32750_
	);
	LUT2 #(
		.INIT('h1)
	) name28704 (
		_w32749_,
		_w32750_,
		_w32751_
	);
	LUT2 #(
		.INIT('h4)
	) name28705 (
		_w29887_,
		_w31134_,
		_w32752_
	);
	LUT2 #(
		.INIT('h2)
	) name28706 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[10]/P0001 ,
		_w31134_,
		_w32753_
	);
	LUT2 #(
		.INIT('h1)
	) name28707 (
		_w32752_,
		_w32753_,
		_w32754_
	);
	LUT2 #(
		.INIT('h4)
	) name28708 (
		_w30547_,
		_w31134_,
		_w32755_
	);
	LUT2 #(
		.INIT('h2)
	) name28709 (
		\core_eu_ea_alu_ea_reg_arrwe_DO_reg[0]/P0001 ,
		_w31134_,
		_w32756_
	);
	LUT2 #(
		.INIT('h1)
	) name28710 (
		_w32755_,
		_w32756_,
		_w32757_
	);
	LUT2 #(
		.INIT('h8)
	) name28711 (
		\bdma_BCTL_reg[3]/NET0131 ,
		_w13757_,
		_w32758_
	);
	LUT2 #(
		.INIT('h1)
	) name28712 (
		\bdma_BRST_s2_reg/NET0131 ,
		\sice_IRST_syn_reg/P0001 ,
		_w32759_
	);
	LUT2 #(
		.INIT('h4)
	) name28713 (
		_w32758_,
		_w32759_,
		_w32760_
	);
	LUT2 #(
		.INIT('h8)
	) name28714 (
		_w10911_,
		_w32048_,
		_w32761_
	);
	LUT2 #(
		.INIT('h2)
	) name28715 (
		_w10638_,
		_w32048_,
		_w32762_
	);
	LUT2 #(
		.INIT('h2)
	) name28716 (
		_w32068_,
		_w32761_,
		_w32763_
	);
	LUT2 #(
		.INIT('h4)
	) name28717 (
		_w32762_,
		_w32763_,
		_w32764_
	);
	LUT2 #(
		.INIT('h4)
	) name28718 (
		_w10663_,
		_w32048_,
		_w32765_
	);
	LUT2 #(
		.INIT('h1)
	) name28719 (
		_w10343_,
		_w32048_,
		_w32766_
	);
	LUT2 #(
		.INIT('h1)
	) name28720 (
		_w32068_,
		_w32765_,
		_w32767_
	);
	LUT2 #(
		.INIT('h4)
	) name28721 (
		_w32766_,
		_w32767_,
		_w32768_
	);
	LUT2 #(
		.INIT('h1)
	) name28722 (
		_w32764_,
		_w32768_,
		_w32769_
	);
	LUT2 #(
		.INIT('h2)
	) name28723 (
		_w32054_,
		_w32769_,
		_w32770_
	);
	LUT2 #(
		.INIT('h1)
	) name28724 (
		_w10324_,
		_w32048_,
		_w32771_
	);
	LUT2 #(
		.INIT('h4)
	) name28725 (
		_w10356_,
		_w32058_,
		_w32772_
	);
	LUT2 #(
		.INIT('h1)
	) name28726 (
		_w10367_,
		_w32772_,
		_w32773_
	);
	LUT2 #(
		.INIT('h2)
	) name28727 (
		_w32048_,
		_w32773_,
		_w32774_
	);
	LUT2 #(
		.INIT('h1)
	) name28728 (
		_w32068_,
		_w32774_,
		_w32775_
	);
	LUT2 #(
		.INIT('h4)
	) name28729 (
		_w32771_,
		_w32775_,
		_w32776_
	);
	LUT2 #(
		.INIT('h1)
	) name28730 (
		_w10414_,
		_w32048_,
		_w32777_
	);
	LUT2 #(
		.INIT('h4)
	) name28731 (
		_w10384_,
		_w32048_,
		_w32778_
	);
	LUT2 #(
		.INIT('h2)
	) name28732 (
		_w32068_,
		_w32777_,
		_w32779_
	);
	LUT2 #(
		.INIT('h4)
	) name28733 (
		_w32778_,
		_w32779_,
		_w32780_
	);
	LUT2 #(
		.INIT('h1)
	) name28734 (
		_w32776_,
		_w32780_,
		_w32781_
	);
	LUT2 #(
		.INIT('h1)
	) name28735 (
		_w32054_,
		_w32781_,
		_w32782_
	);
	LUT2 #(
		.INIT('h1)
	) name28736 (
		_w32770_,
		_w32782_,
		_w32783_
	);
	LUT2 #(
		.INIT('h8)
	) name28737 (
		_w11265_,
		_w32048_,
		_w32784_
	);
	LUT2 #(
		.INIT('h2)
	) name28738 (
		_w11525_,
		_w32048_,
		_w32785_
	);
	LUT2 #(
		.INIT('h2)
	) name28739 (
		_w32068_,
		_w32784_,
		_w32786_
	);
	LUT2 #(
		.INIT('h4)
	) name28740 (
		_w32785_,
		_w32786_,
		_w32787_
	);
	LUT2 #(
		.INIT('h4)
	) name28741 (
		_w10954_,
		_w32048_,
		_w32788_
	);
	LUT2 #(
		.INIT('h1)
	) name28742 (
		_w11280_,
		_w32048_,
		_w32789_
	);
	LUT2 #(
		.INIT('h1)
	) name28743 (
		_w32068_,
		_w32788_,
		_w32790_
	);
	LUT2 #(
		.INIT('h4)
	) name28744 (
		_w32789_,
		_w32790_,
		_w32791_
	);
	LUT2 #(
		.INIT('h1)
	) name28745 (
		_w32787_,
		_w32791_,
		_w32792_
	);
	LUT2 #(
		.INIT('h2)
	) name28746 (
		_w32054_,
		_w32792_,
		_w32793_
	);
	LUT2 #(
		.INIT('h1)
	) name28747 (
		_w11579_,
		_w32048_,
		_w32794_
	);
	LUT2 #(
		.INIT('h4)
	) name28748 (
		_w11540_,
		_w32058_,
		_w32795_
	);
	LUT2 #(
		.INIT('h1)
	) name28749 (
		_w11551_,
		_w32795_,
		_w32796_
	);
	LUT2 #(
		.INIT('h2)
	) name28750 (
		_w32048_,
		_w32796_,
		_w32797_
	);
	LUT2 #(
		.INIT('h1)
	) name28751 (
		_w32068_,
		_w32797_,
		_w32798_
	);
	LUT2 #(
		.INIT('h4)
	) name28752 (
		_w32794_,
		_w32798_,
		_w32799_
	);
	LUT2 #(
		.INIT('h1)
	) name28753 (
		_w10994_,
		_w32048_,
		_w32800_
	);
	LUT2 #(
		.INIT('h4)
	) name28754 (
		_w11023_,
		_w32048_,
		_w32801_
	);
	LUT2 #(
		.INIT('h2)
	) name28755 (
		_w32068_,
		_w32800_,
		_w32802_
	);
	LUT2 #(
		.INIT('h4)
	) name28756 (
		_w32801_,
		_w32802_,
		_w32803_
	);
	LUT2 #(
		.INIT('h1)
	) name28757 (
		_w32799_,
		_w32803_,
		_w32804_
	);
	LUT2 #(
		.INIT('h1)
	) name28758 (
		_w32054_,
		_w32804_,
		_w32805_
	);
	LUT2 #(
		.INIT('h1)
	) name28759 (
		_w32793_,
		_w32805_,
		_w32806_
	);
	LUT2 #(
		.INIT('h8)
	) name28760 (
		_w11525_,
		_w32048_,
		_w32807_
	);
	LUT2 #(
		.INIT('h2)
	) name28761 (
		_w11265_,
		_w32048_,
		_w32808_
	);
	LUT2 #(
		.INIT('h2)
	) name28762 (
		_w32068_,
		_w32808_,
		_w32809_
	);
	LUT2 #(
		.INIT('h4)
	) name28763 (
		_w32807_,
		_w32809_,
		_w32810_
	);
	LUT2 #(
		.INIT('h1)
	) name28764 (
		_w10954_,
		_w32048_,
		_w32811_
	);
	LUT2 #(
		.INIT('h4)
	) name28765 (
		_w11280_,
		_w32048_,
		_w32812_
	);
	LUT2 #(
		.INIT('h1)
	) name28766 (
		_w32068_,
		_w32811_,
		_w32813_
	);
	LUT2 #(
		.INIT('h4)
	) name28767 (
		_w32812_,
		_w32813_,
		_w32814_
	);
	LUT2 #(
		.INIT('h1)
	) name28768 (
		_w32810_,
		_w32814_,
		_w32815_
	);
	LUT2 #(
		.INIT('h2)
	) name28769 (
		_w32054_,
		_w32815_,
		_w32816_
	);
	LUT2 #(
		.INIT('h1)
	) name28770 (
		_w10930_,
		_w32048_,
		_w32817_
	);
	LUT2 #(
		.INIT('h4)
	) name28771 (
		_w10967_,
		_w32058_,
		_w32818_
	);
	LUT2 #(
		.INIT('h1)
	) name28772 (
		_w10978_,
		_w32818_,
		_w32819_
	);
	LUT2 #(
		.INIT('h2)
	) name28773 (
		_w32048_,
		_w32819_,
		_w32820_
	);
	LUT2 #(
		.INIT('h1)
	) name28774 (
		_w32068_,
		_w32820_,
		_w32821_
	);
	LUT2 #(
		.INIT('h4)
	) name28775 (
		_w32817_,
		_w32821_,
		_w32822_
	);
	LUT2 #(
		.INIT('h1)
	) name28776 (
		_w11023_,
		_w32048_,
		_w32823_
	);
	LUT2 #(
		.INIT('h4)
	) name28777 (
		_w10994_,
		_w32048_,
		_w32824_
	);
	LUT2 #(
		.INIT('h2)
	) name28778 (
		_w32068_,
		_w32823_,
		_w32825_
	);
	LUT2 #(
		.INIT('h4)
	) name28779 (
		_w32824_,
		_w32825_,
		_w32826_
	);
	LUT2 #(
		.INIT('h1)
	) name28780 (
		_w32822_,
		_w32826_,
		_w32827_
	);
	LUT2 #(
		.INIT('h1)
	) name28781 (
		_w32054_,
		_w32827_,
		_w32828_
	);
	LUT2 #(
		.INIT('h1)
	) name28782 (
		_w32816_,
		_w32828_,
		_w32829_
	);
	LUT2 #(
		.INIT('h8)
	) name28783 (
		_w10289_,
		_w32048_,
		_w32830_
	);
	LUT2 #(
		.INIT('h2)
	) name28784 (
		_w10069_,
		_w32048_,
		_w32831_
	);
	LUT2 #(
		.INIT('h2)
	) name28785 (
		_w32068_,
		_w32830_,
		_w32832_
	);
	LUT2 #(
		.INIT('h4)
	) name28786 (
		_w32831_,
		_w32832_,
		_w32833_
	);
	LUT2 #(
		.INIT('h4)
	) name28787 (
		_w9752_,
		_w32048_,
		_w32834_
	);
	LUT2 #(
		.INIT('h1)
	) name28788 (
		_w10302_,
		_w32048_,
		_w32835_
	);
	LUT2 #(
		.INIT('h1)
	) name28789 (
		_w32068_,
		_w32834_,
		_w32836_
	);
	LUT2 #(
		.INIT('h4)
	) name28790 (
		_w32835_,
		_w32836_,
		_w32837_
	);
	LUT2 #(
		.INIT('h1)
	) name28791 (
		_w32833_,
		_w32837_,
		_w32838_
	);
	LUT2 #(
		.INIT('h2)
	) name28792 (
		_w32054_,
		_w32838_,
		_w32839_
	);
	LUT2 #(
		.INIT('h1)
	) name28793 (
		_w11720_,
		_w32048_,
		_w32840_
	);
	LUT2 #(
		.INIT('h4)
	) name28794 (
		_w11668_,
		_w32058_,
		_w32841_
	);
	LUT2 #(
		.INIT('h1)
	) name28795 (
		_w11692_,
		_w32841_,
		_w32842_
	);
	LUT2 #(
		.INIT('h2)
	) name28796 (
		_w32048_,
		_w32842_,
		_w32843_
	);
	LUT2 #(
		.INIT('h1)
	) name28797 (
		_w32068_,
		_w32843_,
		_w32844_
	);
	LUT2 #(
		.INIT('h4)
	) name28798 (
		_w32840_,
		_w32844_,
		_w32845_
	);
	LUT2 #(
		.INIT('h1)
	) name28799 (
		_w9786_,
		_w32048_,
		_w32846_
	);
	LUT2 #(
		.INIT('h4)
	) name28800 (
		_w9733_,
		_w32048_,
		_w32847_
	);
	LUT2 #(
		.INIT('h2)
	) name28801 (
		_w32068_,
		_w32846_,
		_w32848_
	);
	LUT2 #(
		.INIT('h4)
	) name28802 (
		_w32847_,
		_w32848_,
		_w32849_
	);
	LUT2 #(
		.INIT('h1)
	) name28803 (
		_w32845_,
		_w32849_,
		_w32850_
	);
	LUT2 #(
		.INIT('h1)
	) name28804 (
		_w32054_,
		_w32850_,
		_w32851_
	);
	LUT2 #(
		.INIT('h1)
	) name28805 (
		_w32839_,
		_w32851_,
		_w32852_
	);
	LUT2 #(
		.INIT('h8)
	) name28806 (
		_w7859_,
		_w32048_,
		_w32853_
	);
	LUT2 #(
		.INIT('h2)
	) name28807 (
		_w8113_,
		_w32048_,
		_w32854_
	);
	LUT2 #(
		.INIT('h2)
	) name28808 (
		_w32068_,
		_w32853_,
		_w32855_
	);
	LUT2 #(
		.INIT('h4)
	) name28809 (
		_w32854_,
		_w32855_,
		_w32856_
	);
	LUT2 #(
		.INIT('h4)
	) name28810 (
		_w7644_,
		_w32048_,
		_w32857_
	);
	LUT2 #(
		.INIT('h1)
	) name28811 (
		_w8224_,
		_w32048_,
		_w32858_
	);
	LUT2 #(
		.INIT('h1)
	) name28812 (
		_w32068_,
		_w32857_,
		_w32859_
	);
	LUT2 #(
		.INIT('h4)
	) name28813 (
		_w32858_,
		_w32859_,
		_w32860_
	);
	LUT2 #(
		.INIT('h1)
	) name28814 (
		_w32856_,
		_w32860_,
		_w32861_
	);
	LUT2 #(
		.INIT('h2)
	) name28815 (
		_w32054_,
		_w32861_,
		_w32862_
	);
	LUT2 #(
		.INIT('h1)
	) name28816 (
		_w8211_,
		_w32048_,
		_w32863_
	);
	LUT2 #(
		.INIT('h4)
	) name28817 (
		_w8121_,
		_w32058_,
		_w32864_
	);
	LUT2 #(
		.INIT('h1)
	) name28818 (
		_w8162_,
		_w32864_,
		_w32865_
	);
	LUT2 #(
		.INIT('h2)
	) name28819 (
		_w32048_,
		_w32865_,
		_w32866_
	);
	LUT2 #(
		.INIT('h1)
	) name28820 (
		_w32068_,
		_w32866_,
		_w32867_
	);
	LUT2 #(
		.INIT('h4)
	) name28821 (
		_w32863_,
		_w32867_,
		_w32868_
	);
	LUT2 #(
		.INIT('h1)
	) name28822 (
		_w8190_,
		_w32048_,
		_w32869_
	);
	LUT2 #(
		.INIT('h4)
	) name28823 (
		_w8149_,
		_w32048_,
		_w32870_
	);
	LUT2 #(
		.INIT('h2)
	) name28824 (
		_w32068_,
		_w32869_,
		_w32871_
	);
	LUT2 #(
		.INIT('h4)
	) name28825 (
		_w32870_,
		_w32871_,
		_w32872_
	);
	LUT2 #(
		.INIT('h1)
	) name28826 (
		_w32868_,
		_w32872_,
		_w32873_
	);
	LUT2 #(
		.INIT('h1)
	) name28827 (
		_w32054_,
		_w32873_,
		_w32874_
	);
	LUT2 #(
		.INIT('h1)
	) name28828 (
		_w32862_,
		_w32874_,
		_w32875_
	);
	LUT2 #(
		.INIT('h8)
	) name28829 (
		_w10638_,
		_w32048_,
		_w32876_
	);
	LUT2 #(
		.INIT('h2)
	) name28830 (
		_w10911_,
		_w32048_,
		_w32877_
	);
	LUT2 #(
		.INIT('h2)
	) name28831 (
		_w32068_,
		_w32876_,
		_w32878_
	);
	LUT2 #(
		.INIT('h4)
	) name28832 (
		_w32877_,
		_w32878_,
		_w32879_
	);
	LUT2 #(
		.INIT('h4)
	) name28833 (
		_w10343_,
		_w32048_,
		_w32880_
	);
	LUT2 #(
		.INIT('h1)
	) name28834 (
		_w10663_,
		_w32048_,
		_w32881_
	);
	LUT2 #(
		.INIT('h1)
	) name28835 (
		_w32068_,
		_w32880_,
		_w32882_
	);
	LUT2 #(
		.INIT('h4)
	) name28836 (
		_w32881_,
		_w32882_,
		_w32883_
	);
	LUT2 #(
		.INIT('h1)
	) name28837 (
		_w32879_,
		_w32883_,
		_w32884_
	);
	LUT2 #(
		.INIT('h2)
	) name28838 (
		_w32054_,
		_w32884_,
		_w32885_
	);
	LUT2 #(
		.INIT('h1)
	) name28839 (
		_w11654_,
		_w32048_,
		_w32886_
	);
	LUT2 #(
		.INIT('h4)
	) name28840 (
		_w11609_,
		_w32058_,
		_w32887_
	);
	LUT2 #(
		.INIT('h1)
	) name28841 (
		_w11620_,
		_w32887_,
		_w32888_
	);
	LUT2 #(
		.INIT('h2)
	) name28842 (
		_w32048_,
		_w32888_,
		_w32889_
	);
	LUT2 #(
		.INIT('h1)
	) name28843 (
		_w32068_,
		_w32889_,
		_w32890_
	);
	LUT2 #(
		.INIT('h4)
	) name28844 (
		_w32886_,
		_w32890_,
		_w32891_
	);
	LUT2 #(
		.INIT('h1)
	) name28845 (
		_w10384_,
		_w32048_,
		_w32892_
	);
	LUT2 #(
		.INIT('h4)
	) name28846 (
		_w10414_,
		_w32048_,
		_w32893_
	);
	LUT2 #(
		.INIT('h2)
	) name28847 (
		_w32068_,
		_w32892_,
		_w32894_
	);
	LUT2 #(
		.INIT('h4)
	) name28848 (
		_w32893_,
		_w32894_,
		_w32895_
	);
	LUT2 #(
		.INIT('h1)
	) name28849 (
		_w32891_,
		_w32895_,
		_w32896_
	);
	LUT2 #(
		.INIT('h1)
	) name28850 (
		_w32054_,
		_w32896_,
		_w32897_
	);
	LUT2 #(
		.INIT('h1)
	) name28851 (
		_w32885_,
		_w32897_,
		_w32898_
	);
	LUT2 #(
		.INIT('h8)
	) name28852 (
		_w9178_,
		_w32048_,
		_w32899_
	);
	LUT2 #(
		.INIT('h2)
	) name28853 (
		_w9435_,
		_w32048_,
		_w32900_
	);
	LUT2 #(
		.INIT('h2)
	) name28854 (
		_w32068_,
		_w32899_,
		_w32901_
	);
	LUT2 #(
		.INIT('h4)
	) name28855 (
		_w32900_,
		_w32901_,
		_w32902_
	);
	LUT2 #(
		.INIT('h1)
	) name28856 (
		_w8926_,
		_w32048_,
		_w32903_
	);
	LUT2 #(
		.INIT('h4)
	) name28857 (
		_w8962_,
		_w32048_,
		_w32904_
	);
	LUT2 #(
		.INIT('h1)
	) name28858 (
		_w32068_,
		_w32903_,
		_w32905_
	);
	LUT2 #(
		.INIT('h4)
	) name28859 (
		_w32904_,
		_w32905_,
		_w32906_
	);
	LUT2 #(
		.INIT('h1)
	) name28860 (
		_w32902_,
		_w32906_,
		_w32907_
	);
	LUT2 #(
		.INIT('h2)
	) name28861 (
		_w32054_,
		_w32907_,
		_w32908_
	);
	LUT2 #(
		.INIT('h1)
	) name28862 (
		_w8945_,
		_w32048_,
		_w32909_
	);
	LUT2 #(
		.INIT('h4)
	) name28863 (
		_w8845_,
		_w32058_,
		_w32910_
	);
	LUT2 #(
		.INIT('h1)
	) name28864 (
		_w8856_,
		_w32910_,
		_w32911_
	);
	LUT2 #(
		.INIT('h2)
	) name28865 (
		_w32048_,
		_w32911_,
		_w32912_
	);
	LUT2 #(
		.INIT('h1)
	) name28866 (
		_w32068_,
		_w32912_,
		_w32913_
	);
	LUT2 #(
		.INIT('h4)
	) name28867 (
		_w32909_,
		_w32913_,
		_w32914_
	);
	LUT2 #(
		.INIT('h1)
	) name28868 (
		_w8903_,
		_w32048_,
		_w32915_
	);
	LUT2 #(
		.INIT('h4)
	) name28869 (
		_w8873_,
		_w32048_,
		_w32916_
	);
	LUT2 #(
		.INIT('h2)
	) name28870 (
		_w32068_,
		_w32915_,
		_w32917_
	);
	LUT2 #(
		.INIT('h4)
	) name28871 (
		_w32916_,
		_w32917_,
		_w32918_
	);
	LUT2 #(
		.INIT('h1)
	) name28872 (
		_w32914_,
		_w32918_,
		_w32919_
	);
	LUT2 #(
		.INIT('h1)
	) name28873 (
		_w32054_,
		_w32919_,
		_w32920_
	);
	LUT2 #(
		.INIT('h1)
	) name28874 (
		_w32908_,
		_w32920_,
		_w32921_
	);
	LUT2 #(
		.INIT('h8)
	) name28875 (
		_w8460_,
		_w32048_,
		_w32922_
	);
	LUT2 #(
		.INIT('h2)
	) name28876 (
		_w8715_,
		_w32048_,
		_w32923_
	);
	LUT2 #(
		.INIT('h2)
	) name28877 (
		_w32068_,
		_w32922_,
		_w32924_
	);
	LUT2 #(
		.INIT('h4)
	) name28878 (
		_w32923_,
		_w32924_,
		_w32925_
	);
	LUT2 #(
		.INIT('h1)
	) name28879 (
		_w8794_,
		_w32048_,
		_w32926_
	);
	LUT2 #(
		.INIT('h4)
	) name28880 (
		_w8246_,
		_w32048_,
		_w32927_
	);
	LUT2 #(
		.INIT('h1)
	) name28881 (
		_w32068_,
		_w32926_,
		_w32928_
	);
	LUT2 #(
		.INIT('h4)
	) name28882 (
		_w32927_,
		_w32928_,
		_w32929_
	);
	LUT2 #(
		.INIT('h1)
	) name28883 (
		_w32925_,
		_w32929_,
		_w32930_
	);
	LUT2 #(
		.INIT('h2)
	) name28884 (
		_w32054_,
		_w32930_,
		_w32931_
	);
	LUT2 #(
		.INIT('h1)
	) name28885 (
		_w8813_,
		_w32048_,
		_w32932_
	);
	LUT2 #(
		.INIT('h4)
	) name28886 (
		_w8723_,
		_w32058_,
		_w32933_
	);
	LUT2 #(
		.INIT('h1)
	) name28887 (
		_w8819_,
		_w32933_,
		_w32934_
	);
	LUT2 #(
		.INIT('h2)
	) name28888 (
		_w32048_,
		_w32934_,
		_w32935_
	);
	LUT2 #(
		.INIT('h1)
	) name28889 (
		_w32068_,
		_w32935_,
		_w32936_
	);
	LUT2 #(
		.INIT('h4)
	) name28890 (
		_w32932_,
		_w32936_,
		_w32937_
	);
	LUT2 #(
		.INIT('h1)
	) name28891 (
		_w8773_,
		_w32048_,
		_w32938_
	);
	LUT2 #(
		.INIT('h4)
	) name28892 (
		_w8750_,
		_w32048_,
		_w32939_
	);
	LUT2 #(
		.INIT('h2)
	) name28893 (
		_w32068_,
		_w32938_,
		_w32940_
	);
	LUT2 #(
		.INIT('h4)
	) name28894 (
		_w32939_,
		_w32940_,
		_w32941_
	);
	LUT2 #(
		.INIT('h1)
	) name28895 (
		_w32937_,
		_w32941_,
		_w32942_
	);
	LUT2 #(
		.INIT('h1)
	) name28896 (
		_w32054_,
		_w32942_,
		_w32943_
	);
	LUT2 #(
		.INIT('h1)
	) name28897 (
		_w32931_,
		_w32943_,
		_w32944_
	);
	LUT2 #(
		.INIT('h1)
	) name28898 (
		_w24649_,
		_w32080_,
		_w32945_
	);
	LUT2 #(
		.INIT('h8)
	) name28899 (
		_w32783_,
		_w32806_,
		_w32946_
	);
	LUT2 #(
		.INIT('h8)
	) name28900 (
		_w32829_,
		_w32898_,
		_w32947_
	);
	LUT2 #(
		.INIT('h8)
	) name28901 (
		_w32921_,
		_w32944_,
		_w32948_
	);
	LUT2 #(
		.INIT('h8)
	) name28902 (
		_w32947_,
		_w32948_,
		_w32949_
	);
	LUT2 #(
		.INIT('h8)
	) name28903 (
		_w32945_,
		_w32946_,
		_w32950_
	);
	LUT2 #(
		.INIT('h8)
	) name28904 (
		_w32852_,
		_w32875_,
		_w32951_
	);
	LUT2 #(
		.INIT('h8)
	) name28905 (
		_w32950_,
		_w32951_,
		_w32952_
	);
	LUT2 #(
		.INIT('h8)
	) name28906 (
		_w32949_,
		_w32952_,
		_w32953_
	);
	LUT2 #(
		.INIT('h2)
	) name28907 (
		_w20386_,
		_w32465_,
		_w32954_
	);
	LUT2 #(
		.INIT('h1)
	) name28908 (
		\idma_DCTL_reg[14]/NET0131 ,
		_w32465_,
		_w32955_
	);
	LUT2 #(
		.INIT('h2)
	) name28909 (
		\idma_PM_1st_reg/NET0131 ,
		_w32955_,
		_w32956_
	);
	LUT2 #(
		.INIT('h1)
	) name28910 (
		_w32954_,
		_w32956_,
		_w32957_
	);
	LUT2 #(
		.INIT('h8)
	) name28911 (
		_w20074_,
		_w32957_,
		_w32958_
	);
	LUT2 #(
		.INIT('h2)
	) name28912 (
		_w4150_,
		_w25780_,
		_w32959_
	);
	LUT2 #(
		.INIT('h8)
	) name28913 (
		\tm_tcr_reg_DO_reg[12]/NET0131 ,
		_w20355_,
		_w32960_
	);
	LUT2 #(
		.INIT('h4)
	) name28914 (
		\tm_tpr_reg_DO_reg[12]/NET0131 ,
		_w22400_,
		_w32961_
	);
	LUT2 #(
		.INIT('h2)
	) name28915 (
		\tm_TCR_TMP_reg[12]/NET0131 ,
		_w25839_,
		_w32962_
	);
	LUT2 #(
		.INIT('h1)
	) name28916 (
		_w22400_,
		_w25840_,
		_w32963_
	);
	LUT2 #(
		.INIT('h4)
	) name28917 (
		_w32962_,
		_w32963_,
		_w32964_
	);
	LUT2 #(
		.INIT('h1)
	) name28918 (
		_w20355_,
		_w32961_,
		_w32965_
	);
	LUT2 #(
		.INIT('h4)
	) name28919 (
		_w32964_,
		_w32965_,
		_w32966_
	);
	LUT2 #(
		.INIT('h1)
	) name28920 (
		_w32960_,
		_w32966_,
		_w32967_
	);
	LUT2 #(
		.INIT('h2)
	) name28921 (
		\sport1_rxctl_LMcnt_reg[4]/NET0131 ,
		_w30753_,
		_w32968_
	);
	LUT2 #(
		.INIT('h2)
	) name28922 (
		_w31705_,
		_w32968_,
		_w32969_
	);
	LUT2 #(
		.INIT('h2)
	) name28923 (
		\sport0_rxctl_LMcnt_reg[4]/NET0131 ,
		_w30777_,
		_w32970_
	);
	LUT2 #(
		.INIT('h2)
	) name28924 (
		_w31868_,
		_w32970_,
		_w32971_
	);
	LUT2 #(
		.INIT('h2)
	) name28925 (
		_w4055_,
		_w6033_,
		_w32972_
	);
	LUT2 #(
		.INIT('h8)
	) name28926 (
		_w5692_,
		_w5974_,
		_w32973_
	);
	LUT2 #(
		.INIT('h4)
	) name28927 (
		_w32972_,
		_w32973_,
		_w32974_
	);
	LUT2 #(
		.INIT('h1)
	) name28928 (
		\core_dag_ilm2reg_IL_E_reg[1]/P0001 ,
		_w5692_,
		_w32975_
	);
	LUT2 #(
		.INIT('h1)
	) name28929 (
		_w32974_,
		_w32975_,
		_w32976_
	);
	LUT2 #(
		.INIT('h2)
	) name28930 (
		_w4055_,
		_w6036_,
		_w32977_
	);
	LUT2 #(
		.INIT('h8)
	) name28931 (
		_w5692_,
		_w5989_,
		_w32978_
	);
	LUT2 #(
		.INIT('h4)
	) name28932 (
		_w32977_,
		_w32978_,
		_w32979_
	);
	LUT2 #(
		.INIT('h1)
	) name28933 (
		\core_dag_ilm2reg_IL_E_reg[0]/P0001 ,
		_w5692_,
		_w32980_
	);
	LUT2 #(
		.INIT('h1)
	) name28934 (
		_w32979_,
		_w32980_,
		_w32981_
	);
	LUT2 #(
		.INIT('h4)
	) name28935 (
		_w32976_,
		_w32981_,
		_w32982_
	);
	LUT2 #(
		.INIT('h8)
	) name28936 (
		_w25955_,
		_w32982_,
		_w32983_
	);
	LUT2 #(
		.INIT('h2)
	) name28937 (
		_w32976_,
		_w32981_,
		_w32984_
	);
	LUT2 #(
		.INIT('h8)
	) name28938 (
		_w25965_,
		_w32984_,
		_w32985_
	);
	LUT2 #(
		.INIT('h1)
	) name28939 (
		_w32976_,
		_w32981_,
		_w32986_
	);
	LUT2 #(
		.INIT('h8)
	) name28940 (
		_w25954_,
		_w32986_,
		_w32987_
	);
	LUT2 #(
		.INIT('h8)
	) name28941 (
		_w32976_,
		_w32981_,
		_w32988_
	);
	LUT2 #(
		.INIT('h8)
	) name28942 (
		_w25959_,
		_w32988_,
		_w32989_
	);
	LUT2 #(
		.INIT('h1)
	) name28943 (
		_w32983_,
		_w32985_,
		_w32990_
	);
	LUT2 #(
		.INIT('h1)
	) name28944 (
		_w32987_,
		_w32989_,
		_w32991_
	);
	LUT2 #(
		.INIT('h8)
	) name28945 (
		_w32990_,
		_w32991_,
		_w32992_
	);
	LUT2 #(
		.INIT('h2)
	) name28946 (
		_w11265_,
		_w32992_,
		_w32993_
	);
	LUT2 #(
		.INIT('h4)
	) name28947 (
		_w25965_,
		_w32984_,
		_w32994_
	);
	LUT2 #(
		.INIT('h8)
	) name28948 (
		\core_dag_ilm2reg_L6_we_DO_reg[7]/NET0131 ,
		_w32994_,
		_w32995_
	);
	LUT2 #(
		.INIT('h4)
	) name28949 (
		_w25954_,
		_w32986_,
		_w32996_
	);
	LUT2 #(
		.INIT('h8)
	) name28950 (
		\core_dag_ilm2reg_L4_we_DO_reg[7]/NET0131 ,
		_w32996_,
		_w32997_
	);
	LUT2 #(
		.INIT('h4)
	) name28951 (
		_w25959_,
		_w32988_,
		_w32998_
	);
	LUT2 #(
		.INIT('h8)
	) name28952 (
		\core_dag_ilm2reg_L7_we_DO_reg[7]/NET0131 ,
		_w32998_,
		_w32999_
	);
	LUT2 #(
		.INIT('h4)
	) name28953 (
		_w25955_,
		_w32982_,
		_w33000_
	);
	LUT2 #(
		.INIT('h8)
	) name28954 (
		\core_dag_ilm2reg_L5_we_DO_reg[7]/NET0131 ,
		_w33000_,
		_w33001_
	);
	LUT2 #(
		.INIT('h1)
	) name28955 (
		_w21579_,
		_w32995_,
		_w33002_
	);
	LUT2 #(
		.INIT('h1)
	) name28956 (
		_w32997_,
		_w32999_,
		_w33003_
	);
	LUT2 #(
		.INIT('h4)
	) name28957 (
		_w33001_,
		_w33003_,
		_w33004_
	);
	LUT2 #(
		.INIT('h8)
	) name28958 (
		_w33002_,
		_w33004_,
		_w33005_
	);
	LUT2 #(
		.INIT('h4)
	) name28959 (
		_w32993_,
		_w33005_,
		_w33006_
	);
	LUT2 #(
		.INIT('h4)
	) name28960 (
		\core_dag_ilm2reg_L_reg[7]/NET0131 ,
		_w21579_,
		_w33007_
	);
	LUT2 #(
		.INIT('h1)
	) name28961 (
		_w33006_,
		_w33007_,
		_w33008_
	);
	LUT2 #(
		.INIT('h2)
	) name28962 (
		_w11525_,
		_w32992_,
		_w33009_
	);
	LUT2 #(
		.INIT('h8)
	) name28963 (
		\core_dag_ilm2reg_L6_we_DO_reg[6]/NET0131 ,
		_w32994_,
		_w33010_
	);
	LUT2 #(
		.INIT('h8)
	) name28964 (
		\core_dag_ilm2reg_L4_we_DO_reg[6]/NET0131 ,
		_w32996_,
		_w33011_
	);
	LUT2 #(
		.INIT('h8)
	) name28965 (
		\core_dag_ilm2reg_L7_we_DO_reg[6]/NET0131 ,
		_w32998_,
		_w33012_
	);
	LUT2 #(
		.INIT('h8)
	) name28966 (
		\core_dag_ilm2reg_L5_we_DO_reg[6]/NET0131 ,
		_w33000_,
		_w33013_
	);
	LUT2 #(
		.INIT('h1)
	) name28967 (
		_w21579_,
		_w33010_,
		_w33014_
	);
	LUT2 #(
		.INIT('h1)
	) name28968 (
		_w33011_,
		_w33012_,
		_w33015_
	);
	LUT2 #(
		.INIT('h4)
	) name28969 (
		_w33013_,
		_w33015_,
		_w33016_
	);
	LUT2 #(
		.INIT('h8)
	) name28970 (
		_w33014_,
		_w33016_,
		_w33017_
	);
	LUT2 #(
		.INIT('h4)
	) name28971 (
		_w33009_,
		_w33017_,
		_w33018_
	);
	LUT2 #(
		.INIT('h4)
	) name28972 (
		\core_dag_ilm2reg_L_reg[6]/NET0131 ,
		_w21579_,
		_w33019_
	);
	LUT2 #(
		.INIT('h1)
	) name28973 (
		_w33018_,
		_w33019_,
		_w33020_
	);
	LUT2 #(
		.INIT('h2)
	) name28974 (
		_w10069_,
		_w32992_,
		_w33021_
	);
	LUT2 #(
		.INIT('h8)
	) name28975 (
		\core_dag_ilm2reg_L4_we_DO_reg[4]/NET0131 ,
		_w32996_,
		_w33022_
	);
	LUT2 #(
		.INIT('h8)
	) name28976 (
		\core_dag_ilm2reg_L6_we_DO_reg[4]/NET0131 ,
		_w32994_,
		_w33023_
	);
	LUT2 #(
		.INIT('h8)
	) name28977 (
		\core_dag_ilm2reg_L5_we_DO_reg[4]/NET0131 ,
		_w33000_,
		_w33024_
	);
	LUT2 #(
		.INIT('h8)
	) name28978 (
		\core_dag_ilm2reg_L7_we_DO_reg[4]/NET0131 ,
		_w32998_,
		_w33025_
	);
	LUT2 #(
		.INIT('h1)
	) name28979 (
		_w21579_,
		_w33022_,
		_w33026_
	);
	LUT2 #(
		.INIT('h1)
	) name28980 (
		_w33023_,
		_w33024_,
		_w33027_
	);
	LUT2 #(
		.INIT('h4)
	) name28981 (
		_w33025_,
		_w33027_,
		_w33028_
	);
	LUT2 #(
		.INIT('h8)
	) name28982 (
		_w33026_,
		_w33028_,
		_w33029_
	);
	LUT2 #(
		.INIT('h4)
	) name28983 (
		_w33021_,
		_w33029_,
		_w33030_
	);
	LUT2 #(
		.INIT('h4)
	) name28984 (
		\core_dag_ilm2reg_L_reg[4]/NET0131 ,
		_w21579_,
		_w33031_
	);
	LUT2 #(
		.INIT('h1)
	) name28985 (
		_w33030_,
		_w33031_,
		_w33032_
	);
	LUT2 #(
		.INIT('h2)
	) name28986 (
		_w8113_,
		_w32992_,
		_w33033_
	);
	LUT2 #(
		.INIT('h8)
	) name28987 (
		\core_dag_ilm2reg_L6_we_DO_reg[3]/NET0131 ,
		_w32994_,
		_w33034_
	);
	LUT2 #(
		.INIT('h8)
	) name28988 (
		\core_dag_ilm2reg_L4_we_DO_reg[3]/NET0131 ,
		_w32996_,
		_w33035_
	);
	LUT2 #(
		.INIT('h8)
	) name28989 (
		\core_dag_ilm2reg_L7_we_DO_reg[3]/NET0131 ,
		_w32998_,
		_w33036_
	);
	LUT2 #(
		.INIT('h8)
	) name28990 (
		\core_dag_ilm2reg_L5_we_DO_reg[3]/NET0131 ,
		_w33000_,
		_w33037_
	);
	LUT2 #(
		.INIT('h1)
	) name28991 (
		_w21579_,
		_w33034_,
		_w33038_
	);
	LUT2 #(
		.INIT('h1)
	) name28992 (
		_w33035_,
		_w33036_,
		_w33039_
	);
	LUT2 #(
		.INIT('h4)
	) name28993 (
		_w33037_,
		_w33039_,
		_w33040_
	);
	LUT2 #(
		.INIT('h8)
	) name28994 (
		_w33038_,
		_w33040_,
		_w33041_
	);
	LUT2 #(
		.INIT('h4)
	) name28995 (
		_w33033_,
		_w33041_,
		_w33042_
	);
	LUT2 #(
		.INIT('h4)
	) name28996 (
		\core_dag_ilm2reg_L_reg[3]/NET0131 ,
		_w21579_,
		_w33043_
	);
	LUT2 #(
		.INIT('h1)
	) name28997 (
		_w33042_,
		_w33043_,
		_w33044_
	);
	LUT2 #(
		.INIT('h2)
	) name28998 (
		_w8715_,
		_w32992_,
		_w33045_
	);
	LUT2 #(
		.INIT('h8)
	) name28999 (
		\core_dag_ilm2reg_L6_we_DO_reg[2]/NET0131 ,
		_w32994_,
		_w33046_
	);
	LUT2 #(
		.INIT('h8)
	) name29000 (
		\core_dag_ilm2reg_L4_we_DO_reg[2]/NET0131 ,
		_w32996_,
		_w33047_
	);
	LUT2 #(
		.INIT('h8)
	) name29001 (
		\core_dag_ilm2reg_L7_we_DO_reg[2]/NET0131 ,
		_w32998_,
		_w33048_
	);
	LUT2 #(
		.INIT('h8)
	) name29002 (
		\core_dag_ilm2reg_L5_we_DO_reg[2]/NET0131 ,
		_w33000_,
		_w33049_
	);
	LUT2 #(
		.INIT('h1)
	) name29003 (
		_w21579_,
		_w33046_,
		_w33050_
	);
	LUT2 #(
		.INIT('h1)
	) name29004 (
		_w33047_,
		_w33048_,
		_w33051_
	);
	LUT2 #(
		.INIT('h4)
	) name29005 (
		_w33049_,
		_w33051_,
		_w33052_
	);
	LUT2 #(
		.INIT('h8)
	) name29006 (
		_w33050_,
		_w33052_,
		_w33053_
	);
	LUT2 #(
		.INIT('h4)
	) name29007 (
		_w33045_,
		_w33053_,
		_w33054_
	);
	LUT2 #(
		.INIT('h4)
	) name29008 (
		\core_dag_ilm2reg_L_reg[2]/NET0131 ,
		_w21579_,
		_w33055_
	);
	LUT2 #(
		.INIT('h1)
	) name29009 (
		_w33054_,
		_w33055_,
		_w33056_
	);
	LUT2 #(
		.INIT('h2)
	) name29010 (
		_w9435_,
		_w32992_,
		_w33057_
	);
	LUT2 #(
		.INIT('h8)
	) name29011 (
		\core_dag_ilm2reg_L4_we_DO_reg[1]/NET0131 ,
		_w32996_,
		_w33058_
	);
	LUT2 #(
		.INIT('h8)
	) name29012 (
		\core_dag_ilm2reg_L6_we_DO_reg[1]/NET0131 ,
		_w32994_,
		_w33059_
	);
	LUT2 #(
		.INIT('h8)
	) name29013 (
		\core_dag_ilm2reg_L5_we_DO_reg[1]/NET0131 ,
		_w33000_,
		_w33060_
	);
	LUT2 #(
		.INIT('h8)
	) name29014 (
		\core_dag_ilm2reg_L7_we_DO_reg[1]/NET0131 ,
		_w32998_,
		_w33061_
	);
	LUT2 #(
		.INIT('h1)
	) name29015 (
		_w21579_,
		_w33058_,
		_w33062_
	);
	LUT2 #(
		.INIT('h1)
	) name29016 (
		_w33059_,
		_w33060_,
		_w33063_
	);
	LUT2 #(
		.INIT('h4)
	) name29017 (
		_w33061_,
		_w33063_,
		_w33064_
	);
	LUT2 #(
		.INIT('h8)
	) name29018 (
		_w33062_,
		_w33064_,
		_w33065_
	);
	LUT2 #(
		.INIT('h4)
	) name29019 (
		_w33057_,
		_w33065_,
		_w33066_
	);
	LUT2 #(
		.INIT('h4)
	) name29020 (
		\core_dag_ilm2reg_L_reg[1]/NET0131 ,
		_w21579_,
		_w33067_
	);
	LUT2 #(
		.INIT('h1)
	) name29021 (
		_w33066_,
		_w33067_,
		_w33068_
	);
	LUT2 #(
		.INIT('h2)
	) name29022 (
		_w7607_,
		_w32992_,
		_w33069_
	);
	LUT2 #(
		.INIT('h8)
	) name29023 (
		\core_dag_ilm2reg_L6_we_DO_reg[0]/NET0131 ,
		_w32994_,
		_w33070_
	);
	LUT2 #(
		.INIT('h8)
	) name29024 (
		\core_dag_ilm2reg_L4_we_DO_reg[0]/NET0131 ,
		_w32996_,
		_w33071_
	);
	LUT2 #(
		.INIT('h8)
	) name29025 (
		\core_dag_ilm2reg_L7_we_DO_reg[0]/NET0131 ,
		_w32998_,
		_w33072_
	);
	LUT2 #(
		.INIT('h8)
	) name29026 (
		\core_dag_ilm2reg_L5_we_DO_reg[0]/NET0131 ,
		_w33000_,
		_w33073_
	);
	LUT2 #(
		.INIT('h1)
	) name29027 (
		_w21579_,
		_w33070_,
		_w33074_
	);
	LUT2 #(
		.INIT('h1)
	) name29028 (
		_w33071_,
		_w33072_,
		_w33075_
	);
	LUT2 #(
		.INIT('h4)
	) name29029 (
		_w33073_,
		_w33075_,
		_w33076_
	);
	LUT2 #(
		.INIT('h8)
	) name29030 (
		_w33074_,
		_w33076_,
		_w33077_
	);
	LUT2 #(
		.INIT('h4)
	) name29031 (
		_w33069_,
		_w33077_,
		_w33078_
	);
	LUT2 #(
		.INIT('h4)
	) name29032 (
		\core_dag_ilm2reg_L_reg[0]/NET0131 ,
		_w21579_,
		_w33079_
	);
	LUT2 #(
		.INIT('h1)
	) name29033 (
		_w33078_,
		_w33079_,
		_w33080_
	);
	LUT2 #(
		.INIT('h1)
	) name29034 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		_w5692_,
		_w33081_
	);
	LUT2 #(
		.INIT('h8)
	) name29035 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w4055_,
		_w33082_
	);
	LUT2 #(
		.INIT('h2)
	) name29036 (
		_w32973_,
		_w33082_,
		_w33083_
	);
	LUT2 #(
		.INIT('h1)
	) name29037 (
		_w33081_,
		_w33083_,
		_w33084_
	);
	LUT2 #(
		.INIT('h1)
	) name29038 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w5692_,
		_w33085_
	);
	LUT2 #(
		.INIT('h8)
	) name29039 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w4055_,
		_w33086_
	);
	LUT2 #(
		.INIT('h2)
	) name29040 (
		_w32978_,
		_w33086_,
		_w33087_
	);
	LUT2 #(
		.INIT('h1)
	) name29041 (
		_w33085_,
		_w33087_,
		_w33088_
	);
	LUT2 #(
		.INIT('h8)
	) name29042 (
		_w33084_,
		_w33088_,
		_w33089_
	);
	LUT2 #(
		.INIT('h8)
	) name29043 (
		_w25976_,
		_w33089_,
		_w33090_
	);
	LUT2 #(
		.INIT('h1)
	) name29044 (
		_w33084_,
		_w33088_,
		_w33091_
	);
	LUT2 #(
		.INIT('h8)
	) name29045 (
		_w25975_,
		_w33091_,
		_w33092_
	);
	LUT2 #(
		.INIT('h2)
	) name29046 (
		_w33084_,
		_w33088_,
		_w33093_
	);
	LUT2 #(
		.INIT('h8)
	) name29047 (
		_w25973_,
		_w33093_,
		_w33094_
	);
	LUT2 #(
		.INIT('h4)
	) name29048 (
		_w33084_,
		_w33088_,
		_w33095_
	);
	LUT2 #(
		.INIT('h8)
	) name29049 (
		_w25974_,
		_w33095_,
		_w33096_
	);
	LUT2 #(
		.INIT('h1)
	) name29050 (
		_w33090_,
		_w33092_,
		_w33097_
	);
	LUT2 #(
		.INIT('h1)
	) name29051 (
		_w33094_,
		_w33096_,
		_w33098_
	);
	LUT2 #(
		.INIT('h8)
	) name29052 (
		_w33097_,
		_w33098_,
		_w33099_
	);
	LUT2 #(
		.INIT('h2)
	) name29053 (
		_w11265_,
		_w33099_,
		_w33100_
	);
	LUT2 #(
		.INIT('h4)
	) name29054 (
		_w25976_,
		_w33089_,
		_w33101_
	);
	LUT2 #(
		.INIT('h8)
	) name29055 (
		\core_dag_ilm1reg_L3_we_DO_reg[7]/NET0131 ,
		_w33101_,
		_w33102_
	);
	LUT2 #(
		.INIT('h4)
	) name29056 (
		_w25975_,
		_w33091_,
		_w33103_
	);
	LUT2 #(
		.INIT('h8)
	) name29057 (
		\core_dag_ilm1reg_L0_we_DO_reg[7]/NET0131 ,
		_w33103_,
		_w33104_
	);
	LUT2 #(
		.INIT('h4)
	) name29058 (
		_w25974_,
		_w33095_,
		_w33105_
	);
	LUT2 #(
		.INIT('h8)
	) name29059 (
		\core_dag_ilm1reg_L1_we_DO_reg[7]/NET0131 ,
		_w33105_,
		_w33106_
	);
	LUT2 #(
		.INIT('h4)
	) name29060 (
		_w25973_,
		_w33093_,
		_w33107_
	);
	LUT2 #(
		.INIT('h8)
	) name29061 (
		\core_dag_ilm1reg_L2_we_DO_reg[7]/NET0131 ,
		_w33107_,
		_w33108_
	);
	LUT2 #(
		.INIT('h1)
	) name29062 (
		_w33102_,
		_w33104_,
		_w33109_
	);
	LUT2 #(
		.INIT('h1)
	) name29063 (
		_w33106_,
		_w33108_,
		_w33110_
	);
	LUT2 #(
		.INIT('h8)
	) name29064 (
		_w33109_,
		_w33110_,
		_w33111_
	);
	LUT2 #(
		.INIT('h4)
	) name29065 (
		_w21592_,
		_w33111_,
		_w33112_
	);
	LUT2 #(
		.INIT('h4)
	) name29066 (
		_w33100_,
		_w33112_,
		_w33113_
	);
	LUT2 #(
		.INIT('h4)
	) name29067 (
		\core_dag_ilm1reg_L_reg[7]/NET0131 ,
		_w21592_,
		_w33114_
	);
	LUT2 #(
		.INIT('h1)
	) name29068 (
		_w33113_,
		_w33114_,
		_w33115_
	);
	LUT2 #(
		.INIT('h2)
	) name29069 (
		_w11525_,
		_w33099_,
		_w33116_
	);
	LUT2 #(
		.INIT('h8)
	) name29070 (
		\core_dag_ilm1reg_L1_we_DO_reg[6]/NET0131 ,
		_w33105_,
		_w33117_
	);
	LUT2 #(
		.INIT('h8)
	) name29071 (
		\core_dag_ilm1reg_L2_we_DO_reg[6]/NET0131 ,
		_w33107_,
		_w33118_
	);
	LUT2 #(
		.INIT('h8)
	) name29072 (
		\core_dag_ilm1reg_L3_we_DO_reg[6]/NET0131 ,
		_w33101_,
		_w33119_
	);
	LUT2 #(
		.INIT('h8)
	) name29073 (
		\core_dag_ilm1reg_L0_we_DO_reg[6]/NET0131 ,
		_w33103_,
		_w33120_
	);
	LUT2 #(
		.INIT('h1)
	) name29074 (
		_w33117_,
		_w33118_,
		_w33121_
	);
	LUT2 #(
		.INIT('h1)
	) name29075 (
		_w33119_,
		_w33120_,
		_w33122_
	);
	LUT2 #(
		.INIT('h8)
	) name29076 (
		_w33121_,
		_w33122_,
		_w33123_
	);
	LUT2 #(
		.INIT('h4)
	) name29077 (
		_w21592_,
		_w33123_,
		_w33124_
	);
	LUT2 #(
		.INIT('h4)
	) name29078 (
		_w33116_,
		_w33124_,
		_w33125_
	);
	LUT2 #(
		.INIT('h4)
	) name29079 (
		\core_dag_ilm1reg_L_reg[6]/NET0131 ,
		_w21592_,
		_w33126_
	);
	LUT2 #(
		.INIT('h1)
	) name29080 (
		_w33125_,
		_w33126_,
		_w33127_
	);
	LUT2 #(
		.INIT('h2)
	) name29081 (
		_w10911_,
		_w33099_,
		_w33128_
	);
	LUT2 #(
		.INIT('h8)
	) name29082 (
		\core_dag_ilm1reg_L1_we_DO_reg[5]/NET0131 ,
		_w33105_,
		_w33129_
	);
	LUT2 #(
		.INIT('h8)
	) name29083 (
		\core_dag_ilm1reg_L2_we_DO_reg[5]/NET0131 ,
		_w33107_,
		_w33130_
	);
	LUT2 #(
		.INIT('h8)
	) name29084 (
		\core_dag_ilm1reg_L3_we_DO_reg[5]/NET0131 ,
		_w33101_,
		_w33131_
	);
	LUT2 #(
		.INIT('h8)
	) name29085 (
		\core_dag_ilm1reg_L0_we_DO_reg[5]/NET0131 ,
		_w33103_,
		_w33132_
	);
	LUT2 #(
		.INIT('h1)
	) name29086 (
		_w33129_,
		_w33130_,
		_w33133_
	);
	LUT2 #(
		.INIT('h1)
	) name29087 (
		_w33131_,
		_w33132_,
		_w33134_
	);
	LUT2 #(
		.INIT('h8)
	) name29088 (
		_w33133_,
		_w33134_,
		_w33135_
	);
	LUT2 #(
		.INIT('h4)
	) name29089 (
		_w21592_,
		_w33135_,
		_w33136_
	);
	LUT2 #(
		.INIT('h4)
	) name29090 (
		_w33128_,
		_w33136_,
		_w33137_
	);
	LUT2 #(
		.INIT('h4)
	) name29091 (
		\core_dag_ilm1reg_L_reg[5]/NET0131 ,
		_w21592_,
		_w33138_
	);
	LUT2 #(
		.INIT('h1)
	) name29092 (
		_w33137_,
		_w33138_,
		_w33139_
	);
	LUT2 #(
		.INIT('h2)
	) name29093 (
		_w10069_,
		_w33099_,
		_w33140_
	);
	LUT2 #(
		.INIT('h8)
	) name29094 (
		\core_dag_ilm1reg_L1_we_DO_reg[4]/NET0131 ,
		_w33105_,
		_w33141_
	);
	LUT2 #(
		.INIT('h8)
	) name29095 (
		\core_dag_ilm1reg_L2_we_DO_reg[4]/NET0131 ,
		_w33107_,
		_w33142_
	);
	LUT2 #(
		.INIT('h8)
	) name29096 (
		\core_dag_ilm1reg_L3_we_DO_reg[4]/NET0131 ,
		_w33101_,
		_w33143_
	);
	LUT2 #(
		.INIT('h8)
	) name29097 (
		\core_dag_ilm1reg_L0_we_DO_reg[4]/NET0131 ,
		_w33103_,
		_w33144_
	);
	LUT2 #(
		.INIT('h1)
	) name29098 (
		_w33141_,
		_w33142_,
		_w33145_
	);
	LUT2 #(
		.INIT('h1)
	) name29099 (
		_w33143_,
		_w33144_,
		_w33146_
	);
	LUT2 #(
		.INIT('h8)
	) name29100 (
		_w33145_,
		_w33146_,
		_w33147_
	);
	LUT2 #(
		.INIT('h4)
	) name29101 (
		_w21592_,
		_w33147_,
		_w33148_
	);
	LUT2 #(
		.INIT('h4)
	) name29102 (
		_w33140_,
		_w33148_,
		_w33149_
	);
	LUT2 #(
		.INIT('h4)
	) name29103 (
		\core_dag_ilm1reg_L_reg[4]/NET0131 ,
		_w21592_,
		_w33150_
	);
	LUT2 #(
		.INIT('h1)
	) name29104 (
		_w33149_,
		_w33150_,
		_w33151_
	);
	LUT2 #(
		.INIT('h2)
	) name29105 (
		_w8113_,
		_w33099_,
		_w33152_
	);
	LUT2 #(
		.INIT('h8)
	) name29106 (
		\core_dag_ilm1reg_L1_we_DO_reg[3]/NET0131 ,
		_w33105_,
		_w33153_
	);
	LUT2 #(
		.INIT('h8)
	) name29107 (
		\core_dag_ilm1reg_L2_we_DO_reg[3]/NET0131 ,
		_w33107_,
		_w33154_
	);
	LUT2 #(
		.INIT('h8)
	) name29108 (
		\core_dag_ilm1reg_L3_we_DO_reg[3]/NET0131 ,
		_w33101_,
		_w33155_
	);
	LUT2 #(
		.INIT('h8)
	) name29109 (
		\core_dag_ilm1reg_L0_we_DO_reg[3]/NET0131 ,
		_w33103_,
		_w33156_
	);
	LUT2 #(
		.INIT('h1)
	) name29110 (
		_w33153_,
		_w33154_,
		_w33157_
	);
	LUT2 #(
		.INIT('h1)
	) name29111 (
		_w33155_,
		_w33156_,
		_w33158_
	);
	LUT2 #(
		.INIT('h8)
	) name29112 (
		_w33157_,
		_w33158_,
		_w33159_
	);
	LUT2 #(
		.INIT('h4)
	) name29113 (
		_w21592_,
		_w33159_,
		_w33160_
	);
	LUT2 #(
		.INIT('h4)
	) name29114 (
		_w33152_,
		_w33160_,
		_w33161_
	);
	LUT2 #(
		.INIT('h4)
	) name29115 (
		\core_dag_ilm1reg_L_reg[3]/NET0131 ,
		_w21592_,
		_w33162_
	);
	LUT2 #(
		.INIT('h1)
	) name29116 (
		_w33161_,
		_w33162_,
		_w33163_
	);
	LUT2 #(
		.INIT('h2)
	) name29117 (
		_w8715_,
		_w33099_,
		_w33164_
	);
	LUT2 #(
		.INIT('h8)
	) name29118 (
		\core_dag_ilm1reg_L1_we_DO_reg[2]/NET0131 ,
		_w33105_,
		_w33165_
	);
	LUT2 #(
		.INIT('h8)
	) name29119 (
		\core_dag_ilm1reg_L2_we_DO_reg[2]/NET0131 ,
		_w33107_,
		_w33166_
	);
	LUT2 #(
		.INIT('h8)
	) name29120 (
		\core_dag_ilm1reg_L3_we_DO_reg[2]/NET0131 ,
		_w33101_,
		_w33167_
	);
	LUT2 #(
		.INIT('h8)
	) name29121 (
		\core_dag_ilm1reg_L0_we_DO_reg[2]/NET0131 ,
		_w33103_,
		_w33168_
	);
	LUT2 #(
		.INIT('h1)
	) name29122 (
		_w33165_,
		_w33166_,
		_w33169_
	);
	LUT2 #(
		.INIT('h1)
	) name29123 (
		_w33167_,
		_w33168_,
		_w33170_
	);
	LUT2 #(
		.INIT('h8)
	) name29124 (
		_w33169_,
		_w33170_,
		_w33171_
	);
	LUT2 #(
		.INIT('h4)
	) name29125 (
		_w21592_,
		_w33171_,
		_w33172_
	);
	LUT2 #(
		.INIT('h4)
	) name29126 (
		_w33164_,
		_w33172_,
		_w33173_
	);
	LUT2 #(
		.INIT('h4)
	) name29127 (
		\core_dag_ilm1reg_L_reg[2]/NET0131 ,
		_w21592_,
		_w33174_
	);
	LUT2 #(
		.INIT('h1)
	) name29128 (
		_w33173_,
		_w33174_,
		_w33175_
	);
	LUT2 #(
		.INIT('h2)
	) name29129 (
		_w9435_,
		_w33099_,
		_w33176_
	);
	LUT2 #(
		.INIT('h8)
	) name29130 (
		\core_dag_ilm1reg_L3_we_DO_reg[1]/NET0131 ,
		_w33101_,
		_w33177_
	);
	LUT2 #(
		.INIT('h8)
	) name29131 (
		\core_dag_ilm1reg_L0_we_DO_reg[1]/NET0131 ,
		_w33103_,
		_w33178_
	);
	LUT2 #(
		.INIT('h8)
	) name29132 (
		\core_dag_ilm1reg_L1_we_DO_reg[1]/NET0131 ,
		_w33105_,
		_w33179_
	);
	LUT2 #(
		.INIT('h8)
	) name29133 (
		\core_dag_ilm1reg_L2_we_DO_reg[1]/NET0131 ,
		_w33107_,
		_w33180_
	);
	LUT2 #(
		.INIT('h1)
	) name29134 (
		_w33177_,
		_w33178_,
		_w33181_
	);
	LUT2 #(
		.INIT('h1)
	) name29135 (
		_w33179_,
		_w33180_,
		_w33182_
	);
	LUT2 #(
		.INIT('h8)
	) name29136 (
		_w33181_,
		_w33182_,
		_w33183_
	);
	LUT2 #(
		.INIT('h4)
	) name29137 (
		_w21592_,
		_w33183_,
		_w33184_
	);
	LUT2 #(
		.INIT('h4)
	) name29138 (
		_w33176_,
		_w33184_,
		_w33185_
	);
	LUT2 #(
		.INIT('h4)
	) name29139 (
		\core_dag_ilm1reg_L_reg[1]/NET0131 ,
		_w21592_,
		_w33186_
	);
	LUT2 #(
		.INIT('h1)
	) name29140 (
		_w33185_,
		_w33186_,
		_w33187_
	);
	LUT2 #(
		.INIT('h2)
	) name29141 (
		_w7607_,
		_w33099_,
		_w33188_
	);
	LUT2 #(
		.INIT('h8)
	) name29142 (
		\core_dag_ilm1reg_L1_we_DO_reg[0]/NET0131 ,
		_w33105_,
		_w33189_
	);
	LUT2 #(
		.INIT('h8)
	) name29143 (
		\core_dag_ilm1reg_L2_we_DO_reg[0]/NET0131 ,
		_w33107_,
		_w33190_
	);
	LUT2 #(
		.INIT('h8)
	) name29144 (
		\core_dag_ilm1reg_L3_we_DO_reg[0]/NET0131 ,
		_w33101_,
		_w33191_
	);
	LUT2 #(
		.INIT('h8)
	) name29145 (
		\core_dag_ilm1reg_L0_we_DO_reg[0]/NET0131 ,
		_w33103_,
		_w33192_
	);
	LUT2 #(
		.INIT('h1)
	) name29146 (
		_w33189_,
		_w33190_,
		_w33193_
	);
	LUT2 #(
		.INIT('h1)
	) name29147 (
		_w33191_,
		_w33192_,
		_w33194_
	);
	LUT2 #(
		.INIT('h8)
	) name29148 (
		_w33193_,
		_w33194_,
		_w33195_
	);
	LUT2 #(
		.INIT('h4)
	) name29149 (
		_w21592_,
		_w33195_,
		_w33196_
	);
	LUT2 #(
		.INIT('h4)
	) name29150 (
		_w33188_,
		_w33196_,
		_w33197_
	);
	LUT2 #(
		.INIT('h4)
	) name29151 (
		\core_dag_ilm1reg_L_reg[0]/NET0131 ,
		_w21592_,
		_w33198_
	);
	LUT2 #(
		.INIT('h1)
	) name29152 (
		_w33197_,
		_w33198_,
		_w33199_
	);
	LUT2 #(
		.INIT('h2)
	) name29153 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w19477_,
		_w33200_
	);
	LUT2 #(
		.INIT('h1)
	) name29154 (
		\core_c_psq_Iflag_reg[12]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w33201_
	);
	LUT2 #(
		.INIT('h4)
	) name29155 (
		\core_c_psq_Iflag_reg[2]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w33202_
	);
	LUT2 #(
		.INIT('h2)
	) name29156 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w33201_,
		_w33203_
	);
	LUT2 #(
		.INIT('h4)
	) name29157 (
		_w33202_,
		_w33203_,
		_w33204_
	);
	LUT2 #(
		.INIT('h4)
	) name29158 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w33204_,
		_w33205_
	);
	LUT2 #(
		.INIT('h4)
	) name29159 (
		\core_c_psq_Iflag_reg[1]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w33206_
	);
	LUT2 #(
		.INIT('h1)
	) name29160 (
		\core_c_psq_Iflag_reg[11]/NET0131 ,
		\memc_usysr_DO_reg[11]/NET0131 ,
		_w33207_
	);
	LUT2 #(
		.INIT('h2)
	) name29161 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w33208_
	);
	LUT2 #(
		.INIT('h4)
	) name29162 (
		_w33206_,
		_w33208_,
		_w33209_
	);
	LUT2 #(
		.INIT('h4)
	) name29163 (
		_w33207_,
		_w33209_,
		_w33210_
	);
	LUT2 #(
		.INIT('h1)
	) name29164 (
		_w33205_,
		_w33210_,
		_w33211_
	);
	LUT2 #(
		.INIT('h8)
	) name29165 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		\core_c_psq_Iflag_reg[0]/NET0131 ,
		_w33212_
	);
	LUT2 #(
		.INIT('h4)
	) name29166 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w33212_,
		_w33213_
	);
	LUT2 #(
		.INIT('h1)
	) name29167 (
		_w19480_,
		_w19486_,
		_w33214_
	);
	LUT2 #(
		.INIT('h8)
	) name29168 (
		_w19495_,
		_w33214_,
		_w33215_
	);
	LUT2 #(
		.INIT('h4)
	) name29169 (
		_w19483_,
		_w33215_,
		_w33216_
	);
	LUT2 #(
		.INIT('h8)
	) name29170 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		\core_c_psq_Iflag_reg[3]/NET0131 ,
		_w33217_
	);
	LUT2 #(
		.INIT('h4)
	) name29171 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w33217_,
		_w33218_
	);
	LUT2 #(
		.INIT('h1)
	) name29172 (
		_w33213_,
		_w33218_,
		_w33219_
	);
	LUT2 #(
		.INIT('h8)
	) name29173 (
		_w33211_,
		_w33219_,
		_w33220_
	);
	LUT2 #(
		.INIT('h8)
	) name29174 (
		_w33216_,
		_w33220_,
		_w33221_
	);
	LUT2 #(
		.INIT('h4)
	) name29175 (
		\core_c_psq_PCS_reg[7]/NET0131 ,
		_w33221_,
		_w33222_
	);
	LUT2 #(
		.INIT('h1)
	) name29176 (
		_w26030_,
		_w33222_,
		_w33223_
	);
	LUT2 #(
		.INIT('h8)
	) name29177 (
		_w19477_,
		_w33223_,
		_w33224_
	);
	LUT2 #(
		.INIT('h8)
	) name29178 (
		_w11741_,
		_w33224_,
		_w33225_
	);
	LUT2 #(
		.INIT('h1)
	) name29179 (
		_w33200_,
		_w33225_,
		_w33226_
	);
	LUT2 #(
		.INIT('h2)
	) name29180 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w11525_,
		_w33227_
	);
	LUT2 #(
		.INIT('h8)
	) name29181 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001 ,
		_w14711_,
		_w33228_
	);
	LUT2 #(
		.INIT('h8)
	) name29182 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001 ,
		_w14706_,
		_w33229_
	);
	LUT2 #(
		.INIT('h8)
	) name29183 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001 ,
		_w14699_,
		_w33230_
	);
	LUT2 #(
		.INIT('h8)
	) name29184 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001 ,
		_w14704_,
		_w33231_
	);
	LUT2 #(
		.INIT('h8)
	) name29185 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][21]/P0001 ,
		_w14708_,
		_w33232_
	);
	LUT2 #(
		.INIT('h8)
	) name29186 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][21]/P0001 ,
		_w14713_,
		_w33233_
	);
	LUT2 #(
		.INIT('h8)
	) name29187 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][21]/P0001 ,
		_w14702_,
		_w33234_
	);
	LUT2 #(
		.INIT('h1)
	) name29188 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w33228_,
		_w33235_
	);
	LUT2 #(
		.INIT('h1)
	) name29189 (
		_w33229_,
		_w33230_,
		_w33236_
	);
	LUT2 #(
		.INIT('h1)
	) name29190 (
		_w33231_,
		_w33232_,
		_w33237_
	);
	LUT2 #(
		.INIT('h1)
	) name29191 (
		_w33233_,
		_w33234_,
		_w33238_
	);
	LUT2 #(
		.INIT('h8)
	) name29192 (
		_w33237_,
		_w33238_,
		_w33239_
	);
	LUT2 #(
		.INIT('h8)
	) name29193 (
		_w33235_,
		_w33236_,
		_w33240_
	);
	LUT2 #(
		.INIT('h8)
	) name29194 (
		_w33239_,
		_w33240_,
		_w33241_
	);
	LUT2 #(
		.INIT('h1)
	) name29195 (
		_w33227_,
		_w33241_,
		_w33242_
	);
	LUT2 #(
		.INIT('h8)
	) name29196 (
		_w32367_,
		_w33242_,
		_w33243_
	);
	LUT2 #(
		.INIT('h4)
	) name29197 (
		\core_c_psq_Iact_E_reg[3]/NET0131 ,
		_w32385_,
		_w33244_
	);
	LUT2 #(
		.INIT('h4)
	) name29198 (
		\core_c_psq_Iact_E_reg[4]/NET0131 ,
		_w33244_,
		_w33245_
	);
	LUT2 #(
		.INIT('h4)
	) name29199 (
		\core_c_psq_Iact_E_reg[5]/NET0131 ,
		_w33245_,
		_w33246_
	);
	LUT2 #(
		.INIT('h2)
	) name29200 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w33246_,
		_w33247_
	);
	LUT2 #(
		.INIT('h2)
	) name29201 (
		_w32364_,
		_w33247_,
		_w33248_
	);
	LUT2 #(
		.INIT('h2)
	) name29202 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w33248_,
		_w33249_
	);
	LUT2 #(
		.INIT('h4)
	) name29203 (
		_w32367_,
		_w33249_,
		_w33250_
	);
	LUT2 #(
		.INIT('h1)
	) name29204 (
		_w33243_,
		_w33250_,
		_w33251_
	);
	LUT2 #(
		.INIT('h2)
	) name29205 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w10911_,
		_w33252_
	);
	LUT2 #(
		.INIT('h8)
	) name29206 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][20]/P0001 ,
		_w14713_,
		_w33253_
	);
	LUT2 #(
		.INIT('h8)
	) name29207 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001 ,
		_w14706_,
		_w33254_
	);
	LUT2 #(
		.INIT('h8)
	) name29208 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][20]/P0001 ,
		_w14708_,
		_w33255_
	);
	LUT2 #(
		.INIT('h8)
	) name29209 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001 ,
		_w14704_,
		_w33256_
	);
	LUT2 #(
		.INIT('h8)
	) name29210 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001 ,
		_w14699_,
		_w33257_
	);
	LUT2 #(
		.INIT('h8)
	) name29211 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001 ,
		_w14711_,
		_w33258_
	);
	LUT2 #(
		.INIT('h8)
	) name29212 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][20]/P0001 ,
		_w14702_,
		_w33259_
	);
	LUT2 #(
		.INIT('h1)
	) name29213 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w33253_,
		_w33260_
	);
	LUT2 #(
		.INIT('h1)
	) name29214 (
		_w33254_,
		_w33255_,
		_w33261_
	);
	LUT2 #(
		.INIT('h1)
	) name29215 (
		_w33256_,
		_w33257_,
		_w33262_
	);
	LUT2 #(
		.INIT('h1)
	) name29216 (
		_w33258_,
		_w33259_,
		_w33263_
	);
	LUT2 #(
		.INIT('h8)
	) name29217 (
		_w33262_,
		_w33263_,
		_w33264_
	);
	LUT2 #(
		.INIT('h8)
	) name29218 (
		_w33260_,
		_w33261_,
		_w33265_
	);
	LUT2 #(
		.INIT('h8)
	) name29219 (
		_w33264_,
		_w33265_,
		_w33266_
	);
	LUT2 #(
		.INIT('h1)
	) name29220 (
		_w33252_,
		_w33266_,
		_w33267_
	);
	LUT2 #(
		.INIT('h8)
	) name29221 (
		_w32367_,
		_w33267_,
		_w33268_
	);
	LUT2 #(
		.INIT('h2)
	) name29222 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w33245_,
		_w33269_
	);
	LUT2 #(
		.INIT('h2)
	) name29223 (
		_w32364_,
		_w33269_,
		_w33270_
	);
	LUT2 #(
		.INIT('h2)
	) name29224 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w33270_,
		_w33271_
	);
	LUT2 #(
		.INIT('h4)
	) name29225 (
		_w32367_,
		_w33271_,
		_w33272_
	);
	LUT2 #(
		.INIT('h1)
	) name29226 (
		_w33268_,
		_w33272_,
		_w33273_
	);
	LUT2 #(
		.INIT('h4)
	) name29227 (
		\core_c_dec_MFPSQ_Ei_reg/NET0131 ,
		_w4117_,
		_w33274_
	);
	LUT2 #(
		.INIT('h8)
	) name29228 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w31966_,
		_w33275_
	);
	LUT2 #(
		.INIT('h8)
	) name29229 (
		_w31981_,
		_w33275_,
		_w33276_
	);
	LUT2 #(
		.INIT('h1)
	) name29230 (
		_w4117_,
		_w33276_,
		_w33277_
	);
	LUT2 #(
		.INIT('h8)
	) name29231 (
		_w31974_,
		_w33275_,
		_w33278_
	);
	LUT2 #(
		.INIT('h8)
	) name29232 (
		_w31969_,
		_w33275_,
		_w33279_
	);
	LUT2 #(
		.INIT('h4)
	) name29233 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w19270_,
		_w33280_
	);
	LUT2 #(
		.INIT('h1)
	) name29234 (
		_w31653_,
		_w33280_,
		_w33281_
	);
	LUT2 #(
		.INIT('h8)
	) name29235 (
		_w31264_,
		_w33281_,
		_w33282_
	);
	LUT2 #(
		.INIT('h8)
	) name29236 (
		_w31978_,
		_w33282_,
		_w33283_
	);
	LUT2 #(
		.INIT('h2)
	) name29237 (
		_w24442_,
		_w25244_,
		_w33284_
	);
	LUT2 #(
		.INIT('h4)
	) name29238 (
		_w32025_,
		_w33284_,
		_w33285_
	);
	LUT2 #(
		.INIT('h1)
	) name29239 (
		_w33278_,
		_w33279_,
		_w33286_
	);
	LUT2 #(
		.INIT('h4)
	) name29240 (
		_w33283_,
		_w33286_,
		_w33287_
	);
	LUT2 #(
		.INIT('h8)
	) name29241 (
		_w33277_,
		_w33285_,
		_w33288_
	);
	LUT2 #(
		.INIT('h8)
	) name29242 (
		_w33287_,
		_w33288_,
		_w33289_
	);
	LUT2 #(
		.INIT('h1)
	) name29243 (
		_w33274_,
		_w33289_,
		_w33290_
	);
	LUT2 #(
		.INIT('h8)
	) name29244 (
		_w13739_,
		_w13764_,
		_w33291_
	);
	LUT2 #(
		.INIT('h4)
	) name29245 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		_w33291_,
		_w33292_
	);
	LUT2 #(
		.INIT('h4)
	) name29246 (
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		_w33292_,
		_w33293_
	);
	LUT2 #(
		.INIT('h4)
	) name29247 (
		\bdma_BWCOUNT_reg[9]/NET0131 ,
		_w33293_,
		_w33294_
	);
	LUT2 #(
		.INIT('h4)
	) name29248 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		_w33294_,
		_w33295_
	);
	LUT2 #(
		.INIT('h4)
	) name29249 (
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		_w33295_,
		_w33296_
	);
	LUT2 #(
		.INIT('h4)
	) name29250 (
		\bdma_BWCOUNT_reg[12]/NET0131 ,
		_w33296_,
		_w33297_
	);
	LUT2 #(
		.INIT('h1)
	) name29251 (
		\bdma_BWCOUNT_reg[13]/NET0131 ,
		_w33297_,
		_w33298_
	);
	LUT2 #(
		.INIT('h8)
	) name29252 (
		\bdma_BWCOUNT_reg[13]/NET0131 ,
		_w33297_,
		_w33299_
	);
	LUT2 #(
		.INIT('h1)
	) name29253 (
		_w33298_,
		_w33299_,
		_w33300_
	);
	LUT2 #(
		.INIT('h1)
	) name29254 (
		_w13763_,
		_w33300_,
		_w33301_
	);
	LUT2 #(
		.INIT('h4)
	) name29255 (
		_w7340_,
		_w13763_,
		_w33302_
	);
	LUT2 #(
		.INIT('h1)
	) name29256 (
		_w33301_,
		_w33302_,
		_w33303_
	);
	LUT2 #(
		.INIT('h8)
	) name29257 (
		\bdma_BEAD_reg[2]/NET0131 ,
		_w20769_,
		_w33304_
	);
	LUT2 #(
		.INIT('h8)
	) name29258 (
		\bdma_BEAD_reg[3]/NET0131 ,
		_w33304_,
		_w33305_
	);
	LUT2 #(
		.INIT('h8)
	) name29259 (
		\bdma_BEAD_reg[4]/NET0131 ,
		_w33305_,
		_w33306_
	);
	LUT2 #(
		.INIT('h8)
	) name29260 (
		\bdma_BEAD_reg[5]/NET0131 ,
		_w33306_,
		_w33307_
	);
	LUT2 #(
		.INIT('h8)
	) name29261 (
		\bdma_BEAD_reg[6]/NET0131 ,
		_w33307_,
		_w33308_
	);
	LUT2 #(
		.INIT('h8)
	) name29262 (
		\bdma_BEAD_reg[7]/NET0131 ,
		_w33308_,
		_w33309_
	);
	LUT2 #(
		.INIT('h8)
	) name29263 (
		\bdma_BEAD_reg[8]/NET0131 ,
		_w33309_,
		_w33310_
	);
	LUT2 #(
		.INIT('h8)
	) name29264 (
		\bdma_BEAD_reg[9]/NET0131 ,
		_w33310_,
		_w33311_
	);
	LUT2 #(
		.INIT('h8)
	) name29265 (
		\bdma_BEAD_reg[10]/NET0131 ,
		_w33311_,
		_w33312_
	);
	LUT2 #(
		.INIT('h8)
	) name29266 (
		\bdma_BEAD_reg[11]/NET0131 ,
		_w33312_,
		_w33313_
	);
	LUT2 #(
		.INIT('h8)
	) name29267 (
		\bdma_BEAD_reg[12]/NET0131 ,
		_w33313_,
		_w33314_
	);
	LUT2 #(
		.INIT('h1)
	) name29268 (
		\bdma_BEAD_reg[12]/NET0131 ,
		_w33313_,
		_w33315_
	);
	LUT2 #(
		.INIT('h1)
	) name29269 (
		_w20765_,
		_w33314_,
		_w33316_
	);
	LUT2 #(
		.INIT('h4)
	) name29270 (
		_w33315_,
		_w33316_,
		_w33317_
	);
	LUT2 #(
		.INIT('h8)
	) name29271 (
		_w9178_,
		_w20765_,
		_w33318_
	);
	LUT2 #(
		.INIT('h1)
	) name29272 (
		_w33317_,
		_w33318_,
		_w33319_
	);
	LUT2 #(
		.INIT('h2)
	) name29273 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 ,
		_w18266_,
		_w33320_
	);
	LUT2 #(
		.INIT('h1)
	) name29274 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[0]/P0001 ,
		_w18271_,
		_w33321_
	);
	LUT2 #(
		.INIT('h2)
	) name29275 (
		_w18271_,
		_w19559_,
		_w33322_
	);
	LUT2 #(
		.INIT('h2)
	) name29276 (
		_w18273_,
		_w33321_,
		_w33323_
	);
	LUT2 #(
		.INIT('h4)
	) name29277 (
		_w33322_,
		_w33323_,
		_w33324_
	);
	LUT2 #(
		.INIT('h1)
	) name29278 (
		_w18270_,
		_w33320_,
		_w33325_
	);
	LUT2 #(
		.INIT('h4)
	) name29279 (
		_w33324_,
		_w33325_,
		_w33326_
	);
	LUT2 #(
		.INIT('h1)
	) name29280 (
		_w18262_,
		_w33326_,
		_w33327_
	);
	LUT2 #(
		.INIT('h2)
	) name29281 (
		_w18262_,
		_w19653_,
		_w33328_
	);
	LUT2 #(
		.INIT('h1)
	) name29282 (
		_w33327_,
		_w33328_,
		_w33329_
	);
	LUT2 #(
		.INIT('h8)
	) name29283 (
		_w14752_,
		_w19653_,
		_w33330_
	);
	LUT2 #(
		.INIT('h8)
	) name29284 (
		_w18328_,
		_w19559_,
		_w33331_
	);
	LUT2 #(
		.INIT('h2)
	) name29285 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[0]/P0001 ,
		_w18330_,
		_w33332_
	);
	LUT2 #(
		.INIT('h2)
	) name29286 (
		_w18334_,
		_w33332_,
		_w33333_
	);
	LUT2 #(
		.INIT('h4)
	) name29287 (
		_w33331_,
		_w33333_,
		_w33334_
	);
	LUT2 #(
		.INIT('h1)
	) name29288 (
		_w33330_,
		_w33334_,
		_w33335_
	);
	LUT2 #(
		.INIT('h2)
	) name29289 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w13778_,
		_w33336_
	);
	LUT2 #(
		.INIT('h1)
	) name29290 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w13784_,
		_w33337_
	);
	LUT2 #(
		.INIT('h1)
	) name29291 (
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		_w13777_,
		_w33338_
	);
	LUT2 #(
		.INIT('h4)
	) name29292 (
		_w27907_,
		_w33338_,
		_w33339_
	);
	LUT2 #(
		.INIT('h4)
	) name29293 (
		_w27911_,
		_w33339_,
		_w33340_
	);
	LUT2 #(
		.INIT('h1)
	) name29294 (
		_w5950_,
		_w27920_,
		_w33341_
	);
	LUT2 #(
		.INIT('h1)
	) name29295 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w33340_,
		_w33342_
	);
	LUT2 #(
		.INIT('h8)
	) name29296 (
		_w33341_,
		_w33342_,
		_w33343_
	);
	LUT2 #(
		.INIT('h1)
	) name29297 (
		_w13779_,
		_w33343_,
		_w33344_
	);
	LUT2 #(
		.INIT('h4)
	) name29298 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w13778_,
		_w33345_
	);
	LUT2 #(
		.INIT('h1)
	) name29299 (
		_w13775_,
		_w33337_,
		_w33346_
	);
	LUT2 #(
		.INIT('h4)
	) name29300 (
		_w33345_,
		_w33346_,
		_w33347_
	);
	LUT2 #(
		.INIT('h4)
	) name29301 (
		_w33344_,
		_w33347_,
		_w33348_
	);
	LUT2 #(
		.INIT('h1)
	) name29302 (
		_w33336_,
		_w33348_,
		_w33349_
	);
	LUT2 #(
		.INIT('h1)
	) name29303 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		_w33344_,
		_w33350_
	);
	LUT2 #(
		.INIT('h8)
	) name29304 (
		\core_c_psq_cntstk_ptr_reg[0]/NET0131 ,
		_w33344_,
		_w33351_
	);
	LUT2 #(
		.INIT('h1)
	) name29305 (
		_w33350_,
		_w33351_,
		_w33352_
	);
	LUT2 #(
		.INIT('h8)
	) name29306 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001 ,
		_w14711_,
		_w33353_
	);
	LUT2 #(
		.INIT('h8)
	) name29307 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001 ,
		_w14704_,
		_w33354_
	);
	LUT2 #(
		.INIT('h8)
	) name29308 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][14]/P0001 ,
		_w14708_,
		_w33355_
	);
	LUT2 #(
		.INIT('h8)
	) name29309 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][14]/P0001 ,
		_w14702_,
		_w33356_
	);
	LUT2 #(
		.INIT('h8)
	) name29310 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001 ,
		_w14699_,
		_w33357_
	);
	LUT2 #(
		.INIT('h8)
	) name29311 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001 ,
		_w14706_,
		_w33358_
	);
	LUT2 #(
		.INIT('h8)
	) name29312 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][14]/P0001 ,
		_w14713_,
		_w33359_
	);
	LUT2 #(
		.INIT('h1)
	) name29313 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w33353_,
		_w33360_
	);
	LUT2 #(
		.INIT('h1)
	) name29314 (
		_w33354_,
		_w33355_,
		_w33361_
	);
	LUT2 #(
		.INIT('h1)
	) name29315 (
		_w33356_,
		_w33357_,
		_w33362_
	);
	LUT2 #(
		.INIT('h1)
	) name29316 (
		_w33358_,
		_w33359_,
		_w33363_
	);
	LUT2 #(
		.INIT('h8)
	) name29317 (
		_w33362_,
		_w33363_,
		_w33364_
	);
	LUT2 #(
		.INIT('h8)
	) name29318 (
		_w33360_,
		_w33361_,
		_w33365_
	);
	LUT2 #(
		.INIT('h8)
	) name29319 (
		_w33364_,
		_w33365_,
		_w33366_
	);
	LUT2 #(
		.INIT('h4)
	) name29320 (
		\core_c_dec_IRE_reg[3]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w33367_
	);
	LUT2 #(
		.INIT('h2)
	) name29321 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w6071_,
		_w33368_
	);
	LUT2 #(
		.INIT('h4)
	) name29322 (
		_w33367_,
		_w33368_,
		_w33369_
	);
	LUT2 #(
		.INIT('h1)
	) name29323 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w33369_,
		_w33370_
	);
	LUT2 #(
		.INIT('h4)
	) name29324 (
		_w33366_,
		_w33370_,
		_w33371_
	);
	LUT2 #(
		.INIT('h8)
	) name29325 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w11525_,
		_w33372_
	);
	LUT2 #(
		.INIT('h1)
	) name29326 (
		_w33371_,
		_w33372_,
		_w33373_
	);
	LUT2 #(
		.INIT('h2)
	) name29327 (
		_w23243_,
		_w33373_,
		_w33374_
	);
	LUT2 #(
		.INIT('h2)
	) name29328 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w23243_,
		_w33375_
	);
	LUT2 #(
		.INIT('h1)
	) name29329 (
		_w33374_,
		_w33375_,
		_w33376_
	);
	LUT2 #(
		.INIT('h4)
	) name29330 (
		\core_c_dec_IRE_reg[15]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w33377_
	);
	LUT2 #(
		.INIT('h8)
	) name29331 (
		\core_c_dec_IRE_reg[14]/NET0131 ,
		\core_c_dec_IRE_reg[15]/NET0131 ,
		_w33378_
	);
	LUT2 #(
		.INIT('h2)
	) name29332 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w33377_,
		_w33379_
	);
	LUT2 #(
		.INIT('h4)
	) name29333 (
		_w33378_,
		_w33379_,
		_w33380_
	);
	LUT2 #(
		.INIT('h8)
	) name29334 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][13]/P0001 ,
		_w14702_,
		_w33381_
	);
	LUT2 #(
		.INIT('h8)
	) name29335 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001 ,
		_w14706_,
		_w33382_
	);
	LUT2 #(
		.INIT('h8)
	) name29336 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001 ,
		_w14711_,
		_w33383_
	);
	LUT2 #(
		.INIT('h8)
	) name29337 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][13]/P0001 ,
		_w14713_,
		_w33384_
	);
	LUT2 #(
		.INIT('h8)
	) name29338 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001 ,
		_w14699_,
		_w33385_
	);
	LUT2 #(
		.INIT('h8)
	) name29339 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][13]/P0001 ,
		_w14708_,
		_w33386_
	);
	LUT2 #(
		.INIT('h8)
	) name29340 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001 ,
		_w14704_,
		_w33387_
	);
	LUT2 #(
		.INIT('h1)
	) name29341 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w33381_,
		_w33388_
	);
	LUT2 #(
		.INIT('h1)
	) name29342 (
		_w33382_,
		_w33383_,
		_w33389_
	);
	LUT2 #(
		.INIT('h1)
	) name29343 (
		_w33384_,
		_w33385_,
		_w33390_
	);
	LUT2 #(
		.INIT('h1)
	) name29344 (
		_w33386_,
		_w33387_,
		_w33391_
	);
	LUT2 #(
		.INIT('h8)
	) name29345 (
		_w33390_,
		_w33391_,
		_w33392_
	);
	LUT2 #(
		.INIT('h8)
	) name29346 (
		_w33388_,
		_w33389_,
		_w33393_
	);
	LUT2 #(
		.INIT('h8)
	) name29347 (
		_w33392_,
		_w33393_,
		_w33394_
	);
	LUT2 #(
		.INIT('h1)
	) name29348 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w33380_,
		_w33395_
	);
	LUT2 #(
		.INIT('h4)
	) name29349 (
		_w33394_,
		_w33395_,
		_w33396_
	);
	LUT2 #(
		.INIT('h8)
	) name29350 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w10911_,
		_w33397_
	);
	LUT2 #(
		.INIT('h1)
	) name29351 (
		_w33396_,
		_w33397_,
		_w33398_
	);
	LUT2 #(
		.INIT('h2)
	) name29352 (
		_w23243_,
		_w33398_,
		_w33399_
	);
	LUT2 #(
		.INIT('h2)
	) name29353 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w23243_,
		_w33400_
	);
	LUT2 #(
		.INIT('h1)
	) name29354 (
		_w33399_,
		_w33400_,
		_w33401_
	);
	LUT2 #(
		.INIT('h4)
	) name29355 (
		\core_c_dec_IRE_reg[13]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w33402_
	);
	LUT2 #(
		.INIT('h8)
	) name29356 (
		\core_c_dec_IRE_reg[10]/NET0131 ,
		\core_c_dec_IRE_reg[13]/NET0131 ,
		_w33403_
	);
	LUT2 #(
		.INIT('h2)
	) name29357 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w33402_,
		_w33404_
	);
	LUT2 #(
		.INIT('h4)
	) name29358 (
		_w33403_,
		_w33404_,
		_w33405_
	);
	LUT2 #(
		.INIT('h8)
	) name29359 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][11]/P0001 ,
		_w14702_,
		_w33406_
	);
	LUT2 #(
		.INIT('h8)
	) name29360 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001 ,
		_w14706_,
		_w33407_
	);
	LUT2 #(
		.INIT('h8)
	) name29361 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][11]/P0001 ,
		_w14713_,
		_w33408_
	);
	LUT2 #(
		.INIT('h8)
	) name29362 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001 ,
		_w14711_,
		_w33409_
	);
	LUT2 #(
		.INIT('h8)
	) name29363 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][11]/P0001 ,
		_w14708_,
		_w33410_
	);
	LUT2 #(
		.INIT('h8)
	) name29364 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001 ,
		_w14699_,
		_w33411_
	);
	LUT2 #(
		.INIT('h8)
	) name29365 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001 ,
		_w14704_,
		_w33412_
	);
	LUT2 #(
		.INIT('h1)
	) name29366 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w33406_,
		_w33413_
	);
	LUT2 #(
		.INIT('h1)
	) name29367 (
		_w33407_,
		_w33408_,
		_w33414_
	);
	LUT2 #(
		.INIT('h1)
	) name29368 (
		_w33409_,
		_w33410_,
		_w33415_
	);
	LUT2 #(
		.INIT('h1)
	) name29369 (
		_w33411_,
		_w33412_,
		_w33416_
	);
	LUT2 #(
		.INIT('h8)
	) name29370 (
		_w33415_,
		_w33416_,
		_w33417_
	);
	LUT2 #(
		.INIT('h8)
	) name29371 (
		_w33413_,
		_w33414_,
		_w33418_
	);
	LUT2 #(
		.INIT('h8)
	) name29372 (
		_w33417_,
		_w33418_,
		_w33419_
	);
	LUT2 #(
		.INIT('h1)
	) name29373 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w33405_,
		_w33420_
	);
	LUT2 #(
		.INIT('h4)
	) name29374 (
		_w33419_,
		_w33420_,
		_w33421_
	);
	LUT2 #(
		.INIT('h8)
	) name29375 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w8113_,
		_w33422_
	);
	LUT2 #(
		.INIT('h1)
	) name29376 (
		_w33421_,
		_w33422_,
		_w33423_
	);
	LUT2 #(
		.INIT('h2)
	) name29377 (
		_w23243_,
		_w33423_,
		_w33424_
	);
	LUT2 #(
		.INIT('h2)
	) name29378 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w23243_,
		_w33425_
	);
	LUT2 #(
		.INIT('h1)
	) name29379 (
		_w33424_,
		_w33425_,
		_w33426_
	);
	LUT2 #(
		.INIT('h8)
	) name29380 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001 ,
		_w14699_,
		_w33427_
	);
	LUT2 #(
		.INIT('h8)
	) name29381 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][10]/P0001 ,
		_w14713_,
		_w33428_
	);
	LUT2 #(
		.INIT('h8)
	) name29382 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][10]/P0001 ,
		_w14702_,
		_w33429_
	);
	LUT2 #(
		.INIT('h8)
	) name29383 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001 ,
		_w14706_,
		_w33430_
	);
	LUT2 #(
		.INIT('h8)
	) name29384 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][10]/P0001 ,
		_w14708_,
		_w33431_
	);
	LUT2 #(
		.INIT('h8)
	) name29385 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001 ,
		_w14704_,
		_w33432_
	);
	LUT2 #(
		.INIT('h8)
	) name29386 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001 ,
		_w14711_,
		_w33433_
	);
	LUT2 #(
		.INIT('h1)
	) name29387 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w33427_,
		_w33434_
	);
	LUT2 #(
		.INIT('h1)
	) name29388 (
		_w33428_,
		_w33429_,
		_w33435_
	);
	LUT2 #(
		.INIT('h1)
	) name29389 (
		_w33430_,
		_w33431_,
		_w33436_
	);
	LUT2 #(
		.INIT('h1)
	) name29390 (
		_w33432_,
		_w33433_,
		_w33437_
	);
	LUT2 #(
		.INIT('h8)
	) name29391 (
		_w33436_,
		_w33437_,
		_w33438_
	);
	LUT2 #(
		.INIT('h8)
	) name29392 (
		_w33434_,
		_w33435_,
		_w33439_
	);
	LUT2 #(
		.INIT('h8)
	) name29393 (
		_w33438_,
		_w33439_,
		_w33440_
	);
	LUT2 #(
		.INIT('h4)
	) name29394 (
		\core_c_dec_IRE_reg[9]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w33441_
	);
	LUT2 #(
		.INIT('h2)
	) name29395 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w13818_,
		_w33442_
	);
	LUT2 #(
		.INIT('h4)
	) name29396 (
		_w33441_,
		_w33442_,
		_w33443_
	);
	LUT2 #(
		.INIT('h1)
	) name29397 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w33443_,
		_w33444_
	);
	LUT2 #(
		.INIT('h4)
	) name29398 (
		_w33440_,
		_w33444_,
		_w33445_
	);
	LUT2 #(
		.INIT('h8)
	) name29399 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w8715_,
		_w33446_
	);
	LUT2 #(
		.INIT('h1)
	) name29400 (
		_w33445_,
		_w33446_,
		_w33447_
	);
	LUT2 #(
		.INIT('h2)
	) name29401 (
		_w23243_,
		_w33447_,
		_w33448_
	);
	LUT2 #(
		.INIT('h2)
	) name29402 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w23243_,
		_w33449_
	);
	LUT2 #(
		.INIT('h1)
	) name29403 (
		_w33448_,
		_w33449_,
		_w33450_
	);
	LUT2 #(
		.INIT('h4)
	) name29404 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w33451_
	);
	LUT2 #(
		.INIT('h8)
	) name29405 (
		\core_c_dec_IRE_reg[5]/NET0131 ,
		\core_c_dec_IRE_reg[6]/NET0131 ,
		_w33452_
	);
	LUT2 #(
		.INIT('h2)
	) name29406 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w33451_,
		_w33453_
	);
	LUT2 #(
		.INIT('h4)
	) name29407 (
		_w33452_,
		_w33453_,
		_w33454_
	);
	LUT2 #(
		.INIT('h8)
	) name29408 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][9]/P0001 ,
		_w14702_,
		_w33455_
	);
	LUT2 #(
		.INIT('h8)
	) name29409 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001 ,
		_w14706_,
		_w33456_
	);
	LUT2 #(
		.INIT('h8)
	) name29410 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001 ,
		_w14711_,
		_w33457_
	);
	LUT2 #(
		.INIT('h8)
	) name29411 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][9]/P0001 ,
		_w14713_,
		_w33458_
	);
	LUT2 #(
		.INIT('h8)
	) name29412 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001 ,
		_w14699_,
		_w33459_
	);
	LUT2 #(
		.INIT('h8)
	) name29413 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][9]/P0001 ,
		_w14708_,
		_w33460_
	);
	LUT2 #(
		.INIT('h8)
	) name29414 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001 ,
		_w14704_,
		_w33461_
	);
	LUT2 #(
		.INIT('h1)
	) name29415 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w33455_,
		_w33462_
	);
	LUT2 #(
		.INIT('h1)
	) name29416 (
		_w33456_,
		_w33457_,
		_w33463_
	);
	LUT2 #(
		.INIT('h1)
	) name29417 (
		_w33458_,
		_w33459_,
		_w33464_
	);
	LUT2 #(
		.INIT('h1)
	) name29418 (
		_w33460_,
		_w33461_,
		_w33465_
	);
	LUT2 #(
		.INIT('h8)
	) name29419 (
		_w33464_,
		_w33465_,
		_w33466_
	);
	LUT2 #(
		.INIT('h8)
	) name29420 (
		_w33462_,
		_w33463_,
		_w33467_
	);
	LUT2 #(
		.INIT('h8)
	) name29421 (
		_w33466_,
		_w33467_,
		_w33468_
	);
	LUT2 #(
		.INIT('h1)
	) name29422 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w33454_,
		_w33469_
	);
	LUT2 #(
		.INIT('h4)
	) name29423 (
		_w33468_,
		_w33469_,
		_w33470_
	);
	LUT2 #(
		.INIT('h8)
	) name29424 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w9435_,
		_w33471_
	);
	LUT2 #(
		.INIT('h1)
	) name29425 (
		_w33470_,
		_w33471_,
		_w33472_
	);
	LUT2 #(
		.INIT('h2)
	) name29426 (
		_w23243_,
		_w33472_,
		_w33473_
	);
	LUT2 #(
		.INIT('h2)
	) name29427 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w23243_,
		_w33474_
	);
	LUT2 #(
		.INIT('h1)
	) name29428 (
		_w33473_,
		_w33474_,
		_w33475_
	);
	LUT2 #(
		.INIT('h2)
	) name29429 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w10289_,
		_w33476_
	);
	LUT2 #(
		.INIT('h8)
	) name29430 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][24]/P0001 ,
		_w14713_,
		_w33477_
	);
	LUT2 #(
		.INIT('h8)
	) name29431 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001 ,
		_w14706_,
		_w33478_
	);
	LUT2 #(
		.INIT('h8)
	) name29432 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][24]/P0001 ,
		_w14708_,
		_w33479_
	);
	LUT2 #(
		.INIT('h8)
	) name29433 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001 ,
		_w14704_,
		_w33480_
	);
	LUT2 #(
		.INIT('h8)
	) name29434 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001 ,
		_w14699_,
		_w33481_
	);
	LUT2 #(
		.INIT('h8)
	) name29435 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001 ,
		_w14711_,
		_w33482_
	);
	LUT2 #(
		.INIT('h8)
	) name29436 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][24]/P0001 ,
		_w14702_,
		_w33483_
	);
	LUT2 #(
		.INIT('h1)
	) name29437 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w33477_,
		_w33484_
	);
	LUT2 #(
		.INIT('h1)
	) name29438 (
		_w33478_,
		_w33479_,
		_w33485_
	);
	LUT2 #(
		.INIT('h1)
	) name29439 (
		_w33480_,
		_w33481_,
		_w33486_
	);
	LUT2 #(
		.INIT('h1)
	) name29440 (
		_w33482_,
		_w33483_,
		_w33487_
	);
	LUT2 #(
		.INIT('h8)
	) name29441 (
		_w33486_,
		_w33487_,
		_w33488_
	);
	LUT2 #(
		.INIT('h8)
	) name29442 (
		_w33484_,
		_w33485_,
		_w33489_
	);
	LUT2 #(
		.INIT('h8)
	) name29443 (
		_w33488_,
		_w33489_,
		_w33490_
	);
	LUT2 #(
		.INIT('h1)
	) name29444 (
		_w33476_,
		_w33490_,
		_w33491_
	);
	LUT2 #(
		.INIT('h8)
	) name29445 (
		_w32367_,
		_w33491_,
		_w33492_
	);
	LUT2 #(
		.INIT('h4)
	) name29446 (
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		_w33246_,
		_w33493_
	);
	LUT2 #(
		.INIT('h4)
	) name29447 (
		\core_c_psq_Iact_E_reg[7]/NET0131 ,
		_w33493_,
		_w33494_
	);
	LUT2 #(
		.INIT('h4)
	) name29448 (
		\core_c_psq_Iact_E_reg[8]/NET0131 ,
		_w33494_,
		_w33495_
	);
	LUT2 #(
		.INIT('h2)
	) name29449 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w33495_,
		_w33496_
	);
	LUT2 #(
		.INIT('h2)
	) name29450 (
		_w32364_,
		_w33496_,
		_w33497_
	);
	LUT2 #(
		.INIT('h2)
	) name29451 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w33497_,
		_w33498_
	);
	LUT2 #(
		.INIT('h4)
	) name29452 (
		_w32367_,
		_w33498_,
		_w33499_
	);
	LUT2 #(
		.INIT('h1)
	) name29453 (
		_w33492_,
		_w33499_,
		_w33500_
	);
	LUT2 #(
		.INIT('h2)
	) name29454 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w9435_,
		_w33501_
	);
	LUT2 #(
		.INIT('h8)
	) name29455 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][16]/P0001 ,
		_w14708_,
		_w33502_
	);
	LUT2 #(
		.INIT('h8)
	) name29456 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][16]/P0001 ,
		_w14713_,
		_w33503_
	);
	LUT2 #(
		.INIT('h8)
	) name29457 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001 ,
		_w14711_,
		_w33504_
	);
	LUT2 #(
		.INIT('h8)
	) name29458 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001 ,
		_w14699_,
		_w33505_
	);
	LUT2 #(
		.INIT('h8)
	) name29459 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001 ,
		_w14704_,
		_w33506_
	);
	LUT2 #(
		.INIT('h8)
	) name29460 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][16]/P0001 ,
		_w14702_,
		_w33507_
	);
	LUT2 #(
		.INIT('h8)
	) name29461 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001 ,
		_w14706_,
		_w33508_
	);
	LUT2 #(
		.INIT('h1)
	) name29462 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w33502_,
		_w33509_
	);
	LUT2 #(
		.INIT('h1)
	) name29463 (
		_w33503_,
		_w33504_,
		_w33510_
	);
	LUT2 #(
		.INIT('h1)
	) name29464 (
		_w33505_,
		_w33506_,
		_w33511_
	);
	LUT2 #(
		.INIT('h1)
	) name29465 (
		_w33507_,
		_w33508_,
		_w33512_
	);
	LUT2 #(
		.INIT('h8)
	) name29466 (
		_w33511_,
		_w33512_,
		_w33513_
	);
	LUT2 #(
		.INIT('h8)
	) name29467 (
		_w33509_,
		_w33510_,
		_w33514_
	);
	LUT2 #(
		.INIT('h8)
	) name29468 (
		_w33513_,
		_w33514_,
		_w33515_
	);
	LUT2 #(
		.INIT('h1)
	) name29469 (
		_w33501_,
		_w33515_,
		_w33516_
	);
	LUT2 #(
		.INIT('h8)
	) name29470 (
		_w32367_,
		_w33516_,
		_w33517_
	);
	LUT2 #(
		.INIT('h8)
	) name29471 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		_w33518_
	);
	LUT2 #(
		.INIT('h2)
	) name29472 (
		_w32364_,
		_w33518_,
		_w33519_
	);
	LUT2 #(
		.INIT('h2)
	) name29473 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w33519_,
		_w33520_
	);
	LUT2 #(
		.INIT('h4)
	) name29474 (
		_w32367_,
		_w33520_,
		_w33521_
	);
	LUT2 #(
		.INIT('h1)
	) name29475 (
		_w33517_,
		_w33521_,
		_w33522_
	);
	LUT2 #(
		.INIT('h4)
	) name29476 (
		_w4117_,
		_w31648_,
		_w33523_
	);
	LUT2 #(
		.INIT('h8)
	) name29477 (
		\core_c_dec_MFSR1_E_reg/P0001 ,
		_w4117_,
		_w33524_
	);
	LUT2 #(
		.INIT('h1)
	) name29478 (
		_w33523_,
		_w33524_,
		_w33525_
	);
	LUT2 #(
		.INIT('h4)
	) name29479 (
		_w4117_,
		_w31649_,
		_w33526_
	);
	LUT2 #(
		.INIT('h8)
	) name29480 (
		\core_c_dec_MFSR0_E_reg/P0001 ,
		_w4117_,
		_w33527_
	);
	LUT2 #(
		.INIT('h1)
	) name29481 (
		_w33526_,
		_w33527_,
		_w33528_
	);
	LUT2 #(
		.INIT('h4)
	) name29482 (
		_w4117_,
		_w31656_,
		_w33529_
	);
	LUT2 #(
		.INIT('h8)
	) name29483 (
		\core_c_dec_MFSI_E_reg/P0001 ,
		_w4117_,
		_w33530_
	);
	LUT2 #(
		.INIT('h1)
	) name29484 (
		_w33529_,
		_w33530_,
		_w33531_
	);
	LUT2 #(
		.INIT('h4)
	) name29485 (
		_w4117_,
		_w31652_,
		_w33532_
	);
	LUT2 #(
		.INIT('h8)
	) name29486 (
		\core_c_dec_MFSE_E_reg/P0001 ,
		_w4117_,
		_w33533_
	);
	LUT2 #(
		.INIT('h1)
	) name29487 (
		_w33532_,
		_w33533_,
		_w33534_
	);
	LUT2 #(
		.INIT('h8)
	) name29488 (
		\core_c_dec_MFMX1_E_reg/P0001 ,
		_w4117_,
		_w33535_
	);
	LUT2 #(
		.INIT('h8)
	) name29489 (
		_w30962_,
		_w32643_,
		_w33536_
	);
	LUT2 #(
		.INIT('h1)
	) name29490 (
		_w33535_,
		_w33536_,
		_w33537_
	);
	LUT2 #(
		.INIT('h4)
	) name29491 (
		_w4117_,
		_w30979_,
		_w33538_
	);
	LUT2 #(
		.INIT('h8)
	) name29492 (
		\core_c_dec_MFMR2_E_reg/P0001 ,
		_w4117_,
		_w33539_
	);
	LUT2 #(
		.INIT('h1)
	) name29493 (
		_w33538_,
		_w33539_,
		_w33540_
	);
	LUT2 #(
		.INIT('h4)
	) name29494 (
		_w4117_,
		_w30982_,
		_w33541_
	);
	LUT2 #(
		.INIT('h8)
	) name29495 (
		\core_c_dec_MFMR1_E_reg/P0001 ,
		_w4117_,
		_w33542_
	);
	LUT2 #(
		.INIT('h1)
	) name29496 (
		_w33541_,
		_w33542_,
		_w33543_
	);
	LUT2 #(
		.INIT('h4)
	) name29497 (
		_w4117_,
		_w30968_,
		_w33544_
	);
	LUT2 #(
		.INIT('h8)
	) name29498 (
		\core_c_dec_MFMR0_E_reg/P0001 ,
		_w4117_,
		_w33545_
	);
	LUT2 #(
		.INIT('h1)
	) name29499 (
		_w33544_,
		_w33545_,
		_w33546_
	);
	LUT2 #(
		.INIT('h8)
	) name29500 (
		\core_c_dec_MFAX1_E_reg/P0001 ,
		_w4117_,
		_w33547_
	);
	LUT2 #(
		.INIT('h8)
	) name29501 (
		_w31650_,
		_w32643_,
		_w33548_
	);
	LUT2 #(
		.INIT('h1)
	) name29502 (
		_w33547_,
		_w33548_,
		_w33549_
	);
	LUT2 #(
		.INIT('h4)
	) name29503 (
		_w4117_,
		_w31260_,
		_w33550_
	);
	LUT2 #(
		.INIT('h8)
	) name29504 (
		\core_c_dec_MFAR_E_reg/P0001 ,
		_w4117_,
		_w33551_
	);
	LUT2 #(
		.INIT('h1)
	) name29505 (
		_w33550_,
		_w33551_,
		_w33552_
	);
	LUT2 #(
		.INIT('h2)
	) name29506 (
		\sport1_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w32612_,
		_w33553_
	);
	LUT2 #(
		.INIT('h8)
	) name29507 (
		_w20407_,
		_w32616_,
		_w33554_
	);
	LUT2 #(
		.INIT('h2)
	) name29508 (
		\sport1_rxctl_Wcnt_reg[7]/NET0131 ,
		_w33554_,
		_w33555_
	);
	LUT2 #(
		.INIT('h8)
	) name29509 (
		_w32612_,
		_w33555_,
		_w33556_
	);
	LUT2 #(
		.INIT('h1)
	) name29510 (
		_w33553_,
		_w33556_,
		_w33557_
	);
	LUT2 #(
		.INIT('h4)
	) name29511 (
		\sport1_rxctl_Wcnt_reg[5]/NET0131 ,
		_w32618_,
		_w33558_
	);
	LUT2 #(
		.INIT('h2)
	) name29512 (
		\sport1_rxctl_Wcnt_reg[6]/NET0131 ,
		_w33558_,
		_w33559_
	);
	LUT2 #(
		.INIT('h1)
	) name29513 (
		_w33554_,
		_w33559_,
		_w33560_
	);
	LUT2 #(
		.INIT('h2)
	) name29514 (
		_w32612_,
		_w33560_,
		_w33561_
	);
	LUT2 #(
		.INIT('h2)
	) name29515 (
		\sport1_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w32612_,
		_w33562_
	);
	LUT2 #(
		.INIT('h1)
	) name29516 (
		_w33561_,
		_w33562_,
		_w33563_
	);
	LUT2 #(
		.INIT('h1)
	) name29517 (
		\sport1_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w32612_,
		_w33564_
	);
	LUT2 #(
		.INIT('h2)
	) name29518 (
		\sport1_rxctl_Wcnt_reg[5]/NET0131 ,
		_w32618_,
		_w33565_
	);
	LUT2 #(
		.INIT('h1)
	) name29519 (
		_w33558_,
		_w33565_,
		_w33566_
	);
	LUT2 #(
		.INIT('h8)
	) name29520 (
		_w32612_,
		_w33566_,
		_w33567_
	);
	LUT2 #(
		.INIT('h1)
	) name29521 (
		_w33564_,
		_w33567_,
		_w33568_
	);
	LUT2 #(
		.INIT('h2)
	) name29522 (
		\sport1_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w32612_,
		_w33569_
	);
	LUT2 #(
		.INIT('h2)
	) name29523 (
		\sport1_rxctl_Wcnt_reg[3]/NET0131 ,
		_w32615_,
		_w33570_
	);
	LUT2 #(
		.INIT('h1)
	) name29524 (
		_w32616_,
		_w33570_,
		_w33571_
	);
	LUT2 #(
		.INIT('h2)
	) name29525 (
		_w32612_,
		_w33571_,
		_w33572_
	);
	LUT2 #(
		.INIT('h1)
	) name29526 (
		_w33569_,
		_w33572_,
		_w33573_
	);
	LUT2 #(
		.INIT('h1)
	) name29527 (
		\sport1_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w32612_,
		_w33574_
	);
	LUT2 #(
		.INIT('h2)
	) name29528 (
		\sport1_rxctl_Wcnt_reg[2]/NET0131 ,
		_w32614_,
		_w33575_
	);
	LUT2 #(
		.INIT('h1)
	) name29529 (
		_w32615_,
		_w33575_,
		_w33576_
	);
	LUT2 #(
		.INIT('h8)
	) name29530 (
		_w32612_,
		_w33576_,
		_w33577_
	);
	LUT2 #(
		.INIT('h1)
	) name29531 (
		_w33574_,
		_w33577_,
		_w33578_
	);
	LUT2 #(
		.INIT('h4)
	) name29532 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		_w32613_,
		_w33579_
	);
	LUT2 #(
		.INIT('h2)
	) name29533 (
		\sport1_rxctl_Wcnt_reg[1]/NET0131 ,
		_w33579_,
		_w33580_
	);
	LUT2 #(
		.INIT('h1)
	) name29534 (
		_w32614_,
		_w33580_,
		_w33581_
	);
	LUT2 #(
		.INIT('h2)
	) name29535 (
		_w32612_,
		_w33581_,
		_w33582_
	);
	LUT2 #(
		.INIT('h2)
	) name29536 (
		\sport1_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w32612_,
		_w33583_
	);
	LUT2 #(
		.INIT('h1)
	) name29537 (
		_w33582_,
		_w33583_,
		_w33584_
	);
	LUT2 #(
		.INIT('h2)
	) name29538 (
		\sport1_rxctl_Wcnt_reg[0]/NET0131 ,
		_w32613_,
		_w33585_
	);
	LUT2 #(
		.INIT('h1)
	) name29539 (
		_w33579_,
		_w33585_,
		_w33586_
	);
	LUT2 #(
		.INIT('h2)
	) name29540 (
		_w32612_,
		_w33586_,
		_w33587_
	);
	LUT2 #(
		.INIT('h2)
	) name29541 (
		\sport1_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w32612_,
		_w33588_
	);
	LUT2 #(
		.INIT('h1)
	) name29542 (
		_w33587_,
		_w33588_,
		_w33589_
	);
	LUT2 #(
		.INIT('h2)
	) name29543 (
		\sport0_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w32658_,
		_w33590_
	);
	LUT2 #(
		.INIT('h8)
	) name29544 (
		_w20429_,
		_w32662_,
		_w33591_
	);
	LUT2 #(
		.INIT('h2)
	) name29545 (
		\sport0_rxctl_Wcnt_reg[7]/NET0131 ,
		_w33591_,
		_w33592_
	);
	LUT2 #(
		.INIT('h8)
	) name29546 (
		_w32658_,
		_w33592_,
		_w33593_
	);
	LUT2 #(
		.INIT('h1)
	) name29547 (
		_w33590_,
		_w33593_,
		_w33594_
	);
	LUT2 #(
		.INIT('h1)
	) name29548 (
		\sport0_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w32658_,
		_w33595_
	);
	LUT2 #(
		.INIT('h2)
	) name29549 (
		\sport0_rxctl_Wcnt_reg[5]/NET0131 ,
		_w32664_,
		_w33596_
	);
	LUT2 #(
		.INIT('h4)
	) name29550 (
		\sport0_rxctl_Wcnt_reg[5]/NET0131 ,
		_w32664_,
		_w33597_
	);
	LUT2 #(
		.INIT('h1)
	) name29551 (
		_w33596_,
		_w33597_,
		_w33598_
	);
	LUT2 #(
		.INIT('h8)
	) name29552 (
		_w32658_,
		_w33598_,
		_w33599_
	);
	LUT2 #(
		.INIT('h1)
	) name29553 (
		_w33595_,
		_w33599_,
		_w33600_
	);
	LUT2 #(
		.INIT('h2)
	) name29554 (
		\sport0_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w32658_,
		_w33601_
	);
	LUT2 #(
		.INIT('h2)
	) name29555 (
		\sport0_rxctl_Wcnt_reg[3]/NET0131 ,
		_w32661_,
		_w33602_
	);
	LUT2 #(
		.INIT('h1)
	) name29556 (
		_w32662_,
		_w33602_,
		_w33603_
	);
	LUT2 #(
		.INIT('h2)
	) name29557 (
		_w32658_,
		_w33603_,
		_w33604_
	);
	LUT2 #(
		.INIT('h1)
	) name29558 (
		_w33601_,
		_w33604_,
		_w33605_
	);
	LUT2 #(
		.INIT('h4)
	) name29559 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		_w32659_,
		_w33606_
	);
	LUT2 #(
		.INIT('h2)
	) name29560 (
		\sport0_rxctl_Wcnt_reg[1]/NET0131 ,
		_w33606_,
		_w33607_
	);
	LUT2 #(
		.INIT('h1)
	) name29561 (
		_w32660_,
		_w33607_,
		_w33608_
	);
	LUT2 #(
		.INIT('h2)
	) name29562 (
		_w32658_,
		_w33608_,
		_w33609_
	);
	LUT2 #(
		.INIT('h2)
	) name29563 (
		\sport0_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w32658_,
		_w33610_
	);
	LUT2 #(
		.INIT('h1)
	) name29564 (
		_w33609_,
		_w33610_,
		_w33611_
	);
	LUT2 #(
		.INIT('h2)
	) name29565 (
		\sport0_rxctl_Wcnt_reg[0]/NET0131 ,
		_w32659_,
		_w33612_
	);
	LUT2 #(
		.INIT('h1)
	) name29566 (
		_w33606_,
		_w33612_,
		_w33613_
	);
	LUT2 #(
		.INIT('h2)
	) name29567 (
		_w32658_,
		_w33613_,
		_w33614_
	);
	LUT2 #(
		.INIT('h2)
	) name29568 (
		\sport0_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w32658_,
		_w33615_
	);
	LUT2 #(
		.INIT('h1)
	) name29569 (
		_w33614_,
		_w33615_,
		_w33616_
	);
	LUT2 #(
		.INIT('h8)
	) name29570 (
		\clkc_oscntr_reg_DO_reg[10]/NET0131 ,
		_w23424_,
		_w33617_
	);
	LUT2 #(
		.INIT('h2)
	) name29571 (
		\clkc_oscntr_reg_DO_reg[11]/NET0131 ,
		_w33617_,
		_w33618_
	);
	LUT2 #(
		.INIT('h4)
	) name29572 (
		\clkc_oscntr_reg_DO_reg[11]/NET0131 ,
		_w33617_,
		_w33619_
	);
	LUT2 #(
		.INIT('h1)
	) name29573 (
		_w33618_,
		_w33619_,
		_w33620_
	);
	LUT2 #(
		.INIT('h1)
	) name29574 (
		\sport0_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w32658_,
		_w33621_
	);
	LUT2 #(
		.INIT('h2)
	) name29575 (
		\sport0_rxctl_Wcnt_reg[2]/NET0131 ,
		_w32660_,
		_w33622_
	);
	LUT2 #(
		.INIT('h1)
	) name29576 (
		_w32661_,
		_w33622_,
		_w33623_
	);
	LUT2 #(
		.INIT('h8)
	) name29577 (
		_w32658_,
		_w33623_,
		_w33624_
	);
	LUT2 #(
		.INIT('h1)
	) name29578 (
		_w33621_,
		_w33624_,
		_w33625_
	);
	LUT2 #(
		.INIT('h2)
	) name29579 (
		\sport0_rxctl_Wcnt_reg[6]/NET0131 ,
		_w33597_,
		_w33626_
	);
	LUT2 #(
		.INIT('h1)
	) name29580 (
		_w33591_,
		_w33626_,
		_w33627_
	);
	LUT2 #(
		.INIT('h2)
	) name29581 (
		_w32658_,
		_w33627_,
		_w33628_
	);
	LUT2 #(
		.INIT('h2)
	) name29582 (
		\sport0_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w32658_,
		_w33629_
	);
	LUT2 #(
		.INIT('h1)
	) name29583 (
		_w33628_,
		_w33629_,
		_w33630_
	);
	LUT2 #(
		.INIT('h1)
	) name29584 (
		\sice_IIRC_reg[16]/NET0131 ,
		_w22581_,
		_w33631_
	);
	LUT2 #(
		.INIT('h1)
	) name29585 (
		_w22582_,
		_w33631_,
		_w33632_
	);
	LUT2 #(
		.INIT('h8)
	) name29586 (
		\core_c_dec_MFAX0_E_reg/P0001 ,
		_w4117_,
		_w33633_
	);
	LUT2 #(
		.INIT('h8)
	) name29587 (
		_w31650_,
		_w32639_,
		_w33634_
	);
	LUT2 #(
		.INIT('h1)
	) name29588 (
		_w33633_,
		_w33634_,
		_w33635_
	);
	LUT2 #(
		.INIT('h2)
	) name29589 (
		_w10289_,
		_w32992_,
		_w33636_
	);
	LUT2 #(
		.INIT('h8)
	) name29590 (
		\core_dag_ilm2reg_L6_we_DO_reg[9]/NET0131 ,
		_w32994_,
		_w33637_
	);
	LUT2 #(
		.INIT('h8)
	) name29591 (
		\core_dag_ilm2reg_L4_we_DO_reg[9]/NET0131 ,
		_w32996_,
		_w33638_
	);
	LUT2 #(
		.INIT('h8)
	) name29592 (
		\core_dag_ilm2reg_L7_we_DO_reg[9]/NET0131 ,
		_w32998_,
		_w33639_
	);
	LUT2 #(
		.INIT('h8)
	) name29593 (
		\core_dag_ilm2reg_L5_we_DO_reg[9]/NET0131 ,
		_w33000_,
		_w33640_
	);
	LUT2 #(
		.INIT('h1)
	) name29594 (
		_w21579_,
		_w33637_,
		_w33641_
	);
	LUT2 #(
		.INIT('h1)
	) name29595 (
		_w33638_,
		_w33639_,
		_w33642_
	);
	LUT2 #(
		.INIT('h4)
	) name29596 (
		_w33640_,
		_w33642_,
		_w33643_
	);
	LUT2 #(
		.INIT('h8)
	) name29597 (
		_w33641_,
		_w33643_,
		_w33644_
	);
	LUT2 #(
		.INIT('h4)
	) name29598 (
		_w33636_,
		_w33644_,
		_w33645_
	);
	LUT2 #(
		.INIT('h4)
	) name29599 (
		\core_dag_ilm2reg_L_reg[9]/NET0131 ,
		_w21579_,
		_w33646_
	);
	LUT2 #(
		.INIT('h1)
	) name29600 (
		_w33645_,
		_w33646_,
		_w33647_
	);
	LUT2 #(
		.INIT('h2)
	) name29601 (
		_w10638_,
		_w32992_,
		_w33648_
	);
	LUT2 #(
		.INIT('h8)
	) name29602 (
		\core_dag_ilm2reg_L6_we_DO_reg[8]/NET0131 ,
		_w32994_,
		_w33649_
	);
	LUT2 #(
		.INIT('h8)
	) name29603 (
		\core_dag_ilm2reg_L4_we_DO_reg[8]/NET0131 ,
		_w32996_,
		_w33650_
	);
	LUT2 #(
		.INIT('h8)
	) name29604 (
		\core_dag_ilm2reg_L7_we_DO_reg[8]/NET0131 ,
		_w32998_,
		_w33651_
	);
	LUT2 #(
		.INIT('h8)
	) name29605 (
		\core_dag_ilm2reg_L5_we_DO_reg[8]/NET0131 ,
		_w33000_,
		_w33652_
	);
	LUT2 #(
		.INIT('h1)
	) name29606 (
		_w21579_,
		_w33649_,
		_w33653_
	);
	LUT2 #(
		.INIT('h1)
	) name29607 (
		_w33650_,
		_w33651_,
		_w33654_
	);
	LUT2 #(
		.INIT('h4)
	) name29608 (
		_w33652_,
		_w33654_,
		_w33655_
	);
	LUT2 #(
		.INIT('h8)
	) name29609 (
		_w33653_,
		_w33655_,
		_w33656_
	);
	LUT2 #(
		.INIT('h4)
	) name29610 (
		_w33648_,
		_w33656_,
		_w33657_
	);
	LUT2 #(
		.INIT('h4)
	) name29611 (
		\core_dag_ilm2reg_L_reg[8]/NET0131 ,
		_w21579_,
		_w33658_
	);
	LUT2 #(
		.INIT('h1)
	) name29612 (
		_w33657_,
		_w33658_,
		_w33659_
	);
	LUT2 #(
		.INIT('h2)
	) name29613 (
		_w9178_,
		_w32992_,
		_w33660_
	);
	LUT2 #(
		.INIT('h8)
	) name29614 (
		\core_dag_ilm2reg_L6_we_DO_reg[12]/NET0131 ,
		_w32994_,
		_w33661_
	);
	LUT2 #(
		.INIT('h8)
	) name29615 (
		\core_dag_ilm2reg_L4_we_DO_reg[12]/NET0131 ,
		_w32996_,
		_w33662_
	);
	LUT2 #(
		.INIT('h8)
	) name29616 (
		\core_dag_ilm2reg_L7_we_DO_reg[12]/NET0131 ,
		_w32998_,
		_w33663_
	);
	LUT2 #(
		.INIT('h8)
	) name29617 (
		\core_dag_ilm2reg_L5_we_DO_reg[12]/NET0131 ,
		_w33000_,
		_w33664_
	);
	LUT2 #(
		.INIT('h1)
	) name29618 (
		_w21579_,
		_w33661_,
		_w33665_
	);
	LUT2 #(
		.INIT('h1)
	) name29619 (
		_w33662_,
		_w33663_,
		_w33666_
	);
	LUT2 #(
		.INIT('h4)
	) name29620 (
		_w33664_,
		_w33666_,
		_w33667_
	);
	LUT2 #(
		.INIT('h8)
	) name29621 (
		_w33665_,
		_w33667_,
		_w33668_
	);
	LUT2 #(
		.INIT('h4)
	) name29622 (
		_w33660_,
		_w33668_,
		_w33669_
	);
	LUT2 #(
		.INIT('h4)
	) name29623 (
		\core_dag_ilm2reg_L_reg[12]/NET0131 ,
		_w21579_,
		_w33670_
	);
	LUT2 #(
		.INIT('h1)
	) name29624 (
		_w33669_,
		_w33670_,
		_w33671_
	);
	LUT2 #(
		.INIT('h2)
	) name29625 (
		_w8460_,
		_w32992_,
		_w33672_
	);
	LUT2 #(
		.INIT('h8)
	) name29626 (
		\core_dag_ilm2reg_L6_we_DO_reg[11]/NET0131 ,
		_w32994_,
		_w33673_
	);
	LUT2 #(
		.INIT('h8)
	) name29627 (
		\core_dag_ilm2reg_L4_we_DO_reg[11]/NET0131 ,
		_w32996_,
		_w33674_
	);
	LUT2 #(
		.INIT('h8)
	) name29628 (
		\core_dag_ilm2reg_L7_we_DO_reg[11]/NET0131 ,
		_w32998_,
		_w33675_
	);
	LUT2 #(
		.INIT('h8)
	) name29629 (
		\core_dag_ilm2reg_L5_we_DO_reg[11]/NET0131 ,
		_w33000_,
		_w33676_
	);
	LUT2 #(
		.INIT('h1)
	) name29630 (
		_w21579_,
		_w33673_,
		_w33677_
	);
	LUT2 #(
		.INIT('h1)
	) name29631 (
		_w33674_,
		_w33675_,
		_w33678_
	);
	LUT2 #(
		.INIT('h4)
	) name29632 (
		_w33676_,
		_w33678_,
		_w33679_
	);
	LUT2 #(
		.INIT('h8)
	) name29633 (
		_w33677_,
		_w33679_,
		_w33680_
	);
	LUT2 #(
		.INIT('h4)
	) name29634 (
		_w33672_,
		_w33680_,
		_w33681_
	);
	LUT2 #(
		.INIT('h4)
	) name29635 (
		\core_dag_ilm2reg_L_reg[11]/NET0131 ,
		_w21579_,
		_w33682_
	);
	LUT2 #(
		.INIT('h1)
	) name29636 (
		_w33681_,
		_w33682_,
		_w33683_
	);
	LUT2 #(
		.INIT('h8)
	) name29637 (
		_w6008_,
		_w32984_,
		_w33684_
	);
	LUT2 #(
		.INIT('h8)
	) name29638 (
		\core_dag_ilm2reg_I6_we_DO_reg[9]/NET0131 ,
		_w33684_,
		_w33685_
	);
	LUT2 #(
		.INIT('h8)
	) name29639 (
		_w6000_,
		_w32988_,
		_w33686_
	);
	LUT2 #(
		.INIT('h8)
	) name29640 (
		\core_dag_ilm2reg_I7_we_DO_reg[9]/NET0131 ,
		_w33686_,
		_w33687_
	);
	LUT2 #(
		.INIT('h8)
	) name29641 (
		_w6015_,
		_w32982_,
		_w33688_
	);
	LUT2 #(
		.INIT('h8)
	) name29642 (
		\core_dag_ilm2reg_I5_we_DO_reg[9]/NET0131 ,
		_w33688_,
		_w33689_
	);
	LUT2 #(
		.INIT('h8)
	) name29643 (
		_w5964_,
		_w32986_,
		_w33690_
	);
	LUT2 #(
		.INIT('h8)
	) name29644 (
		\core_dag_ilm2reg_I4_we_DO_reg[9]/NET0131 ,
		_w33690_,
		_w33691_
	);
	LUT2 #(
		.INIT('h4)
	) name29645 (
		_w6008_,
		_w32984_,
		_w33692_
	);
	LUT2 #(
		.INIT('h4)
	) name29646 (
		_w5964_,
		_w32986_,
		_w33693_
	);
	LUT2 #(
		.INIT('h4)
	) name29647 (
		_w6000_,
		_w32988_,
		_w33694_
	);
	LUT2 #(
		.INIT('h4)
	) name29648 (
		_w6015_,
		_w32982_,
		_w33695_
	);
	LUT2 #(
		.INIT('h1)
	) name29649 (
		_w33692_,
		_w33693_,
		_w33696_
	);
	LUT2 #(
		.INIT('h1)
	) name29650 (
		_w33694_,
		_w33695_,
		_w33697_
	);
	LUT2 #(
		.INIT('h8)
	) name29651 (
		_w33696_,
		_w33697_,
		_w33698_
	);
	LUT2 #(
		.INIT('h2)
	) name29652 (
		_w20755_,
		_w33698_,
		_w33699_
	);
	LUT2 #(
		.INIT('h1)
	) name29653 (
		_w21579_,
		_w33685_,
		_w33700_
	);
	LUT2 #(
		.INIT('h1)
	) name29654 (
		_w33687_,
		_w33689_,
		_w33701_
	);
	LUT2 #(
		.INIT('h4)
	) name29655 (
		_w33691_,
		_w33701_,
		_w33702_
	);
	LUT2 #(
		.INIT('h8)
	) name29656 (
		_w33700_,
		_w33702_,
		_w33703_
	);
	LUT2 #(
		.INIT('h4)
	) name29657 (
		_w33699_,
		_w33703_,
		_w33704_
	);
	LUT2 #(
		.INIT('h4)
	) name29658 (
		\core_dag_ilm2reg_I_reg[9]/NET0131 ,
		_w21579_,
		_w33705_
	);
	LUT2 #(
		.INIT('h1)
	) name29659 (
		_w33704_,
		_w33705_,
		_w33706_
	);
	LUT2 #(
		.INIT('h8)
	) name29660 (
		\core_dag_ilm2reg_I6_we_DO_reg[6]/NET0131 ,
		_w33684_,
		_w33707_
	);
	LUT2 #(
		.INIT('h8)
	) name29661 (
		\core_dag_ilm2reg_I7_we_DO_reg[6]/NET0131 ,
		_w33686_,
		_w33708_
	);
	LUT2 #(
		.INIT('h8)
	) name29662 (
		\core_dag_ilm2reg_I5_we_DO_reg[6]/NET0131 ,
		_w33688_,
		_w33709_
	);
	LUT2 #(
		.INIT('h8)
	) name29663 (
		\core_dag_ilm2reg_I4_we_DO_reg[6]/NET0131 ,
		_w33690_,
		_w33710_
	);
	LUT2 #(
		.INIT('h2)
	) name29664 (
		_w20624_,
		_w33698_,
		_w33711_
	);
	LUT2 #(
		.INIT('h1)
	) name29665 (
		_w21579_,
		_w33707_,
		_w33712_
	);
	LUT2 #(
		.INIT('h1)
	) name29666 (
		_w33708_,
		_w33709_,
		_w33713_
	);
	LUT2 #(
		.INIT('h4)
	) name29667 (
		_w33710_,
		_w33713_,
		_w33714_
	);
	LUT2 #(
		.INIT('h8)
	) name29668 (
		_w33712_,
		_w33714_,
		_w33715_
	);
	LUT2 #(
		.INIT('h4)
	) name29669 (
		_w33711_,
		_w33715_,
		_w33716_
	);
	LUT2 #(
		.INIT('h4)
	) name29670 (
		\core_dag_ilm2reg_I_reg[6]/NET0131 ,
		_w21579_,
		_w33717_
	);
	LUT2 #(
		.INIT('h1)
	) name29671 (
		_w33716_,
		_w33717_,
		_w33718_
	);
	LUT2 #(
		.INIT('h8)
	) name29672 (
		\core_dag_ilm2reg_I6_we_DO_reg[5]/NET0131 ,
		_w33684_,
		_w33719_
	);
	LUT2 #(
		.INIT('h8)
	) name29673 (
		\core_dag_ilm2reg_I7_we_DO_reg[5]/NET0131 ,
		_w33686_,
		_w33720_
	);
	LUT2 #(
		.INIT('h8)
	) name29674 (
		\core_dag_ilm2reg_I5_we_DO_reg[5]/NET0131 ,
		_w33688_,
		_w33721_
	);
	LUT2 #(
		.INIT('h8)
	) name29675 (
		\core_dag_ilm2reg_I4_we_DO_reg[5]/NET0131 ,
		_w33690_,
		_w33722_
	);
	LUT2 #(
		.INIT('h2)
	) name29676 (
		_w20634_,
		_w33698_,
		_w33723_
	);
	LUT2 #(
		.INIT('h1)
	) name29677 (
		_w21579_,
		_w33719_,
		_w33724_
	);
	LUT2 #(
		.INIT('h1)
	) name29678 (
		_w33720_,
		_w33721_,
		_w33725_
	);
	LUT2 #(
		.INIT('h4)
	) name29679 (
		_w33722_,
		_w33725_,
		_w33726_
	);
	LUT2 #(
		.INIT('h8)
	) name29680 (
		_w33724_,
		_w33726_,
		_w33727_
	);
	LUT2 #(
		.INIT('h4)
	) name29681 (
		_w33723_,
		_w33727_,
		_w33728_
	);
	LUT2 #(
		.INIT('h4)
	) name29682 (
		\core_dag_ilm2reg_I_reg[5]/NET0131 ,
		_w21579_,
		_w33729_
	);
	LUT2 #(
		.INIT('h1)
	) name29683 (
		_w33728_,
		_w33729_,
		_w33730_
	);
	LUT2 #(
		.INIT('h8)
	) name29684 (
		\core_dag_ilm2reg_I6_we_DO_reg[4]/NET0131 ,
		_w33684_,
		_w33731_
	);
	LUT2 #(
		.INIT('h8)
	) name29685 (
		\core_dag_ilm2reg_I7_we_DO_reg[4]/NET0131 ,
		_w33686_,
		_w33732_
	);
	LUT2 #(
		.INIT('h8)
	) name29686 (
		\core_dag_ilm2reg_I5_we_DO_reg[4]/NET0131 ,
		_w33688_,
		_w33733_
	);
	LUT2 #(
		.INIT('h8)
	) name29687 (
		\core_dag_ilm2reg_I4_we_DO_reg[4]/NET0131 ,
		_w33690_,
		_w33734_
	);
	LUT2 #(
		.INIT('h2)
	) name29688 (
		_w20644_,
		_w33698_,
		_w33735_
	);
	LUT2 #(
		.INIT('h1)
	) name29689 (
		_w21579_,
		_w33731_,
		_w33736_
	);
	LUT2 #(
		.INIT('h1)
	) name29690 (
		_w33732_,
		_w33733_,
		_w33737_
	);
	LUT2 #(
		.INIT('h4)
	) name29691 (
		_w33734_,
		_w33737_,
		_w33738_
	);
	LUT2 #(
		.INIT('h8)
	) name29692 (
		_w33736_,
		_w33738_,
		_w33739_
	);
	LUT2 #(
		.INIT('h4)
	) name29693 (
		_w33735_,
		_w33739_,
		_w33740_
	);
	LUT2 #(
		.INIT('h4)
	) name29694 (
		\core_dag_ilm2reg_I_reg[4]/NET0131 ,
		_w21579_,
		_w33741_
	);
	LUT2 #(
		.INIT('h1)
	) name29695 (
		_w33740_,
		_w33741_,
		_w33742_
	);
	LUT2 #(
		.INIT('h8)
	) name29696 (
		\core_dag_ilm2reg_I6_we_DO_reg[3]/NET0131 ,
		_w33684_,
		_w33743_
	);
	LUT2 #(
		.INIT('h8)
	) name29697 (
		\core_dag_ilm2reg_I5_we_DO_reg[3]/NET0131 ,
		_w33688_,
		_w33744_
	);
	LUT2 #(
		.INIT('h8)
	) name29698 (
		\core_dag_ilm2reg_I7_we_DO_reg[3]/NET0131 ,
		_w33686_,
		_w33745_
	);
	LUT2 #(
		.INIT('h8)
	) name29699 (
		\core_dag_ilm2reg_I4_we_DO_reg[3]/NET0131 ,
		_w33690_,
		_w33746_
	);
	LUT2 #(
		.INIT('h2)
	) name29700 (
		_w13262_,
		_w33698_,
		_w33747_
	);
	LUT2 #(
		.INIT('h1)
	) name29701 (
		_w21579_,
		_w33743_,
		_w33748_
	);
	LUT2 #(
		.INIT('h1)
	) name29702 (
		_w33744_,
		_w33745_,
		_w33749_
	);
	LUT2 #(
		.INIT('h4)
	) name29703 (
		_w33746_,
		_w33749_,
		_w33750_
	);
	LUT2 #(
		.INIT('h8)
	) name29704 (
		_w33748_,
		_w33750_,
		_w33751_
	);
	LUT2 #(
		.INIT('h4)
	) name29705 (
		_w33747_,
		_w33751_,
		_w33752_
	);
	LUT2 #(
		.INIT('h4)
	) name29706 (
		\core_dag_ilm2reg_I_reg[3]/NET0131 ,
		_w21579_,
		_w33753_
	);
	LUT2 #(
		.INIT('h1)
	) name29707 (
		_w33752_,
		_w33753_,
		_w33754_
	);
	LUT2 #(
		.INIT('h8)
	) name29708 (
		\core_dag_ilm2reg_I6_we_DO_reg[2]/NET0131 ,
		_w33684_,
		_w33755_
	);
	LUT2 #(
		.INIT('h8)
	) name29709 (
		\core_dag_ilm2reg_I7_we_DO_reg[2]/NET0131 ,
		_w33686_,
		_w33756_
	);
	LUT2 #(
		.INIT('h8)
	) name29710 (
		\core_dag_ilm2reg_I5_we_DO_reg[2]/NET0131 ,
		_w33688_,
		_w33757_
	);
	LUT2 #(
		.INIT('h8)
	) name29711 (
		\core_dag_ilm2reg_I4_we_DO_reg[2]/NET0131 ,
		_w33690_,
		_w33758_
	);
	LUT2 #(
		.INIT('h1)
	) name29712 (
		_w20663_,
		_w33698_,
		_w33759_
	);
	LUT2 #(
		.INIT('h1)
	) name29713 (
		_w21579_,
		_w33755_,
		_w33760_
	);
	LUT2 #(
		.INIT('h1)
	) name29714 (
		_w33756_,
		_w33757_,
		_w33761_
	);
	LUT2 #(
		.INIT('h4)
	) name29715 (
		_w33758_,
		_w33761_,
		_w33762_
	);
	LUT2 #(
		.INIT('h8)
	) name29716 (
		_w33760_,
		_w33762_,
		_w33763_
	);
	LUT2 #(
		.INIT('h4)
	) name29717 (
		_w33759_,
		_w33763_,
		_w33764_
	);
	LUT2 #(
		.INIT('h4)
	) name29718 (
		\core_dag_ilm2reg_I_reg[2]/NET0131 ,
		_w21579_,
		_w33765_
	);
	LUT2 #(
		.INIT('h1)
	) name29719 (
		_w33764_,
		_w33765_,
		_w33766_
	);
	LUT2 #(
		.INIT('h8)
	) name29720 (
		\core_dag_ilm2reg_I6_we_DO_reg[1]/NET0131 ,
		_w33684_,
		_w33767_
	);
	LUT2 #(
		.INIT('h8)
	) name29721 (
		\core_dag_ilm2reg_I5_we_DO_reg[1]/NET0131 ,
		_w33688_,
		_w33768_
	);
	LUT2 #(
		.INIT('h8)
	) name29722 (
		\core_dag_ilm2reg_I7_we_DO_reg[1]/NET0131 ,
		_w33686_,
		_w33769_
	);
	LUT2 #(
		.INIT('h8)
	) name29723 (
		\core_dag_ilm2reg_I4_we_DO_reg[1]/NET0131 ,
		_w33690_,
		_w33770_
	);
	LUT2 #(
		.INIT('h1)
	) name29724 (
		_w20674_,
		_w33698_,
		_w33771_
	);
	LUT2 #(
		.INIT('h1)
	) name29725 (
		_w21579_,
		_w33767_,
		_w33772_
	);
	LUT2 #(
		.INIT('h1)
	) name29726 (
		_w33768_,
		_w33769_,
		_w33773_
	);
	LUT2 #(
		.INIT('h4)
	) name29727 (
		_w33770_,
		_w33773_,
		_w33774_
	);
	LUT2 #(
		.INIT('h8)
	) name29728 (
		_w33772_,
		_w33774_,
		_w33775_
	);
	LUT2 #(
		.INIT('h4)
	) name29729 (
		_w33771_,
		_w33775_,
		_w33776_
	);
	LUT2 #(
		.INIT('h4)
	) name29730 (
		\core_dag_ilm2reg_I_reg[1]/NET0131 ,
		_w21579_,
		_w33777_
	);
	LUT2 #(
		.INIT('h1)
	) name29731 (
		_w33776_,
		_w33777_,
		_w33778_
	);
	LUT2 #(
		.INIT('h8)
	) name29732 (
		\core_dag_ilm2reg_I6_we_DO_reg[13]/NET0131 ,
		_w33684_,
		_w33779_
	);
	LUT2 #(
		.INIT('h8)
	) name29733 (
		\core_dag_ilm2reg_I5_we_DO_reg[13]/NET0131 ,
		_w33688_,
		_w33780_
	);
	LUT2 #(
		.INIT('h8)
	) name29734 (
		\core_dag_ilm2reg_I7_we_DO_reg[13]/NET0131 ,
		_w33686_,
		_w33781_
	);
	LUT2 #(
		.INIT('h8)
	) name29735 (
		\core_dag_ilm2reg_I4_we_DO_reg[13]/NET0131 ,
		_w33690_,
		_w33782_
	);
	LUT2 #(
		.INIT('h1)
	) name29736 (
		_w20685_,
		_w33698_,
		_w33783_
	);
	LUT2 #(
		.INIT('h1)
	) name29737 (
		_w21579_,
		_w33779_,
		_w33784_
	);
	LUT2 #(
		.INIT('h1)
	) name29738 (
		_w33780_,
		_w33781_,
		_w33785_
	);
	LUT2 #(
		.INIT('h4)
	) name29739 (
		_w33782_,
		_w33785_,
		_w33786_
	);
	LUT2 #(
		.INIT('h8)
	) name29740 (
		_w33784_,
		_w33786_,
		_w33787_
	);
	LUT2 #(
		.INIT('h4)
	) name29741 (
		_w33783_,
		_w33787_,
		_w33788_
	);
	LUT2 #(
		.INIT('h4)
	) name29742 (
		\core_dag_ilm2reg_I_reg[13]/NET0131 ,
		_w21579_,
		_w33789_
	);
	LUT2 #(
		.INIT('h1)
	) name29743 (
		_w33788_,
		_w33789_,
		_w33790_
	);
	LUT2 #(
		.INIT('h8)
	) name29744 (
		\core_dag_ilm2reg_I6_we_DO_reg[12]/NET0131 ,
		_w33684_,
		_w33791_
	);
	LUT2 #(
		.INIT('h8)
	) name29745 (
		\core_dag_ilm2reg_I7_we_DO_reg[12]/NET0131 ,
		_w33686_,
		_w33792_
	);
	LUT2 #(
		.INIT('h8)
	) name29746 (
		\core_dag_ilm2reg_I5_we_DO_reg[12]/NET0131 ,
		_w33688_,
		_w33793_
	);
	LUT2 #(
		.INIT('h8)
	) name29747 (
		\core_dag_ilm2reg_I4_we_DO_reg[12]/NET0131 ,
		_w33690_,
		_w33794_
	);
	LUT2 #(
		.INIT('h1)
	) name29748 (
		_w20696_,
		_w33698_,
		_w33795_
	);
	LUT2 #(
		.INIT('h1)
	) name29749 (
		_w21579_,
		_w33791_,
		_w33796_
	);
	LUT2 #(
		.INIT('h1)
	) name29750 (
		_w33792_,
		_w33793_,
		_w33797_
	);
	LUT2 #(
		.INIT('h4)
	) name29751 (
		_w33794_,
		_w33797_,
		_w33798_
	);
	LUT2 #(
		.INIT('h8)
	) name29752 (
		_w33796_,
		_w33798_,
		_w33799_
	);
	LUT2 #(
		.INIT('h4)
	) name29753 (
		_w33795_,
		_w33799_,
		_w33800_
	);
	LUT2 #(
		.INIT('h4)
	) name29754 (
		\core_dag_ilm2reg_I_reg[12]/NET0131 ,
		_w21579_,
		_w33801_
	);
	LUT2 #(
		.INIT('h1)
	) name29755 (
		_w33800_,
		_w33801_,
		_w33802_
	);
	LUT2 #(
		.INIT('h8)
	) name29756 (
		\core_dag_ilm2reg_I6_we_DO_reg[0]/NET0131 ,
		_w33684_,
		_w33803_
	);
	LUT2 #(
		.INIT('h8)
	) name29757 (
		\core_dag_ilm2reg_I7_we_DO_reg[0]/NET0131 ,
		_w33686_,
		_w33804_
	);
	LUT2 #(
		.INIT('h8)
	) name29758 (
		\core_dag_ilm2reg_I5_we_DO_reg[0]/NET0131 ,
		_w33688_,
		_w33805_
	);
	LUT2 #(
		.INIT('h8)
	) name29759 (
		\core_dag_ilm2reg_I4_we_DO_reg[0]/NET0131 ,
		_w33690_,
		_w33806_
	);
	LUT2 #(
		.INIT('h1)
	) name29760 (
		_w20729_,
		_w33698_,
		_w33807_
	);
	LUT2 #(
		.INIT('h1)
	) name29761 (
		_w21579_,
		_w33803_,
		_w33808_
	);
	LUT2 #(
		.INIT('h1)
	) name29762 (
		_w33804_,
		_w33805_,
		_w33809_
	);
	LUT2 #(
		.INIT('h4)
	) name29763 (
		_w33806_,
		_w33809_,
		_w33810_
	);
	LUT2 #(
		.INIT('h8)
	) name29764 (
		_w33808_,
		_w33810_,
		_w33811_
	);
	LUT2 #(
		.INIT('h4)
	) name29765 (
		_w33807_,
		_w33811_,
		_w33812_
	);
	LUT2 #(
		.INIT('h4)
	) name29766 (
		\core_dag_ilm2reg_I_reg[0]/NET0131 ,
		_w21579_,
		_w33813_
	);
	LUT2 #(
		.INIT('h1)
	) name29767 (
		_w33812_,
		_w33813_,
		_w33814_
	);
	LUT2 #(
		.INIT('h2)
	) name29768 (
		_w10289_,
		_w33099_,
		_w33815_
	);
	LUT2 #(
		.INIT('h8)
	) name29769 (
		\core_dag_ilm1reg_L1_we_DO_reg[9]/NET0131 ,
		_w33105_,
		_w33816_
	);
	LUT2 #(
		.INIT('h8)
	) name29770 (
		\core_dag_ilm1reg_L2_we_DO_reg[9]/NET0131 ,
		_w33107_,
		_w33817_
	);
	LUT2 #(
		.INIT('h8)
	) name29771 (
		\core_dag_ilm1reg_L3_we_DO_reg[9]/NET0131 ,
		_w33101_,
		_w33818_
	);
	LUT2 #(
		.INIT('h8)
	) name29772 (
		\core_dag_ilm1reg_L0_we_DO_reg[9]/NET0131 ,
		_w33103_,
		_w33819_
	);
	LUT2 #(
		.INIT('h1)
	) name29773 (
		_w33816_,
		_w33817_,
		_w33820_
	);
	LUT2 #(
		.INIT('h1)
	) name29774 (
		_w33818_,
		_w33819_,
		_w33821_
	);
	LUT2 #(
		.INIT('h8)
	) name29775 (
		_w33820_,
		_w33821_,
		_w33822_
	);
	LUT2 #(
		.INIT('h4)
	) name29776 (
		_w21592_,
		_w33822_,
		_w33823_
	);
	LUT2 #(
		.INIT('h4)
	) name29777 (
		_w33815_,
		_w33823_,
		_w33824_
	);
	LUT2 #(
		.INIT('h4)
	) name29778 (
		\core_dag_ilm1reg_L_reg[9]/NET0131 ,
		_w21592_,
		_w33825_
	);
	LUT2 #(
		.INIT('h1)
	) name29779 (
		_w33824_,
		_w33825_,
		_w33826_
	);
	LUT2 #(
		.INIT('h2)
	) name29780 (
		_w10638_,
		_w33099_,
		_w33827_
	);
	LUT2 #(
		.INIT('h8)
	) name29781 (
		\core_dag_ilm1reg_L3_we_DO_reg[8]/NET0131 ,
		_w33101_,
		_w33828_
	);
	LUT2 #(
		.INIT('h8)
	) name29782 (
		\core_dag_ilm1reg_L0_we_DO_reg[8]/NET0131 ,
		_w33103_,
		_w33829_
	);
	LUT2 #(
		.INIT('h8)
	) name29783 (
		\core_dag_ilm1reg_L1_we_DO_reg[8]/NET0131 ,
		_w33105_,
		_w33830_
	);
	LUT2 #(
		.INIT('h8)
	) name29784 (
		\core_dag_ilm1reg_L2_we_DO_reg[8]/NET0131 ,
		_w33107_,
		_w33831_
	);
	LUT2 #(
		.INIT('h1)
	) name29785 (
		_w33828_,
		_w33829_,
		_w33832_
	);
	LUT2 #(
		.INIT('h1)
	) name29786 (
		_w33830_,
		_w33831_,
		_w33833_
	);
	LUT2 #(
		.INIT('h8)
	) name29787 (
		_w33832_,
		_w33833_,
		_w33834_
	);
	LUT2 #(
		.INIT('h4)
	) name29788 (
		_w21592_,
		_w33834_,
		_w33835_
	);
	LUT2 #(
		.INIT('h4)
	) name29789 (
		_w33827_,
		_w33835_,
		_w33836_
	);
	LUT2 #(
		.INIT('h4)
	) name29790 (
		\core_dag_ilm1reg_L_reg[8]/NET0131 ,
		_w21592_,
		_w33837_
	);
	LUT2 #(
		.INIT('h1)
	) name29791 (
		_w33836_,
		_w33837_,
		_w33838_
	);
	LUT2 #(
		.INIT('h2)
	) name29792 (
		_w7340_,
		_w33099_,
		_w33839_
	);
	LUT2 #(
		.INIT('h8)
	) name29793 (
		\core_dag_ilm1reg_L3_we_DO_reg[13]/NET0131 ,
		_w33101_,
		_w33840_
	);
	LUT2 #(
		.INIT('h8)
	) name29794 (
		\core_dag_ilm1reg_L0_we_DO_reg[13]/NET0131 ,
		_w33103_,
		_w33841_
	);
	LUT2 #(
		.INIT('h8)
	) name29795 (
		\core_dag_ilm1reg_L1_we_DO_reg[13]/NET0131 ,
		_w33105_,
		_w33842_
	);
	LUT2 #(
		.INIT('h8)
	) name29796 (
		\core_dag_ilm1reg_L2_we_DO_reg[13]/NET0131 ,
		_w33107_,
		_w33843_
	);
	LUT2 #(
		.INIT('h1)
	) name29797 (
		_w33840_,
		_w33841_,
		_w33844_
	);
	LUT2 #(
		.INIT('h1)
	) name29798 (
		_w33842_,
		_w33843_,
		_w33845_
	);
	LUT2 #(
		.INIT('h8)
	) name29799 (
		_w33844_,
		_w33845_,
		_w33846_
	);
	LUT2 #(
		.INIT('h4)
	) name29800 (
		_w21592_,
		_w33846_,
		_w33847_
	);
	LUT2 #(
		.INIT('h4)
	) name29801 (
		_w33839_,
		_w33847_,
		_w33848_
	);
	LUT2 #(
		.INIT('h4)
	) name29802 (
		\core_dag_ilm1reg_L_reg[13]/NET0131 ,
		_w21592_,
		_w33849_
	);
	LUT2 #(
		.INIT('h1)
	) name29803 (
		_w33848_,
		_w33849_,
		_w33850_
	);
	LUT2 #(
		.INIT('h2)
	) name29804 (
		_w9178_,
		_w33099_,
		_w33851_
	);
	LUT2 #(
		.INIT('h8)
	) name29805 (
		\core_dag_ilm1reg_L3_we_DO_reg[12]/NET0131 ,
		_w33101_,
		_w33852_
	);
	LUT2 #(
		.INIT('h8)
	) name29806 (
		\core_dag_ilm1reg_L0_we_DO_reg[12]/NET0131 ,
		_w33103_,
		_w33853_
	);
	LUT2 #(
		.INIT('h8)
	) name29807 (
		\core_dag_ilm1reg_L1_we_DO_reg[12]/NET0131 ,
		_w33105_,
		_w33854_
	);
	LUT2 #(
		.INIT('h8)
	) name29808 (
		\core_dag_ilm1reg_L2_we_DO_reg[12]/NET0131 ,
		_w33107_,
		_w33855_
	);
	LUT2 #(
		.INIT('h1)
	) name29809 (
		_w33852_,
		_w33853_,
		_w33856_
	);
	LUT2 #(
		.INIT('h1)
	) name29810 (
		_w33854_,
		_w33855_,
		_w33857_
	);
	LUT2 #(
		.INIT('h8)
	) name29811 (
		_w33856_,
		_w33857_,
		_w33858_
	);
	LUT2 #(
		.INIT('h4)
	) name29812 (
		_w21592_,
		_w33858_,
		_w33859_
	);
	LUT2 #(
		.INIT('h4)
	) name29813 (
		_w33851_,
		_w33859_,
		_w33860_
	);
	LUT2 #(
		.INIT('h4)
	) name29814 (
		\core_dag_ilm1reg_L_reg[12]/NET0131 ,
		_w21592_,
		_w33861_
	);
	LUT2 #(
		.INIT('h1)
	) name29815 (
		_w33860_,
		_w33861_,
		_w33862_
	);
	LUT2 #(
		.INIT('h2)
	) name29816 (
		_w8460_,
		_w33099_,
		_w33863_
	);
	LUT2 #(
		.INIT('h8)
	) name29817 (
		\core_dag_ilm1reg_L1_we_DO_reg[11]/NET0131 ,
		_w33105_,
		_w33864_
	);
	LUT2 #(
		.INIT('h8)
	) name29818 (
		\core_dag_ilm1reg_L2_we_DO_reg[11]/NET0131 ,
		_w33107_,
		_w33865_
	);
	LUT2 #(
		.INIT('h8)
	) name29819 (
		\core_dag_ilm1reg_L3_we_DO_reg[11]/NET0131 ,
		_w33101_,
		_w33866_
	);
	LUT2 #(
		.INIT('h8)
	) name29820 (
		\core_dag_ilm1reg_L0_we_DO_reg[11]/NET0131 ,
		_w33103_,
		_w33867_
	);
	LUT2 #(
		.INIT('h1)
	) name29821 (
		_w33864_,
		_w33865_,
		_w33868_
	);
	LUT2 #(
		.INIT('h1)
	) name29822 (
		_w33866_,
		_w33867_,
		_w33869_
	);
	LUT2 #(
		.INIT('h8)
	) name29823 (
		_w33868_,
		_w33869_,
		_w33870_
	);
	LUT2 #(
		.INIT('h4)
	) name29824 (
		_w21592_,
		_w33870_,
		_w33871_
	);
	LUT2 #(
		.INIT('h4)
	) name29825 (
		_w33863_,
		_w33871_,
		_w33872_
	);
	LUT2 #(
		.INIT('h4)
	) name29826 (
		\core_dag_ilm1reg_L_reg[11]/NET0131 ,
		_w21592_,
		_w33873_
	);
	LUT2 #(
		.INIT('h1)
	) name29827 (
		_w33872_,
		_w33873_,
		_w33874_
	);
	LUT2 #(
		.INIT('h2)
	) name29828 (
		_w7859_,
		_w33099_,
		_w33875_
	);
	LUT2 #(
		.INIT('h8)
	) name29829 (
		\core_dag_ilm1reg_L1_we_DO_reg[10]/NET0131 ,
		_w33105_,
		_w33876_
	);
	LUT2 #(
		.INIT('h8)
	) name29830 (
		\core_dag_ilm1reg_L2_we_DO_reg[10]/NET0131 ,
		_w33107_,
		_w33877_
	);
	LUT2 #(
		.INIT('h8)
	) name29831 (
		\core_dag_ilm1reg_L3_we_DO_reg[10]/NET0131 ,
		_w33101_,
		_w33878_
	);
	LUT2 #(
		.INIT('h8)
	) name29832 (
		\core_dag_ilm1reg_L0_we_DO_reg[10]/NET0131 ,
		_w33103_,
		_w33879_
	);
	LUT2 #(
		.INIT('h1)
	) name29833 (
		_w33876_,
		_w33877_,
		_w33880_
	);
	LUT2 #(
		.INIT('h1)
	) name29834 (
		_w33878_,
		_w33879_,
		_w33881_
	);
	LUT2 #(
		.INIT('h8)
	) name29835 (
		_w33880_,
		_w33881_,
		_w33882_
	);
	LUT2 #(
		.INIT('h4)
	) name29836 (
		_w21592_,
		_w33882_,
		_w33883_
	);
	LUT2 #(
		.INIT('h4)
	) name29837 (
		_w33875_,
		_w33883_,
		_w33884_
	);
	LUT2 #(
		.INIT('h4)
	) name29838 (
		\core_dag_ilm1reg_L_reg[10]/NET0131 ,
		_w21592_,
		_w33885_
	);
	LUT2 #(
		.INIT('h1)
	) name29839 (
		_w33884_,
		_w33885_,
		_w33886_
	);
	LUT2 #(
		.INIT('h8)
	) name29840 (
		_w24166_,
		_w33091_,
		_w33887_
	);
	LUT2 #(
		.INIT('h8)
	) name29841 (
		_w24064_,
		_w33089_,
		_w33888_
	);
	LUT2 #(
		.INIT('h8)
	) name29842 (
		_w10398_,
		_w33093_,
		_w33889_
	);
	LUT2 #(
		.INIT('h4)
	) name29843 (
		_w6067_,
		_w33095_,
		_w33890_
	);
	LUT2 #(
		.INIT('h4)
	) name29844 (
		_w6075_,
		_w33089_,
		_w33891_
	);
	LUT2 #(
		.INIT('h4)
	) name29845 (
		_w6058_,
		_w33091_,
		_w33892_
	);
	LUT2 #(
		.INIT('h4)
	) name29846 (
		_w6084_,
		_w33093_,
		_w33893_
	);
	LUT2 #(
		.INIT('h1)
	) name29847 (
		_w33890_,
		_w33891_,
		_w33894_
	);
	LUT2 #(
		.INIT('h1)
	) name29848 (
		_w33892_,
		_w33893_,
		_w33895_
	);
	LUT2 #(
		.INIT('h8)
	) name29849 (
		_w33894_,
		_w33895_,
		_w33896_
	);
	LUT2 #(
		.INIT('h2)
	) name29850 (
		_w24062_,
		_w33896_,
		_w33897_
	);
	LUT2 #(
		.INIT('h8)
	) name29851 (
		_w10402_,
		_w33095_,
		_w33898_
	);
	LUT2 #(
		.INIT('h1)
	) name29852 (
		_w21592_,
		_w33887_,
		_w33899_
	);
	LUT2 #(
		.INIT('h1)
	) name29853 (
		_w33888_,
		_w33889_,
		_w33900_
	);
	LUT2 #(
		.INIT('h4)
	) name29854 (
		_w33898_,
		_w33900_,
		_w33901_
	);
	LUT2 #(
		.INIT('h8)
	) name29855 (
		_w33899_,
		_w33901_,
		_w33902_
	);
	LUT2 #(
		.INIT('h4)
	) name29856 (
		_w33897_,
		_w33902_,
		_w33903_
	);
	LUT2 #(
		.INIT('h4)
	) name29857 (
		\core_dag_ilm1reg_I_reg[8]/NET0131 ,
		_w21592_,
		_w33904_
	);
	LUT2 #(
		.INIT('h1)
	) name29858 (
		_w33903_,
		_w33904_,
		_w33905_
	);
	LUT2 #(
		.INIT('h8)
	) name29859 (
		_w10369_,
		_w33091_,
		_w33906_
	);
	LUT2 #(
		.INIT('h2)
	) name29860 (
		_w24068_,
		_w33896_,
		_w33907_
	);
	LUT2 #(
		.INIT('h8)
	) name29861 (
		_w6075_,
		_w33089_,
		_w33908_
	);
	LUT2 #(
		.INIT('h8)
	) name29862 (
		\core_dag_ilm1reg_I3_we_DO_reg[5]/NET0131 ,
		_w33908_,
		_w33909_
	);
	LUT2 #(
		.INIT('h8)
	) name29863 (
		_w6084_,
		_w33093_,
		_w33910_
	);
	LUT2 #(
		.INIT('h8)
	) name29864 (
		\core_dag_ilm1reg_I2_we_DO_reg[5]/NET0131 ,
		_w33910_,
		_w33911_
	);
	LUT2 #(
		.INIT('h8)
	) name29865 (
		_w24149_,
		_w33095_,
		_w33912_
	);
	LUT2 #(
		.INIT('h1)
	) name29866 (
		_w21592_,
		_w33906_,
		_w33913_
	);
	LUT2 #(
		.INIT('h1)
	) name29867 (
		_w33909_,
		_w33911_,
		_w33914_
	);
	LUT2 #(
		.INIT('h4)
	) name29868 (
		_w33912_,
		_w33914_,
		_w33915_
	);
	LUT2 #(
		.INIT('h8)
	) name29869 (
		_w33913_,
		_w33915_,
		_w33916_
	);
	LUT2 #(
		.INIT('h4)
	) name29870 (
		_w33907_,
		_w33916_,
		_w33917_
	);
	LUT2 #(
		.INIT('h4)
	) name29871 (
		\core_dag_ilm1reg_I_reg[5]/NET0131 ,
		_w21592_,
		_w33918_
	);
	LUT2 #(
		.INIT('h1)
	) name29872 (
		_w33917_,
		_w33918_,
		_w33919_
	);
	LUT2 #(
		.INIT('h2)
	) name29873 (
		_w24074_,
		_w33896_,
		_w33920_
	);
	LUT2 #(
		.INIT('h8)
	) name29874 (
		_w8891_,
		_w33095_,
		_w33921_
	);
	LUT2 #(
		.INIT('h8)
	) name29875 (
		_w6058_,
		_w33091_,
		_w33922_
	);
	LUT2 #(
		.INIT('h8)
	) name29876 (
		\core_dag_ilm1reg_I0_we_DO_reg[1]/NET0131 ,
		_w33922_,
		_w33923_
	);
	LUT2 #(
		.INIT('h8)
	) name29877 (
		\core_dag_ilm1reg_I2_we_DO_reg[1]/NET0131 ,
		_w33910_,
		_w33924_
	);
	LUT2 #(
		.INIT('h8)
	) name29878 (
		\core_dag_ilm1reg_I3_we_DO_reg[1]/NET0131 ,
		_w33908_,
		_w33925_
	);
	LUT2 #(
		.INIT('h1)
	) name29879 (
		_w21592_,
		_w33921_,
		_w33926_
	);
	LUT2 #(
		.INIT('h1)
	) name29880 (
		_w33923_,
		_w33924_,
		_w33927_
	);
	LUT2 #(
		.INIT('h4)
	) name29881 (
		_w33925_,
		_w33927_,
		_w33928_
	);
	LUT2 #(
		.INIT('h8)
	) name29882 (
		_w33926_,
		_w33928_,
		_w33929_
	);
	LUT2 #(
		.INIT('h4)
	) name29883 (
		_w33920_,
		_w33929_,
		_w33930_
	);
	LUT2 #(
		.INIT('h4)
	) name29884 (
		\core_dag_ilm1reg_I_reg[1]/NET0131 ,
		_w21592_,
		_w33931_
	);
	LUT2 #(
		.INIT('h1)
	) name29885 (
		_w33930_,
		_w33931_,
		_w33932_
	);
	LUT2 #(
		.INIT('h8)
	) name29886 (
		_w6136_,
		_w33091_,
		_w33933_
	);
	LUT2 #(
		.INIT('h8)
	) name29887 (
		_w24082_,
		_w33089_,
		_w33934_
	);
	LUT2 #(
		.INIT('h8)
	) name29888 (
		\core_dag_ilm1reg_I2_we_DO_reg[13]/NET0131 ,
		_w33910_,
		_w33935_
	);
	LUT2 #(
		.INIT('h2)
	) name29889 (
		_w24080_,
		_w33896_,
		_w33936_
	);
	LUT2 #(
		.INIT('h8)
	) name29890 (
		_w6067_,
		_w33095_,
		_w33937_
	);
	LUT2 #(
		.INIT('h8)
	) name29891 (
		\core_dag_ilm1reg_I1_we_DO_reg[13]/NET0131 ,
		_w33937_,
		_w33938_
	);
	LUT2 #(
		.INIT('h1)
	) name29892 (
		_w21592_,
		_w33933_,
		_w33939_
	);
	LUT2 #(
		.INIT('h1)
	) name29893 (
		_w33934_,
		_w33935_,
		_w33940_
	);
	LUT2 #(
		.INIT('h4)
	) name29894 (
		_w33938_,
		_w33940_,
		_w33941_
	);
	LUT2 #(
		.INIT('h8)
	) name29895 (
		_w33939_,
		_w33941_,
		_w33942_
	);
	LUT2 #(
		.INIT('h4)
	) name29896 (
		_w33936_,
		_w33942_,
		_w33943_
	);
	LUT2 #(
		.INIT('h4)
	) name29897 (
		\core_dag_ilm1reg_I_reg[13]/NET0131 ,
		_w21592_,
		_w33944_
	);
	LUT2 #(
		.INIT('h1)
	) name29898 (
		_w33943_,
		_w33944_,
		_w33945_
	);
	LUT2 #(
		.INIT('h8)
	) name29899 (
		_w24134_,
		_w33093_,
		_w33946_
	);
	LUT2 #(
		.INIT('h1)
	) name29900 (
		_w24086_,
		_w33896_,
		_w33947_
	);
	LUT2 #(
		.INIT('h8)
	) name29901 (
		\core_dag_ilm1reg_I1_we_DO_reg[12]/NET0131 ,
		_w33937_,
		_w33948_
	);
	LUT2 #(
		.INIT('h8)
	) name29902 (
		_w8869_,
		_w33089_,
		_w33949_
	);
	LUT2 #(
		.INIT('h8)
	) name29903 (
		\core_dag_ilm1reg_I0_we_DO_reg[12]/NET0131 ,
		_w33922_,
		_w33950_
	);
	LUT2 #(
		.INIT('h1)
	) name29904 (
		_w21592_,
		_w33946_,
		_w33951_
	);
	LUT2 #(
		.INIT('h1)
	) name29905 (
		_w33948_,
		_w33949_,
		_w33952_
	);
	LUT2 #(
		.INIT('h4)
	) name29906 (
		_w33950_,
		_w33952_,
		_w33953_
	);
	LUT2 #(
		.INIT('h8)
	) name29907 (
		_w33951_,
		_w33953_,
		_w33954_
	);
	LUT2 #(
		.INIT('h4)
	) name29908 (
		_w33947_,
		_w33954_,
		_w33955_
	);
	LUT2 #(
		.INIT('h4)
	) name29909 (
		\core_dag_ilm1reg_I_reg[12]/NET0131 ,
		_w21592_,
		_w33956_
	);
	LUT2 #(
		.INIT('h1)
	) name29910 (
		_w33955_,
		_w33956_,
		_w33957_
	);
	LUT2 #(
		.INIT('h8)
	) name29911 (
		\core_dag_ilm1reg_I1_we_DO_reg[11]/NET0131 ,
		_w33937_,
		_w33958_
	);
	LUT2 #(
		.INIT('h8)
	) name29912 (
		_w8734_,
		_w33093_,
		_w33959_
	);
	LUT2 #(
		.INIT('h8)
	) name29913 (
		\core_dag_ilm1reg_I3_we_DO_reg[11]/NET0131 ,
		_w33908_,
		_w33960_
	);
	LUT2 #(
		.INIT('h1)
	) name29914 (
		_w24091_,
		_w33896_,
		_w33961_
	);
	LUT2 #(
		.INIT('h8)
	) name29915 (
		\core_dag_ilm1reg_I0_we_DO_reg[11]/NET0131 ,
		_w33922_,
		_w33962_
	);
	LUT2 #(
		.INIT('h1)
	) name29916 (
		_w21592_,
		_w33958_,
		_w33963_
	);
	LUT2 #(
		.INIT('h1)
	) name29917 (
		_w33959_,
		_w33960_,
		_w33964_
	);
	LUT2 #(
		.INIT('h4)
	) name29918 (
		_w33962_,
		_w33964_,
		_w33965_
	);
	LUT2 #(
		.INIT('h8)
	) name29919 (
		_w33963_,
		_w33965_,
		_w33966_
	);
	LUT2 #(
		.INIT('h4)
	) name29920 (
		_w33961_,
		_w33966_,
		_w33967_
	);
	LUT2 #(
		.INIT('h4)
	) name29921 (
		\core_dag_ilm1reg_I_reg[11]/NET0131 ,
		_w21592_,
		_w33968_
	);
	LUT2 #(
		.INIT('h1)
	) name29922 (
		_w33967_,
		_w33968_,
		_w33969_
	);
	LUT2 #(
		.INIT('h8)
	) name29923 (
		\core_dag_ilm1reg_I1_we_DO_reg[10]/NET0131 ,
		_w33937_,
		_w33970_
	);
	LUT2 #(
		.INIT('h8)
	) name29924 (
		_w8133_,
		_w33093_,
		_w33971_
	);
	LUT2 #(
		.INIT('h8)
	) name29925 (
		\core_dag_ilm1reg_I3_we_DO_reg[10]/NET0131 ,
		_w33908_,
		_w33972_
	);
	LUT2 #(
		.INIT('h2)
	) name29926 (
		_w23763_,
		_w33896_,
		_w33973_
	);
	LUT2 #(
		.INIT('h8)
	) name29927 (
		\core_dag_ilm1reg_I0_we_DO_reg[10]/NET0131 ,
		_w33922_,
		_w33974_
	);
	LUT2 #(
		.INIT('h1)
	) name29928 (
		_w21592_,
		_w33970_,
		_w33975_
	);
	LUT2 #(
		.INIT('h1)
	) name29929 (
		_w33971_,
		_w33972_,
		_w33976_
	);
	LUT2 #(
		.INIT('h4)
	) name29930 (
		_w33974_,
		_w33976_,
		_w33977_
	);
	LUT2 #(
		.INIT('h8)
	) name29931 (
		_w33975_,
		_w33977_,
		_w33978_
	);
	LUT2 #(
		.INIT('h4)
	) name29932 (
		_w33973_,
		_w33978_,
		_w33979_
	);
	LUT2 #(
		.INIT('h4)
	) name29933 (
		\core_dag_ilm1reg_I_reg[10]/NET0131 ,
		_w21592_,
		_w33980_
	);
	LUT2 #(
		.INIT('h1)
	) name29934 (
		_w33979_,
		_w33980_,
		_w33981_
	);
	LUT2 #(
		.INIT('h1)
	) name29935 (
		\sice_ICYC_reg[16]/NET0131 ,
		_w20745_,
		_w33982_
	);
	LUT2 #(
		.INIT('h1)
	) name29936 (
		_w20746_,
		_w33982_,
		_w33983_
	);
	LUT2 #(
		.INIT('h2)
	) name29937 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w23920_,
		_w33984_
	);
	LUT2 #(
		.INIT('h4)
	) name29938 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w30142_,
		_w33985_
	);
	LUT2 #(
		.INIT('h1)
	) name29939 (
		_w33984_,
		_w33985_,
		_w33986_
	);
	LUT2 #(
		.INIT('h2)
	) name29940 (
		_w18717_,
		_w33986_,
		_w33987_
	);
	LUT2 #(
		.INIT('h1)
	) name29941 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[12]/P0001 ,
		_w18717_,
		_w33988_
	);
	LUT2 #(
		.INIT('h1)
	) name29942 (
		_w33987_,
		_w33988_,
		_w33989_
	);
	LUT2 #(
		.INIT('h2)
	) name29943 (
		_w17833_,
		_w33986_,
		_w33990_
	);
	LUT2 #(
		.INIT('h1)
	) name29944 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[12]/P0001 ,
		_w17833_,
		_w33991_
	);
	LUT2 #(
		.INIT('h1)
	) name29945 (
		_w33990_,
		_w33991_,
		_w33992_
	);
	LUT2 #(
		.INIT('h2)
	) name29946 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 ,
		_w18266_,
		_w33993_
	);
	LUT2 #(
		.INIT('h1)
	) name29947 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[10]/P0001 ,
		_w18271_,
		_w33994_
	);
	LUT2 #(
		.INIT('h2)
	) name29948 (
		_w18271_,
		_w19848_,
		_w33995_
	);
	LUT2 #(
		.INIT('h2)
	) name29949 (
		_w18273_,
		_w33994_,
		_w33996_
	);
	LUT2 #(
		.INIT('h4)
	) name29950 (
		_w33995_,
		_w33996_,
		_w33997_
	);
	LUT2 #(
		.INIT('h1)
	) name29951 (
		_w18270_,
		_w33993_,
		_w33998_
	);
	LUT2 #(
		.INIT('h4)
	) name29952 (
		_w33997_,
		_w33998_,
		_w33999_
	);
	LUT2 #(
		.INIT('h1)
	) name29953 (
		_w18262_,
		_w33999_,
		_w34000_
	);
	LUT2 #(
		.INIT('h8)
	) name29954 (
		_w18262_,
		_w19643_,
		_w34001_
	);
	LUT2 #(
		.INIT('h1)
	) name29955 (
		_w34000_,
		_w34001_,
		_w34002_
	);
	LUT2 #(
		.INIT('h2)
	) name29956 (
		\sport1_txctl_TXSHT_reg[10]/P0001 ,
		_w22677_,
		_w34003_
	);
	LUT2 #(
		.INIT('h8)
	) name29957 (
		\sport1_txctl_TX_reg[11]/P0001 ,
		_w22677_,
		_w34004_
	);
	LUT2 #(
		.INIT('h1)
	) name29958 (
		_w34003_,
		_w34004_,
		_w34005_
	);
	LUT2 #(
		.INIT('h2)
	) name29959 (
		_w14752_,
		_w19643_,
		_w34006_
	);
	LUT2 #(
		.INIT('h8)
	) name29960 (
		_w18328_,
		_w19848_,
		_w34007_
	);
	LUT2 #(
		.INIT('h2)
	) name29961 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[10]/P0001 ,
		_w18330_,
		_w34008_
	);
	LUT2 #(
		.INIT('h2)
	) name29962 (
		_w18334_,
		_w34008_,
		_w34009_
	);
	LUT2 #(
		.INIT('h4)
	) name29963 (
		_w34007_,
		_w34009_,
		_w34010_
	);
	LUT2 #(
		.INIT('h1)
	) name29964 (
		_w34006_,
		_w34010_,
		_w34011_
	);
	LUT2 #(
		.INIT('h2)
	) name29965 (
		\sport1_rxctl_RCS_reg[1]/NET0131 ,
		_w31705_,
		_w34012_
	);
	LUT2 #(
		.INIT('h2)
	) name29966 (
		\sport0_rxctl_RCS_reg[1]/NET0131 ,
		_w31868_,
		_w34013_
	);
	LUT2 #(
		.INIT('h2)
	) name29967 (
		\sport0_txctl_TXSHT_reg[10]/P0001 ,
		_w19960_,
		_w34014_
	);
	LUT2 #(
		.INIT('h8)
	) name29968 (
		\sport0_txctl_TX_reg[11]/P0001 ,
		_w19960_,
		_w34015_
	);
	LUT2 #(
		.INIT('h1)
	) name29969 (
		_w34014_,
		_w34015_,
		_w34016_
	);
	LUT2 #(
		.INIT('h1)
	) name29970 (
		\sport0_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		_w19538_,
		_w34017_
	);
	LUT2 #(
		.INIT('h1)
	) name29971 (
		_w19544_,
		_w34017_,
		_w34018_
	);
	LUT2 #(
		.INIT('h8)
	) name29972 (
		_w19197_,
		_w34018_,
		_w34019_
	);
	LUT2 #(
		.INIT('h1)
	) name29973 (
		\sport0_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		_w19535_,
		_w34020_
	);
	LUT2 #(
		.INIT('h1)
	) name29974 (
		_w19536_,
		_w34020_,
		_w34021_
	);
	LUT2 #(
		.INIT('h8)
	) name29975 (
		_w19197_,
		_w34021_,
		_w34022_
	);
	LUT2 #(
		.INIT('h4)
	) name29976 (
		\core_c_dec_MFDAG2_Ei_reg/NET0131 ,
		_w4117_,
		_w34023_
	);
	LUT2 #(
		.INIT('h4)
	) name29977 (
		_w30936_,
		_w31263_,
		_w34024_
	);
	LUT2 #(
		.INIT('h8)
	) name29978 (
		_w31265_,
		_w34024_,
		_w34025_
	);
	LUT2 #(
		.INIT('h8)
	) name29979 (
		_w31270_,
		_w34025_,
		_w34026_
	);
	LUT2 #(
		.INIT('h8)
	) name29980 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w34024_,
		_w34027_
	);
	LUT2 #(
		.INIT('h4)
	) name29981 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w34027_,
		_w34028_
	);
	LUT2 #(
		.INIT('h4)
	) name29982 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w34029_
	);
	LUT2 #(
		.INIT('h8)
	) name29983 (
		_w34024_,
		_w34029_,
		_w34030_
	);
	LUT2 #(
		.INIT('h1)
	) name29984 (
		_w34028_,
		_w34030_,
		_w34031_
	);
	LUT2 #(
		.INIT('h2)
	) name29985 (
		_w31271_,
		_w34031_,
		_w34032_
	);
	LUT2 #(
		.INIT('h8)
	) name29986 (
		_w32024_,
		_w34028_,
		_w34033_
	);
	LUT2 #(
		.INIT('h1)
	) name29987 (
		_w4117_,
		_w34033_,
		_w34034_
	);
	LUT2 #(
		.INIT('h8)
	) name29988 (
		_w32024_,
		_w34025_,
		_w34035_
	);
	LUT2 #(
		.INIT('h4)
	) name29989 (
		_w31653_,
		_w31979_,
		_w34036_
	);
	LUT2 #(
		.INIT('h8)
	) name29990 (
		_w6095_,
		_w19298_,
		_w34037_
	);
	LUT2 #(
		.INIT('h4)
	) name29991 (
		_w31269_,
		_w34037_,
		_w34038_
	);
	LUT2 #(
		.INIT('h1)
	) name29992 (
		_w34036_,
		_w34038_,
		_w34039_
	);
	LUT2 #(
		.INIT('h2)
	) name29993 (
		_w34024_,
		_w34039_,
		_w34040_
	);
	LUT2 #(
		.INIT('h2)
	) name29994 (
		_w6091_,
		_w31269_,
		_w34041_
	);
	LUT2 #(
		.INIT('h8)
	) name29995 (
		_w34027_,
		_w34041_,
		_w34042_
	);
	LUT2 #(
		.INIT('h1)
	) name29996 (
		_w34026_,
		_w34035_,
		_w34043_
	);
	LUT2 #(
		.INIT('h4)
	) name29997 (
		_w34042_,
		_w34043_,
		_w34044_
	);
	LUT2 #(
		.INIT('h4)
	) name29998 (
		_w34032_,
		_w34044_,
		_w34045_
	);
	LUT2 #(
		.INIT('h2)
	) name29999 (
		_w34034_,
		_w34040_,
		_w34046_
	);
	LUT2 #(
		.INIT('h8)
	) name30000 (
		_w34045_,
		_w34046_,
		_w34047_
	);
	LUT2 #(
		.INIT('h1)
	) name30001 (
		_w34023_,
		_w34047_,
		_w34048_
	);
	LUT2 #(
		.INIT('h1)
	) name30002 (
		\sport1_cfg_SCLKi_cnt_reg[6]/NET0131 ,
		_w20235_,
		_w34049_
	);
	LUT2 #(
		.INIT('h1)
	) name30003 (
		_w20236_,
		_w34049_,
		_w34050_
	);
	LUT2 #(
		.INIT('h8)
	) name30004 (
		_w19130_,
		_w34050_,
		_w34051_
	);
	LUT2 #(
		.INIT('h1)
	) name30005 (
		\sport1_cfg_SCLKi_cnt_reg[4]/NET0131 ,
		_w20233_,
		_w34052_
	);
	LUT2 #(
		.INIT('h1)
	) name30006 (
		_w20234_,
		_w34052_,
		_w34053_
	);
	LUT2 #(
		.INIT('h8)
	) name30007 (
		_w19130_,
		_w34053_,
		_w34054_
	);
	LUT2 #(
		.INIT('h2)
	) name30008 (
		\core_c_psq_SSTAT_reg[2]/NET0131 ,
		_w13778_,
		_w34055_
	);
	LUT2 #(
		.INIT('h1)
	) name30009 (
		_w33341_,
		_w34055_,
		_w34056_
	);
	LUT2 #(
		.INIT('h8)
	) name30010 (
		_w33337_,
		_w33341_,
		_w34057_
	);
	LUT2 #(
		.INIT('h1)
	) name30011 (
		_w34056_,
		_w34057_,
		_w34058_
	);
	LUT2 #(
		.INIT('h2)
	) name30012 (
		\bdma_BCTL_reg[0]/NET0131 ,
		_w6914_,
		_w34059_
	);
	LUT2 #(
		.INIT('h1)
	) name30013 (
		_w5733_,
		_w34059_,
		_w34060_
	);
	LUT2 #(
		.INIT('h2)
	) name30014 (
		_w19923_,
		_w34060_,
		_w34061_
	);
	LUT2 #(
		.INIT('h4)
	) name30015 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		_w34062_
	);
	LUT2 #(
		.INIT('h1)
	) name30016 (
		_w34061_,
		_w34062_,
		_w34063_
	);
	LUT2 #(
		.INIT('h1)
	) name30017 (
		_w5729_,
		_w34059_,
		_w34064_
	);
	LUT2 #(
		.INIT('h1)
	) name30018 (
		_w13146_,
		_w34064_,
		_w34065_
	);
	LUT2 #(
		.INIT('h2)
	) name30019 (
		_w19923_,
		_w34065_,
		_w34066_
	);
	LUT2 #(
		.INIT('h1)
	) name30020 (
		_w25024_,
		_w34066_,
		_w34067_
	);
	LUT2 #(
		.INIT('h4)
	) name30021 (
		_w34063_,
		_w34067_,
		_w34068_
	);
	LUT2 #(
		.INIT('h2)
	) name30022 (
		\bdma_BRdataBUF_reg[0]/P0001 ,
		_w34068_,
		_w34069_
	);
	LUT2 #(
		.INIT('h8)
	) name30023 (
		\T_ED[0]_pad ,
		_w34061_,
		_w34070_
	);
	LUT2 #(
		.INIT('h8)
	) name30024 (
		_w34067_,
		_w34070_,
		_w34071_
	);
	LUT2 #(
		.INIT('h1)
	) name30025 (
		_w34069_,
		_w34071_,
		_w34072_
	);
	LUT2 #(
		.INIT('h2)
	) name30026 (
		\bdma_BWCOUNT_reg[11]/NET0131 ,
		_w33295_,
		_w34073_
	);
	LUT2 #(
		.INIT('h1)
	) name30027 (
		_w13763_,
		_w33296_,
		_w34074_
	);
	LUT2 #(
		.INIT('h4)
	) name30028 (
		_w34073_,
		_w34074_,
		_w34075_
	);
	LUT2 #(
		.INIT('h4)
	) name30029 (
		_w8460_,
		_w13763_,
		_w34076_
	);
	LUT2 #(
		.INIT('h1)
	) name30030 (
		_w34075_,
		_w34076_,
		_w34077_
	);
	LUT2 #(
		.INIT('h8)
	) name30031 (
		_w7232_,
		_w20764_,
		_w34078_
	);
	LUT2 #(
		.INIT('h2)
	) name30032 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w13755_,
		_w34079_
	);
	LUT2 #(
		.INIT('h8)
	) name30033 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w34079_,
		_w34080_
	);
	LUT2 #(
		.INIT('h8)
	) name30034 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w34080_,
		_w34081_
	);
	LUT2 #(
		.INIT('h8)
	) name30035 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w34081_,
		_w34082_
	);
	LUT2 #(
		.INIT('h8)
	) name30036 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w34082_,
		_w34083_
	);
	LUT2 #(
		.INIT('h8)
	) name30037 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w34083_,
		_w34084_
	);
	LUT2 #(
		.INIT('h8)
	) name30038 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w34084_,
		_w34085_
	);
	LUT2 #(
		.INIT('h8)
	) name30039 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w34085_,
		_w34086_
	);
	LUT2 #(
		.INIT('h8)
	) name30040 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w34086_,
		_w34087_
	);
	LUT2 #(
		.INIT('h8)
	) name30041 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w34087_,
		_w34088_
	);
	LUT2 #(
		.INIT('h8)
	) name30042 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w34088_,
		_w34089_
	);
	LUT2 #(
		.INIT('h8)
	) name30043 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w34089_,
		_w34090_
	);
	LUT2 #(
		.INIT('h1)
	) name30044 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w34090_,
		_w34091_
	);
	LUT2 #(
		.INIT('h8)
	) name30045 (
		\bdma_BIAD_reg[12]/NET0131 ,
		_w34090_,
		_w34092_
	);
	LUT2 #(
		.INIT('h1)
	) name30046 (
		_w34078_,
		_w34091_,
		_w34093_
	);
	LUT2 #(
		.INIT('h4)
	) name30047 (
		_w34092_,
		_w34093_,
		_w34094_
	);
	LUT2 #(
		.INIT('h8)
	) name30048 (
		_w9178_,
		_w34078_,
		_w34095_
	);
	LUT2 #(
		.INIT('h1)
	) name30049 (
		_w34094_,
		_w34095_,
		_w34096_
	);
	LUT2 #(
		.INIT('h1)
	) name30050 (
		\bdma_BIAD_reg[11]/NET0131 ,
		_w34089_,
		_w34097_
	);
	LUT2 #(
		.INIT('h1)
	) name30051 (
		_w34078_,
		_w34090_,
		_w34098_
	);
	LUT2 #(
		.INIT('h4)
	) name30052 (
		_w34097_,
		_w34098_,
		_w34099_
	);
	LUT2 #(
		.INIT('h8)
	) name30053 (
		_w8460_,
		_w34078_,
		_w34100_
	);
	LUT2 #(
		.INIT('h1)
	) name30054 (
		_w34099_,
		_w34100_,
		_w34101_
	);
	LUT2 #(
		.INIT('h2)
	) name30055 (
		\bdma_BEAD_reg[13]/NET0131 ,
		_w33314_,
		_w34102_
	);
	LUT2 #(
		.INIT('h4)
	) name30056 (
		\bdma_BEAD_reg[13]/NET0131 ,
		_w33314_,
		_w34103_
	);
	LUT2 #(
		.INIT('h1)
	) name30057 (
		_w34102_,
		_w34103_,
		_w34104_
	);
	LUT2 #(
		.INIT('h1)
	) name30058 (
		_w20765_,
		_w34104_,
		_w34105_
	);
	LUT2 #(
		.INIT('h8)
	) name30059 (
		_w7340_,
		_w20765_,
		_w34106_
	);
	LUT2 #(
		.INIT('h1)
	) name30060 (
		_w34105_,
		_w34106_,
		_w34107_
	);
	LUT2 #(
		.INIT('h1)
	) name30061 (
		\bdma_BEAD_reg[11]/NET0131 ,
		_w33312_,
		_w34108_
	);
	LUT2 #(
		.INIT('h1)
	) name30062 (
		_w20765_,
		_w33313_,
		_w34109_
	);
	LUT2 #(
		.INIT('h4)
	) name30063 (
		_w34108_,
		_w34109_,
		_w34110_
	);
	LUT2 #(
		.INIT('h8)
	) name30064 (
		_w8460_,
		_w20765_,
		_w34111_
	);
	LUT2 #(
		.INIT('h1)
	) name30065 (
		_w34110_,
		_w34111_,
		_w34112_
	);
	LUT2 #(
		.INIT('h2)
	) name30066 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w10638_,
		_w34113_
	);
	LUT2 #(
		.INIT('h8)
	) name30067 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001 ,
		_w14704_,
		_w34114_
	);
	LUT2 #(
		.INIT('h8)
	) name30068 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001 ,
		_w14699_,
		_w34115_
	);
	LUT2 #(
		.INIT('h8)
	) name30069 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001 ,
		_w14706_,
		_w34116_
	);
	LUT2 #(
		.INIT('h8)
	) name30070 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001 ,
		_w14711_,
		_w34117_
	);
	LUT2 #(
		.INIT('h8)
	) name30071 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][23]/P0001 ,
		_w14713_,
		_w34118_
	);
	LUT2 #(
		.INIT('h8)
	) name30072 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][23]/P0001 ,
		_w14702_,
		_w34119_
	);
	LUT2 #(
		.INIT('h8)
	) name30073 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][23]/P0001 ,
		_w14708_,
		_w34120_
	);
	LUT2 #(
		.INIT('h1)
	) name30074 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w34114_,
		_w34121_
	);
	LUT2 #(
		.INIT('h1)
	) name30075 (
		_w34115_,
		_w34116_,
		_w34122_
	);
	LUT2 #(
		.INIT('h1)
	) name30076 (
		_w34117_,
		_w34118_,
		_w34123_
	);
	LUT2 #(
		.INIT('h1)
	) name30077 (
		_w34119_,
		_w34120_,
		_w34124_
	);
	LUT2 #(
		.INIT('h8)
	) name30078 (
		_w34123_,
		_w34124_,
		_w34125_
	);
	LUT2 #(
		.INIT('h8)
	) name30079 (
		_w34121_,
		_w34122_,
		_w34126_
	);
	LUT2 #(
		.INIT('h8)
	) name30080 (
		_w34125_,
		_w34126_,
		_w34127_
	);
	LUT2 #(
		.INIT('h1)
	) name30081 (
		_w34113_,
		_w34127_,
		_w34128_
	);
	LUT2 #(
		.INIT('h8)
	) name30082 (
		_w32367_,
		_w34128_,
		_w34129_
	);
	LUT2 #(
		.INIT('h2)
	) name30083 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w33494_,
		_w34130_
	);
	LUT2 #(
		.INIT('h2)
	) name30084 (
		_w32364_,
		_w34130_,
		_w34131_
	);
	LUT2 #(
		.INIT('h2)
	) name30085 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w34131_,
		_w34132_
	);
	LUT2 #(
		.INIT('h4)
	) name30086 (
		_w32367_,
		_w34132_,
		_w34133_
	);
	LUT2 #(
		.INIT('h1)
	) name30087 (
		_w34129_,
		_w34133_,
		_w34134_
	);
	LUT2 #(
		.INIT('h2)
	) name30088 (
		\bdma_BRdataBUF_reg[5]/P0001 ,
		_w34068_,
		_w34135_
	);
	LUT2 #(
		.INIT('h2)
	) name30089 (
		\T_ED[5]_pad ,
		_w25024_,
		_w34136_
	);
	LUT2 #(
		.INIT('h8)
	) name30090 (
		_w34061_,
		_w34136_,
		_w34137_
	);
	LUT2 #(
		.INIT('h1)
	) name30091 (
		_w34135_,
		_w34137_,
		_w34138_
	);
	LUT2 #(
		.INIT('h2)
	) name30092 (
		\bdma_BRdataBUF_reg[7]/P0001 ,
		_w34068_,
		_w34139_
	);
	LUT2 #(
		.INIT('h2)
	) name30093 (
		\T_ED[7]_pad ,
		_w25024_,
		_w34140_
	);
	LUT2 #(
		.INIT('h8)
	) name30094 (
		_w34061_,
		_w34140_,
		_w34141_
	);
	LUT2 #(
		.INIT('h1)
	) name30095 (
		_w34139_,
		_w34141_,
		_w34142_
	);
	LUT2 #(
		.INIT('h2)
	) name30096 (
		\bdma_BRdataBUF_reg[4]/P0001 ,
		_w34068_,
		_w34143_
	);
	LUT2 #(
		.INIT('h2)
	) name30097 (
		\T_ED[4]_pad ,
		_w25024_,
		_w34144_
	);
	LUT2 #(
		.INIT('h8)
	) name30098 (
		_w34061_,
		_w34144_,
		_w34145_
	);
	LUT2 #(
		.INIT('h1)
	) name30099 (
		_w34143_,
		_w34145_,
		_w34146_
	);
	LUT2 #(
		.INIT('h2)
	) name30100 (
		\bdma_BRdataBUF_reg[6]/P0001 ,
		_w34068_,
		_w34147_
	);
	LUT2 #(
		.INIT('h2)
	) name30101 (
		\T_ED[6]_pad ,
		_w25024_,
		_w34148_
	);
	LUT2 #(
		.INIT('h8)
	) name30102 (
		_w34061_,
		_w34148_,
		_w34149_
	);
	LUT2 #(
		.INIT('h1)
	) name30103 (
		_w34147_,
		_w34149_,
		_w34150_
	);
	LUT2 #(
		.INIT('h2)
	) name30104 (
		\bdma_BRdataBUF_reg[3]/P0001 ,
		_w34068_,
		_w34151_
	);
	LUT2 #(
		.INIT('h2)
	) name30105 (
		\T_ED[3]_pad ,
		_w25024_,
		_w34152_
	);
	LUT2 #(
		.INIT('h8)
	) name30106 (
		_w34061_,
		_w34152_,
		_w34153_
	);
	LUT2 #(
		.INIT('h1)
	) name30107 (
		_w34151_,
		_w34153_,
		_w34154_
	);
	LUT2 #(
		.INIT('h2)
	) name30108 (
		\bdma_BRdataBUF_reg[2]/P0001 ,
		_w34068_,
		_w34155_
	);
	LUT2 #(
		.INIT('h2)
	) name30109 (
		\T_ED[2]_pad ,
		_w25024_,
		_w34156_
	);
	LUT2 #(
		.INIT('h8)
	) name30110 (
		_w34061_,
		_w34156_,
		_w34157_
	);
	LUT2 #(
		.INIT('h1)
	) name30111 (
		_w34155_,
		_w34157_,
		_w34158_
	);
	LUT2 #(
		.INIT('h2)
	) name30112 (
		\bdma_BRdataBUF_reg[1]/P0001 ,
		_w34068_,
		_w34159_
	);
	LUT2 #(
		.INIT('h2)
	) name30113 (
		\T_ED[1]_pad ,
		_w25024_,
		_w34160_
	);
	LUT2 #(
		.INIT('h8)
	) name30114 (
		_w34061_,
		_w34160_,
		_w34161_
	);
	LUT2 #(
		.INIT('h1)
	) name30115 (
		_w34159_,
		_w34161_,
		_w34162_
	);
	LUT2 #(
		.INIT('h1)
	) name30116 (
		\sice_ICYC_reg[20]/NET0131 ,
		_w20749_,
		_w34163_
	);
	LUT2 #(
		.INIT('h1)
	) name30117 (
		_w20750_,
		_w34163_,
		_w34164_
	);
	LUT2 #(
		.INIT('h8)
	) name30118 (
		\sice_IIRC_reg[21]/NET0131 ,
		_w32042_,
		_w34165_
	);
	LUT2 #(
		.INIT('h8)
	) name30119 (
		\sice_IIRC_reg[22]/NET0131 ,
		_w34165_,
		_w34166_
	);
	LUT2 #(
		.INIT('h1)
	) name30120 (
		\sice_IIRC_reg[23]/NET0131 ,
		_w34166_,
		_w34167_
	);
	LUT2 #(
		.INIT('h8)
	) name30121 (
		\sice_IIRC_reg[23]/NET0131 ,
		_w34166_,
		_w34168_
	);
	LUT2 #(
		.INIT('h1)
	) name30122 (
		_w34167_,
		_w34168_,
		_w34169_
	);
	LUT2 #(
		.INIT('h1)
	) name30123 (
		\clkc_oscntr_reg_DO_reg[10]/NET0131 ,
		_w23424_,
		_w34170_
	);
	LUT2 #(
		.INIT('h1)
	) name30124 (
		_w33617_,
		_w34170_,
		_w34171_
	);
	LUT2 #(
		.INIT('h2)
	) name30125 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w11265_,
		_w34172_
	);
	LUT2 #(
		.INIT('h8)
	) name30126 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001 ,
		_w14706_,
		_w34173_
	);
	LUT2 #(
		.INIT('h8)
	) name30127 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001 ,
		_w14704_,
		_w34174_
	);
	LUT2 #(
		.INIT('h8)
	) name30128 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][22]/P0001 ,
		_w14702_,
		_w34175_
	);
	LUT2 #(
		.INIT('h8)
	) name30129 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][22]/P0001 ,
		_w14713_,
		_w34176_
	);
	LUT2 #(
		.INIT('h8)
	) name30130 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001 ,
		_w14711_,
		_w34177_
	);
	LUT2 #(
		.INIT('h8)
	) name30131 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][22]/P0001 ,
		_w14708_,
		_w34178_
	);
	LUT2 #(
		.INIT('h8)
	) name30132 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001 ,
		_w14699_,
		_w34179_
	);
	LUT2 #(
		.INIT('h1)
	) name30133 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w34173_,
		_w34180_
	);
	LUT2 #(
		.INIT('h1)
	) name30134 (
		_w34174_,
		_w34175_,
		_w34181_
	);
	LUT2 #(
		.INIT('h1)
	) name30135 (
		_w34176_,
		_w34177_,
		_w34182_
	);
	LUT2 #(
		.INIT('h1)
	) name30136 (
		_w34178_,
		_w34179_,
		_w34183_
	);
	LUT2 #(
		.INIT('h8)
	) name30137 (
		_w34182_,
		_w34183_,
		_w34184_
	);
	LUT2 #(
		.INIT('h8)
	) name30138 (
		_w34180_,
		_w34181_,
		_w34185_
	);
	LUT2 #(
		.INIT('h8)
	) name30139 (
		_w34184_,
		_w34185_,
		_w34186_
	);
	LUT2 #(
		.INIT('h1)
	) name30140 (
		_w34172_,
		_w34186_,
		_w34187_
	);
	LUT2 #(
		.INIT('h8)
	) name30141 (
		_w32367_,
		_w34187_,
		_w34188_
	);
	LUT2 #(
		.INIT('h2)
	) name30142 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w33493_,
		_w34189_
	);
	LUT2 #(
		.INIT('h2)
	) name30143 (
		_w32364_,
		_w34189_,
		_w34190_
	);
	LUT2 #(
		.INIT('h2)
	) name30144 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w34190_,
		_w34191_
	);
	LUT2 #(
		.INIT('h4)
	) name30145 (
		_w32367_,
		_w34191_,
		_w34192_
	);
	LUT2 #(
		.INIT('h1)
	) name30146 (
		_w34188_,
		_w34192_,
		_w34193_
	);
	LUT2 #(
		.INIT('h2)
	) name30147 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w8715_,
		_w34194_
	);
	LUT2 #(
		.INIT('h8)
	) name30148 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001 ,
		_w14706_,
		_w34195_
	);
	LUT2 #(
		.INIT('h8)
	) name30149 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001 ,
		_w14704_,
		_w34196_
	);
	LUT2 #(
		.INIT('h8)
	) name30150 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][17]/P0001 ,
		_w14702_,
		_w34197_
	);
	LUT2 #(
		.INIT('h8)
	) name30151 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][17]/P0001 ,
		_w14713_,
		_w34198_
	);
	LUT2 #(
		.INIT('h8)
	) name30152 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001 ,
		_w14711_,
		_w34199_
	);
	LUT2 #(
		.INIT('h8)
	) name30153 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][17]/P0001 ,
		_w14708_,
		_w34200_
	);
	LUT2 #(
		.INIT('h8)
	) name30154 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001 ,
		_w14699_,
		_w34201_
	);
	LUT2 #(
		.INIT('h1)
	) name30155 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w34195_,
		_w34202_
	);
	LUT2 #(
		.INIT('h1)
	) name30156 (
		_w34196_,
		_w34197_,
		_w34203_
	);
	LUT2 #(
		.INIT('h1)
	) name30157 (
		_w34198_,
		_w34199_,
		_w34204_
	);
	LUT2 #(
		.INIT('h1)
	) name30158 (
		_w34200_,
		_w34201_,
		_w34205_
	);
	LUT2 #(
		.INIT('h8)
	) name30159 (
		_w34204_,
		_w34205_,
		_w34206_
	);
	LUT2 #(
		.INIT('h8)
	) name30160 (
		_w34202_,
		_w34203_,
		_w34207_
	);
	LUT2 #(
		.INIT('h8)
	) name30161 (
		_w34206_,
		_w34207_,
		_w34208_
	);
	LUT2 #(
		.INIT('h1)
	) name30162 (
		_w34194_,
		_w34208_,
		_w34209_
	);
	LUT2 #(
		.INIT('h8)
	) name30163 (
		_w32367_,
		_w34209_,
		_w34210_
	);
	LUT2 #(
		.INIT('h2)
	) name30164 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w5299_,
		_w34211_
	);
	LUT2 #(
		.INIT('h2)
	) name30165 (
		_w32364_,
		_w34211_,
		_w34212_
	);
	LUT2 #(
		.INIT('h2)
	) name30166 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w34212_,
		_w34213_
	);
	LUT2 #(
		.INIT('h4)
	) name30167 (
		_w32367_,
		_w34213_,
		_w34214_
	);
	LUT2 #(
		.INIT('h1)
	) name30168 (
		_w34210_,
		_w34214_,
		_w34215_
	);
	LUT2 #(
		.INIT('h1)
	) name30169 (
		\clkc_oscntr_reg_DO_reg[8]/NET0131 ,
		_w23421_,
		_w34216_
	);
	LUT2 #(
		.INIT('h1)
	) name30170 (
		_w23422_,
		_w34216_,
		_w34217_
	);
	LUT2 #(
		.INIT('h2)
	) name30171 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w10069_,
		_w34218_
	);
	LUT2 #(
		.INIT('h8)
	) name30172 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001 ,
		_w14706_,
		_w34219_
	);
	LUT2 #(
		.INIT('h8)
	) name30173 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001 ,
		_w14704_,
		_w34220_
	);
	LUT2 #(
		.INIT('h8)
	) name30174 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][19]/P0001 ,
		_w14702_,
		_w34221_
	);
	LUT2 #(
		.INIT('h8)
	) name30175 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][19]/P0001 ,
		_w14713_,
		_w34222_
	);
	LUT2 #(
		.INIT('h8)
	) name30176 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001 ,
		_w14711_,
		_w34223_
	);
	LUT2 #(
		.INIT('h8)
	) name30177 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][19]/P0001 ,
		_w14708_,
		_w34224_
	);
	LUT2 #(
		.INIT('h8)
	) name30178 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001 ,
		_w14699_,
		_w34225_
	);
	LUT2 #(
		.INIT('h1)
	) name30179 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w34219_,
		_w34226_
	);
	LUT2 #(
		.INIT('h1)
	) name30180 (
		_w34220_,
		_w34221_,
		_w34227_
	);
	LUT2 #(
		.INIT('h1)
	) name30181 (
		_w34222_,
		_w34223_,
		_w34228_
	);
	LUT2 #(
		.INIT('h1)
	) name30182 (
		_w34224_,
		_w34225_,
		_w34229_
	);
	LUT2 #(
		.INIT('h8)
	) name30183 (
		_w34228_,
		_w34229_,
		_w34230_
	);
	LUT2 #(
		.INIT('h8)
	) name30184 (
		_w34226_,
		_w34227_,
		_w34231_
	);
	LUT2 #(
		.INIT('h8)
	) name30185 (
		_w34230_,
		_w34231_,
		_w34232_
	);
	LUT2 #(
		.INIT('h1)
	) name30186 (
		_w34218_,
		_w34232_,
		_w34233_
	);
	LUT2 #(
		.INIT('h8)
	) name30187 (
		_w32367_,
		_w34233_,
		_w34234_
	);
	LUT2 #(
		.INIT('h2)
	) name30188 (
		\core_c_psq_ICNTL_reg_DO_reg[4]/NET0131 ,
		_w33244_,
		_w34235_
	);
	LUT2 #(
		.INIT('h2)
	) name30189 (
		_w32364_,
		_w34235_,
		_w34236_
	);
	LUT2 #(
		.INIT('h2)
	) name30190 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w34236_,
		_w34237_
	);
	LUT2 #(
		.INIT('h4)
	) name30191 (
		_w32367_,
		_w34237_,
		_w34238_
	);
	LUT2 #(
		.INIT('h1)
	) name30192 (
		_w34234_,
		_w34238_,
		_w34239_
	);
	LUT2 #(
		.INIT('h8)
	) name30193 (
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w28876_,
		_w34240_
	);
	LUT2 #(
		.INIT('h1)
	) name30194 (
		\sport0_cfg_FSi_cnt_reg[3]/NET0131 ,
		_w28948_,
		_w34241_
	);
	LUT2 #(
		.INIT('h1)
	) name30195 (
		_w28949_,
		_w34241_,
		_w34242_
	);
	LUT2 #(
		.INIT('h8)
	) name30196 (
		_w28945_,
		_w34242_,
		_w34243_
	);
	LUT2 #(
		.INIT('h1)
	) name30197 (
		_w34240_,
		_w34243_,
		_w34244_
	);
	LUT2 #(
		.INIT('h1)
	) name30198 (
		\sice_ICYC_reg[12]/NET0131 ,
		_w20741_,
		_w34245_
	);
	LUT2 #(
		.INIT('h1)
	) name30199 (
		_w20742_,
		_w34245_,
		_w34246_
	);
	LUT2 #(
		.INIT('h8)
	) name30200 (
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w28786_,
		_w34247_
	);
	LUT2 #(
		.INIT('h1)
	) name30201 (
		\sport1_cfg_FSi_cnt_reg[3]/NET0131 ,
		_w28858_,
		_w34248_
	);
	LUT2 #(
		.INIT('h1)
	) name30202 (
		_w28859_,
		_w34248_,
		_w34249_
	);
	LUT2 #(
		.INIT('h8)
	) name30203 (
		_w28855_,
		_w34249_,
		_w34250_
	);
	LUT2 #(
		.INIT('h1)
	) name30204 (
		_w34247_,
		_w34250_,
		_w34251_
	);
	LUT2 #(
		.INIT('h1)
	) name30205 (
		\sice_IIRC_reg[12]/NET0131 ,
		_w20856_,
		_w34252_
	);
	LUT2 #(
		.INIT('h1)
	) name30206 (
		_w20857_,
		_w34252_,
		_w34253_
	);
	LUT2 #(
		.INIT('h4)
	) name30207 (
		\core_c_dec_Dummy_E_reg/NET0131 ,
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w34254_
	);
	LUT2 #(
		.INIT('h8)
	) name30208 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_dec_IRE_reg[12]/NET0131 ,
		_w34255_
	);
	LUT2 #(
		.INIT('h2)
	) name30209 (
		_w7168_,
		_w29480_,
		_w34256_
	);
	LUT2 #(
		.INIT('h4)
	) name30210 (
		_w7168_,
		_w29480_,
		_w34257_
	);
	LUT2 #(
		.INIT('h8)
	) name30211 (
		_w7983_,
		_w29493_,
		_w34258_
	);
	LUT2 #(
		.INIT('h8)
	) name30212 (
		_w9268_,
		_w26276_,
		_w34259_
	);
	LUT2 #(
		.INIT('h1)
	) name30213 (
		_w9268_,
		_w26276_,
		_w34260_
	);
	LUT2 #(
		.INIT('h2)
	) name30214 (
		_w7365_,
		_w34260_,
		_w34261_
	);
	LUT2 #(
		.INIT('h4)
	) name30215 (
		_w23671_,
		_w34261_,
		_w34262_
	);
	LUT2 #(
		.INIT('h8)
	) name30216 (
		_w8489_,
		_w27488_,
		_w34263_
	);
	LUT2 #(
		.INIT('h1)
	) name30217 (
		_w34259_,
		_w34263_,
		_w34264_
	);
	LUT2 #(
		.INIT('h4)
	) name30218 (
		_w34262_,
		_w34264_,
		_w34265_
	);
	LUT2 #(
		.INIT('h1)
	) name30219 (
		_w7983_,
		_w29493_,
		_w34266_
	);
	LUT2 #(
		.INIT('h1)
	) name30220 (
		_w8489_,
		_w27488_,
		_w34267_
	);
	LUT2 #(
		.INIT('h1)
	) name30221 (
		_w34266_,
		_w34267_,
		_w34268_
	);
	LUT2 #(
		.INIT('h4)
	) name30222 (
		_w34265_,
		_w34268_,
		_w34269_
	);
	LUT2 #(
		.INIT('h1)
	) name30223 (
		_w34257_,
		_w34258_,
		_w34270_
	);
	LUT2 #(
		.INIT('h4)
	) name30224 (
		_w34269_,
		_w34270_,
		_w34271_
	);
	LUT2 #(
		.INIT('h8)
	) name30225 (
		_w23585_,
		_w34255_,
		_w34272_
	);
	LUT2 #(
		.INIT('h8)
	) name30226 (
		_w13803_,
		_w34272_,
		_w34273_
	);
	LUT2 #(
		.INIT('h4)
	) name30227 (
		_w34256_,
		_w34273_,
		_w34274_
	);
	LUT2 #(
		.INIT('h4)
	) name30228 (
		_w34271_,
		_w34274_,
		_w34275_
	);
	LUT2 #(
		.INIT('h1)
	) name30229 (
		_w34254_,
		_w34275_,
		_w34276_
	);
	LUT2 #(
		.INIT('h2)
	) name30230 (
		_w14664_,
		_w34276_,
		_w34277_
	);
	LUT2 #(
		.INIT('h2)
	) name30231 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w9435_,
		_w34278_
	);
	LUT2 #(
		.INIT('h1)
	) name30232 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w26276_,
		_w34279_
	);
	LUT2 #(
		.INIT('h1)
	) name30233 (
		_w34278_,
		_w34279_,
		_w34280_
	);
	LUT2 #(
		.INIT('h2)
	) name30234 (
		_w34277_,
		_w34280_,
		_w34281_
	);
	LUT2 #(
		.INIT('h1)
	) name30235 (
		\core_eu_es_sht_es_reg_SBs_reg[1]/P0001 ,
		_w34277_,
		_w34282_
	);
	LUT2 #(
		.INIT('h1)
	) name30236 (
		_w34281_,
		_w34282_,
		_w34283_
	);
	LUT2 #(
		.INIT('h2)
	) name30237 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w7607_,
		_w34284_
	);
	LUT2 #(
		.INIT('h4)
	) name30238 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w23671_,
		_w34285_
	);
	LUT2 #(
		.INIT('h1)
	) name30239 (
		_w34284_,
		_w34285_,
		_w34286_
	);
	LUT2 #(
		.INIT('h2)
	) name30240 (
		_w34277_,
		_w34286_,
		_w34287_
	);
	LUT2 #(
		.INIT('h1)
	) name30241 (
		\core_eu_es_sht_es_reg_SBs_reg[0]/P0001 ,
		_w34277_,
		_w34288_
	);
	LUT2 #(
		.INIT('h1)
	) name30242 (
		_w34287_,
		_w34288_,
		_w34289_
	);
	LUT2 #(
		.INIT('h2)
	) name30243 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w8113_,
		_w34290_
	);
	LUT2 #(
		.INIT('h1)
	) name30244 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w29493_,
		_w34291_
	);
	LUT2 #(
		.INIT('h1)
	) name30245 (
		_w34290_,
		_w34291_,
		_w34292_
	);
	LUT2 #(
		.INIT('h2)
	) name30246 (
		_w34277_,
		_w34292_,
		_w34293_
	);
	LUT2 #(
		.INIT('h1)
	) name30247 (
		\core_eu_es_sht_es_reg_SBs_reg[3]/P0001 ,
		_w34277_,
		_w34294_
	);
	LUT2 #(
		.INIT('h1)
	) name30248 (
		_w34293_,
		_w34294_,
		_w34295_
	);
	LUT2 #(
		.INIT('h2)
	) name30249 (
		_w13801_,
		_w34276_,
		_w34296_
	);
	LUT2 #(
		.INIT('h4)
	) name30250 (
		_w34292_,
		_w34296_,
		_w34297_
	);
	LUT2 #(
		.INIT('h1)
	) name30251 (
		\core_eu_es_sht_es_reg_SBr_reg[3]/P0001 ,
		_w34296_,
		_w34298_
	);
	LUT2 #(
		.INIT('h1)
	) name30252 (
		_w34297_,
		_w34298_,
		_w34299_
	);
	LUT2 #(
		.INIT('h2)
	) name30253 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w8715_,
		_w34300_
	);
	LUT2 #(
		.INIT('h1)
	) name30254 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w27488_,
		_w34301_
	);
	LUT2 #(
		.INIT('h1)
	) name30255 (
		_w34300_,
		_w34301_,
		_w34302_
	);
	LUT2 #(
		.INIT('h2)
	) name30256 (
		_w34277_,
		_w34302_,
		_w34303_
	);
	LUT2 #(
		.INIT('h1)
	) name30257 (
		\core_eu_es_sht_es_reg_SBs_reg[2]/P0001 ,
		_w34277_,
		_w34304_
	);
	LUT2 #(
		.INIT('h1)
	) name30258 (
		_w34303_,
		_w34304_,
		_w34305_
	);
	LUT2 #(
		.INIT('h2)
	) name30259 (
		_w34296_,
		_w34302_,
		_w34306_
	);
	LUT2 #(
		.INIT('h1)
	) name30260 (
		\core_eu_es_sht_es_reg_SBr_reg[2]/P0001 ,
		_w34296_,
		_w34307_
	);
	LUT2 #(
		.INIT('h1)
	) name30261 (
		_w34306_,
		_w34307_,
		_w34308_
	);
	LUT2 #(
		.INIT('h2)
	) name30262 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w10069_,
		_w34309_
	);
	LUT2 #(
		.INIT('h4)
	) name30263 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w29480_,
		_w34310_
	);
	LUT2 #(
		.INIT('h1)
	) name30264 (
		_w34309_,
		_w34310_,
		_w34311_
	);
	LUT2 #(
		.INIT('h2)
	) name30265 (
		_w34296_,
		_w34311_,
		_w34312_
	);
	LUT2 #(
		.INIT('h1)
	) name30266 (
		\core_eu_es_sht_es_reg_SBr_reg[4]/P0001 ,
		_w34296_,
		_w34313_
	);
	LUT2 #(
		.INIT('h1)
	) name30267 (
		_w34312_,
		_w34313_,
		_w34314_
	);
	LUT2 #(
		.INIT('h4)
	) name30268 (
		_w34280_,
		_w34296_,
		_w34315_
	);
	LUT2 #(
		.INIT('h1)
	) name30269 (
		\core_eu_es_sht_es_reg_SBr_reg[1]/P0001 ,
		_w34296_,
		_w34316_
	);
	LUT2 #(
		.INIT('h1)
	) name30270 (
		_w34315_,
		_w34316_,
		_w34317_
	);
	LUT2 #(
		.INIT('h2)
	) name30271 (
		_w34277_,
		_w34311_,
		_w34318_
	);
	LUT2 #(
		.INIT('h1)
	) name30272 (
		\core_eu_es_sht_es_reg_SBs_reg[4]/P0001 ,
		_w34277_,
		_w34319_
	);
	LUT2 #(
		.INIT('h1)
	) name30273 (
		_w34318_,
		_w34319_,
		_w34320_
	);
	LUT2 #(
		.INIT('h4)
	) name30274 (
		_w34286_,
		_w34296_,
		_w34321_
	);
	LUT2 #(
		.INIT('h1)
	) name30275 (
		\core_eu_es_sht_es_reg_SBr_reg[0]/P0001 ,
		_w34296_,
		_w34322_
	);
	LUT2 #(
		.INIT('h1)
	) name30276 (
		_w34321_,
		_w34322_,
		_w34323_
	);
	LUT2 #(
		.INIT('h2)
	) name30277 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 ,
		_w18266_,
		_w34324_
	);
	LUT2 #(
		.INIT('h1)
	) name30278 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[9]/P0001 ,
		_w18271_,
		_w34325_
	);
	LUT2 #(
		.INIT('h2)
	) name30279 (
		_w18271_,
		_w19504_,
		_w34326_
	);
	LUT2 #(
		.INIT('h2)
	) name30280 (
		_w18273_,
		_w34325_,
		_w34327_
	);
	LUT2 #(
		.INIT('h4)
	) name30281 (
		_w34326_,
		_w34327_,
		_w34328_
	);
	LUT2 #(
		.INIT('h1)
	) name30282 (
		_w18270_,
		_w34324_,
		_w34329_
	);
	LUT2 #(
		.INIT('h4)
	) name30283 (
		_w34328_,
		_w34329_,
		_w34330_
	);
	LUT2 #(
		.INIT('h1)
	) name30284 (
		_w18262_,
		_w34330_,
		_w34331_
	);
	LUT2 #(
		.INIT('h2)
	) name30285 (
		_w18262_,
		_w19646_,
		_w34332_
	);
	LUT2 #(
		.INIT('h1)
	) name30286 (
		_w34331_,
		_w34332_,
		_w34333_
	);
	LUT2 #(
		.INIT('h8)
	) name30287 (
		_w14752_,
		_w19646_,
		_w34334_
	);
	LUT2 #(
		.INIT('h8)
	) name30288 (
		_w18328_,
		_w19504_,
		_w34335_
	);
	LUT2 #(
		.INIT('h2)
	) name30289 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[9]/P0001 ,
		_w18330_,
		_w34336_
	);
	LUT2 #(
		.INIT('h2)
	) name30290 (
		_w18334_,
		_w34336_,
		_w34337_
	);
	LUT2 #(
		.INIT('h4)
	) name30291 (
		_w34335_,
		_w34337_,
		_w34338_
	);
	LUT2 #(
		.INIT('h1)
	) name30292 (
		_w34334_,
		_w34338_,
		_w34339_
	);
	LUT2 #(
		.INIT('h4)
	) name30293 (
		\sport0_rxctl_RXSHT_reg[8]/P0001 ,
		_w20868_,
		_w34340_
	);
	LUT2 #(
		.INIT('h8)
	) name30294 (
		\sport0_rxctl_RX_reg[8]/P0001 ,
		_w20873_,
		_w34341_
	);
	LUT2 #(
		.INIT('h2)
	) name30295 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w20914_,
		_w34342_
	);
	LUT2 #(
		.INIT('h2)
	) name30296 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w34343_
	);
	LUT2 #(
		.INIT('h1)
	) name30297 (
		_w20878_,
		_w34343_,
		_w34344_
	);
	LUT2 #(
		.INIT('h4)
	) name30298 (
		_w34342_,
		_w34344_,
		_w34345_
	);
	LUT2 #(
		.INIT('h1)
	) name30299 (
		_w20905_,
		_w34345_,
		_w34346_
	);
	LUT2 #(
		.INIT('h1)
	) name30300 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w34346_,
		_w34347_
	);
	LUT2 #(
		.INIT('h2)
	) name30301 (
		\sport0_rxctl_RX_reg[0]/P0001 ,
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w34348_
	);
	LUT2 #(
		.INIT('h2)
	) name30302 (
		_w31045_,
		_w34348_,
		_w34349_
	);
	LUT2 #(
		.INIT('h1)
	) name30303 (
		_w34347_,
		_w34349_,
		_w34350_
	);
	LUT2 #(
		.INIT('h2)
	) name30304 (
		_w20882_,
		_w34350_,
		_w34351_
	);
	LUT2 #(
		.INIT('h4)
	) name30305 (
		_w20882_,
		_w31037_,
		_w34352_
	);
	LUT2 #(
		.INIT('h1)
	) name30306 (
		_w34351_,
		_w34352_,
		_w34353_
	);
	LUT2 #(
		.INIT('h8)
	) name30307 (
		_w31031_,
		_w34353_,
		_w34354_
	);
	LUT2 #(
		.INIT('h1)
	) name30308 (
		_w20925_,
		_w20926_,
		_w34355_
	);
	LUT2 #(
		.INIT('h1)
	) name30309 (
		\sport0_rxctl_RX_reg[4]/P0001 ,
		_w34355_,
		_w34356_
	);
	LUT2 #(
		.INIT('h1)
	) name30310 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20931_,
		_w34357_
	);
	LUT2 #(
		.INIT('h4)
	) name30311 (
		_w34356_,
		_w34357_,
		_w34358_
	);
	LUT2 #(
		.INIT('h2)
	) name30312 (
		_w20882_,
		_w34358_,
		_w34359_
	);
	LUT2 #(
		.INIT('h4)
	) name30313 (
		_w20882_,
		_w34350_,
		_w34360_
	);
	LUT2 #(
		.INIT('h1)
	) name30314 (
		_w34359_,
		_w34360_,
		_w34361_
	);
	LUT2 #(
		.INIT('h4)
	) name30315 (
		_w34354_,
		_w34361_,
		_w34362_
	);
	LUT2 #(
		.INIT('h2)
	) name30316 (
		_w34354_,
		_w34361_,
		_w34363_
	);
	LUT2 #(
		.INIT('h1)
	) name30317 (
		_w34362_,
		_w34363_,
		_w34364_
	);
	LUT2 #(
		.INIT('h8)
	) name30318 (
		_w31043_,
		_w34353_,
		_w34365_
	);
	LUT2 #(
		.INIT('h1)
	) name30319 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w34365_,
		_w34366_
	);
	LUT2 #(
		.INIT('h4)
	) name30320 (
		_w34364_,
		_w34366_,
		_w34367_
	);
	LUT2 #(
		.INIT('h2)
	) name30321 (
		_w34364_,
		_w34366_,
		_w34368_
	);
	LUT2 #(
		.INIT('h2)
	) name30322 (
		_w20875_,
		_w34367_,
		_w34369_
	);
	LUT2 #(
		.INIT('h4)
	) name30323 (
		_w34368_,
		_w34369_,
		_w34370_
	);
	LUT2 #(
		.INIT('h4)
	) name30324 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w10638_,
		_w34371_
	);
	LUT2 #(
		.INIT('h1)
	) name30325 (
		_w20868_,
		_w34341_,
		_w34372_
	);
	LUT2 #(
		.INIT('h4)
	) name30326 (
		_w34371_,
		_w34372_,
		_w34373_
	);
	LUT2 #(
		.INIT('h4)
	) name30327 (
		_w34370_,
		_w34373_,
		_w34374_
	);
	LUT2 #(
		.INIT('h1)
	) name30328 (
		_w20871_,
		_w34340_,
		_w34375_
	);
	LUT2 #(
		.INIT('h4)
	) name30329 (
		_w34374_,
		_w34375_,
		_w34376_
	);
	LUT2 #(
		.INIT('h8)
	) name30330 (
		\sport0_rxctl_RX_reg[8]/P0001 ,
		_w20871_,
		_w34377_
	);
	LUT2 #(
		.INIT('h1)
	) name30331 (
		_w34376_,
		_w34377_,
		_w34378_
	);
	LUT2 #(
		.INIT('h4)
	) name30332 (
		_w17796_,
		_w18262_,
		_w34379_
	);
	LUT2 #(
		.INIT('h1)
	) name30333 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 ,
		_w28530_,
		_w34380_
	);
	LUT2 #(
		.INIT('h2)
	) name30334 (
		_w17814_,
		_w19381_,
		_w34381_
	);
	LUT2 #(
		.INIT('h2)
	) name30335 (
		_w28534_,
		_w34381_,
		_w34382_
	);
	LUT2 #(
		.INIT('h1)
	) name30336 (
		_w34380_,
		_w34382_,
		_w34383_
	);
	LUT2 #(
		.INIT('h1)
	) name30337 (
		_w19385_,
		_w34383_,
		_w34384_
	);
	LUT2 #(
		.INIT('h1)
	) name30338 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[2]/P0001 ,
		_w28532_,
		_w34385_
	);
	LUT2 #(
		.INIT('h1)
	) name30339 (
		_w34384_,
		_w34385_,
		_w34386_
	);
	LUT2 #(
		.INIT('h2)
	) name30340 (
		_w28529_,
		_w34386_,
		_w34387_
	);
	LUT2 #(
		.INIT('h1)
	) name30341 (
		_w34379_,
		_w34387_,
		_w34388_
	);
	LUT2 #(
		.INIT('h4)
	) name30342 (
		\sport0_rxctl_RXSHT_reg[10]/P0001 ,
		_w20868_,
		_w34389_
	);
	LUT2 #(
		.INIT('h8)
	) name30343 (
		\sport0_rxctl_RX_reg[10]/P0001 ,
		_w20873_,
		_w34390_
	);
	LUT2 #(
		.INIT('h4)
	) name30344 (
		_w20882_,
		_w34358_,
		_w34391_
	);
	LUT2 #(
		.INIT('h8)
	) name30345 (
		\sport0_rxctl_RX_reg[2]/P0001 ,
		_w31045_,
		_w34392_
	);
	LUT2 #(
		.INIT('h1)
	) name30346 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20961_,
		_w34393_
	);
	LUT2 #(
		.INIT('h4)
	) name30347 (
		_w34392_,
		_w34393_,
		_w34394_
	);
	LUT2 #(
		.INIT('h8)
	) name30348 (
		_w20882_,
		_w34394_,
		_w34395_
	);
	LUT2 #(
		.INIT('h1)
	) name30349 (
		_w34391_,
		_w34395_,
		_w34396_
	);
	LUT2 #(
		.INIT('h8)
	) name30350 (
		_w34363_,
		_w34396_,
		_w34397_
	);
	LUT2 #(
		.INIT('h8)
	) name30351 (
		_w34364_,
		_w34365_,
		_w34398_
	);
	LUT2 #(
		.INIT('h1)
	) name30352 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w34398_,
		_w34399_
	);
	LUT2 #(
		.INIT('h4)
	) name30353 (
		_w20882_,
		_w34394_,
		_w34400_
	);
	LUT2 #(
		.INIT('h4)
	) name30354 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w31033_,
		_w34401_
	);
	LUT2 #(
		.INIT('h8)
	) name30355 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w34401_,
		_w34402_
	);
	LUT2 #(
		.INIT('h1)
	) name30356 (
		_w34400_,
		_w34402_,
		_w34403_
	);
	LUT2 #(
		.INIT('h2)
	) name30357 (
		_w34399_,
		_w34403_,
		_w34404_
	);
	LUT2 #(
		.INIT('h4)
	) name30358 (
		_w34399_,
		_w34403_,
		_w34405_
	);
	LUT2 #(
		.INIT('h1)
	) name30359 (
		_w34404_,
		_w34405_,
		_w34406_
	);
	LUT2 #(
		.INIT('h8)
	) name30360 (
		_w34397_,
		_w34406_,
		_w34407_
	);
	LUT2 #(
		.INIT('h1)
	) name30361 (
		_w34397_,
		_w34406_,
		_w34408_
	);
	LUT2 #(
		.INIT('h2)
	) name30362 (
		_w20875_,
		_w34407_,
		_w34409_
	);
	LUT2 #(
		.INIT('h4)
	) name30363 (
		_w34408_,
		_w34409_,
		_w34410_
	);
	LUT2 #(
		.INIT('h4)
	) name30364 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w7859_,
		_w34411_
	);
	LUT2 #(
		.INIT('h1)
	) name30365 (
		_w20868_,
		_w34390_,
		_w34412_
	);
	LUT2 #(
		.INIT('h4)
	) name30366 (
		_w34411_,
		_w34412_,
		_w34413_
	);
	LUT2 #(
		.INIT('h4)
	) name30367 (
		_w34410_,
		_w34413_,
		_w34414_
	);
	LUT2 #(
		.INIT('h1)
	) name30368 (
		_w20871_,
		_w34389_,
		_w34415_
	);
	LUT2 #(
		.INIT('h4)
	) name30369 (
		_w34414_,
		_w34415_,
		_w34416_
	);
	LUT2 #(
		.INIT('h8)
	) name30370 (
		\sport0_rxctl_RX_reg[10]/P0001 ,
		_w20871_,
		_w34417_
	);
	LUT2 #(
		.INIT('h1)
	) name30371 (
		_w34416_,
		_w34417_,
		_w34418_
	);
	LUT2 #(
		.INIT('h1)
	) name30372 (
		\idma_DCTL_reg[0]/NET0131 ,
		\idma_DCTL_reg[10]/NET0131 ,
		_w34419_
	);
	LUT2 #(
		.INIT('h1)
	) name30373 (
		\idma_DCTL_reg[11]/NET0131 ,
		\idma_DCTL_reg[12]/NET0131 ,
		_w34420_
	);
	LUT2 #(
		.INIT('h1)
	) name30374 (
		\idma_DCTL_reg[13]/NET0131 ,
		\idma_DCTL_reg[1]/NET0131 ,
		_w34421_
	);
	LUT2 #(
		.INIT('h1)
	) name30375 (
		\idma_DCTL_reg[2]/NET0131 ,
		\idma_DCTL_reg[3]/NET0131 ,
		_w34422_
	);
	LUT2 #(
		.INIT('h1)
	) name30376 (
		\idma_DCTL_reg[4]/NET0131 ,
		\idma_DCTL_reg[5]/NET0131 ,
		_w34423_
	);
	LUT2 #(
		.INIT('h1)
	) name30377 (
		\idma_DCTL_reg[6]/NET0131 ,
		\idma_DCTL_reg[7]/NET0131 ,
		_w34424_
	);
	LUT2 #(
		.INIT('h1)
	) name30378 (
		\idma_DCTL_reg[8]/NET0131 ,
		\idma_DCTL_reg[9]/NET0131 ,
		_w34425_
	);
	LUT2 #(
		.INIT('h8)
	) name30379 (
		_w34424_,
		_w34425_,
		_w34426_
	);
	LUT2 #(
		.INIT('h8)
	) name30380 (
		_w34422_,
		_w34423_,
		_w34427_
	);
	LUT2 #(
		.INIT('h8)
	) name30381 (
		_w34420_,
		_w34421_,
		_w34428_
	);
	LUT2 #(
		.INIT('h8)
	) name30382 (
		_w20386_,
		_w34419_,
		_w34429_
	);
	LUT2 #(
		.INIT('h8)
	) name30383 (
		_w34428_,
		_w34429_,
		_w34430_
	);
	LUT2 #(
		.INIT('h8)
	) name30384 (
		_w34426_,
		_w34427_,
		_w34431_
	);
	LUT2 #(
		.INIT('h8)
	) name30385 (
		_w34430_,
		_w34431_,
		_w34432_
	);
	LUT2 #(
		.INIT('h8)
	) name30386 (
		_w32464_,
		_w34432_,
		_w34433_
	);
	LUT2 #(
		.INIT('h1)
	) name30387 (
		_w4060_,
		_w34433_,
		_w34434_
	);
	LUT2 #(
		.INIT('h1)
	) name30388 (
		\clkc_OUTcnt_reg[4]/NET0131 ,
		_w19470_,
		_w34435_
	);
	LUT2 #(
		.INIT('h1)
	) name30389 (
		_w19471_,
		_w34435_,
		_w34436_
	);
	LUT2 #(
		.INIT('h4)
	) name30390 (
		_w19467_,
		_w34436_,
		_w34437_
	);
	LUT2 #(
		.INIT('h1)
	) name30391 (
		\clkc_STDcnt_reg[4]/NET0131 ,
		_w31524_,
		_w34438_
	);
	LUT2 #(
		.INIT('h1)
	) name30392 (
		_w31525_,
		_w34438_,
		_w34439_
	);
	LUT2 #(
		.INIT('h4)
	) name30393 (
		_w31521_,
		_w34439_,
		_w34440_
	);
	LUT2 #(
		.INIT('h2)
	) name30394 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w7607_,
		_w34441_
	);
	LUT2 #(
		.INIT('h8)
	) name30395 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001 ,
		_w14704_,
		_w34442_
	);
	LUT2 #(
		.INIT('h8)
	) name30396 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001 ,
		_w14699_,
		_w34443_
	);
	LUT2 #(
		.INIT('h8)
	) name30397 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001 ,
		_w14706_,
		_w34444_
	);
	LUT2 #(
		.INIT('h8)
	) name30398 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001 ,
		_w14711_,
		_w34445_
	);
	LUT2 #(
		.INIT('h8)
	) name30399 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][15]/P0001 ,
		_w14713_,
		_w34446_
	);
	LUT2 #(
		.INIT('h8)
	) name30400 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][15]/P0001 ,
		_w14702_,
		_w34447_
	);
	LUT2 #(
		.INIT('h8)
	) name30401 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][15]/P0001 ,
		_w14708_,
		_w34448_
	);
	LUT2 #(
		.INIT('h1)
	) name30402 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w34442_,
		_w34449_
	);
	LUT2 #(
		.INIT('h1)
	) name30403 (
		_w34443_,
		_w34444_,
		_w34450_
	);
	LUT2 #(
		.INIT('h1)
	) name30404 (
		_w34445_,
		_w34446_,
		_w34451_
	);
	LUT2 #(
		.INIT('h1)
	) name30405 (
		_w34447_,
		_w34448_,
		_w34452_
	);
	LUT2 #(
		.INIT('h8)
	) name30406 (
		_w34451_,
		_w34452_,
		_w34453_
	);
	LUT2 #(
		.INIT('h8)
	) name30407 (
		_w34449_,
		_w34450_,
		_w34454_
	);
	LUT2 #(
		.INIT('h8)
	) name30408 (
		_w34453_,
		_w34454_,
		_w34455_
	);
	LUT2 #(
		.INIT('h1)
	) name30409 (
		_w34441_,
		_w34455_,
		_w34456_
	);
	LUT2 #(
		.INIT('h2)
	) name30410 (
		_w32366_,
		_w34456_,
		_w34457_
	);
	LUT2 #(
		.INIT('h1)
	) name30411 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w32366_,
		_w34458_
	);
	LUT2 #(
		.INIT('h1)
	) name30412 (
		_w32364_,
		_w34457_,
		_w34459_
	);
	LUT2 #(
		.INIT('h4)
	) name30413 (
		_w34458_,
		_w34459_,
		_w34460_
	);
	LUT2 #(
		.INIT('h8)
	) name30414 (
		\core_c_dec_MTTX1_E_reg/P0001 ,
		_w4117_,
		_w34461_
	);
	LUT2 #(
		.INIT('h2)
	) name30415 (
		_w31995_,
		_w31998_,
		_w34462_
	);
	LUT2 #(
		.INIT('h1)
	) name30416 (
		_w4117_,
		_w32007_,
		_w34463_
	);
	LUT2 #(
		.INIT('h4)
	) name30417 (
		_w32003_,
		_w34463_,
		_w34464_
	);
	LUT2 #(
		.INIT('h8)
	) name30418 (
		_w34462_,
		_w34464_,
		_w34465_
	);
	LUT2 #(
		.INIT('h8)
	) name30419 (
		_w32018_,
		_w34465_,
		_w34466_
	);
	LUT2 #(
		.INIT('h1)
	) name30420 (
		_w34461_,
		_w34466_,
		_w34467_
	);
	LUT2 #(
		.INIT('h2)
	) name30421 (
		_w4116_,
		_w34467_,
		_w34468_
	);
	LUT2 #(
		.INIT('h8)
	) name30422 (
		\core_c_dec_MTTX0_E_reg/P0001 ,
		_w4117_,
		_w34469_
	);
	LUT2 #(
		.INIT('h8)
	) name30423 (
		_w32014_,
		_w34464_,
		_w34470_
	);
	LUT2 #(
		.INIT('h8)
	) name30424 (
		_w32018_,
		_w34470_,
		_w34471_
	);
	LUT2 #(
		.INIT('h1)
	) name30425 (
		_w34469_,
		_w34471_,
		_w34472_
	);
	LUT2 #(
		.INIT('h2)
	) name30426 (
		_w4116_,
		_w34472_,
		_w34473_
	);
	LUT2 #(
		.INIT('h8)
	) name30427 (
		\core_c_dec_MTMreg_E_reg[1]/P0001 ,
		_w4117_,
		_w34474_
	);
	LUT2 #(
		.INIT('h2)
	) name30428 (
		_w31992_,
		_w32000_,
		_w34475_
	);
	LUT2 #(
		.INIT('h4)
	) name30429 (
		_w31995_,
		_w34475_,
		_w34476_
	);
	LUT2 #(
		.INIT('h2)
	) name30430 (
		_w31998_,
		_w32007_,
		_w34477_
	);
	LUT2 #(
		.INIT('h4)
	) name30431 (
		_w32001_,
		_w32003_,
		_w34478_
	);
	LUT2 #(
		.INIT('h4)
	) name30432 (
		_w4117_,
		_w34478_,
		_w34479_
	);
	LUT2 #(
		.INIT('h8)
	) name30433 (
		_w34477_,
		_w34479_,
		_w34480_
	);
	LUT2 #(
		.INIT('h8)
	) name30434 (
		_w34476_,
		_w34480_,
		_w34481_
	);
	LUT2 #(
		.INIT('h1)
	) name30435 (
		_w34474_,
		_w34481_,
		_w34482_
	);
	LUT2 #(
		.INIT('h2)
	) name30436 (
		_w4116_,
		_w34482_,
		_w34483_
	);
	LUT2 #(
		.INIT('h1)
	) name30437 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w23265_,
		_w34484_
	);
	LUT2 #(
		.INIT('h2)
	) name30438 (
		\sport1_txctl_Bcnt_reg[4]/NET0131 ,
		_w22674_,
		_w34485_
	);
	LUT2 #(
		.INIT('h1)
	) name30439 (
		_w22675_,
		_w34485_,
		_w34486_
	);
	LUT2 #(
		.INIT('h8)
	) name30440 (
		_w23265_,
		_w34486_,
		_w34487_
	);
	LUT2 #(
		.INIT('h1)
	) name30441 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w34484_,
		_w34488_
	);
	LUT2 #(
		.INIT('h4)
	) name30442 (
		_w34487_,
		_w34488_,
		_w34489_
	);
	LUT2 #(
		.INIT('h1)
	) name30443 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w23277_,
		_w34490_
	);
	LUT2 #(
		.INIT('h2)
	) name30444 (
		\sport0_txctl_Bcnt_reg[4]/NET0131 ,
		_w19957_,
		_w34491_
	);
	LUT2 #(
		.INIT('h1)
	) name30445 (
		_w19958_,
		_w34491_,
		_w34492_
	);
	LUT2 #(
		.INIT('h8)
	) name30446 (
		_w23277_,
		_w34492_,
		_w34493_
	);
	LUT2 #(
		.INIT('h1)
	) name30447 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w34490_,
		_w34494_
	);
	LUT2 #(
		.INIT('h4)
	) name30448 (
		_w34493_,
		_w34494_,
		_w34495_
	);
	LUT2 #(
		.INIT('h4)
	) name30449 (
		_w10289_,
		_w13763_,
		_w34496_
	);
	LUT2 #(
		.INIT('h2)
	) name30450 (
		\bdma_BWCOUNT_reg[9]/NET0131 ,
		_w33293_,
		_w34497_
	);
	LUT2 #(
		.INIT('h1)
	) name30451 (
		_w13763_,
		_w33294_,
		_w34498_
	);
	LUT2 #(
		.INIT('h4)
	) name30452 (
		_w34497_,
		_w34498_,
		_w34499_
	);
	LUT2 #(
		.INIT('h1)
	) name30453 (
		_w34496_,
		_w34499_,
		_w34500_
	);
	LUT2 #(
		.INIT('h4)
	) name30454 (
		_w10638_,
		_w13763_,
		_w34501_
	);
	LUT2 #(
		.INIT('h2)
	) name30455 (
		\bdma_BWCOUNT_reg[8]/NET0131 ,
		_w33292_,
		_w34502_
	);
	LUT2 #(
		.INIT('h1)
	) name30456 (
		_w13763_,
		_w33293_,
		_w34503_
	);
	LUT2 #(
		.INIT('h4)
	) name30457 (
		_w34502_,
		_w34503_,
		_w34504_
	);
	LUT2 #(
		.INIT('h1)
	) name30458 (
		_w34501_,
		_w34504_,
		_w34505_
	);
	LUT2 #(
		.INIT('h2)
	) name30459 (
		\bdma_BWCOUNT_reg[12]/NET0131 ,
		_w33296_,
		_w34506_
	);
	LUT2 #(
		.INIT('h1)
	) name30460 (
		_w13763_,
		_w33297_,
		_w34507_
	);
	LUT2 #(
		.INIT('h4)
	) name30461 (
		_w34506_,
		_w34507_,
		_w34508_
	);
	LUT2 #(
		.INIT('h4)
	) name30462 (
		_w9178_,
		_w13763_,
		_w34509_
	);
	LUT2 #(
		.INIT('h1)
	) name30463 (
		_w34508_,
		_w34509_,
		_w34510_
	);
	LUT2 #(
		.INIT('h2)
	) name30464 (
		\bdma_BWCOUNT_reg[10]/NET0131 ,
		_w33294_,
		_w34511_
	);
	LUT2 #(
		.INIT('h1)
	) name30465 (
		_w13763_,
		_w33295_,
		_w34512_
	);
	LUT2 #(
		.INIT('h4)
	) name30466 (
		_w34511_,
		_w34512_,
		_w34513_
	);
	LUT2 #(
		.INIT('h4)
	) name30467 (
		_w7859_,
		_w13763_,
		_w34514_
	);
	LUT2 #(
		.INIT('h1)
	) name30468 (
		_w34513_,
		_w34514_,
		_w34515_
	);
	LUT2 #(
		.INIT('h1)
	) name30469 (
		\bdma_BIAD_reg[9]/NET0131 ,
		_w34087_,
		_w34516_
	);
	LUT2 #(
		.INIT('h1)
	) name30470 (
		_w34078_,
		_w34088_,
		_w34517_
	);
	LUT2 #(
		.INIT('h4)
	) name30471 (
		_w34516_,
		_w34517_,
		_w34518_
	);
	LUT2 #(
		.INIT('h8)
	) name30472 (
		_w10289_,
		_w34078_,
		_w34519_
	);
	LUT2 #(
		.INIT('h1)
	) name30473 (
		_w34518_,
		_w34519_,
		_w34520_
	);
	LUT2 #(
		.INIT('h1)
	) name30474 (
		\bdma_BIAD_reg[8]/NET0131 ,
		_w34086_,
		_w34521_
	);
	LUT2 #(
		.INIT('h1)
	) name30475 (
		_w34078_,
		_w34087_,
		_w34522_
	);
	LUT2 #(
		.INIT('h4)
	) name30476 (
		_w34521_,
		_w34522_,
		_w34523_
	);
	LUT2 #(
		.INIT('h8)
	) name30477 (
		_w10638_,
		_w34078_,
		_w34524_
	);
	LUT2 #(
		.INIT('h1)
	) name30478 (
		_w34523_,
		_w34524_,
		_w34525_
	);
	LUT2 #(
		.INIT('h2)
	) name30479 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w34092_,
		_w34526_
	);
	LUT2 #(
		.INIT('h4)
	) name30480 (
		\bdma_BIAD_reg[13]/NET0131 ,
		_w34092_,
		_w34527_
	);
	LUT2 #(
		.INIT('h1)
	) name30481 (
		_w34526_,
		_w34527_,
		_w34528_
	);
	LUT2 #(
		.INIT('h1)
	) name30482 (
		_w34078_,
		_w34528_,
		_w34529_
	);
	LUT2 #(
		.INIT('h8)
	) name30483 (
		_w7340_,
		_w34078_,
		_w34530_
	);
	LUT2 #(
		.INIT('h1)
	) name30484 (
		_w34529_,
		_w34530_,
		_w34531_
	);
	LUT2 #(
		.INIT('h1)
	) name30485 (
		\bdma_BIAD_reg[10]/NET0131 ,
		_w34088_,
		_w34532_
	);
	LUT2 #(
		.INIT('h1)
	) name30486 (
		_w34078_,
		_w34089_,
		_w34533_
	);
	LUT2 #(
		.INIT('h4)
	) name30487 (
		_w34532_,
		_w34533_,
		_w34534_
	);
	LUT2 #(
		.INIT('h8)
	) name30488 (
		_w7859_,
		_w34078_,
		_w34535_
	);
	LUT2 #(
		.INIT('h1)
	) name30489 (
		_w34534_,
		_w34535_,
		_w34536_
	);
	LUT2 #(
		.INIT('h1)
	) name30490 (
		\bdma_BEAD_reg[9]/NET0131 ,
		_w33310_,
		_w34537_
	);
	LUT2 #(
		.INIT('h1)
	) name30491 (
		_w20765_,
		_w33311_,
		_w34538_
	);
	LUT2 #(
		.INIT('h4)
	) name30492 (
		_w34537_,
		_w34538_,
		_w34539_
	);
	LUT2 #(
		.INIT('h8)
	) name30493 (
		_w10289_,
		_w20765_,
		_w34540_
	);
	LUT2 #(
		.INIT('h1)
	) name30494 (
		_w34539_,
		_w34540_,
		_w34541_
	);
	LUT2 #(
		.INIT('h1)
	) name30495 (
		\bdma_BEAD_reg[8]/NET0131 ,
		_w33309_,
		_w34542_
	);
	LUT2 #(
		.INIT('h1)
	) name30496 (
		_w20765_,
		_w33310_,
		_w34543_
	);
	LUT2 #(
		.INIT('h4)
	) name30497 (
		_w34542_,
		_w34543_,
		_w34544_
	);
	LUT2 #(
		.INIT('h8)
	) name30498 (
		_w10638_,
		_w20765_,
		_w34545_
	);
	LUT2 #(
		.INIT('h1)
	) name30499 (
		_w34544_,
		_w34545_,
		_w34546_
	);
	LUT2 #(
		.INIT('h1)
	) name30500 (
		\bdma_BEAD_reg[10]/NET0131 ,
		_w33311_,
		_w34547_
	);
	LUT2 #(
		.INIT('h1)
	) name30501 (
		_w20765_,
		_w33312_,
		_w34548_
	);
	LUT2 #(
		.INIT('h4)
	) name30502 (
		_w34547_,
		_w34548_,
		_w34549_
	);
	LUT2 #(
		.INIT('h8)
	) name30503 (
		_w7859_,
		_w20765_,
		_w34550_
	);
	LUT2 #(
		.INIT('h1)
	) name30504 (
		_w34549_,
		_w34550_,
		_w34551_
	);
	LUT2 #(
		.INIT('h2)
	) name30505 (
		\sport1_txctl_TXSHT_reg[3]/P0001 ,
		_w22677_,
		_w34552_
	);
	LUT2 #(
		.INIT('h8)
	) name30506 (
		\sport1_txctl_TX_reg[4]/P0001 ,
		_w22677_,
		_w34553_
	);
	LUT2 #(
		.INIT('h1)
	) name30507 (
		_w34552_,
		_w34553_,
		_w34554_
	);
	LUT2 #(
		.INIT('h8)
	) name30508 (
		\core_c_dec_MFSPT_Ei_reg/NET0131 ,
		_w4117_,
		_w34555_
	);
	LUT2 #(
		.INIT('h4)
	) name30509 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w31264_,
		_w34556_
	);
	LUT2 #(
		.INIT('h4)
	) name30510 (
		_w31269_,
		_w34556_,
		_w34557_
	);
	LUT2 #(
		.INIT('h8)
	) name30511 (
		_w25864_,
		_w34557_,
		_w34558_
	);
	LUT2 #(
		.INIT('h1)
	) name30512 (
		_w34555_,
		_w34558_,
		_w34559_
	);
	LUT2 #(
		.INIT('h2)
	) name30513 (
		\bdma_BWCOUNT_reg[7]/NET0131 ,
		_w33291_,
		_w34560_
	);
	LUT2 #(
		.INIT('h1)
	) name30514 (
		_w13763_,
		_w33292_,
		_w34561_
	);
	LUT2 #(
		.INIT('h4)
	) name30515 (
		_w34560_,
		_w34561_,
		_w34562_
	);
	LUT2 #(
		.INIT('h4)
	) name30516 (
		_w11265_,
		_w13763_,
		_w34563_
	);
	LUT2 #(
		.INIT('h1)
	) name30517 (
		_w34562_,
		_w34563_,
		_w34564_
	);
	LUT2 #(
		.INIT('h4)
	) name30518 (
		_w11525_,
		_w13763_,
		_w34565_
	);
	LUT2 #(
		.INIT('h2)
	) name30519 (
		\bdma_BWCOUNT_reg[6]/NET0131 ,
		_w13769_,
		_w34566_
	);
	LUT2 #(
		.INIT('h1)
	) name30520 (
		_w13763_,
		_w33291_,
		_w34567_
	);
	LUT2 #(
		.INIT('h4)
	) name30521 (
		_w34566_,
		_w34567_,
		_w34568_
	);
	LUT2 #(
		.INIT('h1)
	) name30522 (
		_w34565_,
		_w34568_,
		_w34569_
	);
	LUT2 #(
		.INIT('h2)
	) name30523 (
		\sport0_txctl_TXSHT_reg[3]/P0001 ,
		_w19960_,
		_w34570_
	);
	LUT2 #(
		.INIT('h8)
	) name30524 (
		\sport0_txctl_TX_reg[4]/P0001 ,
		_w19960_,
		_w34571_
	);
	LUT2 #(
		.INIT('h1)
	) name30525 (
		_w34570_,
		_w34571_,
		_w34572_
	);
	LUT2 #(
		.INIT('h4)
	) name30526 (
		\bdma_BWCOUNT_reg[3]/NET0131 ,
		_w13766_,
		_w34573_
	);
	LUT2 #(
		.INIT('h2)
	) name30527 (
		\bdma_BWCOUNT_reg[4]/NET0131 ,
		_w34573_,
		_w34574_
	);
	LUT2 #(
		.INIT('h1)
	) name30528 (
		_w13763_,
		_w13767_,
		_w34575_
	);
	LUT2 #(
		.INIT('h4)
	) name30529 (
		_w34574_,
		_w34575_,
		_w34576_
	);
	LUT2 #(
		.INIT('h4)
	) name30530 (
		_w10069_,
		_w13763_,
		_w34577_
	);
	LUT2 #(
		.INIT('h1)
	) name30531 (
		_w34576_,
		_w34577_,
		_w34578_
	);
	LUT2 #(
		.INIT('h2)
	) name30532 (
		\bdma_BWCOUNT_reg[3]/NET0131 ,
		_w13766_,
		_w34579_
	);
	LUT2 #(
		.INIT('h1)
	) name30533 (
		_w13763_,
		_w34573_,
		_w34580_
	);
	LUT2 #(
		.INIT('h4)
	) name30534 (
		_w34579_,
		_w34580_,
		_w34581_
	);
	LUT2 #(
		.INIT('h4)
	) name30535 (
		_w8113_,
		_w13763_,
		_w34582_
	);
	LUT2 #(
		.INIT('h1)
	) name30536 (
		_w34581_,
		_w34582_,
		_w34583_
	);
	LUT2 #(
		.INIT('h2)
	) name30537 (
		\bdma_BWCOUNT_reg[2]/NET0131 ,
		_w13765_,
		_w34584_
	);
	LUT2 #(
		.INIT('h1)
	) name30538 (
		_w13763_,
		_w13766_,
		_w34585_
	);
	LUT2 #(
		.INIT('h4)
	) name30539 (
		_w34584_,
		_w34585_,
		_w34586_
	);
	LUT2 #(
		.INIT('h4)
	) name30540 (
		_w8715_,
		_w13763_,
		_w34587_
	);
	LUT2 #(
		.INIT('h1)
	) name30541 (
		_w34586_,
		_w34587_,
		_w34588_
	);
	LUT2 #(
		.INIT('h8)
	) name30542 (
		\bdma_BWCOUNT_reg[0]/NET0131 ,
		_w13755_,
		_w34589_
	);
	LUT2 #(
		.INIT('h1)
	) name30543 (
		_w13763_,
		_w13764_,
		_w34590_
	);
	LUT2 #(
		.INIT('h4)
	) name30544 (
		_w34589_,
		_w34590_,
		_w34591_
	);
	LUT2 #(
		.INIT('h4)
	) name30545 (
		_w7607_,
		_w13763_,
		_w34592_
	);
	LUT2 #(
		.INIT('h1)
	) name30546 (
		_w34591_,
		_w34592_,
		_w34593_
	);
	LUT2 #(
		.INIT('h1)
	) name30547 (
		\bdma_BIAD_reg[6]/NET0131 ,
		_w34084_,
		_w34594_
	);
	LUT2 #(
		.INIT('h1)
	) name30548 (
		_w34078_,
		_w34085_,
		_w34595_
	);
	LUT2 #(
		.INIT('h4)
	) name30549 (
		_w34594_,
		_w34595_,
		_w34596_
	);
	LUT2 #(
		.INIT('h8)
	) name30550 (
		_w11525_,
		_w34078_,
		_w34597_
	);
	LUT2 #(
		.INIT('h1)
	) name30551 (
		_w34596_,
		_w34597_,
		_w34598_
	);
	LUT2 #(
		.INIT('h1)
	) name30552 (
		\bdma_BIAD_reg[7]/NET0131 ,
		_w34085_,
		_w34599_
	);
	LUT2 #(
		.INIT('h1)
	) name30553 (
		_w34078_,
		_w34086_,
		_w34600_
	);
	LUT2 #(
		.INIT('h4)
	) name30554 (
		_w34599_,
		_w34600_,
		_w34601_
	);
	LUT2 #(
		.INIT('h8)
	) name30555 (
		_w11265_,
		_w34078_,
		_w34602_
	);
	LUT2 #(
		.INIT('h1)
	) name30556 (
		_w34601_,
		_w34602_,
		_w34603_
	);
	LUT2 #(
		.INIT('h1)
	) name30557 (
		\bdma_BIAD_reg[5]/NET0131 ,
		_w34083_,
		_w34604_
	);
	LUT2 #(
		.INIT('h1)
	) name30558 (
		_w34078_,
		_w34084_,
		_w34605_
	);
	LUT2 #(
		.INIT('h4)
	) name30559 (
		_w34604_,
		_w34605_,
		_w34606_
	);
	LUT2 #(
		.INIT('h8)
	) name30560 (
		_w10911_,
		_w34078_,
		_w34607_
	);
	LUT2 #(
		.INIT('h1)
	) name30561 (
		_w34606_,
		_w34607_,
		_w34608_
	);
	LUT2 #(
		.INIT('h1)
	) name30562 (
		\bdma_BIAD_reg[4]/NET0131 ,
		_w34082_,
		_w34609_
	);
	LUT2 #(
		.INIT('h1)
	) name30563 (
		_w34078_,
		_w34083_,
		_w34610_
	);
	LUT2 #(
		.INIT('h4)
	) name30564 (
		_w34609_,
		_w34610_,
		_w34611_
	);
	LUT2 #(
		.INIT('h8)
	) name30565 (
		_w10069_,
		_w34078_,
		_w34612_
	);
	LUT2 #(
		.INIT('h1)
	) name30566 (
		_w34611_,
		_w34612_,
		_w34613_
	);
	LUT2 #(
		.INIT('h1)
	) name30567 (
		\bdma_BIAD_reg[3]/NET0131 ,
		_w34081_,
		_w34614_
	);
	LUT2 #(
		.INIT('h1)
	) name30568 (
		_w34078_,
		_w34082_,
		_w34615_
	);
	LUT2 #(
		.INIT('h4)
	) name30569 (
		_w34614_,
		_w34615_,
		_w34616_
	);
	LUT2 #(
		.INIT('h8)
	) name30570 (
		_w8113_,
		_w34078_,
		_w34617_
	);
	LUT2 #(
		.INIT('h1)
	) name30571 (
		_w34616_,
		_w34617_,
		_w34618_
	);
	LUT2 #(
		.INIT('h1)
	) name30572 (
		\bdma_BIAD_reg[2]/NET0131 ,
		_w34080_,
		_w34619_
	);
	LUT2 #(
		.INIT('h1)
	) name30573 (
		_w34078_,
		_w34081_,
		_w34620_
	);
	LUT2 #(
		.INIT('h4)
	) name30574 (
		_w34619_,
		_w34620_,
		_w34621_
	);
	LUT2 #(
		.INIT('h8)
	) name30575 (
		_w8715_,
		_w34078_,
		_w34622_
	);
	LUT2 #(
		.INIT('h1)
	) name30576 (
		_w34621_,
		_w34622_,
		_w34623_
	);
	LUT2 #(
		.INIT('h1)
	) name30577 (
		\bdma_BIAD_reg[1]/NET0131 ,
		_w34079_,
		_w34624_
	);
	LUT2 #(
		.INIT('h1)
	) name30578 (
		_w34078_,
		_w34080_,
		_w34625_
	);
	LUT2 #(
		.INIT('h4)
	) name30579 (
		_w34624_,
		_w34625_,
		_w34626_
	);
	LUT2 #(
		.INIT('h8)
	) name30580 (
		_w9435_,
		_w34078_,
		_w34627_
	);
	LUT2 #(
		.INIT('h1)
	) name30581 (
		_w34626_,
		_w34627_,
		_w34628_
	);
	LUT2 #(
		.INIT('h4)
	) name30582 (
		\bdma_BIAD_reg[0]/NET0131 ,
		_w13755_,
		_w34629_
	);
	LUT2 #(
		.INIT('h1)
	) name30583 (
		_w34078_,
		_w34079_,
		_w34630_
	);
	LUT2 #(
		.INIT('h4)
	) name30584 (
		_w34629_,
		_w34630_,
		_w34631_
	);
	LUT2 #(
		.INIT('h8)
	) name30585 (
		_w7607_,
		_w34078_,
		_w34632_
	);
	LUT2 #(
		.INIT('h1)
	) name30586 (
		_w34631_,
		_w34632_,
		_w34633_
	);
	LUT2 #(
		.INIT('h8)
	) name30587 (
		_w18868_,
		_w32038_,
		_w34634_
	);
	LUT2 #(
		.INIT('h1)
	) name30588 (
		\sice_IIRC_reg[5]/NET0131 ,
		_w34634_,
		_w34635_
	);
	LUT2 #(
		.INIT('h8)
	) name30589 (
		_w18869_,
		_w32038_,
		_w34636_
	);
	LUT2 #(
		.INIT('h1)
	) name30590 (
		_w34635_,
		_w34636_,
		_w34637_
	);
	LUT2 #(
		.INIT('h2)
	) name30591 (
		\sice_IIRC_reg[0]/NET0131 ,
		_w32038_,
		_w34638_
	);
	LUT2 #(
		.INIT('h4)
	) name30592 (
		\sice_IIRC_reg[0]/NET0131 ,
		_w32038_,
		_w34639_
	);
	LUT2 #(
		.INIT('h1)
	) name30593 (
		_w34638_,
		_w34639_,
		_w34640_
	);
	LUT2 #(
		.INIT('h1)
	) name30594 (
		\sice_IIRC_reg[18]/NET0131 ,
		_w32039_,
		_w34641_
	);
	LUT2 #(
		.INIT('h1)
	) name30595 (
		_w32040_,
		_w34641_,
		_w34642_
	);
	LUT2 #(
		.INIT('h1)
	) name30596 (
		\sice_IIRC_reg[19]/NET0131 ,
		_w32040_,
		_w34643_
	);
	LUT2 #(
		.INIT('h1)
	) name30597 (
		_w32041_,
		_w34643_,
		_w34644_
	);
	LUT2 #(
		.INIT('h1)
	) name30598 (
		\sice_IIRC_reg[21]/NET0131 ,
		_w32042_,
		_w34645_
	);
	LUT2 #(
		.INIT('h1)
	) name30599 (
		_w34165_,
		_w34645_,
		_w34646_
	);
	LUT2 #(
		.INIT('h1)
	) name30600 (
		\sice_IIRC_reg[22]/NET0131 ,
		_w34165_,
		_w34647_
	);
	LUT2 #(
		.INIT('h1)
	) name30601 (
		_w34166_,
		_w34647_,
		_w34648_
	);
	LUT2 #(
		.INIT('h1)
	) name30602 (
		\clkc_oscntr_reg_DO_reg[7]/NET0131 ,
		_w23420_,
		_w34649_
	);
	LUT2 #(
		.INIT('h1)
	) name30603 (
		_w23421_,
		_w34649_,
		_w34650_
	);
	LUT2 #(
		.INIT('h2)
	) name30604 (
		_w7340_,
		_w32992_,
		_w34651_
	);
	LUT2 #(
		.INIT('h8)
	) name30605 (
		\core_dag_ilm2reg_L5_we_DO_reg[13]/NET0131 ,
		_w33000_,
		_w34652_
	);
	LUT2 #(
		.INIT('h8)
	) name30606 (
		\core_dag_ilm2reg_L6_we_DO_reg[13]/NET0131 ,
		_w32994_,
		_w34653_
	);
	LUT2 #(
		.INIT('h8)
	) name30607 (
		\core_dag_ilm2reg_L4_we_DO_reg[13]/NET0131 ,
		_w32996_,
		_w34654_
	);
	LUT2 #(
		.INIT('h8)
	) name30608 (
		\core_dag_ilm2reg_L7_we_DO_reg[13]/NET0131 ,
		_w32998_,
		_w34655_
	);
	LUT2 #(
		.INIT('h1)
	) name30609 (
		_w21579_,
		_w34652_,
		_w34656_
	);
	LUT2 #(
		.INIT('h1)
	) name30610 (
		_w34653_,
		_w34654_,
		_w34657_
	);
	LUT2 #(
		.INIT('h4)
	) name30611 (
		_w34655_,
		_w34657_,
		_w34658_
	);
	LUT2 #(
		.INIT('h8)
	) name30612 (
		_w34656_,
		_w34658_,
		_w34659_
	);
	LUT2 #(
		.INIT('h4)
	) name30613 (
		_w34651_,
		_w34659_,
		_w34660_
	);
	LUT2 #(
		.INIT('h4)
	) name30614 (
		\core_dag_ilm2reg_L_reg[13]/NET0131 ,
		_w21579_,
		_w34661_
	);
	LUT2 #(
		.INIT('h1)
	) name30615 (
		_w34660_,
		_w34661_,
		_w34662_
	);
	LUT2 #(
		.INIT('h2)
	) name30616 (
		_w7859_,
		_w32992_,
		_w34663_
	);
	LUT2 #(
		.INIT('h8)
	) name30617 (
		\core_dag_ilm2reg_L5_we_DO_reg[10]/NET0131 ,
		_w33000_,
		_w34664_
	);
	LUT2 #(
		.INIT('h8)
	) name30618 (
		\core_dag_ilm2reg_L6_we_DO_reg[10]/NET0131 ,
		_w32994_,
		_w34665_
	);
	LUT2 #(
		.INIT('h8)
	) name30619 (
		\core_dag_ilm2reg_L4_we_DO_reg[10]/NET0131 ,
		_w32996_,
		_w34666_
	);
	LUT2 #(
		.INIT('h8)
	) name30620 (
		\core_dag_ilm2reg_L7_we_DO_reg[10]/NET0131 ,
		_w32998_,
		_w34667_
	);
	LUT2 #(
		.INIT('h1)
	) name30621 (
		_w21579_,
		_w34664_,
		_w34668_
	);
	LUT2 #(
		.INIT('h1)
	) name30622 (
		_w34665_,
		_w34666_,
		_w34669_
	);
	LUT2 #(
		.INIT('h4)
	) name30623 (
		_w34667_,
		_w34669_,
		_w34670_
	);
	LUT2 #(
		.INIT('h8)
	) name30624 (
		_w34668_,
		_w34670_,
		_w34671_
	);
	LUT2 #(
		.INIT('h4)
	) name30625 (
		_w34663_,
		_w34671_,
		_w34672_
	);
	LUT2 #(
		.INIT('h4)
	) name30626 (
		\core_dag_ilm2reg_L_reg[10]/NET0131 ,
		_w21579_,
		_w34673_
	);
	LUT2 #(
		.INIT('h1)
	) name30627 (
		_w34672_,
		_w34673_,
		_w34674_
	);
	LUT2 #(
		.INIT('h8)
	) name30628 (
		\core_dag_ilm2reg_I6_we_DO_reg[8]/NET0131 ,
		_w33684_,
		_w34675_
	);
	LUT2 #(
		.INIT('h8)
	) name30629 (
		\core_dag_ilm2reg_I7_we_DO_reg[8]/NET0131 ,
		_w33686_,
		_w34676_
	);
	LUT2 #(
		.INIT('h8)
	) name30630 (
		\core_dag_ilm2reg_I4_we_DO_reg[8]/NET0131 ,
		_w33690_,
		_w34677_
	);
	LUT2 #(
		.INIT('h8)
	) name30631 (
		\core_dag_ilm2reg_I5_we_DO_reg[8]/NET0131 ,
		_w33688_,
		_w34678_
	);
	LUT2 #(
		.INIT('h2)
	) name30632 (
		_w20602_,
		_w33698_,
		_w34679_
	);
	LUT2 #(
		.INIT('h1)
	) name30633 (
		_w21579_,
		_w34675_,
		_w34680_
	);
	LUT2 #(
		.INIT('h1)
	) name30634 (
		_w34676_,
		_w34677_,
		_w34681_
	);
	LUT2 #(
		.INIT('h4)
	) name30635 (
		_w34678_,
		_w34681_,
		_w34682_
	);
	LUT2 #(
		.INIT('h8)
	) name30636 (
		_w34680_,
		_w34682_,
		_w34683_
	);
	LUT2 #(
		.INIT('h4)
	) name30637 (
		_w34679_,
		_w34683_,
		_w34684_
	);
	LUT2 #(
		.INIT('h4)
	) name30638 (
		\core_dag_ilm2reg_I_reg[8]/NET0131 ,
		_w21579_,
		_w34685_
	);
	LUT2 #(
		.INIT('h1)
	) name30639 (
		_w34684_,
		_w34685_,
		_w34686_
	);
	LUT2 #(
		.INIT('h8)
	) name30640 (
		\core_dag_ilm2reg_I6_we_DO_reg[11]/NET0131 ,
		_w33684_,
		_w34687_
	);
	LUT2 #(
		.INIT('h8)
	) name30641 (
		\core_dag_ilm2reg_I7_we_DO_reg[11]/NET0131 ,
		_w33686_,
		_w34688_
	);
	LUT2 #(
		.INIT('h8)
	) name30642 (
		\core_dag_ilm2reg_I4_we_DO_reg[11]/NET0131 ,
		_w33690_,
		_w34689_
	);
	LUT2 #(
		.INIT('h8)
	) name30643 (
		\core_dag_ilm2reg_I5_we_DO_reg[11]/NET0131 ,
		_w33688_,
		_w34690_
	);
	LUT2 #(
		.INIT('h1)
	) name30644 (
		_w20707_,
		_w33698_,
		_w34691_
	);
	LUT2 #(
		.INIT('h1)
	) name30645 (
		_w21579_,
		_w34687_,
		_w34692_
	);
	LUT2 #(
		.INIT('h1)
	) name30646 (
		_w34688_,
		_w34689_,
		_w34693_
	);
	LUT2 #(
		.INIT('h4)
	) name30647 (
		_w34690_,
		_w34693_,
		_w34694_
	);
	LUT2 #(
		.INIT('h8)
	) name30648 (
		_w34692_,
		_w34694_,
		_w34695_
	);
	LUT2 #(
		.INIT('h4)
	) name30649 (
		_w34691_,
		_w34695_,
		_w34696_
	);
	LUT2 #(
		.INIT('h4)
	) name30650 (
		\core_dag_ilm2reg_I_reg[11]/NET0131 ,
		_w21579_,
		_w34697_
	);
	LUT2 #(
		.INIT('h1)
	) name30651 (
		_w34696_,
		_w34697_,
		_w34698_
	);
	LUT2 #(
		.INIT('h8)
	) name30652 (
		\core_dag_ilm2reg_I6_we_DO_reg[10]/NET0131 ,
		_w33684_,
		_w34699_
	);
	LUT2 #(
		.INIT('h8)
	) name30653 (
		\core_dag_ilm2reg_I7_we_DO_reg[10]/NET0131 ,
		_w33686_,
		_w34700_
	);
	LUT2 #(
		.INIT('h8)
	) name30654 (
		\core_dag_ilm2reg_I4_we_DO_reg[10]/NET0131 ,
		_w33690_,
		_w34701_
	);
	LUT2 #(
		.INIT('h8)
	) name30655 (
		\core_dag_ilm2reg_I5_we_DO_reg[10]/NET0131 ,
		_w33688_,
		_w34702_
	);
	LUT2 #(
		.INIT('h2)
	) name30656 (
		_w20718_,
		_w33698_,
		_w34703_
	);
	LUT2 #(
		.INIT('h1)
	) name30657 (
		_w21579_,
		_w34699_,
		_w34704_
	);
	LUT2 #(
		.INIT('h1)
	) name30658 (
		_w34700_,
		_w34701_,
		_w34705_
	);
	LUT2 #(
		.INIT('h4)
	) name30659 (
		_w34702_,
		_w34705_,
		_w34706_
	);
	LUT2 #(
		.INIT('h8)
	) name30660 (
		_w34704_,
		_w34706_,
		_w34707_
	);
	LUT2 #(
		.INIT('h4)
	) name30661 (
		_w34703_,
		_w34707_,
		_w34708_
	);
	LUT2 #(
		.INIT('h4)
	) name30662 (
		\core_dag_ilm2reg_I_reg[10]/NET0131 ,
		_w21579_,
		_w34709_
	);
	LUT2 #(
		.INIT('h1)
	) name30663 (
		_w34708_,
		_w34709_,
		_w34710_
	);
	LUT2 #(
		.INIT('h8)
	) name30664 (
		\core_dag_ilm1reg_I2_we_DO_reg[9]/NET0131 ,
		_w33910_,
		_w34711_
	);
	LUT2 #(
		.INIT('h8)
	) name30665 (
		\core_dag_ilm1reg_I1_we_DO_reg[9]/NET0131 ,
		_w33937_,
		_w34712_
	);
	LUT2 #(
		.INIT('h8)
	) name30666 (
		\core_dag_ilm1reg_I0_we_DO_reg[9]/NET0131 ,
		_w33922_,
		_w34713_
	);
	LUT2 #(
		.INIT('h8)
	) name30667 (
		\core_dag_ilm1reg_I3_we_DO_reg[9]/NET0131 ,
		_w33908_,
		_w34714_
	);
	LUT2 #(
		.INIT('h1)
	) name30668 (
		_w24098_,
		_w33896_,
		_w34715_
	);
	LUT2 #(
		.INIT('h1)
	) name30669 (
		_w21592_,
		_w34711_,
		_w34716_
	);
	LUT2 #(
		.INIT('h1)
	) name30670 (
		_w34712_,
		_w34713_,
		_w34717_
	);
	LUT2 #(
		.INIT('h4)
	) name30671 (
		_w34714_,
		_w34717_,
		_w34718_
	);
	LUT2 #(
		.INIT('h8)
	) name30672 (
		_w34716_,
		_w34718_,
		_w34719_
	);
	LUT2 #(
		.INIT('h4)
	) name30673 (
		_w34715_,
		_w34719_,
		_w34720_
	);
	LUT2 #(
		.INIT('h4)
	) name30674 (
		\core_dag_ilm1reg_I_reg[9]/NET0131 ,
		_w21592_,
		_w34721_
	);
	LUT2 #(
		.INIT('h1)
	) name30675 (
		_w34720_,
		_w34721_,
		_w34722_
	);
	LUT2 #(
		.INIT('h2)
	) name30676 (
		_w10911_,
		_w32992_,
		_w34723_
	);
	LUT2 #(
		.INIT('h8)
	) name30677 (
		\core_dag_ilm2reg_L7_we_DO_reg[5]/NET0131 ,
		_w32998_,
		_w34724_
	);
	LUT2 #(
		.INIT('h8)
	) name30678 (
		\core_dag_ilm2reg_L4_we_DO_reg[5]/NET0131 ,
		_w32996_,
		_w34725_
	);
	LUT2 #(
		.INIT('h8)
	) name30679 (
		\core_dag_ilm2reg_L6_we_DO_reg[5]/NET0131 ,
		_w32994_,
		_w34726_
	);
	LUT2 #(
		.INIT('h8)
	) name30680 (
		\core_dag_ilm2reg_L5_we_DO_reg[5]/NET0131 ,
		_w33000_,
		_w34727_
	);
	LUT2 #(
		.INIT('h1)
	) name30681 (
		_w21579_,
		_w34724_,
		_w34728_
	);
	LUT2 #(
		.INIT('h1)
	) name30682 (
		_w34725_,
		_w34726_,
		_w34729_
	);
	LUT2 #(
		.INIT('h4)
	) name30683 (
		_w34727_,
		_w34729_,
		_w34730_
	);
	LUT2 #(
		.INIT('h8)
	) name30684 (
		_w34728_,
		_w34730_,
		_w34731_
	);
	LUT2 #(
		.INIT('h4)
	) name30685 (
		_w34723_,
		_w34731_,
		_w34732_
	);
	LUT2 #(
		.INIT('h4)
	) name30686 (
		\core_dag_ilm2reg_L_reg[5]/NET0131 ,
		_w21579_,
		_w34733_
	);
	LUT2 #(
		.INIT('h1)
	) name30687 (
		_w34732_,
		_w34733_,
		_w34734_
	);
	LUT2 #(
		.INIT('h8)
	) name30688 (
		\core_dag_ilm2reg_I6_we_DO_reg[7]/NET0131 ,
		_w33684_,
		_w34735_
	);
	LUT2 #(
		.INIT('h8)
	) name30689 (
		\core_dag_ilm2reg_I5_we_DO_reg[7]/NET0131 ,
		_w33688_,
		_w34736_
	);
	LUT2 #(
		.INIT('h8)
	) name30690 (
		\core_dag_ilm2reg_I7_we_DO_reg[7]/NET0131 ,
		_w33686_,
		_w34737_
	);
	LUT2 #(
		.INIT('h8)
	) name30691 (
		\core_dag_ilm2reg_I4_we_DO_reg[7]/NET0131 ,
		_w33690_,
		_w34738_
	);
	LUT2 #(
		.INIT('h2)
	) name30692 (
		_w20614_,
		_w33698_,
		_w34739_
	);
	LUT2 #(
		.INIT('h1)
	) name30693 (
		_w21579_,
		_w34735_,
		_w34740_
	);
	LUT2 #(
		.INIT('h1)
	) name30694 (
		_w34736_,
		_w34737_,
		_w34741_
	);
	LUT2 #(
		.INIT('h4)
	) name30695 (
		_w34738_,
		_w34741_,
		_w34742_
	);
	LUT2 #(
		.INIT('h8)
	) name30696 (
		_w34740_,
		_w34742_,
		_w34743_
	);
	LUT2 #(
		.INIT('h4)
	) name30697 (
		_w34739_,
		_w34743_,
		_w34744_
	);
	LUT2 #(
		.INIT('h4)
	) name30698 (
		\core_dag_ilm2reg_I_reg[7]/NET0131 ,
		_w21579_,
		_w34745_
	);
	LUT2 #(
		.INIT('h1)
	) name30699 (
		_w34744_,
		_w34745_,
		_w34746_
	);
	LUT2 #(
		.INIT('h8)
	) name30700 (
		_w24170_,
		_w33091_,
		_w34747_
	);
	LUT2 #(
		.INIT('h8)
	) name30701 (
		\core_dag_ilm1reg_I3_we_DO_reg[7]/NET0131 ,
		_w33908_,
		_w34748_
	);
	LUT2 #(
		.INIT('h8)
	) name30702 (
		\core_dag_ilm1reg_I2_we_DO_reg[7]/NET0131 ,
		_w33910_,
		_w34749_
	);
	LUT2 #(
		.INIT('h8)
	) name30703 (
		\core_dag_ilm1reg_I1_we_DO_reg[7]/NET0131 ,
		_w33937_,
		_w34750_
	);
	LUT2 #(
		.INIT('h1)
	) name30704 (
		_w24106_,
		_w33896_,
		_w34751_
	);
	LUT2 #(
		.INIT('h1)
	) name30705 (
		_w21592_,
		_w34747_,
		_w34752_
	);
	LUT2 #(
		.INIT('h1)
	) name30706 (
		_w34748_,
		_w34749_,
		_w34753_
	);
	LUT2 #(
		.INIT('h4)
	) name30707 (
		_w34750_,
		_w34753_,
		_w34754_
	);
	LUT2 #(
		.INIT('h8)
	) name30708 (
		_w34752_,
		_w34754_,
		_w34755_
	);
	LUT2 #(
		.INIT('h4)
	) name30709 (
		_w34751_,
		_w34755_,
		_w34756_
	);
	LUT2 #(
		.INIT('h4)
	) name30710 (
		\core_dag_ilm1reg_I_reg[7]/NET0131 ,
		_w21592_,
		_w34757_
	);
	LUT2 #(
		.INIT('h1)
	) name30711 (
		_w34756_,
		_w34757_,
		_w34758_
	);
	LUT2 #(
		.INIT('h8)
	) name30712 (
		_w24173_,
		_w33091_,
		_w34759_
	);
	LUT2 #(
		.INIT('h8)
	) name30713 (
		\core_dag_ilm1reg_I3_we_DO_reg[6]/NET0131 ,
		_w33908_,
		_w34760_
	);
	LUT2 #(
		.INIT('h8)
	) name30714 (
		\core_dag_ilm1reg_I2_we_DO_reg[6]/NET0131 ,
		_w33910_,
		_w34761_
	);
	LUT2 #(
		.INIT('h8)
	) name30715 (
		\core_dag_ilm1reg_I1_we_DO_reg[6]/NET0131 ,
		_w33937_,
		_w34762_
	);
	LUT2 #(
		.INIT('h1)
	) name30716 (
		_w24111_,
		_w33896_,
		_w34763_
	);
	LUT2 #(
		.INIT('h1)
	) name30717 (
		_w21592_,
		_w34759_,
		_w34764_
	);
	LUT2 #(
		.INIT('h1)
	) name30718 (
		_w34760_,
		_w34761_,
		_w34765_
	);
	LUT2 #(
		.INIT('h4)
	) name30719 (
		_w34762_,
		_w34765_,
		_w34766_
	);
	LUT2 #(
		.INIT('h8)
	) name30720 (
		_w34764_,
		_w34766_,
		_w34767_
	);
	LUT2 #(
		.INIT('h4)
	) name30721 (
		_w34763_,
		_w34767_,
		_w34768_
	);
	LUT2 #(
		.INIT('h4)
	) name30722 (
		\core_dag_ilm1reg_I_reg[6]/NET0131 ,
		_w21592_,
		_w34769_
	);
	LUT2 #(
		.INIT('h1)
	) name30723 (
		_w34768_,
		_w34769_,
		_w34770_
	);
	LUT2 #(
		.INIT('h8)
	) name30724 (
		\core_dag_ilm1reg_I2_we_DO_reg[4]/NET0131 ,
		_w33910_,
		_w34771_
	);
	LUT2 #(
		.INIT('h8)
	) name30725 (
		\core_dag_ilm1reg_I1_we_DO_reg[4]/NET0131 ,
		_w33937_,
		_w34772_
	);
	LUT2 #(
		.INIT('h8)
	) name30726 (
		\core_dag_ilm1reg_I0_we_DO_reg[4]/NET0131 ,
		_w33922_,
		_w34773_
	);
	LUT2 #(
		.INIT('h8)
	) name30727 (
		\core_dag_ilm1reg_I3_we_DO_reg[4]/NET0131 ,
		_w33908_,
		_w34774_
	);
	LUT2 #(
		.INIT('h1)
	) name30728 (
		_w24118_,
		_w33896_,
		_w34775_
	);
	LUT2 #(
		.INIT('h1)
	) name30729 (
		_w21592_,
		_w34771_,
		_w34776_
	);
	LUT2 #(
		.INIT('h1)
	) name30730 (
		_w34772_,
		_w34773_,
		_w34777_
	);
	LUT2 #(
		.INIT('h4)
	) name30731 (
		_w34774_,
		_w34777_,
		_w34778_
	);
	LUT2 #(
		.INIT('h8)
	) name30732 (
		_w34776_,
		_w34778_,
		_w34779_
	);
	LUT2 #(
		.INIT('h4)
	) name30733 (
		_w34775_,
		_w34779_,
		_w34780_
	);
	LUT2 #(
		.INIT('h4)
	) name30734 (
		\core_dag_ilm1reg_I_reg[4]/NET0131 ,
		_w21592_,
		_w34781_
	);
	LUT2 #(
		.INIT('h1)
	) name30735 (
		_w34780_,
		_w34781_,
		_w34782_
	);
	LUT2 #(
		.INIT('h8)
	) name30736 (
		\core_dag_ilm1reg_I2_we_DO_reg[3]/NET0131 ,
		_w33910_,
		_w34783_
	);
	LUT2 #(
		.INIT('h8)
	) name30737 (
		\core_dag_ilm1reg_I1_we_DO_reg[3]/NET0131 ,
		_w33937_,
		_w34784_
	);
	LUT2 #(
		.INIT('h8)
	) name30738 (
		\core_dag_ilm1reg_I3_we_DO_reg[3]/NET0131 ,
		_w33908_,
		_w34785_
	);
	LUT2 #(
		.INIT('h2)
	) name30739 (
		_w23886_,
		_w33896_,
		_w34786_
	);
	LUT2 #(
		.INIT('h8)
	) name30740 (
		\core_dag_ilm1reg_I0_we_DO_reg[3]/NET0131 ,
		_w33922_,
		_w34787_
	);
	LUT2 #(
		.INIT('h1)
	) name30741 (
		_w21592_,
		_w34783_,
		_w34788_
	);
	LUT2 #(
		.INIT('h1)
	) name30742 (
		_w34784_,
		_w34785_,
		_w34789_
	);
	LUT2 #(
		.INIT('h4)
	) name30743 (
		_w34787_,
		_w34789_,
		_w34790_
	);
	LUT2 #(
		.INIT('h8)
	) name30744 (
		_w34788_,
		_w34790_,
		_w34791_
	);
	LUT2 #(
		.INIT('h4)
	) name30745 (
		_w34786_,
		_w34791_,
		_w34792_
	);
	LUT2 #(
		.INIT('h4)
	) name30746 (
		\core_dag_ilm1reg_I_reg[3]/NET0131 ,
		_w21592_,
		_w34793_
	);
	LUT2 #(
		.INIT('h1)
	) name30747 (
		_w34792_,
		_w34793_,
		_w34794_
	);
	LUT2 #(
		.INIT('h8)
	) name30748 (
		\core_dag_ilm1reg_I0_we_DO_reg[2]/NET0131 ,
		_w33922_,
		_w34795_
	);
	LUT2 #(
		.INIT('h8)
	) name30749 (
		\core_dag_ilm1reg_I1_we_DO_reg[2]/NET0131 ,
		_w33937_,
		_w34796_
	);
	LUT2 #(
		.INIT('h8)
	) name30750 (
		\core_dag_ilm1reg_I2_we_DO_reg[2]/NET0131 ,
		_w33910_,
		_w34797_
	);
	LUT2 #(
		.INIT('h8)
	) name30751 (
		\core_dag_ilm1reg_I3_we_DO_reg[2]/NET0131 ,
		_w33908_,
		_w34798_
	);
	LUT2 #(
		.INIT('h1)
	) name30752 (
		_w24124_,
		_w33896_,
		_w34799_
	);
	LUT2 #(
		.INIT('h1)
	) name30753 (
		_w21592_,
		_w34795_,
		_w34800_
	);
	LUT2 #(
		.INIT('h1)
	) name30754 (
		_w34796_,
		_w34797_,
		_w34801_
	);
	LUT2 #(
		.INIT('h4)
	) name30755 (
		_w34798_,
		_w34801_,
		_w34802_
	);
	LUT2 #(
		.INIT('h8)
	) name30756 (
		_w34800_,
		_w34802_,
		_w34803_
	);
	LUT2 #(
		.INIT('h4)
	) name30757 (
		_w34799_,
		_w34803_,
		_w34804_
	);
	LUT2 #(
		.INIT('h4)
	) name30758 (
		\core_dag_ilm1reg_I_reg[2]/NET0131 ,
		_w21592_,
		_w34805_
	);
	LUT2 #(
		.INIT('h1)
	) name30759 (
		_w34804_,
		_w34805_,
		_w34806_
	);
	LUT2 #(
		.INIT('h8)
	) name30760 (
		\core_dag_ilm1reg_I2_we_DO_reg[0]/NET0131 ,
		_w33910_,
		_w34807_
	);
	LUT2 #(
		.INIT('h8)
	) name30761 (
		\core_dag_ilm1reg_I3_we_DO_reg[0]/NET0131 ,
		_w33908_,
		_w34808_
	);
	LUT2 #(
		.INIT('h8)
	) name30762 (
		\core_dag_ilm1reg_I0_we_DO_reg[0]/NET0131 ,
		_w33922_,
		_w34809_
	);
	LUT2 #(
		.INIT('h8)
	) name30763 (
		\core_dag_ilm1reg_I1_we_DO_reg[0]/NET0131 ,
		_w33937_,
		_w34810_
	);
	LUT2 #(
		.INIT('h1)
	) name30764 (
		_w24143_,
		_w33896_,
		_w34811_
	);
	LUT2 #(
		.INIT('h1)
	) name30765 (
		_w21592_,
		_w34807_,
		_w34812_
	);
	LUT2 #(
		.INIT('h1)
	) name30766 (
		_w34808_,
		_w34809_,
		_w34813_
	);
	LUT2 #(
		.INIT('h4)
	) name30767 (
		_w34810_,
		_w34813_,
		_w34814_
	);
	LUT2 #(
		.INIT('h8)
	) name30768 (
		_w34812_,
		_w34814_,
		_w34815_
	);
	LUT2 #(
		.INIT('h4)
	) name30769 (
		_w34811_,
		_w34815_,
		_w34816_
	);
	LUT2 #(
		.INIT('h4)
	) name30770 (
		\core_dag_ilm1reg_I_reg[0]/NET0131 ,
		_w21592_,
		_w34817_
	);
	LUT2 #(
		.INIT('h1)
	) name30771 (
		_w34816_,
		_w34817_,
		_w34818_
	);
	LUT2 #(
		.INIT('h1)
	) name30772 (
		_w5950_,
		_w27908_,
		_w34819_
	);
	LUT2 #(
		.INIT('h8)
	) name30773 (
		\core_c_psq_cntstk_ptr_reg[2]/NET0131 ,
		_w33341_,
		_w34820_
	);
	LUT2 #(
		.INIT('h2)
	) name30774 (
		\core_c_psq_CNTRval_reg/NET0131 ,
		_w34820_,
		_w34821_
	);
	LUT2 #(
		.INIT('h1)
	) name30775 (
		_w34819_,
		_w34821_,
		_w34822_
	);
	LUT2 #(
		.INIT('h1)
	) name30776 (
		\sice_IIRC_reg[8]/NET0131 ,
		_w18871_,
		_w34823_
	);
	LUT2 #(
		.INIT('h1)
	) name30777 (
		_w20853_,
		_w34823_,
		_w34824_
	);
	LUT2 #(
		.INIT('h8)
	) name30778 (
		\sice_ICS_reg[2]/NET0131 ,
		_w26064_,
		_w34825_
	);
	LUT2 #(
		.INIT('h8)
	) name30779 (
		\sice_SPC_reg[20]/P0001 ,
		_w34825_,
		_w34826_
	);
	LUT2 #(
		.INIT('h4)
	) name30780 (
		_w26336_,
		_w28982_,
		_w34827_
	);
	LUT2 #(
		.INIT('h2)
	) name30781 (
		\sice_SPC_reg[22]/P0001 ,
		_w34825_,
		_w34828_
	);
	LUT2 #(
		.INIT('h1)
	) name30782 (
		_w34826_,
		_w34828_,
		_w34829_
	);
	LUT2 #(
		.INIT('h4)
	) name30783 (
		_w34827_,
		_w34829_,
		_w34830_
	);
	LUT2 #(
		.INIT('h8)
	) name30784 (
		_w23028_,
		_w25053_,
		_w34831_
	);
	LUT2 #(
		.INIT('h8)
	) name30785 (
		\sice_IBR1_reg[15]/P0001 ,
		_w34831_,
		_w34832_
	);
	LUT2 #(
		.INIT('h8)
	) name30786 (
		\sice_IMR2_reg[15]/NET0131 ,
		_w25034_,
		_w34833_
	);
	LUT2 #(
		.INIT('h8)
	) name30787 (
		\sice_DBR1_reg[16]/P0001 ,
		_w25054_,
		_w34834_
	);
	LUT2 #(
		.INIT('h8)
	) name30788 (
		\sice_IIRC_reg[21]/NET0131 ,
		_w24267_,
		_w34835_
	);
	LUT2 #(
		.INIT('h8)
	) name30789 (
		\sice_DMR2_reg[15]/NET0131 ,
		_w25025_,
		_w34836_
	);
	LUT2 #(
		.INIT('h8)
	) name30790 (
		\sice_CLR_I_reg/NET0131 ,
		_w23029_,
		_w34837_
	);
	LUT2 #(
		.INIT('h8)
	) name30791 (
		\sice_idr1_reg_DO_reg[9]/P0001 ,
		_w26968_,
		_w34838_
	);
	LUT2 #(
		.INIT('h8)
	) name30792 (
		\sice_DMR1_reg[15]/NET0131 ,
		_w27903_,
		_w34839_
	);
	LUT2 #(
		.INIT('h8)
	) name30793 (
		\sice_ICYC_reg[21]/NET0131 ,
		_w23409_,
		_w34840_
	);
	LUT2 #(
		.INIT('h8)
	) name30794 (
		_w23027_,
		_w25010_,
		_w34841_
	);
	LUT2 #(
		.INIT('h8)
	) name30795 (
		\sice_IRR_reg[11]/P0001 ,
		_w34841_,
		_w34842_
	);
	LUT2 #(
		.INIT('h8)
	) name30796 (
		\sice_DBR2_reg[16]/P0001 ,
		_w25012_,
		_w34843_
	);
	LUT2 #(
		.INIT('h8)
	) name30797 (
		\core_c_dec_IR_reg[21]/NET0131 ,
		_w28203_,
		_w34844_
	);
	LUT2 #(
		.INIT('h8)
	) name30798 (
		\sice_IBR2_reg[15]/P0001 ,
		_w25074_,
		_w34845_
	);
	LUT2 #(
		.INIT('h8)
	) name30799 (
		_w25033_,
		_w25053_,
		_w34846_
	);
	LUT2 #(
		.INIT('h8)
	) name30800 (
		\sice_IMR1_reg[15]/NET0131 ,
		_w34846_,
		_w34847_
	);
	LUT2 #(
		.INIT('h1)
	) name30801 (
		_w25084_,
		_w34832_,
		_w34848_
	);
	LUT2 #(
		.INIT('h1)
	) name30802 (
		_w34833_,
		_w34834_,
		_w34849_
	);
	LUT2 #(
		.INIT('h1)
	) name30803 (
		_w34835_,
		_w34836_,
		_w34850_
	);
	LUT2 #(
		.INIT('h1)
	) name30804 (
		_w34837_,
		_w34838_,
		_w34851_
	);
	LUT2 #(
		.INIT('h1)
	) name30805 (
		_w34839_,
		_w34840_,
		_w34852_
	);
	LUT2 #(
		.INIT('h1)
	) name30806 (
		_w34842_,
		_w34843_,
		_w34853_
	);
	LUT2 #(
		.INIT('h1)
	) name30807 (
		_w34844_,
		_w34845_,
		_w34854_
	);
	LUT2 #(
		.INIT('h4)
	) name30808 (
		_w34847_,
		_w34854_,
		_w34855_
	);
	LUT2 #(
		.INIT('h8)
	) name30809 (
		_w34852_,
		_w34853_,
		_w34856_
	);
	LUT2 #(
		.INIT('h8)
	) name30810 (
		_w34850_,
		_w34851_,
		_w34857_
	);
	LUT2 #(
		.INIT('h8)
	) name30811 (
		_w34848_,
		_w34849_,
		_w34858_
	);
	LUT2 #(
		.INIT('h8)
	) name30812 (
		_w34857_,
		_w34858_,
		_w34859_
	);
	LUT2 #(
		.INIT('h8)
	) name30813 (
		_w34855_,
		_w34856_,
		_w34860_
	);
	LUT2 #(
		.INIT('h8)
	) name30814 (
		_w34859_,
		_w34860_,
		_w34861_
	);
	LUT2 #(
		.INIT('h8)
	) name30815 (
		_w34827_,
		_w34861_,
		_w34862_
	);
	LUT2 #(
		.INIT('h1)
	) name30816 (
		_w34830_,
		_w34862_,
		_w34863_
	);
	LUT2 #(
		.INIT('h2)
	) name30817 (
		_w18262_,
		_w24721_,
		_w34864_
	);
	LUT2 #(
		.INIT('h1)
	) name30818 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 ,
		_w28530_,
		_w34865_
	);
	LUT2 #(
		.INIT('h4)
	) name30819 (
		_w19381_,
		_w20259_,
		_w34866_
	);
	LUT2 #(
		.INIT('h2)
	) name30820 (
		_w28534_,
		_w34866_,
		_w34867_
	);
	LUT2 #(
		.INIT('h1)
	) name30821 (
		_w34865_,
		_w34867_,
		_w34868_
	);
	LUT2 #(
		.INIT('h1)
	) name30822 (
		_w19385_,
		_w34868_,
		_w34869_
	);
	LUT2 #(
		.INIT('h1)
	) name30823 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[5]/P0001 ,
		_w28532_,
		_w34870_
	);
	LUT2 #(
		.INIT('h1)
	) name30824 (
		_w34869_,
		_w34870_,
		_w34871_
	);
	LUT2 #(
		.INIT('h2)
	) name30825 (
		_w28529_,
		_w34871_,
		_w34872_
	);
	LUT2 #(
		.INIT('h1)
	) name30826 (
		_w34864_,
		_w34872_,
		_w34873_
	);
	LUT2 #(
		.INIT('h2)
	) name30827 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w10069_,
		_w34874_
	);
	LUT2 #(
		.INIT('h8)
	) name30828 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][12]/P0001 ,
		_w14702_,
		_w34875_
	);
	LUT2 #(
		.INIT('h8)
	) name30829 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][12]/P0001 ,
		_w14713_,
		_w34876_
	);
	LUT2 #(
		.INIT('h8)
	) name30830 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001 ,
		_w14704_,
		_w34877_
	);
	LUT2 #(
		.INIT('h8)
	) name30831 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][12]/P0001 ,
		_w14708_,
		_w34878_
	);
	LUT2 #(
		.INIT('h8)
	) name30832 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001 ,
		_w14711_,
		_w34879_
	);
	LUT2 #(
		.INIT('h8)
	) name30833 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001 ,
		_w14699_,
		_w34880_
	);
	LUT2 #(
		.INIT('h8)
	) name30834 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001 ,
		_w14706_,
		_w34881_
	);
	LUT2 #(
		.INIT('h1)
	) name30835 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w34875_,
		_w34882_
	);
	LUT2 #(
		.INIT('h1)
	) name30836 (
		_w34876_,
		_w34877_,
		_w34883_
	);
	LUT2 #(
		.INIT('h1)
	) name30837 (
		_w34878_,
		_w34879_,
		_w34884_
	);
	LUT2 #(
		.INIT('h1)
	) name30838 (
		_w34880_,
		_w34881_,
		_w34885_
	);
	LUT2 #(
		.INIT('h8)
	) name30839 (
		_w34884_,
		_w34885_,
		_w34886_
	);
	LUT2 #(
		.INIT('h8)
	) name30840 (
		_w34882_,
		_w34883_,
		_w34887_
	);
	LUT2 #(
		.INIT('h8)
	) name30841 (
		_w34886_,
		_w34887_,
		_w34888_
	);
	LUT2 #(
		.INIT('h4)
	) name30842 (
		\core_c_dec_IRE_reg[11]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w34889_
	);
	LUT2 #(
		.INIT('h2)
	) name30843 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w34255_,
		_w34890_
	);
	LUT2 #(
		.INIT('h4)
	) name30844 (
		_w34889_,
		_w34890_,
		_w34891_
	);
	LUT2 #(
		.INIT('h1)
	) name30845 (
		_w34888_,
		_w34891_,
		_w34892_
	);
	LUT2 #(
		.INIT('h1)
	) name30846 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w34892_,
		_w34893_
	);
	LUT2 #(
		.INIT('h1)
	) name30847 (
		_w34874_,
		_w34893_,
		_w34894_
	);
	LUT2 #(
		.INIT('h2)
	) name30848 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w7607_,
		_w34895_
	);
	LUT2 #(
		.INIT('h4)
	) name30849 (
		\core_c_dec_IRE_reg[7]/NET0131 ,
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w34896_
	);
	LUT2 #(
		.INIT('h8)
	) name30850 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_IRE_reg[7]/NET0131 ,
		_w34897_
	);
	LUT2 #(
		.INIT('h2)
	) name30851 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w34896_,
		_w34898_
	);
	LUT2 #(
		.INIT('h4)
	) name30852 (
		_w34897_,
		_w34898_,
		_w34899_
	);
	LUT2 #(
		.INIT('h8)
	) name30853 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001 ,
		_w14711_,
		_w34900_
	);
	LUT2 #(
		.INIT('h8)
	) name30854 (
		\core_c_psq_ststk_sts7x23_STcell_reg[1][8]/P0001 ,
		_w14708_,
		_w34901_
	);
	LUT2 #(
		.INIT('h8)
	) name30855 (
		\core_c_psq_ststk_sts7x23_STcell_reg[2][8]/P0001 ,
		_w14713_,
		_w34902_
	);
	LUT2 #(
		.INIT('h8)
	) name30856 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001 ,
		_w14704_,
		_w34903_
	);
	LUT2 #(
		.INIT('h8)
	) name30857 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001 ,
		_w14706_,
		_w34904_
	);
	LUT2 #(
		.INIT('h8)
	) name30858 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001 ,
		_w14699_,
		_w34905_
	);
	LUT2 #(
		.INIT('h8)
	) name30859 (
		\core_c_psq_ststk_sts7x23_STcell_reg[0][8]/P0001 ,
		_w14702_,
		_w34906_
	);
	LUT2 #(
		.INIT('h1)
	) name30860 (
		\core_c_dec_Modctl_Eg_reg/P0001 ,
		_w34900_,
		_w34907_
	);
	LUT2 #(
		.INIT('h1)
	) name30861 (
		_w34901_,
		_w34902_,
		_w34908_
	);
	LUT2 #(
		.INIT('h1)
	) name30862 (
		_w34903_,
		_w34904_,
		_w34909_
	);
	LUT2 #(
		.INIT('h1)
	) name30863 (
		_w34905_,
		_w34906_,
		_w34910_
	);
	LUT2 #(
		.INIT('h8)
	) name30864 (
		_w34909_,
		_w34910_,
		_w34911_
	);
	LUT2 #(
		.INIT('h8)
	) name30865 (
		_w34907_,
		_w34908_,
		_w34912_
	);
	LUT2 #(
		.INIT('h8)
	) name30866 (
		_w34911_,
		_w34912_,
		_w34913_
	);
	LUT2 #(
		.INIT('h1)
	) name30867 (
		_w34899_,
		_w34913_,
		_w34914_
	);
	LUT2 #(
		.INIT('h1)
	) name30868 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w34914_,
		_w34915_
	);
	LUT2 #(
		.INIT('h1)
	) name30869 (
		_w34895_,
		_w34915_,
		_w34916_
	);
	LUT2 #(
		.INIT('h8)
	) name30870 (
		\bdma_WRlat_reg/P0001 ,
		_w13150_,
		_w34917_
	);
	LUT2 #(
		.INIT('h2)
	) name30871 (
		\bdma_WRlat_reg/P0001 ,
		_w34065_,
		_w34918_
	);
	LUT2 #(
		.INIT('h2)
	) name30872 (
		\bdma_WRlat_reg/P0001 ,
		_w34060_,
		_w34919_
	);
	LUT2 #(
		.INIT('h2)
	) name30873 (
		\bdma_BWdataBUF_reg[6]/P0001 ,
		_w34919_,
		_w34920_
	);
	LUT2 #(
		.INIT('h8)
	) name30874 (
		\bdma_BWdataBUF_h_reg[6]/P0001 ,
		_w34919_,
		_w34921_
	);
	LUT2 #(
		.INIT('h1)
	) name30875 (
		_w34920_,
		_w34921_,
		_w34922_
	);
	LUT2 #(
		.INIT('h1)
	) name30876 (
		_w34918_,
		_w34922_,
		_w34923_
	);
	LUT2 #(
		.INIT('h8)
	) name30877 (
		\bdma_BWdataBUF_h_reg[14]/P0001 ,
		_w34918_,
		_w34924_
	);
	LUT2 #(
		.INIT('h1)
	) name30878 (
		_w34923_,
		_w34924_,
		_w34925_
	);
	LUT2 #(
		.INIT('h1)
	) name30879 (
		_w34917_,
		_w34925_,
		_w34926_
	);
	LUT2 #(
		.INIT('h8)
	) name30880 (
		\bdma_BWdataBUF_h_reg[22]/P0001 ,
		_w34917_,
		_w34927_
	);
	LUT2 #(
		.INIT('h1)
	) name30881 (
		_w34926_,
		_w34927_,
		_w34928_
	);
	LUT2 #(
		.INIT('h2)
	) name30882 (
		\bdma_BWdataBUF_reg[5]/P0001 ,
		_w34919_,
		_w34929_
	);
	LUT2 #(
		.INIT('h8)
	) name30883 (
		\bdma_BWdataBUF_h_reg[5]/P0001 ,
		_w34919_,
		_w34930_
	);
	LUT2 #(
		.INIT('h1)
	) name30884 (
		_w34929_,
		_w34930_,
		_w34931_
	);
	LUT2 #(
		.INIT('h1)
	) name30885 (
		_w34918_,
		_w34931_,
		_w34932_
	);
	LUT2 #(
		.INIT('h8)
	) name30886 (
		\bdma_BWdataBUF_h_reg[13]/P0001 ,
		_w34918_,
		_w34933_
	);
	LUT2 #(
		.INIT('h1)
	) name30887 (
		_w34932_,
		_w34933_,
		_w34934_
	);
	LUT2 #(
		.INIT('h1)
	) name30888 (
		_w34917_,
		_w34934_,
		_w34935_
	);
	LUT2 #(
		.INIT('h8)
	) name30889 (
		\bdma_BWdataBUF_h_reg[21]/P0001 ,
		_w34917_,
		_w34936_
	);
	LUT2 #(
		.INIT('h1)
	) name30890 (
		_w34935_,
		_w34936_,
		_w34937_
	);
	LUT2 #(
		.INIT('h2)
	) name30891 (
		\bdma_BWdataBUF_reg[7]/P0001 ,
		_w34919_,
		_w34938_
	);
	LUT2 #(
		.INIT('h8)
	) name30892 (
		\bdma_BWdataBUF_h_reg[7]/P0001 ,
		_w34919_,
		_w34939_
	);
	LUT2 #(
		.INIT('h1)
	) name30893 (
		_w34938_,
		_w34939_,
		_w34940_
	);
	LUT2 #(
		.INIT('h1)
	) name30894 (
		_w34918_,
		_w34940_,
		_w34941_
	);
	LUT2 #(
		.INIT('h8)
	) name30895 (
		\bdma_BWdataBUF_h_reg[15]/P0001 ,
		_w34918_,
		_w34942_
	);
	LUT2 #(
		.INIT('h1)
	) name30896 (
		_w34941_,
		_w34942_,
		_w34943_
	);
	LUT2 #(
		.INIT('h1)
	) name30897 (
		_w34917_,
		_w34943_,
		_w34944_
	);
	LUT2 #(
		.INIT('h8)
	) name30898 (
		\bdma_BWdataBUF_h_reg[23]/P0001 ,
		_w34917_,
		_w34945_
	);
	LUT2 #(
		.INIT('h1)
	) name30899 (
		_w34944_,
		_w34945_,
		_w34946_
	);
	LUT2 #(
		.INIT('h2)
	) name30900 (
		\bdma_BWdataBUF_reg[4]/P0001 ,
		_w34919_,
		_w34947_
	);
	LUT2 #(
		.INIT('h8)
	) name30901 (
		\bdma_BWdataBUF_h_reg[4]/P0001 ,
		_w34919_,
		_w34948_
	);
	LUT2 #(
		.INIT('h1)
	) name30902 (
		_w34947_,
		_w34948_,
		_w34949_
	);
	LUT2 #(
		.INIT('h1)
	) name30903 (
		_w34918_,
		_w34949_,
		_w34950_
	);
	LUT2 #(
		.INIT('h8)
	) name30904 (
		\bdma_BWdataBUF_h_reg[12]/P0001 ,
		_w34918_,
		_w34951_
	);
	LUT2 #(
		.INIT('h1)
	) name30905 (
		_w34950_,
		_w34951_,
		_w34952_
	);
	LUT2 #(
		.INIT('h1)
	) name30906 (
		_w34917_,
		_w34952_,
		_w34953_
	);
	LUT2 #(
		.INIT('h8)
	) name30907 (
		\bdma_BWdataBUF_h_reg[20]/P0001 ,
		_w34917_,
		_w34954_
	);
	LUT2 #(
		.INIT('h1)
	) name30908 (
		_w34953_,
		_w34954_,
		_w34955_
	);
	LUT2 #(
		.INIT('h2)
	) name30909 (
		\bdma_BWdataBUF_reg[3]/P0001 ,
		_w34919_,
		_w34956_
	);
	LUT2 #(
		.INIT('h8)
	) name30910 (
		\bdma_BWdataBUF_h_reg[3]/P0001 ,
		_w34919_,
		_w34957_
	);
	LUT2 #(
		.INIT('h1)
	) name30911 (
		_w34956_,
		_w34957_,
		_w34958_
	);
	LUT2 #(
		.INIT('h1)
	) name30912 (
		_w34918_,
		_w34958_,
		_w34959_
	);
	LUT2 #(
		.INIT('h8)
	) name30913 (
		\bdma_BWdataBUF_h_reg[11]/P0001 ,
		_w34918_,
		_w34960_
	);
	LUT2 #(
		.INIT('h1)
	) name30914 (
		_w34959_,
		_w34960_,
		_w34961_
	);
	LUT2 #(
		.INIT('h1)
	) name30915 (
		_w34917_,
		_w34961_,
		_w34962_
	);
	LUT2 #(
		.INIT('h8)
	) name30916 (
		\bdma_BWdataBUF_h_reg[19]/P0001 ,
		_w34917_,
		_w34963_
	);
	LUT2 #(
		.INIT('h1)
	) name30917 (
		_w34962_,
		_w34963_,
		_w34964_
	);
	LUT2 #(
		.INIT('h2)
	) name30918 (
		\bdma_BWdataBUF_reg[2]/P0001 ,
		_w34919_,
		_w34965_
	);
	LUT2 #(
		.INIT('h8)
	) name30919 (
		\bdma_BWdataBUF_h_reg[2]/P0001 ,
		_w34919_,
		_w34966_
	);
	LUT2 #(
		.INIT('h1)
	) name30920 (
		_w34965_,
		_w34966_,
		_w34967_
	);
	LUT2 #(
		.INIT('h1)
	) name30921 (
		_w34918_,
		_w34967_,
		_w34968_
	);
	LUT2 #(
		.INIT('h8)
	) name30922 (
		\bdma_BWdataBUF_h_reg[10]/P0001 ,
		_w34918_,
		_w34969_
	);
	LUT2 #(
		.INIT('h1)
	) name30923 (
		_w34968_,
		_w34969_,
		_w34970_
	);
	LUT2 #(
		.INIT('h1)
	) name30924 (
		_w34917_,
		_w34970_,
		_w34971_
	);
	LUT2 #(
		.INIT('h8)
	) name30925 (
		\bdma_BWdataBUF_h_reg[18]/P0001 ,
		_w34917_,
		_w34972_
	);
	LUT2 #(
		.INIT('h1)
	) name30926 (
		_w34971_,
		_w34972_,
		_w34973_
	);
	LUT2 #(
		.INIT('h2)
	) name30927 (
		\bdma_BWdataBUF_reg[1]/P0001 ,
		_w34919_,
		_w34974_
	);
	LUT2 #(
		.INIT('h8)
	) name30928 (
		\bdma_BWdataBUF_h_reg[1]/P0001 ,
		_w34919_,
		_w34975_
	);
	LUT2 #(
		.INIT('h1)
	) name30929 (
		_w34974_,
		_w34975_,
		_w34976_
	);
	LUT2 #(
		.INIT('h1)
	) name30930 (
		_w34918_,
		_w34976_,
		_w34977_
	);
	LUT2 #(
		.INIT('h8)
	) name30931 (
		\bdma_BWdataBUF_h_reg[9]/P0001 ,
		_w34918_,
		_w34978_
	);
	LUT2 #(
		.INIT('h1)
	) name30932 (
		_w34977_,
		_w34978_,
		_w34979_
	);
	LUT2 #(
		.INIT('h1)
	) name30933 (
		_w34917_,
		_w34979_,
		_w34980_
	);
	LUT2 #(
		.INIT('h8)
	) name30934 (
		\bdma_BWdataBUF_h_reg[17]/P0001 ,
		_w34917_,
		_w34981_
	);
	LUT2 #(
		.INIT('h1)
	) name30935 (
		_w34980_,
		_w34981_,
		_w34982_
	);
	LUT2 #(
		.INIT('h2)
	) name30936 (
		\bdma_BWdataBUF_reg[0]/P0001 ,
		_w34919_,
		_w34983_
	);
	LUT2 #(
		.INIT('h8)
	) name30937 (
		\bdma_BWdataBUF_h_reg[0]/P0001 ,
		_w34919_,
		_w34984_
	);
	LUT2 #(
		.INIT('h1)
	) name30938 (
		_w34983_,
		_w34984_,
		_w34985_
	);
	LUT2 #(
		.INIT('h1)
	) name30939 (
		_w34918_,
		_w34985_,
		_w34986_
	);
	LUT2 #(
		.INIT('h8)
	) name30940 (
		\bdma_BWdataBUF_h_reg[8]/P0001 ,
		_w34918_,
		_w34987_
	);
	LUT2 #(
		.INIT('h1)
	) name30941 (
		_w34986_,
		_w34987_,
		_w34988_
	);
	LUT2 #(
		.INIT('h1)
	) name30942 (
		_w34917_,
		_w34988_,
		_w34989_
	);
	LUT2 #(
		.INIT('h8)
	) name30943 (
		\bdma_BWdataBUF_h_reg[16]/P0001 ,
		_w34917_,
		_w34990_
	);
	LUT2 #(
		.INIT('h1)
	) name30944 (
		_w34989_,
		_w34990_,
		_w34991_
	);
	LUT2 #(
		.INIT('h8)
	) name30945 (
		\sice_SPC_reg[11]/P0001 ,
		_w34825_,
		_w34992_
	);
	LUT2 #(
		.INIT('h2)
	) name30946 (
		\sice_SPC_reg[13]/P0001 ,
		_w34825_,
		_w34993_
	);
	LUT2 #(
		.INIT('h1)
	) name30947 (
		_w34992_,
		_w34993_,
		_w34994_
	);
	LUT2 #(
		.INIT('h4)
	) name30948 (
		_w34827_,
		_w34994_,
		_w34995_
	);
	LUT2 #(
		.INIT('h8)
	) name30949 (
		\sice_DMR2_reg[6]/NET0131 ,
		_w25025_,
		_w34996_
	);
	LUT2 #(
		.INIT('h8)
	) name30950 (
		\sice_DBR1_reg[7]/P0001 ,
		_w25054_,
		_w34997_
	);
	LUT2 #(
		.INIT('h8)
	) name30951 (
		\sice_ITR_reg[2]/NET0131 ,
		_w25084_,
		_w34998_
	);
	LUT2 #(
		.INIT('h8)
	) name30952 (
		\sice_IMR1_reg[6]/NET0131 ,
		_w34846_,
		_w34999_
	);
	LUT2 #(
		.INIT('h8)
	) name30953 (
		\sice_idr1_reg_DO_reg[0]/P0001 ,
		_w26968_,
		_w35000_
	);
	LUT2 #(
		.INIT('h8)
	) name30954 (
		\sice_DMR1_reg[6]/NET0131 ,
		_w27903_,
		_w35001_
	);
	LUT2 #(
		.INIT('h8)
	) name30955 (
		\sice_IIRC_reg[12]/NET0131 ,
		_w24267_,
		_w35002_
	);
	LUT2 #(
		.INIT('h8)
	) name30956 (
		\sice_IMR2_reg[6]/NET0131 ,
		_w25034_,
		_w35003_
	);
	LUT2 #(
		.INIT('h8)
	) name30957 (
		\sice_IBR1_reg[6]/P0001 ,
		_w34831_,
		_w35004_
	);
	LUT2 #(
		.INIT('h8)
	) name30958 (
		\sice_DBR2_reg[7]/P0001 ,
		_w25012_,
		_w35005_
	);
	LUT2 #(
		.INIT('h8)
	) name30959 (
		\sice_IRR_reg[2]/P0001 ,
		_w34841_,
		_w35006_
	);
	LUT2 #(
		.INIT('h8)
	) name30960 (
		\sice_ICYC_reg[12]/NET0131 ,
		_w23409_,
		_w35007_
	);
	LUT2 #(
		.INIT('h4)
	) name30961 (
		\sice_IAR_reg[2]/NET0131 ,
		_w25083_,
		_w35008_
	);
	LUT2 #(
		.INIT('h8)
	) name30962 (
		\sice_IBR2_reg[6]/P0001 ,
		_w25074_,
		_w35009_
	);
	LUT2 #(
		.INIT('h8)
	) name30963 (
		\core_c_dec_IR_reg[12]/NET0131 ,
		_w28203_,
		_w35010_
	);
	LUT2 #(
		.INIT('h1)
	) name30964 (
		_w34996_,
		_w34997_,
		_w35011_
	);
	LUT2 #(
		.INIT('h1)
	) name30965 (
		_w34999_,
		_w35000_,
		_w35012_
	);
	LUT2 #(
		.INIT('h1)
	) name30966 (
		_w35001_,
		_w35002_,
		_w35013_
	);
	LUT2 #(
		.INIT('h1)
	) name30967 (
		_w35003_,
		_w35004_,
		_w35014_
	);
	LUT2 #(
		.INIT('h1)
	) name30968 (
		_w35005_,
		_w35006_,
		_w35015_
	);
	LUT2 #(
		.INIT('h1)
	) name30969 (
		_w35007_,
		_w35008_,
		_w35016_
	);
	LUT2 #(
		.INIT('h1)
	) name30970 (
		_w35009_,
		_w35010_,
		_w35017_
	);
	LUT2 #(
		.INIT('h8)
	) name30971 (
		_w35016_,
		_w35017_,
		_w35018_
	);
	LUT2 #(
		.INIT('h8)
	) name30972 (
		_w35014_,
		_w35015_,
		_w35019_
	);
	LUT2 #(
		.INIT('h8)
	) name30973 (
		_w35012_,
		_w35013_,
		_w35020_
	);
	LUT2 #(
		.INIT('h4)
	) name30974 (
		_w34998_,
		_w35011_,
		_w35021_
	);
	LUT2 #(
		.INIT('h8)
	) name30975 (
		_w35020_,
		_w35021_,
		_w35022_
	);
	LUT2 #(
		.INIT('h8)
	) name30976 (
		_w35018_,
		_w35019_,
		_w35023_
	);
	LUT2 #(
		.INIT('h8)
	) name30977 (
		_w35022_,
		_w35023_,
		_w35024_
	);
	LUT2 #(
		.INIT('h8)
	) name30978 (
		_w34827_,
		_w35024_,
		_w35025_
	);
	LUT2 #(
		.INIT('h1)
	) name30979 (
		_w34995_,
		_w35025_,
		_w35026_
	);
	LUT2 #(
		.INIT('h8)
	) name30980 (
		\sice_SPC_reg[10]/P0001 ,
		_w34825_,
		_w35027_
	);
	LUT2 #(
		.INIT('h2)
	) name30981 (
		\sice_SPC_reg[12]/P0001 ,
		_w34825_,
		_w35028_
	);
	LUT2 #(
		.INIT('h1)
	) name30982 (
		_w35027_,
		_w35028_,
		_w35029_
	);
	LUT2 #(
		.INIT('h4)
	) name30983 (
		_w34827_,
		_w35029_,
		_w35030_
	);
	LUT2 #(
		.INIT('h8)
	) name30984 (
		\sice_IBR2_reg[5]/P0001 ,
		_w25074_,
		_w35031_
	);
	LUT2 #(
		.INIT('h8)
	) name30985 (
		\sice_IMR2_reg[5]/NET0131 ,
		_w25034_,
		_w35032_
	);
	LUT2 #(
		.INIT('h8)
	) name30986 (
		\sice_ICYC_reg[11]/NET0131 ,
		_w23409_,
		_w35033_
	);
	LUT2 #(
		.INIT('h8)
	) name30987 (
		\sice_ITR_reg[1]/NET0131 ,
		_w25084_,
		_w35034_
	);
	LUT2 #(
		.INIT('h8)
	) name30988 (
		\sice_DBR1_reg[6]/P0001 ,
		_w25054_,
		_w35035_
	);
	LUT2 #(
		.INIT('h8)
	) name30989 (
		\core_c_dec_IR_reg[11]/NET0131 ,
		_w28203_,
		_w35036_
	);
	LUT2 #(
		.INIT('h8)
	) name30990 (
		\sice_IMR1_reg[5]/NET0131 ,
		_w34846_,
		_w35037_
	);
	LUT2 #(
		.INIT('h8)
	) name30991 (
		\sice_DMR2_reg[5]/NET0131 ,
		_w25025_,
		_w35038_
	);
	LUT2 #(
		.INIT('h8)
	) name30992 (
		\sice_IBR1_reg[5]/P0001 ,
		_w34831_,
		_w35039_
	);
	LUT2 #(
		.INIT('h8)
	) name30993 (
		\sice_idr0_reg_DO_reg[11]/P0001 ,
		_w26968_,
		_w35040_
	);
	LUT2 #(
		.INIT('h8)
	) name30994 (
		\sice_DBR2_reg[6]/P0001 ,
		_w25012_,
		_w35041_
	);
	LUT2 #(
		.INIT('h8)
	) name30995 (
		\sice_IIRC_reg[11]/NET0131 ,
		_w24267_,
		_w35042_
	);
	LUT2 #(
		.INIT('h8)
	) name30996 (
		\sice_DMR1_reg[5]/NET0131 ,
		_w27903_,
		_w35043_
	);
	LUT2 #(
		.INIT('h8)
	) name30997 (
		\sice_IRR_reg[1]/P0001 ,
		_w34841_,
		_w35044_
	);
	LUT2 #(
		.INIT('h1)
	) name30998 (
		_w35008_,
		_w35031_,
		_w35045_
	);
	LUT2 #(
		.INIT('h1)
	) name30999 (
		_w35032_,
		_w35033_,
		_w35046_
	);
	LUT2 #(
		.INIT('h1)
	) name31000 (
		_w35035_,
		_w35036_,
		_w35047_
	);
	LUT2 #(
		.INIT('h1)
	) name31001 (
		_w35037_,
		_w35038_,
		_w35048_
	);
	LUT2 #(
		.INIT('h1)
	) name31002 (
		_w35039_,
		_w35040_,
		_w35049_
	);
	LUT2 #(
		.INIT('h1)
	) name31003 (
		_w35041_,
		_w35042_,
		_w35050_
	);
	LUT2 #(
		.INIT('h1)
	) name31004 (
		_w35043_,
		_w35044_,
		_w35051_
	);
	LUT2 #(
		.INIT('h8)
	) name31005 (
		_w35050_,
		_w35051_,
		_w35052_
	);
	LUT2 #(
		.INIT('h8)
	) name31006 (
		_w35048_,
		_w35049_,
		_w35053_
	);
	LUT2 #(
		.INIT('h8)
	) name31007 (
		_w35046_,
		_w35047_,
		_w35054_
	);
	LUT2 #(
		.INIT('h4)
	) name31008 (
		_w35034_,
		_w35045_,
		_w35055_
	);
	LUT2 #(
		.INIT('h8)
	) name31009 (
		_w35054_,
		_w35055_,
		_w35056_
	);
	LUT2 #(
		.INIT('h8)
	) name31010 (
		_w35052_,
		_w35053_,
		_w35057_
	);
	LUT2 #(
		.INIT('h8)
	) name31011 (
		_w35056_,
		_w35057_,
		_w35058_
	);
	LUT2 #(
		.INIT('h8)
	) name31012 (
		_w34827_,
		_w35058_,
		_w35059_
	);
	LUT2 #(
		.INIT('h1)
	) name31013 (
		_w35030_,
		_w35059_,
		_w35060_
	);
	LUT2 #(
		.INIT('h8)
	) name31014 (
		\sice_SPC_reg[9]/P0001 ,
		_w34825_,
		_w35061_
	);
	LUT2 #(
		.INIT('h2)
	) name31015 (
		\sice_SPC_reg[11]/P0001 ,
		_w34825_,
		_w35062_
	);
	LUT2 #(
		.INIT('h1)
	) name31016 (
		_w35061_,
		_w35062_,
		_w35063_
	);
	LUT2 #(
		.INIT('h4)
	) name31017 (
		_w34827_,
		_w35063_,
		_w35064_
	);
	LUT2 #(
		.INIT('h8)
	) name31018 (
		\sice_IBR2_reg[4]/P0001 ,
		_w25074_,
		_w35065_
	);
	LUT2 #(
		.INIT('h8)
	) name31019 (
		\sice_IMR2_reg[4]/NET0131 ,
		_w25034_,
		_w35066_
	);
	LUT2 #(
		.INIT('h8)
	) name31020 (
		\sice_IIRC_reg[10]/NET0131 ,
		_w24267_,
		_w35067_
	);
	LUT2 #(
		.INIT('h8)
	) name31021 (
		\sice_ITR_reg[0]/NET0131 ,
		_w25084_,
		_w35068_
	);
	LUT2 #(
		.INIT('h8)
	) name31022 (
		\sice_DBR1_reg[5]/P0001 ,
		_w25054_,
		_w35069_
	);
	LUT2 #(
		.INIT('h8)
	) name31023 (
		\core_c_dec_IR_reg[10]/NET0131 ,
		_w28203_,
		_w35070_
	);
	LUT2 #(
		.INIT('h8)
	) name31024 (
		\sice_IMR1_reg[4]/NET0131 ,
		_w34846_,
		_w35071_
	);
	LUT2 #(
		.INIT('h8)
	) name31025 (
		\sice_ICYC_reg[10]/NET0131 ,
		_w23409_,
		_w35072_
	);
	LUT2 #(
		.INIT('h8)
	) name31026 (
		\sice_IBR1_reg[4]/P0001 ,
		_w34831_,
		_w35073_
	);
	LUT2 #(
		.INIT('h8)
	) name31027 (
		\sice_idr0_reg_DO_reg[10]/P0001 ,
		_w26968_,
		_w35074_
	);
	LUT2 #(
		.INIT('h8)
	) name31028 (
		\sice_DMR2_reg[4]/NET0131 ,
		_w25025_,
		_w35075_
	);
	LUT2 #(
		.INIT('h8)
	) name31029 (
		\sice_DBR2_reg[5]/P0001 ,
		_w25012_,
		_w35076_
	);
	LUT2 #(
		.INIT('h8)
	) name31030 (
		\sice_DMR1_reg[4]/NET0131 ,
		_w27903_,
		_w35077_
	);
	LUT2 #(
		.INIT('h8)
	) name31031 (
		\sice_IRR_reg[0]/P0001 ,
		_w34841_,
		_w35078_
	);
	LUT2 #(
		.INIT('h1)
	) name31032 (
		_w35008_,
		_w35065_,
		_w35079_
	);
	LUT2 #(
		.INIT('h1)
	) name31033 (
		_w35066_,
		_w35067_,
		_w35080_
	);
	LUT2 #(
		.INIT('h1)
	) name31034 (
		_w35069_,
		_w35070_,
		_w35081_
	);
	LUT2 #(
		.INIT('h1)
	) name31035 (
		_w35071_,
		_w35072_,
		_w35082_
	);
	LUT2 #(
		.INIT('h1)
	) name31036 (
		_w35073_,
		_w35074_,
		_w35083_
	);
	LUT2 #(
		.INIT('h1)
	) name31037 (
		_w35075_,
		_w35076_,
		_w35084_
	);
	LUT2 #(
		.INIT('h1)
	) name31038 (
		_w35077_,
		_w35078_,
		_w35085_
	);
	LUT2 #(
		.INIT('h8)
	) name31039 (
		_w35084_,
		_w35085_,
		_w35086_
	);
	LUT2 #(
		.INIT('h8)
	) name31040 (
		_w35082_,
		_w35083_,
		_w35087_
	);
	LUT2 #(
		.INIT('h8)
	) name31041 (
		_w35080_,
		_w35081_,
		_w35088_
	);
	LUT2 #(
		.INIT('h4)
	) name31042 (
		_w35068_,
		_w35079_,
		_w35089_
	);
	LUT2 #(
		.INIT('h8)
	) name31043 (
		_w35088_,
		_w35089_,
		_w35090_
	);
	LUT2 #(
		.INIT('h8)
	) name31044 (
		_w35086_,
		_w35087_,
		_w35091_
	);
	LUT2 #(
		.INIT('h8)
	) name31045 (
		_w35090_,
		_w35091_,
		_w35092_
	);
	LUT2 #(
		.INIT('h8)
	) name31046 (
		_w34827_,
		_w35092_,
		_w35093_
	);
	LUT2 #(
		.INIT('h1)
	) name31047 (
		_w35064_,
		_w35093_,
		_w35094_
	);
	LUT2 #(
		.INIT('h1)
	) name31048 (
		\sice_ICYC_reg[8]/NET0131 ,
		_w18863_,
		_w35095_
	);
	LUT2 #(
		.INIT('h1)
	) name31049 (
		_w20738_,
		_w35095_,
		_w35096_
	);
	LUT2 #(
		.INIT('h1)
	) name31050 (
		\clkc_oscntr_reg_DO_reg[6]/NET0131 ,
		_w23419_,
		_w35097_
	);
	LUT2 #(
		.INIT('h1)
	) name31051 (
		_w23420_,
		_w35097_,
		_w35098_
	);
	LUT2 #(
		.INIT('h8)
	) name31052 (
		_w18262_,
		_w25069_,
		_w35099_
	);
	LUT2 #(
		.INIT('h1)
	) name31053 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 ,
		_w28530_,
		_w35100_
	);
	LUT2 #(
		.INIT('h4)
	) name31054 (
		_w19381_,
		_w20080_,
		_w35101_
	);
	LUT2 #(
		.INIT('h2)
	) name31055 (
		_w28534_,
		_w35101_,
		_w35102_
	);
	LUT2 #(
		.INIT('h1)
	) name31056 (
		_w35100_,
		_w35102_,
		_w35103_
	);
	LUT2 #(
		.INIT('h1)
	) name31057 (
		_w19385_,
		_w35103_,
		_w35104_
	);
	LUT2 #(
		.INIT('h1)
	) name31058 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[4]/P0001 ,
		_w28532_,
		_w35105_
	);
	LUT2 #(
		.INIT('h1)
	) name31059 (
		_w35104_,
		_w35105_,
		_w35106_
	);
	LUT2 #(
		.INIT('h2)
	) name31060 (
		_w28529_,
		_w35106_,
		_w35107_
	);
	LUT2 #(
		.INIT('h1)
	) name31061 (
		_w35099_,
		_w35107_,
		_w35108_
	);
	LUT2 #(
		.INIT('h2)
	) name31062 (
		_w18262_,
		_w25088_,
		_w35109_
	);
	LUT2 #(
		.INIT('h1)
	) name31063 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 ,
		_w28530_,
		_w35110_
	);
	LUT2 #(
		.INIT('h4)
	) name31064 (
		_w19381_,
		_w19559_,
		_w35111_
	);
	LUT2 #(
		.INIT('h2)
	) name31065 (
		_w28534_,
		_w35111_,
		_w35112_
	);
	LUT2 #(
		.INIT('h1)
	) name31066 (
		_w35110_,
		_w35112_,
		_w35113_
	);
	LUT2 #(
		.INIT('h1)
	) name31067 (
		_w19385_,
		_w35113_,
		_w35114_
	);
	LUT2 #(
		.INIT('h1)
	) name31068 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[0]/P0001 ,
		_w28532_,
		_w35115_
	);
	LUT2 #(
		.INIT('h1)
	) name31069 (
		_w35114_,
		_w35115_,
		_w35116_
	);
	LUT2 #(
		.INIT('h2)
	) name31070 (
		_w28529_,
		_w35116_,
		_w35117_
	);
	LUT2 #(
		.INIT('h1)
	) name31071 (
		_w35109_,
		_w35117_,
		_w35118_
	);
	LUT2 #(
		.INIT('h8)
	) name31072 (
		_w6560_,
		_w6599_,
		_w35119_
	);
	LUT2 #(
		.INIT('h2)
	) name31073 (
		_w8198_,
		_w35119_,
		_w35120_
	);
	LUT2 #(
		.INIT('h2)
	) name31074 (
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w35120_,
		_w35121_
	);
	LUT2 #(
		.INIT('h8)
	) name31075 (
		_w6221_,
		_w6315_,
		_w35122_
	);
	LUT2 #(
		.INIT('h1)
	) name31076 (
		_w7631_,
		_w35122_,
		_w35123_
	);
	LUT2 #(
		.INIT('h1)
	) name31077 (
		\core_dag_ilm1reg_STEALI_E_reg[2]/P0001 ,
		_w35123_,
		_w35124_
	);
	LUT2 #(
		.INIT('h1)
	) name31078 (
		_w35121_,
		_w35124_,
		_w35125_
	);
	LUT2 #(
		.INIT('h8)
	) name31079 (
		\auctl_T0Sack_reg/NET0131 ,
		_w35125_,
		_w35126_
	);
	LUT2 #(
		.INIT('h8)
	) name31080 (
		\auctl_R0Sack_reg/NET0131 ,
		_w35125_,
		_w35127_
	);
	LUT2 #(
		.INIT('h8)
	) name31081 (
		\auctl_T1Sack_reg/NET0131 ,
		_w35125_,
		_w35128_
	);
	LUT2 #(
		.INIT('h8)
	) name31082 (
		\auctl_R1Sack_reg/NET0131 ,
		_w35125_,
		_w35129_
	);
	LUT2 #(
		.INIT('h8)
	) name31083 (
		\core_c_dec_MTIreg_E_reg[4]/P0001 ,
		_w4117_,
		_w35130_
	);
	LUT2 #(
		.INIT('h2)
	) name31084 (
		_w32000_,
		_w32001_,
		_w35131_
	);
	LUT2 #(
		.INIT('h8)
	) name31085 (
		_w31992_,
		_w35131_,
		_w35132_
	);
	LUT2 #(
		.INIT('h4)
	) name31086 (
		_w4117_,
		_w32007_,
		_w35133_
	);
	LUT2 #(
		.INIT('h4)
	) name31087 (
		_w32003_,
		_w35133_,
		_w35134_
	);
	LUT2 #(
		.INIT('h8)
	) name31088 (
		_w32014_,
		_w35134_,
		_w35135_
	);
	LUT2 #(
		.INIT('h8)
	) name31089 (
		_w35132_,
		_w35135_,
		_w35136_
	);
	LUT2 #(
		.INIT('h1)
	) name31090 (
		_w35130_,
		_w35136_,
		_w35137_
	);
	LUT2 #(
		.INIT('h2)
	) name31091 (
		_w4116_,
		_w35137_,
		_w35138_
	);
	LUT2 #(
		.INIT('h1)
	) name31092 (
		\core_c_dec_IRE_reg[0]/NET0131 ,
		\core_c_dec_IRE_reg[1]/NET0131 ,
		_w35139_
	);
	LUT2 #(
		.INIT('h4)
	) name31093 (
		\core_c_dec_IRE_reg[2]/NET0131 ,
		_w35139_,
		_w35140_
	);
	LUT2 #(
		.INIT('h2)
	) name31094 (
		\clkc_SIDLE_s1_reg/NET0131 ,
		\clkc_SIDLE_s2_reg/NET0131 ,
		_w35141_
	);
	LUT2 #(
		.INIT('h4)
	) name31095 (
		_w35140_,
		_w35141_,
		_w35142_
	);
	LUT2 #(
		.INIT('h4)
	) name31096 (
		\clkc_STBY_reg/NET0131 ,
		_w35142_,
		_w35143_
	);
	LUT2 #(
		.INIT('h1)
	) name31097 (
		\clkc_SlowDn_reg/NET0131 ,
		_w35142_,
		_w35144_
	);
	LUT2 #(
		.INIT('h2)
	) name31098 (
		_w23018_,
		_w35143_,
		_w35145_
	);
	LUT2 #(
		.INIT('h4)
	) name31099 (
		_w35144_,
		_w35145_,
		_w35146_
	);
	LUT2 #(
		.INIT('h8)
	) name31100 (
		_w33221_,
		_w35146_,
		_w35147_
	);
	LUT2 #(
		.INIT('h1)
	) name31101 (
		\clkc_STDcnt_reg[7]/NET0131 ,
		_w31527_,
		_w35148_
	);
	LUT2 #(
		.INIT('h1)
	) name31102 (
		_w31521_,
		_w31528_,
		_w35149_
	);
	LUT2 #(
		.INIT('h4)
	) name31103 (
		_w35148_,
		_w35149_,
		_w35150_
	);
	LUT2 #(
		.INIT('h8)
	) name31104 (
		\core_c_dec_MTIreg_E_reg[7]/P0001 ,
		_w4117_,
		_w35151_
	);
	LUT2 #(
		.INIT('h8)
	) name31105 (
		_w34465_,
		_w35132_,
		_w35152_
	);
	LUT2 #(
		.INIT('h1)
	) name31106 (
		_w35151_,
		_w35152_,
		_w35153_
	);
	LUT2 #(
		.INIT('h2)
	) name31107 (
		_w4116_,
		_w35153_,
		_w35154_
	);
	LUT2 #(
		.INIT('h8)
	) name31108 (
		\core_c_dec_MTDMOVL_E_reg/P0001 ,
		_w4117_,
		_w35155_
	);
	LUT2 #(
		.INIT('h8)
	) name31109 (
		_w32020_,
		_w34463_,
		_w35156_
	);
	LUT2 #(
		.INIT('h1)
	) name31110 (
		_w35155_,
		_w35156_,
		_w35157_
	);
	LUT2 #(
		.INIT('h2)
	) name31111 (
		_w4116_,
		_w35157_,
		_w35158_
	);
	LUT2 #(
		.INIT('h4)
	) name31112 (
		\core_c_dec_MTASTAT_E_reg/P0001 ,
		_w4117_,
		_w35159_
	);
	LUT2 #(
		.INIT('h1)
	) name31113 (
		_w4117_,
		_w32017_,
		_w35160_
	);
	LUT2 #(
		.INIT('h2)
	) name31114 (
		_w4116_,
		_w35159_,
		_w35161_
	);
	LUT2 #(
		.INIT('h4)
	) name31115 (
		_w35160_,
		_w35161_,
		_w35162_
	);
	LUT2 #(
		.INIT('h8)
	) name31116 (
		\core_c_dec_MTSB_E_reg/P0001 ,
		_w4117_,
		_w35163_
	);
	LUT2 #(
		.INIT('h8)
	) name31117 (
		_w32004_,
		_w35133_,
		_w35164_
	);
	LUT2 #(
		.INIT('h8)
	) name31118 (
		_w31992_,
		_w31999_,
		_w35165_
	);
	LUT2 #(
		.INIT('h8)
	) name31119 (
		_w35164_,
		_w35165_,
		_w35166_
	);
	LUT2 #(
		.INIT('h1)
	) name31120 (
		_w35163_,
		_w35166_,
		_w35167_
	);
	LUT2 #(
		.INIT('h2)
	) name31121 (
		_w4116_,
		_w35167_,
		_w35168_
	);
	LUT2 #(
		.INIT('h8)
	) name31122 (
		\core_c_dec_MTRX1_E_reg/P0001 ,
		_w4117_,
		_w35169_
	);
	LUT2 #(
		.INIT('h8)
	) name31123 (
		_w34462_,
		_w35134_,
		_w35170_
	);
	LUT2 #(
		.INIT('h8)
	) name31124 (
		_w32018_,
		_w35170_,
		_w35171_
	);
	LUT2 #(
		.INIT('h1)
	) name31125 (
		_w35169_,
		_w35171_,
		_w35172_
	);
	LUT2 #(
		.INIT('h2)
	) name31126 (
		_w4116_,
		_w35172_,
		_w35173_
	);
	LUT2 #(
		.INIT('h8)
	) name31127 (
		\core_c_dec_MTRX0_E_reg/P0001 ,
		_w4117_,
		_w35174_
	);
	LUT2 #(
		.INIT('h8)
	) name31128 (
		_w32018_,
		_w35135_,
		_w35175_
	);
	LUT2 #(
		.INIT('h1)
	) name31129 (
		_w35174_,
		_w35175_,
		_w35176_
	);
	LUT2 #(
		.INIT('h2)
	) name31130 (
		_w4116_,
		_w35176_,
		_w35177_
	);
	LUT2 #(
		.INIT('h8)
	) name31131 (
		\core_c_dec_MTPMOVL_E_reg/P0001 ,
		_w4117_,
		_w35178_
	);
	LUT2 #(
		.INIT('h8)
	) name31132 (
		_w32020_,
		_w35133_,
		_w35179_
	);
	LUT2 #(
		.INIT('h1)
	) name31133 (
		_w35178_,
		_w35179_,
		_w35180_
	);
	LUT2 #(
		.INIT('h2)
	) name31134 (
		_w4116_,
		_w35180_,
		_w35181_
	);
	LUT2 #(
		.INIT('h8)
	) name31135 (
		\core_c_dec_MTOWRCNTR_Eg_reg/P0001 ,
		_w4117_,
		_w35182_
	);
	LUT2 #(
		.INIT('h4)
	) name31136 (
		_w31995_,
		_w31998_,
		_w35183_
	);
	LUT2 #(
		.INIT('h8)
	) name31137 (
		_w11741_,
		_w35183_,
		_w35184_
	);
	LUT2 #(
		.INIT('h4)
	) name31138 (
		_w31992_,
		_w35184_,
		_w35185_
	);
	LUT2 #(
		.INIT('h8)
	) name31139 (
		_w32004_,
		_w34463_,
		_w35186_
	);
	LUT2 #(
		.INIT('h8)
	) name31140 (
		_w35185_,
		_w35186_,
		_w35187_
	);
	LUT2 #(
		.INIT('h1)
	) name31141 (
		_w35182_,
		_w35187_,
		_w35188_
	);
	LUT2 #(
		.INIT('h2)
	) name31142 (
		_w4116_,
		_w35188_,
		_w35189_
	);
	LUT2 #(
		.INIT('h8)
	) name31143 (
		\core_c_dec_MTMreg_E_reg[7]/P0001 ,
		_w4117_,
		_w35190_
	);
	LUT2 #(
		.INIT('h8)
	) name31144 (
		_w34464_,
		_w35132_,
		_w35191_
	);
	LUT2 #(
		.INIT('h8)
	) name31145 (
		_w31999_,
		_w35191_,
		_w35192_
	);
	LUT2 #(
		.INIT('h1)
	) name31146 (
		_w35190_,
		_w35192_,
		_w35193_
	);
	LUT2 #(
		.INIT('h2)
	) name31147 (
		_w4116_,
		_w35193_,
		_w35194_
	);
	LUT2 #(
		.INIT('h8)
	) name31148 (
		\core_c_dec_MTMreg_E_reg[6]/P0001 ,
		_w4117_,
		_w35195_
	);
	LUT2 #(
		.INIT('h8)
	) name31149 (
		_w35132_,
		_w35134_,
		_w35196_
	);
	LUT2 #(
		.INIT('h8)
	) name31150 (
		_w31999_,
		_w35196_,
		_w35197_
	);
	LUT2 #(
		.INIT('h1)
	) name31151 (
		_w35195_,
		_w35197_,
		_w35198_
	);
	LUT2 #(
		.INIT('h2)
	) name31152 (
		_w4116_,
		_w35198_,
		_w35199_
	);
	LUT2 #(
		.INIT('h8)
	) name31153 (
		\core_c_dec_MTMreg_E_reg[5]/P0001 ,
		_w4117_,
		_w35200_
	);
	LUT2 #(
		.INIT('h8)
	) name31154 (
		_w35183_,
		_w35191_,
		_w35201_
	);
	LUT2 #(
		.INIT('h1)
	) name31155 (
		_w35200_,
		_w35201_,
		_w35202_
	);
	LUT2 #(
		.INIT('h2)
	) name31156 (
		_w4116_,
		_w35202_,
		_w35203_
	);
	LUT2 #(
		.INIT('h8)
	) name31157 (
		\core_c_dec_MTMreg_E_reg[4]/P0001 ,
		_w4117_,
		_w35204_
	);
	LUT2 #(
		.INIT('h8)
	) name31158 (
		_w35183_,
		_w35196_,
		_w35205_
	);
	LUT2 #(
		.INIT('h1)
	) name31159 (
		_w35204_,
		_w35205_,
		_w35206_
	);
	LUT2 #(
		.INIT('h2)
	) name31160 (
		_w4116_,
		_w35206_,
		_w35207_
	);
	LUT2 #(
		.INIT('h1)
	) name31161 (
		_w31998_,
		_w32007_,
		_w35208_
	);
	LUT2 #(
		.INIT('h8)
	) name31162 (
		_w34479_,
		_w35208_,
		_w35209_
	);
	LUT2 #(
		.INIT('h8)
	) name31163 (
		_w34476_,
		_w35209_,
		_w35210_
	);
	LUT2 #(
		.INIT('h8)
	) name31164 (
		\core_c_dec_MTMreg_E_reg[3]/P0001 ,
		_w4117_,
		_w35211_
	);
	LUT2 #(
		.INIT('h1)
	) name31165 (
		_w35210_,
		_w35211_,
		_w35212_
	);
	LUT2 #(
		.INIT('h2)
	) name31166 (
		_w4116_,
		_w35212_,
		_w35213_
	);
	LUT2 #(
		.INIT('h4)
	) name31167 (
		_w31998_,
		_w32007_,
		_w35214_
	);
	LUT2 #(
		.INIT('h8)
	) name31168 (
		_w34479_,
		_w35214_,
		_w35215_
	);
	LUT2 #(
		.INIT('h8)
	) name31169 (
		_w34476_,
		_w35215_,
		_w35216_
	);
	LUT2 #(
		.INIT('h8)
	) name31170 (
		\core_c_dec_MTMreg_E_reg[2]/P0001 ,
		_w4117_,
		_w35217_
	);
	LUT2 #(
		.INIT('h1)
	) name31171 (
		_w35216_,
		_w35217_,
		_w35218_
	);
	LUT2 #(
		.INIT('h2)
	) name31172 (
		_w4116_,
		_w35218_,
		_w35219_
	);
	LUT2 #(
		.INIT('h8)
	) name31173 (
		\core_c_dec_MTMreg_E_reg[0]/P0001 ,
		_w4117_,
		_w35220_
	);
	LUT2 #(
		.INIT('h8)
	) name31174 (
		_w34475_,
		_w34479_,
		_w35221_
	);
	LUT2 #(
		.INIT('h8)
	) name31175 (
		_w32007_,
		_w35183_,
		_w35222_
	);
	LUT2 #(
		.INIT('h8)
	) name31176 (
		_w35221_,
		_w35222_,
		_w35223_
	);
	LUT2 #(
		.INIT('h1)
	) name31177 (
		_w35220_,
		_w35223_,
		_w35224_
	);
	LUT2 #(
		.INIT('h2)
	) name31178 (
		_w4116_,
		_w35224_,
		_w35225_
	);
	LUT2 #(
		.INIT('h4)
	) name31179 (
		_w31992_,
		_w35131_,
		_w35226_
	);
	LUT2 #(
		.INIT('h8)
	) name31180 (
		_w34465_,
		_w35226_,
		_w35227_
	);
	LUT2 #(
		.INIT('h8)
	) name31181 (
		\core_c_dec_MTLreg_E_reg[7]/P0001 ,
		_w4117_,
		_w35228_
	);
	LUT2 #(
		.INIT('h1)
	) name31182 (
		_w35227_,
		_w35228_,
		_w35229_
	);
	LUT2 #(
		.INIT('h2)
	) name31183 (
		_w4116_,
		_w35229_,
		_w35230_
	);
	LUT2 #(
		.INIT('h8)
	) name31184 (
		_w35170_,
		_w35226_,
		_w35231_
	);
	LUT2 #(
		.INIT('h8)
	) name31185 (
		\core_c_dec_MTLreg_E_reg[6]/P0001 ,
		_w4117_,
		_w35232_
	);
	LUT2 #(
		.INIT('h1)
	) name31186 (
		_w35231_,
		_w35232_,
		_w35233_
	);
	LUT2 #(
		.INIT('h2)
	) name31187 (
		_w4116_,
		_w35233_,
		_w35234_
	);
	LUT2 #(
		.INIT('h8)
	) name31188 (
		_w34470_,
		_w35226_,
		_w35235_
	);
	LUT2 #(
		.INIT('h8)
	) name31189 (
		\core_c_dec_MTLreg_E_reg[5]/P0001 ,
		_w4117_,
		_w35236_
	);
	LUT2 #(
		.INIT('h1)
	) name31190 (
		_w35235_,
		_w35236_,
		_w35237_
	);
	LUT2 #(
		.INIT('h2)
	) name31191 (
		_w4116_,
		_w35237_,
		_w35238_
	);
	LUT2 #(
		.INIT('h8)
	) name31192 (
		\core_c_dec_MTLreg_E_reg[4]/P0001 ,
		_w4117_,
		_w35239_
	);
	LUT2 #(
		.INIT('h8)
	) name31193 (
		_w35135_,
		_w35226_,
		_w35240_
	);
	LUT2 #(
		.INIT('h1)
	) name31194 (
		_w35239_,
		_w35240_,
		_w35241_
	);
	LUT2 #(
		.INIT('h2)
	) name31195 (
		_w4116_,
		_w35241_,
		_w35242_
	);
	LUT2 #(
		.INIT('h8)
	) name31196 (
		\core_c_dec_MTLreg_E_reg[3]/P0001 ,
		_w4117_,
		_w35243_
	);
	LUT2 #(
		.INIT('h4)
	) name31197 (
		_w4117_,
		_w32019_,
		_w35244_
	);
	LUT2 #(
		.INIT('h8)
	) name31198 (
		_w31995_,
		_w35244_,
		_w35245_
	);
	LUT2 #(
		.INIT('h8)
	) name31199 (
		_w35208_,
		_w35245_,
		_w35246_
	);
	LUT2 #(
		.INIT('h1)
	) name31200 (
		_w35243_,
		_w35246_,
		_w35247_
	);
	LUT2 #(
		.INIT('h2)
	) name31201 (
		_w4116_,
		_w35247_,
		_w35248_
	);
	LUT2 #(
		.INIT('h8)
	) name31202 (
		\core_c_dec_MTLreg_E_reg[2]/P0001 ,
		_w4117_,
		_w35249_
	);
	LUT2 #(
		.INIT('h8)
	) name31203 (
		_w35214_,
		_w35245_,
		_w35250_
	);
	LUT2 #(
		.INIT('h1)
	) name31204 (
		_w35249_,
		_w35250_,
		_w35251_
	);
	LUT2 #(
		.INIT('h2)
	) name31205 (
		_w4116_,
		_w35251_,
		_w35252_
	);
	LUT2 #(
		.INIT('h8)
	) name31206 (
		\core_c_dec_MTLreg_E_reg[1]/P0001 ,
		_w4117_,
		_w35253_
	);
	LUT2 #(
		.INIT('h8)
	) name31207 (
		_w34477_,
		_w35245_,
		_w35254_
	);
	LUT2 #(
		.INIT('h1)
	) name31208 (
		_w35253_,
		_w35254_,
		_w35255_
	);
	LUT2 #(
		.INIT('h2)
	) name31209 (
		_w4116_,
		_w35255_,
		_w35256_
	);
	LUT2 #(
		.INIT('h8)
	) name31210 (
		\core_c_dec_MTLreg_E_reg[0]/P0001 ,
		_w4117_,
		_w35257_
	);
	LUT2 #(
		.INIT('h8)
	) name31211 (
		_w32015_,
		_w35244_,
		_w35258_
	);
	LUT2 #(
		.INIT('h1)
	) name31212 (
		_w35257_,
		_w35258_,
		_w35259_
	);
	LUT2 #(
		.INIT('h2)
	) name31213 (
		_w4116_,
		_w35259_,
		_w35260_
	);
	LUT2 #(
		.INIT('h8)
	) name31214 (
		\core_c_dec_MTIreg_E_reg[6]/P0001 ,
		_w4117_,
		_w35261_
	);
	LUT2 #(
		.INIT('h8)
	) name31215 (
		_w35132_,
		_w35170_,
		_w35262_
	);
	LUT2 #(
		.INIT('h1)
	) name31216 (
		_w35261_,
		_w35262_,
		_w35263_
	);
	LUT2 #(
		.INIT('h2)
	) name31217 (
		_w4116_,
		_w35263_,
		_w35264_
	);
	LUT2 #(
		.INIT('h8)
	) name31218 (
		\core_c_dec_MTIreg_E_reg[5]/P0001 ,
		_w4117_,
		_w35265_
	);
	LUT2 #(
		.INIT('h8)
	) name31219 (
		_w34470_,
		_w35132_,
		_w35266_
	);
	LUT2 #(
		.INIT('h1)
	) name31220 (
		_w35265_,
		_w35266_,
		_w35267_
	);
	LUT2 #(
		.INIT('h2)
	) name31221 (
		_w4116_,
		_w35267_,
		_w35268_
	);
	LUT2 #(
		.INIT('h8)
	) name31222 (
		_w31995_,
		_w34475_,
		_w35269_
	);
	LUT2 #(
		.INIT('h8)
	) name31223 (
		_w35209_,
		_w35269_,
		_w35270_
	);
	LUT2 #(
		.INIT('h8)
	) name31224 (
		\core_c_dec_MTIreg_E_reg[3]/P0001 ,
		_w4117_,
		_w35271_
	);
	LUT2 #(
		.INIT('h1)
	) name31225 (
		_w35270_,
		_w35271_,
		_w35272_
	);
	LUT2 #(
		.INIT('h2)
	) name31226 (
		_w4116_,
		_w35272_,
		_w35273_
	);
	LUT2 #(
		.INIT('h8)
	) name31227 (
		_w35215_,
		_w35269_,
		_w35274_
	);
	LUT2 #(
		.INIT('h8)
	) name31228 (
		\core_c_dec_MTIreg_E_reg[2]/P0001 ,
		_w4117_,
		_w35275_
	);
	LUT2 #(
		.INIT('h1)
	) name31229 (
		_w35274_,
		_w35275_,
		_w35276_
	);
	LUT2 #(
		.INIT('h2)
	) name31230 (
		_w4116_,
		_w35276_,
		_w35277_
	);
	LUT2 #(
		.INIT('h8)
	) name31231 (
		\core_c_dec_MTIreg_E_reg[1]/P0001 ,
		_w4117_,
		_w35278_
	);
	LUT2 #(
		.INIT('h8)
	) name31232 (
		_w34480_,
		_w35269_,
		_w35279_
	);
	LUT2 #(
		.INIT('h1)
	) name31233 (
		_w35278_,
		_w35279_,
		_w35280_
	);
	LUT2 #(
		.INIT('h2)
	) name31234 (
		_w4116_,
		_w35280_,
		_w35281_
	);
	LUT2 #(
		.INIT('h8)
	) name31235 (
		_w14752_,
		_w25069_,
		_w35282_
	);
	LUT2 #(
		.INIT('h1)
	) name31236 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 ,
		_w17799_,
		_w35283_
	);
	LUT2 #(
		.INIT('h4)
	) name31237 (
		_w17809_,
		_w20080_,
		_w35284_
	);
	LUT2 #(
		.INIT('h2)
	) name31238 (
		_w17811_,
		_w35284_,
		_w35285_
	);
	LUT2 #(
		.INIT('h1)
	) name31239 (
		_w35283_,
		_w35285_,
		_w35286_
	);
	LUT2 #(
		.INIT('h1)
	) name31240 (
		_w17823_,
		_w35286_,
		_w35287_
	);
	LUT2 #(
		.INIT('h1)
	) name31241 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[4]/P0001 ,
		_w17808_,
		_w35288_
	);
	LUT2 #(
		.INIT('h1)
	) name31242 (
		_w35287_,
		_w35288_,
		_w35289_
	);
	LUT2 #(
		.INIT('h2)
	) name31243 (
		_w17829_,
		_w35289_,
		_w35290_
	);
	LUT2 #(
		.INIT('h1)
	) name31244 (
		_w35282_,
		_w35290_,
		_w35291_
	);
	LUT2 #(
		.INIT('h8)
	) name31245 (
		\core_c_dec_MTIreg_E_reg[0]/P0001 ,
		_w4117_,
		_w35292_
	);
	LUT2 #(
		.INIT('h8)
	) name31246 (
		_w32015_,
		_w35221_,
		_w35293_
	);
	LUT2 #(
		.INIT('h1)
	) name31247 (
		_w35292_,
		_w35293_,
		_w35294_
	);
	LUT2 #(
		.INIT('h2)
	) name31248 (
		_w4116_,
		_w35294_,
		_w35295_
	);
	LUT2 #(
		.INIT('h8)
	) name31249 (
		\core_c_dec_MTIFC_Eg_reg/P0001 ,
		_w4117_,
		_w35296_
	);
	LUT2 #(
		.INIT('h8)
	) name31250 (
		_w35164_,
		_w35185_,
		_w35297_
	);
	LUT2 #(
		.INIT('h1)
	) name31251 (
		_w35296_,
		_w35297_,
		_w35298_
	);
	LUT2 #(
		.INIT('h2)
	) name31252 (
		_w4116_,
		_w35298_,
		_w35299_
	);
	LUT2 #(
		.INIT('h8)
	) name31253 (
		\core_c_dec_MTIDR_E_reg/P0001 ,
		_w4117_,
		_w35300_
	);
	LUT2 #(
		.INIT('h8)
	) name31254 (
		_w35222_,
		_w35244_,
		_w35301_
	);
	LUT2 #(
		.INIT('h1)
	) name31255 (
		_w35300_,
		_w35301_,
		_w35302_
	);
	LUT2 #(
		.INIT('h2)
	) name31256 (
		_w4116_,
		_w35302_,
		_w35303_
	);
	LUT2 #(
		.INIT('h8)
	) name31257 (
		\core_c_dec_MTICNTL_Eg_reg/P0001 ,
		_w4117_,
		_w35304_
	);
	LUT2 #(
		.INIT('h8)
	) name31258 (
		_w31992_,
		_w35184_,
		_w35305_
	);
	LUT2 #(
		.INIT('h8)
	) name31259 (
		_w35164_,
		_w35305_,
		_w35306_
	);
	LUT2 #(
		.INIT('h1)
	) name31260 (
		_w35304_,
		_w35306_,
		_w35307_
	);
	LUT2 #(
		.INIT('h2)
	) name31261 (
		_w4116_,
		_w35307_,
		_w35308_
	);
	LUT2 #(
		.INIT('h8)
	) name31262 (
		\core_c_dec_MTCNTR_Eg_reg/P0001 ,
		_w4117_,
		_w35309_
	);
	LUT2 #(
		.INIT('h8)
	) name31263 (
		_w35186_,
		_w35305_,
		_w35310_
	);
	LUT2 #(
		.INIT('h1)
	) name31264 (
		_w35309_,
		_w35310_,
		_w35311_
	);
	LUT2 #(
		.INIT('h2)
	) name31265 (
		_w4116_,
		_w35311_,
		_w35312_
	);
	LUT2 #(
		.INIT('h2)
	) name31266 (
		\bdma_BWCOUNT_reg[1]/NET0131 ,
		_w13764_,
		_w35313_
	);
	LUT2 #(
		.INIT('h1)
	) name31267 (
		_w13763_,
		_w13765_,
		_w35314_
	);
	LUT2 #(
		.INIT('h4)
	) name31268 (
		_w35313_,
		_w35314_,
		_w35315_
	);
	LUT2 #(
		.INIT('h4)
	) name31269 (
		_w9435_,
		_w13763_,
		_w35316_
	);
	LUT2 #(
		.INIT('h1)
	) name31270 (
		_w35315_,
		_w35316_,
		_w35317_
	);
	LUT2 #(
		.INIT('h2)
	) name31271 (
		_w13746_,
		_w34589_,
		_w35318_
	);
	LUT2 #(
		.INIT('h4)
	) name31272 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w19205_,
		_w35319_
	);
	LUT2 #(
		.INIT('h4)
	) name31273 (
		_w19205_,
		_w19296_,
		_w35320_
	);
	LUT2 #(
		.INIT('h2)
	) name31274 (
		_w4150_,
		_w35319_,
		_w35321_
	);
	LUT2 #(
		.INIT('h4)
	) name31275 (
		_w35320_,
		_w35321_,
		_w35322_
	);
	LUT2 #(
		.INIT('h2)
	) name31276 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w19848_,
		_w35323_
	);
	LUT2 #(
		.INIT('h4)
	) name31277 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w29942_,
		_w35324_
	);
	LUT2 #(
		.INIT('h1)
	) name31278 (
		_w35323_,
		_w35324_,
		_w35325_
	);
	LUT2 #(
		.INIT('h2)
	) name31279 (
		_w18717_,
		_w35325_,
		_w35326_
	);
	LUT2 #(
		.INIT('h1)
	) name31280 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[10]/P0001 ,
		_w18717_,
		_w35327_
	);
	LUT2 #(
		.INIT('h1)
	) name31281 (
		_w35326_,
		_w35327_,
		_w35328_
	);
	LUT2 #(
		.INIT('h2)
	) name31282 (
		_w17833_,
		_w35325_,
		_w35329_
	);
	LUT2 #(
		.INIT('h1)
	) name31283 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[10]/P0001 ,
		_w17833_,
		_w35330_
	);
	LUT2 #(
		.INIT('h1)
	) name31284 (
		_w35329_,
		_w35330_,
		_w35331_
	);
	LUT2 #(
		.INIT('h2)
	) name31285 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w23860_,
		_w35332_
	);
	LUT2 #(
		.INIT('h4)
	) name31286 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w30441_,
		_w35333_
	);
	LUT2 #(
		.INIT('h1)
	) name31287 (
		_w35332_,
		_w35333_,
		_w35334_
	);
	LUT2 #(
		.INIT('h2)
	) name31288 (
		_w18886_,
		_w35334_,
		_w35335_
	);
	LUT2 #(
		.INIT('h1)
	) name31289 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[8]/P0001 ,
		_w18886_,
		_w35336_
	);
	LUT2 #(
		.INIT('h1)
	) name31290 (
		_w35335_,
		_w35336_,
		_w35337_
	);
	LUT2 #(
		.INIT('h2)
	) name31291 (
		_w19034_,
		_w35334_,
		_w35338_
	);
	LUT2 #(
		.INIT('h1)
	) name31292 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[8]/P0001 ,
		_w19034_,
		_w35339_
	);
	LUT2 #(
		.INIT('h1)
	) name31293 (
		_w35338_,
		_w35339_,
		_w35340_
	);
	LUT2 #(
		.INIT('h2)
	) name31294 (
		_w14752_,
		_w24721_,
		_w35341_
	);
	LUT2 #(
		.INIT('h1)
	) name31295 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 ,
		_w17799_,
		_w35342_
	);
	LUT2 #(
		.INIT('h4)
	) name31296 (
		_w17809_,
		_w20259_,
		_w35343_
	);
	LUT2 #(
		.INIT('h2)
	) name31297 (
		_w17811_,
		_w35343_,
		_w35344_
	);
	LUT2 #(
		.INIT('h1)
	) name31298 (
		_w35342_,
		_w35344_,
		_w35345_
	);
	LUT2 #(
		.INIT('h1)
	) name31299 (
		_w17823_,
		_w35345_,
		_w35346_
	);
	LUT2 #(
		.INIT('h1)
	) name31300 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[5]/P0001 ,
		_w17808_,
		_w35347_
	);
	LUT2 #(
		.INIT('h1)
	) name31301 (
		_w35346_,
		_w35347_,
		_w35348_
	);
	LUT2 #(
		.INIT('h2)
	) name31302 (
		_w17829_,
		_w35348_,
		_w35349_
	);
	LUT2 #(
		.INIT('h1)
	) name31303 (
		_w35341_,
		_w35349_,
		_w35350_
	);
	LUT2 #(
		.INIT('h2)
	) name31304 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 ,
		_w18266_,
		_w35351_
	);
	LUT2 #(
		.INIT('h1)
	) name31305 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[8]/P0001 ,
		_w18271_,
		_w35352_
	);
	LUT2 #(
		.INIT('h2)
	) name31306 (
		_w18271_,
		_w23860_,
		_w35353_
	);
	LUT2 #(
		.INIT('h2)
	) name31307 (
		_w18273_,
		_w35352_,
		_w35354_
	);
	LUT2 #(
		.INIT('h4)
	) name31308 (
		_w35353_,
		_w35354_,
		_w35355_
	);
	LUT2 #(
		.INIT('h1)
	) name31309 (
		_w18270_,
		_w35351_,
		_w35356_
	);
	LUT2 #(
		.INIT('h4)
	) name31310 (
		_w35355_,
		_w35356_,
		_w35357_
	);
	LUT2 #(
		.INIT('h1)
	) name31311 (
		_w18262_,
		_w35357_,
		_w35358_
	);
	LUT2 #(
		.INIT('h8)
	) name31312 (
		_w18262_,
		_w19633_,
		_w35359_
	);
	LUT2 #(
		.INIT('h1)
	) name31313 (
		_w35358_,
		_w35359_,
		_w35360_
	);
	LUT2 #(
		.INIT('h2)
	) name31314 (
		_w14752_,
		_w19633_,
		_w35361_
	);
	LUT2 #(
		.INIT('h8)
	) name31315 (
		_w18328_,
		_w23860_,
		_w35362_
	);
	LUT2 #(
		.INIT('h2)
	) name31316 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[8]/P0001 ,
		_w18330_,
		_w35363_
	);
	LUT2 #(
		.INIT('h2)
	) name31317 (
		_w18334_,
		_w35363_,
		_w35364_
	);
	LUT2 #(
		.INIT('h4)
	) name31318 (
		_w35362_,
		_w35364_,
		_w35365_
	);
	LUT2 #(
		.INIT('h1)
	) name31319 (
		_w35361_,
		_w35365_,
		_w35366_
	);
	LUT2 #(
		.INIT('h2)
	) name31320 (
		\bdma_BWRn_reg/NET0131 ,
		\bdma_WRlat_reg/P0001 ,
		_w35367_
	);
	LUT2 #(
		.INIT('h1)
	) name31321 (
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		_w35368_
	);
	LUT2 #(
		.INIT('h2)
	) name31322 (
		\bdma_BCTL_reg[6]/NET0131 ,
		_w35368_,
		_w35369_
	);
	LUT2 #(
		.INIT('h8)
	) name31323 (
		\bdma_BCTL_reg[7]/NET0131 ,
		_w35369_,
		_w35370_
	);
	LUT2 #(
		.INIT('h2)
	) name31324 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w35370_,
		_w35371_
	);
	LUT2 #(
		.INIT('h4)
	) name31325 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w35370_,
		_w35372_
	);
	LUT2 #(
		.INIT('h4)
	) name31326 (
		\bdma_BCTL_reg[6]/NET0131 ,
		_w35368_,
		_w35373_
	);
	LUT2 #(
		.INIT('h1)
	) name31327 (
		_w35369_,
		_w35373_,
		_w35374_
	);
	LUT2 #(
		.INIT('h2)
	) name31328 (
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w35374_,
		_w35375_
	);
	LUT2 #(
		.INIT('h4)
	) name31329 (
		\bdma_BWcnt_reg[2]/NET0131 ,
		_w35374_,
		_w35376_
	);
	LUT2 #(
		.INIT('h1)
	) name31330 (
		\bdma_BCTL_reg[7]/NET0131 ,
		_w35369_,
		_w35377_
	);
	LUT2 #(
		.INIT('h1)
	) name31331 (
		\bdma_BWcnt_reg[4]/NET0131 ,
		_w35377_,
		_w35378_
	);
	LUT2 #(
		.INIT('h2)
	) name31332 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w35378_,
		_w35379_
	);
	LUT2 #(
		.INIT('h4)
	) name31333 (
		\bdma_BWcnt_reg[3]/NET0131 ,
		_w35378_,
		_w35380_
	);
	LUT2 #(
		.INIT('h8)
	) name31334 (
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BCTL_reg[5]/NET0131 ,
		_w35381_
	);
	LUT2 #(
		.INIT('h1)
	) name31335 (
		_w35368_,
		_w35381_,
		_w35382_
	);
	LUT2 #(
		.INIT('h8)
	) name31336 (
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w35382_,
		_w35383_
	);
	LUT2 #(
		.INIT('h1)
	) name31337 (
		\bdma_BWcnt_reg[1]/NET0131 ,
		_w35382_,
		_w35384_
	);
	LUT2 #(
		.INIT('h1)
	) name31338 (
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w35385_
	);
	LUT2 #(
		.INIT('h8)
	) name31339 (
		\bdma_BCTL_reg[4]/NET0131 ,
		\bdma_BWcnt_reg[0]/NET0131 ,
		_w35386_
	);
	LUT2 #(
		.INIT('h2)
	) name31340 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w35385_,
		_w35387_
	);
	LUT2 #(
		.INIT('h4)
	) name31341 (
		_w35386_,
		_w35387_,
		_w35388_
	);
	LUT2 #(
		.INIT('h4)
	) name31342 (
		_w35383_,
		_w35388_,
		_w35389_
	);
	LUT2 #(
		.INIT('h4)
	) name31343 (
		_w35384_,
		_w35389_,
		_w35390_
	);
	LUT2 #(
		.INIT('h1)
	) name31344 (
		_w35371_,
		_w35372_,
		_w35391_
	);
	LUT2 #(
		.INIT('h1)
	) name31345 (
		_w35375_,
		_w35376_,
		_w35392_
	);
	LUT2 #(
		.INIT('h8)
	) name31346 (
		_w35391_,
		_w35392_,
		_w35393_
	);
	LUT2 #(
		.INIT('h4)
	) name31347 (
		_w35379_,
		_w35390_,
		_w35394_
	);
	LUT2 #(
		.INIT('h4)
	) name31348 (
		_w35380_,
		_w35394_,
		_w35395_
	);
	LUT2 #(
		.INIT('h8)
	) name31349 (
		_w35393_,
		_w35395_,
		_w35396_
	);
	LUT2 #(
		.INIT('h1)
	) name31350 (
		_w35367_,
		_w35396_,
		_w35397_
	);
	LUT2 #(
		.INIT('h4)
	) name31351 (
		\sport0_rxctl_RXSHT_reg[11]/P0001 ,
		_w20868_,
		_w35398_
	);
	LUT2 #(
		.INIT('h8)
	) name31352 (
		\sport0_rxctl_RX_reg[11]/P0001 ,
		_w20873_,
		_w35399_
	);
	LUT2 #(
		.INIT('h1)
	) name31353 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w34401_,
		_w35400_
	);
	LUT2 #(
		.INIT('h2)
	) name31354 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w31046_,
		_w35401_
	);
	LUT2 #(
		.INIT('h1)
	) name31355 (
		_w35400_,
		_w35401_,
		_w35402_
	);
	LUT2 #(
		.INIT('h8)
	) name31356 (
		_w31044_,
		_w35402_,
		_w35403_
	);
	LUT2 #(
		.INIT('h1)
	) name31357 (
		_w31044_,
		_w35402_,
		_w35404_
	);
	LUT2 #(
		.INIT('h2)
	) name31358 (
		_w20875_,
		_w35403_,
		_w35405_
	);
	LUT2 #(
		.INIT('h4)
	) name31359 (
		_w35404_,
		_w35405_,
		_w35406_
	);
	LUT2 #(
		.INIT('h4)
	) name31360 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w8460_,
		_w35407_
	);
	LUT2 #(
		.INIT('h1)
	) name31361 (
		_w20868_,
		_w35399_,
		_w35408_
	);
	LUT2 #(
		.INIT('h4)
	) name31362 (
		_w35407_,
		_w35408_,
		_w35409_
	);
	LUT2 #(
		.INIT('h4)
	) name31363 (
		_w35406_,
		_w35409_,
		_w35410_
	);
	LUT2 #(
		.INIT('h1)
	) name31364 (
		_w20871_,
		_w35398_,
		_w35411_
	);
	LUT2 #(
		.INIT('h4)
	) name31365 (
		_w35410_,
		_w35411_,
		_w35412_
	);
	LUT2 #(
		.INIT('h8)
	) name31366 (
		\sport0_rxctl_RX_reg[11]/P0001 ,
		_w20871_,
		_w35413_
	);
	LUT2 #(
		.INIT('h1)
	) name31367 (
		_w35412_,
		_w35413_,
		_w35414_
	);
	LUT2 #(
		.INIT('h1)
	) name31368 (
		IACKn_pad,
		_w20384_,
		_w35415_
	);
	LUT2 #(
		.INIT('h4)
	) name31369 (
		_w20821_,
		_w35415_,
		_w35416_
	);
	LUT2 #(
		.INIT('h2)
	) name31370 (
		_w32465_,
		_w35416_,
		_w35417_
	);
	LUT2 #(
		.INIT('h1)
	) name31371 (
		_w4117_,
		_w25009_,
		_w35418_
	);
	LUT2 #(
		.INIT('h4)
	) name31372 (
		_w32852_,
		_w35418_,
		_w35419_
	);
	LUT2 #(
		.INIT('h1)
	) name31373 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[9]/NET0131 ,
		_w35418_,
		_w35420_
	);
	LUT2 #(
		.INIT('h1)
	) name31374 (
		_w35419_,
		_w35420_,
		_w35421_
	);
	LUT2 #(
		.INIT('h4)
	) name31375 (
		_w32898_,
		_w35418_,
		_w35422_
	);
	LUT2 #(
		.INIT('h1)
	) name31376 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[8]/NET0131 ,
		_w35418_,
		_w35423_
	);
	LUT2 #(
		.INIT('h1)
	) name31377 (
		_w35422_,
		_w35423_,
		_w35424_
	);
	LUT2 #(
		.INIT('h4)
	) name31378 (
		_w32806_,
		_w35418_,
		_w35425_
	);
	LUT2 #(
		.INIT('h1)
	) name31379 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[7]/NET0131 ,
		_w35418_,
		_w35426_
	);
	LUT2 #(
		.INIT('h1)
	) name31380 (
		_w35425_,
		_w35426_,
		_w35427_
	);
	LUT2 #(
		.INIT('h4)
	) name31381 (
		_w32829_,
		_w35418_,
		_w35428_
	);
	LUT2 #(
		.INIT('h1)
	) name31382 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[6]/NET0131 ,
		_w35418_,
		_w35429_
	);
	LUT2 #(
		.INIT('h1)
	) name31383 (
		_w35428_,
		_w35429_,
		_w35430_
	);
	LUT2 #(
		.INIT('h4)
	) name31384 (
		_w32783_,
		_w35418_,
		_w35431_
	);
	LUT2 #(
		.INIT('h1)
	) name31385 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[5]/NET0131 ,
		_w35418_,
		_w35432_
	);
	LUT2 #(
		.INIT('h1)
	) name31386 (
		_w35431_,
		_w35432_,
		_w35433_
	);
	LUT2 #(
		.INIT('h4)
	) name31387 (
		_w10302_,
		_w32048_,
		_w35434_
	);
	LUT2 #(
		.INIT('h1)
	) name31388 (
		_w9752_,
		_w32048_,
		_w35435_
	);
	LUT2 #(
		.INIT('h2)
	) name31389 (
		_w32054_,
		_w35434_,
		_w35436_
	);
	LUT2 #(
		.INIT('h4)
	) name31390 (
		_w35435_,
		_w35436_,
		_w35437_
	);
	LUT2 #(
		.INIT('h4)
	) name31391 (
		_w9805_,
		_w32058_,
		_w35438_
	);
	LUT2 #(
		.INIT('h1)
	) name31392 (
		_w9767_,
		_w32048_,
		_w35439_
	);
	LUT2 #(
		.INIT('h1)
	) name31393 (
		_w9790_,
		_w35438_,
		_w35440_
	);
	LUT2 #(
		.INIT('h4)
	) name31394 (
		_w32054_,
		_w35440_,
		_w35441_
	);
	LUT2 #(
		.INIT('h4)
	) name31395 (
		_w35439_,
		_w35441_,
		_w35442_
	);
	LUT2 #(
		.INIT('h1)
	) name31396 (
		_w35437_,
		_w35442_,
		_w35443_
	);
	LUT2 #(
		.INIT('h1)
	) name31397 (
		_w32068_,
		_w35443_,
		_w35444_
	);
	LUT2 #(
		.INIT('h1)
	) name31398 (
		_w9733_,
		_w32048_,
		_w35445_
	);
	LUT2 #(
		.INIT('h4)
	) name31399 (
		_w9786_,
		_w32048_,
		_w35446_
	);
	LUT2 #(
		.INIT('h1)
	) name31400 (
		_w32054_,
		_w35445_,
		_w35447_
	);
	LUT2 #(
		.INIT('h4)
	) name31401 (
		_w35446_,
		_w35447_,
		_w35448_
	);
	LUT2 #(
		.INIT('h2)
	) name31402 (
		_w10289_,
		_w32048_,
		_w35449_
	);
	LUT2 #(
		.INIT('h8)
	) name31403 (
		_w10069_,
		_w32048_,
		_w35450_
	);
	LUT2 #(
		.INIT('h2)
	) name31404 (
		_w32054_,
		_w35449_,
		_w35451_
	);
	LUT2 #(
		.INIT('h4)
	) name31405 (
		_w35450_,
		_w35451_,
		_w35452_
	);
	LUT2 #(
		.INIT('h1)
	) name31406 (
		_w35448_,
		_w35452_,
		_w35453_
	);
	LUT2 #(
		.INIT('h2)
	) name31407 (
		_w32068_,
		_w35453_,
		_w35454_
	);
	LUT2 #(
		.INIT('h1)
	) name31408 (
		_w35444_,
		_w35454_,
		_w35455_
	);
	LUT2 #(
		.INIT('h2)
	) name31409 (
		_w35418_,
		_w35455_,
		_w35456_
	);
	LUT2 #(
		.INIT('h1)
	) name31410 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[4]/NET0131 ,
		_w35418_,
		_w35457_
	);
	LUT2 #(
		.INIT('h1)
	) name31411 (
		_w35456_,
		_w35457_,
		_w35458_
	);
	LUT2 #(
		.INIT('h1)
	) name31412 (
		_w7644_,
		_w32048_,
		_w35459_
	);
	LUT2 #(
		.INIT('h4)
	) name31413 (
		_w8224_,
		_w32048_,
		_w35460_
	);
	LUT2 #(
		.INIT('h2)
	) name31414 (
		_w32054_,
		_w35459_,
		_w35461_
	);
	LUT2 #(
		.INIT('h4)
	) name31415 (
		_w35460_,
		_w35461_,
		_w35462_
	);
	LUT2 #(
		.INIT('h4)
	) name31416 (
		_w9666_,
		_w32058_,
		_w35463_
	);
	LUT2 #(
		.INIT('h1)
	) name31417 (
		_w9695_,
		_w32048_,
		_w35464_
	);
	LUT2 #(
		.INIT('h1)
	) name31418 (
		_w9700_,
		_w35463_,
		_w35465_
	);
	LUT2 #(
		.INIT('h4)
	) name31419 (
		_w32054_,
		_w35465_,
		_w35466_
	);
	LUT2 #(
		.INIT('h4)
	) name31420 (
		_w35464_,
		_w35466_,
		_w35467_
	);
	LUT2 #(
		.INIT('h1)
	) name31421 (
		_w35462_,
		_w35467_,
		_w35468_
	);
	LUT2 #(
		.INIT('h1)
	) name31422 (
		_w32068_,
		_w35468_,
		_w35469_
	);
	LUT2 #(
		.INIT('h1)
	) name31423 (
		_w8149_,
		_w32048_,
		_w35470_
	);
	LUT2 #(
		.INIT('h4)
	) name31424 (
		_w8190_,
		_w32048_,
		_w35471_
	);
	LUT2 #(
		.INIT('h1)
	) name31425 (
		_w32054_,
		_w35470_,
		_w35472_
	);
	LUT2 #(
		.INIT('h4)
	) name31426 (
		_w35471_,
		_w35472_,
		_w35473_
	);
	LUT2 #(
		.INIT('h2)
	) name31427 (
		_w7859_,
		_w32048_,
		_w35474_
	);
	LUT2 #(
		.INIT('h8)
	) name31428 (
		_w8113_,
		_w32048_,
		_w35475_
	);
	LUT2 #(
		.INIT('h2)
	) name31429 (
		_w32054_,
		_w35474_,
		_w35476_
	);
	LUT2 #(
		.INIT('h4)
	) name31430 (
		_w35475_,
		_w35476_,
		_w35477_
	);
	LUT2 #(
		.INIT('h1)
	) name31431 (
		_w35473_,
		_w35477_,
		_w35478_
	);
	LUT2 #(
		.INIT('h2)
	) name31432 (
		_w32068_,
		_w35478_,
		_w35479_
	);
	LUT2 #(
		.INIT('h1)
	) name31433 (
		_w35469_,
		_w35479_,
		_w35480_
	);
	LUT2 #(
		.INIT('h2)
	) name31434 (
		_w35418_,
		_w35480_,
		_w35481_
	);
	LUT2 #(
		.INIT('h1)
	) name31435 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[3]/NET0131 ,
		_w35418_,
		_w35482_
	);
	LUT2 #(
		.INIT('h1)
	) name31436 (
		_w35481_,
		_w35482_,
		_w35483_
	);
	LUT2 #(
		.INIT('h4)
	) name31437 (
		_w8794_,
		_w32048_,
		_w35484_
	);
	LUT2 #(
		.INIT('h1)
	) name31438 (
		_w8246_,
		_w32048_,
		_w35485_
	);
	LUT2 #(
		.INIT('h2)
	) name31439 (
		_w32054_,
		_w35484_,
		_w35486_
	);
	LUT2 #(
		.INIT('h4)
	) name31440 (
		_w35485_,
		_w35486_,
		_w35487_
	);
	LUT2 #(
		.INIT('h4)
	) name31441 (
		_w9600_,
		_w32058_,
		_w35488_
	);
	LUT2 #(
		.INIT('h1)
	) name31442 (
		_w9625_,
		_w32048_,
		_w35489_
	);
	LUT2 #(
		.INIT('h1)
	) name31443 (
		_w9633_,
		_w35488_,
		_w35490_
	);
	LUT2 #(
		.INIT('h4)
	) name31444 (
		_w32054_,
		_w35490_,
		_w35491_
	);
	LUT2 #(
		.INIT('h4)
	) name31445 (
		_w35489_,
		_w35491_,
		_w35492_
	);
	LUT2 #(
		.INIT('h1)
	) name31446 (
		_w35487_,
		_w35492_,
		_w35493_
	);
	LUT2 #(
		.INIT('h1)
	) name31447 (
		_w32068_,
		_w35493_,
		_w35494_
	);
	LUT2 #(
		.INIT('h1)
	) name31448 (
		_w8750_,
		_w32048_,
		_w35495_
	);
	LUT2 #(
		.INIT('h4)
	) name31449 (
		_w8773_,
		_w32048_,
		_w35496_
	);
	LUT2 #(
		.INIT('h1)
	) name31450 (
		_w32054_,
		_w35495_,
		_w35497_
	);
	LUT2 #(
		.INIT('h4)
	) name31451 (
		_w35496_,
		_w35497_,
		_w35498_
	);
	LUT2 #(
		.INIT('h2)
	) name31452 (
		_w8460_,
		_w32048_,
		_w35499_
	);
	LUT2 #(
		.INIT('h8)
	) name31453 (
		_w8715_,
		_w32048_,
		_w35500_
	);
	LUT2 #(
		.INIT('h2)
	) name31454 (
		_w32054_,
		_w35499_,
		_w35501_
	);
	LUT2 #(
		.INIT('h4)
	) name31455 (
		_w35500_,
		_w35501_,
		_w35502_
	);
	LUT2 #(
		.INIT('h1)
	) name31456 (
		_w35498_,
		_w35502_,
		_w35503_
	);
	LUT2 #(
		.INIT('h2)
	) name31457 (
		_w32068_,
		_w35503_,
		_w35504_
	);
	LUT2 #(
		.INIT('h1)
	) name31458 (
		_w35494_,
		_w35504_,
		_w35505_
	);
	LUT2 #(
		.INIT('h2)
	) name31459 (
		_w35418_,
		_w35505_,
		_w35506_
	);
	LUT2 #(
		.INIT('h1)
	) name31460 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[2]/NET0131 ,
		_w35418_,
		_w35507_
	);
	LUT2 #(
		.INIT('h1)
	) name31461 (
		_w35506_,
		_w35507_,
		_w35508_
	);
	LUT2 #(
		.INIT('h4)
	) name31462 (
		_w8926_,
		_w32048_,
		_w35509_
	);
	LUT2 #(
		.INIT('h1)
	) name31463 (
		_w8962_,
		_w32048_,
		_w35510_
	);
	LUT2 #(
		.INIT('h2)
	) name31464 (
		_w32054_,
		_w35509_,
		_w35511_
	);
	LUT2 #(
		.INIT('h4)
	) name31465 (
		_w35510_,
		_w35511_,
		_w35512_
	);
	LUT2 #(
		.INIT('h4)
	) name31466 (
		_w9528_,
		_w32058_,
		_w35513_
	);
	LUT2 #(
		.INIT('h1)
	) name31467 (
		_w9559_,
		_w32048_,
		_w35514_
	);
	LUT2 #(
		.INIT('h1)
	) name31468 (
		_w9567_,
		_w35513_,
		_w35515_
	);
	LUT2 #(
		.INIT('h4)
	) name31469 (
		_w32054_,
		_w35515_,
		_w35516_
	);
	LUT2 #(
		.INIT('h4)
	) name31470 (
		_w35514_,
		_w35516_,
		_w35517_
	);
	LUT2 #(
		.INIT('h1)
	) name31471 (
		_w35512_,
		_w35517_,
		_w35518_
	);
	LUT2 #(
		.INIT('h1)
	) name31472 (
		_w32068_,
		_w35518_,
		_w35519_
	);
	LUT2 #(
		.INIT('h1)
	) name31473 (
		_w8873_,
		_w32048_,
		_w35520_
	);
	LUT2 #(
		.INIT('h4)
	) name31474 (
		_w8903_,
		_w32048_,
		_w35521_
	);
	LUT2 #(
		.INIT('h1)
	) name31475 (
		_w32054_,
		_w35520_,
		_w35522_
	);
	LUT2 #(
		.INIT('h4)
	) name31476 (
		_w35521_,
		_w35522_,
		_w35523_
	);
	LUT2 #(
		.INIT('h2)
	) name31477 (
		_w9178_,
		_w32048_,
		_w35524_
	);
	LUT2 #(
		.INIT('h8)
	) name31478 (
		_w9435_,
		_w32048_,
		_w35525_
	);
	LUT2 #(
		.INIT('h2)
	) name31479 (
		_w32054_,
		_w35524_,
		_w35526_
	);
	LUT2 #(
		.INIT('h4)
	) name31480 (
		_w35525_,
		_w35526_,
		_w35527_
	);
	LUT2 #(
		.INIT('h1)
	) name31481 (
		_w35523_,
		_w35527_,
		_w35528_
	);
	LUT2 #(
		.INIT('h2)
	) name31482 (
		_w32068_,
		_w35528_,
		_w35529_
	);
	LUT2 #(
		.INIT('h1)
	) name31483 (
		_w35519_,
		_w35529_,
		_w35530_
	);
	LUT2 #(
		.INIT('h2)
	) name31484 (
		_w35418_,
		_w35530_,
		_w35531_
	);
	LUT2 #(
		.INIT('h1)
	) name31485 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[1]/NET0131 ,
		_w35418_,
		_w35532_
	);
	LUT2 #(
		.INIT('h1)
	) name31486 (
		_w35531_,
		_w35532_,
		_w35533_
	);
	LUT2 #(
		.INIT('h2)
	) name31487 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[13]/NET0131 ,
		_w35418_,
		_w35534_
	);
	LUT2 #(
		.INIT('h4)
	) name31488 (
		_w32080_,
		_w35418_,
		_w35535_
	);
	LUT2 #(
		.INIT('h1)
	) name31489 (
		_w35534_,
		_w35535_,
		_w35536_
	);
	LUT2 #(
		.INIT('h4)
	) name31490 (
		_w32921_,
		_w35418_,
		_w35537_
	);
	LUT2 #(
		.INIT('h1)
	) name31491 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[12]/NET0131 ,
		_w35418_,
		_w35538_
	);
	LUT2 #(
		.INIT('h1)
	) name31492 (
		_w35537_,
		_w35538_,
		_w35539_
	);
	LUT2 #(
		.INIT('h4)
	) name31493 (
		_w32944_,
		_w35418_,
		_w35540_
	);
	LUT2 #(
		.INIT('h1)
	) name31494 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w35418_,
		_w35541_
	);
	LUT2 #(
		.INIT('h1)
	) name31495 (
		_w35540_,
		_w35541_,
		_w35542_
	);
	LUT2 #(
		.INIT('h4)
	) name31496 (
		_w32875_,
		_w35418_,
		_w35543_
	);
	LUT2 #(
		.INIT('h1)
	) name31497 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[10]/NET0131 ,
		_w35418_,
		_w35544_
	);
	LUT2 #(
		.INIT('h1)
	) name31498 (
		_w35543_,
		_w35544_,
		_w35545_
	);
	LUT2 #(
		.INIT('h1)
	) name31499 (
		_w6546_,
		_w32048_,
		_w35546_
	);
	LUT2 #(
		.INIT('h4)
	) name31500 (
		_w7622_,
		_w32048_,
		_w35547_
	);
	LUT2 #(
		.INIT('h2)
	) name31501 (
		_w32054_,
		_w35546_,
		_w35548_
	);
	LUT2 #(
		.INIT('h4)
	) name31502 (
		_w35547_,
		_w35548_,
		_w35549_
	);
	LUT2 #(
		.INIT('h1)
	) name31503 (
		_w6911_,
		_w32048_,
		_w35550_
	);
	LUT2 #(
		.INIT('h4)
	) name31504 (
		_w6980_,
		_w32058_,
		_w35551_
	);
	LUT2 #(
		.INIT('h1)
	) name31505 (
		_w6957_,
		_w35551_,
		_w35552_
	);
	LUT2 #(
		.INIT('h4)
	) name31506 (
		_w32054_,
		_w35552_,
		_w35553_
	);
	LUT2 #(
		.INIT('h4)
	) name31507 (
		_w35550_,
		_w35553_,
		_w35554_
	);
	LUT2 #(
		.INIT('h1)
	) name31508 (
		_w35549_,
		_w35554_,
		_w35555_
	);
	LUT2 #(
		.INIT('h1)
	) name31509 (
		_w32068_,
		_w35555_,
		_w35556_
	);
	LUT2 #(
		.INIT('h1)
	) name31510 (
		_w6158_,
		_w32048_,
		_w35557_
	);
	LUT2 #(
		.INIT('h4)
	) name31511 (
		_w6951_,
		_w32048_,
		_w35558_
	);
	LUT2 #(
		.INIT('h1)
	) name31512 (
		_w32054_,
		_w35557_,
		_w35559_
	);
	LUT2 #(
		.INIT('h4)
	) name31513 (
		_w35558_,
		_w35559_,
		_w35560_
	);
	LUT2 #(
		.INIT('h2)
	) name31514 (
		_w7340_,
		_w32048_,
		_w35561_
	);
	LUT2 #(
		.INIT('h8)
	) name31515 (
		_w7607_,
		_w32048_,
		_w35562_
	);
	LUT2 #(
		.INIT('h2)
	) name31516 (
		_w32054_,
		_w35561_,
		_w35563_
	);
	LUT2 #(
		.INIT('h4)
	) name31517 (
		_w35562_,
		_w35563_,
		_w35564_
	);
	LUT2 #(
		.INIT('h1)
	) name31518 (
		_w35560_,
		_w35564_,
		_w35565_
	);
	LUT2 #(
		.INIT('h2)
	) name31519 (
		_w32068_,
		_w35565_,
		_w35566_
	);
	LUT2 #(
		.INIT('h1)
	) name31520 (
		_w35556_,
		_w35566_,
		_w35567_
	);
	LUT2 #(
		.INIT('h2)
	) name31521 (
		_w35418_,
		_w35567_,
		_w35568_
	);
	LUT2 #(
		.INIT('h1)
	) name31522 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[0]/NET0131 ,
		_w35418_,
		_w35569_
	);
	LUT2 #(
		.INIT('h1)
	) name31523 (
		_w35568_,
		_w35569_,
		_w35570_
	);
	LUT2 #(
		.INIT('h8)
	) name31524 (
		\core_c_dec_MTMSTAT_Eg_reg/P0001 ,
		_w4118_,
		_w35571_
	);
	LUT2 #(
		.INIT('h8)
	) name31525 (
		_w23231_,
		_w32022_,
		_w35572_
	);
	LUT2 #(
		.INIT('h8)
	) name31526 (
		_w31998_,
		_w35572_,
		_w35573_
	);
	LUT2 #(
		.INIT('h1)
	) name31527 (
		_w35571_,
		_w35573_,
		_w35574_
	);
	LUT2 #(
		.INIT('h1)
	) name31528 (
		\bdma_BEAD_reg[7]/NET0131 ,
		_w33308_,
		_w35575_
	);
	LUT2 #(
		.INIT('h1)
	) name31529 (
		_w20765_,
		_w33309_,
		_w35576_
	);
	LUT2 #(
		.INIT('h4)
	) name31530 (
		_w35575_,
		_w35576_,
		_w35577_
	);
	LUT2 #(
		.INIT('h8)
	) name31531 (
		_w11265_,
		_w20765_,
		_w35578_
	);
	LUT2 #(
		.INIT('h1)
	) name31532 (
		_w35577_,
		_w35578_,
		_w35579_
	);
	LUT2 #(
		.INIT('h1)
	) name31533 (
		\bdma_BEAD_reg[6]/NET0131 ,
		_w33307_,
		_w35580_
	);
	LUT2 #(
		.INIT('h1)
	) name31534 (
		_w20765_,
		_w33308_,
		_w35581_
	);
	LUT2 #(
		.INIT('h4)
	) name31535 (
		_w35580_,
		_w35581_,
		_w35582_
	);
	LUT2 #(
		.INIT('h8)
	) name31536 (
		_w11525_,
		_w20765_,
		_w35583_
	);
	LUT2 #(
		.INIT('h1)
	) name31537 (
		_w35582_,
		_w35583_,
		_w35584_
	);
	LUT2 #(
		.INIT('h1)
	) name31538 (
		\bdma_BEAD_reg[5]/NET0131 ,
		_w33306_,
		_w35585_
	);
	LUT2 #(
		.INIT('h1)
	) name31539 (
		_w20765_,
		_w33307_,
		_w35586_
	);
	LUT2 #(
		.INIT('h4)
	) name31540 (
		_w35585_,
		_w35586_,
		_w35587_
	);
	LUT2 #(
		.INIT('h8)
	) name31541 (
		_w10911_,
		_w20765_,
		_w35588_
	);
	LUT2 #(
		.INIT('h1)
	) name31542 (
		_w35587_,
		_w35588_,
		_w35589_
	);
	LUT2 #(
		.INIT('h8)
	) name31543 (
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w28786_,
		_w35590_
	);
	LUT2 #(
		.INIT('h1)
	) name31544 (
		\sport1_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport1_cfg_SP_ENg_reg/NET0131 ,
		_w35591_
	);
	LUT2 #(
		.INIT('h1)
	) name31545 (
		_w28856_,
		_w35591_,
		_w35592_
	);
	LUT2 #(
		.INIT('h8)
	) name31546 (
		_w28855_,
		_w35592_,
		_w35593_
	);
	LUT2 #(
		.INIT('h1)
	) name31547 (
		_w35590_,
		_w35593_,
		_w35594_
	);
	LUT2 #(
		.INIT('h8)
	) name31548 (
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w28876_,
		_w35595_
	);
	LUT2 #(
		.INIT('h1)
	) name31549 (
		\sport0_cfg_FSi_cnt_reg[0]/NET0131 ,
		\sport0_cfg_SP_ENg_reg/NET0131 ,
		_w35596_
	);
	LUT2 #(
		.INIT('h1)
	) name31550 (
		_w28946_,
		_w35596_,
		_w35597_
	);
	LUT2 #(
		.INIT('h8)
	) name31551 (
		_w28945_,
		_w35597_,
		_w35598_
	);
	LUT2 #(
		.INIT('h1)
	) name31552 (
		_w35595_,
		_w35598_,
		_w35599_
	);
	LUT2 #(
		.INIT('h2)
	) name31553 (
		_w14752_,
		_w25088_,
		_w35600_
	);
	LUT2 #(
		.INIT('h1)
	) name31554 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 ,
		_w17799_,
		_w35601_
	);
	LUT2 #(
		.INIT('h4)
	) name31555 (
		_w17809_,
		_w19559_,
		_w35602_
	);
	LUT2 #(
		.INIT('h2)
	) name31556 (
		_w17811_,
		_w35602_,
		_w35603_
	);
	LUT2 #(
		.INIT('h1)
	) name31557 (
		_w35601_,
		_w35603_,
		_w35604_
	);
	LUT2 #(
		.INIT('h1)
	) name31558 (
		_w17823_,
		_w35604_,
		_w35605_
	);
	LUT2 #(
		.INIT('h1)
	) name31559 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[0]/P0001 ,
		_w17808_,
		_w35606_
	);
	LUT2 #(
		.INIT('h1)
	) name31560 (
		_w35605_,
		_w35606_,
		_w35607_
	);
	LUT2 #(
		.INIT('h2)
	) name31561 (
		_w17829_,
		_w35607_,
		_w35608_
	);
	LUT2 #(
		.INIT('h1)
	) name31562 (
		_w35600_,
		_w35608_,
		_w35609_
	);
	LUT2 #(
		.INIT('h1)
	) name31563 (
		\sice_ICYC_reg[23]/NET0131 ,
		_w20785_,
		_w35610_
	);
	LUT2 #(
		.INIT('h1)
	) name31564 (
		_w32035_,
		_w35610_,
		_w35611_
	);
	LUT2 #(
		.INIT('h8)
	) name31565 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w4118_,
		_w35612_
	);
	LUT2 #(
		.INIT('h8)
	) name31566 (
		_w23231_,
		_w32010_,
		_w35613_
	);
	LUT2 #(
		.INIT('h1)
	) name31567 (
		_w35612_,
		_w35613_,
		_w35614_
	);
	LUT2 #(
		.INIT('h8)
	) name31568 (
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w28876_,
		_w35615_
	);
	LUT2 #(
		.INIT('h1)
	) name31569 (
		\sport0_cfg_FSi_cnt_reg[1]/NET0131 ,
		_w28946_,
		_w35616_
	);
	LUT2 #(
		.INIT('h1)
	) name31570 (
		_w28947_,
		_w35616_,
		_w35617_
	);
	LUT2 #(
		.INIT('h8)
	) name31571 (
		_w28945_,
		_w35617_,
		_w35618_
	);
	LUT2 #(
		.INIT('h1)
	) name31572 (
		_w35615_,
		_w35618_,
		_w35619_
	);
	LUT2 #(
		.INIT('h8)
	) name31573 (
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w28786_,
		_w35620_
	);
	LUT2 #(
		.INIT('h1)
	) name31574 (
		\sport1_cfg_FSi_cnt_reg[1]/NET0131 ,
		_w28856_,
		_w35621_
	);
	LUT2 #(
		.INIT('h1)
	) name31575 (
		_w28857_,
		_w35621_,
		_w35622_
	);
	LUT2 #(
		.INIT('h8)
	) name31576 (
		_w28855_,
		_w35622_,
		_w35623_
	);
	LUT2 #(
		.INIT('h1)
	) name31577 (
		_w35620_,
		_w35623_,
		_w35624_
	);
	LUT2 #(
		.INIT('h8)
	) name31578 (
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w28786_,
		_w35625_
	);
	LUT2 #(
		.INIT('h1)
	) name31579 (
		\sport1_cfg_FSi_cnt_reg[2]/NET0131 ,
		_w28857_,
		_w35626_
	);
	LUT2 #(
		.INIT('h1)
	) name31580 (
		_w28858_,
		_w35626_,
		_w35627_
	);
	LUT2 #(
		.INIT('h8)
	) name31581 (
		_w28855_,
		_w35627_,
		_w35628_
	);
	LUT2 #(
		.INIT('h1)
	) name31582 (
		_w35625_,
		_w35628_,
		_w35629_
	);
	LUT2 #(
		.INIT('h8)
	) name31583 (
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w28786_,
		_w35630_
	);
	LUT2 #(
		.INIT('h1)
	) name31584 (
		\sport1_cfg_FSi_cnt_reg[5]/NET0131 ,
		_w28860_,
		_w35631_
	);
	LUT2 #(
		.INIT('h1)
	) name31585 (
		_w28861_,
		_w35631_,
		_w35632_
	);
	LUT2 #(
		.INIT('h8)
	) name31586 (
		_w28855_,
		_w35632_,
		_w35633_
	);
	LUT2 #(
		.INIT('h1)
	) name31587 (
		_w35630_,
		_w35633_,
		_w35634_
	);
	LUT2 #(
		.INIT('h8)
	) name31588 (
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w28786_,
		_w35635_
	);
	LUT2 #(
		.INIT('h1)
	) name31589 (
		\sport1_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w28864_,
		_w35636_
	);
	LUT2 #(
		.INIT('h2)
	) name31590 (
		_w28855_,
		_w28865_,
		_w35637_
	);
	LUT2 #(
		.INIT('h4)
	) name31591 (
		_w35636_,
		_w35637_,
		_w35638_
	);
	LUT2 #(
		.INIT('h1)
	) name31592 (
		_w35635_,
		_w35638_,
		_w35639_
	);
	LUT2 #(
		.INIT('h8)
	) name31593 (
		\sport0_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w28876_,
		_w35640_
	);
	LUT2 #(
		.INIT('h1)
	) name31594 (
		\sport0_cfg_FSi_cnt_reg[13]/NET0131 ,
		_w28958_,
		_w35641_
	);
	LUT2 #(
		.INIT('h2)
	) name31595 (
		_w28945_,
		_w28959_,
		_w35642_
	);
	LUT2 #(
		.INIT('h4)
	) name31596 (
		_w35641_,
		_w35642_,
		_w35643_
	);
	LUT2 #(
		.INIT('h1)
	) name31597 (
		_w35640_,
		_w35643_,
		_w35644_
	);
	LUT2 #(
		.INIT('h8)
	) name31598 (
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w28876_,
		_w35645_
	);
	LUT2 #(
		.INIT('h1)
	) name31599 (
		\sport0_cfg_FSi_cnt_reg[2]/NET0131 ,
		_w28947_,
		_w35646_
	);
	LUT2 #(
		.INIT('h1)
	) name31600 (
		_w28948_,
		_w35646_,
		_w35647_
	);
	LUT2 #(
		.INIT('h8)
	) name31601 (
		_w28945_,
		_w35647_,
		_w35648_
	);
	LUT2 #(
		.INIT('h1)
	) name31602 (
		_w35645_,
		_w35648_,
		_w35649_
	);
	LUT2 #(
		.INIT('h8)
	) name31603 (
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w28876_,
		_w35650_
	);
	LUT2 #(
		.INIT('h1)
	) name31604 (
		\sport0_cfg_FSi_cnt_reg[5]/NET0131 ,
		_w28950_,
		_w35651_
	);
	LUT2 #(
		.INIT('h1)
	) name31605 (
		_w28951_,
		_w35651_,
		_w35652_
	);
	LUT2 #(
		.INIT('h8)
	) name31606 (
		_w28945_,
		_w35652_,
		_w35653_
	);
	LUT2 #(
		.INIT('h1)
	) name31607 (
		_w35650_,
		_w35653_,
		_w35654_
	);
	LUT2 #(
		.INIT('h1)
	) name31608 (
		\sice_ICYC_reg[4]/NET0131 ,
		_w18858_,
		_w35655_
	);
	LUT2 #(
		.INIT('h1)
	) name31609 (
		_w18859_,
		_w35655_,
		_w35656_
	);
	LUT2 #(
		.INIT('h8)
	) name31610 (
		\sport0_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w28876_,
		_w35657_
	);
	LUT2 #(
		.INIT('h1)
	) name31611 (
		\sport0_cfg_FSi_cnt_reg[9]/NET0131 ,
		_w28954_,
		_w35658_
	);
	LUT2 #(
		.INIT('h2)
	) name31612 (
		_w28945_,
		_w28955_,
		_w35659_
	);
	LUT2 #(
		.INIT('h4)
	) name31613 (
		_w35658_,
		_w35659_,
		_w35660_
	);
	LUT2 #(
		.INIT('h1)
	) name31614 (
		_w35657_,
		_w35660_,
		_w35661_
	);
	LUT2 #(
		.INIT('h1)
	) name31615 (
		\clkc_oscntr_reg_DO_reg[4]/NET0131 ,
		_w23417_,
		_w35662_
	);
	LUT2 #(
		.INIT('h1)
	) name31616 (
		_w23418_,
		_w35662_,
		_w35663_
	);
	LUT2 #(
		.INIT('h1)
	) name31617 (
		\sice_IIRC_reg[4]/NET0131 ,
		_w18867_,
		_w35664_
	);
	LUT2 #(
		.INIT('h1)
	) name31618 (
		_w18868_,
		_w35664_,
		_w35665_
	);
	LUT2 #(
		.INIT('h8)
	) name31619 (
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w28786_,
		_w35666_
	);
	LUT2 #(
		.INIT('h1)
	) name31620 (
		\sport1_cfg_FSi_cnt_reg[13]/NET0131 ,
		_w28868_,
		_w35667_
	);
	LUT2 #(
		.INIT('h2)
	) name31621 (
		_w28855_,
		_w28869_,
		_w35668_
	);
	LUT2 #(
		.INIT('h4)
	) name31622 (
		_w35667_,
		_w35668_,
		_w35669_
	);
	LUT2 #(
		.INIT('h1)
	) name31623 (
		_w35666_,
		_w35669_,
		_w35670_
	);
	LUT2 #(
		.INIT('h8)
	) name31624 (
		_w26967_,
		_w34841_,
		_w35671_
	);
	LUT2 #(
		.INIT('h2)
	) name31625 (
		\sice_IRR_reg[4]/P0001 ,
		_w35671_,
		_w35672_
	);
	LUT2 #(
		.INIT('h8)
	) name31626 (
		\sice_SPC_reg[14]/P0001 ,
		_w35671_,
		_w35673_
	);
	LUT2 #(
		.INIT('h1)
	) name31627 (
		_w35672_,
		_w35673_,
		_w35674_
	);
	LUT2 #(
		.INIT('h2)
	) name31628 (
		_w4093_,
		_w35674_,
		_w35675_
	);
	LUT2 #(
		.INIT('h2)
	) name31629 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		_w4093_,
		_w35676_
	);
	LUT2 #(
		.INIT('h1)
	) name31630 (
		_w35675_,
		_w35676_,
		_w35677_
	);
	LUT2 #(
		.INIT('h2)
	) name31631 (
		\sice_IRR_reg[9]/P0001 ,
		_w35671_,
		_w35678_
	);
	LUT2 #(
		.INIT('h8)
	) name31632 (
		\sice_SPC_reg[19]/P0001 ,
		_w35671_,
		_w35679_
	);
	LUT2 #(
		.INIT('h1)
	) name31633 (
		_w35678_,
		_w35679_,
		_w35680_
	);
	LUT2 #(
		.INIT('h2)
	) name31634 (
		_w4093_,
		_w35680_,
		_w35681_
	);
	LUT2 #(
		.INIT('h2)
	) name31635 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		_w4093_,
		_w35682_
	);
	LUT2 #(
		.INIT('h1)
	) name31636 (
		_w35681_,
		_w35682_,
		_w35683_
	);
	LUT2 #(
		.INIT('h2)
	) name31637 (
		\sice_IRR_reg[8]/P0001 ,
		_w35671_,
		_w35684_
	);
	LUT2 #(
		.INIT('h8)
	) name31638 (
		\sice_SPC_reg[18]/P0001 ,
		_w35671_,
		_w35685_
	);
	LUT2 #(
		.INIT('h1)
	) name31639 (
		_w35684_,
		_w35685_,
		_w35686_
	);
	LUT2 #(
		.INIT('h2)
	) name31640 (
		_w4093_,
		_w35686_,
		_w35687_
	);
	LUT2 #(
		.INIT('h2)
	) name31641 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		_w4093_,
		_w35688_
	);
	LUT2 #(
		.INIT('h1)
	) name31642 (
		_w35687_,
		_w35688_,
		_w35689_
	);
	LUT2 #(
		.INIT('h2)
	) name31643 (
		\sice_IRR_reg[7]/P0001 ,
		_w35671_,
		_w35690_
	);
	LUT2 #(
		.INIT('h8)
	) name31644 (
		\sice_SPC_reg[17]/P0001 ,
		_w35671_,
		_w35691_
	);
	LUT2 #(
		.INIT('h1)
	) name31645 (
		_w35690_,
		_w35691_,
		_w35692_
	);
	LUT2 #(
		.INIT('h2)
	) name31646 (
		_w4093_,
		_w35692_,
		_w35693_
	);
	LUT2 #(
		.INIT('h2)
	) name31647 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		_w4093_,
		_w35694_
	);
	LUT2 #(
		.INIT('h1)
	) name31648 (
		_w35693_,
		_w35694_,
		_w35695_
	);
	LUT2 #(
		.INIT('h2)
	) name31649 (
		\sice_IRR_reg[6]/P0001 ,
		_w35671_,
		_w35696_
	);
	LUT2 #(
		.INIT('h8)
	) name31650 (
		\sice_SPC_reg[16]/P0001 ,
		_w35671_,
		_w35697_
	);
	LUT2 #(
		.INIT('h1)
	) name31651 (
		_w35696_,
		_w35697_,
		_w35698_
	);
	LUT2 #(
		.INIT('h2)
	) name31652 (
		_w4093_,
		_w35698_,
		_w35699_
	);
	LUT2 #(
		.INIT('h2)
	) name31653 (
		\core_c_psq_EXA_reg[6]/P0001 ,
		_w4093_,
		_w35700_
	);
	LUT2 #(
		.INIT('h1)
	) name31654 (
		_w35699_,
		_w35700_,
		_w35701_
	);
	LUT2 #(
		.INIT('h2)
	) name31655 (
		\sice_IRR_reg[5]/P0001 ,
		_w35671_,
		_w35702_
	);
	LUT2 #(
		.INIT('h8)
	) name31656 (
		\sice_SPC_reg[15]/P0001 ,
		_w35671_,
		_w35703_
	);
	LUT2 #(
		.INIT('h1)
	) name31657 (
		_w35702_,
		_w35703_,
		_w35704_
	);
	LUT2 #(
		.INIT('h2)
	) name31658 (
		_w4093_,
		_w35704_,
		_w35705_
	);
	LUT2 #(
		.INIT('h2)
	) name31659 (
		\core_c_psq_EXA_reg[5]/P0001 ,
		_w4093_,
		_w35706_
	);
	LUT2 #(
		.INIT('h1)
	) name31660 (
		_w35705_,
		_w35706_,
		_w35707_
	);
	LUT2 #(
		.INIT('h2)
	) name31661 (
		\sice_IRR_reg[3]/P0001 ,
		_w35671_,
		_w35708_
	);
	LUT2 #(
		.INIT('h8)
	) name31662 (
		\sice_SPC_reg[13]/P0001 ,
		_w35671_,
		_w35709_
	);
	LUT2 #(
		.INIT('h1)
	) name31663 (
		_w35708_,
		_w35709_,
		_w35710_
	);
	LUT2 #(
		.INIT('h2)
	) name31664 (
		_w4093_,
		_w35710_,
		_w35711_
	);
	LUT2 #(
		.INIT('h2)
	) name31665 (
		\core_c_psq_EXA_reg[3]/P0001 ,
		_w4093_,
		_w35712_
	);
	LUT2 #(
		.INIT('h1)
	) name31666 (
		_w35711_,
		_w35712_,
		_w35713_
	);
	LUT2 #(
		.INIT('h2)
	) name31667 (
		\sice_IRR_reg[2]/P0001 ,
		_w35671_,
		_w35714_
	);
	LUT2 #(
		.INIT('h8)
	) name31668 (
		\sice_SPC_reg[12]/P0001 ,
		_w35671_,
		_w35715_
	);
	LUT2 #(
		.INIT('h1)
	) name31669 (
		_w35714_,
		_w35715_,
		_w35716_
	);
	LUT2 #(
		.INIT('h2)
	) name31670 (
		_w4093_,
		_w35716_,
		_w35717_
	);
	LUT2 #(
		.INIT('h2)
	) name31671 (
		\core_c_psq_EXA_reg[2]/P0001 ,
		_w4093_,
		_w35718_
	);
	LUT2 #(
		.INIT('h1)
	) name31672 (
		_w35717_,
		_w35718_,
		_w35719_
	);
	LUT2 #(
		.INIT('h2)
	) name31673 (
		\sice_IRR_reg[13]/P0001 ,
		_w35671_,
		_w35720_
	);
	LUT2 #(
		.INIT('h8)
	) name31674 (
		\sice_SPC_reg[23]/P0001 ,
		_w35671_,
		_w35721_
	);
	LUT2 #(
		.INIT('h1)
	) name31675 (
		_w35720_,
		_w35721_,
		_w35722_
	);
	LUT2 #(
		.INIT('h2)
	) name31676 (
		_w4093_,
		_w35722_,
		_w35723_
	);
	LUT2 #(
		.INIT('h2)
	) name31677 (
		\core_c_psq_EXA_reg[13]/P0001 ,
		_w4093_,
		_w35724_
	);
	LUT2 #(
		.INIT('h1)
	) name31678 (
		_w35723_,
		_w35724_,
		_w35725_
	);
	LUT2 #(
		.INIT('h2)
	) name31679 (
		\sice_IRR_reg[1]/P0001 ,
		_w35671_,
		_w35726_
	);
	LUT2 #(
		.INIT('h8)
	) name31680 (
		\sice_SPC_reg[11]/P0001 ,
		_w35671_,
		_w35727_
	);
	LUT2 #(
		.INIT('h1)
	) name31681 (
		_w35726_,
		_w35727_,
		_w35728_
	);
	LUT2 #(
		.INIT('h2)
	) name31682 (
		_w4093_,
		_w35728_,
		_w35729_
	);
	LUT2 #(
		.INIT('h2)
	) name31683 (
		\core_c_psq_EXA_reg[1]/P0001 ,
		_w4093_,
		_w35730_
	);
	LUT2 #(
		.INIT('h1)
	) name31684 (
		_w35729_,
		_w35730_,
		_w35731_
	);
	LUT2 #(
		.INIT('h2)
	) name31685 (
		\sice_IRR_reg[12]/P0001 ,
		_w35671_,
		_w35732_
	);
	LUT2 #(
		.INIT('h8)
	) name31686 (
		\sice_SPC_reg[22]/P0001 ,
		_w35671_,
		_w35733_
	);
	LUT2 #(
		.INIT('h1)
	) name31687 (
		_w35732_,
		_w35733_,
		_w35734_
	);
	LUT2 #(
		.INIT('h2)
	) name31688 (
		_w4093_,
		_w35734_,
		_w35735_
	);
	LUT2 #(
		.INIT('h2)
	) name31689 (
		\core_c_psq_EXA_reg[12]/P0001 ,
		_w4093_,
		_w35736_
	);
	LUT2 #(
		.INIT('h1)
	) name31690 (
		_w35735_,
		_w35736_,
		_w35737_
	);
	LUT2 #(
		.INIT('h2)
	) name31691 (
		\sice_IRR_reg[11]/P0001 ,
		_w35671_,
		_w35738_
	);
	LUT2 #(
		.INIT('h8)
	) name31692 (
		\sice_SPC_reg[21]/P0001 ,
		_w35671_,
		_w35739_
	);
	LUT2 #(
		.INIT('h1)
	) name31693 (
		_w35738_,
		_w35739_,
		_w35740_
	);
	LUT2 #(
		.INIT('h2)
	) name31694 (
		_w4093_,
		_w35740_,
		_w35741_
	);
	LUT2 #(
		.INIT('h2)
	) name31695 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		_w4093_,
		_w35742_
	);
	LUT2 #(
		.INIT('h1)
	) name31696 (
		_w35741_,
		_w35742_,
		_w35743_
	);
	LUT2 #(
		.INIT('h2)
	) name31697 (
		\sice_IRR_reg[10]/P0001 ,
		_w35671_,
		_w35744_
	);
	LUT2 #(
		.INIT('h8)
	) name31698 (
		\sice_SPC_reg[20]/P0001 ,
		_w35671_,
		_w35745_
	);
	LUT2 #(
		.INIT('h1)
	) name31699 (
		_w35744_,
		_w35745_,
		_w35746_
	);
	LUT2 #(
		.INIT('h2)
	) name31700 (
		_w4093_,
		_w35746_,
		_w35747_
	);
	LUT2 #(
		.INIT('h2)
	) name31701 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		_w4093_,
		_w35748_
	);
	LUT2 #(
		.INIT('h1)
	) name31702 (
		_w35747_,
		_w35748_,
		_w35749_
	);
	LUT2 #(
		.INIT('h2)
	) name31703 (
		\sice_IRR_reg[0]/P0001 ,
		_w35671_,
		_w35750_
	);
	LUT2 #(
		.INIT('h8)
	) name31704 (
		\sice_SPC_reg[10]/P0001 ,
		_w35671_,
		_w35751_
	);
	LUT2 #(
		.INIT('h1)
	) name31705 (
		_w35750_,
		_w35751_,
		_w35752_
	);
	LUT2 #(
		.INIT('h2)
	) name31706 (
		_w4093_,
		_w35752_,
		_w35753_
	);
	LUT2 #(
		.INIT('h2)
	) name31707 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		_w4093_,
		_w35754_
	);
	LUT2 #(
		.INIT('h1)
	) name31708 (
		_w35753_,
		_w35754_,
		_w35755_
	);
	LUT2 #(
		.INIT('h8)
	) name31709 (
		_w31264_,
		_w34029_,
		_w35756_
	);
	LUT2 #(
		.INIT('h4)
	) name31710 (
		_w4117_,
		_w31271_,
		_w35757_
	);
	LUT2 #(
		.INIT('h8)
	) name31711 (
		_w35756_,
		_w35757_,
		_w35758_
	);
	LUT2 #(
		.INIT('h8)
	) name31712 (
		\core_c_dec_MFICNTL_E_reg/P0001 ,
		_w4117_,
		_w35759_
	);
	LUT2 #(
		.INIT('h1)
	) name31713 (
		_w35758_,
		_w35759_,
		_w35760_
	);
	LUT2 #(
		.INIT('h2)
	) name31714 (
		\sport0_txctl_TXSHT_reg[13]/P0001 ,
		_w19960_,
		_w35761_
	);
	LUT2 #(
		.INIT('h8)
	) name31715 (
		\sport0_txctl_TX_reg[14]/P0001 ,
		_w19960_,
		_w35762_
	);
	LUT2 #(
		.INIT('h1)
	) name31716 (
		_w35761_,
		_w35762_,
		_w35763_
	);
	LUT2 #(
		.INIT('h2)
	) name31717 (
		\sport0_txctl_TXSHT_reg[9]/P0001 ,
		_w19960_,
		_w35764_
	);
	LUT2 #(
		.INIT('h8)
	) name31718 (
		\sport0_txctl_TX_reg[10]/P0001 ,
		_w19960_,
		_w35765_
	);
	LUT2 #(
		.INIT('h1)
	) name31719 (
		_w35764_,
		_w35765_,
		_w35766_
	);
	LUT2 #(
		.INIT('h2)
	) name31720 (
		\sport0_txctl_TXSHT_reg[8]/P0001 ,
		_w19960_,
		_w35767_
	);
	LUT2 #(
		.INIT('h8)
	) name31721 (
		\sport0_txctl_TX_reg[9]/P0001 ,
		_w19960_,
		_w35768_
	);
	LUT2 #(
		.INIT('h1)
	) name31722 (
		_w35767_,
		_w35768_,
		_w35769_
	);
	LUT2 #(
		.INIT('h2)
	) name31723 (
		\sport0_txctl_TXSHT_reg[7]/P0001 ,
		_w19960_,
		_w35770_
	);
	LUT2 #(
		.INIT('h8)
	) name31724 (
		\sport0_txctl_TX_reg[8]/P0001 ,
		_w19960_,
		_w35771_
	);
	LUT2 #(
		.INIT('h1)
	) name31725 (
		_w35770_,
		_w35771_,
		_w35772_
	);
	LUT2 #(
		.INIT('h2)
	) name31726 (
		\sport1_txctl_TXSHT_reg[8]/P0001 ,
		_w22677_,
		_w35773_
	);
	LUT2 #(
		.INIT('h8)
	) name31727 (
		\sport1_txctl_TX_reg[9]/P0001 ,
		_w22677_,
		_w35774_
	);
	LUT2 #(
		.INIT('h1)
	) name31728 (
		_w35773_,
		_w35774_,
		_w35775_
	);
	LUT2 #(
		.INIT('h2)
	) name31729 (
		\sport0_txctl_TXSHT_reg[5]/P0001 ,
		_w19960_,
		_w35776_
	);
	LUT2 #(
		.INIT('h8)
	) name31730 (
		\sport0_txctl_TX_reg[6]/P0001 ,
		_w19960_,
		_w35777_
	);
	LUT2 #(
		.INIT('h1)
	) name31731 (
		_w35776_,
		_w35777_,
		_w35778_
	);
	LUT2 #(
		.INIT('h2)
	) name31732 (
		\sport1_txctl_TXSHT_reg[7]/P0001 ,
		_w22677_,
		_w35779_
	);
	LUT2 #(
		.INIT('h8)
	) name31733 (
		\sport1_txctl_TX_reg[8]/P0001 ,
		_w22677_,
		_w35780_
	);
	LUT2 #(
		.INIT('h1)
	) name31734 (
		_w35779_,
		_w35780_,
		_w35781_
	);
	LUT2 #(
		.INIT('h1)
	) name31735 (
		\sice_ICYC_reg[15]/NET0131 ,
		_w20744_,
		_w35782_
	);
	LUT2 #(
		.INIT('h1)
	) name31736 (
		_w20745_,
		_w35782_,
		_w35783_
	);
	LUT2 #(
		.INIT('h2)
	) name31737 (
		\sport0_txctl_TXSHT_reg[4]/P0001 ,
		_w19960_,
		_w35784_
	);
	LUT2 #(
		.INIT('h8)
	) name31738 (
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w19960_,
		_w35785_
	);
	LUT2 #(
		.INIT('h1)
	) name31739 (
		_w35784_,
		_w35785_,
		_w35786_
	);
	LUT2 #(
		.INIT('h1)
	) name31740 (
		\sice_IIRC_reg[15]/NET0131 ,
		_w20859_,
		_w35787_
	);
	LUT2 #(
		.INIT('h1)
	) name31741 (
		_w22581_,
		_w35787_,
		_w35788_
	);
	LUT2 #(
		.INIT('h2)
	) name31742 (
		\sport1_txctl_TXSHT_reg[5]/P0001 ,
		_w22677_,
		_w35789_
	);
	LUT2 #(
		.INIT('h8)
	) name31743 (
		\sport1_txctl_TX_reg[6]/P0001 ,
		_w22677_,
		_w35790_
	);
	LUT2 #(
		.INIT('h1)
	) name31744 (
		_w35789_,
		_w35790_,
		_w35791_
	);
	LUT2 #(
		.INIT('h2)
	) name31745 (
		\sport1_txctl_TXSHT_reg[4]/P0001 ,
		_w22677_,
		_w35792_
	);
	LUT2 #(
		.INIT('h8)
	) name31746 (
		\sport1_txctl_TX_reg[5]/P0001 ,
		_w22677_,
		_w35793_
	);
	LUT2 #(
		.INIT('h1)
	) name31747 (
		_w35792_,
		_w35793_,
		_w35794_
	);
	LUT2 #(
		.INIT('h2)
	) name31748 (
		\sport0_txctl_TXSHT_reg[2]/P0001 ,
		_w19960_,
		_w35795_
	);
	LUT2 #(
		.INIT('h8)
	) name31749 (
		\sport0_txctl_TX_reg[3]/P0001 ,
		_w19960_,
		_w35796_
	);
	LUT2 #(
		.INIT('h1)
	) name31750 (
		_w35795_,
		_w35796_,
		_w35797_
	);
	LUT2 #(
		.INIT('h2)
	) name31751 (
		\sice_ICYC_reg[0]/NET0131 ,
		_w32036_,
		_w35798_
	);
	LUT2 #(
		.INIT('h4)
	) name31752 (
		\sice_ICYC_reg[0]/NET0131 ,
		_w32036_,
		_w35799_
	);
	LUT2 #(
		.INIT('h1)
	) name31753 (
		_w35798_,
		_w35799_,
		_w35800_
	);
	LUT2 #(
		.INIT('h2)
	) name31754 (
		\sice_SPC_reg[5]/P0001 ,
		_w26297_,
		_w35801_
	);
	LUT2 #(
		.INIT('h8)
	) name31755 (
		\sice_SPC_reg[4]/P0001 ,
		_w34825_,
		_w35802_
	);
	LUT2 #(
		.INIT('h2)
	) name31756 (
		\sice_SPC_reg[6]/P0001 ,
		_w34825_,
		_w35803_
	);
	LUT2 #(
		.INIT('h1)
	) name31757 (
		_w35802_,
		_w35803_,
		_w35804_
	);
	LUT2 #(
		.INIT('h4)
	) name31758 (
		_w34827_,
		_w35804_,
		_w35805_
	);
	LUT2 #(
		.INIT('h8)
	) name31759 (
		\core_c_dec_IR_reg[5]/NET0131 ,
		_w28203_,
		_w35806_
	);
	LUT2 #(
		.INIT('h8)
	) name31760 (
		\sice_DBR2_reg[0]/P0001 ,
		_w25012_,
		_w35807_
	);
	LUT2 #(
		.INIT('h8)
	) name31761 (
		\sice_ICYC_reg[5]/NET0131 ,
		_w23409_,
		_w35808_
	);
	LUT2 #(
		.INIT('h8)
	) name31762 (
		\sice_idr0_reg_DO_reg[5]/P0001 ,
		_w26968_,
		_w35809_
	);
	LUT2 #(
		.INIT('h8)
	) name31763 (
		\sice_IIRC_reg[5]/NET0131 ,
		_w24267_,
		_w35810_
	);
	LUT2 #(
		.INIT('h8)
	) name31764 (
		\sice_DBR1_reg[0]/P0001 ,
		_w25054_,
		_w35811_
	);
	LUT2 #(
		.INIT('h1)
	) name31765 (
		_w35806_,
		_w35807_,
		_w35812_
	);
	LUT2 #(
		.INIT('h1)
	) name31766 (
		_w35808_,
		_w35809_,
		_w35813_
	);
	LUT2 #(
		.INIT('h1)
	) name31767 (
		_w35810_,
		_w35811_,
		_w35814_
	);
	LUT2 #(
		.INIT('h8)
	) name31768 (
		_w35813_,
		_w35814_,
		_w35815_
	);
	LUT2 #(
		.INIT('h8)
	) name31769 (
		_w35812_,
		_w35815_,
		_w35816_
	);
	LUT2 #(
		.INIT('h8)
	) name31770 (
		_w34827_,
		_w35816_,
		_w35817_
	);
	LUT2 #(
		.INIT('h2)
	) name31771 (
		_w26297_,
		_w35805_,
		_w35818_
	);
	LUT2 #(
		.INIT('h4)
	) name31772 (
		_w35817_,
		_w35818_,
		_w35819_
	);
	LUT2 #(
		.INIT('h1)
	) name31773 (
		_w35801_,
		_w35819_,
		_w35820_
	);
	LUT2 #(
		.INIT('h8)
	) name31774 (
		\sice_SPC_reg[8]/P0001 ,
		_w34825_,
		_w35821_
	);
	LUT2 #(
		.INIT('h2)
	) name31775 (
		\sice_SPC_reg[10]/P0001 ,
		_w34825_,
		_w35822_
	);
	LUT2 #(
		.INIT('h1)
	) name31776 (
		_w35821_,
		_w35822_,
		_w35823_
	);
	LUT2 #(
		.INIT('h4)
	) name31777 (
		_w34827_,
		_w35823_,
		_w35824_
	);
	LUT2 #(
		.INIT('h8)
	) name31778 (
		\core_c_dec_IR_reg[9]/NET0131 ,
		_w28203_,
		_w35825_
	);
	LUT2 #(
		.INIT('h8)
	) name31779 (
		\sice_DBR2_reg[4]/P0001 ,
		_w25012_,
		_w35826_
	);
	LUT2 #(
		.INIT('h8)
	) name31780 (
		\sice_IBR2_reg[3]/P0001 ,
		_w25074_,
		_w35827_
	);
	LUT2 #(
		.INIT('h8)
	) name31781 (
		\sice_IMR1_reg[3]/NET0131 ,
		_w34846_,
		_w35828_
	);
	LUT2 #(
		.INIT('h8)
	) name31782 (
		\sice_DMR2_reg[3]/NET0131 ,
		_w25025_,
		_w35829_
	);
	LUT2 #(
		.INIT('h8)
	) name31783 (
		\sice_IBR1_reg[3]/P0001 ,
		_w34831_,
		_w35830_
	);
	LUT2 #(
		.INIT('h8)
	) name31784 (
		\sice_IIRC_reg[9]/NET0131 ,
		_w24267_,
		_w35831_
	);
	LUT2 #(
		.INIT('h8)
	) name31785 (
		\sice_IMR2_reg[3]/NET0131 ,
		_w25034_,
		_w35832_
	);
	LUT2 #(
		.INIT('h8)
	) name31786 (
		\sice_DBR1_reg[4]/P0001 ,
		_w25054_,
		_w35833_
	);
	LUT2 #(
		.INIT('h8)
	) name31787 (
		\sice_idr0_reg_DO_reg[9]/P0001 ,
		_w26968_,
		_w35834_
	);
	LUT2 #(
		.INIT('h8)
	) name31788 (
		\sice_DMR1_reg[3]/NET0131 ,
		_w27903_,
		_w35835_
	);
	LUT2 #(
		.INIT('h8)
	) name31789 (
		\sice_ICYC_reg[9]/NET0131 ,
		_w23409_,
		_w35836_
	);
	LUT2 #(
		.INIT('h1)
	) name31790 (
		_w35825_,
		_w35826_,
		_w35837_
	);
	LUT2 #(
		.INIT('h1)
	) name31791 (
		_w35827_,
		_w35828_,
		_w35838_
	);
	LUT2 #(
		.INIT('h1)
	) name31792 (
		_w35829_,
		_w35830_,
		_w35839_
	);
	LUT2 #(
		.INIT('h1)
	) name31793 (
		_w35831_,
		_w35832_,
		_w35840_
	);
	LUT2 #(
		.INIT('h1)
	) name31794 (
		_w35833_,
		_w35834_,
		_w35841_
	);
	LUT2 #(
		.INIT('h1)
	) name31795 (
		_w35835_,
		_w35836_,
		_w35842_
	);
	LUT2 #(
		.INIT('h8)
	) name31796 (
		_w35841_,
		_w35842_,
		_w35843_
	);
	LUT2 #(
		.INIT('h8)
	) name31797 (
		_w35839_,
		_w35840_,
		_w35844_
	);
	LUT2 #(
		.INIT('h8)
	) name31798 (
		_w35837_,
		_w35838_,
		_w35845_
	);
	LUT2 #(
		.INIT('h8)
	) name31799 (
		_w35844_,
		_w35845_,
		_w35846_
	);
	LUT2 #(
		.INIT('h8)
	) name31800 (
		_w35843_,
		_w35846_,
		_w35847_
	);
	LUT2 #(
		.INIT('h8)
	) name31801 (
		_w34827_,
		_w35847_,
		_w35848_
	);
	LUT2 #(
		.INIT('h1)
	) name31802 (
		_w35824_,
		_w35848_,
		_w35849_
	);
	LUT2 #(
		.INIT('h2)
	) name31803 (
		\sport0_txctl_TXSHT_reg[1]/P0001 ,
		_w19960_,
		_w35850_
	);
	LUT2 #(
		.INIT('h8)
	) name31804 (
		\sport0_txctl_TX_reg[2]/P0001 ,
		_w19960_,
		_w35851_
	);
	LUT2 #(
		.INIT('h1)
	) name31805 (
		_w35850_,
		_w35851_,
		_w35852_
	);
	LUT2 #(
		.INIT('h8)
	) name31806 (
		\sice_SPC_reg[5]/P0001 ,
		_w34825_,
		_w35853_
	);
	LUT2 #(
		.INIT('h2)
	) name31807 (
		\sice_SPC_reg[7]/P0001 ,
		_w34825_,
		_w35854_
	);
	LUT2 #(
		.INIT('h1)
	) name31808 (
		_w35853_,
		_w35854_,
		_w35855_
	);
	LUT2 #(
		.INIT('h4)
	) name31809 (
		_w34827_,
		_w35855_,
		_w35856_
	);
	LUT2 #(
		.INIT('h8)
	) name31810 (
		\core_c_dec_IR_reg[6]/NET0131 ,
		_w28203_,
		_w35857_
	);
	LUT2 #(
		.INIT('h8)
	) name31811 (
		\sice_DMR1_reg[0]/NET0131 ,
		_w27903_,
		_w35858_
	);
	LUT2 #(
		.INIT('h8)
	) name31812 (
		\sice_DMR2_reg[0]/NET0131 ,
		_w25025_,
		_w35859_
	);
	LUT2 #(
		.INIT('h8)
	) name31813 (
		\sice_DBR1_reg[1]/P0001 ,
		_w25054_,
		_w35860_
	);
	LUT2 #(
		.INIT('h8)
	) name31814 (
		\sice_IMR2_reg[0]/NET0131 ,
		_w25034_,
		_w35861_
	);
	LUT2 #(
		.INIT('h8)
	) name31815 (
		\sice_IBR1_reg[0]/P0001 ,
		_w34831_,
		_w35862_
	);
	LUT2 #(
		.INIT('h8)
	) name31816 (
		\sice_IIRC_reg[6]/NET0131 ,
		_w24267_,
		_w35863_
	);
	LUT2 #(
		.INIT('h8)
	) name31817 (
		\sice_IMR1_reg[0]/NET0131 ,
		_w34846_,
		_w35864_
	);
	LUT2 #(
		.INIT('h8)
	) name31818 (
		\sice_IBR2_reg[0]/P0001 ,
		_w25074_,
		_w35865_
	);
	LUT2 #(
		.INIT('h8)
	) name31819 (
		\sice_idr0_reg_DO_reg[6]/P0001 ,
		_w26968_,
		_w35866_
	);
	LUT2 #(
		.INIT('h8)
	) name31820 (
		\sice_DBR2_reg[1]/P0001 ,
		_w25012_,
		_w35867_
	);
	LUT2 #(
		.INIT('h8)
	) name31821 (
		\sice_ICYC_reg[6]/NET0131 ,
		_w23409_,
		_w35868_
	);
	LUT2 #(
		.INIT('h1)
	) name31822 (
		_w35857_,
		_w35858_,
		_w35869_
	);
	LUT2 #(
		.INIT('h1)
	) name31823 (
		_w35859_,
		_w35860_,
		_w35870_
	);
	LUT2 #(
		.INIT('h1)
	) name31824 (
		_w35861_,
		_w35862_,
		_w35871_
	);
	LUT2 #(
		.INIT('h1)
	) name31825 (
		_w35863_,
		_w35864_,
		_w35872_
	);
	LUT2 #(
		.INIT('h1)
	) name31826 (
		_w35865_,
		_w35866_,
		_w35873_
	);
	LUT2 #(
		.INIT('h1)
	) name31827 (
		_w35867_,
		_w35868_,
		_w35874_
	);
	LUT2 #(
		.INIT('h8)
	) name31828 (
		_w35873_,
		_w35874_,
		_w35875_
	);
	LUT2 #(
		.INIT('h8)
	) name31829 (
		_w35871_,
		_w35872_,
		_w35876_
	);
	LUT2 #(
		.INIT('h8)
	) name31830 (
		_w35869_,
		_w35870_,
		_w35877_
	);
	LUT2 #(
		.INIT('h8)
	) name31831 (
		_w35876_,
		_w35877_,
		_w35878_
	);
	LUT2 #(
		.INIT('h8)
	) name31832 (
		_w35875_,
		_w35878_,
		_w35879_
	);
	LUT2 #(
		.INIT('h8)
	) name31833 (
		_w34827_,
		_w35879_,
		_w35880_
	);
	LUT2 #(
		.INIT('h1)
	) name31834 (
		_w35856_,
		_w35880_,
		_w35881_
	);
	LUT2 #(
		.INIT('h2)
	) name31835 (
		\sport0_txctl_TXSHT_reg[0]/P0001 ,
		_w19960_,
		_w35882_
	);
	LUT2 #(
		.INIT('h8)
	) name31836 (
		\sport0_txctl_TX_reg[1]/P0001 ,
		_w19960_,
		_w35883_
	);
	LUT2 #(
		.INIT('h1)
	) name31837 (
		_w35882_,
		_w35883_,
		_w35884_
	);
	LUT2 #(
		.INIT('h2)
	) name31838 (
		\sport1_txctl_TXSHT_reg[2]/P0001 ,
		_w22677_,
		_w35885_
	);
	LUT2 #(
		.INIT('h8)
	) name31839 (
		\sport1_txctl_TX_reg[3]/P0001 ,
		_w22677_,
		_w35886_
	);
	LUT2 #(
		.INIT('h1)
	) name31840 (
		_w35885_,
		_w35886_,
		_w35887_
	);
	LUT2 #(
		.INIT('h2)
	) name31841 (
		\sport1_txctl_TXSHT_reg[1]/P0001 ,
		_w22677_,
		_w35888_
	);
	LUT2 #(
		.INIT('h8)
	) name31842 (
		\sport1_txctl_TX_reg[2]/P0001 ,
		_w22677_,
		_w35889_
	);
	LUT2 #(
		.INIT('h1)
	) name31843 (
		_w35888_,
		_w35889_,
		_w35890_
	);
	LUT2 #(
		.INIT('h8)
	) name31844 (
		_w18262_,
		_w31574_,
		_w35891_
	);
	LUT2 #(
		.INIT('h1)
	) name31845 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 ,
		_w28530_,
		_w35892_
	);
	LUT2 #(
		.INIT('h4)
	) name31846 (
		_w19381_,
		_w21663_,
		_w35893_
	);
	LUT2 #(
		.INIT('h2)
	) name31847 (
		_w28534_,
		_w35893_,
		_w35894_
	);
	LUT2 #(
		.INIT('h1)
	) name31848 (
		_w35892_,
		_w35894_,
		_w35895_
	);
	LUT2 #(
		.INIT('h1)
	) name31849 (
		_w19385_,
		_w35895_,
		_w35896_
	);
	LUT2 #(
		.INIT('h1)
	) name31850 (
		\core_eu_em_mac_em_reg_mr2swe_DO_reg[3]/P0001 ,
		_w28532_,
		_w35897_
	);
	LUT2 #(
		.INIT('h1)
	) name31851 (
		_w35896_,
		_w35897_,
		_w35898_
	);
	LUT2 #(
		.INIT('h2)
	) name31852 (
		_w28529_,
		_w35898_,
		_w35899_
	);
	LUT2 #(
		.INIT('h1)
	) name31853 (
		_w35891_,
		_w35899_,
		_w35900_
	);
	LUT2 #(
		.INIT('h8)
	) name31854 (
		\sport0_txctl_TX_reg[0]/P0001 ,
		_w19960_,
		_w35901_
	);
	LUT2 #(
		.INIT('h2)
	) name31855 (
		\sport1_txctl_TXSHT_reg[0]/P0001 ,
		_w22677_,
		_w35902_
	);
	LUT2 #(
		.INIT('h8)
	) name31856 (
		\sport1_txctl_TX_reg[1]/P0001 ,
		_w22677_,
		_w35903_
	);
	LUT2 #(
		.INIT('h1)
	) name31857 (
		_w35902_,
		_w35903_,
		_w35904_
	);
	LUT2 #(
		.INIT('h2)
	) name31858 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w5607_,
		_w35905_
	);
	LUT2 #(
		.INIT('h1)
	) name31859 (
		_w5582_,
		_w20208_,
		_w35906_
	);
	LUT2 #(
		.INIT('h2)
	) name31860 (
		_w12442_,
		_w35906_,
		_w35907_
	);
	LUT2 #(
		.INIT('h2)
	) name31861 (
		\memc_Dwrite_E_reg/NET0131 ,
		_w5600_,
		_w35908_
	);
	LUT2 #(
		.INIT('h1)
	) name31862 (
		_w35905_,
		_w35908_,
		_w35909_
	);
	LUT2 #(
		.INIT('h4)
	) name31863 (
		_w35907_,
		_w35909_,
		_w35910_
	);
	LUT2 #(
		.INIT('h1)
	) name31864 (
		_w5581_,
		_w5597_,
		_w35911_
	);
	LUT2 #(
		.INIT('h8)
	) name31865 (
		_w5560_,
		_w35911_,
		_w35912_
	);
	LUT2 #(
		.INIT('h8)
	) name31866 (
		_w5586_,
		_w35912_,
		_w35913_
	);
	LUT2 #(
		.INIT('h8)
	) name31867 (
		\bdma_BCTL_reg[2]/NET0131 ,
		_w35913_,
		_w35914_
	);
	LUT2 #(
		.INIT('h2)
	) name31868 (
		_w5599_,
		_w14732_,
		_w35915_
	);
	LUT2 #(
		.INIT('h4)
	) name31869 (
		_w12442_,
		_w20208_,
		_w35916_
	);
	LUT2 #(
		.INIT('h8)
	) name31870 (
		\memc_Pread_E_reg/NET0131 ,
		_w5606_,
		_w35917_
	);
	LUT2 #(
		.INIT('h1)
	) name31871 (
		_w35913_,
		_w35915_,
		_w35918_
	);
	LUT2 #(
		.INIT('h4)
	) name31872 (
		_w35917_,
		_w35918_,
		_w35919_
	);
	LUT2 #(
		.INIT('h4)
	) name31873 (
		_w35916_,
		_w35919_,
		_w35920_
	);
	LUT2 #(
		.INIT('h1)
	) name31874 (
		_w35914_,
		_w35920_,
		_w35921_
	);
	LUT2 #(
		.INIT('h8)
	) name31875 (
		_w12442_,
		_w20208_,
		_w35922_
	);
	LUT2 #(
		.INIT('h8)
	) name31876 (
		\memc_Pwrite_E_reg/NET0131 ,
		_w5606_,
		_w35923_
	);
	LUT2 #(
		.INIT('h8)
	) name31877 (
		\memc_Dwrite_E_reg/NET0131 ,
		_w5599_,
		_w35924_
	);
	LUT2 #(
		.INIT('h1)
	) name31878 (
		_w35923_,
		_w35924_,
		_w35925_
	);
	LUT2 #(
		.INIT('h4)
	) name31879 (
		_w35922_,
		_w35925_,
		_w35926_
	);
	LUT2 #(
		.INIT('h8)
	) name31880 (
		\sport1_txctl_TX_reg[0]/P0001 ,
		_w22677_,
		_w35927_
	);
	LUT2 #(
		.INIT('h1)
	) name31881 (
		_w5556_,
		_w35912_,
		_w35928_
	);
	LUT2 #(
		.INIT('h2)
	) name31882 (
		\core_c_psq_PCS_reg[12]/NET0131 ,
		\emc_eRDY_reg/NET0131 ,
		_w35929_
	);
	LUT2 #(
		.INIT('h2)
	) name31883 (
		\core_c_psq_PCS_reg[1]/NET0131 ,
		_w4068_,
		_w35930_
	);
	LUT2 #(
		.INIT('h1)
	) name31884 (
		_w35929_,
		_w35930_,
		_w35931_
	);
	LUT2 #(
		.INIT('h8)
	) name31885 (
		_w5700_,
		_w35931_,
		_w35932_
	);
	LUT2 #(
		.INIT('h1)
	) name31886 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w35932_,
		_w35933_
	);
	LUT2 #(
		.INIT('h2)
	) name31887 (
		_w19047_,
		_w35933_,
		_w35934_
	);
	LUT2 #(
		.INIT('h2)
	) name31888 (
		_w4118_,
		_w35934_,
		_w35935_
	);
	LUT2 #(
		.INIT('h2)
	) name31889 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w19504_,
		_w35936_
	);
	LUT2 #(
		.INIT('h4)
	) name31890 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w29555_,
		_w35937_
	);
	LUT2 #(
		.INIT('h1)
	) name31891 (
		_w35936_,
		_w35937_,
		_w35938_
	);
	LUT2 #(
		.INIT('h2)
	) name31892 (
		_w18886_,
		_w35938_,
		_w35939_
	);
	LUT2 #(
		.INIT('h1)
	) name31893 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[9]/P0001 ,
		_w18886_,
		_w35940_
	);
	LUT2 #(
		.INIT('h1)
	) name31894 (
		_w35939_,
		_w35940_,
		_w35941_
	);
	LUT2 #(
		.INIT('h2)
	) name31895 (
		_w19034_,
		_w35938_,
		_w35942_
	);
	LUT2 #(
		.INIT('h1)
	) name31896 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[9]/P0001 ,
		_w19034_,
		_w35943_
	);
	LUT2 #(
		.INIT('h1)
	) name31897 (
		_w35942_,
		_w35943_,
		_w35944_
	);
	LUT2 #(
		.INIT('h2)
	) name31898 (
		_w18513_,
		_w23044_,
		_w35945_
	);
	LUT2 #(
		.INIT('h2)
	) name31899 (
		_w18471_,
		_w35945_,
		_w35946_
	);
	LUT2 #(
		.INIT('h1)
	) name31900 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w35946_,
		_w35947_
	);
	LUT2 #(
		.INIT('h8)
	) name31901 (
		\sport0_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w35946_,
		_w35948_
	);
	LUT2 #(
		.INIT('h2)
	) name31902 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w35947_,
		_w35949_
	);
	LUT2 #(
		.INIT('h4)
	) name31903 (
		_w35948_,
		_w35949_,
		_w35950_
	);
	LUT2 #(
		.INIT('h4)
	) name31904 (
		\sport0_txctl_TX_reg[5]/P0001 ,
		_w18519_,
		_w35951_
	);
	LUT2 #(
		.INIT('h1)
	) name31905 (
		_w10911_,
		_w18519_,
		_w35952_
	);
	LUT2 #(
		.INIT('h1)
	) name31906 (
		\sport0_txctl_ldTX_cmp_reg/P0001 ,
		_w35951_,
		_w35953_
	);
	LUT2 #(
		.INIT('h4)
	) name31907 (
		_w35952_,
		_w35953_,
		_w35954_
	);
	LUT2 #(
		.INIT('h1)
	) name31908 (
		_w35950_,
		_w35954_,
		_w35955_
	);
	LUT2 #(
		.INIT('h8)
	) name31909 (
		\ISCLK0_pad ,
		\sport0_cfg_SCLKi_h_reg/NET0131 ,
		_w35956_
	);
	LUT2 #(
		.INIT('h1)
	) name31910 (
		\T_SCLK0_pad ,
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w35957_
	);
	LUT2 #(
		.INIT('h8)
	) name31911 (
		\T_SCLK0_pad ,
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w35958_
	);
	LUT2 #(
		.INIT('h1)
	) name31912 (
		\ISCLK0_pad ,
		_w35957_,
		_w35959_
	);
	LUT2 #(
		.INIT('h4)
	) name31913 (
		_w35958_,
		_w35959_,
		_w35960_
	);
	LUT2 #(
		.INIT('h1)
	) name31914 (
		_w35956_,
		_w35960_,
		_w35961_
	);
	LUT2 #(
		.INIT('h8)
	) name31915 (
		\ISCLK1_pad ,
		\sport1_cfg_SCLKi_h_reg/NET0131 ,
		_w35962_
	);
	LUT2 #(
		.INIT('h1)
	) name31916 (
		\T_SCLK1_pad ,
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w35963_
	);
	LUT2 #(
		.INIT('h8)
	) name31917 (
		\T_SCLK1_pad ,
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w35964_
	);
	LUT2 #(
		.INIT('h1)
	) name31918 (
		\ISCLK1_pad ,
		_w35963_,
		_w35965_
	);
	LUT2 #(
		.INIT('h4)
	) name31919 (
		_w35964_,
		_w35965_,
		_w35966_
	);
	LUT2 #(
		.INIT('h1)
	) name31920 (
		_w35962_,
		_w35966_,
		_w35967_
	);
	LUT2 #(
		.INIT('h2)
	) name31921 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w23860_,
		_w35968_
	);
	LUT2 #(
		.INIT('h4)
	) name31922 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w30392_,
		_w35969_
	);
	LUT2 #(
		.INIT('h1)
	) name31923 (
		_w35968_,
		_w35969_,
		_w35970_
	);
	LUT2 #(
		.INIT('h2)
	) name31924 (
		_w18717_,
		_w35970_,
		_w35971_
	);
	LUT2 #(
		.INIT('h1)
	) name31925 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[8]/P0001 ,
		_w18717_,
		_w35972_
	);
	LUT2 #(
		.INIT('h1)
	) name31926 (
		_w35971_,
		_w35972_,
		_w35973_
	);
	LUT2 #(
		.INIT('h1)
	) name31927 (
		_w13806_,
		_w19222_,
		_w35974_
	);
	LUT2 #(
		.INIT('h8)
	) name31928 (
		_w13806_,
		_w14540_,
		_w35975_
	);
	LUT2 #(
		.INIT('h1)
	) name31929 (
		_w35974_,
		_w35975_,
		_w35976_
	);
	LUT2 #(
		.INIT('h2)
	) name31930 (
		_w14667_,
		_w35976_,
		_w35977_
	);
	LUT2 #(
		.INIT('h2)
	) name31931 (
		\core_eu_ea_alu_ea_reg_afswe_DO_reg[15]/P0001 ,
		_w14667_,
		_w35978_
	);
	LUT2 #(
		.INIT('h1)
	) name31932 (
		_w35977_,
		_w35978_,
		_w35979_
	);
	LUT2 #(
		.INIT('h2)
	) name31933 (
		_w13805_,
		_w35976_,
		_w35980_
	);
	LUT2 #(
		.INIT('h2)
	) name31934 (
		\core_eu_ea_alu_ea_reg_afrwe_DO_reg[15]/P0001 ,
		_w13805_,
		_w35981_
	);
	LUT2 #(
		.INIT('h1)
	) name31935 (
		_w35980_,
		_w35981_,
		_w35982_
	);
	LUT2 #(
		.INIT('h2)
	) name31936 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w23757_,
		_w35983_
	);
	LUT2 #(
		.INIT('h4)
	) name31937 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w29839_,
		_w35984_
	);
	LUT2 #(
		.INIT('h1)
	) name31938 (
		_w35983_,
		_w35984_,
		_w35985_
	);
	LUT2 #(
		.INIT('h2)
	) name31939 (
		_w18717_,
		_w35985_,
		_w35986_
	);
	LUT2 #(
		.INIT('h1)
	) name31940 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[11]/P0001 ,
		_w18717_,
		_w35987_
	);
	LUT2 #(
		.INIT('h1)
	) name31941 (
		_w35986_,
		_w35987_,
		_w35988_
	);
	LUT2 #(
		.INIT('h2)
	) name31942 (
		_w17833_,
		_w35970_,
		_w35989_
	);
	LUT2 #(
		.INIT('h1)
	) name31943 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[8]/P0001 ,
		_w17833_,
		_w35990_
	);
	LUT2 #(
		.INIT('h1)
	) name31944 (
		_w35989_,
		_w35990_,
		_w35991_
	);
	LUT2 #(
		.INIT('h2)
	) name31945 (
		_w17833_,
		_w35985_,
		_w35992_
	);
	LUT2 #(
		.INIT('h1)
	) name31946 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[11]/P0001 ,
		_w17833_,
		_w35993_
	);
	LUT2 #(
		.INIT('h1)
	) name31947 (
		_w35992_,
		_w35993_,
		_w35994_
	);
	LUT2 #(
		.INIT('h2)
	) name31948 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w17820_,
		_w35995_
	);
	LUT2 #(
		.INIT('h4)
	) name31949 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w29285_,
		_w35996_
	);
	LUT2 #(
		.INIT('h1)
	) name31950 (
		_w35995_,
		_w35996_,
		_w35997_
	);
	LUT2 #(
		.INIT('h2)
	) name31951 (
		_w18886_,
		_w35997_,
		_w35998_
	);
	LUT2 #(
		.INIT('h1)
	) name31952 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[15]/P0001 ,
		_w18886_,
		_w35999_
	);
	LUT2 #(
		.INIT('h1)
	) name31953 (
		_w35998_,
		_w35999_,
		_w36000_
	);
	LUT2 #(
		.INIT('h2)
	) name31954 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w23277_,
		_w36001_
	);
	LUT2 #(
		.INIT('h2)
	) name31955 (
		\sport0_txctl_Bcnt_reg[3]/NET0131 ,
		_w19956_,
		_w36002_
	);
	LUT2 #(
		.INIT('h1)
	) name31956 (
		_w19957_,
		_w36002_,
		_w36003_
	);
	LUT2 #(
		.INIT('h2)
	) name31957 (
		_w23277_,
		_w36003_,
		_w36004_
	);
	LUT2 #(
		.INIT('h1)
	) name31958 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w36001_,
		_w36005_
	);
	LUT2 #(
		.INIT('h4)
	) name31959 (
		_w36004_,
		_w36005_,
		_w36006_
	);
	LUT2 #(
		.INIT('h2)
	) name31960 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w23265_,
		_w36007_
	);
	LUT2 #(
		.INIT('h2)
	) name31961 (
		\sport1_txctl_Bcnt_reg[3]/NET0131 ,
		_w22673_,
		_w36008_
	);
	LUT2 #(
		.INIT('h1)
	) name31962 (
		_w22674_,
		_w36008_,
		_w36009_
	);
	LUT2 #(
		.INIT('h2)
	) name31963 (
		_w23265_,
		_w36009_,
		_w36010_
	);
	LUT2 #(
		.INIT('h1)
	) name31964 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w36007_,
		_w36011_
	);
	LUT2 #(
		.INIT('h4)
	) name31965 (
		_w36010_,
		_w36011_,
		_w36012_
	);
	LUT2 #(
		.INIT('h2)
	) name31966 (
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w23265_,
		_w36013_
	);
	LUT2 #(
		.INIT('h2)
	) name31967 (
		\sport1_txctl_Bcnt_reg[2]/NET0131 ,
		_w22672_,
		_w36014_
	);
	LUT2 #(
		.INIT('h1)
	) name31968 (
		_w22673_,
		_w36014_,
		_w36015_
	);
	LUT2 #(
		.INIT('h2)
	) name31969 (
		_w23265_,
		_w36015_,
		_w36016_
	);
	LUT2 #(
		.INIT('h1)
	) name31970 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w36013_,
		_w36017_
	);
	LUT2 #(
		.INIT('h4)
	) name31971 (
		_w36016_,
		_w36017_,
		_w36018_
	);
	LUT2 #(
		.INIT('h2)
	) name31972 (
		_w19034_,
		_w35997_,
		_w36019_
	);
	LUT2 #(
		.INIT('h1)
	) name31973 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[15]/P0001 ,
		_w19034_,
		_w36020_
	);
	LUT2 #(
		.INIT('h1)
	) name31974 (
		_w36019_,
		_w36020_,
		_w36021_
	);
	LUT2 #(
		.INIT('h2)
	) name31975 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w23265_,
		_w36022_
	);
	LUT2 #(
		.INIT('h8)
	) name31976 (
		\sport1_txctl_Bcnt_reg[0]/NET0131 ,
		\sport1_txctl_Bcnt_reg[1]/NET0131 ,
		_w36023_
	);
	LUT2 #(
		.INIT('h1)
	) name31977 (
		_w22672_,
		_w36023_,
		_w36024_
	);
	LUT2 #(
		.INIT('h2)
	) name31978 (
		_w23265_,
		_w36024_,
		_w36025_
	);
	LUT2 #(
		.INIT('h1)
	) name31979 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w36022_,
		_w36026_
	);
	LUT2 #(
		.INIT('h4)
	) name31980 (
		_w36025_,
		_w36026_,
		_w36027_
	);
	LUT2 #(
		.INIT('h1)
	) name31981 (
		T_IRDn_pad,
		T_ISn_pad,
		_w36028_
	);
	LUT2 #(
		.INIT('h4)
	) name31982 (
		\sport1_txctl_Bcnt_reg[0]/NET0131 ,
		_w23265_,
		_w36029_
	);
	LUT2 #(
		.INIT('h2)
	) name31983 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w23265_,
		_w36030_
	);
	LUT2 #(
		.INIT('h1)
	) name31984 (
		\sport1_rxctl_TAG_SLOT_reg/P0001 ,
		_w36029_,
		_w36031_
	);
	LUT2 #(
		.INIT('h4)
	) name31985 (
		_w36030_,
		_w36031_,
		_w36032_
	);
	LUT2 #(
		.INIT('h2)
	) name31986 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w23277_,
		_w36033_
	);
	LUT2 #(
		.INIT('h8)
	) name31987 (
		\sport0_txctl_Bcnt_reg[0]/NET0131 ,
		\sport0_txctl_Bcnt_reg[1]/NET0131 ,
		_w36034_
	);
	LUT2 #(
		.INIT('h1)
	) name31988 (
		_w19955_,
		_w36034_,
		_w36035_
	);
	LUT2 #(
		.INIT('h2)
	) name31989 (
		_w23277_,
		_w36035_,
		_w36036_
	);
	LUT2 #(
		.INIT('h1)
	) name31990 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w36033_,
		_w36037_
	);
	LUT2 #(
		.INIT('h4)
	) name31991 (
		_w36036_,
		_w36037_,
		_w36038_
	);
	LUT2 #(
		.INIT('h4)
	) name31992 (
		\sport0_txctl_Bcnt_reg[0]/NET0131 ,
		_w23277_,
		_w36039_
	);
	LUT2 #(
		.INIT('h2)
	) name31993 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w23277_,
		_w36040_
	);
	LUT2 #(
		.INIT('h1)
	) name31994 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w36039_,
		_w36041_
	);
	LUT2 #(
		.INIT('h4)
	) name31995 (
		_w36040_,
		_w36041_,
		_w36042_
	);
	LUT2 #(
		.INIT('h2)
	) name31996 (
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w23277_,
		_w36043_
	);
	LUT2 #(
		.INIT('h2)
	) name31997 (
		\sport0_txctl_Bcnt_reg[2]/NET0131 ,
		_w19955_,
		_w36044_
	);
	LUT2 #(
		.INIT('h1)
	) name31998 (
		_w19956_,
		_w36044_,
		_w36045_
	);
	LUT2 #(
		.INIT('h2)
	) name31999 (
		_w23277_,
		_w36045_,
		_w36046_
	);
	LUT2 #(
		.INIT('h1)
	) name32000 (
		\sport0_rxctl_TAG_SLOT_reg/P0001 ,
		_w36043_,
		_w36047_
	);
	LUT2 #(
		.INIT('h4)
	) name32001 (
		_w36046_,
		_w36047_,
		_w36048_
	);
	LUT2 #(
		.INIT('h2)
	) name32002 (
		_w23715_,
		_w33221_,
		_w36049_
	);
	LUT2 #(
		.INIT('h1)
	) name32003 (
		\clkc_OUTcnt_reg[3]/NET0131 ,
		_w19469_,
		_w36050_
	);
	LUT2 #(
		.INIT('h1)
	) name32004 (
		_w19470_,
		_w36050_,
		_w36051_
	);
	LUT2 #(
		.INIT('h4)
	) name32005 (
		_w19467_,
		_w36051_,
		_w36052_
	);
	LUT2 #(
		.INIT('h1)
	) name32006 (
		\clkc_STDcnt_reg[3]/NET0131 ,
		_w31523_,
		_w36053_
	);
	LUT2 #(
		.INIT('h1)
	) name32007 (
		_w31524_,
		_w36053_,
		_w36054_
	);
	LUT2 #(
		.INIT('h4)
	) name32008 (
		_w31521_,
		_w36054_,
		_w36055_
	);
	LUT2 #(
		.INIT('h4)
	) name32009 (
		\core_c_dec_Usecond_E_reg/P0001 ,
		_w4117_,
		_w36056_
	);
	LUT2 #(
		.INIT('h8)
	) name32010 (
		_w6115_,
		_w21249_,
		_w36057_
	);
	LUT2 #(
		.INIT('h4)
	) name32011 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w19529_,
		_w36058_
	);
	LUT2 #(
		.INIT('h2)
	) name32012 (
		_w21256_,
		_w36057_,
		_w36059_
	);
	LUT2 #(
		.INIT('h1)
	) name32013 (
		_w21428_,
		_w36058_,
		_w36060_
	);
	LUT2 #(
		.INIT('h8)
	) name32014 (
		_w36059_,
		_w36060_,
		_w36061_
	);
	LUT2 #(
		.INIT('h8)
	) name32015 (
		_w14729_,
		_w36061_,
		_w36062_
	);
	LUT2 #(
		.INIT('h2)
	) name32016 (
		_w4116_,
		_w36056_,
		_w36063_
	);
	LUT2 #(
		.INIT('h4)
	) name32017 (
		_w36062_,
		_w36063_,
		_w36064_
	);
	LUT2 #(
		.INIT('h1)
	) name32018 (
		\sport0_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		_w19534_,
		_w36065_
	);
	LUT2 #(
		.INIT('h1)
	) name32019 (
		_w19535_,
		_w36065_,
		_w36066_
	);
	LUT2 #(
		.INIT('h8)
	) name32020 (
		_w19197_,
		_w36066_,
		_w36067_
	);
	LUT2 #(
		.INIT('h2)
	) name32021 (
		\idma_WRcyc_reg/NET0131 ,
		_w32460_,
		_w36068_
	);
	LUT2 #(
		.INIT('h8)
	) name32022 (
		_w20382_,
		_w36068_,
		_w36069_
	);
	LUT2 #(
		.INIT('h4)
	) name32023 (
		_w20386_,
		_w20821_,
		_w36070_
	);
	LUT2 #(
		.INIT('h1)
	) name32024 (
		\idma_DSreq_reg/NET0131 ,
		_w36070_,
		_w36071_
	);
	LUT2 #(
		.INIT('h4)
	) name32025 (
		_w36069_,
		_w36071_,
		_w36072_
	);
	LUT2 #(
		.INIT('h8)
	) name32026 (
		_w20070_,
		_w22457_,
		_w36073_
	);
	LUT2 #(
		.INIT('h8)
	) name32027 (
		_w10638_,
		_w36073_,
		_w36074_
	);
	LUT2 #(
		.INIT('h8)
	) name32028 (
		_w12688_,
		_w18946_,
		_w36075_
	);
	LUT2 #(
		.INIT('h2)
	) name32029 (
		\IRFS1_pad ,
		_w36073_,
		_w36076_
	);
	LUT2 #(
		.INIT('h1)
	) name32030 (
		_w36075_,
		_w36076_,
		_w36077_
	);
	LUT2 #(
		.INIT('h4)
	) name32031 (
		_w36074_,
		_w36077_,
		_w36078_
	);
	LUT2 #(
		.INIT('h8)
	) name32032 (
		_w10289_,
		_w36073_,
		_w36079_
	);
	LUT2 #(
		.INIT('h2)
	) name32033 (
		\ITFS1_pad ,
		_w36073_,
		_w36080_
	);
	LUT2 #(
		.INIT('h1)
	) name32034 (
		_w36075_,
		_w36080_,
		_w36081_
	);
	LUT2 #(
		.INIT('h4)
	) name32035 (
		_w36079_,
		_w36081_,
		_w36082_
	);
	LUT2 #(
		.INIT('h8)
	) name32036 (
		_w9435_,
		_w36073_,
		_w36083_
	);
	LUT2 #(
		.INIT('h2)
	) name32037 (
		\sport1_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w36073_,
		_w36084_
	);
	LUT2 #(
		.INIT('h1)
	) name32038 (
		_w36075_,
		_w36084_,
		_w36085_
	);
	LUT2 #(
		.INIT('h4)
	) name32039 (
		_w36083_,
		_w36085_,
		_w36086_
	);
	LUT2 #(
		.INIT('h8)
	) name32040 (
		_w8460_,
		_w36073_,
		_w36087_
	);
	LUT2 #(
		.INIT('h2)
	) name32041 (
		\sport1_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w36073_,
		_w36088_
	);
	LUT2 #(
		.INIT('h1)
	) name32042 (
		_w36075_,
		_w36088_,
		_w36089_
	);
	LUT2 #(
		.INIT('h4)
	) name32043 (
		_w36087_,
		_w36089_,
		_w36090_
	);
	LUT2 #(
		.INIT('h8)
	) name32044 (
		_w7859_,
		_w36073_,
		_w36091_
	);
	LUT2 #(
		.INIT('h2)
	) name32045 (
		\sport1_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w36073_,
		_w36092_
	);
	LUT2 #(
		.INIT('h1)
	) name32046 (
		_w36075_,
		_w36092_,
		_w36093_
	);
	LUT2 #(
		.INIT('h4)
	) name32047 (
		_w36091_,
		_w36093_,
		_w36094_
	);
	LUT2 #(
		.INIT('h8)
	) name32048 (
		_w7607_,
		_w36073_,
		_w36095_
	);
	LUT2 #(
		.INIT('h2)
	) name32049 (
		\sport1_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w36073_,
		_w36096_
	);
	LUT2 #(
		.INIT('h1)
	) name32050 (
		_w36075_,
		_w36096_,
		_w36097_
	);
	LUT2 #(
		.INIT('h4)
	) name32051 (
		_w36095_,
		_w36097_,
		_w36098_
	);
	LUT2 #(
		.INIT('h1)
	) name32052 (
		\sport1_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w18946_,
		_w36099_
	);
	LUT2 #(
		.INIT('h4)
	) name32053 (
		_w8715_,
		_w18948_,
		_w36100_
	);
	LUT2 #(
		.INIT('h1)
	) name32054 (
		_w36099_,
		_w36100_,
		_w36101_
	);
	LUT2 #(
		.INIT('h1)
	) name32055 (
		\sport1_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w18946_,
		_w36102_
	);
	LUT2 #(
		.INIT('h4)
	) name32056 (
		_w8113_,
		_w18948_,
		_w36103_
	);
	LUT2 #(
		.INIT('h1)
	) name32057 (
		_w36102_,
		_w36103_,
		_w36104_
	);
	LUT2 #(
		.INIT('h1)
	) name32058 (
		\sport1_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w18946_,
		_w36105_
	);
	LUT2 #(
		.INIT('h4)
	) name32059 (
		_w12743_,
		_w18948_,
		_w36106_
	);
	LUT2 #(
		.INIT('h1)
	) name32060 (
		_w36105_,
		_w36106_,
		_w36107_
	);
	LUT2 #(
		.INIT('h8)
	) name32061 (
		_w18227_,
		_w20071_,
		_w36108_
	);
	LUT2 #(
		.INIT('h8)
	) name32062 (
		_w11265_,
		_w36108_,
		_w36109_
	);
	LUT2 #(
		.INIT('h2)
	) name32063 (
		\sport1_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w36108_,
		_w36110_
	);
	LUT2 #(
		.INIT('h1)
	) name32064 (
		_w36075_,
		_w36110_,
		_w36111_
	);
	LUT2 #(
		.INIT('h4)
	) name32065 (
		_w36109_,
		_w36111_,
		_w36112_
	);
	LUT2 #(
		.INIT('h8)
	) name32066 (
		_w11525_,
		_w36108_,
		_w36113_
	);
	LUT2 #(
		.INIT('h2)
	) name32067 (
		\sport1_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w36108_,
		_w36114_
	);
	LUT2 #(
		.INIT('h1)
	) name32068 (
		_w36075_,
		_w36114_,
		_w36115_
	);
	LUT2 #(
		.INIT('h4)
	) name32069 (
		_w36113_,
		_w36115_,
		_w36116_
	);
	LUT2 #(
		.INIT('h8)
	) name32070 (
		_w10911_,
		_w36108_,
		_w36117_
	);
	LUT2 #(
		.INIT('h2)
	) name32071 (
		\sport1_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w36108_,
		_w36118_
	);
	LUT2 #(
		.INIT('h1)
	) name32072 (
		_w36075_,
		_w36118_,
		_w36119_
	);
	LUT2 #(
		.INIT('h4)
	) name32073 (
		_w36117_,
		_w36119_,
		_w36120_
	);
	LUT2 #(
		.INIT('h8)
	) name32074 (
		_w10069_,
		_w36108_,
		_w36121_
	);
	LUT2 #(
		.INIT('h2)
	) name32075 (
		\sport1_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w36108_,
		_w36122_
	);
	LUT2 #(
		.INIT('h1)
	) name32076 (
		_w36075_,
		_w36122_,
		_w36123_
	);
	LUT2 #(
		.INIT('h4)
	) name32077 (
		_w36121_,
		_w36123_,
		_w36124_
	);
	LUT2 #(
		.INIT('h8)
	) name32078 (
		_w8113_,
		_w36108_,
		_w36125_
	);
	LUT2 #(
		.INIT('h2)
	) name32079 (
		\sport1_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w36108_,
		_w36126_
	);
	LUT2 #(
		.INIT('h1)
	) name32080 (
		_w36075_,
		_w36126_,
		_w36127_
	);
	LUT2 #(
		.INIT('h4)
	) name32081 (
		_w36125_,
		_w36127_,
		_w36128_
	);
	LUT2 #(
		.INIT('h8)
	) name32082 (
		_w8715_,
		_w36108_,
		_w36129_
	);
	LUT2 #(
		.INIT('h2)
	) name32083 (
		\sport1_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w36108_,
		_w36130_
	);
	LUT2 #(
		.INIT('h1)
	) name32084 (
		_w36075_,
		_w36130_,
		_w36131_
	);
	LUT2 #(
		.INIT('h4)
	) name32085 (
		_w36129_,
		_w36131_,
		_w36132_
	);
	LUT2 #(
		.INIT('h8)
	) name32086 (
		_w9435_,
		_w36108_,
		_w36133_
	);
	LUT2 #(
		.INIT('h2)
	) name32087 (
		\sport1_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w36108_,
		_w36134_
	);
	LUT2 #(
		.INIT('h1)
	) name32088 (
		_w36075_,
		_w36134_,
		_w36135_
	);
	LUT2 #(
		.INIT('h4)
	) name32089 (
		_w36133_,
		_w36135_,
		_w36136_
	);
	LUT2 #(
		.INIT('h8)
	) name32090 (
		_w7607_,
		_w36108_,
		_w36137_
	);
	LUT2 #(
		.INIT('h2)
	) name32091 (
		\sport1_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w36108_,
		_w36138_
	);
	LUT2 #(
		.INIT('h1)
	) name32092 (
		_w36075_,
		_w36138_,
		_w36139_
	);
	LUT2 #(
		.INIT('h4)
	) name32093 (
		_w36137_,
		_w36139_,
		_w36140_
	);
	LUT2 #(
		.INIT('h1)
	) name32094 (
		\sport1_cfg_SCLKi_cnt_reg[3]/NET0131 ,
		_w20232_,
		_w36141_
	);
	LUT2 #(
		.INIT('h1)
	) name32095 (
		_w20233_,
		_w36141_,
		_w36142_
	);
	LUT2 #(
		.INIT('h8)
	) name32096 (
		_w19130_,
		_w36142_,
		_w36143_
	);
	LUT2 #(
		.INIT('h8)
	) name32097 (
		_w10289_,
		_w18229_,
		_w36144_
	);
	LUT2 #(
		.INIT('h2)
	) name32098 (
		\ITFS0_pad ,
		_w18229_,
		_w36145_
	);
	LUT2 #(
		.INIT('h1)
	) name32099 (
		_w18232_,
		_w36145_,
		_w36146_
	);
	LUT2 #(
		.INIT('h4)
	) name32100 (
		_w36144_,
		_w36146_,
		_w36147_
	);
	LUT2 #(
		.INIT('h8)
	) name32101 (
		_w10638_,
		_w18229_,
		_w36148_
	);
	LUT2 #(
		.INIT('h2)
	) name32102 (
		\IRFS0_pad ,
		_w18229_,
		_w36149_
	);
	LUT2 #(
		.INIT('h1)
	) name32103 (
		_w18232_,
		_w36149_,
		_w36150_
	);
	LUT2 #(
		.INIT('h4)
	) name32104 (
		_w36148_,
		_w36150_,
		_w36151_
	);
	LUT2 #(
		.INIT('h8)
	) name32105 (
		_w9435_,
		_w18229_,
		_w36152_
	);
	LUT2 #(
		.INIT('h2)
	) name32106 (
		\sport0_regs_SCTLreg_DO_reg[1]/NET0131 ,
		_w18229_,
		_w36153_
	);
	LUT2 #(
		.INIT('h1)
	) name32107 (
		_w18232_,
		_w36153_,
		_w36154_
	);
	LUT2 #(
		.INIT('h4)
	) name32108 (
		_w36152_,
		_w36154_,
		_w36155_
	);
	LUT2 #(
		.INIT('h8)
	) name32109 (
		_w8460_,
		_w18229_,
		_w36156_
	);
	LUT2 #(
		.INIT('h2)
	) name32110 (
		\sport0_regs_SCTLreg_DO_reg[11]/NET0131 ,
		_w18229_,
		_w36157_
	);
	LUT2 #(
		.INIT('h1)
	) name32111 (
		_w18232_,
		_w36157_,
		_w36158_
	);
	LUT2 #(
		.INIT('h4)
	) name32112 (
		_w36156_,
		_w36158_,
		_w36159_
	);
	LUT2 #(
		.INIT('h8)
	) name32113 (
		_w7859_,
		_w18229_,
		_w36160_
	);
	LUT2 #(
		.INIT('h2)
	) name32114 (
		\sport0_regs_SCTLreg_DO_reg[10]/NET0131 ,
		_w18229_,
		_w36161_
	);
	LUT2 #(
		.INIT('h1)
	) name32115 (
		_w18232_,
		_w36161_,
		_w36162_
	);
	LUT2 #(
		.INIT('h4)
	) name32116 (
		_w36160_,
		_w36162_,
		_w36163_
	);
	LUT2 #(
		.INIT('h8)
	) name32117 (
		_w7607_,
		_w18229_,
		_w36164_
	);
	LUT2 #(
		.INIT('h2)
	) name32118 (
		\sport0_regs_SCTLreg_DO_reg[0]/NET0131 ,
		_w18229_,
		_w36165_
	);
	LUT2 #(
		.INIT('h1)
	) name32119 (
		_w18232_,
		_w36165_,
		_w36166_
	);
	LUT2 #(
		.INIT('h4)
	) name32120 (
		_w36164_,
		_w36166_,
		_w36167_
	);
	LUT2 #(
		.INIT('h1)
	) name32121 (
		\sport0_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w18231_,
		_w36168_
	);
	LUT2 #(
		.INIT('h4)
	) name32122 (
		_w8113_,
		_w19015_,
		_w36169_
	);
	LUT2 #(
		.INIT('h1)
	) name32123 (
		_w36168_,
		_w36169_,
		_w36170_
	);
	LUT2 #(
		.INIT('h1)
	) name32124 (
		\sport0_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w18231_,
		_w36171_
	);
	LUT2 #(
		.INIT('h4)
	) name32125 (
		_w8715_,
		_w19015_,
		_w36172_
	);
	LUT2 #(
		.INIT('h1)
	) name32126 (
		_w36171_,
		_w36172_,
		_w36173_
	);
	LUT2 #(
		.INIT('h1)
	) name32127 (
		\sport0_regs_MWORDreg_DO_reg[10]/NET0131 ,
		_w18231_,
		_w36174_
	);
	LUT2 #(
		.INIT('h4)
	) name32128 (
		_w12743_,
		_w19015_,
		_w36175_
	);
	LUT2 #(
		.INIT('h1)
	) name32129 (
		_w36174_,
		_w36175_,
		_w36176_
	);
	LUT2 #(
		.INIT('h8)
	) name32130 (
		_w11265_,
		_w18652_,
		_w36177_
	);
	LUT2 #(
		.INIT('h2)
	) name32131 (
		\sport0_regs_FSDIVreg_DO_reg[7]/NET0131 ,
		_w18652_,
		_w36178_
	);
	LUT2 #(
		.INIT('h1)
	) name32132 (
		_w18232_,
		_w36178_,
		_w36179_
	);
	LUT2 #(
		.INIT('h4)
	) name32133 (
		_w36177_,
		_w36179_,
		_w36180_
	);
	LUT2 #(
		.INIT('h8)
	) name32134 (
		_w11525_,
		_w18652_,
		_w36181_
	);
	LUT2 #(
		.INIT('h2)
	) name32135 (
		\sport0_regs_FSDIVreg_DO_reg[6]/NET0131 ,
		_w18652_,
		_w36182_
	);
	LUT2 #(
		.INIT('h1)
	) name32136 (
		_w18232_,
		_w36182_,
		_w36183_
	);
	LUT2 #(
		.INIT('h4)
	) name32137 (
		_w36181_,
		_w36183_,
		_w36184_
	);
	LUT2 #(
		.INIT('h8)
	) name32138 (
		_w10911_,
		_w18652_,
		_w36185_
	);
	LUT2 #(
		.INIT('h2)
	) name32139 (
		\sport0_regs_FSDIVreg_DO_reg[5]/NET0131 ,
		_w18652_,
		_w36186_
	);
	LUT2 #(
		.INIT('h1)
	) name32140 (
		_w18232_,
		_w36186_,
		_w36187_
	);
	LUT2 #(
		.INIT('h4)
	) name32141 (
		_w36185_,
		_w36187_,
		_w36188_
	);
	LUT2 #(
		.INIT('h8)
	) name32142 (
		_w10069_,
		_w18652_,
		_w36189_
	);
	LUT2 #(
		.INIT('h2)
	) name32143 (
		\sport0_regs_FSDIVreg_DO_reg[4]/NET0131 ,
		_w18652_,
		_w36190_
	);
	LUT2 #(
		.INIT('h1)
	) name32144 (
		_w18232_,
		_w36190_,
		_w36191_
	);
	LUT2 #(
		.INIT('h4)
	) name32145 (
		_w36189_,
		_w36191_,
		_w36192_
	);
	LUT2 #(
		.INIT('h8)
	) name32146 (
		_w8113_,
		_w18652_,
		_w36193_
	);
	LUT2 #(
		.INIT('h2)
	) name32147 (
		\sport0_regs_FSDIVreg_DO_reg[3]/NET0131 ,
		_w18652_,
		_w36194_
	);
	LUT2 #(
		.INIT('h1)
	) name32148 (
		_w18232_,
		_w36194_,
		_w36195_
	);
	LUT2 #(
		.INIT('h4)
	) name32149 (
		_w36193_,
		_w36195_,
		_w36196_
	);
	LUT2 #(
		.INIT('h8)
	) name32150 (
		_w8715_,
		_w18652_,
		_w36197_
	);
	LUT2 #(
		.INIT('h2)
	) name32151 (
		\sport0_regs_FSDIVreg_DO_reg[2]/NET0131 ,
		_w18652_,
		_w36198_
	);
	LUT2 #(
		.INIT('h1)
	) name32152 (
		_w18232_,
		_w36198_,
		_w36199_
	);
	LUT2 #(
		.INIT('h4)
	) name32153 (
		_w36197_,
		_w36199_,
		_w36200_
	);
	LUT2 #(
		.INIT('h8)
	) name32154 (
		_w9435_,
		_w18652_,
		_w36201_
	);
	LUT2 #(
		.INIT('h2)
	) name32155 (
		\sport0_regs_FSDIVreg_DO_reg[1]/NET0131 ,
		_w18652_,
		_w36202_
	);
	LUT2 #(
		.INIT('h1)
	) name32156 (
		_w18232_,
		_w36202_,
		_w36203_
	);
	LUT2 #(
		.INIT('h4)
	) name32157 (
		_w36201_,
		_w36203_,
		_w36204_
	);
	LUT2 #(
		.INIT('h8)
	) name32158 (
		_w7607_,
		_w18652_,
		_w36205_
	);
	LUT2 #(
		.INIT('h2)
	) name32159 (
		\sport0_regs_FSDIVreg_DO_reg[0]/NET0131 ,
		_w18652_,
		_w36206_
	);
	LUT2 #(
		.INIT('h1)
	) name32160 (
		_w18232_,
		_w36206_,
		_w36207_
	);
	LUT2 #(
		.INIT('h4)
	) name32161 (
		_w36205_,
		_w36207_,
		_w36208_
	);
	LUT2 #(
		.INIT('h8)
	) name32162 (
		_w7232_,
		_w7283_,
		_w36209_
	);
	LUT2 #(
		.INIT('h8)
	) name32163 (
		_w13762_,
		_w36209_,
		_w36210_
	);
	LUT2 #(
		.INIT('h4)
	) name32164 (
		_w25671_,
		_w36210_,
		_w36211_
	);
	LUT2 #(
		.INIT('h2)
	) name32165 (
		\PIO_out[6]_pad ,
		_w36211_,
		_w36212_
	);
	LUT2 #(
		.INIT('h8)
	) name32166 (
		_w11525_,
		_w36211_,
		_w36213_
	);
	LUT2 #(
		.INIT('h1)
	) name32167 (
		_w36212_,
		_w36213_,
		_w36214_
	);
	LUT2 #(
		.INIT('h2)
	) name32168 (
		\PIO_oe[6]_pad ,
		_w36214_,
		_w36215_
	);
	LUT2 #(
		.INIT('h4)
	) name32169 (
		\PIO_oe[6]_pad ,
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w36216_
	);
	LUT2 #(
		.INIT('h1)
	) name32170 (
		_w36215_,
		_w36216_,
		_w36217_
	);
	LUT2 #(
		.INIT('h4)
	) name32171 (
		_w25679_,
		_w36210_,
		_w36218_
	);
	LUT2 #(
		.INIT('h2)
	) name32172 (
		\PIO_out[4]_pad ,
		_w36218_,
		_w36219_
	);
	LUT2 #(
		.INIT('h8)
	) name32173 (
		_w10069_,
		_w36218_,
		_w36220_
	);
	LUT2 #(
		.INIT('h1)
	) name32174 (
		_w36219_,
		_w36220_,
		_w36221_
	);
	LUT2 #(
		.INIT('h2)
	) name32175 (
		\PIO_oe[4]_pad ,
		_w36221_,
		_w36222_
	);
	LUT2 #(
		.INIT('h4)
	) name32176 (
		\PIO_oe[4]_pad ,
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w36223_
	);
	LUT2 #(
		.INIT('h1)
	) name32177 (
		_w36222_,
		_w36223_,
		_w36224_
	);
	LUT2 #(
		.INIT('h4)
	) name32178 (
		_w25666_,
		_w36210_,
		_w36225_
	);
	LUT2 #(
		.INIT('h2)
	) name32179 (
		\PIO_out[2]_pad ,
		_w36225_,
		_w36226_
	);
	LUT2 #(
		.INIT('h8)
	) name32180 (
		_w8715_,
		_w36225_,
		_w36227_
	);
	LUT2 #(
		.INIT('h1)
	) name32181 (
		_w36226_,
		_w36227_,
		_w36228_
	);
	LUT2 #(
		.INIT('h2)
	) name32182 (
		\PIO_oe[2]_pad ,
		_w36228_,
		_w36229_
	);
	LUT2 #(
		.INIT('h4)
	) name32183 (
		\PIO_oe[2]_pad ,
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w36230_
	);
	LUT2 #(
		.INIT('h1)
	) name32184 (
		_w36229_,
		_w36230_,
		_w36231_
	);
	LUT2 #(
		.INIT('h4)
	) name32185 (
		_w25661_,
		_w36210_,
		_w36232_
	);
	LUT2 #(
		.INIT('h2)
	) name32186 (
		\PIO_out[10]_pad ,
		_w36232_,
		_w36233_
	);
	LUT2 #(
		.INIT('h8)
	) name32187 (
		_w12688_,
		_w36232_,
		_w36234_
	);
	LUT2 #(
		.INIT('h1)
	) name32188 (
		_w36233_,
		_w36234_,
		_w36235_
	);
	LUT2 #(
		.INIT('h2)
	) name32189 (
		\PIO_oe[10]_pad ,
		_w36235_,
		_w36236_
	);
	LUT2 #(
		.INIT('h4)
	) name32190 (
		\PIO_oe[10]_pad ,
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w36237_
	);
	LUT2 #(
		.INIT('h1)
	) name32191 (
		_w36236_,
		_w36237_,
		_w36238_
	);
	LUT2 #(
		.INIT('h4)
	) name32192 (
		_w25656_,
		_w36210_,
		_w36239_
	);
	LUT2 #(
		.INIT('h2)
	) name32193 (
		\PIO_out[0]_pad ,
		_w36239_,
		_w36240_
	);
	LUT2 #(
		.INIT('h8)
	) name32194 (
		_w7607_,
		_w36239_,
		_w36241_
	);
	LUT2 #(
		.INIT('h1)
	) name32195 (
		_w36240_,
		_w36241_,
		_w36242_
	);
	LUT2 #(
		.INIT('h2)
	) name32196 (
		\PIO_oe[0]_pad ,
		_w36242_,
		_w36243_
	);
	LUT2 #(
		.INIT('h4)
	) name32197 (
		\PIO_oe[0]_pad ,
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w36244_
	);
	LUT2 #(
		.INIT('h1)
	) name32198 (
		_w36243_,
		_w36244_,
		_w36245_
	);
	LUT2 #(
		.INIT('h2)
	) name32199 (
		\sice_DMR1_reg[8]/NET0131 ,
		_w27904_,
		_w36246_
	);
	LUT2 #(
		.INIT('h8)
	) name32200 (
		\sice_SPC_reg[14]/P0001 ,
		_w27904_,
		_w36247_
	);
	LUT2 #(
		.INIT('h1)
	) name32201 (
		_w36246_,
		_w36247_,
		_w36248_
	);
	LUT2 #(
		.INIT('h8)
	) name32202 (
		\core_c_psq_T_IRQL0p_reg/P0001 ,
		\core_c_psq_irql0_de_OUT_reg/P0001 ,
		_w36249_
	);
	LUT2 #(
		.INIT('h1)
	) name32203 (
		\core_c_psq_T_IRQL0p_reg/P0001 ,
		\core_c_psq_irql0_de_OUT_reg/P0001 ,
		_w36250_
	);
	LUT2 #(
		.INIT('h2)
	) name32204 (
		\core_c_psq_irql0_de_IN_syn_reg/P0001 ,
		_w36250_,
		_w36251_
	);
	LUT2 #(
		.INIT('h1)
	) name32205 (
		_w36249_,
		_w36251_,
		_w36252_
	);
	LUT2 #(
		.INIT('h4)
	) name32206 (
		_w25651_,
		_w36210_,
		_w36253_
	);
	LUT2 #(
		.INIT('h2)
	) name32207 (
		\PIO_out[9]_pad ,
		_w36253_,
		_w36254_
	);
	LUT2 #(
		.INIT('h8)
	) name32208 (
		_w7340_,
		_w36253_,
		_w36255_
	);
	LUT2 #(
		.INIT('h1)
	) name32209 (
		_w36254_,
		_w36255_,
		_w36256_
	);
	LUT2 #(
		.INIT('h2)
	) name32210 (
		\PIO_oe[9]_pad ,
		_w36256_,
		_w36257_
	);
	LUT2 #(
		.INIT('h4)
	) name32211 (
		\PIO_oe[9]_pad ,
		\pio_PIO_RES_reg[9]/NET0131 ,
		_w36258_
	);
	LUT2 #(
		.INIT('h1)
	) name32212 (
		_w36257_,
		_w36258_,
		_w36259_
	);
	LUT2 #(
		.INIT('h2)
	) name32213 (
		\PIO_out[8]_pad ,
		_w36253_,
		_w36260_
	);
	LUT2 #(
		.INIT('h8)
	) name32214 (
		_w9178_,
		_w36253_,
		_w36261_
	);
	LUT2 #(
		.INIT('h1)
	) name32215 (
		_w36260_,
		_w36261_,
		_w36262_
	);
	LUT2 #(
		.INIT('h2)
	) name32216 (
		\PIO_oe[8]_pad ,
		_w36262_,
		_w36263_
	);
	LUT2 #(
		.INIT('h4)
	) name32217 (
		\PIO_oe[8]_pad ,
		\pio_PIO_RES_reg[8]/NET0131 ,
		_w36264_
	);
	LUT2 #(
		.INIT('h1)
	) name32218 (
		_w36263_,
		_w36264_,
		_w36265_
	);
	LUT2 #(
		.INIT('h2)
	) name32219 (
		\PIO_out[5]_pad ,
		_w36218_,
		_w36266_
	);
	LUT2 #(
		.INIT('h8)
	) name32220 (
		_w10911_,
		_w36218_,
		_w36267_
	);
	LUT2 #(
		.INIT('h1)
	) name32221 (
		_w36266_,
		_w36267_,
		_w36268_
	);
	LUT2 #(
		.INIT('h2)
	) name32222 (
		\PIO_oe[5]_pad ,
		_w36268_,
		_w36269_
	);
	LUT2 #(
		.INIT('h4)
	) name32223 (
		\PIO_oe[5]_pad ,
		\pio_PIO_RES_reg[5]/NET0131 ,
		_w36270_
	);
	LUT2 #(
		.INIT('h1)
	) name32224 (
		_w36269_,
		_w36270_,
		_w36271_
	);
	LUT2 #(
		.INIT('h2)
	) name32225 (
		\PIO_out[7]_pad ,
		_w36211_,
		_w36272_
	);
	LUT2 #(
		.INIT('h8)
	) name32226 (
		_w11265_,
		_w36211_,
		_w36273_
	);
	LUT2 #(
		.INIT('h1)
	) name32227 (
		_w36272_,
		_w36273_,
		_w36274_
	);
	LUT2 #(
		.INIT('h2)
	) name32228 (
		\PIO_oe[7]_pad ,
		_w36274_,
		_w36275_
	);
	LUT2 #(
		.INIT('h4)
	) name32229 (
		\PIO_oe[7]_pad ,
		\pio_PIO_RES_reg[7]/NET0131 ,
		_w36276_
	);
	LUT2 #(
		.INIT('h1)
	) name32230 (
		_w36275_,
		_w36276_,
		_w36277_
	);
	LUT2 #(
		.INIT('h2)
	) name32231 (
		\PIO_out[3]_pad ,
		_w36225_,
		_w36278_
	);
	LUT2 #(
		.INIT('h8)
	) name32232 (
		_w8113_,
		_w36225_,
		_w36279_
	);
	LUT2 #(
		.INIT('h1)
	) name32233 (
		_w36278_,
		_w36279_,
		_w36280_
	);
	LUT2 #(
		.INIT('h2)
	) name32234 (
		\PIO_oe[3]_pad ,
		_w36280_,
		_w36281_
	);
	LUT2 #(
		.INIT('h4)
	) name32235 (
		\PIO_oe[3]_pad ,
		\pio_PIO_RES_reg[3]/NET0131 ,
		_w36282_
	);
	LUT2 #(
		.INIT('h1)
	) name32236 (
		_w36281_,
		_w36282_,
		_w36283_
	);
	LUT2 #(
		.INIT('h2)
	) name32237 (
		\PIO_out[1]_pad ,
		_w36239_,
		_w36284_
	);
	LUT2 #(
		.INIT('h8)
	) name32238 (
		_w9435_,
		_w36239_,
		_w36285_
	);
	LUT2 #(
		.INIT('h1)
	) name32239 (
		_w36284_,
		_w36285_,
		_w36286_
	);
	LUT2 #(
		.INIT('h2)
	) name32240 (
		\PIO_oe[1]_pad ,
		_w36286_,
		_w36287_
	);
	LUT2 #(
		.INIT('h4)
	) name32241 (
		\PIO_oe[1]_pad ,
		\pio_PIO_RES_reg[1]/NET0131 ,
		_w36288_
	);
	LUT2 #(
		.INIT('h1)
	) name32242 (
		_w36287_,
		_w36288_,
		_w36289_
	);
	LUT2 #(
		.INIT('h2)
	) name32243 (
		\sice_SPC_reg[7]/P0001 ,
		_w26297_,
		_w36290_
	);
	LUT2 #(
		.INIT('h8)
	) name32244 (
		\sice_SPC_reg[6]/P0001 ,
		_w34825_,
		_w36291_
	);
	LUT2 #(
		.INIT('h2)
	) name32245 (
		\sice_SPC_reg[8]/P0001 ,
		_w34825_,
		_w36292_
	);
	LUT2 #(
		.INIT('h1)
	) name32246 (
		_w36291_,
		_w36292_,
		_w36293_
	);
	LUT2 #(
		.INIT('h4)
	) name32247 (
		_w34827_,
		_w36293_,
		_w36294_
	);
	LUT2 #(
		.INIT('h8)
	) name32248 (
		\sice_DMR1_reg[1]/NET0131 ,
		_w27903_,
		_w36295_
	);
	LUT2 #(
		.INIT('h8)
	) name32249 (
		\sice_IMR2_reg[1]/NET0131 ,
		_w25034_,
		_w36296_
	);
	LUT2 #(
		.INIT('h8)
	) name32250 (
		\sice_IBR1_reg[1]/P0001 ,
		_w34831_,
		_w36297_
	);
	LUT2 #(
		.INIT('h8)
	) name32251 (
		\core_c_dec_IR_reg[7]/NET0131 ,
		_w28203_,
		_w36298_
	);
	LUT2 #(
		.INIT('h8)
	) name32252 (
		\sice_DMR2_reg[1]/NET0131 ,
		_w25025_,
		_w36299_
	);
	LUT2 #(
		.INIT('h8)
	) name32253 (
		\sice_DBR2_reg[2]/P0001 ,
		_w25012_,
		_w36300_
	);
	LUT2 #(
		.INIT('h8)
	) name32254 (
		\sice_idr0_reg_DO_reg[7]/P0001 ,
		_w26968_,
		_w36301_
	);
	LUT2 #(
		.INIT('h8)
	) name32255 (
		\sice_IBR2_reg[1]/P0001 ,
		_w25074_,
		_w36302_
	);
	LUT2 #(
		.INIT('h8)
	) name32256 (
		\sice_DBR1_reg[2]/P0001 ,
		_w25054_,
		_w36303_
	);
	LUT2 #(
		.INIT('h8)
	) name32257 (
		\sice_IMR1_reg[1]/NET0131 ,
		_w34846_,
		_w36304_
	);
	LUT2 #(
		.INIT('h8)
	) name32258 (
		\sice_IIRC_reg[7]/NET0131 ,
		_w24267_,
		_w36305_
	);
	LUT2 #(
		.INIT('h8)
	) name32259 (
		\sice_ICYC_reg[7]/NET0131 ,
		_w23409_,
		_w36306_
	);
	LUT2 #(
		.INIT('h1)
	) name32260 (
		_w36295_,
		_w36296_,
		_w36307_
	);
	LUT2 #(
		.INIT('h1)
	) name32261 (
		_w36297_,
		_w36298_,
		_w36308_
	);
	LUT2 #(
		.INIT('h1)
	) name32262 (
		_w36299_,
		_w36300_,
		_w36309_
	);
	LUT2 #(
		.INIT('h1)
	) name32263 (
		_w36301_,
		_w36302_,
		_w36310_
	);
	LUT2 #(
		.INIT('h1)
	) name32264 (
		_w36303_,
		_w36304_,
		_w36311_
	);
	LUT2 #(
		.INIT('h1)
	) name32265 (
		_w36305_,
		_w36306_,
		_w36312_
	);
	LUT2 #(
		.INIT('h8)
	) name32266 (
		_w36311_,
		_w36312_,
		_w36313_
	);
	LUT2 #(
		.INIT('h8)
	) name32267 (
		_w36309_,
		_w36310_,
		_w36314_
	);
	LUT2 #(
		.INIT('h8)
	) name32268 (
		_w36307_,
		_w36308_,
		_w36315_
	);
	LUT2 #(
		.INIT('h8)
	) name32269 (
		_w36314_,
		_w36315_,
		_w36316_
	);
	LUT2 #(
		.INIT('h8)
	) name32270 (
		_w36313_,
		_w36316_,
		_w36317_
	);
	LUT2 #(
		.INIT('h8)
	) name32271 (
		_w34827_,
		_w36317_,
		_w36318_
	);
	LUT2 #(
		.INIT('h2)
	) name32272 (
		_w26297_,
		_w36294_,
		_w36319_
	);
	LUT2 #(
		.INIT('h4)
	) name32273 (
		_w36318_,
		_w36319_,
		_w36320_
	);
	LUT2 #(
		.INIT('h1)
	) name32274 (
		_w36290_,
		_w36320_,
		_w36321_
	);
	LUT2 #(
		.INIT('h2)
	) name32275 (
		\sice_SPC_reg[8]/P0001 ,
		_w26297_,
		_w36322_
	);
	LUT2 #(
		.INIT('h8)
	) name32276 (
		\sice_SPC_reg[7]/P0001 ,
		_w34825_,
		_w36323_
	);
	LUT2 #(
		.INIT('h2)
	) name32277 (
		\sice_SPC_reg[9]/P0001 ,
		_w34825_,
		_w36324_
	);
	LUT2 #(
		.INIT('h1)
	) name32278 (
		_w36323_,
		_w36324_,
		_w36325_
	);
	LUT2 #(
		.INIT('h4)
	) name32279 (
		_w34827_,
		_w36325_,
		_w36326_
	);
	LUT2 #(
		.INIT('h8)
	) name32280 (
		\sice_DMR1_reg[2]/NET0131 ,
		_w27903_,
		_w36327_
	);
	LUT2 #(
		.INIT('h8)
	) name32281 (
		\sice_IMR2_reg[2]/NET0131 ,
		_w25034_,
		_w36328_
	);
	LUT2 #(
		.INIT('h8)
	) name32282 (
		\sice_IBR1_reg[2]/P0001 ,
		_w34831_,
		_w36329_
	);
	LUT2 #(
		.INIT('h8)
	) name32283 (
		\core_c_dec_IR_reg[8]/NET0131 ,
		_w28203_,
		_w36330_
	);
	LUT2 #(
		.INIT('h8)
	) name32284 (
		\sice_DMR2_reg[2]/NET0131 ,
		_w25025_,
		_w36331_
	);
	LUT2 #(
		.INIT('h8)
	) name32285 (
		\sice_DBR2_reg[3]/P0001 ,
		_w25012_,
		_w36332_
	);
	LUT2 #(
		.INIT('h8)
	) name32286 (
		\sice_idr0_reg_DO_reg[8]/P0001 ,
		_w26968_,
		_w36333_
	);
	LUT2 #(
		.INIT('h8)
	) name32287 (
		\sice_IBR2_reg[2]/P0001 ,
		_w25074_,
		_w36334_
	);
	LUT2 #(
		.INIT('h8)
	) name32288 (
		\sice_DBR1_reg[3]/P0001 ,
		_w25054_,
		_w36335_
	);
	LUT2 #(
		.INIT('h8)
	) name32289 (
		\sice_IMR1_reg[2]/NET0131 ,
		_w34846_,
		_w36336_
	);
	LUT2 #(
		.INIT('h8)
	) name32290 (
		\sice_IIRC_reg[8]/NET0131 ,
		_w24267_,
		_w36337_
	);
	LUT2 #(
		.INIT('h8)
	) name32291 (
		\sice_ICYC_reg[8]/NET0131 ,
		_w23409_,
		_w36338_
	);
	LUT2 #(
		.INIT('h1)
	) name32292 (
		_w36327_,
		_w36328_,
		_w36339_
	);
	LUT2 #(
		.INIT('h1)
	) name32293 (
		_w36329_,
		_w36330_,
		_w36340_
	);
	LUT2 #(
		.INIT('h1)
	) name32294 (
		_w36331_,
		_w36332_,
		_w36341_
	);
	LUT2 #(
		.INIT('h1)
	) name32295 (
		_w36333_,
		_w36334_,
		_w36342_
	);
	LUT2 #(
		.INIT('h1)
	) name32296 (
		_w36335_,
		_w36336_,
		_w36343_
	);
	LUT2 #(
		.INIT('h1)
	) name32297 (
		_w36337_,
		_w36338_,
		_w36344_
	);
	LUT2 #(
		.INIT('h8)
	) name32298 (
		_w36343_,
		_w36344_,
		_w36345_
	);
	LUT2 #(
		.INIT('h8)
	) name32299 (
		_w36341_,
		_w36342_,
		_w36346_
	);
	LUT2 #(
		.INIT('h8)
	) name32300 (
		_w36339_,
		_w36340_,
		_w36347_
	);
	LUT2 #(
		.INIT('h8)
	) name32301 (
		_w36346_,
		_w36347_,
		_w36348_
	);
	LUT2 #(
		.INIT('h8)
	) name32302 (
		_w36345_,
		_w36348_,
		_w36349_
	);
	LUT2 #(
		.INIT('h8)
	) name32303 (
		_w34827_,
		_w36349_,
		_w36350_
	);
	LUT2 #(
		.INIT('h2)
	) name32304 (
		_w26297_,
		_w36326_,
		_w36351_
	);
	LUT2 #(
		.INIT('h4)
	) name32305 (
		_w36350_,
		_w36351_,
		_w36352_
	);
	LUT2 #(
		.INIT('h1)
	) name32306 (
		_w36322_,
		_w36352_,
		_w36353_
	);
	LUT2 #(
		.INIT('h8)
	) name32307 (
		\idma_WRcyc_reg/NET0131 ,
		_w32463_,
		_w36354_
	);
	LUT2 #(
		.INIT('h1)
	) name32308 (
		_w20384_,
		_w36354_,
		_w36355_
	);
	LUT2 #(
		.INIT('h2)
	) name32309 (
		\PIO_out[11]_pad ,
		_w36232_,
		_w36356_
	);
	LUT2 #(
		.INIT('h8)
	) name32310 (
		_w12743_,
		_w36232_,
		_w36357_
	);
	LUT2 #(
		.INIT('h1)
	) name32311 (
		_w36356_,
		_w36357_,
		_w36358_
	);
	LUT2 #(
		.INIT('h2)
	) name32312 (
		\PIO_oe[11]_pad ,
		_w36358_,
		_w36359_
	);
	LUT2 #(
		.INIT('h4)
	) name32313 (
		\PIO_oe[11]_pad ,
		\pio_PIO_RES_reg[11]/NET0131 ,
		_w36360_
	);
	LUT2 #(
		.INIT('h1)
	) name32314 (
		_w36359_,
		_w36360_,
		_w36361_
	);
	LUT2 #(
		.INIT('h2)
	) name32315 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[10]/P0001 ,
		_w18848_,
		_w36362_
	);
	LUT2 #(
		.INIT('h8)
	) name32316 (
		_w20398_,
		_w21422_,
		_w36363_
	);
	LUT2 #(
		.INIT('h8)
	) name32317 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w18847_,
		_w36364_
	);
	LUT2 #(
		.INIT('h8)
	) name32318 (
		_w5123_,
		_w36364_,
		_w36365_
	);
	LUT2 #(
		.INIT('h1)
	) name32319 (
		_w36362_,
		_w36365_,
		_w36366_
	);
	LUT2 #(
		.INIT('h4)
	) name32320 (
		_w36363_,
		_w36366_,
		_w36367_
	);
	LUT2 #(
		.INIT('h1)
	) name32321 (
		_w5951_,
		_w6988_,
		_w36368_
	);
	LUT2 #(
		.INIT('h1)
	) name32322 (
		_w11738_,
		_w36368_,
		_w36369_
	);
	LUT2 #(
		.INIT('h2)
	) name32323 (
		_w11764_,
		_w36369_,
		_w36370_
	);
	LUT2 #(
		.INIT('h8)
	) name32324 (
		_w9513_,
		_w12197_,
		_w36371_
	);
	LUT2 #(
		.INIT('h1)
	) name32325 (
		_w11735_,
		_w36371_,
		_w36372_
	);
	LUT2 #(
		.INIT('h1)
	) name32326 (
		_w36370_,
		_w36372_,
		_w36373_
	);
	LUT2 #(
		.INIT('h8)
	) name32327 (
		_w23032_,
		_w34846_,
		_w36374_
	);
	LUT2 #(
		.INIT('h2)
	) name32328 (
		\core_eu_em_mac_em_dec_emcorepi_DO_reg[1]/P0001 ,
		_w18848_,
		_w36375_
	);
	LUT2 #(
		.INIT('h2)
	) name32329 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w36376_
	);
	LUT2 #(
		.INIT('h1)
	) name32330 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w36376_,
		_w36377_
	);
	LUT2 #(
		.INIT('h8)
	) name32331 (
		_w18848_,
		_w36377_,
		_w36378_
	);
	LUT2 #(
		.INIT('h1)
	) name32332 (
		_w36375_,
		_w36378_,
		_w36379_
	);
	LUT2 #(
		.INIT('h2)
	) name32333 (
		\core_c_psq_Iact_E_reg[2]/NET0131 ,
		_w19477_,
		_w36380_
	);
	LUT2 #(
		.INIT('h2)
	) name32334 (
		_w19477_,
		_w33213_,
		_w36381_
	);
	LUT2 #(
		.INIT('h8)
	) name32335 (
		_w33205_,
		_w33216_,
		_w36382_
	);
	LUT2 #(
		.INIT('h8)
	) name32336 (
		_w36381_,
		_w36382_,
		_w36383_
	);
	LUT2 #(
		.INIT('h1)
	) name32337 (
		_w36380_,
		_w36383_,
		_w36384_
	);
	LUT2 #(
		.INIT('h2)
	) name32338 (
		\clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131 ,
		_w31521_,
		_w36385_
	);
	LUT2 #(
		.INIT('h4)
	) name32339 (
		\clkc_ckSTDCLK_STDCLK_reg_Q_reg/NET0131 ,
		_w31521_,
		_w36386_
	);
	LUT2 #(
		.INIT('h1)
	) name32340 (
		_w36385_,
		_w36386_,
		_w36387_
	);
	LUT2 #(
		.INIT('h8)
	) name32341 (
		_w23032_,
		_w34831_,
		_w36388_
	);
	LUT2 #(
		.INIT('h8)
	) name32342 (
		\sport1_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w23274_,
		_w36389_
	);
	LUT2 #(
		.INIT('h4)
	) name32343 (
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		_w23726_,
		_w36390_
	);
	LUT2 #(
		.INIT('h4)
	) name32344 (
		\sport1_txctl_Wcnt_reg[1]/NET0131 ,
		_w36390_,
		_w36391_
	);
	LUT2 #(
		.INIT('h4)
	) name32345 (
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		_w36391_,
		_w36392_
	);
	LUT2 #(
		.INIT('h4)
	) name32346 (
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		_w36392_,
		_w36393_
	);
	LUT2 #(
		.INIT('h4)
	) name32347 (
		\sport1_txctl_Wcnt_reg[4]/NET0131 ,
		_w36393_,
		_w36394_
	);
	LUT2 #(
		.INIT('h4)
	) name32348 (
		\sport1_txctl_Wcnt_reg[5]/NET0131 ,
		_w36394_,
		_w36395_
	);
	LUT2 #(
		.INIT('h4)
	) name32349 (
		\sport1_txctl_Wcnt_reg[6]/NET0131 ,
		_w36395_,
		_w36396_
	);
	LUT2 #(
		.INIT('h1)
	) name32350 (
		_w23274_,
		_w36396_,
		_w36397_
	);
	LUT2 #(
		.INIT('h8)
	) name32351 (
		\sport1_txctl_Wcnt_reg[7]/NET0131 ,
		_w36397_,
		_w36398_
	);
	LUT2 #(
		.INIT('h1)
	) name32352 (
		_w36389_,
		_w36398_,
		_w36399_
	);
	LUT2 #(
		.INIT('h2)
	) name32353 (
		\sport1_txctl_Wcnt_reg[5]/NET0131 ,
		_w36394_,
		_w36400_
	);
	LUT2 #(
		.INIT('h1)
	) name32354 (
		_w36395_,
		_w36400_,
		_w36401_
	);
	LUT2 #(
		.INIT('h4)
	) name32355 (
		_w23274_,
		_w36401_,
		_w36402_
	);
	LUT2 #(
		.INIT('h4)
	) name32356 (
		\sport1_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w23274_,
		_w36403_
	);
	LUT2 #(
		.INIT('h1)
	) name32357 (
		_w36402_,
		_w36403_,
		_w36404_
	);
	LUT2 #(
		.INIT('h8)
	) name32358 (
		\sport0_regs_MWORDreg_DO_reg[7]/NET0131 ,
		_w23286_,
		_w36405_
	);
	LUT2 #(
		.INIT('h4)
	) name32359 (
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		_w23744_,
		_w36406_
	);
	LUT2 #(
		.INIT('h4)
	) name32360 (
		\sport0_txctl_Wcnt_reg[1]/NET0131 ,
		_w36406_,
		_w36407_
	);
	LUT2 #(
		.INIT('h4)
	) name32361 (
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		_w36407_,
		_w36408_
	);
	LUT2 #(
		.INIT('h4)
	) name32362 (
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		_w36408_,
		_w36409_
	);
	LUT2 #(
		.INIT('h4)
	) name32363 (
		\sport0_txctl_Wcnt_reg[4]/NET0131 ,
		_w36409_,
		_w36410_
	);
	LUT2 #(
		.INIT('h4)
	) name32364 (
		\sport0_txctl_Wcnt_reg[5]/NET0131 ,
		_w36410_,
		_w36411_
	);
	LUT2 #(
		.INIT('h4)
	) name32365 (
		\sport0_txctl_Wcnt_reg[6]/NET0131 ,
		_w36411_,
		_w36412_
	);
	LUT2 #(
		.INIT('h1)
	) name32366 (
		_w23286_,
		_w36412_,
		_w36413_
	);
	LUT2 #(
		.INIT('h8)
	) name32367 (
		\sport0_txctl_Wcnt_reg[7]/NET0131 ,
		_w36413_,
		_w36414_
	);
	LUT2 #(
		.INIT('h1)
	) name32368 (
		_w36405_,
		_w36414_,
		_w36415_
	);
	LUT2 #(
		.INIT('h2)
	) name32369 (
		\sport0_txctl_Wcnt_reg[5]/NET0131 ,
		_w36410_,
		_w36416_
	);
	LUT2 #(
		.INIT('h1)
	) name32370 (
		_w36411_,
		_w36416_,
		_w36417_
	);
	LUT2 #(
		.INIT('h4)
	) name32371 (
		_w23286_,
		_w36417_,
		_w36418_
	);
	LUT2 #(
		.INIT('h4)
	) name32372 (
		\sport0_regs_MWORDreg_DO_reg[5]/NET0131 ,
		_w23286_,
		_w36419_
	);
	LUT2 #(
		.INIT('h1)
	) name32373 (
		_w36418_,
		_w36419_,
		_w36420_
	);
	LUT2 #(
		.INIT('h1)
	) name32374 (
		\idma_WRcnt_reg[2]/NET0131 ,
		_w20459_,
		_w36421_
	);
	LUT2 #(
		.INIT('h8)
	) name32375 (
		\idma_WRcnt_reg[2]/NET0131 ,
		_w20459_,
		_w36422_
	);
	LUT2 #(
		.INIT('h1)
	) name32376 (
		_w36421_,
		_w36422_,
		_w36423_
	);
	LUT2 #(
		.INIT('h1)
	) name32377 (
		_w20455_,
		_w36423_,
		_w36424_
	);
	LUT2 #(
		.INIT('h4)
	) name32378 (
		\memc_usysr_DO_reg[9]/NET0131 ,
		_w20455_,
		_w36425_
	);
	LUT2 #(
		.INIT('h1)
	) name32379 (
		_w36424_,
		_w36425_,
		_w36426_
	);
	LUT2 #(
		.INIT('h1)
	) name32380 (
		_w21137_,
		_w21138_,
		_w36427_
	);
	LUT2 #(
		.INIT('h1)
	) name32381 (
		_w4217_,
		_w36427_,
		_w36428_
	);
	LUT2 #(
		.INIT('h8)
	) name32382 (
		\core_c_dec_IRE_reg[4]/NET0131 ,
		\core_c_dec_Stkctl_Eg_reg/P0001 ,
		_w36429_
	);
	LUT2 #(
		.INIT('h1)
	) name32383 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w36429_,
		_w36430_
	);
	LUT2 #(
		.INIT('h2)
	) name32384 (
		\core_c_dec_RET_Ed_reg/P0001 ,
		_w4184_,
		_w36431_
	);
	LUT2 #(
		.INIT('h2)
	) name32385 (
		_w36430_,
		_w36431_,
		_w36432_
	);
	LUT2 #(
		.INIT('h4)
	) name32386 (
		_w4842_,
		_w36432_,
		_w36433_
	);
	LUT2 #(
		.INIT('h1)
	) name32387 (
		_w5950_,
		_w36433_,
		_w36434_
	);
	LUT2 #(
		.INIT('h4)
	) name32388 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w36434_,
		_w36435_
	);
	LUT2 #(
		.INIT('h1)
	) name32389 (
		\core_c_dec_Call_Ed_reg/P0001 ,
		\core_c_dec_RET_Ed_reg/P0001 ,
		_w36436_
	);
	LUT2 #(
		.INIT('h1)
	) name32390 (
		\core_c_psq_Eqend_Ed_reg/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w36437_
	);
	LUT2 #(
		.INIT('h8)
	) name32391 (
		_w36436_,
		_w36437_,
		_w36438_
	);
	LUT2 #(
		.INIT('h8)
	) name32392 (
		_w21134_,
		_w36438_,
		_w36439_
	);
	LUT2 #(
		.INIT('h8)
	) name32393 (
		_w36430_,
		_w36439_,
		_w36440_
	);
	LUT2 #(
		.INIT('h2)
	) name32394 (
		_w36435_,
		_w36440_,
		_w36441_
	);
	LUT2 #(
		.INIT('h1)
	) name32395 (
		_w36427_,
		_w36441_,
		_w36442_
	);
	LUT2 #(
		.INIT('h1)
	) name32396 (
		_w4208_,
		_w21137_,
		_w36443_
	);
	LUT2 #(
		.INIT('h1)
	) name32397 (
		_w36428_,
		_w36443_,
		_w36444_
	);
	LUT2 #(
		.INIT('h4)
	) name32398 (
		_w36442_,
		_w36444_,
		_w36445_
	);
	LUT2 #(
		.INIT('h2)
	) name32399 (
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w36445_,
		_w36446_
	);
	LUT2 #(
		.INIT('h4)
	) name32400 (
		\core_c_psq_pcstk_ptr_reg[3]/NET0131 ,
		_w36445_,
		_w36447_
	);
	LUT2 #(
		.INIT('h1)
	) name32401 (
		_w36446_,
		_w36447_,
		_w36448_
	);
	LUT2 #(
		.INIT('h1)
	) name32402 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		_w36442_,
		_w36449_
	);
	LUT2 #(
		.INIT('h8)
	) name32403 (
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		_w36427_,
		_w36450_
	);
	LUT2 #(
		.INIT('h1)
	) name32404 (
		_w36449_,
		_w36450_,
		_w36451_
	);
	LUT2 #(
		.INIT('h1)
	) name32405 (
		\core_c_psq_pcstk_ptr_reg[1]/NET0131 ,
		_w36427_,
		_w36452_
	);
	LUT2 #(
		.INIT('h1)
	) name32406 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		_w36452_,
		_w36453_
	);
	LUT2 #(
		.INIT('h1)
	) name32407 (
		_w36451_,
		_w36453_,
		_w36454_
	);
	LUT2 #(
		.INIT('h2)
	) name32408 (
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w36454_,
		_w36455_
	);
	LUT2 #(
		.INIT('h4)
	) name32409 (
		\core_c_psq_pcstk_ptr_reg[2]/NET0131 ,
		_w36454_,
		_w36456_
	);
	LUT2 #(
		.INIT('h1)
	) name32410 (
		_w36455_,
		_w36456_,
		_w36457_
	);
	LUT2 #(
		.INIT('h1)
	) name32411 (
		_w36450_,
		_w36452_,
		_w36458_
	);
	LUT2 #(
		.INIT('h2)
	) name32412 (
		_w36449_,
		_w36458_,
		_w36459_
	);
	LUT2 #(
		.INIT('h4)
	) name32413 (
		_w36449_,
		_w36458_,
		_w36460_
	);
	LUT2 #(
		.INIT('h1)
	) name32414 (
		_w36459_,
		_w36460_,
		_w36461_
	);
	LUT2 #(
		.INIT('h8)
	) name32415 (
		\core_c_psq_pcstk_ptr_reg[0]/NET0131 ,
		_w36442_,
		_w36462_
	);
	LUT2 #(
		.INIT('h1)
	) name32416 (
		_w36449_,
		_w36462_,
		_w36463_
	);
	LUT2 #(
		.INIT('h2)
	) name32417 (
		\core_c_psq_Iact_E_reg[1]/NET0131 ,
		_w19477_,
		_w36464_
	);
	LUT2 #(
		.INIT('h4)
	) name32418 (
		_w33204_,
		_w33210_,
		_w36465_
	);
	LUT2 #(
		.INIT('h8)
	) name32419 (
		_w33216_,
		_w36465_,
		_w36466_
	);
	LUT2 #(
		.INIT('h8)
	) name32420 (
		_w36381_,
		_w36466_,
		_w36467_
	);
	LUT2 #(
		.INIT('h1)
	) name32421 (
		_w36464_,
		_w36467_,
		_w36468_
	);
	LUT2 #(
		.INIT('h2)
	) name32422 (
		\core_c_psq_Iact_E_reg[0]/NET0131 ,
		_w19477_,
		_w36469_
	);
	LUT2 #(
		.INIT('h1)
	) name32423 (
		_w19488_,
		_w33212_,
		_w36470_
	);
	LUT2 #(
		.INIT('h4)
	) name32424 (
		_w19480_,
		_w36470_,
		_w36471_
	);
	LUT2 #(
		.INIT('h8)
	) name32425 (
		_w33218_,
		_w36471_,
		_w36472_
	);
	LUT2 #(
		.INIT('h8)
	) name32426 (
		_w19494_,
		_w36472_,
		_w36473_
	);
	LUT2 #(
		.INIT('h8)
	) name32427 (
		_w33211_,
		_w36473_,
		_w36474_
	);
	LUT2 #(
		.INIT('h8)
	) name32428 (
		_w19487_,
		_w36474_,
		_w36475_
	);
	LUT2 #(
		.INIT('h1)
	) name32429 (
		_w36469_,
		_w36475_,
		_w36476_
	);
	LUT2 #(
		.INIT('h8)
	) name32430 (
		\core_c_dec_MTIMASK_Eg_reg/P0001 ,
		_w4118_,
		_w36477_
	);
	LUT2 #(
		.INIT('h4)
	) name32431 (
		_w31998_,
		_w35572_,
		_w36478_
	);
	LUT2 #(
		.INIT('h1)
	) name32432 (
		_w36477_,
		_w36478_,
		_w36479_
	);
	LUT2 #(
		.INIT('h8)
	) name32433 (
		\core_c_dec_MFTX1_E_reg/P0001 ,
		_w4117_,
		_w36480_
	);
	LUT2 #(
		.INIT('h8)
	) name32434 (
		_w25734_,
		_w34556_,
		_w36481_
	);
	LUT2 #(
		.INIT('h8)
	) name32435 (
		_w32024_,
		_w36481_,
		_w36482_
	);
	LUT2 #(
		.INIT('h1)
	) name32436 (
		_w36480_,
		_w36482_,
		_w36483_
	);
	LUT2 #(
		.INIT('h8)
	) name32437 (
		\core_c_dec_MFTX0_E_reg/P0001 ,
		_w4117_,
		_w36484_
	);
	LUT2 #(
		.INIT('h8)
	) name32438 (
		_w31266_,
		_w32023_,
		_w36485_
	);
	LUT2 #(
		.INIT('h8)
	) name32439 (
		_w26100_,
		_w36485_,
		_w36486_
	);
	LUT2 #(
		.INIT('h1)
	) name32440 (
		_w36484_,
		_w36486_,
		_w36487_
	);
	LUT2 #(
		.INIT('h8)
	) name32441 (
		\core_c_dec_MFSSTAT_E_reg/P0001 ,
		_w4117_,
		_w36488_
	);
	LUT2 #(
		.INIT('h8)
	) name32442 (
		_w31271_,
		_w36481_,
		_w36489_
	);
	LUT2 #(
		.INIT('h1)
	) name32443 (
		_w36488_,
		_w36489_,
		_w36490_
	);
	LUT2 #(
		.INIT('h8)
	) name32444 (
		\core_c_dec_MFRX1_E_reg/P0001 ,
		_w4117_,
		_w36491_
	);
	LUT2 #(
		.INIT('h4)
	) name32445 (
		_w4117_,
		_w34038_,
		_w36492_
	);
	LUT2 #(
		.INIT('h8)
	) name32446 (
		_w31264_,
		_w36492_,
		_w36493_
	);
	LUT2 #(
		.INIT('h1)
	) name32447 (
		_w36491_,
		_w36493_,
		_w36494_
	);
	LUT2 #(
		.INIT('h8)
	) name32448 (
		\core_c_dec_MFRX0_E_reg/P0001 ,
		_w4117_,
		_w36495_
	);
	LUT2 #(
		.INIT('h8)
	) name32449 (
		_w25729_,
		_w36485_,
		_w36496_
	);
	LUT2 #(
		.INIT('h1)
	) name32450 (
		_w36495_,
		_w36496_,
		_w36497_
	);
	LUT2 #(
		.INIT('h1)
	) name32451 (
		_w4117_,
		_w33278_,
		_w36498_
	);
	LUT2 #(
		.INIT('h4)
	) name32452 (
		\core_c_dec_MFPMOVL_E_reg/P0001 ,
		_w4117_,
		_w36499_
	);
	LUT2 #(
		.INIT('h1)
	) name32453 (
		_w36498_,
		_w36499_,
		_w36500_
	);
	LUT2 #(
		.INIT('h8)
	) name32454 (
		\core_c_dec_MFMreg_E_reg[7]/P0001 ,
		_w4117_,
		_w36501_
	);
	LUT2 #(
		.INIT('h8)
	) name32455 (
		_w26100_,
		_w34042_,
		_w36502_
	);
	LUT2 #(
		.INIT('h1)
	) name32456 (
		_w36501_,
		_w36502_,
		_w36503_
	);
	LUT2 #(
		.INIT('h8)
	) name32457 (
		\core_c_dec_MFMreg_E_reg[6]/P0001 ,
		_w4117_,
		_w36504_
	);
	LUT2 #(
		.INIT('h8)
	) name32458 (
		_w25729_,
		_w34042_,
		_w36505_
	);
	LUT2 #(
		.INIT('h1)
	) name32459 (
		_w36504_,
		_w36505_,
		_w36506_
	);
	LUT2 #(
		.INIT('h8)
	) name32460 (
		_w26100_,
		_w31978_,
		_w36507_
	);
	LUT2 #(
		.INIT('h8)
	) name32461 (
		_w34030_,
		_w36507_,
		_w36508_
	);
	LUT2 #(
		.INIT('h8)
	) name32462 (
		\core_c_dec_MFMreg_E_reg[5]/P0001 ,
		_w4117_,
		_w36509_
	);
	LUT2 #(
		.INIT('h1)
	) name32463 (
		_w36508_,
		_w36509_,
		_w36510_
	);
	LUT2 #(
		.INIT('h8)
	) name32464 (
		\core_c_dec_MFMreg_E_reg[4]/P0001 ,
		_w4117_,
		_w36511_
	);
	LUT2 #(
		.INIT('h8)
	) name32465 (
		_w34030_,
		_w35757_,
		_w36512_
	);
	LUT2 #(
		.INIT('h1)
	) name32466 (
		_w36511_,
		_w36512_,
		_w36513_
	);
	LUT2 #(
		.INIT('h8)
	) name32467 (
		\core_c_dec_MFMreg_E_reg[3]/P0001 ,
		_w4117_,
		_w36514_
	);
	LUT2 #(
		.INIT('h2)
	) name32468 (
		_w6091_,
		_w31263_,
		_w36515_
	);
	LUT2 #(
		.INIT('h8)
	) name32469 (
		_w19301_,
		_w31966_,
		_w36516_
	);
	LUT2 #(
		.INIT('h4)
	) name32470 (
		_w4117_,
		_w36516_,
		_w36517_
	);
	LUT2 #(
		.INIT('h8)
	) name32471 (
		_w36515_,
		_w36517_,
		_w36518_
	);
	LUT2 #(
		.INIT('h1)
	) name32472 (
		_w36514_,
		_w36518_,
		_w36519_
	);
	LUT2 #(
		.INIT('h8)
	) name32473 (
		\core_c_dec_MFMreg_E_reg[2]/P0001 ,
		_w4117_,
		_w36520_
	);
	LUT2 #(
		.INIT('h8)
	) name32474 (
		_w19298_,
		_w31966_,
		_w36521_
	);
	LUT2 #(
		.INIT('h4)
	) name32475 (
		_w4117_,
		_w36521_,
		_w36522_
	);
	LUT2 #(
		.INIT('h8)
	) name32476 (
		_w36515_,
		_w36522_,
		_w36523_
	);
	LUT2 #(
		.INIT('h1)
	) name32477 (
		_w36520_,
		_w36523_,
		_w36524_
	);
	LUT2 #(
		.INIT('h8)
	) name32478 (
		\core_c_dec_MFMreg_E_reg[1]/P0001 ,
		_w4117_,
		_w36525_
	);
	LUT2 #(
		.INIT('h8)
	) name32479 (
		_w19267_,
		_w31966_,
		_w36526_
	);
	LUT2 #(
		.INIT('h4)
	) name32480 (
		_w4117_,
		_w36526_,
		_w36527_
	);
	LUT2 #(
		.INIT('h8)
	) name32481 (
		_w36515_,
		_w36527_,
		_w36528_
	);
	LUT2 #(
		.INIT('h1)
	) name32482 (
		_w36525_,
		_w36528_,
		_w36529_
	);
	LUT2 #(
		.INIT('h8)
	) name32483 (
		\core_c_dec_MFMreg_E_reg[0]/P0001 ,
		_w4117_,
		_w36530_
	);
	LUT2 #(
		.INIT('h8)
	) name32484 (
		_w19270_,
		_w31973_,
		_w36531_
	);
	LUT2 #(
		.INIT('h8)
	) name32485 (
		_w25852_,
		_w36531_,
		_w36532_
	);
	LUT2 #(
		.INIT('h1)
	) name32486 (
		_w36530_,
		_w36532_,
		_w36533_
	);
	LUT2 #(
		.INIT('h8)
	) name32487 (
		\core_c_dec_MFMSTAT_E_reg/P0001 ,
		_w4117_,
		_w36534_
	);
	LUT2 #(
		.INIT('h8)
	) name32488 (
		_w31266_,
		_w36507_,
		_w36535_
	);
	LUT2 #(
		.INIT('h1)
	) name32489 (
		_w36534_,
		_w36535_,
		_w36536_
	);
	LUT2 #(
		.INIT('h4)
	) name32490 (
		\core_c_dec_MFLreg_E_reg[7]/P0001 ,
		_w4117_,
		_w36537_
	);
	LUT2 #(
		.INIT('h1)
	) name32491 (
		_w34034_,
		_w36537_,
		_w36538_
	);
	LUT2 #(
		.INIT('h8)
	) name32492 (
		\core_c_dec_MFLreg_E_reg[6]/P0001 ,
		_w4117_,
		_w36539_
	);
	LUT2 #(
		.INIT('h8)
	) name32493 (
		_w34024_,
		_w36492_,
		_w36540_
	);
	LUT2 #(
		.INIT('h1)
	) name32494 (
		_w36539_,
		_w36540_,
		_w36541_
	);
	LUT2 #(
		.INIT('h1)
	) name32495 (
		_w4117_,
		_w34035_,
		_w36542_
	);
	LUT2 #(
		.INIT('h4)
	) name32496 (
		\core_c_dec_MFLreg_E_reg[5]/P0001 ,
		_w4117_,
		_w36543_
	);
	LUT2 #(
		.INIT('h1)
	) name32497 (
		_w36542_,
		_w36543_,
		_w36544_
	);
	LUT2 #(
		.INIT('h8)
	) name32498 (
		\core_c_dec_MFLreg_E_reg[4]/P0001 ,
		_w4117_,
		_w36545_
	);
	LUT2 #(
		.INIT('h8)
	) name32499 (
		_w25864_,
		_w34026_,
		_w36546_
	);
	LUT2 #(
		.INIT('h1)
	) name32500 (
		_w36545_,
		_w36546_,
		_w36547_
	);
	LUT2 #(
		.INIT('h4)
	) name32501 (
		_w4117_,
		_w31982_,
		_w36548_
	);
	LUT2 #(
		.INIT('h8)
	) name32502 (
		\core_c_dec_MFLreg_E_reg[3]/P0001 ,
		_w4117_,
		_w36549_
	);
	LUT2 #(
		.INIT('h1)
	) name32503 (
		_w36548_,
		_w36549_,
		_w36550_
	);
	LUT2 #(
		.INIT('h4)
	) name32504 (
		_w4117_,
		_w31975_,
		_w36551_
	);
	LUT2 #(
		.INIT('h8)
	) name32505 (
		\core_c_dec_MFLreg_E_reg[2]/P0001 ,
		_w4117_,
		_w36552_
	);
	LUT2 #(
		.INIT('h1)
	) name32506 (
		_w36551_,
		_w36552_,
		_w36553_
	);
	LUT2 #(
		.INIT('h4)
	) name32507 (
		\core_c_dec_MFLreg_E_reg[0]/P0001 ,
		_w4117_,
		_w36554_
	);
	LUT2 #(
		.INIT('h1)
	) name32508 (
		_w31971_,
		_w36554_,
		_w36555_
	);
	LUT2 #(
		.INIT('h8)
	) name32509 (
		\core_c_dec_MFIreg_E_reg[7]/P0001 ,
		_w4117_,
		_w36556_
	);
	LUT2 #(
		.INIT('h8)
	) name32510 (
		_w34028_,
		_w36507_,
		_w36557_
	);
	LUT2 #(
		.INIT('h1)
	) name32511 (
		_w36556_,
		_w36557_,
		_w36558_
	);
	LUT2 #(
		.INIT('h8)
	) name32512 (
		\core_c_dec_MFIreg_E_reg[6]/P0001 ,
		_w4117_,
		_w36559_
	);
	LUT2 #(
		.INIT('h8)
	) name32513 (
		_w34028_,
		_w35757_,
		_w36560_
	);
	LUT2 #(
		.INIT('h1)
	) name32514 (
		_w36559_,
		_w36560_,
		_w36561_
	);
	LUT2 #(
		.INIT('h8)
	) name32515 (
		\core_c_dec_MFIreg_E_reg[5]/P0001 ,
		_w4117_,
		_w36562_
	);
	LUT2 #(
		.INIT('h8)
	) name32516 (
		_w34025_,
		_w36507_,
		_w36563_
	);
	LUT2 #(
		.INIT('h1)
	) name32517 (
		_w36562_,
		_w36563_,
		_w36564_
	);
	LUT2 #(
		.INIT('h8)
	) name32518 (
		\core_c_dec_MFIreg_E_reg[4]/P0001 ,
		_w4117_,
		_w36565_
	);
	LUT2 #(
		.INIT('h8)
	) name32519 (
		_w34025_,
		_w35757_,
		_w36566_
	);
	LUT2 #(
		.INIT('h1)
	) name32520 (
		_w36565_,
		_w36566_,
		_w36567_
	);
	LUT2 #(
		.INIT('h8)
	) name32521 (
		\core_c_dec_MFIreg_E_reg[3]/P0001 ,
		_w4117_,
		_w36568_
	);
	LUT2 #(
		.INIT('h2)
	) name32522 (
		_w6093_,
		_w31263_,
		_w36569_
	);
	LUT2 #(
		.INIT('h8)
	) name32523 (
		_w36517_,
		_w36569_,
		_w36570_
	);
	LUT2 #(
		.INIT('h1)
	) name32524 (
		_w36568_,
		_w36570_,
		_w36571_
	);
	LUT2 #(
		.INIT('h8)
	) name32525 (
		\core_c_dec_MFIreg_E_reg[1]/P0001 ,
		_w4117_,
		_w36572_
	);
	LUT2 #(
		.INIT('h8)
	) name32526 (
		_w36527_,
		_w36569_,
		_w36573_
	);
	LUT2 #(
		.INIT('h1)
	) name32527 (
		_w36572_,
		_w36573_,
		_w36574_
	);
	LUT2 #(
		.INIT('h8)
	) name32528 (
		\core_c_dec_MFIreg_E_reg[0]/P0001 ,
		_w4117_,
		_w36575_
	);
	LUT2 #(
		.INIT('h8)
	) name32529 (
		_w31265_,
		_w31973_,
		_w36576_
	);
	LUT2 #(
		.INIT('h8)
	) name32530 (
		_w25729_,
		_w36576_,
		_w36577_
	);
	LUT2 #(
		.INIT('h1)
	) name32531 (
		_w36575_,
		_w36577_,
		_w36578_
	);
	LUT2 #(
		.INIT('h8)
	) name32532 (
		\core_c_dec_MFIMASK_E_reg/P0001 ,
		_w4117_,
		_w36579_
	);
	LUT2 #(
		.INIT('h8)
	) name32533 (
		_w31979_,
		_w36481_,
		_w36580_
	);
	LUT2 #(
		.INIT('h1)
	) name32534 (
		_w36579_,
		_w36580_,
		_w36581_
	);
	LUT2 #(
		.INIT('h4)
	) name32535 (
		_w4117_,
		_w33279_,
		_w36582_
	);
	LUT2 #(
		.INIT('h8)
	) name32536 (
		\core_c_dec_MFIDR_E_reg/P0001 ,
		_w4117_,
		_w36583_
	);
	LUT2 #(
		.INIT('h1)
	) name32537 (
		_w36582_,
		_w36583_,
		_w36584_
	);
	LUT2 #(
		.INIT('h4)
	) name32538 (
		\core_c_dec_MFDMOVL_E_reg/P0001 ,
		_w4117_,
		_w36585_
	);
	LUT2 #(
		.INIT('h1)
	) name32539 (
		_w33277_,
		_w36585_,
		_w36586_
	);
	LUT2 #(
		.INIT('h8)
	) name32540 (
		\core_c_dec_MFASTAT_E_reg/P0001 ,
		_w4117_,
		_w36587_
	);
	LUT2 #(
		.INIT('h8)
	) name32541 (
		_w31266_,
		_w35757_,
		_w36588_
	);
	LUT2 #(
		.INIT('h1)
	) name32542 (
		_w36587_,
		_w36588_,
		_w36589_
	);
	LUT2 #(
		.INIT('h1)
	) name32543 (
		\bdma_BEAD_reg[4]/NET0131 ,
		_w33305_,
		_w36590_
	);
	LUT2 #(
		.INIT('h1)
	) name32544 (
		_w20765_,
		_w33306_,
		_w36591_
	);
	LUT2 #(
		.INIT('h4)
	) name32545 (
		_w36590_,
		_w36591_,
		_w36592_
	);
	LUT2 #(
		.INIT('h8)
	) name32546 (
		_w10069_,
		_w20765_,
		_w36593_
	);
	LUT2 #(
		.INIT('h1)
	) name32547 (
		_w36592_,
		_w36593_,
		_w36594_
	);
	LUT2 #(
		.INIT('h1)
	) name32548 (
		\bdma_BEAD_reg[3]/NET0131 ,
		_w33304_,
		_w36595_
	);
	LUT2 #(
		.INIT('h1)
	) name32549 (
		_w20765_,
		_w33305_,
		_w36596_
	);
	LUT2 #(
		.INIT('h4)
	) name32550 (
		_w36595_,
		_w36596_,
		_w36597_
	);
	LUT2 #(
		.INIT('h8)
	) name32551 (
		_w8113_,
		_w20765_,
		_w36598_
	);
	LUT2 #(
		.INIT('h1)
	) name32552 (
		_w36597_,
		_w36598_,
		_w36599_
	);
	LUT2 #(
		.INIT('h8)
	) name32553 (
		\core_c_dec_MFIreg_E_reg[2]/P0001 ,
		_w4117_,
		_w36600_
	);
	LUT2 #(
		.INIT('h8)
	) name32554 (
		_w36522_,
		_w36569_,
		_w36601_
	);
	LUT2 #(
		.INIT('h1)
	) name32555 (
		_w36600_,
		_w36601_,
		_w36602_
	);
	LUT2 #(
		.INIT('h8)
	) name32556 (
		_w4215_,
		_w36427_,
		_w36603_
	);
	LUT2 #(
		.INIT('h2)
	) name32557 (
		_w4218_,
		_w36427_,
		_w36604_
	);
	LUT2 #(
		.INIT('h8)
	) name32558 (
		_w36441_,
		_w36604_,
		_w36605_
	);
	LUT2 #(
		.INIT('h1)
	) name32559 (
		\core_c_psq_pcstk_ptr_reg[4]/NET0131 ,
		_w36605_,
		_w36606_
	);
	LUT2 #(
		.INIT('h1)
	) name32560 (
		_w36603_,
		_w36606_,
		_w36607_
	);
	LUT2 #(
		.INIT('h1)
	) name32561 (
		\sice_ICYC_reg[19]/NET0131 ,
		_w20748_,
		_w36608_
	);
	LUT2 #(
		.INIT('h1)
	) name32562 (
		_w20749_,
		_w36608_,
		_w36609_
	);
	LUT2 #(
		.INIT('h8)
	) name32563 (
		\core_c_dec_MFtoppcs_Eg_reg/P0001 ,
		_w4118_,
		_w36610_
	);
	LUT2 #(
		.INIT('h8)
	) name32564 (
		_w23231_,
		_w32025_,
		_w36611_
	);
	LUT2 #(
		.INIT('h1)
	) name32565 (
		_w36610_,
		_w36611_,
		_w36612_
	);
	LUT2 #(
		.INIT('h8)
	) name32566 (
		\sice_SPC_reg[22]/P0001 ,
		_w34825_,
		_w36613_
	);
	LUT2 #(
		.INIT('h2)
	) name32567 (
		T_ID_pad,
		_w34825_,
		_w36614_
	);
	LUT2 #(
		.INIT('h1)
	) name32568 (
		_w36613_,
		_w36614_,
		_w36615_
	);
	LUT2 #(
		.INIT('h4)
	) name32569 (
		_w34827_,
		_w36615_,
		_w36616_
	);
	LUT2 #(
		.INIT('h8)
	) name32570 (
		\sice_IMR1_reg[17]/NET0131 ,
		_w34846_,
		_w36617_
	);
	LUT2 #(
		.INIT('h8)
	) name32571 (
		\sice_CMRW_reg/NET0131 ,
		_w23029_,
		_w36618_
	);
	LUT2 #(
		.INIT('h8)
	) name32572 (
		\sice_DMR1_reg[17]/NET0131 ,
		_w27903_,
		_w36619_
	);
	LUT2 #(
		.INIT('h8)
	) name32573 (
		\sice_DBR1_reg[18]/P0001 ,
		_w25054_,
		_w36620_
	);
	LUT2 #(
		.INIT('h8)
	) name32574 (
		\sice_DBR2_reg[18]/P0001 ,
		_w25012_,
		_w36621_
	);
	LUT2 #(
		.INIT('h8)
	) name32575 (
		\sice_IBR2_reg[17]/P0001 ,
		_w25074_,
		_w36622_
	);
	LUT2 #(
		.INIT('h8)
	) name32576 (
		\sice_idr1_reg_DO_reg[11]/P0001 ,
		_w26968_,
		_w36623_
	);
	LUT2 #(
		.INIT('h8)
	) name32577 (
		\emc_eRDY_reg/NET0131 ,
		_w35008_,
		_w36624_
	);
	LUT2 #(
		.INIT('h8)
	) name32578 (
		\core_c_dec_IR_reg[23]/NET0131 ,
		_w28203_,
		_w36625_
	);
	LUT2 #(
		.INIT('h8)
	) name32579 (
		\sice_IRR_reg[13]/P0001 ,
		_w34841_,
		_w36626_
	);
	LUT2 #(
		.INIT('h8)
	) name32580 (
		\sice_IIRC_reg[23]/NET0131 ,
		_w24267_,
		_w36627_
	);
	LUT2 #(
		.INIT('h8)
	) name32581 (
		\sice_IMR2_reg[17]/NET0131 ,
		_w25034_,
		_w36628_
	);
	LUT2 #(
		.INIT('h8)
	) name32582 (
		\sice_ICYC_reg[23]/NET0131 ,
		_w23409_,
		_w36629_
	);
	LUT2 #(
		.INIT('h8)
	) name32583 (
		\sice_IBR1_reg[17]/P0001 ,
		_w34831_,
		_w36630_
	);
	LUT2 #(
		.INIT('h8)
	) name32584 (
		\sice_DMR2_reg[17]/NET0131 ,
		_w25025_,
		_w36631_
	);
	LUT2 #(
		.INIT('h1)
	) name32585 (
		_w25084_,
		_w36617_,
		_w36632_
	);
	LUT2 #(
		.INIT('h1)
	) name32586 (
		_w36618_,
		_w36619_,
		_w36633_
	);
	LUT2 #(
		.INIT('h1)
	) name32587 (
		_w36620_,
		_w36621_,
		_w36634_
	);
	LUT2 #(
		.INIT('h1)
	) name32588 (
		_w36622_,
		_w36623_,
		_w36635_
	);
	LUT2 #(
		.INIT('h1)
	) name32589 (
		_w36625_,
		_w36626_,
		_w36636_
	);
	LUT2 #(
		.INIT('h1)
	) name32590 (
		_w36627_,
		_w36628_,
		_w36637_
	);
	LUT2 #(
		.INIT('h1)
	) name32591 (
		_w36629_,
		_w36630_,
		_w36638_
	);
	LUT2 #(
		.INIT('h4)
	) name32592 (
		_w36631_,
		_w36638_,
		_w36639_
	);
	LUT2 #(
		.INIT('h8)
	) name32593 (
		_w36636_,
		_w36637_,
		_w36640_
	);
	LUT2 #(
		.INIT('h8)
	) name32594 (
		_w36634_,
		_w36635_,
		_w36641_
	);
	LUT2 #(
		.INIT('h8)
	) name32595 (
		_w36632_,
		_w36633_,
		_w36642_
	);
	LUT2 #(
		.INIT('h4)
	) name32596 (
		_w36624_,
		_w36642_,
		_w36643_
	);
	LUT2 #(
		.INIT('h8)
	) name32597 (
		_w36640_,
		_w36641_,
		_w36644_
	);
	LUT2 #(
		.INIT('h8)
	) name32598 (
		_w36639_,
		_w36644_,
		_w36645_
	);
	LUT2 #(
		.INIT('h8)
	) name32599 (
		_w36643_,
		_w36645_,
		_w36646_
	);
	LUT2 #(
		.INIT('h8)
	) name32600 (
		_w34827_,
		_w36646_,
		_w36647_
	);
	LUT2 #(
		.INIT('h1)
	) name32601 (
		_w36616_,
		_w36647_,
		_w36648_
	);
	LUT2 #(
		.INIT('h8)
	) name32602 (
		\sice_SPC_reg[21]/P0001 ,
		_w34825_,
		_w36649_
	);
	LUT2 #(
		.INIT('h2)
	) name32603 (
		\sice_SPC_reg[23]/P0001 ,
		_w34825_,
		_w36650_
	);
	LUT2 #(
		.INIT('h1)
	) name32604 (
		_w36649_,
		_w36650_,
		_w36651_
	);
	LUT2 #(
		.INIT('h4)
	) name32605 (
		_w34827_,
		_w36651_,
		_w36652_
	);
	LUT2 #(
		.INIT('h8)
	) name32606 (
		\sice_IMR1_reg[16]/NET0131 ,
		_w34846_,
		_w36653_
	);
	LUT2 #(
		.INIT('h8)
	) name32607 (
		\sice_IIRC_reg[22]/NET0131 ,
		_w24267_,
		_w36654_
	);
	LUT2 #(
		.INIT('h8)
	) name32608 (
		\sice_DMR1_reg[16]/NET0131 ,
		_w27903_,
		_w36655_
	);
	LUT2 #(
		.INIT('h8)
	) name32609 (
		\sice_DBR1_reg[17]/P0001 ,
		_w25054_,
		_w36656_
	);
	LUT2 #(
		.INIT('h8)
	) name32610 (
		\sice_DBR2_reg[17]/P0001 ,
		_w25012_,
		_w36657_
	);
	LUT2 #(
		.INIT('h8)
	) name32611 (
		\sice_CLR_M_reg/NET0131 ,
		_w23029_,
		_w36658_
	);
	LUT2 #(
		.INIT('h8)
	) name32612 (
		\sice_idr1_reg_DO_reg[10]/P0001 ,
		_w26968_,
		_w36659_
	);
	LUT2 #(
		.INIT('h8)
	) name32613 (
		\sice_IDONE_reg/NET0131 ,
		_w35008_,
		_w36660_
	);
	LUT2 #(
		.INIT('h8)
	) name32614 (
		\core_c_dec_IR_reg[22]/NET0131 ,
		_w28203_,
		_w36661_
	);
	LUT2 #(
		.INIT('h8)
	) name32615 (
		\sice_IRR_reg[12]/P0001 ,
		_w34841_,
		_w36662_
	);
	LUT2 #(
		.INIT('h8)
	) name32616 (
		\sice_ICYC_reg[22]/NET0131 ,
		_w23409_,
		_w36663_
	);
	LUT2 #(
		.INIT('h8)
	) name32617 (
		\sice_IMR2_reg[16]/NET0131 ,
		_w25034_,
		_w36664_
	);
	LUT2 #(
		.INIT('h8)
	) name32618 (
		\sice_IBR2_reg[16]/P0001 ,
		_w25074_,
		_w36665_
	);
	LUT2 #(
		.INIT('h8)
	) name32619 (
		\sice_IBR1_reg[16]/P0001 ,
		_w34831_,
		_w36666_
	);
	LUT2 #(
		.INIT('h8)
	) name32620 (
		\sice_DMR2_reg[16]/NET0131 ,
		_w25025_,
		_w36667_
	);
	LUT2 #(
		.INIT('h1)
	) name32621 (
		_w25084_,
		_w36653_,
		_w36668_
	);
	LUT2 #(
		.INIT('h1)
	) name32622 (
		_w36654_,
		_w36655_,
		_w36669_
	);
	LUT2 #(
		.INIT('h1)
	) name32623 (
		_w36656_,
		_w36657_,
		_w36670_
	);
	LUT2 #(
		.INIT('h1)
	) name32624 (
		_w36658_,
		_w36659_,
		_w36671_
	);
	LUT2 #(
		.INIT('h1)
	) name32625 (
		_w36661_,
		_w36662_,
		_w36672_
	);
	LUT2 #(
		.INIT('h1)
	) name32626 (
		_w36663_,
		_w36664_,
		_w36673_
	);
	LUT2 #(
		.INIT('h1)
	) name32627 (
		_w36665_,
		_w36666_,
		_w36674_
	);
	LUT2 #(
		.INIT('h4)
	) name32628 (
		_w36667_,
		_w36674_,
		_w36675_
	);
	LUT2 #(
		.INIT('h8)
	) name32629 (
		_w36672_,
		_w36673_,
		_w36676_
	);
	LUT2 #(
		.INIT('h8)
	) name32630 (
		_w36670_,
		_w36671_,
		_w36677_
	);
	LUT2 #(
		.INIT('h8)
	) name32631 (
		_w36668_,
		_w36669_,
		_w36678_
	);
	LUT2 #(
		.INIT('h4)
	) name32632 (
		_w36660_,
		_w36678_,
		_w36679_
	);
	LUT2 #(
		.INIT('h8)
	) name32633 (
		_w36676_,
		_w36677_,
		_w36680_
	);
	LUT2 #(
		.INIT('h8)
	) name32634 (
		_w36675_,
		_w36680_,
		_w36681_
	);
	LUT2 #(
		.INIT('h8)
	) name32635 (
		_w36679_,
		_w36681_,
		_w36682_
	);
	LUT2 #(
		.INIT('h8)
	) name32636 (
		_w34827_,
		_w36682_,
		_w36683_
	);
	LUT2 #(
		.INIT('h1)
	) name32637 (
		_w36652_,
		_w36683_,
		_w36684_
	);
	LUT2 #(
		.INIT('h8)
	) name32638 (
		\sice_SPC_reg[19]/P0001 ,
		_w34825_,
		_w36685_
	);
	LUT2 #(
		.INIT('h2)
	) name32639 (
		\sice_SPC_reg[21]/P0001 ,
		_w34825_,
		_w36686_
	);
	LUT2 #(
		.INIT('h1)
	) name32640 (
		_w36685_,
		_w36686_,
		_w36687_
	);
	LUT2 #(
		.INIT('h4)
	) name32641 (
		_w34827_,
		_w36687_,
		_w36688_
	);
	LUT2 #(
		.INIT('h8)
	) name32642 (
		\sice_IMR1_reg[14]/NET0131 ,
		_w34846_,
		_w36689_
	);
	LUT2 #(
		.INIT('h8)
	) name32643 (
		\sice_IIRC_reg[20]/NET0131 ,
		_w24267_,
		_w36690_
	);
	LUT2 #(
		.INIT('h8)
	) name32644 (
		\sice_DMR1_reg[14]/NET0131 ,
		_w27903_,
		_w36691_
	);
	LUT2 #(
		.INIT('h8)
	) name32645 (
		\sice_DBR1_reg[15]/P0001 ,
		_w25054_,
		_w36692_
	);
	LUT2 #(
		.INIT('h8)
	) name32646 (
		\sice_DBR2_reg[15]/P0001 ,
		_w25012_,
		_w36693_
	);
	LUT2 #(
		.INIT('h8)
	) name32647 (
		\sice_GO_NX_reg/NET0131 ,
		_w23029_,
		_w36694_
	);
	LUT2 #(
		.INIT('h8)
	) name32648 (
		\sice_idr1_reg_DO_reg[8]/P0001 ,
		_w26968_,
		_w36695_
	);
	LUT2 #(
		.INIT('h4)
	) name32649 (
		_w4068_,
		_w35008_,
		_w36696_
	);
	LUT2 #(
		.INIT('h8)
	) name32650 (
		\core_c_dec_IR_reg[20]/NET0131 ,
		_w28203_,
		_w36697_
	);
	LUT2 #(
		.INIT('h8)
	) name32651 (
		\sice_IRR_reg[10]/P0001 ,
		_w34841_,
		_w36698_
	);
	LUT2 #(
		.INIT('h8)
	) name32652 (
		\sice_ICYC_reg[20]/NET0131 ,
		_w23409_,
		_w36699_
	);
	LUT2 #(
		.INIT('h8)
	) name32653 (
		\sice_IMR2_reg[14]/NET0131 ,
		_w25034_,
		_w36700_
	);
	LUT2 #(
		.INIT('h8)
	) name32654 (
		\sice_IBR2_reg[14]/P0001 ,
		_w25074_,
		_w36701_
	);
	LUT2 #(
		.INIT('h8)
	) name32655 (
		\sice_IBR1_reg[14]/P0001 ,
		_w34831_,
		_w36702_
	);
	LUT2 #(
		.INIT('h8)
	) name32656 (
		\sice_DMR2_reg[14]/NET0131 ,
		_w25025_,
		_w36703_
	);
	LUT2 #(
		.INIT('h1)
	) name32657 (
		_w25084_,
		_w36689_,
		_w36704_
	);
	LUT2 #(
		.INIT('h1)
	) name32658 (
		_w36690_,
		_w36691_,
		_w36705_
	);
	LUT2 #(
		.INIT('h1)
	) name32659 (
		_w36692_,
		_w36693_,
		_w36706_
	);
	LUT2 #(
		.INIT('h1)
	) name32660 (
		_w36694_,
		_w36695_,
		_w36707_
	);
	LUT2 #(
		.INIT('h1)
	) name32661 (
		_w36697_,
		_w36698_,
		_w36708_
	);
	LUT2 #(
		.INIT('h1)
	) name32662 (
		_w36699_,
		_w36700_,
		_w36709_
	);
	LUT2 #(
		.INIT('h1)
	) name32663 (
		_w36701_,
		_w36702_,
		_w36710_
	);
	LUT2 #(
		.INIT('h4)
	) name32664 (
		_w36703_,
		_w36710_,
		_w36711_
	);
	LUT2 #(
		.INIT('h8)
	) name32665 (
		_w36708_,
		_w36709_,
		_w36712_
	);
	LUT2 #(
		.INIT('h8)
	) name32666 (
		_w36706_,
		_w36707_,
		_w36713_
	);
	LUT2 #(
		.INIT('h8)
	) name32667 (
		_w36704_,
		_w36705_,
		_w36714_
	);
	LUT2 #(
		.INIT('h4)
	) name32668 (
		_w36696_,
		_w36714_,
		_w36715_
	);
	LUT2 #(
		.INIT('h8)
	) name32669 (
		_w36712_,
		_w36713_,
		_w36716_
	);
	LUT2 #(
		.INIT('h8)
	) name32670 (
		_w36711_,
		_w36716_,
		_w36717_
	);
	LUT2 #(
		.INIT('h8)
	) name32671 (
		_w36715_,
		_w36717_,
		_w36718_
	);
	LUT2 #(
		.INIT('h8)
	) name32672 (
		_w34827_,
		_w36718_,
		_w36719_
	);
	LUT2 #(
		.INIT('h1)
	) name32673 (
		_w36688_,
		_w36719_,
		_w36720_
	);
	LUT2 #(
		.INIT('h8)
	) name32674 (
		\sice_SPC_reg[18]/P0001 ,
		_w34825_,
		_w36721_
	);
	LUT2 #(
		.INIT('h2)
	) name32675 (
		\sice_SPC_reg[20]/P0001 ,
		_w34825_,
		_w36722_
	);
	LUT2 #(
		.INIT('h1)
	) name32676 (
		_w36721_,
		_w36722_,
		_w36723_
	);
	LUT2 #(
		.INIT('h4)
	) name32677 (
		_w34827_,
		_w36723_,
		_w36724_
	);
	LUT2 #(
		.INIT('h8)
	) name32678 (
		\sice_IMR1_reg[13]/NET0131 ,
		_w34846_,
		_w36725_
	);
	LUT2 #(
		.INIT('h8)
	) name32679 (
		\sice_IIRC_reg[19]/NET0131 ,
		_w24267_,
		_w36726_
	);
	LUT2 #(
		.INIT('h8)
	) name32680 (
		\sice_DMR1_reg[13]/NET0131 ,
		_w27903_,
		_w36727_
	);
	LUT2 #(
		.INIT('h8)
	) name32681 (
		\sice_DBR1_reg[14]/P0001 ,
		_w25054_,
		_w36728_
	);
	LUT2 #(
		.INIT('h8)
	) name32682 (
		\sice_DBR2_reg[14]/P0001 ,
		_w25012_,
		_w36729_
	);
	LUT2 #(
		.INIT('h4)
	) name32683 (
		_w23018_,
		_w23029_,
		_w36730_
	);
	LUT2 #(
		.INIT('h8)
	) name32684 (
		\sice_idr1_reg_DO_reg[7]/P0001 ,
		_w26968_,
		_w36731_
	);
	LUT2 #(
		.INIT('h8)
	) name32685 (
		\core_c_psq_MGNT_reg/NET0131 ,
		_w35008_,
		_w36732_
	);
	LUT2 #(
		.INIT('h8)
	) name32686 (
		\core_c_dec_IR_reg[19]/NET0131 ,
		_w28203_,
		_w36733_
	);
	LUT2 #(
		.INIT('h8)
	) name32687 (
		\sice_IRR_reg[9]/P0001 ,
		_w34841_,
		_w36734_
	);
	LUT2 #(
		.INIT('h8)
	) name32688 (
		\sice_ICYC_reg[19]/NET0131 ,
		_w23409_,
		_w36735_
	);
	LUT2 #(
		.INIT('h8)
	) name32689 (
		\sice_IMR2_reg[13]/NET0131 ,
		_w25034_,
		_w36736_
	);
	LUT2 #(
		.INIT('h8)
	) name32690 (
		\sice_IBR2_reg[13]/P0001 ,
		_w25074_,
		_w36737_
	);
	LUT2 #(
		.INIT('h8)
	) name32691 (
		\sice_IBR1_reg[13]/P0001 ,
		_w34831_,
		_w36738_
	);
	LUT2 #(
		.INIT('h8)
	) name32692 (
		\sice_DMR2_reg[13]/NET0131 ,
		_w25025_,
		_w36739_
	);
	LUT2 #(
		.INIT('h1)
	) name32693 (
		_w25084_,
		_w36725_,
		_w36740_
	);
	LUT2 #(
		.INIT('h1)
	) name32694 (
		_w36726_,
		_w36727_,
		_w36741_
	);
	LUT2 #(
		.INIT('h1)
	) name32695 (
		_w36728_,
		_w36729_,
		_w36742_
	);
	LUT2 #(
		.INIT('h1)
	) name32696 (
		_w36730_,
		_w36731_,
		_w36743_
	);
	LUT2 #(
		.INIT('h1)
	) name32697 (
		_w36733_,
		_w36734_,
		_w36744_
	);
	LUT2 #(
		.INIT('h1)
	) name32698 (
		_w36735_,
		_w36736_,
		_w36745_
	);
	LUT2 #(
		.INIT('h1)
	) name32699 (
		_w36737_,
		_w36738_,
		_w36746_
	);
	LUT2 #(
		.INIT('h4)
	) name32700 (
		_w36739_,
		_w36746_,
		_w36747_
	);
	LUT2 #(
		.INIT('h8)
	) name32701 (
		_w36744_,
		_w36745_,
		_w36748_
	);
	LUT2 #(
		.INIT('h8)
	) name32702 (
		_w36742_,
		_w36743_,
		_w36749_
	);
	LUT2 #(
		.INIT('h8)
	) name32703 (
		_w36740_,
		_w36741_,
		_w36750_
	);
	LUT2 #(
		.INIT('h4)
	) name32704 (
		_w36732_,
		_w36750_,
		_w36751_
	);
	LUT2 #(
		.INIT('h8)
	) name32705 (
		_w36748_,
		_w36749_,
		_w36752_
	);
	LUT2 #(
		.INIT('h8)
	) name32706 (
		_w36747_,
		_w36752_,
		_w36753_
	);
	LUT2 #(
		.INIT('h8)
	) name32707 (
		_w36751_,
		_w36753_,
		_w36754_
	);
	LUT2 #(
		.INIT('h8)
	) name32708 (
		_w34827_,
		_w36754_,
		_w36755_
	);
	LUT2 #(
		.INIT('h1)
	) name32709 (
		_w36724_,
		_w36755_,
		_w36756_
	);
	LUT2 #(
		.INIT('h8)
	) name32710 (
		\sice_SPC_reg[17]/P0001 ,
		_w34825_,
		_w36757_
	);
	LUT2 #(
		.INIT('h2)
	) name32711 (
		\sice_SPC_reg[19]/P0001 ,
		_w34825_,
		_w36758_
	);
	LUT2 #(
		.INIT('h1)
	) name32712 (
		_w36757_,
		_w36758_,
		_w36759_
	);
	LUT2 #(
		.INIT('h4)
	) name32713 (
		_w34827_,
		_w36759_,
		_w36760_
	);
	LUT2 #(
		.INIT('h8)
	) name32714 (
		\sice_IMR1_reg[12]/NET0131 ,
		_w34846_,
		_w36761_
	);
	LUT2 #(
		.INIT('h8)
	) name32715 (
		\sice_IIRC_reg[18]/NET0131 ,
		_w24267_,
		_w36762_
	);
	LUT2 #(
		.INIT('h8)
	) name32716 (
		\sice_DMR1_reg[12]/NET0131 ,
		_w27903_,
		_w36763_
	);
	LUT2 #(
		.INIT('h8)
	) name32717 (
		\sice_DBR1_reg[13]/P0001 ,
		_w25054_,
		_w36764_
	);
	LUT2 #(
		.INIT('h8)
	) name32718 (
		\sice_DBR2_reg[13]/P0001 ,
		_w25012_,
		_w36765_
	);
	LUT2 #(
		.INIT('h8)
	) name32719 (
		\sice_IRST_reg/NET0131 ,
		_w23029_,
		_w36766_
	);
	LUT2 #(
		.INIT('h8)
	) name32720 (
		\sice_idr1_reg_DO_reg[6]/P0001 ,
		_w26968_,
		_w36767_
	);
	LUT2 #(
		.INIT('h8)
	) name32721 (
		\core_c_psq_PCS_reg[3]/NET0131 ,
		_w35008_,
		_w36768_
	);
	LUT2 #(
		.INIT('h8)
	) name32722 (
		\core_c_dec_IR_reg[18]/NET0131 ,
		_w28203_,
		_w36769_
	);
	LUT2 #(
		.INIT('h8)
	) name32723 (
		\sice_IRR_reg[8]/P0001 ,
		_w34841_,
		_w36770_
	);
	LUT2 #(
		.INIT('h8)
	) name32724 (
		\sice_ICYC_reg[18]/NET0131 ,
		_w23409_,
		_w36771_
	);
	LUT2 #(
		.INIT('h8)
	) name32725 (
		\sice_IMR2_reg[12]/NET0131 ,
		_w25034_,
		_w36772_
	);
	LUT2 #(
		.INIT('h8)
	) name32726 (
		\sice_IBR2_reg[12]/P0001 ,
		_w25074_,
		_w36773_
	);
	LUT2 #(
		.INIT('h8)
	) name32727 (
		\sice_IBR1_reg[12]/P0001 ,
		_w34831_,
		_w36774_
	);
	LUT2 #(
		.INIT('h8)
	) name32728 (
		\sice_DMR2_reg[12]/NET0131 ,
		_w25025_,
		_w36775_
	);
	LUT2 #(
		.INIT('h1)
	) name32729 (
		_w25084_,
		_w36761_,
		_w36776_
	);
	LUT2 #(
		.INIT('h1)
	) name32730 (
		_w36762_,
		_w36763_,
		_w36777_
	);
	LUT2 #(
		.INIT('h1)
	) name32731 (
		_w36764_,
		_w36765_,
		_w36778_
	);
	LUT2 #(
		.INIT('h1)
	) name32732 (
		_w36766_,
		_w36767_,
		_w36779_
	);
	LUT2 #(
		.INIT('h1)
	) name32733 (
		_w36769_,
		_w36770_,
		_w36780_
	);
	LUT2 #(
		.INIT('h1)
	) name32734 (
		_w36771_,
		_w36772_,
		_w36781_
	);
	LUT2 #(
		.INIT('h1)
	) name32735 (
		_w36773_,
		_w36774_,
		_w36782_
	);
	LUT2 #(
		.INIT('h4)
	) name32736 (
		_w36775_,
		_w36782_,
		_w36783_
	);
	LUT2 #(
		.INIT('h8)
	) name32737 (
		_w36780_,
		_w36781_,
		_w36784_
	);
	LUT2 #(
		.INIT('h8)
	) name32738 (
		_w36778_,
		_w36779_,
		_w36785_
	);
	LUT2 #(
		.INIT('h8)
	) name32739 (
		_w36776_,
		_w36777_,
		_w36786_
	);
	LUT2 #(
		.INIT('h4)
	) name32740 (
		_w36768_,
		_w36786_,
		_w36787_
	);
	LUT2 #(
		.INIT('h8)
	) name32741 (
		_w36784_,
		_w36785_,
		_w36788_
	);
	LUT2 #(
		.INIT('h8)
	) name32742 (
		_w36783_,
		_w36788_,
		_w36789_
	);
	LUT2 #(
		.INIT('h8)
	) name32743 (
		_w36787_,
		_w36789_,
		_w36790_
	);
	LUT2 #(
		.INIT('h8)
	) name32744 (
		_w34827_,
		_w36790_,
		_w36791_
	);
	LUT2 #(
		.INIT('h1)
	) name32745 (
		_w36760_,
		_w36791_,
		_w36792_
	);
	LUT2 #(
		.INIT('h8)
	) name32746 (
		\core_c_dec_MFSB_E_reg/P0001 ,
		_w4117_,
		_w36793_
	);
	LUT2 #(
		.INIT('h8)
	) name32747 (
		_w31654_,
		_w35757_,
		_w36794_
	);
	LUT2 #(
		.INIT('h1)
	) name32748 (
		_w36793_,
		_w36794_,
		_w36795_
	);
	LUT2 #(
		.INIT('h4)
	) name32749 (
		_w4117_,
		_w31977_,
		_w36796_
	);
	LUT2 #(
		.INIT('h8)
	) name32750 (
		\core_c_dec_MFLreg_E_reg[1]/P0001 ,
		_w4117_,
		_w36797_
	);
	LUT2 #(
		.INIT('h1)
	) name32751 (
		_w36796_,
		_w36797_,
		_w36798_
	);
	LUT2 #(
		.INIT('h8)
	) name32752 (
		\core_c_dec_MFCNTR_E_reg/P0001 ,
		_w4117_,
		_w36799_
	);
	LUT2 #(
		.INIT('h8)
	) name32753 (
		_w35756_,
		_w36507_,
		_w36800_
	);
	LUT2 #(
		.INIT('h1)
	) name32754 (
		_w36799_,
		_w36800_,
		_w36801_
	);
	LUT2 #(
		.INIT('h8)
	) name32755 (
		\sice_SPC_reg[12]/P0001 ,
		_w34825_,
		_w36802_
	);
	LUT2 #(
		.INIT('h2)
	) name32756 (
		\sice_SPC_reg[14]/P0001 ,
		_w34825_,
		_w36803_
	);
	LUT2 #(
		.INIT('h1)
	) name32757 (
		_w36802_,
		_w36803_,
		_w36804_
	);
	LUT2 #(
		.INIT('h4)
	) name32758 (
		_w34827_,
		_w36804_,
		_w36805_
	);
	LUT2 #(
		.INIT('h8)
	) name32759 (
		\sice_IMR2_reg[7]/NET0131 ,
		_w25034_,
		_w36806_
	);
	LUT2 #(
		.INIT('h8)
	) name32760 (
		\sice_IRR_reg[3]/P0001 ,
		_w34841_,
		_w36807_
	);
	LUT2 #(
		.INIT('h8)
	) name32761 (
		\sice_IBR1_reg[7]/P0001 ,
		_w34831_,
		_w36808_
	);
	LUT2 #(
		.INIT('h8)
	) name32762 (
		\sice_IBR2_reg[7]/P0001 ,
		_w25074_,
		_w36809_
	);
	LUT2 #(
		.INIT('h8)
	) name32763 (
		\core_c_dec_IR_reg[13]/NET0131 ,
		_w28203_,
		_w36810_
	);
	LUT2 #(
		.INIT('h8)
	) name32764 (
		\sice_DMR2_reg[7]/NET0131 ,
		_w25025_,
		_w36811_
	);
	LUT2 #(
		.INIT('h8)
	) name32765 (
		\sice_ICYC_reg[13]/NET0131 ,
		_w23409_,
		_w36812_
	);
	LUT2 #(
		.INIT('h8)
	) name32766 (
		\sice_IMR1_reg[7]/NET0131 ,
		_w34846_,
		_w36813_
	);
	LUT2 #(
		.INIT('h8)
	) name32767 (
		\sice_DMR1_reg[7]/NET0131 ,
		_w27903_,
		_w36814_
	);
	LUT2 #(
		.INIT('h8)
	) name32768 (
		\sice_DBR2_reg[8]/P0001 ,
		_w25012_,
		_w36815_
	);
	LUT2 #(
		.INIT('h8)
	) name32769 (
		\sice_DBR1_reg[8]/P0001 ,
		_w25054_,
		_w36816_
	);
	LUT2 #(
		.INIT('h8)
	) name32770 (
		\sice_IIRC_reg[13]/NET0131 ,
		_w24267_,
		_w36817_
	);
	LUT2 #(
		.INIT('h8)
	) name32771 (
		\sice_idr1_reg_DO_reg[1]/P0001 ,
		_w26968_,
		_w36818_
	);
	LUT2 #(
		.INIT('h1)
	) name32772 (
		_w25083_,
		_w36806_,
		_w36819_
	);
	LUT2 #(
		.INIT('h1)
	) name32773 (
		_w36807_,
		_w36808_,
		_w36820_
	);
	LUT2 #(
		.INIT('h1)
	) name32774 (
		_w36809_,
		_w36810_,
		_w36821_
	);
	LUT2 #(
		.INIT('h1)
	) name32775 (
		_w36811_,
		_w36812_,
		_w36822_
	);
	LUT2 #(
		.INIT('h1)
	) name32776 (
		_w36813_,
		_w36814_,
		_w36823_
	);
	LUT2 #(
		.INIT('h1)
	) name32777 (
		_w36815_,
		_w36816_,
		_w36824_
	);
	LUT2 #(
		.INIT('h1)
	) name32778 (
		_w36817_,
		_w36818_,
		_w36825_
	);
	LUT2 #(
		.INIT('h8)
	) name32779 (
		_w36824_,
		_w36825_,
		_w36826_
	);
	LUT2 #(
		.INIT('h8)
	) name32780 (
		_w36822_,
		_w36823_,
		_w36827_
	);
	LUT2 #(
		.INIT('h8)
	) name32781 (
		_w36820_,
		_w36821_,
		_w36828_
	);
	LUT2 #(
		.INIT('h8)
	) name32782 (
		_w36819_,
		_w36828_,
		_w36829_
	);
	LUT2 #(
		.INIT('h8)
	) name32783 (
		_w36826_,
		_w36827_,
		_w36830_
	);
	LUT2 #(
		.INIT('h8)
	) name32784 (
		_w36829_,
		_w36830_,
		_w36831_
	);
	LUT2 #(
		.INIT('h8)
	) name32785 (
		_w34827_,
		_w36831_,
		_w36832_
	);
	LUT2 #(
		.INIT('h1)
	) name32786 (
		_w36805_,
		_w36832_,
		_w36833_
	);
	LUT2 #(
		.INIT('h8)
	) name32787 (
		\sice_SPC_reg[13]/P0001 ,
		_w34825_,
		_w36834_
	);
	LUT2 #(
		.INIT('h2)
	) name32788 (
		\sice_SPC_reg[15]/P0001 ,
		_w34825_,
		_w36835_
	);
	LUT2 #(
		.INIT('h1)
	) name32789 (
		_w36834_,
		_w36835_,
		_w36836_
	);
	LUT2 #(
		.INIT('h4)
	) name32790 (
		_w34827_,
		_w36836_,
		_w36837_
	);
	LUT2 #(
		.INIT('h8)
	) name32791 (
		\sice_DBR1_reg[9]/P0001 ,
		_w25054_,
		_w36838_
	);
	LUT2 #(
		.INIT('h8)
	) name32792 (
		\sice_IRR_reg[4]/P0001 ,
		_w34841_,
		_w36839_
	);
	LUT2 #(
		.INIT('h8)
	) name32793 (
		\sice_IMR2_reg[8]/NET0131 ,
		_w25034_,
		_w36840_
	);
	LUT2 #(
		.INIT('h8)
	) name32794 (
		\sice_IBR2_reg[8]/P0001 ,
		_w25074_,
		_w36841_
	);
	LUT2 #(
		.INIT('h8)
	) name32795 (
		\core_c_dec_IR_reg[14]/NET0131 ,
		_w28203_,
		_w36842_
	);
	LUT2 #(
		.INIT('h8)
	) name32796 (
		\sice_DMR2_reg[8]/NET0131 ,
		_w25025_,
		_w36843_
	);
	LUT2 #(
		.INIT('h8)
	) name32797 (
		\sice_ICYC_reg[14]/NET0131 ,
		_w23409_,
		_w36844_
	);
	LUT2 #(
		.INIT('h8)
	) name32798 (
		\sice_IMR1_reg[8]/NET0131 ,
		_w34846_,
		_w36845_
	);
	LUT2 #(
		.INIT('h8)
	) name32799 (
		\sice_IBR1_reg[8]/P0001 ,
		_w34831_,
		_w36846_
	);
	LUT2 #(
		.INIT('h8)
	) name32800 (
		\sice_IIRC_reg[14]/NET0131 ,
		_w24267_,
		_w36847_
	);
	LUT2 #(
		.INIT('h8)
	) name32801 (
		\sice_DBR2_reg[9]/P0001 ,
		_w25012_,
		_w36848_
	);
	LUT2 #(
		.INIT('h8)
	) name32802 (
		\sice_DMR1_reg[8]/NET0131 ,
		_w27903_,
		_w36849_
	);
	LUT2 #(
		.INIT('h8)
	) name32803 (
		\sice_idr1_reg_DO_reg[2]/P0001 ,
		_w26968_,
		_w36850_
	);
	LUT2 #(
		.INIT('h1)
	) name32804 (
		_w25083_,
		_w36838_,
		_w36851_
	);
	LUT2 #(
		.INIT('h1)
	) name32805 (
		_w36839_,
		_w36840_,
		_w36852_
	);
	LUT2 #(
		.INIT('h1)
	) name32806 (
		_w36841_,
		_w36842_,
		_w36853_
	);
	LUT2 #(
		.INIT('h1)
	) name32807 (
		_w36843_,
		_w36844_,
		_w36854_
	);
	LUT2 #(
		.INIT('h1)
	) name32808 (
		_w36845_,
		_w36846_,
		_w36855_
	);
	LUT2 #(
		.INIT('h1)
	) name32809 (
		_w36847_,
		_w36848_,
		_w36856_
	);
	LUT2 #(
		.INIT('h1)
	) name32810 (
		_w36849_,
		_w36850_,
		_w36857_
	);
	LUT2 #(
		.INIT('h8)
	) name32811 (
		_w36856_,
		_w36857_,
		_w36858_
	);
	LUT2 #(
		.INIT('h8)
	) name32812 (
		_w36854_,
		_w36855_,
		_w36859_
	);
	LUT2 #(
		.INIT('h8)
	) name32813 (
		_w36852_,
		_w36853_,
		_w36860_
	);
	LUT2 #(
		.INIT('h8)
	) name32814 (
		_w36851_,
		_w36860_,
		_w36861_
	);
	LUT2 #(
		.INIT('h8)
	) name32815 (
		_w36858_,
		_w36859_,
		_w36862_
	);
	LUT2 #(
		.INIT('h8)
	) name32816 (
		_w36861_,
		_w36862_,
		_w36863_
	);
	LUT2 #(
		.INIT('h8)
	) name32817 (
		_w34827_,
		_w36863_,
		_w36864_
	);
	LUT2 #(
		.INIT('h1)
	) name32818 (
		_w36837_,
		_w36864_,
		_w36865_
	);
	LUT2 #(
		.INIT('h8)
	) name32819 (
		\sice_SPC_reg[14]/P0001 ,
		_w34825_,
		_w36866_
	);
	LUT2 #(
		.INIT('h2)
	) name32820 (
		\sice_SPC_reg[16]/P0001 ,
		_w34825_,
		_w36867_
	);
	LUT2 #(
		.INIT('h1)
	) name32821 (
		_w36866_,
		_w36867_,
		_w36868_
	);
	LUT2 #(
		.INIT('h4)
	) name32822 (
		_w34827_,
		_w36868_,
		_w36869_
	);
	LUT2 #(
		.INIT('h8)
	) name32823 (
		\sice_DBR1_reg[10]/P0001 ,
		_w25054_,
		_w36870_
	);
	LUT2 #(
		.INIT('h8)
	) name32824 (
		\sice_IRR_reg[5]/P0001 ,
		_w34841_,
		_w36871_
	);
	LUT2 #(
		.INIT('h8)
	) name32825 (
		\sice_IMR2_reg[9]/NET0131 ,
		_w25034_,
		_w36872_
	);
	LUT2 #(
		.INIT('h8)
	) name32826 (
		\sice_IBR2_reg[9]/P0001 ,
		_w25074_,
		_w36873_
	);
	LUT2 #(
		.INIT('h8)
	) name32827 (
		\core_c_dec_IR_reg[15]/NET0131 ,
		_w28203_,
		_w36874_
	);
	LUT2 #(
		.INIT('h8)
	) name32828 (
		\sice_DMR2_reg[9]/NET0131 ,
		_w25025_,
		_w36875_
	);
	LUT2 #(
		.INIT('h8)
	) name32829 (
		\sice_ICYC_reg[15]/NET0131 ,
		_w23409_,
		_w36876_
	);
	LUT2 #(
		.INIT('h8)
	) name32830 (
		\sice_IMR1_reg[9]/NET0131 ,
		_w34846_,
		_w36877_
	);
	LUT2 #(
		.INIT('h8)
	) name32831 (
		\sice_IBR1_reg[9]/P0001 ,
		_w34831_,
		_w36878_
	);
	LUT2 #(
		.INIT('h8)
	) name32832 (
		\sice_IIRC_reg[15]/NET0131 ,
		_w24267_,
		_w36879_
	);
	LUT2 #(
		.INIT('h8)
	) name32833 (
		\sice_DBR2_reg[10]/P0001 ,
		_w25012_,
		_w36880_
	);
	LUT2 #(
		.INIT('h8)
	) name32834 (
		\sice_DMR1_reg[9]/NET0131 ,
		_w27903_,
		_w36881_
	);
	LUT2 #(
		.INIT('h8)
	) name32835 (
		\sice_idr1_reg_DO_reg[3]/P0001 ,
		_w26968_,
		_w36882_
	);
	LUT2 #(
		.INIT('h1)
	) name32836 (
		_w25083_,
		_w36870_,
		_w36883_
	);
	LUT2 #(
		.INIT('h1)
	) name32837 (
		_w36871_,
		_w36872_,
		_w36884_
	);
	LUT2 #(
		.INIT('h1)
	) name32838 (
		_w36873_,
		_w36874_,
		_w36885_
	);
	LUT2 #(
		.INIT('h1)
	) name32839 (
		_w36875_,
		_w36876_,
		_w36886_
	);
	LUT2 #(
		.INIT('h1)
	) name32840 (
		_w36877_,
		_w36878_,
		_w36887_
	);
	LUT2 #(
		.INIT('h1)
	) name32841 (
		_w36879_,
		_w36880_,
		_w36888_
	);
	LUT2 #(
		.INIT('h1)
	) name32842 (
		_w36881_,
		_w36882_,
		_w36889_
	);
	LUT2 #(
		.INIT('h8)
	) name32843 (
		_w36888_,
		_w36889_,
		_w36890_
	);
	LUT2 #(
		.INIT('h8)
	) name32844 (
		_w36886_,
		_w36887_,
		_w36891_
	);
	LUT2 #(
		.INIT('h8)
	) name32845 (
		_w36884_,
		_w36885_,
		_w36892_
	);
	LUT2 #(
		.INIT('h8)
	) name32846 (
		_w36883_,
		_w36892_,
		_w36893_
	);
	LUT2 #(
		.INIT('h8)
	) name32847 (
		_w36890_,
		_w36891_,
		_w36894_
	);
	LUT2 #(
		.INIT('h8)
	) name32848 (
		_w36893_,
		_w36894_,
		_w36895_
	);
	LUT2 #(
		.INIT('h8)
	) name32849 (
		_w34827_,
		_w36895_,
		_w36896_
	);
	LUT2 #(
		.INIT('h1)
	) name32850 (
		_w36869_,
		_w36896_,
		_w36897_
	);
	LUT2 #(
		.INIT('h1)
	) name32851 (
		\sice_ICYC_reg[11]/NET0131 ,
		_w20740_,
		_w36898_
	);
	LUT2 #(
		.INIT('h1)
	) name32852 (
		_w20741_,
		_w36898_,
		_w36899_
	);
	LUT2 #(
		.INIT('h1)
	) name32853 (
		\sice_IIRC_reg[11]/NET0131 ,
		_w20855_,
		_w36900_
	);
	LUT2 #(
		.INIT('h1)
	) name32854 (
		_w20856_,
		_w36900_,
		_w36901_
	);
	LUT2 #(
		.INIT('h8)
	) name32855 (
		\sice_SPC_reg[16]/P0001 ,
		_w34825_,
		_w36902_
	);
	LUT2 #(
		.INIT('h2)
	) name32856 (
		\sice_SPC_reg[18]/P0001 ,
		_w34825_,
		_w36903_
	);
	LUT2 #(
		.INIT('h1)
	) name32857 (
		_w36902_,
		_w36903_,
		_w36904_
	);
	LUT2 #(
		.INIT('h4)
	) name32858 (
		_w34827_,
		_w36904_,
		_w36905_
	);
	LUT2 #(
		.INIT('h8)
	) name32859 (
		\sice_DBR1_reg[12]/P0001 ,
		_w25054_,
		_w36906_
	);
	LUT2 #(
		.INIT('h8)
	) name32860 (
		\sice_IRR_reg[7]/P0001 ,
		_w34841_,
		_w36907_
	);
	LUT2 #(
		.INIT('h8)
	) name32861 (
		\sice_IMR2_reg[11]/NET0131 ,
		_w25034_,
		_w36908_
	);
	LUT2 #(
		.INIT('h8)
	) name32862 (
		\sice_IBR2_reg[11]/P0001 ,
		_w25074_,
		_w36909_
	);
	LUT2 #(
		.INIT('h8)
	) name32863 (
		\sice_idr1_reg_DO_reg[5]/P0001 ,
		_w26968_,
		_w36910_
	);
	LUT2 #(
		.INIT('h8)
	) name32864 (
		\sice_DMR2_reg[11]/NET0131 ,
		_w25025_,
		_w36911_
	);
	LUT2 #(
		.INIT('h8)
	) name32865 (
		\sice_ICYC_reg[17]/NET0131 ,
		_w23409_,
		_w36912_
	);
	LUT2 #(
		.INIT('h8)
	) name32866 (
		\sice_IMR1_reg[11]/NET0131 ,
		_w34846_,
		_w36913_
	);
	LUT2 #(
		.INIT('h8)
	) name32867 (
		\sice_IBR1_reg[11]/P0001 ,
		_w34831_,
		_w36914_
	);
	LUT2 #(
		.INIT('h8)
	) name32868 (
		\sice_IIRC_reg[17]/NET0131 ,
		_w24267_,
		_w36915_
	);
	LUT2 #(
		.INIT('h8)
	) name32869 (
		\sice_DBR2_reg[12]/P0001 ,
		_w25012_,
		_w36916_
	);
	LUT2 #(
		.INIT('h8)
	) name32870 (
		\sice_DMR1_reg[11]/NET0131 ,
		_w27903_,
		_w36917_
	);
	LUT2 #(
		.INIT('h8)
	) name32871 (
		\core_c_dec_IR_reg[17]/NET0131 ,
		_w28203_,
		_w36918_
	);
	LUT2 #(
		.INIT('h1)
	) name32872 (
		_w25083_,
		_w36906_,
		_w36919_
	);
	LUT2 #(
		.INIT('h1)
	) name32873 (
		_w36907_,
		_w36908_,
		_w36920_
	);
	LUT2 #(
		.INIT('h1)
	) name32874 (
		_w36909_,
		_w36910_,
		_w36921_
	);
	LUT2 #(
		.INIT('h1)
	) name32875 (
		_w36911_,
		_w36912_,
		_w36922_
	);
	LUT2 #(
		.INIT('h1)
	) name32876 (
		_w36913_,
		_w36914_,
		_w36923_
	);
	LUT2 #(
		.INIT('h1)
	) name32877 (
		_w36915_,
		_w36916_,
		_w36924_
	);
	LUT2 #(
		.INIT('h1)
	) name32878 (
		_w36917_,
		_w36918_,
		_w36925_
	);
	LUT2 #(
		.INIT('h8)
	) name32879 (
		_w36924_,
		_w36925_,
		_w36926_
	);
	LUT2 #(
		.INIT('h8)
	) name32880 (
		_w36922_,
		_w36923_,
		_w36927_
	);
	LUT2 #(
		.INIT('h8)
	) name32881 (
		_w36920_,
		_w36921_,
		_w36928_
	);
	LUT2 #(
		.INIT('h8)
	) name32882 (
		_w36919_,
		_w36928_,
		_w36929_
	);
	LUT2 #(
		.INIT('h8)
	) name32883 (
		_w36926_,
		_w36927_,
		_w36930_
	);
	LUT2 #(
		.INIT('h8)
	) name32884 (
		_w36929_,
		_w36930_,
		_w36931_
	);
	LUT2 #(
		.INIT('h8)
	) name32885 (
		_w34827_,
		_w36931_,
		_w36932_
	);
	LUT2 #(
		.INIT('h1)
	) name32886 (
		_w36905_,
		_w36932_,
		_w36933_
	);
	LUT2 #(
		.INIT('h1)
	) name32887 (
		\memc_Dread_E_reg/NET0131 ,
		\memc_Dwrite_E_reg/NET0131 ,
		_w36934_
	);
	LUT2 #(
		.INIT('h2)
	) name32888 (
		_w5435_,
		_w36934_,
		_w36935_
	);
	LUT2 #(
		.INIT('h4)
	) name32889 (
		_w4068_,
		_w36935_,
		_w36936_
	);
	LUT2 #(
		.INIT('h4)
	) name32890 (
		_w19054_,
		_w36936_,
		_w36937_
	);
	LUT2 #(
		.INIT('h2)
	) name32891 (
		\emc_DMcst_reg/NET0131 ,
		_w23398_,
		_w36938_
	);
	LUT2 #(
		.INIT('h8)
	) name32892 (
		_w19054_,
		_w36938_,
		_w36939_
	);
	LUT2 #(
		.INIT('h1)
	) name32893 (
		_w36937_,
		_w36939_,
		_w36940_
	);
	LUT2 #(
		.INIT('h8)
	) name32894 (
		\sice_SPC_reg[15]/P0001 ,
		_w34825_,
		_w36941_
	);
	LUT2 #(
		.INIT('h2)
	) name32895 (
		\sice_SPC_reg[17]/P0001 ,
		_w34825_,
		_w36942_
	);
	LUT2 #(
		.INIT('h1)
	) name32896 (
		_w36941_,
		_w36942_,
		_w36943_
	);
	LUT2 #(
		.INIT('h4)
	) name32897 (
		_w34827_,
		_w36943_,
		_w36944_
	);
	LUT2 #(
		.INIT('h8)
	) name32898 (
		\sice_DBR1_reg[11]/P0001 ,
		_w25054_,
		_w36945_
	);
	LUT2 #(
		.INIT('h8)
	) name32899 (
		\sice_IRR_reg[6]/P0001 ,
		_w34841_,
		_w36946_
	);
	LUT2 #(
		.INIT('h8)
	) name32900 (
		\sice_IMR2_reg[10]/NET0131 ,
		_w25034_,
		_w36947_
	);
	LUT2 #(
		.INIT('h8)
	) name32901 (
		\sice_IBR2_reg[10]/P0001 ,
		_w25074_,
		_w36948_
	);
	LUT2 #(
		.INIT('h8)
	) name32902 (
		\sice_idr1_reg_DO_reg[4]/P0001 ,
		_w26968_,
		_w36949_
	);
	LUT2 #(
		.INIT('h8)
	) name32903 (
		\sice_DMR2_reg[10]/NET0131 ,
		_w25025_,
		_w36950_
	);
	LUT2 #(
		.INIT('h8)
	) name32904 (
		\sice_ICYC_reg[16]/NET0131 ,
		_w23409_,
		_w36951_
	);
	LUT2 #(
		.INIT('h8)
	) name32905 (
		\sice_IMR1_reg[10]/NET0131 ,
		_w34846_,
		_w36952_
	);
	LUT2 #(
		.INIT('h8)
	) name32906 (
		\sice_IBR1_reg[10]/P0001 ,
		_w34831_,
		_w36953_
	);
	LUT2 #(
		.INIT('h8)
	) name32907 (
		\sice_IIRC_reg[16]/NET0131 ,
		_w24267_,
		_w36954_
	);
	LUT2 #(
		.INIT('h8)
	) name32908 (
		\sice_DBR2_reg[11]/P0001 ,
		_w25012_,
		_w36955_
	);
	LUT2 #(
		.INIT('h8)
	) name32909 (
		\sice_DMR1_reg[10]/NET0131 ,
		_w27903_,
		_w36956_
	);
	LUT2 #(
		.INIT('h8)
	) name32910 (
		\core_c_dec_IR_reg[16]/NET0131 ,
		_w28203_,
		_w36957_
	);
	LUT2 #(
		.INIT('h1)
	) name32911 (
		_w25083_,
		_w36945_,
		_w36958_
	);
	LUT2 #(
		.INIT('h1)
	) name32912 (
		_w36946_,
		_w36947_,
		_w36959_
	);
	LUT2 #(
		.INIT('h1)
	) name32913 (
		_w36948_,
		_w36949_,
		_w36960_
	);
	LUT2 #(
		.INIT('h1)
	) name32914 (
		_w36950_,
		_w36951_,
		_w36961_
	);
	LUT2 #(
		.INIT('h1)
	) name32915 (
		_w36952_,
		_w36953_,
		_w36962_
	);
	LUT2 #(
		.INIT('h1)
	) name32916 (
		_w36954_,
		_w36955_,
		_w36963_
	);
	LUT2 #(
		.INIT('h1)
	) name32917 (
		_w36956_,
		_w36957_,
		_w36964_
	);
	LUT2 #(
		.INIT('h8)
	) name32918 (
		_w36963_,
		_w36964_,
		_w36965_
	);
	LUT2 #(
		.INIT('h8)
	) name32919 (
		_w36961_,
		_w36962_,
		_w36966_
	);
	LUT2 #(
		.INIT('h8)
	) name32920 (
		_w36959_,
		_w36960_,
		_w36967_
	);
	LUT2 #(
		.INIT('h8)
	) name32921 (
		_w36958_,
		_w36967_,
		_w36968_
	);
	LUT2 #(
		.INIT('h8)
	) name32922 (
		_w36965_,
		_w36966_,
		_w36969_
	);
	LUT2 #(
		.INIT('h8)
	) name32923 (
		_w36968_,
		_w36969_,
		_w36970_
	);
	LUT2 #(
		.INIT('h8)
	) name32924 (
		_w34827_,
		_w36970_,
		_w36971_
	);
	LUT2 #(
		.INIT('h1)
	) name32925 (
		_w36944_,
		_w36971_,
		_w36972_
	);
	LUT2 #(
		.INIT('h2)
	) name32926 (
		\sice_SPC_reg[4]/P0001 ,
		_w26297_,
		_w36973_
	);
	LUT2 #(
		.INIT('h8)
	) name32927 (
		\sice_SPC_reg[3]/P0001 ,
		_w34825_,
		_w36974_
	);
	LUT2 #(
		.INIT('h2)
	) name32928 (
		\sice_SPC_reg[5]/P0001 ,
		_w34825_,
		_w36975_
	);
	LUT2 #(
		.INIT('h1)
	) name32929 (
		_w36974_,
		_w36975_,
		_w36976_
	);
	LUT2 #(
		.INIT('h4)
	) name32930 (
		_w34827_,
		_w36976_,
		_w36977_
	);
	LUT2 #(
		.INIT('h8)
	) name32931 (
		\sice_idr0_reg_DO_reg[4]/P0001 ,
		_w26968_,
		_w36978_
	);
	LUT2 #(
		.INIT('h8)
	) name32932 (
		\core_c_dec_IR_reg[4]/NET0131 ,
		_w28203_,
		_w36979_
	);
	LUT2 #(
		.INIT('h8)
	) name32933 (
		\sice_ICYC_reg[4]/NET0131 ,
		_w23409_,
		_w36980_
	);
	LUT2 #(
		.INIT('h8)
	) name32934 (
		\sice_IIRC_reg[4]/NET0131 ,
		_w24267_,
		_w36981_
	);
	LUT2 #(
		.INIT('h1)
	) name32935 (
		_w36978_,
		_w36979_,
		_w36982_
	);
	LUT2 #(
		.INIT('h1)
	) name32936 (
		_w36980_,
		_w36981_,
		_w36983_
	);
	LUT2 #(
		.INIT('h8)
	) name32937 (
		_w36982_,
		_w36983_,
		_w36984_
	);
	LUT2 #(
		.INIT('h8)
	) name32938 (
		_w34827_,
		_w36984_,
		_w36985_
	);
	LUT2 #(
		.INIT('h2)
	) name32939 (
		_w26297_,
		_w36977_,
		_w36986_
	);
	LUT2 #(
		.INIT('h4)
	) name32940 (
		_w36985_,
		_w36986_,
		_w36987_
	);
	LUT2 #(
		.INIT('h1)
	) name32941 (
		_w36973_,
		_w36987_,
		_w36988_
	);
	LUT2 #(
		.INIT('h2)
	) name32942 (
		\sice_SPC_reg[3]/P0001 ,
		_w26297_,
		_w36989_
	);
	LUT2 #(
		.INIT('h8)
	) name32943 (
		\sice_SPC_reg[2]/P0001 ,
		_w34825_,
		_w36990_
	);
	LUT2 #(
		.INIT('h2)
	) name32944 (
		\sice_SPC_reg[4]/P0001 ,
		_w34825_,
		_w36991_
	);
	LUT2 #(
		.INIT('h1)
	) name32945 (
		_w36990_,
		_w36991_,
		_w36992_
	);
	LUT2 #(
		.INIT('h4)
	) name32946 (
		_w34827_,
		_w36992_,
		_w36993_
	);
	LUT2 #(
		.INIT('h8)
	) name32947 (
		\sice_idr0_reg_DO_reg[3]/P0001 ,
		_w26968_,
		_w36994_
	);
	LUT2 #(
		.INIT('h8)
	) name32948 (
		\core_c_dec_IR_reg[3]/NET0131 ,
		_w28203_,
		_w36995_
	);
	LUT2 #(
		.INIT('h8)
	) name32949 (
		\sice_ICYC_reg[3]/NET0131 ,
		_w23409_,
		_w36996_
	);
	LUT2 #(
		.INIT('h8)
	) name32950 (
		\sice_IIRC_reg[3]/NET0131 ,
		_w24267_,
		_w36997_
	);
	LUT2 #(
		.INIT('h1)
	) name32951 (
		_w36994_,
		_w36995_,
		_w36998_
	);
	LUT2 #(
		.INIT('h1)
	) name32952 (
		_w36996_,
		_w36997_,
		_w36999_
	);
	LUT2 #(
		.INIT('h8)
	) name32953 (
		_w36998_,
		_w36999_,
		_w37000_
	);
	LUT2 #(
		.INIT('h8)
	) name32954 (
		_w34827_,
		_w37000_,
		_w37001_
	);
	LUT2 #(
		.INIT('h2)
	) name32955 (
		_w26297_,
		_w36993_,
		_w37002_
	);
	LUT2 #(
		.INIT('h4)
	) name32956 (
		_w37001_,
		_w37002_,
		_w37003_
	);
	LUT2 #(
		.INIT('h1)
	) name32957 (
		_w36989_,
		_w37003_,
		_w37004_
	);
	LUT2 #(
		.INIT('h2)
	) name32958 (
		\sice_SPC_reg[2]/P0001 ,
		_w26297_,
		_w37005_
	);
	LUT2 #(
		.INIT('h8)
	) name32959 (
		\sice_SPC_reg[1]/P0001 ,
		_w34825_,
		_w37006_
	);
	LUT2 #(
		.INIT('h2)
	) name32960 (
		\sice_SPC_reg[3]/P0001 ,
		_w34825_,
		_w37007_
	);
	LUT2 #(
		.INIT('h1)
	) name32961 (
		_w37006_,
		_w37007_,
		_w37008_
	);
	LUT2 #(
		.INIT('h4)
	) name32962 (
		_w34827_,
		_w37008_,
		_w37009_
	);
	LUT2 #(
		.INIT('h8)
	) name32963 (
		\sice_idr0_reg_DO_reg[2]/P0001 ,
		_w26968_,
		_w37010_
	);
	LUT2 #(
		.INIT('h8)
	) name32964 (
		\core_c_dec_IR_reg[2]/NET0131 ,
		_w28203_,
		_w37011_
	);
	LUT2 #(
		.INIT('h8)
	) name32965 (
		\sice_ICYC_reg[2]/NET0131 ,
		_w23409_,
		_w37012_
	);
	LUT2 #(
		.INIT('h8)
	) name32966 (
		\sice_IIRC_reg[2]/NET0131 ,
		_w24267_,
		_w37013_
	);
	LUT2 #(
		.INIT('h1)
	) name32967 (
		_w37010_,
		_w37011_,
		_w37014_
	);
	LUT2 #(
		.INIT('h1)
	) name32968 (
		_w37012_,
		_w37013_,
		_w37015_
	);
	LUT2 #(
		.INIT('h8)
	) name32969 (
		_w37014_,
		_w37015_,
		_w37016_
	);
	LUT2 #(
		.INIT('h8)
	) name32970 (
		_w34827_,
		_w37016_,
		_w37017_
	);
	LUT2 #(
		.INIT('h2)
	) name32971 (
		_w26297_,
		_w37009_,
		_w37018_
	);
	LUT2 #(
		.INIT('h4)
	) name32972 (
		_w37017_,
		_w37018_,
		_w37019_
	);
	LUT2 #(
		.INIT('h1)
	) name32973 (
		_w37005_,
		_w37019_,
		_w37020_
	);
	LUT2 #(
		.INIT('h2)
	) name32974 (
		\sice_SPC_reg[1]/P0001 ,
		_w26297_,
		_w37021_
	);
	LUT2 #(
		.INIT('h8)
	) name32975 (
		\sice_SPC_reg[0]/P0001 ,
		_w34825_,
		_w37022_
	);
	LUT2 #(
		.INIT('h2)
	) name32976 (
		\sice_SPC_reg[2]/P0001 ,
		_w34825_,
		_w37023_
	);
	LUT2 #(
		.INIT('h1)
	) name32977 (
		_w37022_,
		_w37023_,
		_w37024_
	);
	LUT2 #(
		.INIT('h4)
	) name32978 (
		_w34827_,
		_w37024_,
		_w37025_
	);
	LUT2 #(
		.INIT('h8)
	) name32979 (
		\sice_idr0_reg_DO_reg[1]/P0001 ,
		_w26968_,
		_w37026_
	);
	LUT2 #(
		.INIT('h8)
	) name32980 (
		\core_c_dec_IR_reg[1]/NET0131 ,
		_w28203_,
		_w37027_
	);
	LUT2 #(
		.INIT('h8)
	) name32981 (
		\sice_ICYC_reg[1]/NET0131 ,
		_w23409_,
		_w37028_
	);
	LUT2 #(
		.INIT('h8)
	) name32982 (
		\sice_IIRC_reg[1]/NET0131 ,
		_w24267_,
		_w37029_
	);
	LUT2 #(
		.INIT('h1)
	) name32983 (
		_w37026_,
		_w37027_,
		_w37030_
	);
	LUT2 #(
		.INIT('h1)
	) name32984 (
		_w37028_,
		_w37029_,
		_w37031_
	);
	LUT2 #(
		.INIT('h8)
	) name32985 (
		_w37030_,
		_w37031_,
		_w37032_
	);
	LUT2 #(
		.INIT('h8)
	) name32986 (
		_w34827_,
		_w37032_,
		_w37033_
	);
	LUT2 #(
		.INIT('h2)
	) name32987 (
		_w26297_,
		_w37025_,
		_w37034_
	);
	LUT2 #(
		.INIT('h4)
	) name32988 (
		_w37033_,
		_w37034_,
		_w37035_
	);
	LUT2 #(
		.INIT('h1)
	) name32989 (
		_w37021_,
		_w37035_,
		_w37036_
	);
	LUT2 #(
		.INIT('h8)
	) name32990 (
		_w14752_,
		_w31574_,
		_w37037_
	);
	LUT2 #(
		.INIT('h1)
	) name32991 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 ,
		_w17799_,
		_w37038_
	);
	LUT2 #(
		.INIT('h4)
	) name32992 (
		_w17809_,
		_w21663_,
		_w37039_
	);
	LUT2 #(
		.INIT('h2)
	) name32993 (
		_w17811_,
		_w37039_,
		_w37040_
	);
	LUT2 #(
		.INIT('h1)
	) name32994 (
		_w37038_,
		_w37040_,
		_w37041_
	);
	LUT2 #(
		.INIT('h1)
	) name32995 (
		_w17823_,
		_w37041_,
		_w37042_
	);
	LUT2 #(
		.INIT('h1)
	) name32996 (
		\core_eu_em_mac_em_reg_mr2rwe_DO_reg[3]/P0001 ,
		_w17808_,
		_w37043_
	);
	LUT2 #(
		.INIT('h1)
	) name32997 (
		_w37042_,
		_w37043_,
		_w37044_
	);
	LUT2 #(
		.INIT('h2)
	) name32998 (
		_w17829_,
		_w37044_,
		_w37045_
	);
	LUT2 #(
		.INIT('h1)
	) name32999 (
		_w37037_,
		_w37045_,
		_w37046_
	);
	LUT2 #(
		.INIT('h1)
	) name33000 (
		\clkc_STDcnt_reg[0]/NET0131 ,
		_w31521_,
		_w37047_
	);
	LUT2 #(
		.INIT('h1)
	) name33001 (
		\clkc_STDcnt_reg[9]/NET0131 ,
		_w31529_,
		_w37048_
	);
	LUT2 #(
		.INIT('h1)
	) name33002 (
		_w31521_,
		_w31530_,
		_w37049_
	);
	LUT2 #(
		.INIT('h4)
	) name33003 (
		_w37048_,
		_w37049_,
		_w37050_
	);
	LUT2 #(
		.INIT('h4)
	) name33004 (
		\sport0_rxctl_RXSHT_reg[7]/P0001 ,
		_w20868_,
		_w37051_
	);
	LUT2 #(
		.INIT('h8)
	) name33005 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w20873_,
		_w37052_
	);
	LUT2 #(
		.INIT('h1)
	) name33006 (
		_w31031_,
		_w34353_,
		_w37053_
	);
	LUT2 #(
		.INIT('h1)
	) name33007 (
		_w34354_,
		_w37053_,
		_w37054_
	);
	LUT2 #(
		.INIT('h2)
	) name33008 (
		_w31044_,
		_w37054_,
		_w37055_
	);
	LUT2 #(
		.INIT('h4)
	) name33009 (
		_w31044_,
		_w37054_,
		_w37056_
	);
	LUT2 #(
		.INIT('h2)
	) name33010 (
		_w20875_,
		_w37055_,
		_w37057_
	);
	LUT2 #(
		.INIT('h4)
	) name33011 (
		_w37056_,
		_w37057_,
		_w37058_
	);
	LUT2 #(
		.INIT('h4)
	) name33012 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w11265_,
		_w37059_
	);
	LUT2 #(
		.INIT('h1)
	) name33013 (
		_w20868_,
		_w37052_,
		_w37060_
	);
	LUT2 #(
		.INIT('h4)
	) name33014 (
		_w37059_,
		_w37060_,
		_w37061_
	);
	LUT2 #(
		.INIT('h4)
	) name33015 (
		_w37058_,
		_w37061_,
		_w37062_
	);
	LUT2 #(
		.INIT('h1)
	) name33016 (
		_w20871_,
		_w37051_,
		_w37063_
	);
	LUT2 #(
		.INIT('h4)
	) name33017 (
		_w37062_,
		_w37063_,
		_w37064_
	);
	LUT2 #(
		.INIT('h8)
	) name33018 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w20871_,
		_w37065_
	);
	LUT2 #(
		.INIT('h1)
	) name33019 (
		_w37064_,
		_w37065_,
		_w37066_
	);
	LUT2 #(
		.INIT('h2)
	) name33020 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w20259_,
		_w37067_
	);
	LUT2 #(
		.INIT('h4)
	) name33021 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w29085_,
		_w37068_
	);
	LUT2 #(
		.INIT('h1)
	) name33022 (
		_w37067_,
		_w37068_,
		_w37069_
	);
	LUT2 #(
		.INIT('h2)
	) name33023 (
		_w18717_,
		_w37069_,
		_w37070_
	);
	LUT2 #(
		.INIT('h1)
	) name33024 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[5]/P0001 ,
		_w18717_,
		_w37071_
	);
	LUT2 #(
		.INIT('h1)
	) name33025 (
		_w37070_,
		_w37071_,
		_w37072_
	);
	LUT2 #(
		.INIT('h2)
	) name33026 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w19559_,
		_w37073_
	);
	LUT2 #(
		.INIT('h4)
	) name33027 (
		\core_c_dec_MTSR1_E_reg/P0001 ,
		_w30613_,
		_w37074_
	);
	LUT2 #(
		.INIT('h1)
	) name33028 (
		_w37073_,
		_w37074_,
		_w37075_
	);
	LUT2 #(
		.INIT('h2)
	) name33029 (
		_w18717_,
		_w37075_,
		_w37076_
	);
	LUT2 #(
		.INIT('h1)
	) name33030 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[0]/P0001 ,
		_w18717_,
		_w37077_
	);
	LUT2 #(
		.INIT('h1)
	) name33031 (
		_w37076_,
		_w37077_,
		_w37078_
	);
	LUT2 #(
		.INIT('h2)
	) name33032 (
		_w17833_,
		_w37075_,
		_w37079_
	);
	LUT2 #(
		.INIT('h1)
	) name33033 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[0]/P0001 ,
		_w17833_,
		_w37080_
	);
	LUT2 #(
		.INIT('h1)
	) name33034 (
		_w37079_,
		_w37080_,
		_w37081_
	);
	LUT2 #(
		.INIT('h2)
	) name33035 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w23920_,
		_w37082_
	);
	LUT2 #(
		.INIT('h4)
	) name33036 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w30089_,
		_w37083_
	);
	LUT2 #(
		.INIT('h1)
	) name33037 (
		_w37082_,
		_w37083_,
		_w37084_
	);
	LUT2 #(
		.INIT('h2)
	) name33038 (
		_w18886_,
		_w37084_,
		_w37085_
	);
	LUT2 #(
		.INIT('h1)
	) name33039 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[12]/P0001 ,
		_w18886_,
		_w37086_
	);
	LUT2 #(
		.INIT('h1)
	) name33040 (
		_w37085_,
		_w37086_,
		_w37087_
	);
	LUT2 #(
		.INIT('h2)
	) name33041 (
		_w19034_,
		_w37084_,
		_w37088_
	);
	LUT2 #(
		.INIT('h1)
	) name33042 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[12]/P0001 ,
		_w19034_,
		_w37089_
	);
	LUT2 #(
		.INIT('h1)
	) name33043 (
		_w37088_,
		_w37089_,
		_w37090_
	);
	LUT2 #(
		.INIT('h2)
	) name33044 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 ,
		_w18266_,
		_w37091_
	);
	LUT2 #(
		.INIT('h1)
	) name33045 (
		\core_eu_em_mac_em_reg_mr0swe_DO_reg[7]/P0001 ,
		_w18271_,
		_w37092_
	);
	LUT2 #(
		.INIT('h2)
	) name33046 (
		_w18271_,
		_w19972_,
		_w37093_
	);
	LUT2 #(
		.INIT('h2)
	) name33047 (
		_w18273_,
		_w37092_,
		_w37094_
	);
	LUT2 #(
		.INIT('h4)
	) name33048 (
		_w37093_,
		_w37094_,
		_w37095_
	);
	LUT2 #(
		.INIT('h1)
	) name33049 (
		_w18270_,
		_w37091_,
		_w37096_
	);
	LUT2 #(
		.INIT('h4)
	) name33050 (
		_w37095_,
		_w37096_,
		_w37097_
	);
	LUT2 #(
		.INIT('h1)
	) name33051 (
		_w18262_,
		_w37097_,
		_w37098_
	);
	LUT2 #(
		.INIT('h2)
	) name33052 (
		_w18262_,
		_w19623_,
		_w37099_
	);
	LUT2 #(
		.INIT('h1)
	) name33053 (
		_w37098_,
		_w37099_,
		_w37100_
	);
	LUT2 #(
		.INIT('h8)
	) name33054 (
		_w14752_,
		_w19623_,
		_w37101_
	);
	LUT2 #(
		.INIT('h8)
	) name33055 (
		_w18328_,
		_w19972_,
		_w37102_
	);
	LUT2 #(
		.INIT('h2)
	) name33056 (
		\core_eu_em_mac_em_reg_mr0rwe_DO_reg[7]/P0001 ,
		_w18330_,
		_w37103_
	);
	LUT2 #(
		.INIT('h2)
	) name33057 (
		_w18334_,
		_w37103_,
		_w37104_
	);
	LUT2 #(
		.INIT('h4)
	) name33058 (
		_w37102_,
		_w37104_,
		_w37105_
	);
	LUT2 #(
		.INIT('h1)
	) name33059 (
		_w37101_,
		_w37105_,
		_w37106_
	);
	LUT2 #(
		.INIT('h4)
	) name33060 (
		\sport0_rxctl_RXSHT_reg[9]/P0001 ,
		_w20868_,
		_w37107_
	);
	LUT2 #(
		.INIT('h8)
	) name33061 (
		\sport0_rxctl_RX_reg[9]/P0001 ,
		_w20873_,
		_w37108_
	);
	LUT2 #(
		.INIT('h1)
	) name33062 (
		_w34363_,
		_w34396_,
		_w37109_
	);
	LUT2 #(
		.INIT('h1)
	) name33063 (
		_w34397_,
		_w37109_,
		_w37110_
	);
	LUT2 #(
		.INIT('h2)
	) name33064 (
		_w34399_,
		_w37110_,
		_w37111_
	);
	LUT2 #(
		.INIT('h4)
	) name33065 (
		_w34399_,
		_w37110_,
		_w37112_
	);
	LUT2 #(
		.INIT('h2)
	) name33066 (
		_w20875_,
		_w37111_,
		_w37113_
	);
	LUT2 #(
		.INIT('h4)
	) name33067 (
		_w37112_,
		_w37113_,
		_w37114_
	);
	LUT2 #(
		.INIT('h4)
	) name33068 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w10289_,
		_w37115_
	);
	LUT2 #(
		.INIT('h1)
	) name33069 (
		_w20868_,
		_w37108_,
		_w37116_
	);
	LUT2 #(
		.INIT('h4)
	) name33070 (
		_w37115_,
		_w37116_,
		_w37117_
	);
	LUT2 #(
		.INIT('h4)
	) name33071 (
		_w37114_,
		_w37117_,
		_w37118_
	);
	LUT2 #(
		.INIT('h1)
	) name33072 (
		_w20871_,
		_w37107_,
		_w37119_
	);
	LUT2 #(
		.INIT('h4)
	) name33073 (
		_w37118_,
		_w37119_,
		_w37120_
	);
	LUT2 #(
		.INIT('h8)
	) name33074 (
		\sport0_rxctl_RX_reg[9]/P0001 ,
		_w20871_,
		_w37121_
	);
	LUT2 #(
		.INIT('h1)
	) name33075 (
		_w37120_,
		_w37121_,
		_w37122_
	);
	LUT2 #(
		.INIT('h2)
	) name33076 (
		_w17833_,
		_w37069_,
		_w37123_
	);
	LUT2 #(
		.INIT('h1)
	) name33077 (
		\core_eu_es_sht_es_reg_sr1rwe_DO_reg[5]/P0001 ,
		_w17833_,
		_w37124_
	);
	LUT2 #(
		.INIT('h1)
	) name33078 (
		_w37123_,
		_w37124_,
		_w37125_
	);
	LUT2 #(
		.INIT('h2)
	) name33079 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w19972_,
		_w37126_
	);
	LUT2 #(
		.INIT('h4)
	) name33080 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w30245_,
		_w37127_
	);
	LUT2 #(
		.INIT('h1)
	) name33081 (
		_w37126_,
		_w37127_,
		_w37128_
	);
	LUT2 #(
		.INIT('h2)
	) name33082 (
		_w18886_,
		_w37128_,
		_w37129_
	);
	LUT2 #(
		.INIT('h1)
	) name33083 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[7]/P0001 ,
		_w18886_,
		_w37130_
	);
	LUT2 #(
		.INIT('h1)
	) name33084 (
		_w37129_,
		_w37130_,
		_w37131_
	);
	LUT2 #(
		.INIT('h2)
	) name33085 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w23757_,
		_w37132_
	);
	LUT2 #(
		.INIT('h4)
	) name33086 (
		\core_c_dec_MTSR0_E_reg/P0001 ,
		_w29776_,
		_w37133_
	);
	LUT2 #(
		.INIT('h1)
	) name33087 (
		_w37132_,
		_w37133_,
		_w37134_
	);
	LUT2 #(
		.INIT('h2)
	) name33088 (
		_w18886_,
		_w37134_,
		_w37135_
	);
	LUT2 #(
		.INIT('h1)
	) name33089 (
		\core_eu_es_sht_es_reg_sr0swe_DO_reg[11]/P0001 ,
		_w18886_,
		_w37136_
	);
	LUT2 #(
		.INIT('h1)
	) name33090 (
		_w37135_,
		_w37136_,
		_w37137_
	);
	LUT2 #(
		.INIT('h2)
	) name33091 (
		_w19034_,
		_w37128_,
		_w37138_
	);
	LUT2 #(
		.INIT('h1)
	) name33092 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[7]/P0001 ,
		_w19034_,
		_w37139_
	);
	LUT2 #(
		.INIT('h1)
	) name33093 (
		_w37138_,
		_w37139_,
		_w37140_
	);
	LUT2 #(
		.INIT('h2)
	) name33094 (
		_w19034_,
		_w37134_,
		_w37141_
	);
	LUT2 #(
		.INIT('h1)
	) name33095 (
		\core_eu_es_sht_es_reg_sr0rwe_DO_reg[11]/P0001 ,
		_w19034_,
		_w37142_
	);
	LUT2 #(
		.INIT('h1)
	) name33096 (
		_w37141_,
		_w37142_,
		_w37143_
	);
	LUT2 #(
		.INIT('h1)
	) name33097 (
		\clkc_STDcnt_reg[5]/NET0131 ,
		_w31525_,
		_w37144_
	);
	LUT2 #(
		.INIT('h1)
	) name33098 (
		_w31521_,
		_w31526_,
		_w37145_
	);
	LUT2 #(
		.INIT('h4)
	) name33099 (
		_w37144_,
		_w37145_,
		_w37146_
	);
	LUT2 #(
		.INIT('h1)
	) name33100 (
		\clkc_STDcnt_reg[2]/NET0131 ,
		_w31522_,
		_w37147_
	);
	LUT2 #(
		.INIT('h1)
	) name33101 (
		_w31523_,
		_w37147_,
		_w37148_
	);
	LUT2 #(
		.INIT('h4)
	) name33102 (
		_w31521_,
		_w37148_,
		_w37149_
	);
	LUT2 #(
		.INIT('h1)
	) name33103 (
		_w25833_,
		_w25835_,
		_w37150_
	);
	LUT2 #(
		.INIT('h4)
	) name33104 (
		_w22424_,
		_w37150_,
		_w37151_
	);
	LUT2 #(
		.INIT('h2)
	) name33105 (
		_w22424_,
		_w37150_,
		_w37152_
	);
	LUT2 #(
		.INIT('h1)
	) name33106 (
		_w37151_,
		_w37152_,
		_w37153_
	);
	LUT2 #(
		.INIT('h2)
	) name33107 (
		_w22411_,
		_w37153_,
		_w37154_
	);
	LUT2 #(
		.INIT('h2)
	) name33108 (
		\tm_TCR_TMP_reg[11]/NET0131 ,
		_w22411_,
		_w37155_
	);
	LUT2 #(
		.INIT('h1)
	) name33109 (
		_w37154_,
		_w37155_,
		_w37156_
	);
	LUT2 #(
		.INIT('h1)
	) name33110 (
		_w22400_,
		_w37156_,
		_w37157_
	);
	LUT2 #(
		.INIT('h8)
	) name33111 (
		\tm_tpr_reg_DO_reg[11]/NET0131 ,
		_w22400_,
		_w37158_
	);
	LUT2 #(
		.INIT('h1)
	) name33112 (
		_w37157_,
		_w37158_,
		_w37159_
	);
	LUT2 #(
		.INIT('h1)
	) name33113 (
		_w20355_,
		_w37159_,
		_w37160_
	);
	LUT2 #(
		.INIT('h8)
	) name33114 (
		\tm_tcr_reg_DO_reg[11]/NET0131 ,
		_w20355_,
		_w37161_
	);
	LUT2 #(
		.INIT('h1)
	) name33115 (
		_w37160_,
		_w37161_,
		_w37162_
	);
	LUT2 #(
		.INIT('h8)
	) name33116 (
		\T_ED[1]_pad ,
		_w34066_,
		_w37163_
	);
	LUT2 #(
		.INIT('h8)
	) name33117 (
		\bdma_BCTL_reg[0]/NET0131 ,
		\bdma_BCTL_reg[1]/NET0131 ,
		_w37164_
	);
	LUT2 #(
		.INIT('h4)
	) name33118 (
		_w34061_,
		_w37164_,
		_w37165_
	);
	LUT2 #(
		.INIT('h1)
	) name33119 (
		_w34066_,
		_w37165_,
		_w37166_
	);
	LUT2 #(
		.INIT('h8)
	) name33120 (
		\bdma_BRdataBUF_reg[9]/P0001 ,
		_w37166_,
		_w37167_
	);
	LUT2 #(
		.INIT('h1)
	) name33121 (
		_w37163_,
		_w37167_,
		_w37168_
	);
	LUT2 #(
		.INIT('h8)
	) name33122 (
		\T_ED[0]_pad ,
		_w34066_,
		_w37169_
	);
	LUT2 #(
		.INIT('h8)
	) name33123 (
		\bdma_BRdataBUF_reg[8]/P0001 ,
		_w37166_,
		_w37170_
	);
	LUT2 #(
		.INIT('h1)
	) name33124 (
		_w37169_,
		_w37170_,
		_w37171_
	);
	LUT2 #(
		.INIT('h8)
	) name33125 (
		\T_ED[7]_pad ,
		_w34066_,
		_w37172_
	);
	LUT2 #(
		.INIT('h8)
	) name33126 (
		\bdma_BRdataBUF_reg[15]/P0001 ,
		_w37166_,
		_w37173_
	);
	LUT2 #(
		.INIT('h1)
	) name33127 (
		_w37172_,
		_w37173_,
		_w37174_
	);
	LUT2 #(
		.INIT('h8)
	) name33128 (
		\T_ED[6]_pad ,
		_w34066_,
		_w37175_
	);
	LUT2 #(
		.INIT('h8)
	) name33129 (
		\bdma_BRdataBUF_reg[14]/P0001 ,
		_w37166_,
		_w37176_
	);
	LUT2 #(
		.INIT('h1)
	) name33130 (
		_w37175_,
		_w37176_,
		_w37177_
	);
	LUT2 #(
		.INIT('h8)
	) name33131 (
		\T_ED[5]_pad ,
		_w34066_,
		_w37178_
	);
	LUT2 #(
		.INIT('h8)
	) name33132 (
		\bdma_BRdataBUF_reg[13]/P0001 ,
		_w37166_,
		_w37179_
	);
	LUT2 #(
		.INIT('h1)
	) name33133 (
		_w37178_,
		_w37179_,
		_w37180_
	);
	LUT2 #(
		.INIT('h8)
	) name33134 (
		\T_ED[4]_pad ,
		_w34066_,
		_w37181_
	);
	LUT2 #(
		.INIT('h8)
	) name33135 (
		\bdma_BRdataBUF_reg[12]/P0001 ,
		_w37166_,
		_w37182_
	);
	LUT2 #(
		.INIT('h1)
	) name33136 (
		_w37181_,
		_w37182_,
		_w37183_
	);
	LUT2 #(
		.INIT('h8)
	) name33137 (
		\T_ED[3]_pad ,
		_w34066_,
		_w37184_
	);
	LUT2 #(
		.INIT('h8)
	) name33138 (
		\bdma_BRdataBUF_reg[11]/P0001 ,
		_w37166_,
		_w37185_
	);
	LUT2 #(
		.INIT('h1)
	) name33139 (
		_w37184_,
		_w37185_,
		_w37186_
	);
	LUT2 #(
		.INIT('h8)
	) name33140 (
		\T_ED[2]_pad ,
		_w34066_,
		_w37187_
	);
	LUT2 #(
		.INIT('h8)
	) name33141 (
		\bdma_BRdataBUF_reg[10]/P0001 ,
		_w37166_,
		_w37188_
	);
	LUT2 #(
		.INIT('h1)
	) name33142 (
		_w37187_,
		_w37188_,
		_w37189_
	);
	LUT2 #(
		.INIT('h2)
	) name33143 (
		\sice_SPC_reg[0]/P0001 ,
		_w26297_,
		_w37190_
	);
	LUT2 #(
		.INIT('h8)
	) name33144 (
		\sice_idr0_reg_DO_reg[0]/P0001 ,
		_w26968_,
		_w37191_
	);
	LUT2 #(
		.INIT('h8)
	) name33145 (
		\sice_ICYC_reg[0]/NET0131 ,
		_w23409_,
		_w37192_
	);
	LUT2 #(
		.INIT('h8)
	) name33146 (
		\sice_IIRC_reg[0]/NET0131 ,
		_w24267_,
		_w37193_
	);
	LUT2 #(
		.INIT('h8)
	) name33147 (
		\core_c_dec_IR_reg[0]/NET0131 ,
		_w28203_,
		_w37194_
	);
	LUT2 #(
		.INIT('h1)
	) name33148 (
		_w37191_,
		_w37192_,
		_w37195_
	);
	LUT2 #(
		.INIT('h1)
	) name33149 (
		_w37193_,
		_w37194_,
		_w37196_
	);
	LUT2 #(
		.INIT('h8)
	) name33150 (
		_w37195_,
		_w37196_,
		_w37197_
	);
	LUT2 #(
		.INIT('h2)
	) name33151 (
		_w34827_,
		_w37197_,
		_w37198_
	);
	LUT2 #(
		.INIT('h2)
	) name33152 (
		\sice_SPC_reg[1]/P0001 ,
		_w28982_,
		_w37199_
	);
	LUT2 #(
		.INIT('h1)
	) name33153 (
		_w37198_,
		_w37199_,
		_w37200_
	);
	LUT2 #(
		.INIT('h2)
	) name33154 (
		_w26297_,
		_w37200_,
		_w37201_
	);
	LUT2 #(
		.INIT('h1)
	) name33155 (
		_w37190_,
		_w37201_,
		_w37202_
	);
	LUT2 #(
		.INIT('h1)
	) name33156 (
		\clkc_STDcnt_reg[0]/NET0131 ,
		\clkc_STDcnt_reg[1]/NET0131 ,
		_w37203_
	);
	LUT2 #(
		.INIT('h1)
	) name33157 (
		_w31522_,
		_w37203_,
		_w37204_
	);
	LUT2 #(
		.INIT('h4)
	) name33158 (
		_w31521_,
		_w37204_,
		_w37205_
	);
	LUT2 #(
		.INIT('h8)
	) name33159 (
		\sport0_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w28944_,
		_w37206_
	);
	LUT2 #(
		.INIT('h8)
	) name33160 (
		\sport1_regs_MWORDreg_DO_reg[9]/NET0131 ,
		_w28854_,
		_w37207_
	);
	LUT2 #(
		.INIT('h8)
	) name33161 (
		\core_c_dec_updMF_E_reg/P0001 ,
		_w4118_,
		_w37208_
	);
	LUT2 #(
		.INIT('h8)
	) name33162 (
		_w18848_,
		_w20378_,
		_w37209_
	);
	LUT2 #(
		.INIT('h1)
	) name33163 (
		_w37208_,
		_w37209_,
		_w37210_
	);
	LUT2 #(
		.INIT('h8)
	) name33164 (
		\core_c_psq_SSTAT_reg[0]/NET0131 ,
		_w21137_,
		_w37211_
	);
	LUT2 #(
		.INIT('h1)
	) name33165 (
		_w36434_,
		_w37211_,
		_w37212_
	);
	LUT2 #(
		.INIT('h4)
	) name33166 (
		_w4218_,
		_w36435_,
		_w37213_
	);
	LUT2 #(
		.INIT('h1)
	) name33167 (
		_w37212_,
		_w37213_,
		_w37214_
	);
	LUT2 #(
		.INIT('h1)
	) name33168 (
		_w36073_,
		_w36075_,
		_w37215_
	);
	LUT2 #(
		.INIT('h8)
	) name33169 (
		\sport1_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w37215_,
		_w37216_
	);
	LUT2 #(
		.INIT('h8)
	) name33170 (
		_w7270_,
		_w18235_,
		_w37217_
	);
	LUT2 #(
		.INIT('h2)
	) name33171 (
		_w36073_,
		_w37217_,
		_w37218_
	);
	LUT2 #(
		.INIT('h8)
	) name33172 (
		_w8113_,
		_w37218_,
		_w37219_
	);
	LUT2 #(
		.INIT('h1)
	) name33173 (
		_w37216_,
		_w37219_,
		_w37220_
	);
	LUT2 #(
		.INIT('h8)
	) name33174 (
		\sport1_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w37215_,
		_w37221_
	);
	LUT2 #(
		.INIT('h8)
	) name33175 (
		_w8715_,
		_w37218_,
		_w37222_
	);
	LUT2 #(
		.INIT('h1)
	) name33176 (
		_w37221_,
		_w37222_,
		_w37223_
	);
	LUT2 #(
		.INIT('h8)
	) name33177 (
		\sport0_regs_SCTLreg_DO_reg[3]/NET0131 ,
		_w18233_,
		_w37224_
	);
	LUT2 #(
		.INIT('h8)
	) name33178 (
		_w8113_,
		_w18237_,
		_w37225_
	);
	LUT2 #(
		.INIT('h1)
	) name33179 (
		_w37224_,
		_w37225_,
		_w37226_
	);
	LUT2 #(
		.INIT('h8)
	) name33180 (
		\sport0_regs_SCTLreg_DO_reg[2]/NET0131 ,
		_w18233_,
		_w37227_
	);
	LUT2 #(
		.INIT('h8)
	) name33181 (
		_w8715_,
		_w18237_,
		_w37228_
	);
	LUT2 #(
		.INIT('h1)
	) name33182 (
		_w37227_,
		_w37228_,
		_w37229_
	);
	LUT2 #(
		.INIT('h4)
	) name33183 (
		\idma_IAL_reg/P0001 ,
		_w12688_,
		_w37230_
	);
	LUT2 #(
		.INIT('h8)
	) name33184 (
		\idma_IADi_reg[14]/P0001 ,
		\idma_IAL_reg/P0001 ,
		_w37231_
	);
	LUT2 #(
		.INIT('h1)
	) name33185 (
		_w37230_,
		_w37231_,
		_w37232_
	);
	LUT2 #(
		.INIT('h2)
	) name33186 (
		_w32455_,
		_w37232_,
		_w37233_
	);
	LUT2 #(
		.INIT('h2)
	) name33187 (
		\idma_DCTL_reg[14]/NET0131 ,
		_w32455_,
		_w37234_
	);
	LUT2 #(
		.INIT('h1)
	) name33188 (
		_w37233_,
		_w37234_,
		_w37235_
	);
	LUT2 #(
		.INIT('h2)
	) name33189 (
		\core_c_psq_Iact_E_reg[6]/NET0131 ,
		_w19477_,
		_w37236_
	);
	LUT2 #(
		.INIT('h4)
	) name33190 (
		_w19488_,
		_w19493_,
		_w37237_
	);
	LUT2 #(
		.INIT('h8)
	) name33191 (
		_w19487_,
		_w37237_,
		_w37238_
	);
	LUT2 #(
		.INIT('h1)
	) name33192 (
		_w37236_,
		_w37238_,
		_w37239_
	);
	LUT2 #(
		.INIT('h8)
	) name33193 (
		\bdma_BEAD_reg[11]/NET0131 ,
		\bdma_BM_cyc_reg/P0001 ,
		_w37240_
	);
	LUT2 #(
		.INIT('h8)
	) name33194 (
		\core_dag_ilm1reg_DMA_pi_DO_reg[11]/NET0131 ,
		_w5602_,
		_w37241_
	);
	LUT2 #(
		.INIT('h8)
	) name33195 (
		\emc_ECMA_reg[11]/P0001 ,
		\emc_ECMcs_reg/NET0131 ,
		_w37242_
	);
	LUT2 #(
		.INIT('h2)
	) name33196 (
		\core_dag_ilm2reg_PMA_pi_DO_reg[11]/NET0131 ,
		_w5608_,
		_w37243_
	);
	LUT2 #(
		.INIT('h1)
	) name33197 (
		_w37241_,
		_w37242_,
		_w37244_
	);
	LUT2 #(
		.INIT('h4)
	) name33198 (
		_w37243_,
		_w37244_,
		_w37245_
	);
	LUT2 #(
		.INIT('h1)
	) name33199 (
		\bdma_BM_cyc_reg/P0001 ,
		_w37245_,
		_w37246_
	);
	LUT2 #(
		.INIT('h1)
	) name33200 (
		_w37240_,
		_w37246_,
		_w37247_
	);
	LUT2 #(
		.INIT('h2)
	) name33201 (
		_w36427_,
		_w36440_,
		_w37248_
	);
	LUT2 #(
		.INIT('h8)
	) name33202 (
		_w4190_,
		_w37248_,
		_w37249_
	);
	LUT2 #(
		.INIT('h2)
	) name33203 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][7]/P0001 ,
		_w37249_,
		_w37250_
	);
	LUT2 #(
		.INIT('h4)
	) name33204 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5355_,
		_w37251_
	);
	LUT2 #(
		.INIT('h8)
	) name33205 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w11265_,
		_w37252_
	);
	LUT2 #(
		.INIT('h1)
	) name33206 (
		_w37251_,
		_w37252_,
		_w37253_
	);
	LUT2 #(
		.INIT('h1)
	) name33207 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37253_,
		_w37254_
	);
	LUT2 #(
		.INIT('h8)
	) name33208 (
		\core_c_psq_EXA_reg[7]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37255_
	);
	LUT2 #(
		.INIT('h1)
	) name33209 (
		_w37254_,
		_w37255_,
		_w37256_
	);
	LUT2 #(
		.INIT('h2)
	) name33210 (
		_w37249_,
		_w37256_,
		_w37257_
	);
	LUT2 #(
		.INIT('h1)
	) name33211 (
		_w37250_,
		_w37257_,
		_w37258_
	);
	LUT2 #(
		.INIT('h2)
	) name33212 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][5]/P0001 ,
		_w37249_,
		_w37259_
	);
	LUT2 #(
		.INIT('h4)
	) name33213 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5304_,
		_w37260_
	);
	LUT2 #(
		.INIT('h8)
	) name33214 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w10911_,
		_w37261_
	);
	LUT2 #(
		.INIT('h1)
	) name33215 (
		_w37260_,
		_w37261_,
		_w37262_
	);
	LUT2 #(
		.INIT('h1)
	) name33216 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37262_,
		_w37263_
	);
	LUT2 #(
		.INIT('h8)
	) name33217 (
		\core_c_psq_EXA_reg[5]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37264_
	);
	LUT2 #(
		.INIT('h1)
	) name33218 (
		_w37263_,
		_w37264_,
		_w37265_
	);
	LUT2 #(
		.INIT('h2)
	) name33219 (
		_w37249_,
		_w37265_,
		_w37266_
	);
	LUT2 #(
		.INIT('h1)
	) name33220 (
		_w37259_,
		_w37266_,
		_w37267_
	);
	LUT2 #(
		.INIT('h2)
	) name33221 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][4]/P0001 ,
		_w37249_,
		_w37268_
	);
	LUT2 #(
		.INIT('h4)
	) name33222 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5270_,
		_w37269_
	);
	LUT2 #(
		.INIT('h8)
	) name33223 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w10069_,
		_w37270_
	);
	LUT2 #(
		.INIT('h1)
	) name33224 (
		_w37269_,
		_w37270_,
		_w37271_
	);
	LUT2 #(
		.INIT('h1)
	) name33225 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37271_,
		_w37272_
	);
	LUT2 #(
		.INIT('h8)
	) name33226 (
		\core_c_psq_EXA_reg[4]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37273_
	);
	LUT2 #(
		.INIT('h1)
	) name33227 (
		_w37272_,
		_w37273_,
		_w37274_
	);
	LUT2 #(
		.INIT('h2)
	) name33228 (
		_w37249_,
		_w37274_,
		_w37275_
	);
	LUT2 #(
		.INIT('h1)
	) name33229 (
		_w37268_,
		_w37275_,
		_w37276_
	);
	LUT2 #(
		.INIT('h2)
	) name33230 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][3]/P0001 ,
		_w37249_,
		_w37277_
	);
	LUT2 #(
		.INIT('h4)
	) name33231 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5233_,
		_w37278_
	);
	LUT2 #(
		.INIT('h8)
	) name33232 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w8113_,
		_w37279_
	);
	LUT2 #(
		.INIT('h1)
	) name33233 (
		_w37278_,
		_w37279_,
		_w37280_
	);
	LUT2 #(
		.INIT('h1)
	) name33234 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37280_,
		_w37281_
	);
	LUT2 #(
		.INIT('h8)
	) name33235 (
		\core_c_psq_EXA_reg[3]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37282_
	);
	LUT2 #(
		.INIT('h1)
	) name33236 (
		_w37281_,
		_w37282_,
		_w37283_
	);
	LUT2 #(
		.INIT('h2)
	) name33237 (
		_w37249_,
		_w37283_,
		_w37284_
	);
	LUT2 #(
		.INIT('h1)
	) name33238 (
		_w37277_,
		_w37284_,
		_w37285_
	);
	LUT2 #(
		.INIT('h2)
	) name33239 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][1]/P0001 ,
		_w37249_,
		_w37286_
	);
	LUT2 #(
		.INIT('h4)
	) name33240 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5158_,
		_w37287_
	);
	LUT2 #(
		.INIT('h8)
	) name33241 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w9435_,
		_w37288_
	);
	LUT2 #(
		.INIT('h1)
	) name33242 (
		_w37287_,
		_w37288_,
		_w37289_
	);
	LUT2 #(
		.INIT('h1)
	) name33243 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37289_,
		_w37290_
	);
	LUT2 #(
		.INIT('h8)
	) name33244 (
		\core_c_psq_EXA_reg[1]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37291_
	);
	LUT2 #(
		.INIT('h1)
	) name33245 (
		_w37290_,
		_w37291_,
		_w37292_
	);
	LUT2 #(
		.INIT('h2)
	) name33246 (
		_w37249_,
		_w37292_,
		_w37293_
	);
	LUT2 #(
		.INIT('h1)
	) name33247 (
		_w37286_,
		_w37293_,
		_w37294_
	);
	LUT2 #(
		.INIT('h2)
	) name33248 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][11]/P0001 ,
		_w37249_,
		_w37295_
	);
	LUT2 #(
		.INIT('h4)
	) name33249 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5131_,
		_w37296_
	);
	LUT2 #(
		.INIT('h8)
	) name33250 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w8460_,
		_w37297_
	);
	LUT2 #(
		.INIT('h1)
	) name33251 (
		_w37296_,
		_w37297_,
		_w37298_
	);
	LUT2 #(
		.INIT('h1)
	) name33252 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37298_,
		_w37299_
	);
	LUT2 #(
		.INIT('h8)
	) name33253 (
		\core_c_psq_EXA_reg[11]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37300_
	);
	LUT2 #(
		.INIT('h1)
	) name33254 (
		_w37299_,
		_w37300_,
		_w37301_
	);
	LUT2 #(
		.INIT('h2)
	) name33255 (
		_w37249_,
		_w37301_,
		_w37302_
	);
	LUT2 #(
		.INIT('h1)
	) name33256 (
		_w37295_,
		_w37302_,
		_w37303_
	);
	LUT2 #(
		.INIT('h2)
	) name33257 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][10]/P0001 ,
		_w37249_,
		_w37304_
	);
	LUT2 #(
		.INIT('h4)
	) name33258 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5093_,
		_w37305_
	);
	LUT2 #(
		.INIT('h8)
	) name33259 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7859_,
		_w37306_
	);
	LUT2 #(
		.INIT('h1)
	) name33260 (
		_w37305_,
		_w37306_,
		_w37307_
	);
	LUT2 #(
		.INIT('h1)
	) name33261 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37307_,
		_w37308_
	);
	LUT2 #(
		.INIT('h8)
	) name33262 (
		\core_c_psq_EXA_reg[10]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37309_
	);
	LUT2 #(
		.INIT('h1)
	) name33263 (
		_w37308_,
		_w37309_,
		_w37310_
	);
	LUT2 #(
		.INIT('h2)
	) name33264 (
		_w37249_,
		_w37310_,
		_w37311_
	);
	LUT2 #(
		.INIT('h1)
	) name33265 (
		_w37304_,
		_w37311_,
		_w37312_
	);
	LUT2 #(
		.INIT('h1)
	) name33266 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		\core_c_psq_EXA_reg[0]/P0001 ,
		_w37313_
	);
	LUT2 #(
		.INIT('h8)
	) name33267 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7607_,
		_w37314_
	);
	LUT2 #(
		.INIT('h1)
	) name33268 (
		_w37313_,
		_w37314_,
		_w37315_
	);
	LUT2 #(
		.INIT('h1)
	) name33269 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37315_,
		_w37316_
	);
	LUT2 #(
		.INIT('h8)
	) name33270 (
		\core_c_psq_EXA_reg[0]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37317_
	);
	LUT2 #(
		.INIT('h1)
	) name33271 (
		_w37316_,
		_w37317_,
		_w37318_
	);
	LUT2 #(
		.INIT('h2)
	) name33272 (
		_w37249_,
		_w37318_,
		_w37319_
	);
	LUT2 #(
		.INIT('h2)
	) name33273 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][0]/P0001 ,
		_w37249_,
		_w37320_
	);
	LUT2 #(
		.INIT('h1)
	) name33274 (
		_w37319_,
		_w37320_,
		_w37321_
	);
	LUT2 #(
		.INIT('h8)
	) name33275 (
		_w4218_,
		_w37248_,
		_w37322_
	);
	LUT2 #(
		.INIT('h2)
	) name33276 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][9]/P0001 ,
		_w37322_,
		_w37323_
	);
	LUT2 #(
		.INIT('h4)
	) name33277 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5409_,
		_w37324_
	);
	LUT2 #(
		.INIT('h8)
	) name33278 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w10289_,
		_w37325_
	);
	LUT2 #(
		.INIT('h1)
	) name33279 (
		_w37324_,
		_w37325_,
		_w37326_
	);
	LUT2 #(
		.INIT('h1)
	) name33280 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37326_,
		_w37327_
	);
	LUT2 #(
		.INIT('h8)
	) name33281 (
		\core_c_psq_EXA_reg[9]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37328_
	);
	LUT2 #(
		.INIT('h1)
	) name33282 (
		_w37327_,
		_w37328_,
		_w37329_
	);
	LUT2 #(
		.INIT('h2)
	) name33283 (
		_w37322_,
		_w37329_,
		_w37330_
	);
	LUT2 #(
		.INIT('h1)
	) name33284 (
		_w37323_,
		_w37330_,
		_w37331_
	);
	LUT2 #(
		.INIT('h2)
	) name33285 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][8]/P0001 ,
		_w37322_,
		_w37332_
	);
	LUT2 #(
		.INIT('h4)
	) name33286 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5382_,
		_w37333_
	);
	LUT2 #(
		.INIT('h8)
	) name33287 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w10638_,
		_w37334_
	);
	LUT2 #(
		.INIT('h1)
	) name33288 (
		_w37333_,
		_w37334_,
		_w37335_
	);
	LUT2 #(
		.INIT('h1)
	) name33289 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37335_,
		_w37336_
	);
	LUT2 #(
		.INIT('h8)
	) name33290 (
		\core_c_psq_EXA_reg[8]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37337_
	);
	LUT2 #(
		.INIT('h1)
	) name33291 (
		_w37336_,
		_w37337_,
		_w37338_
	);
	LUT2 #(
		.INIT('h2)
	) name33292 (
		_w37322_,
		_w37338_,
		_w37339_
	);
	LUT2 #(
		.INIT('h1)
	) name33293 (
		_w37332_,
		_w37339_,
		_w37340_
	);
	LUT2 #(
		.INIT('h2)
	) name33294 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][7]/P0001 ,
		_w37322_,
		_w37341_
	);
	LUT2 #(
		.INIT('h4)
	) name33295 (
		_w37256_,
		_w37322_,
		_w37342_
	);
	LUT2 #(
		.INIT('h1)
	) name33296 (
		_w37341_,
		_w37342_,
		_w37343_
	);
	LUT2 #(
		.INIT('h2)
	) name33297 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][6]/P0001 ,
		_w37322_,
		_w37344_
	);
	LUT2 #(
		.INIT('h4)
	) name33298 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5328_,
		_w37345_
	);
	LUT2 #(
		.INIT('h8)
	) name33299 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w11525_,
		_w37346_
	);
	LUT2 #(
		.INIT('h1)
	) name33300 (
		_w37345_,
		_w37346_,
		_w37347_
	);
	LUT2 #(
		.INIT('h1)
	) name33301 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37347_,
		_w37348_
	);
	LUT2 #(
		.INIT('h8)
	) name33302 (
		\core_c_psq_EXA_reg[6]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37349_
	);
	LUT2 #(
		.INIT('h1)
	) name33303 (
		_w37348_,
		_w37349_,
		_w37350_
	);
	LUT2 #(
		.INIT('h2)
	) name33304 (
		_w37322_,
		_w37350_,
		_w37351_
	);
	LUT2 #(
		.INIT('h1)
	) name33305 (
		_w37344_,
		_w37351_,
		_w37352_
	);
	LUT2 #(
		.INIT('h2)
	) name33306 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][3]/P0001 ,
		_w37322_,
		_w37353_
	);
	LUT2 #(
		.INIT('h4)
	) name33307 (
		_w37283_,
		_w37322_,
		_w37354_
	);
	LUT2 #(
		.INIT('h1)
	) name33308 (
		_w37353_,
		_w37354_,
		_w37355_
	);
	LUT2 #(
		.INIT('h2)
	) name33309 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][2]/P0001 ,
		_w37322_,
		_w37356_
	);
	LUT2 #(
		.INIT('h4)
	) name33310 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5195_,
		_w37357_
	);
	LUT2 #(
		.INIT('h8)
	) name33311 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w8715_,
		_w37358_
	);
	LUT2 #(
		.INIT('h1)
	) name33312 (
		_w37357_,
		_w37358_,
		_w37359_
	);
	LUT2 #(
		.INIT('h1)
	) name33313 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37359_,
		_w37360_
	);
	LUT2 #(
		.INIT('h8)
	) name33314 (
		\core_c_psq_EXA_reg[2]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37361_
	);
	LUT2 #(
		.INIT('h1)
	) name33315 (
		_w37360_,
		_w37361_,
		_w37362_
	);
	LUT2 #(
		.INIT('h2)
	) name33316 (
		_w37322_,
		_w37362_,
		_w37363_
	);
	LUT2 #(
		.INIT('h1)
	) name33317 (
		_w37356_,
		_w37363_,
		_w37364_
	);
	LUT2 #(
		.INIT('h2)
	) name33318 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][1]/P0001 ,
		_w37322_,
		_w37365_
	);
	LUT2 #(
		.INIT('h4)
	) name33319 (
		_w37292_,
		_w37322_,
		_w37366_
	);
	LUT2 #(
		.INIT('h1)
	) name33320 (
		_w37365_,
		_w37366_,
		_w37367_
	);
	LUT2 #(
		.INIT('h2)
	) name33321 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][13]/P0001 ,
		_w37322_,
		_w37368_
	);
	LUT2 #(
		.INIT('h4)
	) name33322 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5649_,
		_w37369_
	);
	LUT2 #(
		.INIT('h8)
	) name33323 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w7340_,
		_w37370_
	);
	LUT2 #(
		.INIT('h1)
	) name33324 (
		_w37369_,
		_w37370_,
		_w37371_
	);
	LUT2 #(
		.INIT('h1)
	) name33325 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37371_,
		_w37372_
	);
	LUT2 #(
		.INIT('h8)
	) name33326 (
		\core_c_psq_EXA_reg[13]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37373_
	);
	LUT2 #(
		.INIT('h1)
	) name33327 (
		_w37372_,
		_w37373_,
		_w37374_
	);
	LUT2 #(
		.INIT('h2)
	) name33328 (
		_w37322_,
		_w37374_,
		_w37375_
	);
	LUT2 #(
		.INIT('h1)
	) name33329 (
		_w37368_,
		_w37375_,
		_w37376_
	);
	LUT2 #(
		.INIT('h2)
	) name33330 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][12]/P0001 ,
		_w37322_,
		_w37377_
	);
	LUT2 #(
		.INIT('h4)
	) name33331 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w5624_,
		_w37378_
	);
	LUT2 #(
		.INIT('h8)
	) name33332 (
		\core_c_dec_MTtoppcs_Eg_reg/P0001 ,
		_w9178_,
		_w37379_
	);
	LUT2 #(
		.INIT('h1)
	) name33333 (
		_w37378_,
		_w37379_,
		_w37380_
	);
	LUT2 #(
		.INIT('h1)
	) name33334 (
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37380_,
		_w37381_
	);
	LUT2 #(
		.INIT('h8)
	) name33335 (
		\core_c_psq_EXA_reg[12]/P0001 ,
		\core_c_psq_TRAP_Eg_reg/NET0131 ,
		_w37382_
	);
	LUT2 #(
		.INIT('h1)
	) name33336 (
		_w37381_,
		_w37382_,
		_w37383_
	);
	LUT2 #(
		.INIT('h2)
	) name33337 (
		_w37322_,
		_w37383_,
		_w37384_
	);
	LUT2 #(
		.INIT('h1)
	) name33338 (
		_w37377_,
		_w37384_,
		_w37385_
	);
	LUT2 #(
		.INIT('h2)
	) name33339 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][11]/P0001 ,
		_w37322_,
		_w37386_
	);
	LUT2 #(
		.INIT('h4)
	) name33340 (
		_w37301_,
		_w37322_,
		_w37387_
	);
	LUT2 #(
		.INIT('h1)
	) name33341 (
		_w37386_,
		_w37387_,
		_w37388_
	);
	LUT2 #(
		.INIT('h2)
	) name33342 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][10]/P0001 ,
		_w37322_,
		_w37389_
	);
	LUT2 #(
		.INIT('h4)
	) name33343 (
		_w37310_,
		_w37322_,
		_w37390_
	);
	LUT2 #(
		.INIT('h1)
	) name33344 (
		_w37389_,
		_w37390_,
		_w37391_
	);
	LUT2 #(
		.INIT('h4)
	) name33345 (
		_w37318_,
		_w37322_,
		_w37392_
	);
	LUT2 #(
		.INIT('h2)
	) name33346 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][0]/P0001 ,
		_w37322_,
		_w37393_
	);
	LUT2 #(
		.INIT('h1)
	) name33347 (
		_w37392_,
		_w37393_,
		_w37394_
	);
	LUT2 #(
		.INIT('h8)
	) name33348 (
		_w4222_,
		_w37248_,
		_w37395_
	);
	LUT2 #(
		.INIT('h2)
	) name33349 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][9]/P0001 ,
		_w37395_,
		_w37396_
	);
	LUT2 #(
		.INIT('h4)
	) name33350 (
		_w37329_,
		_w37395_,
		_w37397_
	);
	LUT2 #(
		.INIT('h1)
	) name33351 (
		_w37396_,
		_w37397_,
		_w37398_
	);
	LUT2 #(
		.INIT('h2)
	) name33352 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][8]/P0001 ,
		_w37395_,
		_w37399_
	);
	LUT2 #(
		.INIT('h4)
	) name33353 (
		_w37338_,
		_w37395_,
		_w37400_
	);
	LUT2 #(
		.INIT('h1)
	) name33354 (
		_w37399_,
		_w37400_,
		_w37401_
	);
	LUT2 #(
		.INIT('h2)
	) name33355 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][7]/P0001 ,
		_w37395_,
		_w37402_
	);
	LUT2 #(
		.INIT('h4)
	) name33356 (
		_w37256_,
		_w37395_,
		_w37403_
	);
	LUT2 #(
		.INIT('h1)
	) name33357 (
		_w37402_,
		_w37403_,
		_w37404_
	);
	LUT2 #(
		.INIT('h2)
	) name33358 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][6]/P0001 ,
		_w37395_,
		_w37405_
	);
	LUT2 #(
		.INIT('h4)
	) name33359 (
		_w37350_,
		_w37395_,
		_w37406_
	);
	LUT2 #(
		.INIT('h1)
	) name33360 (
		_w37405_,
		_w37406_,
		_w37407_
	);
	LUT2 #(
		.INIT('h2)
	) name33361 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][5]/P0001 ,
		_w37395_,
		_w37408_
	);
	LUT2 #(
		.INIT('h4)
	) name33362 (
		_w37265_,
		_w37395_,
		_w37409_
	);
	LUT2 #(
		.INIT('h1)
	) name33363 (
		_w37408_,
		_w37409_,
		_w37410_
	);
	LUT2 #(
		.INIT('h2)
	) name33364 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][4]/P0001 ,
		_w37395_,
		_w37411_
	);
	LUT2 #(
		.INIT('h4)
	) name33365 (
		_w37274_,
		_w37395_,
		_w37412_
	);
	LUT2 #(
		.INIT('h1)
	) name33366 (
		_w37411_,
		_w37412_,
		_w37413_
	);
	LUT2 #(
		.INIT('h2)
	) name33367 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][3]/P0001 ,
		_w37395_,
		_w37414_
	);
	LUT2 #(
		.INIT('h4)
	) name33368 (
		_w37283_,
		_w37395_,
		_w37415_
	);
	LUT2 #(
		.INIT('h1)
	) name33369 (
		_w37414_,
		_w37415_,
		_w37416_
	);
	LUT2 #(
		.INIT('h2)
	) name33370 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][2]/P0001 ,
		_w37395_,
		_w37417_
	);
	LUT2 #(
		.INIT('h4)
	) name33371 (
		_w37362_,
		_w37395_,
		_w37418_
	);
	LUT2 #(
		.INIT('h1)
	) name33372 (
		_w37417_,
		_w37418_,
		_w37419_
	);
	LUT2 #(
		.INIT('h2)
	) name33373 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][1]/P0001 ,
		_w37395_,
		_w37420_
	);
	LUT2 #(
		.INIT('h4)
	) name33374 (
		_w37292_,
		_w37395_,
		_w37421_
	);
	LUT2 #(
		.INIT('h1)
	) name33375 (
		_w37420_,
		_w37421_,
		_w37422_
	);
	LUT2 #(
		.INIT('h2)
	) name33376 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][13]/P0001 ,
		_w37395_,
		_w37423_
	);
	LUT2 #(
		.INIT('h4)
	) name33377 (
		_w37374_,
		_w37395_,
		_w37424_
	);
	LUT2 #(
		.INIT('h1)
	) name33378 (
		_w37423_,
		_w37424_,
		_w37425_
	);
	LUT2 #(
		.INIT('h2)
	) name33379 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][12]/P0001 ,
		_w37395_,
		_w37426_
	);
	LUT2 #(
		.INIT('h4)
	) name33380 (
		_w37383_,
		_w37395_,
		_w37427_
	);
	LUT2 #(
		.INIT('h1)
	) name33381 (
		_w37426_,
		_w37427_,
		_w37428_
	);
	LUT2 #(
		.INIT('h2)
	) name33382 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][11]/P0001 ,
		_w37395_,
		_w37429_
	);
	LUT2 #(
		.INIT('h4)
	) name33383 (
		_w37301_,
		_w37395_,
		_w37430_
	);
	LUT2 #(
		.INIT('h1)
	) name33384 (
		_w37429_,
		_w37430_,
		_w37431_
	);
	LUT2 #(
		.INIT('h2)
	) name33385 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][10]/P0001 ,
		_w37395_,
		_w37432_
	);
	LUT2 #(
		.INIT('h4)
	) name33386 (
		_w37310_,
		_w37395_,
		_w37433_
	);
	LUT2 #(
		.INIT('h1)
	) name33387 (
		_w37432_,
		_w37433_,
		_w37434_
	);
	LUT2 #(
		.INIT('h4)
	) name33388 (
		_w37318_,
		_w37395_,
		_w37435_
	);
	LUT2 #(
		.INIT('h2)
	) name33389 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[15][0]/P0001 ,
		_w37395_,
		_w37436_
	);
	LUT2 #(
		.INIT('h1)
	) name33390 (
		_w37435_,
		_w37436_,
		_w37437_
	);
	LUT2 #(
		.INIT('h8)
	) name33391 (
		_w4224_,
		_w37248_,
		_w37438_
	);
	LUT2 #(
		.INIT('h2)
	) name33392 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][9]/P0001 ,
		_w37438_,
		_w37439_
	);
	LUT2 #(
		.INIT('h4)
	) name33393 (
		_w37329_,
		_w37438_,
		_w37440_
	);
	LUT2 #(
		.INIT('h1)
	) name33394 (
		_w37439_,
		_w37440_,
		_w37441_
	);
	LUT2 #(
		.INIT('h2)
	) name33395 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][8]/P0001 ,
		_w37438_,
		_w37442_
	);
	LUT2 #(
		.INIT('h4)
	) name33396 (
		_w37338_,
		_w37438_,
		_w37443_
	);
	LUT2 #(
		.INIT('h1)
	) name33397 (
		_w37442_,
		_w37443_,
		_w37444_
	);
	LUT2 #(
		.INIT('h2)
	) name33398 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][7]/P0001 ,
		_w37438_,
		_w37445_
	);
	LUT2 #(
		.INIT('h4)
	) name33399 (
		_w37256_,
		_w37438_,
		_w37446_
	);
	LUT2 #(
		.INIT('h1)
	) name33400 (
		_w37445_,
		_w37446_,
		_w37447_
	);
	LUT2 #(
		.INIT('h2)
	) name33401 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][6]/P0001 ,
		_w37438_,
		_w37448_
	);
	LUT2 #(
		.INIT('h4)
	) name33402 (
		_w37350_,
		_w37438_,
		_w37449_
	);
	LUT2 #(
		.INIT('h1)
	) name33403 (
		_w37448_,
		_w37449_,
		_w37450_
	);
	LUT2 #(
		.INIT('h2)
	) name33404 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][5]/P0001 ,
		_w37438_,
		_w37451_
	);
	LUT2 #(
		.INIT('h4)
	) name33405 (
		_w37265_,
		_w37438_,
		_w37452_
	);
	LUT2 #(
		.INIT('h1)
	) name33406 (
		_w37451_,
		_w37452_,
		_w37453_
	);
	LUT2 #(
		.INIT('h2)
	) name33407 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][4]/P0001 ,
		_w37438_,
		_w37454_
	);
	LUT2 #(
		.INIT('h4)
	) name33408 (
		_w37274_,
		_w37438_,
		_w37455_
	);
	LUT2 #(
		.INIT('h1)
	) name33409 (
		_w37454_,
		_w37455_,
		_w37456_
	);
	LUT2 #(
		.INIT('h2)
	) name33410 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][3]/P0001 ,
		_w37438_,
		_w37457_
	);
	LUT2 #(
		.INIT('h4)
	) name33411 (
		_w37283_,
		_w37438_,
		_w37458_
	);
	LUT2 #(
		.INIT('h1)
	) name33412 (
		_w37457_,
		_w37458_,
		_w37459_
	);
	LUT2 #(
		.INIT('h2)
	) name33413 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][2]/P0001 ,
		_w37438_,
		_w37460_
	);
	LUT2 #(
		.INIT('h4)
	) name33414 (
		_w37362_,
		_w37438_,
		_w37461_
	);
	LUT2 #(
		.INIT('h1)
	) name33415 (
		_w37460_,
		_w37461_,
		_w37462_
	);
	LUT2 #(
		.INIT('h2)
	) name33416 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][1]/P0001 ,
		_w37438_,
		_w37463_
	);
	LUT2 #(
		.INIT('h4)
	) name33417 (
		_w37292_,
		_w37438_,
		_w37464_
	);
	LUT2 #(
		.INIT('h1)
	) name33418 (
		_w37463_,
		_w37464_,
		_w37465_
	);
	LUT2 #(
		.INIT('h2)
	) name33419 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][13]/P0001 ,
		_w37438_,
		_w37466_
	);
	LUT2 #(
		.INIT('h4)
	) name33420 (
		_w37374_,
		_w37438_,
		_w37467_
	);
	LUT2 #(
		.INIT('h1)
	) name33421 (
		_w37466_,
		_w37467_,
		_w37468_
	);
	LUT2 #(
		.INIT('h2)
	) name33422 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][12]/P0001 ,
		_w37438_,
		_w37469_
	);
	LUT2 #(
		.INIT('h4)
	) name33423 (
		_w37383_,
		_w37438_,
		_w37470_
	);
	LUT2 #(
		.INIT('h1)
	) name33424 (
		_w37469_,
		_w37470_,
		_w37471_
	);
	LUT2 #(
		.INIT('h2)
	) name33425 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][11]/P0001 ,
		_w37438_,
		_w37472_
	);
	LUT2 #(
		.INIT('h4)
	) name33426 (
		_w37301_,
		_w37438_,
		_w37473_
	);
	LUT2 #(
		.INIT('h1)
	) name33427 (
		_w37472_,
		_w37473_,
		_w37474_
	);
	LUT2 #(
		.INIT('h2)
	) name33428 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][10]/P0001 ,
		_w37438_,
		_w37475_
	);
	LUT2 #(
		.INIT('h4)
	) name33429 (
		_w37310_,
		_w37438_,
		_w37476_
	);
	LUT2 #(
		.INIT('h1)
	) name33430 (
		_w37475_,
		_w37476_,
		_w37477_
	);
	LUT2 #(
		.INIT('h4)
	) name33431 (
		_w37318_,
		_w37438_,
		_w37478_
	);
	LUT2 #(
		.INIT('h2)
	) name33432 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[14][0]/P0001 ,
		_w37438_,
		_w37479_
	);
	LUT2 #(
		.INIT('h1)
	) name33433 (
		_w37478_,
		_w37479_,
		_w37480_
	);
	LUT2 #(
		.INIT('h8)
	) name33434 (
		_w4194_,
		_w37248_,
		_w37481_
	);
	LUT2 #(
		.INIT('h2)
	) name33435 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][9]/P0001 ,
		_w37481_,
		_w37482_
	);
	LUT2 #(
		.INIT('h4)
	) name33436 (
		_w37329_,
		_w37481_,
		_w37483_
	);
	LUT2 #(
		.INIT('h1)
	) name33437 (
		_w37482_,
		_w37483_,
		_w37484_
	);
	LUT2 #(
		.INIT('h2)
	) name33438 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][8]/P0001 ,
		_w37481_,
		_w37485_
	);
	LUT2 #(
		.INIT('h4)
	) name33439 (
		_w37338_,
		_w37481_,
		_w37486_
	);
	LUT2 #(
		.INIT('h1)
	) name33440 (
		_w37485_,
		_w37486_,
		_w37487_
	);
	LUT2 #(
		.INIT('h2)
	) name33441 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][7]/P0001 ,
		_w37481_,
		_w37488_
	);
	LUT2 #(
		.INIT('h4)
	) name33442 (
		_w37256_,
		_w37481_,
		_w37489_
	);
	LUT2 #(
		.INIT('h1)
	) name33443 (
		_w37488_,
		_w37489_,
		_w37490_
	);
	LUT2 #(
		.INIT('h2)
	) name33444 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][6]/P0001 ,
		_w37481_,
		_w37491_
	);
	LUT2 #(
		.INIT('h4)
	) name33445 (
		_w37350_,
		_w37481_,
		_w37492_
	);
	LUT2 #(
		.INIT('h1)
	) name33446 (
		_w37491_,
		_w37492_,
		_w37493_
	);
	LUT2 #(
		.INIT('h2)
	) name33447 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][5]/P0001 ,
		_w37481_,
		_w37494_
	);
	LUT2 #(
		.INIT('h4)
	) name33448 (
		_w37265_,
		_w37481_,
		_w37495_
	);
	LUT2 #(
		.INIT('h1)
	) name33449 (
		_w37494_,
		_w37495_,
		_w37496_
	);
	LUT2 #(
		.INIT('h2)
	) name33450 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][4]/P0001 ,
		_w37481_,
		_w37497_
	);
	LUT2 #(
		.INIT('h4)
	) name33451 (
		_w37274_,
		_w37481_,
		_w37498_
	);
	LUT2 #(
		.INIT('h1)
	) name33452 (
		_w37497_,
		_w37498_,
		_w37499_
	);
	LUT2 #(
		.INIT('h2)
	) name33453 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][3]/P0001 ,
		_w37481_,
		_w37500_
	);
	LUT2 #(
		.INIT('h4)
	) name33454 (
		_w37283_,
		_w37481_,
		_w37501_
	);
	LUT2 #(
		.INIT('h1)
	) name33455 (
		_w37500_,
		_w37501_,
		_w37502_
	);
	LUT2 #(
		.INIT('h2)
	) name33456 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][2]/P0001 ,
		_w37481_,
		_w37503_
	);
	LUT2 #(
		.INIT('h4)
	) name33457 (
		_w37362_,
		_w37481_,
		_w37504_
	);
	LUT2 #(
		.INIT('h1)
	) name33458 (
		_w37503_,
		_w37504_,
		_w37505_
	);
	LUT2 #(
		.INIT('h2)
	) name33459 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][1]/P0001 ,
		_w37481_,
		_w37506_
	);
	LUT2 #(
		.INIT('h4)
	) name33460 (
		_w37292_,
		_w37481_,
		_w37507_
	);
	LUT2 #(
		.INIT('h1)
	) name33461 (
		_w37506_,
		_w37507_,
		_w37508_
	);
	LUT2 #(
		.INIT('h2)
	) name33462 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][13]/P0001 ,
		_w37481_,
		_w37509_
	);
	LUT2 #(
		.INIT('h4)
	) name33463 (
		_w37374_,
		_w37481_,
		_w37510_
	);
	LUT2 #(
		.INIT('h1)
	) name33464 (
		_w37509_,
		_w37510_,
		_w37511_
	);
	LUT2 #(
		.INIT('h2)
	) name33465 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][12]/P0001 ,
		_w37481_,
		_w37512_
	);
	LUT2 #(
		.INIT('h4)
	) name33466 (
		_w37383_,
		_w37481_,
		_w37513_
	);
	LUT2 #(
		.INIT('h1)
	) name33467 (
		_w37512_,
		_w37513_,
		_w37514_
	);
	LUT2 #(
		.INIT('h2)
	) name33468 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][11]/P0001 ,
		_w37481_,
		_w37515_
	);
	LUT2 #(
		.INIT('h4)
	) name33469 (
		_w37301_,
		_w37481_,
		_w37516_
	);
	LUT2 #(
		.INIT('h1)
	) name33470 (
		_w37515_,
		_w37516_,
		_w37517_
	);
	LUT2 #(
		.INIT('h2)
	) name33471 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][10]/P0001 ,
		_w37481_,
		_w37518_
	);
	LUT2 #(
		.INIT('h4)
	) name33472 (
		_w37310_,
		_w37481_,
		_w37519_
	);
	LUT2 #(
		.INIT('h1)
	) name33473 (
		_w37518_,
		_w37519_,
		_w37520_
	);
	LUT2 #(
		.INIT('h4)
	) name33474 (
		_w37318_,
		_w37481_,
		_w37521_
	);
	LUT2 #(
		.INIT('h2)
	) name33475 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[13][0]/P0001 ,
		_w37481_,
		_w37522_
	);
	LUT2 #(
		.INIT('h1)
	) name33476 (
		_w37521_,
		_w37522_,
		_w37523_
	);
	LUT2 #(
		.INIT('h8)
	) name33477 (
		_w4205_,
		_w37248_,
		_w37524_
	);
	LUT2 #(
		.INIT('h2)
	) name33478 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][9]/P0001 ,
		_w37524_,
		_w37525_
	);
	LUT2 #(
		.INIT('h4)
	) name33479 (
		_w37329_,
		_w37524_,
		_w37526_
	);
	LUT2 #(
		.INIT('h1)
	) name33480 (
		_w37525_,
		_w37526_,
		_w37527_
	);
	LUT2 #(
		.INIT('h2)
	) name33481 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][8]/P0001 ,
		_w37524_,
		_w37528_
	);
	LUT2 #(
		.INIT('h4)
	) name33482 (
		_w37338_,
		_w37524_,
		_w37529_
	);
	LUT2 #(
		.INIT('h1)
	) name33483 (
		_w37528_,
		_w37529_,
		_w37530_
	);
	LUT2 #(
		.INIT('h2)
	) name33484 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][7]/P0001 ,
		_w37524_,
		_w37531_
	);
	LUT2 #(
		.INIT('h4)
	) name33485 (
		_w37256_,
		_w37524_,
		_w37532_
	);
	LUT2 #(
		.INIT('h1)
	) name33486 (
		_w37531_,
		_w37532_,
		_w37533_
	);
	LUT2 #(
		.INIT('h2)
	) name33487 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][6]/P0001 ,
		_w37524_,
		_w37534_
	);
	LUT2 #(
		.INIT('h4)
	) name33488 (
		_w37350_,
		_w37524_,
		_w37535_
	);
	LUT2 #(
		.INIT('h1)
	) name33489 (
		_w37534_,
		_w37535_,
		_w37536_
	);
	LUT2 #(
		.INIT('h2)
	) name33490 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][5]/P0001 ,
		_w37524_,
		_w37537_
	);
	LUT2 #(
		.INIT('h4)
	) name33491 (
		_w37265_,
		_w37524_,
		_w37538_
	);
	LUT2 #(
		.INIT('h1)
	) name33492 (
		_w37537_,
		_w37538_,
		_w37539_
	);
	LUT2 #(
		.INIT('h2)
	) name33493 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][4]/P0001 ,
		_w37524_,
		_w37540_
	);
	LUT2 #(
		.INIT('h4)
	) name33494 (
		_w37274_,
		_w37524_,
		_w37541_
	);
	LUT2 #(
		.INIT('h1)
	) name33495 (
		_w37540_,
		_w37541_,
		_w37542_
	);
	LUT2 #(
		.INIT('h2)
	) name33496 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][3]/P0001 ,
		_w37524_,
		_w37543_
	);
	LUT2 #(
		.INIT('h4)
	) name33497 (
		_w37283_,
		_w37524_,
		_w37544_
	);
	LUT2 #(
		.INIT('h1)
	) name33498 (
		_w37543_,
		_w37544_,
		_w37545_
	);
	LUT2 #(
		.INIT('h2)
	) name33499 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][2]/P0001 ,
		_w37524_,
		_w37546_
	);
	LUT2 #(
		.INIT('h4)
	) name33500 (
		_w37362_,
		_w37524_,
		_w37547_
	);
	LUT2 #(
		.INIT('h1)
	) name33501 (
		_w37546_,
		_w37547_,
		_w37548_
	);
	LUT2 #(
		.INIT('h2)
	) name33502 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][1]/P0001 ,
		_w37524_,
		_w37549_
	);
	LUT2 #(
		.INIT('h4)
	) name33503 (
		_w37292_,
		_w37524_,
		_w37550_
	);
	LUT2 #(
		.INIT('h1)
	) name33504 (
		_w37549_,
		_w37550_,
		_w37551_
	);
	LUT2 #(
		.INIT('h2)
	) name33505 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][13]/P0001 ,
		_w37524_,
		_w37552_
	);
	LUT2 #(
		.INIT('h4)
	) name33506 (
		_w37374_,
		_w37524_,
		_w37553_
	);
	LUT2 #(
		.INIT('h1)
	) name33507 (
		_w37552_,
		_w37553_,
		_w37554_
	);
	LUT2 #(
		.INIT('h2)
	) name33508 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][12]/P0001 ,
		_w37524_,
		_w37555_
	);
	LUT2 #(
		.INIT('h4)
	) name33509 (
		_w37383_,
		_w37524_,
		_w37556_
	);
	LUT2 #(
		.INIT('h1)
	) name33510 (
		_w37555_,
		_w37556_,
		_w37557_
	);
	LUT2 #(
		.INIT('h2)
	) name33511 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][11]/P0001 ,
		_w37524_,
		_w37558_
	);
	LUT2 #(
		.INIT('h4)
	) name33512 (
		_w37301_,
		_w37524_,
		_w37559_
	);
	LUT2 #(
		.INIT('h1)
	) name33513 (
		_w37558_,
		_w37559_,
		_w37560_
	);
	LUT2 #(
		.INIT('h2)
	) name33514 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][10]/P0001 ,
		_w37524_,
		_w37561_
	);
	LUT2 #(
		.INIT('h4)
	) name33515 (
		_w37310_,
		_w37524_,
		_w37562_
	);
	LUT2 #(
		.INIT('h1)
	) name33516 (
		_w37561_,
		_w37562_,
		_w37563_
	);
	LUT2 #(
		.INIT('h4)
	) name33517 (
		_w37318_,
		_w37524_,
		_w37564_
	);
	LUT2 #(
		.INIT('h2)
	) name33518 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[12][0]/P0001 ,
		_w37524_,
		_w37565_
	);
	LUT2 #(
		.INIT('h1)
	) name33519 (
		_w37564_,
		_w37565_,
		_w37566_
	);
	LUT2 #(
		.INIT('h8)
	) name33520 (
		_w4202_,
		_w37248_,
		_w37567_
	);
	LUT2 #(
		.INIT('h2)
	) name33521 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][9]/P0001 ,
		_w37567_,
		_w37568_
	);
	LUT2 #(
		.INIT('h4)
	) name33522 (
		_w37329_,
		_w37567_,
		_w37569_
	);
	LUT2 #(
		.INIT('h1)
	) name33523 (
		_w37568_,
		_w37569_,
		_w37570_
	);
	LUT2 #(
		.INIT('h2)
	) name33524 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][8]/P0001 ,
		_w37567_,
		_w37571_
	);
	LUT2 #(
		.INIT('h4)
	) name33525 (
		_w37338_,
		_w37567_,
		_w37572_
	);
	LUT2 #(
		.INIT('h1)
	) name33526 (
		_w37571_,
		_w37572_,
		_w37573_
	);
	LUT2 #(
		.INIT('h2)
	) name33527 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][7]/P0001 ,
		_w37567_,
		_w37574_
	);
	LUT2 #(
		.INIT('h4)
	) name33528 (
		_w37256_,
		_w37567_,
		_w37575_
	);
	LUT2 #(
		.INIT('h1)
	) name33529 (
		_w37574_,
		_w37575_,
		_w37576_
	);
	LUT2 #(
		.INIT('h2)
	) name33530 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][6]/P0001 ,
		_w37567_,
		_w37577_
	);
	LUT2 #(
		.INIT('h4)
	) name33531 (
		_w37350_,
		_w37567_,
		_w37578_
	);
	LUT2 #(
		.INIT('h1)
	) name33532 (
		_w37577_,
		_w37578_,
		_w37579_
	);
	LUT2 #(
		.INIT('h2)
	) name33533 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][5]/P0001 ,
		_w37567_,
		_w37580_
	);
	LUT2 #(
		.INIT('h4)
	) name33534 (
		_w37265_,
		_w37567_,
		_w37581_
	);
	LUT2 #(
		.INIT('h1)
	) name33535 (
		_w37580_,
		_w37581_,
		_w37582_
	);
	LUT2 #(
		.INIT('h2)
	) name33536 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][4]/P0001 ,
		_w37567_,
		_w37583_
	);
	LUT2 #(
		.INIT('h4)
	) name33537 (
		_w37274_,
		_w37567_,
		_w37584_
	);
	LUT2 #(
		.INIT('h1)
	) name33538 (
		_w37583_,
		_w37584_,
		_w37585_
	);
	LUT2 #(
		.INIT('h2)
	) name33539 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][3]/P0001 ,
		_w37567_,
		_w37586_
	);
	LUT2 #(
		.INIT('h4)
	) name33540 (
		_w37283_,
		_w37567_,
		_w37587_
	);
	LUT2 #(
		.INIT('h1)
	) name33541 (
		_w37586_,
		_w37587_,
		_w37588_
	);
	LUT2 #(
		.INIT('h2)
	) name33542 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][2]/P0001 ,
		_w37567_,
		_w37589_
	);
	LUT2 #(
		.INIT('h4)
	) name33543 (
		_w37362_,
		_w37567_,
		_w37590_
	);
	LUT2 #(
		.INIT('h1)
	) name33544 (
		_w37589_,
		_w37590_,
		_w37591_
	);
	LUT2 #(
		.INIT('h2)
	) name33545 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][1]/P0001 ,
		_w37567_,
		_w37592_
	);
	LUT2 #(
		.INIT('h4)
	) name33546 (
		_w37292_,
		_w37567_,
		_w37593_
	);
	LUT2 #(
		.INIT('h1)
	) name33547 (
		_w37592_,
		_w37593_,
		_w37594_
	);
	LUT2 #(
		.INIT('h2)
	) name33548 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][13]/P0001 ,
		_w37567_,
		_w37595_
	);
	LUT2 #(
		.INIT('h4)
	) name33549 (
		_w37374_,
		_w37567_,
		_w37596_
	);
	LUT2 #(
		.INIT('h1)
	) name33550 (
		_w37595_,
		_w37596_,
		_w37597_
	);
	LUT2 #(
		.INIT('h2)
	) name33551 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][12]/P0001 ,
		_w37567_,
		_w37598_
	);
	LUT2 #(
		.INIT('h4)
	) name33552 (
		_w37383_,
		_w37567_,
		_w37599_
	);
	LUT2 #(
		.INIT('h1)
	) name33553 (
		_w37598_,
		_w37599_,
		_w37600_
	);
	LUT2 #(
		.INIT('h2)
	) name33554 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][11]/P0001 ,
		_w37567_,
		_w37601_
	);
	LUT2 #(
		.INIT('h4)
	) name33555 (
		_w37301_,
		_w37567_,
		_w37602_
	);
	LUT2 #(
		.INIT('h1)
	) name33556 (
		_w37601_,
		_w37602_,
		_w37603_
	);
	LUT2 #(
		.INIT('h2)
	) name33557 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][10]/P0001 ,
		_w37567_,
		_w37604_
	);
	LUT2 #(
		.INIT('h4)
	) name33558 (
		_w37310_,
		_w37567_,
		_w37605_
	);
	LUT2 #(
		.INIT('h1)
	) name33559 (
		_w37604_,
		_w37605_,
		_w37606_
	);
	LUT2 #(
		.INIT('h4)
	) name33560 (
		_w37318_,
		_w37567_,
		_w37607_
	);
	LUT2 #(
		.INIT('h2)
	) name33561 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[11][0]/P0001 ,
		_w37567_,
		_w37608_
	);
	LUT2 #(
		.INIT('h1)
	) name33562 (
		_w37607_,
		_w37608_,
		_w37609_
	);
	LUT2 #(
		.INIT('h8)
	) name33563 (
		_w4228_,
		_w37248_,
		_w37610_
	);
	LUT2 #(
		.INIT('h2)
	) name33564 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][9]/P0001 ,
		_w37610_,
		_w37611_
	);
	LUT2 #(
		.INIT('h4)
	) name33565 (
		_w37329_,
		_w37610_,
		_w37612_
	);
	LUT2 #(
		.INIT('h1)
	) name33566 (
		_w37611_,
		_w37612_,
		_w37613_
	);
	LUT2 #(
		.INIT('h2)
	) name33567 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][8]/P0001 ,
		_w37610_,
		_w37614_
	);
	LUT2 #(
		.INIT('h4)
	) name33568 (
		_w37338_,
		_w37610_,
		_w37615_
	);
	LUT2 #(
		.INIT('h1)
	) name33569 (
		_w37614_,
		_w37615_,
		_w37616_
	);
	LUT2 #(
		.INIT('h2)
	) name33570 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][7]/P0001 ,
		_w37610_,
		_w37617_
	);
	LUT2 #(
		.INIT('h4)
	) name33571 (
		_w37256_,
		_w37610_,
		_w37618_
	);
	LUT2 #(
		.INIT('h1)
	) name33572 (
		_w37617_,
		_w37618_,
		_w37619_
	);
	LUT2 #(
		.INIT('h2)
	) name33573 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][6]/P0001 ,
		_w37610_,
		_w37620_
	);
	LUT2 #(
		.INIT('h4)
	) name33574 (
		_w37350_,
		_w37610_,
		_w37621_
	);
	LUT2 #(
		.INIT('h1)
	) name33575 (
		_w37620_,
		_w37621_,
		_w37622_
	);
	LUT2 #(
		.INIT('h2)
	) name33576 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][5]/P0001 ,
		_w37610_,
		_w37623_
	);
	LUT2 #(
		.INIT('h4)
	) name33577 (
		_w37265_,
		_w37610_,
		_w37624_
	);
	LUT2 #(
		.INIT('h1)
	) name33578 (
		_w37623_,
		_w37624_,
		_w37625_
	);
	LUT2 #(
		.INIT('h2)
	) name33579 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][4]/P0001 ,
		_w37610_,
		_w37626_
	);
	LUT2 #(
		.INIT('h4)
	) name33580 (
		_w37274_,
		_w37610_,
		_w37627_
	);
	LUT2 #(
		.INIT('h1)
	) name33581 (
		_w37626_,
		_w37627_,
		_w37628_
	);
	LUT2 #(
		.INIT('h2)
	) name33582 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][3]/P0001 ,
		_w37610_,
		_w37629_
	);
	LUT2 #(
		.INIT('h4)
	) name33583 (
		_w37283_,
		_w37610_,
		_w37630_
	);
	LUT2 #(
		.INIT('h1)
	) name33584 (
		_w37629_,
		_w37630_,
		_w37631_
	);
	LUT2 #(
		.INIT('h2)
	) name33585 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][2]/P0001 ,
		_w37610_,
		_w37632_
	);
	LUT2 #(
		.INIT('h4)
	) name33586 (
		_w37362_,
		_w37610_,
		_w37633_
	);
	LUT2 #(
		.INIT('h1)
	) name33587 (
		_w37632_,
		_w37633_,
		_w37634_
	);
	LUT2 #(
		.INIT('h2)
	) name33588 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][1]/P0001 ,
		_w37610_,
		_w37635_
	);
	LUT2 #(
		.INIT('h4)
	) name33589 (
		_w37292_,
		_w37610_,
		_w37636_
	);
	LUT2 #(
		.INIT('h1)
	) name33590 (
		_w37635_,
		_w37636_,
		_w37637_
	);
	LUT2 #(
		.INIT('h2)
	) name33591 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][13]/P0001 ,
		_w37610_,
		_w37638_
	);
	LUT2 #(
		.INIT('h4)
	) name33592 (
		_w37374_,
		_w37610_,
		_w37639_
	);
	LUT2 #(
		.INIT('h1)
	) name33593 (
		_w37638_,
		_w37639_,
		_w37640_
	);
	LUT2 #(
		.INIT('h2)
	) name33594 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][12]/P0001 ,
		_w37610_,
		_w37641_
	);
	LUT2 #(
		.INIT('h4)
	) name33595 (
		_w37383_,
		_w37610_,
		_w37642_
	);
	LUT2 #(
		.INIT('h1)
	) name33596 (
		_w37641_,
		_w37642_,
		_w37643_
	);
	LUT2 #(
		.INIT('h2)
	) name33597 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][11]/P0001 ,
		_w37610_,
		_w37644_
	);
	LUT2 #(
		.INIT('h4)
	) name33598 (
		_w37301_,
		_w37610_,
		_w37645_
	);
	LUT2 #(
		.INIT('h1)
	) name33599 (
		_w37644_,
		_w37645_,
		_w37646_
	);
	LUT2 #(
		.INIT('h2)
	) name33600 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][10]/P0001 ,
		_w37610_,
		_w37647_
	);
	LUT2 #(
		.INIT('h4)
	) name33601 (
		_w37310_,
		_w37610_,
		_w37648_
	);
	LUT2 #(
		.INIT('h1)
	) name33602 (
		_w37647_,
		_w37648_,
		_w37649_
	);
	LUT2 #(
		.INIT('h4)
	) name33603 (
		_w37318_,
		_w37610_,
		_w37650_
	);
	LUT2 #(
		.INIT('h2)
	) name33604 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[10][0]/P0001 ,
		_w37610_,
		_w37651_
	);
	LUT2 #(
		.INIT('h1)
	) name33605 (
		_w37650_,
		_w37651_,
		_w37652_
	);
	LUT2 #(
		.INIT('h4)
	) name33606 (
		_w36440_,
		_w36603_,
		_w37653_
	);
	LUT2 #(
		.INIT('h2)
	) name33607 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][9]/P0001 ,
		_w37653_,
		_w37654_
	);
	LUT2 #(
		.INIT('h4)
	) name33608 (
		_w37329_,
		_w37653_,
		_w37655_
	);
	LUT2 #(
		.INIT('h1)
	) name33609 (
		_w37654_,
		_w37655_,
		_w37656_
	);
	LUT2 #(
		.INIT('h2)
	) name33610 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][8]/P0001 ,
		_w37653_,
		_w37657_
	);
	LUT2 #(
		.INIT('h4)
	) name33611 (
		_w37338_,
		_w37653_,
		_w37658_
	);
	LUT2 #(
		.INIT('h1)
	) name33612 (
		_w37657_,
		_w37658_,
		_w37659_
	);
	LUT2 #(
		.INIT('h2)
	) name33613 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][7]/P0001 ,
		_w37653_,
		_w37660_
	);
	LUT2 #(
		.INIT('h4)
	) name33614 (
		_w37256_,
		_w37653_,
		_w37661_
	);
	LUT2 #(
		.INIT('h1)
	) name33615 (
		_w37660_,
		_w37661_,
		_w37662_
	);
	LUT2 #(
		.INIT('h2)
	) name33616 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][6]/P0001 ,
		_w37653_,
		_w37663_
	);
	LUT2 #(
		.INIT('h4)
	) name33617 (
		_w37350_,
		_w37653_,
		_w37664_
	);
	LUT2 #(
		.INIT('h1)
	) name33618 (
		_w37663_,
		_w37664_,
		_w37665_
	);
	LUT2 #(
		.INIT('h2)
	) name33619 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][5]/P0001 ,
		_w37653_,
		_w37666_
	);
	LUT2 #(
		.INIT('h4)
	) name33620 (
		_w37265_,
		_w37653_,
		_w37667_
	);
	LUT2 #(
		.INIT('h1)
	) name33621 (
		_w37666_,
		_w37667_,
		_w37668_
	);
	LUT2 #(
		.INIT('h2)
	) name33622 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][4]/P0001 ,
		_w37653_,
		_w37669_
	);
	LUT2 #(
		.INIT('h4)
	) name33623 (
		_w37274_,
		_w37653_,
		_w37670_
	);
	LUT2 #(
		.INIT('h1)
	) name33624 (
		_w37669_,
		_w37670_,
		_w37671_
	);
	LUT2 #(
		.INIT('h2)
	) name33625 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][3]/P0001 ,
		_w37653_,
		_w37672_
	);
	LUT2 #(
		.INIT('h4)
	) name33626 (
		_w37283_,
		_w37653_,
		_w37673_
	);
	LUT2 #(
		.INIT('h1)
	) name33627 (
		_w37672_,
		_w37673_,
		_w37674_
	);
	LUT2 #(
		.INIT('h2)
	) name33628 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][2]/P0001 ,
		_w37653_,
		_w37675_
	);
	LUT2 #(
		.INIT('h4)
	) name33629 (
		_w37362_,
		_w37653_,
		_w37676_
	);
	LUT2 #(
		.INIT('h1)
	) name33630 (
		_w37675_,
		_w37676_,
		_w37677_
	);
	LUT2 #(
		.INIT('h2)
	) name33631 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][1]/P0001 ,
		_w37653_,
		_w37678_
	);
	LUT2 #(
		.INIT('h4)
	) name33632 (
		_w37292_,
		_w37653_,
		_w37679_
	);
	LUT2 #(
		.INIT('h1)
	) name33633 (
		_w37678_,
		_w37679_,
		_w37680_
	);
	LUT2 #(
		.INIT('h2)
	) name33634 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][13]/P0001 ,
		_w37653_,
		_w37681_
	);
	LUT2 #(
		.INIT('h4)
	) name33635 (
		_w37374_,
		_w37653_,
		_w37682_
	);
	LUT2 #(
		.INIT('h1)
	) name33636 (
		_w37681_,
		_w37682_,
		_w37683_
	);
	LUT2 #(
		.INIT('h2)
	) name33637 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][12]/P0001 ,
		_w37653_,
		_w37684_
	);
	LUT2 #(
		.INIT('h4)
	) name33638 (
		_w37383_,
		_w37653_,
		_w37685_
	);
	LUT2 #(
		.INIT('h1)
	) name33639 (
		_w37684_,
		_w37685_,
		_w37686_
	);
	LUT2 #(
		.INIT('h2)
	) name33640 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][11]/P0001 ,
		_w37653_,
		_w37687_
	);
	LUT2 #(
		.INIT('h4)
	) name33641 (
		_w37301_,
		_w37653_,
		_w37688_
	);
	LUT2 #(
		.INIT('h1)
	) name33642 (
		_w37687_,
		_w37688_,
		_w37689_
	);
	LUT2 #(
		.INIT('h2)
	) name33643 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][10]/P0001 ,
		_w37653_,
		_w37690_
	);
	LUT2 #(
		.INIT('h4)
	) name33644 (
		_w37310_,
		_w37653_,
		_w37691_
	);
	LUT2 #(
		.INIT('h1)
	) name33645 (
		_w37690_,
		_w37691_,
		_w37692_
	);
	LUT2 #(
		.INIT('h4)
	) name33646 (
		_w37318_,
		_w37653_,
		_w37693_
	);
	LUT2 #(
		.INIT('h2)
	) name33647 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[0][0]/P0001 ,
		_w37653_,
		_w37694_
	);
	LUT2 #(
		.INIT('h1)
	) name33648 (
		_w37693_,
		_w37694_,
		_w37695_
	);
	LUT2 #(
		.INIT('h2)
	) name33649 (
		\core_c_psq_Iact_E_reg[3]/NET0131 ,
		_w19477_,
		_w37696_
	);
	LUT2 #(
		.INIT('h8)
	) name33650 (
		_w19482_,
		_w33213_,
		_w37697_
	);
	LUT2 #(
		.INIT('h8)
	) name33651 (
		_w33215_,
		_w37697_,
		_w37698_
	);
	LUT2 #(
		.INIT('h8)
	) name33652 (
		_w19477_,
		_w37698_,
		_w37699_
	);
	LUT2 #(
		.INIT('h1)
	) name33653 (
		_w37696_,
		_w37699_,
		_w37700_
	);
	LUT2 #(
		.INIT('h2)
	) name33654 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][6]/P0001 ,
		_w37249_,
		_w37701_
	);
	LUT2 #(
		.INIT('h2)
	) name33655 (
		_w37249_,
		_w37350_,
		_w37702_
	);
	LUT2 #(
		.INIT('h1)
	) name33656 (
		_w37701_,
		_w37702_,
		_w37703_
	);
	LUT2 #(
		.INIT('h4)
	) name33657 (
		\sport1_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w23274_,
		_w37704_
	);
	LUT2 #(
		.INIT('h2)
	) name33658 (
		\sport1_txctl_Wcnt_reg[0]/NET0131 ,
		_w23264_,
		_w37705_
	);
	LUT2 #(
		.INIT('h1)
	) name33659 (
		_w36390_,
		_w37705_,
		_w37706_
	);
	LUT2 #(
		.INIT('h4)
	) name33660 (
		_w23274_,
		_w37706_,
		_w37707_
	);
	LUT2 #(
		.INIT('h1)
	) name33661 (
		_w37704_,
		_w37707_,
		_w37708_
	);
	LUT2 #(
		.INIT('h4)
	) name33662 (
		\sport1_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w23274_,
		_w37709_
	);
	LUT2 #(
		.INIT('h2)
	) name33663 (
		\sport1_txctl_Wcnt_reg[6]/NET0131 ,
		_w36395_,
		_w37710_
	);
	LUT2 #(
		.INIT('h2)
	) name33664 (
		_w36397_,
		_w37710_,
		_w37711_
	);
	LUT2 #(
		.INIT('h1)
	) name33665 (
		_w37709_,
		_w37711_,
		_w37712_
	);
	LUT2 #(
		.INIT('h2)
	) name33666 (
		\sport1_txctl_Wcnt_reg[3]/NET0131 ,
		_w36392_,
		_w37713_
	);
	LUT2 #(
		.INIT('h1)
	) name33667 (
		_w36393_,
		_w37713_,
		_w37714_
	);
	LUT2 #(
		.INIT('h4)
	) name33668 (
		_w23274_,
		_w37714_,
		_w37715_
	);
	LUT2 #(
		.INIT('h4)
	) name33669 (
		\sport1_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w23274_,
		_w37716_
	);
	LUT2 #(
		.INIT('h1)
	) name33670 (
		_w37715_,
		_w37716_,
		_w37717_
	);
	LUT2 #(
		.INIT('h2)
	) name33671 (
		\sport1_txctl_Wcnt_reg[2]/NET0131 ,
		_w36391_,
		_w37718_
	);
	LUT2 #(
		.INIT('h1)
	) name33672 (
		_w36392_,
		_w37718_,
		_w37719_
	);
	LUT2 #(
		.INIT('h4)
	) name33673 (
		_w23274_,
		_w37719_,
		_w37720_
	);
	LUT2 #(
		.INIT('h4)
	) name33674 (
		\sport1_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w23274_,
		_w37721_
	);
	LUT2 #(
		.INIT('h1)
	) name33675 (
		_w37720_,
		_w37721_,
		_w37722_
	);
	LUT2 #(
		.INIT('h4)
	) name33676 (
		\sport0_regs_MWORDreg_DO_reg[6]/NET0131 ,
		_w23286_,
		_w37723_
	);
	LUT2 #(
		.INIT('h2)
	) name33677 (
		\sport0_txctl_Wcnt_reg[6]/NET0131 ,
		_w36411_,
		_w37724_
	);
	LUT2 #(
		.INIT('h2)
	) name33678 (
		_w36413_,
		_w37724_,
		_w37725_
	);
	LUT2 #(
		.INIT('h1)
	) name33679 (
		_w37723_,
		_w37725_,
		_w37726_
	);
	LUT2 #(
		.INIT('h2)
	) name33680 (
		\sport0_txctl_Wcnt_reg[3]/NET0131 ,
		_w36408_,
		_w37727_
	);
	LUT2 #(
		.INIT('h1)
	) name33681 (
		_w36409_,
		_w37727_,
		_w37728_
	);
	LUT2 #(
		.INIT('h4)
	) name33682 (
		_w23286_,
		_w37728_,
		_w37729_
	);
	LUT2 #(
		.INIT('h4)
	) name33683 (
		\sport0_regs_MWORDreg_DO_reg[3]/NET0131 ,
		_w23286_,
		_w37730_
	);
	LUT2 #(
		.INIT('h1)
	) name33684 (
		_w37729_,
		_w37730_,
		_w37731_
	);
	LUT2 #(
		.INIT('h2)
	) name33685 (
		\sport0_txctl_Wcnt_reg[2]/NET0131 ,
		_w36407_,
		_w37732_
	);
	LUT2 #(
		.INIT('h1)
	) name33686 (
		_w36408_,
		_w37732_,
		_w37733_
	);
	LUT2 #(
		.INIT('h4)
	) name33687 (
		_w23286_,
		_w37733_,
		_w37734_
	);
	LUT2 #(
		.INIT('h4)
	) name33688 (
		\sport0_regs_MWORDreg_DO_reg[2]/NET0131 ,
		_w23286_,
		_w37735_
	);
	LUT2 #(
		.INIT('h1)
	) name33689 (
		_w37734_,
		_w37735_,
		_w37736_
	);
	LUT2 #(
		.INIT('h4)
	) name33690 (
		\sport0_regs_MWORDreg_DO_reg[0]/NET0131 ,
		_w23286_,
		_w37737_
	);
	LUT2 #(
		.INIT('h2)
	) name33691 (
		\sport0_txctl_Wcnt_reg[0]/NET0131 ,
		_w23276_,
		_w37738_
	);
	LUT2 #(
		.INIT('h1)
	) name33692 (
		_w36406_,
		_w37738_,
		_w37739_
	);
	LUT2 #(
		.INIT('h4)
	) name33693 (
		_w23286_,
		_w37739_,
		_w37740_
	);
	LUT2 #(
		.INIT('h1)
	) name33694 (
		_w37737_,
		_w37740_,
		_w37741_
	);
	LUT2 #(
		.INIT('h1)
	) name33695 (
		_w20068_,
		_w32454_,
		_w37742_
	);
	LUT2 #(
		.INIT('h4)
	) name33696 (
		_w32483_,
		_w37742_,
		_w37743_
	);
	LUT2 #(
		.INIT('h1)
	) name33697 (
		\idma_DOVL_reg[9]/NET0131 ,
		_w37742_,
		_w37744_
	);
	LUT2 #(
		.INIT('h1)
	) name33698 (
		_w37743_,
		_w37744_,
		_w37745_
	);
	LUT2 #(
		.INIT('h4)
	) name33699 (
		_w32458_,
		_w37742_,
		_w37746_
	);
	LUT2 #(
		.INIT('h1)
	) name33700 (
		\idma_DOVL_reg[8]/NET0131 ,
		_w37742_,
		_w37747_
	);
	LUT2 #(
		.INIT('h1)
	) name33701 (
		_w37746_,
		_w37747_,
		_w37748_
	);
	LUT2 #(
		.INIT('h4)
	) name33702 (
		_w32520_,
		_w37742_,
		_w37749_
	);
	LUT2 #(
		.INIT('h1)
	) name33703 (
		\idma_DOVL_reg[10]/NET0131 ,
		_w37742_,
		_w37750_
	);
	LUT2 #(
		.INIT('h1)
	) name33704 (
		_w37749_,
		_w37750_,
		_w37751_
	);
	LUT2 #(
		.INIT('h4)
	) name33705 (
		_w32512_,
		_w37742_,
		_w37752_
	);
	LUT2 #(
		.INIT('h1)
	) name33706 (
		\idma_DOVL_reg[11]/NET0131 ,
		_w37742_,
		_w37753_
	);
	LUT2 #(
		.INIT('h1)
	) name33707 (
		_w37752_,
		_w37753_,
		_w37754_
	);
	LUT2 #(
		.INIT('h2)
	) name33708 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][12]/P0001 ,
		_w37249_,
		_w37755_
	);
	LUT2 #(
		.INIT('h2)
	) name33709 (
		_w37249_,
		_w37383_,
		_w37756_
	);
	LUT2 #(
		.INIT('h1)
	) name33710 (
		_w37755_,
		_w37756_,
		_w37757_
	);
	LUT2 #(
		.INIT('h2)
	) name33711 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][13]/P0001 ,
		_w37249_,
		_w37758_
	);
	LUT2 #(
		.INIT('h2)
	) name33712 (
		_w37249_,
		_w37374_,
		_w37759_
	);
	LUT2 #(
		.INIT('h1)
	) name33713 (
		_w37758_,
		_w37759_,
		_w37760_
	);
	LUT2 #(
		.INIT('h2)
	) name33714 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][5]/P0001 ,
		_w37322_,
		_w37761_
	);
	LUT2 #(
		.INIT('h4)
	) name33715 (
		_w37265_,
		_w37322_,
		_w37762_
	);
	LUT2 #(
		.INIT('h1)
	) name33716 (
		_w37761_,
		_w37762_,
		_w37763_
	);
	LUT2 #(
		.INIT('h2)
	) name33717 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][2]/P0001 ,
		_w37249_,
		_w37764_
	);
	LUT2 #(
		.INIT('h2)
	) name33718 (
		_w37249_,
		_w37362_,
		_w37765_
	);
	LUT2 #(
		.INIT('h1)
	) name33719 (
		_w37764_,
		_w37765_,
		_w37766_
	);
	LUT2 #(
		.INIT('h8)
	) name33720 (
		_w4220_,
		_w37248_,
		_w37767_
	);
	LUT2 #(
		.INIT('h2)
	) name33721 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][9]/P0001 ,
		_w37767_,
		_w37768_
	);
	LUT2 #(
		.INIT('h4)
	) name33722 (
		_w37329_,
		_w37767_,
		_w37769_
	);
	LUT2 #(
		.INIT('h1)
	) name33723 (
		_w37768_,
		_w37769_,
		_w37770_
	);
	LUT2 #(
		.INIT('h2)
	) name33724 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][8]/P0001 ,
		_w37767_,
		_w37771_
	);
	LUT2 #(
		.INIT('h4)
	) name33725 (
		_w37338_,
		_w37767_,
		_w37772_
	);
	LUT2 #(
		.INIT('h1)
	) name33726 (
		_w37771_,
		_w37772_,
		_w37773_
	);
	LUT2 #(
		.INIT('h2)
	) name33727 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][7]/P0001 ,
		_w37767_,
		_w37774_
	);
	LUT2 #(
		.INIT('h4)
	) name33728 (
		_w37256_,
		_w37767_,
		_w37775_
	);
	LUT2 #(
		.INIT('h1)
	) name33729 (
		_w37774_,
		_w37775_,
		_w37776_
	);
	LUT2 #(
		.INIT('h2)
	) name33730 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][6]/P0001 ,
		_w37767_,
		_w37777_
	);
	LUT2 #(
		.INIT('h4)
	) name33731 (
		_w37350_,
		_w37767_,
		_w37778_
	);
	LUT2 #(
		.INIT('h1)
	) name33732 (
		_w37777_,
		_w37778_,
		_w37779_
	);
	LUT2 #(
		.INIT('h2)
	) name33733 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][5]/P0001 ,
		_w37767_,
		_w37780_
	);
	LUT2 #(
		.INIT('h4)
	) name33734 (
		_w37265_,
		_w37767_,
		_w37781_
	);
	LUT2 #(
		.INIT('h1)
	) name33735 (
		_w37780_,
		_w37781_,
		_w37782_
	);
	LUT2 #(
		.INIT('h2)
	) name33736 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][4]/P0001 ,
		_w37767_,
		_w37783_
	);
	LUT2 #(
		.INIT('h4)
	) name33737 (
		_w37274_,
		_w37767_,
		_w37784_
	);
	LUT2 #(
		.INIT('h1)
	) name33738 (
		_w37783_,
		_w37784_,
		_w37785_
	);
	LUT2 #(
		.INIT('h2)
	) name33739 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][3]/P0001 ,
		_w37767_,
		_w37786_
	);
	LUT2 #(
		.INIT('h4)
	) name33740 (
		_w37283_,
		_w37767_,
		_w37787_
	);
	LUT2 #(
		.INIT('h1)
	) name33741 (
		_w37786_,
		_w37787_,
		_w37788_
	);
	LUT2 #(
		.INIT('h2)
	) name33742 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][2]/P0001 ,
		_w37767_,
		_w37789_
	);
	LUT2 #(
		.INIT('h4)
	) name33743 (
		_w37362_,
		_w37767_,
		_w37790_
	);
	LUT2 #(
		.INIT('h1)
	) name33744 (
		_w37789_,
		_w37790_,
		_w37791_
	);
	LUT2 #(
		.INIT('h2)
	) name33745 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][1]/P0001 ,
		_w37767_,
		_w37792_
	);
	LUT2 #(
		.INIT('h4)
	) name33746 (
		_w37292_,
		_w37767_,
		_w37793_
	);
	LUT2 #(
		.INIT('h1)
	) name33747 (
		_w37792_,
		_w37793_,
		_w37794_
	);
	LUT2 #(
		.INIT('h2)
	) name33748 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][13]/P0001 ,
		_w37767_,
		_w37795_
	);
	LUT2 #(
		.INIT('h4)
	) name33749 (
		_w37374_,
		_w37767_,
		_w37796_
	);
	LUT2 #(
		.INIT('h1)
	) name33750 (
		_w37795_,
		_w37796_,
		_w37797_
	);
	LUT2 #(
		.INIT('h2)
	) name33751 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][12]/P0001 ,
		_w37767_,
		_w37798_
	);
	LUT2 #(
		.INIT('h4)
	) name33752 (
		_w37383_,
		_w37767_,
		_w37799_
	);
	LUT2 #(
		.INIT('h1)
	) name33753 (
		_w37798_,
		_w37799_,
		_w37800_
	);
	LUT2 #(
		.INIT('h2)
	) name33754 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][11]/P0001 ,
		_w37767_,
		_w37801_
	);
	LUT2 #(
		.INIT('h4)
	) name33755 (
		_w37301_,
		_w37767_,
		_w37802_
	);
	LUT2 #(
		.INIT('h1)
	) name33756 (
		_w37801_,
		_w37802_,
		_w37803_
	);
	LUT2 #(
		.INIT('h2)
	) name33757 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][10]/P0001 ,
		_w37767_,
		_w37804_
	);
	LUT2 #(
		.INIT('h4)
	) name33758 (
		_w37310_,
		_w37767_,
		_w37805_
	);
	LUT2 #(
		.INIT('h1)
	) name33759 (
		_w37804_,
		_w37805_,
		_w37806_
	);
	LUT2 #(
		.INIT('h4)
	) name33760 (
		_w37318_,
		_w37767_,
		_w37807_
	);
	LUT2 #(
		.INIT('h2)
	) name33761 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[9][0]/P0001 ,
		_w37767_,
		_w37808_
	);
	LUT2 #(
		.INIT('h1)
	) name33762 (
		_w37807_,
		_w37808_,
		_w37809_
	);
	LUT2 #(
		.INIT('h8)
	) name33763 (
		_w4209_,
		_w37248_,
		_w37810_
	);
	LUT2 #(
		.INIT('h2)
	) name33764 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][9]/P0001 ,
		_w37810_,
		_w37811_
	);
	LUT2 #(
		.INIT('h4)
	) name33765 (
		_w37329_,
		_w37810_,
		_w37812_
	);
	LUT2 #(
		.INIT('h1)
	) name33766 (
		_w37811_,
		_w37812_,
		_w37813_
	);
	LUT2 #(
		.INIT('h2)
	) name33767 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][8]/P0001 ,
		_w37810_,
		_w37814_
	);
	LUT2 #(
		.INIT('h4)
	) name33768 (
		_w37338_,
		_w37810_,
		_w37815_
	);
	LUT2 #(
		.INIT('h1)
	) name33769 (
		_w37814_,
		_w37815_,
		_w37816_
	);
	LUT2 #(
		.INIT('h2)
	) name33770 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][7]/P0001 ,
		_w37810_,
		_w37817_
	);
	LUT2 #(
		.INIT('h4)
	) name33771 (
		_w37256_,
		_w37810_,
		_w37818_
	);
	LUT2 #(
		.INIT('h1)
	) name33772 (
		_w37817_,
		_w37818_,
		_w37819_
	);
	LUT2 #(
		.INIT('h2)
	) name33773 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][6]/P0001 ,
		_w37810_,
		_w37820_
	);
	LUT2 #(
		.INIT('h4)
	) name33774 (
		_w37350_,
		_w37810_,
		_w37821_
	);
	LUT2 #(
		.INIT('h1)
	) name33775 (
		_w37820_,
		_w37821_,
		_w37822_
	);
	LUT2 #(
		.INIT('h2)
	) name33776 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][5]/P0001 ,
		_w37810_,
		_w37823_
	);
	LUT2 #(
		.INIT('h4)
	) name33777 (
		_w37265_,
		_w37810_,
		_w37824_
	);
	LUT2 #(
		.INIT('h1)
	) name33778 (
		_w37823_,
		_w37824_,
		_w37825_
	);
	LUT2 #(
		.INIT('h2)
	) name33779 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][4]/P0001 ,
		_w37810_,
		_w37826_
	);
	LUT2 #(
		.INIT('h4)
	) name33780 (
		_w37274_,
		_w37810_,
		_w37827_
	);
	LUT2 #(
		.INIT('h1)
	) name33781 (
		_w37826_,
		_w37827_,
		_w37828_
	);
	LUT2 #(
		.INIT('h2)
	) name33782 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][3]/P0001 ,
		_w37810_,
		_w37829_
	);
	LUT2 #(
		.INIT('h4)
	) name33783 (
		_w37283_,
		_w37810_,
		_w37830_
	);
	LUT2 #(
		.INIT('h1)
	) name33784 (
		_w37829_,
		_w37830_,
		_w37831_
	);
	LUT2 #(
		.INIT('h2)
	) name33785 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][2]/P0001 ,
		_w37810_,
		_w37832_
	);
	LUT2 #(
		.INIT('h4)
	) name33786 (
		_w37362_,
		_w37810_,
		_w37833_
	);
	LUT2 #(
		.INIT('h1)
	) name33787 (
		_w37832_,
		_w37833_,
		_w37834_
	);
	LUT2 #(
		.INIT('h2)
	) name33788 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][1]/P0001 ,
		_w37810_,
		_w37835_
	);
	LUT2 #(
		.INIT('h4)
	) name33789 (
		_w37292_,
		_w37810_,
		_w37836_
	);
	LUT2 #(
		.INIT('h1)
	) name33790 (
		_w37835_,
		_w37836_,
		_w37837_
	);
	LUT2 #(
		.INIT('h2)
	) name33791 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][13]/P0001 ,
		_w37810_,
		_w37838_
	);
	LUT2 #(
		.INIT('h4)
	) name33792 (
		_w37374_,
		_w37810_,
		_w37839_
	);
	LUT2 #(
		.INIT('h1)
	) name33793 (
		_w37838_,
		_w37839_,
		_w37840_
	);
	LUT2 #(
		.INIT('h2)
	) name33794 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][12]/P0001 ,
		_w37810_,
		_w37841_
	);
	LUT2 #(
		.INIT('h4)
	) name33795 (
		_w37383_,
		_w37810_,
		_w37842_
	);
	LUT2 #(
		.INIT('h1)
	) name33796 (
		_w37841_,
		_w37842_,
		_w37843_
	);
	LUT2 #(
		.INIT('h2)
	) name33797 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][11]/P0001 ,
		_w37810_,
		_w37844_
	);
	LUT2 #(
		.INIT('h4)
	) name33798 (
		_w37301_,
		_w37810_,
		_w37845_
	);
	LUT2 #(
		.INIT('h1)
	) name33799 (
		_w37844_,
		_w37845_,
		_w37846_
	);
	LUT2 #(
		.INIT('h2)
	) name33800 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][10]/P0001 ,
		_w37810_,
		_w37847_
	);
	LUT2 #(
		.INIT('h4)
	) name33801 (
		_w37310_,
		_w37810_,
		_w37848_
	);
	LUT2 #(
		.INIT('h1)
	) name33802 (
		_w37847_,
		_w37848_,
		_w37849_
	);
	LUT2 #(
		.INIT('h4)
	) name33803 (
		_w37318_,
		_w37810_,
		_w37850_
	);
	LUT2 #(
		.INIT('h2)
	) name33804 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[8][0]/P0001 ,
		_w37810_,
		_w37851_
	);
	LUT2 #(
		.INIT('h1)
	) name33805 (
		_w37850_,
		_w37851_,
		_w37852_
	);
	LUT2 #(
		.INIT('h8)
	) name33806 (
		_w4226_,
		_w37248_,
		_w37853_
	);
	LUT2 #(
		.INIT('h2)
	) name33807 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][9]/P0001 ,
		_w37853_,
		_w37854_
	);
	LUT2 #(
		.INIT('h4)
	) name33808 (
		_w37329_,
		_w37853_,
		_w37855_
	);
	LUT2 #(
		.INIT('h1)
	) name33809 (
		_w37854_,
		_w37855_,
		_w37856_
	);
	LUT2 #(
		.INIT('h2)
	) name33810 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][8]/P0001 ,
		_w37853_,
		_w37857_
	);
	LUT2 #(
		.INIT('h4)
	) name33811 (
		_w37338_,
		_w37853_,
		_w37858_
	);
	LUT2 #(
		.INIT('h1)
	) name33812 (
		_w37857_,
		_w37858_,
		_w37859_
	);
	LUT2 #(
		.INIT('h2)
	) name33813 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][7]/P0001 ,
		_w37853_,
		_w37860_
	);
	LUT2 #(
		.INIT('h4)
	) name33814 (
		_w37256_,
		_w37853_,
		_w37861_
	);
	LUT2 #(
		.INIT('h1)
	) name33815 (
		_w37860_,
		_w37861_,
		_w37862_
	);
	LUT2 #(
		.INIT('h2)
	) name33816 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][6]/P0001 ,
		_w37853_,
		_w37863_
	);
	LUT2 #(
		.INIT('h4)
	) name33817 (
		_w37350_,
		_w37853_,
		_w37864_
	);
	LUT2 #(
		.INIT('h1)
	) name33818 (
		_w37863_,
		_w37864_,
		_w37865_
	);
	LUT2 #(
		.INIT('h2)
	) name33819 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][5]/P0001 ,
		_w37853_,
		_w37866_
	);
	LUT2 #(
		.INIT('h4)
	) name33820 (
		_w37265_,
		_w37853_,
		_w37867_
	);
	LUT2 #(
		.INIT('h1)
	) name33821 (
		_w37866_,
		_w37867_,
		_w37868_
	);
	LUT2 #(
		.INIT('h2)
	) name33822 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][4]/P0001 ,
		_w37853_,
		_w37869_
	);
	LUT2 #(
		.INIT('h4)
	) name33823 (
		_w37274_,
		_w37853_,
		_w37870_
	);
	LUT2 #(
		.INIT('h1)
	) name33824 (
		_w37869_,
		_w37870_,
		_w37871_
	);
	LUT2 #(
		.INIT('h2)
	) name33825 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][3]/P0001 ,
		_w37853_,
		_w37872_
	);
	LUT2 #(
		.INIT('h4)
	) name33826 (
		_w37283_,
		_w37853_,
		_w37873_
	);
	LUT2 #(
		.INIT('h1)
	) name33827 (
		_w37872_,
		_w37873_,
		_w37874_
	);
	LUT2 #(
		.INIT('h2)
	) name33828 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][2]/P0001 ,
		_w37853_,
		_w37875_
	);
	LUT2 #(
		.INIT('h4)
	) name33829 (
		_w37362_,
		_w37853_,
		_w37876_
	);
	LUT2 #(
		.INIT('h1)
	) name33830 (
		_w37875_,
		_w37876_,
		_w37877_
	);
	LUT2 #(
		.INIT('h2)
	) name33831 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][1]/P0001 ,
		_w37853_,
		_w37878_
	);
	LUT2 #(
		.INIT('h4)
	) name33832 (
		_w37292_,
		_w37853_,
		_w37879_
	);
	LUT2 #(
		.INIT('h1)
	) name33833 (
		_w37878_,
		_w37879_,
		_w37880_
	);
	LUT2 #(
		.INIT('h2)
	) name33834 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][13]/P0001 ,
		_w37853_,
		_w37881_
	);
	LUT2 #(
		.INIT('h4)
	) name33835 (
		_w37374_,
		_w37853_,
		_w37882_
	);
	LUT2 #(
		.INIT('h1)
	) name33836 (
		_w37881_,
		_w37882_,
		_w37883_
	);
	LUT2 #(
		.INIT('h2)
	) name33837 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][12]/P0001 ,
		_w37853_,
		_w37884_
	);
	LUT2 #(
		.INIT('h4)
	) name33838 (
		_w37383_,
		_w37853_,
		_w37885_
	);
	LUT2 #(
		.INIT('h1)
	) name33839 (
		_w37884_,
		_w37885_,
		_w37886_
	);
	LUT2 #(
		.INIT('h2)
	) name33840 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][11]/P0001 ,
		_w37853_,
		_w37887_
	);
	LUT2 #(
		.INIT('h4)
	) name33841 (
		_w37301_,
		_w37853_,
		_w37888_
	);
	LUT2 #(
		.INIT('h1)
	) name33842 (
		_w37887_,
		_w37888_,
		_w37889_
	);
	LUT2 #(
		.INIT('h2)
	) name33843 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][10]/P0001 ,
		_w37853_,
		_w37890_
	);
	LUT2 #(
		.INIT('h4)
	) name33844 (
		_w37310_,
		_w37853_,
		_w37891_
	);
	LUT2 #(
		.INIT('h1)
	) name33845 (
		_w37890_,
		_w37891_,
		_w37892_
	);
	LUT2 #(
		.INIT('h4)
	) name33846 (
		_w37318_,
		_w37853_,
		_w37893_
	);
	LUT2 #(
		.INIT('h2)
	) name33847 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[7][0]/P0001 ,
		_w37853_,
		_w37894_
	);
	LUT2 #(
		.INIT('h1)
	) name33848 (
		_w37893_,
		_w37894_,
		_w37895_
	);
	LUT2 #(
		.INIT('h8)
	) name33849 (
		_w4213_,
		_w37248_,
		_w37896_
	);
	LUT2 #(
		.INIT('h2)
	) name33850 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][9]/P0001 ,
		_w37896_,
		_w37897_
	);
	LUT2 #(
		.INIT('h4)
	) name33851 (
		_w37329_,
		_w37896_,
		_w37898_
	);
	LUT2 #(
		.INIT('h1)
	) name33852 (
		_w37897_,
		_w37898_,
		_w37899_
	);
	LUT2 #(
		.INIT('h2)
	) name33853 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][8]/P0001 ,
		_w37896_,
		_w37900_
	);
	LUT2 #(
		.INIT('h4)
	) name33854 (
		_w37338_,
		_w37896_,
		_w37901_
	);
	LUT2 #(
		.INIT('h1)
	) name33855 (
		_w37900_,
		_w37901_,
		_w37902_
	);
	LUT2 #(
		.INIT('h2)
	) name33856 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][7]/P0001 ,
		_w37896_,
		_w37903_
	);
	LUT2 #(
		.INIT('h4)
	) name33857 (
		_w37256_,
		_w37896_,
		_w37904_
	);
	LUT2 #(
		.INIT('h1)
	) name33858 (
		_w37903_,
		_w37904_,
		_w37905_
	);
	LUT2 #(
		.INIT('h2)
	) name33859 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][6]/P0001 ,
		_w37896_,
		_w37906_
	);
	LUT2 #(
		.INIT('h4)
	) name33860 (
		_w37350_,
		_w37896_,
		_w37907_
	);
	LUT2 #(
		.INIT('h1)
	) name33861 (
		_w37906_,
		_w37907_,
		_w37908_
	);
	LUT2 #(
		.INIT('h2)
	) name33862 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][4]/P0001 ,
		_w37896_,
		_w37909_
	);
	LUT2 #(
		.INIT('h4)
	) name33863 (
		_w37274_,
		_w37896_,
		_w37910_
	);
	LUT2 #(
		.INIT('h1)
	) name33864 (
		_w37909_,
		_w37910_,
		_w37911_
	);
	LUT2 #(
		.INIT('h2)
	) name33865 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][3]/P0001 ,
		_w37896_,
		_w37912_
	);
	LUT2 #(
		.INIT('h4)
	) name33866 (
		_w37283_,
		_w37896_,
		_w37913_
	);
	LUT2 #(
		.INIT('h1)
	) name33867 (
		_w37912_,
		_w37913_,
		_w37914_
	);
	LUT2 #(
		.INIT('h2)
	) name33868 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][5]/P0001 ,
		_w37896_,
		_w37915_
	);
	LUT2 #(
		.INIT('h4)
	) name33869 (
		_w37265_,
		_w37896_,
		_w37916_
	);
	LUT2 #(
		.INIT('h1)
	) name33870 (
		_w37915_,
		_w37916_,
		_w37917_
	);
	LUT2 #(
		.INIT('h2)
	) name33871 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][2]/P0001 ,
		_w37896_,
		_w37918_
	);
	LUT2 #(
		.INIT('h4)
	) name33872 (
		_w37362_,
		_w37896_,
		_w37919_
	);
	LUT2 #(
		.INIT('h1)
	) name33873 (
		_w37918_,
		_w37919_,
		_w37920_
	);
	LUT2 #(
		.INIT('h2)
	) name33874 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][13]/P0001 ,
		_w37896_,
		_w37921_
	);
	LUT2 #(
		.INIT('h4)
	) name33875 (
		_w37374_,
		_w37896_,
		_w37922_
	);
	LUT2 #(
		.INIT('h1)
	) name33876 (
		_w37921_,
		_w37922_,
		_w37923_
	);
	LUT2 #(
		.INIT('h2)
	) name33877 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][1]/P0001 ,
		_w37896_,
		_w37924_
	);
	LUT2 #(
		.INIT('h4)
	) name33878 (
		_w37292_,
		_w37896_,
		_w37925_
	);
	LUT2 #(
		.INIT('h1)
	) name33879 (
		_w37924_,
		_w37925_,
		_w37926_
	);
	LUT2 #(
		.INIT('h2)
	) name33880 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][12]/P0001 ,
		_w37896_,
		_w37927_
	);
	LUT2 #(
		.INIT('h4)
	) name33881 (
		_w37383_,
		_w37896_,
		_w37928_
	);
	LUT2 #(
		.INIT('h1)
	) name33882 (
		_w37927_,
		_w37928_,
		_w37929_
	);
	LUT2 #(
		.INIT('h2)
	) name33883 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][11]/P0001 ,
		_w37896_,
		_w37930_
	);
	LUT2 #(
		.INIT('h4)
	) name33884 (
		_w37301_,
		_w37896_,
		_w37931_
	);
	LUT2 #(
		.INIT('h1)
	) name33885 (
		_w37930_,
		_w37931_,
		_w37932_
	);
	LUT2 #(
		.INIT('h2)
	) name33886 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][10]/P0001 ,
		_w37896_,
		_w37933_
	);
	LUT2 #(
		.INIT('h4)
	) name33887 (
		_w37310_,
		_w37896_,
		_w37934_
	);
	LUT2 #(
		.INIT('h1)
	) name33888 (
		_w37933_,
		_w37934_,
		_w37935_
	);
	LUT2 #(
		.INIT('h4)
	) name33889 (
		_w37318_,
		_w37896_,
		_w37936_
	);
	LUT2 #(
		.INIT('h2)
	) name33890 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[6][0]/P0001 ,
		_w37896_,
		_w37937_
	);
	LUT2 #(
		.INIT('h1)
	) name33891 (
		_w37936_,
		_w37937_,
		_w37938_
	);
	LUT2 #(
		.INIT('h8)
	) name33892 (
		_w4197_,
		_w37248_,
		_w37939_
	);
	LUT2 #(
		.INIT('h2)
	) name33893 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][9]/P0001 ,
		_w37939_,
		_w37940_
	);
	LUT2 #(
		.INIT('h4)
	) name33894 (
		_w37329_,
		_w37939_,
		_w37941_
	);
	LUT2 #(
		.INIT('h1)
	) name33895 (
		_w37940_,
		_w37941_,
		_w37942_
	);
	LUT2 #(
		.INIT('h2)
	) name33896 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][8]/P0001 ,
		_w37939_,
		_w37943_
	);
	LUT2 #(
		.INIT('h4)
	) name33897 (
		_w37338_,
		_w37939_,
		_w37944_
	);
	LUT2 #(
		.INIT('h1)
	) name33898 (
		_w37943_,
		_w37944_,
		_w37945_
	);
	LUT2 #(
		.INIT('h2)
	) name33899 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][7]/P0001 ,
		_w37939_,
		_w37946_
	);
	LUT2 #(
		.INIT('h4)
	) name33900 (
		_w37256_,
		_w37939_,
		_w37947_
	);
	LUT2 #(
		.INIT('h1)
	) name33901 (
		_w37946_,
		_w37947_,
		_w37948_
	);
	LUT2 #(
		.INIT('h2)
	) name33902 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][6]/P0001 ,
		_w37939_,
		_w37949_
	);
	LUT2 #(
		.INIT('h4)
	) name33903 (
		_w37350_,
		_w37939_,
		_w37950_
	);
	LUT2 #(
		.INIT('h1)
	) name33904 (
		_w37949_,
		_w37950_,
		_w37951_
	);
	LUT2 #(
		.INIT('h2)
	) name33905 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][5]/P0001 ,
		_w37939_,
		_w37952_
	);
	LUT2 #(
		.INIT('h4)
	) name33906 (
		_w37265_,
		_w37939_,
		_w37953_
	);
	LUT2 #(
		.INIT('h1)
	) name33907 (
		_w37952_,
		_w37953_,
		_w37954_
	);
	LUT2 #(
		.INIT('h2)
	) name33908 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][4]/P0001 ,
		_w37939_,
		_w37955_
	);
	LUT2 #(
		.INIT('h4)
	) name33909 (
		_w37274_,
		_w37939_,
		_w37956_
	);
	LUT2 #(
		.INIT('h1)
	) name33910 (
		_w37955_,
		_w37956_,
		_w37957_
	);
	LUT2 #(
		.INIT('h2)
	) name33911 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][3]/P0001 ,
		_w37939_,
		_w37958_
	);
	LUT2 #(
		.INIT('h4)
	) name33912 (
		_w37283_,
		_w37939_,
		_w37959_
	);
	LUT2 #(
		.INIT('h1)
	) name33913 (
		_w37958_,
		_w37959_,
		_w37960_
	);
	LUT2 #(
		.INIT('h2)
	) name33914 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][2]/P0001 ,
		_w37939_,
		_w37961_
	);
	LUT2 #(
		.INIT('h4)
	) name33915 (
		_w37362_,
		_w37939_,
		_w37962_
	);
	LUT2 #(
		.INIT('h1)
	) name33916 (
		_w37961_,
		_w37962_,
		_w37963_
	);
	LUT2 #(
		.INIT('h2)
	) name33917 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][1]/P0001 ,
		_w37939_,
		_w37964_
	);
	LUT2 #(
		.INIT('h4)
	) name33918 (
		_w37292_,
		_w37939_,
		_w37965_
	);
	LUT2 #(
		.INIT('h1)
	) name33919 (
		_w37964_,
		_w37965_,
		_w37966_
	);
	LUT2 #(
		.INIT('h2)
	) name33920 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][13]/P0001 ,
		_w37939_,
		_w37967_
	);
	LUT2 #(
		.INIT('h4)
	) name33921 (
		_w37374_,
		_w37939_,
		_w37968_
	);
	LUT2 #(
		.INIT('h1)
	) name33922 (
		_w37967_,
		_w37968_,
		_w37969_
	);
	LUT2 #(
		.INIT('h2)
	) name33923 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][12]/P0001 ,
		_w37939_,
		_w37970_
	);
	LUT2 #(
		.INIT('h4)
	) name33924 (
		_w37383_,
		_w37939_,
		_w37971_
	);
	LUT2 #(
		.INIT('h1)
	) name33925 (
		_w37970_,
		_w37971_,
		_w37972_
	);
	LUT2 #(
		.INIT('h2)
	) name33926 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][11]/P0001 ,
		_w37939_,
		_w37973_
	);
	LUT2 #(
		.INIT('h4)
	) name33927 (
		_w37301_,
		_w37939_,
		_w37974_
	);
	LUT2 #(
		.INIT('h1)
	) name33928 (
		_w37973_,
		_w37974_,
		_w37975_
	);
	LUT2 #(
		.INIT('h4)
	) name33929 (
		_w37318_,
		_w37939_,
		_w37976_
	);
	LUT2 #(
		.INIT('h2)
	) name33930 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][0]/P0001 ,
		_w37939_,
		_w37977_
	);
	LUT2 #(
		.INIT('h1)
	) name33931 (
		_w37976_,
		_w37977_,
		_w37978_
	);
	LUT2 #(
		.INIT('h2)
	) name33932 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[5][10]/P0001 ,
		_w37939_,
		_w37979_
	);
	LUT2 #(
		.INIT('h4)
	) name33933 (
		_w37310_,
		_w37939_,
		_w37980_
	);
	LUT2 #(
		.INIT('h1)
	) name33934 (
		_w37979_,
		_w37980_,
		_w37981_
	);
	LUT2 #(
		.INIT('h8)
	) name33935 (
		_w4200_,
		_w37248_,
		_w37982_
	);
	LUT2 #(
		.INIT('h2)
	) name33936 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][9]/P0001 ,
		_w37982_,
		_w37983_
	);
	LUT2 #(
		.INIT('h4)
	) name33937 (
		_w37329_,
		_w37982_,
		_w37984_
	);
	LUT2 #(
		.INIT('h1)
	) name33938 (
		_w37983_,
		_w37984_,
		_w37985_
	);
	LUT2 #(
		.INIT('h2)
	) name33939 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][8]/P0001 ,
		_w37982_,
		_w37986_
	);
	LUT2 #(
		.INIT('h4)
	) name33940 (
		_w37338_,
		_w37982_,
		_w37987_
	);
	LUT2 #(
		.INIT('h1)
	) name33941 (
		_w37986_,
		_w37987_,
		_w37988_
	);
	LUT2 #(
		.INIT('h2)
	) name33942 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][7]/P0001 ,
		_w37982_,
		_w37989_
	);
	LUT2 #(
		.INIT('h4)
	) name33943 (
		_w37256_,
		_w37982_,
		_w37990_
	);
	LUT2 #(
		.INIT('h1)
	) name33944 (
		_w37989_,
		_w37990_,
		_w37991_
	);
	LUT2 #(
		.INIT('h2)
	) name33945 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][6]/P0001 ,
		_w37982_,
		_w37992_
	);
	LUT2 #(
		.INIT('h4)
	) name33946 (
		_w37350_,
		_w37982_,
		_w37993_
	);
	LUT2 #(
		.INIT('h1)
	) name33947 (
		_w37992_,
		_w37993_,
		_w37994_
	);
	LUT2 #(
		.INIT('h2)
	) name33948 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][5]/P0001 ,
		_w37982_,
		_w37995_
	);
	LUT2 #(
		.INIT('h4)
	) name33949 (
		_w37265_,
		_w37982_,
		_w37996_
	);
	LUT2 #(
		.INIT('h1)
	) name33950 (
		_w37995_,
		_w37996_,
		_w37997_
	);
	LUT2 #(
		.INIT('h2)
	) name33951 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][4]/P0001 ,
		_w37982_,
		_w37998_
	);
	LUT2 #(
		.INIT('h4)
	) name33952 (
		_w37274_,
		_w37982_,
		_w37999_
	);
	LUT2 #(
		.INIT('h1)
	) name33953 (
		_w37998_,
		_w37999_,
		_w38000_
	);
	LUT2 #(
		.INIT('h2)
	) name33954 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][3]/P0001 ,
		_w37982_,
		_w38001_
	);
	LUT2 #(
		.INIT('h4)
	) name33955 (
		_w37283_,
		_w37982_,
		_w38002_
	);
	LUT2 #(
		.INIT('h1)
	) name33956 (
		_w38001_,
		_w38002_,
		_w38003_
	);
	LUT2 #(
		.INIT('h2)
	) name33957 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][2]/P0001 ,
		_w37982_,
		_w38004_
	);
	LUT2 #(
		.INIT('h4)
	) name33958 (
		_w37362_,
		_w37982_,
		_w38005_
	);
	LUT2 #(
		.INIT('h1)
	) name33959 (
		_w38004_,
		_w38005_,
		_w38006_
	);
	LUT2 #(
		.INIT('h2)
	) name33960 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][1]/P0001 ,
		_w37982_,
		_w38007_
	);
	LUT2 #(
		.INIT('h4)
	) name33961 (
		_w37292_,
		_w37982_,
		_w38008_
	);
	LUT2 #(
		.INIT('h1)
	) name33962 (
		_w38007_,
		_w38008_,
		_w38009_
	);
	LUT2 #(
		.INIT('h2)
	) name33963 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][13]/P0001 ,
		_w37982_,
		_w38010_
	);
	LUT2 #(
		.INIT('h4)
	) name33964 (
		_w37374_,
		_w37982_,
		_w38011_
	);
	LUT2 #(
		.INIT('h1)
	) name33965 (
		_w38010_,
		_w38011_,
		_w38012_
	);
	LUT2 #(
		.INIT('h2)
	) name33966 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][12]/P0001 ,
		_w37982_,
		_w38013_
	);
	LUT2 #(
		.INIT('h4)
	) name33967 (
		_w37383_,
		_w37982_,
		_w38014_
	);
	LUT2 #(
		.INIT('h1)
	) name33968 (
		_w38013_,
		_w38014_,
		_w38015_
	);
	LUT2 #(
		.INIT('h2)
	) name33969 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][11]/P0001 ,
		_w37982_,
		_w38016_
	);
	LUT2 #(
		.INIT('h4)
	) name33970 (
		_w37301_,
		_w37982_,
		_w38017_
	);
	LUT2 #(
		.INIT('h1)
	) name33971 (
		_w38016_,
		_w38017_,
		_w38018_
	);
	LUT2 #(
		.INIT('h2)
	) name33972 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][10]/P0001 ,
		_w37982_,
		_w38019_
	);
	LUT2 #(
		.INIT('h4)
	) name33973 (
		_w37310_,
		_w37982_,
		_w38020_
	);
	LUT2 #(
		.INIT('h1)
	) name33974 (
		_w38019_,
		_w38020_,
		_w38021_
	);
	LUT2 #(
		.INIT('h4)
	) name33975 (
		_w37318_,
		_w37982_,
		_w38022_
	);
	LUT2 #(
		.INIT('h2)
	) name33976 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[4][0]/P0001 ,
		_w37982_,
		_w38023_
	);
	LUT2 #(
		.INIT('h1)
	) name33977 (
		_w38022_,
		_w38023_,
		_w38024_
	);
	LUT2 #(
		.INIT('h8)
	) name33978 (
		_w4211_,
		_w37248_,
		_w38025_
	);
	LUT2 #(
		.INIT('h2)
	) name33979 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][9]/P0001 ,
		_w38025_,
		_w38026_
	);
	LUT2 #(
		.INIT('h4)
	) name33980 (
		_w37329_,
		_w38025_,
		_w38027_
	);
	LUT2 #(
		.INIT('h1)
	) name33981 (
		_w38026_,
		_w38027_,
		_w38028_
	);
	LUT2 #(
		.INIT('h2)
	) name33982 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][8]/P0001 ,
		_w38025_,
		_w38029_
	);
	LUT2 #(
		.INIT('h4)
	) name33983 (
		_w37338_,
		_w38025_,
		_w38030_
	);
	LUT2 #(
		.INIT('h1)
	) name33984 (
		_w38029_,
		_w38030_,
		_w38031_
	);
	LUT2 #(
		.INIT('h2)
	) name33985 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][7]/P0001 ,
		_w38025_,
		_w38032_
	);
	LUT2 #(
		.INIT('h4)
	) name33986 (
		_w37256_,
		_w38025_,
		_w38033_
	);
	LUT2 #(
		.INIT('h1)
	) name33987 (
		_w38032_,
		_w38033_,
		_w38034_
	);
	LUT2 #(
		.INIT('h2)
	) name33988 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[1][4]/P0001 ,
		_w37322_,
		_w38035_
	);
	LUT2 #(
		.INIT('h4)
	) name33989 (
		_w37274_,
		_w37322_,
		_w38036_
	);
	LUT2 #(
		.INIT('h1)
	) name33990 (
		_w38035_,
		_w38036_,
		_w38037_
	);
	LUT2 #(
		.INIT('h2)
	) name33991 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][6]/P0001 ,
		_w38025_,
		_w38038_
	);
	LUT2 #(
		.INIT('h4)
	) name33992 (
		_w37350_,
		_w38025_,
		_w38039_
	);
	LUT2 #(
		.INIT('h1)
	) name33993 (
		_w38038_,
		_w38039_,
		_w38040_
	);
	LUT2 #(
		.INIT('h2)
	) name33994 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][5]/P0001 ,
		_w38025_,
		_w38041_
	);
	LUT2 #(
		.INIT('h4)
	) name33995 (
		_w37265_,
		_w38025_,
		_w38042_
	);
	LUT2 #(
		.INIT('h1)
	) name33996 (
		_w38041_,
		_w38042_,
		_w38043_
	);
	LUT2 #(
		.INIT('h2)
	) name33997 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][4]/P0001 ,
		_w38025_,
		_w38044_
	);
	LUT2 #(
		.INIT('h4)
	) name33998 (
		_w37274_,
		_w38025_,
		_w38045_
	);
	LUT2 #(
		.INIT('h1)
	) name33999 (
		_w38044_,
		_w38045_,
		_w38046_
	);
	LUT2 #(
		.INIT('h2)
	) name34000 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][3]/P0001 ,
		_w38025_,
		_w38047_
	);
	LUT2 #(
		.INIT('h4)
	) name34001 (
		_w37283_,
		_w38025_,
		_w38048_
	);
	LUT2 #(
		.INIT('h1)
	) name34002 (
		_w38047_,
		_w38048_,
		_w38049_
	);
	LUT2 #(
		.INIT('h2)
	) name34003 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][2]/P0001 ,
		_w38025_,
		_w38050_
	);
	LUT2 #(
		.INIT('h4)
	) name34004 (
		_w37362_,
		_w38025_,
		_w38051_
	);
	LUT2 #(
		.INIT('h1)
	) name34005 (
		_w38050_,
		_w38051_,
		_w38052_
	);
	LUT2 #(
		.INIT('h2)
	) name34006 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][1]/P0001 ,
		_w38025_,
		_w38053_
	);
	LUT2 #(
		.INIT('h4)
	) name34007 (
		_w37292_,
		_w38025_,
		_w38054_
	);
	LUT2 #(
		.INIT('h1)
	) name34008 (
		_w38053_,
		_w38054_,
		_w38055_
	);
	LUT2 #(
		.INIT('h2)
	) name34009 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][13]/P0001 ,
		_w38025_,
		_w38056_
	);
	LUT2 #(
		.INIT('h4)
	) name34010 (
		_w37374_,
		_w38025_,
		_w38057_
	);
	LUT2 #(
		.INIT('h1)
	) name34011 (
		_w38056_,
		_w38057_,
		_w38058_
	);
	LUT2 #(
		.INIT('h2)
	) name34012 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][12]/P0001 ,
		_w38025_,
		_w38059_
	);
	LUT2 #(
		.INIT('h4)
	) name34013 (
		_w37383_,
		_w38025_,
		_w38060_
	);
	LUT2 #(
		.INIT('h1)
	) name34014 (
		_w38059_,
		_w38060_,
		_w38061_
	);
	LUT2 #(
		.INIT('h2)
	) name34015 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][11]/P0001 ,
		_w38025_,
		_w38062_
	);
	LUT2 #(
		.INIT('h4)
	) name34016 (
		_w37301_,
		_w38025_,
		_w38063_
	);
	LUT2 #(
		.INIT('h1)
	) name34017 (
		_w38062_,
		_w38063_,
		_w38064_
	);
	LUT2 #(
		.INIT('h2)
	) name34018 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][10]/P0001 ,
		_w38025_,
		_w38065_
	);
	LUT2 #(
		.INIT('h4)
	) name34019 (
		_w37310_,
		_w38025_,
		_w38066_
	);
	LUT2 #(
		.INIT('h1)
	) name34020 (
		_w38065_,
		_w38066_,
		_w38067_
	);
	LUT2 #(
		.INIT('h4)
	) name34021 (
		_w37318_,
		_w38025_,
		_w38068_
	);
	LUT2 #(
		.INIT('h2)
	) name34022 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[3][0]/P0001 ,
		_w38025_,
		_w38069_
	);
	LUT2 #(
		.INIT('h1)
	) name34023 (
		_w38068_,
		_w38069_,
		_w38070_
	);
	LUT2 #(
		.INIT('h2)
	) name34024 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][9]/P0001 ,
		_w37249_,
		_w38071_
	);
	LUT2 #(
		.INIT('h2)
	) name34025 (
		_w37249_,
		_w37329_,
		_w38072_
	);
	LUT2 #(
		.INIT('h1)
	) name34026 (
		_w38071_,
		_w38072_,
		_w38073_
	);
	LUT2 #(
		.INIT('h2)
	) name34027 (
		\core_c_psq_pcstk_cnts16x14_PCcell_reg[2][8]/P0001 ,
		_w37249_,
		_w38074_
	);
	LUT2 #(
		.INIT('h2)
	) name34028 (
		_w37249_,
		_w37338_,
		_w38075_
	);
	LUT2 #(
		.INIT('h1)
	) name34029 (
		_w38074_,
		_w38075_,
		_w38076_
	);
	LUT2 #(
		.INIT('h4)
	) name34030 (
		_w32541_,
		_w37742_,
		_w38077_
	);
	LUT2 #(
		.INIT('h1)
	) name34031 (
		\idma_DOVL_reg[7]/NET0131 ,
		_w37742_,
		_w38078_
	);
	LUT2 #(
		.INIT('h1)
	) name34032 (
		_w38077_,
		_w38078_,
		_w38079_
	);
	LUT2 #(
		.INIT('h4)
	) name34033 (
		_w32557_,
		_w37742_,
		_w38080_
	);
	LUT2 #(
		.INIT('h1)
	) name34034 (
		\idma_DOVL_reg[6]/NET0131 ,
		_w37742_,
		_w38081_
	);
	LUT2 #(
		.INIT('h1)
	) name34035 (
		_w38080_,
		_w38081_,
		_w38082_
	);
	LUT2 #(
		.INIT('h4)
	) name34036 (
		_w32549_,
		_w37742_,
		_w38083_
	);
	LUT2 #(
		.INIT('h1)
	) name34037 (
		\idma_DOVL_reg[5]/NET0131 ,
		_w37742_,
		_w38084_
	);
	LUT2 #(
		.INIT('h1)
	) name34038 (
		_w38083_,
		_w38084_,
		_w38085_
	);
	LUT2 #(
		.INIT('h4)
	) name34039 (
		_w32573_,
		_w37742_,
		_w38086_
	);
	LUT2 #(
		.INIT('h1)
	) name34040 (
		\idma_DOVL_reg[3]/NET0131 ,
		_w37742_,
		_w38087_
	);
	LUT2 #(
		.INIT('h1)
	) name34041 (
		_w38086_,
		_w38087_,
		_w38088_
	);
	LUT2 #(
		.INIT('h4)
	) name34042 (
		_w32565_,
		_w37742_,
		_w38089_
	);
	LUT2 #(
		.INIT('h1)
	) name34043 (
		\idma_DOVL_reg[4]/NET0131 ,
		_w37742_,
		_w38090_
	);
	LUT2 #(
		.INIT('h1)
	) name34044 (
		_w38089_,
		_w38090_,
		_w38091_
	);
	LUT2 #(
		.INIT('h4)
	) name34045 (
		_w32581_,
		_w37742_,
		_w38092_
	);
	LUT2 #(
		.INIT('h1)
	) name34046 (
		\idma_DOVL_reg[2]/NET0131 ,
		_w37742_,
		_w38093_
	);
	LUT2 #(
		.INIT('h1)
	) name34047 (
		_w38092_,
		_w38093_,
		_w38094_
	);
	LUT2 #(
		.INIT('h4)
	) name34048 (
		_w32677_,
		_w37742_,
		_w38095_
	);
	LUT2 #(
		.INIT('h1)
	) name34049 (
		\idma_DOVL_reg[1]/NET0131 ,
		_w37742_,
		_w38096_
	);
	LUT2 #(
		.INIT('h1)
	) name34050 (
		_w38095_,
		_w38096_,
		_w38097_
	);
	LUT2 #(
		.INIT('h4)
	) name34051 (
		_w32589_,
		_w37742_,
		_w38098_
	);
	LUT2 #(
		.INIT('h1)
	) name34052 (
		\idma_DOVL_reg[0]/NET0131 ,
		_w37742_,
		_w38099_
	);
	LUT2 #(
		.INIT('h1)
	) name34053 (
		_w38098_,
		_w38099_,
		_w38100_
	);
	LUT2 #(
		.INIT('h8)
	) name34054 (
		\sport0_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w18233_,
		_w38101_
	);
	LUT2 #(
		.INIT('h8)
	) name34055 (
		_w11265_,
		_w18237_,
		_w38102_
	);
	LUT2 #(
		.INIT('h1)
	) name34056 (
		_w38101_,
		_w38102_,
		_w38103_
	);
	LUT2 #(
		.INIT('h8)
	) name34057 (
		\sport0_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w18233_,
		_w38104_
	);
	LUT2 #(
		.INIT('h8)
	) name34058 (
		_w11525_,
		_w18237_,
		_w38105_
	);
	LUT2 #(
		.INIT('h1)
	) name34059 (
		_w38104_,
		_w38105_,
		_w38106_
	);
	LUT2 #(
		.INIT('h8)
	) name34060 (
		\sport0_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w18233_,
		_w38107_
	);
	LUT2 #(
		.INIT('h8)
	) name34061 (
		_w10911_,
		_w18237_,
		_w38108_
	);
	LUT2 #(
		.INIT('h1)
	) name34062 (
		_w38107_,
		_w38108_,
		_w38109_
	);
	LUT2 #(
		.INIT('h8)
	) name34063 (
		\sport0_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w18233_,
		_w38110_
	);
	LUT2 #(
		.INIT('h8)
	) name34064 (
		_w12743_,
		_w18237_,
		_w38111_
	);
	LUT2 #(
		.INIT('h1)
	) name34065 (
		_w38110_,
		_w38111_,
		_w38112_
	);
	LUT2 #(
		.INIT('h8)
	) name34066 (
		\ISCLK0_pad ,
		_w18233_,
		_w38113_
	);
	LUT2 #(
		.INIT('h8)
	) name34067 (
		_w12688_,
		_w18237_,
		_w38114_
	);
	LUT2 #(
		.INIT('h1)
	) name34068 (
		_w38113_,
		_w38114_,
		_w38115_
	);
	LUT2 #(
		.INIT('h2)
	) name34069 (
		\sport0_txctl_Wcnt_reg[4]/NET0131 ,
		_w36409_,
		_w38116_
	);
	LUT2 #(
		.INIT('h1)
	) name34070 (
		_w36410_,
		_w38116_,
		_w38117_
	);
	LUT2 #(
		.INIT('h4)
	) name34071 (
		_w23286_,
		_w38117_,
		_w38118_
	);
	LUT2 #(
		.INIT('h4)
	) name34072 (
		\sport0_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w23286_,
		_w38119_
	);
	LUT2 #(
		.INIT('h1)
	) name34073 (
		_w38118_,
		_w38119_,
		_w38120_
	);
	LUT2 #(
		.INIT('h2)
	) name34074 (
		\sport1_txctl_Wcnt_reg[4]/NET0131 ,
		_w36393_,
		_w38121_
	);
	LUT2 #(
		.INIT('h1)
	) name34075 (
		_w36394_,
		_w38121_,
		_w38122_
	);
	LUT2 #(
		.INIT('h4)
	) name34076 (
		_w23274_,
		_w38122_,
		_w38123_
	);
	LUT2 #(
		.INIT('h4)
	) name34077 (
		\sport1_regs_MWORDreg_DO_reg[4]/NET0131 ,
		_w23274_,
		_w38124_
	);
	LUT2 #(
		.INIT('h1)
	) name34078 (
		_w38123_,
		_w38124_,
		_w38125_
	);
	LUT2 #(
		.INIT('h1)
	) name34079 (
		\bdma_BEAD_reg[2]/NET0131 ,
		_w20769_,
		_w38126_
	);
	LUT2 #(
		.INIT('h1)
	) name34080 (
		_w20765_,
		_w33304_,
		_w38127_
	);
	LUT2 #(
		.INIT('h4)
	) name34081 (
		_w38126_,
		_w38127_,
		_w38128_
	);
	LUT2 #(
		.INIT('h8)
	) name34082 (
		_w8715_,
		_w20765_,
		_w38129_
	);
	LUT2 #(
		.INIT('h1)
	) name34083 (
		_w38128_,
		_w38129_,
		_w38130_
	);
	LUT2 #(
		.INIT('h2)
	) name34084 (
		\sport1_txctl_Wcnt_reg[1]/NET0131 ,
		_w36390_,
		_w38131_
	);
	LUT2 #(
		.INIT('h1)
	) name34085 (
		_w36391_,
		_w38131_,
		_w38132_
	);
	LUT2 #(
		.INIT('h4)
	) name34086 (
		_w23274_,
		_w38132_,
		_w38133_
	);
	LUT2 #(
		.INIT('h4)
	) name34087 (
		\sport1_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w23274_,
		_w38134_
	);
	LUT2 #(
		.INIT('h1)
	) name34088 (
		_w38133_,
		_w38134_,
		_w38135_
	);
	LUT2 #(
		.INIT('h2)
	) name34089 (
		\sport0_txctl_Wcnt_reg[1]/NET0131 ,
		_w36406_,
		_w38136_
	);
	LUT2 #(
		.INIT('h1)
	) name34090 (
		_w36407_,
		_w38136_,
		_w38137_
	);
	LUT2 #(
		.INIT('h4)
	) name34091 (
		_w23286_,
		_w38137_,
		_w38138_
	);
	LUT2 #(
		.INIT('h4)
	) name34092 (
		\sport0_regs_MWORDreg_DO_reg[1]/NET0131 ,
		_w23286_,
		_w38139_
	);
	LUT2 #(
		.INIT('h1)
	) name34093 (
		_w38138_,
		_w38139_,
		_w38140_
	);
	LUT2 #(
		.INIT('h1)
	) name34094 (
		\idma_RDcnt_reg[2]/NET0131 ,
		_w20828_,
		_w38141_
	);
	LUT2 #(
		.INIT('h8)
	) name34095 (
		\idma_RDcnt_reg[2]/NET0131 ,
		_w20828_,
		_w38142_
	);
	LUT2 #(
		.INIT('h1)
	) name34096 (
		_w38141_,
		_w38142_,
		_w38143_
	);
	LUT2 #(
		.INIT('h1)
	) name34097 (
		_w20824_,
		_w38143_,
		_w38144_
	);
	LUT2 #(
		.INIT('h4)
	) name34098 (
		\memc_usysr_DO_reg[6]/NET0131 ,
		_w20824_,
		_w38145_
	);
	LUT2 #(
		.INIT('h1)
	) name34099 (
		_w38144_,
		_w38145_,
		_w38146_
	);
	LUT2 #(
		.INIT('h8)
	) name34100 (
		\sport1_regs_SCTLreg_DO_reg[7]/NET0131 ,
		_w37215_,
		_w38147_
	);
	LUT2 #(
		.INIT('h8)
	) name34101 (
		_w11265_,
		_w37218_,
		_w38148_
	);
	LUT2 #(
		.INIT('h1)
	) name34102 (
		_w38147_,
		_w38148_,
		_w38149_
	);
	LUT2 #(
		.INIT('h8)
	) name34103 (
		\sport1_regs_SCTLreg_DO_reg[6]/NET0131 ,
		_w37215_,
		_w38150_
	);
	LUT2 #(
		.INIT('h8)
	) name34104 (
		_w11525_,
		_w37218_,
		_w38151_
	);
	LUT2 #(
		.INIT('h1)
	) name34105 (
		_w38150_,
		_w38151_,
		_w38152_
	);
	LUT2 #(
		.INIT('h8)
	) name34106 (
		\sport1_regs_SCTLreg_DO_reg[5]/NET0131 ,
		_w37215_,
		_w38153_
	);
	LUT2 #(
		.INIT('h8)
	) name34107 (
		_w10911_,
		_w37218_,
		_w38154_
	);
	LUT2 #(
		.INIT('h1)
	) name34108 (
		_w38153_,
		_w38154_,
		_w38155_
	);
	LUT2 #(
		.INIT('h8)
	) name34109 (
		\sport1_regs_SCTLreg_DO_reg[4]/NET0131 ,
		_w37215_,
		_w38156_
	);
	LUT2 #(
		.INIT('h8)
	) name34110 (
		_w10069_,
		_w37218_,
		_w38157_
	);
	LUT2 #(
		.INIT('h1)
	) name34111 (
		_w38156_,
		_w38157_,
		_w38158_
	);
	LUT2 #(
		.INIT('h8)
	) name34112 (
		\sport1_regs_SCTLreg_DO_reg[15]/NET0131 ,
		_w37215_,
		_w38159_
	);
	LUT2 #(
		.INIT('h2)
	) name34113 (
		_w12743_,
		_w37217_,
		_w38160_
	);
	LUT2 #(
		.INIT('h8)
	) name34114 (
		_w36073_,
		_w38160_,
		_w38161_
	);
	LUT2 #(
		.INIT('h1)
	) name34115 (
		_w38159_,
		_w38161_,
		_w38162_
	);
	LUT2 #(
		.INIT('h8)
	) name34116 (
		\ISCLK1_pad ,
		_w37215_,
		_w38163_
	);
	LUT2 #(
		.INIT('h2)
	) name34117 (
		_w12688_,
		_w37217_,
		_w38164_
	);
	LUT2 #(
		.INIT('h8)
	) name34118 (
		_w36073_,
		_w38164_,
		_w38165_
	);
	LUT2 #(
		.INIT('h1)
	) name34119 (
		_w38163_,
		_w38165_,
		_w38166_
	);
	LUT2 #(
		.INIT('h8)
	) name34120 (
		\sport1_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w37215_,
		_w38167_
	);
	LUT2 #(
		.INIT('h2)
	) name34121 (
		_w7340_,
		_w37217_,
		_w38168_
	);
	LUT2 #(
		.INIT('h8)
	) name34122 (
		_w36073_,
		_w38168_,
		_w38169_
	);
	LUT2 #(
		.INIT('h1)
	) name34123 (
		_w38167_,
		_w38169_,
		_w38170_
	);
	LUT2 #(
		.INIT('h8)
	) name34124 (
		\sport1_regs_SCTLreg_DO_reg[12]/NET0131 ,
		_w37215_,
		_w38171_
	);
	LUT2 #(
		.INIT('h2)
	) name34125 (
		_w9178_,
		_w37217_,
		_w38172_
	);
	LUT2 #(
		.INIT('h8)
	) name34126 (
		_w36073_,
		_w38172_,
		_w38173_
	);
	LUT2 #(
		.INIT('h1)
	) name34127 (
		_w38171_,
		_w38173_,
		_w38174_
	);
	LUT2 #(
		.INIT('h1)
	) name34128 (
		_w36075_,
		_w36108_,
		_w38175_
	);
	LUT2 #(
		.INIT('h8)
	) name34129 (
		\sport1_regs_FSDIVreg_DO_reg[9]/NET0131 ,
		_w38175_,
		_w38176_
	);
	LUT2 #(
		.INIT('h2)
	) name34130 (
		_w36108_,
		_w37217_,
		_w38177_
	);
	LUT2 #(
		.INIT('h8)
	) name34131 (
		_w10289_,
		_w38177_,
		_w38178_
	);
	LUT2 #(
		.INIT('h1)
	) name34132 (
		_w38176_,
		_w38178_,
		_w38179_
	);
	LUT2 #(
		.INIT('h8)
	) name34133 (
		\sport1_regs_FSDIVreg_DO_reg[8]/NET0131 ,
		_w38175_,
		_w38180_
	);
	LUT2 #(
		.INIT('h8)
	) name34134 (
		_w10638_,
		_w38177_,
		_w38181_
	);
	LUT2 #(
		.INIT('h1)
	) name34135 (
		_w38180_,
		_w38181_,
		_w38182_
	);
	LUT2 #(
		.INIT('h8)
	) name34136 (
		\sport1_regs_FSDIVreg_DO_reg[15]/NET0131 ,
		_w38175_,
		_w38183_
	);
	LUT2 #(
		.INIT('h8)
	) name34137 (
		_w36108_,
		_w38160_,
		_w38184_
	);
	LUT2 #(
		.INIT('h1)
	) name34138 (
		_w38183_,
		_w38184_,
		_w38185_
	);
	LUT2 #(
		.INIT('h8)
	) name34139 (
		\sport1_regs_FSDIVreg_DO_reg[14]/NET0131 ,
		_w38175_,
		_w38186_
	);
	LUT2 #(
		.INIT('h8)
	) name34140 (
		_w36108_,
		_w38164_,
		_w38187_
	);
	LUT2 #(
		.INIT('h1)
	) name34141 (
		_w38186_,
		_w38187_,
		_w38188_
	);
	LUT2 #(
		.INIT('h8)
	) name34142 (
		\sport1_regs_FSDIVreg_DO_reg[13]/NET0131 ,
		_w38175_,
		_w38189_
	);
	LUT2 #(
		.INIT('h8)
	) name34143 (
		_w36108_,
		_w38168_,
		_w38190_
	);
	LUT2 #(
		.INIT('h1)
	) name34144 (
		_w38189_,
		_w38190_,
		_w38191_
	);
	LUT2 #(
		.INIT('h8)
	) name34145 (
		\sport1_regs_FSDIVreg_DO_reg[12]/NET0131 ,
		_w38175_,
		_w38192_
	);
	LUT2 #(
		.INIT('h8)
	) name34146 (
		_w36108_,
		_w38172_,
		_w38193_
	);
	LUT2 #(
		.INIT('h1)
	) name34147 (
		_w38192_,
		_w38193_,
		_w38194_
	);
	LUT2 #(
		.INIT('h8)
	) name34148 (
		\sport1_regs_FSDIVreg_DO_reg[10]/NET0131 ,
		_w38175_,
		_w38195_
	);
	LUT2 #(
		.INIT('h8)
	) name34149 (
		_w7859_,
		_w38177_,
		_w38196_
	);
	LUT2 #(
		.INIT('h1)
	) name34150 (
		_w38195_,
		_w38196_,
		_w38197_
	);
	LUT2 #(
		.INIT('h8)
	) name34151 (
		\sport1_regs_FSDIVreg_DO_reg[11]/NET0131 ,
		_w38175_,
		_w38198_
	);
	LUT2 #(
		.INIT('h8)
	) name34152 (
		_w8460_,
		_w38177_,
		_w38199_
	);
	LUT2 #(
		.INIT('h1)
	) name34153 (
		_w38198_,
		_w38199_,
		_w38200_
	);
	LUT2 #(
		.INIT('h2)
	) name34154 (
		_w14699_,
		_w18220_,
		_w38201_
	);
	LUT2 #(
		.INIT('h2)
	) name34155 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][9]/P0001 ,
		_w38201_,
		_w38202_
	);
	LUT2 #(
		.INIT('h8)
	) name34156 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w38201_,
		_w38203_
	);
	LUT2 #(
		.INIT('h1)
	) name34157 (
		_w38202_,
		_w38203_,
		_w38204_
	);
	LUT2 #(
		.INIT('h2)
	) name34158 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][8]/P0001 ,
		_w38201_,
		_w38205_
	);
	LUT2 #(
		.INIT('h8)
	) name34159 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w38201_,
		_w38206_
	);
	LUT2 #(
		.INIT('h1)
	) name34160 (
		_w38205_,
		_w38206_,
		_w38207_
	);
	LUT2 #(
		.INIT('h2)
	) name34161 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][7]/P0001 ,
		_w38201_,
		_w38208_
	);
	LUT2 #(
		.INIT('h8)
	) name34162 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w38201_,
		_w38209_
	);
	LUT2 #(
		.INIT('h1)
	) name34163 (
		_w38208_,
		_w38209_,
		_w38210_
	);
	LUT2 #(
		.INIT('h2)
	) name34164 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][6]/P0001 ,
		_w38201_,
		_w38211_
	);
	LUT2 #(
		.INIT('h4)
	) name34165 (
		_w4174_,
		_w38201_,
		_w38212_
	);
	LUT2 #(
		.INIT('h1)
	) name34166 (
		_w38211_,
		_w38212_,
		_w38213_
	);
	LUT2 #(
		.INIT('h2)
	) name34167 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][5]/P0001 ,
		_w38201_,
		_w38214_
	);
	LUT2 #(
		.INIT('h8)
	) name34168 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w38201_,
		_w38215_
	);
	LUT2 #(
		.INIT('h1)
	) name34169 (
		_w38214_,
		_w38215_,
		_w38216_
	);
	LUT2 #(
		.INIT('h2)
	) name34170 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][4]/P0001 ,
		_w38201_,
		_w38217_
	);
	LUT2 #(
		.INIT('h8)
	) name34171 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w38201_,
		_w38218_
	);
	LUT2 #(
		.INIT('h1)
	) name34172 (
		_w38217_,
		_w38218_,
		_w38219_
	);
	LUT2 #(
		.INIT('h2)
	) name34173 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][3]/P0001 ,
		_w38201_,
		_w38220_
	);
	LUT2 #(
		.INIT('h8)
	) name34174 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w38201_,
		_w38221_
	);
	LUT2 #(
		.INIT('h1)
	) name34175 (
		_w38220_,
		_w38221_,
		_w38222_
	);
	LUT2 #(
		.INIT('h2)
	) name34176 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][2]/P0001 ,
		_w38201_,
		_w38223_
	);
	LUT2 #(
		.INIT('h8)
	) name34177 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w38201_,
		_w38224_
	);
	LUT2 #(
		.INIT('h1)
	) name34178 (
		_w38223_,
		_w38224_,
		_w38225_
	);
	LUT2 #(
		.INIT('h2)
	) name34179 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][24]/P0001 ,
		_w38201_,
		_w38226_
	);
	LUT2 #(
		.INIT('h8)
	) name34180 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w38201_,
		_w38227_
	);
	LUT2 #(
		.INIT('h1)
	) name34181 (
		_w38226_,
		_w38227_,
		_w38228_
	);
	LUT2 #(
		.INIT('h2)
	) name34182 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][23]/P0001 ,
		_w38201_,
		_w38229_
	);
	LUT2 #(
		.INIT('h8)
	) name34183 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w38201_,
		_w38230_
	);
	LUT2 #(
		.INIT('h1)
	) name34184 (
		_w38229_,
		_w38230_,
		_w38231_
	);
	LUT2 #(
		.INIT('h2)
	) name34185 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][22]/P0001 ,
		_w38201_,
		_w38232_
	);
	LUT2 #(
		.INIT('h8)
	) name34186 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w38201_,
		_w38233_
	);
	LUT2 #(
		.INIT('h1)
	) name34187 (
		_w38232_,
		_w38233_,
		_w38234_
	);
	LUT2 #(
		.INIT('h2)
	) name34188 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][21]/P0001 ,
		_w38201_,
		_w38235_
	);
	LUT2 #(
		.INIT('h8)
	) name34189 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w38201_,
		_w38236_
	);
	LUT2 #(
		.INIT('h1)
	) name34190 (
		_w38235_,
		_w38236_,
		_w38237_
	);
	LUT2 #(
		.INIT('h2)
	) name34191 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][20]/P0001 ,
		_w38201_,
		_w38238_
	);
	LUT2 #(
		.INIT('h8)
	) name34192 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w38201_,
		_w38239_
	);
	LUT2 #(
		.INIT('h1)
	) name34193 (
		_w38238_,
		_w38239_,
		_w38240_
	);
	LUT2 #(
		.INIT('h2)
	) name34194 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][1]/P0001 ,
		_w38201_,
		_w38241_
	);
	LUT2 #(
		.INIT('h8)
	) name34195 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w38201_,
		_w38242_
	);
	LUT2 #(
		.INIT('h1)
	) name34196 (
		_w38241_,
		_w38242_,
		_w38243_
	);
	LUT2 #(
		.INIT('h2)
	) name34197 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][19]/P0001 ,
		_w38201_,
		_w38244_
	);
	LUT2 #(
		.INIT('h8)
	) name34198 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w38201_,
		_w38245_
	);
	LUT2 #(
		.INIT('h1)
	) name34199 (
		_w38244_,
		_w38245_,
		_w38246_
	);
	LUT2 #(
		.INIT('h2)
	) name34200 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][18]/P0001 ,
		_w38201_,
		_w38247_
	);
	LUT2 #(
		.INIT('h8)
	) name34201 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w38201_,
		_w38248_
	);
	LUT2 #(
		.INIT('h1)
	) name34202 (
		_w38247_,
		_w38248_,
		_w38249_
	);
	LUT2 #(
		.INIT('h2)
	) name34203 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][17]/P0001 ,
		_w38201_,
		_w38250_
	);
	LUT2 #(
		.INIT('h8)
	) name34204 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w38201_,
		_w38251_
	);
	LUT2 #(
		.INIT('h1)
	) name34205 (
		_w38250_,
		_w38251_,
		_w38252_
	);
	LUT2 #(
		.INIT('h2)
	) name34206 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][16]/P0001 ,
		_w38201_,
		_w38253_
	);
	LUT2 #(
		.INIT('h8)
	) name34207 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w38201_,
		_w38254_
	);
	LUT2 #(
		.INIT('h1)
	) name34208 (
		_w38253_,
		_w38254_,
		_w38255_
	);
	LUT2 #(
		.INIT('h2)
	) name34209 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][15]/P0001 ,
		_w38201_,
		_w38256_
	);
	LUT2 #(
		.INIT('h8)
	) name34210 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w38201_,
		_w38257_
	);
	LUT2 #(
		.INIT('h1)
	) name34211 (
		_w38256_,
		_w38257_,
		_w38258_
	);
	LUT2 #(
		.INIT('h2)
	) name34212 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][14]/P0001 ,
		_w38201_,
		_w38259_
	);
	LUT2 #(
		.INIT('h8)
	) name34213 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w38201_,
		_w38260_
	);
	LUT2 #(
		.INIT('h1)
	) name34214 (
		_w38259_,
		_w38260_,
		_w38261_
	);
	LUT2 #(
		.INIT('h2)
	) name34215 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][13]/P0001 ,
		_w38201_,
		_w38262_
	);
	LUT2 #(
		.INIT('h8)
	) name34216 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w38201_,
		_w38263_
	);
	LUT2 #(
		.INIT('h1)
	) name34217 (
		_w38262_,
		_w38263_,
		_w38264_
	);
	LUT2 #(
		.INIT('h4)
	) name34218 (
		\sport0_rxctl_RXSHT_reg[6]/P0001 ,
		_w20868_,
		_w38265_
	);
	LUT2 #(
		.INIT('h8)
	) name34219 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20873_,
		_w38266_
	);
	LUT2 #(
		.INIT('h1)
	) name34220 (
		\sport0_rxctl_RX_reg[7]/P0001 ,
		_w31030_,
		_w38267_
	);
	LUT2 #(
		.INIT('h4)
	) name34221 (
		_w31042_,
		_w38267_,
		_w38268_
	);
	LUT2 #(
		.INIT('h2)
	) name34222 (
		_w31042_,
		_w38267_,
		_w38269_
	);
	LUT2 #(
		.INIT('h2)
	) name34223 (
		_w20875_,
		_w38268_,
		_w38270_
	);
	LUT2 #(
		.INIT('h4)
	) name34224 (
		_w38269_,
		_w38270_,
		_w38271_
	);
	LUT2 #(
		.INIT('h4)
	) name34225 (
		\sport0_rxctl_ldRX_cmp_reg/P0001 ,
		_w11525_,
		_w38272_
	);
	LUT2 #(
		.INIT('h1)
	) name34226 (
		_w20868_,
		_w38266_,
		_w38273_
	);
	LUT2 #(
		.INIT('h4)
	) name34227 (
		_w38272_,
		_w38273_,
		_w38274_
	);
	LUT2 #(
		.INIT('h4)
	) name34228 (
		_w38271_,
		_w38274_,
		_w38275_
	);
	LUT2 #(
		.INIT('h1)
	) name34229 (
		_w20871_,
		_w38265_,
		_w38276_
	);
	LUT2 #(
		.INIT('h4)
	) name34230 (
		_w38275_,
		_w38276_,
		_w38277_
	);
	LUT2 #(
		.INIT('h8)
	) name34231 (
		\sport0_rxctl_RX_reg[6]/P0001 ,
		_w20871_,
		_w38278_
	);
	LUT2 #(
		.INIT('h1)
	) name34232 (
		_w38277_,
		_w38278_,
		_w38279_
	);
	LUT2 #(
		.INIT('h2)
	) name34233 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][12]/P0001 ,
		_w38201_,
		_w38280_
	);
	LUT2 #(
		.INIT('h8)
	) name34234 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w38201_,
		_w38281_
	);
	LUT2 #(
		.INIT('h1)
	) name34235 (
		_w38280_,
		_w38281_,
		_w38282_
	);
	LUT2 #(
		.INIT('h2)
	) name34236 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][11]/P0001 ,
		_w38201_,
		_w38283_
	);
	LUT2 #(
		.INIT('h8)
	) name34237 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w38201_,
		_w38284_
	);
	LUT2 #(
		.INIT('h1)
	) name34238 (
		_w38283_,
		_w38284_,
		_w38285_
	);
	LUT2 #(
		.INIT('h2)
	) name34239 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][10]/P0001 ,
		_w38201_,
		_w38286_
	);
	LUT2 #(
		.INIT('h8)
	) name34240 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w38201_,
		_w38287_
	);
	LUT2 #(
		.INIT('h1)
	) name34241 (
		_w38286_,
		_w38287_,
		_w38288_
	);
	LUT2 #(
		.INIT('h2)
	) name34242 (
		\core_c_psq_ststk_sts7x23_STcell_reg[6][0]/P0001 ,
		_w38201_,
		_w38289_
	);
	LUT2 #(
		.INIT('h8)
	) name34243 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w38201_,
		_w38290_
	);
	LUT2 #(
		.INIT('h1)
	) name34244 (
		_w38289_,
		_w38290_,
		_w38291_
	);
	LUT2 #(
		.INIT('h2)
	) name34245 (
		_w14706_,
		_w18220_,
		_w38292_
	);
	LUT2 #(
		.INIT('h2)
	) name34246 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][9]/P0001 ,
		_w38292_,
		_w38293_
	);
	LUT2 #(
		.INIT('h8)
	) name34247 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w38292_,
		_w38294_
	);
	LUT2 #(
		.INIT('h1)
	) name34248 (
		_w38293_,
		_w38294_,
		_w38295_
	);
	LUT2 #(
		.INIT('h2)
	) name34249 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][8]/P0001 ,
		_w38292_,
		_w38296_
	);
	LUT2 #(
		.INIT('h8)
	) name34250 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w38292_,
		_w38297_
	);
	LUT2 #(
		.INIT('h1)
	) name34251 (
		_w38296_,
		_w38297_,
		_w38298_
	);
	LUT2 #(
		.INIT('h2)
	) name34252 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][7]/P0001 ,
		_w38292_,
		_w38299_
	);
	LUT2 #(
		.INIT('h8)
	) name34253 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w38292_,
		_w38300_
	);
	LUT2 #(
		.INIT('h1)
	) name34254 (
		_w38299_,
		_w38300_,
		_w38301_
	);
	LUT2 #(
		.INIT('h2)
	) name34255 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][6]/P0001 ,
		_w38292_,
		_w38302_
	);
	LUT2 #(
		.INIT('h4)
	) name34256 (
		_w4174_,
		_w38292_,
		_w38303_
	);
	LUT2 #(
		.INIT('h1)
	) name34257 (
		_w38302_,
		_w38303_,
		_w38304_
	);
	LUT2 #(
		.INIT('h2)
	) name34258 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][5]/P0001 ,
		_w38292_,
		_w38305_
	);
	LUT2 #(
		.INIT('h8)
	) name34259 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w38292_,
		_w38306_
	);
	LUT2 #(
		.INIT('h1)
	) name34260 (
		_w38305_,
		_w38306_,
		_w38307_
	);
	LUT2 #(
		.INIT('h2)
	) name34261 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][4]/P0001 ,
		_w38292_,
		_w38308_
	);
	LUT2 #(
		.INIT('h8)
	) name34262 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w38292_,
		_w38309_
	);
	LUT2 #(
		.INIT('h1)
	) name34263 (
		_w38308_,
		_w38309_,
		_w38310_
	);
	LUT2 #(
		.INIT('h2)
	) name34264 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][3]/P0001 ,
		_w38292_,
		_w38311_
	);
	LUT2 #(
		.INIT('h8)
	) name34265 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w38292_,
		_w38312_
	);
	LUT2 #(
		.INIT('h1)
	) name34266 (
		_w38311_,
		_w38312_,
		_w38313_
	);
	LUT2 #(
		.INIT('h2)
	) name34267 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][2]/P0001 ,
		_w38292_,
		_w38314_
	);
	LUT2 #(
		.INIT('h8)
	) name34268 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w38292_,
		_w38315_
	);
	LUT2 #(
		.INIT('h1)
	) name34269 (
		_w38314_,
		_w38315_,
		_w38316_
	);
	LUT2 #(
		.INIT('h2)
	) name34270 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][24]/P0001 ,
		_w38292_,
		_w38317_
	);
	LUT2 #(
		.INIT('h8)
	) name34271 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w38292_,
		_w38318_
	);
	LUT2 #(
		.INIT('h1)
	) name34272 (
		_w38317_,
		_w38318_,
		_w38319_
	);
	LUT2 #(
		.INIT('h2)
	) name34273 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][23]/P0001 ,
		_w38292_,
		_w38320_
	);
	LUT2 #(
		.INIT('h8)
	) name34274 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w38292_,
		_w38321_
	);
	LUT2 #(
		.INIT('h1)
	) name34275 (
		_w38320_,
		_w38321_,
		_w38322_
	);
	LUT2 #(
		.INIT('h2)
	) name34276 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][22]/P0001 ,
		_w38292_,
		_w38323_
	);
	LUT2 #(
		.INIT('h8)
	) name34277 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w38292_,
		_w38324_
	);
	LUT2 #(
		.INIT('h1)
	) name34278 (
		_w38323_,
		_w38324_,
		_w38325_
	);
	LUT2 #(
		.INIT('h2)
	) name34279 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][21]/P0001 ,
		_w38292_,
		_w38326_
	);
	LUT2 #(
		.INIT('h8)
	) name34280 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w38292_,
		_w38327_
	);
	LUT2 #(
		.INIT('h1)
	) name34281 (
		_w38326_,
		_w38327_,
		_w38328_
	);
	LUT2 #(
		.INIT('h2)
	) name34282 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][20]/P0001 ,
		_w38292_,
		_w38329_
	);
	LUT2 #(
		.INIT('h8)
	) name34283 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w38292_,
		_w38330_
	);
	LUT2 #(
		.INIT('h1)
	) name34284 (
		_w38329_,
		_w38330_,
		_w38331_
	);
	LUT2 #(
		.INIT('h2)
	) name34285 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][1]/P0001 ,
		_w38292_,
		_w38332_
	);
	LUT2 #(
		.INIT('h8)
	) name34286 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w38292_,
		_w38333_
	);
	LUT2 #(
		.INIT('h1)
	) name34287 (
		_w38332_,
		_w38333_,
		_w38334_
	);
	LUT2 #(
		.INIT('h2)
	) name34288 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][19]/P0001 ,
		_w38292_,
		_w38335_
	);
	LUT2 #(
		.INIT('h8)
	) name34289 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w38292_,
		_w38336_
	);
	LUT2 #(
		.INIT('h1)
	) name34290 (
		_w38335_,
		_w38336_,
		_w38337_
	);
	LUT2 #(
		.INIT('h2)
	) name34291 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][18]/P0001 ,
		_w38292_,
		_w38338_
	);
	LUT2 #(
		.INIT('h8)
	) name34292 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w38292_,
		_w38339_
	);
	LUT2 #(
		.INIT('h1)
	) name34293 (
		_w38338_,
		_w38339_,
		_w38340_
	);
	LUT2 #(
		.INIT('h2)
	) name34294 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][17]/P0001 ,
		_w38292_,
		_w38341_
	);
	LUT2 #(
		.INIT('h8)
	) name34295 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w38292_,
		_w38342_
	);
	LUT2 #(
		.INIT('h1)
	) name34296 (
		_w38341_,
		_w38342_,
		_w38343_
	);
	LUT2 #(
		.INIT('h2)
	) name34297 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][16]/P0001 ,
		_w38292_,
		_w38344_
	);
	LUT2 #(
		.INIT('h8)
	) name34298 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w38292_,
		_w38345_
	);
	LUT2 #(
		.INIT('h1)
	) name34299 (
		_w38344_,
		_w38345_,
		_w38346_
	);
	LUT2 #(
		.INIT('h2)
	) name34300 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][15]/P0001 ,
		_w38292_,
		_w38347_
	);
	LUT2 #(
		.INIT('h8)
	) name34301 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w38292_,
		_w38348_
	);
	LUT2 #(
		.INIT('h1)
	) name34302 (
		_w38347_,
		_w38348_,
		_w38349_
	);
	LUT2 #(
		.INIT('h2)
	) name34303 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][14]/P0001 ,
		_w38292_,
		_w38350_
	);
	LUT2 #(
		.INIT('h8)
	) name34304 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w38292_,
		_w38351_
	);
	LUT2 #(
		.INIT('h1)
	) name34305 (
		_w38350_,
		_w38351_,
		_w38352_
	);
	LUT2 #(
		.INIT('h2)
	) name34306 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][13]/P0001 ,
		_w38292_,
		_w38353_
	);
	LUT2 #(
		.INIT('h8)
	) name34307 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w38292_,
		_w38354_
	);
	LUT2 #(
		.INIT('h1)
	) name34308 (
		_w38353_,
		_w38354_,
		_w38355_
	);
	LUT2 #(
		.INIT('h2)
	) name34309 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][12]/P0001 ,
		_w38292_,
		_w38356_
	);
	LUT2 #(
		.INIT('h8)
	) name34310 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w38292_,
		_w38357_
	);
	LUT2 #(
		.INIT('h1)
	) name34311 (
		_w38356_,
		_w38357_,
		_w38358_
	);
	LUT2 #(
		.INIT('h2)
	) name34312 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][11]/P0001 ,
		_w38292_,
		_w38359_
	);
	LUT2 #(
		.INIT('h8)
	) name34313 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w38292_,
		_w38360_
	);
	LUT2 #(
		.INIT('h1)
	) name34314 (
		_w38359_,
		_w38360_,
		_w38361_
	);
	LUT2 #(
		.INIT('h2)
	) name34315 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][10]/P0001 ,
		_w38292_,
		_w38362_
	);
	LUT2 #(
		.INIT('h8)
	) name34316 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w38292_,
		_w38363_
	);
	LUT2 #(
		.INIT('h1)
	) name34317 (
		_w38362_,
		_w38363_,
		_w38364_
	);
	LUT2 #(
		.INIT('h2)
	) name34318 (
		\core_c_psq_ststk_sts7x23_STcell_reg[5][0]/P0001 ,
		_w38292_,
		_w38365_
	);
	LUT2 #(
		.INIT('h8)
	) name34319 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w38292_,
		_w38366_
	);
	LUT2 #(
		.INIT('h1)
	) name34320 (
		_w38365_,
		_w38366_,
		_w38367_
	);
	LUT2 #(
		.INIT('h4)
	) name34321 (
		\core_c_psq_ststk_ptr_reg[2]/NET0131 ,
		_w18679_,
		_w38368_
	);
	LUT2 #(
		.INIT('h2)
	) name34322 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][9]/P0001 ,
		_w38368_,
		_w38369_
	);
	LUT2 #(
		.INIT('h8)
	) name34323 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w38368_,
		_w38370_
	);
	LUT2 #(
		.INIT('h1)
	) name34324 (
		_w38369_,
		_w38370_,
		_w38371_
	);
	LUT2 #(
		.INIT('h2)
	) name34325 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][8]/P0001 ,
		_w38368_,
		_w38372_
	);
	LUT2 #(
		.INIT('h8)
	) name34326 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w38368_,
		_w38373_
	);
	LUT2 #(
		.INIT('h1)
	) name34327 (
		_w38372_,
		_w38373_,
		_w38374_
	);
	LUT2 #(
		.INIT('h2)
	) name34328 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][7]/P0001 ,
		_w38368_,
		_w38375_
	);
	LUT2 #(
		.INIT('h8)
	) name34329 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w38368_,
		_w38376_
	);
	LUT2 #(
		.INIT('h1)
	) name34330 (
		_w38375_,
		_w38376_,
		_w38377_
	);
	LUT2 #(
		.INIT('h2)
	) name34331 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][6]/P0001 ,
		_w38368_,
		_w38378_
	);
	LUT2 #(
		.INIT('h4)
	) name34332 (
		_w4174_,
		_w38368_,
		_w38379_
	);
	LUT2 #(
		.INIT('h1)
	) name34333 (
		_w38378_,
		_w38379_,
		_w38380_
	);
	LUT2 #(
		.INIT('h2)
	) name34334 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][5]/P0001 ,
		_w38368_,
		_w38381_
	);
	LUT2 #(
		.INIT('h8)
	) name34335 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w38368_,
		_w38382_
	);
	LUT2 #(
		.INIT('h1)
	) name34336 (
		_w38381_,
		_w38382_,
		_w38383_
	);
	LUT2 #(
		.INIT('h2)
	) name34337 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][4]/P0001 ,
		_w38368_,
		_w38384_
	);
	LUT2 #(
		.INIT('h8)
	) name34338 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w38368_,
		_w38385_
	);
	LUT2 #(
		.INIT('h1)
	) name34339 (
		_w38384_,
		_w38385_,
		_w38386_
	);
	LUT2 #(
		.INIT('h2)
	) name34340 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][3]/P0001 ,
		_w38368_,
		_w38387_
	);
	LUT2 #(
		.INIT('h8)
	) name34341 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w38368_,
		_w38388_
	);
	LUT2 #(
		.INIT('h1)
	) name34342 (
		_w38387_,
		_w38388_,
		_w38389_
	);
	LUT2 #(
		.INIT('h2)
	) name34343 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][2]/P0001 ,
		_w38368_,
		_w38390_
	);
	LUT2 #(
		.INIT('h8)
	) name34344 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w38368_,
		_w38391_
	);
	LUT2 #(
		.INIT('h1)
	) name34345 (
		_w38390_,
		_w38391_,
		_w38392_
	);
	LUT2 #(
		.INIT('h2)
	) name34346 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][24]/P0001 ,
		_w38368_,
		_w38393_
	);
	LUT2 #(
		.INIT('h8)
	) name34347 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w38368_,
		_w38394_
	);
	LUT2 #(
		.INIT('h1)
	) name34348 (
		_w38393_,
		_w38394_,
		_w38395_
	);
	LUT2 #(
		.INIT('h2)
	) name34349 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][23]/P0001 ,
		_w38368_,
		_w38396_
	);
	LUT2 #(
		.INIT('h8)
	) name34350 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w38368_,
		_w38397_
	);
	LUT2 #(
		.INIT('h1)
	) name34351 (
		_w38396_,
		_w38397_,
		_w38398_
	);
	LUT2 #(
		.INIT('h2)
	) name34352 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][22]/P0001 ,
		_w38368_,
		_w38399_
	);
	LUT2 #(
		.INIT('h8)
	) name34353 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w38368_,
		_w38400_
	);
	LUT2 #(
		.INIT('h1)
	) name34354 (
		_w38399_,
		_w38400_,
		_w38401_
	);
	LUT2 #(
		.INIT('h2)
	) name34355 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][21]/P0001 ,
		_w38368_,
		_w38402_
	);
	LUT2 #(
		.INIT('h8)
	) name34356 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w38368_,
		_w38403_
	);
	LUT2 #(
		.INIT('h1)
	) name34357 (
		_w38402_,
		_w38403_,
		_w38404_
	);
	LUT2 #(
		.INIT('h2)
	) name34358 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][20]/P0001 ,
		_w38368_,
		_w38405_
	);
	LUT2 #(
		.INIT('h8)
	) name34359 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w38368_,
		_w38406_
	);
	LUT2 #(
		.INIT('h1)
	) name34360 (
		_w38405_,
		_w38406_,
		_w38407_
	);
	LUT2 #(
		.INIT('h2)
	) name34361 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][1]/P0001 ,
		_w38368_,
		_w38408_
	);
	LUT2 #(
		.INIT('h8)
	) name34362 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w38368_,
		_w38409_
	);
	LUT2 #(
		.INIT('h1)
	) name34363 (
		_w38408_,
		_w38409_,
		_w38410_
	);
	LUT2 #(
		.INIT('h2)
	) name34364 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][19]/P0001 ,
		_w38368_,
		_w38411_
	);
	LUT2 #(
		.INIT('h8)
	) name34365 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w38368_,
		_w38412_
	);
	LUT2 #(
		.INIT('h1)
	) name34366 (
		_w38411_,
		_w38412_,
		_w38413_
	);
	LUT2 #(
		.INIT('h2)
	) name34367 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][18]/P0001 ,
		_w38368_,
		_w38414_
	);
	LUT2 #(
		.INIT('h8)
	) name34368 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w38368_,
		_w38415_
	);
	LUT2 #(
		.INIT('h1)
	) name34369 (
		_w38414_,
		_w38415_,
		_w38416_
	);
	LUT2 #(
		.INIT('h2)
	) name34370 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][17]/P0001 ,
		_w38368_,
		_w38417_
	);
	LUT2 #(
		.INIT('h8)
	) name34371 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w38368_,
		_w38418_
	);
	LUT2 #(
		.INIT('h1)
	) name34372 (
		_w38417_,
		_w38418_,
		_w38419_
	);
	LUT2 #(
		.INIT('h2)
	) name34373 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][16]/P0001 ,
		_w38368_,
		_w38420_
	);
	LUT2 #(
		.INIT('h8)
	) name34374 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w38368_,
		_w38421_
	);
	LUT2 #(
		.INIT('h1)
	) name34375 (
		_w38420_,
		_w38421_,
		_w38422_
	);
	LUT2 #(
		.INIT('h2)
	) name34376 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][15]/P0001 ,
		_w38368_,
		_w38423_
	);
	LUT2 #(
		.INIT('h8)
	) name34377 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w38368_,
		_w38424_
	);
	LUT2 #(
		.INIT('h1)
	) name34378 (
		_w38423_,
		_w38424_,
		_w38425_
	);
	LUT2 #(
		.INIT('h2)
	) name34379 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][14]/P0001 ,
		_w38368_,
		_w38426_
	);
	LUT2 #(
		.INIT('h8)
	) name34380 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w38368_,
		_w38427_
	);
	LUT2 #(
		.INIT('h1)
	) name34381 (
		_w38426_,
		_w38427_,
		_w38428_
	);
	LUT2 #(
		.INIT('h2)
	) name34382 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][13]/P0001 ,
		_w38368_,
		_w38429_
	);
	LUT2 #(
		.INIT('h8)
	) name34383 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w38368_,
		_w38430_
	);
	LUT2 #(
		.INIT('h1)
	) name34384 (
		_w38429_,
		_w38430_,
		_w38431_
	);
	LUT2 #(
		.INIT('h2)
	) name34385 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][12]/P0001 ,
		_w38368_,
		_w38432_
	);
	LUT2 #(
		.INIT('h8)
	) name34386 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w38368_,
		_w38433_
	);
	LUT2 #(
		.INIT('h1)
	) name34387 (
		_w38432_,
		_w38433_,
		_w38434_
	);
	LUT2 #(
		.INIT('h2)
	) name34388 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][11]/P0001 ,
		_w38368_,
		_w38435_
	);
	LUT2 #(
		.INIT('h8)
	) name34389 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w38368_,
		_w38436_
	);
	LUT2 #(
		.INIT('h1)
	) name34390 (
		_w38435_,
		_w38436_,
		_w38437_
	);
	LUT2 #(
		.INIT('h2)
	) name34391 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][10]/P0001 ,
		_w38368_,
		_w38438_
	);
	LUT2 #(
		.INIT('h8)
	) name34392 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w38368_,
		_w38439_
	);
	LUT2 #(
		.INIT('h1)
	) name34393 (
		_w38438_,
		_w38439_,
		_w38440_
	);
	LUT2 #(
		.INIT('h2)
	) name34394 (
		\core_c_psq_ststk_sts7x23_STcell_reg[4][0]/P0001 ,
		_w38368_,
		_w38441_
	);
	LUT2 #(
		.INIT('h8)
	) name34395 (
		\core_eu_ec_cun_AZ_reg/P0001 ,
		_w38368_,
		_w38442_
	);
	LUT2 #(
		.INIT('h1)
	) name34396 (
		_w38441_,
		_w38442_,
		_w38443_
	);
	LUT2 #(
		.INIT('h2)
	) name34397 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][9]/P0001 ,
		_w18221_,
		_w38444_
	);
	LUT2 #(
		.INIT('h8)
	) name34398 (
		\core_c_psq_MSTAT_reg_DO_reg[1]/NET0131 ,
		_w18221_,
		_w38445_
	);
	LUT2 #(
		.INIT('h1)
	) name34399 (
		_w38444_,
		_w38445_,
		_w38446_
	);
	LUT2 #(
		.INIT('h2)
	) name34400 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][8]/P0001 ,
		_w18221_,
		_w38447_
	);
	LUT2 #(
		.INIT('h8)
	) name34401 (
		\core_c_psq_MSTAT_reg_DO_reg[0]/P0002 ,
		_w18221_,
		_w38448_
	);
	LUT2 #(
		.INIT('h1)
	) name34402 (
		_w38447_,
		_w38448_,
		_w38449_
	);
	LUT2 #(
		.INIT('h2)
	) name34403 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][7]/P0001 ,
		_w18221_,
		_w38450_
	);
	LUT2 #(
		.INIT('h8)
	) name34404 (
		\core_eu_ec_cun_SS_reg/P0001 ,
		_w18221_,
		_w38451_
	);
	LUT2 #(
		.INIT('h1)
	) name34405 (
		_w38450_,
		_w38451_,
		_w38452_
	);
	LUT2 #(
		.INIT('h2)
	) name34406 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][6]/P0001 ,
		_w18221_,
		_w38453_
	);
	LUT2 #(
		.INIT('h4)
	) name34407 (
		_w4174_,
		_w18221_,
		_w38454_
	);
	LUT2 #(
		.INIT('h1)
	) name34408 (
		_w38453_,
		_w38454_,
		_w38455_
	);
	LUT2 #(
		.INIT('h2)
	) name34409 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][5]/P0001 ,
		_w18221_,
		_w38456_
	);
	LUT2 #(
		.INIT('h8)
	) name34410 (
		\core_eu_ec_cun_AQ_reg/P0001 ,
		_w18221_,
		_w38457_
	);
	LUT2 #(
		.INIT('h1)
	) name34411 (
		_w38456_,
		_w38457_,
		_w38458_
	);
	LUT2 #(
		.INIT('h2)
	) name34412 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][4]/P0001 ,
		_w18221_,
		_w38459_
	);
	LUT2 #(
		.INIT('h8)
	) name34413 (
		\core_eu_ec_cun_AS_reg/P0001 ,
		_w18221_,
		_w38460_
	);
	LUT2 #(
		.INIT('h1)
	) name34414 (
		_w38459_,
		_w38460_,
		_w38461_
	);
	LUT2 #(
		.INIT('h2)
	) name34415 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][3]/P0001 ,
		_w18221_,
		_w38462_
	);
	LUT2 #(
		.INIT('h8)
	) name34416 (
		\core_eu_ec_cun_AC_reg/P0001 ,
		_w18221_,
		_w38463_
	);
	LUT2 #(
		.INIT('h1)
	) name34417 (
		_w38462_,
		_w38463_,
		_w38464_
	);
	LUT2 #(
		.INIT('h2)
	) name34418 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][2]/P0001 ,
		_w18221_,
		_w38465_
	);
	LUT2 #(
		.INIT('h8)
	) name34419 (
		\core_eu_ec_cun_AV_reg/P0001 ,
		_w18221_,
		_w38466_
	);
	LUT2 #(
		.INIT('h1)
	) name34420 (
		_w38465_,
		_w38466_,
		_w38467_
	);
	LUT2 #(
		.INIT('h2)
	) name34421 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][24]/P0001 ,
		_w18221_,
		_w38468_
	);
	LUT2 #(
		.INIT('h8)
	) name34422 (
		\core_c_psq_IMASK_reg[9]/NET0131 ,
		_w18221_,
		_w38469_
	);
	LUT2 #(
		.INIT('h1)
	) name34423 (
		_w38468_,
		_w38469_,
		_w38470_
	);
	LUT2 #(
		.INIT('h2)
	) name34424 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][23]/P0001 ,
		_w18221_,
		_w38471_
	);
	LUT2 #(
		.INIT('h8)
	) name34425 (
		\core_c_psq_IMASK_reg[8]/NET0131 ,
		_w18221_,
		_w38472_
	);
	LUT2 #(
		.INIT('h1)
	) name34426 (
		_w38471_,
		_w38472_,
		_w38473_
	);
	LUT2 #(
		.INIT('h2)
	) name34427 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][22]/P0001 ,
		_w18221_,
		_w38474_
	);
	LUT2 #(
		.INIT('h8)
	) name34428 (
		\core_c_psq_IMASK_reg[7]/NET0131 ,
		_w18221_,
		_w38475_
	);
	LUT2 #(
		.INIT('h1)
	) name34429 (
		_w38474_,
		_w38475_,
		_w38476_
	);
	LUT2 #(
		.INIT('h2)
	) name34430 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][21]/P0001 ,
		_w18221_,
		_w38477_
	);
	LUT2 #(
		.INIT('h8)
	) name34431 (
		\core_c_psq_IMASK_reg[6]/NET0131 ,
		_w18221_,
		_w38478_
	);
	LUT2 #(
		.INIT('h1)
	) name34432 (
		_w38477_,
		_w38478_,
		_w38479_
	);
	LUT2 #(
		.INIT('h2)
	) name34433 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][20]/P0001 ,
		_w18221_,
		_w38480_
	);
	LUT2 #(
		.INIT('h8)
	) name34434 (
		\core_c_psq_IMASK_reg[5]/NET0131 ,
		_w18221_,
		_w38481_
	);
	LUT2 #(
		.INIT('h1)
	) name34435 (
		_w38480_,
		_w38481_,
		_w38482_
	);
	LUT2 #(
		.INIT('h2)
	) name34436 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][1]/P0001 ,
		_w18221_,
		_w38483_
	);
	LUT2 #(
		.INIT('h8)
	) name34437 (
		\core_eu_ec_cun_AN_reg/P0001 ,
		_w18221_,
		_w38484_
	);
	LUT2 #(
		.INIT('h1)
	) name34438 (
		_w38483_,
		_w38484_,
		_w38485_
	);
	LUT2 #(
		.INIT('h2)
	) name34439 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][19]/P0001 ,
		_w18221_,
		_w38486_
	);
	LUT2 #(
		.INIT('h8)
	) name34440 (
		\core_c_psq_IMASK_reg[4]/NET0131 ,
		_w18221_,
		_w38487_
	);
	LUT2 #(
		.INIT('h1)
	) name34441 (
		_w38486_,
		_w38487_,
		_w38488_
	);
	LUT2 #(
		.INIT('h4)
	) name34442 (
		_w18213_,
		_w18717_,
		_w38489_
	);
	LUT2 #(
		.INIT('h1)
	) name34443 (
		\core_eu_es_sht_es_reg_sr1swe_DO_reg[13]/P0001 ,
		_w18717_,
		_w38490_
	);
	LUT2 #(
		.INIT('h1)
	) name34444 (
		_w38489_,
		_w38490_,
		_w38491_
	);
	LUT2 #(
		.INIT('h2)
	) name34445 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][18]/P0001 ,
		_w18221_,
		_w38492_
	);
	LUT2 #(
		.INIT('h8)
	) name34446 (
		\core_c_psq_IMASK_reg[3]/NET0131 ,
		_w18221_,
		_w38493_
	);
	LUT2 #(
		.INIT('h1)
	) name34447 (
		_w38492_,
		_w38493_,
		_w38494_
	);
	LUT2 #(
		.INIT('h2)
	) name34448 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][17]/P0001 ,
		_w18221_,
		_w38495_
	);
	LUT2 #(
		.INIT('h8)
	) name34449 (
		\core_c_psq_IMASK_reg[2]/NET0131 ,
		_w18221_,
		_w38496_
	);
	LUT2 #(
		.INIT('h1)
	) name34450 (
		_w38495_,
		_w38496_,
		_w38497_
	);
	LUT2 #(
		.INIT('h8)
	) name34451 (
		\sport0_regs_SCTLreg_DO_reg[13]/NET0131 ,
		_w18233_,
		_w38498_
	);
	LUT2 #(
		.INIT('h8)
	) name34452 (
		_w7340_,
		_w18237_,
		_w38499_
	);
	LUT2 #(
		.INIT('h1)
	) name34453 (
		_w38498_,
		_w38499_,
		_w38500_
	);
	LUT2 #(
		.INIT('h2)
	) name34454 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][16]/P0001 ,
		_w18221_,
		_w38501_
	);
	LUT2 #(
		.INIT('h8)
	) name34455 (
		\core_c_psq_IMASK_reg[1]/NET0131 ,
		_w18221_,
		_w38502_
	);
	LUT2 #(
		.INIT('h1)
	) name34456 (
		_w38501_,
		_w38502_,
		_w38503_
	);
	LUT2 #(
		.INIT('h2)
	) name34457 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][15]/P0001 ,
		_w18221_,
		_w38504_
	);
	LUT2 #(
		.INIT('h8)
	) name34458 (
		\core_c_psq_IMASK_reg[0]/NET0131 ,
		_w18221_,
		_w38505_
	);
	LUT2 #(
		.INIT('h1)
	) name34459 (
		_w38504_,
		_w38505_,
		_w38506_
	);
	LUT2 #(
		.INIT('h2)
	) name34460 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][14]/P0001 ,
		_w18221_,
		_w38507_
	);
	LUT2 #(
		.INIT('h8)
	) name34461 (
		\core_c_psq_MSTAT_reg_DO_reg[6]/NET0131 ,
		_w18221_,
		_w38508_
	);
	LUT2 #(
		.INIT('h1)
	) name34462 (
		_w38507_,
		_w38508_,
		_w38509_
	);
	LUT2 #(
		.INIT('h2)
	) name34463 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][13]/P0001 ,
		_w18221_,
		_w38510_
	);
	LUT2 #(
		.INIT('h8)
	) name34464 (
		\core_c_psq_MSTAT_reg_DO_reg[5]/NET0131 ,
		_w18221_,
		_w38511_
	);
	LUT2 #(
		.INIT('h1)
	) name34465 (
		_w38510_,
		_w38511_,
		_w38512_
	);
	LUT2 #(
		.INIT('h2)
	) name34466 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][12]/P0001 ,
		_w18221_,
		_w38513_
	);
	LUT2 #(
		.INIT('h8)
	) name34467 (
		\core_c_psq_MSTAT_reg_DO_reg[4]/NET0131 ,
		_w18221_,
		_w38514_
	);
	LUT2 #(
		.INIT('h1)
	) name34468 (
		_w38513_,
		_w38514_,
		_w38515_
	);
	LUT2 #(
		.INIT('h2)
	) name34469 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][11]/P0001 ,
		_w18221_,
		_w38516_
	);
	LUT2 #(
		.INIT('h8)
	) name34470 (
		\core_c_psq_MSTAT_reg_DO_reg[3]/NET0131 ,
		_w18221_,
		_w38517_
	);
	LUT2 #(
		.INIT('h1)
	) name34471 (
		_w38516_,
		_w38517_,
		_w38518_
	);
	LUT2 #(
		.INIT('h2)
	) name34472 (
		\core_c_psq_ststk_sts7x23_STcell_reg[3][10]/P0001 ,
		_w18221_,
		_w38519_
	);
	LUT2 #(
		.INIT('h8)
	) name34473 (
		\core_c_psq_MSTAT_reg_DO_reg[2]/NET0131 ,
		_w18221_,
		_w38520_
	);
	LUT2 #(
		.INIT('h1)
	) name34474 (
		_w38519_,
		_w38520_,
		_w38521_
	);
	LUT2 #(
		.INIT('h1)
	) name34475 (
		_w26090_,
		_w34434_,
		_w38522_
	);
	LUT2 #(
		.INIT('h8)
	) name34476 (
		\T_TMODE[1]_pad ,
		\core_c_dec_PPclr_reg/P0001 ,
		_w38523_
	);
	LUT2 #(
		.INIT('h1)
	) name34477 (
		_w32093_,
		_w38523_,
		_w38524_
	);
	LUT2 #(
		.INIT('h2)
	) name34478 (
		\T_PIOin[0]_pad ,
		_w25656_,
		_w38525_
	);
	LUT2 #(
		.INIT('h8)
	) name34479 (
		\pio_PIO_IN_P_reg[0]/P0001 ,
		_w25656_,
		_w38526_
	);
	LUT2 #(
		.INIT('h1)
	) name34480 (
		_w38525_,
		_w38526_,
		_w38527_
	);
	LUT2 #(
		.INIT('h2)
	) name34481 (
		\T_PIOin[10]_pad ,
		_w25661_,
		_w38528_
	);
	LUT2 #(
		.INIT('h8)
	) name34482 (
		\pio_PIO_IN_P_reg[10]/P0001 ,
		_w25661_,
		_w38529_
	);
	LUT2 #(
		.INIT('h1)
	) name34483 (
		_w38528_,
		_w38529_,
		_w38530_
	);
	LUT2 #(
		.INIT('h2)
	) name34484 (
		\T_PIOin[11]_pad ,
		_w25661_,
		_w38531_
	);
	LUT2 #(
		.INIT('h8)
	) name34485 (
		\pio_PIO_IN_P_reg[11]/P0001 ,
		_w25661_,
		_w38532_
	);
	LUT2 #(
		.INIT('h1)
	) name34486 (
		_w38531_,
		_w38532_,
		_w38533_
	);
	LUT2 #(
		.INIT('h2)
	) name34487 (
		\T_PIOin[1]_pad ,
		_w25656_,
		_w38534_
	);
	LUT2 #(
		.INIT('h8)
	) name34488 (
		\pio_PIO_IN_P_reg[1]/P0001 ,
		_w25656_,
		_w38535_
	);
	LUT2 #(
		.INIT('h1)
	) name34489 (
		_w38534_,
		_w38535_,
		_w38536_
	);
	LUT2 #(
		.INIT('h2)
	) name34490 (
		\T_PIOin[2]_pad ,
		_w25666_,
		_w38537_
	);
	LUT2 #(
		.INIT('h8)
	) name34491 (
		\pio_PIO_IN_P_reg[2]/P0001 ,
		_w25666_,
		_w38538_
	);
	LUT2 #(
		.INIT('h1)
	) name34492 (
		_w38537_,
		_w38538_,
		_w38539_
	);
	LUT2 #(
		.INIT('h2)
	) name34493 (
		\T_PIOin[3]_pad ,
		_w25666_,
		_w38540_
	);
	LUT2 #(
		.INIT('h8)
	) name34494 (
		\pio_PIO_IN_P_reg[3]/P0001 ,
		_w25666_,
		_w38541_
	);
	LUT2 #(
		.INIT('h1)
	) name34495 (
		_w38540_,
		_w38541_,
		_w38542_
	);
	LUT2 #(
		.INIT('h2)
	) name34496 (
		\T_PIOin[4]_pad ,
		_w25679_,
		_w38543_
	);
	LUT2 #(
		.INIT('h8)
	) name34497 (
		\pio_PIO_IN_P_reg[4]/P0001 ,
		_w25679_,
		_w38544_
	);
	LUT2 #(
		.INIT('h1)
	) name34498 (
		_w38543_,
		_w38544_,
		_w38545_
	);
	LUT2 #(
		.INIT('h2)
	) name34499 (
		\T_PIOin[5]_pad ,
		_w25679_,
		_w38546_
	);
	LUT2 #(
		.INIT('h8)
	) name34500 (
		\pio_PIO_IN_P_reg[5]/P0001 ,
		_w25679_,
		_w38547_
	);
	LUT2 #(
		.INIT('h1)
	) name34501 (
		_w38546_,
		_w38547_,
		_w38548_
	);
	LUT2 #(
		.INIT('h2)
	) name34502 (
		\T_PIOin[6]_pad ,
		_w25671_,
		_w38549_
	);
	LUT2 #(
		.INIT('h8)
	) name34503 (
		\pio_PIO_IN_P_reg[6]/P0001 ,
		_w25671_,
		_w38550_
	);
	LUT2 #(
		.INIT('h1)
	) name34504 (
		_w38549_,
		_w38550_,
		_w38551_
	);
	LUT2 #(
		.INIT('h2)
	) name34505 (
		\T_PIOin[7]_pad ,
		_w25671_,
		_w38552_
	);
	LUT2 #(
		.INIT('h8)
	) name34506 (
		\pio_PIO_IN_P_reg[7]/P0001 ,
		_w25671_,
		_w38553_
	);
	LUT2 #(
		.INIT('h1)
	) name34507 (
		_w38552_,
		_w38553_,
		_w38554_
	);
	LUT2 #(
		.INIT('h2)
	) name34508 (
		\T_PIOin[8]_pad ,
		_w25651_,
		_w38555_
	);
	LUT2 #(
		.INIT('h8)
	) name34509 (
		\pio_PIO_IN_P_reg[8]/P0001 ,
		_w25651_,
		_w38556_
	);
	LUT2 #(
		.INIT('h1)
	) name34510 (
		_w38555_,
		_w38556_,
		_w38557_
	);
	LUT2 #(
		.INIT('h2)
	) name34511 (
		\T_PIOin[9]_pad ,
		_w25651_,
		_w38558_
	);
	LUT2 #(
		.INIT('h8)
	) name34512 (
		\pio_PIO_IN_P_reg[9]/P0001 ,
		_w25651_,
		_w38559_
	);
	LUT2 #(
		.INIT('h1)
	) name34513 (
		_w38558_,
		_w38559_,
		_w38560_
	);
	LUT2 #(
		.INIT('h2)
	) name34514 (
		\pio_PIO_RES_reg[0]/NET0131 ,
		_w25656_,
		_w38561_
	);
	LUT2 #(
		.INIT('h8)
	) name34515 (
		\pio_PIO_RES_OUT_reg[0]/P0001 ,
		_w25656_,
		_w38562_
	);
	LUT2 #(
		.INIT('h1)
	) name34516 (
		_w38561_,
		_w38562_,
		_w38563_
	);
	LUT2 #(
		.INIT('h2)
	) name34517 (
		\pio_PIO_RES_reg[10]/NET0131 ,
		_w25661_,
		_w38564_
	);
	LUT2 #(
		.INIT('h8)
	) name34518 (
		\pio_PIO_RES_OUT_reg[10]/P0001 ,
		_w25661_,
		_w38565_
	);
	LUT2 #(
		.INIT('h1)
	) name34519 (
		_w38564_,
		_w38565_,
		_w38566_
	);
	LUT2 #(
		.INIT('h2)
	) name34520 (
		\pio_PIO_RES_reg[2]/NET0131 ,
		_w25666_,
		_w38567_
	);
	LUT2 #(
		.INIT('h8)
	) name34521 (
		\pio_PIO_RES_OUT_reg[2]/P0001 ,
		_w25666_,
		_w38568_
	);
	LUT2 #(
		.INIT('h1)
	) name34522 (
		_w38567_,
		_w38568_,
		_w38569_
	);
	LUT2 #(
		.INIT('h2)
	) name34523 (
		\pio_PIO_RES_reg[4]/NET0131 ,
		_w25679_,
		_w38570_
	);
	LUT2 #(
		.INIT('h8)
	) name34524 (
		\pio_PIO_RES_OUT_reg[4]/P0001 ,
		_w25679_,
		_w38571_
	);
	LUT2 #(
		.INIT('h1)
	) name34525 (
		_w38570_,
		_w38571_,
		_w38572_
	);
	LUT2 #(
		.INIT('h2)
	) name34526 (
		\pio_PIO_RES_reg[6]/NET0131 ,
		_w25671_,
		_w38573_
	);
	LUT2 #(
		.INIT('h8)
	) name34527 (
		\pio_PIO_RES_OUT_reg[6]/P0001 ,
		_w25671_,
		_w38574_
	);
	LUT2 #(
		.INIT('h1)
	) name34528 (
		_w38573_,
		_w38574_,
		_w38575_
	);
	LUT2 #(
		.INIT('h2)
	) name34529 (
		\sice_GO_NXi_reg/NET0131 ,
		_w23033_,
		_w38576_
	);
	LUT2 #(
		.INIT('h8)
	) name34530 (
		\sice_SPC_reg[20]/P0001 ,
		_w23033_,
		_w38577_
	);
	LUT2 #(
		.INIT('h1)
	) name34531 (
		_w38576_,
		_w38577_,
		_w38578_
	);
	LUT2 #(
		.INIT('h4)
	) name34532 (
		_w20442_,
		_w30779_,
		_w38579_
	);
	LUT2 #(
		.INIT('h1)
	) name34533 (
		\sport0_rxctl_RXSHT_reg[0]/P0001 ,
		_w30779_,
		_w38580_
	);
	LUT2 #(
		.INIT('h1)
	) name34534 (
		_w38579_,
		_w38580_,
		_w38581_
	);
	LUT2 #(
		.INIT('h2)
	) name34535 (
		\sport0_rxctl_RXSHT_reg[1]/P0001 ,
		_w30779_,
		_w38582_
	);
	LUT2 #(
		.INIT('h1)
	) name34536 (
		_w30784_,
		_w38582_,
		_w38583_
	);
	LUT2 #(
		.INIT('h4)
	) name34537 (
		_w20420_,
		_w30755_,
		_w38584_
	);
	LUT2 #(
		.INIT('h1)
	) name34538 (
		\sport1_rxctl_RXSHT_reg[0]/P0001 ,
		_w30755_,
		_w38585_
	);
	LUT2 #(
		.INIT('h1)
	) name34539 (
		_w38584_,
		_w38585_,
		_w38586_
	);
	LUT2 #(
		.INIT('h2)
	) name34540 (
		\sport1_rxctl_RXSHT_reg[1]/P0001 ,
		_w30755_,
		_w38587_
	);
	LUT2 #(
		.INIT('h1)
	) name34541 (
		_w30760_,
		_w38587_,
		_w38588_
	);
	assign CLKO_pad = _w4047_ ;
	assign \CMAinx[0]_pad  = _w5073_ ;
	assign \CMAinx[10]_pad  = _w5120_ ;
	assign \CMAinx[11]_pad  = _w5149_ ;
	assign \CMAinx[1]_pad  = _w5176_ ;
	assign \CMAinx[2]_pad  = _w5215_ ;
	assign \CMAinx[3]_pad  = _w5252_ ;
	assign \CMAinx[4]_pad  = _w5286_ ;
	assign \CMAinx[5]_pad  = _w5318_ ;
	assign \CMAinx[6]_pad  = _w5345_ ;
	assign \CMAinx[7]_pad  = _w5372_ ;
	assign \CMAinx[8]_pad  = _w5399_ ;
	assign \CMAinx[9]_pad  = _w5426_ ;
	assign CMSn_pad = _w5613_ ;
	assign CM_cs_pad = _w5725_ ;
	assign \CM_wd[0]_pad  = _w5741_ ;
	assign \CM_wd[10]_pad  = _w5747_ ;
	assign \CM_wd[11]_pad  = _w5753_ ;
	assign \CM_wd[12]_pad  = _w5759_ ;
	assign \CM_wd[13]_pad  = _w5765_ ;
	assign \CM_wd[14]_pad  = _w5771_ ;
	assign \CM_wd[15]_pad  = _w5777_ ;
	assign \CM_wd[16]_pad  = _w5783_ ;
	assign \CM_wd[17]_pad  = _w5789_ ;
	assign \CM_wd[18]_pad  = _w5795_ ;
	assign \CM_wd[19]_pad  = _w5801_ ;
	assign \CM_wd[1]_pad  = _w5807_ ;
	assign \CM_wd[20]_pad  = _w5813_ ;
	assign \CM_wd[21]_pad  = _w5819_ ;
	assign \CM_wd[22]_pad  = _w5825_ ;
	assign \CM_wd[23]_pad  = _w5831_ ;
	assign \CM_wd[2]_pad  = _w5837_ ;
	assign \CM_wd[3]_pad  = _w5843_ ;
	assign \CM_wd[4]_pad  = _w5849_ ;
	assign \CM_wd[5]_pad  = _w5855_ ;
	assign \CM_wd[6]_pad  = _w5861_ ;
	assign \CM_wd[7]_pad  = _w5867_ ;
	assign \CM_wd[8]_pad  = _w5873_ ;
	assign \CM_wd[9]_pad  = _w5879_ ;
	assign CM_web_pad = _w5891_ ;
	assign \CMo_cs0_pad  = _w5924_ ;
	assign \CMo_cs1_pad  = _w5925_ ;
	assign \CMo_cs2_pad  = _w5927_ ;
	assign \CMo_cs3_pad  = _w5928_ ;
	assign \CMo_cs4_pad  = _w5931_ ;
	assign \CMo_cs5_pad  = _w5932_ ;
	assign \CMo_cs6_pad  = _w5934_ ;
	assign \CMo_cs7_pad  = _w5935_ ;
	assign \DMAinx[0]_pad  = _w7628_ ;
	assign \DMAinx[10]_pad  = _w8230_ ;
	assign \DMAinx[11]_pad  = _w8835_ ;
	assign \DMAinx[12]_pad  = _w9440_ ;
	assign \DMAinx[13]_pad  = _w9513_ ;
	assign \DMAinx[1]_pad  = _w9585_ ;
	assign \DMAinx[2]_pad  = _w9651_ ;
	assign \DMAinx[3]_pad  = _w9717_ ;
	assign \DMAinx[4]_pad  = _w10308_ ;
	assign \DMAinx[5]_pad  = _w10916_ ;
	assign \DMAinx[6]_pad  = _w11530_ ;
	assign \DMAinx[7]_pad  = _w11596_ ;
	assign \DMAinx[8]_pad  = _w11660_ ;
	assign \DMAinx[9]_pad  = _w11726_ ;
	assign DMSn_pad = _w5602_ ;
	assign DM_cs_pad = _w11767_ ;
	assign \DM_wd[0]_pad  = _w11780_ ;
	assign \DM_wd[10]_pad  = _w11789_ ;
	assign \DM_wd[11]_pad  = _w11798_ ;
	assign \DM_wd[12]_pad  = _w11807_ ;
	assign \DM_wd[13]_pad  = _w11816_ ;
	assign \DM_wd[14]_pad  = _w11962_ ;
	assign \DM_wd[15]_pad  = _w12104_ ;
	assign \DM_wd[1]_pad  = _w12113_ ;
	assign \DM_wd[2]_pad  = _w12122_ ;
	assign \DM_wd[3]_pad  = _w12131_ ;
	assign \DM_wd[4]_pad  = _w12140_ ;
	assign \DM_wd[5]_pad  = _w12149_ ;
	assign \DM_wd[6]_pad  = _w12158_ ;
	assign \DM_wd[7]_pad  = _w12167_ ;
	assign \DM_wd[8]_pad  = _w12176_ ;
	assign \DM_wd[9]_pad  = _w12185_ ;
	assign \DMo_cs0_pad  = _w12214_ ;
	assign \DMo_cs1_pad  = _w12217_ ;
	assign \DMo_cs2_pad  = _w12220_ ;
	assign \DMo_cs3_pad  = _w12222_ ;
	assign \DMo_cs4_pad  = _w12226_ ;
	assign \DMo_cs5_pad  = _w12229_ ;
	assign \DMo_cs6_pad  = _w12231_ ;
	assign \DMo_cs7_pad  = _w12233_ ;
	assign \DSPCLK_cm1_pad  = _w12245_ ;
	assign \EA_do[0]_pad  = _w12260_ ;
	assign \EA_do[10]_pad  = _w12270_ ;
	assign \EA_do[12]_pad  = _w12296_ ;
	assign \EA_do[13]_pad  = _w12316_ ;
	assign \EA_do[14]_pad  = _w12336_ ;
	assign \EA_do[1]_pad  = _w12348_ ;
	assign \EA_do[2]_pad  = _w12360_ ;
	assign \EA_do[3]_pad  = _w12372_ ;
	assign \EA_do[4]_pad  = _w12384_ ;
	assign \EA_do[5]_pad  = _w12396_ ;
	assign \EA_do[6]_pad  = _w12408_ ;
	assign \EA_do[7]_pad  = _w12420_ ;
	assign \EA_do[8]_pad  = _w12430_ ;
	assign \EA_do[9]_pad  = _w12440_ ;
	assign EA_oe_pad = _w12450_ ;
	assign \ED_do[0]_pad  = _w12527_ ;
	assign \ED_do[10]_pad  = _w12561_ ;
	assign \ED_do[11]_pad  = _w12595_ ;
	assign \ED_do[12]_pad  = _w12629_ ;
	assign \ED_do[13]_pad  = _w12663_ ;
	assign \ED_do[14]_pad  = _w12720_ ;
	assign \ED_do[15]_pad  = _w12774_ ;
	assign \ED_do[1]_pad  = _w12808_ ;
	assign \ED_do[2]_pad  = _w12842_ ;
	assign \ED_do[3]_pad  = _w12876_ ;
	assign \ED_do[4]_pad  = _w12910_ ;
	assign \ED_do[5]_pad  = _w12944_ ;
	assign \ED_do[6]_pad  = _w12978_ ;
	assign \ED_do[7]_pad  = _w13012_ ;
	assign \ED_do[8]_pad  = _w13046_ ;
	assign \ED_do[9]_pad  = _w13080_ ;
	assign \ED_oe_14_8_pad  = _w13081_ ;
	assign \ED_oe_7_0_pad  = _w13082_ ;
	assign \IAD_do[0]_pad  = _w13087_ ;
	assign \IAD_do[10]_pad  = _w13089_ ;
	assign \IAD_do[11]_pad  = _w13091_ ;
	assign \IAD_do[12]_pad  = _w13092_ ;
	assign \IAD_do[13]_pad  = _w13094_ ;
	assign \IAD_do[14]_pad  = _w13095_ ;
	assign \IAD_do[15]_pad  = _w13097_ ;
	assign \IAD_do[1]_pad  = _w13101_ ;
	assign \IAD_do[2]_pad  = _w13105_ ;
	assign \IAD_do[3]_pad  = _w13109_ ;
	assign \IAD_do[4]_pad  = _w13113_ ;
	assign \IAD_do[5]_pad  = _w13117_ ;
	assign \IAD_do[6]_pad  = _w13121_ ;
	assign \IAD_do[7]_pad  = _w13125_ ;
	assign \IAD_do[8]_pad  = _w13126_ ;
	assign \IAD_do[9]_pad  = _w13127_ ;
	assign IAD_oe_pad = _w13128_ ;
	assign IDoe_pad = _w13129_ ;
	assign IOSn_pad = _w5610_ ;
	assign \PMAinx[0]_pad  = _w13173_ ;
	assign \PMAinx[10]_pad  = _w13192_ ;
	assign \PMAinx[11]_pad  = _w13211_ ;
	assign \PMAinx[1]_pad  = _w13230_ ;
	assign \PMAinx[2]_pad  = _w13249_ ;
	assign \PMAinx[3]_pad  = _w13268_ ;
	assign \PMAinx[4]_pad  = _w13287_ ;
	assign \PMAinx[5]_pad  = _w13306_ ;
	assign \PMAinx[6]_pad  = _w13325_ ;
	assign \PMAinx[7]_pad  = _w13344_ ;
	assign \PMAinx[8]_pad  = _w13363_ ;
	assign \PMAinx[9]_pad  = _w13382_ ;
	assign \PM_wd[0]_pad  = _w13392_ ;
	assign \PM_wd[10]_pad  = _w13399_ ;
	assign \PM_wd[11]_pad  = _w13406_ ;
	assign \PM_wd[12]_pad  = _w13413_ ;
	assign \PM_wd[13]_pad  = _w13420_ ;
	assign \PM_wd[14]_pad  = _w13427_ ;
	assign \PM_wd[15]_pad  = _w13434_ ;
	assign \PM_wd[1]_pad  = _w13441_ ;
	assign \PM_wd[2]_pad  = _w13448_ ;
	assign \PM_wd[3]_pad  = _w13455_ ;
	assign \PM_wd[4]_pad  = _w13462_ ;
	assign \PM_wd[5]_pad  = _w13469_ ;
	assign \PM_wd[6]_pad  = _w13476_ ;
	assign \PM_wd[7]_pad  = _w13483_ ;
	assign \PM_wd[8]_pad  = _w13490_ ;
	assign \PM_wd[9]_pad  = _w13497_ ;
	assign \PMo_cs0_pad  = _w13588_ ;
	assign \PMo_cs1_pad  = _w13591_ ;
	assign \PMo_cs2_pad  = _w13594_ ;
	assign \PMo_cs3_pad  = _w13596_ ;
	assign \PMo_cs4_pad  = _w13601_ ;
	assign \PMo_cs5_pad  = _w13604_ ;
	assign \PMo_cs6_pad  = _w13606_ ;
	assign \PMo_cs7_pad  = _w13608_ ;
	assign \PMo_oe0_pad  = 1'b0;
	assign \RFS0_pad  = _w13613_ ;
	assign \RFS1_pad  = _w13618_ ;
	assign \SCLK0_pad  = _w13621_ ;
	assign \SCLK1_pad  = _w13624_ ;
	assign \TD0_pad  = _w13672_ ;
	assign \TD1_pad  = _w13721_ ;
	assign \TFS0_pad  = _w13725_ ;
	assign \TFS1_pad  = _w13729_ ;
	assign \T_ISn_syn_2  = T_ISn_pad;
	assign WRn_pad = _w13732_ ;
	assign XTALoffn_pad = _w12239_ ;
	assign \_al_n0  = 1'b0;
	assign \bdma_BDMA_boot_reg/NET0131_reg_syn_3  = _w13759_ ;
	assign \bdma_BDMA_boot_reg/n0  = _w13734_ ;
	assign \bdma_BM_cyc_reg/P0000  = \bdma_BM_cyc_reg/P0001 ;
	assign \bdma_BWCOUNT_reg[5]/NET0131_reg_syn_3  = _w13774_ ;
	assign \core_c_psq_MGNT_reg/P0001  = \core_c_psq_MGNT_reg/NET0131 ;
	assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[0][5]/P0001_reg_syn_3  = _w13783_ ;
	assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[1][5]/P0001_reg_syn_3  = _w13788_ ;
	assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[2][5]/P0001_reg_syn_3  = _w13793_ ;
	assign \core_c_psq_cntstk_cnts4x14_CNTcell_reg[3][5]/P0001_reg_syn_3  = _w13798_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[12]/P0001_reg_syn_3  = _w14429_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[14]/P0001_reg_syn_3  = _w14556_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[1]/P0001_reg_syn_3  = _w14578_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[2]/P0001_reg_syn_3  = _w14592_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[4]/P0001_reg_syn_3  = _w14615_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[6]/P0001_reg_syn_3  = _w14639_ ;
	assign \core_eu_ea_alu_ea_reg_afrwe_DO_reg[9]/P0001_reg_syn_3  = _w14663_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[12]/P0001_reg_syn_3  = _w14670_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[14]/P0001_reg_syn_3  = _w14673_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[1]/P0001_reg_syn_3  = _w14676_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[2]/P0001_reg_syn_3  = _w14679_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[4]/P0001_reg_syn_3  = _w14682_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[6]/P0001_reg_syn_3  = _w14685_ ;
	assign \core_eu_ea_alu_ea_reg_afswe_DO_reg[9]/P0001_reg_syn_3  = _w14688_ ;
	assign \core_eu_ec_cun_MVi_pre_C_reg/P0001_reg_syn_3  = _w14725_ ;
	assign \core_eu_em_mac_em_reg_Sq_E_reg/P0001_reg_syn_3  = _w14731_ ;
	assign \emc_DMDreg_reg[8]/P0001_reg_syn_3  = _w14740_ ;
	assign \emc_DMDreg_reg[9]/P0001_reg_syn_3  = _w14743_ ;
	assign \emc_ECMcs_reg/P0001  = \emc_ECMcs_reg/NET0131 ;
	assign \emc_PMDreg_reg[8]/P0001_reg_syn_3  = _w14748_ ;
	assign \emc_PMDreg_reg[9]/P0001_reg_syn_3  = _w14751_ ;
	assign \g10/_0_  = _w17831_ ;
	assign \g1000/_0_  = _w18216_ ;
	assign \g10000/_0_  = _w18224_ ;
	assign \g10001/_0_  = _w18239_ ;
	assign \g10002/_0_  = _w18243_ ;
	assign \g10003/_0_  = _w18246_ ;
	assign \g10004/_0_  = _w18249_ ;
	assign \g10005/_0_  = _w18252_ ;
	assign \g10007/_0_  = _w18255_ ;
	assign \g10008/_0_  = _w18258_ ;
	assign \g10009/_0_  = _w18261_ ;
	assign \g1001/_3_  = _w18293_ ;
	assign \g10010/_0_  = _w18296_ ;
	assign \g10011/_0_  = _w18299_ ;
	assign \g10012/_0_  = _w18302_ ;
	assign \g10013/_0_  = _w18305_ ;
	assign \g10014/_0_  = _w18308_ ;
	assign \g10015/_0_  = _w18311_ ;
	assign \g10016/_0_  = _w18314_ ;
	assign \g10017/_0_  = _w18317_ ;
	assign \g10018/_0_  = _w18320_ ;
	assign \g10019/_0_  = _w18323_ ;
	assign \g1002/_3_  = _w18337_ ;
	assign \g10020/_0_  = _w18340_ ;
	assign \g10021/_0_  = _w18343_ ;
	assign \g10022/_0_  = _w18346_ ;
	assign \g10023/_0_  = _w18349_ ;
	assign \g10024/_0_  = _w18352_ ;
	assign \g10025/_0_  = _w18355_ ;
	assign \g10026/_0_  = _w18358_ ;
	assign \g10027/_0_  = _w18361_ ;
	assign \g10028/_0_  = _w18365_ ;
	assign \g10029/_0_  = _w18368_ ;
	assign \g1003/_0_  = _w18524_ ;
	assign \g10030/_0_  = _w18527_ ;
	assign \g10031/_0_  = _w18530_ ;
	assign \g10032/_0_  = _w18533_ ;
	assign \g10033/_0_  = _w18536_ ;
	assign \g10034/_0_  = _w18539_ ;
	assign \g10035/_0_  = _w18542_ ;
	assign \g10036/_0_  = _w18545_ ;
	assign \g10037/_0_  = _w18548_ ;
	assign \g10038/_0_  = _w18551_ ;
	assign \g10039/_0_  = _w18554_ ;
	assign \g10040/_0_  = _w18557_ ;
	assign \g10041/_0_  = _w18560_ ;
	assign \g10042/_0_  = _w18563_ ;
	assign \g10043/_0_  = _w18566_ ;
	assign \g10044/_0_  = _w18569_ ;
	assign \g10045/_0_  = _w18572_ ;
	assign \g10046/_0_  = _w18575_ ;
	assign \g10047/_0_  = _w18578_ ;
	assign \g10048/_0_  = _w18581_ ;
	assign \g10049/_0_  = _w18584_ ;
	assign \g10050/_0_  = _w18587_ ;
	assign \g10051/_0_  = _w18590_ ;
	assign \g10052/_0_  = _w18593_ ;
	assign \g10053/_0_  = _w18597_ ;
	assign \g10054/_0_  = _w18600_ ;
	assign \g10055/_0_  = _w18603_ ;
	assign \g10056/_0_  = _w18606_ ;
	assign \g10057/_0_  = _w18609_ ;
	assign \g10058/_0_  = _w18612_ ;
	assign \g10059/_0_  = _w18615_ ;
	assign \g10060/_0_  = _w18618_ ;
	assign \g10061/_0_  = _w18621_ ;
	assign \g10062/_0_  = _w18624_ ;
	assign \g10063/_0_  = _w18627_ ;
	assign \g10064/_0_  = _w18630_ ;
	assign \g10065/_0_  = _w18633_ ;
	assign \g10066/_0_  = _w18636_ ;
	assign \g10067/_0_  = _w18639_ ;
	assign \g10068/_0_  = _w18642_ ;
	assign \g10069/_0_  = _w18645_ ;
	assign \g10070/_0_  = _w18648_ ;
	assign \g10071/_0_  = _w18651_ ;
	assign \g10072/_0_  = _w18657_ ;
	assign \g10073/_0_  = _w18660_ ;
	assign \g10074/_0_  = _w18663_ ;
	assign \g10075/_0_  = _w18666_ ;
	assign \g10076/_0_  = _w18669_ ;
	assign \g10077/_0_  = _w18672_ ;
	assign \g10078/_0_  = _w18675_ ;
	assign \g10080/_0_  = _w18678_ ;
	assign \g10081/_0_  = _w18687_ ;
	assign \g10083/_0_  = _w18692_ ;
	assign \g10089/_0_  = _w18695_ ;
	assign \g1009/_0_  = _w18701_ ;
	assign \g10090/_0_  = _w18704_ ;
	assign \g10091/_0_  = _w18707_ ;
	assign \g10092/_0_  = _w18710_ ;
	assign \g10093/_0_  = _w18713_ ;
	assign \g10094/_0_  = _w18716_ ;
	assign \g1010/_0_  = _w18836_ ;
	assign \g10108/_3_  = _w18852_ ;
	assign \g1011/_0_  = _w18855_ ;
	assign \g10110/_0_  = _w18864_ ;
	assign \g10111/_0_  = _w18873_ ;
	assign \g10113/_3_  = _w18877_ ;
	assign \g10115/_3_  = _w18881_ ;
	assign \g1013/_0_  = _w18884_ ;
	assign \g1014/_0_  = _w18945_ ;
	assign \g10152/_0_  = _w18950_ ;
	assign \g10153/_0_  = _w18953_ ;
	assign \g10154/_0_  = _w18956_ ;
	assign \g10155/_0_  = _w18959_ ;
	assign \g10156/_0_  = _w18962_ ;
	assign \g10157/_0_  = _w18965_ ;
	assign \g10158/_0_  = _w18968_ ;
	assign \g10159/_0_  = _w18971_ ;
	assign \g1016/_0_  = _w19013_ ;
	assign \g10160/_0_  = _w19017_ ;
	assign \g10161/_0_  = _w19020_ ;
	assign \g10162/_0_  = _w19023_ ;
	assign \g10163/_0_  = _w19027_ ;
	assign \g10164/_0_  = _w19030_ ;
	assign \g10165/_0_  = _w19033_ ;
	assign \g1017/_0_  = _w19037_ ;
	assign \g10170/_3_  = _w19059_ ;
	assign \g1018/_0_  = _w19062_ ;
	assign \g10190/_3_  = _w19064_ ;
	assign \g10194/_3_  = _w19066_ ;
	assign \g10198/_0_  = _w19133_ ;
	assign \g10199/_0_  = _w19200_ ;
	assign \g102/_0_  = _w19363_ ;
	assign \g103/_0_  = _w19392_ ;
	assign \g104/_0_  = _w19402_ ;
	assign \g105/_0_  = _w19409_ ;
	assign \g10598/_0_  = _w19413_ ;
	assign \g106/_0_  = _w19436_ ;
	assign \g10667/_0_  = _w19440_ ;
	assign \g10683/_0_  = _w19476_ ;
	assign \g10685/_0_  = _w19498_ ;
	assign \g107/_0_  = _w19527_ ;
	assign \g10721/_0_  = _w19533_ ;
	assign \g10758/_0_  = _w19540_ ;
	assign \g10765/_0_  = _w19543_ ;
	assign \g10778/_0_  = _w19554_ ;
	assign \g10791/_0_  = _w19555_ ;
	assign \g108/_0_  = _w19694_ ;
	assign \g10887/_0_  = _w19707_ ;
	assign \g1089/_0_  = _w19774_ ;
	assign \g109/_0_  = _w19783_ ;
	assign \g1090/_0_  = _w19845_ ;
	assign \g1091/_0_  = _w19900_ ;
	assign \g1092/_0_  = _w19903_ ;
	assign \g10923/_0_  = _w19906_ ;
	assign \g1093/_0_  = _w19909_ ;
	assign \g10930/_0_  = _w19915_ ;
	assign \g10931/_0_  = _w19918_ ;
	assign \g10936/_0_  = _w19926_ ;
	assign \g1097/_0_  = _w19929_ ;
	assign \g11/_0_  = _w19963_ ;
	assign \g110/_0_  = _w19969_ ;
	assign \g1101/_0_  = _w20035_ ;
	assign \g11013/_0_  = _w20044_ ;
	assign \g1102/_0_  = _w20058_ ;
	assign \g1103/_0_  = _w20061_ ;
	assign \g11032/_0_  = _w20077_ ;
	assign \g1104/_0_  = _w20147_ ;
	assign \g1105/_0_  = _w20197_ ;
	assign \g1107/_0_  = _w20200_ ;
	assign \g11074/_0_  = _w20222_ ;
	assign \g11077/_0_  = _w20225_ ;
	assign \g1108/_0_  = _w20228_ ;
	assign \g1109/_0_  = _w20231_ ;
	assign \g11112/_0_  = _w20242_ ;
	assign \g11115/_0_  = _w20245_ ;
	assign \g11116/_0_  = _w20248_ ;
	assign \g11119/_0_  = _w20255_ ;
	assign \g11120/_0_  = _w20256_ ;
	assign \g1113/_0_  = _w20293_ ;
	assign \g1115/_0_  = _w20331_ ;
	assign \g1116/_0_  = _w20334_ ;
	assign \g1117/_0_  = _w20337_ ;
	assign \g11267/_0_  = _w20340_ ;
	assign \g11281/_0_  = _w20353_ ;
	assign \g11287/_0_  = _w20375_ ;
	assign \g11300/_0_  = _w20380_ ;
	assign \g11323/_0_  = _w20385_ ;
	assign \g11325/_2__syn_2  = _w20396_ ;
	assign \g11345/_2_  = _w20399_ ;
	assign \g11470/_0_  = _w20405_ ;
	assign \g11471/_0_  = _w20423_ ;
	assign \g11472/_0_  = _w20427_ ;
	assign \g11473/_0_  = _w20445_ ;
	assign \g11474/_0_  = _w20449_ ;
	assign \g11476/_0_  = _w20452_ ;
	assign \g11477/_0_  = _w20463_ ;
	assign \g11496/_0_  = _w20482_ ;
	assign \g11497/_0_  = _w20491_ ;
	assign \g11498/_0_  = _w20500_ ;
	assign \g11499/_0_  = _w20506_ ;
	assign \g11500/_0_  = _w20515_ ;
	assign \g11501/_0_  = _w20521_ ;
	assign \g11502/_0_  = _w20530_ ;
	assign \g11503/_0_  = _w20536_ ;
	assign \g11504/_0_  = _w20544_ ;
	assign \g11505/_0_  = _w20552_ ;
	assign \g11506/_0_  = _w20558_ ;
	assign \g11507/_0_  = _w20564_ ;
	assign \g11509/_0_  = _w20567_ ;
	assign \g11510/_0_  = _w20570_ ;
	assign \g11515/_0_  = _w20588_ ;
	assign \g11516/_0_  = _w20591_ ;
	assign \g11520/_0_  = _w20594_ ;
	assign \g11521/_0_  = _w20600_ ;
	assign \g11576/_0_  = _w20612_ ;
	assign \g11577/_0_  = _w20622_ ;
	assign \g11578/_0_  = _w20632_ ;
	assign \g11579/_0_  = _w20642_ ;
	assign \g11580/_0_  = _w20652_ ;
	assign \g11581/_0_  = _w20660_ ;
	assign \g11582/_0_  = _w20671_ ;
	assign \g11583/_0_  = _w20682_ ;
	assign \g11584/_0_  = _w20693_ ;
	assign \g11585/_0_  = _w20704_ ;
	assign \g11586/_0_  = _w20715_ ;
	assign \g11587/_0_  = _w20726_ ;
	assign \g11588/_0_  = _w20737_ ;
	assign \g11589/_0_  = _w20753_ ;
	assign \g11591/_0_  = _w20763_ ;
	assign \g11593/_0_  = _w20773_ ;
	assign \g11595/_0_  = _w20780_ ;
	assign \g11596/_0_  = _w20783_ ;
	assign \g11597/_0_  = _w20786_ ;
	assign \g11605/_0_  = _w20791_ ;
	assign \g11606/_0_  = _w20794_ ;
	assign \g11607/_0_  = _w20797_ ;
	assign \g11608/_0_  = _w20800_ ;
	assign \g11609/_0_  = _w20803_ ;
	assign \g11610/_0_  = _w20806_ ;
	assign \g11611/_0_  = _w20809_ ;
	assign \g11612/_0_  = _w20812_ ;
	assign \g11613/_0_  = _w20815_ ;
	assign \g11615/_0_  = _w20820_ ;
	assign \g11616/_0_  = _w20832_ ;
	assign \g11617/_0_  = _w20837_ ;
	assign \g11651/_3_  = _w20840_ ;
	assign \g11704/_0_  = _w20842_ ;
	assign \g11705/_0_  = _w20844_ ;
	assign \g11709/_0_  = _w20852_ ;
	assign \g11722/_0_  = _w20861_ ;
	assign \g11723/_0_  = _w20863_ ;
	assign \g119/_0_  = _w20867_ ;
	assign \g1192/_0_  = _w20988_ ;
	assign \g11994/_0_  = _w20989_ ;
	assign \g120/_0_  = _w20993_ ;
	assign \g1200/_0_  = _w21051_ ;
	assign \g12003/_0_  = _w21054_ ;
	assign \g1201/_0_  = _w21057_ ;
	assign \g12019/_0_  = _w21060_ ;
	assign \g1203/_3_  = _w21070_ ;
	assign \g1204/_3_  = _w21076_ ;
	assign \g1207/_0_  = _w21129_ ;
	assign \g1208/_0_  = _w21132_ ;
	assign \g12092/_0_  = _w21140_ ;
	assign \g1210/_0_  = _w21179_ ;
	assign \g1211/_0_  = _w21231_ ;
	assign \g1212/_0_  = _w21234_ ;
	assign \g1213/_0_  = _w21237_ ;
	assign \g12145/_0_  = _w21246_ ;
	assign \g12155/_0_  = _w21254_ ;
	assign \g12186/_0_  = _w21261_ ;
	assign \g12187/_0_  = _w21264_ ;
	assign \g12192/_0_  = _w21267_ ;
	assign \g12201/_0_  = _w21276_ ;
	assign \g12202/_0_  = _w21280_ ;
	assign \g12203/_0_  = _w21284_ ;
	assign \g12204/_0_  = _w21287_ ;
	assign \g12207/_0_  = _w21290_ ;
	assign \g12229/_3_  = _w21300_ ;
	assign \g12267/_0_  = _w21301_ ;
	assign \g12276/_0_  = _w21304_ ;
	assign \g12278/_0_  = _w21307_ ;
	assign \g12279/_0_  = _w21310_ ;
	assign \g12280/_0_  = _w21313_ ;
	assign \g12302/_0_  = _w21315_ ;
	assign \g12316/_0_  = _w21322_ ;
	assign \g12317/_0_  = _w21326_ ;
	assign \g12319/_0_  = _w21330_ ;
	assign \g12328/_3_  = _w21339_ ;
	assign \g1233/_0_  = _w10069_ ;
	assign \g12348/_0_  = _w21343_ ;
	assign \g12351/_0_  = _w21347_ ;
	assign \g12352/_0_  = _w21351_ ;
	assign \g12353/_0_  = _w21355_ ;
	assign \g12354/_0_  = _w21359_ ;
	assign \g12355/_0_  = _w21363_ ;
	assign \g1237/_0_  = _w8113_ ;
	assign \g124/_0_  = _w21366_ ;
	assign \g12444/_0_  = _w21371_ ;
	assign \g125/_0_  = _w21374_ ;
	assign \g12637/_0_  = _w21382_ ;
	assign \g12639/_0_  = _w21390_ ;
	assign \g12658/_0_  = _w21399_ ;
	assign \g12659/_0_  = _w21409_ ;
	assign \g12660/_0_  = _w21419_ ;
	assign \g12663/_0_  = _w21425_ ;
	assign \g12664/_0_  = _w21432_ ;
	assign \g12665/_0_  = _w21437_ ;
	assign \g12672/_3_  = _w21446_ ;
	assign \g12673/_3_  = _w21455_ ;
	assign \g12674/_3_  = _w21464_ ;
	assign \g12675/_3_  = _w21473_ ;
	assign \g12676/_3_  = _w21482_ ;
	assign \g12677/_3_  = _w21491_ ;
	assign \g12678/_0_  = _w21496_ ;
	assign \g12679/_3_  = _w21505_ ;
	assign \g12697/_3_  = _w21514_ ;
	assign \g12701/_3_  = _w21523_ ;
	assign \g12711/_2_  = _w21535_ ;
	assign \g12713/_2_  = _w21541_ ;
	assign \g12715/_2_  = _w21549_ ;
	assign \g12717/_2_  = _w21555_ ;
	assign \g12718/_2__syn_2  = _w21562_ ;
	assign \g1272/_0_  = _w21577_ ;
	assign \g12728/_1__syn_2  = _w21579_ ;
	assign \g12730/_3_  = _w21588_ ;
	assign \g12741/_1__syn_2  = _w21592_ ;
	assign \g12746/_0__syn_2  = _w18689_ ;
	assign \g12748/_0_  = _w21598_ ;
	assign \g12749/_0_  = _w21601_ ;
	assign \g12759/_1__syn_2  = _w18233_ ;
	assign \g12760/_0_  = _w21605_ ;
	assign \g12762/_0_  = _w21609_ ;
	assign \g12763/_0_  = _w21612_ ;
	assign \g12764/_0_  = _w21615_ ;
	assign \g12765/_0_  = _w21618_ ;
	assign \g12766/_0_  = _w21621_ ;
	assign \g12767/_0_  = _w21624_ ;
	assign \g12768/_0_  = _w21627_ ;
	assign \g12769/_0_  = _w21630_ ;
	assign \g12770/_0_  = _w21633_ ;
	assign \g12771/_0_  = _w21636_ ;
	assign \g12772/_0_  = _w21639_ ;
	assign \g12773/_0_  = _w21642_ ;
	assign \g12774/_0_  = _w21645_ ;
	assign \g12775/_0_  = _w21648_ ;
	assign \g12776/_0_  = _w21651_ ;
	assign \g12777/_0_  = _w21654_ ;
	assign \g12778/_0_  = _w21657_ ;
	assign \g12779/_0_  = _w21660_ ;
	assign \g1278/_0_  = _w21705_ ;
	assign \g12780/_0_  = _w21709_ ;
	assign \g12781/_0_  = _w21712_ ;
	assign \g12782/_0_  = _w21715_ ;
	assign \g12783/_0_  = _w21718_ ;
	assign \g12784/_0_  = _w21721_ ;
	assign \g12785/_0_  = _w21724_ ;
	assign \g12786/_0_  = _w21727_ ;
	assign \g12787/_0_  = _w21730_ ;
	assign \g12788/_0_  = _w21733_ ;
	assign \g12789/_0_  = _w21736_ ;
	assign \g12790/_0_  = _w21739_ ;
	assign \g12791/_0_  = _w21742_ ;
	assign \g12792/_0_  = _w21745_ ;
	assign \g12793/_0_  = _w21748_ ;
	assign \g12794/_0_  = _w21751_ ;
	assign \g12795/_0_  = _w21754_ ;
	assign \g12796/_0_  = _w21757_ ;
	assign \g12797/_0_  = _w21760_ ;
	assign \g12798/_0_  = _w21764_ ;
	assign \g12799/_0_  = _w21767_ ;
	assign \g12800/_0_  = _w21770_ ;
	assign \g12801/_0_  = _w21773_ ;
	assign \g12802/_0_  = _w21776_ ;
	assign \g12803/_0_  = _w21779_ ;
	assign \g12804/_0_  = _w21782_ ;
	assign \g12805/_0_  = _w21785_ ;
	assign \g12806/_0_  = _w21788_ ;
	assign \g12807/_0_  = _w21791_ ;
	assign \g12808/_0_  = _w21794_ ;
	assign \g12809/_0_  = _w21797_ ;
	assign \g1281/_0_  = _w21803_ ;
	assign \g12810/_0_  = _w21806_ ;
	assign \g12811/_0_  = _w21809_ ;
	assign \g12812/_0_  = _w21812_ ;
	assign \g12813/_0_  = _w21815_ ;
	assign \g12814/_0_  = _w21818_ ;
	assign \g12815/_0_  = _w21821_ ;
	assign \g12816/_0_  = _w21824_ ;
	assign \g12817/_0_  = _w21827_ ;
	assign \g12818/_0_  = _w21830_ ;
	assign \g12819/_0_  = _w21833_ ;
	assign \g1282/_0_  = _w21836_ ;
	assign \g12820/_0_  = _w21839_ ;
	assign \g12821/_0_  = _w21842_ ;
	assign \g12822/_0_  = _w21845_ ;
	assign \g12823/_0_  = _w21848_ ;
	assign \g12824/_0_  = _w21851_ ;
	assign \g12825/_0_  = _w21854_ ;
	assign \g12826/_0_  = _w21857_ ;
	assign \g12827/_0_  = _w21860_ ;
	assign \g12828/_0_  = _w21863_ ;
	assign \g12829/_0_  = _w21866_ ;
	assign \g12830/_0_  = _w21869_ ;
	assign \g12831/_0_  = _w21873_ ;
	assign \g12832/_0_  = _w21879_ ;
	assign \g12833/_0_  = _w21881_ ;
	assign \g12835/_0_  = _w21884_ ;
	assign \g12836/_0_  = _w21887_ ;
	assign \g12838/_0_  = _w21890_ ;
	assign \g12848/_0_  = _w21895_ ;
	assign \g12849/_0_  = _w21899_ ;
	assign \g1285/_0_  = _w21902_ ;
	assign \g12850/_0_  = _w21905_ ;
	assign \g12857/_0_  = _w21909_ ;
	assign \g12858/_0_  = _w21912_ ;
	assign \g12859/_0_  = _w21915_ ;
	assign \g12861/_0_  = _w21918_ ;
	assign \g12862/_0_  = _w21921_ ;
	assign \g12868/_0_  = _w21926_ ;
	assign \g12869/_0_  = _w21929_ ;
	assign \g1287/_0_  = _w21963_ ;
	assign \g12870/_0_  = _w21966_ ;
	assign \g12871/_0_  = _w21969_ ;
	assign \g12872/_0_  = _w21972_ ;
	assign \g12873/_0_  = _w21975_ ;
	assign \g12874/_0_  = _w21979_ ;
	assign \g12875/_0_  = _w21982_ ;
	assign \g12876/_0_  = _w21985_ ;
	assign \g12877/_0_  = _w21988_ ;
	assign \g12878/_0_  = _w22000_ ;
	assign \g12879/_0_  = _w22009_ ;
	assign \g12880/_0_  = _w22018_ ;
	assign \g12881/_0_  = _w22027_ ;
	assign \g12882/_0_  = _w22036_ ;
	assign \g12883/_0_  = _w22045_ ;
	assign \g12884/_0_  = _w22054_ ;
	assign \g12885/_0_  = _w22063_ ;
	assign \g12886/_0_  = _w22072_ ;
	assign \g12887/_0_  = _w22081_ ;
	assign \g12888/_0_  = _w22090_ ;
	assign \g12889/_0_  = _w22099_ ;
	assign \g1289/_0_  = _w22102_ ;
	assign \g12890/_0_  = _w22111_ ;
	assign \g12891/_0_  = _w22120_ ;
	assign \g12894/_0_  = _w22123_ ;
	assign \g12898/_0_  = _w22127_ ;
	assign \g12899/_0_  = _w22130_ ;
	assign \g12900/_0_  = _w22133_ ;
	assign \g12901/_0_  = _w22136_ ;
	assign \g12902/_0_  = _w22139_ ;
	assign \g12903/_0_  = _w22142_ ;
	assign \g12906/_0_  = _w22145_ ;
	assign \g12907/_0_  = _w22148_ ;
	assign \g12908/_0_  = _w22157_ ;
	assign \g12912/_0_  = _w22161_ ;
	assign \g12913/_0_  = _w22164_ ;
	assign \g12914/_0_  = _w22167_ ;
	assign \g12915/_0_  = _w22170_ ;
	assign \g12916/_0_  = _w22173_ ;
	assign \g12917/_0_  = _w22176_ ;
	assign \g12918/_0_  = _w22179_ ;
	assign \g12919/_0_  = _w22182_ ;
	assign \g12920/_0_  = _w22185_ ;
	assign \g12921/_0_  = _w22188_ ;
	assign \g12922/_0_  = _w22191_ ;
	assign \g12923/_0_  = _w22194_ ;
	assign \g12924/_0_  = _w22197_ ;
	assign \g12925/_0_  = _w22200_ ;
	assign \g12926/_0_  = _w22203_ ;
	assign \g12932/_0_  = _w22206_ ;
	assign \g12933/_0_  = _w22209_ ;
	assign \g12936/_0_  = _w22212_ ;
	assign \g12955/_0_  = _w22215_ ;
	assign \g13015/_0_  = _w22218_ ;
	assign \g13016/_0_  = _w22221_ ;
	assign \g13017/_0_  = _w22224_ ;
	assign \g13018/_0_  = _w22227_ ;
	assign \g13019/_0_  = _w22229_ ;
	assign \g13020/_0_  = _w22232_ ;
	assign \g13021/_0_  = _w22235_ ;
	assign \g13024/_0_  = _w22238_ ;
	assign \g13025/_0_  = _w22241_ ;
	assign \g13027/_0_  = _w22244_ ;
	assign \g13028/_0_  = _w22247_ ;
	assign \g13030/_0_  = _w22250_ ;
	assign \g13031/_0_  = _w22253_ ;
	assign \g13033/_0_  = _w22256_ ;
	assign \g13047/_0_  = _w22259_ ;
	assign \g13060/_0_  = _w22262_ ;
	assign \g13062/_0_  = _w22265_ ;
	assign \g13063/_0_  = _w22268_ ;
	assign \g13064/_0_  = _w22271_ ;
	assign \g13067/_0_  = _w22274_ ;
	assign \g13068/_0_  = _w22277_ ;
	assign \g13069/_0_  = _w22280_ ;
	assign \g13070/_0_  = _w22283_ ;
	assign \g13072/_0_  = _w22286_ ;
	assign \g13094/_0_  = _w22288_ ;
	assign \g13104/_0_  = _w22294_ ;
	assign \g13110/_0_  = _w22297_ ;
	assign \g13114/_0_  = _w22301_ ;
	assign \g13115/_0_  = _w22304_ ;
	assign \g13116/_0_  = _w22307_ ;
	assign \g13117/_0_  = _w22310_ ;
	assign \g13118/_0_  = _w22313_ ;
	assign \g13119/_0_  = _w22316_ ;
	assign \g13120/_0_  = _w22319_ ;
	assign \g13121/_0_  = _w22322_ ;
	assign \g13124/_0_  = _w22325_ ;
	assign \g13125/_0_  = _w22328_ ;
	assign \g13127/_0_  = _w22331_ ;
	assign \g13128/_0_  = _w22334_ ;
	assign \g13129/_0_  = _w22337_ ;
	assign \g13130/_0_  = _w22340_ ;
	assign \g13131/_0_  = _w22343_ ;
	assign \g13132/_0_  = _w22346_ ;
	assign \g13133/_0_  = _w22349_ ;
	assign \g13134/_0_  = _w22352_ ;
	assign \g13138/_0_  = _w22355_ ;
	assign \g13139/_0_  = _w22358_ ;
	assign \g13140/_0_  = _w22361_ ;
	assign \g13141/_0_  = _w22364_ ;
	assign \g13142/_0_  = _w22367_ ;
	assign \g13143/_0_  = _w22370_ ;
	assign \g13144/_0_  = _w22373_ ;
	assign \g13146/_0_  = _w22376_ ;
	assign \g13150/_0_  = _w22379_ ;
	assign \g13152/_0_  = _w22382_ ;
	assign \g13154/_0_  = _w22385_ ;
	assign \g13155/_0_  = _w22388_ ;
	assign \g13156/_0_  = _w22391_ ;
	assign \g13157/_0_  = _w22394_ ;
	assign \g13158/_0_  = _w22397_ ;
	assign \g1320/_3_  = _w22432_ ;
	assign \g13266/_0_  = _w22435_ ;
	assign \g13269/_0_  = _w22438_ ;
	assign \g13274/_0_  = _w22441_ ;
	assign \g13277/_0_  = _w22444_ ;
	assign \g13280/_0_  = _w22447_ ;
	assign \g13283/_0_  = _w22450_ ;
	assign \g13294/_0_  = _w22453_ ;
	assign \g13330/_0_  = _w22456_ ;
	assign \g13333/_0_  = _w22461_ ;
	assign \g13334/_0_  = _w22464_ ;
	assign \g13335/_0_  = _w22467_ ;
	assign \g13336/_0_  = _w22470_ ;
	assign \g13337/_0_  = _w22473_ ;
	assign \g13338/_0_  = _w22476_ ;
	assign \g13345/_0_  = _w22480_ ;
	assign \g13346/_0_  = _w22483_ ;
	assign \g13347/_0_  = _w22487_ ;
	assign \g13348/_0_  = _w22490_ ;
	assign \g13349/_0_  = _w22493_ ;
	assign \g13350/_0_  = _w22496_ ;
	assign \g13351/_0_  = _w22499_ ;
	assign \g13352/_0_  = _w22502_ ;
	assign \g13486/_0_  = _w22504_ ;
	assign \g13488/_0_  = _w22506_ ;
	assign \g13508/_0_  = _w22509_ ;
	assign \g13509/_0_  = _w22512_ ;
	assign \g13510/_0_  = _w22515_ ;
	assign \g13511/_0_  = _w22518_ ;
	assign \g13512/_0_  = _w22521_ ;
	assign \g13513/_0_  = _w22524_ ;
	assign \g13514/_0_  = _w22527_ ;
	assign \g13515/_0_  = _w22530_ ;
	assign \g13516/_0_  = _w22533_ ;
	assign \g13517/_0_  = _w22536_ ;
	assign \g13518/_0_  = _w22539_ ;
	assign \g13519/_0_  = _w22542_ ;
	assign \g13520/_0_  = _w22545_ ;
	assign \g13521/_0_  = _w22548_ ;
	assign \g13540/_0_  = _w22551_ ;
	assign \g13541/_0_  = _w22554_ ;
	assign \g13542/_0_  = _w22557_ ;
	assign \g13543/_0_  = _w22560_ ;
	assign \g13544/_0_  = _w22563_ ;
	assign \g13545/_0_  = _w22566_ ;
	assign \g13546/_0_  = _w22569_ ;
	assign \g13547/_0_  = _w22572_ ;
	assign \g13548/_0_  = _w22575_ ;
	assign \g13549/_0_  = _w22578_ ;
	assign \g13550/_0_  = _w22580_ ;
	assign \g13551/_0_  = _w22585_ ;
	assign \g13552/_0_  = _w22587_ ;
	assign \g13553/_0_  = _w22589_ ;
	assign \g13554/_0_  = _w22592_ ;
	assign \g13555/_0_  = _w22595_ ;
	assign \g13556/_0_  = _w22598_ ;
	assign \g13557/_0_  = _w22601_ ;
	assign \g13558/_0_  = _w22604_ ;
	assign \g13559/_0_  = _w22607_ ;
	assign \g13560/_0_  = _w22610_ ;
	assign \g13561/_0_  = _w22613_ ;
	assign \g13562/_0_  = _w22616_ ;
	assign \g13563/_0_  = _w22619_ ;
	assign \g13564/_0_  = _w22622_ ;
	assign \g13565/_0_  = _w22625_ ;
	assign \g13566/_0_  = _w22628_ ;
	assign \g13567/_0_  = _w22631_ ;
	assign \g13568/_0_  = _w22634_ ;
	assign \g13569/_0_  = _w22637_ ;
	assign \g13570/_0_  = _w22640_ ;
	assign \g13571/_0_  = _w22643_ ;
	assign \g13572/_0_  = _w22646_ ;
	assign \g137/_3_  = _w22680_ ;
	assign \g1387/_3_  = _w22690_ ;
	assign \g1388/_3_  = _w22696_ ;
	assign \g1389/_0_  = _w22701_ ;
	assign \g139/_0_  = _w22883_ ;
	assign \g1390/_0_  = _w22916_ ;
	assign \g1393/_0_  = _w22919_ ;
	assign \g140/_0_  = _w22926_ ;
	assign \g141/_0_  = _w22929_ ;
	assign \g14173/_0_  = _w22933_ ;
	assign \g14176/_0_  = _w22936_ ;
	assign \g142/_3_  = _w22961_ ;
	assign \g14273/_1__syn_2  = _w20402_ ;
	assign \g14274/_0_  = _w22962_ ;
	assign \g14280/_0_  = _w22973_ ;
	assign \g14281/_0_  = _w22984_ ;
	assign \g143/_3_  = _w23001_ ;
	assign \g14354/_3__syn_2  = _w13779_ ;
	assign \g14370/_0_  = _w23004_ ;
	assign \g14385/_0_  = _w23008_ ;
	assign \g14386/_0_  = _w23011_ ;
	assign \g144/_3_  = _w23017_ ;
	assign \g14407/_0_  = _w23023_ ;
	assign \g14412/_0_  = _w23026_ ;
	assign \g14435/_0_  = _w23035_ ;
	assign \g14439/_0_  = _w23037_ ;
	assign \g145/_0_  = _w23089_ ;
	assign \g14522/_0_  = _w23091_ ;
	assign \g14528/_0_  = _w23093_ ;
	assign \g14533/_0_  = _w23116_ ;
	assign \g14581/_1_  = _w23117_ ;
	assign \g14582/_0_  = _w23118_ ;
	assign \g146/_3_  = _w23124_ ;
	assign \g14671/_0_  = _w23135_ ;
	assign \g14672/_0_  = _w23146_ ;
	assign \g147/_0_  = _w23188_ ;
	assign \g1473/_0_  = _w23205_ ;
	assign \g148/_0_  = _w23222_ ;
	assign \g14826/_0_  = _w19024_ ;
	assign \g149/_0_  = _w23228_ ;
	assign \g14908/_0_  = _w23234_ ;
	assign \g14911/_0_  = _w23240_ ;
	assign \g14936/_2_  = _w23243_ ;
	assign \g1494/_0_  = _w23259_ ;
	assign \g1495/_0_  = _w23262_ ;
	assign \g14950/_2_  = _w23274_ ;
	assign \g14953/_2_  = _w23286_ ;
	assign \g15003/_0_  = _w23290_ ;
	assign \g15004/_0_  = _w23293_ ;
	assign \g15006/_0_  = _w23296_ ;
	assign \g15007/_0_  = _w23299_ ;
	assign \g15008/_0_  = _w23302_ ;
	assign \g15009/_0_  = _w23305_ ;
	assign \g15010/_0_  = _w23308_ ;
	assign \g15011/_0_  = _w23311_ ;
	assign \g15012/_0_  = _w23314_ ;
	assign \g15013/_0_  = _w23317_ ;
	assign \g15014/_0_  = _w23320_ ;
	assign \g15015/_0_  = _w23323_ ;
	assign \g15016/_0_  = _w23326_ ;
	assign \g15017/_0_  = _w23329_ ;
	assign \g15018/_0_  = _w23332_ ;
	assign \g15019/_0_  = _w23335_ ;
	assign \g15035/_0_  = _w23339_ ;
	assign \g15036/_0_  = _w23342_ ;
	assign \g15038/_0_  = _w23349_ ;
	assign \g15039/_0_  = _w23355_ ;
	assign \g15040/_0_  = _w23361_ ;
	assign \g15041/_0_  = _w23367_ ;
	assign \g15042/_0_  = _w23373_ ;
	assign \g15043/_0_  = _w23379_ ;
	assign \g15044/_0_  = _w23385_ ;
	assign \g15045/_0_  = _w23391_ ;
	assign \g15046/_0_  = _w23397_ ;
	assign \g15056/_00_  = _w23403_ ;
	assign \g151/_0_  = _w23406_ ;
	assign \g15193/_0_  = _w23413_ ;
	assign \g152/_0_  = _w23416_ ;
	assign \g15256/_0_  = _w23425_ ;
	assign \g153/_0_  = _w23428_ ;
	assign \g15393/_0_  = _w23436_ ;
	assign \g15394/_0_  = _w23442_ ;
	assign \g15395/_0_  = _w23448_ ;
	assign \g15396/_0_  = _w23454_ ;
	assign \g15397/_0_  = _w23460_ ;
	assign \g15398/_0_  = _w23466_ ;
	assign \g15399/_0_  = _w23472_ ;
	assign \g154/_0_  = _w23475_ ;
	assign \g15400/_0_  = _w23481_ ;
	assign \g15401/_0_  = _w23487_ ;
	assign \g15402/_0_  = _w23493_ ;
	assign \g15403/_0_  = _w23499_ ;
	assign \g15404/_0_  = _w23505_ ;
	assign \g15405/_0_  = _w23511_ ;
	assign \g15406/_0_  = _w23517_ ;
	assign \g15407/_0_  = _w23523_ ;
	assign \g15408/_0_  = _w23529_ ;
	assign \g15473/_0_  = _w23534_ ;
	assign \g15650/_0_  = _w23536_ ;
	assign \g15651/_0_  = _w23538_ ;
	assign \g15652/_0_  = _w23540_ ;
	assign \g15653/_0_  = _w23542_ ;
	assign \g15662/_0_  = _w23545_ ;
	assign \g15663/_0_  = _w23548_ ;
	assign \g15664/_0_  = _w23551_ ;
	assign \g15665/_0_  = _w23554_ ;
	assign \g15666/_0_  = _w23557_ ;
	assign \g15667/_0_  = _w23560_ ;
	assign \g15668/_0_  = _w23563_ ;
	assign \g15669/_0_  = _w23566_ ;
	assign \g15670/_0_  = _w23569_ ;
	assign \g15671/_0_  = _w23572_ ;
	assign \g15672/_0_  = _w23575_ ;
	assign \g15673/_0_  = _w23578_ ;
	assign \g15674/_0_  = _w23581_ ;
	assign \g15675/_0_  = _w23584_ ;
	assign \g1569/_0_  = _w23676_ ;
	assign \g1570/_0_  = _w23680_ ;
	assign \g1575/_0_  = _w23686_ ;
	assign \g1576/_0_  = _w23689_ ;
	assign \g15922/_1_  = _w23690_ ;
	assign \g15970/_0_  = _w23691_ ;
	assign \g16059/_0_  = _w23694_ ;
	assign \g1606/_3_  = _w23704_ ;
	assign \g16124/_0_  = _w20576_ ;
	assign \g16144/_0_  = _w23706_ ;
	assign \g16202/_0_  = _w23709_ ;
	assign \g16214/_0_  = _w23713_ ;
	assign \g16247/_0_  = _w23719_ ;
	assign \g16257/_0_  = _w23725_ ;
	assign \g16274/_1_  = _w23726_ ;
	assign \g16324/_0_  = _w20787_ ;
	assign \g16343/_1__syn_2  = _w22291_ ;
	assign \g16381/_0_  = _w23730_ ;
	assign \g16383/_0_  = _w23739_ ;
	assign \g16386/_0_  = _w23742_ ;
	assign \g16414/_1__syn_2  = _w21906_ ;
	assign \g16416/_0__syn_2  = _w20864_ ;
	assign \g16448/_0_  = _w23743_ ;
	assign \g16460/_1_  = _w23744_ ;
	assign \g16625/_3_  = _w23033_ ;
	assign \g16662/_0_  = _w23751_ ;
	assign \g16668/_1__syn_2  = _w22477_ ;
	assign \g16692/_0_  = _w23753_ ;
	assign \g16721/_0_  = _w23760_ ;
	assign \g16723/_0_  = _w23765_ ;
	assign \g16725/_0_  = _w23769_ ;
	assign \g16726/_0_  = _w23772_ ;
	assign \g16727/_0_  = _w23775_ ;
	assign \g16728/_0_  = _w23778_ ;
	assign \g16729/_0_  = _w23781_ ;
	assign \g16730/_0_  = _w23785_ ;
	assign \g16731/_0_  = _w23788_ ;
	assign \g16732/_0_  = _w23791_ ;
	assign \g16733/_0_  = _w23794_ ;
	assign \g16734/_0_  = _w23797_ ;
	assign \g16735/_0_  = _w23801_ ;
	assign \g16736/_0_  = _w23804_ ;
	assign \g16737/_0_  = _w23807_ ;
	assign \g16738/_0_  = _w23810_ ;
	assign \g16739/_0_  = _w23813_ ;
	assign \g16740/_0_  = _w23817_ ;
	assign \g16741/_0_  = _w23820_ ;
	assign \g16742/_0_  = _w23823_ ;
	assign \g16743/_0_  = _w23826_ ;
	assign \g16747/_0_  = _w23830_ ;
	assign \g16748/_0_  = _w23833_ ;
	assign \g16749/_0_  = _w23836_ ;
	assign \g16750/_0_  = _w23839_ ;
	assign \g16753/_0_  = _w23842_ ;
	assign \g16754/_0_  = _w23845_ ;
	assign \g16755/_0_  = _w23848_ ;
	assign \g16756/_0_  = _w23851_ ;
	assign \g16757/_0_  = _w23854_ ;
	assign \g16758/_0_  = _w23857_ ;
	assign \g16761/_0_  = _w23863_ ;
	assign \g16765/_0_  = _w23868_ ;
	assign \g16766/_0_  = _w23871_ ;
	assign \g16767/_0_  = _w23874_ ;
	assign \g16768/_0_  = _w23877_ ;
	assign \g16769/_0_  = _w23880_ ;
	assign \g16772/_0_  = _w23883_ ;
	assign \g16785/_0_  = _w23888_ ;
	assign \g16786/_0_  = _w23892_ ;
	assign \g16787/_0_  = _w23895_ ;
	assign \g16788/_0_  = _w23898_ ;
	assign \g16789/_0_  = _w23901_ ;
	assign \g16790/_0_  = _w23904_ ;
	assign \g16791/_0_  = _w23907_ ;
	assign \g16804/_0_  = _w23911_ ;
	assign \g16805/_0_  = _w23914_ ;
	assign \g16806/_0_  = _w23917_ ;
	assign \g16807/_0_  = _w23923_ ;
	assign \g16808/_0_  = _w23926_ ;
	assign \g16809/_0_  = _w23929_ ;
	assign \g16810/_0_  = _w23933_ ;
	assign \g16811/_0_  = _w23936_ ;
	assign \g16812/_0_  = _w23939_ ;
	assign \g16813/_0_  = _w23942_ ;
	assign \g16814/_0_  = _w23945_ ;
	assign \g16815/_0_  = _w23948_ ;
	assign \g16816/_0_  = _w23951_ ;
	assign \g16817/_0_  = _w23954_ ;
	assign \g16819/_0_  = _w23961_ ;
	assign \g16822/_0_  = _w23964_ ;
	assign \g16823/_0_  = _w23967_ ;
	assign \g16824/_0_  = _w23970_ ;
	assign \g16825/_0_  = _w23973_ ;
	assign \g16828/_0_  = _w23976_ ;
	assign \g16829/_0_  = _w23979_ ;
	assign \g16830/_0_  = _w23982_ ;
	assign \g16831/_0_  = _w23985_ ;
	assign \g16832/_0_  = _w23988_ ;
	assign \g16833/_0_  = _w23991_ ;
	assign \g16834/_0_  = _w23994_ ;
	assign \g16835/_0_  = _w23997_ ;
	assign \g16836/_0_  = _w24000_ ;
	assign \g16837/_0_  = _w24007_ ;
	assign \g16840/_0_  = _w24010_ ;
	assign \g16841/_0_  = _w24013_ ;
	assign \g16842/_0_  = _w24016_ ;
	assign \g16843/_0_  = _w24019_ ;
	assign \g16846/_0_  = _w24026_ ;
	assign \g16847/_0_  = _w24029_ ;
	assign \g16848/_0_  = _w24032_ ;
	assign \g16849/_0_  = _w24035_ ;
	assign \g16850/_0_  = _w24038_ ;
	assign \g16851/_0_  = _w24041_ ;
	assign \g16852/_0_  = _w24044_ ;
	assign \g16853/_0_  = _w24047_ ;
	assign \g16854/_0_  = _w24050_ ;
	assign \g16855/_0_  = _w24053_ ;
	assign \g16856/_0_  = _w24056_ ;
	assign \g16857/_0_  = _w24059_ ;
	assign \g16859/_0_  = _w24065_ ;
	assign \g16862/_0_  = _w24071_ ;
	assign \g16865/_0_  = _w24077_ ;
	assign \g16866/_0_  = _w24083_ ;
	assign \g16867/_0_  = _w24088_ ;
	assign \g16868/_0_  = _w24093_ ;
	assign \g16869/_0_  = _w24095_ ;
	assign \g16870/_0_  = _w24101_ ;
	assign \g16871/_0_  = _w24103_ ;
	assign \g16872/_0_  = _w24108_ ;
	assign \g16873/_0_  = _w24113_ ;
	assign \g16874/_0_  = _w24115_ ;
	assign \g16875/_0_  = _w24121_ ;
	assign \g16876/_0_  = _w24126_ ;
	assign \g16877/_0_  = _w24129_ ;
	assign \g16878/_0_  = _w24132_ ;
	assign \g16879/_0_  = _w24135_ ;
	assign \g16880/_0_  = _w24137_ ;
	assign \g16881/_0_  = _w24140_ ;
	assign \g16882/_0_  = _w24146_ ;
	assign \g16884/_0_  = _w24148_ ;
	assign \g16887/_0_  = _w24151_ ;
	assign \g16891/_0_  = _w24153_ ;
	assign \g16892/_0_  = _w24156_ ;
	assign \g16893/_0_  = _w24159_ ;
	assign \g16894/_0_  = _w24161_ ;
	assign \g16895/_0_  = _w24163_ ;
	assign \g16897/_0_  = _w24165_ ;
	assign \g16898/_0_  = _w24168_ ;
	assign \g16899/_0_  = _w24171_ ;
	assign \g16900/_0_  = _w24174_ ;
	assign \g16901/_0_  = _w24176_ ;
	assign \g16902/_0_  = _w24178_ ;
	assign \g16903/_0_  = _w24180_ ;
	assign \g16904/_0_  = _w24183_ ;
	assign \g16905/_0_  = _w24185_ ;
	assign \g16906/_0_  = _w24187_ ;
	assign \g16907/_0_  = _w24189_ ;
	assign \g16908/_0_  = _w24192_ ;
	assign \g16909/_0_  = _w24195_ ;
	assign \g16910/_0_  = _w24197_ ;
	assign \g16912/_0_  = _w24200_ ;
	assign \g16914/_0_  = _w24203_ ;
	assign \g16915/_0_  = _w24206_ ;
	assign \g16950/_0_  = _w24209_ ;
	assign \g16951/_0_  = _w24212_ ;
	assign \g16952/_0_  = _w24215_ ;
	assign \g16953/_0_  = _w24218_ ;
	assign \g16954/_0_  = _w24221_ ;
	assign \g16955/_0_  = _w24224_ ;
	assign \g16956/_0_  = _w24227_ ;
	assign \g16957/_0_  = _w24230_ ;
	assign \g16958/_0_  = _w24233_ ;
	assign \g16959/_0_  = _w24236_ ;
	assign \g16960/_0_  = _w24239_ ;
	assign \g16961/_0_  = _w24242_ ;
	assign \g16962/_0_  = _w24245_ ;
	assign \g16963/_0_  = _w24248_ ;
	assign \g16964/_0_  = _w24251_ ;
	assign \g16965/_0_  = _w24254_ ;
	assign \g16966/_0_  = _w24257_ ;
	assign \g16967/_0_  = _w24260_ ;
	assign \g16968/_0_  = _w24263_ ;
	assign \g16970/_0_  = _w24266_ ;
	assign \g17102/_3_  = _w24270_ ;
	assign \g17106/_0_  = _w24275_ ;
	assign \g17107/_0_  = _w24278_ ;
	assign \g17109/_0_  = _w24281_ ;
	assign \g17110/_0_  = _w24284_ ;
	assign \g17111/_0_  = _w24287_ ;
	assign \g17112/_0_  = _w24290_ ;
	assign \g17115/_0_  = _w24293_ ;
	assign \g17116/_0_  = _w24296_ ;
	assign \g17119/_0_  = _w24299_ ;
	assign \g17120/_0_  = _w24302_ ;
	assign \g17122/_0_  = _w24305_ ;
	assign \g17123/_0_  = _w24308_ ;
	assign \g17124/_0_  = _w24311_ ;
	assign \g17125/_0_  = _w24314_ ;
	assign \g17126/_0_  = _w24317_ ;
	assign \g17127/_0_  = _w24320_ ;
	assign \g17128/_0_  = _w24323_ ;
	assign \g17130/_0_  = _w24326_ ;
	assign \g17131/_0_  = _w24329_ ;
	assign \g17132/_0_  = _w24332_ ;
	assign \g17133/_0_  = _w24335_ ;
	assign \g17134/_0_  = _w24338_ ;
	assign \g17135/_0_  = _w24341_ ;
	assign \g17136/_0_  = _w24344_ ;
	assign \g17137/_0_  = _w24347_ ;
	assign \g17138/_0_  = _w24350_ ;
	assign \g17140/_0_  = _w24353_ ;
	assign \g17141/_0_  = _w24356_ ;
	assign \g17142/_0_  = _w24359_ ;
	assign \g17143/_0_  = _w24362_ ;
	assign \g17144/_0_  = _w24365_ ;
	assign \g17145/_0_  = _w24368_ ;
	assign \g17146/_0_  = _w24371_ ;
	assign \g17147/_0_  = _w24374_ ;
	assign \g17148/_0_  = _w24377_ ;
	assign \g17149/_0_  = _w24380_ ;
	assign \g17150/_0_  = _w24383_ ;
	assign \g17151/_0_  = _w24386_ ;
	assign \g17152/_0_  = _w24389_ ;
	assign \g17153/_0_  = _w24392_ ;
	assign \g17154/_0_  = _w24395_ ;
	assign \g17155/_0_  = _w24398_ ;
	assign \g17157/_0_  = _w24401_ ;
	assign \g17159/_0_  = _w24409_ ;
	assign \g17160/_0_  = _w24412_ ;
	assign \g17161/_0_  = _w24415_ ;
	assign \g17162/_0_  = _w24418_ ;
	assign \g17163/_0_  = _w24425_ ;
	assign \g17164/_0_  = _w24428_ ;
	assign \g17165/_0_  = _w24431_ ;
	assign \g17166/_0_  = _w24434_ ;
	assign \g17168/_0_  = _w24437_ ;
	assign \g17171/_0_  = _w24440_ ;
	assign \g17173/_0_  = _w24445_ ;
	assign \g17177/_0_  = _w24448_ ;
	assign \g17178/_0_  = _w24451_ ;
	assign \g17179/_0_  = _w24454_ ;
	assign \g17180/_0_  = _w24457_ ;
	assign \g17182/_0_  = _w24460_ ;
	assign \g17183/_0_  = _w24463_ ;
	assign \g17184/_0_  = _w24466_ ;
	assign \g17185/_0_  = _w24469_ ;
	assign \g17186/_0_  = _w24472_ ;
	assign \g17188/_0_  = _w24475_ ;
	assign \g17189/_0_  = _w24478_ ;
	assign \g17190/_0_  = _w24481_ ;
	assign \g17191/_0_  = _w24484_ ;
	assign \g17193/_0_  = _w24487_ ;
	assign \g17194/_0_  = _w24490_ ;
	assign \g17195/_0_  = _w24493_ ;
	assign \g17196/_0_  = _w24496_ ;
	assign \g17197/_0_  = _w24499_ ;
	assign \g17198/_0_  = _w24502_ ;
	assign \g17199/_0_  = _w24505_ ;
	assign \g17200/_0_  = _w24508_ ;
	assign \g17201/_0_  = _w24511_ ;
	assign \g17202/_0_  = _w24514_ ;
	assign \g17203/_0_  = _w24520_ ;
	assign \g17204/_0_  = _w24523_ ;
	assign \g17205/_0_  = _w24526_ ;
	assign \g17206/_0_  = _w24529_ ;
	assign \g17207/_0_  = _w24532_ ;
	assign \g17208/_0_  = _w24535_ ;
	assign \g17209/_0_  = _w24538_ ;
	assign \g17210/_0_  = _w24541_ ;
	assign \g17211/_0_  = _w24544_ ;
	assign \g17212/_0_  = _w24547_ ;
	assign \g17213/_0_  = _w24550_ ;
	assign \g17214/_0_  = _w24553_ ;
	assign \g17215/_0_  = _w24556_ ;
	assign \g17216/_0_  = _w24559_ ;
	assign \g17217/_0_  = _w24562_ ;
	assign \g17218/_0_  = _w24565_ ;
	assign \g17219/_0_  = _w24568_ ;
	assign \g17223/_0_  = _w24571_ ;
	assign \g17224/_0_  = _w24574_ ;
	assign \g17225/_0_  = _w24577_ ;
	assign \g17226/_0_  = _w24580_ ;
	assign \g17227/_0_  = _w24583_ ;
	assign \g17228/_0_  = _w24586_ ;
	assign \g17229/_0_  = _w24589_ ;
	assign \g17231/_0_  = _w24592_ ;
	assign \g17232/_0_  = _w24595_ ;
	assign \g17233/_0_  = _w24597_ ;
	assign \g17234/_0_  = _w24600_ ;
	assign \g17237/_0_  = _w24603_ ;
	assign \g17239/_0_  = _w24606_ ;
	assign \g17240/_0_  = _w24609_ ;
	assign \g17243/_0_  = _w24612_ ;
	assign \g17246/_0_  = _w24615_ ;
	assign \g17247/_0_  = _w24618_ ;
	assign \g17248/_0_  = _w24621_ ;
	assign \g17249/_0_  = _w24624_ ;
	assign \g17250/_0_  = _w24627_ ;
	assign \g17251/_0_  = _w24630_ ;
	assign \g17252/_0_  = _w24633_ ;
	assign \g17253/_0_  = _w24636_ ;
	assign \g17254/_0_  = _w24639_ ;
	assign \g17258/_0_  = _w24642_ ;
	assign \g17261/_0_  = _w24651_ ;
	assign \g17262/_0_  = _w24654_ ;
	assign \g17269/_0_  = _w24657_ ;
	assign \g17271/_0_  = _w24660_ ;
	assign \g17274/_0_  = _w24663_ ;
	assign \g17275/_0_  = _w24666_ ;
	assign \g17276/_0_  = _w24669_ ;
	assign \g17277/_0_  = _w24672_ ;
	assign \g17278/_0_  = _w24675_ ;
	assign \g17279/_0_  = _w24678_ ;
	assign \g17280/_0_  = _w24681_ ;
	assign \g17281/_0_  = _w24684_ ;
	assign \g17282/_0_  = _w24687_ ;
	assign \g17283/_0_  = _w24690_ ;
	assign \g17285/_0_  = _w24693_ ;
	assign \g17290/_0_  = _w24696_ ;
	assign \g17292/_0_  = _w24699_ ;
	assign \g17293/_0_  = _w24702_ ;
	assign \g17296/_0_  = _w24705_ ;
	assign \g17297/_0_  = _w24708_ ;
	assign \g17298/_0_  = _w24710_ ;
	assign \g173/_0_  = _w24721_ ;
	assign \g17303/_0_  = _w24724_ ;
	assign \g17304/_0_  = _w24727_ ;
	assign \g17305/_0_  = _w24730_ ;
	assign \g17306/_0_  = _w24733_ ;
	assign \g17307/_0_  = _w24736_ ;
	assign \g17308/_0_  = _w24739_ ;
	assign \g17309/_0_  = _w24742_ ;
	assign \g17310/_0_  = _w24745_ ;
	assign \g17311/_0_  = _w24748_ ;
	assign \g17312/_0_  = _w24751_ ;
	assign \g17314/_0_  = _w24754_ ;
	assign \g17315/_0_  = _w24757_ ;
	assign \g17316/_0_  = _w24760_ ;
	assign \g17317/_0_  = _w24763_ ;
	assign \g17318/_0_  = _w24766_ ;
	assign \g17319/_0_  = _w24769_ ;
	assign \g17320/_0_  = _w24772_ ;
	assign \g17321/_0_  = _w24775_ ;
	assign \g17322/_0_  = _w24778_ ;
	assign \g17323/_0_  = _w24781_ ;
	assign \g17324/_0_  = _w24784_ ;
	assign \g17325/_0_  = _w24787_ ;
	assign \g17326/_0_  = _w24790_ ;
	assign \g17327/_0_  = _w24793_ ;
	assign \g17328/_0_  = _w24796_ ;
	assign \g17329/_0_  = _w24799_ ;
	assign \g17330/_0_  = _w24802_ ;
	assign \g17331/_0_  = _w24805_ ;
	assign \g17332/_0_  = _w24808_ ;
	assign \g17333/_0_  = _w24811_ ;
	assign \g17335/_0_  = _w24814_ ;
	assign \g17336/_0_  = _w24818_ ;
	assign \g17337/_0_  = _w24821_ ;
	assign \g17338/_0_  = _w24824_ ;
	assign \g17339/_0_  = _w24827_ ;
	assign \g17340/_0_  = _w24830_ ;
	assign \g17342/_0_  = _w24833_ ;
	assign \g17343/_0_  = _w24836_ ;
	assign \g17347/_0_  = _w24839_ ;
	assign \g17350/_0_  = _w24842_ ;
	assign \g17354/_0_  = _w24845_ ;
	assign \g17356/_0_  = _w24848_ ;
	assign \g17357/_0_  = _w24851_ ;
	assign \g17358/_0_  = _w24854_ ;
	assign \g17359/_0_  = _w24857_ ;
	assign \g17360/_0_  = _w24860_ ;
	assign \g17415/_0_  = _w24863_ ;
	assign \g17441/_0_  = _w24865_ ;
	assign \g17442/_0_  = _w24867_ ;
	assign \g17451/_0_  = _w24869_ ;
	assign \g17457/_0_  = _w24873_ ;
	assign \g17458/_0_  = _w24876_ ;
	assign \g17459/_0_  = _w24879_ ;
	assign \g17460/_0_  = _w24882_ ;
	assign \g17461/_0_  = _w24885_ ;
	assign \g17462/_0_  = _w24888_ ;
	assign \g17463/_0_  = _w24891_ ;
	assign \g17464/_0_  = _w24894_ ;
	assign \g17465/_0_  = _w24897_ ;
	assign \g17466/_0_  = _w24900_ ;
	assign \g17467/_0_  = _w24903_ ;
	assign \g17468/_0_  = _w24906_ ;
	assign \g17469/_0_  = _w24909_ ;
	assign \g17470/_0_  = _w24912_ ;
	assign \g17471/_0_  = _w24915_ ;
	assign \g17472/_0_  = _w24918_ ;
	assign \g175/_3_  = _w24931_ ;
	assign \g1750/_0_  = _w24946_ ;
	assign \g176/_3_  = _w24965_ ;
	assign \g17619/_0_  = _w24967_ ;
	assign \g17620/_0_  = _w24968_ ;
	assign \g1763/_3_  = _w24978_ ;
	assign \g1764/_3_  = _w24984_ ;
	assign \g1768/_0_  = _w24990_ ;
	assign \g1769/_0_  = _w24993_ ;
	assign \g177/_3_  = _w25006_ ;
	assign \g17737/_0_  = _w25009_ ;
	assign \g17747/_0_  = _w25013_ ;
	assign \g178/_3_  = _w25019_ ;
	assign \g17814/_1_  = _w21314_ ;
	assign \g17815/_0_  = _w25023_ ;
	assign \g17821/_1_  = _w25024_ ;
	assign \g17821/_1__syn_2  = _w25024_ ;
	assign \g17872/_0_  = _w25026_ ;
	assign \g179/_3_  = _w25032_ ;
	assign \g17902/_0_  = _w25035_ ;
	assign \g180/_3_  = _w25041_ ;
	assign \g18020/_1_  = _w25043_ ;
	assign \g18057/_0_  = _w25045_ ;
	assign \g18096/_0_  = _w25049_ ;
	assign \g18099/_0_  = _w25052_ ;
	assign \g18107/_0_  = _w25055_ ;
	assign \g18133/_0_  = _w25059_ ;
	assign \g18140/_1_  = _w23021_ ;
	assign \g18153/_0_  = _w25062_ ;
	assign \g182/_0_  = _w25069_ ;
	assign \g18218/_0_  = _w25073_ ;
	assign \g18244/_0_  = _w25075_ ;
	assign \g18262/_0_  = _w25079_ ;
	assign \g18267/_0_  = _w25082_ ;
	assign \g18387/_1__syn_2  = _w25085_ ;
	assign \g184/_0_  = _w25088_ ;
	assign \g18478/_1_  = _w23343_ ;
	assign \g18585/_3_  = _w22290_ ;
	assign \g18608/_0_  = _w25092_ ;
	assign \g18609/_0_  = _w25096_ ;
	assign \g18613/_0_  = _w25101_ ;
	assign \g18618/_0_  = _w25105_ ;
	assign \g18647/_0_  = _w25109_ ;
	assign \g18687/_2_  = _w20990_ ;
	assign \g18707/_0_  = _w25113_ ;
	assign \g18748/_0_  = _w25117_ ;
	assign \g18753/_0_  = _w25121_ ;
	assign \g18758/_0_  = _w25124_ ;
	assign \g18759/_0_  = _w25128_ ;
	assign \g18760/_0_  = _w25131_ ;
	assign \g18761/_0_  = _w25135_ ;
	assign \g18762/_0_  = _w25138_ ;
	assign \g18763/_0_  = _w25141_ ;
	assign \g18764/_0_  = _w25144_ ;
	assign \g18765/_0_  = _w25147_ ;
	assign \g18766/_0_  = _w25150_ ;
	assign \g18767/_0_  = _w25153_ ;
	assign \g18768/_0_  = _w25156_ ;
	assign \g18770/_0_  = _w25159_ ;
	assign \g18771/_0_  = _w25162_ ;
	assign \g18788/_0_  = _w25165_ ;
	assign \g18796/_0_  = _w25168_ ;
	assign \g18800/_0_  = _w25171_ ;
	assign \g18801/_0_  = _w25174_ ;
	assign \g18802/_0_  = _w25177_ ;
	assign \g18803/_0_  = _w25180_ ;
	assign \g18804/_0_  = _w25183_ ;
	assign \g18805/_0_  = _w25186_ ;
	assign \g18807/_0_  = _w25189_ ;
	assign \g18840/_0_  = _w25196_ ;
	assign \g18843/_0_  = _w25199_ ;
	assign \g18844/_0_  = _w25205_ ;
	assign \g18846/_0_  = _w25210_ ;
	assign \g18847/_0_  = _w25216_ ;
	assign \g18848/_0_  = _w25220_ ;
	assign \g18849/_0_  = _w25224_ ;
	assign \g18850/_0_  = _w25228_ ;
	assign \g18851/_0_  = _w25231_ ;
	assign \g18852/_0_  = _w25234_ ;
	assign \g18853/_0_  = _w25237_ ;
	assign \g18854/_0_  = _w25243_ ;
	assign \g18855/_0_  = _w25247_ ;
	assign \g18856/_0_  = _w20720_ ;
	assign \g18858/_0_  = _w20709_ ;
	assign \g18860/_0_  = _w25251_ ;
	assign \g18861/_0_  = _w25254_ ;
	assign \g18863/_0_  = _w25257_ ;
	assign \g18864/_0_  = _w25260_ ;
	assign \g18866/_0_  = _w25263_ ;
	assign \g18867/_0_  = _w25266_ ;
	assign \g18868/_0_  = _w25269_ ;
	assign \g18869/_0_  = _w25272_ ;
	assign \g18870/_0_  = _w25275_ ;
	assign \g18871/_0_  = _w25278_ ;
	assign \g18872/_0_  = _w25281_ ;
	assign \g18873/_0_  = _w25284_ ;
	assign \g18874/_0_  = _w25287_ ;
	assign \g18875/_0_  = _w25290_ ;
	assign \g18876/_0_  = _w25293_ ;
	assign \g18877/_0_  = _w25296_ ;
	assign \g18878/_0_  = _w25299_ ;
	assign \g18879/_0_  = _w25302_ ;
	assign \g18880/_0_  = _w25305_ ;
	assign \g18881/_0_  = _w25308_ ;
	assign \g18882/_0_  = _w25311_ ;
	assign \g18883/_0_  = _w25314_ ;
	assign \g18888/_0_  = _w25318_ ;
	assign \g18892/_0_  = _w25324_ ;
	assign \g18895/_0_  = _w25330_ ;
	assign \g18896/_0_  = _w25336_ ;
	assign \g18897/_0_  = _w25339_ ;
	assign \g18905/_0_  = _w25343_ ;
	assign \g18908/_0_  = _w25346_ ;
	assign \g18909/_0_  = _w25349_ ;
	assign \g18912/_0_  = _w25352_ ;
	assign \g18918/_0_  = _w25356_ ;
	assign \g18919/_0_  = _w25360_ ;
	assign \g18920/_0_  = _w25363_ ;
	assign \g18921/_0_  = _w25369_ ;
	assign \g18922/_0_  = _w25372_ ;
	assign \g18924/_0_  = _w25378_ ;
	assign \g18925/_0_  = _w25381_ ;
	assign \g18927/_0_  = _w25384_ ;
	assign \g18930/_0_  = _w25387_ ;
	assign \g18966/_0_  = _w25393_ ;
	assign \g18968/_0_  = _w25399_ ;
	assign \g18970/_0_  = _w25402_ ;
	assign \g18974/_0_  = _w25405_ ;
	assign \g18975/_0_  = _w25411_ ;
	assign \g18977/_0_  = _w25417_ ;
	assign \g18981/_0_  = _w20757_ ;
	assign \g18983/_0_  = _w20604_ ;
	assign \g18985/_0_  = _w20616_ ;
	assign \g18987/_0_  = _w20626_ ;
	assign \g18989/_0_  = _w20636_ ;
	assign \g18991/_0_  = _w25421_ ;
	assign \g18992/_0_  = _w25427_ ;
	assign \g18993/_0_  = _w25433_ ;
	assign \g18994/_0_  = _w25436_ ;
	assign \g18995/_0_  = _w25442_ ;
	assign \g18996/_0_  = _w25445_ ;
	assign \g18997/_0_  = _w25451_ ;
	assign \g18998/_0_  = _w25454_ ;
	assign \g18999/_0_  = _w25457_ ;
	assign \g19001/_0_  = _w25460_ ;
	assign \g19003/_0_  = _w25463_ ;
	assign \g19005/_0_  = _w25466_ ;
	assign \g19006/_0_  = _w25472_ ;
	assign \g19014/_0_  = _w20646_ ;
	assign \g19016/_0_  = _w20654_ ;
	assign \g19018/_0_  = _w20665_ ;
	assign \g19020/_0_  = _w20676_ ;
	assign \g19022/_0_  = _w20731_ ;
	assign \g19056/_3_  = _w25476_ ;
	assign \g19058/_3_  = _w25480_ ;
	assign \g19060/_3_  = _w25484_ ;
	assign \g19062/_3_  = _w25488_ ;
	assign \g1910/_0_  = _w25502_ ;
	assign \g19186/_0_  = _w21380_ ;
	assign \g19188/_0_  = _w21388_ ;
	assign \g19235/_0_  = _w25506_ ;
	assign \g19239/_0_  = _w25509_ ;
	assign \g19244/_0_  = _w25512_ ;
	assign \g19253/_0_  = _w25515_ ;
	assign \g19254/_0_  = _w25518_ ;
	assign \g19259/_0_  = _w25521_ ;
	assign \g19261/_0_  = _w25524_ ;
	assign \g19267/_0_  = _w25527_ ;
	assign \g19277/_0_  = _w25531_ ;
	assign \g19278/_0_  = _w25534_ ;
	assign \g19280/_0_  = _w25538_ ;
	assign \g19281/_0_  = _w25541_ ;
	assign \g19282/_0_  = _w25544_ ;
	assign \g19283/_0_  = _w25547_ ;
	assign \g19284/_0_  = _w25550_ ;
	assign \g19285/_0_  = _w25553_ ;
	assign \g19286/_0_  = _w25556_ ;
	assign \g19287/_0_  = _w25559_ ;
	assign \g19288/_0_  = _w25562_ ;
	assign \g19289/_0_  = _w25565_ ;
	assign \g19290/_0_  = _w25568_ ;
	assign \g19291/_0_  = _w25571_ ;
	assign \g19292/_0_  = _w25574_ ;
	assign \g19293/_0_  = _w25577_ ;
	assign \g19294/_0_  = _w25580_ ;
	assign \g19295/_0_  = _w25583_ ;
	assign \g19296/_0_  = _w25586_ ;
	assign \g19297/_0_  = _w25589_ ;
	assign \g19298/_0_  = _w25592_ ;
	assign \g19299/_0_  = _w25595_ ;
	assign \g19300/_0_  = _w25598_ ;
	assign \g19301/_0_  = _w25601_ ;
	assign \g19302/_0_  = _w25604_ ;
	assign \g19303/_0_  = _w25607_ ;
	assign \g19304/_0_  = _w25610_ ;
	assign \g19305/_0_  = _w25613_ ;
	assign \g19306/_0_  = _w25616_ ;
	assign \g19307/_0_  = _w25619_ ;
	assign \g19308/_0_  = _w25622_ ;
	assign \g19315/_0_  = _w25625_ ;
	assign \g19316/_0_  = _w25628_ ;
	assign \g19317/_0_  = _w25631_ ;
	assign \g19318/_0_  = _w25634_ ;
	assign \g19319/_0_  = _w25637_ ;
	assign \g19320/_0_  = _w25640_ ;
	assign \g19321/_0_  = _w25643_ ;
	assign \g19322/_0_  = _w25646_ ;
	assign \g19323/_0_  = _w25649_ ;
	assign \g19325/_3_  = _w25654_ ;
	assign \g19326/_3_  = _w25659_ ;
	assign \g19333/_3_  = _w25664_ ;
	assign \g19341/_3_  = _w25669_ ;
	assign \g19347/_3_  = _w25674_ ;
	assign \g19377/_3_  = _w25677_ ;
	assign \g19381/_3_  = _w25682_ ;
	assign \g19393/_0_  = _w25687_ ;
	assign \g19401/_0_  = _w25693_ ;
	assign \g19402/_0_  = _w25699_ ;
	assign \g195/_2_  = _w13516_ ;
	assign \g19513/_0_  = _w25700_ ;
	assign \g19514/_0_  = _w25701_ ;
	assign \g19515/_0_  = _w25702_ ;
	assign \g19516/_0_  = _w25703_ ;
	assign \g1952/_3_  = _w25711_ ;
	assign \g19529/_0_  = _w25712_ ;
	assign \g19530/_0_  = _w25713_ ;
	assign \g19531/_0_  = _w25714_ ;
	assign \g19532/_0_  = _w25715_ ;
	assign \g19533/_0_  = _w25716_ ;
	assign \g19534/_0_  = _w25717_ ;
	assign \g19535/_0_  = _w25718_ ;
	assign \g19536/_0_  = _w25719_ ;
	assign \g19537/_0_  = _w25720_ ;
	assign \g19539/_0_  = _w25721_ ;
	assign \g19546/_0_  = _w25722_ ;
	assign \g19552/_0_  = _w25723_ ;
	assign \g19553/_0_  = _w25724_ ;
	assign \g19562/_0_  = _w25728_ ;
	assign \g19563/_0_  = _w25732_ ;
	assign \g19564/_0_  = _w25736_ ;
	assign \g19572/_0_  = _w19702_ ;
	assign \g19575/_0_  = _w25737_ ;
	assign \g19615/_0_  = _w25738_ ;
	assign \g19686/_0_  = _w25739_ ;
	assign \g19688/_0_  = _w25740_ ;
	assign \g197/_0_  = _w25792_ ;
	assign \g19729/_0_  = _w25796_ ;
	assign \g19774/_0_  = _w25800_ ;
	assign \g19777/_0_  = _w25804_ ;
	assign \g19791/_0_  = _w25808_ ;
	assign \g19818/_0_  = _w25810_ ;
	assign \g19819/_0_  = _w25811_ ;
	assign \g19828/_0_  = _w25815_ ;
	assign \g19852/_1_  = _w6067_ ;
	assign \g19860/_0_  = _w25819_ ;
	assign \g19861/_0_  = _w25823_ ;
	assign \g19864/_0_  = _w25827_ ;
	assign \g19886/_0_  = _w25828_ ;
	assign \g19887/_0_  = _w25830_ ;
	assign \g199/_0_  = _w25849_ ;
	assign \g19908/_0_  = _w25850_ ;
	assign \g19918/_0_  = _w25854_ ;
	assign \g19927/_0_  = _w25858_ ;
	assign \g19933/_0_  = _w25862_ ;
	assign \g200/_0_  = _w22959_ ;
	assign \g20019/_0_  = _w25866_ ;
	assign \g20046/_0_  = _w25870_ ;
	assign \g20068/_1_  = _w23958_ ;
	assign \g20080/_1_  = _w24004_ ;
	assign \g201/_0_  = _w25900_ ;
	assign \g20137/_0_  = _w25904_ ;
	assign \g20139/_0_  = _w25909_ ;
	assign \g20141/_0_  = _w25913_ ;
	assign \g20152/_1_  = _w6075_ ;
	assign \g20154/_00_  = _w25918_ ;
	assign \g202/_0_  = _w25948_ ;
	assign \g20206/_0_  = _w25953_ ;
	assign \g20211/_2_  = _w25954_ ;
	assign \g20217/_2_  = _w25955_ ;
	assign \g20239/_0_  = _w25958_ ;
	assign \g20265/_2_  = _w25959_ ;
	assign \g20266/_0_  = _w25961_ ;
	assign \g20272/_2_  = _w25964_ ;
	assign \g20278/_2_  = _w25965_ ;
	assign \g20283/_0_  = _w18519_ ;
	assign \g20285/_2_  = _w25968_ ;
	assign \g20288/_2__syn_2  = _w23336_ ;
	assign \g20293/_0_  = _w25972_ ;
	assign \g20295/_2_  = _w20870_ ;
	assign \g203/_0_  = _w22999_ ;
	assign \g20302/_2_  = _w25973_ ;
	assign \g20303/_2_  = _w25974_ ;
	assign \g20304/_2_  = _w25975_ ;
	assign \g20311/_2_  = _w25976_ ;
	assign \g20326/_0_  = _w25980_ ;
	assign \g20330/_0_  = _w25982_ ;
	assign \g2034/_0_  = _w25988_ ;
	assign \g20345/_0_  = _w25992_ ;
	assign \g20346/_0_  = _w25995_ ;
	assign \g2035/_0_  = _w25998_ ;
	assign \g20363/_0_  = _w21241_ ;
	assign \g20364/_0_  = _w26002_ ;
	assign \g204/_0_  = _w26021_ ;
	assign \g2047/_0_  = _w26026_ ;
	assign \g20483/_0_  = _w26029_ ;
	assign \g20493/_00_  = _w26034_ ;
	assign \g205/_0_  = _w26040_ ;
	assign \g20569/_0_  = _w26042_ ;
	assign \g20570/_0_  = _w26044_ ;
	assign \g20571/_0_  = _w26046_ ;
	assign \g206/_0_  = _w26049_ ;
	assign \g20613/_0_  = _w26050_ ;
	assign \g20615/_0_  = _w26051_ ;
	assign \g20657/_1__syn_2  = _w26052_ ;
	assign \g20660/_0_  = _w26053_ ;
	assign \g20685/_0_  = _w26055_ ;
	assign \g207/_0_  = _w26058_ ;
	assign \g20713/_1_  = _w26059_ ;
	assign \g20747/_1_  = _w26060_ ;
	assign \g20784/_0_  = _w23018_ ;
	assign \g20820/_1_  = _w25042_ ;
	assign \g20859/_0_  = _w26063_ ;
	assign \g20873/_2_  = _w26065_ ;
	assign \g20886/_0_  = _w26066_ ;
	assign \g20887/_0_  = _w26067_ ;
	assign \g20891/_2__syn_2  = _w25666_ ;
	assign \g20907/_2_  = _w25071_ ;
	assign \g20936/_2__syn_2  = _w25661_ ;
	assign \g20937/_1_  = _w26068_ ;
	assign \g20955/_0_  = _w26070_ ;
	assign \g20959/_2__syn_2  = _w25656_ ;
	assign \g20967/_0_  = _w26071_ ;
	assign \g20971/_2__syn_2  = _w25679_ ;
	assign \g20974/_1__syn_2  = _w25684_ ;
	assign \g21015/_1_  = _w26073_ ;
	assign \g21051/_2_  = _w25057_ ;
	assign \g21079/_1_  = _w26074_ ;
	assign \g21081/_1_  = _w26075_ ;
	assign \g21087/_2__syn_2  = _w25671_ ;
	assign \g21114/_1_  = _w26076_ ;
	assign \g21116/_1_  = _w26077_ ;
	assign \g21120/_2__syn_2  = _w25651_ ;
	assign \g21147/_0_  = _w26078_ ;
	assign \g21179/_1_  = _w26079_ ;
	assign \g21185/_1_  = _w26080_ ;
	assign \g21223/_0_  = _w26082_ ;
	assign \g21242/_0_  = _w26084_ ;
	assign \g21253/_0_  = _w26085_ ;
	assign \g21257/_0_  = _w26087_ ;
	assign \g21323/_1_  = _w26089_ ;
	assign \g21324/_1_  = _w26090_ ;
	assign \g21366/_0_  = _w26092_ ;
	assign \g21385/_2_  = _w26094_ ;
	assign \g21464/_0_  = _w26096_ ;
	assign \g21475/_3_  = _w26099_ ;
	assign \g21481/_0_  = _w26102_ ;
	assign \g21482/_0_  = _w26104_ ;
	assign \g21494/_3_  = _w26107_ ;
	assign \g21500/_3_  = _w26110_ ;
	assign \g21507/_3_  = _w26113_ ;
	assign \g21511/_3_  = _w26116_ ;
	assign \g21537/_1_  = _w26119_ ;
	assign \g21568/_0_  = _w26122_ ;
	assign \g21591/_0_  = _w26125_ ;
	assign \g21604/_0_  = _w26129_ ;
	assign \g21605/_3_  = _w20602_ ;
	assign \g21606/_0_  = _w26132_ ;
	assign \g21607/_0_  = _w26135_ ;
	assign \g21608/_0_  = _w26138_ ;
	assign \g21609/_0_  = _w26141_ ;
	assign \g21610/_0_  = _w26144_ ;
	assign \g21611/_0_  = _w26147_ ;
	assign \g21612/_0_  = _w26150_ ;
	assign \g21613/_0_  = _w26153_ ;
	assign \g21614/_0_  = _w26156_ ;
	assign \g21615/_0_  = _w26159_ ;
	assign \g21616/_0_  = _w26162_ ;
	assign \g21617/_0_  = _w26165_ ;
	assign \g21618/_0_  = _w26168_ ;
	assign \g21621/_0_  = _w26170_ ;
	assign \g21640/_0_  = _w26173_ ;
	assign \g21678/_0_  = _w26176_ ;
	assign \g21679/_0_  = _w26179_ ;
	assign \g21686/_0_  = _w26182_ ;
	assign \g21692/_3_  = _w24098_ ;
	assign \g21696/_0_  = _w26185_ ;
	assign \g21698/_0_  = _w26188_ ;
	assign \g21702/_3_  = _w20718_ ;
	assign \g21707/_0_  = _w26191_ ;
	assign \g21709/_0_  = _w26194_ ;
	assign \g21728/_0_  = _w26197_ ;
	assign \g21729/_0_  = _w26200_ ;
	assign \g21731/_0_  = _w26203_ ;
	assign \g21732/_0_  = _w26206_ ;
	assign \g21733/_0_  = _w26209_ ;
	assign \g21736/_0_  = _w26212_ ;
	assign \g21744/_3_  = _w20707_ ;
	assign \g21753/_0_  = _w26215_ ;
	assign \g21754/_0_  = _w26218_ ;
	assign \g21755/_0_  = _w26221_ ;
	assign \g21756/_0_  = _w26224_ ;
	assign \g21757/_0_  = _w26227_ ;
	assign \g21759/_0_  = _w26230_ ;
	assign \g21761/_0_  = _w26233_ ;
	assign \g21763/_0_  = _w26236_ ;
	assign \g21764/_0_  = _w26239_ ;
	assign \g21766/_0_  = _w26242_ ;
	assign \g2180/_0_  = _w26259_ ;
	assign \g21853/_3_  = _w23886_ ;
	assign \g21861/_3_  = _w24111_ ;
	assign \g21863/_3_  = _w24118_ ;
	assign \g21869/_3_  = _w20614_ ;
	assign \g2187/_0_  = _w26281_ ;
	assign \g21875/_3_  = _w24124_ ;
	assign \g21877/_3_  = _w24143_ ;
	assign \g21879/_3_  = _w24106_ ;
	assign \g2188/_0_  = _w26284_ ;
	assign \g21900/_0_  = _w26286_ ;
	assign \g22080/_0_  = _w26287_ ;
	assign \g22082/_0_  = _w26288_ ;
	assign \g22135/_0_  = _w26289_ ;
	assign \g22145/_1_  = _w26290_ ;
	assign \g22225/_0_  = _w26291_ ;
	assign \g223/_0_  = _w25004_ ;
	assign \g22354/_0_  = _w26292_ ;
	assign \g224/_0_  = _w24929_ ;
	assign \g22412/_0_  = _w26302_ ;
	assign \g22415/_1__syn_2  = _w23020_ ;
	assign \g225/_0_  = _w24963_ ;
	assign \g2257/_0_  = _w5560_ ;
	assign \g226/_3_  = _w26319_ ;
	assign \g22624/_0_  = _w26320_ ;
	assign \g227/_3_  = _w26326_ ;
	assign \g22702/_0_  = _w26327_ ;
	assign \g22919/_1__syn_2  = _w25989_ ;
	assign \g22933/_0_  = _w26334_ ;
	assign \g22954/_0_  = _w26337_ ;
	assign \g22989/_1_  = _w26338_ ;
	assign \g23529/_0_  = \T_IRQE1n_pad ;
	assign \g23539/_0_  = \T_IRQ2n_pad ;
	assign \g2362/_2_  = _w26396_ ;
	assign \g23766/_0_  = T_PWDn_pad;
	assign \g24/_3_  = _w26399_ ;
	assign \g24018/_0_  = \T_IRQ0n_pad ;
	assign \g2416/_0_  = _w26962_ ;
	assign \g2420/_0_  = _w26966_ ;
	assign \g24213/_0_  = \T_IRQL1n_pad ;
	assign \g24301/_0_  = \T_IRQ1n_pad ;
	assign \g2479/_0_  = _w27036_ ;
	assign \g248/_3_  = _w27055_ ;
	assign \g2480/_0_  = _w27083_ ;
	assign \g2481/_0_  = _w27111_ ;
	assign \g2482/_0_  = _w27139_ ;
	assign \g2483/_0_  = _w27167_ ;
	assign \g2484/_0_  = _w27195_ ;
	assign \g2485/_0_  = _w27223_ ;
	assign \g2486/_0_  = _w27251_ ;
	assign \g2487/_0_  = _w27279_ ;
	assign \g2488/_0_  = _w27307_ ;
	assign \g249/_3_  = _w27313_ ;
	assign \g2490/_0_  = _w27341_ ;
	assign \g2491/_0_  = _w27369_ ;
	assign \g2492/_0_  = _w27397_ ;
	assign \g2493/_0_  = _w27425_ ;
	assign \g2494/_0_  = _w27453_ ;
	assign \g2495/_0_  = _w27481_ ;
	assign \g2496/_0_  = _w27493_ ;
	assign \g2497/_0_  = _w27496_ ;
	assign \g2507/_0_  = _w27506_ ;
	assign \g2508/_0_  = _w27515_ ;
	assign \g2509/_0_  = _w27524_ ;
	assign \g2510/_0_  = _w27533_ ;
	assign \g2511/_0_  = _w27542_ ;
	assign \g2512/_0_  = _w27551_ ;
	assign \g2513/_0_  = _w27560_ ;
	assign \g2514/_0_  = _w27586_ ;
	assign \g2515/_0_  = _w27612_ ;
	assign \g2516/_0_  = _w27621_ ;
	assign \g25237/_0_  = \T_IRQE0n_pad ;
	assign \g2558/_0_  = _w27626_ ;
	assign \g2562/_0_  = _w27652_ ;
	assign \g2563/_0_  = _w27678_ ;
	assign \g2564/_0_  = _w27704_ ;
	assign \g2565/_0_  = _w27730_ ;
	assign \g2566/_0_  = _w27756_ ;
	assign \g2567/_0_  = _w27782_ ;
	assign \g2699/_0_  = _w26394_ ;
	assign \g27/_2_  = _w27786_ ;
	assign \g271/_0_  = _w26317_ ;
	assign \g272/_3_  = _w27805_ ;
	assign \g273/_3_  = _w27818_ ;
	assign \g274/_3_  = _w27824_ ;
	assign \g275/_3_  = _w27830_ ;
	assign \g276/_3_  = _w27840_ ;
	assign \g277/_3_  = _w27846_ ;
	assign \g2787/_3_  = _w27856_ ;
	assign \g2788/_3_  = _w27862_ ;
	assign \g279/_0_  = _w27872_ ;
	assign \g2795/_0_  = _w27878_ ;
	assign \g2796/_0_  = _w27881_ ;
	assign \g280/_0_  = _w27887_ ;
	assign \g2842/_3_  = _w27902_ ;
	assign \g29/_1_  = _w27904_ ;
	assign \g2927/_0_  = _w28157_ ;
	assign \g2978/_0_  = _w28167_ ;
	assign \g2979/_0_  = _w28172_ ;
	assign \g2980/_0_  = _w28177_ ;
	assign \g2981/_0_  = _w28182_ ;
	assign \g2982/_0_  = _w28187_ ;
	assign \g2983/_0_  = _w28192_ ;
	assign \g2984/_0_  = _w28197_ ;
	assign \g2985/_0_  = _w28202_ ;
	assign \g3021/_3_  = _w28210_ ;
	assign \g3022/_3_  = _w28216_ ;
	assign \g3023/_3_  = _w28222_ ;
	assign \g3024/_3_  = _w28228_ ;
	assign \g3025/_3_  = _w28234_ ;
	assign \g3026/_3_  = _w28240_ ;
	assign \g3027/_3_  = _w28246_ ;
	assign \g3028/_3_  = _w28252_ ;
	assign \g3029/_3_  = _w28261_ ;
	assign \g3030/_3_  = _w28270_ ;
	assign \g3031/_3_  = _w28279_ ;
	assign \g3032/_3_  = _w28288_ ;
	assign \g3033/_3_  = _w28297_ ;
	assign \g3034/_3_  = _w28306_ ;
	assign \g3035/_3_  = _w28315_ ;
	assign \g3036/_3_  = _w28324_ ;
	assign \g3037/_3_  = _w28330_ ;
	assign \g3038/_3_  = _w28336_ ;
	assign \g3039/_3_  = _w28342_ ;
	assign \g3040/_3_  = _w28348_ ;
	assign \g3041/_3_  = _w28354_ ;
	assign \g3042/_3_  = _w28360_ ;
	assign \g3049/_0_  = _w28363_ ;
	assign \g3050/_0_  = _w28366_ ;
	assign \g3051/_0_  = _w28369_ ;
	assign \g3052/_0_  = _w28372_ ;
	assign \g3053/_0_  = _w28375_ ;
	assign \g3054/_0_  = _w28378_ ;
	assign \g3058/_0_  = _w28381_ ;
	assign \g3059/_0_  = _w28384_ ;
	assign \g3088/_0_  = _w28393_ ;
	assign \g3089/_0_  = _w28401_ ;
	assign \g3090/_0_  = _w28409_ ;
	assign \g3091/_0_  = _w28417_ ;
	assign \g3092/_0_  = _w28425_ ;
	assign \g3093/_0_  = _w28433_ ;
	assign \g3094/_0_  = _w28441_ ;
	assign \g3095/_0_  = _w28449_ ;
	assign \g314/_0_  = _w27053_ ;
	assign \g3147/_3_  = _w28455_ ;
	assign \g3148/_3_  = _w28461_ ;
	assign \g3189/_0_  = _w28467_ ;
	assign \g3190/_0_  = _w28473_ ;
	assign \g3191/_0_  = _w28479_ ;
	assign \g3192/_0_  = _w28485_ ;
	assign \g3193/_0_  = _w28491_ ;
	assign \g3194/_0_  = _w28497_ ;
	assign \g3195/_0_  = _w28503_ ;
	assign \g3196/_0_  = _w28509_ ;
	assign \g3197/_0_  = _w28515_ ;
	assign \g3198/_0_  = _w28521_ ;
	assign \g3199/_0_  = _w28527_ ;
	assign \g32/_0_  = _w28542_ ;
	assign \g320/_3_  = _w28669_ ;
	assign \g3200/_0_  = _w28675_ ;
	assign \g3201/_0_  = _w28681_ ;
	assign \g3202/_0_  = _w28687_ ;
	assign \g3203/_0_  = _w28693_ ;
	assign \g3204/_0_  = _w28699_ ;
	assign \g321/_3_  = _w28755_ ;
	assign \g325/_3_  = _w28763_ ;
	assign \g3271/_2_  = _w26388_ ;
	assign \g33/_0_  = _w28773_ ;
	assign \g3363/_0_  = _w28785_ ;
	assign \g3413/_0_  = _w28875_ ;
	assign \g3414/_0_  = _w28965_ ;
	assign \g352/_0_  = _w27803_ ;
	assign \g355/_0_  = _w27816_ ;
	assign \g356/_3_  = _w28975_ ;
	assign \g357/_3_  = _w28981_ ;
	assign \g35_dup/_1_  = _w28982_ ;
	assign \g36/_3_  = _w28985_ ;
	assign \g365/_3_  = _w29038_ ;
	assign \g366/_3_  = _w29127_ ;
	assign \g367/_3_  = _w29178_ ;
	assign \g368/_3_  = _w29227_ ;
	assign \g3687/_0_  = _w29232_ ;
	assign \g369/_3_  = _w29340_ ;
	assign \g37/_3_  = _w29343_ ;
	assign \g370/_3_  = _w29364_ ;
	assign \g372/_3_  = _w29385_ ;
	assign \g374/_3_  = _w29406_ ;
	assign \g3740/_0_  = _w29411_ ;
	assign \g375/_3_  = _w29432_ ;
	assign \g376/_3_  = _w29453_ ;
	assign \g3878/_0_  = _w29461_ ;
	assign \g3879/_0_  = _w29466_ ;
	assign \g388/_3_  = _w29476_ ;
	assign \g3880/_0_  = _w29485_ ;
	assign \g3881/_0_  = _w29490_ ;
	assign \g3882/_0_  = _w29498_ ;
	assign \g389/_3_  = _w29504_ ;
	assign \g3894/_0_  = _w29507_ ;
	assign \g3895/_0_  = _w29510_ ;
	assign \g3896/_0_  = _w29513_ ;
	assign \g3897/_0_  = _w29516_ ;
	assign \g3898/_0_  = _w29519_ ;
	assign \g392/_3_  = _w29669_ ;
	assign \g393/_3_  = _w29731_ ;
	assign \g394/_3_  = _w29882_ ;
	assign \g395/_3_  = _w29987_ ;
	assign \g396/_3_  = _w29995_ ;
	assign \g397/_3_  = _w30003_ ;
	assign \g398/_3_  = _w30011_ ;
	assign \g399/_3_  = _w30019_ ;
	assign \g401/_3_  = _w30155_ ;
	assign \g402/_3_  = _w30163_ ;
	assign \g404/_3_  = _w30261_ ;
	assign \g4048/_0_  = _w30266_ ;
	assign \g405/_3_  = _w30324_ ;
	assign \g4050/_0_  = _w30329_ ;
	assign \g406/_3_  = _w30337_ ;
	assign \g407/_3_  = _w30345_ ;
	assign \g410/_3_  = _w30485_ ;
	assign \g411/_3_  = _w30493_ ;
	assign \g412/_3_  = _w30542_ ;
	assign \g413/_3_  = _w30647_ ;
	assign \g415/_3_  = _w30668_ ;
	assign \g416/_3_  = _w30689_ ;
	assign \g42/_0_  = _w30699_ ;
	assign \g4216/_3_  = _w30709_ ;
	assign \g4217/_3_  = _w30718_ ;
	assign \g4218/_3_  = _w30726_ ;
	assign \g4219/_3_  = _w30740_ ;
	assign \g4296/_0_  = _w30764_ ;
	assign \g4297/_0_  = _w30788_ ;
	assign \g4298/_0_  = _w30792_ ;
	assign \g4299/_0_  = _w30796_ ;
	assign \g43/_0_  = _w30804_ ;
	assign \g4300/_0_  = _w30808_ ;
	assign \g4301/_0_  = _w30812_ ;
	assign \g4302/_0_  = _w30816_ ;
	assign \g4303/_0_  = _w30820_ ;
	assign \g4304/_0_  = _w30824_ ;
	assign \g4305/_0_  = _w30828_ ;
	assign \g4306/_0_  = _w30832_ ;
	assign \g4307/_0_  = _w30836_ ;
	assign \g4308/_0_  = _w30840_ ;
	assign \g4309/_0_  = _w30844_ ;
	assign \g4310/_0_  = _w30848_ ;
	assign \g4311/_0_  = _w30852_ ;
	assign \g4312/_0_  = _w30856_ ;
	assign \g4313/_0_  = _w30860_ ;
	assign \g4314/_0_  = _w30864_ ;
	assign \g4315/_0_  = _w30868_ ;
	assign \g4316/_0_  = _w30872_ ;
	assign \g4317/_0_  = _w30876_ ;
	assign \g4318/_0_  = _w30880_ ;
	assign \g4319/_0_  = _w30884_ ;
	assign \g4320/_0_  = _w30888_ ;
	assign \g4321/_0_  = _w30892_ ;
	assign \g4322/_0_  = _w30896_ ;
	assign \g4323/_0_  = _w30900_ ;
	assign \g436/_0_  = _w30904_ ;
	assign \g44/_0_  = _w30914_ ;
	assign \g448/_3_  = _w30922_ ;
	assign \g45/_0_  = _w30932_ ;
	assign \g4587/_0_  = _w30989_ ;
	assign \g4588/_0_  = _w30992_ ;
	assign \g46/_0_  = _w17796_ ;
	assign \g4601/_0_  = _w30997_ ;
	assign \g4602/_0_  = _w31002_ ;
	assign \g4613/_3_  = _w31010_ ;
	assign \g4614/_3_  = _w31019_ ;
	assign \g4615/_3_  = _w31027_ ;
	assign \g463/_0_  = _w31062_ ;
	assign \g465/_0_  = _w31067_ ;
	assign \g4653/_0_  = _w31109_ ;
	assign \g4654/_0_  = _w31118_ ;
	assign \g4655/_0_  = _w31125_ ;
	assign \g4656/_0_  = _w31130_ ;
	assign \g4659/_0_  = _w31133_ ;
	assign \g466/_0_  = _w31137_ ;
	assign \g468/_3_  = _w31147_ ;
	assign \g469/_3_  = _w31153_ ;
	assign \g4697/_0_  = _w31158_ ;
	assign \g47/_3_  = _w31168_ ;
	assign \g470/_0_  = _w31183_ ;
	assign \g471/_0_  = _w31186_ ;
	assign \g4755/_0_  = _w31189_ ;
	assign \g476/_0_  = _w31226_ ;
	assign \g48/_3_  = _w31232_ ;
	assign \g480/_00_  = _w31256_ ;
	assign \g4839/_0_  = _w31276_ ;
	assign \g4840/_0_  = _w31279_ ;
	assign \g485/_3_  = _w31282_ ;
	assign \g4854/_0_  = _w31287_ ;
	assign \g4855/_0_  = _w31292_ ;
	assign \g4859/_0_  = _w31297_ ;
	assign \g486/_3_  = _w31300_ ;
	assign \g4860/_0_  = _w31305_ ;
	assign \g4880/_0_  = _w31353_ ;
	assign \g4881/_0_  = _w31365_ ;
	assign \g4882/_0_  = _w31377_ ;
	assign \g4883/_0_  = _w31389_ ;
	assign \g4884/_0_  = _w31423_ ;
	assign \g4885/_0_  = _w31435_ ;
	assign \g4886/_0_  = _w31447_ ;
	assign \g4887/_0_  = _w31459_ ;
	assign \g4888/_0_  = _w31471_ ;
	assign \g49/_0_  = _w31484_ ;
	assign \g494/_0_  = _w5673_ ;
	assign \g499/_1_  = _w5642_ ;
	assign \g50/_0_  = _w31490_ ;
	assign \g5002/_0_  = _w31534_ ;
	assign \g5003/_0_  = _w31543_ ;
	assign \g5009/_0_  = _w31551_ ;
	assign \g5010/_0_  = _w31558_ ;
	assign \g5011/_0_  = _w31568_ ;
	assign \g5014/_0_  = _w31571_ ;
	assign \g51/_0_  = _w31574_ ;
	assign \g5105/_0_  = _w31577_ ;
	assign \g5129/_2_  = _w31585_ ;
	assign \g5132/_0_  = _w31615_ ;
	assign \g5135/_0_  = _w31645_ ;
	assign \g5168/_0_  = _w31662_ ;
	assign \g5169/_0_  = _w31665_ ;
	assign \g5173/_0_  = _w31670_ ;
	assign \g5224/_0_  = _w31675_ ;
	assign \g5225/_0_  = _w31680_ ;
	assign \g5226/_0_  = _w31685_ ;
	assign \g5227/_0_  = _w31690_ ;
	assign \g5334/_0_  = _w31709_ ;
	assign \g5335/_0_  = _w31715_ ;
	assign \g5336/_0_  = _w31721_ ;
	assign \g5337/_0_  = _w31725_ ;
	assign \g5338/_0_  = _w31734_ ;
	assign \g5339/_0_  = _w31743_ ;
	assign \g5340/_0_  = _w31752_ ;
	assign \g5341/_0_  = _w31761_ ;
	assign \g5342/_0_  = _w31770_ ;
	assign \g5343/_0_  = _w31779_ ;
	assign \g5344/_0_  = _w31788_ ;
	assign \g5345/_0_  = _w31797_ ;
	assign \g5346/_0_  = _w31806_ ;
	assign \g5347/_0_  = _w31815_ ;
	assign \g5348/_0_  = _w31824_ ;
	assign \g5349/_0_  = _w31833_ ;
	assign \g5395/_0_  = _w31836_ ;
	assign \g54/_0_  = _w31839_ ;
	assign \g5434/_0_  = _w31849_ ;
	assign \g5447/_0_  = _w31855_ ;
	assign \g5450/_0_  = _w31874_ ;
	assign \g5451/_0_  = _w31880_ ;
	assign \g5452/_0_  = _w31886_ ;
	assign \g5453/_0_  = _w31892_ ;
	assign \g5454/_0_  = _w31896_ ;
	assign \g5461/_0_  = _w31899_ ;
	assign \g5483/_0_  = _w31907_ ;
	assign \g5484/_0_  = _w31929_ ;
	assign \g5492/_0_  = _w31932_ ;
	assign \g5493/_0_  = _w31938_ ;
	assign \g5496/_3_  = _w31948_ ;
	assign \g5497/_3_  = _w31954_ ;
	assign \g55/_0_  = _w31957_ ;
	assign \g5500/_0_  = _w31964_ ;
	assign \g5502/_0_  = _w31988_ ;
	assign \g5503/_0_  = _w32034_ ;
	assign \g5506/_0_  = _w32044_ ;
	assign \g5511/_0_  = _w32093_ ;
	assign \g5518/_0_  = _w32105_ ;
	assign \g5519/_0_  = _w32117_ ;
	assign \g5520/_0_  = _w32129_ ;
	assign \g5522/_0_  = _w32141_ ;
	assign \g5523/_0_  = _w32153_ ;
	assign \g5524/_0_  = _w32165_ ;
	assign \g5525/_0_  = _w32177_ ;
	assign \g5532/_0_  = _w32182_ ;
	assign \g5533/_0_  = _w32187_ ;
	assign \g5534/_0_  = _w32192_ ;
	assign \g5535/_0_  = _w32197_ ;
	assign \g5536/_0_  = _w32203_ ;
	assign \g5537/_0_  = _w32209_ ;
	assign \g5538/_0_  = _w32215_ ;
	assign \g5546/_0_  = _w32223_ ;
	assign \g5555/_00_  = _w32251_ ;
	assign \g5593/_0_  = _w4148_ ;
	assign \g5614/_2_  = _w6929_ ;
	assign \g567/_0_  = _w32255_ ;
	assign \g5677/_0_  = _w32258_ ;
	assign \g5678/_0_  = _w32261_ ;
	assign \g5682/_0_  = _w32265_ ;
	assign \g5683/_0_  = _w32270_ ;
	assign \g5684/_0_  = _w32274_ ;
	assign \g5686/_0_  = _w32280_ ;
	assign \g5687/_0_  = _w32284_ ;
	assign \g5689/_0_  = _w32289_ ;
	assign \g5690/_0_  = _w32293_ ;
	assign \g5691/_0_  = _w32298_ ;
	assign \g5692/_0_  = _w32302_ ;
	assign \g5698/_0_  = _w32305_ ;
	assign \g5699/_0_  = _w32308_ ;
	assign \g5700/_0_  = _w32312_ ;
	assign \g5701/_0_  = _w32315_ ;
	assign \g5702/_0_  = _w32318_ ;
	assign \g5703/_0_  = _w32319_ ;
	assign \g5704/_0_  = _w32335_ ;
	assign \g5709/_0_  = _w32338_ ;
	assign \g5711/_0_  = _w32341_ ;
	assign \g5714/_0_  = _w32342_ ;
	assign \g572/_0_  = _w32348_ ;
	assign \g5723/_0_  = _w32356_ ;
	assign \g5724/_0_  = _w32363_ ;
	assign \g5725/_0_  = _w32390_ ;
	assign \g573/_0_  = _w32393_ ;
	assign \g5739/_0_  = _w32409_ ;
	assign \g5740/_0_  = _w32419_ ;
	assign \g575/_0_  = _w32422_ ;
	assign \g5756/_0_  = _w32425_ ;
	assign \g5757/_0_  = _w32428_ ;
	assign \g5758/_0_  = _w32431_ ;
	assign \g5759/_0_  = _w32434_ ;
	assign \g576/_0_  = _w32437_ ;
	assign \g5760/_0_  = _w32440_ ;
	assign \g5761/_0_  = _w32443_ ;
	assign \g5762/_0_  = _w32446_ ;
	assign \g5763/_0_  = _w32449_ ;
	assign \g577/_0_  = _w32452_ ;
	assign \g5772/_0_  = _w32480_ ;
	assign \g5773/_0_  = _w32489_ ;
	assign \g5774/_0_  = _w32501_ ;
	assign \g5775/_0_  = _w32509_ ;
	assign \g5776/_0_  = _w32517_ ;
	assign \g5777/_0_  = _w32525_ ;
	assign \g578/_0_  = _w32528_ ;
	assign \g5781/_0_  = _w32538_ ;
	assign \g5783/_0_  = _w32546_ ;
	assign \g5784/_0_  = _w32554_ ;
	assign \g5785/_0_  = _w32562_ ;
	assign \g5786/_0_  = _w32570_ ;
	assign \g5787/_0_  = _w32578_ ;
	assign \g5788/_0_  = _w32586_ ;
	assign \g5789/_0_  = _w32594_ ;
	assign \g579/_0_  = _w32597_ ;
	assign \g5790/_0_  = _w32600_ ;
	assign \g5791/_0_  = _w32603_ ;
	assign \g5792/_0_  = _w32605_ ;
	assign \g5794/_0_  = _w32622_ ;
	assign \g5795/_0_  = _w32625_ ;
	assign \g5796/_0_  = _w32628_ ;
	assign \g580/_0_  = _w32631_ ;
	assign \g5801/_0_  = _w32634_ ;
	assign \g5802/_0_  = _w32637_ ;
	assign \g5803/_0_  = _w32641_ ;
	assign \g5804/_0_  = _w32645_ ;
	assign \g5805/_0_  = _w32648_ ;
	assign \g581/_0_  = _w32651_ ;
	assign \g5814/_0_  = _w32668_ ;
	assign \g582/_0_  = _w32671_ ;
	assign \g583/_0_  = _w32674_ ;
	assign \g5849/_3_  = _w32682_ ;
	assign \g585/_0_  = _w32685_ ;
	assign \g586/_0_  = _w32688_ ;
	assign \g587/_0_  = _w32691_ ;
	assign \g588/_0_  = _w32694_ ;
	assign \g589/_0_  = _w32697_ ;
	assign \g590/_0_  = _w32700_ ;
	assign \g591/_0_  = _w32703_ ;
	assign \g592/_0_  = _w32706_ ;
	assign \g593/_0_  = _w32709_ ;
	assign \g594/_0_  = _w32712_ ;
	assign \g595/_0_  = _w32715_ ;
	assign \g596/_0_  = _w32718_ ;
	assign \g597/_0_  = _w32721_ ;
	assign \g5971/_0_  = _w32724_ ;
	assign \g5972/_0_  = _w32727_ ;
	assign \g5976/_0_  = _w32730_ ;
	assign \g598/_0_  = _w32733_ ;
	assign \g5989/_0_  = _w32736_ ;
	assign \g599/_0_  = _w32739_ ;
	assign \g600/_0_  = _w32742_ ;
	assign \g601/_0_  = _w32745_ ;
	assign \g602/_0_  = _w32748_ ;
	assign \g603/_0_  = _w32751_ ;
	assign \g604/_0_  = _w32754_ ;
	assign \g605/_0_  = _w32757_ ;
	assign \g6092/_0_  = _w32760_ ;
	assign \g6093/_2_  = _w32953_ ;
	assign \g6094/_0_  = _w32958_ ;
	assign \g6114/_0_  = _w32959_ ;
	assign \g614/_3_  = _w32967_ ;
	assign \g6148/_0_  = _w32969_ ;
	assign \g6149/_0_  = _w32971_ ;
	assign \g6171/_0_  = _w33008_ ;
	assign \g6172/_0_  = _w33020_ ;
	assign \g6173/_0_  = _w33032_ ;
	assign \g6174/_0_  = _w33044_ ;
	assign \g6175/_0_  = _w33056_ ;
	assign \g6176/_0_  = _w33068_ ;
	assign \g6177/_0_  = _w33080_ ;
	assign \g6178/_0_  = _w33115_ ;
	assign \g6179/_0_  = _w33127_ ;
	assign \g6180/_0_  = _w33139_ ;
	assign \g6181/_0_  = _w33151_ ;
	assign \g6182/_0_  = _w33163_ ;
	assign \g6183/_0_  = _w33175_ ;
	assign \g6184/_0_  = _w33187_ ;
	assign \g6185/_0_  = _w33199_ ;
	assign \g6186/_0_  = _w33226_ ;
	assign \g6187/_0_  = _w33251_ ;
	assign \g6193/_0_  = _w33273_ ;
	assign \g6196/_0_  = _w33290_ ;
	assign \g6197/_0_  = _w33303_ ;
	assign \g6198/_3_  = _w33319_ ;
	assign \g6200/_2_  = _w31701_ ;
	assign \g6202/_2_  = _w31861_ ;
	assign \g6203/_3_  = _w33329_ ;
	assign \g6204/_3_  = _w33335_ ;
	assign \g6209/_0_  = _w33349_ ;
	assign \g6211/_0_  = _w33352_ ;
	assign \g6215/_0_  = _w33376_ ;
	assign \g6217/_0_  = _w33401_ ;
	assign \g6219/_0_  = _w33426_ ;
	assign \g6220/_0_  = _w33450_ ;
	assign \g6222/_0_  = _w33475_ ;
	assign \g6224/_0_  = _w33500_ ;
	assign \g6228/_0_  = _w33522_ ;
	assign \g6238/_0_  = _w33525_ ;
	assign \g6239/_0_  = _w33528_ ;
	assign \g6240/_0_  = _w33531_ ;
	assign \g6242/_0_  = _w33534_ ;
	assign \g6243/_0_  = _w33537_ ;
	assign \g6244/_0_  = _w33540_ ;
	assign \g6245/_0_  = _w33543_ ;
	assign \g6246/_0_  = _w33546_ ;
	assign \g6248/_0_  = _w33549_ ;
	assign \g6249/_0_  = _w33552_ ;
	assign \g6259/_0_  = _w33557_ ;
	assign \g6260/_0_  = _w33563_ ;
	assign \g6261/_0_  = _w33568_ ;
	assign \g6262/_0_  = _w33573_ ;
	assign \g6263/_0_  = _w33578_ ;
	assign \g6264/_0_  = _w33584_ ;
	assign \g6265/_0_  = _w33589_ ;
	assign \g6266/_0_  = _w33594_ ;
	assign \g6267/_0_  = _w33600_ ;
	assign \g6268/_0_  = _w33605_ ;
	assign \g6269/_0_  = _w33611_ ;
	assign \g6270/_0_  = _w33616_ ;
	assign \g6271/_0_  = _w33620_ ;
	assign \g6272/_0_  = _w33625_ ;
	assign \g6277/_0_  = _w33630_ ;
	assign \g6318/_0_  = _w33632_ ;
	assign \g6326/_0_  = _w33635_ ;
	assign \g6329/_0_  = _w33647_ ;
	assign \g6330/_0_  = _w33659_ ;
	assign \g6331/_0_  = _w33671_ ;
	assign \g6332/_0_  = _w33683_ ;
	assign \g6333/_0_  = _w33706_ ;
	assign \g6334/_0_  = _w33718_ ;
	assign \g6335/_0_  = _w33730_ ;
	assign \g6336/_0_  = _w33742_ ;
	assign \g6337/_0_  = _w33754_ ;
	assign \g6338/_0_  = _w33766_ ;
	assign \g6339/_0_  = _w33778_ ;
	assign \g6340/_0_  = _w33790_ ;
	assign \g6341/_0_  = _w33802_ ;
	assign \g6342/_0_  = _w33814_ ;
	assign \g6343/_0_  = _w33826_ ;
	assign \g6344/_0_  = _w33838_ ;
	assign \g6345/_0_  = _w33850_ ;
	assign \g6346/_0_  = _w33862_ ;
	assign \g6347/_0_  = _w33874_ ;
	assign \g6348/_0_  = _w33886_ ;
	assign \g6349/_0_  = _w33905_ ;
	assign \g6350/_0_  = _w33919_ ;
	assign \g6351/_0_  = _w33932_ ;
	assign \g6352/_0_  = _w33945_ ;
	assign \g6353/_0_  = _w33957_ ;
	assign \g6354/_0_  = _w33969_ ;
	assign \g6355/_0_  = _w33981_ ;
	assign \g6361/_0_  = _w33983_ ;
	assign \g637/_0_  = _w33989_ ;
	assign \g638/_0_  = _w33992_ ;
	assign \g639/_3_  = _w34002_ ;
	assign \g64/_3_  = _w34005_ ;
	assign \g640/_3_  = _w34011_ ;
	assign \g6419/_0_  = _w5681_ ;
	assign \g6442/_0_  = _w12234_ ;
	assign \g6442/_1_  = _w12234_ ;
	assign \g6489/_0_  = _w34012_ ;
	assign \g6490/_0_  = _w34013_ ;
	assign \g65/_3_  = _w34016_ ;
	assign \g6513/_0_  = _w34019_ ;
	assign \g6515/_0_  = _w34022_ ;
	assign \g6571/_0_  = _w34048_ ;
	assign \g6588/_0_  = _w34051_ ;
	assign \g6589/_0_  = _w34054_ ;
	assign \g6638/_0_  = _w34058_ ;
	assign \g6639/_0_  = _w34072_ ;
	assign \g6653/_0_  = _w34077_ ;
	assign \g6654/_3_  = _w34096_ ;
	assign \g6655/_0_  = _w34101_ ;
	assign \g6656/_0_  = _w34107_ ;
	assign \g6657/_0_  = _w34112_ ;
	assign \g6687/_0_  = _w34134_ ;
	assign \g6688/_0_  = _w34138_ ;
	assign \g6689/_0_  = _w34142_ ;
	assign \g6690/_0_  = _w34146_ ;
	assign \g6691/_0_  = _w34150_ ;
	assign \g6692/_0_  = _w34154_ ;
	assign \g6693/_0_  = _w34158_ ;
	assign \g6694/_0_  = _w34162_ ;
	assign \g6701/_0_  = _w34164_ ;
	assign \g6706/_0_  = _w34169_ ;
	assign \g6711/_0_  = _w34171_ ;
	assign \g6727/_0_  = _w34193_ ;
	assign \g6728/_0_  = _w34215_ ;
	assign \g6736/_0_  = _w34217_ ;
	assign \g6739/_0_  = _w34239_ ;
	assign \g6742/_0_  = _w34244_ ;
	assign \g6746/_0_  = _w34246_ ;
	assign \g6752/_0_  = _w34251_ ;
	assign \g6771/_0_  = _w34253_ ;
	assign \g684/_0_  = _w34283_ ;
	assign \g685/_0_  = _w34289_ ;
	assign \g686/_0_  = _w34295_ ;
	assign \g687/_0_  = _w34299_ ;
	assign \g688/_0_  = _w34305_ ;
	assign \g689/_0_  = _w34308_ ;
	assign \g690/_0_  = _w34314_ ;
	assign \g691/_0_  = _w34317_ ;
	assign \g692/_0_  = _w34320_ ;
	assign \g693/_0_  = _w34323_ ;
	assign \g696/_3_  = _w34333_ ;
	assign \g697/_3_  = _w34339_ ;
	assign \g699/_0_  = _w34378_ ;
	assign \g7/_0_  = _w34388_ ;
	assign \g700/_0_  = _w34418_ ;
	assign \g7005/_0_  = _w34434_ ;
	assign \g7056/_0_  = _w34437_ ;
	assign \g7057/_0_  = _w31705_ ;
	assign \g7058/_0_  = _w31868_ ;
	assign \g7060/_0_  = _w34440_ ;
	assign \g7075/_0_  = _w34460_ ;
	assign \g7086/_0_  = _w34468_ ;
	assign \g7087/_0_  = _w34473_ ;
	assign \g7089/_0_  = _w34483_ ;
	assign \g7108/_0_  = _w34489_ ;
	assign \g7109/_0_  = _w34495_ ;
	assign \g7112/_0_  = _w32088_ ;
	assign \g7172/_2_  = _w33344_ ;
	assign \g7210/_2_  = _w32658_ ;
	assign \g7211/_0_  = _w34500_ ;
	assign \g7212/_0_  = _w34505_ ;
	assign \g7213/_0_  = _w34510_ ;
	assign \g7214/_0_  = _w34515_ ;
	assign \g7215/_0_  = _w34520_ ;
	assign \g7216/_0_  = _w34525_ ;
	assign \g7217/_3_  = _w34531_ ;
	assign \g7218/_0_  = _w34536_ ;
	assign \g7219/_0_  = _w34541_ ;
	assign \g7220/_0_  = _w34546_ ;
	assign \g7222/_0_  = _w34551_ ;
	assign \g7227/_2_  = _w32612_ ;
	assign \g723/_3_  = _w34554_ ;
	assign \g7234/_0_  = _w34559_ ;
	assign \g7237/_3_  = _w34564_ ;
	assign \g7238/_3_  = _w34569_ ;
	assign \g7239/_3_  = _w13773_ ;
	assign \g724/_3_  = _w34572_ ;
	assign \g7240/_3_  = _w34578_ ;
	assign \g7241/_3_  = _w34583_ ;
	assign \g7242/_3_  = _w34588_ ;
	assign \g7243/_3_  = _w34593_ ;
	assign \g7244/_0_  = _w34598_ ;
	assign \g7245/_0_  = _w34603_ ;
	assign \g7246/_0_  = _w34608_ ;
	assign \g7247/_0_  = _w34613_ ;
	assign \g7248/_0_  = _w34618_ ;
	assign \g7249/_0_  = _w34623_ ;
	assign \g7250/_0_  = _w34628_ ;
	assign \g7251/_0_  = _w34633_ ;
	assign \g7253/_0_  = _w34637_ ;
	assign \g7254/_0_  = _w34640_ ;
	assign \g7255/_0_  = _w34642_ ;
	assign \g7256/_0_  = _w34644_ ;
	assign \g7257/_0_  = _w34646_ ;
	assign \g7258/_0_  = _w34648_ ;
	assign \g7261/_0_  = _w34650_ ;
	assign \g7264/_0_  = _w34662_ ;
	assign \g7265/_0_  = _w34674_ ;
	assign \g7266/_0_  = _w34686_ ;
	assign \g7267/_0_  = _w34698_ ;
	assign \g7268/_0_  = _w34710_ ;
	assign \g7269/_0_  = _w34722_ ;
	assign \g7278/_0_  = _w34734_ ;
	assign \g7279/_0_  = _w34746_ ;
	assign \g7280/_0_  = _w34758_ ;
	assign \g7281/_0_  = _w34770_ ;
	assign \g7282/_0_  = _w34782_ ;
	assign \g7283/_0_  = _w34794_ ;
	assign \g7284/_0_  = _w34806_ ;
	assign \g7285/_0_  = _w34818_ ;
	assign \g7286/_3_  = _w26973_ ;
	assign \g7288/_3_  = _w34822_ ;
	assign \g7291/_0_  = _w34824_ ;
	assign \g7296/_3_  = _w34863_ ;
	assign \g73/_0_  = _w34873_ ;
	assign \g7302/_3_  = _w34894_ ;
	assign \g7306/_3_  = _w34916_ ;
	assign \g7310/_3_  = _w34928_ ;
	assign \g7311/_3_  = _w34937_ ;
	assign \g7312/_3_  = _w34946_ ;
	assign \g7313/_3_  = _w34955_ ;
	assign \g7314/_3_  = _w34964_ ;
	assign \g7315/_3_  = _w34973_ ;
	assign \g7316/_3_  = _w34982_ ;
	assign \g7317/_3_  = _w34991_ ;
	assign \g7323/_3_  = _w35026_ ;
	assign \g7324/_3_  = _w35060_ ;
	assign \g7325/_3_  = _w35094_ ;
	assign \g7327/_0_  = _w35096_ ;
	assign \g7362/_0_  = _w35098_ ;
	assign \g74/_0_  = _w35108_ ;
	assign \g75/_0_  = _w35118_ ;
	assign \g7512/_0_  = _w13758_ ;
	assign \g7513/_0_  = _w35126_ ;
	assign \g7514/_0_  = _w35127_ ;
	assign \g7515/_0_  = _w35128_ ;
	assign \g7516/_0_  = _w35129_ ;
	assign \g7518/_0_  = _w35138_ ;
	assign \g7528/_0_  = _w35147_ ;
	assign \g7529/_0_  = _w35150_ ;
	assign \g7548/_0_  = _w35154_ ;
	assign \g7549/_0_  = _w35158_ ;
	assign \g7550/_0_  = _w35162_ ;
	assign \g7575/_0_  = _w35168_ ;
	assign \g7576/_0_  = _w35173_ ;
	assign \g7577/_0_  = _w35177_ ;
	assign \g7578/_0_  = _w35181_ ;
	assign \g7579/_0_  = _w35189_ ;
	assign \g7580/_0_  = _w35194_ ;
	assign \g7581/_0_  = _w35199_ ;
	assign \g7582/_0_  = _w35203_ ;
	assign \g7583/_0_  = _w35207_ ;
	assign \g7584/_0_  = _w35213_ ;
	assign \g7585/_0_  = _w35219_ ;
	assign \g7586/_0_  = _w35225_ ;
	assign \g7587/_0_  = _w35230_ ;
	assign \g7588/_0_  = _w35234_ ;
	assign \g7589/_0_  = _w35238_ ;
	assign \g7590/_0_  = _w35242_ ;
	assign \g7591/_0_  = _w35248_ ;
	assign \g7592/_0_  = _w35252_ ;
	assign \g7593/_0_  = _w35256_ ;
	assign \g7594/_0_  = _w35260_ ;
	assign \g7595/_0_  = _w35264_ ;
	assign \g7596/_0_  = _w35268_ ;
	assign \g7597/_0_  = _w35273_ ;
	assign \g7598/_0_  = _w35277_ ;
	assign \g7599/_0_  = _w35281_ ;
	assign \g76/_0_  = _w35291_ ;
	assign \g7600/_0_  = _w35295_ ;
	assign \g7601/_0_  = _w35299_ ;
	assign \g7602/_0_  = _w35303_ ;
	assign \g7603/_0_  = _w35308_ ;
	assign \g7604/_0_  = _w35312_ ;
	assign \g7614/_0_  = _w35317_ ;
	assign \g7618/_0_  = _w35318_ ;
	assign \g762/_0_  = _w35322_ ;
	assign \g7634/_0_  = _w32758_ ;
	assign \g766/_0_  = _w35328_ ;
	assign \g767/_0_  = _w35331_ ;
	assign \g768/_0_  = _w35337_ ;
	assign \g769/_0_  = _w35340_ ;
	assign \g77/_0_  = _w35350_ ;
	assign \g770/_3_  = _w35360_ ;
	assign \g771/_3_  = _w35366_ ;
	assign \g7715/_0_  = _w35397_ ;
	assign \g774/_0_  = _w35414_ ;
	assign \g7746/_0_  = _w35417_ ;
	assign \g7753/_0_  = _w35421_ ;
	assign \g7754/_0_  = _w35424_ ;
	assign \g7755/_0_  = _w35427_ ;
	assign \g7756/_0_  = _w35430_ ;
	assign \g7757/_0_  = _w35433_ ;
	assign \g7758/_0_  = _w35458_ ;
	assign \g7759/_0_  = _w35483_ ;
	assign \g7760/_0_  = _w35508_ ;
	assign \g7761/_0_  = _w35533_ ;
	assign \g7762/_0_  = _w35536_ ;
	assign \g7763/_0_  = _w35539_ ;
	assign \g7764/_0_  = _w35542_ ;
	assign \g7765/_0_  = _w35545_ ;
	assign \g7766/_0_  = _w35570_ ;
	assign \g7778/_0_  = _w35574_ ;
	assign \g7779/_0_  = _w35579_ ;
	assign \g7780/_0_  = _w35584_ ;
	assign \g7781/_0_  = _w35589_ ;
	assign \g7782/_0_  = _w35594_ ;
	assign \g7784/_0_  = _w35599_ ;
	assign \g78/_0_  = _w35609_ ;
	assign \g7800/_0_  = _w35611_ ;
	assign \g7823/_3_  = _w35614_ ;
	assign \g7837/_0_  = _w35619_ ;
	assign \g7841/_0_  = _w35624_ ;
	assign \g7842/_0_  = _w35629_ ;
	assign \g7843/_0_  = _w35634_ ;
	assign \g7844/_0_  = _w35639_ ;
	assign \g7845/_0_  = _w35644_ ;
	assign \g7846/_0_  = _w35649_ ;
	assign \g7847/_0_  = _w35654_ ;
	assign \g7849/_0_  = _w35656_ ;
	assign \g7850/_0_  = _w35661_ ;
	assign \g7852/_0_  = _w35663_ ;
	assign \g7854/_0_  = _w35665_ ;
	assign \g7855/_0_  = _w35670_ ;
	assign \g7857/_0_  = _w35677_ ;
	assign \g7858/_0_  = _w35683_ ;
	assign \g7859/_0_  = _w35689_ ;
	assign \g7860/_0_  = _w35695_ ;
	assign \g7861/_0_  = _w35701_ ;
	assign \g7862/_0_  = _w35707_ ;
	assign \g7863/_0_  = _w35713_ ;
	assign \g7864/_0_  = _w35719_ ;
	assign \g7865/_0_  = _w35725_ ;
	assign \g7866/_0_  = _w35731_ ;
	assign \g7867/_0_  = _w35737_ ;
	assign \g7868/_0_  = _w35743_ ;
	assign \g7869/_0_  = _w35749_ ;
	assign \g7870/_0_  = _w35755_ ;
	assign \g7871/_0_  = _w35760_ ;
	assign \g79211/_3_  = _w35763_ ;
	assign \g79258/_3_  = _w35766_ ;
	assign \g79299/_3_  = _w35769_ ;
	assign \g79316/_2_  = _w13534_ ;
	assign \g79342/_3_  = _w35772_ ;
	assign \g79401/_3_  = _w35775_ ;
	assign \g79452/_3_  = _w35778_ ;
	assign \g79457/_3_  = _w35781_ ;
	assign \g7951/_0_  = _w35783_ ;
	assign \g79541/_3_  = _w35786_ ;
	assign \g7958/_0_  = _w35788_ ;
	assign \g79598/_3_  = _w35791_ ;
	assign \g79654/_3_  = _w35794_ ;
	assign \g79675/_3_  = _w35797_ ;
	assign \g7971/_0_  = _w35800_ ;
	assign \g7972/_0_  = _w35820_ ;
	assign \g7973/_3_  = _w35849_ ;
	assign \g79753/_3_  = _w35852_ ;
	assign \g7976/_3_  = _w35881_ ;
	assign \g79855/_3_  = _w35884_ ;
	assign \g79858/_3_  = _w35887_ ;
	assign \g79997/_3_  = _w35890_ ;
	assign \g8/_0_  = _w35900_ ;
	assign \g80008/_3_  = _w11525_ ;
	assign \g80011/_0_  = _w35901_ ;
	assign \g80104/_0_  = _w19960_ ;
	assign \g80172/_1_  = _w12451_ ;
	assign \g80195/_3_  = _w8715_ ;
	assign \g80238/_3_  = _w35904_ ;
	assign \g80290/_2_  = _w7340_ ;
	assign \g80294/_0_  = _w10911_ ;
	assign \g80302/_0_  = _w11265_ ;
	assign \g80327/_0_  = _w35910_ ;
	assign \g80360/_3_  = _w10289_ ;
	assign \g80373/_0_  = _w35921_ ;
	assign \g80401/_0_  = _w7607_ ;
	assign \g80410/_0_  = _w8460_ ;
	assign \g80475/_0_  = _w7859_ ;
	assign \g80476/_0_  = _w10638_ ;
	assign \g80516/_3_  = _w35926_ ;
	assign \g80536/_0_  = _w35927_ ;
	assign \g80537/_0_  = _w9178_ ;
	assign \g80572/_0_  = _w35908_ ;
	assign \g80573/_0_  = _w35905_ ;
	assign \g80609/_2_  = _w12688_ ;
	assign \g80610/_2_  = _w12743_ ;
	assign \g80676/_0_  = _w22677_ ;
	assign \g80798/_0_  = _w35928_ ;
	assign \g80807/_0_  = _w25905_ ;
	assign \g80890/_2_  = _w5608_ ;
	assign \g80904/_0_  = _w25905_ ;
	assign \g81719/_2_  = _w19941_ ;
	assign \g81746/_0_  = _w5586_ ;
	assign \g81775/_0_  = _w5708_ ;
	assign \g81872/_0_  = _w35935_ ;
	assign \g81961/_0_  = _w4151_ ;
	assign \g81968/_0_  = _w4172_ ;
	assign \g82096/_0_  = _w4150_ ;
	assign \g82123/_0_  = _w4117_ ;
	assign \g82147/_0_  = _w4149_ ;
	assign \g82147/_1_  = _w4149_ ;
	assign \g82335/_0_  = _w5581_ ;
	assign \g82338/_2_  = _w5597_ ;
	assign \g82368/_0_  = _w4094_ ;
	assign \g82460/_2_  = _w22658_ ;
	assign \g82469/_0_  = _w19045_ ;
	assign \g82481/_0_  = _w4093_ ;
	assign \g82625/_1_  = _w12245_ ;
	assign \g82711/_0_  = _w5689_ ;
	assign \g82772/_0_  = _w4116_ ;
	assign \g82946/_0_  = _w22656_ ;
	assign \g82947/_0_  = _w19939_ ;
	assign \g82956/_0_  = _w5679_ ;
	assign \g83003/_0_  = _w4112_ ;
	assign \g83006/_1_  = _w12244_ ;
	assign \g83415/_0_  = _w5700_ ;
	assign \g83498/_0_  = _w4115_ ;
	assign \g837/_0_  = _w35941_ ;
	assign \g838/_0_  = _w35944_ ;
	assign \g83863/_0_  = _w12241_ ;
	assign \g839/_0_  = _w35955_ ;
	assign \g84049/_3_  = _w35961_ ;
	assign \g84050/_3_  = _w35967_ ;
	assign \g84077/_2_  = _w5692_ ;
	assign \g842/_0_  = _w35973_ ;
	assign \g84245/_0_  = _w4071_ ;
	assign \g843/_0_  = _w35979_ ;
	assign \g844/_0_  = _w35982_ ;
	assign \g84448/_0_  = _w6988_ ;
	assign \g84478/_3_  = _w35931_ ;
	assign \g845/_0_  = _w35988_ ;
	assign \g846/_0_  = _w35991_ ;
	assign \g847/_0_  = _w35994_ ;
	assign \g848/_0_  = _w36000_ ;
	assign \g8487/_0_  = _w36006_ ;
	assign \g8488/_0_  = _w36012_ ;
	assign \g8489/_0_  = _w36018_ ;
	assign \g849/_0_  = _w36021_ ;
	assign \g8490/_0_  = _w36027_ ;
	assign \g84904/_0_  = _w36028_ ;
	assign \g8491/_0_  = _w36032_ ;
	assign \g8492/_0_  = _w36038_ ;
	assign \g8493/_0_  = _w36042_ ;
	assign \g8494/_0_  = _w36048_ ;
	assign \g8496/_0_  = _w36049_ ;
	assign \g8517/_0_  = _w36052_ ;
	assign \g8534/_0_  = _w36055_ ;
	assign \g8538/_0_  = _w36064_ ;
	assign \g8540/_0_  = _w36067_ ;
	assign \g8576/_2_  = _w32038_ ;
	assign \g8597/_0_  = _w36072_ ;
	assign \g8598/_0_  = _w36078_ ;
	assign \g8599/_0_  = _w36082_ ;
	assign \g8600/_0_  = _w36086_ ;
	assign \g8601/_0_  = _w36090_ ;
	assign \g8602/_0_  = _w36094_ ;
	assign \g8603/_0_  = _w36098_ ;
	assign \g8605/_0_  = _w36101_ ;
	assign \g8606/_0_  = _w36104_ ;
	assign \g8607/_0_  = _w36107_ ;
	assign \g8608/_0_  = _w36112_ ;
	assign \g8609/_0_  = _w36116_ ;
	assign \g8610/_0_  = _w36120_ ;
	assign \g8611/_0_  = _w36124_ ;
	assign \g8612/_0_  = _w36128_ ;
	assign \g8613/_0_  = _w36132_ ;
	assign \g8614/_0_  = _w36136_ ;
	assign \g8615/_0_  = _w36140_ ;
	assign \g8617/_0_  = _w36143_ ;
	assign \g8643/_0_  = _w36147_ ;
	assign \g8644/_0_  = _w36151_ ;
	assign \g8645/_0_  = _w36155_ ;
	assign \g8646/_0_  = _w36159_ ;
	assign \g8647/_0_  = _w36163_ ;
	assign \g8648/_0_  = _w36167_ ;
	assign \g8650/_0_  = _w36170_ ;
	assign \g8651/_0_  = _w36173_ ;
	assign \g8652/_0_  = _w36176_ ;
	assign \g8653/_0_  = _w36180_ ;
	assign \g8654/_0_  = _w36184_ ;
	assign \g8655/_0_  = _w36188_ ;
	assign \g8656/_0_  = _w36192_ ;
	assign \g8657/_0_  = _w36196_ ;
	assign \g8658/_0_  = _w36200_ ;
	assign \g8659/_0_  = _w36204_ ;
	assign \g8660/_0_  = _w36208_ ;
	assign \g8665/_00_  = _w36217_ ;
	assign \g8666/_00_  = _w36224_ ;
	assign \g8667/_00_  = _w36231_ ;
	assign \g8668/_00_  = _w36238_ ;
	assign \g8669/_00_  = _w36245_ ;
	assign \g86715/_0_  = _w36248_ ;
	assign \g86745/_3_  = _w9435_ ;
	assign \g8691/_0_  = _w36252_ ;
	assign \g8700/_0_  = _w36259_ ;
	assign \g8701/_0_  = _w36265_ ;
	assign \g8702/_0_  = _w36271_ ;
	assign \g8703/_0_  = _w36277_ ;
	assign \g8704/_0_  = _w36283_ ;
	assign \g8705/_0_  = _w36289_ ;
	assign \g87063/_0_  = _w36321_ ;
	assign \g87114/_0_  = _w36353_ ;
	assign \g8712/_0_  = _w36355_ ;
	assign \g8713/_0_  = _w36361_ ;
	assign \g8714/_0_  = _w36367_ ;
	assign \g87171/_1_  = _w36373_ ;
	assign \g87252/_1_  = _w4099_ ;
	assign \g87298/_0_  = _w36374_ ;
	assign \g8730/_0_  = _w36379_ ;
	assign \g8741/_0_  = _w36384_ ;
	assign \g8747/_0_  = _w36387_ ;
	assign \g87480/_0_  = _w36388_ ;
	assign \g87484/_2_  = _w23032_ ;
	assign \g87488/_1__syn_2  = _w26297_ ;
	assign \g8761/_0_  = _w36399_ ;
	assign \g8762/_0_  = _w36404_ ;
	assign \g8763/_0_  = _w36415_ ;
	assign \g8764/_0_  = _w36420_ ;
	assign \g8765/_0_  = _w36426_ ;
	assign \g8775/_0_  = _w36448_ ;
	assign \g8776/_0_  = _w36457_ ;
	assign \g8777/_0_  = _w36461_ ;
	assign \g8778/_0_  = _w36463_ ;
	assign \g8784/_0_  = _w36468_ ;
	assign \g8804/_0_  = _w36476_ ;
	assign \g8807/_0_  = _w36479_ ;
	assign \g8808/_0_  = _w36483_ ;
	assign \g8809/_0_  = _w36487_ ;
	assign \g8810/_0_  = _w36490_ ;
	assign \g8811/_0_  = _w36494_ ;
	assign \g8812/_0_  = _w36497_ ;
	assign \g8813/_0_  = _w36500_ ;
	assign \g8814/_0_  = _w36503_ ;
	assign \g8815/_0_  = _w36506_ ;
	assign \g8816/_0_  = _w36510_ ;
	assign \g8817/_0_  = _w36513_ ;
	assign \g8818/_0_  = _w36519_ ;
	assign \g8819/_0_  = _w36524_ ;
	assign \g8820/_0_  = _w36529_ ;
	assign \g8821/_0_  = _w36533_ ;
	assign \g8822/_0_  = _w36536_ ;
	assign \g8823/_0_  = _w36538_ ;
	assign \g8824/_0_  = _w36541_ ;
	assign \g8825/_0_  = _w36544_ ;
	assign \g8826/_0_  = _w36547_ ;
	assign \g8827/_0_  = _w36550_ ;
	assign \g8828/_0_  = _w36553_ ;
	assign \g8829/_0_  = _w36555_ ;
	assign \g8830/_0_  = _w36558_ ;
	assign \g8831/_0_  = _w36561_ ;
	assign \g8832/_0_  = _w36564_ ;
	assign \g8833/_0_  = _w36567_ ;
	assign \g8834/_0_  = _w36571_ ;
	assign \g8835/_0_  = _w36574_ ;
	assign \g8836/_0_  = _w36578_ ;
	assign \g8837/_0_  = _w36581_ ;
	assign \g8838/_0_  = _w36584_ ;
	assign \g8839/_0_  = _w36586_ ;
	assign \g8840/_0_  = _w36589_ ;
	assign \g8842/_0_  = _w36594_ ;
	assign \g8843/_0_  = _w36599_ ;
	assign \g8846/_0_  = _w36602_ ;
	assign \g8848/_0_  = _w36607_ ;
	assign \g8857/_0_  = _w36609_ ;
	assign \g8895/_0_  = _w36612_ ;
	assign \g8902/_3_  = _w36648_ ;
	assign \g8903/_3_  = _w36684_ ;
	assign \g8904/_3_  = _w36720_ ;
	assign \g8905/_3_  = _w36756_ ;
	assign \g8906/_3_  = _w36792_ ;
	assign \g8909/_0_  = _w36795_ ;
	assign \g8910/_0_  = _w36798_ ;
	assign \g8911/_0_  = _w36801_ ;
	assign \g8924/_3_  = _w36833_ ;
	assign \g8926/_3_  = _w36865_ ;
	assign \g8927/_3_  = _w36897_ ;
	assign \g8943/_0_  = _w36899_ ;
	assign \g8944/_0_  = _w36901_ ;
	assign \g8958/_3_  = _w36933_ ;
	assign \g8960/_00_  = _w36940_ ;
	assign \g8961/_3_  = _w36972_ ;
	assign \g8965/_0_  = _w36988_ ;
	assign \g8966/_0_  = _w37004_ ;
	assign \g8967/_0_  = _w37020_ ;
	assign \g8968/_0_  = _w37036_ ;
	assign \g9/_0_  = _w37046_ ;
	assign \g9123/_0_  = _w32036_ ;
	assign \g9125/_0_  = _w37047_ ;
	assign \g9126/_0_  = _w37050_ ;
	assign \g913/_0_  = _w37066_ ;
	assign \g915/_0_  = _w37072_ ;
	assign \g916/_0_  = _w37078_ ;
	assign \g917/_0_  = _w37081_ ;
	assign \g918/_0_  = _w37087_ ;
	assign \g919/_0_  = _w37090_ ;
	assign \g920/_3_  = _w37100_ ;
	assign \g921/_3_  = _w37106_ ;
	assign \g925/_0_  = _w37122_ ;
	assign \g926/_0_  = _w37125_ ;
	assign \g927/_0_  = _w37131_ ;
	assign \g928/_0_  = _w37137_ ;
	assign \g929/_0_  = _w37140_ ;
	assign \g930/_0_  = _w37143_ ;
	assign \g9336/_0_  = _w37146_ ;
	assign \g9337/_0_  = _w37149_ ;
	assign \g939/_3_  = _w37162_ ;
	assign \g9396/_0_  = _w37168_ ;
	assign \g9397/_0_  = _w37171_ ;
	assign \g9399/_0_  = _w37174_ ;
	assign \g9400/_0_  = _w37177_ ;
	assign \g9401/_0_  = _w37180_ ;
	assign \g9402/_0_  = _w37183_ ;
	assign \g9403/_0_  = _w37186_ ;
	assign \g9404/_0_  = _w37189_ ;
	assign \g9415/_0_  = _w32613_ ;
	assign \g9418/_0_  = _w32659_ ;
	assign \g9419/_0_  = _w37202_ ;
	assign \g9420/_0_  = _w37205_ ;
	assign \g9446/_0_  = _w37206_ ;
	assign \g9465/_0_  = _w37207_ ;
	assign \g9493/_0_  = _w37210_ ;
	assign \g9536/_0_  = _w37214_ ;
	assign \g9537/_0_  = _w37220_ ;
	assign \g9538/_0_  = _w37223_ ;
	assign \g9539/_0_  = _w37226_ ;
	assign \g9540/_0_  = _w37229_ ;
	assign \g9541/_0_  = _w37235_ ;
	assign \g9542/_0_  = _w37239_ ;
	assign \g955/_2_  = _w37247_ ;
	assign \g9561/_0_  = _w37258_ ;
	assign \g9562/_0_  = _w37267_ ;
	assign \g9563/_0_  = _w37276_ ;
	assign \g9564/_0_  = _w37285_ ;
	assign \g9565/_0_  = _w37294_ ;
	assign \g9566/_0_  = _w37303_ ;
	assign \g9567/_0_  = _w37312_ ;
	assign \g9568/_0_  = _w37321_ ;
	assign \g9569/_0_  = _w37331_ ;
	assign \g9570/_0_  = _w37340_ ;
	assign \g9571/_0_  = _w37343_ ;
	assign \g9572/_0_  = _w37352_ ;
	assign \g9573/_0_  = _w37355_ ;
	assign \g9574/_0_  = _w37364_ ;
	assign \g9575/_0_  = _w37367_ ;
	assign \g9576/_0_  = _w37376_ ;
	assign \g9577/_0_  = _w37385_ ;
	assign \g9578/_0_  = _w37388_ ;
	assign \g9579/_0_  = _w37391_ ;
	assign \g9580/_0_  = _w37394_ ;
	assign \g9581/_0_  = _w37398_ ;
	assign \g9582/_0_  = _w37401_ ;
	assign \g9583/_0_  = _w37404_ ;
	assign \g9584/_0_  = _w37407_ ;
	assign \g9585/_0_  = _w37410_ ;
	assign \g9586/_0_  = _w37413_ ;
	assign \g9587/_0_  = _w37416_ ;
	assign \g9588/_0_  = _w37419_ ;
	assign \g9589/_0_  = _w37422_ ;
	assign \g9590/_0_  = _w37425_ ;
	assign \g9591/_0_  = _w37428_ ;
	assign \g9592/_0_  = _w37431_ ;
	assign \g9593/_0_  = _w37434_ ;
	assign \g9594/_0_  = _w37437_ ;
	assign \g9595/_0_  = _w37441_ ;
	assign \g9596/_0_  = _w37444_ ;
	assign \g9597/_0_  = _w37447_ ;
	assign \g9598/_0_  = _w37450_ ;
	assign \g9599/_0_  = _w37453_ ;
	assign \g9600/_0_  = _w37456_ ;
	assign \g9601/_0_  = _w37459_ ;
	assign \g9602/_0_  = _w37462_ ;
	assign \g9603/_0_  = _w37465_ ;
	assign \g9604/_0_  = _w37468_ ;
	assign \g9605/_0_  = _w37471_ ;
	assign \g9606/_0_  = _w37474_ ;
	assign \g9607/_0_  = _w37477_ ;
	assign \g9608/_0_  = _w37480_ ;
	assign \g9609/_0_  = _w37484_ ;
	assign \g9610/_0_  = _w37487_ ;
	assign \g9611/_0_  = _w37490_ ;
	assign \g9612/_0_  = _w37493_ ;
	assign \g9613/_0_  = _w37496_ ;
	assign \g9614/_0_  = _w37499_ ;
	assign \g9615/_0_  = _w37502_ ;
	assign \g9616/_0_  = _w37505_ ;
	assign \g9617/_0_  = _w37508_ ;
	assign \g9618/_0_  = _w37511_ ;
	assign \g9619/_0_  = _w37514_ ;
	assign \g9620/_0_  = _w37517_ ;
	assign \g9621/_0_  = _w37520_ ;
	assign \g9622/_0_  = _w37523_ ;
	assign \g9623/_0_  = _w37527_ ;
	assign \g9624/_0_  = _w37530_ ;
	assign \g9625/_0_  = _w37533_ ;
	assign \g9626/_0_  = _w37536_ ;
	assign \g9627/_0_  = _w37539_ ;
	assign \g9628/_0_  = _w37542_ ;
	assign \g9629/_0_  = _w37545_ ;
	assign \g9630/_0_  = _w37548_ ;
	assign \g9631/_0_  = _w37551_ ;
	assign \g9632/_0_  = _w37554_ ;
	assign \g9633/_0_  = _w37557_ ;
	assign \g9634/_0_  = _w37560_ ;
	assign \g9635/_0_  = _w37563_ ;
	assign \g9636/_0_  = _w37566_ ;
	assign \g9637/_0_  = _w37570_ ;
	assign \g9638/_0_  = _w37573_ ;
	assign \g9639/_0_  = _w37576_ ;
	assign \g9640/_0_  = _w37579_ ;
	assign \g9641/_0_  = _w37582_ ;
	assign \g9642/_0_  = _w37585_ ;
	assign \g9643/_0_  = _w37588_ ;
	assign \g9644/_0_  = _w37591_ ;
	assign \g9645/_0_  = _w37594_ ;
	assign \g9646/_0_  = _w37597_ ;
	assign \g9647/_0_  = _w37600_ ;
	assign \g9648/_0_  = _w37603_ ;
	assign \g9649/_0_  = _w37606_ ;
	assign \g9650/_0_  = _w37609_ ;
	assign \g9651/_0_  = _w37613_ ;
	assign \g9652/_0_  = _w37616_ ;
	assign \g9653/_0_  = _w37619_ ;
	assign \g9654/_0_  = _w37622_ ;
	assign \g9655/_0_  = _w37625_ ;
	assign \g9656/_0_  = _w37628_ ;
	assign \g9657/_0_  = _w37631_ ;
	assign \g9658/_0_  = _w37634_ ;
	assign \g9659/_0_  = _w37637_ ;
	assign \g9660/_0_  = _w37640_ ;
	assign \g9661/_0_  = _w37643_ ;
	assign \g9662/_0_  = _w37646_ ;
	assign \g9663/_0_  = _w37649_ ;
	assign \g9664/_0_  = _w37652_ ;
	assign \g9665/_0_  = _w37656_ ;
	assign \g9666/_0_  = _w37659_ ;
	assign \g9667/_0_  = _w37662_ ;
	assign \g9668/_0_  = _w37665_ ;
	assign \g9669/_0_  = _w37668_ ;
	assign \g9670/_0_  = _w37671_ ;
	assign \g9671/_0_  = _w37674_ ;
	assign \g9672/_0_  = _w37677_ ;
	assign \g9673/_0_  = _w37680_ ;
	assign \g9674/_0_  = _w37683_ ;
	assign \g9675/_0_  = _w37686_ ;
	assign \g9676/_0_  = _w37689_ ;
	assign \g9677/_0_  = _w37692_ ;
	assign \g9678/_0_  = _w37695_ ;
	assign \g9681/_0_  = _w37700_ ;
	assign \g9683/_0_  = _w37703_ ;
	assign \g9689/_0_  = _w37708_ ;
	assign \g9692/_0_  = _w37712_ ;
	assign \g9694/_0_  = _w37717_ ;
	assign \g9695/_0_  = _w37722_ ;
	assign \g9701/_0_  = _w37726_ ;
	assign \g9702/_0_  = _w37731_ ;
	assign \g9703/_0_  = _w37736_ ;
	assign \g9704/_0_  = _w37741_ ;
	assign \g9709/_0_  = _w37745_ ;
	assign \g9710/_0_  = _w37748_ ;
	assign \g9711/_0_  = _w37751_ ;
	assign \g9712/_0_  = _w37754_ ;
	assign \g9720/_0_  = _w37757_ ;
	assign \g9721/_0_  = _w37760_ ;
	assign \g9722/_0_  = _w37763_ ;
	assign \g9726/_0_  = _w37766_ ;
	assign \g9733/_0_  = _w37770_ ;
	assign \g9734/_0_  = _w37773_ ;
	assign \g9735/_0_  = _w37776_ ;
	assign \g9736/_0_  = _w37779_ ;
	assign \g9737/_0_  = _w37782_ ;
	assign \g9738/_0_  = _w37785_ ;
	assign \g9739/_0_  = _w37788_ ;
	assign \g9740/_0_  = _w37791_ ;
	assign \g9741/_0_  = _w37794_ ;
	assign \g9742/_0_  = _w37797_ ;
	assign \g9743/_0_  = _w37800_ ;
	assign \g9744/_0_  = _w37803_ ;
	assign \g9745/_0_  = _w37806_ ;
	assign \g9746/_0_  = _w37809_ ;
	assign \g9747/_0_  = _w37813_ ;
	assign \g9748/_0_  = _w37816_ ;
	assign \g9749/_0_  = _w37819_ ;
	assign \g9750/_0_  = _w37822_ ;
	assign \g9751/_0_  = _w37825_ ;
	assign \g9752/_0_  = _w37828_ ;
	assign \g9753/_0_  = _w37831_ ;
	assign \g9754/_0_  = _w37834_ ;
	assign \g9755/_0_  = _w37837_ ;
	assign \g9756/_0_  = _w37840_ ;
	assign \g9757/_0_  = _w37843_ ;
	assign \g9758/_0_  = _w37846_ ;
	assign \g9759/_0_  = _w37849_ ;
	assign \g9760/_0_  = _w37852_ ;
	assign \g9761/_0_  = _w37856_ ;
	assign \g9762/_0_  = _w37859_ ;
	assign \g9763/_0_  = _w37862_ ;
	assign \g9764/_0_  = _w37865_ ;
	assign \g9765/_0_  = _w37868_ ;
	assign \g9766/_0_  = _w37871_ ;
	assign \g9767/_0_  = _w37874_ ;
	assign \g9768/_0_  = _w37877_ ;
	assign \g9769/_0_  = _w37880_ ;
	assign \g9770/_0_  = _w37883_ ;
	assign \g9771/_0_  = _w37886_ ;
	assign \g9772/_0_  = _w37889_ ;
	assign \g9773/_0_  = _w37892_ ;
	assign \g9774/_0_  = _w37895_ ;
	assign \g9775/_0_  = _w37899_ ;
	assign \g9776/_0_  = _w37902_ ;
	assign \g9777/_0_  = _w37905_ ;
	assign \g9778/_0_  = _w37908_ ;
	assign \g9779/_0_  = _w37911_ ;
	assign \g9780/_0_  = _w37914_ ;
	assign \g9781/_0_  = _w37917_ ;
	assign \g9782/_0_  = _w37920_ ;
	assign \g9783/_0_  = _w37923_ ;
	assign \g9784/_0_  = _w37926_ ;
	assign \g9785/_0_  = _w37929_ ;
	assign \g9786/_0_  = _w37932_ ;
	assign \g9787/_0_  = _w37935_ ;
	assign \g9788/_0_  = _w37938_ ;
	assign \g9789/_0_  = _w37942_ ;
	assign \g9790/_0_  = _w37945_ ;
	assign \g9791/_0_  = _w37948_ ;
	assign \g9792/_0_  = _w37951_ ;
	assign \g9793/_0_  = _w37954_ ;
	assign \g9794/_0_  = _w37957_ ;
	assign \g9795/_0_  = _w37960_ ;
	assign \g9796/_0_  = _w37963_ ;
	assign \g9797/_0_  = _w37966_ ;
	assign \g9798/_0_  = _w37969_ ;
	assign \g9799/_0_  = _w37972_ ;
	assign \g9800/_0_  = _w37975_ ;
	assign \g9801/_0_  = _w37978_ ;
	assign \g9802/_0_  = _w37981_ ;
	assign \g9803/_0_  = _w37985_ ;
	assign \g9804/_0_  = _w37988_ ;
	assign \g9805/_0_  = _w37991_ ;
	assign \g9806/_0_  = _w37994_ ;
	assign \g9807/_0_  = _w37997_ ;
	assign \g9808/_0_  = _w38000_ ;
	assign \g9809/_0_  = _w38003_ ;
	assign \g9810/_0_  = _w38006_ ;
	assign \g9811/_0_  = _w38009_ ;
	assign \g9812/_0_  = _w38012_ ;
	assign \g9813/_0_  = _w38015_ ;
	assign \g9814/_0_  = _w38018_ ;
	assign \g9815/_0_  = _w38021_ ;
	assign \g9816/_0_  = _w38024_ ;
	assign \g9817/_0_  = _w38028_ ;
	assign \g9818/_0_  = _w38031_ ;
	assign \g9819/_0_  = _w38034_ ;
	assign \g9820/_0_  = _w38037_ ;
	assign \g9821/_0_  = _w38040_ ;
	assign \g9822/_0_  = _w38043_ ;
	assign \g9823/_0_  = _w38046_ ;
	assign \g9824/_0_  = _w38049_ ;
	assign \g9825/_0_  = _w38052_ ;
	assign \g9826/_0_  = _w38055_ ;
	assign \g9827/_0_  = _w38058_ ;
	assign \g9828/_0_  = _w38061_ ;
	assign \g9829/_0_  = _w38064_ ;
	assign \g9830/_0_  = _w38067_ ;
	assign \g9831/_0_  = _w38070_ ;
	assign \g9832/_0_  = _w38073_ ;
	assign \g9833/_0_  = _w38076_ ;
	assign \g9835/_0_  = _w38079_ ;
	assign \g9836/_0_  = _w38082_ ;
	assign \g9837/_0_  = _w38085_ ;
	assign \g9838/_0_  = _w38088_ ;
	assign \g9839/_0_  = _w38091_ ;
	assign \g9840/_0_  = _w38094_ ;
	assign \g9841/_0_  = _w38097_ ;
	assign \g9842/_0_  = _w38100_ ;
	assign \g9844/_0_  = _w38103_ ;
	assign \g9845/_0_  = _w38106_ ;
	assign \g9846/_0_  = _w38109_ ;
	assign \g9848/_0_  = _w38112_ ;
	assign \g9849/_0_  = _w38115_ ;
	assign \g9850/_0_  = _w38120_ ;
	assign \g9851/_0_  = _w38125_ ;
	assign \g9853/_0_  = _w38130_ ;
	assign \g9854/_0_  = _w38135_ ;
	assign \g9855/_0_  = _w38140_ ;
	assign \g9856/_0_  = _w38146_ ;
	assign \g9857/_0_  = _w38149_ ;
	assign \g9858/_0_  = _w38152_ ;
	assign \g9859/_0_  = _w38155_ ;
	assign \g9860/_0_  = _w38158_ ;
	assign \g9862/_0_  = _w38162_ ;
	assign \g9863/_0_  = _w38166_ ;
	assign \g9864/_0_  = _w38170_ ;
	assign \g9865/_0_  = _w38174_ ;
	assign \g9867/_0_  = _w38179_ ;
	assign \g9868/_0_  = _w38182_ ;
	assign \g9876/_0_  = _w38185_ ;
	assign \g9877/_0_  = _w38188_ ;
	assign \g9878/_0_  = _w38191_ ;
	assign \g9879/_0_  = _w38194_ ;
	assign \g9880/_0_  = _w38197_ ;
	assign \g9881/_0_  = _w38200_ ;
	assign \g9898/_0_  = _w38204_ ;
	assign \g9900/_0_  = _w38207_ ;
	assign \g9901/_0_  = _w38210_ ;
	assign \g9902/_0_  = _w38213_ ;
	assign \g9903/_0_  = _w38216_ ;
	assign \g9904/_0_  = _w38219_ ;
	assign \g9905/_0_  = _w38222_ ;
	assign \g9906/_0_  = _w38225_ ;
	assign \g9907/_0_  = _w38228_ ;
	assign \g9908/_0_  = _w38231_ ;
	assign \g9909/_0_  = _w38234_ ;
	assign \g9910/_0_  = _w38237_ ;
	assign \g9911/_0_  = _w38240_ ;
	assign \g9912/_0_  = _w38243_ ;
	assign \g9913/_0_  = _w38246_ ;
	assign \g9914/_0_  = _w38249_ ;
	assign \g9915/_0_  = _w38252_ ;
	assign \g9916/_0_  = _w38255_ ;
	assign \g9917/_0_  = _w38258_ ;
	assign \g9918/_0_  = _w38261_ ;
	assign \g9919/_0_  = _w38264_ ;
	assign \g992/_0_  = _w38279_ ;
	assign \g9920/_0_  = _w38282_ ;
	assign \g9921/_0_  = _w38285_ ;
	assign \g9922/_0_  = _w38288_ ;
	assign \g9923/_0_  = _w38291_ ;
	assign \g9924/_0_  = _w38295_ ;
	assign \g9925/_0_  = _w38298_ ;
	assign \g9926/_0_  = _w38301_ ;
	assign \g9927/_0_  = _w38304_ ;
	assign \g9928/_0_  = _w38307_ ;
	assign \g9929/_0_  = _w38310_ ;
	assign \g9930/_0_  = _w38313_ ;
	assign \g9931/_0_  = _w38316_ ;
	assign \g9932/_0_  = _w38319_ ;
	assign \g9933/_0_  = _w38322_ ;
	assign \g9934/_0_  = _w38325_ ;
	assign \g9935/_0_  = _w38328_ ;
	assign \g9936/_0_  = _w38331_ ;
	assign \g9937/_0_  = _w38334_ ;
	assign \g9938/_0_  = _w38337_ ;
	assign \g9939/_0_  = _w38340_ ;
	assign \g9940/_0_  = _w38343_ ;
	assign \g9941/_0_  = _w38346_ ;
	assign \g9942/_0_  = _w38349_ ;
	assign \g9943/_0_  = _w38352_ ;
	assign \g9944/_0_  = _w38355_ ;
	assign \g9945/_0_  = _w38358_ ;
	assign \g9946/_0_  = _w38361_ ;
	assign \g9947/_0_  = _w38364_ ;
	assign \g9948/_0_  = _w38367_ ;
	assign \g9949/_0_  = _w38371_ ;
	assign \g9950/_0_  = _w38374_ ;
	assign \g9951/_0_  = _w38377_ ;
	assign \g9952/_0_  = _w38380_ ;
	assign \g9953/_0_  = _w38383_ ;
	assign \g9954/_0_  = _w38386_ ;
	assign \g9955/_0_  = _w38389_ ;
	assign \g9956/_0_  = _w38392_ ;
	assign \g9957/_0_  = _w38395_ ;
	assign \g9958/_0_  = _w38398_ ;
	assign \g9959/_0_  = _w38401_ ;
	assign \g9960/_0_  = _w38404_ ;
	assign \g9961/_0_  = _w38407_ ;
	assign \g9962/_0_  = _w38410_ ;
	assign \g9963/_0_  = _w38413_ ;
	assign \g9964/_0_  = _w38416_ ;
	assign \g9965/_0_  = _w38419_ ;
	assign \g9966/_0_  = _w38422_ ;
	assign \g9967/_0_  = _w38425_ ;
	assign \g9968/_0_  = _w38428_ ;
	assign \g9969/_0_  = _w38431_ ;
	assign \g9970/_0_  = _w38434_ ;
	assign \g9971/_0_  = _w38437_ ;
	assign \g9972/_0_  = _w38440_ ;
	assign \g9973/_0_  = _w38443_ ;
	assign \g9974/_0_  = _w38446_ ;
	assign \g9975/_0_  = _w38449_ ;
	assign \g9976/_0_  = _w38452_ ;
	assign \g9977/_0_  = _w38455_ ;
	assign \g9978/_0_  = _w38458_ ;
	assign \g9979/_0_  = _w38461_ ;
	assign \g9980/_0_  = _w38464_ ;
	assign \g9981/_0_  = _w38467_ ;
	assign \g9982/_0_  = _w38470_ ;
	assign \g9983/_0_  = _w38473_ ;
	assign \g9984/_0_  = _w38476_ ;
	assign \g9985/_0_  = _w38479_ ;
	assign \g9987/_0_  = _w38482_ ;
	assign \g9988/_0_  = _w38485_ ;
	assign \g9989/_0_  = _w38488_ ;
	assign \g999/_0_  = _w38491_ ;
	assign \g9990/_0_  = _w38494_ ;
	assign \g9991/_0_  = _w38497_ ;
	assign \g9992/_0_  = _w38500_ ;
	assign \g9993/_0_  = _w38503_ ;
	assign \g9994/_0_  = _w38506_ ;
	assign \g9995/_0_  = _w38509_ ;
	assign \g9996/_0_  = _w38512_ ;
	assign \g9997/_0_  = _w38515_ ;
	assign \g9998/_0_  = _w38518_ ;
	assign \g9999/_0_  = _w38521_ ;
	assign \idma_IDMA_boot_reg/NET0131_reg_syn_3  = _w38522_ ;
	assign \memc_EXTC_Eg_reg/NET0131  = _w4068_ ;
	assign \memc_EXTC_Eg_reg/NET0131_reg_syn_3  = _w38524_ ;
	assign \memc_EXTC_Eg_reg/n0  = _w38523_ ;
	assign \pio_PIO_IN_P_reg[0]/P0001_reg_syn_3  = _w38527_ ;
	assign \pio_PIO_IN_P_reg[10]/P0001_reg_syn_3  = _w38530_ ;
	assign \pio_PIO_IN_P_reg[11]/P0001_reg_syn_3  = _w38533_ ;
	assign \pio_PIO_IN_P_reg[1]/P0001_reg_syn_3  = _w38536_ ;
	assign \pio_PIO_IN_P_reg[2]/P0001_reg_syn_3  = _w38539_ ;
	assign \pio_PIO_IN_P_reg[3]/P0001_reg_syn_3  = _w38542_ ;
	assign \pio_PIO_IN_P_reg[4]/P0001_reg_syn_3  = _w38545_ ;
	assign \pio_PIO_IN_P_reg[5]/P0001_reg_syn_3  = _w38548_ ;
	assign \pio_PIO_IN_P_reg[6]/P0001_reg_syn_3  = _w38551_ ;
	assign \pio_PIO_IN_P_reg[7]/P0001_reg_syn_3  = _w38554_ ;
	assign \pio_PIO_IN_P_reg[8]/P0001_reg_syn_3  = _w38557_ ;
	assign \pio_PIO_IN_P_reg[9]/P0001_reg_syn_3  = _w38560_ ;
	assign \pio_PIO_RES_OUT_reg[0]/P0001_reg_syn_3  = _w38563_ ;
	assign \pio_PIO_RES_OUT_reg[10]/P0001_reg_syn_3  = _w38566_ ;
	assign \pio_PIO_RES_OUT_reg[2]/P0001_reg_syn_3  = _w38569_ ;
	assign \pio_PIO_RES_OUT_reg[4]/P0001_reg_syn_3  = _w38572_ ;
	assign \pio_PIO_RES_OUT_reg[6]/P0001_reg_syn_3  = _w38575_ ;
	assign \sice_GO_NXi_reg/NET0131_reg_syn_3  = _w38578_ ;
	assign \sport0_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  = _w38581_ ;
	assign \sport0_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  = _w38583_ ;
	assign \sport1_rxctl_RXSHT_reg[0]/P0001_reg_syn_3  = _w38586_ ;
	assign \sport1_rxctl_RXSHT_reg[1]/P0001_reg_syn_3  = _w38588_ ;
endmodule;