module top( \d_in_reg[0]/NET0131  , \d_in_reg[1]/NET0131  , \d_in_reg[2]/NET0131  , \d_in_reg[3]/NET0131  , \d_in_reg[4]/NET0131  , \d_in_reg[5]/NET0131  , \d_in_reg[6]/NET0131  , \d_in_reg[7]/NET0131  , \d_in_reg[8]/NET0131  , \d_out_reg[0]/NET0131  , \d_out_reg[1]/NET0131  , \d_out_reg[2]/NET0131  , \d_out_reg[3]/NET0131  , \d_out_reg[4]/NET0131  , \d_out_reg[5]/NET0131  , \d_out_reg[6]/NET0131  , \d_out_reg[7]/NET0131  , \old_reg[0]/NET0131  , \old_reg[1]/NET0131  , \old_reg[2]/NET0131  , \old_reg[3]/NET0131  , \old_reg[4]/NET0131  , \old_reg[5]/NET0131  , \old_reg[6]/NET0131  , \old_reg[7]/NET0131  , \stato_reg[0]/NET0131  , \stato_reg[1]/NET0131  , x_pad , y_pad , \_al_n0  , \_al_n1  , \g1026/_0_  , \g1035/_0_  , \g41/_0_  , \g708/_0_  , \g709/_0_  , \g711/_0_  , \g712/_0_  , \g714/_0_  , \g716/_0_  , \g718/_0_  , \g728/_0_  , \g770/_0_  , \g771/_0_  , \g772/_0_  , \g773/_0_  , \g774/_0_  , \g775/_0_  , \g776/_0_  , \g777/_0_  , \g782/_0_  , \g783/_0_  , \g784/_0_  , \g785/_0_  , \g786/_0_  , \g787/_0_  , \g788/_0_  , \g789/_0_  , \g806/_0_  );
  input \d_in_reg[0]/NET0131  ;
  input \d_in_reg[1]/NET0131  ;
  input \d_in_reg[2]/NET0131  ;
  input \d_in_reg[3]/NET0131  ;
  input \d_in_reg[4]/NET0131  ;
  input \d_in_reg[5]/NET0131  ;
  input \d_in_reg[6]/NET0131  ;
  input \d_in_reg[7]/NET0131  ;
  input \d_in_reg[8]/NET0131  ;
  input \d_out_reg[0]/NET0131  ;
  input \d_out_reg[1]/NET0131  ;
  input \d_out_reg[2]/NET0131  ;
  input \d_out_reg[3]/NET0131  ;
  input \d_out_reg[4]/NET0131  ;
  input \d_out_reg[5]/NET0131  ;
  input \d_out_reg[6]/NET0131  ;
  input \d_out_reg[7]/NET0131  ;
  input \old_reg[0]/NET0131  ;
  input \old_reg[1]/NET0131  ;
  input \old_reg[2]/NET0131  ;
  input \old_reg[3]/NET0131  ;
  input \old_reg[4]/NET0131  ;
  input \old_reg[5]/NET0131  ;
  input \old_reg[6]/NET0131  ;
  input \old_reg[7]/NET0131  ;
  input \stato_reg[0]/NET0131  ;
  input \stato_reg[1]/NET0131  ;
  input x_pad ;
  input y_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g1026/_0_  ;
  output \g1035/_0_  ;
  output \g41/_0_  ;
  output \g708/_0_  ;
  output \g709/_0_  ;
  output \g711/_0_  ;
  output \g712/_0_  ;
  output \g714/_0_  ;
  output \g716/_0_  ;
  output \g718/_0_  ;
  output \g728/_0_  ;
  output \g770/_0_  ;
  output \g771/_0_  ;
  output \g772/_0_  ;
  output \g773/_0_  ;
  output \g774/_0_  ;
  output \g775/_0_  ;
  output \g776/_0_  ;
  output \g777/_0_  ;
  output \g782/_0_  ;
  output \g783/_0_  ;
  output \g784/_0_  ;
  output \g785/_0_  ;
  output \g786/_0_  ;
  output \g787/_0_  ;
  output \g788/_0_  ;
  output \g789/_0_  ;
  output \g806/_0_  ;
  wire n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 ;
  assign n30 = ~\d_in_reg[4]/NET0131  & ~\old_reg[3]/NET0131  ;
  assign n31 = \d_in_reg[4]/NET0131  & \old_reg[3]/NET0131  ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = ~\d_in_reg[5]/NET0131  & ~\old_reg[4]/NET0131  ;
  assign n34 = \d_in_reg[5]/NET0131  & \old_reg[4]/NET0131  ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = ~n32 & ~n35 ;
  assign n37 = ~\d_in_reg[8]/NET0131  & ~\old_reg[7]/NET0131  ;
  assign n38 = \d_in_reg[8]/NET0131  & \old_reg[7]/NET0131  ;
  assign n39 = ~n37 & ~n38 ;
  assign n40 = ~\d_in_reg[7]/NET0131  & ~\old_reg[6]/NET0131  ;
  assign n41 = \d_in_reg[7]/NET0131  & \old_reg[6]/NET0131  ;
  assign n42 = ~n40 & ~n41 ;
  assign n43 = ~n39 & ~n42 ;
  assign n44 = n36 & n43 ;
  assign n45 = \d_in_reg[3]/NET0131  & ~\old_reg[2]/NET0131  ;
  assign n46 = ~\d_in_reg[3]/NET0131  & \old_reg[2]/NET0131  ;
  assign n47 = ~n45 & ~n46 ;
  assign n48 = \d_in_reg[6]/NET0131  & ~\old_reg[5]/NET0131  ;
  assign n49 = ~\d_in_reg[6]/NET0131  & \old_reg[5]/NET0131  ;
  assign n50 = ~n48 & ~n49 ;
  assign n51 = n47 & n50 ;
  assign n52 = ~\d_in_reg[2]/NET0131  & ~\old_reg[1]/NET0131  ;
  assign n53 = \d_in_reg[2]/NET0131  & \old_reg[1]/NET0131  ;
  assign n54 = ~n52 & ~n53 ;
  assign n55 = ~\d_in_reg[1]/NET0131  & ~\old_reg[0]/NET0131  ;
  assign n56 = \d_in_reg[1]/NET0131  & \old_reg[0]/NET0131  ;
  assign n57 = ~n55 & ~n56 ;
  assign n58 = ~n54 & ~n57 ;
  assign n59 = n51 & n58 ;
  assign n60 = n44 & n59 ;
  assign n61 = \stato_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n62 = \d_in_reg[0]/NET0131  & n61 ;
  assign n63 = \d_in_reg[1]/NET0131  & n62 ;
  assign n64 = ~n60 & n63 ;
  assign n65 = \d_out_reg[0]/NET0131  & n62 ;
  assign n66 = n60 & n65 ;
  assign n67 = ~n64 & ~n66 ;
  assign n68 = \d_in_reg[0]/NET0131  & ~\stato_reg[0]/NET0131  ;
  assign n69 = \d_out_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n70 = n68 & n69 ;
  assign n71 = ~\d_in_reg[0]/NET0131  & \d_out_reg[0]/NET0131  ;
  assign n72 = \stato_reg[0]/NET0131  & n71 ;
  assign n73 = ~n70 & ~n72 ;
  assign n74 = \stato_reg[0]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n75 = \d_in_reg[0]/NET0131  & \d_in_reg[1]/NET0131  ;
  assign n76 = n74 & n75 ;
  assign n77 = ~\stato_reg[0]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n78 = ~\d_in_reg[0]/NET0131  & \d_out_reg[1]/NET0131  ;
  assign n79 = n77 & n78 ;
  assign n80 = ~n76 & ~n79 ;
  assign n81 = n73 & n80 ;
  assign n82 = n67 & n81 ;
  assign n83 = \d_in_reg[2]/NET0131  & n62 ;
  assign n84 = ~n60 & n83 ;
  assign n85 = \d_out_reg[1]/NET0131  & n62 ;
  assign n86 = n60 & n85 ;
  assign n87 = ~n84 & ~n86 ;
  assign n88 = \d_out_reg[1]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n89 = n68 & n88 ;
  assign n90 = \stato_reg[0]/NET0131  & n78 ;
  assign n91 = ~n89 & ~n90 ;
  assign n92 = \d_in_reg[0]/NET0131  & \d_in_reg[2]/NET0131  ;
  assign n93 = n74 & n92 ;
  assign n94 = ~\d_in_reg[0]/NET0131  & \d_out_reg[2]/NET0131  ;
  assign n95 = n77 & n94 ;
  assign n96 = ~n93 & ~n95 ;
  assign n97 = n91 & n96 ;
  assign n98 = n87 & n97 ;
  assign n99 = \d_in_reg[8]/NET0131  & n62 ;
  assign n100 = ~n60 & n99 ;
  assign n101 = \d_out_reg[7]/NET0131  & n62 ;
  assign n102 = n60 & n101 ;
  assign n103 = ~n100 & ~n102 ;
  assign n104 = \d_out_reg[7]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n105 = n68 & n104 ;
  assign n106 = ~\d_in_reg[0]/NET0131  & \d_out_reg[7]/NET0131  ;
  assign n107 = \stato_reg[0]/NET0131  & n106 ;
  assign n108 = ~n105 & ~n107 ;
  assign n109 = \d_in_reg[0]/NET0131  & \d_in_reg[8]/NET0131  ;
  assign n110 = n74 & n109 ;
  assign n111 = n108 & ~n110 ;
  assign n112 = n103 & n111 ;
  assign n113 = \d_in_reg[0]/NET0131  & \stato_reg[0]/NET0131  ;
  assign n114 = ~\d_in_reg[0]/NET0131  & \stato_reg[0]/NET0131  ;
  assign n115 = ~n77 & ~n114 ;
  assign n116 = x_pad & ~n115 ;
  assign n117 = ~n113 & ~n116 ;
  assign n118 = \stato_reg[1]/NET0131  & ~n116 ;
  assign n119 = n60 & n118 ;
  assign n120 = ~n117 & ~n119 ;
  assign n121 = \d_in_reg[4]/NET0131  & n62 ;
  assign n122 = ~n60 & n121 ;
  assign n123 = \d_out_reg[3]/NET0131  & n62 ;
  assign n124 = n60 & n123 ;
  assign n125 = ~n122 & ~n124 ;
  assign n126 = \d_in_reg[0]/NET0131  & \d_out_reg[3]/NET0131  ;
  assign n127 = n77 & n126 ;
  assign n128 = ~\d_in_reg[0]/NET0131  & \d_out_reg[3]/NET0131  ;
  assign n129 = n61 & n128 ;
  assign n130 = ~n127 & ~n129 ;
  assign n131 = \d_in_reg[0]/NET0131  & \d_in_reg[4]/NET0131  ;
  assign n132 = ~n128 & ~n131 ;
  assign n133 = n74 & ~n132 ;
  assign n134 = ~\d_in_reg[0]/NET0131  & \d_out_reg[4]/NET0131  ;
  assign n135 = n77 & n134 ;
  assign n136 = ~n133 & ~n135 ;
  assign n137 = n130 & n136 ;
  assign n138 = n125 & n137 ;
  assign n139 = \d_in_reg[5]/NET0131  & n62 ;
  assign n140 = ~n60 & n139 ;
  assign n141 = \d_out_reg[4]/NET0131  & n62 ;
  assign n142 = n60 & n141 ;
  assign n143 = ~n140 & ~n142 ;
  assign n144 = \d_out_reg[4]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n145 = n68 & n144 ;
  assign n146 = \stato_reg[0]/NET0131  & n134 ;
  assign n147 = ~n145 & ~n146 ;
  assign n148 = \d_in_reg[0]/NET0131  & \d_in_reg[5]/NET0131  ;
  assign n149 = n74 & n148 ;
  assign n150 = ~\d_in_reg[0]/NET0131  & \d_out_reg[5]/NET0131  ;
  assign n151 = n77 & n150 ;
  assign n152 = ~n149 & ~n151 ;
  assign n153 = n147 & n152 ;
  assign n154 = n143 & n153 ;
  assign n155 = \d_in_reg[6]/NET0131  & n62 ;
  assign n156 = ~n60 & n155 ;
  assign n157 = \d_out_reg[5]/NET0131  & n62 ;
  assign n158 = n60 & n157 ;
  assign n159 = ~n156 & ~n158 ;
  assign n160 = \d_out_reg[5]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n161 = n68 & n160 ;
  assign n162 = \stato_reg[0]/NET0131  & n150 ;
  assign n163 = ~n161 & ~n162 ;
  assign n164 = \d_in_reg[0]/NET0131  & \d_in_reg[6]/NET0131  ;
  assign n165 = n74 & n164 ;
  assign n166 = ~\d_in_reg[0]/NET0131  & \d_out_reg[6]/NET0131  ;
  assign n167 = n77 & n166 ;
  assign n168 = ~n165 & ~n167 ;
  assign n169 = n163 & n168 ;
  assign n170 = n159 & n169 ;
  assign n171 = \d_in_reg[7]/NET0131  & n62 ;
  assign n172 = ~n60 & n171 ;
  assign n173 = \d_out_reg[6]/NET0131  & n62 ;
  assign n174 = n60 & n173 ;
  assign n175 = ~n172 & ~n174 ;
  assign n176 = \d_out_reg[6]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n177 = n68 & n176 ;
  assign n178 = \stato_reg[0]/NET0131  & n166 ;
  assign n179 = ~n177 & ~n178 ;
  assign n180 = \d_in_reg[0]/NET0131  & \d_in_reg[7]/NET0131  ;
  assign n181 = n74 & n180 ;
  assign n182 = n77 & n106 ;
  assign n183 = ~n181 & ~n182 ;
  assign n184 = n179 & n183 ;
  assign n185 = n175 & n184 ;
  assign n186 = \d_in_reg[3]/NET0131  & n62 ;
  assign n187 = ~n60 & n186 ;
  assign n188 = \d_out_reg[2]/NET0131  & n62 ;
  assign n189 = n60 & n188 ;
  assign n190 = ~n187 & ~n189 ;
  assign n191 = \d_out_reg[2]/NET0131  & \stato_reg[1]/NET0131  ;
  assign n192 = n68 & n191 ;
  assign n193 = \stato_reg[0]/NET0131  & n94 ;
  assign n194 = ~n192 & ~n193 ;
  assign n195 = n77 & n128 ;
  assign n196 = \d_in_reg[0]/NET0131  & \d_in_reg[3]/NET0131  ;
  assign n197 = n74 & n196 ;
  assign n198 = ~n195 & ~n197 ;
  assign n199 = n194 & n198 ;
  assign n200 = n190 & n199 ;
  assign n201 = ~\d_in_reg[0]/NET0131  & n77 ;
  assign n202 = ~n113 & ~n201 ;
  assign n203 = \stato_reg[1]/NET0131  & ~n201 ;
  assign n204 = n60 & n203 ;
  assign n205 = ~n202 & ~n204 ;
  assign n206 = ~n60 & n62 ;
  assign n207 = ~\d_in_reg[0]/NET0131  & ~y_pad ;
  assign n208 = n74 & ~n207 ;
  assign n209 = n71 & n77 ;
  assign n210 = ~n208 & ~n209 ;
  assign n211 = ~n206 & n210 ;
  assign n212 = \d_in_reg[2]/NET0131  & ~n115 ;
  assign n213 = \d_in_reg[7]/NET0131  & ~n115 ;
  assign n214 = \d_in_reg[8]/NET0131  & ~n115 ;
  assign n215 = \d_in_reg[1]/NET0131  & ~n115 ;
  assign n216 = \d_in_reg[6]/NET0131  & ~n115 ;
  assign n217 = \d_in_reg[3]/NET0131  & ~n115 ;
  assign n218 = \d_in_reg[4]/NET0131  & ~n115 ;
  assign n219 = \d_in_reg[5]/NET0131  & ~n115 ;
  assign n220 = ~\d_in_reg[0]/NET0131  & \old_reg[5]/NET0131  ;
  assign n221 = ~n164 & ~n220 ;
  assign n222 = \stato_reg[0]/NET0131  & ~n221 ;
  assign n223 = \old_reg[5]/NET0131  & n77 ;
  assign n224 = ~n222 & ~n223 ;
  assign n225 = ~\d_in_reg[0]/NET0131  & \old_reg[6]/NET0131  ;
  assign n226 = ~n180 & ~n225 ;
  assign n227 = \stato_reg[0]/NET0131  & ~n226 ;
  assign n228 = \old_reg[6]/NET0131  & n77 ;
  assign n229 = ~n227 & ~n228 ;
  assign n230 = ~\d_in_reg[0]/NET0131  & \old_reg[7]/NET0131  ;
  assign n231 = ~n109 & ~n230 ;
  assign n232 = \stato_reg[0]/NET0131  & ~n231 ;
  assign n233 = \old_reg[7]/NET0131  & n77 ;
  assign n234 = ~n232 & ~n233 ;
  assign n235 = ~\d_in_reg[0]/NET0131  & \old_reg[0]/NET0131  ;
  assign n236 = ~n75 & ~n235 ;
  assign n237 = \stato_reg[0]/NET0131  & ~n236 ;
  assign n238 = \old_reg[0]/NET0131  & n77 ;
  assign n239 = ~n237 & ~n238 ;
  assign n240 = ~\d_in_reg[0]/NET0131  & \old_reg[1]/NET0131  ;
  assign n241 = ~n92 & ~n240 ;
  assign n242 = \stato_reg[0]/NET0131  & ~n241 ;
  assign n243 = \old_reg[1]/NET0131  & n77 ;
  assign n244 = ~n242 & ~n243 ;
  assign n245 = \d_in_reg[3]/NET0131  & n113 ;
  assign n246 = \old_reg[2]/NET0131  & ~n115 ;
  assign n247 = ~n245 & ~n246 ;
  assign n248 = ~\d_in_reg[0]/NET0131  & \old_reg[3]/NET0131  ;
  assign n249 = ~n131 & ~n248 ;
  assign n250 = \stato_reg[0]/NET0131  & ~n249 ;
  assign n251 = \old_reg[3]/NET0131  & n77 ;
  assign n252 = ~n250 & ~n251 ;
  assign n253 = ~\d_in_reg[0]/NET0131  & \old_reg[4]/NET0131  ;
  assign n254 = ~n148 & ~n253 ;
  assign n255 = \stato_reg[0]/NET0131  & ~n254 ;
  assign n256 = \old_reg[4]/NET0131  & n77 ;
  assign n257 = ~n255 & ~n256 ;
  assign n258 = ~\stato_reg[0]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n259 = ~\d_in_reg[0]/NET0131  & ~\stato_reg[1]/NET0131  ;
  assign n260 = ~n258 & ~n259 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g1026/_0_  = ~n82 ;
  assign \g1035/_0_  = ~n98 ;
  assign \g41/_0_  = ~n112 ;
  assign \g708/_0_  = n120 ;
  assign \g709/_0_  = ~n138 ;
  assign \g711/_0_  = ~n154 ;
  assign \g712/_0_  = ~n170 ;
  assign \g714/_0_  = ~n185 ;
  assign \g716/_0_  = ~n200 ;
  assign \g718/_0_  = ~n205 ;
  assign \g728/_0_  = ~n211 ;
  assign \g770/_0_  = n212 ;
  assign \g771/_0_  = n213 ;
  assign \g772/_0_  = n214 ;
  assign \g773/_0_  = n215 ;
  assign \g774/_0_  = n216 ;
  assign \g775/_0_  = n217 ;
  assign \g776/_0_  = n218 ;
  assign \g777/_0_  = n219 ;
  assign \g782/_0_  = ~n224 ;
  assign \g783/_0_  = ~n229 ;
  assign \g784/_0_  = ~n234 ;
  assign \g785/_0_  = ~n239 ;
  assign \g786/_0_  = ~n244 ;
  assign \g787/_0_  = ~n247 ;
  assign \g788/_0_  = ~n252 ;
  assign \g789/_0_  = ~n257 ;
  assign \g806/_0_  = n260 ;
endmodule
