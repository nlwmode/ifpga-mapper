module top (a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad);
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	output l_pad ;
	output m_pad ;
	output n_pad ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w13_ ;
	wire _w14_ ;
	wire _w15_ ;
	wire _w16_ ;
	wire _w17_ ;
	wire _w18_ ;
	wire _w19_ ;
	wire _w20_ ;
	wire _w21_ ;
	wire _w22_ ;
	wire _w23_ ;
	wire _w24_ ;
	wire _w25_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		f_pad,
		g_pad,
		_w13_
	);
	LUT2 #(
		.INIT('h4)
	) name1 (
		j_pad,
		k_pad,
		_w14_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2 (
		h_pad,
		i_pad,
		j_pad,
		k_pad,
		_w15_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name3 (
		f_pad,
		g_pad,
		h_pad,
		i_pad,
		_w16_
	);
	LUT3 #(
		.INIT('h82)
	) name4 (
		b_pad,
		d_pad,
		e_pad,
		_w17_
	);
	LUT4 #(
		.INIT('hba00)
	) name5 (
		_w13_,
		_w15_,
		_w16_,
		_w17_,
		_w18_
	);
	LUT4 #(
		.INIT('h5155)
	) name6 (
		a_pad,
		b_pad,
		d_pad,
		e_pad,
		_w19_
	);
	LUT2 #(
		.INIT('hb)
	) name7 (
		_w18_,
		_w19_,
		_w20_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		j_pad,
		k_pad,
		_w21_
	);
	LUT2 #(
		.INIT('h2)
	) name9 (
		_w16_,
		_w21_,
		_w22_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name10 (
		f_pad,
		g_pad,
		h_pad,
		i_pad,
		_w23_
	);
	LUT3 #(
		.INIT('h40)
	) name11 (
		_w14_,
		_w17_,
		_w23_,
		_w24_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		_w22_,
		_w24_,
		_w25_
	);
	LUT4 #(
		.INIT('h4d44)
	) name13 (
		f_pad,
		g_pad,
		h_pad,
		i_pad,
		_w26_
	);
	LUT4 #(
		.INIT('h00c4)
	) name14 (
		_w16_,
		_w17_,
		_w21_,
		_w26_,
		_w27_
	);
	LUT4 #(
		.INIT('h3313)
	) name15 (
		b_pad,
		c_pad,
		d_pad,
		e_pad,
		_w28_
	);
	LUT2 #(
		.INIT('hb)
	) name16 (
		_w27_,
		_w28_,
		_w29_
	);
	assign l_pad = _w20_ ;
	assign m_pad = _w25_ ;
	assign n_pad = _w29_ ;
endmodule;