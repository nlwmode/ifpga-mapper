module top (\a0_pad , \a1_pad , \a2_pad , \a3_pad , \a4_pad , a_pad, \b0_pad , \b1_pad , \b2_pad , \b3_pad , \b4_pad , b_pad, \c0_pad , \c1_pad , \c2_pad , \c3_pad , \c4_pad , c_pad, \d0_pad , \d1_pad , \d2_pad , \d3_pad , \d4_pad , d_pad, \e0_pad , \e1_pad , \e2_pad , \e3_pad , \e4_pad , e_pad, \f0_pad , \f1_pad , \f2_pad , \f3_pad , \f4_pad , f_pad, \g0_pad , \g1_pad , \g2_pad , \g3_pad , \g4_pad , g_pad, \h0_pad , \h1_pad , \h2_pad , \h3_pad , \h4_pad , h_pad, \i0_pad , \i1_pad , \i2_pad , \i3_pad , \i4_pad , i_pad, \j0_pad , \j1_pad , \j2_pad , \j3_pad , \j4_pad , j_pad, \k0_pad , \k1_pad , \k2_pad , \k3_pad , k_pad, \l0_pad , \l1_pad , \l2_pad , \l3_pad , \l4_pad , l_pad, \m0_pad , \m1_pad , \m2_pad , \m3_pad , \m6_pad , m_pad, \n0_pad , \n1_pad , \n2_pad , \n3_pad , \n4_pad , n_pad, \o0_pad , \o1_pad , \o2_pad , \o3_pad , o_pad, \p0_pad , \p1_pad , \p2_pad , \p3_pad , p_pad, \q0_pad , \q1_pad , \q2_pad , \q3_pad , q_pad, \r1_pad , \r2_pad , \r3_pad , r_pad, \s0_pad , \s1_pad , \s2_pad , \s3_pad , s_pad, \t0_pad , \t1_pad , \t2_pad , \t3_pad , \t4_pad , t_pad, \u0_pad , \u1_pad , \u2_pad , \u4_pad , u_pad, \v0_pad , \v1_pad , \v2_pad , v_pad, \w0_pad , \w1_pad , \w2_pad , \w3_pad , w_pad, \x0_pad , \x1_pad , \x2_pad , \x3_pad , x_pad, \y0_pad , \y1_pad , \y2_pad , \y3_pad , y_pad, \z0_pad , \z1_pad , \z2_pad , \z3_pad , z_pad, \a5_pad , \a6_pad , \a7_pad , \a8_pad , \a9_pad , \b5_pad , \b6_pad , \b7_pad , \b8_pad , \b9_pad , \c5_pad , \c6_pad , \c7_pad , \c8_pad , \c9_pad , \d5_pad , \d6_pad , \d7_pad , \d8_pad , \d9_pad , \e5_pad , \e6_pad , \e7_pad , \e8_pad , \e9_pad , \f5_pad , \f6_pad , \f7_pad , \f8_pad , \f9_pad , \g5_pad , \g6_pad , \g7_pad , \g8_pad , \g9_pad , \h5_pad , \h6_pad , \h7_pad , \h8_pad , \h9_pad , \i5_pad , \i6_pad , \i7_pad , \i8_pad , \i9_pad , \j5_pad , \j6_pad , \j7_pad , \j8_pad , \j9_pad , \k5_pad , \k6_pad , \k7_pad , \k8_pad , \k9_pad , \l5_pad , \l6_pad , \l7_pad , \l8_pad , \l9_pad , \m7_pad , \m8_pad , \m9_pad , \n5_pad , \n6_pad , \n7_pad , \n8_pad , \n9_pad , \o4_pad , \o5_pad , \o6_pad , \o7_pad , \o8_pad , \o9_pad , \p4_pad , \p5_pad , \p6_pad , \p7_pad , \p8_pad , \p9_pad , \q4_pad , \q5_pad , \q6_pad , \q7_pad , \q8_pad , \q9_pad , \r4_pad , \r5_pad , \r6_pad , \r7_pad , \r8_pad , \r9_pad , \s4_pad , \s6_pad , \s7_pad , \s8_pad , \s9_pad , \t6_pad , \t7_pad , \t8_pad , \t9_pad , \u6_pad , \u7_pad , \u8_pad , \u9_pad , \v4_pad , \v6_pad , \v7_pad , \v8_pad , \v9_pad , \w4_pad , \w5_pad , \w6_pad , \w7_pad , \w8_pad , \w9_pad , \x4_pad , \x5_pad , \x6_pad , \x7_pad , \x8_pad , \y4_pad , \y5_pad , \y6_pad , \y7_pad , \y8_pad , \z4_pad , \z5_pad , \z6_pad , \z7_pad , \z8_pad );
	input \a0_pad  ;
	input \a1_pad  ;
	input \a2_pad  ;
	input \a3_pad  ;
	input \a4_pad  ;
	input a_pad ;
	input \b0_pad  ;
	input \b1_pad  ;
	input \b2_pad  ;
	input \b3_pad  ;
	input \b4_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input \c1_pad  ;
	input \c2_pad  ;
	input \c3_pad  ;
	input \c4_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input \d1_pad  ;
	input \d2_pad  ;
	input \d3_pad  ;
	input \d4_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input \e1_pad  ;
	input \e2_pad  ;
	input \e3_pad  ;
	input \e4_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input \f1_pad  ;
	input \f2_pad  ;
	input \f3_pad  ;
	input \f4_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input \g1_pad  ;
	input \g2_pad  ;
	input \g3_pad  ;
	input \g4_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input \h1_pad  ;
	input \h2_pad  ;
	input \h3_pad  ;
	input \h4_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input \i1_pad  ;
	input \i2_pad  ;
	input \i3_pad  ;
	input \i4_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input \j1_pad  ;
	input \j2_pad  ;
	input \j3_pad  ;
	input \j4_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input \k1_pad  ;
	input \k2_pad  ;
	input \k3_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input \l1_pad  ;
	input \l2_pad  ;
	input \l3_pad  ;
	input \l4_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input \m1_pad  ;
	input \m2_pad  ;
	input \m3_pad  ;
	input \m6_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input \n1_pad  ;
	input \n2_pad  ;
	input \n3_pad  ;
	input \n4_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input \o1_pad  ;
	input \o2_pad  ;
	input \o3_pad  ;
	input o_pad ;
	input \p0_pad  ;
	input \p1_pad  ;
	input \p2_pad  ;
	input \p3_pad  ;
	input p_pad ;
	input \q0_pad  ;
	input \q1_pad  ;
	input \q2_pad  ;
	input \q3_pad  ;
	input q_pad ;
	input \r1_pad  ;
	input \r2_pad  ;
	input \r3_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input \s1_pad  ;
	input \s2_pad  ;
	input \s3_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input \t1_pad  ;
	input \t2_pad  ;
	input \t3_pad  ;
	input \t4_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input \u1_pad  ;
	input \u2_pad  ;
	input \u4_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input v_pad ;
	input \w0_pad  ;
	input \w1_pad  ;
	input \w2_pad  ;
	input \w3_pad  ;
	input w_pad ;
	input \x0_pad  ;
	input \x1_pad  ;
	input \x2_pad  ;
	input \x3_pad  ;
	input x_pad ;
	input \y0_pad  ;
	input \y1_pad  ;
	input \y2_pad  ;
	input \y3_pad  ;
	input y_pad ;
	input \z0_pad  ;
	input \z1_pad  ;
	input \z2_pad  ;
	input \z3_pad  ;
	input z_pad ;
	output \a5_pad  ;
	output \a6_pad  ;
	output \a7_pad  ;
	output \a8_pad  ;
	output \a9_pad  ;
	output \b5_pad  ;
	output \b6_pad  ;
	output \b7_pad  ;
	output \b8_pad  ;
	output \b9_pad  ;
	output \c5_pad  ;
	output \c6_pad  ;
	output \c7_pad  ;
	output \c8_pad  ;
	output \c9_pad  ;
	output \d5_pad  ;
	output \d6_pad  ;
	output \d7_pad  ;
	output \d8_pad  ;
	output \d9_pad  ;
	output \e5_pad  ;
	output \e6_pad  ;
	output \e7_pad  ;
	output \e8_pad  ;
	output \e9_pad  ;
	output \f5_pad  ;
	output \f6_pad  ;
	output \f7_pad  ;
	output \f8_pad  ;
	output \f9_pad  ;
	output \g5_pad  ;
	output \g6_pad  ;
	output \g7_pad  ;
	output \g8_pad  ;
	output \g9_pad  ;
	output \h5_pad  ;
	output \h6_pad  ;
	output \h7_pad  ;
	output \h8_pad  ;
	output \h9_pad  ;
	output \i5_pad  ;
	output \i6_pad  ;
	output \i7_pad  ;
	output \i8_pad  ;
	output \i9_pad  ;
	output \j5_pad  ;
	output \j6_pad  ;
	output \j7_pad  ;
	output \j8_pad  ;
	output \j9_pad  ;
	output \k5_pad  ;
	output \k6_pad  ;
	output \k7_pad  ;
	output \k8_pad  ;
	output \k9_pad  ;
	output \l5_pad  ;
	output \l6_pad  ;
	output \l7_pad  ;
	output \l8_pad  ;
	output \l9_pad  ;
	output \m7_pad  ;
	output \m8_pad  ;
	output \m9_pad  ;
	output \n5_pad  ;
	output \n6_pad  ;
	output \n7_pad  ;
	output \n8_pad  ;
	output \n9_pad  ;
	output \o4_pad  ;
	output \o5_pad  ;
	output \o6_pad  ;
	output \o7_pad  ;
	output \o8_pad  ;
	output \o9_pad  ;
	output \p4_pad  ;
	output \p5_pad  ;
	output \p6_pad  ;
	output \p7_pad  ;
	output \p8_pad  ;
	output \p9_pad  ;
	output \q4_pad  ;
	output \q5_pad  ;
	output \q6_pad  ;
	output \q7_pad  ;
	output \q8_pad  ;
	output \q9_pad  ;
	output \r4_pad  ;
	output \r5_pad  ;
	output \r6_pad  ;
	output \r7_pad  ;
	output \r8_pad  ;
	output \r9_pad  ;
	output \s4_pad  ;
	output \s6_pad  ;
	output \s7_pad  ;
	output \s8_pad  ;
	output \s9_pad  ;
	output \t6_pad  ;
	output \t7_pad  ;
	output \t8_pad  ;
	output \t9_pad  ;
	output \u6_pad  ;
	output \u7_pad  ;
	output \u8_pad  ;
	output \u9_pad  ;
	output \v4_pad  ;
	output \v6_pad  ;
	output \v7_pad  ;
	output \v8_pad  ;
	output \v9_pad  ;
	output \w4_pad  ;
	output \w5_pad  ;
	output \w6_pad  ;
	output \w7_pad  ;
	output \w8_pad  ;
	output \w9_pad  ;
	output \x4_pad  ;
	output \x5_pad  ;
	output \x6_pad  ;
	output \x7_pad  ;
	output \x8_pad  ;
	output \y4_pad  ;
	output \y5_pad  ;
	output \y6_pad  ;
	output \y7_pad  ;
	output \y8_pad  ;
	output \z4_pad  ;
	output \z5_pad  ;
	output \z6_pad  ;
	output \z7_pad  ;
	output \z8_pad  ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w526_ ;
	wire _w525_ ;
	wire _w524_ ;
	wire _w523_ ;
	wire _w522_ ;
	wire _w521_ ;
	wire _w520_ ;
	wire _w519_ ;
	wire _w518_ ;
	wire _w517_ ;
	wire _w516_ ;
	wire _w515_ ;
	wire _w514_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w270_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w162_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w167_ ;
	wire _w40_ ;
	wire _w297_ ;
	wire _w157_ ;
	wire _w163_ ;
	wire _w151_ ;
	wire _w170_ ;
	wire _w179_ ;
	wire _w161_ ;
	wire _w192_ ;
	wire _w152_ ;
	wire _w150_ ;
	wire _w153_ ;
	wire _w154_ ;
	wire _w186_ ;
	wire _w155_ ;
	wire _w156_ ;
	wire _w173_ ;
	wire _w47_ ;
	wire _w304_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w180_ ;
	wire _w54_ ;
	wire _w311_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w187_ ;
	wire _w61_ ;
	wire _w318_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w68_ ;
	wire _w325_ ;
	wire _w195_ ;
	wire _w196_ ;
	wire _w197_ ;
	wire _w198_ ;
	wire _w199_ ;
	wire _w200_ ;
	wire _w74_ ;
	wire _w331_ ;
	wire _w201_ ;
	wire _w202_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	wire _w394_ ;
	wire _w395_ ;
	wire _w396_ ;
	wire _w397_ ;
	wire _w398_ ;
	wire _w399_ ;
	wire _w400_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\g1_pad ,
		_w40_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\h1_pad ,
		_w47_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\i1_pad ,
		_w54_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\j1_pad ,
		_w61_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\k1_pad ,
		_w68_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\l1_pad ,
		_w74_
	);
	LUT2 #(
		.INIT('h9)
	) name6 (
		\k0_pad ,
		\l0_pad ,
		_w150_
	);
	LUT3 #(
		.INIT('h41)
	) name7 (
		\j3_pad ,
		\k0_pad ,
		\l0_pad ,
		_w151_
	);
	LUT4 #(
		.INIT('hf090)
	) name8 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		\r3_pad ,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT3 #(
		.INIT('hf7)
	) name10 (
		\k1_pad ,
		\m1_pad ,
		\m6_pad ,
		_w154_
	);
	LUT2 #(
		.INIT('h2)
	) name11 (
		\o0_pad ,
		\q0_pad ,
		_w155_
	);
	LUT3 #(
		.INIT('h01)
	) name12 (
		\j1_pad ,
		\k1_pad ,
		\l1_pad ,
		_w156_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		\h1_pad ,
		\i1_pad ,
		_w157_
	);
	LUT3 #(
		.INIT('h40)
	) name14 (
		\n0_pad ,
		_w156_,
		_w157_,
		_w158_
	);
	LUT4 #(
		.INIT('h2000)
	) name15 (
		\f0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w159_
	);
	LUT2 #(
		.INIT('h8)
	) name16 (
		\y3_pad ,
		\z3_pad ,
		_w160_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\a4_pad ,
		\b4_pad ,
		_w161_
	);
	LUT3 #(
		.INIT('h01)
	) name18 (
		\a4_pad ,
		\b4_pad ,
		\c4_pad ,
		_w162_
	);
	LUT4 #(
		.INIT('h8aaa)
	) name19 (
		\l4_pad ,
		\x3_pad ,
		_w160_,
		_w162_,
		_w163_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name20 (
		\r1_pad ,
		\s1_pad ,
		_w158_,
		_w163_,
		_w164_
	);
	LUT3 #(
		.INIT('ha8)
	) name21 (
		_w155_,
		_w159_,
		_w164_,
		_w165_
	);
	LUT4 #(
		.INIT('h1000)
	) name22 (
		\m0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w166_
	);
	LUT4 #(
		.INIT('haea2)
	) name23 (
		h_pad,
		\k0_pad ,
		\l0_pad ,
		p_pad,
		_w167_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w166_,
		_w167_,
		_w168_
	);
	LUT4 #(
		.INIT('h00ca)
	) name25 (
		\r2_pad ,
		\s2_pad ,
		_w163_,
		_w166_,
		_w169_
	);
	LUT3 #(
		.INIT('ha8)
	) name26 (
		_w155_,
		_w168_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		\e4_pad ,
		\f4_pad ,
		_w171_
	);
	LUT3 #(
		.INIT('h08)
	) name28 (
		\e4_pad ,
		\f4_pad ,
		\g4_pad ,
		_w172_
	);
	LUT4 #(
		.INIT('h0008)
	) name29 (
		\e4_pad ,
		\f4_pad ,
		\g4_pad ,
		\h4_pad ,
		_w173_
	);
	LUT4 #(
		.INIT('hf531)
	) name30 (
		\h1_pad ,
		\j1_pad ,
		\x0_pad ,
		\z0_pad ,
		_w174_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\a1_pad ,
		\k1_pad ,
		_w175_
	);
	LUT4 #(
		.INIT('haf23)
	) name32 (
		\b1_pad ,
		\i1_pad ,
		\l1_pad ,
		\y0_pad ,
		_w176_
	);
	LUT3 #(
		.INIT('h40)
	) name33 (
		_w175_,
		_w174_,
		_w176_,
		_w177_
	);
	LUT4 #(
		.INIT('h4555)
	) name34 (
		_w173_,
		_w175_,
		_w174_,
		_w176_,
		_w178_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		\m6_pad ,
		_w178_,
		_w179_
	);
	LUT3 #(
		.INIT('h17)
	) name36 (
		\j1_pad ,
		\k1_pad ,
		\l1_pad ,
		_w180_
	);
	LUT4 #(
		.INIT('h6160)
	) name37 (
		\h1_pad ,
		\i1_pad ,
		_w156_,
		_w180_,
		_w181_
	);
	LUT4 #(
		.INIT('h2000)
	) name38 (
		\m6_pad ,
		\s3_pad ,
		_w178_,
		_w181_,
		_w182_
	);
	LUT4 #(
		.INIT('h1333)
	) name39 (
		\m6_pad ,
		\r3_pad ,
		_w178_,
		_w181_,
		_w183_
	);
	LUT3 #(
		.INIT('h02)
	) name40 (
		_w155_,
		_w183_,
		_w182_,
		_w184_
	);
	LUT3 #(
		.INIT('h21)
	) name41 (
		\k0_pad ,
		\k3_pad ,
		\l0_pad ,
		_w185_
	);
	LUT4 #(
		.INIT('hf090)
	) name42 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		\s3_pad ,
		_w186_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w185_,
		_w186_,
		_w187_
	);
	LUT3 #(
		.INIT('hf7)
	) name44 (
		\l1_pad ,
		\m1_pad ,
		\m6_pad ,
		_w188_
	);
	LUT4 #(
		.INIT('h2000)
	) name45 (
		\e0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w189_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name46 (
		\s1_pad ,
		\t1_pad ,
		_w158_,
		_w163_,
		_w190_
	);
	LUT3 #(
		.INIT('ha8)
	) name47 (
		_w155_,
		_w189_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w150_,
		_w166_,
		_w192_
	);
	LUT3 #(
		.INIT('hca)
	) name49 (
		\s2_pad ,
		\t2_pad ,
		_w163_,
		_w193_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name50 (
		i_pad,
		_w150_,
		_w155_,
		_w166_,
		_w194_
	);
	LUT3 #(
		.INIT('he0)
	) name51 (
		_w192_,
		_w193_,
		_w194_,
		_w195_
	);
	LUT4 #(
		.INIT('h2000)
	) name52 (
		\m6_pad ,
		\t3_pad ,
		_w178_,
		_w181_,
		_w196_
	);
	LUT4 #(
		.INIT('h1333)
	) name53 (
		\m6_pad ,
		\s3_pad ,
		_w178_,
		_w181_,
		_w197_
	);
	LUT3 #(
		.INIT('h02)
	) name54 (
		_w155_,
		_w197_,
		_w196_,
		_w198_
	);
	LUT3 #(
		.INIT('h09)
	) name55 (
		\k0_pad ,
		\l0_pad ,
		\l3_pad ,
		_w199_
	);
	LUT4 #(
		.INIT('hf090)
	) name56 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		\t3_pad ,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		_w199_,
		_w200_,
		_w201_
	);
	LUT2 #(
		.INIT('h7)
	) name58 (
		\h1_pad ,
		\l4_pad ,
		_w202_
	);
	LUT4 #(
		.INIT('h2000)
	) name59 (
		\d0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w203_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name60 (
		\t1_pad ,
		\u1_pad ,
		_w158_,
		_w163_,
		_w204_
	);
	LUT3 #(
		.INIT('ha8)
	) name61 (
		_w155_,
		_w203_,
		_w204_,
		_w205_
	);
	LUT3 #(
		.INIT('hca)
	) name62 (
		\t2_pad ,
		\u2_pad ,
		_w163_,
		_w206_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name63 (
		j_pad,
		_w150_,
		_w155_,
		_w166_,
		_w207_
	);
	LUT3 #(
		.INIT('he0)
	) name64 (
		_w192_,
		_w206_,
		_w207_,
		_w208_
	);
	LUT4 #(
		.INIT('h2000)
	) name65 (
		\m6_pad ,
		\t4_pad ,
		_w178_,
		_w181_,
		_w209_
	);
	LUT4 #(
		.INIT('h1333)
	) name66 (
		\m6_pad ,
		\t3_pad ,
		_w178_,
		_w181_,
		_w210_
	);
	LUT3 #(
		.INIT('h02)
	) name67 (
		_w155_,
		_w210_,
		_w209_,
		_w211_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\m0_pad ,
		\m3_pad ,
		_w212_
	);
	LUT2 #(
		.INIT('h7)
	) name69 (
		\i1_pad ,
		\l4_pad ,
		_w213_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		_w155_,
		_w166_,
		_w214_
	);
	LUT4 #(
		.INIT('h0305)
	) name71 (
		\u1_pad ,
		\v1_pad ,
		_w158_,
		_w163_,
		_w215_
	);
	LUT2 #(
		.INIT('h2)
	) name72 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT3 #(
		.INIT('hca)
	) name73 (
		\u2_pad ,
		\v2_pad ,
		_w163_,
		_w217_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name74 (
		k_pad,
		_w150_,
		_w155_,
		_w166_,
		_w218_
	);
	LUT3 #(
		.INIT('he0)
	) name75 (
		_w192_,
		_w217_,
		_w218_,
		_w219_
	);
	LUT4 #(
		.INIT('h2000)
	) name76 (
		\m6_pad ,
		\u4_pad ,
		_w178_,
		_w181_,
		_w220_
	);
	LUT4 #(
		.INIT('h1333)
	) name77 (
		\m6_pad ,
		\t4_pad ,
		_w178_,
		_w181_,
		_w221_
	);
	LUT3 #(
		.INIT('h02)
	) name78 (
		_w155_,
		_w221_,
		_w220_,
		_w222_
	);
	LUT2 #(
		.INIT('h8)
	) name79 (
		\m0_pad ,
		\n3_pad ,
		_w223_
	);
	LUT2 #(
		.INIT('h7)
	) name80 (
		\j1_pad ,
		\l4_pad ,
		_w224_
	);
	LUT4 #(
		.INIT('h0305)
	) name81 (
		\v1_pad ,
		\w1_pad ,
		_w158_,
		_w163_,
		_w225_
	);
	LUT4 #(
		.INIT('h1000)
	) name82 (
		\k0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w226_
	);
	LUT2 #(
		.INIT('h2)
	) name83 (
		_w155_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name84 (
		_w225_,
		_w227_,
		_w228_
	);
	LUT3 #(
		.INIT('hca)
	) name85 (
		\v2_pad ,
		\w2_pad ,
		_w163_,
		_w229_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name86 (
		l_pad,
		_w150_,
		_w155_,
		_w166_,
		_w230_
	);
	LUT3 #(
		.INIT('he0)
	) name87 (
		_w192_,
		_w229_,
		_w230_,
		_w231_
	);
	LUT4 #(
		.INIT('h2000)
	) name88 (
		\m6_pad ,
		\w3_pad ,
		_w178_,
		_w181_,
		_w232_
	);
	LUT4 #(
		.INIT('h1333)
	) name89 (
		\m6_pad ,
		\u4_pad ,
		_w178_,
		_w181_,
		_w233_
	);
	LUT3 #(
		.INIT('h02)
	) name90 (
		_w155_,
		_w233_,
		_w232_,
		_w234_
	);
	LUT2 #(
		.INIT('h8)
	) name91 (
		\m0_pad ,
		\o3_pad ,
		_w235_
	);
	LUT2 #(
		.INIT('h7)
	) name92 (
		\k1_pad ,
		\l4_pad ,
		_w236_
	);
	LUT4 #(
		.INIT('h0305)
	) name93 (
		\w1_pad ,
		\x1_pad ,
		_w158_,
		_w163_,
		_w237_
	);
	LUT4 #(
		.INIT('h1000)
	) name94 (
		\l0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w238_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w155_,
		_w238_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w237_,
		_w239_,
		_w240_
	);
	LUT3 #(
		.INIT('hca)
	) name97 (
		\w2_pad ,
		\x2_pad ,
		_w163_,
		_w241_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name98 (
		m_pad,
		_w150_,
		_w155_,
		_w166_,
		_w242_
	);
	LUT3 #(
		.INIT('he0)
	) name99 (
		_w192_,
		_w241_,
		_w242_,
		_w243_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name100 (
		\m6_pad ,
		\w3_pad ,
		_w178_,
		_w181_,
		_w244_
	);
	LUT3 #(
		.INIT('h20)
	) name101 (
		\h1_pad ,
		\i1_pad ,
		\s0_pad ,
		_w245_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		_w156_,
		_w245_,
		_w246_
	);
	LUT4 #(
		.INIT('h0100)
	) name103 (
		\j1_pad ,
		\k1_pad ,
		\l1_pad ,
		\t0_pad ,
		_w247_
	);
	LUT2 #(
		.INIT('h2)
	) name104 (
		\i1_pad ,
		_w247_,
		_w248_
	);
	LUT4 #(
		.INIT('h8acf)
	) name105 (
		\j1_pad ,
		\l1_pad ,
		\u0_pad ,
		\w0_pad ,
		_w249_
	);
	LUT3 #(
		.INIT('h32)
	) name106 (
		\j1_pad ,
		\k1_pad ,
		\l1_pad ,
		_w250_
	);
	LUT4 #(
		.INIT('h0400)
	) name107 (
		\j1_pad ,
		\k1_pad ,
		\l1_pad ,
		\v0_pad ,
		_w251_
	);
	LUT4 #(
		.INIT('h1011)
	) name108 (
		\i1_pad ,
		_w251_,
		_w249_,
		_w250_,
		_w252_
	);
	LUT4 #(
		.INIT('h3332)
	) name109 (
		\h1_pad ,
		_w246_,
		_w252_,
		_w248_,
		_w253_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name110 (
		_w155_,
		_w179_,
		_w244_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\m0_pad ,
		\p3_pad ,
		_w255_
	);
	LUT2 #(
		.INIT('h7)
	) name112 (
		\l1_pad ,
		\l4_pad ,
		_w256_
	);
	LUT4 #(
		.INIT('h4000)
	) name113 (
		\n0_pad ,
		q_pad,
		_w156_,
		_w157_,
		_w257_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name114 (
		\x1_pad ,
		\y1_pad ,
		_w158_,
		_w163_,
		_w258_
	);
	LUT3 #(
		.INIT('ha8)
	) name115 (
		_w155_,
		_w257_,
		_w258_,
		_w259_
	);
	LUT3 #(
		.INIT('hca)
	) name116 (
		\x2_pad ,
		\y2_pad ,
		_w163_,
		_w260_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name117 (
		n_pad,
		_w150_,
		_w155_,
		_w166_,
		_w261_
	);
	LUT3 #(
		.INIT('he0)
	) name118 (
		_w192_,
		_w260_,
		_w261_,
		_w262_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name119 (
		\n0_pad ,
		_w155_,
		_w156_,
		_w157_,
		_w263_
	);
	LUT2 #(
		.INIT('h2)
	) name120 (
		\l4_pad ,
		\x3_pad ,
		_w264_
	);
	LUT4 #(
		.INIT('hb999)
	) name121 (
		\l4_pad ,
		\x3_pad ,
		_w160_,
		_w162_,
		_w265_
	);
	LUT2 #(
		.INIT('h2)
	) name122 (
		_w263_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\m0_pad ,
		\q3_pad ,
		_w267_
	);
	LUT4 #(
		.INIT('h4000)
	) name124 (
		\n0_pad ,
		r_pad,
		_w156_,
		_w157_,
		_w268_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name125 (
		\y1_pad ,
		\z1_pad ,
		_w158_,
		_w163_,
		_w269_
	);
	LUT3 #(
		.INIT('ha8)
	) name126 (
		_w155_,
		_w268_,
		_w269_,
		_w270_
	);
	LUT3 #(
		.INIT('hca)
	) name127 (
		\y2_pad ,
		\z2_pad ,
		_w163_,
		_w271_
	);
	LUT4 #(
		.INIT('hb0f0)
	) name128 (
		o_pad,
		_w150_,
		_w155_,
		_w166_,
		_w272_
	);
	LUT3 #(
		.INIT('he0)
	) name129 (
		_w192_,
		_w271_,
		_w272_,
		_w273_
	);
	LUT4 #(
		.INIT('hd5aa)
	) name130 (
		\y3_pad ,
		\z3_pad ,
		_w162_,
		_w264_,
		_w274_
	);
	LUT2 #(
		.INIT('hd)
	) name131 (
		_w263_,
		_w274_,
		_w275_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\m0_pad ,
		\r3_pad ,
		_w276_
	);
	LUT4 #(
		.INIT('h4000)
	) name133 (
		\n0_pad ,
		s_pad,
		_w156_,
		_w157_,
		_w277_
	);
	LUT4 #(
		.INIT('h0a0c)
	) name134 (
		\a2_pad ,
		\z1_pad ,
		_w158_,
		_w163_,
		_w278_
	);
	LUT3 #(
		.INIT('ha8)
	) name135 (
		_w155_,
		_w277_,
		_w278_,
		_w279_
	);
	LUT3 #(
		.INIT('h80)
	) name136 (
		p_pad,
		_w150_,
		_w166_,
		_w280_
	);
	LUT4 #(
		.INIT('h020a)
	) name137 (
		\z2_pad ,
		_w150_,
		_w163_,
		_w166_,
		_w281_
	);
	LUT3 #(
		.INIT('ha8)
	) name138 (
		_w155_,
		_w280_,
		_w281_,
		_w282_
	);
	LUT4 #(
		.INIT('h2000)
	) name139 (
		\l4_pad ,
		\x3_pad ,
		\y3_pad ,
		\z3_pad ,
		_w283_
	);
	LUT4 #(
		.INIT('he6cc)
	) name140 (
		\y3_pad ,
		\z3_pad ,
		_w162_,
		_w264_,
		_w284_
	);
	LUT2 #(
		.INIT('hd)
	) name141 (
		_w263_,
		_w284_,
		_w285_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\m0_pad ,
		\s3_pad ,
		_w286_
	);
	LUT4 #(
		.INIT('h4000)
	) name143 (
		\n0_pad ,
		t_pad,
		_w156_,
		_w157_,
		_w287_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name144 (
		\a2_pad ,
		\b2_pad ,
		_w158_,
		_w163_,
		_w288_
	);
	LUT3 #(
		.INIT('ha8)
	) name145 (
		_w155_,
		_w287_,
		_w288_,
		_w289_
	);
	LUT4 #(
		.INIT('h4000)
	) name146 (
		\b3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w290_
	);
	LUT4 #(
		.INIT('h1555)
	) name147 (
		\a3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w291_
	);
	LUT3 #(
		.INIT('h02)
	) name148 (
		_w155_,
		_w291_,
		_w290_,
		_w292_
	);
	LUT2 #(
		.INIT('h4)
	) name149 (
		_w150_,
		_w166_,
		_w293_
	);
	LUT3 #(
		.INIT('h10)
	) name150 (
		\a4_pad ,
		_w162_,
		_w283_,
		_w294_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		\a4_pad ,
		_w283_,
		_w295_
	);
	LUT4 #(
		.INIT('haaa8)
	) name152 (
		_w155_,
		_w158_,
		_w294_,
		_w295_,
		_w296_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w293_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\m0_pad ,
		\t3_pad ,
		_w298_
	);
	LUT4 #(
		.INIT('h4000)
	) name155 (
		\n0_pad ,
		u_pad,
		_w156_,
		_w157_,
		_w299_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name156 (
		\b2_pad ,
		\c2_pad ,
		_w158_,
		_w163_,
		_w300_
	);
	LUT3 #(
		.INIT('ha8)
	) name157 (
		_w155_,
		_w299_,
		_w300_,
		_w301_
	);
	LUT4 #(
		.INIT('h4000)
	) name158 (
		\c3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w302_
	);
	LUT4 #(
		.INIT('h1555)
	) name159 (
		\b3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w303_
	);
	LUT3 #(
		.INIT('h02)
	) name160 (
		_w155_,
		_w303_,
		_w302_,
		_w304_
	);
	LUT4 #(
		.INIT('h88cc)
	) name161 (
		\a4_pad ,
		\b4_pad ,
		\c4_pad ,
		_w283_,
		_w305_
	);
	LUT3 #(
		.INIT('h80)
	) name162 (
		\c4_pad ,
		_w161_,
		_w283_,
		_w306_
	);
	LUT3 #(
		.INIT('h01)
	) name163 (
		_w158_,
		_w305_,
		_w306_,
		_w307_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		_w214_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h2)
	) name165 (
		\g1_pad ,
		\j4_pad ,
		_w309_
	);
	LUT4 #(
		.INIT('h4000)
	) name166 (
		\n0_pad ,
		v_pad,
		_w156_,
		_w157_,
		_w310_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name167 (
		\c2_pad ,
		\d2_pad ,
		_w158_,
		_w163_,
		_w311_
	);
	LUT3 #(
		.INIT('ha8)
	) name168 (
		_w155_,
		_w310_,
		_w311_,
		_w312_
	);
	LUT4 #(
		.INIT('h4000)
	) name169 (
		\d3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w313_
	);
	LUT4 #(
		.INIT('h1555)
	) name170 (
		\c3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w314_
	);
	LUT3 #(
		.INIT('h02)
	) name171 (
		_w155_,
		_w314_,
		_w313_,
		_w315_
	);
	LUT4 #(
		.INIT('hcfc5)
	) name172 (
		\c4_pad ,
		\m0_pad ,
		_w158_,
		_w306_,
		_w316_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		_w155_,
		_w316_,
		_w317_
	);
	LUT4 #(
		.INIT('h4000)
	) name174 (
		\n0_pad ,
		w_pad,
		_w156_,
		_w157_,
		_w318_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name175 (
		\d2_pad ,
		\e2_pad ,
		_w158_,
		_w163_,
		_w319_
	);
	LUT3 #(
		.INIT('ha8)
	) name176 (
		_w155_,
		_w318_,
		_w319_,
		_w320_
	);
	LUT4 #(
		.INIT('h4000)
	) name177 (
		\e3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w321_
	);
	LUT4 #(
		.INIT('h1555)
	) name178 (
		\d3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w322_
	);
	LUT3 #(
		.INIT('h02)
	) name179 (
		_w155_,
		_w322_,
		_w321_,
		_w323_
	);
	LUT4 #(
		.INIT('h1000)
	) name180 (
		\n0_pad ,
		\q0_pad ,
		_w156_,
		_w157_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		\g1_pad ,
		\q0_pad ,
		_w325_
	);
	LUT4 #(
		.INIT('h6a00)
	) name182 (
		\d4_pad ,
		\m6_pad ,
		_w178_,
		_w325_,
		_w326_
	);
	LUT3 #(
		.INIT('ha8)
	) name183 (
		\o0_pad ,
		_w324_,
		_w326_,
		_w327_
	);
	LUT3 #(
		.INIT('hfd)
	) name184 (
		\h1_pad ,
		\m6_pad ,
		\n0_pad ,
		_w328_
	);
	LUT2 #(
		.INIT('h6)
	) name185 (
		\f1_pad ,
		\i4_pad ,
		_w329_
	);
	LUT2 #(
		.INIT('h9)
	) name186 (
		\f1_pad ,
		\i4_pad ,
		_w330_
	);
	LUT4 #(
		.INIT('h4000)
	) name187 (
		\n0_pad ,
		x_pad,
		_w156_,
		_w157_,
		_w331_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name188 (
		\e2_pad ,
		\f2_pad ,
		_w158_,
		_w163_,
		_w332_
	);
	LUT3 #(
		.INIT('ha8)
	) name189 (
		_w155_,
		_w331_,
		_w332_,
		_w333_
	);
	LUT4 #(
		.INIT('h4000)
	) name190 (
		\f3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w334_
	);
	LUT4 #(
		.INIT('h1555)
	) name191 (
		\e3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w335_
	);
	LUT3 #(
		.INIT('h02)
	) name192 (
		_w155_,
		_w335_,
		_w334_,
		_w336_
	);
	LUT4 #(
		.INIT('h4000)
	) name193 (
		\d4_pad ,
		\e4_pad ,
		\m6_pad ,
		_w178_,
		_w337_
	);
	LUT4 #(
		.INIT('h4555)
	) name194 (
		\d4_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w338_
	);
	LUT4 #(
		.INIT('h1555)
	) name195 (
		\e4_pad ,
		\m6_pad ,
		_w178_,
		_w338_,
		_w339_
	);
	LUT3 #(
		.INIT('h04)
	) name196 (
		\g1_pad ,
		\o0_pad ,
		\q0_pad ,
		_w340_
	);
	LUT4 #(
		.INIT('hbf00)
	) name197 (
		\n0_pad ,
		_w156_,
		_w157_,
		_w340_,
		_w341_
	);
	LUT3 #(
		.INIT('h1f)
	) name198 (
		_w337_,
		_w339_,
		_w341_,
		_w342_
	);
	LUT3 #(
		.INIT('hfd)
	) name199 (
		\i1_pad ,
		\m6_pad ,
		\n0_pad ,
		_w343_
	);
	LUT3 #(
		.INIT('h80)
	) name200 (
		\x3_pad ,
		_w160_,
		_w162_,
		_w344_
	);
	LUT4 #(
		.INIT('h4000)
	) name201 (
		\n0_pad ,
		y_pad,
		_w156_,
		_w157_,
		_w345_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name202 (
		\f2_pad ,
		\g2_pad ,
		_w158_,
		_w163_,
		_w346_
	);
	LUT3 #(
		.INIT('ha8)
	) name203 (
		_w155_,
		_w345_,
		_w346_,
		_w347_
	);
	LUT4 #(
		.INIT('h4000)
	) name204 (
		\g3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w348_
	);
	LUT4 #(
		.INIT('h1555)
	) name205 (
		\f3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w349_
	);
	LUT3 #(
		.INIT('h02)
	) name206 (
		_w155_,
		_w349_,
		_w348_,
		_w350_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		\e4_pad ,
		\f4_pad ,
		_w351_
	);
	LUT4 #(
		.INIT('h8000)
	) name208 (
		\m6_pad ,
		_w178_,
		_w338_,
		_w351_,
		_w352_
	);
	LUT4 #(
		.INIT('hff2f)
	) name209 (
		\f4_pad ,
		_w337_,
		_w341_,
		_w352_,
		_w353_
	);
	LUT4 #(
		.INIT('hbe82)
	) name210 (
		\d3_pad ,
		\k0_pad ,
		\l0_pad ,
		\l3_pad ,
		_w354_
	);
	LUT3 #(
		.INIT('he4)
	) name211 (
		\m0_pad ,
		\t3_pad ,
		_w354_,
		_w355_
	);
	LUT3 #(
		.INIT('hfd)
	) name212 (
		\j1_pad ,
		\m6_pad ,
		\n0_pad ,
		_w356_
	);
	LUT2 #(
		.INIT('h2)
	) name213 (
		\n4_pad ,
		_w173_,
		_w357_
	);
	LUT2 #(
		.INIT('h2)
	) name214 (
		\d4_pad ,
		\g1_pad ,
		_w358_
	);
	LUT2 #(
		.INIT('h8)
	) name215 (
		_w173_,
		_w358_,
		_w359_
	);
	LUT4 #(
		.INIT('haa80)
	) name216 (
		_w155_,
		_w177_,
		_w357_,
		_w359_,
		_w360_
	);
	LUT4 #(
		.INIT('h4000)
	) name217 (
		\n0_pad ,
		z_pad,
		_w156_,
		_w157_,
		_w361_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name218 (
		\g2_pad ,
		\h2_pad ,
		_w158_,
		_w163_,
		_w362_
	);
	LUT3 #(
		.INIT('ha8)
	) name219 (
		_w155_,
		_w361_,
		_w362_,
		_w363_
	);
	LUT4 #(
		.INIT('h4000)
	) name220 (
		\h3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w364_
	);
	LUT4 #(
		.INIT('h1555)
	) name221 (
		\g3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w365_
	);
	LUT3 #(
		.INIT('h02)
	) name222 (
		_w155_,
		_w365_,
		_w364_,
		_w366_
	);
	LUT4 #(
		.INIT('h8000)
	) name223 (
		\m6_pad ,
		_w171_,
		_w178_,
		_w338_,
		_w367_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\g4_pad ,
		_w341_,
		_w368_
	);
	LUT3 #(
		.INIT('h60)
	) name225 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		_w369_
	);
	LUT4 #(
		.INIT('h4000)
	) name226 (
		\n0_pad ,
		_w155_,
		_w156_,
		_w157_,
		_w370_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w369_,
		_w370_,
		_w371_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		\g1_pad ,
		\m6_pad ,
		_w372_
	);
	LUT3 #(
		.INIT('h10)
	) name229 (
		\d4_pad ,
		\g1_pad ,
		\m6_pad ,
		_w373_
	);
	LUT2 #(
		.INIT('h8)
	) name230 (
		_w172_,
		_w373_,
		_w374_
	);
	LUT3 #(
		.INIT('h80)
	) name231 (
		_w178_,
		_w263_,
		_w374_,
		_w375_
	);
	LUT4 #(
		.INIT('hefee)
	) name232 (
		_w371_,
		_w375_,
		_w367_,
		_w368_,
		_w376_
	);
	LUT4 #(
		.INIT('hb8e2)
	) name233 (
		\c3_pad ,
		\k0_pad ,
		\k3_pad ,
		\l0_pad ,
		_w377_
	);
	LUT3 #(
		.INIT('he4)
	) name234 (
		\m0_pad ,
		\s3_pad ,
		_w377_,
		_w378_
	);
	LUT3 #(
		.INIT('hfd)
	) name235 (
		\k1_pad ,
		\m6_pad ,
		\n0_pad ,
		_w379_
	);
	LUT4 #(
		.INIT('h0040)
	) name236 (
		\g1_pad ,
		\h1_pad ,
		\o0_pad ,
		\q0_pad ,
		_w380_
	);
	LUT4 #(
		.INIT('h1000)
	) name237 (
		\e1_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name238 (
		\c1_pad ,
		\d1_pad ,
		_w382_
	);
	LUT4 #(
		.INIT('h0010)
	) name239 (
		\c1_pad ,
		\d1_pad ,
		\o0_pad ,
		\q0_pad ,
		_w383_
	);
	LUT3 #(
		.INIT('hea)
	) name240 (
		_w380_,
		_w381_,
		_w383_,
		_w384_
	);
	LUT4 #(
		.INIT('h2000)
	) name241 (
		\a0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w385_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name242 (
		\h2_pad ,
		\i2_pad ,
		_w158_,
		_w163_,
		_w386_
	);
	LUT3 #(
		.INIT('ha8)
	) name243 (
		_w155_,
		_w385_,
		_w386_,
		_w387_
	);
	LUT4 #(
		.INIT('h4000)
	) name244 (
		\i3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w388_
	);
	LUT4 #(
		.INIT('h1555)
	) name245 (
		\h3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w389_
	);
	LUT3 #(
		.INIT('h02)
	) name246 (
		_w155_,
		_w389_,
		_w388_,
		_w390_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		\m0_pad ,
		_w370_,
		_w391_
	);
	LUT2 #(
		.INIT('h8)
	) name248 (
		\h4_pad ,
		_w341_,
		_w392_
	);
	LUT4 #(
		.INIT('hfbf0)
	) name249 (
		\g4_pad ,
		_w367_,
		_w391_,
		_w392_,
		_w393_
	);
	LUT4 #(
		.INIT('hacca)
	) name250 (
		\b3_pad ,
		\j3_pad ,
		\k0_pad ,
		\l0_pad ,
		_w394_
	);
	LUT3 #(
		.INIT('he4)
	) name251 (
		\m0_pad ,
		\r3_pad ,
		_w394_,
		_w395_
	);
	LUT3 #(
		.INIT('hfd)
	) name252 (
		\l1_pad ,
		\m6_pad ,
		\n0_pad ,
		_w396_
	);
	LUT3 #(
		.INIT('he0)
	) name253 (
		\c1_pad ,
		\d1_pad ,
		\e1_pad ,
		_w397_
	);
	LUT4 #(
		.INIT('h0040)
	) name254 (
		\n0_pad ,
		_w156_,
		_w157_,
		_w397_,
		_w398_
	);
	LUT3 #(
		.INIT('h04)
	) name255 (
		\g1_pad ,
		\i1_pad ,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name256 (
		\c1_pad ,
		\d1_pad ,
		_w400_
	);
	LUT2 #(
		.INIT('h8)
	) name257 (
		_w381_,
		_w400_,
		_w401_
	);
	LUT3 #(
		.INIT('ha8)
	) name258 (
		_w155_,
		_w399_,
		_w401_,
		_w402_
	);
	LUT4 #(
		.INIT('h2000)
	) name259 (
		\b0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w403_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name260 (
		\i2_pad ,
		\j2_pad ,
		_w158_,
		_w163_,
		_w404_
	);
	LUT3 #(
		.INIT('ha8)
	) name261 (
		_w155_,
		_w403_,
		_w404_,
		_w405_
	);
	LUT4 #(
		.INIT('h4000)
	) name262 (
		\j3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w406_
	);
	LUT4 #(
		.INIT('h1555)
	) name263 (
		\i3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w407_
	);
	LUT3 #(
		.INIT('h02)
	) name264 (
		_w155_,
		_w407_,
		_w406_,
		_w408_
	);
	LUT4 #(
		.INIT('h0060)
	) name265 (
		\i4_pad ,
		\n1_pad ,
		\o0_pad ,
		\q0_pad ,
		_w409_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		_w163_,
		_w409_,
		_w410_
	);
	LUT4 #(
		.INIT('hacca)
	) name267 (
		\a3_pad ,
		\i3_pad ,
		\k0_pad ,
		\l0_pad ,
		_w411_
	);
	LUT3 #(
		.INIT('he4)
	) name268 (
		\m0_pad ,
		\q3_pad ,
		_w411_,
		_w412_
	);
	LUT3 #(
		.INIT('h04)
	) name269 (
		\g1_pad ,
		\j1_pad ,
		_w398_,
		_w413_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		\c1_pad ,
		\d1_pad ,
		_w414_
	);
	LUT2 #(
		.INIT('h8)
	) name271 (
		_w381_,
		_w414_,
		_w415_
	);
	LUT3 #(
		.INIT('ha8)
	) name272 (
		_w155_,
		_w413_,
		_w415_,
		_w416_
	);
	LUT4 #(
		.INIT('h2000)
	) name273 (
		\c0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w417_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name274 (
		\j2_pad ,
		\k2_pad ,
		_w158_,
		_w163_,
		_w418_
	);
	LUT3 #(
		.INIT('ha8)
	) name275 (
		_w155_,
		_w417_,
		_w418_,
		_w419_
	);
	LUT4 #(
		.INIT('h4000)
	) name276 (
		\k3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w420_
	);
	LUT4 #(
		.INIT('h1555)
	) name277 (
		\j3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w421_
	);
	LUT3 #(
		.INIT('h02)
	) name278 (
		_w155_,
		_w421_,
		_w420_,
		_w422_
	);
	LUT3 #(
		.INIT('h01)
	) name279 (
		\k1_pad ,
		\l1_pad ,
		\u0_pad ,
		_w423_
	);
	LUT2 #(
		.INIT('h8)
	) name280 (
		\m6_pad ,
		\n4_pad ,
		_w424_
	);
	LUT4 #(
		.INIT('h4c00)
	) name281 (
		_w157_,
		_w180_,
		_w423_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w248_,
		_w425_,
		_w426_
	);
	LUT3 #(
		.INIT('hc8)
	) name283 (
		\k1_pad ,
		\l1_pad ,
		\w0_pad ,
		_w427_
	);
	LUT4 #(
		.INIT('h0111)
	) name284 (
		\i1_pad ,
		\j1_pad ,
		\k1_pad ,
		\v0_pad ,
		_w428_
	);
	LUT3 #(
		.INIT('h45)
	) name285 (
		\h1_pad ,
		_w427_,
		_w428_,
		_w429_
	);
	LUT3 #(
		.INIT('ha8)
	) name286 (
		_w178_,
		_w246_,
		_w429_,
		_w430_
	);
	LUT4 #(
		.INIT('h0040)
	) name287 (
		\g1_pad ,
		\j4_pad ,
		\o0_pad ,
		\q0_pad ,
		_w431_
	);
	LUT3 #(
		.INIT('h70)
	) name288 (
		_w426_,
		_w430_,
		_w431_,
		_w432_
	);
	LUT4 #(
		.INIT('h0040)
	) name289 (
		\j4_pad ,
		\n4_pad ,
		\o0_pad ,
		\q0_pad ,
		_w433_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		_w372_,
		_w433_,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		_w178_,
		_w434_,
		_w435_
	);
	LUT2 #(
		.INIT('h4)
	) name292 (
		_w253_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('he)
	) name293 (
		_w432_,
		_w436_,
		_w437_
	);
	LUT4 #(
		.INIT('h0054)
	) name294 (
		\g1_pad ,
		\k1_pad ,
		_w381_,
		_w398_,
		_w438_
	);
	LUT2 #(
		.INIT('h8)
	) name295 (
		\c1_pad ,
		\d1_pad ,
		_w439_
	);
	LUT2 #(
		.INIT('h8)
	) name296 (
		_w381_,
		_w439_,
		_w440_
	);
	LUT3 #(
		.INIT('ha8)
	) name297 (
		_w155_,
		_w438_,
		_w440_,
		_w441_
	);
	LUT4 #(
		.INIT('haaca)
	) name298 (
		a_pad,
		i_pad,
		\k0_pad ,
		\l0_pad ,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w166_,
		_w442_,
		_w443_
	);
	LUT4 #(
		.INIT('h00ca)
	) name300 (
		\k2_pad ,
		\l2_pad ,
		_w163_,
		_w166_,
		_w444_
	);
	LUT3 #(
		.INIT('ha8)
	) name301 (
		_w155_,
		_w443_,
		_w444_,
		_w445_
	);
	LUT4 #(
		.INIT('h4000)
	) name302 (
		\l3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w446_
	);
	LUT4 #(
		.INIT('h1555)
	) name303 (
		\k3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w447_
	);
	LUT3 #(
		.INIT('h02)
	) name304 (
		_w155_,
		_w447_,
		_w446_,
		_w448_
	);
	LUT3 #(
		.INIT('h08)
	) name305 (
		\m1_pad ,
		\o0_pad ,
		\q0_pad ,
		_w449_
	);
	LUT3 #(
		.INIT('h80)
	) name306 (
		_w160_,
		_w162_,
		_w449_,
		_w450_
	);
	LUT4 #(
		.INIT('h4000)
	) name307 (
		\n0_pad ,
		_w156_,
		_w157_,
		_w382_,
		_w451_
	);
	LUT2 #(
		.INIT('h4)
	) name308 (
		\g1_pad ,
		\l1_pad ,
		_w452_
	);
	LUT4 #(
		.INIT('h2220)
	) name309 (
		_w155_,
		_w381_,
		_w451_,
		_w452_,
		_w453_
	);
	LUT4 #(
		.INIT('haaca)
	) name310 (
		b_pad,
		j_pad,
		\k0_pad ,
		\l0_pad ,
		_w454_
	);
	LUT2 #(
		.INIT('h8)
	) name311 (
		_w166_,
		_w454_,
		_w455_
	);
	LUT4 #(
		.INIT('h00ca)
	) name312 (
		\l2_pad ,
		\m2_pad ,
		_w163_,
		_w166_,
		_w456_
	);
	LUT3 #(
		.INIT('ha8)
	) name313 (
		_w155_,
		_w455_,
		_w456_,
		_w457_
	);
	LUT4 #(
		.INIT('h4000)
	) name314 (
		\m3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w458_
	);
	LUT4 #(
		.INIT('h1555)
	) name315 (
		\l3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w459_
	);
	LUT3 #(
		.INIT('h02)
	) name316 (
		_w155_,
		_w459_,
		_w458_,
		_w460_
	);
	LUT4 #(
		.INIT('hbf00)
	) name317 (
		\x3_pad ,
		_w160_,
		_w162_,
		_w449_,
		_w461_
	);
	LUT3 #(
		.INIT('h41)
	) name318 (
		\e3_pad ,
		\k0_pad ,
		\l0_pad ,
		_w462_
	);
	LUT4 #(
		.INIT('hf090)
	) name319 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		\m3_pad ,
		_w463_
	);
	LUT2 #(
		.INIT('h4)
	) name320 (
		_w462_,
		_w463_,
		_w464_
	);
	LUT4 #(
		.INIT('haa80)
	) name321 (
		\m1_pad ,
		_w177_,
		_w357_,
		_w359_,
		_w465_
	);
	LUT3 #(
		.INIT('h45)
	) name322 (
		\m1_pad ,
		\n0_pad ,
		\p0_pad ,
		_w466_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		_w155_,
		_w466_,
		_w467_
	);
	LUT2 #(
		.INIT('h4)
	) name324 (
		_w465_,
		_w467_,
		_w468_
	);
	LUT4 #(
		.INIT('haae2)
	) name325 (
		c_pad,
		\k0_pad ,
		k_pad,
		\l0_pad ,
		_w469_
	);
	LUT2 #(
		.INIT('h8)
	) name326 (
		_w166_,
		_w469_,
		_w470_
	);
	LUT4 #(
		.INIT('h00ca)
	) name327 (
		\m2_pad ,
		\n2_pad ,
		_w163_,
		_w166_,
		_w471_
	);
	LUT3 #(
		.INIT('ha8)
	) name328 (
		_w155_,
		_w470_,
		_w471_,
		_w472_
	);
	LUT4 #(
		.INIT('h2000)
	) name329 (
		\m6_pad ,
		\n3_pad ,
		_w178_,
		_w181_,
		_w473_
	);
	LUT4 #(
		.INIT('h1555)
	) name330 (
		\m3_pad ,
		\m6_pad ,
		_w178_,
		_w181_,
		_w474_
	);
	LUT3 #(
		.INIT('h02)
	) name331 (
		_w155_,
		_w474_,
		_w473_,
		_w475_
	);
	LUT4 #(
		.INIT('ha280)
	) name332 (
		_w155_,
		_w177_,
		_w357_,
		_w359_,
		_w476_
	);
	LUT3 #(
		.INIT('h41)
	) name333 (
		\f3_pad ,
		\k0_pad ,
		\l0_pad ,
		_w477_
	);
	LUT4 #(
		.INIT('hf090)
	) name334 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		\n3_pad ,
		_w478_
	);
	LUT2 #(
		.INIT('h4)
	) name335 (
		_w477_,
		_w478_,
		_w479_
	);
	LUT4 #(
		.INIT('h2aea)
	) name336 (
		\n1_pad ,
		_w160_,
		_w162_,
		_w329_,
		_w480_
	);
	LUT4 #(
		.INIT('h2000)
	) name337 (
		\j0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w481_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name338 (
		\n1_pad ,
		\o1_pad ,
		_w158_,
		_w163_,
		_w482_
	);
	LUT3 #(
		.INIT('ha8)
	) name339 (
		_w155_,
		_w481_,
		_w482_,
		_w483_
	);
	LUT4 #(
		.INIT('haea2)
	) name340 (
		d_pad,
		\k0_pad ,
		\l0_pad ,
		l_pad,
		_w484_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w166_,
		_w484_,
		_w485_
	);
	LUT4 #(
		.INIT('h00ca)
	) name342 (
		\n2_pad ,
		\o2_pad ,
		_w163_,
		_w166_,
		_w486_
	);
	LUT3 #(
		.INIT('ha8)
	) name343 (
		_w155_,
		_w485_,
		_w486_,
		_w487_
	);
	LUT4 #(
		.INIT('h2000)
	) name344 (
		\m6_pad ,
		\o3_pad ,
		_w178_,
		_w181_,
		_w488_
	);
	LUT4 #(
		.INIT('h1333)
	) name345 (
		\m6_pad ,
		\n3_pad ,
		_w178_,
		_w181_,
		_w489_
	);
	LUT3 #(
		.INIT('h02)
	) name346 (
		_w155_,
		_w489_,
		_w488_,
		_w490_
	);
	LUT3 #(
		.INIT('h08)
	) name347 (
		\m6_pad ,
		\o0_pad ,
		\q0_pad ,
		_w491_
	);
	LUT4 #(
		.INIT('hbf00)
	) name348 (
		_w175_,
		_w174_,
		_w176_,
		_w491_,
		_w492_
	);
	LUT3 #(
		.INIT('h41)
	) name349 (
		\g3_pad ,
		\k0_pad ,
		\l0_pad ,
		_w493_
	);
	LUT4 #(
		.INIT('hf090)
	) name350 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		\o3_pad ,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name351 (
		_w493_,
		_w494_,
		_w495_
	);
	LUT3 #(
		.INIT('hf7)
	) name352 (
		\h1_pad ,
		\m1_pad ,
		\m6_pad ,
		_w496_
	);
	LUT4 #(
		.INIT('h2000)
	) name353 (
		\i0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w497_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name354 (
		\o1_pad ,
		\p1_pad ,
		_w158_,
		_w163_,
		_w498_
	);
	LUT3 #(
		.INIT('ha8)
	) name355 (
		_w155_,
		_w497_,
		_w498_,
		_w499_
	);
	LUT4 #(
		.INIT('haea2)
	) name356 (
		e_pad,
		\k0_pad ,
		\l0_pad ,
		m_pad,
		_w500_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		_w166_,
		_w500_,
		_w501_
	);
	LUT4 #(
		.INIT('h00ca)
	) name358 (
		\o2_pad ,
		\p2_pad ,
		_w163_,
		_w166_,
		_w502_
	);
	LUT3 #(
		.INIT('ha8)
	) name359 (
		_w155_,
		_w501_,
		_w502_,
		_w503_
	);
	LUT4 #(
		.INIT('h2000)
	) name360 (
		\m6_pad ,
		\p3_pad ,
		_w178_,
		_w181_,
		_w504_
	);
	LUT4 #(
		.INIT('h1333)
	) name361 (
		\m6_pad ,
		\o3_pad ,
		_w178_,
		_w181_,
		_w505_
	);
	LUT3 #(
		.INIT('h02)
	) name362 (
		_w155_,
		_w505_,
		_w504_,
		_w506_
	);
	LUT3 #(
		.INIT('h41)
	) name363 (
		\h3_pad ,
		\k0_pad ,
		\l0_pad ,
		_w507_
	);
	LUT4 #(
		.INIT('hf090)
	) name364 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		\p3_pad ,
		_w508_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		_w507_,
		_w508_,
		_w509_
	);
	LUT3 #(
		.INIT('hf7)
	) name366 (
		\i1_pad ,
		\m1_pad ,
		\m6_pad ,
		_w510_
	);
	LUT4 #(
		.INIT('h2000)
	) name367 (
		\h0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w511_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name368 (
		\p1_pad ,
		\q1_pad ,
		_w158_,
		_w163_,
		_w512_
	);
	LUT3 #(
		.INIT('ha8)
	) name369 (
		_w155_,
		_w511_,
		_w512_,
		_w513_
	);
	LUT4 #(
		.INIT('haea2)
	) name370 (
		f_pad,
		\k0_pad ,
		\l0_pad ,
		n_pad,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name371 (
		_w166_,
		_w514_,
		_w515_
	);
	LUT4 #(
		.INIT('h00ca)
	) name372 (
		\p2_pad ,
		\q2_pad ,
		_w163_,
		_w166_,
		_w516_
	);
	LUT3 #(
		.INIT('ha8)
	) name373 (
		_w155_,
		_w515_,
		_w516_,
		_w517_
	);
	LUT4 #(
		.INIT('h2000)
	) name374 (
		\m6_pad ,
		\q3_pad ,
		_w178_,
		_w181_,
		_w518_
	);
	LUT4 #(
		.INIT('h1333)
	) name375 (
		\m6_pad ,
		\p3_pad ,
		_w178_,
		_w181_,
		_w519_
	);
	LUT3 #(
		.INIT('h02)
	) name376 (
		_w155_,
		_w519_,
		_w518_,
		_w520_
	);
	LUT3 #(
		.INIT('h41)
	) name377 (
		\i3_pad ,
		\k0_pad ,
		\l0_pad ,
		_w521_
	);
	LUT4 #(
		.INIT('hf090)
	) name378 (
		\k0_pad ,
		\l0_pad ,
		\m0_pad ,
		\q3_pad ,
		_w522_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		_w521_,
		_w522_,
		_w523_
	);
	LUT3 #(
		.INIT('hf7)
	) name380 (
		\j1_pad ,
		\m1_pad ,
		\m6_pad ,
		_w524_
	);
	LUT4 #(
		.INIT('h2000)
	) name381 (
		\g0_pad ,
		\n0_pad ,
		_w156_,
		_w157_,
		_w525_
	);
	LUT4 #(
		.INIT('h0c0a)
	) name382 (
		\q1_pad ,
		\r1_pad ,
		_w158_,
		_w163_,
		_w526_
	);
	LUT3 #(
		.INIT('ha8)
	) name383 (
		_w155_,
		_w525_,
		_w526_,
		_w527_
	);
	LUT4 #(
		.INIT('haea2)
	) name384 (
		g_pad,
		\k0_pad ,
		\l0_pad ,
		o_pad,
		_w528_
	);
	LUT2 #(
		.INIT('h8)
	) name385 (
		_w166_,
		_w528_,
		_w529_
	);
	LUT4 #(
		.INIT('h00ca)
	) name386 (
		\q2_pad ,
		\r2_pad ,
		_w163_,
		_w166_,
		_w530_
	);
	LUT3 #(
		.INIT('ha8)
	) name387 (
		_w155_,
		_w529_,
		_w530_,
		_w531_
	);
	LUT4 #(
		.INIT('h2000)
	) name388 (
		\m6_pad ,
		\r3_pad ,
		_w178_,
		_w181_,
		_w532_
	);
	LUT4 #(
		.INIT('h1333)
	) name389 (
		\m6_pad ,
		\q3_pad ,
		_w178_,
		_w181_,
		_w533_
	);
	LUT3 #(
		.INIT('h02)
	) name390 (
		_w155_,
		_w533_,
		_w532_,
		_w534_
	);
	assign \a5_pad  = _w153_ ;
	assign \a6_pad  = _w154_ ;
	assign \a7_pad  = _w165_ ;
	assign \a8_pad  = _w170_ ;
	assign \a9_pad  = _w184_ ;
	assign \b5_pad  = _w187_ ;
	assign \b6_pad  = _w188_ ;
	assign \b7_pad  = _w191_ ;
	assign \b8_pad  = _w195_ ;
	assign \b9_pad  = _w198_ ;
	assign \c5_pad  = _w201_ ;
	assign \c6_pad  = _w202_ ;
	assign \c7_pad  = _w205_ ;
	assign \c8_pad  = _w208_ ;
	assign \c9_pad  = _w211_ ;
	assign \d5_pad  = _w212_ ;
	assign \d6_pad  = _w213_ ;
	assign \d7_pad  = _w216_ ;
	assign \d8_pad  = _w219_ ;
	assign \d9_pad  = _w222_ ;
	assign \e5_pad  = _w223_ ;
	assign \e6_pad  = _w224_ ;
	assign \e7_pad  = _w228_ ;
	assign \e8_pad  = _w231_ ;
	assign \e9_pad  = _w234_ ;
	assign \f5_pad  = _w235_ ;
	assign \f6_pad  = _w236_ ;
	assign \f7_pad  = _w240_ ;
	assign \f8_pad  = _w243_ ;
	assign \f9_pad  = _w254_ ;
	assign \g5_pad  = _w255_ ;
	assign \g6_pad  = _w256_ ;
	assign \g7_pad  = _w259_ ;
	assign \g8_pad  = _w262_ ;
	assign \g9_pad  = _w266_ ;
	assign \h5_pad  = _w267_ ;
	assign \h6_pad  = _w47_ ;
	assign \h7_pad  = _w270_ ;
	assign \h8_pad  = _w273_ ;
	assign \h9_pad  = _w275_ ;
	assign \i5_pad  = _w276_ ;
	assign \i6_pad  = _w54_ ;
	assign \i7_pad  = _w279_ ;
	assign \i8_pad  = _w282_ ;
	assign \i9_pad  = _w285_ ;
	assign \j5_pad  = _w286_ ;
	assign \j6_pad  = _w61_ ;
	assign \j7_pad  = _w289_ ;
	assign \j8_pad  = _w292_ ;
	assign \j9_pad  = _w297_ ;
	assign \k5_pad  = _w298_ ;
	assign \k6_pad  = _w68_ ;
	assign \k7_pad  = _w301_ ;
	assign \k8_pad  = _w304_ ;
	assign \k9_pad  = _w308_ ;
	assign \l5_pad  = _w309_ ;
	assign \l6_pad  = _w74_ ;
	assign \l7_pad  = _w312_ ;
	assign \l8_pad  = _w315_ ;
	assign \l9_pad  = _w317_ ;
	assign \m7_pad  = _w320_ ;
	assign \m8_pad  = _w323_ ;
	assign \m9_pad  = _w327_ ;
	assign \n5_pad  = _w328_ ;
	assign \n6_pad  = _w330_ ;
	assign \n7_pad  = _w333_ ;
	assign \n8_pad  = _w336_ ;
	assign \n9_pad  = _w342_ ;
	assign \o4_pad  = _w40_ ;
	assign \o5_pad  = _w343_ ;
	assign \o6_pad  = _w344_ ;
	assign \o7_pad  = _w347_ ;
	assign \o8_pad  = _w350_ ;
	assign \o9_pad  = _w353_ ;
	assign \p4_pad  = _w355_ ;
	assign \p5_pad  = _w356_ ;
	assign \p6_pad  = _w360_ ;
	assign \p7_pad  = _w363_ ;
	assign \p8_pad  = _w366_ ;
	assign \p9_pad  = _w376_ ;
	assign \q4_pad  = _w378_ ;
	assign \q5_pad  = _w379_ ;
	assign \q6_pad  = _w384_ ;
	assign \q7_pad  = _w387_ ;
	assign \q8_pad  = _w390_ ;
	assign \q9_pad  = _w393_ ;
	assign \r4_pad  = _w395_ ;
	assign \r5_pad  = _w396_ ;
	assign \r6_pad  = _w402_ ;
	assign \r7_pad  = _w405_ ;
	assign \r8_pad  = _w408_ ;
	assign \r9_pad  = _w410_ ;
	assign \s4_pad  = _w412_ ;
	assign \s6_pad  = _w416_ ;
	assign \s7_pad  = _w419_ ;
	assign \s8_pad  = _w422_ ;
	assign \s9_pad  = _w437_ ;
	assign \t6_pad  = _w441_ ;
	assign \t7_pad  = _w445_ ;
	assign \t8_pad  = _w448_ ;
	assign \t9_pad  = _w450_ ;
	assign \u6_pad  = _w453_ ;
	assign \u7_pad  = _w457_ ;
	assign \u8_pad  = _w460_ ;
	assign \u9_pad  = _w461_ ;
	assign \v4_pad  = _w464_ ;
	assign \v6_pad  = _w468_ ;
	assign \v7_pad  = _w472_ ;
	assign \v8_pad  = _w475_ ;
	assign \v9_pad  = _w476_ ;
	assign \w4_pad  = _w479_ ;
	assign \w5_pad  = _w480_ ;
	assign \w6_pad  = _w483_ ;
	assign \w7_pad  = _w487_ ;
	assign \w8_pad  = _w490_ ;
	assign \w9_pad  = _w492_ ;
	assign \x4_pad  = _w495_ ;
	assign \x5_pad  = _w496_ ;
	assign \x6_pad  = _w499_ ;
	assign \x7_pad  = _w503_ ;
	assign \x8_pad  = _w506_ ;
	assign \y4_pad  = _w509_ ;
	assign \y5_pad  = _w510_ ;
	assign \y6_pad  = _w513_ ;
	assign \y7_pad  = _w517_ ;
	assign \y8_pad  = _w520_ ;
	assign \z4_pad  = _w523_ ;
	assign \z5_pad  = _w524_ ;
	assign \z6_pad  = _w527_ ;
	assign \z7_pad  = _w531_ ;
	assign \z8_pad  = _w534_ ;
endmodule;