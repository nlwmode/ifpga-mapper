module top (\a0_pad , a_pad, b_pad, c_pad, d_pad, e_pad, f_pad, g_pad, h_pad, i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \b0_pad , \c0_pad , \d0_pad , \e0_pad , \f0_pad , \g0_pad , \h0_pad , \i0_pad , \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad );
	input \a0_pad  ;
	input a_pad ;
	input b_pad ;
	input c_pad ;
	input d_pad ;
	input e_pad ;
	input f_pad ;
	input g_pad ;
	input h_pad ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \b0_pad  ;
	output \c0_pad  ;
	output \d0_pad  ;
	output \e0_pad  ;
	output \f0_pad  ;
	output \g0_pad  ;
	output \h0_pad  ;
	output \i0_pad  ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w41_ ;
	wire _w40_ ;
	wire _w39_ ;
	wire _w38_ ;
	wire _w37_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	LUT4 #(
		.INIT('h8000)
	) name0 (
		t_pad,
		u_pad,
		v_pad,
		w_pad,
		_w29_
	);
	LUT3 #(
		.INIT('h80)
	) name1 (
		x_pad,
		y_pad,
		z_pad,
		_w30_
	);
	LUT3 #(
		.INIT('h04)
	) name2 (
		i_pad,
		j_pad,
		k_pad,
		_w31_
	);
	LUT4 #(
		.INIT('h0020)
	) name3 (
		\a0_pad ,
		i_pad,
		j_pad,
		k_pad,
		_w32_
	);
	LUT3 #(
		.INIT('h80)
	) name4 (
		_w29_,
		_w30_,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		a_pad,
		i_pad,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name6 (
		b_pad,
		i_pad,
		_w35_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		c_pad,
		i_pad,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		d_pad,
		i_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		e_pad,
		i_pad,
		_w38_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		f_pad,
		i_pad,
		_w39_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		g_pad,
		i_pad,
		_w40_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		h_pad,
		i_pad,
		_w41_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\a0_pad ,
		l_pad,
		_w42_
	);
	LUT4 #(
		.INIT('h8000)
	) name14 (
		_w29_,
		_w30_,
		_w31_,
		_w42_,
		_w43_
	);
	LUT4 #(
		.INIT('h0004)
	) name15 (
		i_pad,
		j_pad,
		k_pad,
		t_pad,
		_w44_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w34_,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('hb)
	) name17 (
		_w43_,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h6)
	) name18 (
		t_pad,
		u_pad,
		_w47_
	);
	LUT3 #(
		.INIT('h82)
	) name19 (
		m_pad,
		t_pad,
		u_pad,
		_w48_
	);
	LUT4 #(
		.INIT('h8000)
	) name20 (
		_w29_,
		_w30_,
		_w32_,
		_w48_,
		_w49_
	);
	LUT3 #(
		.INIT('h13)
	) name21 (
		_w31_,
		_w35_,
		_w47_,
		_w50_
	);
	LUT2 #(
		.INIT('hb)
	) name22 (
		_w49_,
		_w50_,
		_w51_
	);
	LUT4 #(
		.INIT('h7fd5)
	) name23 (
		n_pad,
		t_pad,
		u_pad,
		v_pad,
		_w52_
	);
	LUT4 #(
		.INIT('h0080)
	) name24 (
		_w29_,
		_w30_,
		_w32_,
		_w52_,
		_w53_
	);
	LUT3 #(
		.INIT('h80)
	) name25 (
		t_pad,
		u_pad,
		v_pad,
		_w54_
	);
	LUT3 #(
		.INIT('h78)
	) name26 (
		t_pad,
		u_pad,
		v_pad,
		_w55_
	);
	LUT3 #(
		.INIT('h13)
	) name27 (
		_w31_,
		_w36_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('hb)
	) name28 (
		_w53_,
		_w56_,
		_w57_
	);
	LUT3 #(
		.INIT('h7d)
	) name29 (
		o_pad,
		w_pad,
		_w54_,
		_w58_
	);
	LUT4 #(
		.INIT('h007f)
	) name30 (
		t_pad,
		u_pad,
		v_pad,
		w_pad,
		_w59_
	);
	LUT4 #(
		.INIT('h0f0b)
	) name31 (
		_w29_,
		_w31_,
		_w37_,
		_w59_,
		_w60_
	);
	LUT3 #(
		.INIT('h2f)
	) name32 (
		_w33_,
		_w58_,
		_w60_,
		_w61_
	);
	LUT3 #(
		.INIT('h7d)
	) name33 (
		p_pad,
		x_pad,
		_w29_,
		_w62_
	);
	LUT4 #(
		.INIT('h0400)
	) name34 (
		i_pad,
		j_pad,
		k_pad,
		x_pad,
		_w63_
	);
	LUT4 #(
		.INIT('h0004)
	) name35 (
		i_pad,
		j_pad,
		k_pad,
		x_pad,
		_w64_
	);
	LUT4 #(
		.INIT('h0123)
	) name36 (
		_w29_,
		_w38_,
		_w63_,
		_w64_,
		_w65_
	);
	LUT3 #(
		.INIT('h2f)
	) name37 (
		_w33_,
		_w62_,
		_w65_,
		_w66_
	);
	LUT4 #(
		.INIT('h7df5)
	) name38 (
		q_pad,
		x_pad,
		y_pad,
		_w29_,
		_w67_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		x_pad,
		y_pad,
		_w68_
	);
	LUT4 #(
		.INIT('h6c00)
	) name40 (
		x_pad,
		y_pad,
		_w29_,
		_w31_,
		_w69_
	);
	LUT4 #(
		.INIT('hffce)
	) name41 (
		_w33_,
		_w39_,
		_w67_,
		_w69_,
		_w70_
	);
	LUT3 #(
		.INIT('h15)
	) name42 (
		z_pad,
		_w29_,
		_w68_,
		_w71_
	);
	LUT3 #(
		.INIT('h70)
	) name43 (
		_w29_,
		_w30_,
		_w31_,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name44 (
		\a0_pad ,
		r_pad,
		_w73_
	);
	LUT4 #(
		.INIT('h8000)
	) name45 (
		_w29_,
		_w30_,
		_w31_,
		_w73_,
		_w74_
	);
	LUT4 #(
		.INIT('hffba)
	) name46 (
		_w40_,
		_w71_,
		_w72_,
		_w74_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		\a0_pad ,
		s_pad,
		_w76_
	);
	LUT3 #(
		.INIT('h80)
	) name48 (
		_w29_,
		_w30_,
		_w76_,
		_w77_
	);
	LUT4 #(
		.INIT('hea00)
	) name49 (
		\a0_pad ,
		_w29_,
		_w30_,
		_w31_,
		_w78_
	);
	LUT3 #(
		.INIT('hba)
	) name50 (
		_w41_,
		_w77_,
		_w78_,
		_w79_
	);
	assign \b0_pad  = _w33_ ;
	assign \c0_pad  = _w34_ ;
	assign \d0_pad  = _w35_ ;
	assign \e0_pad  = _w36_ ;
	assign \f0_pad  = _w37_ ;
	assign \g0_pad  = _w38_ ;
	assign \h0_pad  = _w39_ ;
	assign \i0_pad  = _w40_ ;
	assign \j0_pad  = _w41_ ;
	assign \k0_pad  = _w46_ ;
	assign \l0_pad  = _w51_ ;
	assign \m0_pad  = _w57_ ;
	assign \n0_pad  = _w61_ ;
	assign \o0_pad  = _w66_ ;
	assign \p0_pad  = _w70_ ;
	assign \q0_pad  = _w75_ ;
	assign \r0_pad  = _w79_ ;
endmodule;