module top (\ac97_reset_pad_o__pad , \dma_ack_i[0]_pad , \dma_ack_i[1]_pad , \dma_ack_i[2]_pad , \dma_ack_i[3]_pad , \dma_ack_i[4]_pad , \dma_ack_i[5]_pad , \dma_ack_i[6]_pad , \dma_ack_i[7]_pad , \dma_ack_i[8]_pad , \dma_req_o[0]_pad , \dma_req_o[1]_pad , \dma_req_o[2]_pad , \dma_req_o[3]_pad , \dma_req_o[4]_pad , \dma_req_o[5]_pad , \dma_req_o[6]_pad , \dma_req_o[7]_pad , \dma_req_o[8]_pad , \in_valid_s_reg[0]/NET0131 , \in_valid_s_reg[1]/NET0131 , \in_valid_s_reg[2]/NET0131 , suspended_o_pad, \u0_slt0_r_reg[0]/P0001 , \u0_slt0_r_reg[10]/P0001 , \u0_slt0_r_reg[11]/P0001 , \u0_slt0_r_reg[12]/P0001 , \u0_slt0_r_reg[13]/P0001 , \u0_slt0_r_reg[14]/P0001 , \u0_slt0_r_reg[1]/P0001 , \u0_slt0_r_reg[2]/P0001 , \u0_slt0_r_reg[3]/P0001 , \u0_slt0_r_reg[4]/P0001 , \u0_slt0_r_reg[5]/P0001 , \u0_slt0_r_reg[6]/P0001 , \u0_slt0_r_reg[7]/P0001 , \u0_slt0_r_reg[8]/P0001 , \u0_slt0_r_reg[9]/P0001 , \u0_slt1_r_reg[0]/P0001 , \u0_slt1_r_reg[10]/P0001 , \u0_slt1_r_reg[11]/P0001 , \u0_slt1_r_reg[12]/P0001 , \u0_slt1_r_reg[13]/P0001 , \u0_slt1_r_reg[14]/P0001 , \u0_slt1_r_reg[15]/P0001 , \u0_slt1_r_reg[16]/P0001 , \u0_slt1_r_reg[17]/P0001 , \u0_slt1_r_reg[18]/P0001 , \u0_slt1_r_reg[19]/P0001 , \u0_slt1_r_reg[1]/P0001 , \u0_slt1_r_reg[2]/P0001 , \u0_slt1_r_reg[3]/P0001 , \u0_slt1_r_reg[4]/P0001 , \u0_slt1_r_reg[5]/P0001 , \u0_slt1_r_reg[6]/P0001 , \u0_slt1_r_reg[7]/P0001 , \u0_slt1_r_reg[8]/P0001 , \u0_slt1_r_reg[9]/P0001 , \u0_slt2_r_reg[0]/P0001 , \u0_slt2_r_reg[10]/P0001 , \u0_slt2_r_reg[11]/P0001 , \u0_slt2_r_reg[12]/P0001 , \u0_slt2_r_reg[13]/P0001 , \u0_slt2_r_reg[14]/P0001 , \u0_slt2_r_reg[15]/P0001 , \u0_slt2_r_reg[16]/P0001 , \u0_slt2_r_reg[17]/P0001 , \u0_slt2_r_reg[18]/P0001 , \u0_slt2_r_reg[19]/P0001 , \u0_slt2_r_reg[1]/P0001 , \u0_slt2_r_reg[2]/P0001 , \u0_slt2_r_reg[3]/P0001 , \u0_slt2_r_reg[4]/P0001 , \u0_slt2_r_reg[5]/P0001 , \u0_slt2_r_reg[6]/P0001 , \u0_slt2_r_reg[7]/P0001 , \u0_slt2_r_reg[8]/P0001 , \u0_slt2_r_reg[9]/P0001 , \u0_slt3_r_reg[0]/P0001 , \u0_slt3_r_reg[10]/P0001 , \u0_slt3_r_reg[11]/P0001 , \u0_slt3_r_reg[12]/P0001 , \u0_slt3_r_reg[13]/P0001 , \u0_slt3_r_reg[14]/P0001 , \u0_slt3_r_reg[15]/P0001 , \u0_slt3_r_reg[16]/P0001 , \u0_slt3_r_reg[17]/P0001 , \u0_slt3_r_reg[18]/P0001 , \u0_slt3_r_reg[19]/P0001 , \u0_slt3_r_reg[1]/P0001 , \u0_slt3_r_reg[2]/P0001 , \u0_slt3_r_reg[3]/P0001 , \u0_slt3_r_reg[4]/P0001 , \u0_slt3_r_reg[5]/P0001 , \u0_slt3_r_reg[6]/P0001 , \u0_slt3_r_reg[7]/P0001 , \u0_slt3_r_reg[8]/P0001 , \u0_slt3_r_reg[9]/P0001 , \u0_slt4_r_reg[0]/P0001 , \u0_slt4_r_reg[10]/P0001 , \u0_slt4_r_reg[11]/P0001 , \u0_slt4_r_reg[12]/P0001 , \u0_slt4_r_reg[13]/P0001 , \u0_slt4_r_reg[14]/P0001 , \u0_slt4_r_reg[15]/P0001 , \u0_slt4_r_reg[16]/P0001 , \u0_slt4_r_reg[17]/P0001 , \u0_slt4_r_reg[18]/P0001 , \u0_slt4_r_reg[19]/P0001 , \u0_slt4_r_reg[1]/P0001 , \u0_slt4_r_reg[2]/P0001 , \u0_slt4_r_reg[3]/P0001 , \u0_slt4_r_reg[4]/P0001 , \u0_slt4_r_reg[5]/P0001 , \u0_slt4_r_reg[6]/P0001 , \u0_slt4_r_reg[7]/P0001 , \u0_slt4_r_reg[8]/P0001 , \u0_slt4_r_reg[9]/P0001 , \u0_slt5_r_reg[0]/P0001 , \u0_slt5_r_reg[10]/P0001 , \u0_slt5_r_reg[11]/P0001 , \u0_slt5_r_reg[12]/P0001 , \u0_slt5_r_reg[13]/P0001 , \u0_slt5_r_reg[14]/P0001 , \u0_slt5_r_reg[15]/P0001 , \u0_slt5_r_reg[16]/P0001 , \u0_slt5_r_reg[17]/P0001 , \u0_slt5_r_reg[18]/P0001 , \u0_slt5_r_reg[19]/P0001 , \u0_slt5_r_reg[1]/P0001 , \u0_slt5_r_reg[2]/P0001 , \u0_slt5_r_reg[3]/P0001 , \u0_slt5_r_reg[4]/P0001 , \u0_slt5_r_reg[5]/P0001 , \u0_slt5_r_reg[6]/P0001 , \u0_slt5_r_reg[7]/P0001 , \u0_slt5_r_reg[8]/P0001 , \u0_slt5_r_reg[9]/P0001 , \u0_slt6_r_reg[0]/P0001 , \u0_slt6_r_reg[10]/P0001 , \u0_slt6_r_reg[11]/P0001 , \u0_slt6_r_reg[12]/P0001 , \u0_slt6_r_reg[13]/P0001 , \u0_slt6_r_reg[14]/P0001 , \u0_slt6_r_reg[15]/P0001 , \u0_slt6_r_reg[16]/P0001 , \u0_slt6_r_reg[17]/P0001 , \u0_slt6_r_reg[18]/P0001 , \u0_slt6_r_reg[19]/P0001 , \u0_slt6_r_reg[1]/P0001 , \u0_slt6_r_reg[2]/P0001 , \u0_slt6_r_reg[3]/P0001 , \u0_slt6_r_reg[4]/P0001 , \u0_slt6_r_reg[5]/P0001 , \u0_slt6_r_reg[6]/P0001 , \u0_slt6_r_reg[7]/P0001 , \u0_slt6_r_reg[8]/P0001 , \u0_slt6_r_reg[9]/P0001 , \u0_slt7_r_reg[0]/P0001 , \u0_slt7_r_reg[10]/P0001 , \u0_slt7_r_reg[11]/P0001 , \u0_slt7_r_reg[12]/P0001 , \u0_slt7_r_reg[13]/P0001 , \u0_slt7_r_reg[14]/P0001 , \u0_slt7_r_reg[15]/P0001 , \u0_slt7_r_reg[16]/P0001 , \u0_slt7_r_reg[17]/P0001 , \u0_slt7_r_reg[18]/P0001 , \u0_slt7_r_reg[19]/P0001 , \u0_slt7_r_reg[1]/P0001 , \u0_slt7_r_reg[2]/P0001 , \u0_slt7_r_reg[3]/P0001 , \u0_slt7_r_reg[4]/P0001 , \u0_slt7_r_reg[5]/P0001 , \u0_slt7_r_reg[6]/P0001 , \u0_slt7_r_reg[7]/P0001 , \u0_slt7_r_reg[8]/P0001 , \u0_slt7_r_reg[9]/P0001 , \u0_slt8_r_reg[0]/P0001 , \u0_slt8_r_reg[10]/P0001 , \u0_slt8_r_reg[11]/P0001 , \u0_slt8_r_reg[12]/P0001 , \u0_slt8_r_reg[13]/P0001 , \u0_slt8_r_reg[14]/P0001 , \u0_slt8_r_reg[15]/P0001 , \u0_slt8_r_reg[16]/P0001 , \u0_slt8_r_reg[17]/P0001 , \u0_slt8_r_reg[18]/P0001 , \u0_slt8_r_reg[19]/P0001 , \u0_slt8_r_reg[1]/P0001 , \u0_slt8_r_reg[2]/P0001 , \u0_slt8_r_reg[3]/P0001 , \u0_slt8_r_reg[4]/P0001 , \u0_slt8_r_reg[5]/P0001 , \u0_slt8_r_reg[6]/P0001 , \u0_slt8_r_reg[7]/P0001 , \u0_slt8_r_reg[8]/P0001 , \u0_slt8_r_reg[9]/P0001 , \u0_slt9_r_reg[0]/P0001 , \u0_slt9_r_reg[10]/P0001 , \u0_slt9_r_reg[11]/P0001 , \u0_slt9_r_reg[12]/P0001 , \u0_slt9_r_reg[13]/P0001 , \u0_slt9_r_reg[14]/P0001 , \u0_slt9_r_reg[15]/P0001 , \u0_slt9_r_reg[16]/P0001 , \u0_slt9_r_reg[17]/P0001 , \u0_slt9_r_reg[18]/P0001 , \u0_slt9_r_reg[19]/P0001 , \u0_slt9_r_reg[1]/P0001 , \u0_slt9_r_reg[2]/P0001 , \u0_slt9_r_reg[3]/P0001 , \u0_slt9_r_reg[4]/P0001 , \u0_slt9_r_reg[5]/P0001 , \u0_slt9_r_reg[6]/P0001 , \u0_slt9_r_reg[7]/P0001 , \u0_slt9_r_reg[8]/P0001 , \u0_slt9_r_reg[9]/P0001 , \u10_din_tmp1_reg[0]/P0001 , \u10_din_tmp1_reg[10]/P0001 , \u10_din_tmp1_reg[11]/P0001 , \u10_din_tmp1_reg[12]/P0001 , \u10_din_tmp1_reg[13]/P0001 , \u10_din_tmp1_reg[14]/P0001 , \u10_din_tmp1_reg[15]/P0001 , \u10_din_tmp1_reg[1]/P0001 , \u10_din_tmp1_reg[2]/P0001 , \u10_din_tmp1_reg[3]/P0001 , \u10_din_tmp1_reg[4]/P0001 , \u10_din_tmp1_reg[5]/P0001 , \u10_din_tmp1_reg[6]/P0001 , \u10_din_tmp1_reg[7]/P0001 , \u10_din_tmp1_reg[8]/P0001 , \u10_din_tmp1_reg[9]/P0001 , \u10_dout_reg[0]/P0001 , \u10_dout_reg[10]/P0001 , \u10_dout_reg[11]/P0001 , \u10_dout_reg[12]/P0001 , \u10_dout_reg[13]/P0001 , \u10_dout_reg[14]/P0001 , \u10_dout_reg[15]/P0001 , \u10_dout_reg[16]/P0001 , \u10_dout_reg[17]/P0001 , \u10_dout_reg[18]/P0001 , \u10_dout_reg[19]/P0001 , \u10_dout_reg[1]/P0001 , \u10_dout_reg[20]/P0001 , \u10_dout_reg[21]/P0001 , \u10_dout_reg[22]/P0001 , \u10_dout_reg[23]/P0001 , \u10_dout_reg[24]/P0001 , \u10_dout_reg[25]/P0001 , \u10_dout_reg[26]/P0001 , \u10_dout_reg[27]/P0001 , \u10_dout_reg[28]/P0001 , \u10_dout_reg[29]/P0001 , \u10_dout_reg[2]/P0001 , \u10_dout_reg[30]/P0001 , \u10_dout_reg[31]/P0001 , \u10_dout_reg[3]/P0001 , \u10_dout_reg[4]/P0001 , \u10_dout_reg[5]/P0001 , \u10_dout_reg[6]/P0001 , \u10_dout_reg[7]/P0001 , \u10_dout_reg[8]/P0001 , \u10_dout_reg[9]/P0001 , \u10_empty_reg/P0001 , \u10_full_reg/NET0131 , \u10_mem_reg[0][0]/P0001 , \u10_mem_reg[0][10]/P0001 , \u10_mem_reg[0][11]/P0001 , \u10_mem_reg[0][12]/P0001 , \u10_mem_reg[0][13]/P0001 , \u10_mem_reg[0][14]/P0001 , \u10_mem_reg[0][15]/P0001 , \u10_mem_reg[0][16]/P0001 , \u10_mem_reg[0][17]/P0001 , \u10_mem_reg[0][18]/P0001 , \u10_mem_reg[0][19]/P0001 , \u10_mem_reg[0][1]/P0001 , \u10_mem_reg[0][20]/P0001 , \u10_mem_reg[0][21]/P0001 , \u10_mem_reg[0][22]/P0001 , \u10_mem_reg[0][23]/P0001 , \u10_mem_reg[0][24]/P0001 , \u10_mem_reg[0][25]/P0001 , \u10_mem_reg[0][26]/P0001 , \u10_mem_reg[0][27]/P0001 , \u10_mem_reg[0][28]/P0001 , \u10_mem_reg[0][29]/P0001 , \u10_mem_reg[0][2]/P0001 , \u10_mem_reg[0][30]/P0001 , \u10_mem_reg[0][31]/P0001 , \u10_mem_reg[0][3]/P0001 , \u10_mem_reg[0][4]/P0001 , \u10_mem_reg[0][5]/P0001 , \u10_mem_reg[0][6]/P0001 , \u10_mem_reg[0][7]/P0001 , \u10_mem_reg[0][8]/P0001 , \u10_mem_reg[0][9]/P0001 , \u10_mem_reg[1][0]/P0001 , \u10_mem_reg[1][10]/P0001 , \u10_mem_reg[1][11]/P0001 , \u10_mem_reg[1][12]/P0001 , \u10_mem_reg[1][13]/P0001 , \u10_mem_reg[1][14]/P0001 , \u10_mem_reg[1][15]/P0001 , \u10_mem_reg[1][16]/P0001 , \u10_mem_reg[1][17]/P0001 , \u10_mem_reg[1][18]/P0001 , \u10_mem_reg[1][19]/P0001 , \u10_mem_reg[1][1]/P0001 , \u10_mem_reg[1][20]/P0001 , \u10_mem_reg[1][21]/P0001 , \u10_mem_reg[1][22]/P0001 , \u10_mem_reg[1][23]/P0001 , \u10_mem_reg[1][24]/P0001 , \u10_mem_reg[1][25]/P0001 , \u10_mem_reg[1][26]/P0001 , \u10_mem_reg[1][27]/P0001 , \u10_mem_reg[1][28]/P0001 , \u10_mem_reg[1][29]/P0001 , \u10_mem_reg[1][2]/P0001 , \u10_mem_reg[1][30]/P0001 , \u10_mem_reg[1][31]/P0001 , \u10_mem_reg[1][3]/P0001 , \u10_mem_reg[1][4]/P0001 , \u10_mem_reg[1][5]/P0001 , \u10_mem_reg[1][6]/P0001 , \u10_mem_reg[1][7]/P0001 , \u10_mem_reg[1][8]/P0001 , \u10_mem_reg[1][9]/P0001 , \u10_mem_reg[2][0]/P0001 , \u10_mem_reg[2][10]/P0001 , \u10_mem_reg[2][11]/P0001 , \u10_mem_reg[2][12]/P0001 , \u10_mem_reg[2][13]/P0001 , \u10_mem_reg[2][14]/P0001 , \u10_mem_reg[2][15]/P0001 , \u10_mem_reg[2][16]/P0001 , \u10_mem_reg[2][17]/P0001 , \u10_mem_reg[2][18]/P0001 , \u10_mem_reg[2][19]/P0001 , \u10_mem_reg[2][1]/P0001 , \u10_mem_reg[2][20]/P0001 , \u10_mem_reg[2][21]/P0001 , \u10_mem_reg[2][22]/P0001 , \u10_mem_reg[2][23]/P0001 , \u10_mem_reg[2][24]/P0001 , \u10_mem_reg[2][25]/P0001 , \u10_mem_reg[2][26]/P0001 , \u10_mem_reg[2][27]/P0001 , \u10_mem_reg[2][28]/P0001 , \u10_mem_reg[2][29]/P0001 , \u10_mem_reg[2][2]/P0001 , \u10_mem_reg[2][30]/P0001 , \u10_mem_reg[2][31]/P0001 , \u10_mem_reg[2][3]/P0001 , \u10_mem_reg[2][4]/P0001 , \u10_mem_reg[2][5]/P0001 , \u10_mem_reg[2][6]/P0001 , \u10_mem_reg[2][7]/P0001 , \u10_mem_reg[2][8]/P0001 , \u10_mem_reg[2][9]/P0001 , \u10_mem_reg[3][0]/P0001 , \u10_mem_reg[3][10]/P0001 , \u10_mem_reg[3][11]/P0001 , \u10_mem_reg[3][12]/P0001 , \u10_mem_reg[3][13]/P0001 , \u10_mem_reg[3][14]/P0001 , \u10_mem_reg[3][15]/P0001 , \u10_mem_reg[3][16]/P0001 , \u10_mem_reg[3][17]/P0001 , \u10_mem_reg[3][18]/P0001 , \u10_mem_reg[3][19]/P0001 , \u10_mem_reg[3][1]/P0001 , \u10_mem_reg[3][20]/P0001 , \u10_mem_reg[3][21]/P0001 , \u10_mem_reg[3][22]/P0001 , \u10_mem_reg[3][23]/P0001 , \u10_mem_reg[3][24]/P0001 , \u10_mem_reg[3][25]/P0001 , \u10_mem_reg[3][26]/P0001 , \u10_mem_reg[3][27]/P0001 , \u10_mem_reg[3][28]/P0001 , \u10_mem_reg[3][29]/P0001 , \u10_mem_reg[3][2]/P0001 , \u10_mem_reg[3][30]/P0001 , \u10_mem_reg[3][31]/P0001 , \u10_mem_reg[3][3]/P0001 , \u10_mem_reg[3][4]/P0001 , \u10_mem_reg[3][5]/P0001 , \u10_mem_reg[3][6]/P0001 , \u10_mem_reg[3][7]/P0001 , \u10_mem_reg[3][8]/P0001 , \u10_mem_reg[3][9]/P0001 , \u10_rp_reg[0]/P0001 , \u10_rp_reg[1]/P0001 , \u10_rp_reg[2]/P0001 , \u10_status_reg[0]/P0001 , \u10_status_reg[1]/P0001 , \u10_wp_reg[0]/NET0131 , \u10_wp_reg[1]/P0001 , \u10_wp_reg[2]/P0001 , \u10_wp_reg[3]/P0001 , \u11_din_tmp1_reg[0]/P0001 , \u11_din_tmp1_reg[10]/P0001 , \u11_din_tmp1_reg[11]/P0001 , \u11_din_tmp1_reg[12]/P0001 , \u11_din_tmp1_reg[13]/P0001 , \u11_din_tmp1_reg[14]/P0001 , \u11_din_tmp1_reg[15]/P0001 , \u11_din_tmp1_reg[1]/P0001 , \u11_din_tmp1_reg[2]/P0001 , \u11_din_tmp1_reg[3]/P0001 , \u11_din_tmp1_reg[4]/P0001 , \u11_din_tmp1_reg[5]/P0001 , \u11_din_tmp1_reg[6]/P0001 , \u11_din_tmp1_reg[7]/P0001 , \u11_din_tmp1_reg[8]/P0001 , \u11_din_tmp1_reg[9]/P0001 , \u11_dout_reg[0]/P0001 , \u11_dout_reg[10]/P0001 , \u11_dout_reg[11]/P0001 , \u11_dout_reg[12]/P0001 , \u11_dout_reg[13]/P0001 , \u11_dout_reg[14]/P0001 , \u11_dout_reg[15]/P0001 , \u11_dout_reg[16]/P0001 , \u11_dout_reg[17]/P0001 , \u11_dout_reg[18]/P0001 , \u11_dout_reg[19]/P0001 , \u11_dout_reg[1]/P0001 , \u11_dout_reg[20]/P0001 , \u11_dout_reg[21]/P0001 , \u11_dout_reg[22]/P0001 , \u11_dout_reg[23]/P0001 , \u11_dout_reg[24]/P0001 , \u11_dout_reg[25]/P0001 , \u11_dout_reg[26]/P0001 , \u11_dout_reg[27]/P0001 , \u11_dout_reg[28]/P0001 , \u11_dout_reg[29]/P0001 , \u11_dout_reg[2]/P0001 , \u11_dout_reg[30]/P0001 , \u11_dout_reg[31]/P0001 , \u11_dout_reg[3]/P0001 , \u11_dout_reg[4]/P0001 , \u11_dout_reg[5]/P0001 , \u11_dout_reg[6]/P0001 , \u11_dout_reg[7]/P0001 , \u11_dout_reg[8]/P0001 , \u11_dout_reg[9]/P0001 , \u11_empty_reg/P0001 , \u11_full_reg/NET0131 , \u11_mem_reg[0][0]/P0001 , \u11_mem_reg[0][10]/P0001 , \u11_mem_reg[0][11]/P0001 , \u11_mem_reg[0][12]/P0001 , \u11_mem_reg[0][13]/P0001 , \u11_mem_reg[0][14]/P0001 , \u11_mem_reg[0][15]/P0001 , \u11_mem_reg[0][16]/P0001 , \u11_mem_reg[0][17]/P0001 , \u11_mem_reg[0][18]/P0001 , \u11_mem_reg[0][19]/P0001 , \u11_mem_reg[0][1]/P0001 , \u11_mem_reg[0][20]/P0001 , \u11_mem_reg[0][21]/P0001 , \u11_mem_reg[0][22]/P0001 , \u11_mem_reg[0][23]/P0001 , \u11_mem_reg[0][24]/P0001 , \u11_mem_reg[0][25]/P0001 , \u11_mem_reg[0][26]/P0001 , \u11_mem_reg[0][27]/P0001 , \u11_mem_reg[0][28]/P0001 , \u11_mem_reg[0][29]/P0001 , \u11_mem_reg[0][2]/P0001 , \u11_mem_reg[0][30]/P0001 , \u11_mem_reg[0][31]/P0001 , \u11_mem_reg[0][3]/P0001 , \u11_mem_reg[0][4]/P0001 , \u11_mem_reg[0][5]/P0001 , \u11_mem_reg[0][6]/P0001 , \u11_mem_reg[0][7]/P0001 , \u11_mem_reg[0][8]/P0001 , \u11_mem_reg[0][9]/P0001 , \u11_mem_reg[1][0]/P0001 , \u11_mem_reg[1][10]/P0001 , \u11_mem_reg[1][11]/P0001 , \u11_mem_reg[1][12]/P0001 , \u11_mem_reg[1][13]/P0001 , \u11_mem_reg[1][14]/P0001 , \u11_mem_reg[1][15]/P0001 , \u11_mem_reg[1][16]/P0001 , \u11_mem_reg[1][17]/P0001 , \u11_mem_reg[1][18]/P0001 , \u11_mem_reg[1][19]/P0001 , \u11_mem_reg[1][1]/P0001 , \u11_mem_reg[1][20]/P0001 , \u11_mem_reg[1][21]/P0001 , \u11_mem_reg[1][22]/P0001 , \u11_mem_reg[1][23]/P0001 , \u11_mem_reg[1][24]/P0001 , \u11_mem_reg[1][25]/P0001 , \u11_mem_reg[1][26]/P0001 , \u11_mem_reg[1][27]/P0001 , \u11_mem_reg[1][28]/P0001 , \u11_mem_reg[1][29]/P0001 , \u11_mem_reg[1][2]/P0001 , \u11_mem_reg[1][30]/P0001 , \u11_mem_reg[1][31]/P0001 , \u11_mem_reg[1][3]/P0001 , \u11_mem_reg[1][4]/P0001 , \u11_mem_reg[1][5]/P0001 , \u11_mem_reg[1][6]/P0001 , \u11_mem_reg[1][7]/P0001 , \u11_mem_reg[1][8]/P0001 , \u11_mem_reg[1][9]/P0001 , \u11_mem_reg[2][0]/P0001 , \u11_mem_reg[2][10]/P0001 , \u11_mem_reg[2][11]/P0001 , \u11_mem_reg[2][12]/P0001 , \u11_mem_reg[2][13]/P0001 , \u11_mem_reg[2][14]/P0001 , \u11_mem_reg[2][15]/P0001 , \u11_mem_reg[2][16]/P0001 , \u11_mem_reg[2][17]/P0001 , \u11_mem_reg[2][18]/P0001 , \u11_mem_reg[2][19]/P0001 , \u11_mem_reg[2][1]/P0001 , \u11_mem_reg[2][20]/P0001 , \u11_mem_reg[2][21]/P0001 , \u11_mem_reg[2][22]/P0001 , \u11_mem_reg[2][23]/P0001 , \u11_mem_reg[2][24]/P0001 , \u11_mem_reg[2][25]/P0001 , \u11_mem_reg[2][26]/P0001 , \u11_mem_reg[2][27]/P0001 , \u11_mem_reg[2][28]/P0001 , \u11_mem_reg[2][29]/P0001 , \u11_mem_reg[2][2]/P0001 , \u11_mem_reg[2][30]/P0001 , \u11_mem_reg[2][31]/P0001 , \u11_mem_reg[2][3]/P0001 , \u11_mem_reg[2][4]/P0001 , \u11_mem_reg[2][5]/P0001 , \u11_mem_reg[2][6]/P0001 , \u11_mem_reg[2][7]/P0001 , \u11_mem_reg[2][8]/P0001 , \u11_mem_reg[2][9]/P0001 , \u11_mem_reg[3][0]/P0001 , \u11_mem_reg[3][10]/P0001 , \u11_mem_reg[3][11]/P0001 , \u11_mem_reg[3][12]/P0001 , \u11_mem_reg[3][13]/P0001 , \u11_mem_reg[3][14]/P0001 , \u11_mem_reg[3][15]/P0001 , \u11_mem_reg[3][16]/P0001 , \u11_mem_reg[3][17]/P0001 , \u11_mem_reg[3][18]/P0001 , \u11_mem_reg[3][19]/P0001 , \u11_mem_reg[3][1]/P0001 , \u11_mem_reg[3][20]/P0001 , \u11_mem_reg[3][21]/P0001 , \u11_mem_reg[3][22]/P0001 , \u11_mem_reg[3][23]/P0001 , \u11_mem_reg[3][24]/P0001 , \u11_mem_reg[3][25]/P0001 , \u11_mem_reg[3][26]/P0001 , \u11_mem_reg[3][27]/P0001 , \u11_mem_reg[3][28]/P0001 , \u11_mem_reg[3][29]/P0001 , \u11_mem_reg[3][2]/P0001 , \u11_mem_reg[3][30]/P0001 , \u11_mem_reg[3][31]/P0001 , \u11_mem_reg[3][3]/P0001 , \u11_mem_reg[3][4]/P0001 , \u11_mem_reg[3][5]/P0001 , \u11_mem_reg[3][6]/P0001 , \u11_mem_reg[3][7]/P0001 , \u11_mem_reg[3][8]/P0001 , \u11_mem_reg[3][9]/P0001 , \u11_rp_reg[0]/P0001 , \u11_rp_reg[1]/P0001 , \u11_rp_reg[2]/P0001 , \u11_status_reg[0]/P0001 , \u11_status_reg[1]/P0001 , \u11_wp_reg[0]/NET0131 , \u11_wp_reg[1]/P0001 , \u11_wp_reg[2]/P0001 , \u11_wp_reg[3]/P0001 , \u12_dout_reg[0]/P0001 , \u12_dout_reg[10]/P0001 , \u12_dout_reg[11]/P0001 , \u12_dout_reg[12]/P0001 , \u12_dout_reg[13]/P0001 , \u12_dout_reg[14]/P0001 , \u12_dout_reg[15]/P0001 , \u12_dout_reg[16]/P0001 , \u12_dout_reg[17]/P0001 , \u12_dout_reg[18]/P0001 , \u12_dout_reg[19]/P0001 , \u12_dout_reg[1]/P0001 , \u12_dout_reg[20]/P0001 , \u12_dout_reg[21]/P0001 , \u12_dout_reg[22]/P0001 , \u12_dout_reg[23]/P0001 , \u12_dout_reg[24]/P0001 , \u12_dout_reg[25]/P0001 , \u12_dout_reg[26]/P0001 , \u12_dout_reg[27]/P0001 , \u12_dout_reg[28]/P0001 , \u12_dout_reg[29]/P0001 , \u12_dout_reg[2]/P0001 , \u12_dout_reg[30]/P0001 , \u12_dout_reg[31]/P0001 , \u12_dout_reg[3]/P0001 , \u12_dout_reg[4]/P0001 , \u12_dout_reg[5]/P0001 , \u12_dout_reg[6]/P0001 , \u12_dout_reg[7]/P0001 , \u12_dout_reg[8]/P0001 , \u12_dout_reg[9]/P0001 , \u12_i3_re_reg/NET0131 , \u12_i4_re_reg/P0001 , \u12_i6_re_reg/NET0131 , \u12_o3_we_reg/P0001 , \u12_o4_we_reg/P0001 , \u12_o6_we_reg/P0001 , \u12_o7_we_reg/P0001 , \u12_o8_we_reg/P0001 , \u12_o9_we_reg/P0001 , \u12_re1_reg/P0001 , \u12_re2_reg/NET0131 , \u12_rf_we_reg/P0001 , \u12_we1_reg/P0001 , \u12_we2_reg/P0001 , \u13_ac97_rst_force_reg/P0001 , \u13_crac_dout_r_reg[0]/P0001 , \u13_crac_dout_r_reg[10]/P0001 , \u13_crac_dout_r_reg[11]/P0001 , \u13_crac_dout_r_reg[12]/P0001 , \u13_crac_dout_r_reg[13]/P0001 , \u13_crac_dout_r_reg[14]/P0001 , \u13_crac_dout_r_reg[15]/P0001 , \u13_crac_dout_r_reg[1]/P0001 , \u13_crac_dout_r_reg[2]/P0001 , \u13_crac_dout_r_reg[3]/P0001 , \u13_crac_dout_r_reg[4]/P0001 , \u13_crac_dout_r_reg[5]/P0001 , \u13_crac_dout_r_reg[6]/P0001 , \u13_crac_dout_r_reg[7]/P0001 , \u13_crac_dout_r_reg[8]/P0001 , \u13_crac_dout_r_reg[9]/P0001 , \u13_crac_r_reg[0]/NET0131 , \u13_crac_r_reg[1]/NET0131 , \u13_crac_r_reg[2]/NET0131 , \u13_crac_r_reg[3]/NET0131 , \u13_crac_r_reg[4]/NET0131 , \u13_crac_r_reg[5]/NET0131 , \u13_crac_r_reg[6]/NET0131 , \u13_crac_r_reg[7]/NET0131 , \u13_icc_r_reg[0]/NET0131 , \u13_icc_r_reg[10]/NET0131 , \u13_icc_r_reg[11]/NET0131 , \u13_icc_r_reg[12]/NET0131 , \u13_icc_r_reg[13]/NET0131 , \u13_icc_r_reg[14]/NET0131 , \u13_icc_r_reg[15]/NET0131 , \u13_icc_r_reg[16]/NET0131 , \u13_icc_r_reg[17]/NET0131 , \u13_icc_r_reg[18]/NET0131 , \u13_icc_r_reg[19]/NET0131 , \u13_icc_r_reg[1]/NET0131 , \u13_icc_r_reg[20]/NET0131 , \u13_icc_r_reg[21]/NET0131 , \u13_icc_r_reg[22]/NET0131 , \u13_icc_r_reg[23]/NET0131 , \u13_icc_r_reg[2]/NET0131 , \u13_icc_r_reg[3]/NET0131 , \u13_icc_r_reg[4]/NET0131 , \u13_icc_r_reg[5]/NET0131 , \u13_icc_r_reg[6]/NET0131 , \u13_icc_r_reg[7]/NET0131 , \u13_icc_r_reg[8]/NET0131 , \u13_icc_r_reg[9]/NET0131 , \u13_intm_r_reg[0]/NET0131 , \u13_intm_r_reg[10]/NET0131 , \u13_intm_r_reg[11]/NET0131 , \u13_intm_r_reg[12]/NET0131 , \u13_intm_r_reg[13]/NET0131 , \u13_intm_r_reg[14]/NET0131 , \u13_intm_r_reg[15]/NET0131 , \u13_intm_r_reg[16]/NET0131 , \u13_intm_r_reg[17]/NET0131 , \u13_intm_r_reg[18]/NET0131 , \u13_intm_r_reg[19]/NET0131 , \u13_intm_r_reg[1]/NET0131 , \u13_intm_r_reg[20]/NET0131 , \u13_intm_r_reg[21]/NET0131 , \u13_intm_r_reg[22]/NET0131 , \u13_intm_r_reg[23]/NET0131 , \u13_intm_r_reg[24]/NET0131 , \u13_intm_r_reg[25]/NET0131 , \u13_intm_r_reg[26]/NET0131 , \u13_intm_r_reg[27]/NET0131 , \u13_intm_r_reg[28]/NET0131 , \u13_intm_r_reg[2]/NET0131 , \u13_intm_r_reg[3]/NET0131 , \u13_intm_r_reg[4]/NET0131 , \u13_intm_r_reg[5]/NET0131 , \u13_intm_r_reg[6]/NET0131 , \u13_intm_r_reg[7]/NET0131 , \u13_intm_r_reg[8]/NET0131 , \u13_intm_r_reg[9]/NET0131 , \u13_ints_r_reg[0]/NET0131 , \u13_ints_r_reg[10]/NET0131 , \u13_ints_r_reg[11]/NET0131 , \u13_ints_r_reg[12]/NET0131 , \u13_ints_r_reg[13]/NET0131 , \u13_ints_r_reg[14]/NET0131 , \u13_ints_r_reg[15]/NET0131 , \u13_ints_r_reg[16]/NET0131 , \u13_ints_r_reg[17]/NET0131 , \u13_ints_r_reg[18]/NET0131 , \u13_ints_r_reg[19]/NET0131 , \u13_ints_r_reg[1]/NET0131 , \u13_ints_r_reg[20]/NET0131 , \u13_ints_r_reg[21]/NET0131 , \u13_ints_r_reg[22]/NET0131 , \u13_ints_r_reg[23]/NET0131 , \u13_ints_r_reg[24]/NET0131 , \u13_ints_r_reg[25]/NET0131 , \u13_ints_r_reg[26]/NET0131 , \u13_ints_r_reg[27]/NET0131 , \u13_ints_r_reg[28]/NET0131 , \u13_ints_r_reg[2]/NET0131 , \u13_ints_r_reg[3]/NET0131 , \u13_ints_r_reg[4]/NET0131 , \u13_ints_r_reg[5]/NET0131 , \u13_ints_r_reg[6]/NET0131 , \u13_ints_r_reg[7]/NET0131 , \u13_ints_r_reg[8]/NET0131 , \u13_ints_r_reg[9]/NET0131 , \u13_occ0_r_reg[0]/NET0131 , \u13_occ0_r_reg[10]/NET0131 , \u13_occ0_r_reg[11]/NET0131 , \u13_occ0_r_reg[12]/NET0131 , \u13_occ0_r_reg[13]/NET0131 , \u13_occ0_r_reg[14]/NET0131 , \u13_occ0_r_reg[15]/NET0131 , \u13_occ0_r_reg[16]/NET0131 , \u13_occ0_r_reg[17]/NET0131 , \u13_occ0_r_reg[18]/NET0131 , \u13_occ0_r_reg[19]/NET0131 , \u13_occ0_r_reg[1]/NET0131 , \u13_occ0_r_reg[20]/NET0131 , \u13_occ0_r_reg[21]/NET0131 , \u13_occ0_r_reg[22]/NET0131 , \u13_occ0_r_reg[23]/NET0131 , \u13_occ0_r_reg[24]/NET0131 , \u13_occ0_r_reg[25]/NET0131 , \u13_occ0_r_reg[26]/NET0131 , \u13_occ0_r_reg[27]/NET0131 , \u13_occ0_r_reg[28]/NET0131 , \u13_occ0_r_reg[29]/NET0131 , \u13_occ0_r_reg[2]/NET0131 , \u13_occ0_r_reg[30]/NET0131 , \u13_occ0_r_reg[31]/NET0131 , \u13_occ0_r_reg[3]/NET0131 , \u13_occ0_r_reg[4]/NET0131 , \u13_occ0_r_reg[5]/NET0131 , \u13_occ0_r_reg[6]/NET0131 , \u13_occ0_r_reg[7]/NET0131 , \u13_occ0_r_reg[8]/NET0131 , \u13_occ0_r_reg[9]/NET0131 , \u13_occ1_r_reg[0]/NET0131 , \u13_occ1_r_reg[10]/NET0131 , \u13_occ1_r_reg[11]/NET0131 , \u13_occ1_r_reg[12]/NET0131 , \u13_occ1_r_reg[13]/NET0131 , \u13_occ1_r_reg[14]/NET0131 , \u13_occ1_r_reg[15]/NET0131 , \u13_occ1_r_reg[1]/NET0131 , \u13_occ1_r_reg[2]/NET0131 , \u13_occ1_r_reg[3]/NET0131 , \u13_occ1_r_reg[4]/NET0131 , \u13_occ1_r_reg[5]/NET0131 , \u13_occ1_r_reg[6]/NET0131 , \u13_occ1_r_reg[7]/NET0131 , \u13_occ1_r_reg[8]/NET0131 , \u13_occ1_r_reg[9]/NET0131 , \u13_resume_req_reg/P0001 , \u14_crac_valid_r_reg/P0001 , \u14_crac_wr_r_reg/P0001 , \u14_u0_en_out_l2_reg/P0001 , \u14_u0_en_out_l_reg/NET0131 , \u14_u0_full_empty_r_reg/P0001 , \u14_u1_en_out_l2_reg/P0001 , \u14_u1_en_out_l_reg/NET0131 , \u14_u1_full_empty_r_reg/P0001 , \u14_u2_en_out_l2_reg/P0001 , \u14_u2_en_out_l_reg/NET0131 , \u14_u2_full_empty_r_reg/P0001 , \u14_u3_en_out_l2_reg/P0001 , \u14_u3_en_out_l_reg/NET0131 , \u14_u3_full_empty_r_reg/P0001 , \u14_u4_en_out_l2_reg/P0001 , \u14_u4_en_out_l_reg/NET0131 , \u14_u4_full_empty_r_reg/P0001 , \u14_u5_en_out_l2_reg/P0001 , \u14_u5_en_out_l_reg/NET0131 , \u14_u5_full_empty_r_reg/P0001 , \u14_u6_en_out_l2_reg/P0001 , \u14_u6_en_out_l_reg/NET0131 , \u14_u6_full_empty_r_reg/P0001 , \u14_u7_en_out_l2_reg/P0001 , \u14_u7_en_out_l_reg/NET0131 , \u14_u7_full_empty_r_reg/P0001 , \u14_u8_en_out_l2_reg/P0001 , \u14_u8_en_out_l_reg/NET0131 , \u14_u8_full_empty_r_reg/P0001 , \u15_crac_din_reg[0]/NET0131 , \u15_crac_din_reg[10]/NET0131 , \u15_crac_din_reg[11]/NET0131 , \u15_crac_din_reg[12]/NET0131 , \u15_crac_din_reg[13]/NET0131 , \u15_crac_din_reg[14]/NET0131 , \u15_crac_din_reg[15]/NET0131 , \u15_crac_din_reg[1]/NET0131 , \u15_crac_din_reg[2]/NET0131 , \u15_crac_din_reg[3]/NET0131 , \u15_crac_din_reg[4]/NET0131 , \u15_crac_din_reg[5]/NET0131 , \u15_crac_din_reg[6]/NET0131 , \u15_crac_din_reg[7]/NET0131 , \u15_crac_din_reg[8]/NET0131 , \u15_crac_din_reg[9]/NET0131 , \u15_crac_rd_done_reg/P0001 , \u15_crac_rd_reg/NET0131 , \u15_crac_we_r_reg/P0001 , \u15_crac_wr_reg/NET0131 , \u15_rdd1_reg/NET0131 , \u15_rdd2_reg/NET0131 , \u15_rdd3_reg/NET0131 , \u15_valid_r_reg/P0001 , \u16_u0_dma_req_r1_reg/P0001 , \u16_u1_dma_req_r1_reg/P0001 , \u16_u2_dma_req_r1_reg/P0001 , \u16_u3_dma_req_r1_reg/P0001 , \u16_u4_dma_req_r1_reg/P0001 , \u16_u5_dma_req_r1_reg/P0001 , \u16_u6_dma_req_r1_reg/P0001 , \u16_u7_dma_req_r1_reg/P0001 , \u16_u8_dma_req_r1_reg/P0001 , \u17_int_set_reg[0]/NET0131 , \u17_int_set_reg[1]/NET0131 , \u17_int_set_reg[2]/NET0131 , \u18_int_set_reg[0]/NET0131 , \u18_int_set_reg[1]/NET0131 , \u18_int_set_reg[2]/NET0131 , \u19_int_set_reg[0]/NET0131 , \u19_int_set_reg[1]/NET0131 , \u19_int_set_reg[2]/NET0131 , \u1_slt0_reg[11]/P0001 , \u1_slt0_reg[12]/P0001 , \u1_slt0_reg[15]/P0001 , \u1_slt0_reg[9]/P0001 , \u1_slt1_reg[10]/P0001 , \u1_slt1_reg[11]/P0001 , \u1_slt1_reg[5]/P0001 , \u1_slt1_reg[6]/P0001 , \u1_slt1_reg[7]/P0001 , \u1_slt1_reg[8]/P0001 , \u1_slt3_reg[0]/P0001 , \u1_slt3_reg[10]/P0001 , \u1_slt3_reg[11]/P0001 , \u1_slt3_reg[12]/P0001 , \u1_slt3_reg[13]/P0001 , \u1_slt3_reg[14]/P0001 , \u1_slt3_reg[15]/P0001 , \u1_slt3_reg[16]/P0001 , \u1_slt3_reg[17]/P0001 , \u1_slt3_reg[18]/P0001 , \u1_slt3_reg[19]/P0001 , \u1_slt3_reg[1]/P0001 , \u1_slt3_reg[2]/P0001 , \u1_slt3_reg[3]/P0001 , \u1_slt3_reg[4]/P0001 , \u1_slt3_reg[5]/P0001 , \u1_slt3_reg[6]/P0001 , \u1_slt3_reg[7]/P0001 , \u1_slt3_reg[8]/P0001 , \u1_slt3_reg[9]/P0001 , \u1_slt4_reg[0]/P0001 , \u1_slt4_reg[10]/P0001 , \u1_slt4_reg[11]/P0001 , \u1_slt4_reg[12]/P0001 , \u1_slt4_reg[13]/P0001 , \u1_slt4_reg[14]/P0001 , \u1_slt4_reg[15]/P0001 , \u1_slt4_reg[16]/P0001 , \u1_slt4_reg[17]/P0001 , \u1_slt4_reg[18]/P0001 , \u1_slt4_reg[19]/P0001 , \u1_slt4_reg[1]/P0001 , \u1_slt4_reg[2]/P0001 , \u1_slt4_reg[3]/P0001 , \u1_slt4_reg[4]/P0001 , \u1_slt4_reg[5]/P0001 , \u1_slt4_reg[6]/P0001 , \u1_slt4_reg[7]/P0001 , \u1_slt4_reg[8]/P0001 , \u1_slt4_reg[9]/P0001 , \u1_slt6_reg[0]/P0001 , \u1_slt6_reg[10]/P0001 , \u1_slt6_reg[11]/P0001 , \u1_slt6_reg[12]/P0001 , \u1_slt6_reg[13]/P0001 , \u1_slt6_reg[14]/P0001 , \u1_slt6_reg[15]/P0001 , \u1_slt6_reg[16]/P0001 , \u1_slt6_reg[17]/P0001 , \u1_slt6_reg[18]/P0001 , \u1_slt6_reg[19]/P0001 , \u1_slt6_reg[1]/P0001 , \u1_slt6_reg[2]/P0001 , \u1_slt6_reg[3]/P0001 , \u1_slt6_reg[4]/P0001 , \u1_slt6_reg[5]/P0001 , \u1_slt6_reg[6]/P0001 , \u1_slt6_reg[7]/P0001 , \u1_slt6_reg[8]/P0001 , \u1_slt6_reg[9]/P0001 , \u1_sr_reg[10]/P0001 , \u1_sr_reg[11]/P0001 , \u1_sr_reg[12]/P0001 , \u1_sr_reg[15]/P0001 , \u1_sr_reg[5]/P0001 , \u1_sr_reg[6]/P0001 , \u1_sr_reg[7]/P0001 , \u1_sr_reg[8]/P0001 , \u1_sr_reg[9]/P0001 , \u20_int_set_reg[0]/NET0131 , \u20_int_set_reg[1]/NET0131 , \u20_int_set_reg[2]/NET0131 , \u21_int_set_reg[0]/NET0131 , \u21_int_set_reg[1]/NET0131 , \u21_int_set_reg[2]/NET0131 , \u22_int_set_reg[0]/NET0131 , \u22_int_set_reg[1]/NET0131 , \u22_int_set_reg[2]/NET0131 , \u23_int_set_reg[0]/NET0131 , \u23_int_set_reg[1]/NET0131 , \u23_int_set_reg[2]/NET0131 , \u24_int_set_reg[0]/NET0131 , \u24_int_set_reg[1]/NET0131 , \u24_int_set_reg[2]/NET0131 , \u25_int_set_reg[0]/NET0131 , \u25_int_set_reg[1]/NET0131 , \u25_int_set_reg[2]/NET0131 , \u26_cnt_reg[0]/NET0131 , \u26_cnt_reg[1]/NET0131 , \u26_cnt_reg[2]/NET0131 , \u26_ps_cnt_reg[0]/NET0131 , \u26_ps_cnt_reg[1]/NET0131 , \u26_ps_cnt_reg[2]/NET0131 , \u26_ps_cnt_reg[3]/NET0131 , \u26_ps_cnt_reg[4]/NET0131 , \u26_ps_cnt_reg[5]/NET0131 , \u2_bit_clk_e_reg/P0001 , \u2_bit_clk_r1_reg/P0001 , \u2_bit_clk_r_reg/P0001 , \u2_cnt_reg[0]/NET0131 , \u2_cnt_reg[1]/NET0131 , \u2_cnt_reg[2]/NET0131 , \u2_cnt_reg[3]/NET0131 , \u2_cnt_reg[4]/NET0131 , \u2_cnt_reg[5]/NET0131 , \u2_cnt_reg[6]/NET0131 , \u2_cnt_reg[7]/NET0131 , \u2_ld_reg/P0001 , \u2_out_le_reg[0]/P0001 , \u2_out_le_reg[1]/P0001 , \u2_res_cnt_reg[0]/P0001 , \u2_res_cnt_reg[1]/P0001 , \u2_res_cnt_reg[2]/P0001 , \u2_res_cnt_reg[3]/P0001 , \u2_sync_beat_reg/P0001 , \u2_sync_resume_reg/NET0131 , \u2_to_cnt_reg[0]/NET0131 , \u2_to_cnt_reg[1]/NET0131 , \u2_to_cnt_reg[2]/NET0131 , \u2_to_cnt_reg[3]/NET0131 , \u2_to_cnt_reg[4]/NET0131 , \u2_to_cnt_reg[5]/NET0131 , \u3_dout_reg[0]/P0001 , \u3_dout_reg[10]/P0001 , \u3_dout_reg[11]/P0001 , \u3_dout_reg[12]/P0001 , \u3_dout_reg[13]/P0001 , \u3_dout_reg[14]/P0001 , \u3_dout_reg[15]/P0001 , \u3_dout_reg[16]/P0001 , \u3_dout_reg[17]/P0001 , \u3_dout_reg[18]/P0001 , \u3_dout_reg[19]/P0001 , \u3_dout_reg[1]/P0001 , \u3_dout_reg[2]/P0001 , \u3_dout_reg[3]/P0001 , \u3_dout_reg[4]/P0001 , \u3_dout_reg[5]/P0001 , \u3_dout_reg[6]/P0001 , \u3_dout_reg[7]/P0001 , \u3_dout_reg[8]/P0001 , \u3_dout_reg[9]/P0001 , \u3_empty_reg/NET0131 , \u3_mem_reg[0][0]/NET0131 , \u3_mem_reg[0][10]/NET0131 , \u3_mem_reg[0][11]/NET0131 , \u3_mem_reg[0][12]/NET0131 , \u3_mem_reg[0][13]/NET0131 , \u3_mem_reg[0][14]/NET0131 , \u3_mem_reg[0][15]/NET0131 , \u3_mem_reg[0][16]/NET0131 , \u3_mem_reg[0][17]/NET0131 , \u3_mem_reg[0][18]/NET0131 , \u3_mem_reg[0][19]/NET0131 , \u3_mem_reg[0][1]/NET0131 , \u3_mem_reg[0][20]/NET0131 , \u3_mem_reg[0][21]/NET0131 , \u3_mem_reg[0][22]/NET0131 , \u3_mem_reg[0][23]/NET0131 , \u3_mem_reg[0][24]/NET0131 , \u3_mem_reg[0][25]/NET0131 , \u3_mem_reg[0][26]/NET0131 , \u3_mem_reg[0][27]/NET0131 , \u3_mem_reg[0][28]/NET0131 , \u3_mem_reg[0][29]/NET0131 , \u3_mem_reg[0][2]/NET0131 , \u3_mem_reg[0][30]/NET0131 , \u3_mem_reg[0][31]/NET0131 , \u3_mem_reg[0][3]/NET0131 , \u3_mem_reg[0][4]/NET0131 , \u3_mem_reg[0][5]/NET0131 , \u3_mem_reg[0][6]/NET0131 , \u3_mem_reg[0][7]/NET0131 , \u3_mem_reg[0][8]/NET0131 , \u3_mem_reg[0][9]/NET0131 , \u3_mem_reg[1][0]/NET0131 , \u3_mem_reg[1][10]/NET0131 , \u3_mem_reg[1][11]/NET0131 , \u3_mem_reg[1][12]/NET0131 , \u3_mem_reg[1][13]/NET0131 , \u3_mem_reg[1][14]/NET0131 , \u3_mem_reg[1][15]/NET0131 , \u3_mem_reg[1][16]/NET0131 , \u3_mem_reg[1][17]/NET0131 , \u3_mem_reg[1][18]/NET0131 , \u3_mem_reg[1][19]/NET0131 , \u3_mem_reg[1][1]/NET0131 , \u3_mem_reg[1][20]/NET0131 , \u3_mem_reg[1][21]/NET0131 , \u3_mem_reg[1][22]/NET0131 , \u3_mem_reg[1][23]/NET0131 , \u3_mem_reg[1][24]/NET0131 , \u3_mem_reg[1][25]/NET0131 , \u3_mem_reg[1][26]/NET0131 , \u3_mem_reg[1][27]/NET0131 , \u3_mem_reg[1][28]/NET0131 , \u3_mem_reg[1][29]/NET0131 , \u3_mem_reg[1][2]/NET0131 , \u3_mem_reg[1][30]/NET0131 , \u3_mem_reg[1][31]/NET0131 , \u3_mem_reg[1][3]/NET0131 , \u3_mem_reg[1][4]/NET0131 , \u3_mem_reg[1][5]/NET0131 , \u3_mem_reg[1][6]/NET0131 , \u3_mem_reg[1][7]/NET0131 , \u3_mem_reg[1][8]/NET0131 , \u3_mem_reg[1][9]/NET0131 , \u3_mem_reg[2][0]/NET0131 , \u3_mem_reg[2][10]/NET0131 , \u3_mem_reg[2][11]/NET0131 , \u3_mem_reg[2][12]/NET0131 , \u3_mem_reg[2][13]/NET0131 , \u3_mem_reg[2][14]/NET0131 , \u3_mem_reg[2][15]/NET0131 , \u3_mem_reg[2][16]/NET0131 , \u3_mem_reg[2][17]/NET0131 , \u3_mem_reg[2][18]/NET0131 , \u3_mem_reg[2][19]/NET0131 , \u3_mem_reg[2][1]/NET0131 , \u3_mem_reg[2][20]/NET0131 , \u3_mem_reg[2][21]/NET0131 , \u3_mem_reg[2][22]/NET0131 , \u3_mem_reg[2][23]/NET0131 , \u3_mem_reg[2][24]/NET0131 , \u3_mem_reg[2][25]/NET0131 , \u3_mem_reg[2][26]/NET0131 , \u3_mem_reg[2][27]/NET0131 , \u3_mem_reg[2][28]/NET0131 , \u3_mem_reg[2][29]/NET0131 , \u3_mem_reg[2][2]/NET0131 , \u3_mem_reg[2][30]/NET0131 , \u3_mem_reg[2][31]/NET0131 , \u3_mem_reg[2][3]/NET0131 , \u3_mem_reg[2][4]/NET0131 , \u3_mem_reg[2][5]/NET0131 , \u3_mem_reg[2][6]/NET0131 , \u3_mem_reg[2][7]/NET0131 , \u3_mem_reg[2][8]/NET0131 , \u3_mem_reg[2][9]/NET0131 , \u3_mem_reg[3][0]/NET0131 , \u3_mem_reg[3][10]/NET0131 , \u3_mem_reg[3][11]/NET0131 , \u3_mem_reg[3][12]/NET0131 , \u3_mem_reg[3][13]/NET0131 , \u3_mem_reg[3][14]/NET0131 , \u3_mem_reg[3][15]/NET0131 , \u3_mem_reg[3][16]/NET0131 , \u3_mem_reg[3][17]/NET0131 , \u3_mem_reg[3][18]/NET0131 , \u3_mem_reg[3][19]/NET0131 , \u3_mem_reg[3][1]/NET0131 , \u3_mem_reg[3][20]/NET0131 , \u3_mem_reg[3][21]/NET0131 , \u3_mem_reg[3][22]/NET0131 , \u3_mem_reg[3][23]/NET0131 , \u3_mem_reg[3][24]/NET0131 , \u3_mem_reg[3][25]/NET0131 , \u3_mem_reg[3][26]/NET0131 , \u3_mem_reg[3][27]/NET0131 , \u3_mem_reg[3][28]/NET0131 , \u3_mem_reg[3][29]/NET0131 , \u3_mem_reg[3][2]/NET0131 , \u3_mem_reg[3][30]/NET0131 , \u3_mem_reg[3][31]/NET0131 , \u3_mem_reg[3][3]/NET0131 , \u3_mem_reg[3][4]/NET0131 , \u3_mem_reg[3][5]/NET0131 , \u3_mem_reg[3][6]/NET0131 , \u3_mem_reg[3][7]/NET0131 , \u3_mem_reg[3][8]/NET0131 , \u3_mem_reg[3][9]/NET0131 , \u3_rp_reg[0]/P0001 , \u3_rp_reg[1]/NET0131 , \u3_rp_reg[2]/NET0131 , \u3_rp_reg[3]/NET0131 , \u3_status_reg[0]/P0001 , \u3_status_reg[1]/P0001 , \u3_wp_reg[0]/P0001 , \u3_wp_reg[1]/NET0131 , \u3_wp_reg[2]/P0001 , \u4_dout_reg[0]/P0001 , \u4_dout_reg[10]/P0001 , \u4_dout_reg[11]/P0001 , \u4_dout_reg[12]/P0001 , \u4_dout_reg[13]/P0001 , \u4_dout_reg[14]/P0001 , \u4_dout_reg[15]/P0001 , \u4_dout_reg[16]/P0001 , \u4_dout_reg[17]/P0001 , \u4_dout_reg[18]/P0001 , \u4_dout_reg[19]/P0001 , \u4_dout_reg[1]/P0001 , \u4_dout_reg[2]/P0001 , \u4_dout_reg[3]/P0001 , \u4_dout_reg[4]/P0001 , \u4_dout_reg[5]/P0001 , \u4_dout_reg[6]/P0001 , \u4_dout_reg[7]/P0001 , \u4_dout_reg[8]/P0001 , \u4_dout_reg[9]/P0001 , \u4_empty_reg/NET0131 , \u4_mem_reg[0][0]/NET0131 , \u4_mem_reg[0][10]/NET0131 , \u4_mem_reg[0][11]/NET0131 , \u4_mem_reg[0][12]/NET0131 , \u4_mem_reg[0][13]/NET0131 , \u4_mem_reg[0][14]/NET0131 , \u4_mem_reg[0][15]/NET0131 , \u4_mem_reg[0][16]/NET0131 , \u4_mem_reg[0][17]/NET0131 , \u4_mem_reg[0][18]/NET0131 , \u4_mem_reg[0][19]/NET0131 , \u4_mem_reg[0][1]/NET0131 , \u4_mem_reg[0][20]/NET0131 , \u4_mem_reg[0][21]/NET0131 , \u4_mem_reg[0][22]/NET0131 , \u4_mem_reg[0][23]/NET0131 , \u4_mem_reg[0][24]/NET0131 , \u4_mem_reg[0][25]/NET0131 , \u4_mem_reg[0][26]/NET0131 , \u4_mem_reg[0][27]/NET0131 , \u4_mem_reg[0][28]/NET0131 , \u4_mem_reg[0][29]/NET0131 , \u4_mem_reg[0][2]/NET0131 , \u4_mem_reg[0][30]/NET0131 , \u4_mem_reg[0][31]/NET0131 , \u4_mem_reg[0][3]/NET0131 , \u4_mem_reg[0][4]/NET0131 , \u4_mem_reg[0][5]/NET0131 , \u4_mem_reg[0][6]/NET0131 , \u4_mem_reg[0][7]/NET0131 , \u4_mem_reg[0][8]/NET0131 , \u4_mem_reg[0][9]/NET0131 , \u4_mem_reg[1][0]/NET0131 , \u4_mem_reg[1][10]/NET0131 , \u4_mem_reg[1][11]/NET0131 , \u4_mem_reg[1][12]/NET0131 , \u4_mem_reg[1][13]/NET0131 , \u4_mem_reg[1][14]/NET0131 , \u4_mem_reg[1][15]/NET0131 , \u4_mem_reg[1][16]/NET0131 , \u4_mem_reg[1][17]/NET0131 , \u4_mem_reg[1][18]/NET0131 , \u4_mem_reg[1][19]/NET0131 , \u4_mem_reg[1][1]/NET0131 , \u4_mem_reg[1][20]/NET0131 , \u4_mem_reg[1][21]/NET0131 , \u4_mem_reg[1][22]/NET0131 , \u4_mem_reg[1][23]/NET0131 , \u4_mem_reg[1][24]/NET0131 , \u4_mem_reg[1][25]/NET0131 , \u4_mem_reg[1][26]/NET0131 , \u4_mem_reg[1][27]/NET0131 , \u4_mem_reg[1][28]/NET0131 , \u4_mem_reg[1][29]/NET0131 , \u4_mem_reg[1][2]/NET0131 , \u4_mem_reg[1][30]/NET0131 , \u4_mem_reg[1][31]/NET0131 , \u4_mem_reg[1][3]/NET0131 , \u4_mem_reg[1][4]/NET0131 , \u4_mem_reg[1][5]/NET0131 , \u4_mem_reg[1][6]/NET0131 , \u4_mem_reg[1][7]/NET0131 , \u4_mem_reg[1][8]/NET0131 , \u4_mem_reg[1][9]/NET0131 , \u4_mem_reg[2][0]/NET0131 , \u4_mem_reg[2][10]/NET0131 , \u4_mem_reg[2][11]/NET0131 , \u4_mem_reg[2][12]/NET0131 , \u4_mem_reg[2][13]/NET0131 , \u4_mem_reg[2][14]/NET0131 , \u4_mem_reg[2][15]/NET0131 , \u4_mem_reg[2][16]/NET0131 , \u4_mem_reg[2][17]/NET0131 , \u4_mem_reg[2][18]/NET0131 , \u4_mem_reg[2][19]/NET0131 , \u4_mem_reg[2][1]/NET0131 , \u4_mem_reg[2][20]/NET0131 , \u4_mem_reg[2][21]/NET0131 , \u4_mem_reg[2][22]/NET0131 , \u4_mem_reg[2][23]/NET0131 , \u4_mem_reg[2][24]/NET0131 , \u4_mem_reg[2][25]/NET0131 , \u4_mem_reg[2][26]/NET0131 , \u4_mem_reg[2][27]/NET0131 , \u4_mem_reg[2][28]/NET0131 , \u4_mem_reg[2][29]/NET0131 , \u4_mem_reg[2][2]/NET0131 , \u4_mem_reg[2][30]/NET0131 , \u4_mem_reg[2][31]/NET0131 , \u4_mem_reg[2][3]/NET0131 , \u4_mem_reg[2][4]/NET0131 , \u4_mem_reg[2][5]/NET0131 , \u4_mem_reg[2][6]/NET0131 , \u4_mem_reg[2][7]/NET0131 , \u4_mem_reg[2][8]/NET0131 , \u4_mem_reg[2][9]/NET0131 , \u4_mem_reg[3][0]/NET0131 , \u4_mem_reg[3][10]/NET0131 , \u4_mem_reg[3][11]/NET0131 , \u4_mem_reg[3][12]/NET0131 , \u4_mem_reg[3][13]/NET0131 , \u4_mem_reg[3][14]/NET0131 , \u4_mem_reg[3][15]/NET0131 , \u4_mem_reg[3][16]/NET0131 , \u4_mem_reg[3][17]/NET0131 , \u4_mem_reg[3][18]/NET0131 , \u4_mem_reg[3][19]/NET0131 , \u4_mem_reg[3][1]/NET0131 , \u4_mem_reg[3][20]/NET0131 , \u4_mem_reg[3][21]/NET0131 , \u4_mem_reg[3][22]/NET0131 , \u4_mem_reg[3][23]/NET0131 , \u4_mem_reg[3][24]/NET0131 , \u4_mem_reg[3][25]/NET0131 , \u4_mem_reg[3][26]/NET0131 , \u4_mem_reg[3][27]/NET0131 , \u4_mem_reg[3][28]/NET0131 , \u4_mem_reg[3][29]/NET0131 , \u4_mem_reg[3][2]/NET0131 , \u4_mem_reg[3][30]/NET0131 , \u4_mem_reg[3][31]/NET0131 , \u4_mem_reg[3][3]/NET0131 , \u4_mem_reg[3][4]/NET0131 , \u4_mem_reg[3][5]/NET0131 , \u4_mem_reg[3][6]/NET0131 , \u4_mem_reg[3][7]/NET0131 , \u4_mem_reg[3][8]/NET0131 , \u4_mem_reg[3][9]/NET0131 , \u4_rp_reg[0]/P0001 , \u4_rp_reg[1]/NET0131 , \u4_rp_reg[2]/NET0131 , \u4_rp_reg[3]/NET0131 , \u4_status_reg[0]/P0001 , \u4_status_reg[1]/P0001 , \u4_wp_reg[0]/P0001 , \u4_wp_reg[1]/NET0131 , \u4_wp_reg[2]/P0001 , \u5_dout_reg[0]/P0001 , \u5_dout_reg[10]/P0001 , \u5_dout_reg[11]/P0001 , \u5_dout_reg[12]/P0001 , \u5_dout_reg[13]/P0001 , \u5_dout_reg[14]/P0001 , \u5_dout_reg[15]/P0001 , \u5_dout_reg[16]/P0001 , \u5_dout_reg[17]/P0001 , \u5_dout_reg[18]/P0001 , \u5_dout_reg[19]/P0001 , \u5_dout_reg[1]/P0001 , \u5_dout_reg[2]/P0001 , \u5_dout_reg[3]/P0001 , \u5_dout_reg[4]/P0001 , \u5_dout_reg[5]/P0001 , \u5_dout_reg[6]/P0001 , \u5_dout_reg[7]/P0001 , \u5_dout_reg[8]/P0001 , \u5_dout_reg[9]/P0001 , \u5_empty_reg/NET0131 , \u5_mem_reg[0][0]/NET0131 , \u5_mem_reg[0][10]/NET0131 , \u5_mem_reg[0][11]/NET0131 , \u5_mem_reg[0][12]/NET0131 , \u5_mem_reg[0][13]/NET0131 , \u5_mem_reg[0][14]/NET0131 , \u5_mem_reg[0][15]/NET0131 , \u5_mem_reg[0][16]/NET0131 , \u5_mem_reg[0][17]/NET0131 , \u5_mem_reg[0][18]/NET0131 , \u5_mem_reg[0][19]/NET0131 , \u5_mem_reg[0][1]/NET0131 , \u5_mem_reg[0][20]/NET0131 , \u5_mem_reg[0][21]/NET0131 , \u5_mem_reg[0][22]/NET0131 , \u5_mem_reg[0][23]/NET0131 , \u5_mem_reg[0][24]/NET0131 , \u5_mem_reg[0][25]/NET0131 , \u5_mem_reg[0][26]/NET0131 , \u5_mem_reg[0][27]/NET0131 , \u5_mem_reg[0][28]/NET0131 , \u5_mem_reg[0][29]/NET0131 , \u5_mem_reg[0][2]/NET0131 , \u5_mem_reg[0][30]/NET0131 , \u5_mem_reg[0][31]/NET0131 , \u5_mem_reg[0][3]/NET0131 , \u5_mem_reg[0][4]/NET0131 , \u5_mem_reg[0][5]/NET0131 , \u5_mem_reg[0][6]/NET0131 , \u5_mem_reg[0][7]/NET0131 , \u5_mem_reg[0][8]/NET0131 , \u5_mem_reg[0][9]/NET0131 , \u5_mem_reg[1][0]/NET0131 , \u5_mem_reg[1][10]/NET0131 , \u5_mem_reg[1][11]/NET0131 , \u5_mem_reg[1][12]/NET0131 , \u5_mem_reg[1][13]/NET0131 , \u5_mem_reg[1][14]/NET0131 , \u5_mem_reg[1][15]/NET0131 , \u5_mem_reg[1][16]/NET0131 , \u5_mem_reg[1][17]/NET0131 , \u5_mem_reg[1][18]/NET0131 , \u5_mem_reg[1][19]/NET0131 , \u5_mem_reg[1][1]/NET0131 , \u5_mem_reg[1][20]/NET0131 , \u5_mem_reg[1][21]/NET0131 , \u5_mem_reg[1][22]/NET0131 , \u5_mem_reg[1][23]/NET0131 , \u5_mem_reg[1][24]/NET0131 , \u5_mem_reg[1][25]/NET0131 , \u5_mem_reg[1][26]/NET0131 , \u5_mem_reg[1][27]/NET0131 , \u5_mem_reg[1][28]/NET0131 , \u5_mem_reg[1][29]/NET0131 , \u5_mem_reg[1][2]/NET0131 , \u5_mem_reg[1][30]/NET0131 , \u5_mem_reg[1][31]/NET0131 , \u5_mem_reg[1][3]/NET0131 , \u5_mem_reg[1][4]/NET0131 , \u5_mem_reg[1][5]/NET0131 , \u5_mem_reg[1][6]/NET0131 , \u5_mem_reg[1][7]/NET0131 , \u5_mem_reg[1][8]/NET0131 , \u5_mem_reg[1][9]/NET0131 , \u5_mem_reg[2][0]/NET0131 , \u5_mem_reg[2][10]/NET0131 , \u5_mem_reg[2][11]/NET0131 , \u5_mem_reg[2][12]/NET0131 , \u5_mem_reg[2][13]/NET0131 , \u5_mem_reg[2][14]/NET0131 , \u5_mem_reg[2][15]/NET0131 , \u5_mem_reg[2][16]/NET0131 , \u5_mem_reg[2][17]/NET0131 , \u5_mem_reg[2][18]/NET0131 , \u5_mem_reg[2][19]/NET0131 , \u5_mem_reg[2][1]/NET0131 , \u5_mem_reg[2][20]/NET0131 , \u5_mem_reg[2][21]/NET0131 , \u5_mem_reg[2][22]/NET0131 , \u5_mem_reg[2][23]/NET0131 , \u5_mem_reg[2][24]/NET0131 , \u5_mem_reg[2][25]/NET0131 , \u5_mem_reg[2][26]/NET0131 , \u5_mem_reg[2][27]/NET0131 , \u5_mem_reg[2][28]/NET0131 , \u5_mem_reg[2][29]/NET0131 , \u5_mem_reg[2][2]/NET0131 , \u5_mem_reg[2][30]/NET0131 , \u5_mem_reg[2][31]/NET0131 , \u5_mem_reg[2][3]/NET0131 , \u5_mem_reg[2][4]/NET0131 , \u5_mem_reg[2][5]/NET0131 , \u5_mem_reg[2][6]/NET0131 , \u5_mem_reg[2][7]/NET0131 , \u5_mem_reg[2][8]/NET0131 , \u5_mem_reg[2][9]/NET0131 , \u5_mem_reg[3][0]/NET0131 , \u5_mem_reg[3][10]/NET0131 , \u5_mem_reg[3][11]/NET0131 , \u5_mem_reg[3][12]/NET0131 , \u5_mem_reg[3][13]/NET0131 , \u5_mem_reg[3][14]/NET0131 , \u5_mem_reg[3][15]/NET0131 , \u5_mem_reg[3][16]/NET0131 , \u5_mem_reg[3][17]/NET0131 , \u5_mem_reg[3][18]/NET0131 , \u5_mem_reg[3][19]/NET0131 , \u5_mem_reg[3][1]/NET0131 , \u5_mem_reg[3][20]/NET0131 , \u5_mem_reg[3][21]/NET0131 , \u5_mem_reg[3][22]/NET0131 , \u5_mem_reg[3][23]/NET0131 , \u5_mem_reg[3][24]/NET0131 , \u5_mem_reg[3][25]/NET0131 , \u5_mem_reg[3][26]/NET0131 , \u5_mem_reg[3][27]/NET0131 , \u5_mem_reg[3][28]/NET0131 , \u5_mem_reg[3][29]/NET0131 , \u5_mem_reg[3][2]/NET0131 , \u5_mem_reg[3][30]/NET0131 , \u5_mem_reg[3][31]/NET0131 , \u5_mem_reg[3][3]/NET0131 , \u5_mem_reg[3][4]/NET0131 , \u5_mem_reg[3][5]/NET0131 , \u5_mem_reg[3][6]/NET0131 , \u5_mem_reg[3][7]/NET0131 , \u5_mem_reg[3][8]/NET0131 , \u5_mem_reg[3][9]/NET0131 , \u5_rp_reg[0]/P0001 , \u5_rp_reg[1]/NET0131 , \u5_rp_reg[2]/NET0131 , \u5_rp_reg[3]/NET0131 , \u5_status_reg[0]/P0001 , \u5_status_reg[1]/P0001 , \u5_wp_reg[0]/P0001 , \u5_wp_reg[1]/NET0131 , \u5_wp_reg[2]/P0001 , \u6_dout_reg[0]/P0001 , \u6_dout_reg[10]/P0001 , \u6_dout_reg[11]/P0001 , \u6_dout_reg[12]/P0001 , \u6_dout_reg[13]/P0001 , \u6_dout_reg[14]/P0001 , \u6_dout_reg[15]/P0001 , \u6_dout_reg[16]/P0001 , \u6_dout_reg[17]/P0001 , \u6_dout_reg[18]/P0001 , \u6_dout_reg[19]/P0001 , \u6_dout_reg[1]/P0001 , \u6_dout_reg[2]/P0001 , \u6_dout_reg[3]/P0001 , \u6_dout_reg[4]/P0001 , \u6_dout_reg[5]/P0001 , \u6_dout_reg[6]/P0001 , \u6_dout_reg[7]/P0001 , \u6_dout_reg[8]/P0001 , \u6_dout_reg[9]/P0001 , \u6_empty_reg/NET0131 , \u6_mem_reg[0][0]/NET0131 , \u6_mem_reg[0][10]/NET0131 , \u6_mem_reg[0][11]/NET0131 , \u6_mem_reg[0][12]/NET0131 , \u6_mem_reg[0][13]/NET0131 , \u6_mem_reg[0][14]/NET0131 , \u6_mem_reg[0][15]/NET0131 , \u6_mem_reg[0][16]/NET0131 , \u6_mem_reg[0][17]/NET0131 , \u6_mem_reg[0][18]/NET0131 , \u6_mem_reg[0][19]/NET0131 , \u6_mem_reg[0][1]/NET0131 , \u6_mem_reg[0][20]/NET0131 , \u6_mem_reg[0][21]/NET0131 , \u6_mem_reg[0][22]/NET0131 , \u6_mem_reg[0][23]/NET0131 , \u6_mem_reg[0][24]/NET0131 , \u6_mem_reg[0][25]/NET0131 , \u6_mem_reg[0][26]/NET0131 , \u6_mem_reg[0][27]/NET0131 , \u6_mem_reg[0][28]/NET0131 , \u6_mem_reg[0][29]/NET0131 , \u6_mem_reg[0][2]/NET0131 , \u6_mem_reg[0][30]/NET0131 , \u6_mem_reg[0][31]/NET0131 , \u6_mem_reg[0][3]/NET0131 , \u6_mem_reg[0][4]/NET0131 , \u6_mem_reg[0][5]/NET0131 , \u6_mem_reg[0][6]/NET0131 , \u6_mem_reg[0][7]/NET0131 , \u6_mem_reg[0][8]/NET0131 , \u6_mem_reg[0][9]/NET0131 , \u6_mem_reg[1][0]/NET0131 , \u6_mem_reg[1][10]/NET0131 , \u6_mem_reg[1][11]/NET0131 , \u6_mem_reg[1][12]/NET0131 , \u6_mem_reg[1][13]/NET0131 , \u6_mem_reg[1][14]/NET0131 , \u6_mem_reg[1][15]/NET0131 , \u6_mem_reg[1][16]/NET0131 , \u6_mem_reg[1][17]/NET0131 , \u6_mem_reg[1][18]/NET0131 , \u6_mem_reg[1][19]/NET0131 , \u6_mem_reg[1][1]/NET0131 , \u6_mem_reg[1][20]/NET0131 , \u6_mem_reg[1][21]/NET0131 , \u6_mem_reg[1][22]/NET0131 , \u6_mem_reg[1][23]/NET0131 , \u6_mem_reg[1][24]/NET0131 , \u6_mem_reg[1][25]/NET0131 , \u6_mem_reg[1][26]/NET0131 , \u6_mem_reg[1][27]/NET0131 , \u6_mem_reg[1][28]/NET0131 , \u6_mem_reg[1][29]/NET0131 , \u6_mem_reg[1][2]/NET0131 , \u6_mem_reg[1][30]/NET0131 , \u6_mem_reg[1][31]/NET0131 , \u6_mem_reg[1][3]/NET0131 , \u6_mem_reg[1][4]/NET0131 , \u6_mem_reg[1][5]/NET0131 , \u6_mem_reg[1][6]/NET0131 , \u6_mem_reg[1][7]/NET0131 , \u6_mem_reg[1][8]/NET0131 , \u6_mem_reg[1][9]/NET0131 , \u6_mem_reg[2][0]/NET0131 , \u6_mem_reg[2][10]/NET0131 , \u6_mem_reg[2][11]/NET0131 , \u6_mem_reg[2][12]/NET0131 , \u6_mem_reg[2][13]/NET0131 , \u6_mem_reg[2][14]/NET0131 , \u6_mem_reg[2][15]/NET0131 , \u6_mem_reg[2][16]/NET0131 , \u6_mem_reg[2][17]/NET0131 , \u6_mem_reg[2][18]/NET0131 , \u6_mem_reg[2][19]/NET0131 , \u6_mem_reg[2][1]/NET0131 , \u6_mem_reg[2][20]/NET0131 , \u6_mem_reg[2][21]/NET0131 , \u6_mem_reg[2][22]/NET0131 , \u6_mem_reg[2][23]/NET0131 , \u6_mem_reg[2][24]/NET0131 , \u6_mem_reg[2][25]/NET0131 , \u6_mem_reg[2][26]/NET0131 , \u6_mem_reg[2][27]/NET0131 , \u6_mem_reg[2][28]/NET0131 , \u6_mem_reg[2][29]/NET0131 , \u6_mem_reg[2][2]/NET0131 , \u6_mem_reg[2][30]/NET0131 , \u6_mem_reg[2][31]/NET0131 , \u6_mem_reg[2][3]/NET0131 , \u6_mem_reg[2][4]/NET0131 , \u6_mem_reg[2][5]/NET0131 , \u6_mem_reg[2][6]/NET0131 , \u6_mem_reg[2][7]/NET0131 , \u6_mem_reg[2][8]/NET0131 , \u6_mem_reg[2][9]/NET0131 , \u6_mem_reg[3][0]/NET0131 , \u6_mem_reg[3][10]/NET0131 , \u6_mem_reg[3][11]/NET0131 , \u6_mem_reg[3][12]/NET0131 , \u6_mem_reg[3][13]/NET0131 , \u6_mem_reg[3][14]/NET0131 , \u6_mem_reg[3][15]/NET0131 , \u6_mem_reg[3][16]/NET0131 , \u6_mem_reg[3][17]/NET0131 , \u6_mem_reg[3][18]/NET0131 , \u6_mem_reg[3][19]/NET0131 , \u6_mem_reg[3][1]/NET0131 , \u6_mem_reg[3][20]/NET0131 , \u6_mem_reg[3][21]/NET0131 , \u6_mem_reg[3][22]/NET0131 , \u6_mem_reg[3][23]/NET0131 , \u6_mem_reg[3][24]/NET0131 , \u6_mem_reg[3][25]/NET0131 , \u6_mem_reg[3][26]/NET0131 , \u6_mem_reg[3][27]/NET0131 , \u6_mem_reg[3][28]/NET0131 , \u6_mem_reg[3][29]/NET0131 , \u6_mem_reg[3][2]/NET0131 , \u6_mem_reg[3][30]/NET0131 , \u6_mem_reg[3][31]/NET0131 , \u6_mem_reg[3][3]/NET0131 , \u6_mem_reg[3][4]/NET0131 , \u6_mem_reg[3][5]/NET0131 , \u6_mem_reg[3][6]/NET0131 , \u6_mem_reg[3][7]/NET0131 , \u6_mem_reg[3][8]/NET0131 , \u6_mem_reg[3][9]/NET0131 , \u6_rp_reg[0]/P0001 , \u6_rp_reg[1]/NET0131 , \u6_rp_reg[2]/NET0131 , \u6_rp_reg[3]/NET0131 , \u6_status_reg[0]/P0001 , \u6_status_reg[1]/P0001 , \u6_wp_reg[0]/P0001 , \u6_wp_reg[1]/NET0131 , \u6_wp_reg[2]/P0001 , \u7_dout_reg[0]/P0001 , \u7_dout_reg[10]/P0001 , \u7_dout_reg[11]/P0001 , \u7_dout_reg[12]/P0001 , \u7_dout_reg[13]/P0001 , \u7_dout_reg[14]/P0001 , \u7_dout_reg[15]/P0001 , \u7_dout_reg[16]/P0001 , \u7_dout_reg[17]/P0001 , \u7_dout_reg[18]/P0001 , \u7_dout_reg[19]/P0001 , \u7_dout_reg[1]/P0001 , \u7_dout_reg[2]/P0001 , \u7_dout_reg[3]/P0001 , \u7_dout_reg[4]/P0001 , \u7_dout_reg[5]/P0001 , \u7_dout_reg[6]/P0001 , \u7_dout_reg[7]/P0001 , \u7_dout_reg[8]/P0001 , \u7_dout_reg[9]/P0001 , \u7_empty_reg/NET0131 , \u7_mem_reg[0][0]/NET0131 , \u7_mem_reg[0][10]/NET0131 , \u7_mem_reg[0][11]/NET0131 , \u7_mem_reg[0][12]/NET0131 , \u7_mem_reg[0][13]/NET0131 , \u7_mem_reg[0][14]/NET0131 , \u7_mem_reg[0][15]/NET0131 , \u7_mem_reg[0][16]/NET0131 , \u7_mem_reg[0][17]/NET0131 , \u7_mem_reg[0][18]/NET0131 , \u7_mem_reg[0][19]/NET0131 , \u7_mem_reg[0][1]/NET0131 , \u7_mem_reg[0][20]/NET0131 , \u7_mem_reg[0][21]/NET0131 , \u7_mem_reg[0][22]/NET0131 , \u7_mem_reg[0][23]/NET0131 , \u7_mem_reg[0][24]/NET0131 , \u7_mem_reg[0][25]/NET0131 , \u7_mem_reg[0][26]/NET0131 , \u7_mem_reg[0][27]/NET0131 , \u7_mem_reg[0][28]/NET0131 , \u7_mem_reg[0][29]/NET0131 , \u7_mem_reg[0][2]/NET0131 , \u7_mem_reg[0][30]/NET0131 , \u7_mem_reg[0][31]/NET0131 , \u7_mem_reg[0][3]/NET0131 , \u7_mem_reg[0][4]/NET0131 , \u7_mem_reg[0][5]/NET0131 , \u7_mem_reg[0][6]/NET0131 , \u7_mem_reg[0][7]/NET0131 , \u7_mem_reg[0][8]/NET0131 , \u7_mem_reg[0][9]/NET0131 , \u7_mem_reg[1][0]/NET0131 , \u7_mem_reg[1][10]/NET0131 , \u7_mem_reg[1][11]/NET0131 , \u7_mem_reg[1][12]/NET0131 , \u7_mem_reg[1][13]/NET0131 , \u7_mem_reg[1][14]/NET0131 , \u7_mem_reg[1][15]/NET0131 , \u7_mem_reg[1][16]/NET0131 , \u7_mem_reg[1][17]/NET0131 , \u7_mem_reg[1][18]/NET0131 , \u7_mem_reg[1][19]/NET0131 , \u7_mem_reg[1][1]/NET0131 , \u7_mem_reg[1][20]/NET0131 , \u7_mem_reg[1][21]/NET0131 , \u7_mem_reg[1][22]/NET0131 , \u7_mem_reg[1][23]/NET0131 , \u7_mem_reg[1][24]/NET0131 , \u7_mem_reg[1][25]/NET0131 , \u7_mem_reg[1][26]/NET0131 , \u7_mem_reg[1][27]/NET0131 , \u7_mem_reg[1][28]/NET0131 , \u7_mem_reg[1][29]/NET0131 , \u7_mem_reg[1][2]/NET0131 , \u7_mem_reg[1][30]/NET0131 , \u7_mem_reg[1][31]/NET0131 , \u7_mem_reg[1][3]/NET0131 , \u7_mem_reg[1][4]/NET0131 , \u7_mem_reg[1][5]/NET0131 , \u7_mem_reg[1][6]/NET0131 , \u7_mem_reg[1][7]/NET0131 , \u7_mem_reg[1][8]/NET0131 , \u7_mem_reg[1][9]/NET0131 , \u7_mem_reg[2][0]/NET0131 , \u7_mem_reg[2][10]/NET0131 , \u7_mem_reg[2][11]/NET0131 , \u7_mem_reg[2][12]/NET0131 , \u7_mem_reg[2][13]/NET0131 , \u7_mem_reg[2][14]/NET0131 , \u7_mem_reg[2][15]/NET0131 , \u7_mem_reg[2][16]/NET0131 , \u7_mem_reg[2][17]/NET0131 , \u7_mem_reg[2][18]/NET0131 , \u7_mem_reg[2][19]/NET0131 , \u7_mem_reg[2][1]/NET0131 , \u7_mem_reg[2][20]/NET0131 , \u7_mem_reg[2][21]/NET0131 , \u7_mem_reg[2][22]/NET0131 , \u7_mem_reg[2][23]/NET0131 , \u7_mem_reg[2][24]/NET0131 , \u7_mem_reg[2][25]/NET0131 , \u7_mem_reg[2][26]/NET0131 , \u7_mem_reg[2][27]/NET0131 , \u7_mem_reg[2][28]/NET0131 , \u7_mem_reg[2][29]/NET0131 , \u7_mem_reg[2][2]/NET0131 , \u7_mem_reg[2][30]/NET0131 , \u7_mem_reg[2][31]/NET0131 , \u7_mem_reg[2][3]/NET0131 , \u7_mem_reg[2][4]/NET0131 , \u7_mem_reg[2][5]/NET0131 , \u7_mem_reg[2][6]/NET0131 , \u7_mem_reg[2][7]/NET0131 , \u7_mem_reg[2][8]/NET0131 , \u7_mem_reg[2][9]/NET0131 , \u7_mem_reg[3][0]/NET0131 , \u7_mem_reg[3][10]/NET0131 , \u7_mem_reg[3][11]/NET0131 , \u7_mem_reg[3][12]/NET0131 , \u7_mem_reg[3][13]/NET0131 , \u7_mem_reg[3][14]/NET0131 , \u7_mem_reg[3][15]/NET0131 , \u7_mem_reg[3][16]/NET0131 , \u7_mem_reg[3][17]/NET0131 , \u7_mem_reg[3][18]/NET0131 , \u7_mem_reg[3][19]/NET0131 , \u7_mem_reg[3][1]/NET0131 , \u7_mem_reg[3][20]/NET0131 , \u7_mem_reg[3][21]/NET0131 , \u7_mem_reg[3][22]/NET0131 , \u7_mem_reg[3][23]/NET0131 , \u7_mem_reg[3][24]/NET0131 , \u7_mem_reg[3][25]/NET0131 , \u7_mem_reg[3][26]/NET0131 , \u7_mem_reg[3][27]/NET0131 , \u7_mem_reg[3][28]/NET0131 , \u7_mem_reg[3][29]/NET0131 , \u7_mem_reg[3][2]/NET0131 , \u7_mem_reg[3][30]/NET0131 , \u7_mem_reg[3][31]/NET0131 , \u7_mem_reg[3][3]/NET0131 , \u7_mem_reg[3][4]/NET0131 , \u7_mem_reg[3][5]/NET0131 , \u7_mem_reg[3][6]/NET0131 , \u7_mem_reg[3][7]/NET0131 , \u7_mem_reg[3][8]/NET0131 , \u7_mem_reg[3][9]/NET0131 , \u7_rp_reg[0]/P0001 , \u7_rp_reg[1]/NET0131 , \u7_rp_reg[2]/NET0131 , \u7_rp_reg[3]/NET0131 , \u7_status_reg[0]/P0001 , \u7_status_reg[1]/P0001 , \u7_wp_reg[0]/P0001 , \u7_wp_reg[1]/NET0131 , \u7_wp_reg[2]/P0001 , \u8_dout_reg[0]/P0001 , \u8_dout_reg[10]/P0001 , \u8_dout_reg[11]/P0001 , \u8_dout_reg[12]/P0001 , \u8_dout_reg[13]/P0001 , \u8_dout_reg[14]/P0001 , \u8_dout_reg[15]/P0001 , \u8_dout_reg[16]/P0001 , \u8_dout_reg[17]/P0001 , \u8_dout_reg[18]/P0001 , \u8_dout_reg[19]/P0001 , \u8_dout_reg[1]/P0001 , \u8_dout_reg[2]/P0001 , \u8_dout_reg[3]/P0001 , \u8_dout_reg[4]/P0001 , \u8_dout_reg[5]/P0001 , \u8_dout_reg[6]/P0001 , \u8_dout_reg[7]/P0001 , \u8_dout_reg[8]/P0001 , \u8_dout_reg[9]/P0001 , \u8_empty_reg/NET0131 , \u8_mem_reg[0][0]/NET0131 , \u8_mem_reg[0][10]/NET0131 , \u8_mem_reg[0][11]/NET0131 , \u8_mem_reg[0][12]/NET0131 , \u8_mem_reg[0][13]/NET0131 , \u8_mem_reg[0][14]/NET0131 , \u8_mem_reg[0][15]/NET0131 , \u8_mem_reg[0][16]/NET0131 , \u8_mem_reg[0][17]/NET0131 , \u8_mem_reg[0][18]/NET0131 , \u8_mem_reg[0][19]/NET0131 , \u8_mem_reg[0][1]/NET0131 , \u8_mem_reg[0][20]/NET0131 , \u8_mem_reg[0][21]/NET0131 , \u8_mem_reg[0][22]/NET0131 , \u8_mem_reg[0][23]/NET0131 , \u8_mem_reg[0][24]/NET0131 , \u8_mem_reg[0][25]/NET0131 , \u8_mem_reg[0][26]/NET0131 , \u8_mem_reg[0][27]/NET0131 , \u8_mem_reg[0][28]/NET0131 , \u8_mem_reg[0][29]/NET0131 , \u8_mem_reg[0][2]/NET0131 , \u8_mem_reg[0][30]/NET0131 , \u8_mem_reg[0][31]/NET0131 , \u8_mem_reg[0][3]/NET0131 , \u8_mem_reg[0][4]/NET0131 , \u8_mem_reg[0][5]/NET0131 , \u8_mem_reg[0][6]/NET0131 , \u8_mem_reg[0][7]/NET0131 , \u8_mem_reg[0][8]/NET0131 , \u8_mem_reg[0][9]/NET0131 , \u8_mem_reg[1][0]/NET0131 , \u8_mem_reg[1][10]/NET0131 , \u8_mem_reg[1][11]/NET0131 , \u8_mem_reg[1][12]/NET0131 , \u8_mem_reg[1][13]/NET0131 , \u8_mem_reg[1][14]/NET0131 , \u8_mem_reg[1][15]/NET0131 , \u8_mem_reg[1][16]/NET0131 , \u8_mem_reg[1][17]/NET0131 , \u8_mem_reg[1][18]/NET0131 , \u8_mem_reg[1][19]/NET0131 , \u8_mem_reg[1][1]/NET0131 , \u8_mem_reg[1][20]/NET0131 , \u8_mem_reg[1][21]/NET0131 , \u8_mem_reg[1][22]/NET0131 , \u8_mem_reg[1][23]/NET0131 , \u8_mem_reg[1][24]/NET0131 , \u8_mem_reg[1][25]/NET0131 , \u8_mem_reg[1][26]/NET0131 , \u8_mem_reg[1][27]/NET0131 , \u8_mem_reg[1][28]/NET0131 , \u8_mem_reg[1][29]/NET0131 , \u8_mem_reg[1][2]/NET0131 , \u8_mem_reg[1][30]/NET0131 , \u8_mem_reg[1][31]/NET0131 , \u8_mem_reg[1][3]/NET0131 , \u8_mem_reg[1][4]/NET0131 , \u8_mem_reg[1][5]/NET0131 , \u8_mem_reg[1][6]/NET0131 , \u8_mem_reg[1][7]/NET0131 , \u8_mem_reg[1][8]/NET0131 , \u8_mem_reg[1][9]/NET0131 , \u8_mem_reg[2][0]/NET0131 , \u8_mem_reg[2][10]/NET0131 , \u8_mem_reg[2][11]/NET0131 , \u8_mem_reg[2][12]/NET0131 , \u8_mem_reg[2][13]/NET0131 , \u8_mem_reg[2][14]/NET0131 , \u8_mem_reg[2][15]/NET0131 , \u8_mem_reg[2][16]/NET0131 , \u8_mem_reg[2][17]/NET0131 , \u8_mem_reg[2][18]/NET0131 , \u8_mem_reg[2][19]/NET0131 , \u8_mem_reg[2][1]/NET0131 , \u8_mem_reg[2][20]/NET0131 , \u8_mem_reg[2][21]/NET0131 , \u8_mem_reg[2][22]/NET0131 , \u8_mem_reg[2][23]/NET0131 , \u8_mem_reg[2][24]/NET0131 , \u8_mem_reg[2][25]/NET0131 , \u8_mem_reg[2][26]/NET0131 , \u8_mem_reg[2][27]/NET0131 , \u8_mem_reg[2][28]/NET0131 , \u8_mem_reg[2][29]/NET0131 , \u8_mem_reg[2][2]/NET0131 , \u8_mem_reg[2][30]/NET0131 , \u8_mem_reg[2][31]/NET0131 , \u8_mem_reg[2][3]/NET0131 , \u8_mem_reg[2][4]/NET0131 , \u8_mem_reg[2][5]/NET0131 , \u8_mem_reg[2][6]/NET0131 , \u8_mem_reg[2][7]/NET0131 , \u8_mem_reg[2][8]/NET0131 , \u8_mem_reg[2][9]/NET0131 , \u8_mem_reg[3][0]/NET0131 , \u8_mem_reg[3][10]/NET0131 , \u8_mem_reg[3][11]/NET0131 , \u8_mem_reg[3][12]/NET0131 , \u8_mem_reg[3][13]/NET0131 , \u8_mem_reg[3][14]/NET0131 , \u8_mem_reg[3][15]/NET0131 , \u8_mem_reg[3][16]/NET0131 , \u8_mem_reg[3][17]/NET0131 , \u8_mem_reg[3][18]/NET0131 , \u8_mem_reg[3][19]/NET0131 , \u8_mem_reg[3][1]/NET0131 , \u8_mem_reg[3][20]/NET0131 , \u8_mem_reg[3][21]/NET0131 , \u8_mem_reg[3][22]/NET0131 , \u8_mem_reg[3][23]/NET0131 , \u8_mem_reg[3][24]/NET0131 , \u8_mem_reg[3][25]/NET0131 , \u8_mem_reg[3][26]/NET0131 , \u8_mem_reg[3][27]/NET0131 , \u8_mem_reg[3][28]/NET0131 , \u8_mem_reg[3][29]/NET0131 , \u8_mem_reg[3][2]/NET0131 , \u8_mem_reg[3][30]/NET0131 , \u8_mem_reg[3][31]/NET0131 , \u8_mem_reg[3][3]/NET0131 , \u8_mem_reg[3][4]/NET0131 , \u8_mem_reg[3][5]/NET0131 , \u8_mem_reg[3][6]/NET0131 , \u8_mem_reg[3][7]/NET0131 , \u8_mem_reg[3][8]/NET0131 , \u8_mem_reg[3][9]/NET0131 , \u8_rp_reg[0]/P0001 , \u8_rp_reg[1]/NET0131 , \u8_rp_reg[2]/NET0131 , \u8_rp_reg[3]/NET0131 , \u8_status_reg[0]/P0001 , \u8_status_reg[1]/P0001 , \u8_wp_reg[0]/P0001 , \u8_wp_reg[1]/NET0131 , \u8_wp_reg[2]/P0001 , \u9_din_tmp1_reg[0]/P0001 , \u9_din_tmp1_reg[10]/P0001 , \u9_din_tmp1_reg[11]/P0001 , \u9_din_tmp1_reg[12]/P0001 , \u9_din_tmp1_reg[13]/P0001 , \u9_din_tmp1_reg[14]/P0001 , \u9_din_tmp1_reg[15]/P0001 , \u9_din_tmp1_reg[1]/P0001 , \u9_din_tmp1_reg[2]/P0001 , \u9_din_tmp1_reg[3]/P0001 , \u9_din_tmp1_reg[4]/P0001 , \u9_din_tmp1_reg[5]/P0001 , \u9_din_tmp1_reg[6]/P0001 , \u9_din_tmp1_reg[7]/P0001 , \u9_din_tmp1_reg[8]/P0001 , \u9_din_tmp1_reg[9]/P0001 , \u9_dout_reg[0]/P0001 , \u9_dout_reg[10]/P0001 , \u9_dout_reg[11]/P0001 , \u9_dout_reg[12]/P0001 , \u9_dout_reg[13]/P0001 , \u9_dout_reg[14]/P0001 , \u9_dout_reg[15]/P0001 , \u9_dout_reg[16]/P0001 , \u9_dout_reg[17]/P0001 , \u9_dout_reg[18]/P0001 , \u9_dout_reg[19]/P0001 , \u9_dout_reg[1]/P0001 , \u9_dout_reg[20]/P0001 , \u9_dout_reg[21]/P0001 , \u9_dout_reg[22]/P0001 , \u9_dout_reg[23]/P0001 , \u9_dout_reg[24]/P0001 , \u9_dout_reg[25]/P0001 , \u9_dout_reg[26]/P0001 , \u9_dout_reg[27]/P0001 , \u9_dout_reg[28]/P0001 , \u9_dout_reg[29]/P0001 , \u9_dout_reg[2]/P0001 , \u9_dout_reg[30]/P0001 , \u9_dout_reg[31]/P0001 , \u9_dout_reg[3]/P0001 , \u9_dout_reg[4]/P0001 , \u9_dout_reg[5]/P0001 , \u9_dout_reg[6]/P0001 , \u9_dout_reg[7]/P0001 , \u9_dout_reg[8]/P0001 , \u9_dout_reg[9]/P0001 , \u9_empty_reg/P0001 , \u9_full_reg/NET0131 , \u9_mem_reg[0][0]/P0001 , \u9_mem_reg[0][10]/P0001 , \u9_mem_reg[0][11]/P0001 , \u9_mem_reg[0][12]/P0001 , \u9_mem_reg[0][13]/P0001 , \u9_mem_reg[0][14]/P0001 , \u9_mem_reg[0][15]/P0001 , \u9_mem_reg[0][16]/P0001 , \u9_mem_reg[0][17]/P0001 , \u9_mem_reg[0][18]/P0001 , \u9_mem_reg[0][19]/P0001 , \u9_mem_reg[0][1]/P0001 , \u9_mem_reg[0][20]/P0001 , \u9_mem_reg[0][21]/P0001 , \u9_mem_reg[0][22]/P0001 , \u9_mem_reg[0][23]/P0001 , \u9_mem_reg[0][24]/P0001 , \u9_mem_reg[0][25]/P0001 , \u9_mem_reg[0][26]/P0001 , \u9_mem_reg[0][27]/P0001 , \u9_mem_reg[0][28]/P0001 , \u9_mem_reg[0][29]/P0001 , \u9_mem_reg[0][2]/P0001 , \u9_mem_reg[0][30]/P0001 , \u9_mem_reg[0][31]/P0001 , \u9_mem_reg[0][3]/P0001 , \u9_mem_reg[0][4]/P0001 , \u9_mem_reg[0][5]/P0001 , \u9_mem_reg[0][6]/P0001 , \u9_mem_reg[0][7]/P0001 , \u9_mem_reg[0][8]/P0001 , \u9_mem_reg[0][9]/P0001 , \u9_mem_reg[1][0]/P0001 , \u9_mem_reg[1][10]/P0001 , \u9_mem_reg[1][11]/P0001 , \u9_mem_reg[1][12]/P0001 , \u9_mem_reg[1][13]/P0001 , \u9_mem_reg[1][14]/P0001 , \u9_mem_reg[1][15]/P0001 , \u9_mem_reg[1][16]/P0001 , \u9_mem_reg[1][17]/P0001 , \u9_mem_reg[1][18]/P0001 , \u9_mem_reg[1][19]/P0001 , \u9_mem_reg[1][1]/P0001 , \u9_mem_reg[1][20]/P0001 , \u9_mem_reg[1][21]/P0001 , \u9_mem_reg[1][22]/P0001 , \u9_mem_reg[1][23]/P0001 , \u9_mem_reg[1][24]/P0001 , \u9_mem_reg[1][25]/P0001 , \u9_mem_reg[1][26]/P0001 , \u9_mem_reg[1][27]/P0001 , \u9_mem_reg[1][28]/P0001 , \u9_mem_reg[1][29]/P0001 , \u9_mem_reg[1][2]/P0001 , \u9_mem_reg[1][30]/P0001 , \u9_mem_reg[1][31]/P0001 , \u9_mem_reg[1][3]/P0001 , \u9_mem_reg[1][4]/P0001 , \u9_mem_reg[1][5]/P0001 , \u9_mem_reg[1][6]/P0001 , \u9_mem_reg[1][7]/P0001 , \u9_mem_reg[1][8]/P0001 , \u9_mem_reg[1][9]/P0001 , \u9_mem_reg[2][0]/P0001 , \u9_mem_reg[2][10]/P0001 , \u9_mem_reg[2][11]/P0001 , \u9_mem_reg[2][12]/P0001 , \u9_mem_reg[2][13]/P0001 , \u9_mem_reg[2][14]/P0001 , \u9_mem_reg[2][15]/P0001 , \u9_mem_reg[2][16]/P0001 , \u9_mem_reg[2][17]/P0001 , \u9_mem_reg[2][18]/P0001 , \u9_mem_reg[2][19]/P0001 , \u9_mem_reg[2][1]/P0001 , \u9_mem_reg[2][20]/P0001 , \u9_mem_reg[2][21]/P0001 , \u9_mem_reg[2][22]/P0001 , \u9_mem_reg[2][23]/P0001 , \u9_mem_reg[2][24]/P0001 , \u9_mem_reg[2][25]/P0001 , \u9_mem_reg[2][26]/P0001 , \u9_mem_reg[2][27]/P0001 , \u9_mem_reg[2][28]/P0001 , \u9_mem_reg[2][29]/P0001 , \u9_mem_reg[2][2]/P0001 , \u9_mem_reg[2][30]/P0001 , \u9_mem_reg[2][31]/P0001 , \u9_mem_reg[2][3]/P0001 , \u9_mem_reg[2][4]/P0001 , \u9_mem_reg[2][5]/P0001 , \u9_mem_reg[2][6]/P0001 , \u9_mem_reg[2][7]/P0001 , \u9_mem_reg[2][8]/P0001 , \u9_mem_reg[2][9]/P0001 , \u9_mem_reg[3][0]/P0001 , \u9_mem_reg[3][10]/P0001 , \u9_mem_reg[3][11]/P0001 , \u9_mem_reg[3][12]/P0001 , \u9_mem_reg[3][13]/P0001 , \u9_mem_reg[3][14]/P0001 , \u9_mem_reg[3][15]/P0001 , \u9_mem_reg[3][16]/P0001 , \u9_mem_reg[3][17]/P0001 , \u9_mem_reg[3][18]/P0001 , \u9_mem_reg[3][19]/P0001 , \u9_mem_reg[3][1]/P0001 , \u9_mem_reg[3][20]/P0001 , \u9_mem_reg[3][21]/P0001 , \u9_mem_reg[3][22]/P0001 , \u9_mem_reg[3][23]/P0001 , \u9_mem_reg[3][24]/P0001 , \u9_mem_reg[3][25]/P0001 , \u9_mem_reg[3][26]/P0001 , \u9_mem_reg[3][27]/P0001 , \u9_mem_reg[3][28]/P0001 , \u9_mem_reg[3][29]/P0001 , \u9_mem_reg[3][2]/P0001 , \u9_mem_reg[3][30]/P0001 , \u9_mem_reg[3][31]/P0001 , \u9_mem_reg[3][3]/P0001 , \u9_mem_reg[3][4]/P0001 , \u9_mem_reg[3][5]/P0001 , \u9_mem_reg[3][6]/P0001 , \u9_mem_reg[3][7]/P0001 , \u9_mem_reg[3][8]/P0001 , \u9_mem_reg[3][9]/P0001 , \u9_rp_reg[0]/P0001 , \u9_rp_reg[1]/P0001 , \u9_rp_reg[2]/P0001 , \u9_status_reg[0]/P0001 , \u9_status_reg[1]/P0001 , \u9_wp_reg[0]/NET0131 , \u9_wp_reg[1]/P0001 , \u9_wp_reg[2]/P0001 , \u9_wp_reg[3]/P0001 , \valid_s_reg/NET0131 , wb_ack_o_pad, \wb_addr_i[29]_pad , \wb_addr_i[2]_pad , \wb_addr_i[30]_pad , \wb_addr_i[31]_pad , \wb_addr_i[3]_pad , \wb_addr_i[4]_pad , \wb_addr_i[5]_pad , \wb_addr_i[6]_pad , wb_cyc_i_pad, wb_stb_i_pad, wb_we_i_pad, \_al_n1 , \g16/_0_ , \g23/_0_ , \g29500/_0_ , \g29503/_3_ , \g29505/_3_ , \g29507/_3_ , \g29509/_3_ , \g29511/_0_ , \g29513/_3_ , \g29515/_3_ , \g29517/_3_ , \g29519/_0_ , \g29522/_0_ , \g29524/_0_ , \g29526/_0_ , \g29528/_0_ , \g29530/_0_ , \g29532/_0_ , \g29534/_3_ , \g29536/_3_ , \g29538/_3_ , \g29540/_3_ , \g29542/_3_ , \g29544/_3_ , \g29546/_3_ , \g29548/_3_ , \g29550/_0_ , \g29552/_0_ , \g29554/_0_ , \g29556/_0_ , \g29558/_0_ , \g29560/_0_ , \g29562/_0_ , \g29564/_0_ , \g29566/_0_ , \g29568/_0_ , \g29570/_0_ , \g29572/_0_ , \g29574/_3_ , \g29576/_3_ , \g29578/_3_ , \g29580/_3_ , \g29582/_3_ , \g29584/_3_ , \g29586/_3_ , \g29588/_3_ , \g29590/_3_ , \g29592/_3_ , \g29594/_3_ , \g29596/_3_ , \g29598/_3_ , \g29600/_3_ , \g29602/_3_ , \g29604/_3_ , \g29606/_0_ , \g29608/_0_ , \g29610/_0_ , \g29612/_0_ , \g29614/_3_ , \g29616/_3_ , \g29618/_3_ , \g29620/_3_ , \g29622/_3_ , \g29624/_3_ , \g29626/_3_ , \g29628/_3_ , \g29630/_3_ , \g29632/_3_ , \g29634/_3_ , \g29636/_3_ , \g29638/_3_ , \g29640/_3_ , \g29642/_3_ , \g29644/_3_ , \g29646/_3_ , \g29648/_3_ , \g29650/_3_ , \g29652/_3_ , \g29654/_3_ , \g29656/_3_ , \g29658/_3_ , \g29660/_3_ , \g29662/_3_ , \g29664/_3_ , \g29666/_3_ , \g29668/_3_ , \g29670/_3_ , \g29672/_3_ , \g29674/_3_ , \g29676/_3_ , \g29678/_3_ , \g29680/_3_ , \g29682/_3_ , \g29684/_3_ , \g29686/_3_ , \g29688/_3_ , \g29690/_3_ , \g29692/_3_ , \g29694/_0_ , \g29696/_0_ , \g29698/_0_ , \g29700/_0_ , \g29702/_0_ , \g29704/_0_ , \g29706/_0_ , \g29708/_0_ , \g29710/_0_ , \g29712/_0_ , \g29714/_0_ , \g29716/_0_ , \g29718/_0_ , \g29720/_0_ , \g29722/_0_ , \g29724/_0_ , \g29726/_0_ , \g29728/_0_ , \g29730/_0_ , \g29732/_0_ , \g29734/_3_ , \g29736/_3_ , \g29738/_3_ , \g29740/_3_ , \g29742/_3_ , \g29744/_3_ , \g29746/_3_ , \g29748/_3_ , \g29750/_3_ , \g29752/_3_ , \g29754/_3_ , \g29756/_3_ , \g29758/_3_ , \g29760/_3_ , \g29762/_3_ , \g29764/_3_ , \g29766/_3_ , \g29768/_3_ , \g29770/_3_ , \g29772/_3_ , \g29774/_3_ , \g29776/_3_ , \g29778/_3_ , \g29780/_3_ , \g29782/_3_ , \g29784/_3_ , \g29786/_3_ , \g29788/_3_ , \g29790/_3_ , \g29792/_3_ , \g29794/_3_ , \g29796/_3_ , \g29798/_3_ , \g29800/_3_ , \g29802/_3_ , \g29804/_3_ , \g29806/_3_ , \g29808/_3_ , \g29810/_3_ , \g29812/_3_ , \g29814/_3_ , \g29816/_3_ , \g29818/_3_ , \g29820/_3_ , \g29822/_3_ , \g29824/_3_ , \g29826/_3_ , \g29828/_3_ , \g29830/_3_ , \g29832/_3_ , \g29834/_3_ , \g29836/_3_ , \g29838/_3_ , \g29840/_3_ , \g29842/_3_ , \g29844/_3_ , \g29846/_3_ , \g29848/_3_ , \g29850/_3_ , \g29852/_3_ , \g29854/_3_ , \g29856/_3_ , \g29858/_3_ , \g29860/_3_ , \g29862/_3_ , \g29864/_3_ , \g29866/_3_ , \g29868/_3_ , \g29870/_3_ , \g29872/_3_ , \g29874/_3_ , \g29876/_3_ , \g29878/_3_ , \g29880/_3_ , \g29904/_0_ , \g29905/_0_ , \g29906/_0_ , \g29907/_0_ , \g29908/_0_ , \g29909/_0_ , \g29914/_3_ , \g29952/_0_ , \g29953/_0_ , \g29954/_0_ , \g29955/_0_ , \g29956/_0_ , \g29957/_0_ , \g29975/_0_ , \g29976/_0_ , \g29977/_0_ , \g29978/_0_ , \g29979/_0_ , \g29980/_0_ , \g29989/_3_ , \g30020/_0_ , \g30021/_0_ , \g30045/_0_ , \g30046/_0_ , \g30047/_0_ , \g30048/_0_ , \g30049/_0_ , \g30050/_0_ , \g30051/_0_ , \g30052/_0_ , \g30053/_0_ , \g30054/_0_ , \g30062/_0_ , \g30063/_0_ , \g30064/_0_ , \g30065/_0_ , \g30066/_0_ , \g30067/_0_ , \g30068/_0_ , \g30069/_0_ , \g30070/_0_ , \g30071/_0_ , \g30072/_0_ , \g30073/_0_ , \g30074/_0_ , \g30075/_0_ , \g30136/_3_ , \g30707/_0_ , \g30708/_0_ , \g30711/_0_ , \g30714/_0_ , \g30715/_0_ , \g30720/_0_ , \g30725/_0_ , \g30741/_0_ , \g30742/_0_ , \g30743/_0_ , \g30744/_0_ , \g30745/_0_ , \g30746/_0_ , \g30747/_0_ , \g30748/_0_ , \g30749/_0_ , \g30750/_0_ , \g30751/_0_ , \g30752/_0_ , \g30789/_0_ , \g30790/_0_ , \g30791/_0_ , \g30792/_0_ , \g30793/_0_ , \g30794/_0_ , \g30795/_0_ , \g30796/_0_ , \g30797/_0_ , \g30798/_0_ , \g30799/_0_ , \g30800/_0_ , \g30801/_0_ , \g30802/_0_ , \g30803/_0_ , \g30804/_0_ , \g30805/_0_ , \g30806/_0_ , \g30807/_0_ , \g30808/_0_ , \g30809/_0_ , \g30810/_0_ , \g30811/_0_ , \g30812/_0_ , \g30813/_0_ , \g30814/_0_ , \g30815/_0_ , \g30816/_0_ , \g30817/_0_ , \g30818/_0_ , \g30819/_0_ , \g30820/_0_ , \g30821/_0_ , \g30822/_0_ , \g30823/_0_ , \g30824/_0_ , \g30825/_0_ , \g30826/_0_ , \g30827/_0_ , \g30828/_0_ , \g30829/_0_ , \g30830/_0_ , \g30831/_0_ , \g30832/_0_ , \g30833/_0_ , \g30834/_0_ , \g30835/_0_ , \g30836/_0_ , \g30837/_0_ , \g30838/_0_ , \g30839/_0_ , \g30840/_0_ , \g30841/_0_ , \g30842/_0_ , \g30843/_0_ , \g30844/_0_ , \g30845/_0_ , \g30846/_0_ , \g30847/_0_ , \g30848/_0_ , \g30849/_0_ , \g30850/_0_ , \g30851/_0_ , \g30852/_0_ , \g30853/_0_ , \g30854/_0_ , \g30855/_0_ , \g30856/_0_ , \g30857/_0_ , \g30858/_0_ , \g30859/_0_ , \g30860/_0_ , \g30861/_0_ , \g30862/_0_ , \g30863/_0_ , \g30864/_0_ , \g30865/_0_ , \g30866/_0_ , \g30867/_0_ , \g30868/_0_ , \g30869/_0_ , \g30870/_0_ , \g30871/_0_ , \g30872/_0_ , \g30873/_0_ , \g30874/_0_ , \g30875/_0_ , \g30876/_0_ , \g30877/_0_ , \g30878/_0_ , \g30879/_0_ , \g30880/_0_ , \g30881/_0_ , \g30882/_0_ , \g30883/_0_ , \g30884/_0_ , \g30885/_0_ , \g30886/_0_ , \g30887/_0_ , \g30888/_0_ , \g30889/_0_ , \g30890/_0_ , \g30891/_0_ , \g30892/_0_ , \g30893/_0_ , \g30894/_0_ , \g30895/_0_ , \g30896/_0_ , \g30897/_0_ , \g30898/_0_ , \g30899/_0_ , \g30900/_0_ , \g30901/_0_ , \g30902/_0_ , \g30906/_0_ , \g30907/_0_ , \g30908/_0_ , \g30909/_0_ , \g30910/_0_ , \g30911/_0_ , \g30918/_0_ , \g30919/_0_ , \g30920/_0_ , \g30921/_0_ , \g30922/_0_ , \g30923/_0_ , \g30924/_0_ , \g30925/_0_ , \g30926/_0_ , \g30946/_0_ , \g30947/_0_ , \g30948/_0_ , \g30949/_0_ , \g30950/_0_ , \g30951/_0_ , \g30952/_0_ , \g30953/_0_ , \g30954/_0_ , \g30955/_0_ , \g30956/_0_ , \g30957/_0_ , \g30958/_0_ , \g30959/_0_ , \g30960/_0_ , \g30961/_0_ , \g30962/_0_ , \g30963/_0_ , \g30964/_0_ , \g30965/_0_ , \g30966/_0_ , \g30967/_0_ , \g30968/_0_ , \g30969/_0_ , \g30970/_0_ , \g30971/_0_ , \g30972/_0_ , \g30973/_0_ , \g30974/_0_ , \g30975/_0_ , \g30976/_0_ , \g30977/_0_ , \g30978/_0_ , \g30979/_0_ , \g30980/_0_ , \g30981/_0_ , \g30982/_0_ , \g30983/_0_ , \g30984/_0_ , \g30985/_0_ , \g30986/_0_ , \g30987/_0_ , \g30988/_0_ , \g30989/_0_ , \g30990/_0_ , \g30991/_0_ , \g30992/_0_ , \g30993/_0_ , \g30994/_0_ , \g30995/_0_ , \g30996/_0_ , \g30997/_0_ , \g30998/_0_ , \g30999/_0_ , \g31000/_0_ , \g31001/_0_ , \g31002/_0_ , \g31003/_0_ , \g31004/_0_ , \g31005/_0_ , \g31006/_0_ , \g31007/_0_ , \g31008/_0_ , \g31009/_0_ , \g31010/_0_ , \g31011/_0_ , \g31012/_0_ , \g31013/_0_ , \g31014/_0_ , \g31015/_0_ , \g31016/_0_ , \g31017/_0_ , \g31018/_0_ , \g31019/_0_ , \g31020/_0_ , \g31021/_0_ , \g31022/_0_ , \g31023/_0_ , \g31024/_0_ , \g31025/_0_ , \g31026/_0_ , \g31027/_0_ , \g31028/_0_ , \g31029/_0_ , \g31030/_0_ , \g31031/_0_ , \g31032/_0_ , \g31033/_0_ , \g31034/_0_ , \g31035/_0_ , \g31036/_0_ , \g31037/_0_ , \g31038/_0_ , \g31039/_0_ , \g31040/_0_ , \g31041/_0_ , \g31042/_0_ , \g31043/_0_ , \g31044/_0_ , \g31045/_0_ , \g31046/_0_ , \g31047/_0_ , \g31048/_0_ , \g31049/_0_ , \g31050/_0_ , \g31051/_0_ , \g31052/_0_ , \g31053/_0_ , \g31054/_0_ , \g31055/_0_ , \g31056/_0_ , \g31057/_0_ , \g31058/_0_ , \g31059/_0_ , \g31060/_0_ , \g31061/_0_ , \g31062/_0_ , \g31063/_0_ , \g31064/_0_ , \g31065/_0_ , \g31066/_0_ , \g31067/_0_ , \g31068/_0_ , \g31069/_0_ , \g31070/_0_ , \g31071/_0_ , \g31072/_0_ , \g31073/_0_ , \g31074/_0_ , \g31075/_0_ , \g31076/_0_ , \g31077/_0_ , \g31084/u3_syn_4 , \g31085/u3_syn_4 , \g31096/u3_syn_4 , \g31115/u3_syn_4 , \g31136/u3_syn_4 , \g31158/u3_syn_4 , \g31176/u3_syn_4 , \g31193/u3_syn_4 , \g31195/u3_syn_4 , \g31247/u3_syn_4 , \g31280/u3_syn_4 , \g31285/u3_syn_4 , \g31568/_0_ , \g31631/_0_ , \g31672/_0_ , \g31731/_0_ , \g31732/_0_ , \g31742/_2_ , \g31744/_2_ , \g31746/_2_ , \g31748/_2_ , \g31751/_2_ , \g31754/_2_ , \g31756/_2_ , \g31758/_2_ , \g31760/_2_ , \g31761/_0_ , \g31789/_0_ , \g31807/_3_ , \g31825/_3_ , \g32607/_0_ , \g32608/_0_ , \g32609/_0_ , \g32610/_0_ , \g32611/_0_ , \g32612/_0_ , \g32613/_0_ , \g32614/_0_ , \g32615/_0_ , \g32616/_0_ , \g32617/_0_ , \g32618/_0_ , \g32645/_0__syn_2 , \g32687/_0__syn_2 , \g32749/_0__syn_2 , \g32757/_0_ , \g32758/_0_ , \g32759/_0_ , \g32760/_0_ , \g32761/_0_ , \g32762/_0_ , \g32763/_0_ , \g32764/_0_ , \g32765/_0_ , \g32769/_0_ , \g32835/_1_ , \g32839/_0_ , \g32844/_0_ , \g32901/_1_ , \g32902/_0_ , \g32963/_1_ , \g32972/_0_ , \g32977/_0_ , \g32979/_0_ , \g32980/_0_ , \g32981/_0_ , \g32982/_0_ , \g32983/_0_ , \g32987/_0_ , \g33018/_0_ , \g33019/_0_ , \g33088/_0_ , \g33261/_0_ , \g33264/_0_ , \g33275/_0_ , \g33276/_0_ , \g33277/_0_ , \g33371/_0_ , \g33382/_0_ , \g33401/_0_ , \g33402/_0_ , \g33403/_0_ , \g33404/_0_ , \g33405/_0_ , \g33406/_0_ , \g33407/_0_ , \g33408/_0_ , \g33409/_0_ , \g33410/_0_ , \g33411/_0_ , \g33412/_0_ , \g33413/_0_ , \g33414/_0_ , \g33415/_0_ , \g33416/_0_ , \g33417/_0_ , \g33418/_0_ , \g33419/_0_ , \g33420/_0_ , \g33421/_0_ , \g33422/_0_ , \g33423/_0_ , \g33424/_0_ , \g33425/_0_ , \g33426/_0_ , \g33427/_0_ , \g33428/_0_ , \g33429/_0_ , \g33430/_0_ , \g33431/_0_ , \g33432/_0_ , \g33433/_0_ , \g33434/_0_ , \g33435/_0_ , \g33436/_0_ , \g33437/_0_ , \g33438/_0_ , \g33439/_0_ , \g33440/_0_ , \g33441/_0_ , \g33442/_0_ , \g33443/_0_ , \g33444/_0_ , \g33445/_0_ , \g33446/_0_ , \g33447/_0_ , \g33448/_0_ , \g33449/_0_ , \g33450/_0_ , \g33451/_0_ , \g33452/_0_ , \g33453/_0_ , \g33454/_0_ , \g33455/_0_ , \g33456/_0_ , \g33457/_0_ , \g33458/_0_ , \g33459/_0_ , \g33460/_0_ , \g33461/_0_ , \g33462/_0_ , \g33463/_0_ , \g33464/_0_ , \g33465/_0_ , \g33466/_0_ , \g33467/_0_ , \g33468/_0_ , \g33469/_0_ , \g33470/_0_ , \g33471/_0_ , \g33472/_0_ , \g33473/_0_ , \g33474/_0_ , \g33475/_0_ , \g33476/_0_ , \g33477/_0_ , \g33478/_0_ , \g33479/_0_ , \g33480/_0_ , \g33481/_0_ , \g33482/_0_ , \g33483/_0_ , \g33484/_0_ , \g33485/_0_ , \g33486/_0_ , \g33487/_0_ , \g33488/_0_ , \g33489/_0_ , \g33490/_0_ , \g33491/_0_ , \g33492/_0_ , \g33493/_0_ , \g33494/_0_ , \g33495/_0_ , \g33496/_0_ , \g33497/_0_ , \g33498/_0_ , \g33499/_0_ , \g33500/_0_ , \g33501/_0_ , \g33502/_0_ , \g33503/_0_ , \g33504/_0_ , \g33505/_0_ , \g33506/_0_ , \g33507/_0_ , \g33508/_0_ , \g33509/_0_ , \g33510/_0_ , \g33511/_0_ , \g33512/_0_ , \g33513/_0_ , \g33514/_0_ , \g33515/_0_ , \g33516/_0_ , \g33517/_0_ , \g33518/_0_ , \g33519/_0_ , \g33520/_0_ , \g33521/_0_ , \g33522/_0_ , \g33523/_0_ , \g33524/_0_ , \g33525/_0_ , \g33526/_0_ , \g33527/_0_ , \g33528/_0_ , \g33529/_0_ , \g33530/_0_ , \g33531/_0_ , \g33532/_0_ , \g33533/_0_ , \g33534/_0_ , \g33535/_0_ , \g33536/_0_ , \g33537/_0_ , \g33538/_0_ , \g33539/_0_ , \g33540/_0_ , \g33541/_0_ , \g33542/_0_ , \g33543/_0_ , \g33544/_0_ , \g33545/_0_ , \g33546/_0_ , \g33547/_0_ , \g33548/_0_ , \g33549/_0_ , \g33550/_0_ , \g33551/_0_ , \g33552/_0_ , \g33553/_0_ , \g33554/_0_ , \g33555/_0_ , \g33556/_0_ , \g33557/_0_ , \g33558/_0_ , \g33559/_0_ , \g33560/_0_ , \g33561/_0_ , \g33562/_0_ , \g33563/_0_ , \g33564/_0_ , \g33565/_0_ , \g33566/_0_ , \g33567/_0_ , \g33568/_0_ , \g33569/_0_ , \g33570/_0_ , \g33571/_0_ , \g33572/_0_ , \g33573/_0_ , \g33574/_0_ , \g33575/_0_ , \g33576/_0_ , \g33577/_0_ , \g33578/_0_ , \g33579/_0_ , \g33580/_0_ , \g33581/_0_ , \g33582/_0_ , \g33583/_0_ , \g33584/_0_ , \g33585/_0_ , \g33586/_0_ , \g33587/_0_ , \g33588/_0_ , \g33589/_0_ , \g33590/_0_ , \g33591/_0_ , \g33592/_0_ , \g33593/_0_ , \g33594/_0_ , \g33595/_0_ , \g33596/_0_ , \g33597/_0_ , \g33598/_0_ , \g33599/_0_ , \g33600/_0_ , \g33601/_0_ , \g33602/_0_ , \g33603/_0_ , \g33604/_0_ , \g33605/_0_ , \g33606/_0_ , \g33607/_0_ , \g33608/_0_ , \g33609/_0_ , \g33610/_0_ , \g33611/_0_ , \g33612/_0_ , \g33613/_0_ , \g33614/_0_ , \g33615/_0_ , \g33616/_0_ , \g33617/_0_ , \g33618/_0_ , \g33619/_0_ , \g33620/_0_ , \g33621/_0_ , \g33622/_0_ , \g33623/_0_ , \g33624/_0_ , \g33625/_0_ , \g33626/_0_ , \g33627/_0_ , \g33628/_0_ , \g33629/_0_ , \g33630/_0_ , \g33631/_0_ , \g33632/_0_ , \g33633/_0_ , \g33634/_0_ , \g33635/_0_ , \g33636/_0_ , \g33637/_0_ , \g33638/_0_ , \g33639/_0_ , \g33640/_0_ , \g33641/_0_ , \g33642/_0_ , \g33643/_0_ , \g33644/_0_ , \g33645/_0_ , \g33646/_0_ , \g33647/_0_ , \g33648/_0_ , \g33649/_0_ , \g33650/_0_ , \g33651/_0_ , \g33652/_0_ , \g33653/_0_ , \g33654/_0_ , \g33655/_0_ , \g33656/_0_ , \g33657/_0_ , \g33658/_0_ , \g33659/_0_ , \g33660/_0_ , \g33661/_0_ , \g33662/_0_ , \g33663/_0_ , \g33664/_0_ , \g33665/_0_ , \g33666/_0_ , \g33667/_0_ , \g33668/_0_ , \g33669/_0_ , \g33670/_0_ , \g33671/_0_ , \g33672/_0_ , \g33673/_0_ , \g33674/_0_ , \g33675/_0_ , \g33676/_0_ , \g33677/_0_ , \g33678/_0_ , \g33679/_0_ , \g33680/_0_ , \g33681/_0_ , \g33682/_0_ , \g33683/_0_ , \g33684/_0_ , \g33685/_0_ , \g33686/_0_ , \g33687/_0_ , \g33688/_0_ , \g33689/_0_ , \g33690/_0_ , \g33691/_0_ , \g33692/_0_ , \g33693/_0_ , \g33694/_0_ , \g33695/_0_ , \g33696/_0_ , \g33697/_0_ , \g33698/_0_ , \g33699/_0_ , \g33700/_0_ , \g33701/_0_ , \g33702/_0_ , \g33703/_0_ , \g33704/_0_ , \g33705/_0_ , \g33706/_0_ , \g33707/_0_ , \g33708/_0_ , \g33709/_0_ , \g33710/_0_ , \g33711/_0_ , \g33712/_0_ , \g33713/_0_ , \g33714/_0_ , \g33715/_0_ , \g33716/_0_ , \g33717/_0_ , \g33718/_0_ , \g33719/_0_ , \g33720/_0_ , \g33721/_0_ , \g33722/_0_ , \g33723/_0_ , \g33724/_0_ , \g33725/_0_ , \g33726/_0_ , \g33727/_0_ , \g33728/_0_ , \g33729/_0_ , \g33730/_0_ , \g33731/_0_ , \g33732/_0_ , \g33733/_0_ , \g33734/_0_ , \g33735/_0_ , \g33736/_0_ , \g33737/_0_ , \g33738/_0_ , \g33739/_0_ , \g33740/_0_ , \g33741/_0_ , \g33742/_0_ , \g33743/_0_ , \g33744/_0_ , \g33745/_0_ , \g33746/_0_ , \g33747/_0_ , \g33748/_0_ , \g33749/_0_ , \g33750/_0_ , \g33751/_0_ , \g33752/_0_ , \g33753/_0_ , \g33754/_0_ , \g33755/_0_ , \g33756/_0_ , \g33757/_0_ , \g33758/_0_ , \g33759/_0_ , \g33760/_0_ , \g33761/_0_ , \g33762/_0_ , \g33763/_0_ , \g33764/_0_ , \g33765/_0_ , \g33766/_0_ , \g33767/_0_ , \g33768/_0_ , \g33769/_0_ , \g33770/_0_ , \g33771/_0_ , \g33772/_0_ , \g33773/_0_ , \g33774/_0_ , \g33775/_0_ , \g33776/_0_ , \g33777/_0_ , \g33778/_0_ , \g33779/_0_ , \g33780/_0_ , \g33781/_0_ , \g33782/_0_ , \g33783/_0_ , \g33784/_0_ , \g33785/_0_ , \g33786/_0_ , \g33787/_0_ , \g33788/_0_ , \g33789/_0_ , \g33790/_0_ , \g33791/_0_ , \g33792/_0_ , \g33793/_0_ , \g33794/_0_ , \g33795/_0_ , \g33796/_0_ , \g33797/_0_ , \g33798/_0_ , \g33799/_0_ , \g33800/_0_ , \g33801/_0_ , \g33802/_0_ , \g33803/_0_ , \g33804/_0_ , \g33805/_0_ , \g33806/_0_ , \g33807/_0_ , \g33808/_0_ , \g33809/_0_ , \g33810/_0_ , \g33811/_0_ , \g33812/_0_ , \g33813/_0_ , \g33814/_0_ , \g33815/_0_ , \g33816/_0_ , \g33817/_0_ , \g33818/_0_ , \g33819/_0_ , \g33820/_0_ , \g33821/_0_ , \g33822/_0_ , \g33823/_0_ , \g33824/_0_ , \g33825/_0_ , \g33826/_0_ , \g33827/_0_ , \g33828/_0_ , \g33829/_0_ , \g33830/_0_ , \g33831/_0_ , \g33832/_0_ , \g33833/_0_ , \g33834/_0_ , \g33835/_0_ , \g33836/_0_ , \g33837/_0_ , \g33838/_0_ , \g33839/_0_ , \g33840/_0_ , \g33841/_0_ , \g33842/_0_ , \g33843/_0_ , \g33844/_0_ , \g33845/_0_ , \g33846/_0_ , \g33847/_0_ , \g33848/_0_ , \g33849/_0_ , \g33850/_0_ , \g33851/_0_ , \g33852/_0_ , \g33853/_0_ , \g33854/_0_ , \g33855/_0_ , \g33856/_0_ , \g33857/_0_ , \g33858/_0_ , \g33859/_0_ , \g33860/_0_ , \g33861/_0_ , \g33862/_0_ , \g33863/_0_ , \g33864/_0_ , \g33865/_0_ , \g33866/_0_ , \g33867/_0_ , \g33868/_0_ , \g33869/_0_ , \g33870/_0_ , \g33871/_0_ , \g33872/_0_ , \g33873/_0_ , \g33874/_0_ , \g33875/_0_ , \g33876/_0_ , \g33877/_0_ , \g33878/_0_ , \g33879/_0_ , \g33880/_0_ , \g33881/_0_ , \g33882/_0_ , \g33883/_0_ , \g33884/_0_ , \g33885/_0_ , \g33886/_0_ , \g33887/_0_ , \g33888/_0_ , \g33889/_0_ , \g33890/_0_ , \g33891/_0_ , \g33892/_0_ , \g33893/_0_ , \g33894/_0_ , \g33895/_0_ , \g33896/_0_ , \g33897/_0_ , \g33898/_0_ , \g33899/_0_ , \g33900/_0_ , \g33901/_0_ , \g33902/_0_ , \g33903/_0_ , \g33904/_0_ , \g33905/_0_ , \g33906/_0_ , \g33907/_0_ , \g33908/_0_ , \g33909/_0_ , \g33910/_0_ , \g33911/_0_ , \g33912/_0_ , \g33913/_0_ , \g33914/_0_ , \g33915/_0_ , \g33916/_0_ , \g33917/_0_ , \g33918/_0_ , \g33919/_0_ , \g33920/_0_ , \g33921/_0_ , \g33922/_0_ , \g33923/_0_ , \g33924/_0_ , \g33925/_0_ , \g33926/_0_ , \g33927/_0_ , \g33928/_0_ , \g33929/_0_ , \g33930/_0_ , \g33931/_0_ , \g33932/_0_ , \g33933/_0_ , \g33934/_0_ , \g33935/_0_ , \g33936/_0_ , \g33937/_0_ , \g33938/_0_ , \g33939/_0_ , \g33940/_0_ , \g33941/_0_ , \g33942/_0_ , \g33943/_0_ , \g33944/_0_ , \g33945/_0_ , \g33946/_0_ , \g33947/_0_ , \g33948/_0_ , \g33949/_0_ , \g33950/_0_ , \g33951/_0_ , \g33952/_0_ , \g33953/_0_ , \g33954/_0_ , \g33955/_0_ , \g33956/_0_ , \g33957/_0_ , \g33958/_0_ , \g33959/_0_ , \g33960/_0_ , \g33961/_0_ , \g33962/_0_ , \g33963/_0_ , \g33964/_0_ , \g33965/_0_ , \g33966/_0_ , \g33967/_0_ , \g33968/_0_ , \g33969/_0_ , \g33970/_0_ , \g33971/_0_ , \g33972/_0_ , \g33973/_0_ , \g33974/_0_ , \g33975/_0_ , \g33976/_0_ , \g33977/u3_syn_4 , \g33981/u3_syn_4 , \g34014/u3_syn_4 , \g34047/u3_syn_4 , \g34084/u3_syn_4 , \g34123/u3_syn_4 , \g34306/_0_ , \g34316/_0_ , \g34324/_0_ , \g34326/_0_ , \g34328/_0_ , \g34331/_0_ , \g34333/_0_ , \g34344/_0_ , \g34347/_0_ , \g34351/_0_ , \g34361/_0_ , \g34368/_0_ , \g34377/_0_ , \g34385/_0_ , \g34393/_0_ , \g34414/_1_ , \g34451/_1_ , \g34476/_1_ , \g34487/_0_ , \g34490/_1_ , \g34715/_0_ , \g34878/_0_ , \g34882/_0_ , \g34883/_0_ , \g34893/_0_ , \g34896/_0_ , \g34898/_0_ , \g34899/_0_ , \g34916/_3_ , \g35264/_0_ , \g35265/_0_ , \g35266/_0_ , \g35267/_0_ , \g35268/_0_ , \g35269/_0_ , \g35270/_0_ , \g35271/_0_ , \g35272/_0_ , \g35273/_0_ , \g35274/_0_ , \g35275/_0_ , \g35276/_0_ , \g35277/_0_ , \g35278/_0_ , \g35279/_0_ , \g35283/_0_ , \g35287/_0_ , \g35294/_0_ , \g35300/_0_ , \g35304/_0_ , \g35308/_0_ , \g35312/_0_ , \g35316/_0_ , \g35318/_0_ , \g35326/_0_ , \g35334/_0_ , \g35336/_0_ , \g35337/_0_ , \g35338/_0_ , \g35357/_0_ , \g35358/_0_ , \g35359/_0_ , \g35419/_0_ , \g35438/_0_ , \g35439/_0_ , \g35440/_0_ , \g35441/_0_ , \g35442/_0_ , \g35444/_0_ , \g35445/_0_ , \g35446/_0_ , \g35447/_0_ , \g35448/_0_ , \g35449/_0_ , \g35450/_0_ , \g35451/_0_ , \g35452/_0_ , \g35463/_0_ , \g35464/_0_ , \g35466/_0_ , \g35485/_2_ , \g35495/_0_ , \g35496/_0_ , \g35499/_0_ , \g35500/_0_ , \g35501/_0_ , \g35502/_0_ , \g35563/_0_ , \g35633/_0_ , \g35717/_0_ , \g35718/_0_ , \g35719/_0_ , \g35809/_0_ , \g35810/_0_ , \g35811/_0_ , \g35812/_0_ , \g35813/_0_ , \g35814/_0_ , \g35815/_0_ , \g35816/_0_ , \g35817/_0_ , \g35818/_0_ , \g35819/_0_ , \g35820/_0_ , \g35821/_0_ , \g35822/_0_ , \g35823/_0_ , \g35824/_0_ , \g35825/_0_ , \g35826/_0_ , \g35827/_0_ , \g35830/_0_ , \g35833/_0_ , \g35835/_0_ , \g35836/_0_ , \g35837/_0_ , \g35839/_0_ , \g35840/_0_ , \g35841/_0_ , \g35843/_0_ , \g35844/_0_ , \g35845/_0_ , \g35853/_0_ , \g35854/_0_ , \g35855/_0_ , \g35856/_0_ , \g36306/_0_ , \g36414/_0_ , \g36415/_0_ , \g36449/_0_ , \g36550/_0_ , \g36551/_0_ , \g36553/_0_ , \g36560/_0_ , \g36562/_3_ , \g36563/_0_ , \g36612/_0_ , \g36614/_2_ , \g36695/_0_ , \g36784/_0_ , \g36785/_0_ , \g36786/_0_ , \g36787/_0_ , \g36788/_0_ , \g36789/_0_ , \g36790/_0_ , \g36791/_0_ , \g36792/_0_ , \g36793/_0_ , \g36794/_0_ , \g36796/_0_ , \g36797/_0_ , \g36798/_0_ , \g36799/_0_ , \g36800/_0_ , \g36801/_0_ , \g36802/_0_ , \g36803/_0_ , \g36804/_0_ , \g36805/_0_ , \g36806/_0_ , \g36807/_0_ , \g36808/_0_ , \g36809/_0_ , \g36810/_0_ , \g36811/_0_ , \g36813/_0_ , \g36814/_0_ , \g36815/_0_ , \g36820/_0_ , \g36825/_0_ , \g36832/_0_ , \g36846/_0_ , \g36855/_0_ , \g36857/_0_ , \g36859/_0_ , \g36860/_0_ , \g36861/_0_ , \g36862/_0_ , \g36863/_0_ , \g36864/_0_ , \g36867/_0_ , \g36870/_0_ , \g36871/_0_ , \g36877/_0_ , \g36879/_0_ , \g36892/_0_ , \g36893/_0_ , \g36901/_0_ , \g36909/_0_ , \g36914/_0_ , \g36919/_0_ , \g36922/_0_ , \g36923/_0_ , \g36927/_0_ , \g36930/_0_ , \g36931/_0_ , \g36933/_0_ , \g36934/_0_ , \g36935/_0_ , \g36936/_0_ , \g36937/_0_ , \g36938/_0_ , \g36939/_0_ , \g36940/_0_ , \g36941/_0_ , \g36943/_0_ , \g36944/_0_ , \g36945/_0_ , \g36946/_0_ , \g36947/_0_ , \g36948/_0_ , \g36949/_0_ , \g36950/_0_ , \g36951/_0_ , \g36952/_0_ , \g36953/_0_ , \g36954/_0_ , \g36957/_0_ , \g36958/_0_ , \g36959/_0_ , \g36960/_0_ , \g36961/_0_ , \g36962/_0_ , \g36963/_0_ , \g36970/_0_ , \g36977/_0_ , \g36986/_0_ , \g36991/_0_ , \g36994/_0_ , \g37015/_0_ , \g37057/_0_ , \g37073/_0_ , \g37128/_0_ , \g37129/_0_ , \g37138/_0_ , \g37139/_0_ , \g37140/_0_ , \g37141/_0_ , \g37142/_0_ , \g37143/_0_ , \g37144/_0_ , \g37145/_0_ , \g37146/_0_ , \g37147/_0_ , \g37148/_0_ , \g37149/_0_ , \g37150/_0_ , \g37151/_0_ , \g37152/_0_ , \g37153/_0_ , \g37154/_0_ , \g37155/_0_ , \g37156/_0_ , \g37157/_0_ , \g37158/_0_ , \g37159/_0_ , \g37160/_0_ , \g37161/_0_ , \g37162/_0_ , \g37163/_0_ , \g37164/_0_ , \g37165/_0_ , \g37166/_0_ , \g37167/_0_ , \g37168/_0_ , \g37169/_0_ , \g37170/_0_ , \g37171/_0_ , \g37172/_0_ , \g37173/_0_ , \g37174/_0_ , \g37175/_0_ , \g37176/_0_ , \g37177/_0_ , \g37178/_0_ , \g37179/_0_ , \g37180/_0_ , \g37181/_0_ , \g37182/_0_ , \g37183/_0_ , \g37184/_0_ , \g37185/_0_ , \g37187/_0_ , \g37188/_0_ , \g37190/_0_ , \g37191/_0_ , \g37192/_0_ , \g37193/_0_ , \g37194/_0_ , \g37372/_3_ , \g37377/_0_ , \g37378/_0_ , \g37379/_0_ , \g37380/_0_ , \g37381/_0_ , \g37382/_0_ , \g37383/_0_ , \g37384/_0_ , \g37385/_0_ , \g37386/_0_ , \g37387/_0_ , \g37388/_0_ , \g37389/_0_ , \g37390/_0_ , \g37391/_0_ , \g37392/_0_ , \g37393/_0_ , \g37394/_0_ , \g37395/_0_ , \g37396/_0_ , \g37397/_0_ , \g37398/_0_ , \g37399/_0_ , \g37400/_0_ , \g37401/_0_ , \g37402/_0_ , \g37403/_0_ , \g37404/_0_ , \g37405/_0_ , \g37406/_0_ , \g37407/_0_ , \g37408/_0_ , \g37409/_0_ , \g37410/_0_ , \g37411/_0_ , \g37412/_0_ , \g37413/_0_ , \g37576/_3_ , \g37590/_2_ , \g40278/_0_ , \g40379/_0_ , \g40389/_2_ , \g40390/_2_ , \g40391/_0_ , \g40393/_2_ , \g40395/_0_ , \g40397/_0_ , \g40400/_0_ , \g40402/_0_ , \g45458/_0_ , \g45675/_0_ , \g45677/_0_ , \g45678/_0_ , \g45682/_0_ , sync_pad_o_pad, \u14_u0_full_empty_r_reg/P0001_reg_syn_3 , \u14_u1_full_empty_r_reg/P0001_reg_syn_3 , \u14_u2_full_empty_r_reg/P0001_reg_syn_3 , \u14_u3_full_empty_r_reg/P0001_reg_syn_3 , \u14_u4_full_empty_r_reg/P0001_reg_syn_3 , \u14_u5_full_empty_r_reg/P0001_reg_syn_3 , \u14_u6_full_empty_r_reg/P0001_reg_syn_3 , \u14_u7_full_empty_r_reg/P0001_reg_syn_3 , \u14_u8_full_empty_r_reg/P0001_reg_syn_3 , \u1_slt0_reg[11]/P0001_reg_syn_3 , \u1_slt0_reg[12]/P0001_reg_syn_3 , \u1_slt0_reg[15]/P0001_reg_syn_3 , \u1_slt0_reg[9]/P0001_reg_syn_3 , \u1_slt1_reg[10]/P0001_reg_syn_3 , \u1_slt1_reg[11]/P0001_reg_syn_3 , \u1_slt1_reg[5]/P0001_reg_syn_3 , \u1_slt1_reg[6]/P0001_reg_syn_3 , \u1_slt1_reg[7]/P0001_reg_syn_3 , \u1_slt1_reg[8]/P0001_reg_syn_3 , wb_err_o_pad);
	input \ac97_reset_pad_o__pad  ;
	input \dma_ack_i[0]_pad  ;
	input \dma_ack_i[1]_pad  ;
	input \dma_ack_i[2]_pad  ;
	input \dma_ack_i[3]_pad  ;
	input \dma_ack_i[4]_pad  ;
	input \dma_ack_i[5]_pad  ;
	input \dma_ack_i[6]_pad  ;
	input \dma_ack_i[7]_pad  ;
	input \dma_ack_i[8]_pad  ;
	input \dma_req_o[0]_pad  ;
	input \dma_req_o[1]_pad  ;
	input \dma_req_o[2]_pad  ;
	input \dma_req_o[3]_pad  ;
	input \dma_req_o[4]_pad  ;
	input \dma_req_o[5]_pad  ;
	input \dma_req_o[6]_pad  ;
	input \dma_req_o[7]_pad  ;
	input \dma_req_o[8]_pad  ;
	input \in_valid_s_reg[0]/NET0131  ;
	input \in_valid_s_reg[1]/NET0131  ;
	input \in_valid_s_reg[2]/NET0131  ;
	input suspended_o_pad ;
	input \u0_slt0_r_reg[0]/P0001  ;
	input \u0_slt0_r_reg[10]/P0001  ;
	input \u0_slt0_r_reg[11]/P0001  ;
	input \u0_slt0_r_reg[12]/P0001  ;
	input \u0_slt0_r_reg[13]/P0001  ;
	input \u0_slt0_r_reg[14]/P0001  ;
	input \u0_slt0_r_reg[1]/P0001  ;
	input \u0_slt0_r_reg[2]/P0001  ;
	input \u0_slt0_r_reg[3]/P0001  ;
	input \u0_slt0_r_reg[4]/P0001  ;
	input \u0_slt0_r_reg[5]/P0001  ;
	input \u0_slt0_r_reg[6]/P0001  ;
	input \u0_slt0_r_reg[7]/P0001  ;
	input \u0_slt0_r_reg[8]/P0001  ;
	input \u0_slt0_r_reg[9]/P0001  ;
	input \u0_slt1_r_reg[0]/P0001  ;
	input \u0_slt1_r_reg[10]/P0001  ;
	input \u0_slt1_r_reg[11]/P0001  ;
	input \u0_slt1_r_reg[12]/P0001  ;
	input \u0_slt1_r_reg[13]/P0001  ;
	input \u0_slt1_r_reg[14]/P0001  ;
	input \u0_slt1_r_reg[15]/P0001  ;
	input \u0_slt1_r_reg[16]/P0001  ;
	input \u0_slt1_r_reg[17]/P0001  ;
	input \u0_slt1_r_reg[18]/P0001  ;
	input \u0_slt1_r_reg[19]/P0001  ;
	input \u0_slt1_r_reg[1]/P0001  ;
	input \u0_slt1_r_reg[2]/P0001  ;
	input \u0_slt1_r_reg[3]/P0001  ;
	input \u0_slt1_r_reg[4]/P0001  ;
	input \u0_slt1_r_reg[5]/P0001  ;
	input \u0_slt1_r_reg[6]/P0001  ;
	input \u0_slt1_r_reg[7]/P0001  ;
	input \u0_slt1_r_reg[8]/P0001  ;
	input \u0_slt1_r_reg[9]/P0001  ;
	input \u0_slt2_r_reg[0]/P0001  ;
	input \u0_slt2_r_reg[10]/P0001  ;
	input \u0_slt2_r_reg[11]/P0001  ;
	input \u0_slt2_r_reg[12]/P0001  ;
	input \u0_slt2_r_reg[13]/P0001  ;
	input \u0_slt2_r_reg[14]/P0001  ;
	input \u0_slt2_r_reg[15]/P0001  ;
	input \u0_slt2_r_reg[16]/P0001  ;
	input \u0_slt2_r_reg[17]/P0001  ;
	input \u0_slt2_r_reg[18]/P0001  ;
	input \u0_slt2_r_reg[19]/P0001  ;
	input \u0_slt2_r_reg[1]/P0001  ;
	input \u0_slt2_r_reg[2]/P0001  ;
	input \u0_slt2_r_reg[3]/P0001  ;
	input \u0_slt2_r_reg[4]/P0001  ;
	input \u0_slt2_r_reg[5]/P0001  ;
	input \u0_slt2_r_reg[6]/P0001  ;
	input \u0_slt2_r_reg[7]/P0001  ;
	input \u0_slt2_r_reg[8]/P0001  ;
	input \u0_slt2_r_reg[9]/P0001  ;
	input \u0_slt3_r_reg[0]/P0001  ;
	input \u0_slt3_r_reg[10]/P0001  ;
	input \u0_slt3_r_reg[11]/P0001  ;
	input \u0_slt3_r_reg[12]/P0001  ;
	input \u0_slt3_r_reg[13]/P0001  ;
	input \u0_slt3_r_reg[14]/P0001  ;
	input \u0_slt3_r_reg[15]/P0001  ;
	input \u0_slt3_r_reg[16]/P0001  ;
	input \u0_slt3_r_reg[17]/P0001  ;
	input \u0_slt3_r_reg[18]/P0001  ;
	input \u0_slt3_r_reg[19]/P0001  ;
	input \u0_slt3_r_reg[1]/P0001  ;
	input \u0_slt3_r_reg[2]/P0001  ;
	input \u0_slt3_r_reg[3]/P0001  ;
	input \u0_slt3_r_reg[4]/P0001  ;
	input \u0_slt3_r_reg[5]/P0001  ;
	input \u0_slt3_r_reg[6]/P0001  ;
	input \u0_slt3_r_reg[7]/P0001  ;
	input \u0_slt3_r_reg[8]/P0001  ;
	input \u0_slt3_r_reg[9]/P0001  ;
	input \u0_slt4_r_reg[0]/P0001  ;
	input \u0_slt4_r_reg[10]/P0001  ;
	input \u0_slt4_r_reg[11]/P0001  ;
	input \u0_slt4_r_reg[12]/P0001  ;
	input \u0_slt4_r_reg[13]/P0001  ;
	input \u0_slt4_r_reg[14]/P0001  ;
	input \u0_slt4_r_reg[15]/P0001  ;
	input \u0_slt4_r_reg[16]/P0001  ;
	input \u0_slt4_r_reg[17]/P0001  ;
	input \u0_slt4_r_reg[18]/P0001  ;
	input \u0_slt4_r_reg[19]/P0001  ;
	input \u0_slt4_r_reg[1]/P0001  ;
	input \u0_slt4_r_reg[2]/P0001  ;
	input \u0_slt4_r_reg[3]/P0001  ;
	input \u0_slt4_r_reg[4]/P0001  ;
	input \u0_slt4_r_reg[5]/P0001  ;
	input \u0_slt4_r_reg[6]/P0001  ;
	input \u0_slt4_r_reg[7]/P0001  ;
	input \u0_slt4_r_reg[8]/P0001  ;
	input \u0_slt4_r_reg[9]/P0001  ;
	input \u0_slt5_r_reg[0]/P0001  ;
	input \u0_slt5_r_reg[10]/P0001  ;
	input \u0_slt5_r_reg[11]/P0001  ;
	input \u0_slt5_r_reg[12]/P0001  ;
	input \u0_slt5_r_reg[13]/P0001  ;
	input \u0_slt5_r_reg[14]/P0001  ;
	input \u0_slt5_r_reg[15]/P0001  ;
	input \u0_slt5_r_reg[16]/P0001  ;
	input \u0_slt5_r_reg[17]/P0001  ;
	input \u0_slt5_r_reg[18]/P0001  ;
	input \u0_slt5_r_reg[19]/P0001  ;
	input \u0_slt5_r_reg[1]/P0001  ;
	input \u0_slt5_r_reg[2]/P0001  ;
	input \u0_slt5_r_reg[3]/P0001  ;
	input \u0_slt5_r_reg[4]/P0001  ;
	input \u0_slt5_r_reg[5]/P0001  ;
	input \u0_slt5_r_reg[6]/P0001  ;
	input \u0_slt5_r_reg[7]/P0001  ;
	input \u0_slt5_r_reg[8]/P0001  ;
	input \u0_slt5_r_reg[9]/P0001  ;
	input \u0_slt6_r_reg[0]/P0001  ;
	input \u0_slt6_r_reg[10]/P0001  ;
	input \u0_slt6_r_reg[11]/P0001  ;
	input \u0_slt6_r_reg[12]/P0001  ;
	input \u0_slt6_r_reg[13]/P0001  ;
	input \u0_slt6_r_reg[14]/P0001  ;
	input \u0_slt6_r_reg[15]/P0001  ;
	input \u0_slt6_r_reg[16]/P0001  ;
	input \u0_slt6_r_reg[17]/P0001  ;
	input \u0_slt6_r_reg[18]/P0001  ;
	input \u0_slt6_r_reg[19]/P0001  ;
	input \u0_slt6_r_reg[1]/P0001  ;
	input \u0_slt6_r_reg[2]/P0001  ;
	input \u0_slt6_r_reg[3]/P0001  ;
	input \u0_slt6_r_reg[4]/P0001  ;
	input \u0_slt6_r_reg[5]/P0001  ;
	input \u0_slt6_r_reg[6]/P0001  ;
	input \u0_slt6_r_reg[7]/P0001  ;
	input \u0_slt6_r_reg[8]/P0001  ;
	input \u0_slt6_r_reg[9]/P0001  ;
	input \u0_slt7_r_reg[0]/P0001  ;
	input \u0_slt7_r_reg[10]/P0001  ;
	input \u0_slt7_r_reg[11]/P0001  ;
	input \u0_slt7_r_reg[12]/P0001  ;
	input \u0_slt7_r_reg[13]/P0001  ;
	input \u0_slt7_r_reg[14]/P0001  ;
	input \u0_slt7_r_reg[15]/P0001  ;
	input \u0_slt7_r_reg[16]/P0001  ;
	input \u0_slt7_r_reg[17]/P0001  ;
	input \u0_slt7_r_reg[18]/P0001  ;
	input \u0_slt7_r_reg[19]/P0001  ;
	input \u0_slt7_r_reg[1]/P0001  ;
	input \u0_slt7_r_reg[2]/P0001  ;
	input \u0_slt7_r_reg[3]/P0001  ;
	input \u0_slt7_r_reg[4]/P0001  ;
	input \u0_slt7_r_reg[5]/P0001  ;
	input \u0_slt7_r_reg[6]/P0001  ;
	input \u0_slt7_r_reg[7]/P0001  ;
	input \u0_slt7_r_reg[8]/P0001  ;
	input \u0_slt7_r_reg[9]/P0001  ;
	input \u0_slt8_r_reg[0]/P0001  ;
	input \u0_slt8_r_reg[10]/P0001  ;
	input \u0_slt8_r_reg[11]/P0001  ;
	input \u0_slt8_r_reg[12]/P0001  ;
	input \u0_slt8_r_reg[13]/P0001  ;
	input \u0_slt8_r_reg[14]/P0001  ;
	input \u0_slt8_r_reg[15]/P0001  ;
	input \u0_slt8_r_reg[16]/P0001  ;
	input \u0_slt8_r_reg[17]/P0001  ;
	input \u0_slt8_r_reg[18]/P0001  ;
	input \u0_slt8_r_reg[19]/P0001  ;
	input \u0_slt8_r_reg[1]/P0001  ;
	input \u0_slt8_r_reg[2]/P0001  ;
	input \u0_slt8_r_reg[3]/P0001  ;
	input \u0_slt8_r_reg[4]/P0001  ;
	input \u0_slt8_r_reg[5]/P0001  ;
	input \u0_slt8_r_reg[6]/P0001  ;
	input \u0_slt8_r_reg[7]/P0001  ;
	input \u0_slt8_r_reg[8]/P0001  ;
	input \u0_slt8_r_reg[9]/P0001  ;
	input \u0_slt9_r_reg[0]/P0001  ;
	input \u0_slt9_r_reg[10]/P0001  ;
	input \u0_slt9_r_reg[11]/P0001  ;
	input \u0_slt9_r_reg[12]/P0001  ;
	input \u0_slt9_r_reg[13]/P0001  ;
	input \u0_slt9_r_reg[14]/P0001  ;
	input \u0_slt9_r_reg[15]/P0001  ;
	input \u0_slt9_r_reg[16]/P0001  ;
	input \u0_slt9_r_reg[17]/P0001  ;
	input \u0_slt9_r_reg[18]/P0001  ;
	input \u0_slt9_r_reg[19]/P0001  ;
	input \u0_slt9_r_reg[1]/P0001  ;
	input \u0_slt9_r_reg[2]/P0001  ;
	input \u0_slt9_r_reg[3]/P0001  ;
	input \u0_slt9_r_reg[4]/P0001  ;
	input \u0_slt9_r_reg[5]/P0001  ;
	input \u0_slt9_r_reg[6]/P0001  ;
	input \u0_slt9_r_reg[7]/P0001  ;
	input \u0_slt9_r_reg[8]/P0001  ;
	input \u0_slt9_r_reg[9]/P0001  ;
	input \u10_din_tmp1_reg[0]/P0001  ;
	input \u10_din_tmp1_reg[10]/P0001  ;
	input \u10_din_tmp1_reg[11]/P0001  ;
	input \u10_din_tmp1_reg[12]/P0001  ;
	input \u10_din_tmp1_reg[13]/P0001  ;
	input \u10_din_tmp1_reg[14]/P0001  ;
	input \u10_din_tmp1_reg[15]/P0001  ;
	input \u10_din_tmp1_reg[1]/P0001  ;
	input \u10_din_tmp1_reg[2]/P0001  ;
	input \u10_din_tmp1_reg[3]/P0001  ;
	input \u10_din_tmp1_reg[4]/P0001  ;
	input \u10_din_tmp1_reg[5]/P0001  ;
	input \u10_din_tmp1_reg[6]/P0001  ;
	input \u10_din_tmp1_reg[7]/P0001  ;
	input \u10_din_tmp1_reg[8]/P0001  ;
	input \u10_din_tmp1_reg[9]/P0001  ;
	input \u10_dout_reg[0]/P0001  ;
	input \u10_dout_reg[10]/P0001  ;
	input \u10_dout_reg[11]/P0001  ;
	input \u10_dout_reg[12]/P0001  ;
	input \u10_dout_reg[13]/P0001  ;
	input \u10_dout_reg[14]/P0001  ;
	input \u10_dout_reg[15]/P0001  ;
	input \u10_dout_reg[16]/P0001  ;
	input \u10_dout_reg[17]/P0001  ;
	input \u10_dout_reg[18]/P0001  ;
	input \u10_dout_reg[19]/P0001  ;
	input \u10_dout_reg[1]/P0001  ;
	input \u10_dout_reg[20]/P0001  ;
	input \u10_dout_reg[21]/P0001  ;
	input \u10_dout_reg[22]/P0001  ;
	input \u10_dout_reg[23]/P0001  ;
	input \u10_dout_reg[24]/P0001  ;
	input \u10_dout_reg[25]/P0001  ;
	input \u10_dout_reg[26]/P0001  ;
	input \u10_dout_reg[27]/P0001  ;
	input \u10_dout_reg[28]/P0001  ;
	input \u10_dout_reg[29]/P0001  ;
	input \u10_dout_reg[2]/P0001  ;
	input \u10_dout_reg[30]/P0001  ;
	input \u10_dout_reg[31]/P0001  ;
	input \u10_dout_reg[3]/P0001  ;
	input \u10_dout_reg[4]/P0001  ;
	input \u10_dout_reg[5]/P0001  ;
	input \u10_dout_reg[6]/P0001  ;
	input \u10_dout_reg[7]/P0001  ;
	input \u10_dout_reg[8]/P0001  ;
	input \u10_dout_reg[9]/P0001  ;
	input \u10_empty_reg/P0001  ;
	input \u10_full_reg/NET0131  ;
	input \u10_mem_reg[0][0]/P0001  ;
	input \u10_mem_reg[0][10]/P0001  ;
	input \u10_mem_reg[0][11]/P0001  ;
	input \u10_mem_reg[0][12]/P0001  ;
	input \u10_mem_reg[0][13]/P0001  ;
	input \u10_mem_reg[0][14]/P0001  ;
	input \u10_mem_reg[0][15]/P0001  ;
	input \u10_mem_reg[0][16]/P0001  ;
	input \u10_mem_reg[0][17]/P0001  ;
	input \u10_mem_reg[0][18]/P0001  ;
	input \u10_mem_reg[0][19]/P0001  ;
	input \u10_mem_reg[0][1]/P0001  ;
	input \u10_mem_reg[0][20]/P0001  ;
	input \u10_mem_reg[0][21]/P0001  ;
	input \u10_mem_reg[0][22]/P0001  ;
	input \u10_mem_reg[0][23]/P0001  ;
	input \u10_mem_reg[0][24]/P0001  ;
	input \u10_mem_reg[0][25]/P0001  ;
	input \u10_mem_reg[0][26]/P0001  ;
	input \u10_mem_reg[0][27]/P0001  ;
	input \u10_mem_reg[0][28]/P0001  ;
	input \u10_mem_reg[0][29]/P0001  ;
	input \u10_mem_reg[0][2]/P0001  ;
	input \u10_mem_reg[0][30]/P0001  ;
	input \u10_mem_reg[0][31]/P0001  ;
	input \u10_mem_reg[0][3]/P0001  ;
	input \u10_mem_reg[0][4]/P0001  ;
	input \u10_mem_reg[0][5]/P0001  ;
	input \u10_mem_reg[0][6]/P0001  ;
	input \u10_mem_reg[0][7]/P0001  ;
	input \u10_mem_reg[0][8]/P0001  ;
	input \u10_mem_reg[0][9]/P0001  ;
	input \u10_mem_reg[1][0]/P0001  ;
	input \u10_mem_reg[1][10]/P0001  ;
	input \u10_mem_reg[1][11]/P0001  ;
	input \u10_mem_reg[1][12]/P0001  ;
	input \u10_mem_reg[1][13]/P0001  ;
	input \u10_mem_reg[1][14]/P0001  ;
	input \u10_mem_reg[1][15]/P0001  ;
	input \u10_mem_reg[1][16]/P0001  ;
	input \u10_mem_reg[1][17]/P0001  ;
	input \u10_mem_reg[1][18]/P0001  ;
	input \u10_mem_reg[1][19]/P0001  ;
	input \u10_mem_reg[1][1]/P0001  ;
	input \u10_mem_reg[1][20]/P0001  ;
	input \u10_mem_reg[1][21]/P0001  ;
	input \u10_mem_reg[1][22]/P0001  ;
	input \u10_mem_reg[1][23]/P0001  ;
	input \u10_mem_reg[1][24]/P0001  ;
	input \u10_mem_reg[1][25]/P0001  ;
	input \u10_mem_reg[1][26]/P0001  ;
	input \u10_mem_reg[1][27]/P0001  ;
	input \u10_mem_reg[1][28]/P0001  ;
	input \u10_mem_reg[1][29]/P0001  ;
	input \u10_mem_reg[1][2]/P0001  ;
	input \u10_mem_reg[1][30]/P0001  ;
	input \u10_mem_reg[1][31]/P0001  ;
	input \u10_mem_reg[1][3]/P0001  ;
	input \u10_mem_reg[1][4]/P0001  ;
	input \u10_mem_reg[1][5]/P0001  ;
	input \u10_mem_reg[1][6]/P0001  ;
	input \u10_mem_reg[1][7]/P0001  ;
	input \u10_mem_reg[1][8]/P0001  ;
	input \u10_mem_reg[1][9]/P0001  ;
	input \u10_mem_reg[2][0]/P0001  ;
	input \u10_mem_reg[2][10]/P0001  ;
	input \u10_mem_reg[2][11]/P0001  ;
	input \u10_mem_reg[2][12]/P0001  ;
	input \u10_mem_reg[2][13]/P0001  ;
	input \u10_mem_reg[2][14]/P0001  ;
	input \u10_mem_reg[2][15]/P0001  ;
	input \u10_mem_reg[2][16]/P0001  ;
	input \u10_mem_reg[2][17]/P0001  ;
	input \u10_mem_reg[2][18]/P0001  ;
	input \u10_mem_reg[2][19]/P0001  ;
	input \u10_mem_reg[2][1]/P0001  ;
	input \u10_mem_reg[2][20]/P0001  ;
	input \u10_mem_reg[2][21]/P0001  ;
	input \u10_mem_reg[2][22]/P0001  ;
	input \u10_mem_reg[2][23]/P0001  ;
	input \u10_mem_reg[2][24]/P0001  ;
	input \u10_mem_reg[2][25]/P0001  ;
	input \u10_mem_reg[2][26]/P0001  ;
	input \u10_mem_reg[2][27]/P0001  ;
	input \u10_mem_reg[2][28]/P0001  ;
	input \u10_mem_reg[2][29]/P0001  ;
	input \u10_mem_reg[2][2]/P0001  ;
	input \u10_mem_reg[2][30]/P0001  ;
	input \u10_mem_reg[2][31]/P0001  ;
	input \u10_mem_reg[2][3]/P0001  ;
	input \u10_mem_reg[2][4]/P0001  ;
	input \u10_mem_reg[2][5]/P0001  ;
	input \u10_mem_reg[2][6]/P0001  ;
	input \u10_mem_reg[2][7]/P0001  ;
	input \u10_mem_reg[2][8]/P0001  ;
	input \u10_mem_reg[2][9]/P0001  ;
	input \u10_mem_reg[3][0]/P0001  ;
	input \u10_mem_reg[3][10]/P0001  ;
	input \u10_mem_reg[3][11]/P0001  ;
	input \u10_mem_reg[3][12]/P0001  ;
	input \u10_mem_reg[3][13]/P0001  ;
	input \u10_mem_reg[3][14]/P0001  ;
	input \u10_mem_reg[3][15]/P0001  ;
	input \u10_mem_reg[3][16]/P0001  ;
	input \u10_mem_reg[3][17]/P0001  ;
	input \u10_mem_reg[3][18]/P0001  ;
	input \u10_mem_reg[3][19]/P0001  ;
	input \u10_mem_reg[3][1]/P0001  ;
	input \u10_mem_reg[3][20]/P0001  ;
	input \u10_mem_reg[3][21]/P0001  ;
	input \u10_mem_reg[3][22]/P0001  ;
	input \u10_mem_reg[3][23]/P0001  ;
	input \u10_mem_reg[3][24]/P0001  ;
	input \u10_mem_reg[3][25]/P0001  ;
	input \u10_mem_reg[3][26]/P0001  ;
	input \u10_mem_reg[3][27]/P0001  ;
	input \u10_mem_reg[3][28]/P0001  ;
	input \u10_mem_reg[3][29]/P0001  ;
	input \u10_mem_reg[3][2]/P0001  ;
	input \u10_mem_reg[3][30]/P0001  ;
	input \u10_mem_reg[3][31]/P0001  ;
	input \u10_mem_reg[3][3]/P0001  ;
	input \u10_mem_reg[3][4]/P0001  ;
	input \u10_mem_reg[3][5]/P0001  ;
	input \u10_mem_reg[3][6]/P0001  ;
	input \u10_mem_reg[3][7]/P0001  ;
	input \u10_mem_reg[3][8]/P0001  ;
	input \u10_mem_reg[3][9]/P0001  ;
	input \u10_rp_reg[0]/P0001  ;
	input \u10_rp_reg[1]/P0001  ;
	input \u10_rp_reg[2]/P0001  ;
	input \u10_status_reg[0]/P0001  ;
	input \u10_status_reg[1]/P0001  ;
	input \u10_wp_reg[0]/NET0131  ;
	input \u10_wp_reg[1]/P0001  ;
	input \u10_wp_reg[2]/P0001  ;
	input \u10_wp_reg[3]/P0001  ;
	input \u11_din_tmp1_reg[0]/P0001  ;
	input \u11_din_tmp1_reg[10]/P0001  ;
	input \u11_din_tmp1_reg[11]/P0001  ;
	input \u11_din_tmp1_reg[12]/P0001  ;
	input \u11_din_tmp1_reg[13]/P0001  ;
	input \u11_din_tmp1_reg[14]/P0001  ;
	input \u11_din_tmp1_reg[15]/P0001  ;
	input \u11_din_tmp1_reg[1]/P0001  ;
	input \u11_din_tmp1_reg[2]/P0001  ;
	input \u11_din_tmp1_reg[3]/P0001  ;
	input \u11_din_tmp1_reg[4]/P0001  ;
	input \u11_din_tmp1_reg[5]/P0001  ;
	input \u11_din_tmp1_reg[6]/P0001  ;
	input \u11_din_tmp1_reg[7]/P0001  ;
	input \u11_din_tmp1_reg[8]/P0001  ;
	input \u11_din_tmp1_reg[9]/P0001  ;
	input \u11_dout_reg[0]/P0001  ;
	input \u11_dout_reg[10]/P0001  ;
	input \u11_dout_reg[11]/P0001  ;
	input \u11_dout_reg[12]/P0001  ;
	input \u11_dout_reg[13]/P0001  ;
	input \u11_dout_reg[14]/P0001  ;
	input \u11_dout_reg[15]/P0001  ;
	input \u11_dout_reg[16]/P0001  ;
	input \u11_dout_reg[17]/P0001  ;
	input \u11_dout_reg[18]/P0001  ;
	input \u11_dout_reg[19]/P0001  ;
	input \u11_dout_reg[1]/P0001  ;
	input \u11_dout_reg[20]/P0001  ;
	input \u11_dout_reg[21]/P0001  ;
	input \u11_dout_reg[22]/P0001  ;
	input \u11_dout_reg[23]/P0001  ;
	input \u11_dout_reg[24]/P0001  ;
	input \u11_dout_reg[25]/P0001  ;
	input \u11_dout_reg[26]/P0001  ;
	input \u11_dout_reg[27]/P0001  ;
	input \u11_dout_reg[28]/P0001  ;
	input \u11_dout_reg[29]/P0001  ;
	input \u11_dout_reg[2]/P0001  ;
	input \u11_dout_reg[30]/P0001  ;
	input \u11_dout_reg[31]/P0001  ;
	input \u11_dout_reg[3]/P0001  ;
	input \u11_dout_reg[4]/P0001  ;
	input \u11_dout_reg[5]/P0001  ;
	input \u11_dout_reg[6]/P0001  ;
	input \u11_dout_reg[7]/P0001  ;
	input \u11_dout_reg[8]/P0001  ;
	input \u11_dout_reg[9]/P0001  ;
	input \u11_empty_reg/P0001  ;
	input \u11_full_reg/NET0131  ;
	input \u11_mem_reg[0][0]/P0001  ;
	input \u11_mem_reg[0][10]/P0001  ;
	input \u11_mem_reg[0][11]/P0001  ;
	input \u11_mem_reg[0][12]/P0001  ;
	input \u11_mem_reg[0][13]/P0001  ;
	input \u11_mem_reg[0][14]/P0001  ;
	input \u11_mem_reg[0][15]/P0001  ;
	input \u11_mem_reg[0][16]/P0001  ;
	input \u11_mem_reg[0][17]/P0001  ;
	input \u11_mem_reg[0][18]/P0001  ;
	input \u11_mem_reg[0][19]/P0001  ;
	input \u11_mem_reg[0][1]/P0001  ;
	input \u11_mem_reg[0][20]/P0001  ;
	input \u11_mem_reg[0][21]/P0001  ;
	input \u11_mem_reg[0][22]/P0001  ;
	input \u11_mem_reg[0][23]/P0001  ;
	input \u11_mem_reg[0][24]/P0001  ;
	input \u11_mem_reg[0][25]/P0001  ;
	input \u11_mem_reg[0][26]/P0001  ;
	input \u11_mem_reg[0][27]/P0001  ;
	input \u11_mem_reg[0][28]/P0001  ;
	input \u11_mem_reg[0][29]/P0001  ;
	input \u11_mem_reg[0][2]/P0001  ;
	input \u11_mem_reg[0][30]/P0001  ;
	input \u11_mem_reg[0][31]/P0001  ;
	input \u11_mem_reg[0][3]/P0001  ;
	input \u11_mem_reg[0][4]/P0001  ;
	input \u11_mem_reg[0][5]/P0001  ;
	input \u11_mem_reg[0][6]/P0001  ;
	input \u11_mem_reg[0][7]/P0001  ;
	input \u11_mem_reg[0][8]/P0001  ;
	input \u11_mem_reg[0][9]/P0001  ;
	input \u11_mem_reg[1][0]/P0001  ;
	input \u11_mem_reg[1][10]/P0001  ;
	input \u11_mem_reg[1][11]/P0001  ;
	input \u11_mem_reg[1][12]/P0001  ;
	input \u11_mem_reg[1][13]/P0001  ;
	input \u11_mem_reg[1][14]/P0001  ;
	input \u11_mem_reg[1][15]/P0001  ;
	input \u11_mem_reg[1][16]/P0001  ;
	input \u11_mem_reg[1][17]/P0001  ;
	input \u11_mem_reg[1][18]/P0001  ;
	input \u11_mem_reg[1][19]/P0001  ;
	input \u11_mem_reg[1][1]/P0001  ;
	input \u11_mem_reg[1][20]/P0001  ;
	input \u11_mem_reg[1][21]/P0001  ;
	input \u11_mem_reg[1][22]/P0001  ;
	input \u11_mem_reg[1][23]/P0001  ;
	input \u11_mem_reg[1][24]/P0001  ;
	input \u11_mem_reg[1][25]/P0001  ;
	input \u11_mem_reg[1][26]/P0001  ;
	input \u11_mem_reg[1][27]/P0001  ;
	input \u11_mem_reg[1][28]/P0001  ;
	input \u11_mem_reg[1][29]/P0001  ;
	input \u11_mem_reg[1][2]/P0001  ;
	input \u11_mem_reg[1][30]/P0001  ;
	input \u11_mem_reg[1][31]/P0001  ;
	input \u11_mem_reg[1][3]/P0001  ;
	input \u11_mem_reg[1][4]/P0001  ;
	input \u11_mem_reg[1][5]/P0001  ;
	input \u11_mem_reg[1][6]/P0001  ;
	input \u11_mem_reg[1][7]/P0001  ;
	input \u11_mem_reg[1][8]/P0001  ;
	input \u11_mem_reg[1][9]/P0001  ;
	input \u11_mem_reg[2][0]/P0001  ;
	input \u11_mem_reg[2][10]/P0001  ;
	input \u11_mem_reg[2][11]/P0001  ;
	input \u11_mem_reg[2][12]/P0001  ;
	input \u11_mem_reg[2][13]/P0001  ;
	input \u11_mem_reg[2][14]/P0001  ;
	input \u11_mem_reg[2][15]/P0001  ;
	input \u11_mem_reg[2][16]/P0001  ;
	input \u11_mem_reg[2][17]/P0001  ;
	input \u11_mem_reg[2][18]/P0001  ;
	input \u11_mem_reg[2][19]/P0001  ;
	input \u11_mem_reg[2][1]/P0001  ;
	input \u11_mem_reg[2][20]/P0001  ;
	input \u11_mem_reg[2][21]/P0001  ;
	input \u11_mem_reg[2][22]/P0001  ;
	input \u11_mem_reg[2][23]/P0001  ;
	input \u11_mem_reg[2][24]/P0001  ;
	input \u11_mem_reg[2][25]/P0001  ;
	input \u11_mem_reg[2][26]/P0001  ;
	input \u11_mem_reg[2][27]/P0001  ;
	input \u11_mem_reg[2][28]/P0001  ;
	input \u11_mem_reg[2][29]/P0001  ;
	input \u11_mem_reg[2][2]/P0001  ;
	input \u11_mem_reg[2][30]/P0001  ;
	input \u11_mem_reg[2][31]/P0001  ;
	input \u11_mem_reg[2][3]/P0001  ;
	input \u11_mem_reg[2][4]/P0001  ;
	input \u11_mem_reg[2][5]/P0001  ;
	input \u11_mem_reg[2][6]/P0001  ;
	input \u11_mem_reg[2][7]/P0001  ;
	input \u11_mem_reg[2][8]/P0001  ;
	input \u11_mem_reg[2][9]/P0001  ;
	input \u11_mem_reg[3][0]/P0001  ;
	input \u11_mem_reg[3][10]/P0001  ;
	input \u11_mem_reg[3][11]/P0001  ;
	input \u11_mem_reg[3][12]/P0001  ;
	input \u11_mem_reg[3][13]/P0001  ;
	input \u11_mem_reg[3][14]/P0001  ;
	input \u11_mem_reg[3][15]/P0001  ;
	input \u11_mem_reg[3][16]/P0001  ;
	input \u11_mem_reg[3][17]/P0001  ;
	input \u11_mem_reg[3][18]/P0001  ;
	input \u11_mem_reg[3][19]/P0001  ;
	input \u11_mem_reg[3][1]/P0001  ;
	input \u11_mem_reg[3][20]/P0001  ;
	input \u11_mem_reg[3][21]/P0001  ;
	input \u11_mem_reg[3][22]/P0001  ;
	input \u11_mem_reg[3][23]/P0001  ;
	input \u11_mem_reg[3][24]/P0001  ;
	input \u11_mem_reg[3][25]/P0001  ;
	input \u11_mem_reg[3][26]/P0001  ;
	input \u11_mem_reg[3][27]/P0001  ;
	input \u11_mem_reg[3][28]/P0001  ;
	input \u11_mem_reg[3][29]/P0001  ;
	input \u11_mem_reg[3][2]/P0001  ;
	input \u11_mem_reg[3][30]/P0001  ;
	input \u11_mem_reg[3][31]/P0001  ;
	input \u11_mem_reg[3][3]/P0001  ;
	input \u11_mem_reg[3][4]/P0001  ;
	input \u11_mem_reg[3][5]/P0001  ;
	input \u11_mem_reg[3][6]/P0001  ;
	input \u11_mem_reg[3][7]/P0001  ;
	input \u11_mem_reg[3][8]/P0001  ;
	input \u11_mem_reg[3][9]/P0001  ;
	input \u11_rp_reg[0]/P0001  ;
	input \u11_rp_reg[1]/P0001  ;
	input \u11_rp_reg[2]/P0001  ;
	input \u11_status_reg[0]/P0001  ;
	input \u11_status_reg[1]/P0001  ;
	input \u11_wp_reg[0]/NET0131  ;
	input \u11_wp_reg[1]/P0001  ;
	input \u11_wp_reg[2]/P0001  ;
	input \u11_wp_reg[3]/P0001  ;
	input \u12_dout_reg[0]/P0001  ;
	input \u12_dout_reg[10]/P0001  ;
	input \u12_dout_reg[11]/P0001  ;
	input \u12_dout_reg[12]/P0001  ;
	input \u12_dout_reg[13]/P0001  ;
	input \u12_dout_reg[14]/P0001  ;
	input \u12_dout_reg[15]/P0001  ;
	input \u12_dout_reg[16]/P0001  ;
	input \u12_dout_reg[17]/P0001  ;
	input \u12_dout_reg[18]/P0001  ;
	input \u12_dout_reg[19]/P0001  ;
	input \u12_dout_reg[1]/P0001  ;
	input \u12_dout_reg[20]/P0001  ;
	input \u12_dout_reg[21]/P0001  ;
	input \u12_dout_reg[22]/P0001  ;
	input \u12_dout_reg[23]/P0001  ;
	input \u12_dout_reg[24]/P0001  ;
	input \u12_dout_reg[25]/P0001  ;
	input \u12_dout_reg[26]/P0001  ;
	input \u12_dout_reg[27]/P0001  ;
	input \u12_dout_reg[28]/P0001  ;
	input \u12_dout_reg[29]/P0001  ;
	input \u12_dout_reg[2]/P0001  ;
	input \u12_dout_reg[30]/P0001  ;
	input \u12_dout_reg[31]/P0001  ;
	input \u12_dout_reg[3]/P0001  ;
	input \u12_dout_reg[4]/P0001  ;
	input \u12_dout_reg[5]/P0001  ;
	input \u12_dout_reg[6]/P0001  ;
	input \u12_dout_reg[7]/P0001  ;
	input \u12_dout_reg[8]/P0001  ;
	input \u12_dout_reg[9]/P0001  ;
	input \u12_i3_re_reg/NET0131  ;
	input \u12_i4_re_reg/P0001  ;
	input \u12_i6_re_reg/NET0131  ;
	input \u12_o3_we_reg/P0001  ;
	input \u12_o4_we_reg/P0001  ;
	input \u12_o6_we_reg/P0001  ;
	input \u12_o7_we_reg/P0001  ;
	input \u12_o8_we_reg/P0001  ;
	input \u12_o9_we_reg/P0001  ;
	input \u12_re1_reg/P0001  ;
	input \u12_re2_reg/NET0131  ;
	input \u12_rf_we_reg/P0001  ;
	input \u12_we1_reg/P0001  ;
	input \u12_we2_reg/P0001  ;
	input \u13_ac97_rst_force_reg/P0001  ;
	input \u13_crac_dout_r_reg[0]/P0001  ;
	input \u13_crac_dout_r_reg[10]/P0001  ;
	input \u13_crac_dout_r_reg[11]/P0001  ;
	input \u13_crac_dout_r_reg[12]/P0001  ;
	input \u13_crac_dout_r_reg[13]/P0001  ;
	input \u13_crac_dout_r_reg[14]/P0001  ;
	input \u13_crac_dout_r_reg[15]/P0001  ;
	input \u13_crac_dout_r_reg[1]/P0001  ;
	input \u13_crac_dout_r_reg[2]/P0001  ;
	input \u13_crac_dout_r_reg[3]/P0001  ;
	input \u13_crac_dout_r_reg[4]/P0001  ;
	input \u13_crac_dout_r_reg[5]/P0001  ;
	input \u13_crac_dout_r_reg[6]/P0001  ;
	input \u13_crac_dout_r_reg[7]/P0001  ;
	input \u13_crac_dout_r_reg[8]/P0001  ;
	input \u13_crac_dout_r_reg[9]/P0001  ;
	input \u13_crac_r_reg[0]/NET0131  ;
	input \u13_crac_r_reg[1]/NET0131  ;
	input \u13_crac_r_reg[2]/NET0131  ;
	input \u13_crac_r_reg[3]/NET0131  ;
	input \u13_crac_r_reg[4]/NET0131  ;
	input \u13_crac_r_reg[5]/NET0131  ;
	input \u13_crac_r_reg[6]/NET0131  ;
	input \u13_crac_r_reg[7]/NET0131  ;
	input \u13_icc_r_reg[0]/NET0131  ;
	input \u13_icc_r_reg[10]/NET0131  ;
	input \u13_icc_r_reg[11]/NET0131  ;
	input \u13_icc_r_reg[12]/NET0131  ;
	input \u13_icc_r_reg[13]/NET0131  ;
	input \u13_icc_r_reg[14]/NET0131  ;
	input \u13_icc_r_reg[15]/NET0131  ;
	input \u13_icc_r_reg[16]/NET0131  ;
	input \u13_icc_r_reg[17]/NET0131  ;
	input \u13_icc_r_reg[18]/NET0131  ;
	input \u13_icc_r_reg[19]/NET0131  ;
	input \u13_icc_r_reg[1]/NET0131  ;
	input \u13_icc_r_reg[20]/NET0131  ;
	input \u13_icc_r_reg[21]/NET0131  ;
	input \u13_icc_r_reg[22]/NET0131  ;
	input \u13_icc_r_reg[23]/NET0131  ;
	input \u13_icc_r_reg[2]/NET0131  ;
	input \u13_icc_r_reg[3]/NET0131  ;
	input \u13_icc_r_reg[4]/NET0131  ;
	input \u13_icc_r_reg[5]/NET0131  ;
	input \u13_icc_r_reg[6]/NET0131  ;
	input \u13_icc_r_reg[7]/NET0131  ;
	input \u13_icc_r_reg[8]/NET0131  ;
	input \u13_icc_r_reg[9]/NET0131  ;
	input \u13_intm_r_reg[0]/NET0131  ;
	input \u13_intm_r_reg[10]/NET0131  ;
	input \u13_intm_r_reg[11]/NET0131  ;
	input \u13_intm_r_reg[12]/NET0131  ;
	input \u13_intm_r_reg[13]/NET0131  ;
	input \u13_intm_r_reg[14]/NET0131  ;
	input \u13_intm_r_reg[15]/NET0131  ;
	input \u13_intm_r_reg[16]/NET0131  ;
	input \u13_intm_r_reg[17]/NET0131  ;
	input \u13_intm_r_reg[18]/NET0131  ;
	input \u13_intm_r_reg[19]/NET0131  ;
	input \u13_intm_r_reg[1]/NET0131  ;
	input \u13_intm_r_reg[20]/NET0131  ;
	input \u13_intm_r_reg[21]/NET0131  ;
	input \u13_intm_r_reg[22]/NET0131  ;
	input \u13_intm_r_reg[23]/NET0131  ;
	input \u13_intm_r_reg[24]/NET0131  ;
	input \u13_intm_r_reg[25]/NET0131  ;
	input \u13_intm_r_reg[26]/NET0131  ;
	input \u13_intm_r_reg[27]/NET0131  ;
	input \u13_intm_r_reg[28]/NET0131  ;
	input \u13_intm_r_reg[2]/NET0131  ;
	input \u13_intm_r_reg[3]/NET0131  ;
	input \u13_intm_r_reg[4]/NET0131  ;
	input \u13_intm_r_reg[5]/NET0131  ;
	input \u13_intm_r_reg[6]/NET0131  ;
	input \u13_intm_r_reg[7]/NET0131  ;
	input \u13_intm_r_reg[8]/NET0131  ;
	input \u13_intm_r_reg[9]/NET0131  ;
	input \u13_ints_r_reg[0]/NET0131  ;
	input \u13_ints_r_reg[10]/NET0131  ;
	input \u13_ints_r_reg[11]/NET0131  ;
	input \u13_ints_r_reg[12]/NET0131  ;
	input \u13_ints_r_reg[13]/NET0131  ;
	input \u13_ints_r_reg[14]/NET0131  ;
	input \u13_ints_r_reg[15]/NET0131  ;
	input \u13_ints_r_reg[16]/NET0131  ;
	input \u13_ints_r_reg[17]/NET0131  ;
	input \u13_ints_r_reg[18]/NET0131  ;
	input \u13_ints_r_reg[19]/NET0131  ;
	input \u13_ints_r_reg[1]/NET0131  ;
	input \u13_ints_r_reg[20]/NET0131  ;
	input \u13_ints_r_reg[21]/NET0131  ;
	input \u13_ints_r_reg[22]/NET0131  ;
	input \u13_ints_r_reg[23]/NET0131  ;
	input \u13_ints_r_reg[24]/NET0131  ;
	input \u13_ints_r_reg[25]/NET0131  ;
	input \u13_ints_r_reg[26]/NET0131  ;
	input \u13_ints_r_reg[27]/NET0131  ;
	input \u13_ints_r_reg[28]/NET0131  ;
	input \u13_ints_r_reg[2]/NET0131  ;
	input \u13_ints_r_reg[3]/NET0131  ;
	input \u13_ints_r_reg[4]/NET0131  ;
	input \u13_ints_r_reg[5]/NET0131  ;
	input \u13_ints_r_reg[6]/NET0131  ;
	input \u13_ints_r_reg[7]/NET0131  ;
	input \u13_ints_r_reg[8]/NET0131  ;
	input \u13_ints_r_reg[9]/NET0131  ;
	input \u13_occ0_r_reg[0]/NET0131  ;
	input \u13_occ0_r_reg[10]/NET0131  ;
	input \u13_occ0_r_reg[11]/NET0131  ;
	input \u13_occ0_r_reg[12]/NET0131  ;
	input \u13_occ0_r_reg[13]/NET0131  ;
	input \u13_occ0_r_reg[14]/NET0131  ;
	input \u13_occ0_r_reg[15]/NET0131  ;
	input \u13_occ0_r_reg[16]/NET0131  ;
	input \u13_occ0_r_reg[17]/NET0131  ;
	input \u13_occ0_r_reg[18]/NET0131  ;
	input \u13_occ0_r_reg[19]/NET0131  ;
	input \u13_occ0_r_reg[1]/NET0131  ;
	input \u13_occ0_r_reg[20]/NET0131  ;
	input \u13_occ0_r_reg[21]/NET0131  ;
	input \u13_occ0_r_reg[22]/NET0131  ;
	input \u13_occ0_r_reg[23]/NET0131  ;
	input \u13_occ0_r_reg[24]/NET0131  ;
	input \u13_occ0_r_reg[25]/NET0131  ;
	input \u13_occ0_r_reg[26]/NET0131  ;
	input \u13_occ0_r_reg[27]/NET0131  ;
	input \u13_occ0_r_reg[28]/NET0131  ;
	input \u13_occ0_r_reg[29]/NET0131  ;
	input \u13_occ0_r_reg[2]/NET0131  ;
	input \u13_occ0_r_reg[30]/NET0131  ;
	input \u13_occ0_r_reg[31]/NET0131  ;
	input \u13_occ0_r_reg[3]/NET0131  ;
	input \u13_occ0_r_reg[4]/NET0131  ;
	input \u13_occ0_r_reg[5]/NET0131  ;
	input \u13_occ0_r_reg[6]/NET0131  ;
	input \u13_occ0_r_reg[7]/NET0131  ;
	input \u13_occ0_r_reg[8]/NET0131  ;
	input \u13_occ0_r_reg[9]/NET0131  ;
	input \u13_occ1_r_reg[0]/NET0131  ;
	input \u13_occ1_r_reg[10]/NET0131  ;
	input \u13_occ1_r_reg[11]/NET0131  ;
	input \u13_occ1_r_reg[12]/NET0131  ;
	input \u13_occ1_r_reg[13]/NET0131  ;
	input \u13_occ1_r_reg[14]/NET0131  ;
	input \u13_occ1_r_reg[15]/NET0131  ;
	input \u13_occ1_r_reg[1]/NET0131  ;
	input \u13_occ1_r_reg[2]/NET0131  ;
	input \u13_occ1_r_reg[3]/NET0131  ;
	input \u13_occ1_r_reg[4]/NET0131  ;
	input \u13_occ1_r_reg[5]/NET0131  ;
	input \u13_occ1_r_reg[6]/NET0131  ;
	input \u13_occ1_r_reg[7]/NET0131  ;
	input \u13_occ1_r_reg[8]/NET0131  ;
	input \u13_occ1_r_reg[9]/NET0131  ;
	input \u13_resume_req_reg/P0001  ;
	input \u14_crac_valid_r_reg/P0001  ;
	input \u14_crac_wr_r_reg/P0001  ;
	input \u14_u0_en_out_l2_reg/P0001  ;
	input \u14_u0_en_out_l_reg/NET0131  ;
	input \u14_u0_full_empty_r_reg/P0001  ;
	input \u14_u1_en_out_l2_reg/P0001  ;
	input \u14_u1_en_out_l_reg/NET0131  ;
	input \u14_u1_full_empty_r_reg/P0001  ;
	input \u14_u2_en_out_l2_reg/P0001  ;
	input \u14_u2_en_out_l_reg/NET0131  ;
	input \u14_u2_full_empty_r_reg/P0001  ;
	input \u14_u3_en_out_l2_reg/P0001  ;
	input \u14_u3_en_out_l_reg/NET0131  ;
	input \u14_u3_full_empty_r_reg/P0001  ;
	input \u14_u4_en_out_l2_reg/P0001  ;
	input \u14_u4_en_out_l_reg/NET0131  ;
	input \u14_u4_full_empty_r_reg/P0001  ;
	input \u14_u5_en_out_l2_reg/P0001  ;
	input \u14_u5_en_out_l_reg/NET0131  ;
	input \u14_u5_full_empty_r_reg/P0001  ;
	input \u14_u6_en_out_l2_reg/P0001  ;
	input \u14_u6_en_out_l_reg/NET0131  ;
	input \u14_u6_full_empty_r_reg/P0001  ;
	input \u14_u7_en_out_l2_reg/P0001  ;
	input \u14_u7_en_out_l_reg/NET0131  ;
	input \u14_u7_full_empty_r_reg/P0001  ;
	input \u14_u8_en_out_l2_reg/P0001  ;
	input \u14_u8_en_out_l_reg/NET0131  ;
	input \u14_u8_full_empty_r_reg/P0001  ;
	input \u15_crac_din_reg[0]/NET0131  ;
	input \u15_crac_din_reg[10]/NET0131  ;
	input \u15_crac_din_reg[11]/NET0131  ;
	input \u15_crac_din_reg[12]/NET0131  ;
	input \u15_crac_din_reg[13]/NET0131  ;
	input \u15_crac_din_reg[14]/NET0131  ;
	input \u15_crac_din_reg[15]/NET0131  ;
	input \u15_crac_din_reg[1]/NET0131  ;
	input \u15_crac_din_reg[2]/NET0131  ;
	input \u15_crac_din_reg[3]/NET0131  ;
	input \u15_crac_din_reg[4]/NET0131  ;
	input \u15_crac_din_reg[5]/NET0131  ;
	input \u15_crac_din_reg[6]/NET0131  ;
	input \u15_crac_din_reg[7]/NET0131  ;
	input \u15_crac_din_reg[8]/NET0131  ;
	input \u15_crac_din_reg[9]/NET0131  ;
	input \u15_crac_rd_done_reg/P0001  ;
	input \u15_crac_rd_reg/NET0131  ;
	input \u15_crac_we_r_reg/P0001  ;
	input \u15_crac_wr_reg/NET0131  ;
	input \u15_rdd1_reg/NET0131  ;
	input \u15_rdd2_reg/NET0131  ;
	input \u15_rdd3_reg/NET0131  ;
	input \u15_valid_r_reg/P0001  ;
	input \u16_u0_dma_req_r1_reg/P0001  ;
	input \u16_u1_dma_req_r1_reg/P0001  ;
	input \u16_u2_dma_req_r1_reg/P0001  ;
	input \u16_u3_dma_req_r1_reg/P0001  ;
	input \u16_u4_dma_req_r1_reg/P0001  ;
	input \u16_u5_dma_req_r1_reg/P0001  ;
	input \u16_u6_dma_req_r1_reg/P0001  ;
	input \u16_u7_dma_req_r1_reg/P0001  ;
	input \u16_u8_dma_req_r1_reg/P0001  ;
	input \u17_int_set_reg[0]/NET0131  ;
	input \u17_int_set_reg[1]/NET0131  ;
	input \u17_int_set_reg[2]/NET0131  ;
	input \u18_int_set_reg[0]/NET0131  ;
	input \u18_int_set_reg[1]/NET0131  ;
	input \u18_int_set_reg[2]/NET0131  ;
	input \u19_int_set_reg[0]/NET0131  ;
	input \u19_int_set_reg[1]/NET0131  ;
	input \u19_int_set_reg[2]/NET0131  ;
	input \u1_slt0_reg[11]/P0001  ;
	input \u1_slt0_reg[12]/P0001  ;
	input \u1_slt0_reg[15]/P0001  ;
	input \u1_slt0_reg[9]/P0001  ;
	input \u1_slt1_reg[10]/P0001  ;
	input \u1_slt1_reg[11]/P0001  ;
	input \u1_slt1_reg[5]/P0001  ;
	input \u1_slt1_reg[6]/P0001  ;
	input \u1_slt1_reg[7]/P0001  ;
	input \u1_slt1_reg[8]/P0001  ;
	input \u1_slt3_reg[0]/P0001  ;
	input \u1_slt3_reg[10]/P0001  ;
	input \u1_slt3_reg[11]/P0001  ;
	input \u1_slt3_reg[12]/P0001  ;
	input \u1_slt3_reg[13]/P0001  ;
	input \u1_slt3_reg[14]/P0001  ;
	input \u1_slt3_reg[15]/P0001  ;
	input \u1_slt3_reg[16]/P0001  ;
	input \u1_slt3_reg[17]/P0001  ;
	input \u1_slt3_reg[18]/P0001  ;
	input \u1_slt3_reg[19]/P0001  ;
	input \u1_slt3_reg[1]/P0001  ;
	input \u1_slt3_reg[2]/P0001  ;
	input \u1_slt3_reg[3]/P0001  ;
	input \u1_slt3_reg[4]/P0001  ;
	input \u1_slt3_reg[5]/P0001  ;
	input \u1_slt3_reg[6]/P0001  ;
	input \u1_slt3_reg[7]/P0001  ;
	input \u1_slt3_reg[8]/P0001  ;
	input \u1_slt3_reg[9]/P0001  ;
	input \u1_slt4_reg[0]/P0001  ;
	input \u1_slt4_reg[10]/P0001  ;
	input \u1_slt4_reg[11]/P0001  ;
	input \u1_slt4_reg[12]/P0001  ;
	input \u1_slt4_reg[13]/P0001  ;
	input \u1_slt4_reg[14]/P0001  ;
	input \u1_slt4_reg[15]/P0001  ;
	input \u1_slt4_reg[16]/P0001  ;
	input \u1_slt4_reg[17]/P0001  ;
	input \u1_slt4_reg[18]/P0001  ;
	input \u1_slt4_reg[19]/P0001  ;
	input \u1_slt4_reg[1]/P0001  ;
	input \u1_slt4_reg[2]/P0001  ;
	input \u1_slt4_reg[3]/P0001  ;
	input \u1_slt4_reg[4]/P0001  ;
	input \u1_slt4_reg[5]/P0001  ;
	input \u1_slt4_reg[6]/P0001  ;
	input \u1_slt4_reg[7]/P0001  ;
	input \u1_slt4_reg[8]/P0001  ;
	input \u1_slt4_reg[9]/P0001  ;
	input \u1_slt6_reg[0]/P0001  ;
	input \u1_slt6_reg[10]/P0001  ;
	input \u1_slt6_reg[11]/P0001  ;
	input \u1_slt6_reg[12]/P0001  ;
	input \u1_slt6_reg[13]/P0001  ;
	input \u1_slt6_reg[14]/P0001  ;
	input \u1_slt6_reg[15]/P0001  ;
	input \u1_slt6_reg[16]/P0001  ;
	input \u1_slt6_reg[17]/P0001  ;
	input \u1_slt6_reg[18]/P0001  ;
	input \u1_slt6_reg[19]/P0001  ;
	input \u1_slt6_reg[1]/P0001  ;
	input \u1_slt6_reg[2]/P0001  ;
	input \u1_slt6_reg[3]/P0001  ;
	input \u1_slt6_reg[4]/P0001  ;
	input \u1_slt6_reg[5]/P0001  ;
	input \u1_slt6_reg[6]/P0001  ;
	input \u1_slt6_reg[7]/P0001  ;
	input \u1_slt6_reg[8]/P0001  ;
	input \u1_slt6_reg[9]/P0001  ;
	input \u1_sr_reg[10]/P0001  ;
	input \u1_sr_reg[11]/P0001  ;
	input \u1_sr_reg[12]/P0001  ;
	input \u1_sr_reg[15]/P0001  ;
	input \u1_sr_reg[5]/P0001  ;
	input \u1_sr_reg[6]/P0001  ;
	input \u1_sr_reg[7]/P0001  ;
	input \u1_sr_reg[8]/P0001  ;
	input \u1_sr_reg[9]/P0001  ;
	input \u20_int_set_reg[0]/NET0131  ;
	input \u20_int_set_reg[1]/NET0131  ;
	input \u20_int_set_reg[2]/NET0131  ;
	input \u21_int_set_reg[0]/NET0131  ;
	input \u21_int_set_reg[1]/NET0131  ;
	input \u21_int_set_reg[2]/NET0131  ;
	input \u22_int_set_reg[0]/NET0131  ;
	input \u22_int_set_reg[1]/NET0131  ;
	input \u22_int_set_reg[2]/NET0131  ;
	input \u23_int_set_reg[0]/NET0131  ;
	input \u23_int_set_reg[1]/NET0131  ;
	input \u23_int_set_reg[2]/NET0131  ;
	input \u24_int_set_reg[0]/NET0131  ;
	input \u24_int_set_reg[1]/NET0131  ;
	input \u24_int_set_reg[2]/NET0131  ;
	input \u25_int_set_reg[0]/NET0131  ;
	input \u25_int_set_reg[1]/NET0131  ;
	input \u25_int_set_reg[2]/NET0131  ;
	input \u26_cnt_reg[0]/NET0131  ;
	input \u26_cnt_reg[1]/NET0131  ;
	input \u26_cnt_reg[2]/NET0131  ;
	input \u26_ps_cnt_reg[0]/NET0131  ;
	input \u26_ps_cnt_reg[1]/NET0131  ;
	input \u26_ps_cnt_reg[2]/NET0131  ;
	input \u26_ps_cnt_reg[3]/NET0131  ;
	input \u26_ps_cnt_reg[4]/NET0131  ;
	input \u26_ps_cnt_reg[5]/NET0131  ;
	input \u2_bit_clk_e_reg/P0001  ;
	input \u2_bit_clk_r1_reg/P0001  ;
	input \u2_bit_clk_r_reg/P0001  ;
	input \u2_cnt_reg[0]/NET0131  ;
	input \u2_cnt_reg[1]/NET0131  ;
	input \u2_cnt_reg[2]/NET0131  ;
	input \u2_cnt_reg[3]/NET0131  ;
	input \u2_cnt_reg[4]/NET0131  ;
	input \u2_cnt_reg[5]/NET0131  ;
	input \u2_cnt_reg[6]/NET0131  ;
	input \u2_cnt_reg[7]/NET0131  ;
	input \u2_ld_reg/P0001  ;
	input \u2_out_le_reg[0]/P0001  ;
	input \u2_out_le_reg[1]/P0001  ;
	input \u2_res_cnt_reg[0]/P0001  ;
	input \u2_res_cnt_reg[1]/P0001  ;
	input \u2_res_cnt_reg[2]/P0001  ;
	input \u2_res_cnt_reg[3]/P0001  ;
	input \u2_sync_beat_reg/P0001  ;
	input \u2_sync_resume_reg/NET0131  ;
	input \u2_to_cnt_reg[0]/NET0131  ;
	input \u2_to_cnt_reg[1]/NET0131  ;
	input \u2_to_cnt_reg[2]/NET0131  ;
	input \u2_to_cnt_reg[3]/NET0131  ;
	input \u2_to_cnt_reg[4]/NET0131  ;
	input \u2_to_cnt_reg[5]/NET0131  ;
	input \u3_dout_reg[0]/P0001  ;
	input \u3_dout_reg[10]/P0001  ;
	input \u3_dout_reg[11]/P0001  ;
	input \u3_dout_reg[12]/P0001  ;
	input \u3_dout_reg[13]/P0001  ;
	input \u3_dout_reg[14]/P0001  ;
	input \u3_dout_reg[15]/P0001  ;
	input \u3_dout_reg[16]/P0001  ;
	input \u3_dout_reg[17]/P0001  ;
	input \u3_dout_reg[18]/P0001  ;
	input \u3_dout_reg[19]/P0001  ;
	input \u3_dout_reg[1]/P0001  ;
	input \u3_dout_reg[2]/P0001  ;
	input \u3_dout_reg[3]/P0001  ;
	input \u3_dout_reg[4]/P0001  ;
	input \u3_dout_reg[5]/P0001  ;
	input \u3_dout_reg[6]/P0001  ;
	input \u3_dout_reg[7]/P0001  ;
	input \u3_dout_reg[8]/P0001  ;
	input \u3_dout_reg[9]/P0001  ;
	input \u3_empty_reg/NET0131  ;
	input \u3_mem_reg[0][0]/NET0131  ;
	input \u3_mem_reg[0][10]/NET0131  ;
	input \u3_mem_reg[0][11]/NET0131  ;
	input \u3_mem_reg[0][12]/NET0131  ;
	input \u3_mem_reg[0][13]/NET0131  ;
	input \u3_mem_reg[0][14]/NET0131  ;
	input \u3_mem_reg[0][15]/NET0131  ;
	input \u3_mem_reg[0][16]/NET0131  ;
	input \u3_mem_reg[0][17]/NET0131  ;
	input \u3_mem_reg[0][18]/NET0131  ;
	input \u3_mem_reg[0][19]/NET0131  ;
	input \u3_mem_reg[0][1]/NET0131  ;
	input \u3_mem_reg[0][20]/NET0131  ;
	input \u3_mem_reg[0][21]/NET0131  ;
	input \u3_mem_reg[0][22]/NET0131  ;
	input \u3_mem_reg[0][23]/NET0131  ;
	input \u3_mem_reg[0][24]/NET0131  ;
	input \u3_mem_reg[0][25]/NET0131  ;
	input \u3_mem_reg[0][26]/NET0131  ;
	input \u3_mem_reg[0][27]/NET0131  ;
	input \u3_mem_reg[0][28]/NET0131  ;
	input \u3_mem_reg[0][29]/NET0131  ;
	input \u3_mem_reg[0][2]/NET0131  ;
	input \u3_mem_reg[0][30]/NET0131  ;
	input \u3_mem_reg[0][31]/NET0131  ;
	input \u3_mem_reg[0][3]/NET0131  ;
	input \u3_mem_reg[0][4]/NET0131  ;
	input \u3_mem_reg[0][5]/NET0131  ;
	input \u3_mem_reg[0][6]/NET0131  ;
	input \u3_mem_reg[0][7]/NET0131  ;
	input \u3_mem_reg[0][8]/NET0131  ;
	input \u3_mem_reg[0][9]/NET0131  ;
	input \u3_mem_reg[1][0]/NET0131  ;
	input \u3_mem_reg[1][10]/NET0131  ;
	input \u3_mem_reg[1][11]/NET0131  ;
	input \u3_mem_reg[1][12]/NET0131  ;
	input \u3_mem_reg[1][13]/NET0131  ;
	input \u3_mem_reg[1][14]/NET0131  ;
	input \u3_mem_reg[1][15]/NET0131  ;
	input \u3_mem_reg[1][16]/NET0131  ;
	input \u3_mem_reg[1][17]/NET0131  ;
	input \u3_mem_reg[1][18]/NET0131  ;
	input \u3_mem_reg[1][19]/NET0131  ;
	input \u3_mem_reg[1][1]/NET0131  ;
	input \u3_mem_reg[1][20]/NET0131  ;
	input \u3_mem_reg[1][21]/NET0131  ;
	input \u3_mem_reg[1][22]/NET0131  ;
	input \u3_mem_reg[1][23]/NET0131  ;
	input \u3_mem_reg[1][24]/NET0131  ;
	input \u3_mem_reg[1][25]/NET0131  ;
	input \u3_mem_reg[1][26]/NET0131  ;
	input \u3_mem_reg[1][27]/NET0131  ;
	input \u3_mem_reg[1][28]/NET0131  ;
	input \u3_mem_reg[1][29]/NET0131  ;
	input \u3_mem_reg[1][2]/NET0131  ;
	input \u3_mem_reg[1][30]/NET0131  ;
	input \u3_mem_reg[1][31]/NET0131  ;
	input \u3_mem_reg[1][3]/NET0131  ;
	input \u3_mem_reg[1][4]/NET0131  ;
	input \u3_mem_reg[1][5]/NET0131  ;
	input \u3_mem_reg[1][6]/NET0131  ;
	input \u3_mem_reg[1][7]/NET0131  ;
	input \u3_mem_reg[1][8]/NET0131  ;
	input \u3_mem_reg[1][9]/NET0131  ;
	input \u3_mem_reg[2][0]/NET0131  ;
	input \u3_mem_reg[2][10]/NET0131  ;
	input \u3_mem_reg[2][11]/NET0131  ;
	input \u3_mem_reg[2][12]/NET0131  ;
	input \u3_mem_reg[2][13]/NET0131  ;
	input \u3_mem_reg[2][14]/NET0131  ;
	input \u3_mem_reg[2][15]/NET0131  ;
	input \u3_mem_reg[2][16]/NET0131  ;
	input \u3_mem_reg[2][17]/NET0131  ;
	input \u3_mem_reg[2][18]/NET0131  ;
	input \u3_mem_reg[2][19]/NET0131  ;
	input \u3_mem_reg[2][1]/NET0131  ;
	input \u3_mem_reg[2][20]/NET0131  ;
	input \u3_mem_reg[2][21]/NET0131  ;
	input \u3_mem_reg[2][22]/NET0131  ;
	input \u3_mem_reg[2][23]/NET0131  ;
	input \u3_mem_reg[2][24]/NET0131  ;
	input \u3_mem_reg[2][25]/NET0131  ;
	input \u3_mem_reg[2][26]/NET0131  ;
	input \u3_mem_reg[2][27]/NET0131  ;
	input \u3_mem_reg[2][28]/NET0131  ;
	input \u3_mem_reg[2][29]/NET0131  ;
	input \u3_mem_reg[2][2]/NET0131  ;
	input \u3_mem_reg[2][30]/NET0131  ;
	input \u3_mem_reg[2][31]/NET0131  ;
	input \u3_mem_reg[2][3]/NET0131  ;
	input \u3_mem_reg[2][4]/NET0131  ;
	input \u3_mem_reg[2][5]/NET0131  ;
	input \u3_mem_reg[2][6]/NET0131  ;
	input \u3_mem_reg[2][7]/NET0131  ;
	input \u3_mem_reg[2][8]/NET0131  ;
	input \u3_mem_reg[2][9]/NET0131  ;
	input \u3_mem_reg[3][0]/NET0131  ;
	input \u3_mem_reg[3][10]/NET0131  ;
	input \u3_mem_reg[3][11]/NET0131  ;
	input \u3_mem_reg[3][12]/NET0131  ;
	input \u3_mem_reg[3][13]/NET0131  ;
	input \u3_mem_reg[3][14]/NET0131  ;
	input \u3_mem_reg[3][15]/NET0131  ;
	input \u3_mem_reg[3][16]/NET0131  ;
	input \u3_mem_reg[3][17]/NET0131  ;
	input \u3_mem_reg[3][18]/NET0131  ;
	input \u3_mem_reg[3][19]/NET0131  ;
	input \u3_mem_reg[3][1]/NET0131  ;
	input \u3_mem_reg[3][20]/NET0131  ;
	input \u3_mem_reg[3][21]/NET0131  ;
	input \u3_mem_reg[3][22]/NET0131  ;
	input \u3_mem_reg[3][23]/NET0131  ;
	input \u3_mem_reg[3][24]/NET0131  ;
	input \u3_mem_reg[3][25]/NET0131  ;
	input \u3_mem_reg[3][26]/NET0131  ;
	input \u3_mem_reg[3][27]/NET0131  ;
	input \u3_mem_reg[3][28]/NET0131  ;
	input \u3_mem_reg[3][29]/NET0131  ;
	input \u3_mem_reg[3][2]/NET0131  ;
	input \u3_mem_reg[3][30]/NET0131  ;
	input \u3_mem_reg[3][31]/NET0131  ;
	input \u3_mem_reg[3][3]/NET0131  ;
	input \u3_mem_reg[3][4]/NET0131  ;
	input \u3_mem_reg[3][5]/NET0131  ;
	input \u3_mem_reg[3][6]/NET0131  ;
	input \u3_mem_reg[3][7]/NET0131  ;
	input \u3_mem_reg[3][8]/NET0131  ;
	input \u3_mem_reg[3][9]/NET0131  ;
	input \u3_rp_reg[0]/P0001  ;
	input \u3_rp_reg[1]/NET0131  ;
	input \u3_rp_reg[2]/NET0131  ;
	input \u3_rp_reg[3]/NET0131  ;
	input \u3_status_reg[0]/P0001  ;
	input \u3_status_reg[1]/P0001  ;
	input \u3_wp_reg[0]/P0001  ;
	input \u3_wp_reg[1]/NET0131  ;
	input \u3_wp_reg[2]/P0001  ;
	input \u4_dout_reg[0]/P0001  ;
	input \u4_dout_reg[10]/P0001  ;
	input \u4_dout_reg[11]/P0001  ;
	input \u4_dout_reg[12]/P0001  ;
	input \u4_dout_reg[13]/P0001  ;
	input \u4_dout_reg[14]/P0001  ;
	input \u4_dout_reg[15]/P0001  ;
	input \u4_dout_reg[16]/P0001  ;
	input \u4_dout_reg[17]/P0001  ;
	input \u4_dout_reg[18]/P0001  ;
	input \u4_dout_reg[19]/P0001  ;
	input \u4_dout_reg[1]/P0001  ;
	input \u4_dout_reg[2]/P0001  ;
	input \u4_dout_reg[3]/P0001  ;
	input \u4_dout_reg[4]/P0001  ;
	input \u4_dout_reg[5]/P0001  ;
	input \u4_dout_reg[6]/P0001  ;
	input \u4_dout_reg[7]/P0001  ;
	input \u4_dout_reg[8]/P0001  ;
	input \u4_dout_reg[9]/P0001  ;
	input \u4_empty_reg/NET0131  ;
	input \u4_mem_reg[0][0]/NET0131  ;
	input \u4_mem_reg[0][10]/NET0131  ;
	input \u4_mem_reg[0][11]/NET0131  ;
	input \u4_mem_reg[0][12]/NET0131  ;
	input \u4_mem_reg[0][13]/NET0131  ;
	input \u4_mem_reg[0][14]/NET0131  ;
	input \u4_mem_reg[0][15]/NET0131  ;
	input \u4_mem_reg[0][16]/NET0131  ;
	input \u4_mem_reg[0][17]/NET0131  ;
	input \u4_mem_reg[0][18]/NET0131  ;
	input \u4_mem_reg[0][19]/NET0131  ;
	input \u4_mem_reg[0][1]/NET0131  ;
	input \u4_mem_reg[0][20]/NET0131  ;
	input \u4_mem_reg[0][21]/NET0131  ;
	input \u4_mem_reg[0][22]/NET0131  ;
	input \u4_mem_reg[0][23]/NET0131  ;
	input \u4_mem_reg[0][24]/NET0131  ;
	input \u4_mem_reg[0][25]/NET0131  ;
	input \u4_mem_reg[0][26]/NET0131  ;
	input \u4_mem_reg[0][27]/NET0131  ;
	input \u4_mem_reg[0][28]/NET0131  ;
	input \u4_mem_reg[0][29]/NET0131  ;
	input \u4_mem_reg[0][2]/NET0131  ;
	input \u4_mem_reg[0][30]/NET0131  ;
	input \u4_mem_reg[0][31]/NET0131  ;
	input \u4_mem_reg[0][3]/NET0131  ;
	input \u4_mem_reg[0][4]/NET0131  ;
	input \u4_mem_reg[0][5]/NET0131  ;
	input \u4_mem_reg[0][6]/NET0131  ;
	input \u4_mem_reg[0][7]/NET0131  ;
	input \u4_mem_reg[0][8]/NET0131  ;
	input \u4_mem_reg[0][9]/NET0131  ;
	input \u4_mem_reg[1][0]/NET0131  ;
	input \u4_mem_reg[1][10]/NET0131  ;
	input \u4_mem_reg[1][11]/NET0131  ;
	input \u4_mem_reg[1][12]/NET0131  ;
	input \u4_mem_reg[1][13]/NET0131  ;
	input \u4_mem_reg[1][14]/NET0131  ;
	input \u4_mem_reg[1][15]/NET0131  ;
	input \u4_mem_reg[1][16]/NET0131  ;
	input \u4_mem_reg[1][17]/NET0131  ;
	input \u4_mem_reg[1][18]/NET0131  ;
	input \u4_mem_reg[1][19]/NET0131  ;
	input \u4_mem_reg[1][1]/NET0131  ;
	input \u4_mem_reg[1][20]/NET0131  ;
	input \u4_mem_reg[1][21]/NET0131  ;
	input \u4_mem_reg[1][22]/NET0131  ;
	input \u4_mem_reg[1][23]/NET0131  ;
	input \u4_mem_reg[1][24]/NET0131  ;
	input \u4_mem_reg[1][25]/NET0131  ;
	input \u4_mem_reg[1][26]/NET0131  ;
	input \u4_mem_reg[1][27]/NET0131  ;
	input \u4_mem_reg[1][28]/NET0131  ;
	input \u4_mem_reg[1][29]/NET0131  ;
	input \u4_mem_reg[1][2]/NET0131  ;
	input \u4_mem_reg[1][30]/NET0131  ;
	input \u4_mem_reg[1][31]/NET0131  ;
	input \u4_mem_reg[1][3]/NET0131  ;
	input \u4_mem_reg[1][4]/NET0131  ;
	input \u4_mem_reg[1][5]/NET0131  ;
	input \u4_mem_reg[1][6]/NET0131  ;
	input \u4_mem_reg[1][7]/NET0131  ;
	input \u4_mem_reg[1][8]/NET0131  ;
	input \u4_mem_reg[1][9]/NET0131  ;
	input \u4_mem_reg[2][0]/NET0131  ;
	input \u4_mem_reg[2][10]/NET0131  ;
	input \u4_mem_reg[2][11]/NET0131  ;
	input \u4_mem_reg[2][12]/NET0131  ;
	input \u4_mem_reg[2][13]/NET0131  ;
	input \u4_mem_reg[2][14]/NET0131  ;
	input \u4_mem_reg[2][15]/NET0131  ;
	input \u4_mem_reg[2][16]/NET0131  ;
	input \u4_mem_reg[2][17]/NET0131  ;
	input \u4_mem_reg[2][18]/NET0131  ;
	input \u4_mem_reg[2][19]/NET0131  ;
	input \u4_mem_reg[2][1]/NET0131  ;
	input \u4_mem_reg[2][20]/NET0131  ;
	input \u4_mem_reg[2][21]/NET0131  ;
	input \u4_mem_reg[2][22]/NET0131  ;
	input \u4_mem_reg[2][23]/NET0131  ;
	input \u4_mem_reg[2][24]/NET0131  ;
	input \u4_mem_reg[2][25]/NET0131  ;
	input \u4_mem_reg[2][26]/NET0131  ;
	input \u4_mem_reg[2][27]/NET0131  ;
	input \u4_mem_reg[2][28]/NET0131  ;
	input \u4_mem_reg[2][29]/NET0131  ;
	input \u4_mem_reg[2][2]/NET0131  ;
	input \u4_mem_reg[2][30]/NET0131  ;
	input \u4_mem_reg[2][31]/NET0131  ;
	input \u4_mem_reg[2][3]/NET0131  ;
	input \u4_mem_reg[2][4]/NET0131  ;
	input \u4_mem_reg[2][5]/NET0131  ;
	input \u4_mem_reg[2][6]/NET0131  ;
	input \u4_mem_reg[2][7]/NET0131  ;
	input \u4_mem_reg[2][8]/NET0131  ;
	input \u4_mem_reg[2][9]/NET0131  ;
	input \u4_mem_reg[3][0]/NET0131  ;
	input \u4_mem_reg[3][10]/NET0131  ;
	input \u4_mem_reg[3][11]/NET0131  ;
	input \u4_mem_reg[3][12]/NET0131  ;
	input \u4_mem_reg[3][13]/NET0131  ;
	input \u4_mem_reg[3][14]/NET0131  ;
	input \u4_mem_reg[3][15]/NET0131  ;
	input \u4_mem_reg[3][16]/NET0131  ;
	input \u4_mem_reg[3][17]/NET0131  ;
	input \u4_mem_reg[3][18]/NET0131  ;
	input \u4_mem_reg[3][19]/NET0131  ;
	input \u4_mem_reg[3][1]/NET0131  ;
	input \u4_mem_reg[3][20]/NET0131  ;
	input \u4_mem_reg[3][21]/NET0131  ;
	input \u4_mem_reg[3][22]/NET0131  ;
	input \u4_mem_reg[3][23]/NET0131  ;
	input \u4_mem_reg[3][24]/NET0131  ;
	input \u4_mem_reg[3][25]/NET0131  ;
	input \u4_mem_reg[3][26]/NET0131  ;
	input \u4_mem_reg[3][27]/NET0131  ;
	input \u4_mem_reg[3][28]/NET0131  ;
	input \u4_mem_reg[3][29]/NET0131  ;
	input \u4_mem_reg[3][2]/NET0131  ;
	input \u4_mem_reg[3][30]/NET0131  ;
	input \u4_mem_reg[3][31]/NET0131  ;
	input \u4_mem_reg[3][3]/NET0131  ;
	input \u4_mem_reg[3][4]/NET0131  ;
	input \u4_mem_reg[3][5]/NET0131  ;
	input \u4_mem_reg[3][6]/NET0131  ;
	input \u4_mem_reg[3][7]/NET0131  ;
	input \u4_mem_reg[3][8]/NET0131  ;
	input \u4_mem_reg[3][9]/NET0131  ;
	input \u4_rp_reg[0]/P0001  ;
	input \u4_rp_reg[1]/NET0131  ;
	input \u4_rp_reg[2]/NET0131  ;
	input \u4_rp_reg[3]/NET0131  ;
	input \u4_status_reg[0]/P0001  ;
	input \u4_status_reg[1]/P0001  ;
	input \u4_wp_reg[0]/P0001  ;
	input \u4_wp_reg[1]/NET0131  ;
	input \u4_wp_reg[2]/P0001  ;
	input \u5_dout_reg[0]/P0001  ;
	input \u5_dout_reg[10]/P0001  ;
	input \u5_dout_reg[11]/P0001  ;
	input \u5_dout_reg[12]/P0001  ;
	input \u5_dout_reg[13]/P0001  ;
	input \u5_dout_reg[14]/P0001  ;
	input \u5_dout_reg[15]/P0001  ;
	input \u5_dout_reg[16]/P0001  ;
	input \u5_dout_reg[17]/P0001  ;
	input \u5_dout_reg[18]/P0001  ;
	input \u5_dout_reg[19]/P0001  ;
	input \u5_dout_reg[1]/P0001  ;
	input \u5_dout_reg[2]/P0001  ;
	input \u5_dout_reg[3]/P0001  ;
	input \u5_dout_reg[4]/P0001  ;
	input \u5_dout_reg[5]/P0001  ;
	input \u5_dout_reg[6]/P0001  ;
	input \u5_dout_reg[7]/P0001  ;
	input \u5_dout_reg[8]/P0001  ;
	input \u5_dout_reg[9]/P0001  ;
	input \u5_empty_reg/NET0131  ;
	input \u5_mem_reg[0][0]/NET0131  ;
	input \u5_mem_reg[0][10]/NET0131  ;
	input \u5_mem_reg[0][11]/NET0131  ;
	input \u5_mem_reg[0][12]/NET0131  ;
	input \u5_mem_reg[0][13]/NET0131  ;
	input \u5_mem_reg[0][14]/NET0131  ;
	input \u5_mem_reg[0][15]/NET0131  ;
	input \u5_mem_reg[0][16]/NET0131  ;
	input \u5_mem_reg[0][17]/NET0131  ;
	input \u5_mem_reg[0][18]/NET0131  ;
	input \u5_mem_reg[0][19]/NET0131  ;
	input \u5_mem_reg[0][1]/NET0131  ;
	input \u5_mem_reg[0][20]/NET0131  ;
	input \u5_mem_reg[0][21]/NET0131  ;
	input \u5_mem_reg[0][22]/NET0131  ;
	input \u5_mem_reg[0][23]/NET0131  ;
	input \u5_mem_reg[0][24]/NET0131  ;
	input \u5_mem_reg[0][25]/NET0131  ;
	input \u5_mem_reg[0][26]/NET0131  ;
	input \u5_mem_reg[0][27]/NET0131  ;
	input \u5_mem_reg[0][28]/NET0131  ;
	input \u5_mem_reg[0][29]/NET0131  ;
	input \u5_mem_reg[0][2]/NET0131  ;
	input \u5_mem_reg[0][30]/NET0131  ;
	input \u5_mem_reg[0][31]/NET0131  ;
	input \u5_mem_reg[0][3]/NET0131  ;
	input \u5_mem_reg[0][4]/NET0131  ;
	input \u5_mem_reg[0][5]/NET0131  ;
	input \u5_mem_reg[0][6]/NET0131  ;
	input \u5_mem_reg[0][7]/NET0131  ;
	input \u5_mem_reg[0][8]/NET0131  ;
	input \u5_mem_reg[0][9]/NET0131  ;
	input \u5_mem_reg[1][0]/NET0131  ;
	input \u5_mem_reg[1][10]/NET0131  ;
	input \u5_mem_reg[1][11]/NET0131  ;
	input \u5_mem_reg[1][12]/NET0131  ;
	input \u5_mem_reg[1][13]/NET0131  ;
	input \u5_mem_reg[1][14]/NET0131  ;
	input \u5_mem_reg[1][15]/NET0131  ;
	input \u5_mem_reg[1][16]/NET0131  ;
	input \u5_mem_reg[1][17]/NET0131  ;
	input \u5_mem_reg[1][18]/NET0131  ;
	input \u5_mem_reg[1][19]/NET0131  ;
	input \u5_mem_reg[1][1]/NET0131  ;
	input \u5_mem_reg[1][20]/NET0131  ;
	input \u5_mem_reg[1][21]/NET0131  ;
	input \u5_mem_reg[1][22]/NET0131  ;
	input \u5_mem_reg[1][23]/NET0131  ;
	input \u5_mem_reg[1][24]/NET0131  ;
	input \u5_mem_reg[1][25]/NET0131  ;
	input \u5_mem_reg[1][26]/NET0131  ;
	input \u5_mem_reg[1][27]/NET0131  ;
	input \u5_mem_reg[1][28]/NET0131  ;
	input \u5_mem_reg[1][29]/NET0131  ;
	input \u5_mem_reg[1][2]/NET0131  ;
	input \u5_mem_reg[1][30]/NET0131  ;
	input \u5_mem_reg[1][31]/NET0131  ;
	input \u5_mem_reg[1][3]/NET0131  ;
	input \u5_mem_reg[1][4]/NET0131  ;
	input \u5_mem_reg[1][5]/NET0131  ;
	input \u5_mem_reg[1][6]/NET0131  ;
	input \u5_mem_reg[1][7]/NET0131  ;
	input \u5_mem_reg[1][8]/NET0131  ;
	input \u5_mem_reg[1][9]/NET0131  ;
	input \u5_mem_reg[2][0]/NET0131  ;
	input \u5_mem_reg[2][10]/NET0131  ;
	input \u5_mem_reg[2][11]/NET0131  ;
	input \u5_mem_reg[2][12]/NET0131  ;
	input \u5_mem_reg[2][13]/NET0131  ;
	input \u5_mem_reg[2][14]/NET0131  ;
	input \u5_mem_reg[2][15]/NET0131  ;
	input \u5_mem_reg[2][16]/NET0131  ;
	input \u5_mem_reg[2][17]/NET0131  ;
	input \u5_mem_reg[2][18]/NET0131  ;
	input \u5_mem_reg[2][19]/NET0131  ;
	input \u5_mem_reg[2][1]/NET0131  ;
	input \u5_mem_reg[2][20]/NET0131  ;
	input \u5_mem_reg[2][21]/NET0131  ;
	input \u5_mem_reg[2][22]/NET0131  ;
	input \u5_mem_reg[2][23]/NET0131  ;
	input \u5_mem_reg[2][24]/NET0131  ;
	input \u5_mem_reg[2][25]/NET0131  ;
	input \u5_mem_reg[2][26]/NET0131  ;
	input \u5_mem_reg[2][27]/NET0131  ;
	input \u5_mem_reg[2][28]/NET0131  ;
	input \u5_mem_reg[2][29]/NET0131  ;
	input \u5_mem_reg[2][2]/NET0131  ;
	input \u5_mem_reg[2][30]/NET0131  ;
	input \u5_mem_reg[2][31]/NET0131  ;
	input \u5_mem_reg[2][3]/NET0131  ;
	input \u5_mem_reg[2][4]/NET0131  ;
	input \u5_mem_reg[2][5]/NET0131  ;
	input \u5_mem_reg[2][6]/NET0131  ;
	input \u5_mem_reg[2][7]/NET0131  ;
	input \u5_mem_reg[2][8]/NET0131  ;
	input \u5_mem_reg[2][9]/NET0131  ;
	input \u5_mem_reg[3][0]/NET0131  ;
	input \u5_mem_reg[3][10]/NET0131  ;
	input \u5_mem_reg[3][11]/NET0131  ;
	input \u5_mem_reg[3][12]/NET0131  ;
	input \u5_mem_reg[3][13]/NET0131  ;
	input \u5_mem_reg[3][14]/NET0131  ;
	input \u5_mem_reg[3][15]/NET0131  ;
	input \u5_mem_reg[3][16]/NET0131  ;
	input \u5_mem_reg[3][17]/NET0131  ;
	input \u5_mem_reg[3][18]/NET0131  ;
	input \u5_mem_reg[3][19]/NET0131  ;
	input \u5_mem_reg[3][1]/NET0131  ;
	input \u5_mem_reg[3][20]/NET0131  ;
	input \u5_mem_reg[3][21]/NET0131  ;
	input \u5_mem_reg[3][22]/NET0131  ;
	input \u5_mem_reg[3][23]/NET0131  ;
	input \u5_mem_reg[3][24]/NET0131  ;
	input \u5_mem_reg[3][25]/NET0131  ;
	input \u5_mem_reg[3][26]/NET0131  ;
	input \u5_mem_reg[3][27]/NET0131  ;
	input \u5_mem_reg[3][28]/NET0131  ;
	input \u5_mem_reg[3][29]/NET0131  ;
	input \u5_mem_reg[3][2]/NET0131  ;
	input \u5_mem_reg[3][30]/NET0131  ;
	input \u5_mem_reg[3][31]/NET0131  ;
	input \u5_mem_reg[3][3]/NET0131  ;
	input \u5_mem_reg[3][4]/NET0131  ;
	input \u5_mem_reg[3][5]/NET0131  ;
	input \u5_mem_reg[3][6]/NET0131  ;
	input \u5_mem_reg[3][7]/NET0131  ;
	input \u5_mem_reg[3][8]/NET0131  ;
	input \u5_mem_reg[3][9]/NET0131  ;
	input \u5_rp_reg[0]/P0001  ;
	input \u5_rp_reg[1]/NET0131  ;
	input \u5_rp_reg[2]/NET0131  ;
	input \u5_rp_reg[3]/NET0131  ;
	input \u5_status_reg[0]/P0001  ;
	input \u5_status_reg[1]/P0001  ;
	input \u5_wp_reg[0]/P0001  ;
	input \u5_wp_reg[1]/NET0131  ;
	input \u5_wp_reg[2]/P0001  ;
	input \u6_dout_reg[0]/P0001  ;
	input \u6_dout_reg[10]/P0001  ;
	input \u6_dout_reg[11]/P0001  ;
	input \u6_dout_reg[12]/P0001  ;
	input \u6_dout_reg[13]/P0001  ;
	input \u6_dout_reg[14]/P0001  ;
	input \u6_dout_reg[15]/P0001  ;
	input \u6_dout_reg[16]/P0001  ;
	input \u6_dout_reg[17]/P0001  ;
	input \u6_dout_reg[18]/P0001  ;
	input \u6_dout_reg[19]/P0001  ;
	input \u6_dout_reg[1]/P0001  ;
	input \u6_dout_reg[2]/P0001  ;
	input \u6_dout_reg[3]/P0001  ;
	input \u6_dout_reg[4]/P0001  ;
	input \u6_dout_reg[5]/P0001  ;
	input \u6_dout_reg[6]/P0001  ;
	input \u6_dout_reg[7]/P0001  ;
	input \u6_dout_reg[8]/P0001  ;
	input \u6_dout_reg[9]/P0001  ;
	input \u6_empty_reg/NET0131  ;
	input \u6_mem_reg[0][0]/NET0131  ;
	input \u6_mem_reg[0][10]/NET0131  ;
	input \u6_mem_reg[0][11]/NET0131  ;
	input \u6_mem_reg[0][12]/NET0131  ;
	input \u6_mem_reg[0][13]/NET0131  ;
	input \u6_mem_reg[0][14]/NET0131  ;
	input \u6_mem_reg[0][15]/NET0131  ;
	input \u6_mem_reg[0][16]/NET0131  ;
	input \u6_mem_reg[0][17]/NET0131  ;
	input \u6_mem_reg[0][18]/NET0131  ;
	input \u6_mem_reg[0][19]/NET0131  ;
	input \u6_mem_reg[0][1]/NET0131  ;
	input \u6_mem_reg[0][20]/NET0131  ;
	input \u6_mem_reg[0][21]/NET0131  ;
	input \u6_mem_reg[0][22]/NET0131  ;
	input \u6_mem_reg[0][23]/NET0131  ;
	input \u6_mem_reg[0][24]/NET0131  ;
	input \u6_mem_reg[0][25]/NET0131  ;
	input \u6_mem_reg[0][26]/NET0131  ;
	input \u6_mem_reg[0][27]/NET0131  ;
	input \u6_mem_reg[0][28]/NET0131  ;
	input \u6_mem_reg[0][29]/NET0131  ;
	input \u6_mem_reg[0][2]/NET0131  ;
	input \u6_mem_reg[0][30]/NET0131  ;
	input \u6_mem_reg[0][31]/NET0131  ;
	input \u6_mem_reg[0][3]/NET0131  ;
	input \u6_mem_reg[0][4]/NET0131  ;
	input \u6_mem_reg[0][5]/NET0131  ;
	input \u6_mem_reg[0][6]/NET0131  ;
	input \u6_mem_reg[0][7]/NET0131  ;
	input \u6_mem_reg[0][8]/NET0131  ;
	input \u6_mem_reg[0][9]/NET0131  ;
	input \u6_mem_reg[1][0]/NET0131  ;
	input \u6_mem_reg[1][10]/NET0131  ;
	input \u6_mem_reg[1][11]/NET0131  ;
	input \u6_mem_reg[1][12]/NET0131  ;
	input \u6_mem_reg[1][13]/NET0131  ;
	input \u6_mem_reg[1][14]/NET0131  ;
	input \u6_mem_reg[1][15]/NET0131  ;
	input \u6_mem_reg[1][16]/NET0131  ;
	input \u6_mem_reg[1][17]/NET0131  ;
	input \u6_mem_reg[1][18]/NET0131  ;
	input \u6_mem_reg[1][19]/NET0131  ;
	input \u6_mem_reg[1][1]/NET0131  ;
	input \u6_mem_reg[1][20]/NET0131  ;
	input \u6_mem_reg[1][21]/NET0131  ;
	input \u6_mem_reg[1][22]/NET0131  ;
	input \u6_mem_reg[1][23]/NET0131  ;
	input \u6_mem_reg[1][24]/NET0131  ;
	input \u6_mem_reg[1][25]/NET0131  ;
	input \u6_mem_reg[1][26]/NET0131  ;
	input \u6_mem_reg[1][27]/NET0131  ;
	input \u6_mem_reg[1][28]/NET0131  ;
	input \u6_mem_reg[1][29]/NET0131  ;
	input \u6_mem_reg[1][2]/NET0131  ;
	input \u6_mem_reg[1][30]/NET0131  ;
	input \u6_mem_reg[1][31]/NET0131  ;
	input \u6_mem_reg[1][3]/NET0131  ;
	input \u6_mem_reg[1][4]/NET0131  ;
	input \u6_mem_reg[1][5]/NET0131  ;
	input \u6_mem_reg[1][6]/NET0131  ;
	input \u6_mem_reg[1][7]/NET0131  ;
	input \u6_mem_reg[1][8]/NET0131  ;
	input \u6_mem_reg[1][9]/NET0131  ;
	input \u6_mem_reg[2][0]/NET0131  ;
	input \u6_mem_reg[2][10]/NET0131  ;
	input \u6_mem_reg[2][11]/NET0131  ;
	input \u6_mem_reg[2][12]/NET0131  ;
	input \u6_mem_reg[2][13]/NET0131  ;
	input \u6_mem_reg[2][14]/NET0131  ;
	input \u6_mem_reg[2][15]/NET0131  ;
	input \u6_mem_reg[2][16]/NET0131  ;
	input \u6_mem_reg[2][17]/NET0131  ;
	input \u6_mem_reg[2][18]/NET0131  ;
	input \u6_mem_reg[2][19]/NET0131  ;
	input \u6_mem_reg[2][1]/NET0131  ;
	input \u6_mem_reg[2][20]/NET0131  ;
	input \u6_mem_reg[2][21]/NET0131  ;
	input \u6_mem_reg[2][22]/NET0131  ;
	input \u6_mem_reg[2][23]/NET0131  ;
	input \u6_mem_reg[2][24]/NET0131  ;
	input \u6_mem_reg[2][25]/NET0131  ;
	input \u6_mem_reg[2][26]/NET0131  ;
	input \u6_mem_reg[2][27]/NET0131  ;
	input \u6_mem_reg[2][28]/NET0131  ;
	input \u6_mem_reg[2][29]/NET0131  ;
	input \u6_mem_reg[2][2]/NET0131  ;
	input \u6_mem_reg[2][30]/NET0131  ;
	input \u6_mem_reg[2][31]/NET0131  ;
	input \u6_mem_reg[2][3]/NET0131  ;
	input \u6_mem_reg[2][4]/NET0131  ;
	input \u6_mem_reg[2][5]/NET0131  ;
	input \u6_mem_reg[2][6]/NET0131  ;
	input \u6_mem_reg[2][7]/NET0131  ;
	input \u6_mem_reg[2][8]/NET0131  ;
	input \u6_mem_reg[2][9]/NET0131  ;
	input \u6_mem_reg[3][0]/NET0131  ;
	input \u6_mem_reg[3][10]/NET0131  ;
	input \u6_mem_reg[3][11]/NET0131  ;
	input \u6_mem_reg[3][12]/NET0131  ;
	input \u6_mem_reg[3][13]/NET0131  ;
	input \u6_mem_reg[3][14]/NET0131  ;
	input \u6_mem_reg[3][15]/NET0131  ;
	input \u6_mem_reg[3][16]/NET0131  ;
	input \u6_mem_reg[3][17]/NET0131  ;
	input \u6_mem_reg[3][18]/NET0131  ;
	input \u6_mem_reg[3][19]/NET0131  ;
	input \u6_mem_reg[3][1]/NET0131  ;
	input \u6_mem_reg[3][20]/NET0131  ;
	input \u6_mem_reg[3][21]/NET0131  ;
	input \u6_mem_reg[3][22]/NET0131  ;
	input \u6_mem_reg[3][23]/NET0131  ;
	input \u6_mem_reg[3][24]/NET0131  ;
	input \u6_mem_reg[3][25]/NET0131  ;
	input \u6_mem_reg[3][26]/NET0131  ;
	input \u6_mem_reg[3][27]/NET0131  ;
	input \u6_mem_reg[3][28]/NET0131  ;
	input \u6_mem_reg[3][29]/NET0131  ;
	input \u6_mem_reg[3][2]/NET0131  ;
	input \u6_mem_reg[3][30]/NET0131  ;
	input \u6_mem_reg[3][31]/NET0131  ;
	input \u6_mem_reg[3][3]/NET0131  ;
	input \u6_mem_reg[3][4]/NET0131  ;
	input \u6_mem_reg[3][5]/NET0131  ;
	input \u6_mem_reg[3][6]/NET0131  ;
	input \u6_mem_reg[3][7]/NET0131  ;
	input \u6_mem_reg[3][8]/NET0131  ;
	input \u6_mem_reg[3][9]/NET0131  ;
	input \u6_rp_reg[0]/P0001  ;
	input \u6_rp_reg[1]/NET0131  ;
	input \u6_rp_reg[2]/NET0131  ;
	input \u6_rp_reg[3]/NET0131  ;
	input \u6_status_reg[0]/P0001  ;
	input \u6_status_reg[1]/P0001  ;
	input \u6_wp_reg[0]/P0001  ;
	input \u6_wp_reg[1]/NET0131  ;
	input \u6_wp_reg[2]/P0001  ;
	input \u7_dout_reg[0]/P0001  ;
	input \u7_dout_reg[10]/P0001  ;
	input \u7_dout_reg[11]/P0001  ;
	input \u7_dout_reg[12]/P0001  ;
	input \u7_dout_reg[13]/P0001  ;
	input \u7_dout_reg[14]/P0001  ;
	input \u7_dout_reg[15]/P0001  ;
	input \u7_dout_reg[16]/P0001  ;
	input \u7_dout_reg[17]/P0001  ;
	input \u7_dout_reg[18]/P0001  ;
	input \u7_dout_reg[19]/P0001  ;
	input \u7_dout_reg[1]/P0001  ;
	input \u7_dout_reg[2]/P0001  ;
	input \u7_dout_reg[3]/P0001  ;
	input \u7_dout_reg[4]/P0001  ;
	input \u7_dout_reg[5]/P0001  ;
	input \u7_dout_reg[6]/P0001  ;
	input \u7_dout_reg[7]/P0001  ;
	input \u7_dout_reg[8]/P0001  ;
	input \u7_dout_reg[9]/P0001  ;
	input \u7_empty_reg/NET0131  ;
	input \u7_mem_reg[0][0]/NET0131  ;
	input \u7_mem_reg[0][10]/NET0131  ;
	input \u7_mem_reg[0][11]/NET0131  ;
	input \u7_mem_reg[0][12]/NET0131  ;
	input \u7_mem_reg[0][13]/NET0131  ;
	input \u7_mem_reg[0][14]/NET0131  ;
	input \u7_mem_reg[0][15]/NET0131  ;
	input \u7_mem_reg[0][16]/NET0131  ;
	input \u7_mem_reg[0][17]/NET0131  ;
	input \u7_mem_reg[0][18]/NET0131  ;
	input \u7_mem_reg[0][19]/NET0131  ;
	input \u7_mem_reg[0][1]/NET0131  ;
	input \u7_mem_reg[0][20]/NET0131  ;
	input \u7_mem_reg[0][21]/NET0131  ;
	input \u7_mem_reg[0][22]/NET0131  ;
	input \u7_mem_reg[0][23]/NET0131  ;
	input \u7_mem_reg[0][24]/NET0131  ;
	input \u7_mem_reg[0][25]/NET0131  ;
	input \u7_mem_reg[0][26]/NET0131  ;
	input \u7_mem_reg[0][27]/NET0131  ;
	input \u7_mem_reg[0][28]/NET0131  ;
	input \u7_mem_reg[0][29]/NET0131  ;
	input \u7_mem_reg[0][2]/NET0131  ;
	input \u7_mem_reg[0][30]/NET0131  ;
	input \u7_mem_reg[0][31]/NET0131  ;
	input \u7_mem_reg[0][3]/NET0131  ;
	input \u7_mem_reg[0][4]/NET0131  ;
	input \u7_mem_reg[0][5]/NET0131  ;
	input \u7_mem_reg[0][6]/NET0131  ;
	input \u7_mem_reg[0][7]/NET0131  ;
	input \u7_mem_reg[0][8]/NET0131  ;
	input \u7_mem_reg[0][9]/NET0131  ;
	input \u7_mem_reg[1][0]/NET0131  ;
	input \u7_mem_reg[1][10]/NET0131  ;
	input \u7_mem_reg[1][11]/NET0131  ;
	input \u7_mem_reg[1][12]/NET0131  ;
	input \u7_mem_reg[1][13]/NET0131  ;
	input \u7_mem_reg[1][14]/NET0131  ;
	input \u7_mem_reg[1][15]/NET0131  ;
	input \u7_mem_reg[1][16]/NET0131  ;
	input \u7_mem_reg[1][17]/NET0131  ;
	input \u7_mem_reg[1][18]/NET0131  ;
	input \u7_mem_reg[1][19]/NET0131  ;
	input \u7_mem_reg[1][1]/NET0131  ;
	input \u7_mem_reg[1][20]/NET0131  ;
	input \u7_mem_reg[1][21]/NET0131  ;
	input \u7_mem_reg[1][22]/NET0131  ;
	input \u7_mem_reg[1][23]/NET0131  ;
	input \u7_mem_reg[1][24]/NET0131  ;
	input \u7_mem_reg[1][25]/NET0131  ;
	input \u7_mem_reg[1][26]/NET0131  ;
	input \u7_mem_reg[1][27]/NET0131  ;
	input \u7_mem_reg[1][28]/NET0131  ;
	input \u7_mem_reg[1][29]/NET0131  ;
	input \u7_mem_reg[1][2]/NET0131  ;
	input \u7_mem_reg[1][30]/NET0131  ;
	input \u7_mem_reg[1][31]/NET0131  ;
	input \u7_mem_reg[1][3]/NET0131  ;
	input \u7_mem_reg[1][4]/NET0131  ;
	input \u7_mem_reg[1][5]/NET0131  ;
	input \u7_mem_reg[1][6]/NET0131  ;
	input \u7_mem_reg[1][7]/NET0131  ;
	input \u7_mem_reg[1][8]/NET0131  ;
	input \u7_mem_reg[1][9]/NET0131  ;
	input \u7_mem_reg[2][0]/NET0131  ;
	input \u7_mem_reg[2][10]/NET0131  ;
	input \u7_mem_reg[2][11]/NET0131  ;
	input \u7_mem_reg[2][12]/NET0131  ;
	input \u7_mem_reg[2][13]/NET0131  ;
	input \u7_mem_reg[2][14]/NET0131  ;
	input \u7_mem_reg[2][15]/NET0131  ;
	input \u7_mem_reg[2][16]/NET0131  ;
	input \u7_mem_reg[2][17]/NET0131  ;
	input \u7_mem_reg[2][18]/NET0131  ;
	input \u7_mem_reg[2][19]/NET0131  ;
	input \u7_mem_reg[2][1]/NET0131  ;
	input \u7_mem_reg[2][20]/NET0131  ;
	input \u7_mem_reg[2][21]/NET0131  ;
	input \u7_mem_reg[2][22]/NET0131  ;
	input \u7_mem_reg[2][23]/NET0131  ;
	input \u7_mem_reg[2][24]/NET0131  ;
	input \u7_mem_reg[2][25]/NET0131  ;
	input \u7_mem_reg[2][26]/NET0131  ;
	input \u7_mem_reg[2][27]/NET0131  ;
	input \u7_mem_reg[2][28]/NET0131  ;
	input \u7_mem_reg[2][29]/NET0131  ;
	input \u7_mem_reg[2][2]/NET0131  ;
	input \u7_mem_reg[2][30]/NET0131  ;
	input \u7_mem_reg[2][31]/NET0131  ;
	input \u7_mem_reg[2][3]/NET0131  ;
	input \u7_mem_reg[2][4]/NET0131  ;
	input \u7_mem_reg[2][5]/NET0131  ;
	input \u7_mem_reg[2][6]/NET0131  ;
	input \u7_mem_reg[2][7]/NET0131  ;
	input \u7_mem_reg[2][8]/NET0131  ;
	input \u7_mem_reg[2][9]/NET0131  ;
	input \u7_mem_reg[3][0]/NET0131  ;
	input \u7_mem_reg[3][10]/NET0131  ;
	input \u7_mem_reg[3][11]/NET0131  ;
	input \u7_mem_reg[3][12]/NET0131  ;
	input \u7_mem_reg[3][13]/NET0131  ;
	input \u7_mem_reg[3][14]/NET0131  ;
	input \u7_mem_reg[3][15]/NET0131  ;
	input \u7_mem_reg[3][16]/NET0131  ;
	input \u7_mem_reg[3][17]/NET0131  ;
	input \u7_mem_reg[3][18]/NET0131  ;
	input \u7_mem_reg[3][19]/NET0131  ;
	input \u7_mem_reg[3][1]/NET0131  ;
	input \u7_mem_reg[3][20]/NET0131  ;
	input \u7_mem_reg[3][21]/NET0131  ;
	input \u7_mem_reg[3][22]/NET0131  ;
	input \u7_mem_reg[3][23]/NET0131  ;
	input \u7_mem_reg[3][24]/NET0131  ;
	input \u7_mem_reg[3][25]/NET0131  ;
	input \u7_mem_reg[3][26]/NET0131  ;
	input \u7_mem_reg[3][27]/NET0131  ;
	input \u7_mem_reg[3][28]/NET0131  ;
	input \u7_mem_reg[3][29]/NET0131  ;
	input \u7_mem_reg[3][2]/NET0131  ;
	input \u7_mem_reg[3][30]/NET0131  ;
	input \u7_mem_reg[3][31]/NET0131  ;
	input \u7_mem_reg[3][3]/NET0131  ;
	input \u7_mem_reg[3][4]/NET0131  ;
	input \u7_mem_reg[3][5]/NET0131  ;
	input \u7_mem_reg[3][6]/NET0131  ;
	input \u7_mem_reg[3][7]/NET0131  ;
	input \u7_mem_reg[3][8]/NET0131  ;
	input \u7_mem_reg[3][9]/NET0131  ;
	input \u7_rp_reg[0]/P0001  ;
	input \u7_rp_reg[1]/NET0131  ;
	input \u7_rp_reg[2]/NET0131  ;
	input \u7_rp_reg[3]/NET0131  ;
	input \u7_status_reg[0]/P0001  ;
	input \u7_status_reg[1]/P0001  ;
	input \u7_wp_reg[0]/P0001  ;
	input \u7_wp_reg[1]/NET0131  ;
	input \u7_wp_reg[2]/P0001  ;
	input \u8_dout_reg[0]/P0001  ;
	input \u8_dout_reg[10]/P0001  ;
	input \u8_dout_reg[11]/P0001  ;
	input \u8_dout_reg[12]/P0001  ;
	input \u8_dout_reg[13]/P0001  ;
	input \u8_dout_reg[14]/P0001  ;
	input \u8_dout_reg[15]/P0001  ;
	input \u8_dout_reg[16]/P0001  ;
	input \u8_dout_reg[17]/P0001  ;
	input \u8_dout_reg[18]/P0001  ;
	input \u8_dout_reg[19]/P0001  ;
	input \u8_dout_reg[1]/P0001  ;
	input \u8_dout_reg[2]/P0001  ;
	input \u8_dout_reg[3]/P0001  ;
	input \u8_dout_reg[4]/P0001  ;
	input \u8_dout_reg[5]/P0001  ;
	input \u8_dout_reg[6]/P0001  ;
	input \u8_dout_reg[7]/P0001  ;
	input \u8_dout_reg[8]/P0001  ;
	input \u8_dout_reg[9]/P0001  ;
	input \u8_empty_reg/NET0131  ;
	input \u8_mem_reg[0][0]/NET0131  ;
	input \u8_mem_reg[0][10]/NET0131  ;
	input \u8_mem_reg[0][11]/NET0131  ;
	input \u8_mem_reg[0][12]/NET0131  ;
	input \u8_mem_reg[0][13]/NET0131  ;
	input \u8_mem_reg[0][14]/NET0131  ;
	input \u8_mem_reg[0][15]/NET0131  ;
	input \u8_mem_reg[0][16]/NET0131  ;
	input \u8_mem_reg[0][17]/NET0131  ;
	input \u8_mem_reg[0][18]/NET0131  ;
	input \u8_mem_reg[0][19]/NET0131  ;
	input \u8_mem_reg[0][1]/NET0131  ;
	input \u8_mem_reg[0][20]/NET0131  ;
	input \u8_mem_reg[0][21]/NET0131  ;
	input \u8_mem_reg[0][22]/NET0131  ;
	input \u8_mem_reg[0][23]/NET0131  ;
	input \u8_mem_reg[0][24]/NET0131  ;
	input \u8_mem_reg[0][25]/NET0131  ;
	input \u8_mem_reg[0][26]/NET0131  ;
	input \u8_mem_reg[0][27]/NET0131  ;
	input \u8_mem_reg[0][28]/NET0131  ;
	input \u8_mem_reg[0][29]/NET0131  ;
	input \u8_mem_reg[0][2]/NET0131  ;
	input \u8_mem_reg[0][30]/NET0131  ;
	input \u8_mem_reg[0][31]/NET0131  ;
	input \u8_mem_reg[0][3]/NET0131  ;
	input \u8_mem_reg[0][4]/NET0131  ;
	input \u8_mem_reg[0][5]/NET0131  ;
	input \u8_mem_reg[0][6]/NET0131  ;
	input \u8_mem_reg[0][7]/NET0131  ;
	input \u8_mem_reg[0][8]/NET0131  ;
	input \u8_mem_reg[0][9]/NET0131  ;
	input \u8_mem_reg[1][0]/NET0131  ;
	input \u8_mem_reg[1][10]/NET0131  ;
	input \u8_mem_reg[1][11]/NET0131  ;
	input \u8_mem_reg[1][12]/NET0131  ;
	input \u8_mem_reg[1][13]/NET0131  ;
	input \u8_mem_reg[1][14]/NET0131  ;
	input \u8_mem_reg[1][15]/NET0131  ;
	input \u8_mem_reg[1][16]/NET0131  ;
	input \u8_mem_reg[1][17]/NET0131  ;
	input \u8_mem_reg[1][18]/NET0131  ;
	input \u8_mem_reg[1][19]/NET0131  ;
	input \u8_mem_reg[1][1]/NET0131  ;
	input \u8_mem_reg[1][20]/NET0131  ;
	input \u8_mem_reg[1][21]/NET0131  ;
	input \u8_mem_reg[1][22]/NET0131  ;
	input \u8_mem_reg[1][23]/NET0131  ;
	input \u8_mem_reg[1][24]/NET0131  ;
	input \u8_mem_reg[1][25]/NET0131  ;
	input \u8_mem_reg[1][26]/NET0131  ;
	input \u8_mem_reg[1][27]/NET0131  ;
	input \u8_mem_reg[1][28]/NET0131  ;
	input \u8_mem_reg[1][29]/NET0131  ;
	input \u8_mem_reg[1][2]/NET0131  ;
	input \u8_mem_reg[1][30]/NET0131  ;
	input \u8_mem_reg[1][31]/NET0131  ;
	input \u8_mem_reg[1][3]/NET0131  ;
	input \u8_mem_reg[1][4]/NET0131  ;
	input \u8_mem_reg[1][5]/NET0131  ;
	input \u8_mem_reg[1][6]/NET0131  ;
	input \u8_mem_reg[1][7]/NET0131  ;
	input \u8_mem_reg[1][8]/NET0131  ;
	input \u8_mem_reg[1][9]/NET0131  ;
	input \u8_mem_reg[2][0]/NET0131  ;
	input \u8_mem_reg[2][10]/NET0131  ;
	input \u8_mem_reg[2][11]/NET0131  ;
	input \u8_mem_reg[2][12]/NET0131  ;
	input \u8_mem_reg[2][13]/NET0131  ;
	input \u8_mem_reg[2][14]/NET0131  ;
	input \u8_mem_reg[2][15]/NET0131  ;
	input \u8_mem_reg[2][16]/NET0131  ;
	input \u8_mem_reg[2][17]/NET0131  ;
	input \u8_mem_reg[2][18]/NET0131  ;
	input \u8_mem_reg[2][19]/NET0131  ;
	input \u8_mem_reg[2][1]/NET0131  ;
	input \u8_mem_reg[2][20]/NET0131  ;
	input \u8_mem_reg[2][21]/NET0131  ;
	input \u8_mem_reg[2][22]/NET0131  ;
	input \u8_mem_reg[2][23]/NET0131  ;
	input \u8_mem_reg[2][24]/NET0131  ;
	input \u8_mem_reg[2][25]/NET0131  ;
	input \u8_mem_reg[2][26]/NET0131  ;
	input \u8_mem_reg[2][27]/NET0131  ;
	input \u8_mem_reg[2][28]/NET0131  ;
	input \u8_mem_reg[2][29]/NET0131  ;
	input \u8_mem_reg[2][2]/NET0131  ;
	input \u8_mem_reg[2][30]/NET0131  ;
	input \u8_mem_reg[2][31]/NET0131  ;
	input \u8_mem_reg[2][3]/NET0131  ;
	input \u8_mem_reg[2][4]/NET0131  ;
	input \u8_mem_reg[2][5]/NET0131  ;
	input \u8_mem_reg[2][6]/NET0131  ;
	input \u8_mem_reg[2][7]/NET0131  ;
	input \u8_mem_reg[2][8]/NET0131  ;
	input \u8_mem_reg[2][9]/NET0131  ;
	input \u8_mem_reg[3][0]/NET0131  ;
	input \u8_mem_reg[3][10]/NET0131  ;
	input \u8_mem_reg[3][11]/NET0131  ;
	input \u8_mem_reg[3][12]/NET0131  ;
	input \u8_mem_reg[3][13]/NET0131  ;
	input \u8_mem_reg[3][14]/NET0131  ;
	input \u8_mem_reg[3][15]/NET0131  ;
	input \u8_mem_reg[3][16]/NET0131  ;
	input \u8_mem_reg[3][17]/NET0131  ;
	input \u8_mem_reg[3][18]/NET0131  ;
	input \u8_mem_reg[3][19]/NET0131  ;
	input \u8_mem_reg[3][1]/NET0131  ;
	input \u8_mem_reg[3][20]/NET0131  ;
	input \u8_mem_reg[3][21]/NET0131  ;
	input \u8_mem_reg[3][22]/NET0131  ;
	input \u8_mem_reg[3][23]/NET0131  ;
	input \u8_mem_reg[3][24]/NET0131  ;
	input \u8_mem_reg[3][25]/NET0131  ;
	input \u8_mem_reg[3][26]/NET0131  ;
	input \u8_mem_reg[3][27]/NET0131  ;
	input \u8_mem_reg[3][28]/NET0131  ;
	input \u8_mem_reg[3][29]/NET0131  ;
	input \u8_mem_reg[3][2]/NET0131  ;
	input \u8_mem_reg[3][30]/NET0131  ;
	input \u8_mem_reg[3][31]/NET0131  ;
	input \u8_mem_reg[3][3]/NET0131  ;
	input \u8_mem_reg[3][4]/NET0131  ;
	input \u8_mem_reg[3][5]/NET0131  ;
	input \u8_mem_reg[3][6]/NET0131  ;
	input \u8_mem_reg[3][7]/NET0131  ;
	input \u8_mem_reg[3][8]/NET0131  ;
	input \u8_mem_reg[3][9]/NET0131  ;
	input \u8_rp_reg[0]/P0001  ;
	input \u8_rp_reg[1]/NET0131  ;
	input \u8_rp_reg[2]/NET0131  ;
	input \u8_rp_reg[3]/NET0131  ;
	input \u8_status_reg[0]/P0001  ;
	input \u8_status_reg[1]/P0001  ;
	input \u8_wp_reg[0]/P0001  ;
	input \u8_wp_reg[1]/NET0131  ;
	input \u8_wp_reg[2]/P0001  ;
	input \u9_din_tmp1_reg[0]/P0001  ;
	input \u9_din_tmp1_reg[10]/P0001  ;
	input \u9_din_tmp1_reg[11]/P0001  ;
	input \u9_din_tmp1_reg[12]/P0001  ;
	input \u9_din_tmp1_reg[13]/P0001  ;
	input \u9_din_tmp1_reg[14]/P0001  ;
	input \u9_din_tmp1_reg[15]/P0001  ;
	input \u9_din_tmp1_reg[1]/P0001  ;
	input \u9_din_tmp1_reg[2]/P0001  ;
	input \u9_din_tmp1_reg[3]/P0001  ;
	input \u9_din_tmp1_reg[4]/P0001  ;
	input \u9_din_tmp1_reg[5]/P0001  ;
	input \u9_din_tmp1_reg[6]/P0001  ;
	input \u9_din_tmp1_reg[7]/P0001  ;
	input \u9_din_tmp1_reg[8]/P0001  ;
	input \u9_din_tmp1_reg[9]/P0001  ;
	input \u9_dout_reg[0]/P0001  ;
	input \u9_dout_reg[10]/P0001  ;
	input \u9_dout_reg[11]/P0001  ;
	input \u9_dout_reg[12]/P0001  ;
	input \u9_dout_reg[13]/P0001  ;
	input \u9_dout_reg[14]/P0001  ;
	input \u9_dout_reg[15]/P0001  ;
	input \u9_dout_reg[16]/P0001  ;
	input \u9_dout_reg[17]/P0001  ;
	input \u9_dout_reg[18]/P0001  ;
	input \u9_dout_reg[19]/P0001  ;
	input \u9_dout_reg[1]/P0001  ;
	input \u9_dout_reg[20]/P0001  ;
	input \u9_dout_reg[21]/P0001  ;
	input \u9_dout_reg[22]/P0001  ;
	input \u9_dout_reg[23]/P0001  ;
	input \u9_dout_reg[24]/P0001  ;
	input \u9_dout_reg[25]/P0001  ;
	input \u9_dout_reg[26]/P0001  ;
	input \u9_dout_reg[27]/P0001  ;
	input \u9_dout_reg[28]/P0001  ;
	input \u9_dout_reg[29]/P0001  ;
	input \u9_dout_reg[2]/P0001  ;
	input \u9_dout_reg[30]/P0001  ;
	input \u9_dout_reg[31]/P0001  ;
	input \u9_dout_reg[3]/P0001  ;
	input \u9_dout_reg[4]/P0001  ;
	input \u9_dout_reg[5]/P0001  ;
	input \u9_dout_reg[6]/P0001  ;
	input \u9_dout_reg[7]/P0001  ;
	input \u9_dout_reg[8]/P0001  ;
	input \u9_dout_reg[9]/P0001  ;
	input \u9_empty_reg/P0001  ;
	input \u9_full_reg/NET0131  ;
	input \u9_mem_reg[0][0]/P0001  ;
	input \u9_mem_reg[0][10]/P0001  ;
	input \u9_mem_reg[0][11]/P0001  ;
	input \u9_mem_reg[0][12]/P0001  ;
	input \u9_mem_reg[0][13]/P0001  ;
	input \u9_mem_reg[0][14]/P0001  ;
	input \u9_mem_reg[0][15]/P0001  ;
	input \u9_mem_reg[0][16]/P0001  ;
	input \u9_mem_reg[0][17]/P0001  ;
	input \u9_mem_reg[0][18]/P0001  ;
	input \u9_mem_reg[0][19]/P0001  ;
	input \u9_mem_reg[0][1]/P0001  ;
	input \u9_mem_reg[0][20]/P0001  ;
	input \u9_mem_reg[0][21]/P0001  ;
	input \u9_mem_reg[0][22]/P0001  ;
	input \u9_mem_reg[0][23]/P0001  ;
	input \u9_mem_reg[0][24]/P0001  ;
	input \u9_mem_reg[0][25]/P0001  ;
	input \u9_mem_reg[0][26]/P0001  ;
	input \u9_mem_reg[0][27]/P0001  ;
	input \u9_mem_reg[0][28]/P0001  ;
	input \u9_mem_reg[0][29]/P0001  ;
	input \u9_mem_reg[0][2]/P0001  ;
	input \u9_mem_reg[0][30]/P0001  ;
	input \u9_mem_reg[0][31]/P0001  ;
	input \u9_mem_reg[0][3]/P0001  ;
	input \u9_mem_reg[0][4]/P0001  ;
	input \u9_mem_reg[0][5]/P0001  ;
	input \u9_mem_reg[0][6]/P0001  ;
	input \u9_mem_reg[0][7]/P0001  ;
	input \u9_mem_reg[0][8]/P0001  ;
	input \u9_mem_reg[0][9]/P0001  ;
	input \u9_mem_reg[1][0]/P0001  ;
	input \u9_mem_reg[1][10]/P0001  ;
	input \u9_mem_reg[1][11]/P0001  ;
	input \u9_mem_reg[1][12]/P0001  ;
	input \u9_mem_reg[1][13]/P0001  ;
	input \u9_mem_reg[1][14]/P0001  ;
	input \u9_mem_reg[1][15]/P0001  ;
	input \u9_mem_reg[1][16]/P0001  ;
	input \u9_mem_reg[1][17]/P0001  ;
	input \u9_mem_reg[1][18]/P0001  ;
	input \u9_mem_reg[1][19]/P0001  ;
	input \u9_mem_reg[1][1]/P0001  ;
	input \u9_mem_reg[1][20]/P0001  ;
	input \u9_mem_reg[1][21]/P0001  ;
	input \u9_mem_reg[1][22]/P0001  ;
	input \u9_mem_reg[1][23]/P0001  ;
	input \u9_mem_reg[1][24]/P0001  ;
	input \u9_mem_reg[1][25]/P0001  ;
	input \u9_mem_reg[1][26]/P0001  ;
	input \u9_mem_reg[1][27]/P0001  ;
	input \u9_mem_reg[1][28]/P0001  ;
	input \u9_mem_reg[1][29]/P0001  ;
	input \u9_mem_reg[1][2]/P0001  ;
	input \u9_mem_reg[1][30]/P0001  ;
	input \u9_mem_reg[1][31]/P0001  ;
	input \u9_mem_reg[1][3]/P0001  ;
	input \u9_mem_reg[1][4]/P0001  ;
	input \u9_mem_reg[1][5]/P0001  ;
	input \u9_mem_reg[1][6]/P0001  ;
	input \u9_mem_reg[1][7]/P0001  ;
	input \u9_mem_reg[1][8]/P0001  ;
	input \u9_mem_reg[1][9]/P0001  ;
	input \u9_mem_reg[2][0]/P0001  ;
	input \u9_mem_reg[2][10]/P0001  ;
	input \u9_mem_reg[2][11]/P0001  ;
	input \u9_mem_reg[2][12]/P0001  ;
	input \u9_mem_reg[2][13]/P0001  ;
	input \u9_mem_reg[2][14]/P0001  ;
	input \u9_mem_reg[2][15]/P0001  ;
	input \u9_mem_reg[2][16]/P0001  ;
	input \u9_mem_reg[2][17]/P0001  ;
	input \u9_mem_reg[2][18]/P0001  ;
	input \u9_mem_reg[2][19]/P0001  ;
	input \u9_mem_reg[2][1]/P0001  ;
	input \u9_mem_reg[2][20]/P0001  ;
	input \u9_mem_reg[2][21]/P0001  ;
	input \u9_mem_reg[2][22]/P0001  ;
	input \u9_mem_reg[2][23]/P0001  ;
	input \u9_mem_reg[2][24]/P0001  ;
	input \u9_mem_reg[2][25]/P0001  ;
	input \u9_mem_reg[2][26]/P0001  ;
	input \u9_mem_reg[2][27]/P0001  ;
	input \u9_mem_reg[2][28]/P0001  ;
	input \u9_mem_reg[2][29]/P0001  ;
	input \u9_mem_reg[2][2]/P0001  ;
	input \u9_mem_reg[2][30]/P0001  ;
	input \u9_mem_reg[2][31]/P0001  ;
	input \u9_mem_reg[2][3]/P0001  ;
	input \u9_mem_reg[2][4]/P0001  ;
	input \u9_mem_reg[2][5]/P0001  ;
	input \u9_mem_reg[2][6]/P0001  ;
	input \u9_mem_reg[2][7]/P0001  ;
	input \u9_mem_reg[2][8]/P0001  ;
	input \u9_mem_reg[2][9]/P0001  ;
	input \u9_mem_reg[3][0]/P0001  ;
	input \u9_mem_reg[3][10]/P0001  ;
	input \u9_mem_reg[3][11]/P0001  ;
	input \u9_mem_reg[3][12]/P0001  ;
	input \u9_mem_reg[3][13]/P0001  ;
	input \u9_mem_reg[3][14]/P0001  ;
	input \u9_mem_reg[3][15]/P0001  ;
	input \u9_mem_reg[3][16]/P0001  ;
	input \u9_mem_reg[3][17]/P0001  ;
	input \u9_mem_reg[3][18]/P0001  ;
	input \u9_mem_reg[3][19]/P0001  ;
	input \u9_mem_reg[3][1]/P0001  ;
	input \u9_mem_reg[3][20]/P0001  ;
	input \u9_mem_reg[3][21]/P0001  ;
	input \u9_mem_reg[3][22]/P0001  ;
	input \u9_mem_reg[3][23]/P0001  ;
	input \u9_mem_reg[3][24]/P0001  ;
	input \u9_mem_reg[3][25]/P0001  ;
	input \u9_mem_reg[3][26]/P0001  ;
	input \u9_mem_reg[3][27]/P0001  ;
	input \u9_mem_reg[3][28]/P0001  ;
	input \u9_mem_reg[3][29]/P0001  ;
	input \u9_mem_reg[3][2]/P0001  ;
	input \u9_mem_reg[3][30]/P0001  ;
	input \u9_mem_reg[3][31]/P0001  ;
	input \u9_mem_reg[3][3]/P0001  ;
	input \u9_mem_reg[3][4]/P0001  ;
	input \u9_mem_reg[3][5]/P0001  ;
	input \u9_mem_reg[3][6]/P0001  ;
	input \u9_mem_reg[3][7]/P0001  ;
	input \u9_mem_reg[3][8]/P0001  ;
	input \u9_mem_reg[3][9]/P0001  ;
	input \u9_rp_reg[0]/P0001  ;
	input \u9_rp_reg[1]/P0001  ;
	input \u9_rp_reg[2]/P0001  ;
	input \u9_status_reg[0]/P0001  ;
	input \u9_status_reg[1]/P0001  ;
	input \u9_wp_reg[0]/NET0131  ;
	input \u9_wp_reg[1]/P0001  ;
	input \u9_wp_reg[2]/P0001  ;
	input \u9_wp_reg[3]/P0001  ;
	input \valid_s_reg/NET0131  ;
	input wb_ack_o_pad ;
	input \wb_addr_i[29]_pad  ;
	input \wb_addr_i[2]_pad  ;
	input \wb_addr_i[30]_pad  ;
	input \wb_addr_i[31]_pad  ;
	input \wb_addr_i[3]_pad  ;
	input \wb_addr_i[4]_pad  ;
	input \wb_addr_i[5]_pad  ;
	input \wb_addr_i[6]_pad  ;
	input wb_cyc_i_pad ;
	input wb_stb_i_pad ;
	input wb_we_i_pad ;
	output \_al_n1  ;
	output \g16/_0_  ;
	output \g23/_0_  ;
	output \g29500/_0_  ;
	output \g29503/_3_  ;
	output \g29505/_3_  ;
	output \g29507/_3_  ;
	output \g29509/_3_  ;
	output \g29511/_0_  ;
	output \g29513/_3_  ;
	output \g29515/_3_  ;
	output \g29517/_3_  ;
	output \g29519/_0_  ;
	output \g29522/_0_  ;
	output \g29524/_0_  ;
	output \g29526/_0_  ;
	output \g29528/_0_  ;
	output \g29530/_0_  ;
	output \g29532/_0_  ;
	output \g29534/_3_  ;
	output \g29536/_3_  ;
	output \g29538/_3_  ;
	output \g29540/_3_  ;
	output \g29542/_3_  ;
	output \g29544/_3_  ;
	output \g29546/_3_  ;
	output \g29548/_3_  ;
	output \g29550/_0_  ;
	output \g29552/_0_  ;
	output \g29554/_0_  ;
	output \g29556/_0_  ;
	output \g29558/_0_  ;
	output \g29560/_0_  ;
	output \g29562/_0_  ;
	output \g29564/_0_  ;
	output \g29566/_0_  ;
	output \g29568/_0_  ;
	output \g29570/_0_  ;
	output \g29572/_0_  ;
	output \g29574/_3_  ;
	output \g29576/_3_  ;
	output \g29578/_3_  ;
	output \g29580/_3_  ;
	output \g29582/_3_  ;
	output \g29584/_3_  ;
	output \g29586/_3_  ;
	output \g29588/_3_  ;
	output \g29590/_3_  ;
	output \g29592/_3_  ;
	output \g29594/_3_  ;
	output \g29596/_3_  ;
	output \g29598/_3_  ;
	output \g29600/_3_  ;
	output \g29602/_3_  ;
	output \g29604/_3_  ;
	output \g29606/_0_  ;
	output \g29608/_0_  ;
	output \g29610/_0_  ;
	output \g29612/_0_  ;
	output \g29614/_3_  ;
	output \g29616/_3_  ;
	output \g29618/_3_  ;
	output \g29620/_3_  ;
	output \g29622/_3_  ;
	output \g29624/_3_  ;
	output \g29626/_3_  ;
	output \g29628/_3_  ;
	output \g29630/_3_  ;
	output \g29632/_3_  ;
	output \g29634/_3_  ;
	output \g29636/_3_  ;
	output \g29638/_3_  ;
	output \g29640/_3_  ;
	output \g29642/_3_  ;
	output \g29644/_3_  ;
	output \g29646/_3_  ;
	output \g29648/_3_  ;
	output \g29650/_3_  ;
	output \g29652/_3_  ;
	output \g29654/_3_  ;
	output \g29656/_3_  ;
	output \g29658/_3_  ;
	output \g29660/_3_  ;
	output \g29662/_3_  ;
	output \g29664/_3_  ;
	output \g29666/_3_  ;
	output \g29668/_3_  ;
	output \g29670/_3_  ;
	output \g29672/_3_  ;
	output \g29674/_3_  ;
	output \g29676/_3_  ;
	output \g29678/_3_  ;
	output \g29680/_3_  ;
	output \g29682/_3_  ;
	output \g29684/_3_  ;
	output \g29686/_3_  ;
	output \g29688/_3_  ;
	output \g29690/_3_  ;
	output \g29692/_3_  ;
	output \g29694/_0_  ;
	output \g29696/_0_  ;
	output \g29698/_0_  ;
	output \g29700/_0_  ;
	output \g29702/_0_  ;
	output \g29704/_0_  ;
	output \g29706/_0_  ;
	output \g29708/_0_  ;
	output \g29710/_0_  ;
	output \g29712/_0_  ;
	output \g29714/_0_  ;
	output \g29716/_0_  ;
	output \g29718/_0_  ;
	output \g29720/_0_  ;
	output \g29722/_0_  ;
	output \g29724/_0_  ;
	output \g29726/_0_  ;
	output \g29728/_0_  ;
	output \g29730/_0_  ;
	output \g29732/_0_  ;
	output \g29734/_3_  ;
	output \g29736/_3_  ;
	output \g29738/_3_  ;
	output \g29740/_3_  ;
	output \g29742/_3_  ;
	output \g29744/_3_  ;
	output \g29746/_3_  ;
	output \g29748/_3_  ;
	output \g29750/_3_  ;
	output \g29752/_3_  ;
	output \g29754/_3_  ;
	output \g29756/_3_  ;
	output \g29758/_3_  ;
	output \g29760/_3_  ;
	output \g29762/_3_  ;
	output \g29764/_3_  ;
	output \g29766/_3_  ;
	output \g29768/_3_  ;
	output \g29770/_3_  ;
	output \g29772/_3_  ;
	output \g29774/_3_  ;
	output \g29776/_3_  ;
	output \g29778/_3_  ;
	output \g29780/_3_  ;
	output \g29782/_3_  ;
	output \g29784/_3_  ;
	output \g29786/_3_  ;
	output \g29788/_3_  ;
	output \g29790/_3_  ;
	output \g29792/_3_  ;
	output \g29794/_3_  ;
	output \g29796/_3_  ;
	output \g29798/_3_  ;
	output \g29800/_3_  ;
	output \g29802/_3_  ;
	output \g29804/_3_  ;
	output \g29806/_3_  ;
	output \g29808/_3_  ;
	output \g29810/_3_  ;
	output \g29812/_3_  ;
	output \g29814/_3_  ;
	output \g29816/_3_  ;
	output \g29818/_3_  ;
	output \g29820/_3_  ;
	output \g29822/_3_  ;
	output \g29824/_3_  ;
	output \g29826/_3_  ;
	output \g29828/_3_  ;
	output \g29830/_3_  ;
	output \g29832/_3_  ;
	output \g29834/_3_  ;
	output \g29836/_3_  ;
	output \g29838/_3_  ;
	output \g29840/_3_  ;
	output \g29842/_3_  ;
	output \g29844/_3_  ;
	output \g29846/_3_  ;
	output \g29848/_3_  ;
	output \g29850/_3_  ;
	output \g29852/_3_  ;
	output \g29854/_3_  ;
	output \g29856/_3_  ;
	output \g29858/_3_  ;
	output \g29860/_3_  ;
	output \g29862/_3_  ;
	output \g29864/_3_  ;
	output \g29866/_3_  ;
	output \g29868/_3_  ;
	output \g29870/_3_  ;
	output \g29872/_3_  ;
	output \g29874/_3_  ;
	output \g29876/_3_  ;
	output \g29878/_3_  ;
	output \g29880/_3_  ;
	output \g29904/_0_  ;
	output \g29905/_0_  ;
	output \g29906/_0_  ;
	output \g29907/_0_  ;
	output \g29908/_0_  ;
	output \g29909/_0_  ;
	output \g29914/_3_  ;
	output \g29952/_0_  ;
	output \g29953/_0_  ;
	output \g29954/_0_  ;
	output \g29955/_0_  ;
	output \g29956/_0_  ;
	output \g29957/_0_  ;
	output \g29975/_0_  ;
	output \g29976/_0_  ;
	output \g29977/_0_  ;
	output \g29978/_0_  ;
	output \g29979/_0_  ;
	output \g29980/_0_  ;
	output \g29989/_3_  ;
	output \g30020/_0_  ;
	output \g30021/_0_  ;
	output \g30045/_0_  ;
	output \g30046/_0_  ;
	output \g30047/_0_  ;
	output \g30048/_0_  ;
	output \g30049/_0_  ;
	output \g30050/_0_  ;
	output \g30051/_0_  ;
	output \g30052/_0_  ;
	output \g30053/_0_  ;
	output \g30054/_0_  ;
	output \g30062/_0_  ;
	output \g30063/_0_  ;
	output \g30064/_0_  ;
	output \g30065/_0_  ;
	output \g30066/_0_  ;
	output \g30067/_0_  ;
	output \g30068/_0_  ;
	output \g30069/_0_  ;
	output \g30070/_0_  ;
	output \g30071/_0_  ;
	output \g30072/_0_  ;
	output \g30073/_0_  ;
	output \g30074/_0_  ;
	output \g30075/_0_  ;
	output \g30136/_3_  ;
	output \g30707/_0_  ;
	output \g30708/_0_  ;
	output \g30711/_0_  ;
	output \g30714/_0_  ;
	output \g30715/_0_  ;
	output \g30720/_0_  ;
	output \g30725/_0_  ;
	output \g30741/_0_  ;
	output \g30742/_0_  ;
	output \g30743/_0_  ;
	output \g30744/_0_  ;
	output \g30745/_0_  ;
	output \g30746/_0_  ;
	output \g30747/_0_  ;
	output \g30748/_0_  ;
	output \g30749/_0_  ;
	output \g30750/_0_  ;
	output \g30751/_0_  ;
	output \g30752/_0_  ;
	output \g30789/_0_  ;
	output \g30790/_0_  ;
	output \g30791/_0_  ;
	output \g30792/_0_  ;
	output \g30793/_0_  ;
	output \g30794/_0_  ;
	output \g30795/_0_  ;
	output \g30796/_0_  ;
	output \g30797/_0_  ;
	output \g30798/_0_  ;
	output \g30799/_0_  ;
	output \g30800/_0_  ;
	output \g30801/_0_  ;
	output \g30802/_0_  ;
	output \g30803/_0_  ;
	output \g30804/_0_  ;
	output \g30805/_0_  ;
	output \g30806/_0_  ;
	output \g30807/_0_  ;
	output \g30808/_0_  ;
	output \g30809/_0_  ;
	output \g30810/_0_  ;
	output \g30811/_0_  ;
	output \g30812/_0_  ;
	output \g30813/_0_  ;
	output \g30814/_0_  ;
	output \g30815/_0_  ;
	output \g30816/_0_  ;
	output \g30817/_0_  ;
	output \g30818/_0_  ;
	output \g30819/_0_  ;
	output \g30820/_0_  ;
	output \g30821/_0_  ;
	output \g30822/_0_  ;
	output \g30823/_0_  ;
	output \g30824/_0_  ;
	output \g30825/_0_  ;
	output \g30826/_0_  ;
	output \g30827/_0_  ;
	output \g30828/_0_  ;
	output \g30829/_0_  ;
	output \g30830/_0_  ;
	output \g30831/_0_  ;
	output \g30832/_0_  ;
	output \g30833/_0_  ;
	output \g30834/_0_  ;
	output \g30835/_0_  ;
	output \g30836/_0_  ;
	output \g30837/_0_  ;
	output \g30838/_0_  ;
	output \g30839/_0_  ;
	output \g30840/_0_  ;
	output \g30841/_0_  ;
	output \g30842/_0_  ;
	output \g30843/_0_  ;
	output \g30844/_0_  ;
	output \g30845/_0_  ;
	output \g30846/_0_  ;
	output \g30847/_0_  ;
	output \g30848/_0_  ;
	output \g30849/_0_  ;
	output \g30850/_0_  ;
	output \g30851/_0_  ;
	output \g30852/_0_  ;
	output \g30853/_0_  ;
	output \g30854/_0_  ;
	output \g30855/_0_  ;
	output \g30856/_0_  ;
	output \g30857/_0_  ;
	output \g30858/_0_  ;
	output \g30859/_0_  ;
	output \g30860/_0_  ;
	output \g30861/_0_  ;
	output \g30862/_0_  ;
	output \g30863/_0_  ;
	output \g30864/_0_  ;
	output \g30865/_0_  ;
	output \g30866/_0_  ;
	output \g30867/_0_  ;
	output \g30868/_0_  ;
	output \g30869/_0_  ;
	output \g30870/_0_  ;
	output \g30871/_0_  ;
	output \g30872/_0_  ;
	output \g30873/_0_  ;
	output \g30874/_0_  ;
	output \g30875/_0_  ;
	output \g30876/_0_  ;
	output \g30877/_0_  ;
	output \g30878/_0_  ;
	output \g30879/_0_  ;
	output \g30880/_0_  ;
	output \g30881/_0_  ;
	output \g30882/_0_  ;
	output \g30883/_0_  ;
	output \g30884/_0_  ;
	output \g30885/_0_  ;
	output \g30886/_0_  ;
	output \g30887/_0_  ;
	output \g30888/_0_  ;
	output \g30889/_0_  ;
	output \g30890/_0_  ;
	output \g30891/_0_  ;
	output \g30892/_0_  ;
	output \g30893/_0_  ;
	output \g30894/_0_  ;
	output \g30895/_0_  ;
	output \g30896/_0_  ;
	output \g30897/_0_  ;
	output \g30898/_0_  ;
	output \g30899/_0_  ;
	output \g30900/_0_  ;
	output \g30901/_0_  ;
	output \g30902/_0_  ;
	output \g30906/_0_  ;
	output \g30907/_0_  ;
	output \g30908/_0_  ;
	output \g30909/_0_  ;
	output \g30910/_0_  ;
	output \g30911/_0_  ;
	output \g30918/_0_  ;
	output \g30919/_0_  ;
	output \g30920/_0_  ;
	output \g30921/_0_  ;
	output \g30922/_0_  ;
	output \g30923/_0_  ;
	output \g30924/_0_  ;
	output \g30925/_0_  ;
	output \g30926/_0_  ;
	output \g30946/_0_  ;
	output \g30947/_0_  ;
	output \g30948/_0_  ;
	output \g30949/_0_  ;
	output \g30950/_0_  ;
	output \g30951/_0_  ;
	output \g30952/_0_  ;
	output \g30953/_0_  ;
	output \g30954/_0_  ;
	output \g30955/_0_  ;
	output \g30956/_0_  ;
	output \g30957/_0_  ;
	output \g30958/_0_  ;
	output \g30959/_0_  ;
	output \g30960/_0_  ;
	output \g30961/_0_  ;
	output \g30962/_0_  ;
	output \g30963/_0_  ;
	output \g30964/_0_  ;
	output \g30965/_0_  ;
	output \g30966/_0_  ;
	output \g30967/_0_  ;
	output \g30968/_0_  ;
	output \g30969/_0_  ;
	output \g30970/_0_  ;
	output \g30971/_0_  ;
	output \g30972/_0_  ;
	output \g30973/_0_  ;
	output \g30974/_0_  ;
	output \g30975/_0_  ;
	output \g30976/_0_  ;
	output \g30977/_0_  ;
	output \g30978/_0_  ;
	output \g30979/_0_  ;
	output \g30980/_0_  ;
	output \g30981/_0_  ;
	output \g30982/_0_  ;
	output \g30983/_0_  ;
	output \g30984/_0_  ;
	output \g30985/_0_  ;
	output \g30986/_0_  ;
	output \g30987/_0_  ;
	output \g30988/_0_  ;
	output \g30989/_0_  ;
	output \g30990/_0_  ;
	output \g30991/_0_  ;
	output \g30992/_0_  ;
	output \g30993/_0_  ;
	output \g30994/_0_  ;
	output \g30995/_0_  ;
	output \g30996/_0_  ;
	output \g30997/_0_  ;
	output \g30998/_0_  ;
	output \g30999/_0_  ;
	output \g31000/_0_  ;
	output \g31001/_0_  ;
	output \g31002/_0_  ;
	output \g31003/_0_  ;
	output \g31004/_0_  ;
	output \g31005/_0_  ;
	output \g31006/_0_  ;
	output \g31007/_0_  ;
	output \g31008/_0_  ;
	output \g31009/_0_  ;
	output \g31010/_0_  ;
	output \g31011/_0_  ;
	output \g31012/_0_  ;
	output \g31013/_0_  ;
	output \g31014/_0_  ;
	output \g31015/_0_  ;
	output \g31016/_0_  ;
	output \g31017/_0_  ;
	output \g31018/_0_  ;
	output \g31019/_0_  ;
	output \g31020/_0_  ;
	output \g31021/_0_  ;
	output \g31022/_0_  ;
	output \g31023/_0_  ;
	output \g31024/_0_  ;
	output \g31025/_0_  ;
	output \g31026/_0_  ;
	output \g31027/_0_  ;
	output \g31028/_0_  ;
	output \g31029/_0_  ;
	output \g31030/_0_  ;
	output \g31031/_0_  ;
	output \g31032/_0_  ;
	output \g31033/_0_  ;
	output \g31034/_0_  ;
	output \g31035/_0_  ;
	output \g31036/_0_  ;
	output \g31037/_0_  ;
	output \g31038/_0_  ;
	output \g31039/_0_  ;
	output \g31040/_0_  ;
	output \g31041/_0_  ;
	output \g31042/_0_  ;
	output \g31043/_0_  ;
	output \g31044/_0_  ;
	output \g31045/_0_  ;
	output \g31046/_0_  ;
	output \g31047/_0_  ;
	output \g31048/_0_  ;
	output \g31049/_0_  ;
	output \g31050/_0_  ;
	output \g31051/_0_  ;
	output \g31052/_0_  ;
	output \g31053/_0_  ;
	output \g31054/_0_  ;
	output \g31055/_0_  ;
	output \g31056/_0_  ;
	output \g31057/_0_  ;
	output \g31058/_0_  ;
	output \g31059/_0_  ;
	output \g31060/_0_  ;
	output \g31061/_0_  ;
	output \g31062/_0_  ;
	output \g31063/_0_  ;
	output \g31064/_0_  ;
	output \g31065/_0_  ;
	output \g31066/_0_  ;
	output \g31067/_0_  ;
	output \g31068/_0_  ;
	output \g31069/_0_  ;
	output \g31070/_0_  ;
	output \g31071/_0_  ;
	output \g31072/_0_  ;
	output \g31073/_0_  ;
	output \g31074/_0_  ;
	output \g31075/_0_  ;
	output \g31076/_0_  ;
	output \g31077/_0_  ;
	output \g31084/u3_syn_4  ;
	output \g31085/u3_syn_4  ;
	output \g31096/u3_syn_4  ;
	output \g31115/u3_syn_4  ;
	output \g31136/u3_syn_4  ;
	output \g31158/u3_syn_4  ;
	output \g31176/u3_syn_4  ;
	output \g31193/u3_syn_4  ;
	output \g31195/u3_syn_4  ;
	output \g31247/u3_syn_4  ;
	output \g31280/u3_syn_4  ;
	output \g31285/u3_syn_4  ;
	output \g31568/_0_  ;
	output \g31631/_0_  ;
	output \g31672/_0_  ;
	output \g31731/_0_  ;
	output \g31732/_0_  ;
	output \g31742/_2_  ;
	output \g31744/_2_  ;
	output \g31746/_2_  ;
	output \g31748/_2_  ;
	output \g31751/_2_  ;
	output \g31754/_2_  ;
	output \g31756/_2_  ;
	output \g31758/_2_  ;
	output \g31760/_2_  ;
	output \g31761/_0_  ;
	output \g31789/_0_  ;
	output \g31807/_3_  ;
	output \g31825/_3_  ;
	output \g32607/_0_  ;
	output \g32608/_0_  ;
	output \g32609/_0_  ;
	output \g32610/_0_  ;
	output \g32611/_0_  ;
	output \g32612/_0_  ;
	output \g32613/_0_  ;
	output \g32614/_0_  ;
	output \g32615/_0_  ;
	output \g32616/_0_  ;
	output \g32617/_0_  ;
	output \g32618/_0_  ;
	output \g32645/_0__syn_2  ;
	output \g32687/_0__syn_2  ;
	output \g32749/_0__syn_2  ;
	output \g32757/_0_  ;
	output \g32758/_0_  ;
	output \g32759/_0_  ;
	output \g32760/_0_  ;
	output \g32761/_0_  ;
	output \g32762/_0_  ;
	output \g32763/_0_  ;
	output \g32764/_0_  ;
	output \g32765/_0_  ;
	output \g32769/_0_  ;
	output \g32835/_1_  ;
	output \g32839/_0_  ;
	output \g32844/_0_  ;
	output \g32901/_1_  ;
	output \g32902/_0_  ;
	output \g32963/_1_  ;
	output \g32972/_0_  ;
	output \g32977/_0_  ;
	output \g32979/_0_  ;
	output \g32980/_0_  ;
	output \g32981/_0_  ;
	output \g32982/_0_  ;
	output \g32983/_0_  ;
	output \g32987/_0_  ;
	output \g33018/_0_  ;
	output \g33019/_0_  ;
	output \g33088/_0_  ;
	output \g33261/_0_  ;
	output \g33264/_0_  ;
	output \g33275/_0_  ;
	output \g33276/_0_  ;
	output \g33277/_0_  ;
	output \g33371/_0_  ;
	output \g33382/_0_  ;
	output \g33401/_0_  ;
	output \g33402/_0_  ;
	output \g33403/_0_  ;
	output \g33404/_0_  ;
	output \g33405/_0_  ;
	output \g33406/_0_  ;
	output \g33407/_0_  ;
	output \g33408/_0_  ;
	output \g33409/_0_  ;
	output \g33410/_0_  ;
	output \g33411/_0_  ;
	output \g33412/_0_  ;
	output \g33413/_0_  ;
	output \g33414/_0_  ;
	output \g33415/_0_  ;
	output \g33416/_0_  ;
	output \g33417/_0_  ;
	output \g33418/_0_  ;
	output \g33419/_0_  ;
	output \g33420/_0_  ;
	output \g33421/_0_  ;
	output \g33422/_0_  ;
	output \g33423/_0_  ;
	output \g33424/_0_  ;
	output \g33425/_0_  ;
	output \g33426/_0_  ;
	output \g33427/_0_  ;
	output \g33428/_0_  ;
	output \g33429/_0_  ;
	output \g33430/_0_  ;
	output \g33431/_0_  ;
	output \g33432/_0_  ;
	output \g33433/_0_  ;
	output \g33434/_0_  ;
	output \g33435/_0_  ;
	output \g33436/_0_  ;
	output \g33437/_0_  ;
	output \g33438/_0_  ;
	output \g33439/_0_  ;
	output \g33440/_0_  ;
	output \g33441/_0_  ;
	output \g33442/_0_  ;
	output \g33443/_0_  ;
	output \g33444/_0_  ;
	output \g33445/_0_  ;
	output \g33446/_0_  ;
	output \g33447/_0_  ;
	output \g33448/_0_  ;
	output \g33449/_0_  ;
	output \g33450/_0_  ;
	output \g33451/_0_  ;
	output \g33452/_0_  ;
	output \g33453/_0_  ;
	output \g33454/_0_  ;
	output \g33455/_0_  ;
	output \g33456/_0_  ;
	output \g33457/_0_  ;
	output \g33458/_0_  ;
	output \g33459/_0_  ;
	output \g33460/_0_  ;
	output \g33461/_0_  ;
	output \g33462/_0_  ;
	output \g33463/_0_  ;
	output \g33464/_0_  ;
	output \g33465/_0_  ;
	output \g33466/_0_  ;
	output \g33467/_0_  ;
	output \g33468/_0_  ;
	output \g33469/_0_  ;
	output \g33470/_0_  ;
	output \g33471/_0_  ;
	output \g33472/_0_  ;
	output \g33473/_0_  ;
	output \g33474/_0_  ;
	output \g33475/_0_  ;
	output \g33476/_0_  ;
	output \g33477/_0_  ;
	output \g33478/_0_  ;
	output \g33479/_0_  ;
	output \g33480/_0_  ;
	output \g33481/_0_  ;
	output \g33482/_0_  ;
	output \g33483/_0_  ;
	output \g33484/_0_  ;
	output \g33485/_0_  ;
	output \g33486/_0_  ;
	output \g33487/_0_  ;
	output \g33488/_0_  ;
	output \g33489/_0_  ;
	output \g33490/_0_  ;
	output \g33491/_0_  ;
	output \g33492/_0_  ;
	output \g33493/_0_  ;
	output \g33494/_0_  ;
	output \g33495/_0_  ;
	output \g33496/_0_  ;
	output \g33497/_0_  ;
	output \g33498/_0_  ;
	output \g33499/_0_  ;
	output \g33500/_0_  ;
	output \g33501/_0_  ;
	output \g33502/_0_  ;
	output \g33503/_0_  ;
	output \g33504/_0_  ;
	output \g33505/_0_  ;
	output \g33506/_0_  ;
	output \g33507/_0_  ;
	output \g33508/_0_  ;
	output \g33509/_0_  ;
	output \g33510/_0_  ;
	output \g33511/_0_  ;
	output \g33512/_0_  ;
	output \g33513/_0_  ;
	output \g33514/_0_  ;
	output \g33515/_0_  ;
	output \g33516/_0_  ;
	output \g33517/_0_  ;
	output \g33518/_0_  ;
	output \g33519/_0_  ;
	output \g33520/_0_  ;
	output \g33521/_0_  ;
	output \g33522/_0_  ;
	output \g33523/_0_  ;
	output \g33524/_0_  ;
	output \g33525/_0_  ;
	output \g33526/_0_  ;
	output \g33527/_0_  ;
	output \g33528/_0_  ;
	output \g33529/_0_  ;
	output \g33530/_0_  ;
	output \g33531/_0_  ;
	output \g33532/_0_  ;
	output \g33533/_0_  ;
	output \g33534/_0_  ;
	output \g33535/_0_  ;
	output \g33536/_0_  ;
	output \g33537/_0_  ;
	output \g33538/_0_  ;
	output \g33539/_0_  ;
	output \g33540/_0_  ;
	output \g33541/_0_  ;
	output \g33542/_0_  ;
	output \g33543/_0_  ;
	output \g33544/_0_  ;
	output \g33545/_0_  ;
	output \g33546/_0_  ;
	output \g33547/_0_  ;
	output \g33548/_0_  ;
	output \g33549/_0_  ;
	output \g33550/_0_  ;
	output \g33551/_0_  ;
	output \g33552/_0_  ;
	output \g33553/_0_  ;
	output \g33554/_0_  ;
	output \g33555/_0_  ;
	output \g33556/_0_  ;
	output \g33557/_0_  ;
	output \g33558/_0_  ;
	output \g33559/_0_  ;
	output \g33560/_0_  ;
	output \g33561/_0_  ;
	output \g33562/_0_  ;
	output \g33563/_0_  ;
	output \g33564/_0_  ;
	output \g33565/_0_  ;
	output \g33566/_0_  ;
	output \g33567/_0_  ;
	output \g33568/_0_  ;
	output \g33569/_0_  ;
	output \g33570/_0_  ;
	output \g33571/_0_  ;
	output \g33572/_0_  ;
	output \g33573/_0_  ;
	output \g33574/_0_  ;
	output \g33575/_0_  ;
	output \g33576/_0_  ;
	output \g33577/_0_  ;
	output \g33578/_0_  ;
	output \g33579/_0_  ;
	output \g33580/_0_  ;
	output \g33581/_0_  ;
	output \g33582/_0_  ;
	output \g33583/_0_  ;
	output \g33584/_0_  ;
	output \g33585/_0_  ;
	output \g33586/_0_  ;
	output \g33587/_0_  ;
	output \g33588/_0_  ;
	output \g33589/_0_  ;
	output \g33590/_0_  ;
	output \g33591/_0_  ;
	output \g33592/_0_  ;
	output \g33593/_0_  ;
	output \g33594/_0_  ;
	output \g33595/_0_  ;
	output \g33596/_0_  ;
	output \g33597/_0_  ;
	output \g33598/_0_  ;
	output \g33599/_0_  ;
	output \g33600/_0_  ;
	output \g33601/_0_  ;
	output \g33602/_0_  ;
	output \g33603/_0_  ;
	output \g33604/_0_  ;
	output \g33605/_0_  ;
	output \g33606/_0_  ;
	output \g33607/_0_  ;
	output \g33608/_0_  ;
	output \g33609/_0_  ;
	output \g33610/_0_  ;
	output \g33611/_0_  ;
	output \g33612/_0_  ;
	output \g33613/_0_  ;
	output \g33614/_0_  ;
	output \g33615/_0_  ;
	output \g33616/_0_  ;
	output \g33617/_0_  ;
	output \g33618/_0_  ;
	output \g33619/_0_  ;
	output \g33620/_0_  ;
	output \g33621/_0_  ;
	output \g33622/_0_  ;
	output \g33623/_0_  ;
	output \g33624/_0_  ;
	output \g33625/_0_  ;
	output \g33626/_0_  ;
	output \g33627/_0_  ;
	output \g33628/_0_  ;
	output \g33629/_0_  ;
	output \g33630/_0_  ;
	output \g33631/_0_  ;
	output \g33632/_0_  ;
	output \g33633/_0_  ;
	output \g33634/_0_  ;
	output \g33635/_0_  ;
	output \g33636/_0_  ;
	output \g33637/_0_  ;
	output \g33638/_0_  ;
	output \g33639/_0_  ;
	output \g33640/_0_  ;
	output \g33641/_0_  ;
	output \g33642/_0_  ;
	output \g33643/_0_  ;
	output \g33644/_0_  ;
	output \g33645/_0_  ;
	output \g33646/_0_  ;
	output \g33647/_0_  ;
	output \g33648/_0_  ;
	output \g33649/_0_  ;
	output \g33650/_0_  ;
	output \g33651/_0_  ;
	output \g33652/_0_  ;
	output \g33653/_0_  ;
	output \g33654/_0_  ;
	output \g33655/_0_  ;
	output \g33656/_0_  ;
	output \g33657/_0_  ;
	output \g33658/_0_  ;
	output \g33659/_0_  ;
	output \g33660/_0_  ;
	output \g33661/_0_  ;
	output \g33662/_0_  ;
	output \g33663/_0_  ;
	output \g33664/_0_  ;
	output \g33665/_0_  ;
	output \g33666/_0_  ;
	output \g33667/_0_  ;
	output \g33668/_0_  ;
	output \g33669/_0_  ;
	output \g33670/_0_  ;
	output \g33671/_0_  ;
	output \g33672/_0_  ;
	output \g33673/_0_  ;
	output \g33674/_0_  ;
	output \g33675/_0_  ;
	output \g33676/_0_  ;
	output \g33677/_0_  ;
	output \g33678/_0_  ;
	output \g33679/_0_  ;
	output \g33680/_0_  ;
	output \g33681/_0_  ;
	output \g33682/_0_  ;
	output \g33683/_0_  ;
	output \g33684/_0_  ;
	output \g33685/_0_  ;
	output \g33686/_0_  ;
	output \g33687/_0_  ;
	output \g33688/_0_  ;
	output \g33689/_0_  ;
	output \g33690/_0_  ;
	output \g33691/_0_  ;
	output \g33692/_0_  ;
	output \g33693/_0_  ;
	output \g33694/_0_  ;
	output \g33695/_0_  ;
	output \g33696/_0_  ;
	output \g33697/_0_  ;
	output \g33698/_0_  ;
	output \g33699/_0_  ;
	output \g33700/_0_  ;
	output \g33701/_0_  ;
	output \g33702/_0_  ;
	output \g33703/_0_  ;
	output \g33704/_0_  ;
	output \g33705/_0_  ;
	output \g33706/_0_  ;
	output \g33707/_0_  ;
	output \g33708/_0_  ;
	output \g33709/_0_  ;
	output \g33710/_0_  ;
	output \g33711/_0_  ;
	output \g33712/_0_  ;
	output \g33713/_0_  ;
	output \g33714/_0_  ;
	output \g33715/_0_  ;
	output \g33716/_0_  ;
	output \g33717/_0_  ;
	output \g33718/_0_  ;
	output \g33719/_0_  ;
	output \g33720/_0_  ;
	output \g33721/_0_  ;
	output \g33722/_0_  ;
	output \g33723/_0_  ;
	output \g33724/_0_  ;
	output \g33725/_0_  ;
	output \g33726/_0_  ;
	output \g33727/_0_  ;
	output \g33728/_0_  ;
	output \g33729/_0_  ;
	output \g33730/_0_  ;
	output \g33731/_0_  ;
	output \g33732/_0_  ;
	output \g33733/_0_  ;
	output \g33734/_0_  ;
	output \g33735/_0_  ;
	output \g33736/_0_  ;
	output \g33737/_0_  ;
	output \g33738/_0_  ;
	output \g33739/_0_  ;
	output \g33740/_0_  ;
	output \g33741/_0_  ;
	output \g33742/_0_  ;
	output \g33743/_0_  ;
	output \g33744/_0_  ;
	output \g33745/_0_  ;
	output \g33746/_0_  ;
	output \g33747/_0_  ;
	output \g33748/_0_  ;
	output \g33749/_0_  ;
	output \g33750/_0_  ;
	output \g33751/_0_  ;
	output \g33752/_0_  ;
	output \g33753/_0_  ;
	output \g33754/_0_  ;
	output \g33755/_0_  ;
	output \g33756/_0_  ;
	output \g33757/_0_  ;
	output \g33758/_0_  ;
	output \g33759/_0_  ;
	output \g33760/_0_  ;
	output \g33761/_0_  ;
	output \g33762/_0_  ;
	output \g33763/_0_  ;
	output \g33764/_0_  ;
	output \g33765/_0_  ;
	output \g33766/_0_  ;
	output \g33767/_0_  ;
	output \g33768/_0_  ;
	output \g33769/_0_  ;
	output \g33770/_0_  ;
	output \g33771/_0_  ;
	output \g33772/_0_  ;
	output \g33773/_0_  ;
	output \g33774/_0_  ;
	output \g33775/_0_  ;
	output \g33776/_0_  ;
	output \g33777/_0_  ;
	output \g33778/_0_  ;
	output \g33779/_0_  ;
	output \g33780/_0_  ;
	output \g33781/_0_  ;
	output \g33782/_0_  ;
	output \g33783/_0_  ;
	output \g33784/_0_  ;
	output \g33785/_0_  ;
	output \g33786/_0_  ;
	output \g33787/_0_  ;
	output \g33788/_0_  ;
	output \g33789/_0_  ;
	output \g33790/_0_  ;
	output \g33791/_0_  ;
	output \g33792/_0_  ;
	output \g33793/_0_  ;
	output \g33794/_0_  ;
	output \g33795/_0_  ;
	output \g33796/_0_  ;
	output \g33797/_0_  ;
	output \g33798/_0_  ;
	output \g33799/_0_  ;
	output \g33800/_0_  ;
	output \g33801/_0_  ;
	output \g33802/_0_  ;
	output \g33803/_0_  ;
	output \g33804/_0_  ;
	output \g33805/_0_  ;
	output \g33806/_0_  ;
	output \g33807/_0_  ;
	output \g33808/_0_  ;
	output \g33809/_0_  ;
	output \g33810/_0_  ;
	output \g33811/_0_  ;
	output \g33812/_0_  ;
	output \g33813/_0_  ;
	output \g33814/_0_  ;
	output \g33815/_0_  ;
	output \g33816/_0_  ;
	output \g33817/_0_  ;
	output \g33818/_0_  ;
	output \g33819/_0_  ;
	output \g33820/_0_  ;
	output \g33821/_0_  ;
	output \g33822/_0_  ;
	output \g33823/_0_  ;
	output \g33824/_0_  ;
	output \g33825/_0_  ;
	output \g33826/_0_  ;
	output \g33827/_0_  ;
	output \g33828/_0_  ;
	output \g33829/_0_  ;
	output \g33830/_0_  ;
	output \g33831/_0_  ;
	output \g33832/_0_  ;
	output \g33833/_0_  ;
	output \g33834/_0_  ;
	output \g33835/_0_  ;
	output \g33836/_0_  ;
	output \g33837/_0_  ;
	output \g33838/_0_  ;
	output \g33839/_0_  ;
	output \g33840/_0_  ;
	output \g33841/_0_  ;
	output \g33842/_0_  ;
	output \g33843/_0_  ;
	output \g33844/_0_  ;
	output \g33845/_0_  ;
	output \g33846/_0_  ;
	output \g33847/_0_  ;
	output \g33848/_0_  ;
	output \g33849/_0_  ;
	output \g33850/_0_  ;
	output \g33851/_0_  ;
	output \g33852/_0_  ;
	output \g33853/_0_  ;
	output \g33854/_0_  ;
	output \g33855/_0_  ;
	output \g33856/_0_  ;
	output \g33857/_0_  ;
	output \g33858/_0_  ;
	output \g33859/_0_  ;
	output \g33860/_0_  ;
	output \g33861/_0_  ;
	output \g33862/_0_  ;
	output \g33863/_0_  ;
	output \g33864/_0_  ;
	output \g33865/_0_  ;
	output \g33866/_0_  ;
	output \g33867/_0_  ;
	output \g33868/_0_  ;
	output \g33869/_0_  ;
	output \g33870/_0_  ;
	output \g33871/_0_  ;
	output \g33872/_0_  ;
	output \g33873/_0_  ;
	output \g33874/_0_  ;
	output \g33875/_0_  ;
	output \g33876/_0_  ;
	output \g33877/_0_  ;
	output \g33878/_0_  ;
	output \g33879/_0_  ;
	output \g33880/_0_  ;
	output \g33881/_0_  ;
	output \g33882/_0_  ;
	output \g33883/_0_  ;
	output \g33884/_0_  ;
	output \g33885/_0_  ;
	output \g33886/_0_  ;
	output \g33887/_0_  ;
	output \g33888/_0_  ;
	output \g33889/_0_  ;
	output \g33890/_0_  ;
	output \g33891/_0_  ;
	output \g33892/_0_  ;
	output \g33893/_0_  ;
	output \g33894/_0_  ;
	output \g33895/_0_  ;
	output \g33896/_0_  ;
	output \g33897/_0_  ;
	output \g33898/_0_  ;
	output \g33899/_0_  ;
	output \g33900/_0_  ;
	output \g33901/_0_  ;
	output \g33902/_0_  ;
	output \g33903/_0_  ;
	output \g33904/_0_  ;
	output \g33905/_0_  ;
	output \g33906/_0_  ;
	output \g33907/_0_  ;
	output \g33908/_0_  ;
	output \g33909/_0_  ;
	output \g33910/_0_  ;
	output \g33911/_0_  ;
	output \g33912/_0_  ;
	output \g33913/_0_  ;
	output \g33914/_0_  ;
	output \g33915/_0_  ;
	output \g33916/_0_  ;
	output \g33917/_0_  ;
	output \g33918/_0_  ;
	output \g33919/_0_  ;
	output \g33920/_0_  ;
	output \g33921/_0_  ;
	output \g33922/_0_  ;
	output \g33923/_0_  ;
	output \g33924/_0_  ;
	output \g33925/_0_  ;
	output \g33926/_0_  ;
	output \g33927/_0_  ;
	output \g33928/_0_  ;
	output \g33929/_0_  ;
	output \g33930/_0_  ;
	output \g33931/_0_  ;
	output \g33932/_0_  ;
	output \g33933/_0_  ;
	output \g33934/_0_  ;
	output \g33935/_0_  ;
	output \g33936/_0_  ;
	output \g33937/_0_  ;
	output \g33938/_0_  ;
	output \g33939/_0_  ;
	output \g33940/_0_  ;
	output \g33941/_0_  ;
	output \g33942/_0_  ;
	output \g33943/_0_  ;
	output \g33944/_0_  ;
	output \g33945/_0_  ;
	output \g33946/_0_  ;
	output \g33947/_0_  ;
	output \g33948/_0_  ;
	output \g33949/_0_  ;
	output \g33950/_0_  ;
	output \g33951/_0_  ;
	output \g33952/_0_  ;
	output \g33953/_0_  ;
	output \g33954/_0_  ;
	output \g33955/_0_  ;
	output \g33956/_0_  ;
	output \g33957/_0_  ;
	output \g33958/_0_  ;
	output \g33959/_0_  ;
	output \g33960/_0_  ;
	output \g33961/_0_  ;
	output \g33962/_0_  ;
	output \g33963/_0_  ;
	output \g33964/_0_  ;
	output \g33965/_0_  ;
	output \g33966/_0_  ;
	output \g33967/_0_  ;
	output \g33968/_0_  ;
	output \g33969/_0_  ;
	output \g33970/_0_  ;
	output \g33971/_0_  ;
	output \g33972/_0_  ;
	output \g33973/_0_  ;
	output \g33974/_0_  ;
	output \g33975/_0_  ;
	output \g33976/_0_  ;
	output \g33977/u3_syn_4  ;
	output \g33981/u3_syn_4  ;
	output \g34014/u3_syn_4  ;
	output \g34047/u3_syn_4  ;
	output \g34084/u3_syn_4  ;
	output \g34123/u3_syn_4  ;
	output \g34306/_0_  ;
	output \g34316/_0_  ;
	output \g34324/_0_  ;
	output \g34326/_0_  ;
	output \g34328/_0_  ;
	output \g34331/_0_  ;
	output \g34333/_0_  ;
	output \g34344/_0_  ;
	output \g34347/_0_  ;
	output \g34351/_0_  ;
	output \g34361/_0_  ;
	output \g34368/_0_  ;
	output \g34377/_0_  ;
	output \g34385/_0_  ;
	output \g34393/_0_  ;
	output \g34414/_1_  ;
	output \g34451/_1_  ;
	output \g34476/_1_  ;
	output \g34487/_0_  ;
	output \g34490/_1_  ;
	output \g34715/_0_  ;
	output \g34878/_0_  ;
	output \g34882/_0_  ;
	output \g34883/_0_  ;
	output \g34893/_0_  ;
	output \g34896/_0_  ;
	output \g34898/_0_  ;
	output \g34899/_0_  ;
	output \g34916/_3_  ;
	output \g35264/_0_  ;
	output \g35265/_0_  ;
	output \g35266/_0_  ;
	output \g35267/_0_  ;
	output \g35268/_0_  ;
	output \g35269/_0_  ;
	output \g35270/_0_  ;
	output \g35271/_0_  ;
	output \g35272/_0_  ;
	output \g35273/_0_  ;
	output \g35274/_0_  ;
	output \g35275/_0_  ;
	output \g35276/_0_  ;
	output \g35277/_0_  ;
	output \g35278/_0_  ;
	output \g35279/_0_  ;
	output \g35283/_0_  ;
	output \g35287/_0_  ;
	output \g35294/_0_  ;
	output \g35300/_0_  ;
	output \g35304/_0_  ;
	output \g35308/_0_  ;
	output \g35312/_0_  ;
	output \g35316/_0_  ;
	output \g35318/_0_  ;
	output \g35326/_0_  ;
	output \g35334/_0_  ;
	output \g35336/_0_  ;
	output \g35337/_0_  ;
	output \g35338/_0_  ;
	output \g35357/_0_  ;
	output \g35358/_0_  ;
	output \g35359/_0_  ;
	output \g35419/_0_  ;
	output \g35438/_0_  ;
	output \g35439/_0_  ;
	output \g35440/_0_  ;
	output \g35441/_0_  ;
	output \g35442/_0_  ;
	output \g35444/_0_  ;
	output \g35445/_0_  ;
	output \g35446/_0_  ;
	output \g35447/_0_  ;
	output \g35448/_0_  ;
	output \g35449/_0_  ;
	output \g35450/_0_  ;
	output \g35451/_0_  ;
	output \g35452/_0_  ;
	output \g35463/_0_  ;
	output \g35464/_0_  ;
	output \g35466/_0_  ;
	output \g35485/_2_  ;
	output \g35495/_0_  ;
	output \g35496/_0_  ;
	output \g35499/_0_  ;
	output \g35500/_0_  ;
	output \g35501/_0_  ;
	output \g35502/_0_  ;
	output \g35563/_0_  ;
	output \g35633/_0_  ;
	output \g35717/_0_  ;
	output \g35718/_0_  ;
	output \g35719/_0_  ;
	output \g35809/_0_  ;
	output \g35810/_0_  ;
	output \g35811/_0_  ;
	output \g35812/_0_  ;
	output \g35813/_0_  ;
	output \g35814/_0_  ;
	output \g35815/_0_  ;
	output \g35816/_0_  ;
	output \g35817/_0_  ;
	output \g35818/_0_  ;
	output \g35819/_0_  ;
	output \g35820/_0_  ;
	output \g35821/_0_  ;
	output \g35822/_0_  ;
	output \g35823/_0_  ;
	output \g35824/_0_  ;
	output \g35825/_0_  ;
	output \g35826/_0_  ;
	output \g35827/_0_  ;
	output \g35830/_0_  ;
	output \g35833/_0_  ;
	output \g35835/_0_  ;
	output \g35836/_0_  ;
	output \g35837/_0_  ;
	output \g35839/_0_  ;
	output \g35840/_0_  ;
	output \g35841/_0_  ;
	output \g35843/_0_  ;
	output \g35844/_0_  ;
	output \g35845/_0_  ;
	output \g35853/_0_  ;
	output \g35854/_0_  ;
	output \g35855/_0_  ;
	output \g35856/_0_  ;
	output \g36306/_0_  ;
	output \g36414/_0_  ;
	output \g36415/_0_  ;
	output \g36449/_0_  ;
	output \g36550/_0_  ;
	output \g36551/_0_  ;
	output \g36553/_0_  ;
	output \g36560/_0_  ;
	output \g36562/_3_  ;
	output \g36563/_0_  ;
	output \g36612/_0_  ;
	output \g36614/_2_  ;
	output \g36695/_0_  ;
	output \g36784/_0_  ;
	output \g36785/_0_  ;
	output \g36786/_0_  ;
	output \g36787/_0_  ;
	output \g36788/_0_  ;
	output \g36789/_0_  ;
	output \g36790/_0_  ;
	output \g36791/_0_  ;
	output \g36792/_0_  ;
	output \g36793/_0_  ;
	output \g36794/_0_  ;
	output \g36796/_0_  ;
	output \g36797/_0_  ;
	output \g36798/_0_  ;
	output \g36799/_0_  ;
	output \g36800/_0_  ;
	output \g36801/_0_  ;
	output \g36802/_0_  ;
	output \g36803/_0_  ;
	output \g36804/_0_  ;
	output \g36805/_0_  ;
	output \g36806/_0_  ;
	output \g36807/_0_  ;
	output \g36808/_0_  ;
	output \g36809/_0_  ;
	output \g36810/_0_  ;
	output \g36811/_0_  ;
	output \g36813/_0_  ;
	output \g36814/_0_  ;
	output \g36815/_0_  ;
	output \g36820/_0_  ;
	output \g36825/_0_  ;
	output \g36832/_0_  ;
	output \g36846/_0_  ;
	output \g36855/_0_  ;
	output \g36857/_0_  ;
	output \g36859/_0_  ;
	output \g36860/_0_  ;
	output \g36861/_0_  ;
	output \g36862/_0_  ;
	output \g36863/_0_  ;
	output \g36864/_0_  ;
	output \g36867/_0_  ;
	output \g36870/_0_  ;
	output \g36871/_0_  ;
	output \g36877/_0_  ;
	output \g36879/_0_  ;
	output \g36892/_0_  ;
	output \g36893/_0_  ;
	output \g36901/_0_  ;
	output \g36909/_0_  ;
	output \g36914/_0_  ;
	output \g36919/_0_  ;
	output \g36922/_0_  ;
	output \g36923/_0_  ;
	output \g36927/_0_  ;
	output \g36930/_0_  ;
	output \g36931/_0_  ;
	output \g36933/_0_  ;
	output \g36934/_0_  ;
	output \g36935/_0_  ;
	output \g36936/_0_  ;
	output \g36937/_0_  ;
	output \g36938/_0_  ;
	output \g36939/_0_  ;
	output \g36940/_0_  ;
	output \g36941/_0_  ;
	output \g36943/_0_  ;
	output \g36944/_0_  ;
	output \g36945/_0_  ;
	output \g36946/_0_  ;
	output \g36947/_0_  ;
	output \g36948/_0_  ;
	output \g36949/_0_  ;
	output \g36950/_0_  ;
	output \g36951/_0_  ;
	output \g36952/_0_  ;
	output \g36953/_0_  ;
	output \g36954/_0_  ;
	output \g36957/_0_  ;
	output \g36958/_0_  ;
	output \g36959/_0_  ;
	output \g36960/_0_  ;
	output \g36961/_0_  ;
	output \g36962/_0_  ;
	output \g36963/_0_  ;
	output \g36970/_0_  ;
	output \g36977/_0_  ;
	output \g36986/_0_  ;
	output \g36991/_0_  ;
	output \g36994/_0_  ;
	output \g37015/_0_  ;
	output \g37057/_0_  ;
	output \g37073/_0_  ;
	output \g37128/_0_  ;
	output \g37129/_0_  ;
	output \g37138/_0_  ;
	output \g37139/_0_  ;
	output \g37140/_0_  ;
	output \g37141/_0_  ;
	output \g37142/_0_  ;
	output \g37143/_0_  ;
	output \g37144/_0_  ;
	output \g37145/_0_  ;
	output \g37146/_0_  ;
	output \g37147/_0_  ;
	output \g37148/_0_  ;
	output \g37149/_0_  ;
	output \g37150/_0_  ;
	output \g37151/_0_  ;
	output \g37152/_0_  ;
	output \g37153/_0_  ;
	output \g37154/_0_  ;
	output \g37155/_0_  ;
	output \g37156/_0_  ;
	output \g37157/_0_  ;
	output \g37158/_0_  ;
	output \g37159/_0_  ;
	output \g37160/_0_  ;
	output \g37161/_0_  ;
	output \g37162/_0_  ;
	output \g37163/_0_  ;
	output \g37164/_0_  ;
	output \g37165/_0_  ;
	output \g37166/_0_  ;
	output \g37167/_0_  ;
	output \g37168/_0_  ;
	output \g37169/_0_  ;
	output \g37170/_0_  ;
	output \g37171/_0_  ;
	output \g37172/_0_  ;
	output \g37173/_0_  ;
	output \g37174/_0_  ;
	output \g37175/_0_  ;
	output \g37176/_0_  ;
	output \g37177/_0_  ;
	output \g37178/_0_  ;
	output \g37179/_0_  ;
	output \g37180/_0_  ;
	output \g37181/_0_  ;
	output \g37182/_0_  ;
	output \g37183/_0_  ;
	output \g37184/_0_  ;
	output \g37185/_0_  ;
	output \g37187/_0_  ;
	output \g37188/_0_  ;
	output \g37190/_0_  ;
	output \g37191/_0_  ;
	output \g37192/_0_  ;
	output \g37193/_0_  ;
	output \g37194/_0_  ;
	output \g37372/_3_  ;
	output \g37377/_0_  ;
	output \g37378/_0_  ;
	output \g37379/_0_  ;
	output \g37380/_0_  ;
	output \g37381/_0_  ;
	output \g37382/_0_  ;
	output \g37383/_0_  ;
	output \g37384/_0_  ;
	output \g37385/_0_  ;
	output \g37386/_0_  ;
	output \g37387/_0_  ;
	output \g37388/_0_  ;
	output \g37389/_0_  ;
	output \g37390/_0_  ;
	output \g37391/_0_  ;
	output \g37392/_0_  ;
	output \g37393/_0_  ;
	output \g37394/_0_  ;
	output \g37395/_0_  ;
	output \g37396/_0_  ;
	output \g37397/_0_  ;
	output \g37398/_0_  ;
	output \g37399/_0_  ;
	output \g37400/_0_  ;
	output \g37401/_0_  ;
	output \g37402/_0_  ;
	output \g37403/_0_  ;
	output \g37404/_0_  ;
	output \g37405/_0_  ;
	output \g37406/_0_  ;
	output \g37407/_0_  ;
	output \g37408/_0_  ;
	output \g37409/_0_  ;
	output \g37410/_0_  ;
	output \g37411/_0_  ;
	output \g37412/_0_  ;
	output \g37413/_0_  ;
	output \g37576/_3_  ;
	output \g37590/_2_  ;
	output \g40278/_0_  ;
	output \g40379/_0_  ;
	output \g40389/_2_  ;
	output \g40390/_2_  ;
	output \g40391/_0_  ;
	output \g40393/_2_  ;
	output \g40395/_0_  ;
	output \g40397/_0_  ;
	output \g40400/_0_  ;
	output \g40402/_0_  ;
	output \g45458/_0_  ;
	output \g45675/_0_  ;
	output \g45677/_0_  ;
	output \g45678/_0_  ;
	output \g45682/_0_  ;
	output sync_pad_o_pad ;
	output \u14_u0_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u1_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u2_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u3_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u4_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u5_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u6_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u7_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u14_u8_full_empty_r_reg/P0001_reg_syn_3  ;
	output \u1_slt0_reg[11]/P0001_reg_syn_3  ;
	output \u1_slt0_reg[12]/P0001_reg_syn_3  ;
	output \u1_slt0_reg[15]/P0001_reg_syn_3  ;
	output \u1_slt0_reg[9]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[10]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[11]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[5]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[6]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[7]/P0001_reg_syn_3  ;
	output \u1_slt1_reg[8]/P0001_reg_syn_3  ;
	output wb_err_o_pad ;
	wire _w10251_ ;
	wire _w10250_ ;
	wire _w10249_ ;
	wire _w10248_ ;
	wire _w10247_ ;
	wire _w10246_ ;
	wire _w10245_ ;
	wire _w10244_ ;
	wire _w10243_ ;
	wire _w10242_ ;
	wire _w10241_ ;
	wire _w10240_ ;
	wire _w10239_ ;
	wire _w10238_ ;
	wire _w10237_ ;
	wire _w10236_ ;
	wire _w10235_ ;
	wire _w10234_ ;
	wire _w10233_ ;
	wire _w10232_ ;
	wire _w10231_ ;
	wire _w10230_ ;
	wire _w10229_ ;
	wire _w10228_ ;
	wire _w10227_ ;
	wire _w10226_ ;
	wire _w10225_ ;
	wire _w10224_ ;
	wire _w10223_ ;
	wire _w10222_ ;
	wire _w10221_ ;
	wire _w10220_ ;
	wire _w10219_ ;
	wire _w10218_ ;
	wire _w10217_ ;
	wire _w10216_ ;
	wire _w10215_ ;
	wire _w10214_ ;
	wire _w10213_ ;
	wire _w10212_ ;
	wire _w10211_ ;
	wire _w10210_ ;
	wire _w10209_ ;
	wire _w10208_ ;
	wire _w10207_ ;
	wire _w10206_ ;
	wire _w10205_ ;
	wire _w10204_ ;
	wire _w10203_ ;
	wire _w10202_ ;
	wire _w10201_ ;
	wire _w10200_ ;
	wire _w10199_ ;
	wire _w10198_ ;
	wire _w10197_ ;
	wire _w10196_ ;
	wire _w10195_ ;
	wire _w10194_ ;
	wire _w10193_ ;
	wire _w10192_ ;
	wire _w10191_ ;
	wire _w10190_ ;
	wire _w10189_ ;
	wire _w10188_ ;
	wire _w10187_ ;
	wire _w10186_ ;
	wire _w10185_ ;
	wire _w10184_ ;
	wire _w10183_ ;
	wire _w10182_ ;
	wire _w10181_ ;
	wire _w10180_ ;
	wire _w10179_ ;
	wire _w10178_ ;
	wire _w10177_ ;
	wire _w10176_ ;
	wire _w10175_ ;
	wire _w10174_ ;
	wire _w10173_ ;
	wire _w10172_ ;
	wire _w10171_ ;
	wire _w10170_ ;
	wire _w10169_ ;
	wire _w10168_ ;
	wire _w10167_ ;
	wire _w10166_ ;
	wire _w10165_ ;
	wire _w10164_ ;
	wire _w10163_ ;
	wire _w10162_ ;
	wire _w10161_ ;
	wire _w10160_ ;
	wire _w10159_ ;
	wire _w10158_ ;
	wire _w10157_ ;
	wire _w10156_ ;
	wire _w10155_ ;
	wire _w10154_ ;
	wire _w10153_ ;
	wire _w10152_ ;
	wire _w10151_ ;
	wire _w10150_ ;
	wire _w10149_ ;
	wire _w10148_ ;
	wire _w10147_ ;
	wire _w10146_ ;
	wire _w10145_ ;
	wire _w10144_ ;
	wire _w10143_ ;
	wire _w10142_ ;
	wire _w10141_ ;
	wire _w10140_ ;
	wire _w10139_ ;
	wire _w10138_ ;
	wire _w10137_ ;
	wire _w10136_ ;
	wire _w10135_ ;
	wire _w10134_ ;
	wire _w10133_ ;
	wire _w10132_ ;
	wire _w10131_ ;
	wire _w10130_ ;
	wire _w10129_ ;
	wire _w10128_ ;
	wire _w10127_ ;
	wire _w10126_ ;
	wire _w10125_ ;
	wire _w10124_ ;
	wire _w10123_ ;
	wire _w10122_ ;
	wire _w10121_ ;
	wire _w10120_ ;
	wire _w10119_ ;
	wire _w10118_ ;
	wire _w10117_ ;
	wire _w10116_ ;
	wire _w10115_ ;
	wire _w10114_ ;
	wire _w10113_ ;
	wire _w10112_ ;
	wire _w10111_ ;
	wire _w10110_ ;
	wire _w10109_ ;
	wire _w10108_ ;
	wire _w10107_ ;
	wire _w10106_ ;
	wire _w10105_ ;
	wire _w10104_ ;
	wire _w10103_ ;
	wire _w10102_ ;
	wire _w10101_ ;
	wire _w10100_ ;
	wire _w10099_ ;
	wire _w10098_ ;
	wire _w10097_ ;
	wire _w10096_ ;
	wire _w10095_ ;
	wire _w10094_ ;
	wire _w10093_ ;
	wire _w10092_ ;
	wire _w10091_ ;
	wire _w10090_ ;
	wire _w10089_ ;
	wire _w10088_ ;
	wire _w10087_ ;
	wire _w10086_ ;
	wire _w10085_ ;
	wire _w10084_ ;
	wire _w10083_ ;
	wire _w10082_ ;
	wire _w10081_ ;
	wire _w10080_ ;
	wire _w10079_ ;
	wire _w10078_ ;
	wire _w10077_ ;
	wire _w10076_ ;
	wire _w10075_ ;
	wire _w10074_ ;
	wire _w10073_ ;
	wire _w10072_ ;
	wire _w10071_ ;
	wire _w10070_ ;
	wire _w10069_ ;
	wire _w10068_ ;
	wire _w10067_ ;
	wire _w10066_ ;
	wire _w10065_ ;
	wire _w10064_ ;
	wire _w10063_ ;
	wire _w10062_ ;
	wire _w10061_ ;
	wire _w10060_ ;
	wire _w10059_ ;
	wire _w10058_ ;
	wire _w10057_ ;
	wire _w10056_ ;
	wire _w10055_ ;
	wire _w10054_ ;
	wire _w10053_ ;
	wire _w10052_ ;
	wire _w10051_ ;
	wire _w10050_ ;
	wire _w10049_ ;
	wire _w10048_ ;
	wire _w10047_ ;
	wire _w10046_ ;
	wire _w10045_ ;
	wire _w10044_ ;
	wire _w10043_ ;
	wire _w10042_ ;
	wire _w10041_ ;
	wire _w10040_ ;
	wire _w10039_ ;
	wire _w10038_ ;
	wire _w10037_ ;
	wire _w10036_ ;
	wire _w10035_ ;
	wire _w10034_ ;
	wire _w10033_ ;
	wire _w10032_ ;
	wire _w10031_ ;
	wire _w10030_ ;
	wire _w10029_ ;
	wire _w10028_ ;
	wire _w10027_ ;
	wire _w10026_ ;
	wire _w10025_ ;
	wire _w10024_ ;
	wire _w10023_ ;
	wire _w10022_ ;
	wire _w10021_ ;
	wire _w10020_ ;
	wire _w10019_ ;
	wire _w10018_ ;
	wire _w10017_ ;
	wire _w10016_ ;
	wire _w10015_ ;
	wire _w10014_ ;
	wire _w10013_ ;
	wire _w10012_ ;
	wire _w10011_ ;
	wire _w10010_ ;
	wire _w10009_ ;
	wire _w10008_ ;
	wire _w10007_ ;
	wire _w10006_ ;
	wire _w10005_ ;
	wire _w10004_ ;
	wire _w10003_ ;
	wire _w10002_ ;
	wire _w10001_ ;
	wire _w10000_ ;
	wire _w9999_ ;
	wire _w9998_ ;
	wire _w9997_ ;
	wire _w9996_ ;
	wire _w9995_ ;
	wire _w9994_ ;
	wire _w9993_ ;
	wire _w9992_ ;
	wire _w9991_ ;
	wire _w9990_ ;
	wire _w9989_ ;
	wire _w9988_ ;
	wire _w9987_ ;
	wire _w9986_ ;
	wire _w9985_ ;
	wire _w9984_ ;
	wire _w9983_ ;
	wire _w9982_ ;
	wire _w9981_ ;
	wire _w9980_ ;
	wire _w9979_ ;
	wire _w9978_ ;
	wire _w9977_ ;
	wire _w9976_ ;
	wire _w9975_ ;
	wire _w9974_ ;
	wire _w9973_ ;
	wire _w9972_ ;
	wire _w9971_ ;
	wire _w9970_ ;
	wire _w9969_ ;
	wire _w9968_ ;
	wire _w9967_ ;
	wire _w9966_ ;
	wire _w9965_ ;
	wire _w9964_ ;
	wire _w9963_ ;
	wire _w9962_ ;
	wire _w9961_ ;
	wire _w9960_ ;
	wire _w9959_ ;
	wire _w9958_ ;
	wire _w9957_ ;
	wire _w9956_ ;
	wire _w9955_ ;
	wire _w9954_ ;
	wire _w9953_ ;
	wire _w9952_ ;
	wire _w9951_ ;
	wire _w9950_ ;
	wire _w9949_ ;
	wire _w9948_ ;
	wire _w9947_ ;
	wire _w9946_ ;
	wire _w9945_ ;
	wire _w9944_ ;
	wire _w9943_ ;
	wire _w9942_ ;
	wire _w9941_ ;
	wire _w9940_ ;
	wire _w9939_ ;
	wire _w9938_ ;
	wire _w9937_ ;
	wire _w9936_ ;
	wire _w9935_ ;
	wire _w9934_ ;
	wire _w9933_ ;
	wire _w9932_ ;
	wire _w9931_ ;
	wire _w9930_ ;
	wire _w9929_ ;
	wire _w9928_ ;
	wire _w9927_ ;
	wire _w9926_ ;
	wire _w9925_ ;
	wire _w9924_ ;
	wire _w9923_ ;
	wire _w9922_ ;
	wire _w9921_ ;
	wire _w9920_ ;
	wire _w9919_ ;
	wire _w9918_ ;
	wire _w9917_ ;
	wire _w9916_ ;
	wire _w9915_ ;
	wire _w9914_ ;
	wire _w9913_ ;
	wire _w9912_ ;
	wire _w9911_ ;
	wire _w9910_ ;
	wire _w9909_ ;
	wire _w9908_ ;
	wire _w9907_ ;
	wire _w9906_ ;
	wire _w9905_ ;
	wire _w9904_ ;
	wire _w9903_ ;
	wire _w9902_ ;
	wire _w9901_ ;
	wire _w9900_ ;
	wire _w9899_ ;
	wire _w9898_ ;
	wire _w9897_ ;
	wire _w9896_ ;
	wire _w9895_ ;
	wire _w9894_ ;
	wire _w9893_ ;
	wire _w9892_ ;
	wire _w9891_ ;
	wire _w9890_ ;
	wire _w9889_ ;
	wire _w9888_ ;
	wire _w9887_ ;
	wire _w9886_ ;
	wire _w9885_ ;
	wire _w9884_ ;
	wire _w9883_ ;
	wire _w9882_ ;
	wire _w9881_ ;
	wire _w9880_ ;
	wire _w9879_ ;
	wire _w9878_ ;
	wire _w9877_ ;
	wire _w9876_ ;
	wire _w9875_ ;
	wire _w9874_ ;
	wire _w9873_ ;
	wire _w9872_ ;
	wire _w9871_ ;
	wire _w9870_ ;
	wire _w9869_ ;
	wire _w9868_ ;
	wire _w9867_ ;
	wire _w9866_ ;
	wire _w9865_ ;
	wire _w9864_ ;
	wire _w9863_ ;
	wire _w9862_ ;
	wire _w9861_ ;
	wire _w9860_ ;
	wire _w9859_ ;
	wire _w9858_ ;
	wire _w9857_ ;
	wire _w9856_ ;
	wire _w9855_ ;
	wire _w9854_ ;
	wire _w9853_ ;
	wire _w9852_ ;
	wire _w9851_ ;
	wire _w9850_ ;
	wire _w9849_ ;
	wire _w9848_ ;
	wire _w9847_ ;
	wire _w9846_ ;
	wire _w9845_ ;
	wire _w9844_ ;
	wire _w9843_ ;
	wire _w9842_ ;
	wire _w9841_ ;
	wire _w9840_ ;
	wire _w9839_ ;
	wire _w9838_ ;
	wire _w9837_ ;
	wire _w9836_ ;
	wire _w9835_ ;
	wire _w9834_ ;
	wire _w9833_ ;
	wire _w9832_ ;
	wire _w9831_ ;
	wire _w9830_ ;
	wire _w9829_ ;
	wire _w9828_ ;
	wire _w9827_ ;
	wire _w9826_ ;
	wire _w9825_ ;
	wire _w9824_ ;
	wire _w9823_ ;
	wire _w9822_ ;
	wire _w9821_ ;
	wire _w9820_ ;
	wire _w9819_ ;
	wire _w9818_ ;
	wire _w9817_ ;
	wire _w9816_ ;
	wire _w9815_ ;
	wire _w9814_ ;
	wire _w9813_ ;
	wire _w9812_ ;
	wire _w9811_ ;
	wire _w9810_ ;
	wire _w9809_ ;
	wire _w9808_ ;
	wire _w9807_ ;
	wire _w9806_ ;
	wire _w9805_ ;
	wire _w9804_ ;
	wire _w9803_ ;
	wire _w9802_ ;
	wire _w9801_ ;
	wire _w9800_ ;
	wire _w9799_ ;
	wire _w9798_ ;
	wire _w9797_ ;
	wire _w9796_ ;
	wire _w9795_ ;
	wire _w9794_ ;
	wire _w9793_ ;
	wire _w9792_ ;
	wire _w9791_ ;
	wire _w9790_ ;
	wire _w9789_ ;
	wire _w9788_ ;
	wire _w9787_ ;
	wire _w9786_ ;
	wire _w9785_ ;
	wire _w9784_ ;
	wire _w9783_ ;
	wire _w9782_ ;
	wire _w9781_ ;
	wire _w9780_ ;
	wire _w9779_ ;
	wire _w9778_ ;
	wire _w9777_ ;
	wire _w9776_ ;
	wire _w9775_ ;
	wire _w9774_ ;
	wire _w9773_ ;
	wire _w9772_ ;
	wire _w9771_ ;
	wire _w9770_ ;
	wire _w9769_ ;
	wire _w9768_ ;
	wire _w9767_ ;
	wire _w9766_ ;
	wire _w9765_ ;
	wire _w9764_ ;
	wire _w9763_ ;
	wire _w9762_ ;
	wire _w9761_ ;
	wire _w9760_ ;
	wire _w9759_ ;
	wire _w9758_ ;
	wire _w9757_ ;
	wire _w9756_ ;
	wire _w9755_ ;
	wire _w9754_ ;
	wire _w9753_ ;
	wire _w9752_ ;
	wire _w9751_ ;
	wire _w9750_ ;
	wire _w9749_ ;
	wire _w9748_ ;
	wire _w9747_ ;
	wire _w9746_ ;
	wire _w9745_ ;
	wire _w9744_ ;
	wire _w9743_ ;
	wire _w9742_ ;
	wire _w9741_ ;
	wire _w9740_ ;
	wire _w9739_ ;
	wire _w9738_ ;
	wire _w9737_ ;
	wire _w9736_ ;
	wire _w9735_ ;
	wire _w9734_ ;
	wire _w9733_ ;
	wire _w9732_ ;
	wire _w9731_ ;
	wire _w9730_ ;
	wire _w9729_ ;
	wire _w9728_ ;
	wire _w9727_ ;
	wire _w9726_ ;
	wire _w9725_ ;
	wire _w9724_ ;
	wire _w9723_ ;
	wire _w9722_ ;
	wire _w9721_ ;
	wire _w9720_ ;
	wire _w9719_ ;
	wire _w9718_ ;
	wire _w9717_ ;
	wire _w9716_ ;
	wire _w9715_ ;
	wire _w9714_ ;
	wire _w9713_ ;
	wire _w9712_ ;
	wire _w9711_ ;
	wire _w9710_ ;
	wire _w9709_ ;
	wire _w9708_ ;
	wire _w9707_ ;
	wire _w9706_ ;
	wire _w9705_ ;
	wire _w9704_ ;
	wire _w9703_ ;
	wire _w9702_ ;
	wire _w9701_ ;
	wire _w9700_ ;
	wire _w9699_ ;
	wire _w9698_ ;
	wire _w9697_ ;
	wire _w9696_ ;
	wire _w9695_ ;
	wire _w9694_ ;
	wire _w9693_ ;
	wire _w9692_ ;
	wire _w9691_ ;
	wire _w9690_ ;
	wire _w9689_ ;
	wire _w9688_ ;
	wire _w9687_ ;
	wire _w9686_ ;
	wire _w9685_ ;
	wire _w9684_ ;
	wire _w9683_ ;
	wire _w9682_ ;
	wire _w9681_ ;
	wire _w9680_ ;
	wire _w9679_ ;
	wire _w9678_ ;
	wire _w9677_ ;
	wire _w9676_ ;
	wire _w9675_ ;
	wire _w9674_ ;
	wire _w9673_ ;
	wire _w9672_ ;
	wire _w9671_ ;
	wire _w9670_ ;
	wire _w9669_ ;
	wire _w9668_ ;
	wire _w9667_ ;
	wire _w9666_ ;
	wire _w9665_ ;
	wire _w9664_ ;
	wire _w9663_ ;
	wire _w9662_ ;
	wire _w9661_ ;
	wire _w9660_ ;
	wire _w9659_ ;
	wire _w9658_ ;
	wire _w9657_ ;
	wire _w9656_ ;
	wire _w9655_ ;
	wire _w9654_ ;
	wire _w9653_ ;
	wire _w9652_ ;
	wire _w9651_ ;
	wire _w9650_ ;
	wire _w9649_ ;
	wire _w9648_ ;
	wire _w9647_ ;
	wire _w9646_ ;
	wire _w9645_ ;
	wire _w9644_ ;
	wire _w9643_ ;
	wire _w9642_ ;
	wire _w9641_ ;
	wire _w9640_ ;
	wire _w9639_ ;
	wire _w9638_ ;
	wire _w9637_ ;
	wire _w9636_ ;
	wire _w9635_ ;
	wire _w9634_ ;
	wire _w9633_ ;
	wire _w9632_ ;
	wire _w9631_ ;
	wire _w9630_ ;
	wire _w9629_ ;
	wire _w9628_ ;
	wire _w9627_ ;
	wire _w9626_ ;
	wire _w9625_ ;
	wire _w9624_ ;
	wire _w9623_ ;
	wire _w9622_ ;
	wire _w9621_ ;
	wire _w9620_ ;
	wire _w9619_ ;
	wire _w9618_ ;
	wire _w9617_ ;
	wire _w9616_ ;
	wire _w9615_ ;
	wire _w9614_ ;
	wire _w9613_ ;
	wire _w9612_ ;
	wire _w9611_ ;
	wire _w9610_ ;
	wire _w9609_ ;
	wire _w9608_ ;
	wire _w9607_ ;
	wire _w9606_ ;
	wire _w9605_ ;
	wire _w9604_ ;
	wire _w9603_ ;
	wire _w9602_ ;
	wire _w9601_ ;
	wire _w9600_ ;
	wire _w9599_ ;
	wire _w9598_ ;
	wire _w9597_ ;
	wire _w9596_ ;
	wire _w9595_ ;
	wire _w9594_ ;
	wire _w9593_ ;
	wire _w9592_ ;
	wire _w9591_ ;
	wire _w9590_ ;
	wire _w9589_ ;
	wire _w9588_ ;
	wire _w9587_ ;
	wire _w9586_ ;
	wire _w9585_ ;
	wire _w9584_ ;
	wire _w9583_ ;
	wire _w9582_ ;
	wire _w9581_ ;
	wire _w9580_ ;
	wire _w9579_ ;
	wire _w9578_ ;
	wire _w9577_ ;
	wire _w9576_ ;
	wire _w9575_ ;
	wire _w9574_ ;
	wire _w9573_ ;
	wire _w9572_ ;
	wire _w9571_ ;
	wire _w9570_ ;
	wire _w9569_ ;
	wire _w9568_ ;
	wire _w9567_ ;
	wire _w9566_ ;
	wire _w9565_ ;
	wire _w9564_ ;
	wire _w9563_ ;
	wire _w9562_ ;
	wire _w9561_ ;
	wire _w9560_ ;
	wire _w9559_ ;
	wire _w9558_ ;
	wire _w9557_ ;
	wire _w9556_ ;
	wire _w9555_ ;
	wire _w9554_ ;
	wire _w9553_ ;
	wire _w9552_ ;
	wire _w9551_ ;
	wire _w9550_ ;
	wire _w9549_ ;
	wire _w9548_ ;
	wire _w9547_ ;
	wire _w9546_ ;
	wire _w9545_ ;
	wire _w9544_ ;
	wire _w9543_ ;
	wire _w9542_ ;
	wire _w9541_ ;
	wire _w9540_ ;
	wire _w9539_ ;
	wire _w9538_ ;
	wire _w9537_ ;
	wire _w9536_ ;
	wire _w9535_ ;
	wire _w9534_ ;
	wire _w9533_ ;
	wire _w9532_ ;
	wire _w9531_ ;
	wire _w9530_ ;
	wire _w9529_ ;
	wire _w9528_ ;
	wire _w9527_ ;
	wire _w9526_ ;
	wire _w9525_ ;
	wire _w9524_ ;
	wire _w9523_ ;
	wire _w9522_ ;
	wire _w9521_ ;
	wire _w9520_ ;
	wire _w9519_ ;
	wire _w9518_ ;
	wire _w9517_ ;
	wire _w9516_ ;
	wire _w9515_ ;
	wire _w9514_ ;
	wire _w9513_ ;
	wire _w9512_ ;
	wire _w9511_ ;
	wire _w9510_ ;
	wire _w9509_ ;
	wire _w9508_ ;
	wire _w9507_ ;
	wire _w9506_ ;
	wire _w9505_ ;
	wire _w9504_ ;
	wire _w9503_ ;
	wire _w9502_ ;
	wire _w9501_ ;
	wire _w9500_ ;
	wire _w9499_ ;
	wire _w9498_ ;
	wire _w9497_ ;
	wire _w9496_ ;
	wire _w9495_ ;
	wire _w9494_ ;
	wire _w9493_ ;
	wire _w9492_ ;
	wire _w9491_ ;
	wire _w9490_ ;
	wire _w9489_ ;
	wire _w9488_ ;
	wire _w9487_ ;
	wire _w9486_ ;
	wire _w9485_ ;
	wire _w9484_ ;
	wire _w9483_ ;
	wire _w9482_ ;
	wire _w9481_ ;
	wire _w9480_ ;
	wire _w9479_ ;
	wire _w9478_ ;
	wire _w9477_ ;
	wire _w9476_ ;
	wire _w9475_ ;
	wire _w9474_ ;
	wire _w9473_ ;
	wire _w9472_ ;
	wire _w9471_ ;
	wire _w9470_ ;
	wire _w9469_ ;
	wire _w9468_ ;
	wire _w9467_ ;
	wire _w9466_ ;
	wire _w9465_ ;
	wire _w9464_ ;
	wire _w9463_ ;
	wire _w9462_ ;
	wire _w9461_ ;
	wire _w9460_ ;
	wire _w9459_ ;
	wire _w9458_ ;
	wire _w9457_ ;
	wire _w9456_ ;
	wire _w9455_ ;
	wire _w9454_ ;
	wire _w9453_ ;
	wire _w9452_ ;
	wire _w9451_ ;
	wire _w9450_ ;
	wire _w9449_ ;
	wire _w9448_ ;
	wire _w9447_ ;
	wire _w9446_ ;
	wire _w9445_ ;
	wire _w9444_ ;
	wire _w9443_ ;
	wire _w9442_ ;
	wire _w9441_ ;
	wire _w9440_ ;
	wire _w9439_ ;
	wire _w9438_ ;
	wire _w9437_ ;
	wire _w9436_ ;
	wire _w9435_ ;
	wire _w9434_ ;
	wire _w9433_ ;
	wire _w9432_ ;
	wire _w9431_ ;
	wire _w9430_ ;
	wire _w9429_ ;
	wire _w9428_ ;
	wire _w9427_ ;
	wire _w9426_ ;
	wire _w9425_ ;
	wire _w9424_ ;
	wire _w9423_ ;
	wire _w9422_ ;
	wire _w9421_ ;
	wire _w9420_ ;
	wire _w9419_ ;
	wire _w9418_ ;
	wire _w9417_ ;
	wire _w9416_ ;
	wire _w9415_ ;
	wire _w9414_ ;
	wire _w9413_ ;
	wire _w9412_ ;
	wire _w9411_ ;
	wire _w9410_ ;
	wire _w9409_ ;
	wire _w9408_ ;
	wire _w9407_ ;
	wire _w9406_ ;
	wire _w9405_ ;
	wire _w9404_ ;
	wire _w9403_ ;
	wire _w9402_ ;
	wire _w9401_ ;
	wire _w9400_ ;
	wire _w9399_ ;
	wire _w9398_ ;
	wire _w9397_ ;
	wire _w9396_ ;
	wire _w9395_ ;
	wire _w9394_ ;
	wire _w9393_ ;
	wire _w9392_ ;
	wire _w9391_ ;
	wire _w9390_ ;
	wire _w9389_ ;
	wire _w9388_ ;
	wire _w9387_ ;
	wire _w9386_ ;
	wire _w9385_ ;
	wire _w9384_ ;
	wire _w9383_ ;
	wire _w9382_ ;
	wire _w9381_ ;
	wire _w9380_ ;
	wire _w9379_ ;
	wire _w9378_ ;
	wire _w9377_ ;
	wire _w9376_ ;
	wire _w9375_ ;
	wire _w9374_ ;
	wire _w9373_ ;
	wire _w9372_ ;
	wire _w9371_ ;
	wire _w9370_ ;
	wire _w9369_ ;
	wire _w9368_ ;
	wire _w9367_ ;
	wire _w9366_ ;
	wire _w9365_ ;
	wire _w9364_ ;
	wire _w9363_ ;
	wire _w9362_ ;
	wire _w9361_ ;
	wire _w9360_ ;
	wire _w9359_ ;
	wire _w9358_ ;
	wire _w9357_ ;
	wire _w9356_ ;
	wire _w9355_ ;
	wire _w9354_ ;
	wire _w9353_ ;
	wire _w9352_ ;
	wire _w9351_ ;
	wire _w9350_ ;
	wire _w9349_ ;
	wire _w9348_ ;
	wire _w9347_ ;
	wire _w9346_ ;
	wire _w9345_ ;
	wire _w9344_ ;
	wire _w9343_ ;
	wire _w9342_ ;
	wire _w9341_ ;
	wire _w9340_ ;
	wire _w9339_ ;
	wire _w9338_ ;
	wire _w9337_ ;
	wire _w9336_ ;
	wire _w9335_ ;
	wire _w9334_ ;
	wire _w9333_ ;
	wire _w9332_ ;
	wire _w9331_ ;
	wire _w9330_ ;
	wire _w9329_ ;
	wire _w9328_ ;
	wire _w9327_ ;
	wire _w9326_ ;
	wire _w9325_ ;
	wire _w9324_ ;
	wire _w9323_ ;
	wire _w9322_ ;
	wire _w9321_ ;
	wire _w9320_ ;
	wire _w9319_ ;
	wire _w9318_ ;
	wire _w9317_ ;
	wire _w9316_ ;
	wire _w9315_ ;
	wire _w9314_ ;
	wire _w9313_ ;
	wire _w9312_ ;
	wire _w9311_ ;
	wire _w9310_ ;
	wire _w9309_ ;
	wire _w9308_ ;
	wire _w9307_ ;
	wire _w9306_ ;
	wire _w9305_ ;
	wire _w9304_ ;
	wire _w9303_ ;
	wire _w9302_ ;
	wire _w9301_ ;
	wire _w9300_ ;
	wire _w9299_ ;
	wire _w9298_ ;
	wire _w9297_ ;
	wire _w9296_ ;
	wire _w9295_ ;
	wire _w9294_ ;
	wire _w9293_ ;
	wire _w9292_ ;
	wire _w9291_ ;
	wire _w9290_ ;
	wire _w9289_ ;
	wire _w9288_ ;
	wire _w9287_ ;
	wire _w9286_ ;
	wire _w9285_ ;
	wire _w9284_ ;
	wire _w9283_ ;
	wire _w9282_ ;
	wire _w9281_ ;
	wire _w9280_ ;
	wire _w9279_ ;
	wire _w9278_ ;
	wire _w9277_ ;
	wire _w9276_ ;
	wire _w9275_ ;
	wire _w9274_ ;
	wire _w9273_ ;
	wire _w9272_ ;
	wire _w9271_ ;
	wire _w9270_ ;
	wire _w9269_ ;
	wire _w9268_ ;
	wire _w9267_ ;
	wire _w9266_ ;
	wire _w9265_ ;
	wire _w9264_ ;
	wire _w9263_ ;
	wire _w9262_ ;
	wire _w9261_ ;
	wire _w9260_ ;
	wire _w9259_ ;
	wire _w9258_ ;
	wire _w9257_ ;
	wire _w9256_ ;
	wire _w9255_ ;
	wire _w9254_ ;
	wire _w9253_ ;
	wire _w9252_ ;
	wire _w9251_ ;
	wire _w9250_ ;
	wire _w9249_ ;
	wire _w9248_ ;
	wire _w9247_ ;
	wire _w9246_ ;
	wire _w9245_ ;
	wire _w9244_ ;
	wire _w9243_ ;
	wire _w9242_ ;
	wire _w9241_ ;
	wire _w9240_ ;
	wire _w9239_ ;
	wire _w9238_ ;
	wire _w9237_ ;
	wire _w9236_ ;
	wire _w9235_ ;
	wire _w9234_ ;
	wire _w9233_ ;
	wire _w9232_ ;
	wire _w9231_ ;
	wire _w9230_ ;
	wire _w9229_ ;
	wire _w9228_ ;
	wire _w9227_ ;
	wire _w9226_ ;
	wire _w9225_ ;
	wire _w9224_ ;
	wire _w9223_ ;
	wire _w9222_ ;
	wire _w9221_ ;
	wire _w9220_ ;
	wire _w9219_ ;
	wire _w9218_ ;
	wire _w9217_ ;
	wire _w9216_ ;
	wire _w9215_ ;
	wire _w9214_ ;
	wire _w9213_ ;
	wire _w9212_ ;
	wire _w9211_ ;
	wire _w9210_ ;
	wire _w9209_ ;
	wire _w9208_ ;
	wire _w9207_ ;
	wire _w9206_ ;
	wire _w9205_ ;
	wire _w9204_ ;
	wire _w9203_ ;
	wire _w9202_ ;
	wire _w9201_ ;
	wire _w9200_ ;
	wire _w9199_ ;
	wire _w9198_ ;
	wire _w9197_ ;
	wire _w9196_ ;
	wire _w9195_ ;
	wire _w9194_ ;
	wire _w9193_ ;
	wire _w9192_ ;
	wire _w9191_ ;
	wire _w9190_ ;
	wire _w9189_ ;
	wire _w9188_ ;
	wire _w9187_ ;
	wire _w9186_ ;
	wire _w9185_ ;
	wire _w9184_ ;
	wire _w9183_ ;
	wire _w9182_ ;
	wire _w9181_ ;
	wire _w9180_ ;
	wire _w9179_ ;
	wire _w9178_ ;
	wire _w9177_ ;
	wire _w9176_ ;
	wire _w9175_ ;
	wire _w9174_ ;
	wire _w9173_ ;
	wire _w9172_ ;
	wire _w9171_ ;
	wire _w9170_ ;
	wire _w9169_ ;
	wire _w9168_ ;
	wire _w9167_ ;
	wire _w9166_ ;
	wire _w9165_ ;
	wire _w9164_ ;
	wire _w9163_ ;
	wire _w9162_ ;
	wire _w9161_ ;
	wire _w9160_ ;
	wire _w9159_ ;
	wire _w9158_ ;
	wire _w9157_ ;
	wire _w9156_ ;
	wire _w9155_ ;
	wire _w9154_ ;
	wire _w9153_ ;
	wire _w9152_ ;
	wire _w9151_ ;
	wire _w9150_ ;
	wire _w9149_ ;
	wire _w9148_ ;
	wire _w9147_ ;
	wire _w9146_ ;
	wire _w9145_ ;
	wire _w9144_ ;
	wire _w9143_ ;
	wire _w9142_ ;
	wire _w9141_ ;
	wire _w9140_ ;
	wire _w9139_ ;
	wire _w9138_ ;
	wire _w9137_ ;
	wire _w9136_ ;
	wire _w9135_ ;
	wire _w9134_ ;
	wire _w9133_ ;
	wire _w9132_ ;
	wire _w9131_ ;
	wire _w9130_ ;
	wire _w9129_ ;
	wire _w9128_ ;
	wire _w9127_ ;
	wire _w9126_ ;
	wire _w9125_ ;
	wire _w9124_ ;
	wire _w9123_ ;
	wire _w9122_ ;
	wire _w9121_ ;
	wire _w9120_ ;
	wire _w9119_ ;
	wire _w9118_ ;
	wire _w9117_ ;
	wire _w9116_ ;
	wire _w9115_ ;
	wire _w9114_ ;
	wire _w9113_ ;
	wire _w9112_ ;
	wire _w9111_ ;
	wire _w9110_ ;
	wire _w9109_ ;
	wire _w9108_ ;
	wire _w9107_ ;
	wire _w9106_ ;
	wire _w9105_ ;
	wire _w9104_ ;
	wire _w9103_ ;
	wire _w9102_ ;
	wire _w9101_ ;
	wire _w9100_ ;
	wire _w9099_ ;
	wire _w9098_ ;
	wire _w9097_ ;
	wire _w9096_ ;
	wire _w9095_ ;
	wire _w9094_ ;
	wire _w9093_ ;
	wire _w9092_ ;
	wire _w9091_ ;
	wire _w9090_ ;
	wire _w9089_ ;
	wire _w9088_ ;
	wire _w9087_ ;
	wire _w9086_ ;
	wire _w9085_ ;
	wire _w9084_ ;
	wire _w9083_ ;
	wire _w9082_ ;
	wire _w9081_ ;
	wire _w9080_ ;
	wire _w9079_ ;
	wire _w9078_ ;
	wire _w9077_ ;
	wire _w9076_ ;
	wire _w9075_ ;
	wire _w9074_ ;
	wire _w9073_ ;
	wire _w9072_ ;
	wire _w9071_ ;
	wire _w9070_ ;
	wire _w9069_ ;
	wire _w9068_ ;
	wire _w9067_ ;
	wire _w9066_ ;
	wire _w9065_ ;
	wire _w9064_ ;
	wire _w9063_ ;
	wire _w9062_ ;
	wire _w9061_ ;
	wire _w9060_ ;
	wire _w9059_ ;
	wire _w9058_ ;
	wire _w9057_ ;
	wire _w9056_ ;
	wire _w9055_ ;
	wire _w9054_ ;
	wire _w9053_ ;
	wire _w9052_ ;
	wire _w9051_ ;
	wire _w9050_ ;
	wire _w9049_ ;
	wire _w9048_ ;
	wire _w9047_ ;
	wire _w9046_ ;
	wire _w9045_ ;
	wire _w9044_ ;
	wire _w9043_ ;
	wire _w9042_ ;
	wire _w9041_ ;
	wire _w9040_ ;
	wire _w9039_ ;
	wire _w9038_ ;
	wire _w9037_ ;
	wire _w9036_ ;
	wire _w9035_ ;
	wire _w9034_ ;
	wire _w9033_ ;
	wire _w9032_ ;
	wire _w9031_ ;
	wire _w9030_ ;
	wire _w9029_ ;
	wire _w9028_ ;
	wire _w9027_ ;
	wire _w9026_ ;
	wire _w9025_ ;
	wire _w9024_ ;
	wire _w9023_ ;
	wire _w9022_ ;
	wire _w9021_ ;
	wire _w9020_ ;
	wire _w9019_ ;
	wire _w9018_ ;
	wire _w9017_ ;
	wire _w9016_ ;
	wire _w9015_ ;
	wire _w9014_ ;
	wire _w9013_ ;
	wire _w9012_ ;
	wire _w9011_ ;
	wire _w9010_ ;
	wire _w9009_ ;
	wire _w9008_ ;
	wire _w9007_ ;
	wire _w9006_ ;
	wire _w9005_ ;
	wire _w9004_ ;
	wire _w9003_ ;
	wire _w9002_ ;
	wire _w9001_ ;
	wire _w9000_ ;
	wire _w8999_ ;
	wire _w8998_ ;
	wire _w8997_ ;
	wire _w8996_ ;
	wire _w8995_ ;
	wire _w8994_ ;
	wire _w8993_ ;
	wire _w8992_ ;
	wire _w8991_ ;
	wire _w8990_ ;
	wire _w8989_ ;
	wire _w8988_ ;
	wire _w8987_ ;
	wire _w8986_ ;
	wire _w8985_ ;
	wire _w8984_ ;
	wire _w8983_ ;
	wire _w8982_ ;
	wire _w8981_ ;
	wire _w8980_ ;
	wire _w8979_ ;
	wire _w8978_ ;
	wire _w8977_ ;
	wire _w8976_ ;
	wire _w8975_ ;
	wire _w8974_ ;
	wire _w8973_ ;
	wire _w8972_ ;
	wire _w8971_ ;
	wire _w8970_ ;
	wire _w8969_ ;
	wire _w8968_ ;
	wire _w8967_ ;
	wire _w8966_ ;
	wire _w8965_ ;
	wire _w8964_ ;
	wire _w8963_ ;
	wire _w8962_ ;
	wire _w8961_ ;
	wire _w8960_ ;
	wire _w8959_ ;
	wire _w8958_ ;
	wire _w8957_ ;
	wire _w8956_ ;
	wire _w8955_ ;
	wire _w8954_ ;
	wire _w8953_ ;
	wire _w8952_ ;
	wire _w8951_ ;
	wire _w8950_ ;
	wire _w8949_ ;
	wire _w8948_ ;
	wire _w8947_ ;
	wire _w8946_ ;
	wire _w8945_ ;
	wire _w8944_ ;
	wire _w8943_ ;
	wire _w8942_ ;
	wire _w8941_ ;
	wire _w8940_ ;
	wire _w8939_ ;
	wire _w8938_ ;
	wire _w8937_ ;
	wire _w8936_ ;
	wire _w8935_ ;
	wire _w8934_ ;
	wire _w8933_ ;
	wire _w8932_ ;
	wire _w8931_ ;
	wire _w8930_ ;
	wire _w8929_ ;
	wire _w8928_ ;
	wire _w8927_ ;
	wire _w8926_ ;
	wire _w8925_ ;
	wire _w8924_ ;
	wire _w8923_ ;
	wire _w8922_ ;
	wire _w8921_ ;
	wire _w8920_ ;
	wire _w8919_ ;
	wire _w8918_ ;
	wire _w8917_ ;
	wire _w8916_ ;
	wire _w8915_ ;
	wire _w8914_ ;
	wire _w8913_ ;
	wire _w8912_ ;
	wire _w8911_ ;
	wire _w8910_ ;
	wire _w8909_ ;
	wire _w8908_ ;
	wire _w8907_ ;
	wire _w8906_ ;
	wire _w8905_ ;
	wire _w8904_ ;
	wire _w8903_ ;
	wire _w8902_ ;
	wire _w8901_ ;
	wire _w8900_ ;
	wire _w8899_ ;
	wire _w8898_ ;
	wire _w8897_ ;
	wire _w8896_ ;
	wire _w8895_ ;
	wire _w8894_ ;
	wire _w8893_ ;
	wire _w8892_ ;
	wire _w8891_ ;
	wire _w8890_ ;
	wire _w8889_ ;
	wire _w8888_ ;
	wire _w8887_ ;
	wire _w8886_ ;
	wire _w8885_ ;
	wire _w8884_ ;
	wire _w8883_ ;
	wire _w8882_ ;
	wire _w8881_ ;
	wire _w8880_ ;
	wire _w8879_ ;
	wire _w8878_ ;
	wire _w8877_ ;
	wire _w8876_ ;
	wire _w8875_ ;
	wire _w8874_ ;
	wire _w8873_ ;
	wire _w8872_ ;
	wire _w8871_ ;
	wire _w8870_ ;
	wire _w8869_ ;
	wire _w8868_ ;
	wire _w8867_ ;
	wire _w8866_ ;
	wire _w8865_ ;
	wire _w8864_ ;
	wire _w8863_ ;
	wire _w8862_ ;
	wire _w8861_ ;
	wire _w8860_ ;
	wire _w8859_ ;
	wire _w8858_ ;
	wire _w8857_ ;
	wire _w8856_ ;
	wire _w8855_ ;
	wire _w8854_ ;
	wire _w8853_ ;
	wire _w8852_ ;
	wire _w8851_ ;
	wire _w8850_ ;
	wire _w8849_ ;
	wire _w8848_ ;
	wire _w8847_ ;
	wire _w8846_ ;
	wire _w8845_ ;
	wire _w8844_ ;
	wire _w8843_ ;
	wire _w8842_ ;
	wire _w8841_ ;
	wire _w8840_ ;
	wire _w8839_ ;
	wire _w8838_ ;
	wire _w8837_ ;
	wire _w8836_ ;
	wire _w8835_ ;
	wire _w8834_ ;
	wire _w8833_ ;
	wire _w8832_ ;
	wire _w8831_ ;
	wire _w8830_ ;
	wire _w8829_ ;
	wire _w8828_ ;
	wire _w8827_ ;
	wire _w8826_ ;
	wire _w8825_ ;
	wire _w8824_ ;
	wire _w8823_ ;
	wire _w8822_ ;
	wire _w8821_ ;
	wire _w8820_ ;
	wire _w8819_ ;
	wire _w8818_ ;
	wire _w8817_ ;
	wire _w8816_ ;
	wire _w8815_ ;
	wire _w8814_ ;
	wire _w8813_ ;
	wire _w8812_ ;
	wire _w8811_ ;
	wire _w8810_ ;
	wire _w8809_ ;
	wire _w8808_ ;
	wire _w8807_ ;
	wire _w8806_ ;
	wire _w8805_ ;
	wire _w8804_ ;
	wire _w8803_ ;
	wire _w8802_ ;
	wire _w8801_ ;
	wire _w8800_ ;
	wire _w8799_ ;
	wire _w8798_ ;
	wire _w8797_ ;
	wire _w8796_ ;
	wire _w8795_ ;
	wire _w8794_ ;
	wire _w8793_ ;
	wire _w8792_ ;
	wire _w8791_ ;
	wire _w8790_ ;
	wire _w8789_ ;
	wire _w8788_ ;
	wire _w8787_ ;
	wire _w8786_ ;
	wire _w8785_ ;
	wire _w8784_ ;
	wire _w8783_ ;
	wire _w8782_ ;
	wire _w8781_ ;
	wire _w8780_ ;
	wire _w8779_ ;
	wire _w8778_ ;
	wire _w8777_ ;
	wire _w8776_ ;
	wire _w8775_ ;
	wire _w8774_ ;
	wire _w8773_ ;
	wire _w8772_ ;
	wire _w8771_ ;
	wire _w8770_ ;
	wire _w8769_ ;
	wire _w8768_ ;
	wire _w8767_ ;
	wire _w8766_ ;
	wire _w8765_ ;
	wire _w8764_ ;
	wire _w8763_ ;
	wire _w8762_ ;
	wire _w8761_ ;
	wire _w8760_ ;
	wire _w8759_ ;
	wire _w8758_ ;
	wire _w8757_ ;
	wire _w8756_ ;
	wire _w8755_ ;
	wire _w8754_ ;
	wire _w8753_ ;
	wire _w8752_ ;
	wire _w8751_ ;
	wire _w8750_ ;
	wire _w8749_ ;
	wire _w8748_ ;
	wire _w8747_ ;
	wire _w8746_ ;
	wire _w8745_ ;
	wire _w8744_ ;
	wire _w8743_ ;
	wire _w8742_ ;
	wire _w8741_ ;
	wire _w8740_ ;
	wire _w8739_ ;
	wire _w8738_ ;
	wire _w8737_ ;
	wire _w8736_ ;
	wire _w8735_ ;
	wire _w8734_ ;
	wire _w8733_ ;
	wire _w8732_ ;
	wire _w8731_ ;
	wire _w8730_ ;
	wire _w8729_ ;
	wire _w8728_ ;
	wire _w8727_ ;
	wire _w8726_ ;
	wire _w8725_ ;
	wire _w8724_ ;
	wire _w8723_ ;
	wire _w8722_ ;
	wire _w8721_ ;
	wire _w8720_ ;
	wire _w8719_ ;
	wire _w8718_ ;
	wire _w8717_ ;
	wire _w8716_ ;
	wire _w8715_ ;
	wire _w8714_ ;
	wire _w8713_ ;
	wire _w8712_ ;
	wire _w8711_ ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2616_ ;
	wire _w2615_ ;
	wire _w2614_ ;
	wire _w2613_ ;
	wire _w2612_ ;
	wire _w2611_ ;
	wire _w2610_ ;
	wire _w2609_ ;
	wire _w2608_ ;
	wire _w2607_ ;
	wire _w2606_ ;
	wire _w2605_ ;
	wire _w2604_ ;
	wire _w2603_ ;
	wire _w2602_ ;
	wire _w2601_ ;
	wire _w2600_ ;
	wire _w2599_ ;
	wire _w2598_ ;
	wire _w2597_ ;
	wire _w2596_ ;
	wire _w2595_ ;
	wire _w2594_ ;
	wire _w2593_ ;
	wire _w2592_ ;
	wire _w2591_ ;
	wire _w2590_ ;
	wire _w2589_ ;
	wire _w2588_ ;
	wire _w2587_ ;
	wire _w2586_ ;
	wire _w2585_ ;
	wire _w2584_ ;
	wire _w2583_ ;
	wire _w2582_ ;
	wire _w2581_ ;
	wire _w2580_ ;
	wire _w2579_ ;
	wire _w2578_ ;
	wire _w2577_ ;
	wire _w2576_ ;
	wire _w2575_ ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2690_ ;
	wire _w2691_ ;
	wire _w2692_ ;
	wire _w2693_ ;
	wire _w2694_ ;
	wire _w2695_ ;
	wire _w2696_ ;
	wire _w2697_ ;
	wire _w2698_ ;
	wire _w2699_ ;
	wire _w2700_ ;
	wire _w2701_ ;
	wire _w2702_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2776_ ;
	wire _w2777_ ;
	wire _w2778_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2898_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2901_ ;
	wire _w2902_ ;
	wire _w2903_ ;
	wire _w2904_ ;
	wire _w2905_ ;
	wire _w2906_ ;
	wire _w2907_ ;
	wire _w2908_ ;
	wire _w2909_ ;
	wire _w2910_ ;
	wire _w2911_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2914_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2993_ ;
	wire _w2994_ ;
	wire _w2995_ ;
	wire _w2996_ ;
	wire _w2997_ ;
	wire _w2998_ ;
	wire _w2999_ ;
	wire _w3000_ ;
	wire _w3001_ ;
	wire _w3002_ ;
	wire _w3003_ ;
	wire _w3004_ ;
	wire _w3005_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3072_ ;
	wire _w3073_ ;
	wire _w3074_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3177_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3195_ ;
	wire _w3196_ ;
	wire _w3197_ ;
	wire _w3198_ ;
	wire _w3199_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3202_ ;
	wire _w3203_ ;
	wire _w3204_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3210_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3217_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	wire _w6595_ ;
	wire _w6596_ ;
	wire _w6597_ ;
	wire _w6598_ ;
	wire _w6599_ ;
	wire _w6600_ ;
	wire _w6601_ ;
	wire _w6602_ ;
	wire _w6603_ ;
	wire _w6604_ ;
	wire _w6605_ ;
	wire _w6606_ ;
	wire _w6607_ ;
	wire _w6608_ ;
	wire _w6609_ ;
	wire _w6610_ ;
	wire _w6611_ ;
	wire _w6612_ ;
	wire _w6613_ ;
	wire _w6614_ ;
	wire _w6615_ ;
	wire _w6616_ ;
	wire _w6617_ ;
	wire _w6618_ ;
	wire _w6619_ ;
	wire _w6620_ ;
	wire _w6621_ ;
	wire _w6622_ ;
	wire _w6623_ ;
	wire _w6624_ ;
	wire _w6625_ ;
	wire _w6626_ ;
	wire _w6627_ ;
	wire _w6628_ ;
	wire _w6629_ ;
	wire _w6630_ ;
	wire _w6631_ ;
	wire _w6632_ ;
	wire _w6633_ ;
	wire _w6634_ ;
	wire _w6635_ ;
	wire _w6636_ ;
	wire _w6637_ ;
	wire _w6638_ ;
	wire _w6639_ ;
	wire _w6640_ ;
	wire _w6641_ ;
	wire _w6642_ ;
	wire _w6643_ ;
	wire _w6644_ ;
	wire _w6645_ ;
	wire _w6646_ ;
	wire _w6647_ ;
	wire _w6648_ ;
	wire _w6649_ ;
	wire _w6650_ ;
	wire _w6651_ ;
	wire _w6652_ ;
	wire _w6653_ ;
	wire _w6654_ ;
	wire _w6655_ ;
	wire _w6656_ ;
	wire _w6657_ ;
	wire _w6658_ ;
	wire _w6659_ ;
	wire _w6660_ ;
	wire _w6661_ ;
	wire _w6662_ ;
	wire _w6663_ ;
	wire _w6664_ ;
	wire _w6665_ ;
	wire _w6666_ ;
	wire _w6667_ ;
	wire _w6668_ ;
	wire _w6669_ ;
	wire _w6670_ ;
	wire _w6671_ ;
	wire _w6672_ ;
	wire _w6673_ ;
	wire _w6674_ ;
	wire _w6675_ ;
	wire _w6676_ ;
	wire _w6677_ ;
	wire _w6678_ ;
	wire _w6679_ ;
	wire _w6680_ ;
	wire _w6681_ ;
	wire _w6682_ ;
	wire _w6683_ ;
	wire _w6684_ ;
	wire _w6685_ ;
	wire _w6686_ ;
	wire _w6687_ ;
	wire _w6688_ ;
	wire _w6689_ ;
	wire _w6690_ ;
	wire _w6691_ ;
	wire _w6692_ ;
	wire _w6693_ ;
	wire _w6694_ ;
	wire _w6695_ ;
	wire _w6696_ ;
	wire _w6697_ ;
	wire _w6698_ ;
	wire _w6699_ ;
	wire _w6700_ ;
	wire _w6701_ ;
	wire _w6702_ ;
	wire _w6703_ ;
	wire _w6704_ ;
	wire _w6705_ ;
	wire _w6706_ ;
	wire _w6707_ ;
	wire _w6708_ ;
	wire _w6709_ ;
	wire _w6710_ ;
	wire _w6711_ ;
	wire _w6712_ ;
	wire _w6713_ ;
	wire _w6714_ ;
	wire _w6715_ ;
	wire _w6716_ ;
	wire _w6717_ ;
	wire _w6718_ ;
	wire _w6719_ ;
	wire _w6720_ ;
	wire _w6721_ ;
	wire _w6722_ ;
	wire _w6723_ ;
	wire _w6724_ ;
	wire _w6725_ ;
	wire _w6726_ ;
	wire _w6727_ ;
	wire _w6728_ ;
	wire _w6729_ ;
	wire _w6730_ ;
	wire _w6731_ ;
	wire _w6732_ ;
	wire _w6733_ ;
	wire _w6734_ ;
	wire _w6735_ ;
	wire _w6736_ ;
	wire _w6737_ ;
	wire _w6738_ ;
	wire _w6739_ ;
	wire _w6740_ ;
	wire _w6741_ ;
	wire _w6742_ ;
	wire _w6743_ ;
	wire _w6744_ ;
	wire _w6745_ ;
	wire _w6746_ ;
	wire _w6747_ ;
	wire _w6748_ ;
	wire _w6749_ ;
	wire _w6750_ ;
	wire _w6751_ ;
	wire _w6752_ ;
	wire _w6753_ ;
	wire _w6754_ ;
	wire _w6755_ ;
	wire _w6756_ ;
	wire _w6757_ ;
	wire _w6758_ ;
	wire _w6759_ ;
	wire _w6760_ ;
	wire _w6761_ ;
	wire _w6762_ ;
	wire _w6763_ ;
	wire _w6764_ ;
	wire _w6765_ ;
	wire _w6766_ ;
	wire _w6767_ ;
	wire _w6768_ ;
	wire _w6769_ ;
	wire _w6770_ ;
	wire _w6771_ ;
	wire _w6772_ ;
	wire _w6773_ ;
	wire _w6774_ ;
	wire _w6775_ ;
	wire _w6776_ ;
	wire _w6777_ ;
	wire _w6778_ ;
	wire _w6779_ ;
	wire _w6780_ ;
	wire _w6781_ ;
	wire _w6782_ ;
	wire _w6783_ ;
	wire _w6784_ ;
	wire _w6785_ ;
	wire _w6786_ ;
	wire _w6787_ ;
	wire _w6788_ ;
	wire _w6789_ ;
	wire _w6790_ ;
	wire _w6791_ ;
	wire _w6792_ ;
	wire _w6793_ ;
	wire _w6794_ ;
	wire _w6795_ ;
	wire _w6796_ ;
	wire _w6797_ ;
	wire _w6798_ ;
	wire _w6799_ ;
	wire _w6800_ ;
	wire _w6801_ ;
	wire _w6802_ ;
	wire _w6803_ ;
	wire _w6804_ ;
	wire _w6805_ ;
	wire _w6806_ ;
	wire _w6807_ ;
	wire _w6808_ ;
	wire _w6809_ ;
	wire _w6810_ ;
	wire _w6811_ ;
	wire _w6812_ ;
	wire _w6813_ ;
	wire _w6814_ ;
	wire _w6815_ ;
	wire _w6816_ ;
	wire _w6817_ ;
	wire _w6818_ ;
	wire _w6819_ ;
	wire _w6820_ ;
	wire _w6821_ ;
	wire _w6822_ ;
	wire _w6823_ ;
	wire _w6824_ ;
	wire _w6825_ ;
	wire _w6826_ ;
	wire _w6827_ ;
	wire _w6828_ ;
	wire _w6829_ ;
	wire _w6830_ ;
	wire _w6831_ ;
	wire _w6832_ ;
	wire _w6833_ ;
	wire _w6834_ ;
	wire _w6835_ ;
	wire _w6836_ ;
	wire _w6837_ ;
	wire _w6838_ ;
	wire _w6839_ ;
	wire _w6840_ ;
	wire _w6841_ ;
	wire _w6842_ ;
	wire _w6843_ ;
	wire _w6844_ ;
	wire _w6845_ ;
	wire _w6846_ ;
	wire _w6847_ ;
	wire _w6848_ ;
	wire _w6849_ ;
	wire _w6850_ ;
	wire _w6851_ ;
	wire _w6852_ ;
	wire _w6853_ ;
	wire _w6854_ ;
	wire _w6855_ ;
	wire _w6856_ ;
	wire _w6857_ ;
	wire _w6858_ ;
	wire _w6859_ ;
	wire _w6860_ ;
	wire _w6861_ ;
	wire _w6862_ ;
	wire _w6863_ ;
	wire _w6864_ ;
	wire _w6865_ ;
	wire _w6866_ ;
	wire _w6867_ ;
	wire _w6868_ ;
	wire _w6869_ ;
	wire _w6870_ ;
	wire _w6871_ ;
	wire _w6872_ ;
	wire _w6873_ ;
	wire _w6874_ ;
	wire _w6875_ ;
	wire _w6876_ ;
	wire _w6877_ ;
	wire _w6878_ ;
	wire _w6879_ ;
	wire _w6880_ ;
	wire _w6881_ ;
	wire _w6882_ ;
	wire _w6883_ ;
	wire _w6884_ ;
	wire _w6885_ ;
	wire _w6886_ ;
	wire _w6887_ ;
	wire _w6888_ ;
	wire _w6889_ ;
	wire _w6890_ ;
	wire _w6891_ ;
	wire _w6892_ ;
	wire _w6893_ ;
	wire _w6894_ ;
	wire _w6895_ ;
	wire _w6896_ ;
	wire _w6897_ ;
	wire _w6898_ ;
	wire _w6899_ ;
	wire _w6900_ ;
	wire _w6901_ ;
	wire _w6902_ ;
	wire _w6903_ ;
	wire _w6904_ ;
	wire _w6905_ ;
	wire _w6906_ ;
	wire _w6907_ ;
	wire _w6908_ ;
	wire _w6909_ ;
	wire _w6910_ ;
	wire _w6911_ ;
	wire _w6912_ ;
	wire _w6913_ ;
	wire _w6914_ ;
	wire _w6915_ ;
	wire _w6916_ ;
	wire _w6917_ ;
	wire _w6918_ ;
	wire _w6919_ ;
	wire _w6920_ ;
	wire _w6921_ ;
	wire _w6922_ ;
	wire _w6923_ ;
	wire _w6924_ ;
	wire _w6925_ ;
	wire _w6926_ ;
	wire _w6927_ ;
	wire _w6928_ ;
	wire _w6929_ ;
	wire _w6930_ ;
	wire _w6931_ ;
	wire _w6932_ ;
	wire _w6933_ ;
	wire _w6934_ ;
	wire _w6935_ ;
	wire _w6936_ ;
	wire _w6937_ ;
	wire _w6938_ ;
	wire _w6939_ ;
	wire _w6940_ ;
	wire _w6941_ ;
	wire _w6942_ ;
	wire _w6943_ ;
	wire _w6944_ ;
	wire _w6945_ ;
	wire _w6946_ ;
	wire _w6947_ ;
	wire _w6948_ ;
	wire _w6949_ ;
	wire _w6950_ ;
	wire _w6951_ ;
	wire _w6952_ ;
	wire _w6953_ ;
	wire _w6954_ ;
	wire _w6955_ ;
	wire _w6956_ ;
	wire _w6957_ ;
	wire _w6958_ ;
	wire _w6959_ ;
	wire _w6960_ ;
	wire _w6961_ ;
	wire _w6962_ ;
	wire _w6963_ ;
	wire _w6964_ ;
	wire _w6965_ ;
	wire _w6966_ ;
	wire _w6967_ ;
	wire _w6968_ ;
	wire _w6969_ ;
	wire _w6970_ ;
	wire _w6971_ ;
	wire _w6972_ ;
	wire _w6973_ ;
	wire _w6974_ ;
	wire _w6975_ ;
	wire _w6976_ ;
	wire _w6977_ ;
	wire _w6978_ ;
	wire _w6979_ ;
	wire _w6980_ ;
	wire _w6981_ ;
	wire _w6982_ ;
	wire _w6983_ ;
	wire _w6984_ ;
	wire _w6985_ ;
	wire _w6986_ ;
	wire _w6987_ ;
	wire _w6988_ ;
	wire _w6989_ ;
	wire _w6990_ ;
	wire _w6991_ ;
	wire _w6992_ ;
	wire _w6993_ ;
	wire _w6994_ ;
	wire _w6995_ ;
	wire _w6996_ ;
	wire _w6997_ ;
	wire _w6998_ ;
	wire _w6999_ ;
	wire _w7000_ ;
	wire _w7001_ ;
	wire _w7002_ ;
	wire _w7003_ ;
	wire _w7004_ ;
	wire _w7005_ ;
	wire _w7006_ ;
	wire _w7007_ ;
	wire _w7008_ ;
	wire _w7009_ ;
	wire _w7010_ ;
	wire _w7011_ ;
	wire _w7012_ ;
	wire _w7013_ ;
	wire _w7014_ ;
	wire _w7015_ ;
	wire _w7016_ ;
	wire _w7017_ ;
	wire _w7018_ ;
	wire _w7019_ ;
	wire _w7020_ ;
	wire _w7021_ ;
	wire _w7022_ ;
	wire _w7023_ ;
	wire _w7024_ ;
	wire _w7025_ ;
	wire _w7026_ ;
	wire _w7027_ ;
	wire _w7028_ ;
	wire _w7029_ ;
	wire _w7030_ ;
	wire _w7031_ ;
	wire _w7032_ ;
	wire _w7033_ ;
	wire _w7034_ ;
	wire _w7035_ ;
	wire _w7036_ ;
	wire _w7037_ ;
	wire _w7038_ ;
	wire _w7039_ ;
	wire _w7040_ ;
	wire _w7041_ ;
	wire _w7042_ ;
	wire _w7043_ ;
	wire _w7044_ ;
	wire _w7045_ ;
	wire _w7046_ ;
	wire _w7047_ ;
	wire _w7048_ ;
	wire _w7049_ ;
	wire _w7050_ ;
	wire _w7051_ ;
	wire _w7052_ ;
	wire _w7053_ ;
	wire _w7054_ ;
	wire _w7055_ ;
	wire _w7056_ ;
	wire _w7057_ ;
	wire _w7058_ ;
	wire _w7059_ ;
	wire _w7060_ ;
	wire _w7061_ ;
	wire _w7062_ ;
	wire _w7063_ ;
	wire _w7064_ ;
	wire _w7065_ ;
	wire _w7066_ ;
	wire _w7067_ ;
	wire _w7068_ ;
	wire _w7069_ ;
	wire _w7070_ ;
	wire _w7071_ ;
	wire _w7072_ ;
	wire _w7073_ ;
	wire _w7074_ ;
	wire _w7075_ ;
	wire _w7076_ ;
	wire _w7077_ ;
	wire _w7078_ ;
	wire _w7079_ ;
	wire _w7080_ ;
	wire _w7081_ ;
	wire _w7082_ ;
	wire _w7083_ ;
	wire _w7084_ ;
	wire _w7085_ ;
	wire _w7086_ ;
	wire _w7087_ ;
	wire _w7088_ ;
	wire _w7089_ ;
	wire _w7090_ ;
	wire _w7091_ ;
	wire _w7092_ ;
	wire _w7093_ ;
	wire _w7094_ ;
	wire _w7095_ ;
	wire _w7096_ ;
	wire _w7097_ ;
	wire _w7098_ ;
	wire _w7099_ ;
	wire _w7100_ ;
	wire _w7101_ ;
	wire _w7102_ ;
	wire _w7103_ ;
	wire _w7104_ ;
	wire _w7105_ ;
	wire _w7106_ ;
	wire _w7107_ ;
	wire _w7108_ ;
	wire _w7109_ ;
	wire _w7110_ ;
	wire _w7111_ ;
	wire _w7112_ ;
	wire _w7113_ ;
	wire _w7114_ ;
	wire _w7115_ ;
	wire _w7116_ ;
	wire _w7117_ ;
	wire _w7118_ ;
	wire _w7119_ ;
	wire _w7120_ ;
	wire _w7121_ ;
	wire _w7122_ ;
	wire _w7123_ ;
	wire _w7124_ ;
	wire _w7125_ ;
	wire _w7126_ ;
	wire _w7127_ ;
	wire _w7128_ ;
	wire _w7129_ ;
	wire _w7130_ ;
	wire _w7131_ ;
	wire _w7132_ ;
	wire _w7133_ ;
	wire _w7134_ ;
	wire _w7135_ ;
	wire _w7136_ ;
	wire _w7137_ ;
	wire _w7138_ ;
	wire _w7139_ ;
	wire _w7140_ ;
	wire _w7141_ ;
	wire _w7142_ ;
	wire _w7143_ ;
	wire _w7144_ ;
	wire _w7145_ ;
	wire _w7146_ ;
	wire _w7147_ ;
	wire _w7148_ ;
	wire _w7149_ ;
	wire _w7150_ ;
	wire _w7151_ ;
	wire _w7152_ ;
	wire _w7153_ ;
	wire _w7154_ ;
	wire _w7155_ ;
	wire _w7156_ ;
	wire _w7157_ ;
	wire _w7158_ ;
	wire _w7159_ ;
	wire _w7160_ ;
	wire _w7161_ ;
	wire _w7162_ ;
	wire _w7163_ ;
	wire _w7164_ ;
	wire _w7165_ ;
	wire _w7166_ ;
	wire _w7167_ ;
	wire _w7168_ ;
	wire _w7169_ ;
	wire _w7170_ ;
	wire _w7171_ ;
	wire _w7172_ ;
	wire _w7173_ ;
	wire _w7174_ ;
	wire _w7175_ ;
	wire _w7176_ ;
	wire _w7177_ ;
	wire _w7178_ ;
	wire _w7179_ ;
	wire _w7180_ ;
	wire _w7181_ ;
	wire _w7182_ ;
	wire _w7183_ ;
	wire _w7184_ ;
	wire _w7185_ ;
	wire _w7186_ ;
	wire _w7187_ ;
	wire _w7188_ ;
	wire _w7189_ ;
	wire _w7190_ ;
	wire _w7191_ ;
	wire _w7192_ ;
	wire _w7193_ ;
	wire _w7194_ ;
	wire _w7195_ ;
	wire _w7196_ ;
	wire _w7197_ ;
	wire _w7198_ ;
	wire _w7199_ ;
	wire _w7200_ ;
	wire _w7201_ ;
	wire _w7202_ ;
	wire _w7203_ ;
	wire _w7204_ ;
	wire _w7205_ ;
	wire _w7206_ ;
	wire _w7207_ ;
	wire _w7208_ ;
	wire _w7209_ ;
	wire _w7210_ ;
	wire _w7211_ ;
	wire _w7212_ ;
	wire _w7213_ ;
	wire _w7214_ ;
	wire _w7215_ ;
	wire _w7216_ ;
	wire _w7217_ ;
	wire _w7218_ ;
	wire _w7219_ ;
	wire _w7220_ ;
	wire _w7221_ ;
	wire _w7222_ ;
	wire _w7223_ ;
	wire _w7224_ ;
	wire _w7225_ ;
	wire _w7226_ ;
	wire _w7227_ ;
	wire _w7228_ ;
	wire _w7229_ ;
	wire _w7230_ ;
	wire _w7231_ ;
	wire _w7232_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\dma_ack_i[8]_pad ,
		\dma_req_o[8]_pad ,
		_w2146_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\u11_status_reg[1]/P0001 ,
		\u13_icc_r_reg[21]/NET0131 ,
		_w2147_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\u11_status_reg[0]/P0001 ,
		\u13_icc_r_reg[20]/NET0131 ,
		_w2148_
	);
	LUT2 #(
		.INIT('h4)
	) name3 (
		_w2147_,
		_w2148_,
		_w2149_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\u11_status_reg[1]/P0001 ,
		\u13_icc_r_reg[21]/NET0131 ,
		_w2150_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		\u11_full_reg/NET0131 ,
		_w2150_,
		_w2151_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		_w2149_,
		_w2151_,
		_w2152_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w2152_,
		_w2153_
	);
	LUT2 #(
		.INIT('h4)
	) name8 (
		\dma_ack_i[8]_pad ,
		\u13_icc_r_reg[22]/NET0131 ,
		_w2154_
	);
	LUT2 #(
		.INIT('h8)
	) name9 (
		_w2153_,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\u16_u8_dma_req_r1_reg/P0001 ,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w2146_,
		_w2156_,
		_w2157_
	);
	LUT2 #(
		.INIT('h8)
	) name12 (
		\u14_u5_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2158_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\u14_u5_en_out_l2_reg/P0001 ,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h1)
	) name14 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\u13_occ1_r_reg[11]/NET0131 ,
		_w2160_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		\u8_rp_reg[0]/P0001 ,
		_w2160_,
		_w2161_
	);
	LUT2 #(
		.INIT('h2)
	) name16 (
		_w2159_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h8)
	) name17 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w2163_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		_w2162_,
		_w2163_,
		_w2164_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		\u8_rp_reg[3]/NET0131 ,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		\u8_rp_reg[3]/NET0131 ,
		_w2164_,
		_w2166_
	);
	LUT2 #(
		.INIT('h2)
	) name21 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2165_,
		_w2167_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w2166_,
		_w2167_,
		_w2168_
	);
	LUT2 #(
		.INIT('h1)
	) name23 (
		\u0_slt0_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2169_
	);
	LUT2 #(
		.INIT('h4)
	) name24 (
		\u14_crac_wr_r_reg/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2170_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\u14_crac_valid_r_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		\u14_u1_en_out_l_reg/NET0131 ,
		\u14_u2_en_out_l_reg/NET0131 ,
		_w2172_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		\u14_u3_en_out_l_reg/NET0131 ,
		\u14_u4_en_out_l_reg/NET0131 ,
		_w2173_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\u14_u5_en_out_l_reg/NET0131 ,
		_w2173_,
		_w2174_
	);
	LUT2 #(
		.INIT('h8)
	) name29 (
		_w2171_,
		_w2172_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w2170_,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('h8)
	) name31 (
		_w2174_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w2169_,
		_w2177_,
		_w2178_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		\u14_crac_valid_r_reg/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2179_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\u0_slt0_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2180_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w2179_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		\u0_slt0_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2182_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w2170_,
		_w2182_,
		_w2183_
	);
	LUT2 #(
		.INIT('h2)
	) name38 (
		\u0_slt0_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2184_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		\u14_u0_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2185_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w2184_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		\u14_u1_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2187_
	);
	LUT2 #(
		.INIT('h2)
	) name42 (
		\u0_slt0_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2188_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w2187_,
		_w2188_,
		_w2189_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\u0_slt0_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2190_
	);
	LUT2 #(
		.INIT('h8)
	) name45 (
		\u14_u2_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2191_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		\u0_slt0_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2192_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w2191_,
		_w2192_,
		_w2193_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		\u14_u3_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2194_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		\u0_slt0_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2195_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w2194_,
		_w2195_,
		_w2196_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		\u14_u4_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2197_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\u0_slt0_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2198_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w2197_,
		_w2198_,
		_w2199_
	);
	LUT2 #(
		.INIT('h2)
	) name54 (
		\u0_slt0_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2200_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		\u14_u5_en_out_l_reg/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2201_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w2200_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\u0_slt0_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2203_
	);
	LUT2 #(
		.INIT('h2)
	) name58 (
		\u0_slt0_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2204_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		\u0_slt0_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2205_
	);
	LUT2 #(
		.INIT('h2)
	) name60 (
		\u0_slt0_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2206_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\u0_slt0_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2207_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\u0_slt1_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2208_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\u13_crac_r_reg[7]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2209_
	);
	LUT2 #(
		.INIT('h2)
	) name64 (
		\u0_slt1_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2210_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		_w2209_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\u13_crac_r_reg[6]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2212_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\u0_slt1_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2213_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w2212_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\u13_crac_r_reg[5]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2215_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\u0_slt1_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2216_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w2215_,
		_w2216_,
		_w2217_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		\u13_crac_r_reg[4]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2218_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\u0_slt1_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2219_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w2218_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		\u13_crac_r_reg[3]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2221_
	);
	LUT2 #(
		.INIT('h2)
	) name76 (
		\u0_slt1_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2222_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		\u13_crac_r_reg[2]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2224_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\u0_slt1_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2225_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w2224_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\u13_crac_r_reg[1]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2227_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\u0_slt1_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2228_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w2227_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h8)
	) name84 (
		\u13_crac_r_reg[0]/NET0131 ,
		\u2_ld_reg/P0001 ,
		_w2230_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		\u0_slt1_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2231_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w2230_,
		_w2231_,
		_w2232_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		\u0_slt1_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2233_
	);
	LUT2 #(
		.INIT('h2)
	) name88 (
		\u0_slt1_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2234_
	);
	LUT2 #(
		.INIT('h2)
	) name89 (
		\u0_slt1_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2235_
	);
	LUT2 #(
		.INIT('h2)
	) name90 (
		\u0_slt1_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2236_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\u0_slt1_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2237_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\u0_slt1_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2238_
	);
	LUT2 #(
		.INIT('h2)
	) name93 (
		\u0_slt1_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		\u0_slt1_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2240_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\u0_slt1_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2241_
	);
	LUT2 #(
		.INIT('h2)
	) name96 (
		\u0_slt1_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2242_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\u0_slt1_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2243_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\u0_slt2_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2244_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\u13_crac_dout_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2245_
	);
	LUT2 #(
		.INIT('h2)
	) name100 (
		\u0_slt2_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2246_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w2245_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\u13_crac_dout_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2248_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		\u0_slt2_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2249_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w2248_,
		_w2249_,
		_w2250_
	);
	LUT2 #(
		.INIT('h8)
	) name105 (
		\u13_crac_dout_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2251_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		\u0_slt2_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2252_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w2251_,
		_w2252_,
		_w2253_
	);
	LUT2 #(
		.INIT('h8)
	) name108 (
		\u13_crac_dout_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2254_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		\u0_slt2_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2255_
	);
	LUT2 #(
		.INIT('h1)
	) name110 (
		_w2254_,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h8)
	) name111 (
		\u13_crac_dout_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2257_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		\u0_slt2_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2258_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		_w2257_,
		_w2258_,
		_w2259_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\u13_crac_dout_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2260_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		\u0_slt2_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2261_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w2260_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h8)
	) name117 (
		\u13_crac_dout_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2263_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		\u0_slt2_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2264_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w2263_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		\u13_crac_dout_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2266_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		\u0_slt2_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2267_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w2266_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\u13_crac_dout_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2269_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		\u0_slt2_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2270_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w2269_,
		_w2270_,
		_w2271_
	);
	LUT2 #(
		.INIT('h8)
	) name126 (
		\u13_crac_dout_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2272_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		\u0_slt2_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2273_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\u13_crac_dout_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2275_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\u0_slt2_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2276_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w2275_,
		_w2276_,
		_w2277_
	);
	LUT2 #(
		.INIT('h8)
	) name132 (
		\u13_crac_dout_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2278_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		\u0_slt2_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name134 (
		_w2278_,
		_w2279_,
		_w2280_
	);
	LUT2 #(
		.INIT('h8)
	) name135 (
		\u13_crac_dout_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2281_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		\u0_slt2_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2282_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w2281_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\u13_crac_dout_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2284_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\u0_slt2_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2285_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		_w2284_,
		_w2285_,
		_w2286_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		\u13_crac_dout_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2287_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		\u0_slt2_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2288_
	);
	LUT2 #(
		.INIT('h1)
	) name143 (
		_w2287_,
		_w2288_,
		_w2289_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		\u13_crac_dout_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2290_
	);
	LUT2 #(
		.INIT('h2)
	) name145 (
		\u0_slt2_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2291_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		_w2290_,
		_w2291_,
		_w2292_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\u0_slt2_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2293_
	);
	LUT2 #(
		.INIT('h2)
	) name148 (
		\u0_slt2_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name149 (
		\u0_slt2_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2295_
	);
	LUT2 #(
		.INIT('h2)
	) name150 (
		\u0_slt3_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2296_
	);
	LUT2 #(
		.INIT('h8)
	) name151 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[19]/P0001 ,
		_w2297_
	);
	LUT2 #(
		.INIT('h2)
	) name152 (
		\u0_slt3_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2298_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w2297_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[18]/P0001 ,
		_w2300_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\u0_slt3_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w2300_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[17]/P0001 ,
		_w2303_
	);
	LUT2 #(
		.INIT('h2)
	) name158 (
		\u0_slt3_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2304_
	);
	LUT2 #(
		.INIT('h1)
	) name159 (
		_w2303_,
		_w2304_,
		_w2305_
	);
	LUT2 #(
		.INIT('h8)
	) name160 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[16]/P0001 ,
		_w2306_
	);
	LUT2 #(
		.INIT('h2)
	) name161 (
		\u0_slt3_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2307_
	);
	LUT2 #(
		.INIT('h1)
	) name162 (
		_w2306_,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[15]/P0001 ,
		_w2309_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		\u0_slt3_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2310_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w2309_,
		_w2310_,
		_w2311_
	);
	LUT2 #(
		.INIT('h8)
	) name166 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[14]/P0001 ,
		_w2312_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		\u0_slt3_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2313_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w2312_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[13]/P0001 ,
		_w2315_
	);
	LUT2 #(
		.INIT('h2)
	) name170 (
		\u0_slt3_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2316_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h8)
	) name172 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[12]/P0001 ,
		_w2318_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\u0_slt3_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2319_
	);
	LUT2 #(
		.INIT('h1)
	) name174 (
		_w2318_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h8)
	) name175 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[11]/P0001 ,
		_w2321_
	);
	LUT2 #(
		.INIT('h2)
	) name176 (
		\u0_slt3_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2322_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w2321_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[10]/P0001 ,
		_w2324_
	);
	LUT2 #(
		.INIT('h2)
	) name179 (
		\u0_slt3_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[9]/P0001 ,
		_w2327_
	);
	LUT2 #(
		.INIT('h2)
	) name182 (
		\u0_slt3_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w2327_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h8)
	) name184 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[8]/P0001 ,
		_w2330_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\u0_slt3_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2331_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w2330_,
		_w2331_,
		_w2332_
	);
	LUT2 #(
		.INIT('h8)
	) name187 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[7]/P0001 ,
		_w2333_
	);
	LUT2 #(
		.INIT('h2)
	) name188 (
		\u0_slt3_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2334_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w2333_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[6]/P0001 ,
		_w2336_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		\u0_slt3_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2337_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w2336_,
		_w2337_,
		_w2338_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[5]/P0001 ,
		_w2339_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		\u0_slt3_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2340_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w2339_,
		_w2340_,
		_w2341_
	);
	LUT2 #(
		.INIT('h8)
	) name196 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[4]/P0001 ,
		_w2342_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		\u0_slt3_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w2342_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h8)
	) name199 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[3]/P0001 ,
		_w2345_
	);
	LUT2 #(
		.INIT('h2)
	) name200 (
		\u0_slt3_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2346_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		_w2345_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[2]/P0001 ,
		_w2348_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\u0_slt3_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w2348_,
		_w2349_,
		_w2350_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[1]/P0001 ,
		_w2351_
	);
	LUT2 #(
		.INIT('h2)
	) name206 (
		\u0_slt3_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2352_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		_w2351_,
		_w2352_,
		_w2353_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\u2_ld_reg/P0001 ,
		\u3_dout_reg[0]/P0001 ,
		_w2354_
	);
	LUT2 #(
		.INIT('h2)
	) name209 (
		\u0_slt4_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2355_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		_w2354_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h8)
	) name211 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[19]/P0001 ,
		_w2357_
	);
	LUT2 #(
		.INIT('h2)
	) name212 (
		\u0_slt4_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2358_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w2357_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[18]/P0001 ,
		_w2360_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		\u0_slt4_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2361_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w2360_,
		_w2361_,
		_w2362_
	);
	LUT2 #(
		.INIT('h8)
	) name217 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[17]/P0001 ,
		_w2363_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		\u0_slt4_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2364_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w2363_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h8)
	) name220 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[16]/P0001 ,
		_w2366_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\u0_slt4_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2367_
	);
	LUT2 #(
		.INIT('h1)
	) name222 (
		_w2366_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h8)
	) name223 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[15]/P0001 ,
		_w2369_
	);
	LUT2 #(
		.INIT('h2)
	) name224 (
		\u0_slt4_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2370_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w2369_,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[14]/P0001 ,
		_w2372_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		\u0_slt4_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2373_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w2372_,
		_w2373_,
		_w2374_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[13]/P0001 ,
		_w2375_
	);
	LUT2 #(
		.INIT('h2)
	) name230 (
		\u0_slt4_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2376_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w2375_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h8)
	) name232 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[12]/P0001 ,
		_w2378_
	);
	LUT2 #(
		.INIT('h2)
	) name233 (
		\u0_slt4_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2379_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w2378_,
		_w2379_,
		_w2380_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[11]/P0001 ,
		_w2381_
	);
	LUT2 #(
		.INIT('h2)
	) name236 (
		\u0_slt4_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2382_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w2381_,
		_w2382_,
		_w2383_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[10]/P0001 ,
		_w2384_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		\u0_slt4_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2385_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w2384_,
		_w2385_,
		_w2386_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[9]/P0001 ,
		_w2387_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		\u0_slt4_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2388_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w2387_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h8)
	) name244 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[8]/P0001 ,
		_w2390_
	);
	LUT2 #(
		.INIT('h2)
	) name245 (
		\u0_slt4_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w2390_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[7]/P0001 ,
		_w2393_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		\u0_slt4_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		_w2393_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[6]/P0001 ,
		_w2396_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\u0_slt4_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2397_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w2396_,
		_w2397_,
		_w2398_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[5]/P0001 ,
		_w2399_
	);
	LUT2 #(
		.INIT('h2)
	) name254 (
		\u0_slt4_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2400_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		_w2399_,
		_w2400_,
		_w2401_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[4]/P0001 ,
		_w2402_
	);
	LUT2 #(
		.INIT('h2)
	) name257 (
		\u0_slt4_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2403_
	);
	LUT2 #(
		.INIT('h1)
	) name258 (
		_w2402_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h8)
	) name259 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[3]/P0001 ,
		_w2405_
	);
	LUT2 #(
		.INIT('h2)
	) name260 (
		\u0_slt4_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2406_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w2405_,
		_w2406_,
		_w2407_
	);
	LUT2 #(
		.INIT('h8)
	) name262 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[2]/P0001 ,
		_w2408_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\u0_slt4_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2409_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w2408_,
		_w2409_,
		_w2410_
	);
	LUT2 #(
		.INIT('h8)
	) name265 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[1]/P0001 ,
		_w2411_
	);
	LUT2 #(
		.INIT('h2)
	) name266 (
		\u0_slt4_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2412_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w2411_,
		_w2412_,
		_w2413_
	);
	LUT2 #(
		.INIT('h8)
	) name268 (
		\u2_ld_reg/P0001 ,
		\u4_dout_reg[0]/P0001 ,
		_w2414_
	);
	LUT2 #(
		.INIT('h2)
	) name269 (
		\u0_slt5_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2415_
	);
	LUT2 #(
		.INIT('h1)
	) name270 (
		_w2414_,
		_w2415_,
		_w2416_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		\u0_slt5_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2417_
	);
	LUT2 #(
		.INIT('h2)
	) name272 (
		\u0_slt5_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2418_
	);
	LUT2 #(
		.INIT('h2)
	) name273 (
		\u0_slt5_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2419_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		\u0_slt5_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2420_
	);
	LUT2 #(
		.INIT('h2)
	) name275 (
		\u0_slt5_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2421_
	);
	LUT2 #(
		.INIT('h2)
	) name276 (
		\u0_slt5_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2422_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\u0_slt5_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name278 (
		\u0_slt5_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2424_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		\u0_slt5_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2425_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\u0_slt5_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2426_
	);
	LUT2 #(
		.INIT('h2)
	) name281 (
		\u0_slt5_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2427_
	);
	LUT2 #(
		.INIT('h2)
	) name282 (
		\u0_slt5_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2428_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		\u0_slt5_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2429_
	);
	LUT2 #(
		.INIT('h2)
	) name284 (
		\u0_slt5_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2430_
	);
	LUT2 #(
		.INIT('h2)
	) name285 (
		\u0_slt5_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2431_
	);
	LUT2 #(
		.INIT('h2)
	) name286 (
		\u0_slt5_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2432_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\u0_slt5_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2433_
	);
	LUT2 #(
		.INIT('h2)
	) name288 (
		\u0_slt5_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2434_
	);
	LUT2 #(
		.INIT('h2)
	) name289 (
		\u0_slt5_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2435_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		\u0_slt6_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2436_
	);
	LUT2 #(
		.INIT('h8)
	) name291 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[19]/P0001 ,
		_w2437_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		\u0_slt6_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2438_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w2437_,
		_w2438_,
		_w2439_
	);
	LUT2 #(
		.INIT('h8)
	) name294 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[18]/P0001 ,
		_w2440_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		\u0_slt6_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2441_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w2440_,
		_w2441_,
		_w2442_
	);
	LUT2 #(
		.INIT('h8)
	) name297 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[17]/P0001 ,
		_w2443_
	);
	LUT2 #(
		.INIT('h2)
	) name298 (
		\u0_slt6_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w2443_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h8)
	) name300 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[16]/P0001 ,
		_w2446_
	);
	LUT2 #(
		.INIT('h2)
	) name301 (
		\u0_slt6_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2447_
	);
	LUT2 #(
		.INIT('h1)
	) name302 (
		_w2446_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('h8)
	) name303 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[15]/P0001 ,
		_w2449_
	);
	LUT2 #(
		.INIT('h2)
	) name304 (
		\u0_slt6_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w2449_,
		_w2450_,
		_w2451_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[14]/P0001 ,
		_w2452_
	);
	LUT2 #(
		.INIT('h2)
	) name307 (
		\u0_slt6_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2453_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w2452_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[13]/P0001 ,
		_w2455_
	);
	LUT2 #(
		.INIT('h2)
	) name310 (
		\u0_slt6_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2456_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w2455_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h8)
	) name312 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[12]/P0001 ,
		_w2458_
	);
	LUT2 #(
		.INIT('h2)
	) name313 (
		\u0_slt6_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2459_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w2458_,
		_w2459_,
		_w2460_
	);
	LUT2 #(
		.INIT('h8)
	) name315 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[11]/P0001 ,
		_w2461_
	);
	LUT2 #(
		.INIT('h2)
	) name316 (
		\u0_slt6_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2462_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w2461_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[10]/P0001 ,
		_w2464_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		\u0_slt6_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2465_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w2464_,
		_w2465_,
		_w2466_
	);
	LUT2 #(
		.INIT('h8)
	) name321 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[9]/P0001 ,
		_w2467_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		\u0_slt6_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2468_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w2467_,
		_w2468_,
		_w2469_
	);
	LUT2 #(
		.INIT('h8)
	) name324 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[8]/P0001 ,
		_w2470_
	);
	LUT2 #(
		.INIT('h2)
	) name325 (
		\u0_slt6_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2471_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w2470_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h8)
	) name327 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[7]/P0001 ,
		_w2473_
	);
	LUT2 #(
		.INIT('h2)
	) name328 (
		\u0_slt6_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2474_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		_w2473_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[6]/P0001 ,
		_w2476_
	);
	LUT2 #(
		.INIT('h2)
	) name331 (
		\u0_slt6_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2477_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w2476_,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[5]/P0001 ,
		_w2479_
	);
	LUT2 #(
		.INIT('h2)
	) name334 (
		\u0_slt6_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2480_
	);
	LUT2 #(
		.INIT('h1)
	) name335 (
		_w2479_,
		_w2480_,
		_w2481_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[4]/P0001 ,
		_w2482_
	);
	LUT2 #(
		.INIT('h2)
	) name337 (
		\u0_slt6_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2483_
	);
	LUT2 #(
		.INIT('h1)
	) name338 (
		_w2482_,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h8)
	) name339 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[3]/P0001 ,
		_w2485_
	);
	LUT2 #(
		.INIT('h2)
	) name340 (
		\u0_slt6_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2486_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT2 #(
		.INIT('h8)
	) name342 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[2]/P0001 ,
		_w2488_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		\u0_slt6_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2489_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w2488_,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h8)
	) name345 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[1]/P0001 ,
		_w2491_
	);
	LUT2 #(
		.INIT('h2)
	) name346 (
		\u0_slt6_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2492_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w2491_,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h8)
	) name348 (
		\u2_ld_reg/P0001 ,
		\u5_dout_reg[0]/P0001 ,
		_w2494_
	);
	LUT2 #(
		.INIT('h2)
	) name349 (
		\u0_slt7_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2495_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w2494_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h8)
	) name351 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[19]/P0001 ,
		_w2497_
	);
	LUT2 #(
		.INIT('h2)
	) name352 (
		\u0_slt7_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2498_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		_w2497_,
		_w2498_,
		_w2499_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[18]/P0001 ,
		_w2500_
	);
	LUT2 #(
		.INIT('h2)
	) name355 (
		\u0_slt7_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2501_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w2500_,
		_w2501_,
		_w2502_
	);
	LUT2 #(
		.INIT('h8)
	) name357 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[17]/P0001 ,
		_w2503_
	);
	LUT2 #(
		.INIT('h2)
	) name358 (
		\u0_slt7_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2504_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w2503_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[16]/P0001 ,
		_w2506_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		\u0_slt7_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w2506_,
		_w2507_,
		_w2508_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[15]/P0001 ,
		_w2509_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		\u0_slt7_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2510_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w2509_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h8)
	) name366 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[14]/P0001 ,
		_w2512_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\u0_slt7_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2513_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w2512_,
		_w2513_,
		_w2514_
	);
	LUT2 #(
		.INIT('h8)
	) name369 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[13]/P0001 ,
		_w2515_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\u0_slt7_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2516_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w2515_,
		_w2516_,
		_w2517_
	);
	LUT2 #(
		.INIT('h8)
	) name372 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[12]/P0001 ,
		_w2518_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\u0_slt7_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2519_
	);
	LUT2 #(
		.INIT('h1)
	) name374 (
		_w2518_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h8)
	) name375 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[11]/P0001 ,
		_w2521_
	);
	LUT2 #(
		.INIT('h2)
	) name376 (
		\u0_slt7_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2522_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		_w2521_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[10]/P0001 ,
		_w2524_
	);
	LUT2 #(
		.INIT('h2)
	) name379 (
		\u0_slt7_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2525_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w2524_,
		_w2525_,
		_w2526_
	);
	LUT2 #(
		.INIT('h8)
	) name381 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[9]/P0001 ,
		_w2527_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\u0_slt7_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2528_
	);
	LUT2 #(
		.INIT('h1)
	) name383 (
		_w2527_,
		_w2528_,
		_w2529_
	);
	LUT2 #(
		.INIT('h8)
	) name384 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[8]/P0001 ,
		_w2530_
	);
	LUT2 #(
		.INIT('h2)
	) name385 (
		\u0_slt7_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2531_
	);
	LUT2 #(
		.INIT('h1)
	) name386 (
		_w2530_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h8)
	) name387 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[7]/P0001 ,
		_w2533_
	);
	LUT2 #(
		.INIT('h2)
	) name388 (
		\u0_slt7_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2534_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w2533_,
		_w2534_,
		_w2535_
	);
	LUT2 #(
		.INIT('h8)
	) name390 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[6]/P0001 ,
		_w2536_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		\u0_slt7_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w2536_,
		_w2537_,
		_w2538_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[5]/P0001 ,
		_w2539_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		\u0_slt7_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2540_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w2539_,
		_w2540_,
		_w2541_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[4]/P0001 ,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name397 (
		\u0_slt7_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2543_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w2542_,
		_w2543_,
		_w2544_
	);
	LUT2 #(
		.INIT('h8)
	) name399 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[3]/P0001 ,
		_w2545_
	);
	LUT2 #(
		.INIT('h2)
	) name400 (
		\u0_slt7_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2546_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		_w2545_,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[2]/P0001 ,
		_w2548_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		\u0_slt7_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2549_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w2548_,
		_w2549_,
		_w2550_
	);
	LUT2 #(
		.INIT('h8)
	) name405 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[1]/P0001 ,
		_w2551_
	);
	LUT2 #(
		.INIT('h2)
	) name406 (
		\u0_slt7_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2552_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w2551_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h8)
	) name408 (
		\u2_ld_reg/P0001 ,
		\u6_dout_reg[0]/P0001 ,
		_w2554_
	);
	LUT2 #(
		.INIT('h2)
	) name409 (
		\u0_slt8_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2555_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w2554_,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[19]/P0001 ,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		\u0_slt8_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2558_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w2557_,
		_w2558_,
		_w2559_
	);
	LUT2 #(
		.INIT('h8)
	) name414 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[18]/P0001 ,
		_w2560_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		\u0_slt8_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2561_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w2560_,
		_w2561_,
		_w2562_
	);
	LUT2 #(
		.INIT('h8)
	) name417 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[17]/P0001 ,
		_w2563_
	);
	LUT2 #(
		.INIT('h2)
	) name418 (
		\u0_slt8_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2564_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w2563_,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('h8)
	) name420 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[16]/P0001 ,
		_w2566_
	);
	LUT2 #(
		.INIT('h2)
	) name421 (
		\u0_slt8_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name422 (
		_w2566_,
		_w2567_,
		_w2568_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[15]/P0001 ,
		_w2569_
	);
	LUT2 #(
		.INIT('h2)
	) name424 (
		\u0_slt8_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2570_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		_w2569_,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[14]/P0001 ,
		_w2572_
	);
	LUT2 #(
		.INIT('h2)
	) name427 (
		\u0_slt8_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2573_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w2572_,
		_w2573_,
		_w2574_
	);
	LUT2 #(
		.INIT('h8)
	) name429 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[13]/P0001 ,
		_w2575_
	);
	LUT2 #(
		.INIT('h2)
	) name430 (
		\u0_slt8_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2576_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w2575_,
		_w2576_,
		_w2577_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[12]/P0001 ,
		_w2578_
	);
	LUT2 #(
		.INIT('h2)
	) name433 (
		\u0_slt8_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2579_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w2578_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[11]/P0001 ,
		_w2581_
	);
	LUT2 #(
		.INIT('h2)
	) name436 (
		\u0_slt8_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2582_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w2581_,
		_w2582_,
		_w2583_
	);
	LUT2 #(
		.INIT('h8)
	) name438 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[10]/P0001 ,
		_w2584_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		\u0_slt8_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2585_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		_w2584_,
		_w2585_,
		_w2586_
	);
	LUT2 #(
		.INIT('h8)
	) name441 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[9]/P0001 ,
		_w2587_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		\u0_slt8_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2588_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		_w2587_,
		_w2588_,
		_w2589_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[8]/P0001 ,
		_w2590_
	);
	LUT2 #(
		.INIT('h2)
	) name445 (
		\u0_slt8_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2591_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		_w2590_,
		_w2591_,
		_w2592_
	);
	LUT2 #(
		.INIT('h8)
	) name447 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[7]/P0001 ,
		_w2593_
	);
	LUT2 #(
		.INIT('h2)
	) name448 (
		\u0_slt8_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w2593_,
		_w2594_,
		_w2595_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[6]/P0001 ,
		_w2596_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		\u0_slt8_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2597_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w2596_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h8)
	) name453 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[5]/P0001 ,
		_w2599_
	);
	LUT2 #(
		.INIT('h2)
	) name454 (
		\u0_slt8_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2600_
	);
	LUT2 #(
		.INIT('h1)
	) name455 (
		_w2599_,
		_w2600_,
		_w2601_
	);
	LUT2 #(
		.INIT('h8)
	) name456 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[4]/P0001 ,
		_w2602_
	);
	LUT2 #(
		.INIT('h2)
	) name457 (
		\u0_slt8_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2603_
	);
	LUT2 #(
		.INIT('h1)
	) name458 (
		_w2602_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h8)
	) name459 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[3]/P0001 ,
		_w2605_
	);
	LUT2 #(
		.INIT('h2)
	) name460 (
		\u0_slt8_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2606_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w2605_,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h8)
	) name462 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[2]/P0001 ,
		_w2608_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		\u0_slt8_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2609_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w2608_,
		_w2609_,
		_w2610_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[1]/P0001 ,
		_w2611_
	);
	LUT2 #(
		.INIT('h2)
	) name466 (
		\u0_slt8_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2612_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w2611_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		\u2_ld_reg/P0001 ,
		\u7_dout_reg[0]/P0001 ,
		_w2614_
	);
	LUT2 #(
		.INIT('h2)
	) name469 (
		\u0_slt9_r_reg[19]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2615_
	);
	LUT2 #(
		.INIT('h1)
	) name470 (
		_w2614_,
		_w2615_,
		_w2616_
	);
	LUT2 #(
		.INIT('h8)
	) name471 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[19]/P0001 ,
		_w2617_
	);
	LUT2 #(
		.INIT('h2)
	) name472 (
		\u0_slt9_r_reg[18]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2618_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		_w2617_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[18]/P0001 ,
		_w2620_
	);
	LUT2 #(
		.INIT('h2)
	) name475 (
		\u0_slt9_r_reg[17]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2621_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h8)
	) name477 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[17]/P0001 ,
		_w2623_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		\u0_slt9_r_reg[16]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2624_
	);
	LUT2 #(
		.INIT('h1)
	) name479 (
		_w2623_,
		_w2624_,
		_w2625_
	);
	LUT2 #(
		.INIT('h8)
	) name480 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[16]/P0001 ,
		_w2626_
	);
	LUT2 #(
		.INIT('h2)
	) name481 (
		\u0_slt9_r_reg[15]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2627_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w2626_,
		_w2627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[15]/P0001 ,
		_w2629_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\u0_slt9_r_reg[14]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2630_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w2629_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h8)
	) name486 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[14]/P0001 ,
		_w2632_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		\u0_slt9_r_reg[13]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w2632_,
		_w2633_,
		_w2634_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[13]/P0001 ,
		_w2635_
	);
	LUT2 #(
		.INIT('h2)
	) name490 (
		\u0_slt9_r_reg[12]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2636_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w2635_,
		_w2636_,
		_w2637_
	);
	LUT2 #(
		.INIT('h8)
	) name492 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[12]/P0001 ,
		_w2638_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		\u0_slt9_r_reg[11]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2639_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		_w2638_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h8)
	) name495 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[11]/P0001 ,
		_w2641_
	);
	LUT2 #(
		.INIT('h2)
	) name496 (
		\u0_slt9_r_reg[10]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2642_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		_w2641_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[10]/P0001 ,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name499 (
		\u0_slt9_r_reg[9]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w2644_,
		_w2645_,
		_w2646_
	);
	LUT2 #(
		.INIT('h8)
	) name501 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[9]/P0001 ,
		_w2647_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		\u0_slt9_r_reg[8]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2648_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		_w2647_,
		_w2648_,
		_w2649_
	);
	LUT2 #(
		.INIT('h8)
	) name504 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[8]/P0001 ,
		_w2650_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		\u0_slt9_r_reg[7]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2651_
	);
	LUT2 #(
		.INIT('h1)
	) name506 (
		_w2650_,
		_w2651_,
		_w2652_
	);
	LUT2 #(
		.INIT('h8)
	) name507 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[7]/P0001 ,
		_w2653_
	);
	LUT2 #(
		.INIT('h2)
	) name508 (
		\u0_slt9_r_reg[6]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w2653_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h8)
	) name510 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[6]/P0001 ,
		_w2656_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		\u0_slt9_r_reg[5]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2657_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w2656_,
		_w2657_,
		_w2658_
	);
	LUT2 #(
		.INIT('h4)
	) name513 (
		\dma_ack_i[0]_pad ,
		\dma_req_o[0]_pad ,
		_w2659_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		\u13_occ0_r_reg[5]/NET0131 ,
		\u3_status_reg[1]/P0001 ,
		_w2660_
	);
	LUT2 #(
		.INIT('h8)
	) name515 (
		\u13_occ0_r_reg[5]/NET0131 ,
		\u3_status_reg[1]/P0001 ,
		_w2661_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		\u13_occ0_r_reg[4]/NET0131 ,
		\u3_status_reg[0]/P0001 ,
		_w2662_
	);
	LUT2 #(
		.INIT('h4)
	) name517 (
		_w2661_,
		_w2662_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		\u3_empty_reg/NET0131 ,
		_w2660_,
		_w2664_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		_w2663_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h2)
	) name520 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h4)
	) name521 (
		\dma_ack_i[0]_pad ,
		\u13_occ0_r_reg[6]/NET0131 ,
		_w2667_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		_w2666_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h8)
	) name523 (
		\u16_u0_dma_req_r1_reg/P0001 ,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w2659_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h4)
	) name525 (
		\dma_ack_i[1]_pad ,
		\dma_req_o[1]_pad ,
		_w2671_
	);
	LUT2 #(
		.INIT('h1)
	) name526 (
		\u13_occ0_r_reg[13]/NET0131 ,
		\u4_status_reg[1]/P0001 ,
		_w2672_
	);
	LUT2 #(
		.INIT('h8)
	) name527 (
		\u13_occ0_r_reg[13]/NET0131 ,
		\u4_status_reg[1]/P0001 ,
		_w2673_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		\u13_occ0_r_reg[12]/NET0131 ,
		\u4_status_reg[0]/P0001 ,
		_w2674_
	);
	LUT2 #(
		.INIT('h4)
	) name529 (
		_w2673_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h1)
	) name530 (
		\u4_empty_reg/NET0131 ,
		_w2672_,
		_w2676_
	);
	LUT2 #(
		.INIT('h4)
	) name531 (
		_w2675_,
		_w2676_,
		_w2677_
	);
	LUT2 #(
		.INIT('h2)
	) name532 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2677_,
		_w2678_
	);
	LUT2 #(
		.INIT('h4)
	) name533 (
		\dma_ack_i[1]_pad ,
		\u13_occ0_r_reg[14]/NET0131 ,
		_w2679_
	);
	LUT2 #(
		.INIT('h8)
	) name534 (
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT2 #(
		.INIT('h8)
	) name535 (
		\u16_u1_dma_req_r1_reg/P0001 ,
		_w2680_,
		_w2681_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w2671_,
		_w2681_,
		_w2682_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		\dma_ack_i[2]_pad ,
		\dma_req_o[2]_pad ,
		_w2683_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		\u13_occ0_r_reg[21]/NET0131 ,
		\u5_status_reg[1]/P0001 ,
		_w2684_
	);
	LUT2 #(
		.INIT('h8)
	) name539 (
		\u13_occ0_r_reg[21]/NET0131 ,
		\u5_status_reg[1]/P0001 ,
		_w2685_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		\u13_occ0_r_reg[20]/NET0131 ,
		\u5_status_reg[0]/P0001 ,
		_w2686_
	);
	LUT2 #(
		.INIT('h4)
	) name541 (
		_w2685_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h1)
	) name542 (
		\u5_empty_reg/NET0131 ,
		_w2684_,
		_w2688_
	);
	LUT2 #(
		.INIT('h4)
	) name543 (
		_w2687_,
		_w2688_,
		_w2689_
	);
	LUT2 #(
		.INIT('h2)
	) name544 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2689_,
		_w2690_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\dma_ack_i[2]_pad ,
		\u13_occ0_r_reg[22]/NET0131 ,
		_w2691_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		_w2690_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h8)
	) name547 (
		\u16_u2_dma_req_r1_reg/P0001 ,
		_w2692_,
		_w2693_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w2683_,
		_w2693_,
		_w2694_
	);
	LUT2 #(
		.INIT('h4)
	) name549 (
		\dma_ack_i[3]_pad ,
		\dma_req_o[3]_pad ,
		_w2695_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		\u13_occ0_r_reg[29]/NET0131 ,
		\u6_status_reg[1]/P0001 ,
		_w2696_
	);
	LUT2 #(
		.INIT('h8)
	) name551 (
		\u13_occ0_r_reg[29]/NET0131 ,
		\u6_status_reg[1]/P0001 ,
		_w2697_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		\u13_occ0_r_reg[28]/NET0131 ,
		\u6_status_reg[0]/P0001 ,
		_w2698_
	);
	LUT2 #(
		.INIT('h4)
	) name553 (
		_w2697_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h1)
	) name554 (
		\u6_empty_reg/NET0131 ,
		_w2696_,
		_w2700_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		\dma_ack_i[3]_pad ,
		\u13_occ0_r_reg[30]/NET0131 ,
		_w2703_
	);
	LUT2 #(
		.INIT('h8)
	) name558 (
		_w2702_,
		_w2703_,
		_w2704_
	);
	LUT2 #(
		.INIT('h8)
	) name559 (
		\u16_u3_dma_req_r1_reg/P0001 ,
		_w2704_,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w2695_,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('h4)
	) name561 (
		\dma_ack_i[4]_pad ,
		\dma_req_o[4]_pad ,
		_w2707_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		\u13_occ1_r_reg[5]/NET0131 ,
		\u7_status_reg[1]/P0001 ,
		_w2708_
	);
	LUT2 #(
		.INIT('h8)
	) name563 (
		\u13_occ1_r_reg[5]/NET0131 ,
		\u7_status_reg[1]/P0001 ,
		_w2709_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		\u13_occ1_r_reg[4]/NET0131 ,
		\u7_status_reg[0]/P0001 ,
		_w2710_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w2709_,
		_w2710_,
		_w2711_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		\u7_empty_reg/NET0131 ,
		_w2708_,
		_w2712_
	);
	LUT2 #(
		.INIT('h4)
	) name567 (
		_w2711_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h2)
	) name568 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2713_,
		_w2714_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		\dma_ack_i[4]_pad ,
		\u13_occ1_r_reg[6]/NET0131 ,
		_w2715_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		_w2714_,
		_w2715_,
		_w2716_
	);
	LUT2 #(
		.INIT('h8)
	) name571 (
		\u16_u4_dma_req_r1_reg/P0001 ,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w2707_,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h4)
	) name573 (
		\dma_ack_i[5]_pad ,
		\dma_req_o[5]_pad ,
		_w2719_
	);
	LUT2 #(
		.INIT('h1)
	) name574 (
		\u13_occ1_r_reg[13]/NET0131 ,
		\u8_status_reg[1]/P0001 ,
		_w2720_
	);
	LUT2 #(
		.INIT('h8)
	) name575 (
		\u13_occ1_r_reg[13]/NET0131 ,
		\u8_status_reg[1]/P0001 ,
		_w2721_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		\u13_occ1_r_reg[12]/NET0131 ,
		\u8_status_reg[0]/P0001 ,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		_w2721_,
		_w2722_,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		\u8_empty_reg/NET0131 ,
		_w2720_,
		_w2724_
	);
	LUT2 #(
		.INIT('h4)
	) name579 (
		_w2723_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h4)
	) name581 (
		\dma_ack_i[5]_pad ,
		\u13_occ1_r_reg[14]/NET0131 ,
		_w2727_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		_w2726_,
		_w2727_,
		_w2728_
	);
	LUT2 #(
		.INIT('h8)
	) name583 (
		\u16_u5_dma_req_r1_reg/P0001 ,
		_w2728_,
		_w2729_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w2719_,
		_w2729_,
		_w2730_
	);
	LUT2 #(
		.INIT('h8)
	) name585 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[5]/P0001 ,
		_w2731_
	);
	LUT2 #(
		.INIT('h2)
	) name586 (
		\u0_slt9_r_reg[4]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2732_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		_w2731_,
		_w2732_,
		_w2733_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		\u13_ints_r_reg[11]/NET0131 ,
		\u20_int_set_reg[0]/NET0131 ,
		_w2734_
	);
	LUT2 #(
		.INIT('h8)
	) name589 (
		wb_cyc_i_pad,
		wb_stb_i_pad,
		_w2735_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		\u12_re2_reg/NET0131 ,
		wb_we_i_pad,
		_w2736_
	);
	LUT2 #(
		.INIT('h8)
	) name591 (
		_w2735_,
		_w2736_,
		_w2737_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		\u12_re1_reg/P0001 ,
		_w2737_,
		_w2738_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w2739_
	);
	LUT2 #(
		.INIT('h4)
	) name594 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w2740_
	);
	LUT2 #(
		.INIT('h8)
	) name595 (
		\wb_addr_i[4]_pad ,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		_w2739_,
		_w2741_,
		_w2742_
	);
	LUT2 #(
		.INIT('h8)
	) name597 (
		_w2738_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name598 (
		_w2734_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h1)
	) name599 (
		\u13_ints_r_reg[14]/NET0131 ,
		\u21_int_set_reg[0]/NET0131 ,
		_w2745_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w2743_,
		_w2745_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		\u13_ints_r_reg[17]/NET0131 ,
		\u22_int_set_reg[0]/NET0131 ,
		_w2747_
	);
	LUT2 #(
		.INIT('h1)
	) name602 (
		_w2743_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		\u13_ints_r_reg[2]/NET0131 ,
		\u17_int_set_reg[0]/NET0131 ,
		_w2749_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w2743_,
		_w2749_,
		_w2750_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		\u13_ints_r_reg[5]/NET0131 ,
		\u18_int_set_reg[0]/NET0131 ,
		_w2751_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		_w2743_,
		_w2751_,
		_w2752_
	);
	LUT2 #(
		.INIT('h1)
	) name607 (
		\u13_ints_r_reg[8]/NET0131 ,
		\u19_int_set_reg[0]/NET0131 ,
		_w2753_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w2743_,
		_w2753_,
		_w2754_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[4]/P0001 ,
		_w2755_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		\u0_slt9_r_reg[3]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2756_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w2755_,
		_w2756_,
		_w2757_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		\u14_u1_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2758_
	);
	LUT2 #(
		.INIT('h4)
	) name613 (
		\u14_u1_en_out_l2_reg/P0001 ,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h1)
	) name614 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\u13_occ0_r_reg[11]/NET0131 ,
		_w2760_
	);
	LUT2 #(
		.INIT('h4)
	) name615 (
		\u4_rp_reg[0]/P0001 ,
		_w2760_,
		_w2761_
	);
	LUT2 #(
		.INIT('h2)
	) name616 (
		_w2759_,
		_w2761_,
		_w2762_
	);
	LUT2 #(
		.INIT('h8)
	) name617 (
		\u4_rp_reg[1]/NET0131 ,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h1)
	) name618 (
		\u4_rp_reg[2]/NET0131 ,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h8)
	) name619 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2765_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w2762_,
		_w2765_,
		_w2766_
	);
	LUT2 #(
		.INIT('h2)
	) name621 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		_w2764_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h8)
	) name623 (
		\u14_u2_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2769_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		\u14_u2_en_out_l2_reg/P0001 ,
		_w2769_,
		_w2770_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		\u13_occ0_r_reg[18]/NET0131 ,
		\u13_occ0_r_reg[19]/NET0131 ,
		_w2771_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		\u5_rp_reg[0]/P0001 ,
		_w2771_,
		_w2772_
	);
	LUT2 #(
		.INIT('h2)
	) name627 (
		_w2770_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h8)
	) name628 (
		\u5_rp_reg[1]/NET0131 ,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		\u5_rp_reg[2]/NET0131 ,
		_w2774_,
		_w2775_
	);
	LUT2 #(
		.INIT('h8)
	) name630 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2776_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		_w2773_,
		_w2776_,
		_w2777_
	);
	LUT2 #(
		.INIT('h2)
	) name632 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h4)
	) name633 (
		_w2775_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		\u8_rp_reg[1]/NET0131 ,
		_w2162_,
		_w2780_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		\u8_rp_reg[2]/NET0131 ,
		_w2780_,
		_w2781_
	);
	LUT2 #(
		.INIT('h2)
	) name636 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2164_,
		_w2782_
	);
	LUT2 #(
		.INIT('h4)
	) name637 (
		_w2781_,
		_w2782_,
		_w2783_
	);
	LUT2 #(
		.INIT('h1)
	) name638 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		_w2784_
	);
	LUT2 #(
		.INIT('h4)
	) name639 (
		\u3_rp_reg[0]/P0001 ,
		_w2784_,
		_w2785_
	);
	LUT2 #(
		.INIT('h4)
	) name640 (
		\u14_u0_en_out_l2_reg/P0001 ,
		\u14_u0_en_out_l_reg/NET0131 ,
		_w2786_
	);
	LUT2 #(
		.INIT('h8)
	) name641 (
		\valid_s_reg/NET0131 ,
		_w2786_,
		_w2787_
	);
	LUT2 #(
		.INIT('h4)
	) name642 (
		_w2785_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		\u3_rp_reg[1]/NET0131 ,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		\u3_rp_reg[2]/NET0131 ,
		_w2789_,
		_w2790_
	);
	LUT2 #(
		.INIT('h8)
	) name645 (
		\u3_rp_reg[2]/NET0131 ,
		_w2789_,
		_w2791_
	);
	LUT2 #(
		.INIT('h2)
	) name646 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w2790_,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name647 (
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h8)
	) name648 (
		\u14_u3_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2794_
	);
	LUT2 #(
		.INIT('h4)
	) name649 (
		\u14_u3_en_out_l2_reg/P0001 ,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h1)
	) name650 (
		\u13_occ0_r_reg[26]/NET0131 ,
		\u13_occ0_r_reg[27]/NET0131 ,
		_w2796_
	);
	LUT2 #(
		.INIT('h4)
	) name651 (
		\u6_rp_reg[0]/P0001 ,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		_w2795_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h8)
	) name653 (
		\u6_rp_reg[1]/NET0131 ,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		\u6_rp_reg[2]/NET0131 ,
		_w2799_,
		_w2800_
	);
	LUT2 #(
		.INIT('h8)
	) name655 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2801_
	);
	LUT2 #(
		.INIT('h8)
	) name656 (
		_w2798_,
		_w2801_,
		_w2802_
	);
	LUT2 #(
		.INIT('h2)
	) name657 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w2800_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		_w2805_
	);
	LUT2 #(
		.INIT('h4)
	) name660 (
		\u7_rp_reg[0]/P0001 ,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h8)
	) name661 (
		\u14_u4_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w2807_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		\u14_u4_en_out_l2_reg/P0001 ,
		_w2807_,
		_w2808_
	);
	LUT2 #(
		.INIT('h4)
	) name663 (
		_w2806_,
		_w2808_,
		_w2809_
	);
	LUT2 #(
		.INIT('h8)
	) name664 (
		\u7_rp_reg[1]/NET0131 ,
		_w2809_,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		\u7_rp_reg[2]/NET0131 ,
		_w2810_,
		_w2811_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		\u7_rp_reg[2]/NET0131 ,
		_w2810_,
		_w2812_
	);
	LUT2 #(
		.INIT('h2)
	) name667 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2811_,
		_w2813_
	);
	LUT2 #(
		.INIT('h4)
	) name668 (
		_w2812_,
		_w2813_,
		_w2814_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		\u3_rp_reg[3]/NET0131 ,
		_w2791_,
		_w2815_
	);
	LUT2 #(
		.INIT('h8)
	) name670 (
		\u3_rp_reg[3]/NET0131 ,
		_w2791_,
		_w2816_
	);
	LUT2 #(
		.INIT('h2)
	) name671 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w2815_,
		_w2817_
	);
	LUT2 #(
		.INIT('h4)
	) name672 (
		_w2816_,
		_w2817_,
		_w2818_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		\u4_rp_reg[3]/NET0131 ,
		_w2766_,
		_w2819_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		\u4_rp_reg[3]/NET0131 ,
		_w2766_,
		_w2820_
	);
	LUT2 #(
		.INIT('h2)
	) name675 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2819_,
		_w2821_
	);
	LUT2 #(
		.INIT('h4)
	) name676 (
		_w2820_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		\u13_ints_r_reg[20]/NET0131 ,
		\u23_int_set_reg[0]/NET0131 ,
		_w2823_
	);
	LUT2 #(
		.INIT('h1)
	) name678 (
		_w2743_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		\u13_ints_r_reg[23]/NET0131 ,
		\u24_int_set_reg[0]/NET0131 ,
		_w2825_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		_w2743_,
		_w2825_,
		_w2826_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		\u13_ints_r_reg[26]/NET0131 ,
		\u25_int_set_reg[0]/NET0131 ,
		_w2827_
	);
	LUT2 #(
		.INIT('h1)
	) name682 (
		_w2743_,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		\u5_rp_reg[3]/NET0131 ,
		_w2777_,
		_w2829_
	);
	LUT2 #(
		.INIT('h8)
	) name684 (
		\u5_rp_reg[3]/NET0131 ,
		_w2777_,
		_w2830_
	);
	LUT2 #(
		.INIT('h2)
	) name685 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2829_,
		_w2831_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		_w2830_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h1)
	) name687 (
		\u6_rp_reg[3]/NET0131 ,
		_w2802_,
		_w2833_
	);
	LUT2 #(
		.INIT('h8)
	) name688 (
		\u6_rp_reg[3]/NET0131 ,
		_w2802_,
		_w2834_
	);
	LUT2 #(
		.INIT('h2)
	) name689 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2833_,
		_w2835_
	);
	LUT2 #(
		.INIT('h4)
	) name690 (
		_w2834_,
		_w2835_,
		_w2836_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		\u7_rp_reg[3]/NET0131 ,
		_w2812_,
		_w2837_
	);
	LUT2 #(
		.INIT('h8)
	) name692 (
		\u7_rp_reg[3]/NET0131 ,
		_w2812_,
		_w2838_
	);
	LUT2 #(
		.INIT('h2)
	) name693 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2837_,
		_w2839_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		_w2838_,
		_w2839_,
		_w2840_
	);
	LUT2 #(
		.INIT('h1)
	) name695 (
		\u8_rp_reg[1]/NET0131 ,
		_w2162_,
		_w2841_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2780_,
		_w2842_
	);
	LUT2 #(
		.INIT('h4)
	) name697 (
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h1)
	) name698 (
		\u3_rp_reg[1]/NET0131 ,
		_w2788_,
		_w2844_
	);
	LUT2 #(
		.INIT('h2)
	) name699 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w2789_,
		_w2845_
	);
	LUT2 #(
		.INIT('h4)
	) name700 (
		_w2844_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		\u4_rp_reg[1]/NET0131 ,
		_w2762_,
		_w2847_
	);
	LUT2 #(
		.INIT('h2)
	) name702 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2763_,
		_w2848_
	);
	LUT2 #(
		.INIT('h4)
	) name703 (
		_w2847_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		\u5_rp_reg[1]/NET0131 ,
		_w2773_,
		_w2850_
	);
	LUT2 #(
		.INIT('h2)
	) name705 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2774_,
		_w2851_
	);
	LUT2 #(
		.INIT('h4)
	) name706 (
		_w2850_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		\u6_rp_reg[1]/NET0131 ,
		_w2798_,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name708 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2799_,
		_w2854_
	);
	LUT2 #(
		.INIT('h4)
	) name709 (
		_w2853_,
		_w2854_,
		_w2855_
	);
	LUT2 #(
		.INIT('h1)
	) name710 (
		\u7_rp_reg[1]/NET0131 ,
		_w2809_,
		_w2856_
	);
	LUT2 #(
		.INIT('h2)
	) name711 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2810_,
		_w2857_
	);
	LUT2 #(
		.INIT('h4)
	) name712 (
		_w2856_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h8)
	) name713 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[3]/P0001 ,
		_w2859_
	);
	LUT2 #(
		.INIT('h2)
	) name714 (
		\u0_slt9_r_reg[2]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w2860_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w2859_,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h8)
	) name716 (
		suspended_o_pad,
		\u13_resume_req_reg/P0001 ,
		_w2862_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		\u2_sync_resume_reg/NET0131 ,
		_w2862_,
		_w2863_
	);
	LUT2 #(
		.INIT('h2)
	) name718 (
		\u2_res_cnt_reg[0]/P0001 ,
		\u2_res_cnt_reg[1]/P0001 ,
		_w2864_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		\u2_res_cnt_reg[2]/P0001 ,
		\u2_res_cnt_reg[3]/P0001 ,
		_w2865_
	);
	LUT2 #(
		.INIT('h8)
	) name720 (
		_w2864_,
		_w2865_,
		_w2866_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		_w2863_,
		_w2866_,
		_w2867_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		_w2159_,
		_w2160_,
		_w2868_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		\u8_rp_reg[0]/P0001 ,
		_w2868_,
		_w2869_
	);
	LUT2 #(
		.INIT('h8)
	) name724 (
		\u8_rp_reg[0]/P0001 ,
		_w2868_,
		_w2870_
	);
	LUT2 #(
		.INIT('h2)
	) name725 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2869_,
		_w2871_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		_w2870_,
		_w2871_,
		_w2872_
	);
	LUT2 #(
		.INIT('h8)
	) name727 (
		_w2784_,
		_w2787_,
		_w2873_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		\u3_rp_reg[0]/P0001 ,
		_w2873_,
		_w2874_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		\u3_rp_reg[0]/P0001 ,
		_w2873_,
		_w2875_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w2874_,
		_w2876_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w2875_,
		_w2876_,
		_w2877_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		_w2759_,
		_w2760_,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name733 (
		\u4_rp_reg[0]/P0001 ,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('h8)
	) name734 (
		\u4_rp_reg[0]/P0001 ,
		_w2878_,
		_w2880_
	);
	LUT2 #(
		.INIT('h2)
	) name735 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2879_,
		_w2881_
	);
	LUT2 #(
		.INIT('h4)
	) name736 (
		_w2880_,
		_w2881_,
		_w2882_
	);
	LUT2 #(
		.INIT('h8)
	) name737 (
		_w2770_,
		_w2771_,
		_w2883_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		\u5_rp_reg[0]/P0001 ,
		_w2883_,
		_w2884_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		\u5_rp_reg[0]/P0001 ,
		_w2883_,
		_w2885_
	);
	LUT2 #(
		.INIT('h2)
	) name740 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2884_,
		_w2886_
	);
	LUT2 #(
		.INIT('h4)
	) name741 (
		_w2885_,
		_w2886_,
		_w2887_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		_w2795_,
		_w2796_,
		_w2888_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		\u6_rp_reg[0]/P0001 ,
		_w2888_,
		_w2889_
	);
	LUT2 #(
		.INIT('h8)
	) name744 (
		\u6_rp_reg[0]/P0001 ,
		_w2888_,
		_w2890_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2889_,
		_w2891_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		_w2890_,
		_w2891_,
		_w2892_
	);
	LUT2 #(
		.INIT('h8)
	) name747 (
		_w2805_,
		_w2808_,
		_w2893_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		\u7_rp_reg[0]/P0001 ,
		_w2893_,
		_w2894_
	);
	LUT2 #(
		.INIT('h8)
	) name749 (
		\u7_rp_reg[0]/P0001 ,
		_w2893_,
		_w2895_
	);
	LUT2 #(
		.INIT('h2)
	) name750 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2894_,
		_w2896_
	);
	LUT2 #(
		.INIT('h4)
	) name751 (
		_w2895_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h2)
	) name752 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2759_,
		_w2898_
	);
	LUT2 #(
		.INIT('h8)
	) name753 (
		\u4_dout_reg[0]/P0001 ,
		_w2898_,
		_w2899_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		\u4_mem_reg[3][0]/NET0131 ,
		_w2765_,
		_w2900_
	);
	LUT2 #(
		.INIT('h4)
	) name755 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2901_
	);
	LUT2 #(
		.INIT('h8)
	) name756 (
		\u4_mem_reg[2][0]/NET0131 ,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h2)
	) name757 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2903_
	);
	LUT2 #(
		.INIT('h8)
	) name758 (
		\u4_mem_reg[1][0]/NET0131 ,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_rp_reg[2]/NET0131 ,
		_w2905_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		\u4_mem_reg[0][0]/NET0131 ,
		_w2905_,
		_w2906_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		_w2900_,
		_w2902_,
		_w2907_
	);
	LUT2 #(
		.INIT('h1)
	) name762 (
		_w2904_,
		_w2906_,
		_w2908_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		_w2907_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\u13_occ0_r_reg[11]/NET0131 ,
		_w2910_
	);
	LUT2 #(
		.INIT('h8)
	) name765 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w2910_,
		_w2911_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		_w2759_,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h4)
	) name767 (
		_w2909_,
		_w2912_,
		_w2913_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		_w2899_,
		_w2913_,
		_w2914_
	);
	LUT2 #(
		.INIT('h8)
	) name769 (
		\u4_dout_reg[1]/P0001 ,
		_w2898_,
		_w2915_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		\u4_mem_reg[3][1]/NET0131 ,
		_w2765_,
		_w2916_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		\u4_mem_reg[2][1]/NET0131 ,
		_w2901_,
		_w2917_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		\u4_mem_reg[1][1]/NET0131 ,
		_w2903_,
		_w2918_
	);
	LUT2 #(
		.INIT('h8)
	) name773 (
		\u4_mem_reg[0][1]/NET0131 ,
		_w2905_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w2916_,
		_w2917_,
		_w2920_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w2918_,
		_w2919_,
		_w2921_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		_w2920_,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h2)
	) name777 (
		_w2912_,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name778 (
		_w2915_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h2)
	) name779 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2770_,
		_w2925_
	);
	LUT2 #(
		.INIT('h8)
	) name780 (
		\u5_dout_reg[0]/P0001 ,
		_w2925_,
		_w2926_
	);
	LUT2 #(
		.INIT('h8)
	) name781 (
		\u5_mem_reg[3][0]/NET0131 ,
		_w2776_,
		_w2927_
	);
	LUT2 #(
		.INIT('h2)
	) name782 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2928_
	);
	LUT2 #(
		.INIT('h8)
	) name783 (
		\u5_mem_reg[1][0]/NET0131 ,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h4)
	) name784 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2930_
	);
	LUT2 #(
		.INIT('h8)
	) name785 (
		\u5_mem_reg[2][0]/NET0131 ,
		_w2930_,
		_w2931_
	);
	LUT2 #(
		.INIT('h1)
	) name786 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_rp_reg[2]/NET0131 ,
		_w2932_
	);
	LUT2 #(
		.INIT('h8)
	) name787 (
		\u5_mem_reg[0][0]/NET0131 ,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		_w2927_,
		_w2929_,
		_w2934_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		_w2931_,
		_w2933_,
		_w2935_
	);
	LUT2 #(
		.INIT('h8)
	) name790 (
		_w2934_,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('h4)
	) name791 (
		\u13_occ0_r_reg[18]/NET0131 ,
		\u13_occ0_r_reg[19]/NET0131 ,
		_w2937_
	);
	LUT2 #(
		.INIT('h8)
	) name792 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h8)
	) name793 (
		_w2770_,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h4)
	) name794 (
		_w2936_,
		_w2939_,
		_w2940_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w2926_,
		_w2940_,
		_w2941_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		\u5_dout_reg[1]/P0001 ,
		_w2925_,
		_w2942_
	);
	LUT2 #(
		.INIT('h8)
	) name797 (
		\u5_mem_reg[3][1]/NET0131 ,
		_w2776_,
		_w2943_
	);
	LUT2 #(
		.INIT('h8)
	) name798 (
		\u5_mem_reg[1][1]/NET0131 ,
		_w2928_,
		_w2944_
	);
	LUT2 #(
		.INIT('h8)
	) name799 (
		\u5_mem_reg[2][1]/NET0131 ,
		_w2930_,
		_w2945_
	);
	LUT2 #(
		.INIT('h8)
	) name800 (
		\u5_mem_reg[0][1]/NET0131 ,
		_w2932_,
		_w2946_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		_w2943_,
		_w2944_,
		_w2947_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		_w2945_,
		_w2946_,
		_w2948_
	);
	LUT2 #(
		.INIT('h8)
	) name803 (
		_w2947_,
		_w2948_,
		_w2949_
	);
	LUT2 #(
		.INIT('h2)
	) name804 (
		_w2939_,
		_w2949_,
		_w2950_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		_w2942_,
		_w2950_,
		_w2951_
	);
	LUT2 #(
		.INIT('h2)
	) name806 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2795_,
		_w2952_
	);
	LUT2 #(
		.INIT('h8)
	) name807 (
		\u6_dout_reg[0]/P0001 ,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h8)
	) name808 (
		\u6_mem_reg[3][0]/NET0131 ,
		_w2801_,
		_w2954_
	);
	LUT2 #(
		.INIT('h4)
	) name809 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2955_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		\u6_mem_reg[2][0]/NET0131 ,
		_w2955_,
		_w2956_
	);
	LUT2 #(
		.INIT('h2)
	) name811 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2957_
	);
	LUT2 #(
		.INIT('h8)
	) name812 (
		\u6_mem_reg[1][0]/NET0131 ,
		_w2957_,
		_w2958_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_rp_reg[2]/NET0131 ,
		_w2959_
	);
	LUT2 #(
		.INIT('h8)
	) name814 (
		\u6_mem_reg[0][0]/NET0131 ,
		_w2959_,
		_w2960_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w2954_,
		_w2956_,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w2958_,
		_w2960_,
		_w2962_
	);
	LUT2 #(
		.INIT('h8)
	) name817 (
		_w2961_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h4)
	) name818 (
		\u13_occ0_r_reg[26]/NET0131 ,
		\u13_occ0_r_reg[27]/NET0131 ,
		_w2964_
	);
	LUT2 #(
		.INIT('h8)
	) name819 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w2964_,
		_w2965_
	);
	LUT2 #(
		.INIT('h8)
	) name820 (
		_w2795_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h4)
	) name821 (
		_w2963_,
		_w2966_,
		_w2967_
	);
	LUT2 #(
		.INIT('h1)
	) name822 (
		_w2953_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h8)
	) name823 (
		\u6_dout_reg[1]/P0001 ,
		_w2952_,
		_w2969_
	);
	LUT2 #(
		.INIT('h8)
	) name824 (
		\u6_mem_reg[2][1]/NET0131 ,
		_w2955_,
		_w2970_
	);
	LUT2 #(
		.INIT('h8)
	) name825 (
		\u6_mem_reg[1][1]/NET0131 ,
		_w2957_,
		_w2971_
	);
	LUT2 #(
		.INIT('h8)
	) name826 (
		\u6_mem_reg[3][1]/NET0131 ,
		_w2801_,
		_w2972_
	);
	LUT2 #(
		.INIT('h8)
	) name827 (
		\u6_mem_reg[0][1]/NET0131 ,
		_w2959_,
		_w2973_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w2970_,
		_w2971_,
		_w2974_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w2972_,
		_w2973_,
		_w2975_
	);
	LUT2 #(
		.INIT('h8)
	) name830 (
		_w2974_,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		_w2966_,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		_w2969_,
		_w2977_,
		_w2978_
	);
	LUT2 #(
		.INIT('h2)
	) name833 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2808_,
		_w2979_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		\u7_dout_reg[0]/P0001 ,
		_w2979_,
		_w2980_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2981_
	);
	LUT2 #(
		.INIT('h8)
	) name836 (
		\u7_mem_reg[3][0]/NET0131 ,
		_w2981_,
		_w2982_
	);
	LUT2 #(
		.INIT('h4)
	) name837 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2983_
	);
	LUT2 #(
		.INIT('h8)
	) name838 (
		\u7_mem_reg[2][0]/NET0131 ,
		_w2983_,
		_w2984_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2985_
	);
	LUT2 #(
		.INIT('h8)
	) name840 (
		\u7_mem_reg[1][0]/NET0131 ,
		_w2985_,
		_w2986_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_rp_reg[2]/NET0131 ,
		_w2987_
	);
	LUT2 #(
		.INIT('h8)
	) name842 (
		\u7_mem_reg[0][0]/NET0131 ,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w2982_,
		_w2984_,
		_w2989_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		_w2986_,
		_w2988_,
		_w2990_
	);
	LUT2 #(
		.INIT('h8)
	) name845 (
		_w2989_,
		_w2990_,
		_w2991_
	);
	LUT2 #(
		.INIT('h4)
	) name846 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		_w2992_
	);
	LUT2 #(
		.INIT('h8)
	) name847 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w2992_,
		_w2993_
	);
	LUT2 #(
		.INIT('h8)
	) name848 (
		_w2808_,
		_w2993_,
		_w2994_
	);
	LUT2 #(
		.INIT('h4)
	) name849 (
		_w2991_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h1)
	) name850 (
		_w2980_,
		_w2995_,
		_w2996_
	);
	LUT2 #(
		.INIT('h8)
	) name851 (
		\u7_dout_reg[1]/P0001 ,
		_w2979_,
		_w2997_
	);
	LUT2 #(
		.INIT('h8)
	) name852 (
		\u7_mem_reg[3][1]/NET0131 ,
		_w2981_,
		_w2998_
	);
	LUT2 #(
		.INIT('h8)
	) name853 (
		\u7_mem_reg[2][1]/NET0131 ,
		_w2983_,
		_w2999_
	);
	LUT2 #(
		.INIT('h8)
	) name854 (
		\u7_mem_reg[1][1]/NET0131 ,
		_w2985_,
		_w3000_
	);
	LUT2 #(
		.INIT('h8)
	) name855 (
		\u7_mem_reg[0][1]/NET0131 ,
		_w2987_,
		_w3001_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w2998_,
		_w2999_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		_w3000_,
		_w3001_,
		_w3003_
	);
	LUT2 #(
		.INIT('h8)
	) name858 (
		_w3002_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h2)
	) name859 (
		_w2994_,
		_w3004_,
		_w3005_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w2997_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('h2)
	) name861 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w2787_,
		_w3007_
	);
	LUT2 #(
		.INIT('h8)
	) name862 (
		\u3_dout_reg[0]/P0001 ,
		_w3007_,
		_w3008_
	);
	LUT2 #(
		.INIT('h8)
	) name863 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3009_
	);
	LUT2 #(
		.INIT('h8)
	) name864 (
		\u3_mem_reg[3][0]/NET0131 ,
		_w3009_,
		_w3010_
	);
	LUT2 #(
		.INIT('h4)
	) name865 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3011_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\u3_mem_reg[2][0]/NET0131 ,
		_w3011_,
		_w3012_
	);
	LUT2 #(
		.INIT('h2)
	) name867 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3013_
	);
	LUT2 #(
		.INIT('h8)
	) name868 (
		\u3_mem_reg[1][0]/NET0131 ,
		_w3013_,
		_w3014_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_rp_reg[2]/NET0131 ,
		_w3015_
	);
	LUT2 #(
		.INIT('h8)
	) name870 (
		\u3_mem_reg[0][0]/NET0131 ,
		_w3015_,
		_w3016_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		_w3010_,
		_w3012_,
		_w3017_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w3014_,
		_w3016_,
		_w3018_
	);
	LUT2 #(
		.INIT('h8)
	) name873 (
		_w3017_,
		_w3018_,
		_w3019_
	);
	LUT2 #(
		.INIT('h4)
	) name874 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		_w3020_
	);
	LUT2 #(
		.INIT('h8)
	) name875 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w3020_,
		_w3021_
	);
	LUT2 #(
		.INIT('h8)
	) name876 (
		_w2787_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h4)
	) name877 (
		_w3019_,
		_w3022_,
		_w3023_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w3008_,
		_w3023_,
		_w3024_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w2159_,
		_w3025_
	);
	LUT2 #(
		.INIT('h8)
	) name880 (
		\u8_dout_reg[0]/P0001 ,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h8)
	) name881 (
		\u8_mem_reg[3][0]/NET0131 ,
		_w2163_,
		_w3027_
	);
	LUT2 #(
		.INIT('h4)
	) name882 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3028_
	);
	LUT2 #(
		.INIT('h8)
	) name883 (
		\u8_mem_reg[2][0]/NET0131 ,
		_w3028_,
		_w3029_
	);
	LUT2 #(
		.INIT('h2)
	) name884 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3030_
	);
	LUT2 #(
		.INIT('h8)
	) name885 (
		\u8_mem_reg[1][0]/NET0131 ,
		_w3030_,
		_w3031_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_rp_reg[2]/NET0131 ,
		_w3032_
	);
	LUT2 #(
		.INIT('h8)
	) name887 (
		\u8_mem_reg[0][0]/NET0131 ,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h1)
	) name888 (
		_w3027_,
		_w3029_,
		_w3034_
	);
	LUT2 #(
		.INIT('h1)
	) name889 (
		_w3031_,
		_w3033_,
		_w3035_
	);
	LUT2 #(
		.INIT('h8)
	) name890 (
		_w3034_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h4)
	) name891 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\u13_occ1_r_reg[11]/NET0131 ,
		_w3037_
	);
	LUT2 #(
		.INIT('h8)
	) name892 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w3037_,
		_w3038_
	);
	LUT2 #(
		.INIT('h8)
	) name893 (
		_w2159_,
		_w3038_,
		_w3039_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		_w3036_,
		_w3039_,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w3026_,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h8)
	) name896 (
		\u3_dout_reg[1]/P0001 ,
		_w3007_,
		_w3042_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		\u3_mem_reg[1][1]/NET0131 ,
		_w3013_,
		_w3043_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		\u3_mem_reg[2][1]/NET0131 ,
		_w3011_,
		_w3044_
	);
	LUT2 #(
		.INIT('h8)
	) name899 (
		\u3_mem_reg[3][1]/NET0131 ,
		_w3009_,
		_w3045_
	);
	LUT2 #(
		.INIT('h8)
	) name900 (
		\u3_mem_reg[0][1]/NET0131 ,
		_w3015_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w3043_,
		_w3044_,
		_w3047_
	);
	LUT2 #(
		.INIT('h1)
	) name902 (
		_w3045_,
		_w3046_,
		_w3048_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		_w3047_,
		_w3048_,
		_w3049_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		_w3022_,
		_w3049_,
		_w3050_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		_w3042_,
		_w3050_,
		_w3051_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		\u8_dout_reg[1]/P0001 ,
		_w3025_,
		_w3052_
	);
	LUT2 #(
		.INIT('h8)
	) name907 (
		\u8_mem_reg[3][1]/NET0131 ,
		_w2163_,
		_w3053_
	);
	LUT2 #(
		.INIT('h8)
	) name908 (
		\u8_mem_reg[2][1]/NET0131 ,
		_w3028_,
		_w3054_
	);
	LUT2 #(
		.INIT('h8)
	) name909 (
		\u8_mem_reg[1][1]/NET0131 ,
		_w3030_,
		_w3055_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		\u8_mem_reg[0][1]/NET0131 ,
		_w3032_,
		_w3056_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w3053_,
		_w3054_,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w3055_,
		_w3056_,
		_w3058_
	);
	LUT2 #(
		.INIT('h8)
	) name913 (
		_w3057_,
		_w3058_,
		_w3059_
	);
	LUT2 #(
		.INIT('h2)
	) name914 (
		_w3039_,
		_w3059_,
		_w3060_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w3052_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h8)
	) name916 (
		\in_valid_s_reg[2]/NET0131 ,
		\u14_u8_en_out_l_reg/NET0131 ,
		_w3062_
	);
	LUT2 #(
		.INIT('h4)
	) name917 (
		\u14_u8_en_out_l2_reg/P0001 ,
		_w3062_,
		_w3063_
	);
	LUT2 #(
		.INIT('h1)
	) name918 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w3064_
	);
	LUT2 #(
		.INIT('h4)
	) name919 (
		\u11_wp_reg[0]/NET0131 ,
		_w3064_,
		_w3065_
	);
	LUT2 #(
		.INIT('h2)
	) name920 (
		_w3063_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h8)
	) name921 (
		\u11_wp_reg[1]/P0001 ,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		\u11_wp_reg[2]/P0001 ,
		_w3067_,
		_w3068_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		\u11_wp_reg[2]/P0001 ,
		_w3067_,
		_w3069_
	);
	LUT2 #(
		.INIT('h2)
	) name924 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w3068_,
		_w3070_
	);
	LUT2 #(
		.INIT('h4)
	) name925 (
		_w3069_,
		_w3070_,
		_w3071_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		\u4_dout_reg[10]/P0001 ,
		_w2759_,
		_w3072_
	);
	LUT2 #(
		.INIT('h8)
	) name927 (
		\u4_mem_reg[3][6]/NET0131 ,
		_w2765_,
		_w3073_
	);
	LUT2 #(
		.INIT('h8)
	) name928 (
		\u4_mem_reg[2][6]/NET0131 ,
		_w2901_,
		_w3074_
	);
	LUT2 #(
		.INIT('h8)
	) name929 (
		\u4_mem_reg[0][6]/NET0131 ,
		_w2905_,
		_w3075_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		\u4_mem_reg[1][6]/NET0131 ,
		_w2903_,
		_w3076_
	);
	LUT2 #(
		.INIT('h1)
	) name931 (
		_w3073_,
		_w3074_,
		_w3077_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w3075_,
		_w3076_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name933 (
		_w3077_,
		_w3078_,
		_w3079_
	);
	LUT2 #(
		.INIT('h4)
	) name934 (
		\u4_rp_reg[0]/P0001 ,
		_w3079_,
		_w3080_
	);
	LUT2 #(
		.INIT('h8)
	) name935 (
		\u4_mem_reg[2][22]/NET0131 ,
		_w2901_,
		_w3081_
	);
	LUT2 #(
		.INIT('h8)
	) name936 (
		\u4_mem_reg[3][22]/NET0131 ,
		_w2765_,
		_w3082_
	);
	LUT2 #(
		.INIT('h8)
	) name937 (
		\u4_mem_reg[1][22]/NET0131 ,
		_w2903_,
		_w3083_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		\u4_mem_reg[0][22]/NET0131 ,
		_w2905_,
		_w3084_
	);
	LUT2 #(
		.INIT('h2)
	) name939 (
		\u4_rp_reg[0]/P0001 ,
		_w3081_,
		_w3085_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w3082_,
		_w3083_,
		_w3086_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w3084_,
		_w3086_,
		_w3087_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		_w3085_,
		_w3087_,
		_w3088_
	);
	LUT2 #(
		.INIT('h2)
	) name943 (
		_w2760_,
		_w3080_,
		_w3089_
	);
	LUT2 #(
		.INIT('h4)
	) name944 (
		_w3088_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h8)
	) name945 (
		\u4_mem_reg[3][10]/NET0131 ,
		_w2765_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name946 (
		\u4_mem_reg[2][10]/NET0131 ,
		_w2901_,
		_w3092_
	);
	LUT2 #(
		.INIT('h8)
	) name947 (
		\u4_mem_reg[0][10]/NET0131 ,
		_w2905_,
		_w3093_
	);
	LUT2 #(
		.INIT('h8)
	) name948 (
		\u4_mem_reg[1][10]/NET0131 ,
		_w2903_,
		_w3094_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w3091_,
		_w3092_,
		_w3095_
	);
	LUT2 #(
		.INIT('h1)
	) name950 (
		_w3093_,
		_w3094_,
		_w3096_
	);
	LUT2 #(
		.INIT('h8)
	) name951 (
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h2)
	) name952 (
		_w2910_,
		_w3097_,
		_w3098_
	);
	LUT2 #(
		.INIT('h2)
	) name953 (
		\u13_occ0_r_reg[10]/NET0131 ,
		\u13_occ0_r_reg[11]/NET0131 ,
		_w3099_
	);
	LUT2 #(
		.INIT('h8)
	) name954 (
		\u4_mem_reg[3][8]/NET0131 ,
		_w2765_,
		_w3100_
	);
	LUT2 #(
		.INIT('h8)
	) name955 (
		\u4_mem_reg[2][8]/NET0131 ,
		_w2901_,
		_w3101_
	);
	LUT2 #(
		.INIT('h8)
	) name956 (
		\u4_mem_reg[0][8]/NET0131 ,
		_w2905_,
		_w3102_
	);
	LUT2 #(
		.INIT('h8)
	) name957 (
		\u4_mem_reg[1][8]/NET0131 ,
		_w2903_,
		_w3103_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w3100_,
		_w3101_,
		_w3104_
	);
	LUT2 #(
		.INIT('h1)
	) name959 (
		_w3102_,
		_w3103_,
		_w3105_
	);
	LUT2 #(
		.INIT('h8)
	) name960 (
		_w3104_,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('h2)
	) name961 (
		_w3099_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h2)
	) name962 (
		_w2759_,
		_w3098_,
		_w3108_
	);
	LUT2 #(
		.INIT('h4)
	) name963 (
		_w3107_,
		_w3108_,
		_w3109_
	);
	LUT2 #(
		.INIT('h4)
	) name964 (
		_w3090_,
		_w3109_,
		_w3110_
	);
	LUT2 #(
		.INIT('h2)
	) name965 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3072_,
		_w3111_
	);
	LUT2 #(
		.INIT('h4)
	) name966 (
		_w3110_,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		\u4_dout_reg[11]/P0001 ,
		_w2759_,
		_w3113_
	);
	LUT2 #(
		.INIT('h8)
	) name968 (
		\u4_mem_reg[1][7]/NET0131 ,
		_w2903_,
		_w3114_
	);
	LUT2 #(
		.INIT('h8)
	) name969 (
		\u4_mem_reg[2][7]/NET0131 ,
		_w2901_,
		_w3115_
	);
	LUT2 #(
		.INIT('h8)
	) name970 (
		\u4_mem_reg[3][7]/NET0131 ,
		_w2765_,
		_w3116_
	);
	LUT2 #(
		.INIT('h8)
	) name971 (
		\u4_mem_reg[0][7]/NET0131 ,
		_w2905_,
		_w3117_
	);
	LUT2 #(
		.INIT('h1)
	) name972 (
		_w3114_,
		_w3115_,
		_w3118_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w3116_,
		_w3117_,
		_w3119_
	);
	LUT2 #(
		.INIT('h8)
	) name974 (
		_w3118_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h4)
	) name975 (
		\u4_rp_reg[0]/P0001 ,
		_w3120_,
		_w3121_
	);
	LUT2 #(
		.INIT('h8)
	) name976 (
		\u4_mem_reg[2][23]/NET0131 ,
		_w2901_,
		_w3122_
	);
	LUT2 #(
		.INIT('h8)
	) name977 (
		\u4_mem_reg[3][23]/NET0131 ,
		_w2765_,
		_w3123_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		\u4_mem_reg[1][23]/NET0131 ,
		_w2903_,
		_w3124_
	);
	LUT2 #(
		.INIT('h8)
	) name979 (
		\u4_mem_reg[0][23]/NET0131 ,
		_w2905_,
		_w3125_
	);
	LUT2 #(
		.INIT('h2)
	) name980 (
		\u4_rp_reg[0]/P0001 ,
		_w3122_,
		_w3126_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w3123_,
		_w3124_,
		_w3127_
	);
	LUT2 #(
		.INIT('h4)
	) name982 (
		_w3125_,
		_w3127_,
		_w3128_
	);
	LUT2 #(
		.INIT('h8)
	) name983 (
		_w3126_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h2)
	) name984 (
		_w2760_,
		_w3121_,
		_w3130_
	);
	LUT2 #(
		.INIT('h4)
	) name985 (
		_w3129_,
		_w3130_,
		_w3131_
	);
	LUT2 #(
		.INIT('h8)
	) name986 (
		\u4_mem_reg[3][11]/NET0131 ,
		_w2765_,
		_w3132_
	);
	LUT2 #(
		.INIT('h8)
	) name987 (
		\u4_mem_reg[1][11]/NET0131 ,
		_w2903_,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name988 (
		\u4_mem_reg[2][11]/NET0131 ,
		_w2901_,
		_w3134_
	);
	LUT2 #(
		.INIT('h8)
	) name989 (
		\u4_mem_reg[0][11]/NET0131 ,
		_w2905_,
		_w3135_
	);
	LUT2 #(
		.INIT('h1)
	) name990 (
		_w3132_,
		_w3133_,
		_w3136_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		_w3134_,
		_w3135_,
		_w3137_
	);
	LUT2 #(
		.INIT('h8)
	) name992 (
		_w3136_,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h2)
	) name993 (
		_w2910_,
		_w3138_,
		_w3139_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		\u4_mem_reg[1][9]/NET0131 ,
		_w2903_,
		_w3140_
	);
	LUT2 #(
		.INIT('h8)
	) name995 (
		\u4_mem_reg[3][9]/NET0131 ,
		_w2765_,
		_w3141_
	);
	LUT2 #(
		.INIT('h8)
	) name996 (
		\u4_mem_reg[2][9]/NET0131 ,
		_w2901_,
		_w3142_
	);
	LUT2 #(
		.INIT('h8)
	) name997 (
		\u4_mem_reg[0][9]/NET0131 ,
		_w2905_,
		_w3143_
	);
	LUT2 #(
		.INIT('h1)
	) name998 (
		_w3140_,
		_w3141_,
		_w3144_
	);
	LUT2 #(
		.INIT('h1)
	) name999 (
		_w3142_,
		_w3143_,
		_w3145_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		_w3144_,
		_w3145_,
		_w3146_
	);
	LUT2 #(
		.INIT('h2)
	) name1001 (
		_w3099_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h2)
	) name1002 (
		_w2759_,
		_w3139_,
		_w3148_
	);
	LUT2 #(
		.INIT('h4)
	) name1003 (
		_w3147_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		_w3131_,
		_w3149_,
		_w3150_
	);
	LUT2 #(
		.INIT('h2)
	) name1005 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3113_,
		_w3151_
	);
	LUT2 #(
		.INIT('h4)
	) name1006 (
		_w3150_,
		_w3151_,
		_w3152_
	);
	LUT2 #(
		.INIT('h1)
	) name1007 (
		\u4_dout_reg[12]/P0001 ,
		_w2759_,
		_w3153_
	);
	LUT2 #(
		.INIT('h4)
	) name1008 (
		\u4_rp_reg[0]/P0001 ,
		_w3106_,
		_w3154_
	);
	LUT2 #(
		.INIT('h8)
	) name1009 (
		\u4_mem_reg[2][24]/NET0131 ,
		_w2901_,
		_w3155_
	);
	LUT2 #(
		.INIT('h8)
	) name1010 (
		\u4_mem_reg[3][24]/NET0131 ,
		_w2765_,
		_w3156_
	);
	LUT2 #(
		.INIT('h8)
	) name1011 (
		\u4_mem_reg[1][24]/NET0131 ,
		_w2903_,
		_w3157_
	);
	LUT2 #(
		.INIT('h8)
	) name1012 (
		\u4_mem_reg[0][24]/NET0131 ,
		_w2905_,
		_w3158_
	);
	LUT2 #(
		.INIT('h2)
	) name1013 (
		\u4_rp_reg[0]/P0001 ,
		_w3155_,
		_w3159_
	);
	LUT2 #(
		.INIT('h1)
	) name1014 (
		_w3156_,
		_w3157_,
		_w3160_
	);
	LUT2 #(
		.INIT('h4)
	) name1015 (
		_w3158_,
		_w3160_,
		_w3161_
	);
	LUT2 #(
		.INIT('h8)
	) name1016 (
		_w3159_,
		_w3161_,
		_w3162_
	);
	LUT2 #(
		.INIT('h2)
	) name1017 (
		_w2760_,
		_w3154_,
		_w3163_
	);
	LUT2 #(
		.INIT('h4)
	) name1018 (
		_w3162_,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h8)
	) name1019 (
		\u4_mem_reg[3][12]/NET0131 ,
		_w2765_,
		_w3165_
	);
	LUT2 #(
		.INIT('h8)
	) name1020 (
		\u4_mem_reg[2][12]/NET0131 ,
		_w2901_,
		_w3166_
	);
	LUT2 #(
		.INIT('h8)
	) name1021 (
		\u4_mem_reg[0][12]/NET0131 ,
		_w2905_,
		_w3167_
	);
	LUT2 #(
		.INIT('h8)
	) name1022 (
		\u4_mem_reg[1][12]/NET0131 ,
		_w2903_,
		_w3168_
	);
	LUT2 #(
		.INIT('h1)
	) name1023 (
		_w3165_,
		_w3166_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w3167_,
		_w3168_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		_w3169_,
		_w3170_,
		_w3171_
	);
	LUT2 #(
		.INIT('h2)
	) name1026 (
		_w2910_,
		_w3171_,
		_w3172_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		_w3097_,
		_w3099_,
		_w3173_
	);
	LUT2 #(
		.INIT('h2)
	) name1028 (
		_w2759_,
		_w3172_,
		_w3174_
	);
	LUT2 #(
		.INIT('h4)
	) name1029 (
		_w3173_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h4)
	) name1030 (
		_w3164_,
		_w3175_,
		_w3176_
	);
	LUT2 #(
		.INIT('h2)
	) name1031 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3153_,
		_w3177_
	);
	LUT2 #(
		.INIT('h4)
	) name1032 (
		_w3176_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h1)
	) name1033 (
		\u4_dout_reg[13]/P0001 ,
		_w2759_,
		_w3179_
	);
	LUT2 #(
		.INIT('h4)
	) name1034 (
		\u4_rp_reg[0]/P0001 ,
		_w3146_,
		_w3180_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		\u4_mem_reg[2][25]/NET0131 ,
		_w2901_,
		_w3181_
	);
	LUT2 #(
		.INIT('h8)
	) name1036 (
		\u4_mem_reg[3][25]/NET0131 ,
		_w2765_,
		_w3182_
	);
	LUT2 #(
		.INIT('h8)
	) name1037 (
		\u4_mem_reg[1][25]/NET0131 ,
		_w2903_,
		_w3183_
	);
	LUT2 #(
		.INIT('h8)
	) name1038 (
		\u4_mem_reg[0][25]/NET0131 ,
		_w2905_,
		_w3184_
	);
	LUT2 #(
		.INIT('h2)
	) name1039 (
		\u4_rp_reg[0]/P0001 ,
		_w3181_,
		_w3185_
	);
	LUT2 #(
		.INIT('h1)
	) name1040 (
		_w3182_,
		_w3183_,
		_w3186_
	);
	LUT2 #(
		.INIT('h4)
	) name1041 (
		_w3184_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('h8)
	) name1042 (
		_w3185_,
		_w3187_,
		_w3188_
	);
	LUT2 #(
		.INIT('h2)
	) name1043 (
		_w2760_,
		_w3180_,
		_w3189_
	);
	LUT2 #(
		.INIT('h4)
	) name1044 (
		_w3188_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h8)
	) name1045 (
		\u4_mem_reg[1][13]/NET0131 ,
		_w2903_,
		_w3191_
	);
	LUT2 #(
		.INIT('h8)
	) name1046 (
		\u4_mem_reg[3][13]/NET0131 ,
		_w2765_,
		_w3192_
	);
	LUT2 #(
		.INIT('h8)
	) name1047 (
		\u4_mem_reg[2][13]/NET0131 ,
		_w2901_,
		_w3193_
	);
	LUT2 #(
		.INIT('h8)
	) name1048 (
		\u4_mem_reg[0][13]/NET0131 ,
		_w2905_,
		_w3194_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		_w3191_,
		_w3192_,
		_w3195_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		_w3193_,
		_w3194_,
		_w3196_
	);
	LUT2 #(
		.INIT('h8)
	) name1051 (
		_w3195_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h2)
	) name1052 (
		_w2910_,
		_w3197_,
		_w3198_
	);
	LUT2 #(
		.INIT('h2)
	) name1053 (
		_w3099_,
		_w3138_,
		_w3199_
	);
	LUT2 #(
		.INIT('h2)
	) name1054 (
		_w2759_,
		_w3198_,
		_w3200_
	);
	LUT2 #(
		.INIT('h4)
	) name1055 (
		_w3199_,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('h4)
	) name1056 (
		_w3190_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h2)
	) name1057 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3179_,
		_w3203_
	);
	LUT2 #(
		.INIT('h4)
	) name1058 (
		_w3202_,
		_w3203_,
		_w3204_
	);
	LUT2 #(
		.INIT('h1)
	) name1059 (
		\u4_dout_reg[14]/P0001 ,
		_w2759_,
		_w3205_
	);
	LUT2 #(
		.INIT('h4)
	) name1060 (
		\u4_rp_reg[0]/P0001 ,
		_w3097_,
		_w3206_
	);
	LUT2 #(
		.INIT('h8)
	) name1061 (
		\u4_mem_reg[2][26]/NET0131 ,
		_w2901_,
		_w3207_
	);
	LUT2 #(
		.INIT('h8)
	) name1062 (
		\u4_mem_reg[3][26]/NET0131 ,
		_w2765_,
		_w3208_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		\u4_mem_reg[1][26]/NET0131 ,
		_w2903_,
		_w3209_
	);
	LUT2 #(
		.INIT('h8)
	) name1064 (
		\u4_mem_reg[0][26]/NET0131 ,
		_w2905_,
		_w3210_
	);
	LUT2 #(
		.INIT('h2)
	) name1065 (
		\u4_rp_reg[0]/P0001 ,
		_w3207_,
		_w3211_
	);
	LUT2 #(
		.INIT('h1)
	) name1066 (
		_w3208_,
		_w3209_,
		_w3212_
	);
	LUT2 #(
		.INIT('h4)
	) name1067 (
		_w3210_,
		_w3212_,
		_w3213_
	);
	LUT2 #(
		.INIT('h8)
	) name1068 (
		_w3211_,
		_w3213_,
		_w3214_
	);
	LUT2 #(
		.INIT('h2)
	) name1069 (
		_w2760_,
		_w3206_,
		_w3215_
	);
	LUT2 #(
		.INIT('h4)
	) name1070 (
		_w3214_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h8)
	) name1071 (
		\u4_mem_reg[1][14]/NET0131 ,
		_w2903_,
		_w3217_
	);
	LUT2 #(
		.INIT('h8)
	) name1072 (
		\u4_mem_reg[2][14]/NET0131 ,
		_w2901_,
		_w3218_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		\u4_mem_reg[0][14]/NET0131 ,
		_w2905_,
		_w3219_
	);
	LUT2 #(
		.INIT('h8)
	) name1074 (
		\u4_mem_reg[3][14]/NET0131 ,
		_w2765_,
		_w3220_
	);
	LUT2 #(
		.INIT('h1)
	) name1075 (
		_w3217_,
		_w3218_,
		_w3221_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w3219_,
		_w3220_,
		_w3222_
	);
	LUT2 #(
		.INIT('h8)
	) name1077 (
		_w3221_,
		_w3222_,
		_w3223_
	);
	LUT2 #(
		.INIT('h2)
	) name1078 (
		_w2910_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('h2)
	) name1079 (
		_w3099_,
		_w3171_,
		_w3225_
	);
	LUT2 #(
		.INIT('h2)
	) name1080 (
		_w2759_,
		_w3224_,
		_w3226_
	);
	LUT2 #(
		.INIT('h4)
	) name1081 (
		_w3225_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h4)
	) name1082 (
		_w3216_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h2)
	) name1083 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3205_,
		_w3229_
	);
	LUT2 #(
		.INIT('h4)
	) name1084 (
		_w3228_,
		_w3229_,
		_w3230_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		\u4_dout_reg[15]/P0001 ,
		_w2759_,
		_w3231_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		\u4_rp_reg[0]/P0001 ,
		_w3138_,
		_w3232_
	);
	LUT2 #(
		.INIT('h8)
	) name1087 (
		\u4_mem_reg[2][27]/NET0131 ,
		_w2901_,
		_w3233_
	);
	LUT2 #(
		.INIT('h8)
	) name1088 (
		\u4_mem_reg[1][27]/NET0131 ,
		_w2903_,
		_w3234_
	);
	LUT2 #(
		.INIT('h8)
	) name1089 (
		\u4_mem_reg[3][27]/NET0131 ,
		_w2765_,
		_w3235_
	);
	LUT2 #(
		.INIT('h8)
	) name1090 (
		\u4_mem_reg[0][27]/NET0131 ,
		_w2905_,
		_w3236_
	);
	LUT2 #(
		.INIT('h2)
	) name1091 (
		\u4_rp_reg[0]/P0001 ,
		_w3233_,
		_w3237_
	);
	LUT2 #(
		.INIT('h1)
	) name1092 (
		_w3234_,
		_w3235_,
		_w3238_
	);
	LUT2 #(
		.INIT('h4)
	) name1093 (
		_w3236_,
		_w3238_,
		_w3239_
	);
	LUT2 #(
		.INIT('h8)
	) name1094 (
		_w3237_,
		_w3239_,
		_w3240_
	);
	LUT2 #(
		.INIT('h2)
	) name1095 (
		_w2760_,
		_w3232_,
		_w3241_
	);
	LUT2 #(
		.INIT('h4)
	) name1096 (
		_w3240_,
		_w3241_,
		_w3242_
	);
	LUT2 #(
		.INIT('h8)
	) name1097 (
		\u4_mem_reg[2][15]/NET0131 ,
		_w2901_,
		_w3243_
	);
	LUT2 #(
		.INIT('h8)
	) name1098 (
		\u4_mem_reg[0][15]/NET0131 ,
		_w2905_,
		_w3244_
	);
	LUT2 #(
		.INIT('h8)
	) name1099 (
		\u4_mem_reg[1][15]/NET0131 ,
		_w2903_,
		_w3245_
	);
	LUT2 #(
		.INIT('h8)
	) name1100 (
		\u4_mem_reg[3][15]/NET0131 ,
		_w2765_,
		_w3246_
	);
	LUT2 #(
		.INIT('h1)
	) name1101 (
		_w3243_,
		_w3244_,
		_w3247_
	);
	LUT2 #(
		.INIT('h1)
	) name1102 (
		_w3245_,
		_w3246_,
		_w3248_
	);
	LUT2 #(
		.INIT('h8)
	) name1103 (
		_w3247_,
		_w3248_,
		_w3249_
	);
	LUT2 #(
		.INIT('h2)
	) name1104 (
		_w2910_,
		_w3249_,
		_w3250_
	);
	LUT2 #(
		.INIT('h2)
	) name1105 (
		_w3099_,
		_w3197_,
		_w3251_
	);
	LUT2 #(
		.INIT('h2)
	) name1106 (
		_w2759_,
		_w3250_,
		_w3252_
	);
	LUT2 #(
		.INIT('h4)
	) name1107 (
		_w3251_,
		_w3252_,
		_w3253_
	);
	LUT2 #(
		.INIT('h4)
	) name1108 (
		_w3242_,
		_w3253_,
		_w3254_
	);
	LUT2 #(
		.INIT('h2)
	) name1109 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3231_,
		_w3255_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		_w3254_,
		_w3255_,
		_w3256_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		\u4_dout_reg[16]/P0001 ,
		_w2759_,
		_w3257_
	);
	LUT2 #(
		.INIT('h4)
	) name1112 (
		\u4_rp_reg[0]/P0001 ,
		_w3171_,
		_w3258_
	);
	LUT2 #(
		.INIT('h8)
	) name1113 (
		\u4_mem_reg[2][28]/NET0131 ,
		_w2901_,
		_w3259_
	);
	LUT2 #(
		.INIT('h8)
	) name1114 (
		\u4_mem_reg[1][28]/NET0131 ,
		_w2903_,
		_w3260_
	);
	LUT2 #(
		.INIT('h8)
	) name1115 (
		\u4_mem_reg[3][28]/NET0131 ,
		_w2765_,
		_w3261_
	);
	LUT2 #(
		.INIT('h8)
	) name1116 (
		\u4_mem_reg[0][28]/NET0131 ,
		_w2905_,
		_w3262_
	);
	LUT2 #(
		.INIT('h2)
	) name1117 (
		\u4_rp_reg[0]/P0001 ,
		_w3259_,
		_w3263_
	);
	LUT2 #(
		.INIT('h1)
	) name1118 (
		_w3260_,
		_w3261_,
		_w3264_
	);
	LUT2 #(
		.INIT('h4)
	) name1119 (
		_w3262_,
		_w3264_,
		_w3265_
	);
	LUT2 #(
		.INIT('h8)
	) name1120 (
		_w3263_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h2)
	) name1121 (
		_w2760_,
		_w3258_,
		_w3267_
	);
	LUT2 #(
		.INIT('h4)
	) name1122 (
		_w3266_,
		_w3267_,
		_w3268_
	);
	LUT2 #(
		.INIT('h8)
	) name1123 (
		\u4_mem_reg[3][16]/NET0131 ,
		_w2765_,
		_w3269_
	);
	LUT2 #(
		.INIT('h8)
	) name1124 (
		\u4_mem_reg[2][16]/NET0131 ,
		_w2901_,
		_w3270_
	);
	LUT2 #(
		.INIT('h8)
	) name1125 (
		\u4_mem_reg[0][16]/NET0131 ,
		_w2905_,
		_w3271_
	);
	LUT2 #(
		.INIT('h8)
	) name1126 (
		\u4_mem_reg[1][16]/NET0131 ,
		_w2903_,
		_w3272_
	);
	LUT2 #(
		.INIT('h1)
	) name1127 (
		_w3269_,
		_w3270_,
		_w3273_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w3271_,
		_w3272_,
		_w3274_
	);
	LUT2 #(
		.INIT('h8)
	) name1129 (
		_w3273_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h2)
	) name1130 (
		_w2910_,
		_w3275_,
		_w3276_
	);
	LUT2 #(
		.INIT('h2)
	) name1131 (
		_w3099_,
		_w3223_,
		_w3277_
	);
	LUT2 #(
		.INIT('h2)
	) name1132 (
		_w2759_,
		_w3276_,
		_w3278_
	);
	LUT2 #(
		.INIT('h4)
	) name1133 (
		_w3277_,
		_w3278_,
		_w3279_
	);
	LUT2 #(
		.INIT('h4)
	) name1134 (
		_w3268_,
		_w3279_,
		_w3280_
	);
	LUT2 #(
		.INIT('h2)
	) name1135 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3257_,
		_w3281_
	);
	LUT2 #(
		.INIT('h4)
	) name1136 (
		_w3280_,
		_w3281_,
		_w3282_
	);
	LUT2 #(
		.INIT('h1)
	) name1137 (
		\u4_dout_reg[17]/P0001 ,
		_w2759_,
		_w3283_
	);
	LUT2 #(
		.INIT('h4)
	) name1138 (
		\u4_rp_reg[0]/P0001 ,
		_w3197_,
		_w3284_
	);
	LUT2 #(
		.INIT('h8)
	) name1139 (
		\u4_mem_reg[2][29]/NET0131 ,
		_w2901_,
		_w3285_
	);
	LUT2 #(
		.INIT('h8)
	) name1140 (
		\u4_mem_reg[3][29]/NET0131 ,
		_w2765_,
		_w3286_
	);
	LUT2 #(
		.INIT('h8)
	) name1141 (
		\u4_mem_reg[1][29]/NET0131 ,
		_w2903_,
		_w3287_
	);
	LUT2 #(
		.INIT('h8)
	) name1142 (
		\u4_mem_reg[0][29]/NET0131 ,
		_w2905_,
		_w3288_
	);
	LUT2 #(
		.INIT('h2)
	) name1143 (
		\u4_rp_reg[0]/P0001 ,
		_w3285_,
		_w3289_
	);
	LUT2 #(
		.INIT('h1)
	) name1144 (
		_w3286_,
		_w3287_,
		_w3290_
	);
	LUT2 #(
		.INIT('h4)
	) name1145 (
		_w3288_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('h8)
	) name1146 (
		_w3289_,
		_w3291_,
		_w3292_
	);
	LUT2 #(
		.INIT('h2)
	) name1147 (
		_w2760_,
		_w3284_,
		_w3293_
	);
	LUT2 #(
		.INIT('h4)
	) name1148 (
		_w3292_,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('h8)
	) name1149 (
		\u4_mem_reg[3][17]/NET0131 ,
		_w2765_,
		_w3295_
	);
	LUT2 #(
		.INIT('h8)
	) name1150 (
		\u4_mem_reg[2][17]/NET0131 ,
		_w2901_,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		\u4_mem_reg[1][17]/NET0131 ,
		_w2903_,
		_w3297_
	);
	LUT2 #(
		.INIT('h8)
	) name1152 (
		\u4_mem_reg[0][17]/NET0131 ,
		_w2905_,
		_w3298_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		_w3295_,
		_w3296_,
		_w3299_
	);
	LUT2 #(
		.INIT('h1)
	) name1154 (
		_w3297_,
		_w3298_,
		_w3300_
	);
	LUT2 #(
		.INIT('h8)
	) name1155 (
		_w3299_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h2)
	) name1156 (
		_w2910_,
		_w3301_,
		_w3302_
	);
	LUT2 #(
		.INIT('h2)
	) name1157 (
		_w3099_,
		_w3249_,
		_w3303_
	);
	LUT2 #(
		.INIT('h2)
	) name1158 (
		_w2759_,
		_w3302_,
		_w3304_
	);
	LUT2 #(
		.INIT('h4)
	) name1159 (
		_w3303_,
		_w3304_,
		_w3305_
	);
	LUT2 #(
		.INIT('h4)
	) name1160 (
		_w3294_,
		_w3305_,
		_w3306_
	);
	LUT2 #(
		.INIT('h2)
	) name1161 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3283_,
		_w3307_
	);
	LUT2 #(
		.INIT('h4)
	) name1162 (
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h8)
	) name1163 (
		\in_valid_s_reg[0]/NET0131 ,
		\u14_u6_en_out_l_reg/NET0131 ,
		_w3309_
	);
	LUT2 #(
		.INIT('h4)
	) name1164 (
		\u14_u6_en_out_l2_reg/P0001 ,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h1)
	) name1165 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		_w3311_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		\u9_wp_reg[0]/NET0131 ,
		_w3311_,
		_w3312_
	);
	LUT2 #(
		.INIT('h2)
	) name1167 (
		_w3310_,
		_w3312_,
		_w3313_
	);
	LUT2 #(
		.INIT('h8)
	) name1168 (
		\u9_wp_reg[1]/P0001 ,
		_w3313_,
		_w3314_
	);
	LUT2 #(
		.INIT('h8)
	) name1169 (
		\u9_wp_reg[2]/P0001 ,
		_w3314_,
		_w3315_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		\u9_wp_reg[2]/P0001 ,
		_w3314_,
		_w3316_
	);
	LUT2 #(
		.INIT('h2)
	) name1171 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w3315_,
		_w3317_
	);
	LUT2 #(
		.INIT('h4)
	) name1172 (
		_w3316_,
		_w3317_,
		_w3318_
	);
	LUT2 #(
		.INIT('h1)
	) name1173 (
		\u4_dout_reg[18]/P0001 ,
		_w2759_,
		_w3319_
	);
	LUT2 #(
		.INIT('h4)
	) name1174 (
		\u4_rp_reg[0]/P0001 ,
		_w3223_,
		_w3320_
	);
	LUT2 #(
		.INIT('h8)
	) name1175 (
		\u4_mem_reg[2][30]/NET0131 ,
		_w2901_,
		_w3321_
	);
	LUT2 #(
		.INIT('h8)
	) name1176 (
		\u4_mem_reg[3][30]/NET0131 ,
		_w2765_,
		_w3322_
	);
	LUT2 #(
		.INIT('h8)
	) name1177 (
		\u4_mem_reg[1][30]/NET0131 ,
		_w2903_,
		_w3323_
	);
	LUT2 #(
		.INIT('h8)
	) name1178 (
		\u4_mem_reg[0][30]/NET0131 ,
		_w2905_,
		_w3324_
	);
	LUT2 #(
		.INIT('h2)
	) name1179 (
		\u4_rp_reg[0]/P0001 ,
		_w3321_,
		_w3325_
	);
	LUT2 #(
		.INIT('h1)
	) name1180 (
		_w3322_,
		_w3323_,
		_w3326_
	);
	LUT2 #(
		.INIT('h4)
	) name1181 (
		_w3324_,
		_w3326_,
		_w3327_
	);
	LUT2 #(
		.INIT('h8)
	) name1182 (
		_w3325_,
		_w3327_,
		_w3328_
	);
	LUT2 #(
		.INIT('h2)
	) name1183 (
		_w2760_,
		_w3320_,
		_w3329_
	);
	LUT2 #(
		.INIT('h4)
	) name1184 (
		_w3328_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h8)
	) name1185 (
		\u4_mem_reg[1][18]/NET0131 ,
		_w2903_,
		_w3331_
	);
	LUT2 #(
		.INIT('h8)
	) name1186 (
		\u4_mem_reg[3][18]/NET0131 ,
		_w2765_,
		_w3332_
	);
	LUT2 #(
		.INIT('h8)
	) name1187 (
		\u4_mem_reg[2][18]/NET0131 ,
		_w2901_,
		_w3333_
	);
	LUT2 #(
		.INIT('h8)
	) name1188 (
		\u4_mem_reg[0][18]/NET0131 ,
		_w2905_,
		_w3334_
	);
	LUT2 #(
		.INIT('h1)
	) name1189 (
		_w3331_,
		_w3332_,
		_w3335_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		_w3333_,
		_w3334_,
		_w3336_
	);
	LUT2 #(
		.INIT('h8)
	) name1191 (
		_w3335_,
		_w3336_,
		_w3337_
	);
	LUT2 #(
		.INIT('h2)
	) name1192 (
		_w2910_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h2)
	) name1193 (
		_w3099_,
		_w3275_,
		_w3339_
	);
	LUT2 #(
		.INIT('h2)
	) name1194 (
		_w2759_,
		_w3338_,
		_w3340_
	);
	LUT2 #(
		.INIT('h4)
	) name1195 (
		_w3339_,
		_w3340_,
		_w3341_
	);
	LUT2 #(
		.INIT('h4)
	) name1196 (
		_w3330_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h2)
	) name1197 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3319_,
		_w3343_
	);
	LUT2 #(
		.INIT('h4)
	) name1198 (
		_w3342_,
		_w3343_,
		_w3344_
	);
	LUT2 #(
		.INIT('h1)
	) name1199 (
		\u4_dout_reg[19]/P0001 ,
		_w2759_,
		_w3345_
	);
	LUT2 #(
		.INIT('h4)
	) name1200 (
		\u4_rp_reg[0]/P0001 ,
		_w3249_,
		_w3346_
	);
	LUT2 #(
		.INIT('h8)
	) name1201 (
		\u4_mem_reg[2][31]/NET0131 ,
		_w2901_,
		_w3347_
	);
	LUT2 #(
		.INIT('h8)
	) name1202 (
		\u4_mem_reg[3][31]/NET0131 ,
		_w2765_,
		_w3348_
	);
	LUT2 #(
		.INIT('h8)
	) name1203 (
		\u4_mem_reg[1][31]/NET0131 ,
		_w2903_,
		_w3349_
	);
	LUT2 #(
		.INIT('h8)
	) name1204 (
		\u4_mem_reg[0][31]/NET0131 ,
		_w2905_,
		_w3350_
	);
	LUT2 #(
		.INIT('h2)
	) name1205 (
		\u4_rp_reg[0]/P0001 ,
		_w3347_,
		_w3351_
	);
	LUT2 #(
		.INIT('h1)
	) name1206 (
		_w3348_,
		_w3349_,
		_w3352_
	);
	LUT2 #(
		.INIT('h4)
	) name1207 (
		_w3350_,
		_w3352_,
		_w3353_
	);
	LUT2 #(
		.INIT('h8)
	) name1208 (
		_w3351_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h2)
	) name1209 (
		_w2760_,
		_w3346_,
		_w3355_
	);
	LUT2 #(
		.INIT('h4)
	) name1210 (
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h8)
	) name1211 (
		\u4_mem_reg[3][19]/NET0131 ,
		_w2765_,
		_w3357_
	);
	LUT2 #(
		.INIT('h8)
	) name1212 (
		\u4_mem_reg[2][19]/NET0131 ,
		_w2901_,
		_w3358_
	);
	LUT2 #(
		.INIT('h8)
	) name1213 (
		\u4_mem_reg[1][19]/NET0131 ,
		_w2903_,
		_w3359_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		\u4_mem_reg[0][19]/NET0131 ,
		_w2905_,
		_w3360_
	);
	LUT2 #(
		.INIT('h1)
	) name1215 (
		_w3357_,
		_w3358_,
		_w3361_
	);
	LUT2 #(
		.INIT('h1)
	) name1216 (
		_w3359_,
		_w3360_,
		_w3362_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		_w3361_,
		_w3362_,
		_w3363_
	);
	LUT2 #(
		.INIT('h2)
	) name1218 (
		_w2910_,
		_w3363_,
		_w3364_
	);
	LUT2 #(
		.INIT('h2)
	) name1219 (
		_w3099_,
		_w3301_,
		_w3365_
	);
	LUT2 #(
		.INIT('h2)
	) name1220 (
		_w2759_,
		_w3364_,
		_w3366_
	);
	LUT2 #(
		.INIT('h4)
	) name1221 (
		_w3365_,
		_w3366_,
		_w3367_
	);
	LUT2 #(
		.INIT('h4)
	) name1222 (
		_w3356_,
		_w3367_,
		_w3368_
	);
	LUT2 #(
		.INIT('h2)
	) name1223 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3345_,
		_w3369_
	);
	LUT2 #(
		.INIT('h4)
	) name1224 (
		_w3368_,
		_w3369_,
		_w3370_
	);
	LUT2 #(
		.INIT('h1)
	) name1225 (
		\u4_dout_reg[2]/P0001 ,
		_w2759_,
		_w3371_
	);
	LUT2 #(
		.INIT('h4)
	) name1226 (
		_w2909_,
		_w3099_,
		_w3372_
	);
	LUT2 #(
		.INIT('h8)
	) name1227 (
		\u4_mem_reg[1][2]/NET0131 ,
		_w2903_,
		_w3373_
	);
	LUT2 #(
		.INIT('h8)
	) name1228 (
		\u4_mem_reg[0][2]/NET0131 ,
		_w2905_,
		_w3374_
	);
	LUT2 #(
		.INIT('h8)
	) name1229 (
		\u4_mem_reg[2][2]/NET0131 ,
		_w2901_,
		_w3375_
	);
	LUT2 #(
		.INIT('h8)
	) name1230 (
		\u4_mem_reg[3][2]/NET0131 ,
		_w2765_,
		_w3376_
	);
	LUT2 #(
		.INIT('h1)
	) name1231 (
		_w3373_,
		_w3374_,
		_w3377_
	);
	LUT2 #(
		.INIT('h1)
	) name1232 (
		_w3375_,
		_w3376_,
		_w3378_
	);
	LUT2 #(
		.INIT('h8)
	) name1233 (
		_w3377_,
		_w3378_,
		_w3379_
	);
	LUT2 #(
		.INIT('h2)
	) name1234 (
		_w2910_,
		_w3379_,
		_w3380_
	);
	LUT2 #(
		.INIT('h2)
	) name1235 (
		_w2759_,
		_w3372_,
		_w3381_
	);
	LUT2 #(
		.INIT('h4)
	) name1236 (
		_w3380_,
		_w3381_,
		_w3382_
	);
	LUT2 #(
		.INIT('h2)
	) name1237 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3371_,
		_w3383_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		_w3382_,
		_w3383_,
		_w3384_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		\u4_dout_reg[3]/P0001 ,
		_w2759_,
		_w3385_
	);
	LUT2 #(
		.INIT('h8)
	) name1240 (
		\u4_mem_reg[2][3]/NET0131 ,
		_w2901_,
		_w3386_
	);
	LUT2 #(
		.INIT('h8)
	) name1241 (
		\u4_mem_reg[3][3]/NET0131 ,
		_w2765_,
		_w3387_
	);
	LUT2 #(
		.INIT('h8)
	) name1242 (
		\u4_mem_reg[1][3]/NET0131 ,
		_w2903_,
		_w3388_
	);
	LUT2 #(
		.INIT('h8)
	) name1243 (
		\u4_mem_reg[0][3]/NET0131 ,
		_w2905_,
		_w3389_
	);
	LUT2 #(
		.INIT('h1)
	) name1244 (
		_w3386_,
		_w3387_,
		_w3390_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		_w3388_,
		_w3389_,
		_w3391_
	);
	LUT2 #(
		.INIT('h8)
	) name1246 (
		_w3390_,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h2)
	) name1247 (
		_w2910_,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h4)
	) name1248 (
		_w2922_,
		_w3099_,
		_w3394_
	);
	LUT2 #(
		.INIT('h2)
	) name1249 (
		_w2759_,
		_w3393_,
		_w3395_
	);
	LUT2 #(
		.INIT('h4)
	) name1250 (
		_w3394_,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h2)
	) name1251 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3385_,
		_w3397_
	);
	LUT2 #(
		.INIT('h4)
	) name1252 (
		_w3396_,
		_w3397_,
		_w3398_
	);
	LUT2 #(
		.INIT('h1)
	) name1253 (
		\u4_dout_reg[4]/P0001 ,
		_w2759_,
		_w3399_
	);
	LUT2 #(
		.INIT('h4)
	) name1254 (
		\u4_rp_reg[0]/P0001 ,
		_w2909_,
		_w3400_
	);
	LUT2 #(
		.INIT('h8)
	) name1255 (
		\u4_rp_reg[0]/P0001 ,
		_w3275_,
		_w3401_
	);
	LUT2 #(
		.INIT('h2)
	) name1256 (
		_w2760_,
		_w3400_,
		_w3402_
	);
	LUT2 #(
		.INIT('h4)
	) name1257 (
		_w3401_,
		_w3402_,
		_w3403_
	);
	LUT2 #(
		.INIT('h8)
	) name1258 (
		\u4_mem_reg[3][4]/NET0131 ,
		_w2765_,
		_w3404_
	);
	LUT2 #(
		.INIT('h8)
	) name1259 (
		\u4_mem_reg[2][4]/NET0131 ,
		_w2901_,
		_w3405_
	);
	LUT2 #(
		.INIT('h8)
	) name1260 (
		\u4_mem_reg[0][4]/NET0131 ,
		_w2905_,
		_w3406_
	);
	LUT2 #(
		.INIT('h8)
	) name1261 (
		\u4_mem_reg[1][4]/NET0131 ,
		_w2903_,
		_w3407_
	);
	LUT2 #(
		.INIT('h1)
	) name1262 (
		_w3404_,
		_w3405_,
		_w3408_
	);
	LUT2 #(
		.INIT('h1)
	) name1263 (
		_w3406_,
		_w3407_,
		_w3409_
	);
	LUT2 #(
		.INIT('h8)
	) name1264 (
		_w3408_,
		_w3409_,
		_w3410_
	);
	LUT2 #(
		.INIT('h2)
	) name1265 (
		_w2910_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h2)
	) name1266 (
		_w3099_,
		_w3379_,
		_w3412_
	);
	LUT2 #(
		.INIT('h2)
	) name1267 (
		_w2759_,
		_w3411_,
		_w3413_
	);
	LUT2 #(
		.INIT('h4)
	) name1268 (
		_w3412_,
		_w3413_,
		_w3414_
	);
	LUT2 #(
		.INIT('h4)
	) name1269 (
		_w3403_,
		_w3414_,
		_w3415_
	);
	LUT2 #(
		.INIT('h2)
	) name1270 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3399_,
		_w3416_
	);
	LUT2 #(
		.INIT('h4)
	) name1271 (
		_w3415_,
		_w3416_,
		_w3417_
	);
	LUT2 #(
		.INIT('h1)
	) name1272 (
		\u4_dout_reg[5]/P0001 ,
		_w2759_,
		_w3418_
	);
	LUT2 #(
		.INIT('h4)
	) name1273 (
		\u4_rp_reg[0]/P0001 ,
		_w2922_,
		_w3419_
	);
	LUT2 #(
		.INIT('h8)
	) name1274 (
		\u4_rp_reg[0]/P0001 ,
		_w3301_,
		_w3420_
	);
	LUT2 #(
		.INIT('h2)
	) name1275 (
		_w2760_,
		_w3419_,
		_w3421_
	);
	LUT2 #(
		.INIT('h4)
	) name1276 (
		_w3420_,
		_w3421_,
		_w3422_
	);
	LUT2 #(
		.INIT('h8)
	) name1277 (
		\u4_mem_reg[2][5]/NET0131 ,
		_w2901_,
		_w3423_
	);
	LUT2 #(
		.INIT('h8)
	) name1278 (
		\u4_mem_reg[1][5]/NET0131 ,
		_w2903_,
		_w3424_
	);
	LUT2 #(
		.INIT('h8)
	) name1279 (
		\u4_mem_reg[3][5]/NET0131 ,
		_w2765_,
		_w3425_
	);
	LUT2 #(
		.INIT('h8)
	) name1280 (
		\u4_mem_reg[0][5]/NET0131 ,
		_w2905_,
		_w3426_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w3423_,
		_w3424_,
		_w3427_
	);
	LUT2 #(
		.INIT('h1)
	) name1282 (
		_w3425_,
		_w3426_,
		_w3428_
	);
	LUT2 #(
		.INIT('h8)
	) name1283 (
		_w3427_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h2)
	) name1284 (
		_w2910_,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h2)
	) name1285 (
		_w3099_,
		_w3392_,
		_w3431_
	);
	LUT2 #(
		.INIT('h2)
	) name1286 (
		_w2759_,
		_w3430_,
		_w3432_
	);
	LUT2 #(
		.INIT('h4)
	) name1287 (
		_w3431_,
		_w3432_,
		_w3433_
	);
	LUT2 #(
		.INIT('h4)
	) name1288 (
		_w3422_,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h2)
	) name1289 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3418_,
		_w3435_
	);
	LUT2 #(
		.INIT('h4)
	) name1290 (
		_w3434_,
		_w3435_,
		_w3436_
	);
	LUT2 #(
		.INIT('h1)
	) name1291 (
		\u4_dout_reg[6]/P0001 ,
		_w2759_,
		_w3437_
	);
	LUT2 #(
		.INIT('h4)
	) name1292 (
		\u4_rp_reg[0]/P0001 ,
		_w3379_,
		_w3438_
	);
	LUT2 #(
		.INIT('h8)
	) name1293 (
		\u4_rp_reg[0]/P0001 ,
		_w3337_,
		_w3439_
	);
	LUT2 #(
		.INIT('h2)
	) name1294 (
		_w2760_,
		_w3438_,
		_w3440_
	);
	LUT2 #(
		.INIT('h4)
	) name1295 (
		_w3439_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h2)
	) name1296 (
		_w2910_,
		_w3079_,
		_w3442_
	);
	LUT2 #(
		.INIT('h2)
	) name1297 (
		_w3099_,
		_w3410_,
		_w3443_
	);
	LUT2 #(
		.INIT('h2)
	) name1298 (
		_w2759_,
		_w3442_,
		_w3444_
	);
	LUT2 #(
		.INIT('h4)
	) name1299 (
		_w3443_,
		_w3444_,
		_w3445_
	);
	LUT2 #(
		.INIT('h4)
	) name1300 (
		_w3441_,
		_w3445_,
		_w3446_
	);
	LUT2 #(
		.INIT('h2)
	) name1301 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3437_,
		_w3447_
	);
	LUT2 #(
		.INIT('h4)
	) name1302 (
		_w3446_,
		_w3447_,
		_w3448_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		\u4_dout_reg[7]/P0001 ,
		_w2759_,
		_w3449_
	);
	LUT2 #(
		.INIT('h4)
	) name1304 (
		\u4_rp_reg[0]/P0001 ,
		_w3392_,
		_w3450_
	);
	LUT2 #(
		.INIT('h8)
	) name1305 (
		\u4_rp_reg[0]/P0001 ,
		_w3363_,
		_w3451_
	);
	LUT2 #(
		.INIT('h2)
	) name1306 (
		_w2760_,
		_w3450_,
		_w3452_
	);
	LUT2 #(
		.INIT('h4)
	) name1307 (
		_w3451_,
		_w3452_,
		_w3453_
	);
	LUT2 #(
		.INIT('h2)
	) name1308 (
		_w2910_,
		_w3120_,
		_w3454_
	);
	LUT2 #(
		.INIT('h2)
	) name1309 (
		_w3099_,
		_w3429_,
		_w3455_
	);
	LUT2 #(
		.INIT('h2)
	) name1310 (
		_w2759_,
		_w3454_,
		_w3456_
	);
	LUT2 #(
		.INIT('h4)
	) name1311 (
		_w3455_,
		_w3456_,
		_w3457_
	);
	LUT2 #(
		.INIT('h4)
	) name1312 (
		_w3453_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h2)
	) name1313 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3449_,
		_w3459_
	);
	LUT2 #(
		.INIT('h4)
	) name1314 (
		_w3458_,
		_w3459_,
		_w3460_
	);
	LUT2 #(
		.INIT('h1)
	) name1315 (
		\u4_dout_reg[8]/P0001 ,
		_w2759_,
		_w3461_
	);
	LUT2 #(
		.INIT('h4)
	) name1316 (
		\u4_rp_reg[0]/P0001 ,
		_w3410_,
		_w3462_
	);
	LUT2 #(
		.INIT('h8)
	) name1317 (
		\u4_mem_reg[2][20]/NET0131 ,
		_w2901_,
		_w3463_
	);
	LUT2 #(
		.INIT('h8)
	) name1318 (
		\u4_mem_reg[3][20]/NET0131 ,
		_w2765_,
		_w3464_
	);
	LUT2 #(
		.INIT('h8)
	) name1319 (
		\u4_mem_reg[1][20]/NET0131 ,
		_w2903_,
		_w3465_
	);
	LUT2 #(
		.INIT('h8)
	) name1320 (
		\u4_mem_reg[0][20]/NET0131 ,
		_w2905_,
		_w3466_
	);
	LUT2 #(
		.INIT('h2)
	) name1321 (
		\u4_rp_reg[0]/P0001 ,
		_w3463_,
		_w3467_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w3464_,
		_w3465_,
		_w3468_
	);
	LUT2 #(
		.INIT('h4)
	) name1323 (
		_w3466_,
		_w3468_,
		_w3469_
	);
	LUT2 #(
		.INIT('h8)
	) name1324 (
		_w3467_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h2)
	) name1325 (
		_w2760_,
		_w3462_,
		_w3471_
	);
	LUT2 #(
		.INIT('h4)
	) name1326 (
		_w3470_,
		_w3471_,
		_w3472_
	);
	LUT2 #(
		.INIT('h2)
	) name1327 (
		_w2910_,
		_w3106_,
		_w3473_
	);
	LUT2 #(
		.INIT('h4)
	) name1328 (
		_w3079_,
		_w3099_,
		_w3474_
	);
	LUT2 #(
		.INIT('h2)
	) name1329 (
		_w2759_,
		_w3473_,
		_w3475_
	);
	LUT2 #(
		.INIT('h4)
	) name1330 (
		_w3474_,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h4)
	) name1331 (
		_w3472_,
		_w3476_,
		_w3477_
	);
	LUT2 #(
		.INIT('h2)
	) name1332 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3461_,
		_w3478_
	);
	LUT2 #(
		.INIT('h4)
	) name1333 (
		_w3477_,
		_w3478_,
		_w3479_
	);
	LUT2 #(
		.INIT('h1)
	) name1334 (
		\u4_dout_reg[9]/P0001 ,
		_w2759_,
		_w3480_
	);
	LUT2 #(
		.INIT('h4)
	) name1335 (
		\u4_rp_reg[0]/P0001 ,
		_w3429_,
		_w3481_
	);
	LUT2 #(
		.INIT('h8)
	) name1336 (
		\u4_mem_reg[2][21]/NET0131 ,
		_w2901_,
		_w3482_
	);
	LUT2 #(
		.INIT('h8)
	) name1337 (
		\u4_mem_reg[3][21]/NET0131 ,
		_w2765_,
		_w3483_
	);
	LUT2 #(
		.INIT('h8)
	) name1338 (
		\u4_mem_reg[1][21]/NET0131 ,
		_w2903_,
		_w3484_
	);
	LUT2 #(
		.INIT('h8)
	) name1339 (
		\u4_mem_reg[0][21]/NET0131 ,
		_w2905_,
		_w3485_
	);
	LUT2 #(
		.INIT('h2)
	) name1340 (
		\u4_rp_reg[0]/P0001 ,
		_w3482_,
		_w3486_
	);
	LUT2 #(
		.INIT('h1)
	) name1341 (
		_w3483_,
		_w3484_,
		_w3487_
	);
	LUT2 #(
		.INIT('h4)
	) name1342 (
		_w3485_,
		_w3487_,
		_w3488_
	);
	LUT2 #(
		.INIT('h8)
	) name1343 (
		_w3486_,
		_w3488_,
		_w3489_
	);
	LUT2 #(
		.INIT('h2)
	) name1344 (
		_w2760_,
		_w3481_,
		_w3490_
	);
	LUT2 #(
		.INIT('h4)
	) name1345 (
		_w3489_,
		_w3490_,
		_w3491_
	);
	LUT2 #(
		.INIT('h2)
	) name1346 (
		_w2910_,
		_w3146_,
		_w3492_
	);
	LUT2 #(
		.INIT('h2)
	) name1347 (
		_w3099_,
		_w3120_,
		_w3493_
	);
	LUT2 #(
		.INIT('h2)
	) name1348 (
		_w2759_,
		_w3492_,
		_w3494_
	);
	LUT2 #(
		.INIT('h4)
	) name1349 (
		_w3493_,
		_w3494_,
		_w3495_
	);
	LUT2 #(
		.INIT('h4)
	) name1350 (
		_w3491_,
		_w3495_,
		_w3496_
	);
	LUT2 #(
		.INIT('h2)
	) name1351 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w3480_,
		_w3497_
	);
	LUT2 #(
		.INIT('h4)
	) name1352 (
		_w3496_,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h8)
	) name1353 (
		\in_valid_s_reg[1]/NET0131 ,
		\u14_u7_en_out_l_reg/NET0131 ,
		_w3499_
	);
	LUT2 #(
		.INIT('h4)
	) name1354 (
		\u14_u7_en_out_l2_reg/P0001 ,
		_w3499_,
		_w3500_
	);
	LUT2 #(
		.INIT('h1)
	) name1355 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w3501_
	);
	LUT2 #(
		.INIT('h4)
	) name1356 (
		\u10_wp_reg[0]/NET0131 ,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h2)
	) name1357 (
		_w3500_,
		_w3502_,
		_w3503_
	);
	LUT2 #(
		.INIT('h8)
	) name1358 (
		\u10_wp_reg[1]/P0001 ,
		_w3503_,
		_w3504_
	);
	LUT2 #(
		.INIT('h8)
	) name1359 (
		\u10_wp_reg[2]/P0001 ,
		_w3504_,
		_w3505_
	);
	LUT2 #(
		.INIT('h1)
	) name1360 (
		\u10_wp_reg[2]/P0001 ,
		_w3504_,
		_w3506_
	);
	LUT2 #(
		.INIT('h2)
	) name1361 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w3505_,
		_w3507_
	);
	LUT2 #(
		.INIT('h4)
	) name1362 (
		_w3506_,
		_w3507_,
		_w3508_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		\u5_dout_reg[10]/P0001 ,
		_w2770_,
		_w3509_
	);
	LUT2 #(
		.INIT('h8)
	) name1364 (
		\u5_mem_reg[1][6]/NET0131 ,
		_w2928_,
		_w3510_
	);
	LUT2 #(
		.INIT('h8)
	) name1365 (
		\u5_mem_reg[2][6]/NET0131 ,
		_w2930_,
		_w3511_
	);
	LUT2 #(
		.INIT('h8)
	) name1366 (
		\u5_mem_reg[3][6]/NET0131 ,
		_w2776_,
		_w3512_
	);
	LUT2 #(
		.INIT('h8)
	) name1367 (
		\u5_mem_reg[0][6]/NET0131 ,
		_w2932_,
		_w3513_
	);
	LUT2 #(
		.INIT('h1)
	) name1368 (
		_w3510_,
		_w3511_,
		_w3514_
	);
	LUT2 #(
		.INIT('h1)
	) name1369 (
		_w3512_,
		_w3513_,
		_w3515_
	);
	LUT2 #(
		.INIT('h8)
	) name1370 (
		_w3514_,
		_w3515_,
		_w3516_
	);
	LUT2 #(
		.INIT('h4)
	) name1371 (
		\u5_rp_reg[0]/P0001 ,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h8)
	) name1372 (
		\u5_mem_reg[2][22]/NET0131 ,
		_w2930_,
		_w3518_
	);
	LUT2 #(
		.INIT('h8)
	) name1373 (
		\u5_mem_reg[3][22]/NET0131 ,
		_w2776_,
		_w3519_
	);
	LUT2 #(
		.INIT('h8)
	) name1374 (
		\u5_mem_reg[1][22]/NET0131 ,
		_w2928_,
		_w3520_
	);
	LUT2 #(
		.INIT('h8)
	) name1375 (
		\u5_mem_reg[0][22]/NET0131 ,
		_w2932_,
		_w3521_
	);
	LUT2 #(
		.INIT('h2)
	) name1376 (
		\u5_rp_reg[0]/P0001 ,
		_w3518_,
		_w3522_
	);
	LUT2 #(
		.INIT('h1)
	) name1377 (
		_w3519_,
		_w3520_,
		_w3523_
	);
	LUT2 #(
		.INIT('h4)
	) name1378 (
		_w3521_,
		_w3523_,
		_w3524_
	);
	LUT2 #(
		.INIT('h8)
	) name1379 (
		_w3522_,
		_w3524_,
		_w3525_
	);
	LUT2 #(
		.INIT('h2)
	) name1380 (
		_w2771_,
		_w3517_,
		_w3526_
	);
	LUT2 #(
		.INIT('h4)
	) name1381 (
		_w3525_,
		_w3526_,
		_w3527_
	);
	LUT2 #(
		.INIT('h8)
	) name1382 (
		\u5_mem_reg[2][10]/NET0131 ,
		_w2930_,
		_w3528_
	);
	LUT2 #(
		.INIT('h8)
	) name1383 (
		\u5_mem_reg[1][10]/NET0131 ,
		_w2928_,
		_w3529_
	);
	LUT2 #(
		.INIT('h8)
	) name1384 (
		\u5_mem_reg[3][10]/NET0131 ,
		_w2776_,
		_w3530_
	);
	LUT2 #(
		.INIT('h8)
	) name1385 (
		\u5_mem_reg[0][10]/NET0131 ,
		_w2932_,
		_w3531_
	);
	LUT2 #(
		.INIT('h1)
	) name1386 (
		_w3528_,
		_w3529_,
		_w3532_
	);
	LUT2 #(
		.INIT('h1)
	) name1387 (
		_w3530_,
		_w3531_,
		_w3533_
	);
	LUT2 #(
		.INIT('h8)
	) name1388 (
		_w3532_,
		_w3533_,
		_w3534_
	);
	LUT2 #(
		.INIT('h2)
	) name1389 (
		_w2937_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('h2)
	) name1390 (
		\u13_occ0_r_reg[18]/NET0131 ,
		\u13_occ0_r_reg[19]/NET0131 ,
		_w3536_
	);
	LUT2 #(
		.INIT('h8)
	) name1391 (
		\u5_mem_reg[2][8]/NET0131 ,
		_w2930_,
		_w3537_
	);
	LUT2 #(
		.INIT('h8)
	) name1392 (
		\u5_mem_reg[1][8]/NET0131 ,
		_w2928_,
		_w3538_
	);
	LUT2 #(
		.INIT('h8)
	) name1393 (
		\u5_mem_reg[3][8]/NET0131 ,
		_w2776_,
		_w3539_
	);
	LUT2 #(
		.INIT('h8)
	) name1394 (
		\u5_mem_reg[0][8]/NET0131 ,
		_w2932_,
		_w3540_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w3537_,
		_w3538_,
		_w3541_
	);
	LUT2 #(
		.INIT('h1)
	) name1396 (
		_w3539_,
		_w3540_,
		_w3542_
	);
	LUT2 #(
		.INIT('h8)
	) name1397 (
		_w3541_,
		_w3542_,
		_w3543_
	);
	LUT2 #(
		.INIT('h2)
	) name1398 (
		_w3536_,
		_w3543_,
		_w3544_
	);
	LUT2 #(
		.INIT('h2)
	) name1399 (
		_w2770_,
		_w3535_,
		_w3545_
	);
	LUT2 #(
		.INIT('h4)
	) name1400 (
		_w3544_,
		_w3545_,
		_w3546_
	);
	LUT2 #(
		.INIT('h4)
	) name1401 (
		_w3527_,
		_w3546_,
		_w3547_
	);
	LUT2 #(
		.INIT('h2)
	) name1402 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3509_,
		_w3548_
	);
	LUT2 #(
		.INIT('h4)
	) name1403 (
		_w3547_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h1)
	) name1404 (
		\u5_dout_reg[11]/P0001 ,
		_w2770_,
		_w3550_
	);
	LUT2 #(
		.INIT('h8)
	) name1405 (
		\u5_mem_reg[2][7]/NET0131 ,
		_w2930_,
		_w3551_
	);
	LUT2 #(
		.INIT('h8)
	) name1406 (
		\u5_mem_reg[1][7]/NET0131 ,
		_w2928_,
		_w3552_
	);
	LUT2 #(
		.INIT('h8)
	) name1407 (
		\u5_mem_reg[3][7]/NET0131 ,
		_w2776_,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name1408 (
		\u5_mem_reg[0][7]/NET0131 ,
		_w2932_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name1409 (
		_w3551_,
		_w3552_,
		_w3555_
	);
	LUT2 #(
		.INIT('h1)
	) name1410 (
		_w3553_,
		_w3554_,
		_w3556_
	);
	LUT2 #(
		.INIT('h8)
	) name1411 (
		_w3555_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h4)
	) name1412 (
		\u5_rp_reg[0]/P0001 ,
		_w3557_,
		_w3558_
	);
	LUT2 #(
		.INIT('h8)
	) name1413 (
		\u5_mem_reg[2][23]/NET0131 ,
		_w2930_,
		_w3559_
	);
	LUT2 #(
		.INIT('h8)
	) name1414 (
		\u5_mem_reg[3][23]/NET0131 ,
		_w2776_,
		_w3560_
	);
	LUT2 #(
		.INIT('h8)
	) name1415 (
		\u5_mem_reg[1][23]/NET0131 ,
		_w2928_,
		_w3561_
	);
	LUT2 #(
		.INIT('h8)
	) name1416 (
		\u5_mem_reg[0][23]/NET0131 ,
		_w2932_,
		_w3562_
	);
	LUT2 #(
		.INIT('h2)
	) name1417 (
		\u5_rp_reg[0]/P0001 ,
		_w3559_,
		_w3563_
	);
	LUT2 #(
		.INIT('h1)
	) name1418 (
		_w3560_,
		_w3561_,
		_w3564_
	);
	LUT2 #(
		.INIT('h4)
	) name1419 (
		_w3562_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h8)
	) name1420 (
		_w3563_,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('h2)
	) name1421 (
		_w2771_,
		_w3558_,
		_w3567_
	);
	LUT2 #(
		.INIT('h4)
	) name1422 (
		_w3566_,
		_w3567_,
		_w3568_
	);
	LUT2 #(
		.INIT('h8)
	) name1423 (
		\u5_mem_reg[2][11]/NET0131 ,
		_w2930_,
		_w3569_
	);
	LUT2 #(
		.INIT('h8)
	) name1424 (
		\u5_mem_reg[1][11]/NET0131 ,
		_w2928_,
		_w3570_
	);
	LUT2 #(
		.INIT('h8)
	) name1425 (
		\u5_mem_reg[3][11]/NET0131 ,
		_w2776_,
		_w3571_
	);
	LUT2 #(
		.INIT('h8)
	) name1426 (
		\u5_mem_reg[0][11]/NET0131 ,
		_w2932_,
		_w3572_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		_w3569_,
		_w3570_,
		_w3573_
	);
	LUT2 #(
		.INIT('h1)
	) name1428 (
		_w3571_,
		_w3572_,
		_w3574_
	);
	LUT2 #(
		.INIT('h8)
	) name1429 (
		_w3573_,
		_w3574_,
		_w3575_
	);
	LUT2 #(
		.INIT('h2)
	) name1430 (
		_w2937_,
		_w3575_,
		_w3576_
	);
	LUT2 #(
		.INIT('h8)
	) name1431 (
		\u5_mem_reg[1][9]/NET0131 ,
		_w2928_,
		_w3577_
	);
	LUT2 #(
		.INIT('h8)
	) name1432 (
		\u5_mem_reg[2][9]/NET0131 ,
		_w2930_,
		_w3578_
	);
	LUT2 #(
		.INIT('h8)
	) name1433 (
		\u5_mem_reg[3][9]/NET0131 ,
		_w2776_,
		_w3579_
	);
	LUT2 #(
		.INIT('h8)
	) name1434 (
		\u5_mem_reg[0][9]/NET0131 ,
		_w2932_,
		_w3580_
	);
	LUT2 #(
		.INIT('h1)
	) name1435 (
		_w3577_,
		_w3578_,
		_w3581_
	);
	LUT2 #(
		.INIT('h1)
	) name1436 (
		_w3579_,
		_w3580_,
		_w3582_
	);
	LUT2 #(
		.INIT('h8)
	) name1437 (
		_w3581_,
		_w3582_,
		_w3583_
	);
	LUT2 #(
		.INIT('h2)
	) name1438 (
		_w3536_,
		_w3583_,
		_w3584_
	);
	LUT2 #(
		.INIT('h2)
	) name1439 (
		_w2770_,
		_w3576_,
		_w3585_
	);
	LUT2 #(
		.INIT('h4)
	) name1440 (
		_w3584_,
		_w3585_,
		_w3586_
	);
	LUT2 #(
		.INIT('h4)
	) name1441 (
		_w3568_,
		_w3586_,
		_w3587_
	);
	LUT2 #(
		.INIT('h2)
	) name1442 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3550_,
		_w3588_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		_w3587_,
		_w3588_,
		_w3589_
	);
	LUT2 #(
		.INIT('h1)
	) name1444 (
		\u5_dout_reg[12]/P0001 ,
		_w2770_,
		_w3590_
	);
	LUT2 #(
		.INIT('h4)
	) name1445 (
		\u5_rp_reg[0]/P0001 ,
		_w3543_,
		_w3591_
	);
	LUT2 #(
		.INIT('h8)
	) name1446 (
		\u5_mem_reg[2][24]/NET0131 ,
		_w2930_,
		_w3592_
	);
	LUT2 #(
		.INIT('h8)
	) name1447 (
		\u5_mem_reg[3][24]/NET0131 ,
		_w2776_,
		_w3593_
	);
	LUT2 #(
		.INIT('h8)
	) name1448 (
		\u5_mem_reg[1][24]/NET0131 ,
		_w2928_,
		_w3594_
	);
	LUT2 #(
		.INIT('h8)
	) name1449 (
		\u5_mem_reg[0][24]/NET0131 ,
		_w2932_,
		_w3595_
	);
	LUT2 #(
		.INIT('h2)
	) name1450 (
		\u5_rp_reg[0]/P0001 ,
		_w3592_,
		_w3596_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w3593_,
		_w3594_,
		_w3597_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		_w3595_,
		_w3597_,
		_w3598_
	);
	LUT2 #(
		.INIT('h8)
	) name1453 (
		_w3596_,
		_w3598_,
		_w3599_
	);
	LUT2 #(
		.INIT('h2)
	) name1454 (
		_w2771_,
		_w3591_,
		_w3600_
	);
	LUT2 #(
		.INIT('h4)
	) name1455 (
		_w3599_,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h8)
	) name1456 (
		\u5_mem_reg[1][12]/NET0131 ,
		_w2928_,
		_w3602_
	);
	LUT2 #(
		.INIT('h8)
	) name1457 (
		\u5_mem_reg[2][12]/NET0131 ,
		_w2930_,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name1458 (
		\u5_mem_reg[3][12]/NET0131 ,
		_w2776_,
		_w3604_
	);
	LUT2 #(
		.INIT('h8)
	) name1459 (
		\u5_mem_reg[0][12]/NET0131 ,
		_w2932_,
		_w3605_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w3602_,
		_w3603_,
		_w3606_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w3604_,
		_w3605_,
		_w3607_
	);
	LUT2 #(
		.INIT('h8)
	) name1462 (
		_w3606_,
		_w3607_,
		_w3608_
	);
	LUT2 #(
		.INIT('h2)
	) name1463 (
		_w2937_,
		_w3608_,
		_w3609_
	);
	LUT2 #(
		.INIT('h4)
	) name1464 (
		_w3534_,
		_w3536_,
		_w3610_
	);
	LUT2 #(
		.INIT('h2)
	) name1465 (
		_w2770_,
		_w3609_,
		_w3611_
	);
	LUT2 #(
		.INIT('h4)
	) name1466 (
		_w3610_,
		_w3611_,
		_w3612_
	);
	LUT2 #(
		.INIT('h4)
	) name1467 (
		_w3601_,
		_w3612_,
		_w3613_
	);
	LUT2 #(
		.INIT('h2)
	) name1468 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3590_,
		_w3614_
	);
	LUT2 #(
		.INIT('h4)
	) name1469 (
		_w3613_,
		_w3614_,
		_w3615_
	);
	LUT2 #(
		.INIT('h1)
	) name1470 (
		\u5_dout_reg[13]/P0001 ,
		_w2770_,
		_w3616_
	);
	LUT2 #(
		.INIT('h4)
	) name1471 (
		\u5_rp_reg[0]/P0001 ,
		_w3583_,
		_w3617_
	);
	LUT2 #(
		.INIT('h8)
	) name1472 (
		\u5_mem_reg[2][25]/NET0131 ,
		_w2930_,
		_w3618_
	);
	LUT2 #(
		.INIT('h8)
	) name1473 (
		\u5_mem_reg[3][25]/NET0131 ,
		_w2776_,
		_w3619_
	);
	LUT2 #(
		.INIT('h8)
	) name1474 (
		\u5_mem_reg[1][25]/NET0131 ,
		_w2928_,
		_w3620_
	);
	LUT2 #(
		.INIT('h8)
	) name1475 (
		\u5_mem_reg[0][25]/NET0131 ,
		_w2932_,
		_w3621_
	);
	LUT2 #(
		.INIT('h2)
	) name1476 (
		\u5_rp_reg[0]/P0001 ,
		_w3618_,
		_w3622_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		_w3619_,
		_w3620_,
		_w3623_
	);
	LUT2 #(
		.INIT('h4)
	) name1478 (
		_w3621_,
		_w3623_,
		_w3624_
	);
	LUT2 #(
		.INIT('h8)
	) name1479 (
		_w3622_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('h2)
	) name1480 (
		_w2771_,
		_w3617_,
		_w3626_
	);
	LUT2 #(
		.INIT('h4)
	) name1481 (
		_w3625_,
		_w3626_,
		_w3627_
	);
	LUT2 #(
		.INIT('h8)
	) name1482 (
		\u5_mem_reg[1][13]/NET0131 ,
		_w2928_,
		_w3628_
	);
	LUT2 #(
		.INIT('h8)
	) name1483 (
		\u5_mem_reg[2][13]/NET0131 ,
		_w2930_,
		_w3629_
	);
	LUT2 #(
		.INIT('h8)
	) name1484 (
		\u5_mem_reg[3][13]/NET0131 ,
		_w2776_,
		_w3630_
	);
	LUT2 #(
		.INIT('h8)
	) name1485 (
		\u5_mem_reg[0][13]/NET0131 ,
		_w2932_,
		_w3631_
	);
	LUT2 #(
		.INIT('h1)
	) name1486 (
		_w3628_,
		_w3629_,
		_w3632_
	);
	LUT2 #(
		.INIT('h1)
	) name1487 (
		_w3630_,
		_w3631_,
		_w3633_
	);
	LUT2 #(
		.INIT('h8)
	) name1488 (
		_w3632_,
		_w3633_,
		_w3634_
	);
	LUT2 #(
		.INIT('h2)
	) name1489 (
		_w2937_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h2)
	) name1490 (
		_w3536_,
		_w3575_,
		_w3636_
	);
	LUT2 #(
		.INIT('h2)
	) name1491 (
		_w2770_,
		_w3635_,
		_w3637_
	);
	LUT2 #(
		.INIT('h4)
	) name1492 (
		_w3636_,
		_w3637_,
		_w3638_
	);
	LUT2 #(
		.INIT('h4)
	) name1493 (
		_w3627_,
		_w3638_,
		_w3639_
	);
	LUT2 #(
		.INIT('h2)
	) name1494 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3616_,
		_w3640_
	);
	LUT2 #(
		.INIT('h4)
	) name1495 (
		_w3639_,
		_w3640_,
		_w3641_
	);
	LUT2 #(
		.INIT('h1)
	) name1496 (
		\u5_dout_reg[14]/P0001 ,
		_w2770_,
		_w3642_
	);
	LUT2 #(
		.INIT('h4)
	) name1497 (
		\u5_rp_reg[0]/P0001 ,
		_w3534_,
		_w3643_
	);
	LUT2 #(
		.INIT('h8)
	) name1498 (
		\u5_mem_reg[2][26]/NET0131 ,
		_w2930_,
		_w3644_
	);
	LUT2 #(
		.INIT('h8)
	) name1499 (
		\u5_mem_reg[3][26]/NET0131 ,
		_w2776_,
		_w3645_
	);
	LUT2 #(
		.INIT('h8)
	) name1500 (
		\u5_mem_reg[1][26]/NET0131 ,
		_w2928_,
		_w3646_
	);
	LUT2 #(
		.INIT('h8)
	) name1501 (
		\u5_mem_reg[0][26]/NET0131 ,
		_w2932_,
		_w3647_
	);
	LUT2 #(
		.INIT('h2)
	) name1502 (
		\u5_rp_reg[0]/P0001 ,
		_w3644_,
		_w3648_
	);
	LUT2 #(
		.INIT('h1)
	) name1503 (
		_w3645_,
		_w3646_,
		_w3649_
	);
	LUT2 #(
		.INIT('h4)
	) name1504 (
		_w3647_,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h8)
	) name1505 (
		_w3648_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h2)
	) name1506 (
		_w2771_,
		_w3643_,
		_w3652_
	);
	LUT2 #(
		.INIT('h4)
	) name1507 (
		_w3651_,
		_w3652_,
		_w3653_
	);
	LUT2 #(
		.INIT('h8)
	) name1508 (
		\u5_mem_reg[2][14]/NET0131 ,
		_w2930_,
		_w3654_
	);
	LUT2 #(
		.INIT('h8)
	) name1509 (
		\u5_mem_reg[3][14]/NET0131 ,
		_w2776_,
		_w3655_
	);
	LUT2 #(
		.INIT('h8)
	) name1510 (
		\u5_mem_reg[0][14]/NET0131 ,
		_w2932_,
		_w3656_
	);
	LUT2 #(
		.INIT('h8)
	) name1511 (
		\u5_mem_reg[1][14]/NET0131 ,
		_w2928_,
		_w3657_
	);
	LUT2 #(
		.INIT('h1)
	) name1512 (
		_w3654_,
		_w3655_,
		_w3658_
	);
	LUT2 #(
		.INIT('h1)
	) name1513 (
		_w3656_,
		_w3657_,
		_w3659_
	);
	LUT2 #(
		.INIT('h8)
	) name1514 (
		_w3658_,
		_w3659_,
		_w3660_
	);
	LUT2 #(
		.INIT('h2)
	) name1515 (
		_w2937_,
		_w3660_,
		_w3661_
	);
	LUT2 #(
		.INIT('h2)
	) name1516 (
		_w3536_,
		_w3608_,
		_w3662_
	);
	LUT2 #(
		.INIT('h2)
	) name1517 (
		_w2770_,
		_w3661_,
		_w3663_
	);
	LUT2 #(
		.INIT('h4)
	) name1518 (
		_w3662_,
		_w3663_,
		_w3664_
	);
	LUT2 #(
		.INIT('h4)
	) name1519 (
		_w3653_,
		_w3664_,
		_w3665_
	);
	LUT2 #(
		.INIT('h2)
	) name1520 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3642_,
		_w3666_
	);
	LUT2 #(
		.INIT('h4)
	) name1521 (
		_w3665_,
		_w3666_,
		_w3667_
	);
	LUT2 #(
		.INIT('h1)
	) name1522 (
		\u5_dout_reg[15]/P0001 ,
		_w2770_,
		_w3668_
	);
	LUT2 #(
		.INIT('h4)
	) name1523 (
		\u5_rp_reg[0]/P0001 ,
		_w3575_,
		_w3669_
	);
	LUT2 #(
		.INIT('h8)
	) name1524 (
		\u5_mem_reg[2][27]/NET0131 ,
		_w2930_,
		_w3670_
	);
	LUT2 #(
		.INIT('h8)
	) name1525 (
		\u5_mem_reg[3][27]/NET0131 ,
		_w2776_,
		_w3671_
	);
	LUT2 #(
		.INIT('h8)
	) name1526 (
		\u5_mem_reg[1][27]/NET0131 ,
		_w2928_,
		_w3672_
	);
	LUT2 #(
		.INIT('h8)
	) name1527 (
		\u5_mem_reg[0][27]/NET0131 ,
		_w2932_,
		_w3673_
	);
	LUT2 #(
		.INIT('h2)
	) name1528 (
		\u5_rp_reg[0]/P0001 ,
		_w3670_,
		_w3674_
	);
	LUT2 #(
		.INIT('h1)
	) name1529 (
		_w3671_,
		_w3672_,
		_w3675_
	);
	LUT2 #(
		.INIT('h4)
	) name1530 (
		_w3673_,
		_w3675_,
		_w3676_
	);
	LUT2 #(
		.INIT('h8)
	) name1531 (
		_w3674_,
		_w3676_,
		_w3677_
	);
	LUT2 #(
		.INIT('h2)
	) name1532 (
		_w2771_,
		_w3669_,
		_w3678_
	);
	LUT2 #(
		.INIT('h4)
	) name1533 (
		_w3677_,
		_w3678_,
		_w3679_
	);
	LUT2 #(
		.INIT('h8)
	) name1534 (
		\u5_mem_reg[1][15]/NET0131 ,
		_w2928_,
		_w3680_
	);
	LUT2 #(
		.INIT('h8)
	) name1535 (
		\u5_mem_reg[3][15]/NET0131 ,
		_w2776_,
		_w3681_
	);
	LUT2 #(
		.INIT('h8)
	) name1536 (
		\u5_mem_reg[2][15]/NET0131 ,
		_w2930_,
		_w3682_
	);
	LUT2 #(
		.INIT('h8)
	) name1537 (
		\u5_mem_reg[0][15]/NET0131 ,
		_w2932_,
		_w3683_
	);
	LUT2 #(
		.INIT('h1)
	) name1538 (
		_w3680_,
		_w3681_,
		_w3684_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		_w3682_,
		_w3683_,
		_w3685_
	);
	LUT2 #(
		.INIT('h8)
	) name1540 (
		_w3684_,
		_w3685_,
		_w3686_
	);
	LUT2 #(
		.INIT('h2)
	) name1541 (
		_w2937_,
		_w3686_,
		_w3687_
	);
	LUT2 #(
		.INIT('h2)
	) name1542 (
		_w3536_,
		_w3634_,
		_w3688_
	);
	LUT2 #(
		.INIT('h2)
	) name1543 (
		_w2770_,
		_w3687_,
		_w3689_
	);
	LUT2 #(
		.INIT('h4)
	) name1544 (
		_w3688_,
		_w3689_,
		_w3690_
	);
	LUT2 #(
		.INIT('h4)
	) name1545 (
		_w3679_,
		_w3690_,
		_w3691_
	);
	LUT2 #(
		.INIT('h2)
	) name1546 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3668_,
		_w3692_
	);
	LUT2 #(
		.INIT('h4)
	) name1547 (
		_w3691_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h1)
	) name1548 (
		\u5_dout_reg[16]/P0001 ,
		_w2770_,
		_w3694_
	);
	LUT2 #(
		.INIT('h4)
	) name1549 (
		\u5_rp_reg[0]/P0001 ,
		_w3608_,
		_w3695_
	);
	LUT2 #(
		.INIT('h8)
	) name1550 (
		\u5_mem_reg[2][28]/NET0131 ,
		_w2930_,
		_w3696_
	);
	LUT2 #(
		.INIT('h8)
	) name1551 (
		\u5_mem_reg[3][28]/NET0131 ,
		_w2776_,
		_w3697_
	);
	LUT2 #(
		.INIT('h8)
	) name1552 (
		\u5_mem_reg[1][28]/NET0131 ,
		_w2928_,
		_w3698_
	);
	LUT2 #(
		.INIT('h8)
	) name1553 (
		\u5_mem_reg[0][28]/NET0131 ,
		_w2932_,
		_w3699_
	);
	LUT2 #(
		.INIT('h2)
	) name1554 (
		\u5_rp_reg[0]/P0001 ,
		_w3696_,
		_w3700_
	);
	LUT2 #(
		.INIT('h1)
	) name1555 (
		_w3697_,
		_w3698_,
		_w3701_
	);
	LUT2 #(
		.INIT('h4)
	) name1556 (
		_w3699_,
		_w3701_,
		_w3702_
	);
	LUT2 #(
		.INIT('h8)
	) name1557 (
		_w3700_,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h2)
	) name1558 (
		_w2771_,
		_w3695_,
		_w3704_
	);
	LUT2 #(
		.INIT('h4)
	) name1559 (
		_w3703_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h8)
	) name1560 (
		\u5_mem_reg[1][16]/NET0131 ,
		_w2928_,
		_w3706_
	);
	LUT2 #(
		.INIT('h8)
	) name1561 (
		\u5_mem_reg[3][16]/NET0131 ,
		_w2776_,
		_w3707_
	);
	LUT2 #(
		.INIT('h8)
	) name1562 (
		\u5_mem_reg[2][16]/NET0131 ,
		_w2930_,
		_w3708_
	);
	LUT2 #(
		.INIT('h8)
	) name1563 (
		\u5_mem_reg[0][16]/NET0131 ,
		_w2932_,
		_w3709_
	);
	LUT2 #(
		.INIT('h1)
	) name1564 (
		_w3706_,
		_w3707_,
		_w3710_
	);
	LUT2 #(
		.INIT('h1)
	) name1565 (
		_w3708_,
		_w3709_,
		_w3711_
	);
	LUT2 #(
		.INIT('h8)
	) name1566 (
		_w3710_,
		_w3711_,
		_w3712_
	);
	LUT2 #(
		.INIT('h2)
	) name1567 (
		_w2937_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		_w3536_,
		_w3660_,
		_w3714_
	);
	LUT2 #(
		.INIT('h2)
	) name1569 (
		_w2770_,
		_w3713_,
		_w3715_
	);
	LUT2 #(
		.INIT('h4)
	) name1570 (
		_w3714_,
		_w3715_,
		_w3716_
	);
	LUT2 #(
		.INIT('h4)
	) name1571 (
		_w3705_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h2)
	) name1572 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3694_,
		_w3718_
	);
	LUT2 #(
		.INIT('h4)
	) name1573 (
		_w3717_,
		_w3718_,
		_w3719_
	);
	LUT2 #(
		.INIT('h1)
	) name1574 (
		\u5_dout_reg[17]/P0001 ,
		_w2770_,
		_w3720_
	);
	LUT2 #(
		.INIT('h4)
	) name1575 (
		\u5_rp_reg[0]/P0001 ,
		_w3634_,
		_w3721_
	);
	LUT2 #(
		.INIT('h8)
	) name1576 (
		\u5_mem_reg[2][29]/NET0131 ,
		_w2930_,
		_w3722_
	);
	LUT2 #(
		.INIT('h8)
	) name1577 (
		\u5_mem_reg[3][29]/NET0131 ,
		_w2776_,
		_w3723_
	);
	LUT2 #(
		.INIT('h8)
	) name1578 (
		\u5_mem_reg[1][29]/NET0131 ,
		_w2928_,
		_w3724_
	);
	LUT2 #(
		.INIT('h8)
	) name1579 (
		\u5_mem_reg[0][29]/NET0131 ,
		_w2932_,
		_w3725_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		\u5_rp_reg[0]/P0001 ,
		_w3722_,
		_w3726_
	);
	LUT2 #(
		.INIT('h1)
	) name1581 (
		_w3723_,
		_w3724_,
		_w3727_
	);
	LUT2 #(
		.INIT('h4)
	) name1582 (
		_w3725_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h8)
	) name1583 (
		_w3726_,
		_w3728_,
		_w3729_
	);
	LUT2 #(
		.INIT('h2)
	) name1584 (
		_w2771_,
		_w3721_,
		_w3730_
	);
	LUT2 #(
		.INIT('h4)
	) name1585 (
		_w3729_,
		_w3730_,
		_w3731_
	);
	LUT2 #(
		.INIT('h8)
	) name1586 (
		\u5_mem_reg[2][17]/NET0131 ,
		_w2930_,
		_w3732_
	);
	LUT2 #(
		.INIT('h8)
	) name1587 (
		\u5_mem_reg[3][17]/NET0131 ,
		_w2776_,
		_w3733_
	);
	LUT2 #(
		.INIT('h8)
	) name1588 (
		\u5_mem_reg[1][17]/NET0131 ,
		_w2928_,
		_w3734_
	);
	LUT2 #(
		.INIT('h8)
	) name1589 (
		\u5_mem_reg[0][17]/NET0131 ,
		_w2932_,
		_w3735_
	);
	LUT2 #(
		.INIT('h1)
	) name1590 (
		_w3732_,
		_w3733_,
		_w3736_
	);
	LUT2 #(
		.INIT('h1)
	) name1591 (
		_w3734_,
		_w3735_,
		_w3737_
	);
	LUT2 #(
		.INIT('h8)
	) name1592 (
		_w3736_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h2)
	) name1593 (
		_w2937_,
		_w3738_,
		_w3739_
	);
	LUT2 #(
		.INIT('h2)
	) name1594 (
		_w3536_,
		_w3686_,
		_w3740_
	);
	LUT2 #(
		.INIT('h2)
	) name1595 (
		_w2770_,
		_w3739_,
		_w3741_
	);
	LUT2 #(
		.INIT('h4)
	) name1596 (
		_w3740_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h4)
	) name1597 (
		_w3731_,
		_w3742_,
		_w3743_
	);
	LUT2 #(
		.INIT('h2)
	) name1598 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3720_,
		_w3744_
	);
	LUT2 #(
		.INIT('h4)
	) name1599 (
		_w3743_,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('h1)
	) name1600 (
		\u5_dout_reg[18]/P0001 ,
		_w2770_,
		_w3746_
	);
	LUT2 #(
		.INIT('h4)
	) name1601 (
		\u5_rp_reg[0]/P0001 ,
		_w3660_,
		_w3747_
	);
	LUT2 #(
		.INIT('h8)
	) name1602 (
		\u5_mem_reg[2][30]/NET0131 ,
		_w2930_,
		_w3748_
	);
	LUT2 #(
		.INIT('h8)
	) name1603 (
		\u5_mem_reg[3][30]/NET0131 ,
		_w2776_,
		_w3749_
	);
	LUT2 #(
		.INIT('h8)
	) name1604 (
		\u5_mem_reg[1][30]/NET0131 ,
		_w2928_,
		_w3750_
	);
	LUT2 #(
		.INIT('h8)
	) name1605 (
		\u5_mem_reg[0][30]/NET0131 ,
		_w2932_,
		_w3751_
	);
	LUT2 #(
		.INIT('h2)
	) name1606 (
		\u5_rp_reg[0]/P0001 ,
		_w3748_,
		_w3752_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w3749_,
		_w3750_,
		_w3753_
	);
	LUT2 #(
		.INIT('h4)
	) name1608 (
		_w3751_,
		_w3753_,
		_w3754_
	);
	LUT2 #(
		.INIT('h8)
	) name1609 (
		_w3752_,
		_w3754_,
		_w3755_
	);
	LUT2 #(
		.INIT('h2)
	) name1610 (
		_w2771_,
		_w3747_,
		_w3756_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		_w3755_,
		_w3756_,
		_w3757_
	);
	LUT2 #(
		.INIT('h8)
	) name1612 (
		\u5_mem_reg[1][18]/NET0131 ,
		_w2928_,
		_w3758_
	);
	LUT2 #(
		.INIT('h8)
	) name1613 (
		\u5_mem_reg[2][18]/NET0131 ,
		_w2930_,
		_w3759_
	);
	LUT2 #(
		.INIT('h8)
	) name1614 (
		\u5_mem_reg[3][18]/NET0131 ,
		_w2776_,
		_w3760_
	);
	LUT2 #(
		.INIT('h8)
	) name1615 (
		\u5_mem_reg[0][18]/NET0131 ,
		_w2932_,
		_w3761_
	);
	LUT2 #(
		.INIT('h1)
	) name1616 (
		_w3758_,
		_w3759_,
		_w3762_
	);
	LUT2 #(
		.INIT('h1)
	) name1617 (
		_w3760_,
		_w3761_,
		_w3763_
	);
	LUT2 #(
		.INIT('h8)
	) name1618 (
		_w3762_,
		_w3763_,
		_w3764_
	);
	LUT2 #(
		.INIT('h2)
	) name1619 (
		_w2937_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h2)
	) name1620 (
		_w3536_,
		_w3712_,
		_w3766_
	);
	LUT2 #(
		.INIT('h2)
	) name1621 (
		_w2770_,
		_w3765_,
		_w3767_
	);
	LUT2 #(
		.INIT('h4)
	) name1622 (
		_w3766_,
		_w3767_,
		_w3768_
	);
	LUT2 #(
		.INIT('h4)
	) name1623 (
		_w3757_,
		_w3768_,
		_w3769_
	);
	LUT2 #(
		.INIT('h2)
	) name1624 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3746_,
		_w3770_
	);
	LUT2 #(
		.INIT('h4)
	) name1625 (
		_w3769_,
		_w3770_,
		_w3771_
	);
	LUT2 #(
		.INIT('h1)
	) name1626 (
		\u5_dout_reg[19]/P0001 ,
		_w2770_,
		_w3772_
	);
	LUT2 #(
		.INIT('h4)
	) name1627 (
		\u5_rp_reg[0]/P0001 ,
		_w3686_,
		_w3773_
	);
	LUT2 #(
		.INIT('h8)
	) name1628 (
		\u5_mem_reg[2][31]/NET0131 ,
		_w2930_,
		_w3774_
	);
	LUT2 #(
		.INIT('h8)
	) name1629 (
		\u5_mem_reg[3][31]/NET0131 ,
		_w2776_,
		_w3775_
	);
	LUT2 #(
		.INIT('h8)
	) name1630 (
		\u5_mem_reg[1][31]/NET0131 ,
		_w2928_,
		_w3776_
	);
	LUT2 #(
		.INIT('h8)
	) name1631 (
		\u5_mem_reg[0][31]/NET0131 ,
		_w2932_,
		_w3777_
	);
	LUT2 #(
		.INIT('h2)
	) name1632 (
		\u5_rp_reg[0]/P0001 ,
		_w3774_,
		_w3778_
	);
	LUT2 #(
		.INIT('h1)
	) name1633 (
		_w3775_,
		_w3776_,
		_w3779_
	);
	LUT2 #(
		.INIT('h4)
	) name1634 (
		_w3777_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('h8)
	) name1635 (
		_w3778_,
		_w3780_,
		_w3781_
	);
	LUT2 #(
		.INIT('h2)
	) name1636 (
		_w2771_,
		_w3773_,
		_w3782_
	);
	LUT2 #(
		.INIT('h4)
	) name1637 (
		_w3781_,
		_w3782_,
		_w3783_
	);
	LUT2 #(
		.INIT('h8)
	) name1638 (
		\u5_mem_reg[2][19]/NET0131 ,
		_w2930_,
		_w3784_
	);
	LUT2 #(
		.INIT('h8)
	) name1639 (
		\u5_mem_reg[3][19]/NET0131 ,
		_w2776_,
		_w3785_
	);
	LUT2 #(
		.INIT('h8)
	) name1640 (
		\u5_mem_reg[1][19]/NET0131 ,
		_w2928_,
		_w3786_
	);
	LUT2 #(
		.INIT('h8)
	) name1641 (
		\u5_mem_reg[0][19]/NET0131 ,
		_w2932_,
		_w3787_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		_w3784_,
		_w3785_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name1643 (
		_w3786_,
		_w3787_,
		_w3789_
	);
	LUT2 #(
		.INIT('h8)
	) name1644 (
		_w3788_,
		_w3789_,
		_w3790_
	);
	LUT2 #(
		.INIT('h2)
	) name1645 (
		_w2937_,
		_w3790_,
		_w3791_
	);
	LUT2 #(
		.INIT('h2)
	) name1646 (
		_w3536_,
		_w3738_,
		_w3792_
	);
	LUT2 #(
		.INIT('h2)
	) name1647 (
		_w2770_,
		_w3791_,
		_w3793_
	);
	LUT2 #(
		.INIT('h4)
	) name1648 (
		_w3792_,
		_w3793_,
		_w3794_
	);
	LUT2 #(
		.INIT('h4)
	) name1649 (
		_w3783_,
		_w3794_,
		_w3795_
	);
	LUT2 #(
		.INIT('h2)
	) name1650 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3772_,
		_w3796_
	);
	LUT2 #(
		.INIT('h4)
	) name1651 (
		_w3795_,
		_w3796_,
		_w3797_
	);
	LUT2 #(
		.INIT('h1)
	) name1652 (
		\u5_dout_reg[2]/P0001 ,
		_w2770_,
		_w3798_
	);
	LUT2 #(
		.INIT('h4)
	) name1653 (
		_w2936_,
		_w3536_,
		_w3799_
	);
	LUT2 #(
		.INIT('h8)
	) name1654 (
		\u5_mem_reg[1][2]/NET0131 ,
		_w2928_,
		_w3800_
	);
	LUT2 #(
		.INIT('h8)
	) name1655 (
		\u5_mem_reg[0][2]/NET0131 ,
		_w2932_,
		_w3801_
	);
	LUT2 #(
		.INIT('h8)
	) name1656 (
		\u5_mem_reg[2][2]/NET0131 ,
		_w2930_,
		_w3802_
	);
	LUT2 #(
		.INIT('h8)
	) name1657 (
		\u5_mem_reg[3][2]/NET0131 ,
		_w2776_,
		_w3803_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		_w3800_,
		_w3801_,
		_w3804_
	);
	LUT2 #(
		.INIT('h1)
	) name1659 (
		_w3802_,
		_w3803_,
		_w3805_
	);
	LUT2 #(
		.INIT('h8)
	) name1660 (
		_w3804_,
		_w3805_,
		_w3806_
	);
	LUT2 #(
		.INIT('h2)
	) name1661 (
		_w2937_,
		_w3806_,
		_w3807_
	);
	LUT2 #(
		.INIT('h2)
	) name1662 (
		_w2770_,
		_w3799_,
		_w3808_
	);
	LUT2 #(
		.INIT('h4)
	) name1663 (
		_w3807_,
		_w3808_,
		_w3809_
	);
	LUT2 #(
		.INIT('h2)
	) name1664 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3798_,
		_w3810_
	);
	LUT2 #(
		.INIT('h4)
	) name1665 (
		_w3809_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h1)
	) name1666 (
		\u5_dout_reg[3]/P0001 ,
		_w2770_,
		_w3812_
	);
	LUT2 #(
		.INIT('h4)
	) name1667 (
		_w2949_,
		_w3536_,
		_w3813_
	);
	LUT2 #(
		.INIT('h8)
	) name1668 (
		\u5_mem_reg[3][3]/NET0131 ,
		_w2776_,
		_w3814_
	);
	LUT2 #(
		.INIT('h8)
	) name1669 (
		\u5_mem_reg[2][3]/NET0131 ,
		_w2930_,
		_w3815_
	);
	LUT2 #(
		.INIT('h8)
	) name1670 (
		\u5_mem_reg[1][3]/NET0131 ,
		_w2928_,
		_w3816_
	);
	LUT2 #(
		.INIT('h8)
	) name1671 (
		\u5_mem_reg[0][3]/NET0131 ,
		_w2932_,
		_w3817_
	);
	LUT2 #(
		.INIT('h1)
	) name1672 (
		_w3814_,
		_w3815_,
		_w3818_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		_w3816_,
		_w3817_,
		_w3819_
	);
	LUT2 #(
		.INIT('h8)
	) name1674 (
		_w3818_,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h2)
	) name1675 (
		_w2937_,
		_w3820_,
		_w3821_
	);
	LUT2 #(
		.INIT('h2)
	) name1676 (
		_w2770_,
		_w3813_,
		_w3822_
	);
	LUT2 #(
		.INIT('h4)
	) name1677 (
		_w3821_,
		_w3822_,
		_w3823_
	);
	LUT2 #(
		.INIT('h2)
	) name1678 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3812_,
		_w3824_
	);
	LUT2 #(
		.INIT('h4)
	) name1679 (
		_w3823_,
		_w3824_,
		_w3825_
	);
	LUT2 #(
		.INIT('h1)
	) name1680 (
		\u5_dout_reg[4]/P0001 ,
		_w2770_,
		_w3826_
	);
	LUT2 #(
		.INIT('h4)
	) name1681 (
		\u5_rp_reg[0]/P0001 ,
		_w2936_,
		_w3827_
	);
	LUT2 #(
		.INIT('h8)
	) name1682 (
		\u5_rp_reg[0]/P0001 ,
		_w3712_,
		_w3828_
	);
	LUT2 #(
		.INIT('h2)
	) name1683 (
		_w2771_,
		_w3827_,
		_w3829_
	);
	LUT2 #(
		.INIT('h4)
	) name1684 (
		_w3828_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h8)
	) name1685 (
		\u5_mem_reg[3][4]/NET0131 ,
		_w2776_,
		_w3831_
	);
	LUT2 #(
		.INIT('h8)
	) name1686 (
		\u5_mem_reg[1][4]/NET0131 ,
		_w2928_,
		_w3832_
	);
	LUT2 #(
		.INIT('h8)
	) name1687 (
		\u5_mem_reg[2][4]/NET0131 ,
		_w2930_,
		_w3833_
	);
	LUT2 #(
		.INIT('h8)
	) name1688 (
		\u5_mem_reg[0][4]/NET0131 ,
		_w2932_,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		_w3831_,
		_w3832_,
		_w3835_
	);
	LUT2 #(
		.INIT('h1)
	) name1690 (
		_w3833_,
		_w3834_,
		_w3836_
	);
	LUT2 #(
		.INIT('h8)
	) name1691 (
		_w3835_,
		_w3836_,
		_w3837_
	);
	LUT2 #(
		.INIT('h2)
	) name1692 (
		_w2937_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h2)
	) name1693 (
		_w3536_,
		_w3806_,
		_w3839_
	);
	LUT2 #(
		.INIT('h2)
	) name1694 (
		_w2770_,
		_w3838_,
		_w3840_
	);
	LUT2 #(
		.INIT('h4)
	) name1695 (
		_w3839_,
		_w3840_,
		_w3841_
	);
	LUT2 #(
		.INIT('h4)
	) name1696 (
		_w3830_,
		_w3841_,
		_w3842_
	);
	LUT2 #(
		.INIT('h2)
	) name1697 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3826_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name1698 (
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h1)
	) name1699 (
		\u5_dout_reg[5]/P0001 ,
		_w2770_,
		_w3845_
	);
	LUT2 #(
		.INIT('h4)
	) name1700 (
		\u5_rp_reg[0]/P0001 ,
		_w2949_,
		_w3846_
	);
	LUT2 #(
		.INIT('h8)
	) name1701 (
		\u5_rp_reg[0]/P0001 ,
		_w3738_,
		_w3847_
	);
	LUT2 #(
		.INIT('h2)
	) name1702 (
		_w2771_,
		_w3846_,
		_w3848_
	);
	LUT2 #(
		.INIT('h4)
	) name1703 (
		_w3847_,
		_w3848_,
		_w3849_
	);
	LUT2 #(
		.INIT('h8)
	) name1704 (
		\u5_mem_reg[1][5]/NET0131 ,
		_w2928_,
		_w3850_
	);
	LUT2 #(
		.INIT('h8)
	) name1705 (
		\u5_mem_reg[2][5]/NET0131 ,
		_w2930_,
		_w3851_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		\u5_mem_reg[3][5]/NET0131 ,
		_w2776_,
		_w3852_
	);
	LUT2 #(
		.INIT('h8)
	) name1707 (
		\u5_mem_reg[0][5]/NET0131 ,
		_w2932_,
		_w3853_
	);
	LUT2 #(
		.INIT('h1)
	) name1708 (
		_w3850_,
		_w3851_,
		_w3854_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w3852_,
		_w3853_,
		_w3855_
	);
	LUT2 #(
		.INIT('h8)
	) name1710 (
		_w3854_,
		_w3855_,
		_w3856_
	);
	LUT2 #(
		.INIT('h2)
	) name1711 (
		_w2937_,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('h2)
	) name1712 (
		_w3536_,
		_w3820_,
		_w3858_
	);
	LUT2 #(
		.INIT('h2)
	) name1713 (
		_w2770_,
		_w3857_,
		_w3859_
	);
	LUT2 #(
		.INIT('h4)
	) name1714 (
		_w3858_,
		_w3859_,
		_w3860_
	);
	LUT2 #(
		.INIT('h4)
	) name1715 (
		_w3849_,
		_w3860_,
		_w3861_
	);
	LUT2 #(
		.INIT('h2)
	) name1716 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3845_,
		_w3862_
	);
	LUT2 #(
		.INIT('h4)
	) name1717 (
		_w3861_,
		_w3862_,
		_w3863_
	);
	LUT2 #(
		.INIT('h1)
	) name1718 (
		\u5_dout_reg[6]/P0001 ,
		_w2770_,
		_w3864_
	);
	LUT2 #(
		.INIT('h4)
	) name1719 (
		\u5_rp_reg[0]/P0001 ,
		_w3806_,
		_w3865_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		\u5_rp_reg[0]/P0001 ,
		_w3764_,
		_w3866_
	);
	LUT2 #(
		.INIT('h2)
	) name1721 (
		_w2771_,
		_w3865_,
		_w3867_
	);
	LUT2 #(
		.INIT('h4)
	) name1722 (
		_w3866_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h2)
	) name1723 (
		_w2937_,
		_w3516_,
		_w3869_
	);
	LUT2 #(
		.INIT('h2)
	) name1724 (
		_w3536_,
		_w3837_,
		_w3870_
	);
	LUT2 #(
		.INIT('h2)
	) name1725 (
		_w2770_,
		_w3869_,
		_w3871_
	);
	LUT2 #(
		.INIT('h4)
	) name1726 (
		_w3870_,
		_w3871_,
		_w3872_
	);
	LUT2 #(
		.INIT('h4)
	) name1727 (
		_w3868_,
		_w3872_,
		_w3873_
	);
	LUT2 #(
		.INIT('h2)
	) name1728 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3864_,
		_w3874_
	);
	LUT2 #(
		.INIT('h4)
	) name1729 (
		_w3873_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h1)
	) name1730 (
		\u5_dout_reg[7]/P0001 ,
		_w2770_,
		_w3876_
	);
	LUT2 #(
		.INIT('h4)
	) name1731 (
		\u5_rp_reg[0]/P0001 ,
		_w3820_,
		_w3877_
	);
	LUT2 #(
		.INIT('h8)
	) name1732 (
		\u5_rp_reg[0]/P0001 ,
		_w3790_,
		_w3878_
	);
	LUT2 #(
		.INIT('h2)
	) name1733 (
		_w2771_,
		_w3877_,
		_w3879_
	);
	LUT2 #(
		.INIT('h4)
	) name1734 (
		_w3878_,
		_w3879_,
		_w3880_
	);
	LUT2 #(
		.INIT('h2)
	) name1735 (
		_w2937_,
		_w3557_,
		_w3881_
	);
	LUT2 #(
		.INIT('h2)
	) name1736 (
		_w3536_,
		_w3856_,
		_w3882_
	);
	LUT2 #(
		.INIT('h2)
	) name1737 (
		_w2770_,
		_w3881_,
		_w3883_
	);
	LUT2 #(
		.INIT('h4)
	) name1738 (
		_w3882_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('h4)
	) name1739 (
		_w3880_,
		_w3884_,
		_w3885_
	);
	LUT2 #(
		.INIT('h2)
	) name1740 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3876_,
		_w3886_
	);
	LUT2 #(
		.INIT('h4)
	) name1741 (
		_w3885_,
		_w3886_,
		_w3887_
	);
	LUT2 #(
		.INIT('h1)
	) name1742 (
		\u5_dout_reg[8]/P0001 ,
		_w2770_,
		_w3888_
	);
	LUT2 #(
		.INIT('h4)
	) name1743 (
		\u5_rp_reg[0]/P0001 ,
		_w3837_,
		_w3889_
	);
	LUT2 #(
		.INIT('h8)
	) name1744 (
		\u5_mem_reg[2][20]/NET0131 ,
		_w2930_,
		_w3890_
	);
	LUT2 #(
		.INIT('h8)
	) name1745 (
		\u5_mem_reg[3][20]/NET0131 ,
		_w2776_,
		_w3891_
	);
	LUT2 #(
		.INIT('h8)
	) name1746 (
		\u5_mem_reg[1][20]/NET0131 ,
		_w2928_,
		_w3892_
	);
	LUT2 #(
		.INIT('h8)
	) name1747 (
		\u5_mem_reg[0][20]/NET0131 ,
		_w2932_,
		_w3893_
	);
	LUT2 #(
		.INIT('h2)
	) name1748 (
		\u5_rp_reg[0]/P0001 ,
		_w3890_,
		_w3894_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		_w3891_,
		_w3892_,
		_w3895_
	);
	LUT2 #(
		.INIT('h4)
	) name1750 (
		_w3893_,
		_w3895_,
		_w3896_
	);
	LUT2 #(
		.INIT('h8)
	) name1751 (
		_w3894_,
		_w3896_,
		_w3897_
	);
	LUT2 #(
		.INIT('h2)
	) name1752 (
		_w2771_,
		_w3889_,
		_w3898_
	);
	LUT2 #(
		.INIT('h4)
	) name1753 (
		_w3897_,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h2)
	) name1754 (
		_w2937_,
		_w3543_,
		_w3900_
	);
	LUT2 #(
		.INIT('h4)
	) name1755 (
		_w3516_,
		_w3536_,
		_w3901_
	);
	LUT2 #(
		.INIT('h2)
	) name1756 (
		_w2770_,
		_w3900_,
		_w3902_
	);
	LUT2 #(
		.INIT('h4)
	) name1757 (
		_w3901_,
		_w3902_,
		_w3903_
	);
	LUT2 #(
		.INIT('h4)
	) name1758 (
		_w3899_,
		_w3903_,
		_w3904_
	);
	LUT2 #(
		.INIT('h2)
	) name1759 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3888_,
		_w3905_
	);
	LUT2 #(
		.INIT('h4)
	) name1760 (
		_w3904_,
		_w3905_,
		_w3906_
	);
	LUT2 #(
		.INIT('h1)
	) name1761 (
		\u5_dout_reg[9]/P0001 ,
		_w2770_,
		_w3907_
	);
	LUT2 #(
		.INIT('h4)
	) name1762 (
		\u5_rp_reg[0]/P0001 ,
		_w3856_,
		_w3908_
	);
	LUT2 #(
		.INIT('h8)
	) name1763 (
		\u5_mem_reg[2][21]/NET0131 ,
		_w2930_,
		_w3909_
	);
	LUT2 #(
		.INIT('h8)
	) name1764 (
		\u5_mem_reg[3][21]/NET0131 ,
		_w2776_,
		_w3910_
	);
	LUT2 #(
		.INIT('h8)
	) name1765 (
		\u5_mem_reg[1][21]/NET0131 ,
		_w2928_,
		_w3911_
	);
	LUT2 #(
		.INIT('h8)
	) name1766 (
		\u5_mem_reg[0][21]/NET0131 ,
		_w2932_,
		_w3912_
	);
	LUT2 #(
		.INIT('h2)
	) name1767 (
		\u5_rp_reg[0]/P0001 ,
		_w3909_,
		_w3913_
	);
	LUT2 #(
		.INIT('h1)
	) name1768 (
		_w3910_,
		_w3911_,
		_w3914_
	);
	LUT2 #(
		.INIT('h4)
	) name1769 (
		_w3912_,
		_w3914_,
		_w3915_
	);
	LUT2 #(
		.INIT('h8)
	) name1770 (
		_w3913_,
		_w3915_,
		_w3916_
	);
	LUT2 #(
		.INIT('h2)
	) name1771 (
		_w2771_,
		_w3908_,
		_w3917_
	);
	LUT2 #(
		.INIT('h4)
	) name1772 (
		_w3916_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h2)
	) name1773 (
		_w2937_,
		_w3583_,
		_w3919_
	);
	LUT2 #(
		.INIT('h2)
	) name1774 (
		_w3536_,
		_w3557_,
		_w3920_
	);
	LUT2 #(
		.INIT('h2)
	) name1775 (
		_w2770_,
		_w3919_,
		_w3921_
	);
	LUT2 #(
		.INIT('h4)
	) name1776 (
		_w3920_,
		_w3921_,
		_w3922_
	);
	LUT2 #(
		.INIT('h4)
	) name1777 (
		_w3918_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h2)
	) name1778 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w3907_,
		_w3924_
	);
	LUT2 #(
		.INIT('h4)
	) name1779 (
		_w3923_,
		_w3924_,
		_w3925_
	);
	LUT2 #(
		.INIT('h1)
	) name1780 (
		\u6_dout_reg[10]/P0001 ,
		_w2795_,
		_w3926_
	);
	LUT2 #(
		.INIT('h8)
	) name1781 (
		\u6_mem_reg[3][6]/NET0131 ,
		_w2801_,
		_w3927_
	);
	LUT2 #(
		.INIT('h8)
	) name1782 (
		\u6_mem_reg[2][6]/NET0131 ,
		_w2955_,
		_w3928_
	);
	LUT2 #(
		.INIT('h8)
	) name1783 (
		\u6_mem_reg[0][6]/NET0131 ,
		_w2959_,
		_w3929_
	);
	LUT2 #(
		.INIT('h8)
	) name1784 (
		\u6_mem_reg[1][6]/NET0131 ,
		_w2957_,
		_w3930_
	);
	LUT2 #(
		.INIT('h1)
	) name1785 (
		_w3927_,
		_w3928_,
		_w3931_
	);
	LUT2 #(
		.INIT('h1)
	) name1786 (
		_w3929_,
		_w3930_,
		_w3932_
	);
	LUT2 #(
		.INIT('h8)
	) name1787 (
		_w3931_,
		_w3932_,
		_w3933_
	);
	LUT2 #(
		.INIT('h4)
	) name1788 (
		\u6_rp_reg[0]/P0001 ,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h8)
	) name1789 (
		\u6_mem_reg[2][22]/NET0131 ,
		_w2955_,
		_w3935_
	);
	LUT2 #(
		.INIT('h8)
	) name1790 (
		\u6_mem_reg[1][22]/NET0131 ,
		_w2957_,
		_w3936_
	);
	LUT2 #(
		.INIT('h8)
	) name1791 (
		\u6_mem_reg[3][22]/NET0131 ,
		_w2801_,
		_w3937_
	);
	LUT2 #(
		.INIT('h8)
	) name1792 (
		\u6_mem_reg[0][22]/NET0131 ,
		_w2959_,
		_w3938_
	);
	LUT2 #(
		.INIT('h2)
	) name1793 (
		\u6_rp_reg[0]/P0001 ,
		_w3935_,
		_w3939_
	);
	LUT2 #(
		.INIT('h1)
	) name1794 (
		_w3936_,
		_w3937_,
		_w3940_
	);
	LUT2 #(
		.INIT('h4)
	) name1795 (
		_w3938_,
		_w3940_,
		_w3941_
	);
	LUT2 #(
		.INIT('h8)
	) name1796 (
		_w3939_,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h2)
	) name1797 (
		_w2796_,
		_w3934_,
		_w3943_
	);
	LUT2 #(
		.INIT('h4)
	) name1798 (
		_w3942_,
		_w3943_,
		_w3944_
	);
	LUT2 #(
		.INIT('h8)
	) name1799 (
		\u6_mem_reg[1][10]/NET0131 ,
		_w2957_,
		_w3945_
	);
	LUT2 #(
		.INIT('h8)
	) name1800 (
		\u6_mem_reg[3][10]/NET0131 ,
		_w2801_,
		_w3946_
	);
	LUT2 #(
		.INIT('h8)
	) name1801 (
		\u6_mem_reg[0][10]/NET0131 ,
		_w2959_,
		_w3947_
	);
	LUT2 #(
		.INIT('h8)
	) name1802 (
		\u6_mem_reg[2][10]/NET0131 ,
		_w2955_,
		_w3948_
	);
	LUT2 #(
		.INIT('h1)
	) name1803 (
		_w3945_,
		_w3946_,
		_w3949_
	);
	LUT2 #(
		.INIT('h1)
	) name1804 (
		_w3947_,
		_w3948_,
		_w3950_
	);
	LUT2 #(
		.INIT('h8)
	) name1805 (
		_w3949_,
		_w3950_,
		_w3951_
	);
	LUT2 #(
		.INIT('h2)
	) name1806 (
		_w2964_,
		_w3951_,
		_w3952_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		\u13_occ0_r_reg[26]/NET0131 ,
		\u13_occ0_r_reg[27]/NET0131 ,
		_w3953_
	);
	LUT2 #(
		.INIT('h8)
	) name1808 (
		\u6_mem_reg[3][8]/NET0131 ,
		_w2801_,
		_w3954_
	);
	LUT2 #(
		.INIT('h8)
	) name1809 (
		\u6_mem_reg[2][8]/NET0131 ,
		_w2955_,
		_w3955_
	);
	LUT2 #(
		.INIT('h8)
	) name1810 (
		\u6_mem_reg[0][8]/NET0131 ,
		_w2959_,
		_w3956_
	);
	LUT2 #(
		.INIT('h8)
	) name1811 (
		\u6_mem_reg[1][8]/NET0131 ,
		_w2957_,
		_w3957_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w3954_,
		_w3955_,
		_w3958_
	);
	LUT2 #(
		.INIT('h1)
	) name1813 (
		_w3956_,
		_w3957_,
		_w3959_
	);
	LUT2 #(
		.INIT('h8)
	) name1814 (
		_w3958_,
		_w3959_,
		_w3960_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		_w3953_,
		_w3960_,
		_w3961_
	);
	LUT2 #(
		.INIT('h2)
	) name1816 (
		_w2795_,
		_w3952_,
		_w3962_
	);
	LUT2 #(
		.INIT('h4)
	) name1817 (
		_w3961_,
		_w3962_,
		_w3963_
	);
	LUT2 #(
		.INIT('h4)
	) name1818 (
		_w3944_,
		_w3963_,
		_w3964_
	);
	LUT2 #(
		.INIT('h2)
	) name1819 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3926_,
		_w3965_
	);
	LUT2 #(
		.INIT('h4)
	) name1820 (
		_w3964_,
		_w3965_,
		_w3966_
	);
	LUT2 #(
		.INIT('h1)
	) name1821 (
		\u6_dout_reg[11]/P0001 ,
		_w2795_,
		_w3967_
	);
	LUT2 #(
		.INIT('h8)
	) name1822 (
		\u6_mem_reg[3][7]/NET0131 ,
		_w2801_,
		_w3968_
	);
	LUT2 #(
		.INIT('h8)
	) name1823 (
		\u6_mem_reg[2][7]/NET0131 ,
		_w2955_,
		_w3969_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		\u6_mem_reg[0][7]/NET0131 ,
		_w2959_,
		_w3970_
	);
	LUT2 #(
		.INIT('h8)
	) name1825 (
		\u6_mem_reg[1][7]/NET0131 ,
		_w2957_,
		_w3971_
	);
	LUT2 #(
		.INIT('h1)
	) name1826 (
		_w3968_,
		_w3969_,
		_w3972_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w3970_,
		_w3971_,
		_w3973_
	);
	LUT2 #(
		.INIT('h8)
	) name1828 (
		_w3972_,
		_w3973_,
		_w3974_
	);
	LUT2 #(
		.INIT('h4)
	) name1829 (
		\u6_rp_reg[0]/P0001 ,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('h8)
	) name1830 (
		\u6_mem_reg[2][23]/NET0131 ,
		_w2955_,
		_w3976_
	);
	LUT2 #(
		.INIT('h8)
	) name1831 (
		\u6_mem_reg[1][23]/NET0131 ,
		_w2957_,
		_w3977_
	);
	LUT2 #(
		.INIT('h8)
	) name1832 (
		\u6_mem_reg[3][23]/NET0131 ,
		_w2801_,
		_w3978_
	);
	LUT2 #(
		.INIT('h8)
	) name1833 (
		\u6_mem_reg[0][23]/NET0131 ,
		_w2959_,
		_w3979_
	);
	LUT2 #(
		.INIT('h2)
	) name1834 (
		\u6_rp_reg[0]/P0001 ,
		_w3976_,
		_w3980_
	);
	LUT2 #(
		.INIT('h1)
	) name1835 (
		_w3977_,
		_w3978_,
		_w3981_
	);
	LUT2 #(
		.INIT('h4)
	) name1836 (
		_w3979_,
		_w3981_,
		_w3982_
	);
	LUT2 #(
		.INIT('h8)
	) name1837 (
		_w3980_,
		_w3982_,
		_w3983_
	);
	LUT2 #(
		.INIT('h2)
	) name1838 (
		_w2796_,
		_w3975_,
		_w3984_
	);
	LUT2 #(
		.INIT('h4)
	) name1839 (
		_w3983_,
		_w3984_,
		_w3985_
	);
	LUT2 #(
		.INIT('h8)
	) name1840 (
		\u6_mem_reg[3][11]/NET0131 ,
		_w2801_,
		_w3986_
	);
	LUT2 #(
		.INIT('h8)
	) name1841 (
		\u6_mem_reg[2][11]/NET0131 ,
		_w2955_,
		_w3987_
	);
	LUT2 #(
		.INIT('h8)
	) name1842 (
		\u6_mem_reg[0][11]/NET0131 ,
		_w2959_,
		_w3988_
	);
	LUT2 #(
		.INIT('h8)
	) name1843 (
		\u6_mem_reg[1][11]/NET0131 ,
		_w2957_,
		_w3989_
	);
	LUT2 #(
		.INIT('h1)
	) name1844 (
		_w3986_,
		_w3987_,
		_w3990_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		_w3988_,
		_w3989_,
		_w3991_
	);
	LUT2 #(
		.INIT('h8)
	) name1846 (
		_w3990_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h2)
	) name1847 (
		_w2964_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h8)
	) name1848 (
		\u6_mem_reg[3][9]/NET0131 ,
		_w2801_,
		_w3994_
	);
	LUT2 #(
		.INIT('h8)
	) name1849 (
		\u6_mem_reg[1][9]/NET0131 ,
		_w2957_,
		_w3995_
	);
	LUT2 #(
		.INIT('h8)
	) name1850 (
		\u6_mem_reg[2][9]/NET0131 ,
		_w2955_,
		_w3996_
	);
	LUT2 #(
		.INIT('h8)
	) name1851 (
		\u6_mem_reg[0][9]/NET0131 ,
		_w2959_,
		_w3997_
	);
	LUT2 #(
		.INIT('h1)
	) name1852 (
		_w3994_,
		_w3995_,
		_w3998_
	);
	LUT2 #(
		.INIT('h1)
	) name1853 (
		_w3996_,
		_w3997_,
		_w3999_
	);
	LUT2 #(
		.INIT('h8)
	) name1854 (
		_w3998_,
		_w3999_,
		_w4000_
	);
	LUT2 #(
		.INIT('h2)
	) name1855 (
		_w3953_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('h2)
	) name1856 (
		_w2795_,
		_w3993_,
		_w4002_
	);
	LUT2 #(
		.INIT('h4)
	) name1857 (
		_w4001_,
		_w4002_,
		_w4003_
	);
	LUT2 #(
		.INIT('h4)
	) name1858 (
		_w3985_,
		_w4003_,
		_w4004_
	);
	LUT2 #(
		.INIT('h2)
	) name1859 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w3967_,
		_w4005_
	);
	LUT2 #(
		.INIT('h4)
	) name1860 (
		_w4004_,
		_w4005_,
		_w4006_
	);
	LUT2 #(
		.INIT('h1)
	) name1861 (
		\u6_dout_reg[12]/P0001 ,
		_w2795_,
		_w4007_
	);
	LUT2 #(
		.INIT('h4)
	) name1862 (
		\u6_rp_reg[0]/P0001 ,
		_w3960_,
		_w4008_
	);
	LUT2 #(
		.INIT('h8)
	) name1863 (
		\u6_mem_reg[2][24]/NET0131 ,
		_w2955_,
		_w4009_
	);
	LUT2 #(
		.INIT('h8)
	) name1864 (
		\u6_mem_reg[1][24]/NET0131 ,
		_w2957_,
		_w4010_
	);
	LUT2 #(
		.INIT('h8)
	) name1865 (
		\u6_mem_reg[3][24]/NET0131 ,
		_w2801_,
		_w4011_
	);
	LUT2 #(
		.INIT('h8)
	) name1866 (
		\u6_mem_reg[0][24]/NET0131 ,
		_w2959_,
		_w4012_
	);
	LUT2 #(
		.INIT('h2)
	) name1867 (
		\u6_rp_reg[0]/P0001 ,
		_w4009_,
		_w4013_
	);
	LUT2 #(
		.INIT('h1)
	) name1868 (
		_w4010_,
		_w4011_,
		_w4014_
	);
	LUT2 #(
		.INIT('h4)
	) name1869 (
		_w4012_,
		_w4014_,
		_w4015_
	);
	LUT2 #(
		.INIT('h8)
	) name1870 (
		_w4013_,
		_w4015_,
		_w4016_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		_w2796_,
		_w4008_,
		_w4017_
	);
	LUT2 #(
		.INIT('h4)
	) name1872 (
		_w4016_,
		_w4017_,
		_w4018_
	);
	LUT2 #(
		.INIT('h8)
	) name1873 (
		\u6_mem_reg[3][12]/NET0131 ,
		_w2801_,
		_w4019_
	);
	LUT2 #(
		.INIT('h8)
	) name1874 (
		\u6_mem_reg[1][12]/NET0131 ,
		_w2957_,
		_w4020_
	);
	LUT2 #(
		.INIT('h8)
	) name1875 (
		\u6_mem_reg[0][12]/NET0131 ,
		_w2959_,
		_w4021_
	);
	LUT2 #(
		.INIT('h8)
	) name1876 (
		\u6_mem_reg[2][12]/NET0131 ,
		_w2955_,
		_w4022_
	);
	LUT2 #(
		.INIT('h1)
	) name1877 (
		_w4019_,
		_w4020_,
		_w4023_
	);
	LUT2 #(
		.INIT('h1)
	) name1878 (
		_w4021_,
		_w4022_,
		_w4024_
	);
	LUT2 #(
		.INIT('h8)
	) name1879 (
		_w4023_,
		_w4024_,
		_w4025_
	);
	LUT2 #(
		.INIT('h2)
	) name1880 (
		_w2964_,
		_w4025_,
		_w4026_
	);
	LUT2 #(
		.INIT('h4)
	) name1881 (
		_w3951_,
		_w3953_,
		_w4027_
	);
	LUT2 #(
		.INIT('h2)
	) name1882 (
		_w2795_,
		_w4026_,
		_w4028_
	);
	LUT2 #(
		.INIT('h4)
	) name1883 (
		_w4027_,
		_w4028_,
		_w4029_
	);
	LUT2 #(
		.INIT('h4)
	) name1884 (
		_w4018_,
		_w4029_,
		_w4030_
	);
	LUT2 #(
		.INIT('h2)
	) name1885 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4007_,
		_w4031_
	);
	LUT2 #(
		.INIT('h4)
	) name1886 (
		_w4030_,
		_w4031_,
		_w4032_
	);
	LUT2 #(
		.INIT('h1)
	) name1887 (
		\u6_dout_reg[13]/P0001 ,
		_w2795_,
		_w4033_
	);
	LUT2 #(
		.INIT('h4)
	) name1888 (
		\u6_rp_reg[0]/P0001 ,
		_w4000_,
		_w4034_
	);
	LUT2 #(
		.INIT('h8)
	) name1889 (
		\u6_mem_reg[2][25]/NET0131 ,
		_w2955_,
		_w4035_
	);
	LUT2 #(
		.INIT('h8)
	) name1890 (
		\u6_mem_reg[1][25]/NET0131 ,
		_w2957_,
		_w4036_
	);
	LUT2 #(
		.INIT('h8)
	) name1891 (
		\u6_mem_reg[3][25]/NET0131 ,
		_w2801_,
		_w4037_
	);
	LUT2 #(
		.INIT('h8)
	) name1892 (
		\u6_mem_reg[0][25]/NET0131 ,
		_w2959_,
		_w4038_
	);
	LUT2 #(
		.INIT('h2)
	) name1893 (
		\u6_rp_reg[0]/P0001 ,
		_w4035_,
		_w4039_
	);
	LUT2 #(
		.INIT('h1)
	) name1894 (
		_w4036_,
		_w4037_,
		_w4040_
	);
	LUT2 #(
		.INIT('h4)
	) name1895 (
		_w4038_,
		_w4040_,
		_w4041_
	);
	LUT2 #(
		.INIT('h8)
	) name1896 (
		_w4039_,
		_w4041_,
		_w4042_
	);
	LUT2 #(
		.INIT('h2)
	) name1897 (
		_w2796_,
		_w4034_,
		_w4043_
	);
	LUT2 #(
		.INIT('h4)
	) name1898 (
		_w4042_,
		_w4043_,
		_w4044_
	);
	LUT2 #(
		.INIT('h8)
	) name1899 (
		\u6_mem_reg[3][13]/NET0131 ,
		_w2801_,
		_w4045_
	);
	LUT2 #(
		.INIT('h8)
	) name1900 (
		\u6_mem_reg[2][13]/NET0131 ,
		_w2955_,
		_w4046_
	);
	LUT2 #(
		.INIT('h8)
	) name1901 (
		\u6_mem_reg[0][13]/NET0131 ,
		_w2959_,
		_w4047_
	);
	LUT2 #(
		.INIT('h8)
	) name1902 (
		\u6_mem_reg[1][13]/NET0131 ,
		_w2957_,
		_w4048_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		_w4045_,
		_w4046_,
		_w4049_
	);
	LUT2 #(
		.INIT('h1)
	) name1904 (
		_w4047_,
		_w4048_,
		_w4050_
	);
	LUT2 #(
		.INIT('h8)
	) name1905 (
		_w4049_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h2)
	) name1906 (
		_w2964_,
		_w4051_,
		_w4052_
	);
	LUT2 #(
		.INIT('h2)
	) name1907 (
		_w3953_,
		_w3992_,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name1908 (
		_w2795_,
		_w4052_,
		_w4054_
	);
	LUT2 #(
		.INIT('h4)
	) name1909 (
		_w4053_,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('h4)
	) name1910 (
		_w4044_,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h2)
	) name1911 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4033_,
		_w4057_
	);
	LUT2 #(
		.INIT('h4)
	) name1912 (
		_w4056_,
		_w4057_,
		_w4058_
	);
	LUT2 #(
		.INIT('h1)
	) name1913 (
		\u6_dout_reg[14]/P0001 ,
		_w2795_,
		_w4059_
	);
	LUT2 #(
		.INIT('h4)
	) name1914 (
		\u6_rp_reg[0]/P0001 ,
		_w3951_,
		_w4060_
	);
	LUT2 #(
		.INIT('h8)
	) name1915 (
		\u6_mem_reg[2][26]/NET0131 ,
		_w2955_,
		_w4061_
	);
	LUT2 #(
		.INIT('h8)
	) name1916 (
		\u6_mem_reg[1][26]/NET0131 ,
		_w2957_,
		_w4062_
	);
	LUT2 #(
		.INIT('h8)
	) name1917 (
		\u6_mem_reg[3][26]/NET0131 ,
		_w2801_,
		_w4063_
	);
	LUT2 #(
		.INIT('h8)
	) name1918 (
		\u6_mem_reg[0][26]/NET0131 ,
		_w2959_,
		_w4064_
	);
	LUT2 #(
		.INIT('h2)
	) name1919 (
		\u6_rp_reg[0]/P0001 ,
		_w4061_,
		_w4065_
	);
	LUT2 #(
		.INIT('h1)
	) name1920 (
		_w4062_,
		_w4063_,
		_w4066_
	);
	LUT2 #(
		.INIT('h4)
	) name1921 (
		_w4064_,
		_w4066_,
		_w4067_
	);
	LUT2 #(
		.INIT('h8)
	) name1922 (
		_w4065_,
		_w4067_,
		_w4068_
	);
	LUT2 #(
		.INIT('h2)
	) name1923 (
		_w2796_,
		_w4060_,
		_w4069_
	);
	LUT2 #(
		.INIT('h4)
	) name1924 (
		_w4068_,
		_w4069_,
		_w4070_
	);
	LUT2 #(
		.INIT('h8)
	) name1925 (
		\u6_mem_reg[1][14]/NET0131 ,
		_w2957_,
		_w4071_
	);
	LUT2 #(
		.INIT('h8)
	) name1926 (
		\u6_mem_reg[0][14]/NET0131 ,
		_w2959_,
		_w4072_
	);
	LUT2 #(
		.INIT('h8)
	) name1927 (
		\u6_mem_reg[3][14]/NET0131 ,
		_w2801_,
		_w4073_
	);
	LUT2 #(
		.INIT('h8)
	) name1928 (
		\u6_mem_reg[2][14]/NET0131 ,
		_w2955_,
		_w4074_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		_w4071_,
		_w4072_,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name1930 (
		_w4073_,
		_w4074_,
		_w4076_
	);
	LUT2 #(
		.INIT('h8)
	) name1931 (
		_w4075_,
		_w4076_,
		_w4077_
	);
	LUT2 #(
		.INIT('h2)
	) name1932 (
		_w2964_,
		_w4077_,
		_w4078_
	);
	LUT2 #(
		.INIT('h2)
	) name1933 (
		_w3953_,
		_w4025_,
		_w4079_
	);
	LUT2 #(
		.INIT('h2)
	) name1934 (
		_w2795_,
		_w4078_,
		_w4080_
	);
	LUT2 #(
		.INIT('h4)
	) name1935 (
		_w4079_,
		_w4080_,
		_w4081_
	);
	LUT2 #(
		.INIT('h4)
	) name1936 (
		_w4070_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h2)
	) name1937 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4059_,
		_w4083_
	);
	LUT2 #(
		.INIT('h4)
	) name1938 (
		_w4082_,
		_w4083_,
		_w4084_
	);
	LUT2 #(
		.INIT('h1)
	) name1939 (
		\u6_dout_reg[15]/P0001 ,
		_w2795_,
		_w4085_
	);
	LUT2 #(
		.INIT('h4)
	) name1940 (
		\u6_rp_reg[0]/P0001 ,
		_w3992_,
		_w4086_
	);
	LUT2 #(
		.INIT('h8)
	) name1941 (
		\u6_mem_reg[2][27]/NET0131 ,
		_w2955_,
		_w4087_
	);
	LUT2 #(
		.INIT('h8)
	) name1942 (
		\u6_mem_reg[3][27]/NET0131 ,
		_w2801_,
		_w4088_
	);
	LUT2 #(
		.INIT('h8)
	) name1943 (
		\u6_mem_reg[1][27]/NET0131 ,
		_w2957_,
		_w4089_
	);
	LUT2 #(
		.INIT('h8)
	) name1944 (
		\u6_mem_reg[0][27]/NET0131 ,
		_w2959_,
		_w4090_
	);
	LUT2 #(
		.INIT('h2)
	) name1945 (
		\u6_rp_reg[0]/P0001 ,
		_w4087_,
		_w4091_
	);
	LUT2 #(
		.INIT('h1)
	) name1946 (
		_w4088_,
		_w4089_,
		_w4092_
	);
	LUT2 #(
		.INIT('h4)
	) name1947 (
		_w4090_,
		_w4092_,
		_w4093_
	);
	LUT2 #(
		.INIT('h8)
	) name1948 (
		_w4091_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h2)
	) name1949 (
		_w2796_,
		_w4086_,
		_w4095_
	);
	LUT2 #(
		.INIT('h4)
	) name1950 (
		_w4094_,
		_w4095_,
		_w4096_
	);
	LUT2 #(
		.INIT('h8)
	) name1951 (
		\u6_mem_reg[3][15]/NET0131 ,
		_w2801_,
		_w4097_
	);
	LUT2 #(
		.INIT('h8)
	) name1952 (
		\u6_mem_reg[2][15]/NET0131 ,
		_w2955_,
		_w4098_
	);
	LUT2 #(
		.INIT('h8)
	) name1953 (
		\u6_mem_reg[0][15]/NET0131 ,
		_w2959_,
		_w4099_
	);
	LUT2 #(
		.INIT('h8)
	) name1954 (
		\u6_mem_reg[1][15]/NET0131 ,
		_w2957_,
		_w4100_
	);
	LUT2 #(
		.INIT('h1)
	) name1955 (
		_w4097_,
		_w4098_,
		_w4101_
	);
	LUT2 #(
		.INIT('h1)
	) name1956 (
		_w4099_,
		_w4100_,
		_w4102_
	);
	LUT2 #(
		.INIT('h8)
	) name1957 (
		_w4101_,
		_w4102_,
		_w4103_
	);
	LUT2 #(
		.INIT('h2)
	) name1958 (
		_w2964_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h2)
	) name1959 (
		_w3953_,
		_w4051_,
		_w4105_
	);
	LUT2 #(
		.INIT('h2)
	) name1960 (
		_w2795_,
		_w4104_,
		_w4106_
	);
	LUT2 #(
		.INIT('h4)
	) name1961 (
		_w4105_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h4)
	) name1962 (
		_w4096_,
		_w4107_,
		_w4108_
	);
	LUT2 #(
		.INIT('h2)
	) name1963 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4085_,
		_w4109_
	);
	LUT2 #(
		.INIT('h4)
	) name1964 (
		_w4108_,
		_w4109_,
		_w4110_
	);
	LUT2 #(
		.INIT('h1)
	) name1965 (
		\u6_dout_reg[16]/P0001 ,
		_w2795_,
		_w4111_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		\u6_rp_reg[0]/P0001 ,
		_w4025_,
		_w4112_
	);
	LUT2 #(
		.INIT('h8)
	) name1967 (
		\u6_mem_reg[2][28]/NET0131 ,
		_w2955_,
		_w4113_
	);
	LUT2 #(
		.INIT('h8)
	) name1968 (
		\u6_mem_reg[1][28]/NET0131 ,
		_w2957_,
		_w4114_
	);
	LUT2 #(
		.INIT('h8)
	) name1969 (
		\u6_mem_reg[3][28]/NET0131 ,
		_w2801_,
		_w4115_
	);
	LUT2 #(
		.INIT('h8)
	) name1970 (
		\u6_mem_reg[0][28]/NET0131 ,
		_w2959_,
		_w4116_
	);
	LUT2 #(
		.INIT('h2)
	) name1971 (
		\u6_rp_reg[0]/P0001 ,
		_w4113_,
		_w4117_
	);
	LUT2 #(
		.INIT('h1)
	) name1972 (
		_w4114_,
		_w4115_,
		_w4118_
	);
	LUT2 #(
		.INIT('h4)
	) name1973 (
		_w4116_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h8)
	) name1974 (
		_w4117_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h2)
	) name1975 (
		_w2796_,
		_w4112_,
		_w4121_
	);
	LUT2 #(
		.INIT('h4)
	) name1976 (
		_w4120_,
		_w4121_,
		_w4122_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		\u6_mem_reg[1][16]/NET0131 ,
		_w2957_,
		_w4123_
	);
	LUT2 #(
		.INIT('h8)
	) name1978 (
		\u6_mem_reg[0][16]/NET0131 ,
		_w2959_,
		_w4124_
	);
	LUT2 #(
		.INIT('h8)
	) name1979 (
		\u6_mem_reg[2][16]/NET0131 ,
		_w2955_,
		_w4125_
	);
	LUT2 #(
		.INIT('h8)
	) name1980 (
		\u6_mem_reg[3][16]/NET0131 ,
		_w2801_,
		_w4126_
	);
	LUT2 #(
		.INIT('h1)
	) name1981 (
		_w4123_,
		_w4124_,
		_w4127_
	);
	LUT2 #(
		.INIT('h1)
	) name1982 (
		_w4125_,
		_w4126_,
		_w4128_
	);
	LUT2 #(
		.INIT('h8)
	) name1983 (
		_w4127_,
		_w4128_,
		_w4129_
	);
	LUT2 #(
		.INIT('h2)
	) name1984 (
		_w2964_,
		_w4129_,
		_w4130_
	);
	LUT2 #(
		.INIT('h2)
	) name1985 (
		_w3953_,
		_w4077_,
		_w4131_
	);
	LUT2 #(
		.INIT('h2)
	) name1986 (
		_w2795_,
		_w4130_,
		_w4132_
	);
	LUT2 #(
		.INIT('h4)
	) name1987 (
		_w4131_,
		_w4132_,
		_w4133_
	);
	LUT2 #(
		.INIT('h4)
	) name1988 (
		_w4122_,
		_w4133_,
		_w4134_
	);
	LUT2 #(
		.INIT('h2)
	) name1989 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4111_,
		_w4135_
	);
	LUT2 #(
		.INIT('h4)
	) name1990 (
		_w4134_,
		_w4135_,
		_w4136_
	);
	LUT2 #(
		.INIT('h1)
	) name1991 (
		\u6_dout_reg[17]/P0001 ,
		_w2795_,
		_w4137_
	);
	LUT2 #(
		.INIT('h4)
	) name1992 (
		\u6_rp_reg[0]/P0001 ,
		_w4051_,
		_w4138_
	);
	LUT2 #(
		.INIT('h8)
	) name1993 (
		\u6_mem_reg[2][29]/NET0131 ,
		_w2955_,
		_w4139_
	);
	LUT2 #(
		.INIT('h8)
	) name1994 (
		\u6_mem_reg[3][29]/NET0131 ,
		_w2801_,
		_w4140_
	);
	LUT2 #(
		.INIT('h8)
	) name1995 (
		\u6_mem_reg[1][29]/NET0131 ,
		_w2957_,
		_w4141_
	);
	LUT2 #(
		.INIT('h8)
	) name1996 (
		\u6_mem_reg[0][29]/NET0131 ,
		_w2959_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name1997 (
		\u6_rp_reg[0]/P0001 ,
		_w4139_,
		_w4143_
	);
	LUT2 #(
		.INIT('h1)
	) name1998 (
		_w4140_,
		_w4141_,
		_w4144_
	);
	LUT2 #(
		.INIT('h4)
	) name1999 (
		_w4142_,
		_w4144_,
		_w4145_
	);
	LUT2 #(
		.INIT('h8)
	) name2000 (
		_w4143_,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h2)
	) name2001 (
		_w2796_,
		_w4138_,
		_w4147_
	);
	LUT2 #(
		.INIT('h4)
	) name2002 (
		_w4146_,
		_w4147_,
		_w4148_
	);
	LUT2 #(
		.INIT('h8)
	) name2003 (
		\u6_mem_reg[3][17]/NET0131 ,
		_w2801_,
		_w4149_
	);
	LUT2 #(
		.INIT('h8)
	) name2004 (
		\u6_mem_reg[1][17]/NET0131 ,
		_w2957_,
		_w4150_
	);
	LUT2 #(
		.INIT('h8)
	) name2005 (
		\u6_mem_reg[2][17]/NET0131 ,
		_w2955_,
		_w4151_
	);
	LUT2 #(
		.INIT('h8)
	) name2006 (
		\u6_mem_reg[0][17]/NET0131 ,
		_w2959_,
		_w4152_
	);
	LUT2 #(
		.INIT('h1)
	) name2007 (
		_w4149_,
		_w4150_,
		_w4153_
	);
	LUT2 #(
		.INIT('h1)
	) name2008 (
		_w4151_,
		_w4152_,
		_w4154_
	);
	LUT2 #(
		.INIT('h8)
	) name2009 (
		_w4153_,
		_w4154_,
		_w4155_
	);
	LUT2 #(
		.INIT('h2)
	) name2010 (
		_w2964_,
		_w4155_,
		_w4156_
	);
	LUT2 #(
		.INIT('h2)
	) name2011 (
		_w3953_,
		_w4103_,
		_w4157_
	);
	LUT2 #(
		.INIT('h2)
	) name2012 (
		_w2795_,
		_w4156_,
		_w4158_
	);
	LUT2 #(
		.INIT('h4)
	) name2013 (
		_w4157_,
		_w4158_,
		_w4159_
	);
	LUT2 #(
		.INIT('h4)
	) name2014 (
		_w4148_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h2)
	) name2015 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4137_,
		_w4161_
	);
	LUT2 #(
		.INIT('h4)
	) name2016 (
		_w4160_,
		_w4161_,
		_w4162_
	);
	LUT2 #(
		.INIT('h1)
	) name2017 (
		\u6_dout_reg[18]/P0001 ,
		_w2795_,
		_w4163_
	);
	LUT2 #(
		.INIT('h4)
	) name2018 (
		\u6_rp_reg[0]/P0001 ,
		_w4077_,
		_w4164_
	);
	LUT2 #(
		.INIT('h8)
	) name2019 (
		\u6_mem_reg[2][30]/NET0131 ,
		_w2955_,
		_w4165_
	);
	LUT2 #(
		.INIT('h8)
	) name2020 (
		\u6_mem_reg[3][30]/NET0131 ,
		_w2801_,
		_w4166_
	);
	LUT2 #(
		.INIT('h8)
	) name2021 (
		\u6_mem_reg[1][30]/NET0131 ,
		_w2957_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name2022 (
		\u6_mem_reg[0][30]/NET0131 ,
		_w2959_,
		_w4168_
	);
	LUT2 #(
		.INIT('h2)
	) name2023 (
		\u6_rp_reg[0]/P0001 ,
		_w4165_,
		_w4169_
	);
	LUT2 #(
		.INIT('h1)
	) name2024 (
		_w4166_,
		_w4167_,
		_w4170_
	);
	LUT2 #(
		.INIT('h4)
	) name2025 (
		_w4168_,
		_w4170_,
		_w4171_
	);
	LUT2 #(
		.INIT('h8)
	) name2026 (
		_w4169_,
		_w4171_,
		_w4172_
	);
	LUT2 #(
		.INIT('h2)
	) name2027 (
		_w2796_,
		_w4164_,
		_w4173_
	);
	LUT2 #(
		.INIT('h4)
	) name2028 (
		_w4172_,
		_w4173_,
		_w4174_
	);
	LUT2 #(
		.INIT('h8)
	) name2029 (
		\u6_mem_reg[1][18]/NET0131 ,
		_w2957_,
		_w4175_
	);
	LUT2 #(
		.INIT('h8)
	) name2030 (
		\u6_mem_reg[3][18]/NET0131 ,
		_w2801_,
		_w4176_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		\u6_mem_reg[2][18]/NET0131 ,
		_w2955_,
		_w4177_
	);
	LUT2 #(
		.INIT('h8)
	) name2032 (
		\u6_mem_reg[0][18]/NET0131 ,
		_w2959_,
		_w4178_
	);
	LUT2 #(
		.INIT('h1)
	) name2033 (
		_w4175_,
		_w4176_,
		_w4179_
	);
	LUT2 #(
		.INIT('h1)
	) name2034 (
		_w4177_,
		_w4178_,
		_w4180_
	);
	LUT2 #(
		.INIT('h8)
	) name2035 (
		_w4179_,
		_w4180_,
		_w4181_
	);
	LUT2 #(
		.INIT('h2)
	) name2036 (
		_w2964_,
		_w4181_,
		_w4182_
	);
	LUT2 #(
		.INIT('h2)
	) name2037 (
		_w3953_,
		_w4129_,
		_w4183_
	);
	LUT2 #(
		.INIT('h2)
	) name2038 (
		_w2795_,
		_w4182_,
		_w4184_
	);
	LUT2 #(
		.INIT('h4)
	) name2039 (
		_w4183_,
		_w4184_,
		_w4185_
	);
	LUT2 #(
		.INIT('h4)
	) name2040 (
		_w4174_,
		_w4185_,
		_w4186_
	);
	LUT2 #(
		.INIT('h2)
	) name2041 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4163_,
		_w4187_
	);
	LUT2 #(
		.INIT('h4)
	) name2042 (
		_w4186_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('h1)
	) name2043 (
		\u6_dout_reg[19]/P0001 ,
		_w2795_,
		_w4189_
	);
	LUT2 #(
		.INIT('h4)
	) name2044 (
		\u6_rp_reg[0]/P0001 ,
		_w4103_,
		_w4190_
	);
	LUT2 #(
		.INIT('h8)
	) name2045 (
		\u6_mem_reg[2][31]/NET0131 ,
		_w2955_,
		_w4191_
	);
	LUT2 #(
		.INIT('h8)
	) name2046 (
		\u6_mem_reg[3][31]/NET0131 ,
		_w2801_,
		_w4192_
	);
	LUT2 #(
		.INIT('h8)
	) name2047 (
		\u6_mem_reg[1][31]/NET0131 ,
		_w2957_,
		_w4193_
	);
	LUT2 #(
		.INIT('h8)
	) name2048 (
		\u6_mem_reg[0][31]/NET0131 ,
		_w2959_,
		_w4194_
	);
	LUT2 #(
		.INIT('h2)
	) name2049 (
		\u6_rp_reg[0]/P0001 ,
		_w4191_,
		_w4195_
	);
	LUT2 #(
		.INIT('h1)
	) name2050 (
		_w4192_,
		_w4193_,
		_w4196_
	);
	LUT2 #(
		.INIT('h4)
	) name2051 (
		_w4194_,
		_w4196_,
		_w4197_
	);
	LUT2 #(
		.INIT('h8)
	) name2052 (
		_w4195_,
		_w4197_,
		_w4198_
	);
	LUT2 #(
		.INIT('h2)
	) name2053 (
		_w2796_,
		_w4190_,
		_w4199_
	);
	LUT2 #(
		.INIT('h4)
	) name2054 (
		_w4198_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h8)
	) name2055 (
		\u6_mem_reg[2][19]/NET0131 ,
		_w2955_,
		_w4201_
	);
	LUT2 #(
		.INIT('h8)
	) name2056 (
		\u6_mem_reg[3][19]/NET0131 ,
		_w2801_,
		_w4202_
	);
	LUT2 #(
		.INIT('h8)
	) name2057 (
		\u6_mem_reg[1][19]/NET0131 ,
		_w2957_,
		_w4203_
	);
	LUT2 #(
		.INIT('h8)
	) name2058 (
		\u6_mem_reg[0][19]/NET0131 ,
		_w2959_,
		_w4204_
	);
	LUT2 #(
		.INIT('h1)
	) name2059 (
		_w4201_,
		_w4202_,
		_w4205_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		_w4203_,
		_w4204_,
		_w4206_
	);
	LUT2 #(
		.INIT('h8)
	) name2061 (
		_w4205_,
		_w4206_,
		_w4207_
	);
	LUT2 #(
		.INIT('h2)
	) name2062 (
		_w2964_,
		_w4207_,
		_w4208_
	);
	LUT2 #(
		.INIT('h2)
	) name2063 (
		_w3953_,
		_w4155_,
		_w4209_
	);
	LUT2 #(
		.INIT('h2)
	) name2064 (
		_w2795_,
		_w4208_,
		_w4210_
	);
	LUT2 #(
		.INIT('h4)
	) name2065 (
		_w4209_,
		_w4210_,
		_w4211_
	);
	LUT2 #(
		.INIT('h4)
	) name2066 (
		_w4200_,
		_w4211_,
		_w4212_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4189_,
		_w4213_
	);
	LUT2 #(
		.INIT('h4)
	) name2068 (
		_w4212_,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		\u6_dout_reg[2]/P0001 ,
		_w2795_,
		_w4215_
	);
	LUT2 #(
		.INIT('h4)
	) name2070 (
		_w2963_,
		_w3953_,
		_w4216_
	);
	LUT2 #(
		.INIT('h8)
	) name2071 (
		\u6_mem_reg[3][2]/NET0131 ,
		_w2801_,
		_w4217_
	);
	LUT2 #(
		.INIT('h8)
	) name2072 (
		\u6_mem_reg[2][2]/NET0131 ,
		_w2955_,
		_w4218_
	);
	LUT2 #(
		.INIT('h8)
	) name2073 (
		\u6_mem_reg[1][2]/NET0131 ,
		_w2957_,
		_w4219_
	);
	LUT2 #(
		.INIT('h8)
	) name2074 (
		\u6_mem_reg[0][2]/NET0131 ,
		_w2959_,
		_w4220_
	);
	LUT2 #(
		.INIT('h1)
	) name2075 (
		_w4217_,
		_w4218_,
		_w4221_
	);
	LUT2 #(
		.INIT('h1)
	) name2076 (
		_w4219_,
		_w4220_,
		_w4222_
	);
	LUT2 #(
		.INIT('h8)
	) name2077 (
		_w4221_,
		_w4222_,
		_w4223_
	);
	LUT2 #(
		.INIT('h2)
	) name2078 (
		_w2964_,
		_w4223_,
		_w4224_
	);
	LUT2 #(
		.INIT('h2)
	) name2079 (
		_w2795_,
		_w4216_,
		_w4225_
	);
	LUT2 #(
		.INIT('h4)
	) name2080 (
		_w4224_,
		_w4225_,
		_w4226_
	);
	LUT2 #(
		.INIT('h2)
	) name2081 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4215_,
		_w4227_
	);
	LUT2 #(
		.INIT('h4)
	) name2082 (
		_w4226_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h1)
	) name2083 (
		\u6_dout_reg[3]/P0001 ,
		_w2795_,
		_w4229_
	);
	LUT2 #(
		.INIT('h4)
	) name2084 (
		_w2976_,
		_w3953_,
		_w4230_
	);
	LUT2 #(
		.INIT('h8)
	) name2085 (
		\u6_mem_reg[3][3]/NET0131 ,
		_w2801_,
		_w4231_
	);
	LUT2 #(
		.INIT('h8)
	) name2086 (
		\u6_mem_reg[1][3]/NET0131 ,
		_w2957_,
		_w4232_
	);
	LUT2 #(
		.INIT('h8)
	) name2087 (
		\u6_mem_reg[2][3]/NET0131 ,
		_w2955_,
		_w4233_
	);
	LUT2 #(
		.INIT('h8)
	) name2088 (
		\u6_mem_reg[0][3]/NET0131 ,
		_w2959_,
		_w4234_
	);
	LUT2 #(
		.INIT('h1)
	) name2089 (
		_w4231_,
		_w4232_,
		_w4235_
	);
	LUT2 #(
		.INIT('h1)
	) name2090 (
		_w4233_,
		_w4234_,
		_w4236_
	);
	LUT2 #(
		.INIT('h8)
	) name2091 (
		_w4235_,
		_w4236_,
		_w4237_
	);
	LUT2 #(
		.INIT('h2)
	) name2092 (
		_w2964_,
		_w4237_,
		_w4238_
	);
	LUT2 #(
		.INIT('h2)
	) name2093 (
		_w2795_,
		_w4230_,
		_w4239_
	);
	LUT2 #(
		.INIT('h4)
	) name2094 (
		_w4238_,
		_w4239_,
		_w4240_
	);
	LUT2 #(
		.INIT('h2)
	) name2095 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4229_,
		_w4241_
	);
	LUT2 #(
		.INIT('h4)
	) name2096 (
		_w4240_,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h1)
	) name2097 (
		\u6_dout_reg[4]/P0001 ,
		_w2795_,
		_w4243_
	);
	LUT2 #(
		.INIT('h4)
	) name2098 (
		\u6_rp_reg[0]/P0001 ,
		_w2963_,
		_w4244_
	);
	LUT2 #(
		.INIT('h8)
	) name2099 (
		\u6_rp_reg[0]/P0001 ,
		_w4129_,
		_w4245_
	);
	LUT2 #(
		.INIT('h2)
	) name2100 (
		_w2796_,
		_w4244_,
		_w4246_
	);
	LUT2 #(
		.INIT('h4)
	) name2101 (
		_w4245_,
		_w4246_,
		_w4247_
	);
	LUT2 #(
		.INIT('h8)
	) name2102 (
		\u6_mem_reg[3][4]/NET0131 ,
		_w2801_,
		_w4248_
	);
	LUT2 #(
		.INIT('h8)
	) name2103 (
		\u6_mem_reg[2][4]/NET0131 ,
		_w2955_,
		_w4249_
	);
	LUT2 #(
		.INIT('h8)
	) name2104 (
		\u6_mem_reg[0][4]/NET0131 ,
		_w2959_,
		_w4250_
	);
	LUT2 #(
		.INIT('h8)
	) name2105 (
		\u6_mem_reg[1][4]/NET0131 ,
		_w2957_,
		_w4251_
	);
	LUT2 #(
		.INIT('h1)
	) name2106 (
		_w4248_,
		_w4249_,
		_w4252_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		_w4250_,
		_w4251_,
		_w4253_
	);
	LUT2 #(
		.INIT('h8)
	) name2108 (
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h2)
	) name2109 (
		_w2964_,
		_w4254_,
		_w4255_
	);
	LUT2 #(
		.INIT('h2)
	) name2110 (
		_w3953_,
		_w4223_,
		_w4256_
	);
	LUT2 #(
		.INIT('h2)
	) name2111 (
		_w2795_,
		_w4255_,
		_w4257_
	);
	LUT2 #(
		.INIT('h4)
	) name2112 (
		_w4256_,
		_w4257_,
		_w4258_
	);
	LUT2 #(
		.INIT('h4)
	) name2113 (
		_w4247_,
		_w4258_,
		_w4259_
	);
	LUT2 #(
		.INIT('h2)
	) name2114 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4243_,
		_w4260_
	);
	LUT2 #(
		.INIT('h4)
	) name2115 (
		_w4259_,
		_w4260_,
		_w4261_
	);
	LUT2 #(
		.INIT('h1)
	) name2116 (
		\u6_dout_reg[5]/P0001 ,
		_w2795_,
		_w4262_
	);
	LUT2 #(
		.INIT('h4)
	) name2117 (
		\u6_rp_reg[0]/P0001 ,
		_w2976_,
		_w4263_
	);
	LUT2 #(
		.INIT('h8)
	) name2118 (
		\u6_rp_reg[0]/P0001 ,
		_w4155_,
		_w4264_
	);
	LUT2 #(
		.INIT('h2)
	) name2119 (
		_w2796_,
		_w4263_,
		_w4265_
	);
	LUT2 #(
		.INIT('h4)
	) name2120 (
		_w4264_,
		_w4265_,
		_w4266_
	);
	LUT2 #(
		.INIT('h8)
	) name2121 (
		\u6_mem_reg[3][5]/NET0131 ,
		_w2801_,
		_w4267_
	);
	LUT2 #(
		.INIT('h8)
	) name2122 (
		\u6_mem_reg[2][5]/NET0131 ,
		_w2955_,
		_w4268_
	);
	LUT2 #(
		.INIT('h8)
	) name2123 (
		\u6_mem_reg[0][5]/NET0131 ,
		_w2959_,
		_w4269_
	);
	LUT2 #(
		.INIT('h8)
	) name2124 (
		\u6_mem_reg[1][5]/NET0131 ,
		_w2957_,
		_w4270_
	);
	LUT2 #(
		.INIT('h1)
	) name2125 (
		_w4267_,
		_w4268_,
		_w4271_
	);
	LUT2 #(
		.INIT('h1)
	) name2126 (
		_w4269_,
		_w4270_,
		_w4272_
	);
	LUT2 #(
		.INIT('h8)
	) name2127 (
		_w4271_,
		_w4272_,
		_w4273_
	);
	LUT2 #(
		.INIT('h2)
	) name2128 (
		_w2964_,
		_w4273_,
		_w4274_
	);
	LUT2 #(
		.INIT('h2)
	) name2129 (
		_w3953_,
		_w4237_,
		_w4275_
	);
	LUT2 #(
		.INIT('h2)
	) name2130 (
		_w2795_,
		_w4274_,
		_w4276_
	);
	LUT2 #(
		.INIT('h4)
	) name2131 (
		_w4275_,
		_w4276_,
		_w4277_
	);
	LUT2 #(
		.INIT('h4)
	) name2132 (
		_w4266_,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h2)
	) name2133 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4262_,
		_w4279_
	);
	LUT2 #(
		.INIT('h4)
	) name2134 (
		_w4278_,
		_w4279_,
		_w4280_
	);
	LUT2 #(
		.INIT('h1)
	) name2135 (
		\u6_dout_reg[6]/P0001 ,
		_w2795_,
		_w4281_
	);
	LUT2 #(
		.INIT('h4)
	) name2136 (
		\u6_rp_reg[0]/P0001 ,
		_w4223_,
		_w4282_
	);
	LUT2 #(
		.INIT('h8)
	) name2137 (
		\u6_rp_reg[0]/P0001 ,
		_w4181_,
		_w4283_
	);
	LUT2 #(
		.INIT('h2)
	) name2138 (
		_w2796_,
		_w4282_,
		_w4284_
	);
	LUT2 #(
		.INIT('h4)
	) name2139 (
		_w4283_,
		_w4284_,
		_w4285_
	);
	LUT2 #(
		.INIT('h2)
	) name2140 (
		_w2964_,
		_w3933_,
		_w4286_
	);
	LUT2 #(
		.INIT('h2)
	) name2141 (
		_w3953_,
		_w4254_,
		_w4287_
	);
	LUT2 #(
		.INIT('h2)
	) name2142 (
		_w2795_,
		_w4286_,
		_w4288_
	);
	LUT2 #(
		.INIT('h4)
	) name2143 (
		_w4287_,
		_w4288_,
		_w4289_
	);
	LUT2 #(
		.INIT('h4)
	) name2144 (
		_w4285_,
		_w4289_,
		_w4290_
	);
	LUT2 #(
		.INIT('h2)
	) name2145 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4281_,
		_w4291_
	);
	LUT2 #(
		.INIT('h4)
	) name2146 (
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h1)
	) name2147 (
		\u6_dout_reg[7]/P0001 ,
		_w2795_,
		_w4293_
	);
	LUT2 #(
		.INIT('h4)
	) name2148 (
		\u6_rp_reg[0]/P0001 ,
		_w4237_,
		_w4294_
	);
	LUT2 #(
		.INIT('h8)
	) name2149 (
		\u6_rp_reg[0]/P0001 ,
		_w4207_,
		_w4295_
	);
	LUT2 #(
		.INIT('h2)
	) name2150 (
		_w2796_,
		_w4294_,
		_w4296_
	);
	LUT2 #(
		.INIT('h4)
	) name2151 (
		_w4295_,
		_w4296_,
		_w4297_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		_w2964_,
		_w3974_,
		_w4298_
	);
	LUT2 #(
		.INIT('h2)
	) name2153 (
		_w3953_,
		_w4273_,
		_w4299_
	);
	LUT2 #(
		.INIT('h2)
	) name2154 (
		_w2795_,
		_w4298_,
		_w4300_
	);
	LUT2 #(
		.INIT('h4)
	) name2155 (
		_w4299_,
		_w4300_,
		_w4301_
	);
	LUT2 #(
		.INIT('h4)
	) name2156 (
		_w4297_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('h2)
	) name2157 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4293_,
		_w4303_
	);
	LUT2 #(
		.INIT('h4)
	) name2158 (
		_w4302_,
		_w4303_,
		_w4304_
	);
	LUT2 #(
		.INIT('h1)
	) name2159 (
		\u6_dout_reg[8]/P0001 ,
		_w2795_,
		_w4305_
	);
	LUT2 #(
		.INIT('h4)
	) name2160 (
		\u6_rp_reg[0]/P0001 ,
		_w4254_,
		_w4306_
	);
	LUT2 #(
		.INIT('h8)
	) name2161 (
		\u6_mem_reg[2][20]/NET0131 ,
		_w2955_,
		_w4307_
	);
	LUT2 #(
		.INIT('h8)
	) name2162 (
		\u6_mem_reg[3][20]/NET0131 ,
		_w2801_,
		_w4308_
	);
	LUT2 #(
		.INIT('h8)
	) name2163 (
		\u6_mem_reg[1][20]/NET0131 ,
		_w2957_,
		_w4309_
	);
	LUT2 #(
		.INIT('h8)
	) name2164 (
		\u6_mem_reg[0][20]/NET0131 ,
		_w2959_,
		_w4310_
	);
	LUT2 #(
		.INIT('h2)
	) name2165 (
		\u6_rp_reg[0]/P0001 ,
		_w4307_,
		_w4311_
	);
	LUT2 #(
		.INIT('h1)
	) name2166 (
		_w4308_,
		_w4309_,
		_w4312_
	);
	LUT2 #(
		.INIT('h4)
	) name2167 (
		_w4310_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h8)
	) name2168 (
		_w4311_,
		_w4313_,
		_w4314_
	);
	LUT2 #(
		.INIT('h2)
	) name2169 (
		_w2796_,
		_w4306_,
		_w4315_
	);
	LUT2 #(
		.INIT('h4)
	) name2170 (
		_w4314_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h2)
	) name2171 (
		_w2964_,
		_w3960_,
		_w4317_
	);
	LUT2 #(
		.INIT('h4)
	) name2172 (
		_w3933_,
		_w3953_,
		_w4318_
	);
	LUT2 #(
		.INIT('h2)
	) name2173 (
		_w2795_,
		_w4317_,
		_w4319_
	);
	LUT2 #(
		.INIT('h4)
	) name2174 (
		_w4318_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h4)
	) name2175 (
		_w4316_,
		_w4320_,
		_w4321_
	);
	LUT2 #(
		.INIT('h2)
	) name2176 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4305_,
		_w4322_
	);
	LUT2 #(
		.INIT('h4)
	) name2177 (
		_w4321_,
		_w4322_,
		_w4323_
	);
	LUT2 #(
		.INIT('h1)
	) name2178 (
		\u6_dout_reg[9]/P0001 ,
		_w2795_,
		_w4324_
	);
	LUT2 #(
		.INIT('h4)
	) name2179 (
		\u6_rp_reg[0]/P0001 ,
		_w4273_,
		_w4325_
	);
	LUT2 #(
		.INIT('h8)
	) name2180 (
		\u6_mem_reg[2][21]/NET0131 ,
		_w2955_,
		_w4326_
	);
	LUT2 #(
		.INIT('h8)
	) name2181 (
		\u6_mem_reg[1][21]/NET0131 ,
		_w2957_,
		_w4327_
	);
	LUT2 #(
		.INIT('h8)
	) name2182 (
		\u6_mem_reg[3][21]/NET0131 ,
		_w2801_,
		_w4328_
	);
	LUT2 #(
		.INIT('h8)
	) name2183 (
		\u6_mem_reg[0][21]/NET0131 ,
		_w2959_,
		_w4329_
	);
	LUT2 #(
		.INIT('h2)
	) name2184 (
		\u6_rp_reg[0]/P0001 ,
		_w4326_,
		_w4330_
	);
	LUT2 #(
		.INIT('h1)
	) name2185 (
		_w4327_,
		_w4328_,
		_w4331_
	);
	LUT2 #(
		.INIT('h4)
	) name2186 (
		_w4329_,
		_w4331_,
		_w4332_
	);
	LUT2 #(
		.INIT('h8)
	) name2187 (
		_w4330_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h2)
	) name2188 (
		_w2796_,
		_w4325_,
		_w4334_
	);
	LUT2 #(
		.INIT('h4)
	) name2189 (
		_w4333_,
		_w4334_,
		_w4335_
	);
	LUT2 #(
		.INIT('h2)
	) name2190 (
		_w2964_,
		_w4000_,
		_w4336_
	);
	LUT2 #(
		.INIT('h2)
	) name2191 (
		_w3953_,
		_w3974_,
		_w4337_
	);
	LUT2 #(
		.INIT('h2)
	) name2192 (
		_w2795_,
		_w4336_,
		_w4338_
	);
	LUT2 #(
		.INIT('h4)
	) name2193 (
		_w4337_,
		_w4338_,
		_w4339_
	);
	LUT2 #(
		.INIT('h4)
	) name2194 (
		_w4335_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h2)
	) name2195 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w4324_,
		_w4341_
	);
	LUT2 #(
		.INIT('h4)
	) name2196 (
		_w4340_,
		_w4341_,
		_w4342_
	);
	LUT2 #(
		.INIT('h1)
	) name2197 (
		\u7_dout_reg[10]/P0001 ,
		_w2808_,
		_w4343_
	);
	LUT2 #(
		.INIT('h8)
	) name2198 (
		\u7_mem_reg[2][6]/NET0131 ,
		_w2983_,
		_w4344_
	);
	LUT2 #(
		.INIT('h8)
	) name2199 (
		\u7_mem_reg[3][6]/NET0131 ,
		_w2981_,
		_w4345_
	);
	LUT2 #(
		.INIT('h8)
	) name2200 (
		\u7_mem_reg[0][6]/NET0131 ,
		_w2987_,
		_w4346_
	);
	LUT2 #(
		.INIT('h8)
	) name2201 (
		\u7_mem_reg[1][6]/NET0131 ,
		_w2985_,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name2202 (
		_w4344_,
		_w4345_,
		_w4348_
	);
	LUT2 #(
		.INIT('h1)
	) name2203 (
		_w4346_,
		_w4347_,
		_w4349_
	);
	LUT2 #(
		.INIT('h8)
	) name2204 (
		_w4348_,
		_w4349_,
		_w4350_
	);
	LUT2 #(
		.INIT('h2)
	) name2205 (
		_w2806_,
		_w4350_,
		_w4351_
	);
	LUT2 #(
		.INIT('h2)
	) name2206 (
		\u13_occ1_r_reg[2]/NET0131 ,
		\u13_occ1_r_reg[3]/NET0131 ,
		_w4352_
	);
	LUT2 #(
		.INIT('h8)
	) name2207 (
		\u7_mem_reg[3][8]/NET0131 ,
		_w2981_,
		_w4353_
	);
	LUT2 #(
		.INIT('h8)
	) name2208 (
		\u7_mem_reg[2][8]/NET0131 ,
		_w2983_,
		_w4354_
	);
	LUT2 #(
		.INIT('h8)
	) name2209 (
		\u7_mem_reg[1][8]/NET0131 ,
		_w2985_,
		_w4355_
	);
	LUT2 #(
		.INIT('h8)
	) name2210 (
		\u7_mem_reg[0][8]/NET0131 ,
		_w2987_,
		_w4356_
	);
	LUT2 #(
		.INIT('h1)
	) name2211 (
		_w4353_,
		_w4354_,
		_w4357_
	);
	LUT2 #(
		.INIT('h1)
	) name2212 (
		_w4355_,
		_w4356_,
		_w4358_
	);
	LUT2 #(
		.INIT('h8)
	) name2213 (
		_w4357_,
		_w4358_,
		_w4359_
	);
	LUT2 #(
		.INIT('h2)
	) name2214 (
		_w4352_,
		_w4359_,
		_w4360_
	);
	LUT2 #(
		.INIT('h8)
	) name2215 (
		\u7_rp_reg[0]/P0001 ,
		_w2805_,
		_w4361_
	);
	LUT2 #(
		.INIT('h8)
	) name2216 (
		\u7_mem_reg[3][22]/NET0131 ,
		_w2981_,
		_w4362_
	);
	LUT2 #(
		.INIT('h8)
	) name2217 (
		\u7_mem_reg[0][22]/NET0131 ,
		_w2987_,
		_w4363_
	);
	LUT2 #(
		.INIT('h8)
	) name2218 (
		\u7_mem_reg[1][22]/NET0131 ,
		_w2985_,
		_w4364_
	);
	LUT2 #(
		.INIT('h8)
	) name2219 (
		\u7_mem_reg[2][22]/NET0131 ,
		_w2983_,
		_w4365_
	);
	LUT2 #(
		.INIT('h1)
	) name2220 (
		_w4362_,
		_w4363_,
		_w4366_
	);
	LUT2 #(
		.INIT('h1)
	) name2221 (
		_w4364_,
		_w4365_,
		_w4367_
	);
	LUT2 #(
		.INIT('h8)
	) name2222 (
		_w4366_,
		_w4367_,
		_w4368_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		_w4361_,
		_w4368_,
		_w4369_
	);
	LUT2 #(
		.INIT('h8)
	) name2224 (
		\u7_mem_reg[3][10]/NET0131 ,
		_w2981_,
		_w4370_
	);
	LUT2 #(
		.INIT('h8)
	) name2225 (
		\u7_mem_reg[2][10]/NET0131 ,
		_w2983_,
		_w4371_
	);
	LUT2 #(
		.INIT('h8)
	) name2226 (
		\u7_mem_reg[1][10]/NET0131 ,
		_w2985_,
		_w4372_
	);
	LUT2 #(
		.INIT('h8)
	) name2227 (
		\u7_mem_reg[0][10]/NET0131 ,
		_w2987_,
		_w4373_
	);
	LUT2 #(
		.INIT('h1)
	) name2228 (
		_w4370_,
		_w4371_,
		_w4374_
	);
	LUT2 #(
		.INIT('h1)
	) name2229 (
		_w4372_,
		_w4373_,
		_w4375_
	);
	LUT2 #(
		.INIT('h8)
	) name2230 (
		_w4374_,
		_w4375_,
		_w4376_
	);
	LUT2 #(
		.INIT('h2)
	) name2231 (
		_w2992_,
		_w4376_,
		_w4377_
	);
	LUT2 #(
		.INIT('h2)
	) name2232 (
		_w2808_,
		_w4351_,
		_w4378_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w4360_,
		_w4369_,
		_w4379_
	);
	LUT2 #(
		.INIT('h4)
	) name2234 (
		_w4377_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h8)
	) name2235 (
		_w4378_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h2)
	) name2236 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4343_,
		_w4382_
	);
	LUT2 #(
		.INIT('h4)
	) name2237 (
		_w4381_,
		_w4382_,
		_w4383_
	);
	LUT2 #(
		.INIT('h1)
	) name2238 (
		\u7_dout_reg[11]/P0001 ,
		_w2808_,
		_w4384_
	);
	LUT2 #(
		.INIT('h8)
	) name2239 (
		\u7_mem_reg[1][11]/NET0131 ,
		_w2985_,
		_w4385_
	);
	LUT2 #(
		.INIT('h8)
	) name2240 (
		\u7_mem_reg[2][11]/NET0131 ,
		_w2983_,
		_w4386_
	);
	LUT2 #(
		.INIT('h8)
	) name2241 (
		\u7_mem_reg[0][11]/NET0131 ,
		_w2987_,
		_w4387_
	);
	LUT2 #(
		.INIT('h8)
	) name2242 (
		\u7_mem_reg[3][11]/NET0131 ,
		_w2981_,
		_w4388_
	);
	LUT2 #(
		.INIT('h1)
	) name2243 (
		_w4385_,
		_w4386_,
		_w4389_
	);
	LUT2 #(
		.INIT('h1)
	) name2244 (
		_w4387_,
		_w4388_,
		_w4390_
	);
	LUT2 #(
		.INIT('h8)
	) name2245 (
		_w4389_,
		_w4390_,
		_w4391_
	);
	LUT2 #(
		.INIT('h2)
	) name2246 (
		_w2992_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h8)
	) name2247 (
		\u7_mem_reg[1][7]/NET0131 ,
		_w2985_,
		_w4393_
	);
	LUT2 #(
		.INIT('h8)
	) name2248 (
		\u7_mem_reg[3][7]/NET0131 ,
		_w2981_,
		_w4394_
	);
	LUT2 #(
		.INIT('h8)
	) name2249 (
		\u7_mem_reg[2][7]/NET0131 ,
		_w2983_,
		_w4395_
	);
	LUT2 #(
		.INIT('h8)
	) name2250 (
		\u7_mem_reg[0][7]/NET0131 ,
		_w2987_,
		_w4396_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		_w4393_,
		_w4394_,
		_w4397_
	);
	LUT2 #(
		.INIT('h1)
	) name2252 (
		_w4395_,
		_w4396_,
		_w4398_
	);
	LUT2 #(
		.INIT('h8)
	) name2253 (
		_w4397_,
		_w4398_,
		_w4399_
	);
	LUT2 #(
		.INIT('h2)
	) name2254 (
		_w2806_,
		_w4399_,
		_w4400_
	);
	LUT2 #(
		.INIT('h8)
	) name2255 (
		\u7_mem_reg[2][23]/NET0131 ,
		_w2983_,
		_w4401_
	);
	LUT2 #(
		.INIT('h8)
	) name2256 (
		\u7_mem_reg[0][23]/NET0131 ,
		_w2987_,
		_w4402_
	);
	LUT2 #(
		.INIT('h8)
	) name2257 (
		\u7_mem_reg[1][23]/NET0131 ,
		_w2985_,
		_w4403_
	);
	LUT2 #(
		.INIT('h8)
	) name2258 (
		\u7_mem_reg[3][23]/NET0131 ,
		_w2981_,
		_w4404_
	);
	LUT2 #(
		.INIT('h1)
	) name2259 (
		_w4401_,
		_w4402_,
		_w4405_
	);
	LUT2 #(
		.INIT('h1)
	) name2260 (
		_w4403_,
		_w4404_,
		_w4406_
	);
	LUT2 #(
		.INIT('h8)
	) name2261 (
		_w4405_,
		_w4406_,
		_w4407_
	);
	LUT2 #(
		.INIT('h2)
	) name2262 (
		_w4361_,
		_w4407_,
		_w4408_
	);
	LUT2 #(
		.INIT('h8)
	) name2263 (
		\u7_mem_reg[3][9]/NET0131 ,
		_w2981_,
		_w4409_
	);
	LUT2 #(
		.INIT('h8)
	) name2264 (
		\u7_mem_reg[0][9]/NET0131 ,
		_w2987_,
		_w4410_
	);
	LUT2 #(
		.INIT('h8)
	) name2265 (
		\u7_mem_reg[2][9]/NET0131 ,
		_w2983_,
		_w4411_
	);
	LUT2 #(
		.INIT('h8)
	) name2266 (
		\u7_mem_reg[1][9]/NET0131 ,
		_w2985_,
		_w4412_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		_w4409_,
		_w4410_,
		_w4413_
	);
	LUT2 #(
		.INIT('h1)
	) name2268 (
		_w4411_,
		_w4412_,
		_w4414_
	);
	LUT2 #(
		.INIT('h8)
	) name2269 (
		_w4413_,
		_w4414_,
		_w4415_
	);
	LUT2 #(
		.INIT('h2)
	) name2270 (
		_w4352_,
		_w4415_,
		_w4416_
	);
	LUT2 #(
		.INIT('h2)
	) name2271 (
		_w2808_,
		_w4392_,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name2272 (
		_w4400_,
		_w4408_,
		_w4418_
	);
	LUT2 #(
		.INIT('h4)
	) name2273 (
		_w4416_,
		_w4418_,
		_w4419_
	);
	LUT2 #(
		.INIT('h8)
	) name2274 (
		_w4417_,
		_w4419_,
		_w4420_
	);
	LUT2 #(
		.INIT('h2)
	) name2275 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4384_,
		_w4421_
	);
	LUT2 #(
		.INIT('h4)
	) name2276 (
		_w4420_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h1)
	) name2277 (
		\u13_icc_r_reg[5]/NET0131 ,
		\u9_status_reg[1]/P0001 ,
		_w4423_
	);
	LUT2 #(
		.INIT('h8)
	) name2278 (
		\u13_icc_r_reg[5]/NET0131 ,
		\u9_status_reg[1]/P0001 ,
		_w4424_
	);
	LUT2 #(
		.INIT('h1)
	) name2279 (
		\u13_icc_r_reg[4]/NET0131 ,
		\u9_status_reg[0]/P0001 ,
		_w4425_
	);
	LUT2 #(
		.INIT('h4)
	) name2280 (
		_w4424_,
		_w4425_,
		_w4426_
	);
	LUT2 #(
		.INIT('h1)
	) name2281 (
		\u9_full_reg/NET0131 ,
		_w4423_,
		_w4427_
	);
	LUT2 #(
		.INIT('h4)
	) name2282 (
		_w4426_,
		_w4427_,
		_w4428_
	);
	LUT2 #(
		.INIT('h2)
	) name2283 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w4428_,
		_w4429_
	);
	LUT2 #(
		.INIT('h1)
	) name2284 (
		\u7_dout_reg[12]/P0001 ,
		_w2808_,
		_w4430_
	);
	LUT2 #(
		.INIT('h4)
	) name2285 (
		\u7_rp_reg[0]/P0001 ,
		_w4359_,
		_w4431_
	);
	LUT2 #(
		.INIT('h8)
	) name2286 (
		\u7_mem_reg[2][24]/NET0131 ,
		_w2983_,
		_w4432_
	);
	LUT2 #(
		.INIT('h8)
	) name2287 (
		\u7_mem_reg[3][24]/NET0131 ,
		_w2981_,
		_w4433_
	);
	LUT2 #(
		.INIT('h8)
	) name2288 (
		\u7_mem_reg[1][24]/NET0131 ,
		_w2985_,
		_w4434_
	);
	LUT2 #(
		.INIT('h8)
	) name2289 (
		\u7_mem_reg[0][24]/NET0131 ,
		_w2987_,
		_w4435_
	);
	LUT2 #(
		.INIT('h2)
	) name2290 (
		\u7_rp_reg[0]/P0001 ,
		_w4432_,
		_w4436_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		_w4433_,
		_w4434_,
		_w4437_
	);
	LUT2 #(
		.INIT('h4)
	) name2292 (
		_w4435_,
		_w4437_,
		_w4438_
	);
	LUT2 #(
		.INIT('h8)
	) name2293 (
		_w4436_,
		_w4438_,
		_w4439_
	);
	LUT2 #(
		.INIT('h2)
	) name2294 (
		_w2805_,
		_w4431_,
		_w4440_
	);
	LUT2 #(
		.INIT('h4)
	) name2295 (
		_w4439_,
		_w4440_,
		_w4441_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		\u7_mem_reg[3][12]/NET0131 ,
		_w2981_,
		_w4442_
	);
	LUT2 #(
		.INIT('h8)
	) name2297 (
		\u7_mem_reg[2][12]/NET0131 ,
		_w2983_,
		_w4443_
	);
	LUT2 #(
		.INIT('h8)
	) name2298 (
		\u7_mem_reg[1][12]/NET0131 ,
		_w2985_,
		_w4444_
	);
	LUT2 #(
		.INIT('h8)
	) name2299 (
		\u7_mem_reg[0][12]/NET0131 ,
		_w2987_,
		_w4445_
	);
	LUT2 #(
		.INIT('h1)
	) name2300 (
		_w4442_,
		_w4443_,
		_w4446_
	);
	LUT2 #(
		.INIT('h1)
	) name2301 (
		_w4444_,
		_w4445_,
		_w4447_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		_w4446_,
		_w4447_,
		_w4448_
	);
	LUT2 #(
		.INIT('h2)
	) name2303 (
		_w2992_,
		_w4448_,
		_w4449_
	);
	LUT2 #(
		.INIT('h2)
	) name2304 (
		_w4352_,
		_w4376_,
		_w4450_
	);
	LUT2 #(
		.INIT('h2)
	) name2305 (
		_w2808_,
		_w4449_,
		_w4451_
	);
	LUT2 #(
		.INIT('h4)
	) name2306 (
		_w4450_,
		_w4451_,
		_w4452_
	);
	LUT2 #(
		.INIT('h4)
	) name2307 (
		_w4441_,
		_w4452_,
		_w4453_
	);
	LUT2 #(
		.INIT('h2)
	) name2308 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4430_,
		_w4454_
	);
	LUT2 #(
		.INIT('h4)
	) name2309 (
		_w4453_,
		_w4454_,
		_w4455_
	);
	LUT2 #(
		.INIT('h8)
	) name2310 (
		\u10_status_reg[1]/P0001 ,
		\u13_icc_r_reg[13]/NET0131 ,
		_w4456_
	);
	LUT2 #(
		.INIT('h1)
	) name2311 (
		\u10_status_reg[0]/P0001 ,
		\u13_icc_r_reg[12]/NET0131 ,
		_w4457_
	);
	LUT2 #(
		.INIT('h4)
	) name2312 (
		_w4456_,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h1)
	) name2313 (
		\u10_status_reg[1]/P0001 ,
		\u13_icc_r_reg[13]/NET0131 ,
		_w4459_
	);
	LUT2 #(
		.INIT('h1)
	) name2314 (
		\u10_full_reg/NET0131 ,
		_w4459_,
		_w4460_
	);
	LUT2 #(
		.INIT('h4)
	) name2315 (
		_w4458_,
		_w4460_,
		_w4461_
	);
	LUT2 #(
		.INIT('h2)
	) name2316 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h1)
	) name2317 (
		\u7_dout_reg[13]/P0001 ,
		_w2808_,
		_w4463_
	);
	LUT2 #(
		.INIT('h2)
	) name2318 (
		_w4352_,
		_w4391_,
		_w4464_
	);
	LUT2 #(
		.INIT('h8)
	) name2319 (
		\u7_mem_reg[3][13]/NET0131 ,
		_w2981_,
		_w4465_
	);
	LUT2 #(
		.INIT('h8)
	) name2320 (
		\u7_mem_reg[2][13]/NET0131 ,
		_w2983_,
		_w4466_
	);
	LUT2 #(
		.INIT('h8)
	) name2321 (
		\u7_mem_reg[1][13]/NET0131 ,
		_w2985_,
		_w4467_
	);
	LUT2 #(
		.INIT('h8)
	) name2322 (
		\u7_mem_reg[0][13]/NET0131 ,
		_w2987_,
		_w4468_
	);
	LUT2 #(
		.INIT('h1)
	) name2323 (
		_w4465_,
		_w4466_,
		_w4469_
	);
	LUT2 #(
		.INIT('h1)
	) name2324 (
		_w4467_,
		_w4468_,
		_w4470_
	);
	LUT2 #(
		.INIT('h8)
	) name2325 (
		_w4469_,
		_w4470_,
		_w4471_
	);
	LUT2 #(
		.INIT('h2)
	) name2326 (
		_w2992_,
		_w4471_,
		_w4472_
	);
	LUT2 #(
		.INIT('h4)
	) name2327 (
		\u7_rp_reg[0]/P0001 ,
		_w4415_,
		_w4473_
	);
	LUT2 #(
		.INIT('h8)
	) name2328 (
		\u7_mem_reg[2][25]/NET0131 ,
		_w2983_,
		_w4474_
	);
	LUT2 #(
		.INIT('h8)
	) name2329 (
		\u7_mem_reg[3][25]/NET0131 ,
		_w2981_,
		_w4475_
	);
	LUT2 #(
		.INIT('h8)
	) name2330 (
		\u7_mem_reg[1][25]/NET0131 ,
		_w2985_,
		_w4476_
	);
	LUT2 #(
		.INIT('h8)
	) name2331 (
		\u7_mem_reg[0][25]/NET0131 ,
		_w2987_,
		_w4477_
	);
	LUT2 #(
		.INIT('h2)
	) name2332 (
		\u7_rp_reg[0]/P0001 ,
		_w4474_,
		_w4478_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		_w4475_,
		_w4476_,
		_w4479_
	);
	LUT2 #(
		.INIT('h4)
	) name2334 (
		_w4477_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h8)
	) name2335 (
		_w4478_,
		_w4480_,
		_w4481_
	);
	LUT2 #(
		.INIT('h2)
	) name2336 (
		_w2805_,
		_w4473_,
		_w4482_
	);
	LUT2 #(
		.INIT('h4)
	) name2337 (
		_w4481_,
		_w4482_,
		_w4483_
	);
	LUT2 #(
		.INIT('h2)
	) name2338 (
		_w2808_,
		_w4464_,
		_w4484_
	);
	LUT2 #(
		.INIT('h4)
	) name2339 (
		_w4472_,
		_w4484_,
		_w4485_
	);
	LUT2 #(
		.INIT('h4)
	) name2340 (
		_w4483_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h2)
	) name2341 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4463_,
		_w4487_
	);
	LUT2 #(
		.INIT('h4)
	) name2342 (
		_w4486_,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h1)
	) name2343 (
		\u7_dout_reg[14]/P0001 ,
		_w2808_,
		_w4489_
	);
	LUT2 #(
		.INIT('h4)
	) name2344 (
		\u7_rp_reg[0]/P0001 ,
		_w4376_,
		_w4490_
	);
	LUT2 #(
		.INIT('h8)
	) name2345 (
		\u7_mem_reg[2][26]/NET0131 ,
		_w2983_,
		_w4491_
	);
	LUT2 #(
		.INIT('h8)
	) name2346 (
		\u7_mem_reg[3][26]/NET0131 ,
		_w2981_,
		_w4492_
	);
	LUT2 #(
		.INIT('h8)
	) name2347 (
		\u7_mem_reg[1][26]/NET0131 ,
		_w2985_,
		_w4493_
	);
	LUT2 #(
		.INIT('h8)
	) name2348 (
		\u7_mem_reg[0][26]/NET0131 ,
		_w2987_,
		_w4494_
	);
	LUT2 #(
		.INIT('h2)
	) name2349 (
		\u7_rp_reg[0]/P0001 ,
		_w4491_,
		_w4495_
	);
	LUT2 #(
		.INIT('h1)
	) name2350 (
		_w4492_,
		_w4493_,
		_w4496_
	);
	LUT2 #(
		.INIT('h4)
	) name2351 (
		_w4494_,
		_w4496_,
		_w4497_
	);
	LUT2 #(
		.INIT('h8)
	) name2352 (
		_w4495_,
		_w4497_,
		_w4498_
	);
	LUT2 #(
		.INIT('h2)
	) name2353 (
		_w2805_,
		_w4490_,
		_w4499_
	);
	LUT2 #(
		.INIT('h4)
	) name2354 (
		_w4498_,
		_w4499_,
		_w4500_
	);
	LUT2 #(
		.INIT('h8)
	) name2355 (
		\u7_mem_reg[3][14]/NET0131 ,
		_w2981_,
		_w4501_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		\u7_mem_reg[2][14]/NET0131 ,
		_w2983_,
		_w4502_
	);
	LUT2 #(
		.INIT('h8)
	) name2357 (
		\u7_mem_reg[1][14]/NET0131 ,
		_w2985_,
		_w4503_
	);
	LUT2 #(
		.INIT('h8)
	) name2358 (
		\u7_mem_reg[0][14]/NET0131 ,
		_w2987_,
		_w4504_
	);
	LUT2 #(
		.INIT('h1)
	) name2359 (
		_w4501_,
		_w4502_,
		_w4505_
	);
	LUT2 #(
		.INIT('h1)
	) name2360 (
		_w4503_,
		_w4504_,
		_w4506_
	);
	LUT2 #(
		.INIT('h8)
	) name2361 (
		_w4505_,
		_w4506_,
		_w4507_
	);
	LUT2 #(
		.INIT('h2)
	) name2362 (
		_w2992_,
		_w4507_,
		_w4508_
	);
	LUT2 #(
		.INIT('h2)
	) name2363 (
		_w4352_,
		_w4448_,
		_w4509_
	);
	LUT2 #(
		.INIT('h2)
	) name2364 (
		_w2808_,
		_w4508_,
		_w4510_
	);
	LUT2 #(
		.INIT('h4)
	) name2365 (
		_w4509_,
		_w4510_,
		_w4511_
	);
	LUT2 #(
		.INIT('h4)
	) name2366 (
		_w4500_,
		_w4511_,
		_w4512_
	);
	LUT2 #(
		.INIT('h2)
	) name2367 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4489_,
		_w4513_
	);
	LUT2 #(
		.INIT('h4)
	) name2368 (
		_w4512_,
		_w4513_,
		_w4514_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		\u7_dout_reg[15]/P0001 ,
		_w2808_,
		_w4515_
	);
	LUT2 #(
		.INIT('h2)
	) name2370 (
		_w2806_,
		_w4391_,
		_w4516_
	);
	LUT2 #(
		.INIT('h2)
	) name2371 (
		_w4352_,
		_w4471_,
		_w4517_
	);
	LUT2 #(
		.INIT('h8)
	) name2372 (
		\u7_mem_reg[1][27]/NET0131 ,
		_w2985_,
		_w4518_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		\u7_mem_reg[0][27]/NET0131 ,
		_w2987_,
		_w4519_
	);
	LUT2 #(
		.INIT('h8)
	) name2374 (
		\u7_mem_reg[2][27]/NET0131 ,
		_w2983_,
		_w4520_
	);
	LUT2 #(
		.INIT('h8)
	) name2375 (
		\u7_mem_reg[3][27]/NET0131 ,
		_w2981_,
		_w4521_
	);
	LUT2 #(
		.INIT('h1)
	) name2376 (
		_w4518_,
		_w4519_,
		_w4522_
	);
	LUT2 #(
		.INIT('h1)
	) name2377 (
		_w4520_,
		_w4521_,
		_w4523_
	);
	LUT2 #(
		.INIT('h8)
	) name2378 (
		_w4522_,
		_w4523_,
		_w4524_
	);
	LUT2 #(
		.INIT('h2)
	) name2379 (
		_w4361_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h8)
	) name2380 (
		\u7_mem_reg[1][15]/NET0131 ,
		_w2985_,
		_w4526_
	);
	LUT2 #(
		.INIT('h8)
	) name2381 (
		\u7_mem_reg[3][15]/NET0131 ,
		_w2981_,
		_w4527_
	);
	LUT2 #(
		.INIT('h8)
	) name2382 (
		\u7_mem_reg[2][15]/NET0131 ,
		_w2983_,
		_w4528_
	);
	LUT2 #(
		.INIT('h8)
	) name2383 (
		\u7_mem_reg[0][15]/NET0131 ,
		_w2987_,
		_w4529_
	);
	LUT2 #(
		.INIT('h1)
	) name2384 (
		_w4526_,
		_w4527_,
		_w4530_
	);
	LUT2 #(
		.INIT('h1)
	) name2385 (
		_w4528_,
		_w4529_,
		_w4531_
	);
	LUT2 #(
		.INIT('h8)
	) name2386 (
		_w4530_,
		_w4531_,
		_w4532_
	);
	LUT2 #(
		.INIT('h2)
	) name2387 (
		_w2992_,
		_w4532_,
		_w4533_
	);
	LUT2 #(
		.INIT('h2)
	) name2388 (
		_w2808_,
		_w4516_,
		_w4534_
	);
	LUT2 #(
		.INIT('h1)
	) name2389 (
		_w4517_,
		_w4525_,
		_w4535_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		_w4533_,
		_w4535_,
		_w4536_
	);
	LUT2 #(
		.INIT('h8)
	) name2391 (
		_w4534_,
		_w4536_,
		_w4537_
	);
	LUT2 #(
		.INIT('h2)
	) name2392 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4515_,
		_w4538_
	);
	LUT2 #(
		.INIT('h4)
	) name2393 (
		_w4537_,
		_w4538_,
		_w4539_
	);
	LUT2 #(
		.INIT('h1)
	) name2394 (
		\u7_dout_reg[16]/P0001 ,
		_w2808_,
		_w4540_
	);
	LUT2 #(
		.INIT('h4)
	) name2395 (
		\u7_rp_reg[0]/P0001 ,
		_w4448_,
		_w4541_
	);
	LUT2 #(
		.INIT('h8)
	) name2396 (
		\u7_mem_reg[2][28]/NET0131 ,
		_w2983_,
		_w4542_
	);
	LUT2 #(
		.INIT('h8)
	) name2397 (
		\u7_mem_reg[3][28]/NET0131 ,
		_w2981_,
		_w4543_
	);
	LUT2 #(
		.INIT('h8)
	) name2398 (
		\u7_mem_reg[1][28]/NET0131 ,
		_w2985_,
		_w4544_
	);
	LUT2 #(
		.INIT('h8)
	) name2399 (
		\u7_mem_reg[0][28]/NET0131 ,
		_w2987_,
		_w4545_
	);
	LUT2 #(
		.INIT('h2)
	) name2400 (
		\u7_rp_reg[0]/P0001 ,
		_w4542_,
		_w4546_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		_w4543_,
		_w4544_,
		_w4547_
	);
	LUT2 #(
		.INIT('h4)
	) name2402 (
		_w4545_,
		_w4547_,
		_w4548_
	);
	LUT2 #(
		.INIT('h8)
	) name2403 (
		_w4546_,
		_w4548_,
		_w4549_
	);
	LUT2 #(
		.INIT('h2)
	) name2404 (
		_w2805_,
		_w4541_,
		_w4550_
	);
	LUT2 #(
		.INIT('h4)
	) name2405 (
		_w4549_,
		_w4550_,
		_w4551_
	);
	LUT2 #(
		.INIT('h8)
	) name2406 (
		\u7_mem_reg[3][16]/NET0131 ,
		_w2981_,
		_w4552_
	);
	LUT2 #(
		.INIT('h8)
	) name2407 (
		\u7_mem_reg[2][16]/NET0131 ,
		_w2983_,
		_w4553_
	);
	LUT2 #(
		.INIT('h8)
	) name2408 (
		\u7_mem_reg[1][16]/NET0131 ,
		_w2985_,
		_w4554_
	);
	LUT2 #(
		.INIT('h8)
	) name2409 (
		\u7_mem_reg[0][16]/NET0131 ,
		_w2987_,
		_w4555_
	);
	LUT2 #(
		.INIT('h1)
	) name2410 (
		_w4552_,
		_w4553_,
		_w4556_
	);
	LUT2 #(
		.INIT('h1)
	) name2411 (
		_w4554_,
		_w4555_,
		_w4557_
	);
	LUT2 #(
		.INIT('h8)
	) name2412 (
		_w4556_,
		_w4557_,
		_w4558_
	);
	LUT2 #(
		.INIT('h2)
	) name2413 (
		_w2992_,
		_w4558_,
		_w4559_
	);
	LUT2 #(
		.INIT('h2)
	) name2414 (
		_w4352_,
		_w4507_,
		_w4560_
	);
	LUT2 #(
		.INIT('h2)
	) name2415 (
		_w2808_,
		_w4559_,
		_w4561_
	);
	LUT2 #(
		.INIT('h4)
	) name2416 (
		_w4560_,
		_w4561_,
		_w4562_
	);
	LUT2 #(
		.INIT('h4)
	) name2417 (
		_w4551_,
		_w4562_,
		_w4563_
	);
	LUT2 #(
		.INIT('h2)
	) name2418 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4540_,
		_w4564_
	);
	LUT2 #(
		.INIT('h4)
	) name2419 (
		_w4563_,
		_w4564_,
		_w4565_
	);
	LUT2 #(
		.INIT('h1)
	) name2420 (
		\u7_dout_reg[17]/P0001 ,
		_w2808_,
		_w4566_
	);
	LUT2 #(
		.INIT('h4)
	) name2421 (
		\u7_rp_reg[0]/P0001 ,
		_w4471_,
		_w4567_
	);
	LUT2 #(
		.INIT('h8)
	) name2422 (
		\u7_mem_reg[2][29]/NET0131 ,
		_w2983_,
		_w4568_
	);
	LUT2 #(
		.INIT('h8)
	) name2423 (
		\u7_mem_reg[3][29]/NET0131 ,
		_w2981_,
		_w4569_
	);
	LUT2 #(
		.INIT('h8)
	) name2424 (
		\u7_mem_reg[1][29]/NET0131 ,
		_w2985_,
		_w4570_
	);
	LUT2 #(
		.INIT('h8)
	) name2425 (
		\u7_mem_reg[0][29]/NET0131 ,
		_w2987_,
		_w4571_
	);
	LUT2 #(
		.INIT('h2)
	) name2426 (
		\u7_rp_reg[0]/P0001 ,
		_w4568_,
		_w4572_
	);
	LUT2 #(
		.INIT('h1)
	) name2427 (
		_w4569_,
		_w4570_,
		_w4573_
	);
	LUT2 #(
		.INIT('h4)
	) name2428 (
		_w4571_,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h8)
	) name2429 (
		_w4572_,
		_w4574_,
		_w4575_
	);
	LUT2 #(
		.INIT('h2)
	) name2430 (
		_w2805_,
		_w4567_,
		_w4576_
	);
	LUT2 #(
		.INIT('h4)
	) name2431 (
		_w4575_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h8)
	) name2432 (
		\u7_mem_reg[1][17]/NET0131 ,
		_w2985_,
		_w4578_
	);
	LUT2 #(
		.INIT('h8)
	) name2433 (
		\u7_mem_reg[3][17]/NET0131 ,
		_w2981_,
		_w4579_
	);
	LUT2 #(
		.INIT('h8)
	) name2434 (
		\u7_mem_reg[2][17]/NET0131 ,
		_w2983_,
		_w4580_
	);
	LUT2 #(
		.INIT('h8)
	) name2435 (
		\u7_mem_reg[0][17]/NET0131 ,
		_w2987_,
		_w4581_
	);
	LUT2 #(
		.INIT('h1)
	) name2436 (
		_w4578_,
		_w4579_,
		_w4582_
	);
	LUT2 #(
		.INIT('h1)
	) name2437 (
		_w4580_,
		_w4581_,
		_w4583_
	);
	LUT2 #(
		.INIT('h8)
	) name2438 (
		_w4582_,
		_w4583_,
		_w4584_
	);
	LUT2 #(
		.INIT('h2)
	) name2439 (
		_w2992_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h2)
	) name2440 (
		_w4352_,
		_w4532_,
		_w4586_
	);
	LUT2 #(
		.INIT('h2)
	) name2441 (
		_w2808_,
		_w4585_,
		_w4587_
	);
	LUT2 #(
		.INIT('h4)
	) name2442 (
		_w4586_,
		_w4587_,
		_w4588_
	);
	LUT2 #(
		.INIT('h4)
	) name2443 (
		_w4577_,
		_w4588_,
		_w4589_
	);
	LUT2 #(
		.INIT('h2)
	) name2444 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4566_,
		_w4590_
	);
	LUT2 #(
		.INIT('h4)
	) name2445 (
		_w4589_,
		_w4590_,
		_w4591_
	);
	LUT2 #(
		.INIT('h1)
	) name2446 (
		\u7_dout_reg[18]/P0001 ,
		_w2808_,
		_w4592_
	);
	LUT2 #(
		.INIT('h4)
	) name2447 (
		\u7_rp_reg[0]/P0001 ,
		_w4507_,
		_w4593_
	);
	LUT2 #(
		.INIT('h8)
	) name2448 (
		\u7_mem_reg[2][30]/NET0131 ,
		_w2983_,
		_w4594_
	);
	LUT2 #(
		.INIT('h8)
	) name2449 (
		\u7_mem_reg[3][30]/NET0131 ,
		_w2981_,
		_w4595_
	);
	LUT2 #(
		.INIT('h8)
	) name2450 (
		\u7_mem_reg[1][30]/NET0131 ,
		_w2985_,
		_w4596_
	);
	LUT2 #(
		.INIT('h8)
	) name2451 (
		\u7_mem_reg[0][30]/NET0131 ,
		_w2987_,
		_w4597_
	);
	LUT2 #(
		.INIT('h2)
	) name2452 (
		\u7_rp_reg[0]/P0001 ,
		_w4594_,
		_w4598_
	);
	LUT2 #(
		.INIT('h1)
	) name2453 (
		_w4595_,
		_w4596_,
		_w4599_
	);
	LUT2 #(
		.INIT('h4)
	) name2454 (
		_w4597_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h8)
	) name2455 (
		_w4598_,
		_w4600_,
		_w4601_
	);
	LUT2 #(
		.INIT('h2)
	) name2456 (
		_w2805_,
		_w4593_,
		_w4602_
	);
	LUT2 #(
		.INIT('h4)
	) name2457 (
		_w4601_,
		_w4602_,
		_w4603_
	);
	LUT2 #(
		.INIT('h8)
	) name2458 (
		\u7_mem_reg[2][18]/NET0131 ,
		_w2983_,
		_w4604_
	);
	LUT2 #(
		.INIT('h8)
	) name2459 (
		\u7_mem_reg[1][18]/NET0131 ,
		_w2985_,
		_w4605_
	);
	LUT2 #(
		.INIT('h8)
	) name2460 (
		\u7_mem_reg[3][18]/NET0131 ,
		_w2981_,
		_w4606_
	);
	LUT2 #(
		.INIT('h8)
	) name2461 (
		\u7_mem_reg[0][18]/NET0131 ,
		_w2987_,
		_w4607_
	);
	LUT2 #(
		.INIT('h1)
	) name2462 (
		_w4604_,
		_w4605_,
		_w4608_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		_w4606_,
		_w4607_,
		_w4609_
	);
	LUT2 #(
		.INIT('h8)
	) name2464 (
		_w4608_,
		_w4609_,
		_w4610_
	);
	LUT2 #(
		.INIT('h2)
	) name2465 (
		_w2992_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h2)
	) name2466 (
		_w4352_,
		_w4558_,
		_w4612_
	);
	LUT2 #(
		.INIT('h2)
	) name2467 (
		_w2808_,
		_w4611_,
		_w4613_
	);
	LUT2 #(
		.INIT('h4)
	) name2468 (
		_w4612_,
		_w4613_,
		_w4614_
	);
	LUT2 #(
		.INIT('h4)
	) name2469 (
		_w4603_,
		_w4614_,
		_w4615_
	);
	LUT2 #(
		.INIT('h2)
	) name2470 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4592_,
		_w4616_
	);
	LUT2 #(
		.INIT('h4)
	) name2471 (
		_w4615_,
		_w4616_,
		_w4617_
	);
	LUT2 #(
		.INIT('h1)
	) name2472 (
		\u7_dout_reg[19]/P0001 ,
		_w2808_,
		_w4618_
	);
	LUT2 #(
		.INIT('h4)
	) name2473 (
		\u7_rp_reg[0]/P0001 ,
		_w4532_,
		_w4619_
	);
	LUT2 #(
		.INIT('h8)
	) name2474 (
		\u7_mem_reg[2][31]/NET0131 ,
		_w2983_,
		_w4620_
	);
	LUT2 #(
		.INIT('h8)
	) name2475 (
		\u7_mem_reg[3][31]/NET0131 ,
		_w2981_,
		_w4621_
	);
	LUT2 #(
		.INIT('h8)
	) name2476 (
		\u7_mem_reg[1][31]/NET0131 ,
		_w2985_,
		_w4622_
	);
	LUT2 #(
		.INIT('h8)
	) name2477 (
		\u7_mem_reg[0][31]/NET0131 ,
		_w2987_,
		_w4623_
	);
	LUT2 #(
		.INIT('h2)
	) name2478 (
		\u7_rp_reg[0]/P0001 ,
		_w4620_,
		_w4624_
	);
	LUT2 #(
		.INIT('h1)
	) name2479 (
		_w4621_,
		_w4622_,
		_w4625_
	);
	LUT2 #(
		.INIT('h4)
	) name2480 (
		_w4623_,
		_w4625_,
		_w4626_
	);
	LUT2 #(
		.INIT('h8)
	) name2481 (
		_w4624_,
		_w4626_,
		_w4627_
	);
	LUT2 #(
		.INIT('h2)
	) name2482 (
		_w2805_,
		_w4619_,
		_w4628_
	);
	LUT2 #(
		.INIT('h4)
	) name2483 (
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT2 #(
		.INIT('h8)
	) name2484 (
		\u7_mem_reg[3][19]/NET0131 ,
		_w2981_,
		_w4630_
	);
	LUT2 #(
		.INIT('h8)
	) name2485 (
		\u7_mem_reg[0][19]/NET0131 ,
		_w2987_,
		_w4631_
	);
	LUT2 #(
		.INIT('h8)
	) name2486 (
		\u7_mem_reg[1][19]/NET0131 ,
		_w2985_,
		_w4632_
	);
	LUT2 #(
		.INIT('h8)
	) name2487 (
		\u7_mem_reg[2][19]/NET0131 ,
		_w2983_,
		_w4633_
	);
	LUT2 #(
		.INIT('h1)
	) name2488 (
		_w4630_,
		_w4631_,
		_w4634_
	);
	LUT2 #(
		.INIT('h1)
	) name2489 (
		_w4632_,
		_w4633_,
		_w4635_
	);
	LUT2 #(
		.INIT('h8)
	) name2490 (
		_w4634_,
		_w4635_,
		_w4636_
	);
	LUT2 #(
		.INIT('h2)
	) name2491 (
		_w2992_,
		_w4636_,
		_w4637_
	);
	LUT2 #(
		.INIT('h2)
	) name2492 (
		_w4352_,
		_w4584_,
		_w4638_
	);
	LUT2 #(
		.INIT('h2)
	) name2493 (
		_w2808_,
		_w4637_,
		_w4639_
	);
	LUT2 #(
		.INIT('h4)
	) name2494 (
		_w4638_,
		_w4639_,
		_w4640_
	);
	LUT2 #(
		.INIT('h4)
	) name2495 (
		_w4629_,
		_w4640_,
		_w4641_
	);
	LUT2 #(
		.INIT('h2)
	) name2496 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4618_,
		_w4642_
	);
	LUT2 #(
		.INIT('h4)
	) name2497 (
		_w4641_,
		_w4642_,
		_w4643_
	);
	LUT2 #(
		.INIT('h1)
	) name2498 (
		\u7_dout_reg[2]/P0001 ,
		_w2808_,
		_w4644_
	);
	LUT2 #(
		.INIT('h4)
	) name2499 (
		_w2991_,
		_w4352_,
		_w4645_
	);
	LUT2 #(
		.INIT('h8)
	) name2500 (
		\u7_mem_reg[3][2]/NET0131 ,
		_w2981_,
		_w4646_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		\u7_mem_reg[2][2]/NET0131 ,
		_w2983_,
		_w4647_
	);
	LUT2 #(
		.INIT('h8)
	) name2502 (
		\u7_mem_reg[1][2]/NET0131 ,
		_w2985_,
		_w4648_
	);
	LUT2 #(
		.INIT('h8)
	) name2503 (
		\u7_mem_reg[0][2]/NET0131 ,
		_w2987_,
		_w4649_
	);
	LUT2 #(
		.INIT('h1)
	) name2504 (
		_w4646_,
		_w4647_,
		_w4650_
	);
	LUT2 #(
		.INIT('h1)
	) name2505 (
		_w4648_,
		_w4649_,
		_w4651_
	);
	LUT2 #(
		.INIT('h8)
	) name2506 (
		_w4650_,
		_w4651_,
		_w4652_
	);
	LUT2 #(
		.INIT('h2)
	) name2507 (
		_w2992_,
		_w4652_,
		_w4653_
	);
	LUT2 #(
		.INIT('h2)
	) name2508 (
		_w2808_,
		_w4645_,
		_w4654_
	);
	LUT2 #(
		.INIT('h4)
	) name2509 (
		_w4653_,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h2)
	) name2510 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4644_,
		_w4656_
	);
	LUT2 #(
		.INIT('h4)
	) name2511 (
		_w4655_,
		_w4656_,
		_w4657_
	);
	LUT2 #(
		.INIT('h1)
	) name2512 (
		\u7_dout_reg[3]/P0001 ,
		_w2808_,
		_w4658_
	);
	LUT2 #(
		.INIT('h8)
	) name2513 (
		\u7_mem_reg[1][3]/NET0131 ,
		_w2985_,
		_w4659_
	);
	LUT2 #(
		.INIT('h8)
	) name2514 (
		\u7_mem_reg[3][3]/NET0131 ,
		_w2981_,
		_w4660_
	);
	LUT2 #(
		.INIT('h8)
	) name2515 (
		\u7_mem_reg[2][3]/NET0131 ,
		_w2983_,
		_w4661_
	);
	LUT2 #(
		.INIT('h8)
	) name2516 (
		\u7_mem_reg[0][3]/NET0131 ,
		_w2987_,
		_w4662_
	);
	LUT2 #(
		.INIT('h1)
	) name2517 (
		_w4659_,
		_w4660_,
		_w4663_
	);
	LUT2 #(
		.INIT('h1)
	) name2518 (
		_w4661_,
		_w4662_,
		_w4664_
	);
	LUT2 #(
		.INIT('h8)
	) name2519 (
		_w4663_,
		_w4664_,
		_w4665_
	);
	LUT2 #(
		.INIT('h2)
	) name2520 (
		_w2992_,
		_w4665_,
		_w4666_
	);
	LUT2 #(
		.INIT('h4)
	) name2521 (
		_w3004_,
		_w4352_,
		_w4667_
	);
	LUT2 #(
		.INIT('h2)
	) name2522 (
		_w2808_,
		_w4666_,
		_w4668_
	);
	LUT2 #(
		.INIT('h4)
	) name2523 (
		_w4667_,
		_w4668_,
		_w4669_
	);
	LUT2 #(
		.INIT('h2)
	) name2524 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4658_,
		_w4670_
	);
	LUT2 #(
		.INIT('h4)
	) name2525 (
		_w4669_,
		_w4670_,
		_w4671_
	);
	LUT2 #(
		.INIT('h1)
	) name2526 (
		\u7_dout_reg[4]/P0001 ,
		_w2808_,
		_w4672_
	);
	LUT2 #(
		.INIT('h4)
	) name2527 (
		\u7_rp_reg[0]/P0001 ,
		_w2991_,
		_w4673_
	);
	LUT2 #(
		.INIT('h8)
	) name2528 (
		\u7_rp_reg[0]/P0001 ,
		_w4558_,
		_w4674_
	);
	LUT2 #(
		.INIT('h2)
	) name2529 (
		_w2805_,
		_w4673_,
		_w4675_
	);
	LUT2 #(
		.INIT('h4)
	) name2530 (
		_w4674_,
		_w4675_,
		_w4676_
	);
	LUT2 #(
		.INIT('h8)
	) name2531 (
		\u7_mem_reg[1][4]/NET0131 ,
		_w2985_,
		_w4677_
	);
	LUT2 #(
		.INIT('h8)
	) name2532 (
		\u7_mem_reg[2][4]/NET0131 ,
		_w2983_,
		_w4678_
	);
	LUT2 #(
		.INIT('h8)
	) name2533 (
		\u7_mem_reg[3][4]/NET0131 ,
		_w2981_,
		_w4679_
	);
	LUT2 #(
		.INIT('h8)
	) name2534 (
		\u7_mem_reg[0][4]/NET0131 ,
		_w2987_,
		_w4680_
	);
	LUT2 #(
		.INIT('h1)
	) name2535 (
		_w4677_,
		_w4678_,
		_w4681_
	);
	LUT2 #(
		.INIT('h1)
	) name2536 (
		_w4679_,
		_w4680_,
		_w4682_
	);
	LUT2 #(
		.INIT('h8)
	) name2537 (
		_w4681_,
		_w4682_,
		_w4683_
	);
	LUT2 #(
		.INIT('h2)
	) name2538 (
		_w2992_,
		_w4683_,
		_w4684_
	);
	LUT2 #(
		.INIT('h2)
	) name2539 (
		_w4352_,
		_w4652_,
		_w4685_
	);
	LUT2 #(
		.INIT('h2)
	) name2540 (
		_w2808_,
		_w4684_,
		_w4686_
	);
	LUT2 #(
		.INIT('h4)
	) name2541 (
		_w4685_,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('h4)
	) name2542 (
		_w4676_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h2)
	) name2543 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4672_,
		_w4689_
	);
	LUT2 #(
		.INIT('h4)
	) name2544 (
		_w4688_,
		_w4689_,
		_w4690_
	);
	LUT2 #(
		.INIT('h1)
	) name2545 (
		\u7_dout_reg[5]/P0001 ,
		_w2808_,
		_w4691_
	);
	LUT2 #(
		.INIT('h4)
	) name2546 (
		\u7_rp_reg[0]/P0001 ,
		_w3004_,
		_w4692_
	);
	LUT2 #(
		.INIT('h8)
	) name2547 (
		\u7_rp_reg[0]/P0001 ,
		_w4584_,
		_w4693_
	);
	LUT2 #(
		.INIT('h2)
	) name2548 (
		_w2805_,
		_w4692_,
		_w4694_
	);
	LUT2 #(
		.INIT('h4)
	) name2549 (
		_w4693_,
		_w4694_,
		_w4695_
	);
	LUT2 #(
		.INIT('h8)
	) name2550 (
		\u7_mem_reg[3][5]/NET0131 ,
		_w2981_,
		_w4696_
	);
	LUT2 #(
		.INIT('h8)
	) name2551 (
		\u7_mem_reg[0][5]/NET0131 ,
		_w2987_,
		_w4697_
	);
	LUT2 #(
		.INIT('h8)
	) name2552 (
		\u7_mem_reg[2][5]/NET0131 ,
		_w2983_,
		_w4698_
	);
	LUT2 #(
		.INIT('h8)
	) name2553 (
		\u7_mem_reg[1][5]/NET0131 ,
		_w2985_,
		_w4699_
	);
	LUT2 #(
		.INIT('h1)
	) name2554 (
		_w4696_,
		_w4697_,
		_w4700_
	);
	LUT2 #(
		.INIT('h1)
	) name2555 (
		_w4698_,
		_w4699_,
		_w4701_
	);
	LUT2 #(
		.INIT('h8)
	) name2556 (
		_w4700_,
		_w4701_,
		_w4702_
	);
	LUT2 #(
		.INIT('h2)
	) name2557 (
		_w2992_,
		_w4702_,
		_w4703_
	);
	LUT2 #(
		.INIT('h2)
	) name2558 (
		_w4352_,
		_w4665_,
		_w4704_
	);
	LUT2 #(
		.INIT('h2)
	) name2559 (
		_w2808_,
		_w4703_,
		_w4705_
	);
	LUT2 #(
		.INIT('h4)
	) name2560 (
		_w4704_,
		_w4705_,
		_w4706_
	);
	LUT2 #(
		.INIT('h4)
	) name2561 (
		_w4695_,
		_w4706_,
		_w4707_
	);
	LUT2 #(
		.INIT('h2)
	) name2562 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4691_,
		_w4708_
	);
	LUT2 #(
		.INIT('h4)
	) name2563 (
		_w4707_,
		_w4708_,
		_w4709_
	);
	LUT2 #(
		.INIT('h1)
	) name2564 (
		\u7_dout_reg[6]/P0001 ,
		_w2808_,
		_w4710_
	);
	LUT2 #(
		.INIT('h2)
	) name2565 (
		_w2992_,
		_w4350_,
		_w4711_
	);
	LUT2 #(
		.INIT('h2)
	) name2566 (
		_w4352_,
		_w4683_,
		_w4712_
	);
	LUT2 #(
		.INIT('h4)
	) name2567 (
		\u7_rp_reg[0]/P0001 ,
		_w4652_,
		_w4713_
	);
	LUT2 #(
		.INIT('h8)
	) name2568 (
		\u7_rp_reg[0]/P0001 ,
		_w4610_,
		_w4714_
	);
	LUT2 #(
		.INIT('h2)
	) name2569 (
		_w2805_,
		_w4713_,
		_w4715_
	);
	LUT2 #(
		.INIT('h4)
	) name2570 (
		_w4714_,
		_w4715_,
		_w4716_
	);
	LUT2 #(
		.INIT('h2)
	) name2571 (
		_w2808_,
		_w4711_,
		_w4717_
	);
	LUT2 #(
		.INIT('h4)
	) name2572 (
		_w4712_,
		_w4717_,
		_w4718_
	);
	LUT2 #(
		.INIT('h4)
	) name2573 (
		_w4716_,
		_w4718_,
		_w4719_
	);
	LUT2 #(
		.INIT('h2)
	) name2574 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4710_,
		_w4720_
	);
	LUT2 #(
		.INIT('h4)
	) name2575 (
		_w4719_,
		_w4720_,
		_w4721_
	);
	LUT2 #(
		.INIT('h1)
	) name2576 (
		\u7_dout_reg[7]/P0001 ,
		_w2808_,
		_w4722_
	);
	LUT2 #(
		.INIT('h2)
	) name2577 (
		_w2992_,
		_w4399_,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name2578 (
		_w4352_,
		_w4702_,
		_w4724_
	);
	LUT2 #(
		.INIT('h4)
	) name2579 (
		\u7_rp_reg[0]/P0001 ,
		_w4665_,
		_w4725_
	);
	LUT2 #(
		.INIT('h8)
	) name2580 (
		\u7_rp_reg[0]/P0001 ,
		_w4636_,
		_w4726_
	);
	LUT2 #(
		.INIT('h2)
	) name2581 (
		_w2805_,
		_w4725_,
		_w4727_
	);
	LUT2 #(
		.INIT('h4)
	) name2582 (
		_w4726_,
		_w4727_,
		_w4728_
	);
	LUT2 #(
		.INIT('h2)
	) name2583 (
		_w2808_,
		_w4723_,
		_w4729_
	);
	LUT2 #(
		.INIT('h4)
	) name2584 (
		_w4724_,
		_w4729_,
		_w4730_
	);
	LUT2 #(
		.INIT('h4)
	) name2585 (
		_w4728_,
		_w4730_,
		_w4731_
	);
	LUT2 #(
		.INIT('h2)
	) name2586 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4722_,
		_w4732_
	);
	LUT2 #(
		.INIT('h4)
	) name2587 (
		_w4731_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h1)
	) name2588 (
		\u7_dout_reg[8]/P0001 ,
		_w2808_,
		_w4734_
	);
	LUT2 #(
		.INIT('h4)
	) name2589 (
		_w4350_,
		_w4352_,
		_w4735_
	);
	LUT2 #(
		.INIT('h2)
	) name2590 (
		_w2992_,
		_w4359_,
		_w4736_
	);
	LUT2 #(
		.INIT('h4)
	) name2591 (
		\u7_rp_reg[0]/P0001 ,
		_w4683_,
		_w4737_
	);
	LUT2 #(
		.INIT('h8)
	) name2592 (
		\u7_mem_reg[2][20]/NET0131 ,
		_w2983_,
		_w4738_
	);
	LUT2 #(
		.INIT('h8)
	) name2593 (
		\u7_mem_reg[3][20]/NET0131 ,
		_w2981_,
		_w4739_
	);
	LUT2 #(
		.INIT('h8)
	) name2594 (
		\u7_mem_reg[1][20]/NET0131 ,
		_w2985_,
		_w4740_
	);
	LUT2 #(
		.INIT('h8)
	) name2595 (
		\u7_mem_reg[0][20]/NET0131 ,
		_w2987_,
		_w4741_
	);
	LUT2 #(
		.INIT('h2)
	) name2596 (
		\u7_rp_reg[0]/P0001 ,
		_w4738_,
		_w4742_
	);
	LUT2 #(
		.INIT('h1)
	) name2597 (
		_w4739_,
		_w4740_,
		_w4743_
	);
	LUT2 #(
		.INIT('h4)
	) name2598 (
		_w4741_,
		_w4743_,
		_w4744_
	);
	LUT2 #(
		.INIT('h8)
	) name2599 (
		_w4742_,
		_w4744_,
		_w4745_
	);
	LUT2 #(
		.INIT('h2)
	) name2600 (
		_w2805_,
		_w4737_,
		_w4746_
	);
	LUT2 #(
		.INIT('h4)
	) name2601 (
		_w4745_,
		_w4746_,
		_w4747_
	);
	LUT2 #(
		.INIT('h2)
	) name2602 (
		_w2808_,
		_w4735_,
		_w4748_
	);
	LUT2 #(
		.INIT('h4)
	) name2603 (
		_w4736_,
		_w4748_,
		_w4749_
	);
	LUT2 #(
		.INIT('h4)
	) name2604 (
		_w4747_,
		_w4749_,
		_w4750_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4734_,
		_w4751_
	);
	LUT2 #(
		.INIT('h4)
	) name2606 (
		_w4750_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h1)
	) name2607 (
		\u7_dout_reg[9]/P0001 ,
		_w2808_,
		_w4753_
	);
	LUT2 #(
		.INIT('h2)
	) name2608 (
		_w4352_,
		_w4399_,
		_w4754_
	);
	LUT2 #(
		.INIT('h2)
	) name2609 (
		_w2992_,
		_w4415_,
		_w4755_
	);
	LUT2 #(
		.INIT('h4)
	) name2610 (
		\u7_rp_reg[0]/P0001 ,
		_w4702_,
		_w4756_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		\u7_mem_reg[2][21]/NET0131 ,
		_w2983_,
		_w4757_
	);
	LUT2 #(
		.INIT('h8)
	) name2612 (
		\u7_mem_reg[3][21]/NET0131 ,
		_w2981_,
		_w4758_
	);
	LUT2 #(
		.INIT('h8)
	) name2613 (
		\u7_mem_reg[1][21]/NET0131 ,
		_w2985_,
		_w4759_
	);
	LUT2 #(
		.INIT('h8)
	) name2614 (
		\u7_mem_reg[0][21]/NET0131 ,
		_w2987_,
		_w4760_
	);
	LUT2 #(
		.INIT('h2)
	) name2615 (
		\u7_rp_reg[0]/P0001 ,
		_w4757_,
		_w4761_
	);
	LUT2 #(
		.INIT('h1)
	) name2616 (
		_w4758_,
		_w4759_,
		_w4762_
	);
	LUT2 #(
		.INIT('h4)
	) name2617 (
		_w4760_,
		_w4762_,
		_w4763_
	);
	LUT2 #(
		.INIT('h8)
	) name2618 (
		_w4761_,
		_w4763_,
		_w4764_
	);
	LUT2 #(
		.INIT('h2)
	) name2619 (
		_w2805_,
		_w4756_,
		_w4765_
	);
	LUT2 #(
		.INIT('h4)
	) name2620 (
		_w4764_,
		_w4765_,
		_w4766_
	);
	LUT2 #(
		.INIT('h2)
	) name2621 (
		_w2808_,
		_w4754_,
		_w4767_
	);
	LUT2 #(
		.INIT('h4)
	) name2622 (
		_w4755_,
		_w4767_,
		_w4768_
	);
	LUT2 #(
		.INIT('h4)
	) name2623 (
		_w4766_,
		_w4768_,
		_w4769_
	);
	LUT2 #(
		.INIT('h2)
	) name2624 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w4753_,
		_w4770_
	);
	LUT2 #(
		.INIT('h4)
	) name2625 (
		_w4769_,
		_w4770_,
		_w4771_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		\u3_dout_reg[10]/P0001 ,
		_w2787_,
		_w4772_
	);
	LUT2 #(
		.INIT('h8)
	) name2627 (
		\u3_mem_reg[3][6]/NET0131 ,
		_w3009_,
		_w4773_
	);
	LUT2 #(
		.INIT('h8)
	) name2628 (
		\u3_mem_reg[2][6]/NET0131 ,
		_w3011_,
		_w4774_
	);
	LUT2 #(
		.INIT('h8)
	) name2629 (
		\u3_mem_reg[1][6]/NET0131 ,
		_w3013_,
		_w4775_
	);
	LUT2 #(
		.INIT('h8)
	) name2630 (
		\u3_mem_reg[0][6]/NET0131 ,
		_w3015_,
		_w4776_
	);
	LUT2 #(
		.INIT('h1)
	) name2631 (
		_w4773_,
		_w4774_,
		_w4777_
	);
	LUT2 #(
		.INIT('h1)
	) name2632 (
		_w4775_,
		_w4776_,
		_w4778_
	);
	LUT2 #(
		.INIT('h8)
	) name2633 (
		_w4777_,
		_w4778_,
		_w4779_
	);
	LUT2 #(
		.INIT('h4)
	) name2634 (
		\u3_rp_reg[0]/P0001 ,
		_w4779_,
		_w4780_
	);
	LUT2 #(
		.INIT('h8)
	) name2635 (
		\u3_mem_reg[2][22]/NET0131 ,
		_w3011_,
		_w4781_
	);
	LUT2 #(
		.INIT('h8)
	) name2636 (
		\u3_mem_reg[3][22]/NET0131 ,
		_w3009_,
		_w4782_
	);
	LUT2 #(
		.INIT('h8)
	) name2637 (
		\u3_mem_reg[1][22]/NET0131 ,
		_w3013_,
		_w4783_
	);
	LUT2 #(
		.INIT('h8)
	) name2638 (
		\u3_mem_reg[0][22]/NET0131 ,
		_w3015_,
		_w4784_
	);
	LUT2 #(
		.INIT('h2)
	) name2639 (
		\u3_rp_reg[0]/P0001 ,
		_w4781_,
		_w4785_
	);
	LUT2 #(
		.INIT('h1)
	) name2640 (
		_w4782_,
		_w4783_,
		_w4786_
	);
	LUT2 #(
		.INIT('h4)
	) name2641 (
		_w4784_,
		_w4786_,
		_w4787_
	);
	LUT2 #(
		.INIT('h8)
	) name2642 (
		_w4785_,
		_w4787_,
		_w4788_
	);
	LUT2 #(
		.INIT('h2)
	) name2643 (
		_w2784_,
		_w4780_,
		_w4789_
	);
	LUT2 #(
		.INIT('h4)
	) name2644 (
		_w4788_,
		_w4789_,
		_w4790_
	);
	LUT2 #(
		.INIT('h8)
	) name2645 (
		\u3_mem_reg[3][10]/NET0131 ,
		_w3009_,
		_w4791_
	);
	LUT2 #(
		.INIT('h8)
	) name2646 (
		\u3_mem_reg[2][10]/NET0131 ,
		_w3011_,
		_w4792_
	);
	LUT2 #(
		.INIT('h8)
	) name2647 (
		\u3_mem_reg[0][10]/NET0131 ,
		_w3015_,
		_w4793_
	);
	LUT2 #(
		.INIT('h8)
	) name2648 (
		\u3_mem_reg[1][10]/NET0131 ,
		_w3013_,
		_w4794_
	);
	LUT2 #(
		.INIT('h1)
	) name2649 (
		_w4791_,
		_w4792_,
		_w4795_
	);
	LUT2 #(
		.INIT('h1)
	) name2650 (
		_w4793_,
		_w4794_,
		_w4796_
	);
	LUT2 #(
		.INIT('h8)
	) name2651 (
		_w4795_,
		_w4796_,
		_w4797_
	);
	LUT2 #(
		.INIT('h2)
	) name2652 (
		_w3020_,
		_w4797_,
		_w4798_
	);
	LUT2 #(
		.INIT('h2)
	) name2653 (
		\u13_occ0_r_reg[2]/NET0131 ,
		\u13_occ0_r_reg[3]/NET0131 ,
		_w4799_
	);
	LUT2 #(
		.INIT('h8)
	) name2654 (
		\u3_mem_reg[3][8]/NET0131 ,
		_w3009_,
		_w4800_
	);
	LUT2 #(
		.INIT('h8)
	) name2655 (
		\u3_mem_reg[2][8]/NET0131 ,
		_w3011_,
		_w4801_
	);
	LUT2 #(
		.INIT('h8)
	) name2656 (
		\u3_mem_reg[1][8]/NET0131 ,
		_w3013_,
		_w4802_
	);
	LUT2 #(
		.INIT('h8)
	) name2657 (
		\u3_mem_reg[0][8]/NET0131 ,
		_w3015_,
		_w4803_
	);
	LUT2 #(
		.INIT('h1)
	) name2658 (
		_w4800_,
		_w4801_,
		_w4804_
	);
	LUT2 #(
		.INIT('h1)
	) name2659 (
		_w4802_,
		_w4803_,
		_w4805_
	);
	LUT2 #(
		.INIT('h8)
	) name2660 (
		_w4804_,
		_w4805_,
		_w4806_
	);
	LUT2 #(
		.INIT('h2)
	) name2661 (
		_w4799_,
		_w4806_,
		_w4807_
	);
	LUT2 #(
		.INIT('h2)
	) name2662 (
		_w2787_,
		_w4798_,
		_w4808_
	);
	LUT2 #(
		.INIT('h4)
	) name2663 (
		_w4807_,
		_w4808_,
		_w4809_
	);
	LUT2 #(
		.INIT('h4)
	) name2664 (
		_w4790_,
		_w4809_,
		_w4810_
	);
	LUT2 #(
		.INIT('h2)
	) name2665 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w4772_,
		_w4811_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		_w4810_,
		_w4811_,
		_w4812_
	);
	LUT2 #(
		.INIT('h1)
	) name2667 (
		\u3_dout_reg[11]/P0001 ,
		_w2787_,
		_w4813_
	);
	LUT2 #(
		.INIT('h8)
	) name2668 (
		\u3_mem_reg[2][9]/NET0131 ,
		_w3011_,
		_w4814_
	);
	LUT2 #(
		.INIT('h8)
	) name2669 (
		\u3_mem_reg[3][9]/NET0131 ,
		_w3009_,
		_w4815_
	);
	LUT2 #(
		.INIT('h8)
	) name2670 (
		\u3_mem_reg[1][9]/NET0131 ,
		_w3013_,
		_w4816_
	);
	LUT2 #(
		.INIT('h8)
	) name2671 (
		\u3_mem_reg[0][9]/NET0131 ,
		_w3015_,
		_w4817_
	);
	LUT2 #(
		.INIT('h1)
	) name2672 (
		_w4814_,
		_w4815_,
		_w4818_
	);
	LUT2 #(
		.INIT('h1)
	) name2673 (
		_w4816_,
		_w4817_,
		_w4819_
	);
	LUT2 #(
		.INIT('h8)
	) name2674 (
		_w4818_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h2)
	) name2675 (
		_w4799_,
		_w4820_,
		_w4821_
	);
	LUT2 #(
		.INIT('h8)
	) name2676 (
		\u3_mem_reg[3][11]/NET0131 ,
		_w3009_,
		_w4822_
	);
	LUT2 #(
		.INIT('h8)
	) name2677 (
		\u3_mem_reg[2][11]/NET0131 ,
		_w3011_,
		_w4823_
	);
	LUT2 #(
		.INIT('h8)
	) name2678 (
		\u3_mem_reg[0][11]/NET0131 ,
		_w3015_,
		_w4824_
	);
	LUT2 #(
		.INIT('h8)
	) name2679 (
		\u3_mem_reg[1][11]/NET0131 ,
		_w3013_,
		_w4825_
	);
	LUT2 #(
		.INIT('h1)
	) name2680 (
		_w4822_,
		_w4823_,
		_w4826_
	);
	LUT2 #(
		.INIT('h1)
	) name2681 (
		_w4824_,
		_w4825_,
		_w4827_
	);
	LUT2 #(
		.INIT('h8)
	) name2682 (
		_w4826_,
		_w4827_,
		_w4828_
	);
	LUT2 #(
		.INIT('h2)
	) name2683 (
		_w3020_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h8)
	) name2684 (
		\u3_mem_reg[2][7]/NET0131 ,
		_w3011_,
		_w4830_
	);
	LUT2 #(
		.INIT('h8)
	) name2685 (
		\u3_mem_reg[0][7]/NET0131 ,
		_w3015_,
		_w4831_
	);
	LUT2 #(
		.INIT('h8)
	) name2686 (
		\u3_mem_reg[3][7]/NET0131 ,
		_w3009_,
		_w4832_
	);
	LUT2 #(
		.INIT('h8)
	) name2687 (
		\u3_mem_reg[1][7]/NET0131 ,
		_w3013_,
		_w4833_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		_w4830_,
		_w4831_,
		_w4834_
	);
	LUT2 #(
		.INIT('h1)
	) name2689 (
		_w4832_,
		_w4833_,
		_w4835_
	);
	LUT2 #(
		.INIT('h8)
	) name2690 (
		_w4834_,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('h2)
	) name2691 (
		_w2785_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('h8)
	) name2692 (
		\u3_rp_reg[0]/P0001 ,
		_w2784_,
		_w4838_
	);
	LUT2 #(
		.INIT('h8)
	) name2693 (
		\u3_mem_reg[2][23]/NET0131 ,
		_w3011_,
		_w4839_
	);
	LUT2 #(
		.INIT('h8)
	) name2694 (
		\u3_mem_reg[0][23]/NET0131 ,
		_w3015_,
		_w4840_
	);
	LUT2 #(
		.INIT('h8)
	) name2695 (
		\u3_mem_reg[3][23]/NET0131 ,
		_w3009_,
		_w4841_
	);
	LUT2 #(
		.INIT('h8)
	) name2696 (
		\u3_mem_reg[1][23]/NET0131 ,
		_w3013_,
		_w4842_
	);
	LUT2 #(
		.INIT('h1)
	) name2697 (
		_w4839_,
		_w4840_,
		_w4843_
	);
	LUT2 #(
		.INIT('h1)
	) name2698 (
		_w4841_,
		_w4842_,
		_w4844_
	);
	LUT2 #(
		.INIT('h8)
	) name2699 (
		_w4843_,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('h2)
	) name2700 (
		_w4838_,
		_w4845_,
		_w4846_
	);
	LUT2 #(
		.INIT('h2)
	) name2701 (
		_w2787_,
		_w4821_,
		_w4847_
	);
	LUT2 #(
		.INIT('h1)
	) name2702 (
		_w4829_,
		_w4837_,
		_w4848_
	);
	LUT2 #(
		.INIT('h4)
	) name2703 (
		_w4846_,
		_w4848_,
		_w4849_
	);
	LUT2 #(
		.INIT('h8)
	) name2704 (
		_w4847_,
		_w4849_,
		_w4850_
	);
	LUT2 #(
		.INIT('h2)
	) name2705 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w4813_,
		_w4851_
	);
	LUT2 #(
		.INIT('h4)
	) name2706 (
		_w4850_,
		_w4851_,
		_w4852_
	);
	LUT2 #(
		.INIT('h1)
	) name2707 (
		\u3_dout_reg[12]/P0001 ,
		_w2787_,
		_w4853_
	);
	LUT2 #(
		.INIT('h4)
	) name2708 (
		\u3_rp_reg[0]/P0001 ,
		_w4806_,
		_w4854_
	);
	LUT2 #(
		.INIT('h8)
	) name2709 (
		\u3_mem_reg[2][24]/NET0131 ,
		_w3011_,
		_w4855_
	);
	LUT2 #(
		.INIT('h8)
	) name2710 (
		\u3_mem_reg[3][24]/NET0131 ,
		_w3009_,
		_w4856_
	);
	LUT2 #(
		.INIT('h8)
	) name2711 (
		\u3_mem_reg[1][24]/NET0131 ,
		_w3013_,
		_w4857_
	);
	LUT2 #(
		.INIT('h8)
	) name2712 (
		\u3_mem_reg[0][24]/NET0131 ,
		_w3015_,
		_w4858_
	);
	LUT2 #(
		.INIT('h2)
	) name2713 (
		\u3_rp_reg[0]/P0001 ,
		_w4855_,
		_w4859_
	);
	LUT2 #(
		.INIT('h1)
	) name2714 (
		_w4856_,
		_w4857_,
		_w4860_
	);
	LUT2 #(
		.INIT('h4)
	) name2715 (
		_w4858_,
		_w4860_,
		_w4861_
	);
	LUT2 #(
		.INIT('h8)
	) name2716 (
		_w4859_,
		_w4861_,
		_w4862_
	);
	LUT2 #(
		.INIT('h2)
	) name2717 (
		_w2784_,
		_w4854_,
		_w4863_
	);
	LUT2 #(
		.INIT('h4)
	) name2718 (
		_w4862_,
		_w4863_,
		_w4864_
	);
	LUT2 #(
		.INIT('h8)
	) name2719 (
		\u3_mem_reg[2][12]/NET0131 ,
		_w3011_,
		_w4865_
	);
	LUT2 #(
		.INIT('h8)
	) name2720 (
		\u3_mem_reg[3][12]/NET0131 ,
		_w3009_,
		_w4866_
	);
	LUT2 #(
		.INIT('h8)
	) name2721 (
		\u3_mem_reg[1][12]/NET0131 ,
		_w3013_,
		_w4867_
	);
	LUT2 #(
		.INIT('h8)
	) name2722 (
		\u3_mem_reg[0][12]/NET0131 ,
		_w3015_,
		_w4868_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		_w4865_,
		_w4866_,
		_w4869_
	);
	LUT2 #(
		.INIT('h1)
	) name2724 (
		_w4867_,
		_w4868_,
		_w4870_
	);
	LUT2 #(
		.INIT('h8)
	) name2725 (
		_w4869_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('h2)
	) name2726 (
		_w3020_,
		_w4871_,
		_w4872_
	);
	LUT2 #(
		.INIT('h4)
	) name2727 (
		_w4797_,
		_w4799_,
		_w4873_
	);
	LUT2 #(
		.INIT('h2)
	) name2728 (
		_w2787_,
		_w4872_,
		_w4874_
	);
	LUT2 #(
		.INIT('h4)
	) name2729 (
		_w4873_,
		_w4874_,
		_w4875_
	);
	LUT2 #(
		.INIT('h4)
	) name2730 (
		_w4864_,
		_w4875_,
		_w4876_
	);
	LUT2 #(
		.INIT('h2)
	) name2731 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w4853_,
		_w4877_
	);
	LUT2 #(
		.INIT('h4)
	) name2732 (
		_w4876_,
		_w4877_,
		_w4878_
	);
	LUT2 #(
		.INIT('h1)
	) name2733 (
		\u3_dout_reg[13]/P0001 ,
		_w2787_,
		_w4879_
	);
	LUT2 #(
		.INIT('h2)
	) name2734 (
		_w2785_,
		_w4820_,
		_w4880_
	);
	LUT2 #(
		.INIT('h8)
	) name2735 (
		\u3_mem_reg[3][13]/NET0131 ,
		_w3009_,
		_w4881_
	);
	LUT2 #(
		.INIT('h8)
	) name2736 (
		\u3_mem_reg[1][13]/NET0131 ,
		_w3013_,
		_w4882_
	);
	LUT2 #(
		.INIT('h8)
	) name2737 (
		\u3_mem_reg[2][13]/NET0131 ,
		_w3011_,
		_w4883_
	);
	LUT2 #(
		.INIT('h8)
	) name2738 (
		\u3_mem_reg[0][13]/NET0131 ,
		_w3015_,
		_w4884_
	);
	LUT2 #(
		.INIT('h1)
	) name2739 (
		_w4881_,
		_w4882_,
		_w4885_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		_w4883_,
		_w4884_,
		_w4886_
	);
	LUT2 #(
		.INIT('h8)
	) name2741 (
		_w4885_,
		_w4886_,
		_w4887_
	);
	LUT2 #(
		.INIT('h2)
	) name2742 (
		_w3020_,
		_w4887_,
		_w4888_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		\u3_mem_reg[3][25]/NET0131 ,
		_w3009_,
		_w4889_
	);
	LUT2 #(
		.INIT('h8)
	) name2744 (
		\u3_mem_reg[1][25]/NET0131 ,
		_w3013_,
		_w4890_
	);
	LUT2 #(
		.INIT('h8)
	) name2745 (
		\u3_mem_reg[0][25]/NET0131 ,
		_w3015_,
		_w4891_
	);
	LUT2 #(
		.INIT('h8)
	) name2746 (
		\u3_mem_reg[2][25]/NET0131 ,
		_w3011_,
		_w4892_
	);
	LUT2 #(
		.INIT('h1)
	) name2747 (
		_w4889_,
		_w4890_,
		_w4893_
	);
	LUT2 #(
		.INIT('h1)
	) name2748 (
		_w4891_,
		_w4892_,
		_w4894_
	);
	LUT2 #(
		.INIT('h8)
	) name2749 (
		_w4893_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h2)
	) name2750 (
		_w4838_,
		_w4895_,
		_w4896_
	);
	LUT2 #(
		.INIT('h2)
	) name2751 (
		_w4799_,
		_w4828_,
		_w4897_
	);
	LUT2 #(
		.INIT('h2)
	) name2752 (
		_w2787_,
		_w4880_,
		_w4898_
	);
	LUT2 #(
		.INIT('h1)
	) name2753 (
		_w4888_,
		_w4896_,
		_w4899_
	);
	LUT2 #(
		.INIT('h4)
	) name2754 (
		_w4897_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('h8)
	) name2755 (
		_w4898_,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('h2)
	) name2756 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w4879_,
		_w4902_
	);
	LUT2 #(
		.INIT('h4)
	) name2757 (
		_w4901_,
		_w4902_,
		_w4903_
	);
	LUT2 #(
		.INIT('h1)
	) name2758 (
		\u3_dout_reg[14]/P0001 ,
		_w2787_,
		_w4904_
	);
	LUT2 #(
		.INIT('h4)
	) name2759 (
		\u3_rp_reg[0]/P0001 ,
		_w4797_,
		_w4905_
	);
	LUT2 #(
		.INIT('h8)
	) name2760 (
		\u3_mem_reg[2][26]/NET0131 ,
		_w3011_,
		_w4906_
	);
	LUT2 #(
		.INIT('h8)
	) name2761 (
		\u3_mem_reg[3][26]/NET0131 ,
		_w3009_,
		_w4907_
	);
	LUT2 #(
		.INIT('h8)
	) name2762 (
		\u3_mem_reg[1][26]/NET0131 ,
		_w3013_,
		_w4908_
	);
	LUT2 #(
		.INIT('h8)
	) name2763 (
		\u3_mem_reg[0][26]/NET0131 ,
		_w3015_,
		_w4909_
	);
	LUT2 #(
		.INIT('h2)
	) name2764 (
		\u3_rp_reg[0]/P0001 ,
		_w4906_,
		_w4910_
	);
	LUT2 #(
		.INIT('h1)
	) name2765 (
		_w4907_,
		_w4908_,
		_w4911_
	);
	LUT2 #(
		.INIT('h4)
	) name2766 (
		_w4909_,
		_w4911_,
		_w4912_
	);
	LUT2 #(
		.INIT('h8)
	) name2767 (
		_w4910_,
		_w4912_,
		_w4913_
	);
	LUT2 #(
		.INIT('h2)
	) name2768 (
		_w2784_,
		_w4905_,
		_w4914_
	);
	LUT2 #(
		.INIT('h4)
	) name2769 (
		_w4913_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('h8)
	) name2770 (
		\u3_mem_reg[1][14]/NET0131 ,
		_w3013_,
		_w4916_
	);
	LUT2 #(
		.INIT('h8)
	) name2771 (
		\u3_mem_reg[3][14]/NET0131 ,
		_w3009_,
		_w4917_
	);
	LUT2 #(
		.INIT('h8)
	) name2772 (
		\u3_mem_reg[0][14]/NET0131 ,
		_w3015_,
		_w4918_
	);
	LUT2 #(
		.INIT('h8)
	) name2773 (
		\u3_mem_reg[2][14]/NET0131 ,
		_w3011_,
		_w4919_
	);
	LUT2 #(
		.INIT('h1)
	) name2774 (
		_w4916_,
		_w4917_,
		_w4920_
	);
	LUT2 #(
		.INIT('h1)
	) name2775 (
		_w4918_,
		_w4919_,
		_w4921_
	);
	LUT2 #(
		.INIT('h8)
	) name2776 (
		_w4920_,
		_w4921_,
		_w4922_
	);
	LUT2 #(
		.INIT('h2)
	) name2777 (
		_w3020_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h2)
	) name2778 (
		_w4799_,
		_w4871_,
		_w4924_
	);
	LUT2 #(
		.INIT('h2)
	) name2779 (
		_w2787_,
		_w4923_,
		_w4925_
	);
	LUT2 #(
		.INIT('h4)
	) name2780 (
		_w4924_,
		_w4925_,
		_w4926_
	);
	LUT2 #(
		.INIT('h4)
	) name2781 (
		_w4915_,
		_w4926_,
		_w4927_
	);
	LUT2 #(
		.INIT('h2)
	) name2782 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w4904_,
		_w4928_
	);
	LUT2 #(
		.INIT('h4)
	) name2783 (
		_w4927_,
		_w4928_,
		_w4929_
	);
	LUT2 #(
		.INIT('h1)
	) name2784 (
		\u3_dout_reg[15]/P0001 ,
		_w2787_,
		_w4930_
	);
	LUT2 #(
		.INIT('h2)
	) name2785 (
		_w4799_,
		_w4887_,
		_w4931_
	);
	LUT2 #(
		.INIT('h8)
	) name2786 (
		\u3_mem_reg[3][15]/NET0131 ,
		_w3009_,
		_w4932_
	);
	LUT2 #(
		.INIT('h8)
	) name2787 (
		\u3_mem_reg[2][15]/NET0131 ,
		_w3011_,
		_w4933_
	);
	LUT2 #(
		.INIT('h8)
	) name2788 (
		\u3_mem_reg[1][15]/NET0131 ,
		_w3013_,
		_w4934_
	);
	LUT2 #(
		.INIT('h8)
	) name2789 (
		\u3_mem_reg[0][15]/NET0131 ,
		_w3015_,
		_w4935_
	);
	LUT2 #(
		.INIT('h1)
	) name2790 (
		_w4932_,
		_w4933_,
		_w4936_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		_w4934_,
		_w4935_,
		_w4937_
	);
	LUT2 #(
		.INIT('h8)
	) name2792 (
		_w4936_,
		_w4937_,
		_w4938_
	);
	LUT2 #(
		.INIT('h2)
	) name2793 (
		_w3020_,
		_w4938_,
		_w4939_
	);
	LUT2 #(
		.INIT('h4)
	) name2794 (
		\u3_rp_reg[0]/P0001 ,
		_w4828_,
		_w4940_
	);
	LUT2 #(
		.INIT('h8)
	) name2795 (
		\u3_mem_reg[2][27]/NET0131 ,
		_w3011_,
		_w4941_
	);
	LUT2 #(
		.INIT('h8)
	) name2796 (
		\u3_mem_reg[3][27]/NET0131 ,
		_w3009_,
		_w4942_
	);
	LUT2 #(
		.INIT('h8)
	) name2797 (
		\u3_mem_reg[1][27]/NET0131 ,
		_w3013_,
		_w4943_
	);
	LUT2 #(
		.INIT('h8)
	) name2798 (
		\u3_mem_reg[0][27]/NET0131 ,
		_w3015_,
		_w4944_
	);
	LUT2 #(
		.INIT('h2)
	) name2799 (
		\u3_rp_reg[0]/P0001 ,
		_w4941_,
		_w4945_
	);
	LUT2 #(
		.INIT('h1)
	) name2800 (
		_w4942_,
		_w4943_,
		_w4946_
	);
	LUT2 #(
		.INIT('h4)
	) name2801 (
		_w4944_,
		_w4946_,
		_w4947_
	);
	LUT2 #(
		.INIT('h8)
	) name2802 (
		_w4945_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h2)
	) name2803 (
		_w2784_,
		_w4940_,
		_w4949_
	);
	LUT2 #(
		.INIT('h4)
	) name2804 (
		_w4948_,
		_w4949_,
		_w4950_
	);
	LUT2 #(
		.INIT('h2)
	) name2805 (
		_w2787_,
		_w4931_,
		_w4951_
	);
	LUT2 #(
		.INIT('h4)
	) name2806 (
		_w4939_,
		_w4951_,
		_w4952_
	);
	LUT2 #(
		.INIT('h4)
	) name2807 (
		_w4950_,
		_w4952_,
		_w4953_
	);
	LUT2 #(
		.INIT('h2)
	) name2808 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w4930_,
		_w4954_
	);
	LUT2 #(
		.INIT('h4)
	) name2809 (
		_w4953_,
		_w4954_,
		_w4955_
	);
	LUT2 #(
		.INIT('h1)
	) name2810 (
		\u3_dout_reg[16]/P0001 ,
		_w2787_,
		_w4956_
	);
	LUT2 #(
		.INIT('h4)
	) name2811 (
		\u3_rp_reg[0]/P0001 ,
		_w4871_,
		_w4957_
	);
	LUT2 #(
		.INIT('h8)
	) name2812 (
		\u3_mem_reg[2][28]/NET0131 ,
		_w3011_,
		_w4958_
	);
	LUT2 #(
		.INIT('h8)
	) name2813 (
		\u3_mem_reg[3][28]/NET0131 ,
		_w3009_,
		_w4959_
	);
	LUT2 #(
		.INIT('h8)
	) name2814 (
		\u3_mem_reg[1][28]/NET0131 ,
		_w3013_,
		_w4960_
	);
	LUT2 #(
		.INIT('h8)
	) name2815 (
		\u3_mem_reg[0][28]/NET0131 ,
		_w3015_,
		_w4961_
	);
	LUT2 #(
		.INIT('h2)
	) name2816 (
		\u3_rp_reg[0]/P0001 ,
		_w4958_,
		_w4962_
	);
	LUT2 #(
		.INIT('h1)
	) name2817 (
		_w4959_,
		_w4960_,
		_w4963_
	);
	LUT2 #(
		.INIT('h4)
	) name2818 (
		_w4961_,
		_w4963_,
		_w4964_
	);
	LUT2 #(
		.INIT('h8)
	) name2819 (
		_w4962_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h2)
	) name2820 (
		_w2784_,
		_w4957_,
		_w4966_
	);
	LUT2 #(
		.INIT('h4)
	) name2821 (
		_w4965_,
		_w4966_,
		_w4967_
	);
	LUT2 #(
		.INIT('h8)
	) name2822 (
		\u3_mem_reg[3][16]/NET0131 ,
		_w3009_,
		_w4968_
	);
	LUT2 #(
		.INIT('h8)
	) name2823 (
		\u3_mem_reg[2][16]/NET0131 ,
		_w3011_,
		_w4969_
	);
	LUT2 #(
		.INIT('h8)
	) name2824 (
		\u3_mem_reg[1][16]/NET0131 ,
		_w3013_,
		_w4970_
	);
	LUT2 #(
		.INIT('h8)
	) name2825 (
		\u3_mem_reg[0][16]/NET0131 ,
		_w3015_,
		_w4971_
	);
	LUT2 #(
		.INIT('h1)
	) name2826 (
		_w4968_,
		_w4969_,
		_w4972_
	);
	LUT2 #(
		.INIT('h1)
	) name2827 (
		_w4970_,
		_w4971_,
		_w4973_
	);
	LUT2 #(
		.INIT('h8)
	) name2828 (
		_w4972_,
		_w4973_,
		_w4974_
	);
	LUT2 #(
		.INIT('h2)
	) name2829 (
		_w3020_,
		_w4974_,
		_w4975_
	);
	LUT2 #(
		.INIT('h2)
	) name2830 (
		_w4799_,
		_w4922_,
		_w4976_
	);
	LUT2 #(
		.INIT('h2)
	) name2831 (
		_w2787_,
		_w4975_,
		_w4977_
	);
	LUT2 #(
		.INIT('h4)
	) name2832 (
		_w4976_,
		_w4977_,
		_w4978_
	);
	LUT2 #(
		.INIT('h4)
	) name2833 (
		_w4967_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h2)
	) name2834 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w4956_,
		_w4980_
	);
	LUT2 #(
		.INIT('h4)
	) name2835 (
		_w4979_,
		_w4980_,
		_w4981_
	);
	LUT2 #(
		.INIT('h1)
	) name2836 (
		\u3_dout_reg[17]/P0001 ,
		_w2787_,
		_w4982_
	);
	LUT2 #(
		.INIT('h2)
	) name2837 (
		_w4799_,
		_w4938_,
		_w4983_
	);
	LUT2 #(
		.INIT('h2)
	) name2838 (
		_w2785_,
		_w4887_,
		_w4984_
	);
	LUT2 #(
		.INIT('h8)
	) name2839 (
		\u3_mem_reg[3][29]/NET0131 ,
		_w3009_,
		_w4985_
	);
	LUT2 #(
		.INIT('h8)
	) name2840 (
		\u3_mem_reg[0][29]/NET0131 ,
		_w3015_,
		_w4986_
	);
	LUT2 #(
		.INIT('h8)
	) name2841 (
		\u3_mem_reg[2][29]/NET0131 ,
		_w3011_,
		_w4987_
	);
	LUT2 #(
		.INIT('h8)
	) name2842 (
		\u3_mem_reg[1][29]/NET0131 ,
		_w3013_,
		_w4988_
	);
	LUT2 #(
		.INIT('h1)
	) name2843 (
		_w4985_,
		_w4986_,
		_w4989_
	);
	LUT2 #(
		.INIT('h1)
	) name2844 (
		_w4987_,
		_w4988_,
		_w4990_
	);
	LUT2 #(
		.INIT('h8)
	) name2845 (
		_w4989_,
		_w4990_,
		_w4991_
	);
	LUT2 #(
		.INIT('h2)
	) name2846 (
		_w4838_,
		_w4991_,
		_w4992_
	);
	LUT2 #(
		.INIT('h8)
	) name2847 (
		\u3_mem_reg[1][17]/NET0131 ,
		_w3013_,
		_w4993_
	);
	LUT2 #(
		.INIT('h8)
	) name2848 (
		\u3_mem_reg[3][17]/NET0131 ,
		_w3009_,
		_w4994_
	);
	LUT2 #(
		.INIT('h8)
	) name2849 (
		\u3_mem_reg[2][17]/NET0131 ,
		_w3011_,
		_w4995_
	);
	LUT2 #(
		.INIT('h8)
	) name2850 (
		\u3_mem_reg[0][17]/NET0131 ,
		_w3015_,
		_w4996_
	);
	LUT2 #(
		.INIT('h1)
	) name2851 (
		_w4993_,
		_w4994_,
		_w4997_
	);
	LUT2 #(
		.INIT('h1)
	) name2852 (
		_w4995_,
		_w4996_,
		_w4998_
	);
	LUT2 #(
		.INIT('h8)
	) name2853 (
		_w4997_,
		_w4998_,
		_w4999_
	);
	LUT2 #(
		.INIT('h2)
	) name2854 (
		_w3020_,
		_w4999_,
		_w5000_
	);
	LUT2 #(
		.INIT('h2)
	) name2855 (
		_w2787_,
		_w4983_,
		_w5001_
	);
	LUT2 #(
		.INIT('h1)
	) name2856 (
		_w4984_,
		_w4992_,
		_w5002_
	);
	LUT2 #(
		.INIT('h4)
	) name2857 (
		_w5000_,
		_w5002_,
		_w5003_
	);
	LUT2 #(
		.INIT('h8)
	) name2858 (
		_w5001_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h2)
	) name2859 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w4982_,
		_w5005_
	);
	LUT2 #(
		.INIT('h4)
	) name2860 (
		_w5004_,
		_w5005_,
		_w5006_
	);
	LUT2 #(
		.INIT('h1)
	) name2861 (
		\u3_dout_reg[18]/P0001 ,
		_w2787_,
		_w5007_
	);
	LUT2 #(
		.INIT('h4)
	) name2862 (
		\u3_rp_reg[0]/P0001 ,
		_w4922_,
		_w5008_
	);
	LUT2 #(
		.INIT('h8)
	) name2863 (
		\u3_mem_reg[2][30]/NET0131 ,
		_w3011_,
		_w5009_
	);
	LUT2 #(
		.INIT('h8)
	) name2864 (
		\u3_mem_reg[3][30]/NET0131 ,
		_w3009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h8)
	) name2865 (
		\u3_mem_reg[1][30]/NET0131 ,
		_w3013_,
		_w5011_
	);
	LUT2 #(
		.INIT('h8)
	) name2866 (
		\u3_mem_reg[0][30]/NET0131 ,
		_w3015_,
		_w5012_
	);
	LUT2 #(
		.INIT('h2)
	) name2867 (
		\u3_rp_reg[0]/P0001 ,
		_w5009_,
		_w5013_
	);
	LUT2 #(
		.INIT('h1)
	) name2868 (
		_w5010_,
		_w5011_,
		_w5014_
	);
	LUT2 #(
		.INIT('h4)
	) name2869 (
		_w5012_,
		_w5014_,
		_w5015_
	);
	LUT2 #(
		.INIT('h8)
	) name2870 (
		_w5013_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h2)
	) name2871 (
		_w2784_,
		_w5008_,
		_w5017_
	);
	LUT2 #(
		.INIT('h4)
	) name2872 (
		_w5016_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h8)
	) name2873 (
		\u3_mem_reg[1][18]/NET0131 ,
		_w3013_,
		_w5019_
	);
	LUT2 #(
		.INIT('h8)
	) name2874 (
		\u3_mem_reg[3][18]/NET0131 ,
		_w3009_,
		_w5020_
	);
	LUT2 #(
		.INIT('h8)
	) name2875 (
		\u3_mem_reg[2][18]/NET0131 ,
		_w3011_,
		_w5021_
	);
	LUT2 #(
		.INIT('h8)
	) name2876 (
		\u3_mem_reg[0][18]/NET0131 ,
		_w3015_,
		_w5022_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		_w5019_,
		_w5020_,
		_w5023_
	);
	LUT2 #(
		.INIT('h1)
	) name2878 (
		_w5021_,
		_w5022_,
		_w5024_
	);
	LUT2 #(
		.INIT('h8)
	) name2879 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h2)
	) name2880 (
		_w3020_,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h2)
	) name2881 (
		_w4799_,
		_w4974_,
		_w5027_
	);
	LUT2 #(
		.INIT('h2)
	) name2882 (
		_w2787_,
		_w5026_,
		_w5028_
	);
	LUT2 #(
		.INIT('h4)
	) name2883 (
		_w5027_,
		_w5028_,
		_w5029_
	);
	LUT2 #(
		.INIT('h4)
	) name2884 (
		_w5018_,
		_w5029_,
		_w5030_
	);
	LUT2 #(
		.INIT('h2)
	) name2885 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5007_,
		_w5031_
	);
	LUT2 #(
		.INIT('h4)
	) name2886 (
		_w5030_,
		_w5031_,
		_w5032_
	);
	LUT2 #(
		.INIT('h1)
	) name2887 (
		\u8_dout_reg[10]/P0001 ,
		_w2159_,
		_w5033_
	);
	LUT2 #(
		.INIT('h8)
	) name2888 (
		\u8_mem_reg[3][6]/NET0131 ,
		_w2163_,
		_w5034_
	);
	LUT2 #(
		.INIT('h8)
	) name2889 (
		\u8_mem_reg[2][6]/NET0131 ,
		_w3028_,
		_w5035_
	);
	LUT2 #(
		.INIT('h8)
	) name2890 (
		\u8_mem_reg[0][6]/NET0131 ,
		_w3032_,
		_w5036_
	);
	LUT2 #(
		.INIT('h8)
	) name2891 (
		\u8_mem_reg[1][6]/NET0131 ,
		_w3030_,
		_w5037_
	);
	LUT2 #(
		.INIT('h1)
	) name2892 (
		_w5034_,
		_w5035_,
		_w5038_
	);
	LUT2 #(
		.INIT('h1)
	) name2893 (
		_w5036_,
		_w5037_,
		_w5039_
	);
	LUT2 #(
		.INIT('h8)
	) name2894 (
		_w5038_,
		_w5039_,
		_w5040_
	);
	LUT2 #(
		.INIT('h4)
	) name2895 (
		\u8_rp_reg[0]/P0001 ,
		_w5040_,
		_w5041_
	);
	LUT2 #(
		.INIT('h8)
	) name2896 (
		\u8_mem_reg[2][22]/NET0131 ,
		_w3028_,
		_w5042_
	);
	LUT2 #(
		.INIT('h8)
	) name2897 (
		\u8_mem_reg[3][22]/NET0131 ,
		_w2163_,
		_w5043_
	);
	LUT2 #(
		.INIT('h8)
	) name2898 (
		\u8_mem_reg[1][22]/NET0131 ,
		_w3030_,
		_w5044_
	);
	LUT2 #(
		.INIT('h8)
	) name2899 (
		\u8_mem_reg[0][22]/NET0131 ,
		_w3032_,
		_w5045_
	);
	LUT2 #(
		.INIT('h2)
	) name2900 (
		\u8_rp_reg[0]/P0001 ,
		_w5042_,
		_w5046_
	);
	LUT2 #(
		.INIT('h1)
	) name2901 (
		_w5043_,
		_w5044_,
		_w5047_
	);
	LUT2 #(
		.INIT('h4)
	) name2902 (
		_w5045_,
		_w5047_,
		_w5048_
	);
	LUT2 #(
		.INIT('h8)
	) name2903 (
		_w5046_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h2)
	) name2904 (
		_w2160_,
		_w5041_,
		_w5050_
	);
	LUT2 #(
		.INIT('h4)
	) name2905 (
		_w5049_,
		_w5050_,
		_w5051_
	);
	LUT2 #(
		.INIT('h8)
	) name2906 (
		\u8_mem_reg[3][10]/NET0131 ,
		_w2163_,
		_w5052_
	);
	LUT2 #(
		.INIT('h8)
	) name2907 (
		\u8_mem_reg[2][10]/NET0131 ,
		_w3028_,
		_w5053_
	);
	LUT2 #(
		.INIT('h8)
	) name2908 (
		\u8_mem_reg[0][10]/NET0131 ,
		_w3032_,
		_w5054_
	);
	LUT2 #(
		.INIT('h8)
	) name2909 (
		\u8_mem_reg[1][10]/NET0131 ,
		_w3030_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name2910 (
		_w5052_,
		_w5053_,
		_w5056_
	);
	LUT2 #(
		.INIT('h1)
	) name2911 (
		_w5054_,
		_w5055_,
		_w5057_
	);
	LUT2 #(
		.INIT('h8)
	) name2912 (
		_w5056_,
		_w5057_,
		_w5058_
	);
	LUT2 #(
		.INIT('h2)
	) name2913 (
		_w3037_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h2)
	) name2914 (
		\u13_occ1_r_reg[10]/NET0131 ,
		\u13_occ1_r_reg[11]/NET0131 ,
		_w5060_
	);
	LUT2 #(
		.INIT('h8)
	) name2915 (
		\u8_mem_reg[3][8]/NET0131 ,
		_w2163_,
		_w5061_
	);
	LUT2 #(
		.INIT('h8)
	) name2916 (
		\u8_mem_reg[2][8]/NET0131 ,
		_w3028_,
		_w5062_
	);
	LUT2 #(
		.INIT('h8)
	) name2917 (
		\u8_mem_reg[0][8]/NET0131 ,
		_w3032_,
		_w5063_
	);
	LUT2 #(
		.INIT('h8)
	) name2918 (
		\u8_mem_reg[1][8]/NET0131 ,
		_w3030_,
		_w5064_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w5061_,
		_w5062_,
		_w5065_
	);
	LUT2 #(
		.INIT('h1)
	) name2920 (
		_w5063_,
		_w5064_,
		_w5066_
	);
	LUT2 #(
		.INIT('h8)
	) name2921 (
		_w5065_,
		_w5066_,
		_w5067_
	);
	LUT2 #(
		.INIT('h2)
	) name2922 (
		_w5060_,
		_w5067_,
		_w5068_
	);
	LUT2 #(
		.INIT('h2)
	) name2923 (
		_w2159_,
		_w5059_,
		_w5069_
	);
	LUT2 #(
		.INIT('h4)
	) name2924 (
		_w5068_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h4)
	) name2925 (
		_w5051_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h2)
	) name2926 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5033_,
		_w5072_
	);
	LUT2 #(
		.INIT('h4)
	) name2927 (
		_w5071_,
		_w5072_,
		_w5073_
	);
	LUT2 #(
		.INIT('h1)
	) name2928 (
		\u3_dout_reg[19]/P0001 ,
		_w2787_,
		_w5074_
	);
	LUT2 #(
		.INIT('h4)
	) name2929 (
		\u3_rp_reg[0]/P0001 ,
		_w4938_,
		_w5075_
	);
	LUT2 #(
		.INIT('h8)
	) name2930 (
		\u3_mem_reg[2][31]/NET0131 ,
		_w3011_,
		_w5076_
	);
	LUT2 #(
		.INIT('h8)
	) name2931 (
		\u3_mem_reg[3][31]/NET0131 ,
		_w3009_,
		_w5077_
	);
	LUT2 #(
		.INIT('h8)
	) name2932 (
		\u3_mem_reg[1][31]/NET0131 ,
		_w3013_,
		_w5078_
	);
	LUT2 #(
		.INIT('h8)
	) name2933 (
		\u3_mem_reg[0][31]/NET0131 ,
		_w3015_,
		_w5079_
	);
	LUT2 #(
		.INIT('h2)
	) name2934 (
		\u3_rp_reg[0]/P0001 ,
		_w5076_,
		_w5080_
	);
	LUT2 #(
		.INIT('h1)
	) name2935 (
		_w5077_,
		_w5078_,
		_w5081_
	);
	LUT2 #(
		.INIT('h4)
	) name2936 (
		_w5079_,
		_w5081_,
		_w5082_
	);
	LUT2 #(
		.INIT('h8)
	) name2937 (
		_w5080_,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('h2)
	) name2938 (
		_w2784_,
		_w5075_,
		_w5084_
	);
	LUT2 #(
		.INIT('h4)
	) name2939 (
		_w5083_,
		_w5084_,
		_w5085_
	);
	LUT2 #(
		.INIT('h8)
	) name2940 (
		\u3_mem_reg[2][19]/NET0131 ,
		_w3011_,
		_w5086_
	);
	LUT2 #(
		.INIT('h8)
	) name2941 (
		\u3_mem_reg[0][19]/NET0131 ,
		_w3015_,
		_w5087_
	);
	LUT2 #(
		.INIT('h8)
	) name2942 (
		\u3_mem_reg[1][19]/NET0131 ,
		_w3013_,
		_w5088_
	);
	LUT2 #(
		.INIT('h8)
	) name2943 (
		\u3_mem_reg[3][19]/NET0131 ,
		_w3009_,
		_w5089_
	);
	LUT2 #(
		.INIT('h1)
	) name2944 (
		_w5086_,
		_w5087_,
		_w5090_
	);
	LUT2 #(
		.INIT('h1)
	) name2945 (
		_w5088_,
		_w5089_,
		_w5091_
	);
	LUT2 #(
		.INIT('h8)
	) name2946 (
		_w5090_,
		_w5091_,
		_w5092_
	);
	LUT2 #(
		.INIT('h2)
	) name2947 (
		_w3020_,
		_w5092_,
		_w5093_
	);
	LUT2 #(
		.INIT('h2)
	) name2948 (
		_w4799_,
		_w4999_,
		_w5094_
	);
	LUT2 #(
		.INIT('h2)
	) name2949 (
		_w2787_,
		_w5093_,
		_w5095_
	);
	LUT2 #(
		.INIT('h4)
	) name2950 (
		_w5094_,
		_w5095_,
		_w5096_
	);
	LUT2 #(
		.INIT('h4)
	) name2951 (
		_w5085_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h2)
	) name2952 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5074_,
		_w5098_
	);
	LUT2 #(
		.INIT('h4)
	) name2953 (
		_w5097_,
		_w5098_,
		_w5099_
	);
	LUT2 #(
		.INIT('h1)
	) name2954 (
		\u8_dout_reg[11]/P0001 ,
		_w2159_,
		_w5100_
	);
	LUT2 #(
		.INIT('h8)
	) name2955 (
		\u8_mem_reg[3][7]/NET0131 ,
		_w2163_,
		_w5101_
	);
	LUT2 #(
		.INIT('h8)
	) name2956 (
		\u8_mem_reg[2][7]/NET0131 ,
		_w3028_,
		_w5102_
	);
	LUT2 #(
		.INIT('h8)
	) name2957 (
		\u8_mem_reg[0][7]/NET0131 ,
		_w3032_,
		_w5103_
	);
	LUT2 #(
		.INIT('h8)
	) name2958 (
		\u8_mem_reg[1][7]/NET0131 ,
		_w3030_,
		_w5104_
	);
	LUT2 #(
		.INIT('h1)
	) name2959 (
		_w5101_,
		_w5102_,
		_w5105_
	);
	LUT2 #(
		.INIT('h1)
	) name2960 (
		_w5103_,
		_w5104_,
		_w5106_
	);
	LUT2 #(
		.INIT('h8)
	) name2961 (
		_w5105_,
		_w5106_,
		_w5107_
	);
	LUT2 #(
		.INIT('h4)
	) name2962 (
		\u8_rp_reg[0]/P0001 ,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h8)
	) name2963 (
		\u8_mem_reg[2][23]/NET0131 ,
		_w3028_,
		_w5109_
	);
	LUT2 #(
		.INIT('h8)
	) name2964 (
		\u8_mem_reg[3][23]/NET0131 ,
		_w2163_,
		_w5110_
	);
	LUT2 #(
		.INIT('h8)
	) name2965 (
		\u8_mem_reg[1][23]/NET0131 ,
		_w3030_,
		_w5111_
	);
	LUT2 #(
		.INIT('h8)
	) name2966 (
		\u8_mem_reg[0][23]/NET0131 ,
		_w3032_,
		_w5112_
	);
	LUT2 #(
		.INIT('h2)
	) name2967 (
		\u8_rp_reg[0]/P0001 ,
		_w5109_,
		_w5113_
	);
	LUT2 #(
		.INIT('h1)
	) name2968 (
		_w5110_,
		_w5111_,
		_w5114_
	);
	LUT2 #(
		.INIT('h4)
	) name2969 (
		_w5112_,
		_w5114_,
		_w5115_
	);
	LUT2 #(
		.INIT('h8)
	) name2970 (
		_w5113_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('h2)
	) name2971 (
		_w2160_,
		_w5108_,
		_w5117_
	);
	LUT2 #(
		.INIT('h4)
	) name2972 (
		_w5116_,
		_w5117_,
		_w5118_
	);
	LUT2 #(
		.INIT('h8)
	) name2973 (
		\u8_mem_reg[3][11]/NET0131 ,
		_w2163_,
		_w5119_
	);
	LUT2 #(
		.INIT('h8)
	) name2974 (
		\u8_mem_reg[2][11]/NET0131 ,
		_w3028_,
		_w5120_
	);
	LUT2 #(
		.INIT('h8)
	) name2975 (
		\u8_mem_reg[0][11]/NET0131 ,
		_w3032_,
		_w5121_
	);
	LUT2 #(
		.INIT('h8)
	) name2976 (
		\u8_mem_reg[1][11]/NET0131 ,
		_w3030_,
		_w5122_
	);
	LUT2 #(
		.INIT('h1)
	) name2977 (
		_w5119_,
		_w5120_,
		_w5123_
	);
	LUT2 #(
		.INIT('h1)
	) name2978 (
		_w5121_,
		_w5122_,
		_w5124_
	);
	LUT2 #(
		.INIT('h8)
	) name2979 (
		_w5123_,
		_w5124_,
		_w5125_
	);
	LUT2 #(
		.INIT('h2)
	) name2980 (
		_w3037_,
		_w5125_,
		_w5126_
	);
	LUT2 #(
		.INIT('h8)
	) name2981 (
		\u8_mem_reg[3][9]/NET0131 ,
		_w2163_,
		_w5127_
	);
	LUT2 #(
		.INIT('h8)
	) name2982 (
		\u8_mem_reg[1][9]/NET0131 ,
		_w3030_,
		_w5128_
	);
	LUT2 #(
		.INIT('h8)
	) name2983 (
		\u8_mem_reg[0][9]/NET0131 ,
		_w3032_,
		_w5129_
	);
	LUT2 #(
		.INIT('h8)
	) name2984 (
		\u8_mem_reg[2][9]/NET0131 ,
		_w3028_,
		_w5130_
	);
	LUT2 #(
		.INIT('h1)
	) name2985 (
		_w5127_,
		_w5128_,
		_w5131_
	);
	LUT2 #(
		.INIT('h1)
	) name2986 (
		_w5129_,
		_w5130_,
		_w5132_
	);
	LUT2 #(
		.INIT('h8)
	) name2987 (
		_w5131_,
		_w5132_,
		_w5133_
	);
	LUT2 #(
		.INIT('h2)
	) name2988 (
		_w5060_,
		_w5133_,
		_w5134_
	);
	LUT2 #(
		.INIT('h2)
	) name2989 (
		_w2159_,
		_w5126_,
		_w5135_
	);
	LUT2 #(
		.INIT('h4)
	) name2990 (
		_w5134_,
		_w5135_,
		_w5136_
	);
	LUT2 #(
		.INIT('h4)
	) name2991 (
		_w5118_,
		_w5136_,
		_w5137_
	);
	LUT2 #(
		.INIT('h2)
	) name2992 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5100_,
		_w5138_
	);
	LUT2 #(
		.INIT('h4)
	) name2993 (
		_w5137_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h1)
	) name2994 (
		\u8_dout_reg[12]/P0001 ,
		_w2159_,
		_w5140_
	);
	LUT2 #(
		.INIT('h4)
	) name2995 (
		\u8_rp_reg[0]/P0001 ,
		_w5067_,
		_w5141_
	);
	LUT2 #(
		.INIT('h8)
	) name2996 (
		\u8_mem_reg[2][24]/NET0131 ,
		_w3028_,
		_w5142_
	);
	LUT2 #(
		.INIT('h8)
	) name2997 (
		\u8_mem_reg[3][24]/NET0131 ,
		_w2163_,
		_w5143_
	);
	LUT2 #(
		.INIT('h8)
	) name2998 (
		\u8_mem_reg[1][24]/NET0131 ,
		_w3030_,
		_w5144_
	);
	LUT2 #(
		.INIT('h8)
	) name2999 (
		\u8_mem_reg[0][24]/NET0131 ,
		_w3032_,
		_w5145_
	);
	LUT2 #(
		.INIT('h2)
	) name3000 (
		\u8_rp_reg[0]/P0001 ,
		_w5142_,
		_w5146_
	);
	LUT2 #(
		.INIT('h1)
	) name3001 (
		_w5143_,
		_w5144_,
		_w5147_
	);
	LUT2 #(
		.INIT('h4)
	) name3002 (
		_w5145_,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h8)
	) name3003 (
		_w5146_,
		_w5148_,
		_w5149_
	);
	LUT2 #(
		.INIT('h2)
	) name3004 (
		_w2160_,
		_w5141_,
		_w5150_
	);
	LUT2 #(
		.INIT('h4)
	) name3005 (
		_w5149_,
		_w5150_,
		_w5151_
	);
	LUT2 #(
		.INIT('h8)
	) name3006 (
		\u8_mem_reg[3][12]/NET0131 ,
		_w2163_,
		_w5152_
	);
	LUT2 #(
		.INIT('h8)
	) name3007 (
		\u8_mem_reg[1][12]/NET0131 ,
		_w3030_,
		_w5153_
	);
	LUT2 #(
		.INIT('h8)
	) name3008 (
		\u8_mem_reg[0][12]/NET0131 ,
		_w3032_,
		_w5154_
	);
	LUT2 #(
		.INIT('h8)
	) name3009 (
		\u8_mem_reg[2][12]/NET0131 ,
		_w3028_,
		_w5155_
	);
	LUT2 #(
		.INIT('h1)
	) name3010 (
		_w5152_,
		_w5153_,
		_w5156_
	);
	LUT2 #(
		.INIT('h1)
	) name3011 (
		_w5154_,
		_w5155_,
		_w5157_
	);
	LUT2 #(
		.INIT('h8)
	) name3012 (
		_w5156_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h2)
	) name3013 (
		_w3037_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h4)
	) name3014 (
		_w5058_,
		_w5060_,
		_w5160_
	);
	LUT2 #(
		.INIT('h2)
	) name3015 (
		_w2159_,
		_w5159_,
		_w5161_
	);
	LUT2 #(
		.INIT('h4)
	) name3016 (
		_w5160_,
		_w5161_,
		_w5162_
	);
	LUT2 #(
		.INIT('h4)
	) name3017 (
		_w5151_,
		_w5162_,
		_w5163_
	);
	LUT2 #(
		.INIT('h2)
	) name3018 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5140_,
		_w5164_
	);
	LUT2 #(
		.INIT('h4)
	) name3019 (
		_w5163_,
		_w5164_,
		_w5165_
	);
	LUT2 #(
		.INIT('h1)
	) name3020 (
		\u3_dout_reg[2]/P0001 ,
		_w2787_,
		_w5166_
	);
	LUT2 #(
		.INIT('h4)
	) name3021 (
		_w3019_,
		_w4799_,
		_w5167_
	);
	LUT2 #(
		.INIT('h8)
	) name3022 (
		\u3_mem_reg[3][2]/NET0131 ,
		_w3009_,
		_w5168_
	);
	LUT2 #(
		.INIT('h8)
	) name3023 (
		\u3_mem_reg[2][2]/NET0131 ,
		_w3011_,
		_w5169_
	);
	LUT2 #(
		.INIT('h8)
	) name3024 (
		\u3_mem_reg[1][2]/NET0131 ,
		_w3013_,
		_w5170_
	);
	LUT2 #(
		.INIT('h8)
	) name3025 (
		\u3_mem_reg[0][2]/NET0131 ,
		_w3015_,
		_w5171_
	);
	LUT2 #(
		.INIT('h1)
	) name3026 (
		_w5168_,
		_w5169_,
		_w5172_
	);
	LUT2 #(
		.INIT('h1)
	) name3027 (
		_w5170_,
		_w5171_,
		_w5173_
	);
	LUT2 #(
		.INIT('h8)
	) name3028 (
		_w5172_,
		_w5173_,
		_w5174_
	);
	LUT2 #(
		.INIT('h2)
	) name3029 (
		_w3020_,
		_w5174_,
		_w5175_
	);
	LUT2 #(
		.INIT('h2)
	) name3030 (
		_w2787_,
		_w5167_,
		_w5176_
	);
	LUT2 #(
		.INIT('h4)
	) name3031 (
		_w5175_,
		_w5176_,
		_w5177_
	);
	LUT2 #(
		.INIT('h2)
	) name3032 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5166_,
		_w5178_
	);
	LUT2 #(
		.INIT('h4)
	) name3033 (
		_w5177_,
		_w5178_,
		_w5179_
	);
	LUT2 #(
		.INIT('h1)
	) name3034 (
		\u8_dout_reg[13]/P0001 ,
		_w2159_,
		_w5180_
	);
	LUT2 #(
		.INIT('h4)
	) name3035 (
		\u8_rp_reg[0]/P0001 ,
		_w5133_,
		_w5181_
	);
	LUT2 #(
		.INIT('h8)
	) name3036 (
		\u8_mem_reg[2][25]/NET0131 ,
		_w3028_,
		_w5182_
	);
	LUT2 #(
		.INIT('h8)
	) name3037 (
		\u8_mem_reg[3][25]/NET0131 ,
		_w2163_,
		_w5183_
	);
	LUT2 #(
		.INIT('h8)
	) name3038 (
		\u8_mem_reg[1][25]/NET0131 ,
		_w3030_,
		_w5184_
	);
	LUT2 #(
		.INIT('h8)
	) name3039 (
		\u8_mem_reg[0][25]/NET0131 ,
		_w3032_,
		_w5185_
	);
	LUT2 #(
		.INIT('h2)
	) name3040 (
		\u8_rp_reg[0]/P0001 ,
		_w5182_,
		_w5186_
	);
	LUT2 #(
		.INIT('h1)
	) name3041 (
		_w5183_,
		_w5184_,
		_w5187_
	);
	LUT2 #(
		.INIT('h4)
	) name3042 (
		_w5185_,
		_w5187_,
		_w5188_
	);
	LUT2 #(
		.INIT('h8)
	) name3043 (
		_w5186_,
		_w5188_,
		_w5189_
	);
	LUT2 #(
		.INIT('h2)
	) name3044 (
		_w2160_,
		_w5181_,
		_w5190_
	);
	LUT2 #(
		.INIT('h4)
	) name3045 (
		_w5189_,
		_w5190_,
		_w5191_
	);
	LUT2 #(
		.INIT('h8)
	) name3046 (
		\u8_mem_reg[3][13]/NET0131 ,
		_w2163_,
		_w5192_
	);
	LUT2 #(
		.INIT('h8)
	) name3047 (
		\u8_mem_reg[2][13]/NET0131 ,
		_w3028_,
		_w5193_
	);
	LUT2 #(
		.INIT('h8)
	) name3048 (
		\u8_mem_reg[0][13]/NET0131 ,
		_w3032_,
		_w5194_
	);
	LUT2 #(
		.INIT('h8)
	) name3049 (
		\u8_mem_reg[1][13]/NET0131 ,
		_w3030_,
		_w5195_
	);
	LUT2 #(
		.INIT('h1)
	) name3050 (
		_w5192_,
		_w5193_,
		_w5196_
	);
	LUT2 #(
		.INIT('h1)
	) name3051 (
		_w5194_,
		_w5195_,
		_w5197_
	);
	LUT2 #(
		.INIT('h8)
	) name3052 (
		_w5196_,
		_w5197_,
		_w5198_
	);
	LUT2 #(
		.INIT('h2)
	) name3053 (
		_w3037_,
		_w5198_,
		_w5199_
	);
	LUT2 #(
		.INIT('h2)
	) name3054 (
		_w5060_,
		_w5125_,
		_w5200_
	);
	LUT2 #(
		.INIT('h2)
	) name3055 (
		_w2159_,
		_w5199_,
		_w5201_
	);
	LUT2 #(
		.INIT('h4)
	) name3056 (
		_w5200_,
		_w5201_,
		_w5202_
	);
	LUT2 #(
		.INIT('h4)
	) name3057 (
		_w5191_,
		_w5202_,
		_w5203_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5180_,
		_w5204_
	);
	LUT2 #(
		.INIT('h4)
	) name3059 (
		_w5203_,
		_w5204_,
		_w5205_
	);
	LUT2 #(
		.INIT('h1)
	) name3060 (
		\u3_dout_reg[3]/P0001 ,
		_w2787_,
		_w5206_
	);
	LUT2 #(
		.INIT('h4)
	) name3061 (
		_w3049_,
		_w4799_,
		_w5207_
	);
	LUT2 #(
		.INIT('h8)
	) name3062 (
		\u3_mem_reg[1][3]/NET0131 ,
		_w3013_,
		_w5208_
	);
	LUT2 #(
		.INIT('h8)
	) name3063 (
		\u3_mem_reg[3][3]/NET0131 ,
		_w3009_,
		_w5209_
	);
	LUT2 #(
		.INIT('h8)
	) name3064 (
		\u3_mem_reg[2][3]/NET0131 ,
		_w3011_,
		_w5210_
	);
	LUT2 #(
		.INIT('h8)
	) name3065 (
		\u3_mem_reg[0][3]/NET0131 ,
		_w3015_,
		_w5211_
	);
	LUT2 #(
		.INIT('h1)
	) name3066 (
		_w5208_,
		_w5209_,
		_w5212_
	);
	LUT2 #(
		.INIT('h1)
	) name3067 (
		_w5210_,
		_w5211_,
		_w5213_
	);
	LUT2 #(
		.INIT('h8)
	) name3068 (
		_w5212_,
		_w5213_,
		_w5214_
	);
	LUT2 #(
		.INIT('h2)
	) name3069 (
		_w3020_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h2)
	) name3070 (
		_w2787_,
		_w5207_,
		_w5216_
	);
	LUT2 #(
		.INIT('h4)
	) name3071 (
		_w5215_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h2)
	) name3072 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5206_,
		_w5218_
	);
	LUT2 #(
		.INIT('h4)
	) name3073 (
		_w5217_,
		_w5218_,
		_w5219_
	);
	LUT2 #(
		.INIT('h1)
	) name3074 (
		\u8_dout_reg[14]/P0001 ,
		_w2159_,
		_w5220_
	);
	LUT2 #(
		.INIT('h4)
	) name3075 (
		\u8_rp_reg[0]/P0001 ,
		_w5058_,
		_w5221_
	);
	LUT2 #(
		.INIT('h8)
	) name3076 (
		\u8_mem_reg[2][26]/NET0131 ,
		_w3028_,
		_w5222_
	);
	LUT2 #(
		.INIT('h8)
	) name3077 (
		\u8_mem_reg[3][26]/NET0131 ,
		_w2163_,
		_w5223_
	);
	LUT2 #(
		.INIT('h8)
	) name3078 (
		\u8_mem_reg[1][26]/NET0131 ,
		_w3030_,
		_w5224_
	);
	LUT2 #(
		.INIT('h8)
	) name3079 (
		\u8_mem_reg[0][26]/NET0131 ,
		_w3032_,
		_w5225_
	);
	LUT2 #(
		.INIT('h2)
	) name3080 (
		\u8_rp_reg[0]/P0001 ,
		_w5222_,
		_w5226_
	);
	LUT2 #(
		.INIT('h1)
	) name3081 (
		_w5223_,
		_w5224_,
		_w5227_
	);
	LUT2 #(
		.INIT('h4)
	) name3082 (
		_w5225_,
		_w5227_,
		_w5228_
	);
	LUT2 #(
		.INIT('h8)
	) name3083 (
		_w5226_,
		_w5228_,
		_w5229_
	);
	LUT2 #(
		.INIT('h2)
	) name3084 (
		_w2160_,
		_w5221_,
		_w5230_
	);
	LUT2 #(
		.INIT('h4)
	) name3085 (
		_w5229_,
		_w5230_,
		_w5231_
	);
	LUT2 #(
		.INIT('h8)
	) name3086 (
		\u8_mem_reg[3][14]/NET0131 ,
		_w2163_,
		_w5232_
	);
	LUT2 #(
		.INIT('h8)
	) name3087 (
		\u8_mem_reg[2][14]/NET0131 ,
		_w3028_,
		_w5233_
	);
	LUT2 #(
		.INIT('h8)
	) name3088 (
		\u8_mem_reg[0][14]/NET0131 ,
		_w3032_,
		_w5234_
	);
	LUT2 #(
		.INIT('h8)
	) name3089 (
		\u8_mem_reg[1][14]/NET0131 ,
		_w3030_,
		_w5235_
	);
	LUT2 #(
		.INIT('h1)
	) name3090 (
		_w5232_,
		_w5233_,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name3091 (
		_w5234_,
		_w5235_,
		_w5237_
	);
	LUT2 #(
		.INIT('h8)
	) name3092 (
		_w5236_,
		_w5237_,
		_w5238_
	);
	LUT2 #(
		.INIT('h2)
	) name3093 (
		_w3037_,
		_w5238_,
		_w5239_
	);
	LUT2 #(
		.INIT('h2)
	) name3094 (
		_w5060_,
		_w5158_,
		_w5240_
	);
	LUT2 #(
		.INIT('h2)
	) name3095 (
		_w2159_,
		_w5239_,
		_w5241_
	);
	LUT2 #(
		.INIT('h4)
	) name3096 (
		_w5240_,
		_w5241_,
		_w5242_
	);
	LUT2 #(
		.INIT('h4)
	) name3097 (
		_w5231_,
		_w5242_,
		_w5243_
	);
	LUT2 #(
		.INIT('h2)
	) name3098 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5220_,
		_w5244_
	);
	LUT2 #(
		.INIT('h4)
	) name3099 (
		_w5243_,
		_w5244_,
		_w5245_
	);
	LUT2 #(
		.INIT('h1)
	) name3100 (
		\u3_dout_reg[4]/P0001 ,
		_w2787_,
		_w5246_
	);
	LUT2 #(
		.INIT('h4)
	) name3101 (
		\u3_rp_reg[0]/P0001 ,
		_w3019_,
		_w5247_
	);
	LUT2 #(
		.INIT('h8)
	) name3102 (
		\u3_rp_reg[0]/P0001 ,
		_w4974_,
		_w5248_
	);
	LUT2 #(
		.INIT('h2)
	) name3103 (
		_w2784_,
		_w5247_,
		_w5249_
	);
	LUT2 #(
		.INIT('h4)
	) name3104 (
		_w5248_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h8)
	) name3105 (
		\u3_mem_reg[3][4]/NET0131 ,
		_w3009_,
		_w5251_
	);
	LUT2 #(
		.INIT('h8)
	) name3106 (
		\u3_mem_reg[2][4]/NET0131 ,
		_w3011_,
		_w5252_
	);
	LUT2 #(
		.INIT('h8)
	) name3107 (
		\u3_mem_reg[0][4]/NET0131 ,
		_w3015_,
		_w5253_
	);
	LUT2 #(
		.INIT('h8)
	) name3108 (
		\u3_mem_reg[1][4]/NET0131 ,
		_w3013_,
		_w5254_
	);
	LUT2 #(
		.INIT('h1)
	) name3109 (
		_w5251_,
		_w5252_,
		_w5255_
	);
	LUT2 #(
		.INIT('h1)
	) name3110 (
		_w5253_,
		_w5254_,
		_w5256_
	);
	LUT2 #(
		.INIT('h8)
	) name3111 (
		_w5255_,
		_w5256_,
		_w5257_
	);
	LUT2 #(
		.INIT('h2)
	) name3112 (
		_w3020_,
		_w5257_,
		_w5258_
	);
	LUT2 #(
		.INIT('h2)
	) name3113 (
		_w4799_,
		_w5174_,
		_w5259_
	);
	LUT2 #(
		.INIT('h2)
	) name3114 (
		_w2787_,
		_w5258_,
		_w5260_
	);
	LUT2 #(
		.INIT('h4)
	) name3115 (
		_w5259_,
		_w5260_,
		_w5261_
	);
	LUT2 #(
		.INIT('h4)
	) name3116 (
		_w5250_,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('h2)
	) name3117 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5246_,
		_w5263_
	);
	LUT2 #(
		.INIT('h4)
	) name3118 (
		_w5262_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h1)
	) name3119 (
		\u8_dout_reg[15]/P0001 ,
		_w2159_,
		_w5265_
	);
	LUT2 #(
		.INIT('h4)
	) name3120 (
		\u8_rp_reg[0]/P0001 ,
		_w5125_,
		_w5266_
	);
	LUT2 #(
		.INIT('h8)
	) name3121 (
		\u8_mem_reg[2][27]/NET0131 ,
		_w3028_,
		_w5267_
	);
	LUT2 #(
		.INIT('h8)
	) name3122 (
		\u8_mem_reg[3][27]/NET0131 ,
		_w2163_,
		_w5268_
	);
	LUT2 #(
		.INIT('h8)
	) name3123 (
		\u8_mem_reg[1][27]/NET0131 ,
		_w3030_,
		_w5269_
	);
	LUT2 #(
		.INIT('h8)
	) name3124 (
		\u8_mem_reg[0][27]/NET0131 ,
		_w3032_,
		_w5270_
	);
	LUT2 #(
		.INIT('h2)
	) name3125 (
		\u8_rp_reg[0]/P0001 ,
		_w5267_,
		_w5271_
	);
	LUT2 #(
		.INIT('h1)
	) name3126 (
		_w5268_,
		_w5269_,
		_w5272_
	);
	LUT2 #(
		.INIT('h4)
	) name3127 (
		_w5270_,
		_w5272_,
		_w5273_
	);
	LUT2 #(
		.INIT('h8)
	) name3128 (
		_w5271_,
		_w5273_,
		_w5274_
	);
	LUT2 #(
		.INIT('h2)
	) name3129 (
		_w2160_,
		_w5266_,
		_w5275_
	);
	LUT2 #(
		.INIT('h4)
	) name3130 (
		_w5274_,
		_w5275_,
		_w5276_
	);
	LUT2 #(
		.INIT('h8)
	) name3131 (
		\u8_mem_reg[3][15]/NET0131 ,
		_w2163_,
		_w5277_
	);
	LUT2 #(
		.INIT('h8)
	) name3132 (
		\u8_mem_reg[2][15]/NET0131 ,
		_w3028_,
		_w5278_
	);
	LUT2 #(
		.INIT('h8)
	) name3133 (
		\u8_mem_reg[0][15]/NET0131 ,
		_w3032_,
		_w5279_
	);
	LUT2 #(
		.INIT('h8)
	) name3134 (
		\u8_mem_reg[1][15]/NET0131 ,
		_w3030_,
		_w5280_
	);
	LUT2 #(
		.INIT('h1)
	) name3135 (
		_w5277_,
		_w5278_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name3136 (
		_w5279_,
		_w5280_,
		_w5282_
	);
	LUT2 #(
		.INIT('h8)
	) name3137 (
		_w5281_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h2)
	) name3138 (
		_w3037_,
		_w5283_,
		_w5284_
	);
	LUT2 #(
		.INIT('h2)
	) name3139 (
		_w5060_,
		_w5198_,
		_w5285_
	);
	LUT2 #(
		.INIT('h2)
	) name3140 (
		_w2159_,
		_w5284_,
		_w5286_
	);
	LUT2 #(
		.INIT('h4)
	) name3141 (
		_w5285_,
		_w5286_,
		_w5287_
	);
	LUT2 #(
		.INIT('h4)
	) name3142 (
		_w5276_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h2)
	) name3143 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5265_,
		_w5289_
	);
	LUT2 #(
		.INIT('h4)
	) name3144 (
		_w5288_,
		_w5289_,
		_w5290_
	);
	LUT2 #(
		.INIT('h1)
	) name3145 (
		\u3_dout_reg[5]/P0001 ,
		_w2787_,
		_w5291_
	);
	LUT2 #(
		.INIT('h4)
	) name3146 (
		\u3_rp_reg[0]/P0001 ,
		_w3049_,
		_w5292_
	);
	LUT2 #(
		.INIT('h8)
	) name3147 (
		\u3_rp_reg[0]/P0001 ,
		_w4999_,
		_w5293_
	);
	LUT2 #(
		.INIT('h2)
	) name3148 (
		_w2784_,
		_w5292_,
		_w5294_
	);
	LUT2 #(
		.INIT('h4)
	) name3149 (
		_w5293_,
		_w5294_,
		_w5295_
	);
	LUT2 #(
		.INIT('h8)
	) name3150 (
		\u3_mem_reg[3][5]/NET0131 ,
		_w3009_,
		_w5296_
	);
	LUT2 #(
		.INIT('h8)
	) name3151 (
		\u3_mem_reg[2][5]/NET0131 ,
		_w3011_,
		_w5297_
	);
	LUT2 #(
		.INIT('h8)
	) name3152 (
		\u3_mem_reg[1][5]/NET0131 ,
		_w3013_,
		_w5298_
	);
	LUT2 #(
		.INIT('h8)
	) name3153 (
		\u3_mem_reg[0][5]/NET0131 ,
		_w3015_,
		_w5299_
	);
	LUT2 #(
		.INIT('h1)
	) name3154 (
		_w5296_,
		_w5297_,
		_w5300_
	);
	LUT2 #(
		.INIT('h1)
	) name3155 (
		_w5298_,
		_w5299_,
		_w5301_
	);
	LUT2 #(
		.INIT('h8)
	) name3156 (
		_w5300_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h2)
	) name3157 (
		_w3020_,
		_w5302_,
		_w5303_
	);
	LUT2 #(
		.INIT('h2)
	) name3158 (
		_w4799_,
		_w5214_,
		_w5304_
	);
	LUT2 #(
		.INIT('h2)
	) name3159 (
		_w2787_,
		_w5303_,
		_w5305_
	);
	LUT2 #(
		.INIT('h4)
	) name3160 (
		_w5304_,
		_w5305_,
		_w5306_
	);
	LUT2 #(
		.INIT('h4)
	) name3161 (
		_w5295_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('h2)
	) name3162 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5291_,
		_w5308_
	);
	LUT2 #(
		.INIT('h4)
	) name3163 (
		_w5307_,
		_w5308_,
		_w5309_
	);
	LUT2 #(
		.INIT('h1)
	) name3164 (
		\u8_dout_reg[16]/P0001 ,
		_w2159_,
		_w5310_
	);
	LUT2 #(
		.INIT('h4)
	) name3165 (
		\u8_rp_reg[0]/P0001 ,
		_w5158_,
		_w5311_
	);
	LUT2 #(
		.INIT('h8)
	) name3166 (
		\u8_mem_reg[2][28]/NET0131 ,
		_w3028_,
		_w5312_
	);
	LUT2 #(
		.INIT('h8)
	) name3167 (
		\u8_mem_reg[3][28]/NET0131 ,
		_w2163_,
		_w5313_
	);
	LUT2 #(
		.INIT('h8)
	) name3168 (
		\u8_mem_reg[1][28]/NET0131 ,
		_w3030_,
		_w5314_
	);
	LUT2 #(
		.INIT('h8)
	) name3169 (
		\u8_mem_reg[0][28]/NET0131 ,
		_w3032_,
		_w5315_
	);
	LUT2 #(
		.INIT('h2)
	) name3170 (
		\u8_rp_reg[0]/P0001 ,
		_w5312_,
		_w5316_
	);
	LUT2 #(
		.INIT('h1)
	) name3171 (
		_w5313_,
		_w5314_,
		_w5317_
	);
	LUT2 #(
		.INIT('h4)
	) name3172 (
		_w5315_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h8)
	) name3173 (
		_w5316_,
		_w5318_,
		_w5319_
	);
	LUT2 #(
		.INIT('h2)
	) name3174 (
		_w2160_,
		_w5311_,
		_w5320_
	);
	LUT2 #(
		.INIT('h4)
	) name3175 (
		_w5319_,
		_w5320_,
		_w5321_
	);
	LUT2 #(
		.INIT('h8)
	) name3176 (
		\u8_mem_reg[2][16]/NET0131 ,
		_w3028_,
		_w5322_
	);
	LUT2 #(
		.INIT('h8)
	) name3177 (
		\u8_mem_reg[0][16]/NET0131 ,
		_w3032_,
		_w5323_
	);
	LUT2 #(
		.INIT('h8)
	) name3178 (
		\u8_mem_reg[1][16]/NET0131 ,
		_w3030_,
		_w5324_
	);
	LUT2 #(
		.INIT('h8)
	) name3179 (
		\u8_mem_reg[3][16]/NET0131 ,
		_w2163_,
		_w5325_
	);
	LUT2 #(
		.INIT('h1)
	) name3180 (
		_w5322_,
		_w5323_,
		_w5326_
	);
	LUT2 #(
		.INIT('h1)
	) name3181 (
		_w5324_,
		_w5325_,
		_w5327_
	);
	LUT2 #(
		.INIT('h8)
	) name3182 (
		_w5326_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h2)
	) name3183 (
		_w3037_,
		_w5328_,
		_w5329_
	);
	LUT2 #(
		.INIT('h2)
	) name3184 (
		_w5060_,
		_w5238_,
		_w5330_
	);
	LUT2 #(
		.INIT('h2)
	) name3185 (
		_w2159_,
		_w5329_,
		_w5331_
	);
	LUT2 #(
		.INIT('h4)
	) name3186 (
		_w5330_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h4)
	) name3187 (
		_w5321_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h2)
	) name3188 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5310_,
		_w5334_
	);
	LUT2 #(
		.INIT('h4)
	) name3189 (
		_w5333_,
		_w5334_,
		_w5335_
	);
	LUT2 #(
		.INIT('h1)
	) name3190 (
		\u8_dout_reg[17]/P0001 ,
		_w2159_,
		_w5336_
	);
	LUT2 #(
		.INIT('h4)
	) name3191 (
		\u8_rp_reg[0]/P0001 ,
		_w5198_,
		_w5337_
	);
	LUT2 #(
		.INIT('h8)
	) name3192 (
		\u8_mem_reg[2][29]/NET0131 ,
		_w3028_,
		_w5338_
	);
	LUT2 #(
		.INIT('h8)
	) name3193 (
		\u8_mem_reg[3][29]/NET0131 ,
		_w2163_,
		_w5339_
	);
	LUT2 #(
		.INIT('h8)
	) name3194 (
		\u8_mem_reg[1][29]/NET0131 ,
		_w3030_,
		_w5340_
	);
	LUT2 #(
		.INIT('h8)
	) name3195 (
		\u8_mem_reg[0][29]/NET0131 ,
		_w3032_,
		_w5341_
	);
	LUT2 #(
		.INIT('h2)
	) name3196 (
		\u8_rp_reg[0]/P0001 ,
		_w5338_,
		_w5342_
	);
	LUT2 #(
		.INIT('h1)
	) name3197 (
		_w5339_,
		_w5340_,
		_w5343_
	);
	LUT2 #(
		.INIT('h4)
	) name3198 (
		_w5341_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h8)
	) name3199 (
		_w5342_,
		_w5344_,
		_w5345_
	);
	LUT2 #(
		.INIT('h2)
	) name3200 (
		_w2160_,
		_w5337_,
		_w5346_
	);
	LUT2 #(
		.INIT('h4)
	) name3201 (
		_w5345_,
		_w5346_,
		_w5347_
	);
	LUT2 #(
		.INIT('h8)
	) name3202 (
		\u8_mem_reg[3][17]/NET0131 ,
		_w2163_,
		_w5348_
	);
	LUT2 #(
		.INIT('h8)
	) name3203 (
		\u8_mem_reg[2][17]/NET0131 ,
		_w3028_,
		_w5349_
	);
	LUT2 #(
		.INIT('h8)
	) name3204 (
		\u8_mem_reg[0][17]/NET0131 ,
		_w3032_,
		_w5350_
	);
	LUT2 #(
		.INIT('h8)
	) name3205 (
		\u8_mem_reg[1][17]/NET0131 ,
		_w3030_,
		_w5351_
	);
	LUT2 #(
		.INIT('h1)
	) name3206 (
		_w5348_,
		_w5349_,
		_w5352_
	);
	LUT2 #(
		.INIT('h1)
	) name3207 (
		_w5350_,
		_w5351_,
		_w5353_
	);
	LUT2 #(
		.INIT('h8)
	) name3208 (
		_w5352_,
		_w5353_,
		_w5354_
	);
	LUT2 #(
		.INIT('h2)
	) name3209 (
		_w3037_,
		_w5354_,
		_w5355_
	);
	LUT2 #(
		.INIT('h2)
	) name3210 (
		_w5060_,
		_w5283_,
		_w5356_
	);
	LUT2 #(
		.INIT('h2)
	) name3211 (
		_w2159_,
		_w5355_,
		_w5357_
	);
	LUT2 #(
		.INIT('h4)
	) name3212 (
		_w5356_,
		_w5357_,
		_w5358_
	);
	LUT2 #(
		.INIT('h4)
	) name3213 (
		_w5347_,
		_w5358_,
		_w5359_
	);
	LUT2 #(
		.INIT('h2)
	) name3214 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5336_,
		_w5360_
	);
	LUT2 #(
		.INIT('h4)
	) name3215 (
		_w5359_,
		_w5360_,
		_w5361_
	);
	LUT2 #(
		.INIT('h1)
	) name3216 (
		\u3_dout_reg[6]/P0001 ,
		_w2787_,
		_w5362_
	);
	LUT2 #(
		.INIT('h4)
	) name3217 (
		\u3_rp_reg[0]/P0001 ,
		_w5174_,
		_w5363_
	);
	LUT2 #(
		.INIT('h8)
	) name3218 (
		\u3_rp_reg[0]/P0001 ,
		_w5025_,
		_w5364_
	);
	LUT2 #(
		.INIT('h2)
	) name3219 (
		_w2784_,
		_w5363_,
		_w5365_
	);
	LUT2 #(
		.INIT('h4)
	) name3220 (
		_w5364_,
		_w5365_,
		_w5366_
	);
	LUT2 #(
		.INIT('h2)
	) name3221 (
		_w3020_,
		_w4779_,
		_w5367_
	);
	LUT2 #(
		.INIT('h2)
	) name3222 (
		_w4799_,
		_w5257_,
		_w5368_
	);
	LUT2 #(
		.INIT('h2)
	) name3223 (
		_w2787_,
		_w5367_,
		_w5369_
	);
	LUT2 #(
		.INIT('h4)
	) name3224 (
		_w5368_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h4)
	) name3225 (
		_w5366_,
		_w5370_,
		_w5371_
	);
	LUT2 #(
		.INIT('h2)
	) name3226 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5362_,
		_w5372_
	);
	LUT2 #(
		.INIT('h4)
	) name3227 (
		_w5371_,
		_w5372_,
		_w5373_
	);
	LUT2 #(
		.INIT('h1)
	) name3228 (
		\u3_dout_reg[7]/P0001 ,
		_w2787_,
		_w5374_
	);
	LUT2 #(
		.INIT('h4)
	) name3229 (
		\u3_rp_reg[0]/P0001 ,
		_w5214_,
		_w5375_
	);
	LUT2 #(
		.INIT('h8)
	) name3230 (
		\u3_rp_reg[0]/P0001 ,
		_w5092_,
		_w5376_
	);
	LUT2 #(
		.INIT('h2)
	) name3231 (
		_w2784_,
		_w5375_,
		_w5377_
	);
	LUT2 #(
		.INIT('h4)
	) name3232 (
		_w5376_,
		_w5377_,
		_w5378_
	);
	LUT2 #(
		.INIT('h2)
	) name3233 (
		_w3020_,
		_w4836_,
		_w5379_
	);
	LUT2 #(
		.INIT('h2)
	) name3234 (
		_w4799_,
		_w5302_,
		_w5380_
	);
	LUT2 #(
		.INIT('h2)
	) name3235 (
		_w2787_,
		_w5379_,
		_w5381_
	);
	LUT2 #(
		.INIT('h4)
	) name3236 (
		_w5380_,
		_w5381_,
		_w5382_
	);
	LUT2 #(
		.INIT('h4)
	) name3237 (
		_w5378_,
		_w5382_,
		_w5383_
	);
	LUT2 #(
		.INIT('h2)
	) name3238 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5374_,
		_w5384_
	);
	LUT2 #(
		.INIT('h4)
	) name3239 (
		_w5383_,
		_w5384_,
		_w5385_
	);
	LUT2 #(
		.INIT('h1)
	) name3240 (
		\u8_dout_reg[18]/P0001 ,
		_w2159_,
		_w5386_
	);
	LUT2 #(
		.INIT('h4)
	) name3241 (
		\u8_rp_reg[0]/P0001 ,
		_w5238_,
		_w5387_
	);
	LUT2 #(
		.INIT('h8)
	) name3242 (
		\u8_mem_reg[2][30]/NET0131 ,
		_w3028_,
		_w5388_
	);
	LUT2 #(
		.INIT('h8)
	) name3243 (
		\u8_mem_reg[3][30]/NET0131 ,
		_w2163_,
		_w5389_
	);
	LUT2 #(
		.INIT('h8)
	) name3244 (
		\u8_mem_reg[1][30]/NET0131 ,
		_w3030_,
		_w5390_
	);
	LUT2 #(
		.INIT('h8)
	) name3245 (
		\u8_mem_reg[0][30]/NET0131 ,
		_w3032_,
		_w5391_
	);
	LUT2 #(
		.INIT('h2)
	) name3246 (
		\u8_rp_reg[0]/P0001 ,
		_w5388_,
		_w5392_
	);
	LUT2 #(
		.INIT('h1)
	) name3247 (
		_w5389_,
		_w5390_,
		_w5393_
	);
	LUT2 #(
		.INIT('h4)
	) name3248 (
		_w5391_,
		_w5393_,
		_w5394_
	);
	LUT2 #(
		.INIT('h8)
	) name3249 (
		_w5392_,
		_w5394_,
		_w5395_
	);
	LUT2 #(
		.INIT('h2)
	) name3250 (
		_w2160_,
		_w5387_,
		_w5396_
	);
	LUT2 #(
		.INIT('h4)
	) name3251 (
		_w5395_,
		_w5396_,
		_w5397_
	);
	LUT2 #(
		.INIT('h8)
	) name3252 (
		\u8_mem_reg[2][18]/NET0131 ,
		_w3028_,
		_w5398_
	);
	LUT2 #(
		.INIT('h8)
	) name3253 (
		\u8_mem_reg[3][18]/NET0131 ,
		_w2163_,
		_w5399_
	);
	LUT2 #(
		.INIT('h8)
	) name3254 (
		\u8_mem_reg[1][18]/NET0131 ,
		_w3030_,
		_w5400_
	);
	LUT2 #(
		.INIT('h8)
	) name3255 (
		\u8_mem_reg[0][18]/NET0131 ,
		_w3032_,
		_w5401_
	);
	LUT2 #(
		.INIT('h1)
	) name3256 (
		_w5398_,
		_w5399_,
		_w5402_
	);
	LUT2 #(
		.INIT('h1)
	) name3257 (
		_w5400_,
		_w5401_,
		_w5403_
	);
	LUT2 #(
		.INIT('h8)
	) name3258 (
		_w5402_,
		_w5403_,
		_w5404_
	);
	LUT2 #(
		.INIT('h2)
	) name3259 (
		_w3037_,
		_w5404_,
		_w5405_
	);
	LUT2 #(
		.INIT('h2)
	) name3260 (
		_w5060_,
		_w5328_,
		_w5406_
	);
	LUT2 #(
		.INIT('h2)
	) name3261 (
		_w2159_,
		_w5405_,
		_w5407_
	);
	LUT2 #(
		.INIT('h4)
	) name3262 (
		_w5406_,
		_w5407_,
		_w5408_
	);
	LUT2 #(
		.INIT('h4)
	) name3263 (
		_w5397_,
		_w5408_,
		_w5409_
	);
	LUT2 #(
		.INIT('h2)
	) name3264 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5386_,
		_w5410_
	);
	LUT2 #(
		.INIT('h4)
	) name3265 (
		_w5409_,
		_w5410_,
		_w5411_
	);
	LUT2 #(
		.INIT('h1)
	) name3266 (
		\u3_dout_reg[8]/P0001 ,
		_w2787_,
		_w5412_
	);
	LUT2 #(
		.INIT('h4)
	) name3267 (
		\u3_rp_reg[0]/P0001 ,
		_w5257_,
		_w5413_
	);
	LUT2 #(
		.INIT('h8)
	) name3268 (
		\u3_mem_reg[2][20]/NET0131 ,
		_w3011_,
		_w5414_
	);
	LUT2 #(
		.INIT('h8)
	) name3269 (
		\u3_mem_reg[3][20]/NET0131 ,
		_w3009_,
		_w5415_
	);
	LUT2 #(
		.INIT('h8)
	) name3270 (
		\u3_mem_reg[1][20]/NET0131 ,
		_w3013_,
		_w5416_
	);
	LUT2 #(
		.INIT('h8)
	) name3271 (
		\u3_mem_reg[0][20]/NET0131 ,
		_w3015_,
		_w5417_
	);
	LUT2 #(
		.INIT('h2)
	) name3272 (
		\u3_rp_reg[0]/P0001 ,
		_w5414_,
		_w5418_
	);
	LUT2 #(
		.INIT('h1)
	) name3273 (
		_w5415_,
		_w5416_,
		_w5419_
	);
	LUT2 #(
		.INIT('h4)
	) name3274 (
		_w5417_,
		_w5419_,
		_w5420_
	);
	LUT2 #(
		.INIT('h8)
	) name3275 (
		_w5418_,
		_w5420_,
		_w5421_
	);
	LUT2 #(
		.INIT('h2)
	) name3276 (
		_w2784_,
		_w5413_,
		_w5422_
	);
	LUT2 #(
		.INIT('h4)
	) name3277 (
		_w5421_,
		_w5422_,
		_w5423_
	);
	LUT2 #(
		.INIT('h2)
	) name3278 (
		_w3020_,
		_w4806_,
		_w5424_
	);
	LUT2 #(
		.INIT('h4)
	) name3279 (
		_w4779_,
		_w4799_,
		_w5425_
	);
	LUT2 #(
		.INIT('h2)
	) name3280 (
		_w2787_,
		_w5424_,
		_w5426_
	);
	LUT2 #(
		.INIT('h4)
	) name3281 (
		_w5425_,
		_w5426_,
		_w5427_
	);
	LUT2 #(
		.INIT('h4)
	) name3282 (
		_w5423_,
		_w5427_,
		_w5428_
	);
	LUT2 #(
		.INIT('h2)
	) name3283 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5412_,
		_w5429_
	);
	LUT2 #(
		.INIT('h4)
	) name3284 (
		_w5428_,
		_w5429_,
		_w5430_
	);
	LUT2 #(
		.INIT('h1)
	) name3285 (
		\u8_dout_reg[19]/P0001 ,
		_w2159_,
		_w5431_
	);
	LUT2 #(
		.INIT('h4)
	) name3286 (
		\u8_rp_reg[0]/P0001 ,
		_w5283_,
		_w5432_
	);
	LUT2 #(
		.INIT('h8)
	) name3287 (
		\u8_mem_reg[2][31]/NET0131 ,
		_w3028_,
		_w5433_
	);
	LUT2 #(
		.INIT('h8)
	) name3288 (
		\u8_mem_reg[3][31]/NET0131 ,
		_w2163_,
		_w5434_
	);
	LUT2 #(
		.INIT('h8)
	) name3289 (
		\u8_mem_reg[1][31]/NET0131 ,
		_w3030_,
		_w5435_
	);
	LUT2 #(
		.INIT('h8)
	) name3290 (
		\u8_mem_reg[0][31]/NET0131 ,
		_w3032_,
		_w5436_
	);
	LUT2 #(
		.INIT('h2)
	) name3291 (
		\u8_rp_reg[0]/P0001 ,
		_w5433_,
		_w5437_
	);
	LUT2 #(
		.INIT('h1)
	) name3292 (
		_w5434_,
		_w5435_,
		_w5438_
	);
	LUT2 #(
		.INIT('h4)
	) name3293 (
		_w5436_,
		_w5438_,
		_w5439_
	);
	LUT2 #(
		.INIT('h8)
	) name3294 (
		_w5437_,
		_w5439_,
		_w5440_
	);
	LUT2 #(
		.INIT('h2)
	) name3295 (
		_w2160_,
		_w5432_,
		_w5441_
	);
	LUT2 #(
		.INIT('h4)
	) name3296 (
		_w5440_,
		_w5441_,
		_w5442_
	);
	LUT2 #(
		.INIT('h8)
	) name3297 (
		\u8_mem_reg[1][19]/NET0131 ,
		_w3030_,
		_w5443_
	);
	LUT2 #(
		.INIT('h8)
	) name3298 (
		\u8_mem_reg[3][19]/NET0131 ,
		_w2163_,
		_w5444_
	);
	LUT2 #(
		.INIT('h8)
	) name3299 (
		\u8_mem_reg[2][19]/NET0131 ,
		_w3028_,
		_w5445_
	);
	LUT2 #(
		.INIT('h8)
	) name3300 (
		\u8_mem_reg[0][19]/NET0131 ,
		_w3032_,
		_w5446_
	);
	LUT2 #(
		.INIT('h1)
	) name3301 (
		_w5443_,
		_w5444_,
		_w5447_
	);
	LUT2 #(
		.INIT('h1)
	) name3302 (
		_w5445_,
		_w5446_,
		_w5448_
	);
	LUT2 #(
		.INIT('h8)
	) name3303 (
		_w5447_,
		_w5448_,
		_w5449_
	);
	LUT2 #(
		.INIT('h2)
	) name3304 (
		_w3037_,
		_w5449_,
		_w5450_
	);
	LUT2 #(
		.INIT('h2)
	) name3305 (
		_w5060_,
		_w5354_,
		_w5451_
	);
	LUT2 #(
		.INIT('h2)
	) name3306 (
		_w2159_,
		_w5450_,
		_w5452_
	);
	LUT2 #(
		.INIT('h4)
	) name3307 (
		_w5451_,
		_w5452_,
		_w5453_
	);
	LUT2 #(
		.INIT('h4)
	) name3308 (
		_w5442_,
		_w5453_,
		_w5454_
	);
	LUT2 #(
		.INIT('h2)
	) name3309 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5431_,
		_w5455_
	);
	LUT2 #(
		.INIT('h4)
	) name3310 (
		_w5454_,
		_w5455_,
		_w5456_
	);
	LUT2 #(
		.INIT('h1)
	) name3311 (
		\u3_dout_reg[9]/P0001 ,
		_w2787_,
		_w5457_
	);
	LUT2 #(
		.INIT('h2)
	) name3312 (
		_w3020_,
		_w4820_,
		_w5458_
	);
	LUT2 #(
		.INIT('h2)
	) name3313 (
		_w4799_,
		_w4836_,
		_w5459_
	);
	LUT2 #(
		.INIT('h4)
	) name3314 (
		\u3_rp_reg[0]/P0001 ,
		_w5302_,
		_w5460_
	);
	LUT2 #(
		.INIT('h8)
	) name3315 (
		\u3_mem_reg[2][21]/NET0131 ,
		_w3011_,
		_w5461_
	);
	LUT2 #(
		.INIT('h8)
	) name3316 (
		\u3_mem_reg[3][21]/NET0131 ,
		_w3009_,
		_w5462_
	);
	LUT2 #(
		.INIT('h8)
	) name3317 (
		\u3_mem_reg[1][21]/NET0131 ,
		_w3013_,
		_w5463_
	);
	LUT2 #(
		.INIT('h8)
	) name3318 (
		\u3_mem_reg[0][21]/NET0131 ,
		_w3015_,
		_w5464_
	);
	LUT2 #(
		.INIT('h2)
	) name3319 (
		\u3_rp_reg[0]/P0001 ,
		_w5461_,
		_w5465_
	);
	LUT2 #(
		.INIT('h1)
	) name3320 (
		_w5462_,
		_w5463_,
		_w5466_
	);
	LUT2 #(
		.INIT('h4)
	) name3321 (
		_w5464_,
		_w5466_,
		_w5467_
	);
	LUT2 #(
		.INIT('h8)
	) name3322 (
		_w5465_,
		_w5467_,
		_w5468_
	);
	LUT2 #(
		.INIT('h2)
	) name3323 (
		_w2784_,
		_w5460_,
		_w5469_
	);
	LUT2 #(
		.INIT('h4)
	) name3324 (
		_w5468_,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h2)
	) name3325 (
		_w2787_,
		_w5458_,
		_w5471_
	);
	LUT2 #(
		.INIT('h4)
	) name3326 (
		_w5459_,
		_w5471_,
		_w5472_
	);
	LUT2 #(
		.INIT('h4)
	) name3327 (
		_w5470_,
		_w5472_,
		_w5473_
	);
	LUT2 #(
		.INIT('h2)
	) name3328 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w5457_,
		_w5474_
	);
	LUT2 #(
		.INIT('h4)
	) name3329 (
		_w5473_,
		_w5474_,
		_w5475_
	);
	LUT2 #(
		.INIT('h1)
	) name3330 (
		\u8_dout_reg[2]/P0001 ,
		_w2159_,
		_w5476_
	);
	LUT2 #(
		.INIT('h4)
	) name3331 (
		_w3036_,
		_w5060_,
		_w5477_
	);
	LUT2 #(
		.INIT('h8)
	) name3332 (
		\u8_mem_reg[3][2]/NET0131 ,
		_w2163_,
		_w5478_
	);
	LUT2 #(
		.INIT('h8)
	) name3333 (
		\u8_mem_reg[0][2]/NET0131 ,
		_w3032_,
		_w5479_
	);
	LUT2 #(
		.INIT('h8)
	) name3334 (
		\u8_mem_reg[1][2]/NET0131 ,
		_w3030_,
		_w5480_
	);
	LUT2 #(
		.INIT('h8)
	) name3335 (
		\u8_mem_reg[2][2]/NET0131 ,
		_w3028_,
		_w5481_
	);
	LUT2 #(
		.INIT('h1)
	) name3336 (
		_w5478_,
		_w5479_,
		_w5482_
	);
	LUT2 #(
		.INIT('h1)
	) name3337 (
		_w5480_,
		_w5481_,
		_w5483_
	);
	LUT2 #(
		.INIT('h8)
	) name3338 (
		_w5482_,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h2)
	) name3339 (
		_w3037_,
		_w5484_,
		_w5485_
	);
	LUT2 #(
		.INIT('h2)
	) name3340 (
		_w2159_,
		_w5477_,
		_w5486_
	);
	LUT2 #(
		.INIT('h4)
	) name3341 (
		_w5485_,
		_w5486_,
		_w5487_
	);
	LUT2 #(
		.INIT('h2)
	) name3342 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5476_,
		_w5488_
	);
	LUT2 #(
		.INIT('h4)
	) name3343 (
		_w5487_,
		_w5488_,
		_w5489_
	);
	LUT2 #(
		.INIT('h1)
	) name3344 (
		\u8_dout_reg[3]/P0001 ,
		_w2159_,
		_w5490_
	);
	LUT2 #(
		.INIT('h4)
	) name3345 (
		_w3059_,
		_w5060_,
		_w5491_
	);
	LUT2 #(
		.INIT('h8)
	) name3346 (
		\u8_mem_reg[3][3]/NET0131 ,
		_w2163_,
		_w5492_
	);
	LUT2 #(
		.INIT('h8)
	) name3347 (
		\u8_mem_reg[0][3]/NET0131 ,
		_w3032_,
		_w5493_
	);
	LUT2 #(
		.INIT('h8)
	) name3348 (
		\u8_mem_reg[2][3]/NET0131 ,
		_w3028_,
		_w5494_
	);
	LUT2 #(
		.INIT('h8)
	) name3349 (
		\u8_mem_reg[1][3]/NET0131 ,
		_w3030_,
		_w5495_
	);
	LUT2 #(
		.INIT('h1)
	) name3350 (
		_w5492_,
		_w5493_,
		_w5496_
	);
	LUT2 #(
		.INIT('h1)
	) name3351 (
		_w5494_,
		_w5495_,
		_w5497_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		_w5496_,
		_w5497_,
		_w5498_
	);
	LUT2 #(
		.INIT('h2)
	) name3353 (
		_w3037_,
		_w5498_,
		_w5499_
	);
	LUT2 #(
		.INIT('h2)
	) name3354 (
		_w2159_,
		_w5491_,
		_w5500_
	);
	LUT2 #(
		.INIT('h4)
	) name3355 (
		_w5499_,
		_w5500_,
		_w5501_
	);
	LUT2 #(
		.INIT('h2)
	) name3356 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5490_,
		_w5502_
	);
	LUT2 #(
		.INIT('h4)
	) name3357 (
		_w5501_,
		_w5502_,
		_w5503_
	);
	LUT2 #(
		.INIT('h1)
	) name3358 (
		\u8_dout_reg[4]/P0001 ,
		_w2159_,
		_w5504_
	);
	LUT2 #(
		.INIT('h4)
	) name3359 (
		\u8_rp_reg[0]/P0001 ,
		_w3036_,
		_w5505_
	);
	LUT2 #(
		.INIT('h8)
	) name3360 (
		\u8_rp_reg[0]/P0001 ,
		_w5328_,
		_w5506_
	);
	LUT2 #(
		.INIT('h2)
	) name3361 (
		_w2160_,
		_w5505_,
		_w5507_
	);
	LUT2 #(
		.INIT('h4)
	) name3362 (
		_w5506_,
		_w5507_,
		_w5508_
	);
	LUT2 #(
		.INIT('h8)
	) name3363 (
		\u8_mem_reg[3][4]/NET0131 ,
		_w2163_,
		_w5509_
	);
	LUT2 #(
		.INIT('h8)
	) name3364 (
		\u8_mem_reg[2][4]/NET0131 ,
		_w3028_,
		_w5510_
	);
	LUT2 #(
		.INIT('h8)
	) name3365 (
		\u8_mem_reg[0][4]/NET0131 ,
		_w3032_,
		_w5511_
	);
	LUT2 #(
		.INIT('h8)
	) name3366 (
		\u8_mem_reg[1][4]/NET0131 ,
		_w3030_,
		_w5512_
	);
	LUT2 #(
		.INIT('h1)
	) name3367 (
		_w5509_,
		_w5510_,
		_w5513_
	);
	LUT2 #(
		.INIT('h1)
	) name3368 (
		_w5511_,
		_w5512_,
		_w5514_
	);
	LUT2 #(
		.INIT('h8)
	) name3369 (
		_w5513_,
		_w5514_,
		_w5515_
	);
	LUT2 #(
		.INIT('h2)
	) name3370 (
		_w3037_,
		_w5515_,
		_w5516_
	);
	LUT2 #(
		.INIT('h2)
	) name3371 (
		_w5060_,
		_w5484_,
		_w5517_
	);
	LUT2 #(
		.INIT('h2)
	) name3372 (
		_w2159_,
		_w5516_,
		_w5518_
	);
	LUT2 #(
		.INIT('h4)
	) name3373 (
		_w5517_,
		_w5518_,
		_w5519_
	);
	LUT2 #(
		.INIT('h4)
	) name3374 (
		_w5508_,
		_w5519_,
		_w5520_
	);
	LUT2 #(
		.INIT('h2)
	) name3375 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5504_,
		_w5521_
	);
	LUT2 #(
		.INIT('h4)
	) name3376 (
		_w5520_,
		_w5521_,
		_w5522_
	);
	LUT2 #(
		.INIT('h1)
	) name3377 (
		\u8_dout_reg[5]/P0001 ,
		_w2159_,
		_w5523_
	);
	LUT2 #(
		.INIT('h4)
	) name3378 (
		\u8_rp_reg[0]/P0001 ,
		_w3059_,
		_w5524_
	);
	LUT2 #(
		.INIT('h8)
	) name3379 (
		\u8_rp_reg[0]/P0001 ,
		_w5354_,
		_w5525_
	);
	LUT2 #(
		.INIT('h2)
	) name3380 (
		_w2160_,
		_w5524_,
		_w5526_
	);
	LUT2 #(
		.INIT('h4)
	) name3381 (
		_w5525_,
		_w5526_,
		_w5527_
	);
	LUT2 #(
		.INIT('h8)
	) name3382 (
		\u8_mem_reg[3][5]/NET0131 ,
		_w2163_,
		_w5528_
	);
	LUT2 #(
		.INIT('h8)
	) name3383 (
		\u8_mem_reg[2][5]/NET0131 ,
		_w3028_,
		_w5529_
	);
	LUT2 #(
		.INIT('h8)
	) name3384 (
		\u8_mem_reg[1][5]/NET0131 ,
		_w3030_,
		_w5530_
	);
	LUT2 #(
		.INIT('h8)
	) name3385 (
		\u8_mem_reg[0][5]/NET0131 ,
		_w3032_,
		_w5531_
	);
	LUT2 #(
		.INIT('h1)
	) name3386 (
		_w5528_,
		_w5529_,
		_w5532_
	);
	LUT2 #(
		.INIT('h1)
	) name3387 (
		_w5530_,
		_w5531_,
		_w5533_
	);
	LUT2 #(
		.INIT('h8)
	) name3388 (
		_w5532_,
		_w5533_,
		_w5534_
	);
	LUT2 #(
		.INIT('h2)
	) name3389 (
		_w3037_,
		_w5534_,
		_w5535_
	);
	LUT2 #(
		.INIT('h2)
	) name3390 (
		_w5060_,
		_w5498_,
		_w5536_
	);
	LUT2 #(
		.INIT('h2)
	) name3391 (
		_w2159_,
		_w5535_,
		_w5537_
	);
	LUT2 #(
		.INIT('h4)
	) name3392 (
		_w5536_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h4)
	) name3393 (
		_w5527_,
		_w5538_,
		_w5539_
	);
	LUT2 #(
		.INIT('h2)
	) name3394 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5523_,
		_w5540_
	);
	LUT2 #(
		.INIT('h4)
	) name3395 (
		_w5539_,
		_w5540_,
		_w5541_
	);
	LUT2 #(
		.INIT('h1)
	) name3396 (
		\u8_dout_reg[6]/P0001 ,
		_w2159_,
		_w5542_
	);
	LUT2 #(
		.INIT('h4)
	) name3397 (
		\u8_rp_reg[0]/P0001 ,
		_w5484_,
		_w5543_
	);
	LUT2 #(
		.INIT('h8)
	) name3398 (
		\u8_rp_reg[0]/P0001 ,
		_w5404_,
		_w5544_
	);
	LUT2 #(
		.INIT('h2)
	) name3399 (
		_w2160_,
		_w5543_,
		_w5545_
	);
	LUT2 #(
		.INIT('h4)
	) name3400 (
		_w5544_,
		_w5545_,
		_w5546_
	);
	LUT2 #(
		.INIT('h2)
	) name3401 (
		_w3037_,
		_w5040_,
		_w5547_
	);
	LUT2 #(
		.INIT('h2)
	) name3402 (
		_w5060_,
		_w5515_,
		_w5548_
	);
	LUT2 #(
		.INIT('h2)
	) name3403 (
		_w2159_,
		_w5547_,
		_w5549_
	);
	LUT2 #(
		.INIT('h4)
	) name3404 (
		_w5548_,
		_w5549_,
		_w5550_
	);
	LUT2 #(
		.INIT('h4)
	) name3405 (
		_w5546_,
		_w5550_,
		_w5551_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5542_,
		_w5552_
	);
	LUT2 #(
		.INIT('h4)
	) name3407 (
		_w5551_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h1)
	) name3408 (
		\u8_dout_reg[7]/P0001 ,
		_w2159_,
		_w5554_
	);
	LUT2 #(
		.INIT('h4)
	) name3409 (
		\u8_rp_reg[0]/P0001 ,
		_w5498_,
		_w5555_
	);
	LUT2 #(
		.INIT('h8)
	) name3410 (
		\u8_rp_reg[0]/P0001 ,
		_w5449_,
		_w5556_
	);
	LUT2 #(
		.INIT('h2)
	) name3411 (
		_w2160_,
		_w5555_,
		_w5557_
	);
	LUT2 #(
		.INIT('h4)
	) name3412 (
		_w5556_,
		_w5557_,
		_w5558_
	);
	LUT2 #(
		.INIT('h2)
	) name3413 (
		_w3037_,
		_w5107_,
		_w5559_
	);
	LUT2 #(
		.INIT('h2)
	) name3414 (
		_w5060_,
		_w5534_,
		_w5560_
	);
	LUT2 #(
		.INIT('h2)
	) name3415 (
		_w2159_,
		_w5559_,
		_w5561_
	);
	LUT2 #(
		.INIT('h4)
	) name3416 (
		_w5560_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h4)
	) name3417 (
		_w5558_,
		_w5562_,
		_w5563_
	);
	LUT2 #(
		.INIT('h2)
	) name3418 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5554_,
		_w5564_
	);
	LUT2 #(
		.INIT('h4)
	) name3419 (
		_w5563_,
		_w5564_,
		_w5565_
	);
	LUT2 #(
		.INIT('h1)
	) name3420 (
		\u8_dout_reg[8]/P0001 ,
		_w2159_,
		_w5566_
	);
	LUT2 #(
		.INIT('h4)
	) name3421 (
		\u8_rp_reg[0]/P0001 ,
		_w5515_,
		_w5567_
	);
	LUT2 #(
		.INIT('h8)
	) name3422 (
		\u8_mem_reg[2][20]/NET0131 ,
		_w3028_,
		_w5568_
	);
	LUT2 #(
		.INIT('h8)
	) name3423 (
		\u8_mem_reg[3][20]/NET0131 ,
		_w2163_,
		_w5569_
	);
	LUT2 #(
		.INIT('h8)
	) name3424 (
		\u8_mem_reg[1][20]/NET0131 ,
		_w3030_,
		_w5570_
	);
	LUT2 #(
		.INIT('h8)
	) name3425 (
		\u8_mem_reg[0][20]/NET0131 ,
		_w3032_,
		_w5571_
	);
	LUT2 #(
		.INIT('h2)
	) name3426 (
		\u8_rp_reg[0]/P0001 ,
		_w5568_,
		_w5572_
	);
	LUT2 #(
		.INIT('h1)
	) name3427 (
		_w5569_,
		_w5570_,
		_w5573_
	);
	LUT2 #(
		.INIT('h4)
	) name3428 (
		_w5571_,
		_w5573_,
		_w5574_
	);
	LUT2 #(
		.INIT('h8)
	) name3429 (
		_w5572_,
		_w5574_,
		_w5575_
	);
	LUT2 #(
		.INIT('h2)
	) name3430 (
		_w2160_,
		_w5567_,
		_w5576_
	);
	LUT2 #(
		.INIT('h4)
	) name3431 (
		_w5575_,
		_w5576_,
		_w5577_
	);
	LUT2 #(
		.INIT('h2)
	) name3432 (
		_w3037_,
		_w5067_,
		_w5578_
	);
	LUT2 #(
		.INIT('h4)
	) name3433 (
		_w5040_,
		_w5060_,
		_w5579_
	);
	LUT2 #(
		.INIT('h2)
	) name3434 (
		_w2159_,
		_w5578_,
		_w5580_
	);
	LUT2 #(
		.INIT('h4)
	) name3435 (
		_w5579_,
		_w5580_,
		_w5581_
	);
	LUT2 #(
		.INIT('h4)
	) name3436 (
		_w5577_,
		_w5581_,
		_w5582_
	);
	LUT2 #(
		.INIT('h2)
	) name3437 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5566_,
		_w5583_
	);
	LUT2 #(
		.INIT('h4)
	) name3438 (
		_w5582_,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h1)
	) name3439 (
		\u8_dout_reg[9]/P0001 ,
		_w2159_,
		_w5585_
	);
	LUT2 #(
		.INIT('h4)
	) name3440 (
		\u8_rp_reg[0]/P0001 ,
		_w5534_,
		_w5586_
	);
	LUT2 #(
		.INIT('h8)
	) name3441 (
		\u8_mem_reg[2][21]/NET0131 ,
		_w3028_,
		_w5587_
	);
	LUT2 #(
		.INIT('h8)
	) name3442 (
		\u8_mem_reg[3][21]/NET0131 ,
		_w2163_,
		_w5588_
	);
	LUT2 #(
		.INIT('h8)
	) name3443 (
		\u8_mem_reg[1][21]/NET0131 ,
		_w3030_,
		_w5589_
	);
	LUT2 #(
		.INIT('h8)
	) name3444 (
		\u8_mem_reg[0][21]/NET0131 ,
		_w3032_,
		_w5590_
	);
	LUT2 #(
		.INIT('h2)
	) name3445 (
		\u8_rp_reg[0]/P0001 ,
		_w5587_,
		_w5591_
	);
	LUT2 #(
		.INIT('h1)
	) name3446 (
		_w5588_,
		_w5589_,
		_w5592_
	);
	LUT2 #(
		.INIT('h4)
	) name3447 (
		_w5590_,
		_w5592_,
		_w5593_
	);
	LUT2 #(
		.INIT('h8)
	) name3448 (
		_w5591_,
		_w5593_,
		_w5594_
	);
	LUT2 #(
		.INIT('h2)
	) name3449 (
		_w2160_,
		_w5586_,
		_w5595_
	);
	LUT2 #(
		.INIT('h4)
	) name3450 (
		_w5594_,
		_w5595_,
		_w5596_
	);
	LUT2 #(
		.INIT('h2)
	) name3451 (
		_w3037_,
		_w5133_,
		_w5597_
	);
	LUT2 #(
		.INIT('h2)
	) name3452 (
		_w5060_,
		_w5107_,
		_w5598_
	);
	LUT2 #(
		.INIT('h2)
	) name3453 (
		_w2159_,
		_w5597_,
		_w5599_
	);
	LUT2 #(
		.INIT('h4)
	) name3454 (
		_w5598_,
		_w5599_,
		_w5600_
	);
	LUT2 #(
		.INIT('h4)
	) name3455 (
		_w5596_,
		_w5600_,
		_w5601_
	);
	LUT2 #(
		.INIT('h2)
	) name3456 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w5585_,
		_w5602_
	);
	LUT2 #(
		.INIT('h4)
	) name3457 (
		_w5601_,
		_w5602_,
		_w5603_
	);
	LUT2 #(
		.INIT('h1)
	) name3458 (
		\u11_wp_reg[1]/P0001 ,
		_w3066_,
		_w5604_
	);
	LUT2 #(
		.INIT('h2)
	) name3459 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w3067_,
		_w5605_
	);
	LUT2 #(
		.INIT('h4)
	) name3460 (
		_w5604_,
		_w5605_,
		_w5606_
	);
	LUT2 #(
		.INIT('h1)
	) name3461 (
		\u9_wp_reg[1]/P0001 ,
		_w3313_,
		_w5607_
	);
	LUT2 #(
		.INIT('h2)
	) name3462 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w3314_,
		_w5608_
	);
	LUT2 #(
		.INIT('h4)
	) name3463 (
		_w5607_,
		_w5608_,
		_w5609_
	);
	LUT2 #(
		.INIT('h1)
	) name3464 (
		\u10_wp_reg[1]/P0001 ,
		_w3503_,
		_w5610_
	);
	LUT2 #(
		.INIT('h2)
	) name3465 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w3504_,
		_w5611_
	);
	LUT2 #(
		.INIT('h4)
	) name3466 (
		_w5610_,
		_w5611_,
		_w5612_
	);
	LUT2 #(
		.INIT('h1)
	) name3467 (
		\u11_wp_reg[3]/P0001 ,
		_w3068_,
		_w5613_
	);
	LUT2 #(
		.INIT('h8)
	) name3468 (
		\u11_wp_reg[3]/P0001 ,
		_w3068_,
		_w5614_
	);
	LUT2 #(
		.INIT('h2)
	) name3469 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w5613_,
		_w5615_
	);
	LUT2 #(
		.INIT('h4)
	) name3470 (
		_w5614_,
		_w5615_,
		_w5616_
	);
	LUT2 #(
		.INIT('h1)
	) name3471 (
		\u9_wp_reg[3]/P0001 ,
		_w3315_,
		_w5617_
	);
	LUT2 #(
		.INIT('h8)
	) name3472 (
		\u9_wp_reg[3]/P0001 ,
		_w3315_,
		_w5618_
	);
	LUT2 #(
		.INIT('h2)
	) name3473 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w5617_,
		_w5619_
	);
	LUT2 #(
		.INIT('h4)
	) name3474 (
		_w5618_,
		_w5619_,
		_w5620_
	);
	LUT2 #(
		.INIT('h1)
	) name3475 (
		\u10_wp_reg[3]/P0001 ,
		_w3505_,
		_w5621_
	);
	LUT2 #(
		.INIT('h8)
	) name3476 (
		\u10_wp_reg[3]/P0001 ,
		_w3505_,
		_w5622_
	);
	LUT2 #(
		.INIT('h2)
	) name3477 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w5621_,
		_w5623_
	);
	LUT2 #(
		.INIT('h4)
	) name3478 (
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h2)
	) name3479 (
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		_w5625_
	);
	LUT2 #(
		.INIT('h1)
	) name3480 (
		\u26_ps_cnt_reg[2]/NET0131 ,
		\u26_ps_cnt_reg[3]/NET0131 ,
		_w5626_
	);
	LUT2 #(
		.INIT('h8)
	) name3481 (
		\u26_ps_cnt_reg[4]/NET0131 ,
		\u26_ps_cnt_reg[5]/NET0131 ,
		_w5627_
	);
	LUT2 #(
		.INIT('h8)
	) name3482 (
		_w5626_,
		_w5627_,
		_w5628_
	);
	LUT2 #(
		.INIT('h8)
	) name3483 (
		_w5625_,
		_w5628_,
		_w5629_
	);
	LUT2 #(
		.INIT('h1)
	) name3484 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w5629_,
		_w5630_
	);
	LUT2 #(
		.INIT('h4)
	) name3485 (
		\u26_ps_cnt_reg[0]/NET0131 ,
		_w5630_,
		_w5631_
	);
	LUT2 #(
		.INIT('h4)
	) name3486 (
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		_w5632_
	);
	LUT2 #(
		.INIT('h1)
	) name3487 (
		_w5625_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h2)
	) name3488 (
		_w5630_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h8)
	) name3489 (
		\u26_ps_cnt_reg[0]/NET0131 ,
		\u26_ps_cnt_reg[1]/NET0131 ,
		_w5635_
	);
	LUT2 #(
		.INIT('h8)
	) name3490 (
		\u26_ps_cnt_reg[2]/NET0131 ,
		_w5635_,
		_w5636_
	);
	LUT2 #(
		.INIT('h1)
	) name3491 (
		\u26_ps_cnt_reg[2]/NET0131 ,
		_w5635_,
		_w5637_
	);
	LUT2 #(
		.INIT('h1)
	) name3492 (
		_w5636_,
		_w5637_,
		_w5638_
	);
	LUT2 #(
		.INIT('h8)
	) name3493 (
		_w5630_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('h1)
	) name3494 (
		\u26_ps_cnt_reg[3]/NET0131 ,
		_w5636_,
		_w5640_
	);
	LUT2 #(
		.INIT('h8)
	) name3495 (
		\u26_ps_cnt_reg[3]/NET0131 ,
		_w5636_,
		_w5641_
	);
	LUT2 #(
		.INIT('h1)
	) name3496 (
		_w5640_,
		_w5641_,
		_w5642_
	);
	LUT2 #(
		.INIT('h8)
	) name3497 (
		_w5630_,
		_w5642_,
		_w5643_
	);
	LUT2 #(
		.INIT('h8)
	) name3498 (
		\u26_ps_cnt_reg[4]/NET0131 ,
		_w5641_,
		_w5644_
	);
	LUT2 #(
		.INIT('h1)
	) name3499 (
		\u26_ps_cnt_reg[4]/NET0131 ,
		_w5641_,
		_w5645_
	);
	LUT2 #(
		.INIT('h2)
	) name3500 (
		_w5630_,
		_w5644_,
		_w5646_
	);
	LUT2 #(
		.INIT('h4)
	) name3501 (
		_w5645_,
		_w5646_,
		_w5647_
	);
	LUT2 #(
		.INIT('h1)
	) name3502 (
		\u26_ps_cnt_reg[5]/NET0131 ,
		_w5644_,
		_w5648_
	);
	LUT2 #(
		.INIT('h8)
	) name3503 (
		\u26_ps_cnt_reg[5]/NET0131 ,
		_w5644_,
		_w5649_
	);
	LUT2 #(
		.INIT('h2)
	) name3504 (
		_w5630_,
		_w5648_,
		_w5650_
	);
	LUT2 #(
		.INIT('h4)
	) name3505 (
		_w5649_,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h8)
	) name3506 (
		_w3063_,
		_w3064_,
		_w5652_
	);
	LUT2 #(
		.INIT('h1)
	) name3507 (
		\u11_wp_reg[0]/NET0131 ,
		_w5652_,
		_w5653_
	);
	LUT2 #(
		.INIT('h8)
	) name3508 (
		\u11_wp_reg[0]/NET0131 ,
		_w5652_,
		_w5654_
	);
	LUT2 #(
		.INIT('h2)
	) name3509 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w5653_,
		_w5655_
	);
	LUT2 #(
		.INIT('h4)
	) name3510 (
		_w5654_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h8)
	) name3511 (
		_w3310_,
		_w3311_,
		_w5657_
	);
	LUT2 #(
		.INIT('h1)
	) name3512 (
		\u9_wp_reg[0]/NET0131 ,
		_w5657_,
		_w5658_
	);
	LUT2 #(
		.INIT('h8)
	) name3513 (
		\u9_wp_reg[0]/NET0131 ,
		_w5657_,
		_w5659_
	);
	LUT2 #(
		.INIT('h2)
	) name3514 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w5658_,
		_w5660_
	);
	LUT2 #(
		.INIT('h4)
	) name3515 (
		_w5659_,
		_w5660_,
		_w5661_
	);
	LUT2 #(
		.INIT('h8)
	) name3516 (
		_w3500_,
		_w3501_,
		_w5662_
	);
	LUT2 #(
		.INIT('h1)
	) name3517 (
		\u10_wp_reg[0]/NET0131 ,
		_w5662_,
		_w5663_
	);
	LUT2 #(
		.INIT('h8)
	) name3518 (
		\u10_wp_reg[0]/NET0131 ,
		_w5662_,
		_w5664_
	);
	LUT2 #(
		.INIT('h2)
	) name3519 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w5663_,
		_w5665_
	);
	LUT2 #(
		.INIT('h4)
	) name3520 (
		_w5664_,
		_w5665_,
		_w5666_
	);
	LUT2 #(
		.INIT('h4)
	) name3521 (
		\u10_wp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w5667_
	);
	LUT2 #(
		.INIT('h8)
	) name3522 (
		_w3503_,
		_w5667_,
		_w5668_
	);
	LUT2 #(
		.INIT('h2)
	) name3523 (
		\u10_mem_reg[2][18]/P0001 ,
		_w5668_,
		_w5669_
	);
	LUT2 #(
		.INIT('h8)
	) name3524 (
		\u1_slt4_reg[6]/P0001 ,
		_w3501_,
		_w5670_
	);
	LUT2 #(
		.INIT('h4)
	) name3525 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w5671_
	);
	LUT2 #(
		.INIT('h8)
	) name3526 (
		\u1_slt4_reg[18]/P0001 ,
		_w5671_,
		_w5672_
	);
	LUT2 #(
		.INIT('h1)
	) name3527 (
		_w5670_,
		_w5672_,
		_w5673_
	);
	LUT2 #(
		.INIT('h2)
	) name3528 (
		_w5668_,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h1)
	) name3529 (
		_w5669_,
		_w5674_,
		_w5675_
	);
	LUT2 #(
		.INIT('h2)
	) name3530 (
		\u10_mem_reg[2][19]/P0001 ,
		_w5668_,
		_w5676_
	);
	LUT2 #(
		.INIT('h8)
	) name3531 (
		\u1_slt4_reg[7]/P0001 ,
		_w3501_,
		_w5677_
	);
	LUT2 #(
		.INIT('h8)
	) name3532 (
		\u1_slt4_reg[19]/P0001 ,
		_w5671_,
		_w5678_
	);
	LUT2 #(
		.INIT('h1)
	) name3533 (
		_w5677_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h2)
	) name3534 (
		_w5668_,
		_w5679_,
		_w5680_
	);
	LUT2 #(
		.INIT('h1)
	) name3535 (
		_w5676_,
		_w5680_,
		_w5681_
	);
	LUT2 #(
		.INIT('h2)
	) name3536 (
		\u10_mem_reg[2][20]/P0001 ,
		_w5668_,
		_w5682_
	);
	LUT2 #(
		.INIT('h8)
	) name3537 (
		\u1_slt4_reg[8]/P0001 ,
		_w3501_,
		_w5683_
	);
	LUT2 #(
		.INIT('h8)
	) name3538 (
		_w5668_,
		_w5683_,
		_w5684_
	);
	LUT2 #(
		.INIT('h1)
	) name3539 (
		_w5682_,
		_w5684_,
		_w5685_
	);
	LUT2 #(
		.INIT('h2)
	) name3540 (
		\u10_mem_reg[2][21]/P0001 ,
		_w5668_,
		_w5686_
	);
	LUT2 #(
		.INIT('h8)
	) name3541 (
		\u1_slt4_reg[9]/P0001 ,
		_w3501_,
		_w5687_
	);
	LUT2 #(
		.INIT('h8)
	) name3542 (
		_w5668_,
		_w5687_,
		_w5688_
	);
	LUT2 #(
		.INIT('h1)
	) name3543 (
		_w5686_,
		_w5688_,
		_w5689_
	);
	LUT2 #(
		.INIT('h2)
	) name3544 (
		\u10_mem_reg[2][22]/P0001 ,
		_w5668_,
		_w5690_
	);
	LUT2 #(
		.INIT('h8)
	) name3545 (
		\u1_slt4_reg[10]/P0001 ,
		_w3501_,
		_w5691_
	);
	LUT2 #(
		.INIT('h8)
	) name3546 (
		_w5668_,
		_w5691_,
		_w5692_
	);
	LUT2 #(
		.INIT('h1)
	) name3547 (
		_w5690_,
		_w5692_,
		_w5693_
	);
	LUT2 #(
		.INIT('h2)
	) name3548 (
		\u10_mem_reg[2][23]/P0001 ,
		_w5668_,
		_w5694_
	);
	LUT2 #(
		.INIT('h8)
	) name3549 (
		\u1_slt4_reg[11]/P0001 ,
		_w3501_,
		_w5695_
	);
	LUT2 #(
		.INIT('h8)
	) name3550 (
		_w5668_,
		_w5695_,
		_w5696_
	);
	LUT2 #(
		.INIT('h1)
	) name3551 (
		_w5694_,
		_w5696_,
		_w5697_
	);
	LUT2 #(
		.INIT('h1)
	) name3552 (
		\u9_wp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w5698_
	);
	LUT2 #(
		.INIT('h8)
	) name3553 (
		_w3313_,
		_w5698_,
		_w5699_
	);
	LUT2 #(
		.INIT('h8)
	) name3554 (
		\u1_slt3_reg[6]/P0001 ,
		_w3311_,
		_w5700_
	);
	LUT2 #(
		.INIT('h4)
	) name3555 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		_w5701_
	);
	LUT2 #(
		.INIT('h8)
	) name3556 (
		\u1_slt3_reg[18]/P0001 ,
		_w5701_,
		_w5702_
	);
	LUT2 #(
		.INIT('h1)
	) name3557 (
		_w5700_,
		_w5702_,
		_w5703_
	);
	LUT2 #(
		.INIT('h2)
	) name3558 (
		_w5699_,
		_w5703_,
		_w5704_
	);
	LUT2 #(
		.INIT('h2)
	) name3559 (
		\u9_mem_reg[0][18]/P0001 ,
		_w5699_,
		_w5705_
	);
	LUT2 #(
		.INIT('h1)
	) name3560 (
		_w5704_,
		_w5705_,
		_w5706_
	);
	LUT2 #(
		.INIT('h8)
	) name3561 (
		\u1_slt3_reg[7]/P0001 ,
		_w3311_,
		_w5707_
	);
	LUT2 #(
		.INIT('h8)
	) name3562 (
		\u1_slt3_reg[19]/P0001 ,
		_w5701_,
		_w5708_
	);
	LUT2 #(
		.INIT('h1)
	) name3563 (
		_w5707_,
		_w5708_,
		_w5709_
	);
	LUT2 #(
		.INIT('h2)
	) name3564 (
		_w5699_,
		_w5709_,
		_w5710_
	);
	LUT2 #(
		.INIT('h2)
	) name3565 (
		\u9_mem_reg[0][19]/P0001 ,
		_w5699_,
		_w5711_
	);
	LUT2 #(
		.INIT('h1)
	) name3566 (
		_w5710_,
		_w5711_,
		_w5712_
	);
	LUT2 #(
		.INIT('h2)
	) name3567 (
		\u10_mem_reg[2][24]/P0001 ,
		_w5668_,
		_w5713_
	);
	LUT2 #(
		.INIT('h8)
	) name3568 (
		\u1_slt4_reg[12]/P0001 ,
		_w3501_,
		_w5714_
	);
	LUT2 #(
		.INIT('h8)
	) name3569 (
		_w5668_,
		_w5714_,
		_w5715_
	);
	LUT2 #(
		.INIT('h1)
	) name3570 (
		_w5713_,
		_w5715_,
		_w5716_
	);
	LUT2 #(
		.INIT('h2)
	) name3571 (
		\u10_mem_reg[2][25]/P0001 ,
		_w5668_,
		_w5717_
	);
	LUT2 #(
		.INIT('h8)
	) name3572 (
		\u1_slt4_reg[13]/P0001 ,
		_w3501_,
		_w5718_
	);
	LUT2 #(
		.INIT('h8)
	) name3573 (
		_w5668_,
		_w5718_,
		_w5719_
	);
	LUT2 #(
		.INIT('h1)
	) name3574 (
		_w5717_,
		_w5719_,
		_w5720_
	);
	LUT2 #(
		.INIT('h2)
	) name3575 (
		\u10_mem_reg[2][26]/P0001 ,
		_w5668_,
		_w5721_
	);
	LUT2 #(
		.INIT('h8)
	) name3576 (
		\u1_slt4_reg[14]/P0001 ,
		_w3501_,
		_w5722_
	);
	LUT2 #(
		.INIT('h8)
	) name3577 (
		_w5668_,
		_w5722_,
		_w5723_
	);
	LUT2 #(
		.INIT('h1)
	) name3578 (
		_w5721_,
		_w5723_,
		_w5724_
	);
	LUT2 #(
		.INIT('h2)
	) name3579 (
		\u10_mem_reg[2][27]/P0001 ,
		_w5668_,
		_w5725_
	);
	LUT2 #(
		.INIT('h8)
	) name3580 (
		\u1_slt4_reg[15]/P0001 ,
		_w3501_,
		_w5726_
	);
	LUT2 #(
		.INIT('h8)
	) name3581 (
		_w5668_,
		_w5726_,
		_w5727_
	);
	LUT2 #(
		.INIT('h1)
	) name3582 (
		_w5725_,
		_w5727_,
		_w5728_
	);
	LUT2 #(
		.INIT('h2)
	) name3583 (
		\u10_mem_reg[2][28]/P0001 ,
		_w5668_,
		_w5729_
	);
	LUT2 #(
		.INIT('h8)
	) name3584 (
		\u1_slt4_reg[16]/P0001 ,
		_w3501_,
		_w5730_
	);
	LUT2 #(
		.INIT('h8)
	) name3585 (
		_w5668_,
		_w5730_,
		_w5731_
	);
	LUT2 #(
		.INIT('h1)
	) name3586 (
		_w5729_,
		_w5731_,
		_w5732_
	);
	LUT2 #(
		.INIT('h4)
	) name3587 (
		\u9_wp_reg[2]/P0001 ,
		_w3314_,
		_w5733_
	);
	LUT2 #(
		.INIT('h4)
	) name3588 (
		_w5703_,
		_w5733_,
		_w5734_
	);
	LUT2 #(
		.INIT('h2)
	) name3589 (
		\u9_mem_reg[1][18]/P0001 ,
		_w5733_,
		_w5735_
	);
	LUT2 #(
		.INIT('h1)
	) name3590 (
		_w5734_,
		_w5735_,
		_w5736_
	);
	LUT2 #(
		.INIT('h4)
	) name3591 (
		_w5709_,
		_w5733_,
		_w5737_
	);
	LUT2 #(
		.INIT('h2)
	) name3592 (
		\u9_mem_reg[1][19]/P0001 ,
		_w5733_,
		_w5738_
	);
	LUT2 #(
		.INIT('h1)
	) name3593 (
		_w5737_,
		_w5738_,
		_w5739_
	);
	LUT2 #(
		.INIT('h2)
	) name3594 (
		\u9_mem_reg[1][20]/P0001 ,
		_w5733_,
		_w5740_
	);
	LUT2 #(
		.INIT('h8)
	) name3595 (
		\u1_slt3_reg[8]/P0001 ,
		_w3311_,
		_w5741_
	);
	LUT2 #(
		.INIT('h8)
	) name3596 (
		_w5733_,
		_w5741_,
		_w5742_
	);
	LUT2 #(
		.INIT('h1)
	) name3597 (
		_w5740_,
		_w5742_,
		_w5743_
	);
	LUT2 #(
		.INIT('h2)
	) name3598 (
		\u9_mem_reg[1][21]/P0001 ,
		_w5733_,
		_w5744_
	);
	LUT2 #(
		.INIT('h8)
	) name3599 (
		\u1_slt3_reg[9]/P0001 ,
		_w3311_,
		_w5745_
	);
	LUT2 #(
		.INIT('h8)
	) name3600 (
		_w5733_,
		_w5745_,
		_w5746_
	);
	LUT2 #(
		.INIT('h1)
	) name3601 (
		_w5744_,
		_w5746_,
		_w5747_
	);
	LUT2 #(
		.INIT('h2)
	) name3602 (
		\u10_mem_reg[2][29]/P0001 ,
		_w5668_,
		_w5748_
	);
	LUT2 #(
		.INIT('h8)
	) name3603 (
		\u1_slt4_reg[17]/P0001 ,
		_w3501_,
		_w5749_
	);
	LUT2 #(
		.INIT('h8)
	) name3604 (
		_w5668_,
		_w5749_,
		_w5750_
	);
	LUT2 #(
		.INIT('h1)
	) name3605 (
		_w5748_,
		_w5750_,
		_w5751_
	);
	LUT2 #(
		.INIT('h2)
	) name3606 (
		\u9_mem_reg[1][22]/P0001 ,
		_w5733_,
		_w5752_
	);
	LUT2 #(
		.INIT('h8)
	) name3607 (
		\u1_slt3_reg[10]/P0001 ,
		_w3311_,
		_w5753_
	);
	LUT2 #(
		.INIT('h8)
	) name3608 (
		_w5733_,
		_w5753_,
		_w5754_
	);
	LUT2 #(
		.INIT('h1)
	) name3609 (
		_w5752_,
		_w5754_,
		_w5755_
	);
	LUT2 #(
		.INIT('h2)
	) name3610 (
		\u9_mem_reg[1][23]/P0001 ,
		_w5733_,
		_w5756_
	);
	LUT2 #(
		.INIT('h8)
	) name3611 (
		\u1_slt3_reg[11]/P0001 ,
		_w3311_,
		_w5757_
	);
	LUT2 #(
		.INIT('h8)
	) name3612 (
		_w5733_,
		_w5757_,
		_w5758_
	);
	LUT2 #(
		.INIT('h1)
	) name3613 (
		_w5756_,
		_w5758_,
		_w5759_
	);
	LUT2 #(
		.INIT('h2)
	) name3614 (
		\u9_mem_reg[1][24]/P0001 ,
		_w5733_,
		_w5760_
	);
	LUT2 #(
		.INIT('h8)
	) name3615 (
		\u1_slt3_reg[12]/P0001 ,
		_w3311_,
		_w5761_
	);
	LUT2 #(
		.INIT('h8)
	) name3616 (
		_w5733_,
		_w5761_,
		_w5762_
	);
	LUT2 #(
		.INIT('h1)
	) name3617 (
		_w5760_,
		_w5762_,
		_w5763_
	);
	LUT2 #(
		.INIT('h2)
	) name3618 (
		\u9_mem_reg[1][25]/P0001 ,
		_w5733_,
		_w5764_
	);
	LUT2 #(
		.INIT('h8)
	) name3619 (
		\u1_slt3_reg[13]/P0001 ,
		_w3311_,
		_w5765_
	);
	LUT2 #(
		.INIT('h8)
	) name3620 (
		_w5733_,
		_w5765_,
		_w5766_
	);
	LUT2 #(
		.INIT('h1)
	) name3621 (
		_w5764_,
		_w5766_,
		_w5767_
	);
	LUT2 #(
		.INIT('h2)
	) name3622 (
		\u9_mem_reg[1][26]/P0001 ,
		_w5733_,
		_w5768_
	);
	LUT2 #(
		.INIT('h8)
	) name3623 (
		\u1_slt3_reg[14]/P0001 ,
		_w3311_,
		_w5769_
	);
	LUT2 #(
		.INIT('h8)
	) name3624 (
		_w5733_,
		_w5769_,
		_w5770_
	);
	LUT2 #(
		.INIT('h1)
	) name3625 (
		_w5768_,
		_w5770_,
		_w5771_
	);
	LUT2 #(
		.INIT('h2)
	) name3626 (
		\u9_mem_reg[1][27]/P0001 ,
		_w5733_,
		_w5772_
	);
	LUT2 #(
		.INIT('h8)
	) name3627 (
		\u1_slt3_reg[15]/P0001 ,
		_w3311_,
		_w5773_
	);
	LUT2 #(
		.INIT('h8)
	) name3628 (
		_w5733_,
		_w5773_,
		_w5774_
	);
	LUT2 #(
		.INIT('h1)
	) name3629 (
		_w5772_,
		_w5774_,
		_w5775_
	);
	LUT2 #(
		.INIT('h2)
	) name3630 (
		\u9_mem_reg[1][28]/P0001 ,
		_w5733_,
		_w5776_
	);
	LUT2 #(
		.INIT('h8)
	) name3631 (
		\u1_slt3_reg[16]/P0001 ,
		_w3311_,
		_w5777_
	);
	LUT2 #(
		.INIT('h8)
	) name3632 (
		_w5733_,
		_w5777_,
		_w5778_
	);
	LUT2 #(
		.INIT('h1)
	) name3633 (
		_w5776_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h2)
	) name3634 (
		\u9_mem_reg[1][29]/P0001 ,
		_w5733_,
		_w5780_
	);
	LUT2 #(
		.INIT('h8)
	) name3635 (
		\u1_slt3_reg[17]/P0001 ,
		_w3311_,
		_w5781_
	);
	LUT2 #(
		.INIT('h8)
	) name3636 (
		_w5733_,
		_w5781_,
		_w5782_
	);
	LUT2 #(
		.INIT('h1)
	) name3637 (
		_w5780_,
		_w5782_,
		_w5783_
	);
	LUT2 #(
		.INIT('h2)
	) name3638 (
		\u9_mem_reg[1][30]/P0001 ,
		_w5733_,
		_w5784_
	);
	LUT2 #(
		.INIT('h8)
	) name3639 (
		\u1_slt3_reg[18]/P0001 ,
		_w3311_,
		_w5785_
	);
	LUT2 #(
		.INIT('h8)
	) name3640 (
		_w5733_,
		_w5785_,
		_w5786_
	);
	LUT2 #(
		.INIT('h1)
	) name3641 (
		_w5784_,
		_w5786_,
		_w5787_
	);
	LUT2 #(
		.INIT('h2)
	) name3642 (
		\u9_mem_reg[1][31]/P0001 ,
		_w5733_,
		_w5788_
	);
	LUT2 #(
		.INIT('h8)
	) name3643 (
		\u1_slt3_reg[19]/P0001 ,
		_w3311_,
		_w5789_
	);
	LUT2 #(
		.INIT('h8)
	) name3644 (
		_w5733_,
		_w5789_,
		_w5790_
	);
	LUT2 #(
		.INIT('h1)
	) name3645 (
		_w5788_,
		_w5790_,
		_w5791_
	);
	LUT2 #(
		.INIT('h2)
	) name3646 (
		\u10_mem_reg[2][30]/P0001 ,
		_w5668_,
		_w5792_
	);
	LUT2 #(
		.INIT('h8)
	) name3647 (
		\u1_slt4_reg[18]/P0001 ,
		_w3501_,
		_w5793_
	);
	LUT2 #(
		.INIT('h8)
	) name3648 (
		_w5668_,
		_w5793_,
		_w5794_
	);
	LUT2 #(
		.INIT('h1)
	) name3649 (
		_w5792_,
		_w5794_,
		_w5795_
	);
	LUT2 #(
		.INIT('h2)
	) name3650 (
		\u10_mem_reg[2][31]/P0001 ,
		_w5668_,
		_w5796_
	);
	LUT2 #(
		.INIT('h8)
	) name3651 (
		\u1_slt4_reg[19]/P0001 ,
		_w3501_,
		_w5797_
	);
	LUT2 #(
		.INIT('h8)
	) name3652 (
		_w5668_,
		_w5797_,
		_w5798_
	);
	LUT2 #(
		.INIT('h1)
	) name3653 (
		_w5796_,
		_w5798_,
		_w5799_
	);
	LUT2 #(
		.INIT('h4)
	) name3654 (
		\u9_wp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w5800_
	);
	LUT2 #(
		.INIT('h8)
	) name3655 (
		_w3313_,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h2)
	) name3656 (
		\u9_mem_reg[2][18]/P0001 ,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h4)
	) name3657 (
		_w5703_,
		_w5801_,
		_w5803_
	);
	LUT2 #(
		.INIT('h1)
	) name3658 (
		_w5802_,
		_w5803_,
		_w5804_
	);
	LUT2 #(
		.INIT('h2)
	) name3659 (
		\u9_mem_reg[2][19]/P0001 ,
		_w5801_,
		_w5805_
	);
	LUT2 #(
		.INIT('h4)
	) name3660 (
		_w5709_,
		_w5801_,
		_w5806_
	);
	LUT2 #(
		.INIT('h1)
	) name3661 (
		_w5805_,
		_w5806_,
		_w5807_
	);
	LUT2 #(
		.INIT('h2)
	) name3662 (
		\u9_mem_reg[2][20]/P0001 ,
		_w5801_,
		_w5808_
	);
	LUT2 #(
		.INIT('h8)
	) name3663 (
		_w5741_,
		_w5801_,
		_w5809_
	);
	LUT2 #(
		.INIT('h1)
	) name3664 (
		_w5808_,
		_w5809_,
		_w5810_
	);
	LUT2 #(
		.INIT('h2)
	) name3665 (
		\u9_mem_reg[2][21]/P0001 ,
		_w5801_,
		_w5811_
	);
	LUT2 #(
		.INIT('h8)
	) name3666 (
		_w5745_,
		_w5801_,
		_w5812_
	);
	LUT2 #(
		.INIT('h1)
	) name3667 (
		_w5811_,
		_w5812_,
		_w5813_
	);
	LUT2 #(
		.INIT('h2)
	) name3668 (
		\u9_mem_reg[2][22]/P0001 ,
		_w5801_,
		_w5814_
	);
	LUT2 #(
		.INIT('h8)
	) name3669 (
		_w5753_,
		_w5801_,
		_w5815_
	);
	LUT2 #(
		.INIT('h1)
	) name3670 (
		_w5814_,
		_w5815_,
		_w5816_
	);
	LUT2 #(
		.INIT('h2)
	) name3671 (
		\u9_mem_reg[2][23]/P0001 ,
		_w5801_,
		_w5817_
	);
	LUT2 #(
		.INIT('h8)
	) name3672 (
		_w5757_,
		_w5801_,
		_w5818_
	);
	LUT2 #(
		.INIT('h1)
	) name3673 (
		_w5817_,
		_w5818_,
		_w5819_
	);
	LUT2 #(
		.INIT('h2)
	) name3674 (
		\u9_mem_reg[2][24]/P0001 ,
		_w5801_,
		_w5820_
	);
	LUT2 #(
		.INIT('h8)
	) name3675 (
		_w5761_,
		_w5801_,
		_w5821_
	);
	LUT2 #(
		.INIT('h1)
	) name3676 (
		_w5820_,
		_w5821_,
		_w5822_
	);
	LUT2 #(
		.INIT('h2)
	) name3677 (
		\u9_mem_reg[2][25]/P0001 ,
		_w5801_,
		_w5823_
	);
	LUT2 #(
		.INIT('h8)
	) name3678 (
		_w5765_,
		_w5801_,
		_w5824_
	);
	LUT2 #(
		.INIT('h1)
	) name3679 (
		_w5823_,
		_w5824_,
		_w5825_
	);
	LUT2 #(
		.INIT('h2)
	) name3680 (
		\u9_mem_reg[2][26]/P0001 ,
		_w5801_,
		_w5826_
	);
	LUT2 #(
		.INIT('h8)
	) name3681 (
		_w5769_,
		_w5801_,
		_w5827_
	);
	LUT2 #(
		.INIT('h1)
	) name3682 (
		_w5826_,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h2)
	) name3683 (
		\u9_mem_reg[2][27]/P0001 ,
		_w5801_,
		_w5829_
	);
	LUT2 #(
		.INIT('h8)
	) name3684 (
		_w5773_,
		_w5801_,
		_w5830_
	);
	LUT2 #(
		.INIT('h1)
	) name3685 (
		_w5829_,
		_w5830_,
		_w5831_
	);
	LUT2 #(
		.INIT('h2)
	) name3686 (
		\u9_mem_reg[2][28]/P0001 ,
		_w5801_,
		_w5832_
	);
	LUT2 #(
		.INIT('h8)
	) name3687 (
		_w5777_,
		_w5801_,
		_w5833_
	);
	LUT2 #(
		.INIT('h1)
	) name3688 (
		_w5832_,
		_w5833_,
		_w5834_
	);
	LUT2 #(
		.INIT('h2)
	) name3689 (
		\u9_mem_reg[2][29]/P0001 ,
		_w5801_,
		_w5835_
	);
	LUT2 #(
		.INIT('h8)
	) name3690 (
		_w5781_,
		_w5801_,
		_w5836_
	);
	LUT2 #(
		.INIT('h1)
	) name3691 (
		_w5835_,
		_w5836_,
		_w5837_
	);
	LUT2 #(
		.INIT('h2)
	) name3692 (
		\u9_mem_reg[2][30]/P0001 ,
		_w5801_,
		_w5838_
	);
	LUT2 #(
		.INIT('h8)
	) name3693 (
		_w5785_,
		_w5801_,
		_w5839_
	);
	LUT2 #(
		.INIT('h1)
	) name3694 (
		_w5838_,
		_w5839_,
		_w5840_
	);
	LUT2 #(
		.INIT('h2)
	) name3695 (
		\u9_mem_reg[2][31]/P0001 ,
		_w5801_,
		_w5841_
	);
	LUT2 #(
		.INIT('h8)
	) name3696 (
		_w5789_,
		_w5801_,
		_w5842_
	);
	LUT2 #(
		.INIT('h1)
	) name3697 (
		_w5841_,
		_w5842_,
		_w5843_
	);
	LUT2 #(
		.INIT('h2)
	) name3698 (
		_w3315_,
		_w5703_,
		_w5844_
	);
	LUT2 #(
		.INIT('h2)
	) name3699 (
		\u9_mem_reg[3][18]/P0001 ,
		_w3315_,
		_w5845_
	);
	LUT2 #(
		.INIT('h1)
	) name3700 (
		_w5844_,
		_w5845_,
		_w5846_
	);
	LUT2 #(
		.INIT('h2)
	) name3701 (
		_w3315_,
		_w5709_,
		_w5847_
	);
	LUT2 #(
		.INIT('h2)
	) name3702 (
		\u9_mem_reg[3][19]/P0001 ,
		_w3315_,
		_w5848_
	);
	LUT2 #(
		.INIT('h1)
	) name3703 (
		_w5847_,
		_w5848_,
		_w5849_
	);
	LUT2 #(
		.INIT('h2)
	) name3704 (
		\u9_mem_reg[3][20]/P0001 ,
		_w3315_,
		_w5850_
	);
	LUT2 #(
		.INIT('h8)
	) name3705 (
		_w3315_,
		_w5741_,
		_w5851_
	);
	LUT2 #(
		.INIT('h1)
	) name3706 (
		_w5850_,
		_w5851_,
		_w5852_
	);
	LUT2 #(
		.INIT('h2)
	) name3707 (
		\u9_mem_reg[3][21]/P0001 ,
		_w3315_,
		_w5853_
	);
	LUT2 #(
		.INIT('h8)
	) name3708 (
		_w3315_,
		_w5745_,
		_w5854_
	);
	LUT2 #(
		.INIT('h1)
	) name3709 (
		_w5853_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h2)
	) name3710 (
		\u9_mem_reg[3][22]/P0001 ,
		_w3315_,
		_w5856_
	);
	LUT2 #(
		.INIT('h8)
	) name3711 (
		_w3315_,
		_w5753_,
		_w5857_
	);
	LUT2 #(
		.INIT('h1)
	) name3712 (
		_w5856_,
		_w5857_,
		_w5858_
	);
	LUT2 #(
		.INIT('h2)
	) name3713 (
		\u9_mem_reg[3][23]/P0001 ,
		_w3315_,
		_w5859_
	);
	LUT2 #(
		.INIT('h8)
	) name3714 (
		_w3315_,
		_w5757_,
		_w5860_
	);
	LUT2 #(
		.INIT('h1)
	) name3715 (
		_w5859_,
		_w5860_,
		_w5861_
	);
	LUT2 #(
		.INIT('h2)
	) name3716 (
		\u9_mem_reg[3][24]/P0001 ,
		_w3315_,
		_w5862_
	);
	LUT2 #(
		.INIT('h8)
	) name3717 (
		_w3315_,
		_w5761_,
		_w5863_
	);
	LUT2 #(
		.INIT('h1)
	) name3718 (
		_w5862_,
		_w5863_,
		_w5864_
	);
	LUT2 #(
		.INIT('h2)
	) name3719 (
		\u9_mem_reg[3][25]/P0001 ,
		_w3315_,
		_w5865_
	);
	LUT2 #(
		.INIT('h8)
	) name3720 (
		_w3315_,
		_w5765_,
		_w5866_
	);
	LUT2 #(
		.INIT('h1)
	) name3721 (
		_w5865_,
		_w5866_,
		_w5867_
	);
	LUT2 #(
		.INIT('h2)
	) name3722 (
		\u9_mem_reg[3][26]/P0001 ,
		_w3315_,
		_w5868_
	);
	LUT2 #(
		.INIT('h8)
	) name3723 (
		_w3315_,
		_w5769_,
		_w5869_
	);
	LUT2 #(
		.INIT('h1)
	) name3724 (
		_w5868_,
		_w5869_,
		_w5870_
	);
	LUT2 #(
		.INIT('h2)
	) name3725 (
		\u9_mem_reg[3][27]/P0001 ,
		_w3315_,
		_w5871_
	);
	LUT2 #(
		.INIT('h8)
	) name3726 (
		_w3315_,
		_w5773_,
		_w5872_
	);
	LUT2 #(
		.INIT('h1)
	) name3727 (
		_w5871_,
		_w5872_,
		_w5873_
	);
	LUT2 #(
		.INIT('h2)
	) name3728 (
		\u9_mem_reg[3][28]/P0001 ,
		_w3315_,
		_w5874_
	);
	LUT2 #(
		.INIT('h8)
	) name3729 (
		_w3315_,
		_w5777_,
		_w5875_
	);
	LUT2 #(
		.INIT('h1)
	) name3730 (
		_w5874_,
		_w5875_,
		_w5876_
	);
	LUT2 #(
		.INIT('h2)
	) name3731 (
		\u9_mem_reg[3][29]/P0001 ,
		_w3315_,
		_w5877_
	);
	LUT2 #(
		.INIT('h8)
	) name3732 (
		_w3315_,
		_w5781_,
		_w5878_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		_w5877_,
		_w5878_,
		_w5879_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		\u9_mem_reg[3][30]/P0001 ,
		_w3315_,
		_w5880_
	);
	LUT2 #(
		.INIT('h8)
	) name3735 (
		_w3315_,
		_w5785_,
		_w5881_
	);
	LUT2 #(
		.INIT('h1)
	) name3736 (
		_w5880_,
		_w5881_,
		_w5882_
	);
	LUT2 #(
		.INIT('h2)
	) name3737 (
		\u9_mem_reg[3][31]/P0001 ,
		_w3315_,
		_w5883_
	);
	LUT2 #(
		.INIT('h8)
	) name3738 (
		_w3315_,
		_w5789_,
		_w5884_
	);
	LUT2 #(
		.INIT('h1)
	) name3739 (
		_w5883_,
		_w5884_,
		_w5885_
	);
	LUT2 #(
		.INIT('h2)
	) name3740 (
		_w3505_,
		_w5673_,
		_w5886_
	);
	LUT2 #(
		.INIT('h2)
	) name3741 (
		\u10_mem_reg[3][18]/P0001 ,
		_w3505_,
		_w5887_
	);
	LUT2 #(
		.INIT('h1)
	) name3742 (
		_w5886_,
		_w5887_,
		_w5888_
	);
	LUT2 #(
		.INIT('h2)
	) name3743 (
		_w3505_,
		_w5679_,
		_w5889_
	);
	LUT2 #(
		.INIT('h2)
	) name3744 (
		\u10_mem_reg[3][19]/P0001 ,
		_w3505_,
		_w5890_
	);
	LUT2 #(
		.INIT('h1)
	) name3745 (
		_w5889_,
		_w5890_,
		_w5891_
	);
	LUT2 #(
		.INIT('h2)
	) name3746 (
		\u10_mem_reg[3][20]/P0001 ,
		_w3505_,
		_w5892_
	);
	LUT2 #(
		.INIT('h8)
	) name3747 (
		_w3505_,
		_w5683_,
		_w5893_
	);
	LUT2 #(
		.INIT('h1)
	) name3748 (
		_w5892_,
		_w5893_,
		_w5894_
	);
	LUT2 #(
		.INIT('h2)
	) name3749 (
		\u10_mem_reg[3][21]/P0001 ,
		_w3505_,
		_w5895_
	);
	LUT2 #(
		.INIT('h8)
	) name3750 (
		_w3505_,
		_w5687_,
		_w5896_
	);
	LUT2 #(
		.INIT('h1)
	) name3751 (
		_w5895_,
		_w5896_,
		_w5897_
	);
	LUT2 #(
		.INIT('h2)
	) name3752 (
		\u10_mem_reg[3][22]/P0001 ,
		_w3505_,
		_w5898_
	);
	LUT2 #(
		.INIT('h8)
	) name3753 (
		_w3505_,
		_w5691_,
		_w5899_
	);
	LUT2 #(
		.INIT('h1)
	) name3754 (
		_w5898_,
		_w5899_,
		_w5900_
	);
	LUT2 #(
		.INIT('h2)
	) name3755 (
		\u10_mem_reg[3][23]/P0001 ,
		_w3505_,
		_w5901_
	);
	LUT2 #(
		.INIT('h8)
	) name3756 (
		_w3505_,
		_w5695_,
		_w5902_
	);
	LUT2 #(
		.INIT('h1)
	) name3757 (
		_w5901_,
		_w5902_,
		_w5903_
	);
	LUT2 #(
		.INIT('h2)
	) name3758 (
		\u10_mem_reg[3][24]/P0001 ,
		_w3505_,
		_w5904_
	);
	LUT2 #(
		.INIT('h8)
	) name3759 (
		_w3505_,
		_w5714_,
		_w5905_
	);
	LUT2 #(
		.INIT('h1)
	) name3760 (
		_w5904_,
		_w5905_,
		_w5906_
	);
	LUT2 #(
		.INIT('h2)
	) name3761 (
		\u10_mem_reg[3][25]/P0001 ,
		_w3505_,
		_w5907_
	);
	LUT2 #(
		.INIT('h8)
	) name3762 (
		_w3505_,
		_w5718_,
		_w5908_
	);
	LUT2 #(
		.INIT('h1)
	) name3763 (
		_w5907_,
		_w5908_,
		_w5909_
	);
	LUT2 #(
		.INIT('h2)
	) name3764 (
		\u10_mem_reg[3][26]/P0001 ,
		_w3505_,
		_w5910_
	);
	LUT2 #(
		.INIT('h8)
	) name3765 (
		_w3505_,
		_w5722_,
		_w5911_
	);
	LUT2 #(
		.INIT('h1)
	) name3766 (
		_w5910_,
		_w5911_,
		_w5912_
	);
	LUT2 #(
		.INIT('h2)
	) name3767 (
		\u10_mem_reg[3][27]/P0001 ,
		_w3505_,
		_w5913_
	);
	LUT2 #(
		.INIT('h8)
	) name3768 (
		_w3505_,
		_w5726_,
		_w5914_
	);
	LUT2 #(
		.INIT('h1)
	) name3769 (
		_w5913_,
		_w5914_,
		_w5915_
	);
	LUT2 #(
		.INIT('h2)
	) name3770 (
		\u10_mem_reg[3][28]/P0001 ,
		_w3505_,
		_w5916_
	);
	LUT2 #(
		.INIT('h8)
	) name3771 (
		_w3505_,
		_w5730_,
		_w5917_
	);
	LUT2 #(
		.INIT('h1)
	) name3772 (
		_w5916_,
		_w5917_,
		_w5918_
	);
	LUT2 #(
		.INIT('h2)
	) name3773 (
		\u10_mem_reg[3][29]/P0001 ,
		_w3505_,
		_w5919_
	);
	LUT2 #(
		.INIT('h8)
	) name3774 (
		_w3505_,
		_w5749_,
		_w5920_
	);
	LUT2 #(
		.INIT('h1)
	) name3775 (
		_w5919_,
		_w5920_,
		_w5921_
	);
	LUT2 #(
		.INIT('h2)
	) name3776 (
		\u10_mem_reg[3][30]/P0001 ,
		_w3505_,
		_w5922_
	);
	LUT2 #(
		.INIT('h8)
	) name3777 (
		_w3505_,
		_w5793_,
		_w5923_
	);
	LUT2 #(
		.INIT('h1)
	) name3778 (
		_w5922_,
		_w5923_,
		_w5924_
	);
	LUT2 #(
		.INIT('h2)
	) name3779 (
		\u10_mem_reg[3][31]/P0001 ,
		_w3505_,
		_w5925_
	);
	LUT2 #(
		.INIT('h8)
	) name3780 (
		_w3505_,
		_w5797_,
		_w5926_
	);
	LUT2 #(
		.INIT('h1)
	) name3781 (
		_w5925_,
		_w5926_,
		_w5927_
	);
	LUT2 #(
		.INIT('h1)
	) name3782 (
		\u10_wp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w5928_
	);
	LUT2 #(
		.INIT('h8)
	) name3783 (
		_w3503_,
		_w5928_,
		_w5929_
	);
	LUT2 #(
		.INIT('h2)
	) name3784 (
		\u10_mem_reg[0][18]/P0001 ,
		_w5929_,
		_w5930_
	);
	LUT2 #(
		.INIT('h4)
	) name3785 (
		_w5673_,
		_w5929_,
		_w5931_
	);
	LUT2 #(
		.INIT('h1)
	) name3786 (
		_w5930_,
		_w5931_,
		_w5932_
	);
	LUT2 #(
		.INIT('h1)
	) name3787 (
		\u11_wp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w5933_
	);
	LUT2 #(
		.INIT('h8)
	) name3788 (
		_w3066_,
		_w5933_,
		_w5934_
	);
	LUT2 #(
		.INIT('h8)
	) name3789 (
		\u1_slt6_reg[6]/P0001 ,
		_w3064_,
		_w5935_
	);
	LUT2 #(
		.INIT('h4)
	) name3790 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w5936_
	);
	LUT2 #(
		.INIT('h8)
	) name3791 (
		\u1_slt6_reg[18]/P0001 ,
		_w5936_,
		_w5937_
	);
	LUT2 #(
		.INIT('h1)
	) name3792 (
		_w5935_,
		_w5937_,
		_w5938_
	);
	LUT2 #(
		.INIT('h2)
	) name3793 (
		_w5934_,
		_w5938_,
		_w5939_
	);
	LUT2 #(
		.INIT('h2)
	) name3794 (
		\u11_mem_reg[0][18]/P0001 ,
		_w5934_,
		_w5940_
	);
	LUT2 #(
		.INIT('h1)
	) name3795 (
		_w5939_,
		_w5940_,
		_w5941_
	);
	LUT2 #(
		.INIT('h8)
	) name3796 (
		\u1_slt6_reg[7]/P0001 ,
		_w3064_,
		_w5942_
	);
	LUT2 #(
		.INIT('h8)
	) name3797 (
		\u1_slt6_reg[19]/P0001 ,
		_w5936_,
		_w5943_
	);
	LUT2 #(
		.INIT('h1)
	) name3798 (
		_w5942_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h2)
	) name3799 (
		_w5934_,
		_w5944_,
		_w5945_
	);
	LUT2 #(
		.INIT('h2)
	) name3800 (
		\u11_mem_reg[0][19]/P0001 ,
		_w5934_,
		_w5946_
	);
	LUT2 #(
		.INIT('h1)
	) name3801 (
		_w5945_,
		_w5946_,
		_w5947_
	);
	LUT2 #(
		.INIT('h2)
	) name3802 (
		\u10_mem_reg[0][19]/P0001 ,
		_w5929_,
		_w5948_
	);
	LUT2 #(
		.INIT('h4)
	) name3803 (
		_w5679_,
		_w5929_,
		_w5949_
	);
	LUT2 #(
		.INIT('h1)
	) name3804 (
		_w5948_,
		_w5949_,
		_w5950_
	);
	LUT2 #(
		.INIT('h4)
	) name3805 (
		\u11_wp_reg[2]/P0001 ,
		_w3067_,
		_w5951_
	);
	LUT2 #(
		.INIT('h4)
	) name3806 (
		_w5938_,
		_w5951_,
		_w5952_
	);
	LUT2 #(
		.INIT('h2)
	) name3807 (
		\u11_mem_reg[1][18]/P0001 ,
		_w5951_,
		_w5953_
	);
	LUT2 #(
		.INIT('h1)
	) name3808 (
		_w5952_,
		_w5953_,
		_w5954_
	);
	LUT2 #(
		.INIT('h4)
	) name3809 (
		_w5944_,
		_w5951_,
		_w5955_
	);
	LUT2 #(
		.INIT('h2)
	) name3810 (
		\u11_mem_reg[1][19]/P0001 ,
		_w5951_,
		_w5956_
	);
	LUT2 #(
		.INIT('h1)
	) name3811 (
		_w5955_,
		_w5956_,
		_w5957_
	);
	LUT2 #(
		.INIT('h2)
	) name3812 (
		\u11_mem_reg[1][20]/P0001 ,
		_w5951_,
		_w5958_
	);
	LUT2 #(
		.INIT('h8)
	) name3813 (
		\u1_slt6_reg[8]/P0001 ,
		_w3064_,
		_w5959_
	);
	LUT2 #(
		.INIT('h8)
	) name3814 (
		_w5951_,
		_w5959_,
		_w5960_
	);
	LUT2 #(
		.INIT('h1)
	) name3815 (
		_w5958_,
		_w5960_,
		_w5961_
	);
	LUT2 #(
		.INIT('h2)
	) name3816 (
		\u11_mem_reg[1][21]/P0001 ,
		_w5951_,
		_w5962_
	);
	LUT2 #(
		.INIT('h8)
	) name3817 (
		\u1_slt6_reg[9]/P0001 ,
		_w3064_,
		_w5963_
	);
	LUT2 #(
		.INIT('h8)
	) name3818 (
		_w5951_,
		_w5963_,
		_w5964_
	);
	LUT2 #(
		.INIT('h1)
	) name3819 (
		_w5962_,
		_w5964_,
		_w5965_
	);
	LUT2 #(
		.INIT('h2)
	) name3820 (
		\u11_mem_reg[1][22]/P0001 ,
		_w5951_,
		_w5966_
	);
	LUT2 #(
		.INIT('h8)
	) name3821 (
		\u1_slt6_reg[10]/P0001 ,
		_w3064_,
		_w5967_
	);
	LUT2 #(
		.INIT('h8)
	) name3822 (
		_w5951_,
		_w5967_,
		_w5968_
	);
	LUT2 #(
		.INIT('h1)
	) name3823 (
		_w5966_,
		_w5968_,
		_w5969_
	);
	LUT2 #(
		.INIT('h2)
	) name3824 (
		\u11_mem_reg[1][23]/P0001 ,
		_w5951_,
		_w5970_
	);
	LUT2 #(
		.INIT('h8)
	) name3825 (
		\u1_slt6_reg[11]/P0001 ,
		_w3064_,
		_w5971_
	);
	LUT2 #(
		.INIT('h8)
	) name3826 (
		_w5951_,
		_w5971_,
		_w5972_
	);
	LUT2 #(
		.INIT('h1)
	) name3827 (
		_w5970_,
		_w5972_,
		_w5973_
	);
	LUT2 #(
		.INIT('h2)
	) name3828 (
		\u11_mem_reg[1][24]/P0001 ,
		_w5951_,
		_w5974_
	);
	LUT2 #(
		.INIT('h8)
	) name3829 (
		\u1_slt6_reg[12]/P0001 ,
		_w3064_,
		_w5975_
	);
	LUT2 #(
		.INIT('h8)
	) name3830 (
		_w5951_,
		_w5975_,
		_w5976_
	);
	LUT2 #(
		.INIT('h1)
	) name3831 (
		_w5974_,
		_w5976_,
		_w5977_
	);
	LUT2 #(
		.INIT('h2)
	) name3832 (
		\u11_mem_reg[1][25]/P0001 ,
		_w5951_,
		_w5978_
	);
	LUT2 #(
		.INIT('h8)
	) name3833 (
		\u1_slt6_reg[13]/P0001 ,
		_w3064_,
		_w5979_
	);
	LUT2 #(
		.INIT('h8)
	) name3834 (
		_w5951_,
		_w5979_,
		_w5980_
	);
	LUT2 #(
		.INIT('h1)
	) name3835 (
		_w5978_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h2)
	) name3836 (
		\u11_mem_reg[1][26]/P0001 ,
		_w5951_,
		_w5982_
	);
	LUT2 #(
		.INIT('h8)
	) name3837 (
		\u1_slt6_reg[14]/P0001 ,
		_w3064_,
		_w5983_
	);
	LUT2 #(
		.INIT('h8)
	) name3838 (
		_w5951_,
		_w5983_,
		_w5984_
	);
	LUT2 #(
		.INIT('h1)
	) name3839 (
		_w5982_,
		_w5984_,
		_w5985_
	);
	LUT2 #(
		.INIT('h2)
	) name3840 (
		\u11_mem_reg[1][27]/P0001 ,
		_w5951_,
		_w5986_
	);
	LUT2 #(
		.INIT('h8)
	) name3841 (
		\u1_slt6_reg[15]/P0001 ,
		_w3064_,
		_w5987_
	);
	LUT2 #(
		.INIT('h8)
	) name3842 (
		_w5951_,
		_w5987_,
		_w5988_
	);
	LUT2 #(
		.INIT('h1)
	) name3843 (
		_w5986_,
		_w5988_,
		_w5989_
	);
	LUT2 #(
		.INIT('h2)
	) name3844 (
		\u11_mem_reg[1][28]/P0001 ,
		_w5951_,
		_w5990_
	);
	LUT2 #(
		.INIT('h8)
	) name3845 (
		\u1_slt6_reg[16]/P0001 ,
		_w3064_,
		_w5991_
	);
	LUT2 #(
		.INIT('h8)
	) name3846 (
		_w5951_,
		_w5991_,
		_w5992_
	);
	LUT2 #(
		.INIT('h1)
	) name3847 (
		_w5990_,
		_w5992_,
		_w5993_
	);
	LUT2 #(
		.INIT('h2)
	) name3848 (
		\u11_mem_reg[1][29]/P0001 ,
		_w5951_,
		_w5994_
	);
	LUT2 #(
		.INIT('h8)
	) name3849 (
		\u1_slt6_reg[17]/P0001 ,
		_w3064_,
		_w5995_
	);
	LUT2 #(
		.INIT('h8)
	) name3850 (
		_w5951_,
		_w5995_,
		_w5996_
	);
	LUT2 #(
		.INIT('h1)
	) name3851 (
		_w5994_,
		_w5996_,
		_w5997_
	);
	LUT2 #(
		.INIT('h2)
	) name3852 (
		\u11_mem_reg[1][30]/P0001 ,
		_w5951_,
		_w5998_
	);
	LUT2 #(
		.INIT('h8)
	) name3853 (
		\u1_slt6_reg[18]/P0001 ,
		_w3064_,
		_w5999_
	);
	LUT2 #(
		.INIT('h8)
	) name3854 (
		_w5951_,
		_w5999_,
		_w6000_
	);
	LUT2 #(
		.INIT('h1)
	) name3855 (
		_w5998_,
		_w6000_,
		_w6001_
	);
	LUT2 #(
		.INIT('h2)
	) name3856 (
		\u11_mem_reg[1][31]/P0001 ,
		_w5951_,
		_w6002_
	);
	LUT2 #(
		.INIT('h8)
	) name3857 (
		\u1_slt6_reg[19]/P0001 ,
		_w3064_,
		_w6003_
	);
	LUT2 #(
		.INIT('h8)
	) name3858 (
		_w5951_,
		_w6003_,
		_w6004_
	);
	LUT2 #(
		.INIT('h1)
	) name3859 (
		_w6002_,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h4)
	) name3860 (
		\u11_wp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w6006_
	);
	LUT2 #(
		.INIT('h8)
	) name3861 (
		_w3066_,
		_w6006_,
		_w6007_
	);
	LUT2 #(
		.INIT('h2)
	) name3862 (
		\u11_mem_reg[2][18]/P0001 ,
		_w6007_,
		_w6008_
	);
	LUT2 #(
		.INIT('h4)
	) name3863 (
		_w5938_,
		_w6007_,
		_w6009_
	);
	LUT2 #(
		.INIT('h1)
	) name3864 (
		_w6008_,
		_w6009_,
		_w6010_
	);
	LUT2 #(
		.INIT('h2)
	) name3865 (
		\u11_mem_reg[2][19]/P0001 ,
		_w6007_,
		_w6011_
	);
	LUT2 #(
		.INIT('h4)
	) name3866 (
		_w5944_,
		_w6007_,
		_w6012_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w6011_,
		_w6012_,
		_w6013_
	);
	LUT2 #(
		.INIT('h2)
	) name3868 (
		\u11_mem_reg[2][20]/P0001 ,
		_w6007_,
		_w6014_
	);
	LUT2 #(
		.INIT('h8)
	) name3869 (
		_w5959_,
		_w6007_,
		_w6015_
	);
	LUT2 #(
		.INIT('h1)
	) name3870 (
		_w6014_,
		_w6015_,
		_w6016_
	);
	LUT2 #(
		.INIT('h2)
	) name3871 (
		\u11_mem_reg[2][21]/P0001 ,
		_w6007_,
		_w6017_
	);
	LUT2 #(
		.INIT('h8)
	) name3872 (
		_w5963_,
		_w6007_,
		_w6018_
	);
	LUT2 #(
		.INIT('h1)
	) name3873 (
		_w6017_,
		_w6018_,
		_w6019_
	);
	LUT2 #(
		.INIT('h2)
	) name3874 (
		\u11_mem_reg[2][22]/P0001 ,
		_w6007_,
		_w6020_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		_w5967_,
		_w6007_,
		_w6021_
	);
	LUT2 #(
		.INIT('h1)
	) name3876 (
		_w6020_,
		_w6021_,
		_w6022_
	);
	LUT2 #(
		.INIT('h2)
	) name3877 (
		\u11_mem_reg[2][23]/P0001 ,
		_w6007_,
		_w6023_
	);
	LUT2 #(
		.INIT('h8)
	) name3878 (
		_w5971_,
		_w6007_,
		_w6024_
	);
	LUT2 #(
		.INIT('h1)
	) name3879 (
		_w6023_,
		_w6024_,
		_w6025_
	);
	LUT2 #(
		.INIT('h2)
	) name3880 (
		\u11_mem_reg[2][24]/P0001 ,
		_w6007_,
		_w6026_
	);
	LUT2 #(
		.INIT('h8)
	) name3881 (
		_w5975_,
		_w6007_,
		_w6027_
	);
	LUT2 #(
		.INIT('h1)
	) name3882 (
		_w6026_,
		_w6027_,
		_w6028_
	);
	LUT2 #(
		.INIT('h2)
	) name3883 (
		\u11_mem_reg[2][25]/P0001 ,
		_w6007_,
		_w6029_
	);
	LUT2 #(
		.INIT('h8)
	) name3884 (
		_w5979_,
		_w6007_,
		_w6030_
	);
	LUT2 #(
		.INIT('h1)
	) name3885 (
		_w6029_,
		_w6030_,
		_w6031_
	);
	LUT2 #(
		.INIT('h4)
	) name3886 (
		\u10_wp_reg[2]/P0001 ,
		_w3504_,
		_w6032_
	);
	LUT2 #(
		.INIT('h4)
	) name3887 (
		_w5673_,
		_w6032_,
		_w6033_
	);
	LUT2 #(
		.INIT('h2)
	) name3888 (
		\u10_mem_reg[1][18]/P0001 ,
		_w6032_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name3889 (
		_w6033_,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h2)
	) name3890 (
		\u11_mem_reg[2][26]/P0001 ,
		_w6007_,
		_w6036_
	);
	LUT2 #(
		.INIT('h8)
	) name3891 (
		_w5983_,
		_w6007_,
		_w6037_
	);
	LUT2 #(
		.INIT('h1)
	) name3892 (
		_w6036_,
		_w6037_,
		_w6038_
	);
	LUT2 #(
		.INIT('h2)
	) name3893 (
		\u11_mem_reg[2][27]/P0001 ,
		_w6007_,
		_w6039_
	);
	LUT2 #(
		.INIT('h8)
	) name3894 (
		_w5987_,
		_w6007_,
		_w6040_
	);
	LUT2 #(
		.INIT('h1)
	) name3895 (
		_w6039_,
		_w6040_,
		_w6041_
	);
	LUT2 #(
		.INIT('h4)
	) name3896 (
		_w5679_,
		_w6032_,
		_w6042_
	);
	LUT2 #(
		.INIT('h2)
	) name3897 (
		\u10_mem_reg[1][19]/P0001 ,
		_w6032_,
		_w6043_
	);
	LUT2 #(
		.INIT('h1)
	) name3898 (
		_w6042_,
		_w6043_,
		_w6044_
	);
	LUT2 #(
		.INIT('h2)
	) name3899 (
		\u11_mem_reg[2][28]/P0001 ,
		_w6007_,
		_w6045_
	);
	LUT2 #(
		.INIT('h8)
	) name3900 (
		_w5991_,
		_w6007_,
		_w6046_
	);
	LUT2 #(
		.INIT('h1)
	) name3901 (
		_w6045_,
		_w6046_,
		_w6047_
	);
	LUT2 #(
		.INIT('h2)
	) name3902 (
		\u11_mem_reg[2][29]/P0001 ,
		_w6007_,
		_w6048_
	);
	LUT2 #(
		.INIT('h8)
	) name3903 (
		_w5995_,
		_w6007_,
		_w6049_
	);
	LUT2 #(
		.INIT('h1)
	) name3904 (
		_w6048_,
		_w6049_,
		_w6050_
	);
	LUT2 #(
		.INIT('h2)
	) name3905 (
		\u11_mem_reg[2][30]/P0001 ,
		_w6007_,
		_w6051_
	);
	LUT2 #(
		.INIT('h8)
	) name3906 (
		_w5999_,
		_w6007_,
		_w6052_
	);
	LUT2 #(
		.INIT('h1)
	) name3907 (
		_w6051_,
		_w6052_,
		_w6053_
	);
	LUT2 #(
		.INIT('h2)
	) name3908 (
		\u10_mem_reg[1][20]/P0001 ,
		_w6032_,
		_w6054_
	);
	LUT2 #(
		.INIT('h8)
	) name3909 (
		_w5683_,
		_w6032_,
		_w6055_
	);
	LUT2 #(
		.INIT('h1)
	) name3910 (
		_w6054_,
		_w6055_,
		_w6056_
	);
	LUT2 #(
		.INIT('h2)
	) name3911 (
		\u11_mem_reg[2][31]/P0001 ,
		_w6007_,
		_w6057_
	);
	LUT2 #(
		.INIT('h8)
	) name3912 (
		_w6003_,
		_w6007_,
		_w6058_
	);
	LUT2 #(
		.INIT('h1)
	) name3913 (
		_w6057_,
		_w6058_,
		_w6059_
	);
	LUT2 #(
		.INIT('h2)
	) name3914 (
		\u10_mem_reg[1][21]/P0001 ,
		_w6032_,
		_w6060_
	);
	LUT2 #(
		.INIT('h8)
	) name3915 (
		_w5687_,
		_w6032_,
		_w6061_
	);
	LUT2 #(
		.INIT('h1)
	) name3916 (
		_w6060_,
		_w6061_,
		_w6062_
	);
	LUT2 #(
		.INIT('h2)
	) name3917 (
		\u10_mem_reg[1][22]/P0001 ,
		_w6032_,
		_w6063_
	);
	LUT2 #(
		.INIT('h8)
	) name3918 (
		_w5691_,
		_w6032_,
		_w6064_
	);
	LUT2 #(
		.INIT('h1)
	) name3919 (
		_w6063_,
		_w6064_,
		_w6065_
	);
	LUT2 #(
		.INIT('h2)
	) name3920 (
		\u10_mem_reg[1][23]/P0001 ,
		_w6032_,
		_w6066_
	);
	LUT2 #(
		.INIT('h8)
	) name3921 (
		_w5695_,
		_w6032_,
		_w6067_
	);
	LUT2 #(
		.INIT('h1)
	) name3922 (
		_w6066_,
		_w6067_,
		_w6068_
	);
	LUT2 #(
		.INIT('h2)
	) name3923 (
		\u10_mem_reg[1][24]/P0001 ,
		_w6032_,
		_w6069_
	);
	LUT2 #(
		.INIT('h8)
	) name3924 (
		_w5714_,
		_w6032_,
		_w6070_
	);
	LUT2 #(
		.INIT('h1)
	) name3925 (
		_w6069_,
		_w6070_,
		_w6071_
	);
	LUT2 #(
		.INIT('h2)
	) name3926 (
		\u10_mem_reg[1][25]/P0001 ,
		_w6032_,
		_w6072_
	);
	LUT2 #(
		.INIT('h8)
	) name3927 (
		_w5718_,
		_w6032_,
		_w6073_
	);
	LUT2 #(
		.INIT('h1)
	) name3928 (
		_w6072_,
		_w6073_,
		_w6074_
	);
	LUT2 #(
		.INIT('h2)
	) name3929 (
		\u10_mem_reg[1][26]/P0001 ,
		_w6032_,
		_w6075_
	);
	LUT2 #(
		.INIT('h8)
	) name3930 (
		_w5722_,
		_w6032_,
		_w6076_
	);
	LUT2 #(
		.INIT('h1)
	) name3931 (
		_w6075_,
		_w6076_,
		_w6077_
	);
	LUT2 #(
		.INIT('h2)
	) name3932 (
		\u10_mem_reg[1][27]/P0001 ,
		_w6032_,
		_w6078_
	);
	LUT2 #(
		.INIT('h8)
	) name3933 (
		_w5726_,
		_w6032_,
		_w6079_
	);
	LUT2 #(
		.INIT('h1)
	) name3934 (
		_w6078_,
		_w6079_,
		_w6080_
	);
	LUT2 #(
		.INIT('h2)
	) name3935 (
		\u10_mem_reg[1][28]/P0001 ,
		_w6032_,
		_w6081_
	);
	LUT2 #(
		.INIT('h8)
	) name3936 (
		_w5730_,
		_w6032_,
		_w6082_
	);
	LUT2 #(
		.INIT('h1)
	) name3937 (
		_w6081_,
		_w6082_,
		_w6083_
	);
	LUT2 #(
		.INIT('h2)
	) name3938 (
		\u10_mem_reg[1][29]/P0001 ,
		_w6032_,
		_w6084_
	);
	LUT2 #(
		.INIT('h8)
	) name3939 (
		_w5749_,
		_w6032_,
		_w6085_
	);
	LUT2 #(
		.INIT('h1)
	) name3940 (
		_w6084_,
		_w6085_,
		_w6086_
	);
	LUT2 #(
		.INIT('h2)
	) name3941 (
		_w3068_,
		_w5938_,
		_w6087_
	);
	LUT2 #(
		.INIT('h2)
	) name3942 (
		\u11_mem_reg[3][18]/P0001 ,
		_w3068_,
		_w6088_
	);
	LUT2 #(
		.INIT('h1)
	) name3943 (
		_w6087_,
		_w6088_,
		_w6089_
	);
	LUT2 #(
		.INIT('h2)
	) name3944 (
		_w3068_,
		_w5944_,
		_w6090_
	);
	LUT2 #(
		.INIT('h2)
	) name3945 (
		\u11_mem_reg[3][19]/P0001 ,
		_w3068_,
		_w6091_
	);
	LUT2 #(
		.INIT('h1)
	) name3946 (
		_w6090_,
		_w6091_,
		_w6092_
	);
	LUT2 #(
		.INIT('h2)
	) name3947 (
		\u11_mem_reg[3][20]/P0001 ,
		_w3068_,
		_w6093_
	);
	LUT2 #(
		.INIT('h8)
	) name3948 (
		_w3068_,
		_w5959_,
		_w6094_
	);
	LUT2 #(
		.INIT('h1)
	) name3949 (
		_w6093_,
		_w6094_,
		_w6095_
	);
	LUT2 #(
		.INIT('h2)
	) name3950 (
		\u10_mem_reg[1][30]/P0001 ,
		_w6032_,
		_w6096_
	);
	LUT2 #(
		.INIT('h8)
	) name3951 (
		_w5793_,
		_w6032_,
		_w6097_
	);
	LUT2 #(
		.INIT('h1)
	) name3952 (
		_w6096_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h2)
	) name3953 (
		\u11_mem_reg[3][21]/P0001 ,
		_w3068_,
		_w6099_
	);
	LUT2 #(
		.INIT('h8)
	) name3954 (
		_w3068_,
		_w5963_,
		_w6100_
	);
	LUT2 #(
		.INIT('h1)
	) name3955 (
		_w6099_,
		_w6100_,
		_w6101_
	);
	LUT2 #(
		.INIT('h2)
	) name3956 (
		\u11_mem_reg[3][22]/P0001 ,
		_w3068_,
		_w6102_
	);
	LUT2 #(
		.INIT('h8)
	) name3957 (
		_w3068_,
		_w5967_,
		_w6103_
	);
	LUT2 #(
		.INIT('h1)
	) name3958 (
		_w6102_,
		_w6103_,
		_w6104_
	);
	LUT2 #(
		.INIT('h2)
	) name3959 (
		\u10_mem_reg[1][31]/P0001 ,
		_w6032_,
		_w6105_
	);
	LUT2 #(
		.INIT('h8)
	) name3960 (
		_w5797_,
		_w6032_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name3961 (
		_w6105_,
		_w6106_,
		_w6107_
	);
	LUT2 #(
		.INIT('h2)
	) name3962 (
		\u11_mem_reg[3][23]/P0001 ,
		_w3068_,
		_w6108_
	);
	LUT2 #(
		.INIT('h8)
	) name3963 (
		_w3068_,
		_w5971_,
		_w6109_
	);
	LUT2 #(
		.INIT('h1)
	) name3964 (
		_w6108_,
		_w6109_,
		_w6110_
	);
	LUT2 #(
		.INIT('h2)
	) name3965 (
		\u11_mem_reg[3][24]/P0001 ,
		_w3068_,
		_w6111_
	);
	LUT2 #(
		.INIT('h8)
	) name3966 (
		_w3068_,
		_w5975_,
		_w6112_
	);
	LUT2 #(
		.INIT('h1)
	) name3967 (
		_w6111_,
		_w6112_,
		_w6113_
	);
	LUT2 #(
		.INIT('h2)
	) name3968 (
		\u11_mem_reg[3][25]/P0001 ,
		_w3068_,
		_w6114_
	);
	LUT2 #(
		.INIT('h8)
	) name3969 (
		_w3068_,
		_w5979_,
		_w6115_
	);
	LUT2 #(
		.INIT('h1)
	) name3970 (
		_w6114_,
		_w6115_,
		_w6116_
	);
	LUT2 #(
		.INIT('h2)
	) name3971 (
		\u11_mem_reg[3][26]/P0001 ,
		_w3068_,
		_w6117_
	);
	LUT2 #(
		.INIT('h8)
	) name3972 (
		_w3068_,
		_w5983_,
		_w6118_
	);
	LUT2 #(
		.INIT('h1)
	) name3973 (
		_w6117_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h2)
	) name3974 (
		\u11_mem_reg[3][27]/P0001 ,
		_w3068_,
		_w6120_
	);
	LUT2 #(
		.INIT('h8)
	) name3975 (
		_w3068_,
		_w5987_,
		_w6121_
	);
	LUT2 #(
		.INIT('h1)
	) name3976 (
		_w6120_,
		_w6121_,
		_w6122_
	);
	LUT2 #(
		.INIT('h2)
	) name3977 (
		\u11_mem_reg[3][28]/P0001 ,
		_w3068_,
		_w6123_
	);
	LUT2 #(
		.INIT('h8)
	) name3978 (
		_w3068_,
		_w5991_,
		_w6124_
	);
	LUT2 #(
		.INIT('h1)
	) name3979 (
		_w6123_,
		_w6124_,
		_w6125_
	);
	LUT2 #(
		.INIT('h2)
	) name3980 (
		\u11_mem_reg[3][29]/P0001 ,
		_w3068_,
		_w6126_
	);
	LUT2 #(
		.INIT('h8)
	) name3981 (
		_w3068_,
		_w5995_,
		_w6127_
	);
	LUT2 #(
		.INIT('h1)
	) name3982 (
		_w6126_,
		_w6127_,
		_w6128_
	);
	LUT2 #(
		.INIT('h2)
	) name3983 (
		\u11_mem_reg[3][30]/P0001 ,
		_w3068_,
		_w6129_
	);
	LUT2 #(
		.INIT('h8)
	) name3984 (
		_w3068_,
		_w5999_,
		_w6130_
	);
	LUT2 #(
		.INIT('h1)
	) name3985 (
		_w6129_,
		_w6130_,
		_w6131_
	);
	LUT2 #(
		.INIT('h2)
	) name3986 (
		\u11_mem_reg[3][31]/P0001 ,
		_w3068_,
		_w6132_
	);
	LUT2 #(
		.INIT('h8)
	) name3987 (
		_w3068_,
		_w6003_,
		_w6133_
	);
	LUT2 #(
		.INIT('h1)
	) name3988 (
		_w6132_,
		_w6133_,
		_w6134_
	);
	LUT2 #(
		.INIT('h2)
	) name3989 (
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w6135_
	);
	LUT2 #(
		.INIT('h8)
	) name3990 (
		\u15_crac_wr_reg/NET0131 ,
		_w6135_,
		_w6136_
	);
	LUT2 #(
		.INIT('h1)
	) name3991 (
		\u13_ints_r_reg[1]/NET0131 ,
		_w6136_,
		_w6137_
	);
	LUT2 #(
		.INIT('h1)
	) name3992 (
		_w2743_,
		_w6137_,
		_w6138_
	);
	LUT2 #(
		.INIT('h2)
	) name3993 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w6139_
	);
	LUT2 #(
		.INIT('h8)
	) name3994 (
		\wb_addr_i[3]_pad ,
		\wb_addr_i[4]_pad ,
		_w6140_
	);
	LUT2 #(
		.INIT('h8)
	) name3995 (
		_w6139_,
		_w6140_,
		_w6141_
	);
	LUT2 #(
		.INIT('h1)
	) name3996 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w6142_
	);
	LUT2 #(
		.INIT('h4)
	) name3997 (
		\wb_addr_i[4]_pad ,
		_w6142_,
		_w6143_
	);
	LUT2 #(
		.INIT('h4)
	) name3998 (
		\wb_addr_i[5]_pad ,
		\wb_addr_i[6]_pad ,
		_w6144_
	);
	LUT2 #(
		.INIT('h8)
	) name3999 (
		_w6143_,
		_w6144_,
		_w6145_
	);
	LUT2 #(
		.INIT('h1)
	) name4000 (
		_w6141_,
		_w6145_,
		_w6146_
	);
	LUT2 #(
		.INIT('h4)
	) name4001 (
		\wb_addr_i[4]_pad ,
		_w2740_,
		_w6147_
	);
	LUT2 #(
		.INIT('h8)
	) name4002 (
		\u13_occ1_r_reg[1]/NET0131 ,
		_w6147_,
		_w6148_
	);
	LUT2 #(
		.INIT('h8)
	) name4003 (
		\u13_ints_r_reg[1]/NET0131 ,
		_w2741_,
		_w6149_
	);
	LUT2 #(
		.INIT('h2)
	) name4004 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w6150_
	);
	LUT2 #(
		.INIT('h4)
	) name4005 (
		\wb_addr_i[4]_pad ,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h8)
	) name4006 (
		\u13_occ0_r_reg[1]/NET0131 ,
		_w6151_,
		_w6152_
	);
	LUT2 #(
		.INIT('h8)
	) name4007 (
		\wb_addr_i[4]_pad ,
		_w6150_,
		_w6153_
	);
	LUT2 #(
		.INIT('h8)
	) name4008 (
		\u13_intm_r_reg[1]/NET0131 ,
		_w6153_,
		_w6154_
	);
	LUT2 #(
		.INIT('h8)
	) name4009 (
		suspended_o_pad,
		_w6143_,
		_w6155_
	);
	LUT2 #(
		.INIT('h8)
	) name4010 (
		\wb_addr_i[2]_pad ,
		\wb_addr_i[3]_pad ,
		_w6156_
	);
	LUT2 #(
		.INIT('h4)
	) name4011 (
		\wb_addr_i[4]_pad ,
		_w6156_,
		_w6157_
	);
	LUT2 #(
		.INIT('h8)
	) name4012 (
		\u13_icc_r_reg[1]/NET0131 ,
		_w6157_,
		_w6158_
	);
	LUT2 #(
		.INIT('h8)
	) name4013 (
		\wb_addr_i[4]_pad ,
		_w6142_,
		_w6159_
	);
	LUT2 #(
		.INIT('h8)
	) name4014 (
		\u15_crac_din_reg[1]/NET0131 ,
		_w6159_,
		_w6160_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w6148_,
		_w6149_,
		_w6161_
	);
	LUT2 #(
		.INIT('h1)
	) name4016 (
		_w6152_,
		_w6154_,
		_w6162_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		_w6155_,
		_w6158_,
		_w6163_
	);
	LUT2 #(
		.INIT('h4)
	) name4018 (
		_w6160_,
		_w6163_,
		_w6164_
	);
	LUT2 #(
		.INIT('h8)
	) name4019 (
		_w6161_,
		_w6162_,
		_w6165_
	);
	LUT2 #(
		.INIT('h8)
	) name4020 (
		_w6164_,
		_w6165_,
		_w6166_
	);
	LUT2 #(
		.INIT('h2)
	) name4021 (
		_w6146_,
		_w6166_,
		_w6167_
	);
	LUT2 #(
		.INIT('h4)
	) name4022 (
		\wb_addr_i[2]_pad ,
		_w6141_,
		_w6168_
	);
	LUT2 #(
		.INIT('h8)
	) name4023 (
		\u9_dout_reg[1]/P0001 ,
		_w6168_,
		_w6169_
	);
	LUT2 #(
		.INIT('h8)
	) name4024 (
		\wb_addr_i[2]_pad ,
		_w6141_,
		_w6170_
	);
	LUT2 #(
		.INIT('h8)
	) name4025 (
		\u10_dout_reg[1]/P0001 ,
		_w6170_,
		_w6171_
	);
	LUT2 #(
		.INIT('h8)
	) name4026 (
		\u11_dout_reg[1]/P0001 ,
		_w6145_,
		_w6172_
	);
	LUT2 #(
		.INIT('h1)
	) name4027 (
		_w6169_,
		_w6171_,
		_w6173_
	);
	LUT2 #(
		.INIT('h4)
	) name4028 (
		_w6172_,
		_w6173_,
		_w6174_
	);
	LUT2 #(
		.INIT('h4)
	) name4029 (
		_w6167_,
		_w6174_,
		_w6175_
	);
	LUT2 #(
		.INIT('h8)
	) name4030 (
		\u26_cnt_reg[0]/NET0131 ,
		_w5629_,
		_w6176_
	);
	LUT2 #(
		.INIT('h1)
	) name4031 (
		\u26_cnt_reg[0]/NET0131 ,
		\u26_cnt_reg[1]/NET0131 ,
		_w6177_
	);
	LUT2 #(
		.INIT('h8)
	) name4032 (
		\u26_cnt_reg[2]/NET0131 ,
		_w6177_,
		_w6178_
	);
	LUT2 #(
		.INIT('h2)
	) name4033 (
		_w5629_,
		_w6178_,
		_w6179_
	);
	LUT2 #(
		.INIT('h1)
	) name4034 (
		\u26_cnt_reg[0]/NET0131 ,
		_w6179_,
		_w6180_
	);
	LUT2 #(
		.INIT('h1)
	) name4035 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w6176_,
		_w6181_
	);
	LUT2 #(
		.INIT('h4)
	) name4036 (
		_w6180_,
		_w6181_,
		_w6182_
	);
	LUT2 #(
		.INIT('h1)
	) name4037 (
		\u26_cnt_reg[1]/NET0131 ,
		_w6176_,
		_w6183_
	);
	LUT2 #(
		.INIT('h8)
	) name4038 (
		\u26_cnt_reg[1]/NET0131 ,
		_w6176_,
		_w6184_
	);
	LUT2 #(
		.INIT('h1)
	) name4039 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w6183_,
		_w6185_
	);
	LUT2 #(
		.INIT('h4)
	) name4040 (
		_w6184_,
		_w6185_,
		_w6186_
	);
	LUT2 #(
		.INIT('h1)
	) name4041 (
		\u26_cnt_reg[2]/NET0131 ,
		_w6184_,
		_w6187_
	);
	LUT2 #(
		.INIT('h8)
	) name4042 (
		\u26_cnt_reg[2]/NET0131 ,
		_w6184_,
		_w6188_
	);
	LUT2 #(
		.INIT('h1)
	) name4043 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w6187_,
		_w6189_
	);
	LUT2 #(
		.INIT('h4)
	) name4044 (
		_w6188_,
		_w6189_,
		_w6190_
	);
	LUT2 #(
		.INIT('h8)
	) name4045 (
		\u3_empty_reg/NET0131 ,
		_w2787_,
		_w6191_
	);
	LUT2 #(
		.INIT('h1)
	) name4046 (
		\u17_int_set_reg[1]/NET0131 ,
		_w6191_,
		_w6192_
	);
	LUT2 #(
		.INIT('h8)
	) name4047 (
		\u4_empty_reg/NET0131 ,
		_w2759_,
		_w6193_
	);
	LUT2 #(
		.INIT('h1)
	) name4048 (
		\u18_int_set_reg[1]/NET0131 ,
		_w6193_,
		_w6194_
	);
	LUT2 #(
		.INIT('h8)
	) name4049 (
		\u5_empty_reg/NET0131 ,
		_w2770_,
		_w6195_
	);
	LUT2 #(
		.INIT('h1)
	) name4050 (
		\u19_int_set_reg[1]/NET0131 ,
		_w6195_,
		_w6196_
	);
	LUT2 #(
		.INIT('h8)
	) name4051 (
		\u6_empty_reg/NET0131 ,
		_w2795_,
		_w6197_
	);
	LUT2 #(
		.INIT('h1)
	) name4052 (
		\u20_int_set_reg[1]/NET0131 ,
		_w6197_,
		_w6198_
	);
	LUT2 #(
		.INIT('h8)
	) name4053 (
		\u7_empty_reg/NET0131 ,
		_w2808_,
		_w6199_
	);
	LUT2 #(
		.INIT('h1)
	) name4054 (
		\u21_int_set_reg[1]/NET0131 ,
		_w6199_,
		_w6200_
	);
	LUT2 #(
		.INIT('h8)
	) name4055 (
		\u8_empty_reg/NET0131 ,
		_w2159_,
		_w6201_
	);
	LUT2 #(
		.INIT('h1)
	) name4056 (
		\u22_int_set_reg[1]/NET0131 ,
		_w6201_,
		_w6202_
	);
	LUT2 #(
		.INIT('h8)
	) name4057 (
		\u9_full_reg/NET0131 ,
		_w3310_,
		_w6203_
	);
	LUT2 #(
		.INIT('h1)
	) name4058 (
		\u23_int_set_reg[2]/NET0131 ,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h8)
	) name4059 (
		\u10_full_reg/NET0131 ,
		_w3500_,
		_w6205_
	);
	LUT2 #(
		.INIT('h1)
	) name4060 (
		\u24_int_set_reg[2]/NET0131 ,
		_w6205_,
		_w6206_
	);
	LUT2 #(
		.INIT('h8)
	) name4061 (
		\u11_full_reg/NET0131 ,
		_w3063_,
		_w6207_
	);
	LUT2 #(
		.INIT('h1)
	) name4062 (
		\u25_int_set_reg[2]/NET0131 ,
		_w6207_,
		_w6208_
	);
	LUT2 #(
		.INIT('h1)
	) name4063 (
		\ac97_reset_pad_o__pad ,
		_w6178_,
		_w6209_
	);
	LUT2 #(
		.INIT('h1)
	) name4064 (
		\u13_ac97_rst_force_reg/P0001 ,
		_w6209_,
		_w6210_
	);
	LUT2 #(
		.INIT('h4)
	) name4065 (
		\u13_crac_r_reg[7]/NET0131 ,
		\u15_crac_we_r_reg/P0001 ,
		_w6211_
	);
	LUT2 #(
		.INIT('h2)
	) name4066 (
		\u15_crac_wr_reg/NET0131 ,
		_w6135_,
		_w6212_
	);
	LUT2 #(
		.INIT('h1)
	) name4067 (
		_w6211_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h8)
	) name4068 (
		\u13_crac_r_reg[7]/NET0131 ,
		\u15_crac_we_r_reg/P0001 ,
		_w6214_
	);
	LUT2 #(
		.INIT('h4)
	) name4069 (
		\u15_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w6215_
	);
	LUT2 #(
		.INIT('h8)
	) name4070 (
		\u15_rdd1_reg/NET0131 ,
		_w6215_,
		_w6216_
	);
	LUT2 #(
		.INIT('h2)
	) name4071 (
		\u15_crac_rd_reg/NET0131 ,
		_w6216_,
		_w6217_
	);
	LUT2 #(
		.INIT('h1)
	) name4072 (
		_w6214_,
		_w6217_,
		_w6218_
	);
	LUT2 #(
		.INIT('h8)
	) name4073 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[2]/P0001 ,
		_w6219_
	);
	LUT2 #(
		.INIT('h2)
	) name4074 (
		\u0_slt9_r_reg[1]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w6220_
	);
	LUT2 #(
		.INIT('h1)
	) name4075 (
		_w6219_,
		_w6220_,
		_w6221_
	);
	LUT2 #(
		.INIT('h1)
	) name4076 (
		\u3_rp_reg[3]/NET0131 ,
		\u3_wp_reg[2]/P0001 ,
		_w6222_
	);
	LUT2 #(
		.INIT('h8)
	) name4077 (
		\u3_rp_reg[3]/NET0131 ,
		\u3_wp_reg[2]/P0001 ,
		_w6223_
	);
	LUT2 #(
		.INIT('h1)
	) name4078 (
		_w6222_,
		_w6223_,
		_w6224_
	);
	LUT2 #(
		.INIT('h4)
	) name4079 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		_w6225_
	);
	LUT2 #(
		.INIT('h2)
	) name4080 (
		\u3_rp_reg[2]/NET0131 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6226_
	);
	LUT2 #(
		.INIT('h4)
	) name4081 (
		\u3_rp_reg[2]/NET0131 ,
		\u3_wp_reg[1]/NET0131 ,
		_w6227_
	);
	LUT2 #(
		.INIT('h1)
	) name4082 (
		_w6226_,
		_w6227_,
		_w6228_
	);
	LUT2 #(
		.INIT('h4)
	) name4083 (
		_w6225_,
		_w6228_,
		_w6229_
	);
	LUT2 #(
		.INIT('h2)
	) name4084 (
		\u3_rp_reg[1]/NET0131 ,
		\u3_wp_reg[0]/P0001 ,
		_w6230_
	);
	LUT2 #(
		.INIT('h2)
	) name4085 (
		\u12_o3_we_reg/P0001 ,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h8)
	) name4086 (
		_w6224_,
		_w6231_,
		_w6232_
	);
	LUT2 #(
		.INIT('h8)
	) name4087 (
		_w6229_,
		_w6232_,
		_w6233_
	);
	LUT2 #(
		.INIT('h1)
	) name4088 (
		\u17_int_set_reg[2]/NET0131 ,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h2)
	) name4089 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		_w6235_
	);
	LUT2 #(
		.INIT('h4)
	) name4090 (
		\u4_rp_reg[1]/NET0131 ,
		\u4_wp_reg[0]/P0001 ,
		_w6236_
	);
	LUT2 #(
		.INIT('h2)
	) name4091 (
		\u4_rp_reg[2]/NET0131 ,
		\u4_wp_reg[1]/NET0131 ,
		_w6237_
	);
	LUT2 #(
		.INIT('h4)
	) name4092 (
		\u4_rp_reg[2]/NET0131 ,
		\u4_wp_reg[1]/NET0131 ,
		_w6238_
	);
	LUT2 #(
		.INIT('h1)
	) name4093 (
		_w6237_,
		_w6238_,
		_w6239_
	);
	LUT2 #(
		.INIT('h4)
	) name4094 (
		_w6236_,
		_w6239_,
		_w6240_
	);
	LUT2 #(
		.INIT('h1)
	) name4095 (
		\u4_rp_reg[3]/NET0131 ,
		\u4_wp_reg[2]/P0001 ,
		_w6241_
	);
	LUT2 #(
		.INIT('h8)
	) name4096 (
		\u4_rp_reg[3]/NET0131 ,
		\u4_wp_reg[2]/P0001 ,
		_w6242_
	);
	LUT2 #(
		.INIT('h1)
	) name4097 (
		_w6241_,
		_w6242_,
		_w6243_
	);
	LUT2 #(
		.INIT('h2)
	) name4098 (
		\u12_o4_we_reg/P0001 ,
		_w6235_,
		_w6244_
	);
	LUT2 #(
		.INIT('h8)
	) name4099 (
		_w6243_,
		_w6244_,
		_w6245_
	);
	LUT2 #(
		.INIT('h8)
	) name4100 (
		_w6240_,
		_w6245_,
		_w6246_
	);
	LUT2 #(
		.INIT('h1)
	) name4101 (
		\u18_int_set_reg[2]/NET0131 ,
		_w6246_,
		_w6247_
	);
	LUT2 #(
		.INIT('h2)
	) name4102 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		_w6248_
	);
	LUT2 #(
		.INIT('h4)
	) name4103 (
		\u5_rp_reg[1]/NET0131 ,
		\u5_wp_reg[0]/P0001 ,
		_w6249_
	);
	LUT2 #(
		.INIT('h2)
	) name4104 (
		\u5_rp_reg[2]/NET0131 ,
		\u5_wp_reg[1]/NET0131 ,
		_w6250_
	);
	LUT2 #(
		.INIT('h4)
	) name4105 (
		\u5_rp_reg[2]/NET0131 ,
		\u5_wp_reg[1]/NET0131 ,
		_w6251_
	);
	LUT2 #(
		.INIT('h1)
	) name4106 (
		_w6250_,
		_w6251_,
		_w6252_
	);
	LUT2 #(
		.INIT('h4)
	) name4107 (
		_w6249_,
		_w6252_,
		_w6253_
	);
	LUT2 #(
		.INIT('h1)
	) name4108 (
		\u5_rp_reg[3]/NET0131 ,
		\u5_wp_reg[2]/P0001 ,
		_w6254_
	);
	LUT2 #(
		.INIT('h8)
	) name4109 (
		\u5_rp_reg[3]/NET0131 ,
		\u5_wp_reg[2]/P0001 ,
		_w6255_
	);
	LUT2 #(
		.INIT('h1)
	) name4110 (
		_w6254_,
		_w6255_,
		_w6256_
	);
	LUT2 #(
		.INIT('h2)
	) name4111 (
		\u12_o6_we_reg/P0001 ,
		_w6248_,
		_w6257_
	);
	LUT2 #(
		.INIT('h8)
	) name4112 (
		_w6256_,
		_w6257_,
		_w6258_
	);
	LUT2 #(
		.INIT('h8)
	) name4113 (
		_w6253_,
		_w6258_,
		_w6259_
	);
	LUT2 #(
		.INIT('h1)
	) name4114 (
		\u19_int_set_reg[2]/NET0131 ,
		_w6259_,
		_w6260_
	);
	LUT2 #(
		.INIT('h4)
	) name4115 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		_w6261_
	);
	LUT2 #(
		.INIT('h2)
	) name4116 (
		\u6_rp_reg[1]/NET0131 ,
		\u6_wp_reg[0]/P0001 ,
		_w6262_
	);
	LUT2 #(
		.INIT('h1)
	) name4117 (
		_w6261_,
		_w6262_,
		_w6263_
	);
	LUT2 #(
		.INIT('h2)
	) name4118 (
		\u6_rp_reg[2]/NET0131 ,
		\u6_wp_reg[1]/NET0131 ,
		_w6264_
	);
	LUT2 #(
		.INIT('h4)
	) name4119 (
		\u6_rp_reg[2]/NET0131 ,
		\u6_wp_reg[1]/NET0131 ,
		_w6265_
	);
	LUT2 #(
		.INIT('h1)
	) name4120 (
		_w6264_,
		_w6265_,
		_w6266_
	);
	LUT2 #(
		.INIT('h8)
	) name4121 (
		_w6263_,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h1)
	) name4122 (
		\u6_rp_reg[3]/NET0131 ,
		\u6_wp_reg[2]/P0001 ,
		_w6268_
	);
	LUT2 #(
		.INIT('h8)
	) name4123 (
		\u6_rp_reg[3]/NET0131 ,
		\u6_wp_reg[2]/P0001 ,
		_w6269_
	);
	LUT2 #(
		.INIT('h1)
	) name4124 (
		_w6268_,
		_w6269_,
		_w6270_
	);
	LUT2 #(
		.INIT('h8)
	) name4125 (
		\u12_o7_we_reg/P0001 ,
		_w6270_,
		_w6271_
	);
	LUT2 #(
		.INIT('h8)
	) name4126 (
		_w6267_,
		_w6271_,
		_w6272_
	);
	LUT2 #(
		.INIT('h1)
	) name4127 (
		\u20_int_set_reg[2]/NET0131 ,
		_w6272_,
		_w6273_
	);
	LUT2 #(
		.INIT('h1)
	) name4128 (
		\u7_rp_reg[3]/NET0131 ,
		\u7_wp_reg[2]/P0001 ,
		_w6274_
	);
	LUT2 #(
		.INIT('h8)
	) name4129 (
		\u7_rp_reg[3]/NET0131 ,
		\u7_wp_reg[2]/P0001 ,
		_w6275_
	);
	LUT2 #(
		.INIT('h1)
	) name4130 (
		_w6274_,
		_w6275_,
		_w6276_
	);
	LUT2 #(
		.INIT('h4)
	) name4131 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		_w6277_
	);
	LUT2 #(
		.INIT('h2)
	) name4132 (
		\u7_rp_reg[2]/NET0131 ,
		\u7_wp_reg[1]/NET0131 ,
		_w6278_
	);
	LUT2 #(
		.INIT('h4)
	) name4133 (
		\u7_rp_reg[2]/NET0131 ,
		\u7_wp_reg[1]/NET0131 ,
		_w6279_
	);
	LUT2 #(
		.INIT('h1)
	) name4134 (
		_w6278_,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h4)
	) name4135 (
		_w6277_,
		_w6280_,
		_w6281_
	);
	LUT2 #(
		.INIT('h2)
	) name4136 (
		\u7_rp_reg[1]/NET0131 ,
		\u7_wp_reg[0]/P0001 ,
		_w6282_
	);
	LUT2 #(
		.INIT('h2)
	) name4137 (
		\u12_o8_we_reg/P0001 ,
		_w6282_,
		_w6283_
	);
	LUT2 #(
		.INIT('h8)
	) name4138 (
		_w6276_,
		_w6283_,
		_w6284_
	);
	LUT2 #(
		.INIT('h8)
	) name4139 (
		_w6281_,
		_w6284_,
		_w6285_
	);
	LUT2 #(
		.INIT('h1)
	) name4140 (
		\u21_int_set_reg[2]/NET0131 ,
		_w6285_,
		_w6286_
	);
	LUT2 #(
		.INIT('h4)
	) name4141 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		_w6287_
	);
	LUT2 #(
		.INIT('h2)
	) name4142 (
		\u8_rp_reg[1]/NET0131 ,
		\u8_wp_reg[0]/P0001 ,
		_w6288_
	);
	LUT2 #(
		.INIT('h1)
	) name4143 (
		_w6287_,
		_w6288_,
		_w6289_
	);
	LUT2 #(
		.INIT('h2)
	) name4144 (
		\u8_rp_reg[2]/NET0131 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6290_
	);
	LUT2 #(
		.INIT('h4)
	) name4145 (
		\u8_rp_reg[2]/NET0131 ,
		\u8_wp_reg[1]/NET0131 ,
		_w6291_
	);
	LUT2 #(
		.INIT('h1)
	) name4146 (
		_w6290_,
		_w6291_,
		_w6292_
	);
	LUT2 #(
		.INIT('h8)
	) name4147 (
		_w6289_,
		_w6292_,
		_w6293_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		\u8_rp_reg[3]/NET0131 ,
		\u8_wp_reg[2]/P0001 ,
		_w6294_
	);
	LUT2 #(
		.INIT('h8)
	) name4149 (
		\u8_rp_reg[3]/NET0131 ,
		\u8_wp_reg[2]/P0001 ,
		_w6295_
	);
	LUT2 #(
		.INIT('h1)
	) name4150 (
		_w6294_,
		_w6295_,
		_w6296_
	);
	LUT2 #(
		.INIT('h8)
	) name4151 (
		\u12_o9_we_reg/P0001 ,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h8)
	) name4152 (
		_w6293_,
		_w6297_,
		_w6298_
	);
	LUT2 #(
		.INIT('h1)
	) name4153 (
		\u22_int_set_reg[2]/NET0131 ,
		_w6298_,
		_w6299_
	);
	LUT2 #(
		.INIT('h8)
	) name4154 (
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		_w6300_
	);
	LUT2 #(
		.INIT('h8)
	) name4155 (
		\u8_wp_reg[1]/NET0131 ,
		_w6300_,
		_w6301_
	);
	LUT2 #(
		.INIT('h1)
	) name4156 (
		\u8_wp_reg[2]/P0001 ,
		_w6301_,
		_w6302_
	);
	LUT2 #(
		.INIT('h8)
	) name4157 (
		\u8_wp_reg[2]/P0001 ,
		_w6301_,
		_w6303_
	);
	LUT2 #(
		.INIT('h2)
	) name4158 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w6302_,
		_w6304_
	);
	LUT2 #(
		.INIT('h4)
	) name4159 (
		_w6303_,
		_w6304_,
		_w6305_
	);
	LUT2 #(
		.INIT('h8)
	) name4160 (
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		_w6306_
	);
	LUT2 #(
		.INIT('h8)
	) name4161 (
		\u4_wp_reg[1]/NET0131 ,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h1)
	) name4162 (
		\u4_wp_reg[2]/P0001 ,
		_w6307_,
		_w6308_
	);
	LUT2 #(
		.INIT('h8)
	) name4163 (
		\u4_wp_reg[2]/P0001 ,
		_w6307_,
		_w6309_
	);
	LUT2 #(
		.INIT('h2)
	) name4164 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w6308_,
		_w6310_
	);
	LUT2 #(
		.INIT('h4)
	) name4165 (
		_w6309_,
		_w6310_,
		_w6311_
	);
	LUT2 #(
		.INIT('h8)
	) name4166 (
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		_w6312_
	);
	LUT2 #(
		.INIT('h8)
	) name4167 (
		\u5_wp_reg[1]/NET0131 ,
		_w6312_,
		_w6313_
	);
	LUT2 #(
		.INIT('h1)
	) name4168 (
		\u5_wp_reg[2]/P0001 ,
		_w6313_,
		_w6314_
	);
	LUT2 #(
		.INIT('h8)
	) name4169 (
		\u5_wp_reg[2]/P0001 ,
		_w6313_,
		_w6315_
	);
	LUT2 #(
		.INIT('h2)
	) name4170 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w6314_,
		_w6316_
	);
	LUT2 #(
		.INIT('h4)
	) name4171 (
		_w6315_,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h8)
	) name4172 (
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		_w6318_
	);
	LUT2 #(
		.INIT('h8)
	) name4173 (
		\u3_wp_reg[1]/NET0131 ,
		_w6318_,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name4174 (
		\u3_wp_reg[2]/P0001 ,
		_w6319_,
		_w6320_
	);
	LUT2 #(
		.INIT('h8)
	) name4175 (
		\u3_wp_reg[2]/P0001 ,
		_w6319_,
		_w6321_
	);
	LUT2 #(
		.INIT('h2)
	) name4176 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w6320_,
		_w6322_
	);
	LUT2 #(
		.INIT('h4)
	) name4177 (
		_w6321_,
		_w6322_,
		_w6323_
	);
	LUT2 #(
		.INIT('h8)
	) name4178 (
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		_w6324_
	);
	LUT2 #(
		.INIT('h8)
	) name4179 (
		\u6_wp_reg[1]/NET0131 ,
		_w6324_,
		_w6325_
	);
	LUT2 #(
		.INIT('h1)
	) name4180 (
		\u6_wp_reg[2]/P0001 ,
		_w6325_,
		_w6326_
	);
	LUT2 #(
		.INIT('h8)
	) name4181 (
		\u6_wp_reg[2]/P0001 ,
		_w6325_,
		_w6327_
	);
	LUT2 #(
		.INIT('h2)
	) name4182 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w6326_,
		_w6328_
	);
	LUT2 #(
		.INIT('h4)
	) name4183 (
		_w6327_,
		_w6328_,
		_w6329_
	);
	LUT2 #(
		.INIT('h8)
	) name4184 (
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		_w6330_
	);
	LUT2 #(
		.INIT('h8)
	) name4185 (
		\u7_wp_reg[1]/NET0131 ,
		_w6330_,
		_w6331_
	);
	LUT2 #(
		.INIT('h1)
	) name4186 (
		\u7_wp_reg[2]/P0001 ,
		_w6331_,
		_w6332_
	);
	LUT2 #(
		.INIT('h8)
	) name4187 (
		\u7_wp_reg[2]/P0001 ,
		_w6331_,
		_w6333_
	);
	LUT2 #(
		.INIT('h2)
	) name4188 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w6332_,
		_w6334_
	);
	LUT2 #(
		.INIT('h4)
	) name4189 (
		_w6333_,
		_w6334_,
		_w6335_
	);
	LUT2 #(
		.INIT('h4)
	) name4190 (
		\u11_wp_reg[0]/NET0131 ,
		_w3063_,
		_w6336_
	);
	LUT2 #(
		.INIT('h4)
	) name4191 (
		\u9_wp_reg[0]/NET0131 ,
		_w3310_,
		_w6337_
	);
	LUT2 #(
		.INIT('h4)
	) name4192 (
		\u10_wp_reg[0]/NET0131 ,
		_w3500_,
		_w6338_
	);
	LUT2 #(
		.INIT('h8)
	) name4193 (
		\u14_u0_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6339_
	);
	LUT2 #(
		.INIT('h1)
	) name4194 (
		\u14_u0_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6340_
	);
	LUT2 #(
		.INIT('h8)
	) name4195 (
		\u13_occ0_r_reg[1]/NET0131 ,
		\u1_slt1_reg[11]/P0001 ,
		_w6341_
	);
	LUT2 #(
		.INIT('h2)
	) name4196 (
		\u13_occ0_r_reg[0]/NET0131 ,
		\u14_u0_full_empty_r_reg/P0001 ,
		_w6342_
	);
	LUT2 #(
		.INIT('h8)
	) name4197 (
		\u1_slt0_reg[15]/P0001 ,
		_w6342_,
		_w6343_
	);
	LUT2 #(
		.INIT('h1)
	) name4198 (
		_w6340_,
		_w6341_,
		_w6344_
	);
	LUT2 #(
		.INIT('h8)
	) name4199 (
		_w6343_,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h1)
	) name4200 (
		_w6339_,
		_w6345_,
		_w6346_
	);
	LUT2 #(
		.INIT('h1)
	) name4201 (
		\u14_u1_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6347_
	);
	LUT2 #(
		.INIT('h8)
	) name4202 (
		\u13_occ0_r_reg[9]/NET0131 ,
		\u1_slt1_reg[10]/P0001 ,
		_w6348_
	);
	LUT2 #(
		.INIT('h2)
	) name4203 (
		\u13_occ0_r_reg[8]/NET0131 ,
		\u14_u1_full_empty_r_reg/P0001 ,
		_w6349_
	);
	LUT2 #(
		.INIT('h8)
	) name4204 (
		\u1_slt0_reg[15]/P0001 ,
		_w6349_,
		_w6350_
	);
	LUT2 #(
		.INIT('h1)
	) name4205 (
		_w6347_,
		_w6348_,
		_w6351_
	);
	LUT2 #(
		.INIT('h8)
	) name4206 (
		_w6350_,
		_w6351_,
		_w6352_
	);
	LUT2 #(
		.INIT('h1)
	) name4207 (
		_w2758_,
		_w6352_,
		_w6353_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		\u14_u2_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6354_
	);
	LUT2 #(
		.INIT('h8)
	) name4209 (
		\u13_occ0_r_reg[17]/NET0131 ,
		\u1_slt1_reg[8]/P0001 ,
		_w6355_
	);
	LUT2 #(
		.INIT('h2)
	) name4210 (
		\u13_occ0_r_reg[16]/NET0131 ,
		\u14_u2_full_empty_r_reg/P0001 ,
		_w6356_
	);
	LUT2 #(
		.INIT('h8)
	) name4211 (
		\u1_slt0_reg[15]/P0001 ,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h1)
	) name4212 (
		_w6354_,
		_w6355_,
		_w6358_
	);
	LUT2 #(
		.INIT('h8)
	) name4213 (
		_w6357_,
		_w6358_,
		_w6359_
	);
	LUT2 #(
		.INIT('h1)
	) name4214 (
		_w2769_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h1)
	) name4215 (
		\u14_u3_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6361_
	);
	LUT2 #(
		.INIT('h8)
	) name4216 (
		\u13_occ0_r_reg[25]/NET0131 ,
		\u1_slt1_reg[7]/P0001 ,
		_w6362_
	);
	LUT2 #(
		.INIT('h2)
	) name4217 (
		\u13_occ0_r_reg[24]/NET0131 ,
		\u14_u3_full_empty_r_reg/P0001 ,
		_w6363_
	);
	LUT2 #(
		.INIT('h8)
	) name4218 (
		\u1_slt0_reg[15]/P0001 ,
		_w6363_,
		_w6364_
	);
	LUT2 #(
		.INIT('h1)
	) name4219 (
		_w6361_,
		_w6362_,
		_w6365_
	);
	LUT2 #(
		.INIT('h8)
	) name4220 (
		_w6364_,
		_w6365_,
		_w6366_
	);
	LUT2 #(
		.INIT('h1)
	) name4221 (
		_w2794_,
		_w6366_,
		_w6367_
	);
	LUT2 #(
		.INIT('h1)
	) name4222 (
		\u14_u4_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6368_
	);
	LUT2 #(
		.INIT('h8)
	) name4223 (
		\u13_occ1_r_reg[1]/NET0131 ,
		\u1_slt1_reg[6]/P0001 ,
		_w6369_
	);
	LUT2 #(
		.INIT('h2)
	) name4224 (
		\u13_occ1_r_reg[0]/NET0131 ,
		\u14_u4_full_empty_r_reg/P0001 ,
		_w6370_
	);
	LUT2 #(
		.INIT('h8)
	) name4225 (
		\u1_slt0_reg[15]/P0001 ,
		_w6370_,
		_w6371_
	);
	LUT2 #(
		.INIT('h1)
	) name4226 (
		_w6368_,
		_w6369_,
		_w6372_
	);
	LUT2 #(
		.INIT('h8)
	) name4227 (
		_w6371_,
		_w6372_,
		_w6373_
	);
	LUT2 #(
		.INIT('h1)
	) name4228 (
		_w2807_,
		_w6373_,
		_w6374_
	);
	LUT2 #(
		.INIT('h1)
	) name4229 (
		\u14_u5_en_out_l_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6375_
	);
	LUT2 #(
		.INIT('h8)
	) name4230 (
		\u13_occ1_r_reg[9]/NET0131 ,
		\u1_slt1_reg[5]/P0001 ,
		_w6376_
	);
	LUT2 #(
		.INIT('h2)
	) name4231 (
		\u13_occ1_r_reg[8]/NET0131 ,
		\u14_u5_full_empty_r_reg/P0001 ,
		_w6377_
	);
	LUT2 #(
		.INIT('h8)
	) name4232 (
		\u1_slt0_reg[15]/P0001 ,
		_w6377_,
		_w6378_
	);
	LUT2 #(
		.INIT('h1)
	) name4233 (
		_w6375_,
		_w6376_,
		_w6379_
	);
	LUT2 #(
		.INIT('h8)
	) name4234 (
		_w6378_,
		_w6379_,
		_w6380_
	);
	LUT2 #(
		.INIT('h1)
	) name4235 (
		_w2158_,
		_w6380_,
		_w6381_
	);
	LUT2 #(
		.INIT('h1)
	) name4236 (
		\in_valid_s_reg[0]/NET0131 ,
		\u14_u6_en_out_l_reg/NET0131 ,
		_w6382_
	);
	LUT2 #(
		.INIT('h2)
	) name4237 (
		\u13_icc_r_reg[1]/NET0131 ,
		\u1_slt0_reg[12]/P0001 ,
		_w6383_
	);
	LUT2 #(
		.INIT('h2)
	) name4238 (
		\u13_icc_r_reg[0]/NET0131 ,
		\u14_u6_full_empty_r_reg/P0001 ,
		_w6384_
	);
	LUT2 #(
		.INIT('h8)
	) name4239 (
		\u1_slt0_reg[15]/P0001 ,
		_w6384_,
		_w6385_
	);
	LUT2 #(
		.INIT('h1)
	) name4240 (
		_w6382_,
		_w6383_,
		_w6386_
	);
	LUT2 #(
		.INIT('h8)
	) name4241 (
		_w6385_,
		_w6386_,
		_w6387_
	);
	LUT2 #(
		.INIT('h1)
	) name4242 (
		_w3309_,
		_w6387_,
		_w6388_
	);
	LUT2 #(
		.INIT('h1)
	) name4243 (
		\in_valid_s_reg[1]/NET0131 ,
		\u14_u7_en_out_l_reg/NET0131 ,
		_w6389_
	);
	LUT2 #(
		.INIT('h2)
	) name4244 (
		\u13_icc_r_reg[9]/NET0131 ,
		\u1_slt0_reg[11]/P0001 ,
		_w6390_
	);
	LUT2 #(
		.INIT('h2)
	) name4245 (
		\u13_icc_r_reg[8]/NET0131 ,
		\u14_u7_full_empty_r_reg/P0001 ,
		_w6391_
	);
	LUT2 #(
		.INIT('h8)
	) name4246 (
		\u1_slt0_reg[15]/P0001 ,
		_w6391_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name4247 (
		_w6389_,
		_w6390_,
		_w6393_
	);
	LUT2 #(
		.INIT('h8)
	) name4248 (
		_w6392_,
		_w6393_,
		_w6394_
	);
	LUT2 #(
		.INIT('h1)
	) name4249 (
		_w3499_,
		_w6394_,
		_w6395_
	);
	LUT2 #(
		.INIT('h1)
	) name4250 (
		\in_valid_s_reg[2]/NET0131 ,
		\u14_u8_en_out_l_reg/NET0131 ,
		_w6396_
	);
	LUT2 #(
		.INIT('h2)
	) name4251 (
		\u13_icc_r_reg[17]/NET0131 ,
		\u1_slt0_reg[9]/P0001 ,
		_w6397_
	);
	LUT2 #(
		.INIT('h2)
	) name4252 (
		\u13_icc_r_reg[16]/NET0131 ,
		\u14_u8_full_empty_r_reg/P0001 ,
		_w6398_
	);
	LUT2 #(
		.INIT('h8)
	) name4253 (
		\u1_slt0_reg[15]/P0001 ,
		_w6398_,
		_w6399_
	);
	LUT2 #(
		.INIT('h1)
	) name4254 (
		_w6396_,
		_w6397_,
		_w6400_
	);
	LUT2 #(
		.INIT('h8)
	) name4255 (
		_w6399_,
		_w6400_,
		_w6401_
	);
	LUT2 #(
		.INIT('h1)
	) name4256 (
		_w3062_,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h2)
	) name4257 (
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		_w6403_
	);
	LUT2 #(
		.INIT('h4)
	) name4258 (
		\u12_o9_we_reg/P0001 ,
		\u8_wp_reg[0]/P0001 ,
		_w6404_
	);
	LUT2 #(
		.INIT('h1)
	) name4259 (
		_w6403_,
		_w6404_,
		_w6405_
	);
	LUT2 #(
		.INIT('h2)
	) name4260 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w6405_,
		_w6406_
	);
	LUT2 #(
		.INIT('h2)
	) name4261 (
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		_w6407_
	);
	LUT2 #(
		.INIT('h4)
	) name4262 (
		\u12_o3_we_reg/P0001 ,
		\u3_wp_reg[0]/P0001 ,
		_w6408_
	);
	LUT2 #(
		.INIT('h1)
	) name4263 (
		_w6407_,
		_w6408_,
		_w6409_
	);
	LUT2 #(
		.INIT('h2)
	) name4264 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w6409_,
		_w6410_
	);
	LUT2 #(
		.INIT('h2)
	) name4265 (
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		_w6411_
	);
	LUT2 #(
		.INIT('h4)
	) name4266 (
		\u12_o4_we_reg/P0001 ,
		\u4_wp_reg[0]/P0001 ,
		_w6412_
	);
	LUT2 #(
		.INIT('h1)
	) name4267 (
		_w6411_,
		_w6412_,
		_w6413_
	);
	LUT2 #(
		.INIT('h2)
	) name4268 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w6413_,
		_w6414_
	);
	LUT2 #(
		.INIT('h2)
	) name4269 (
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		_w6415_
	);
	LUT2 #(
		.INIT('h4)
	) name4270 (
		\u12_o6_we_reg/P0001 ,
		\u5_wp_reg[0]/P0001 ,
		_w6416_
	);
	LUT2 #(
		.INIT('h1)
	) name4271 (
		_w6415_,
		_w6416_,
		_w6417_
	);
	LUT2 #(
		.INIT('h2)
	) name4272 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w6417_,
		_w6418_
	);
	LUT2 #(
		.INIT('h2)
	) name4273 (
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		_w6419_
	);
	LUT2 #(
		.INIT('h4)
	) name4274 (
		\u12_o7_we_reg/P0001 ,
		\u6_wp_reg[0]/P0001 ,
		_w6420_
	);
	LUT2 #(
		.INIT('h1)
	) name4275 (
		_w6419_,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('h2)
	) name4276 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w6421_,
		_w6422_
	);
	LUT2 #(
		.INIT('h2)
	) name4277 (
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		_w6423_
	);
	LUT2 #(
		.INIT('h4)
	) name4278 (
		\u12_o8_we_reg/P0001 ,
		\u7_wp_reg[0]/P0001 ,
		_w6424_
	);
	LUT2 #(
		.INIT('h1)
	) name4279 (
		_w6423_,
		_w6424_,
		_w6425_
	);
	LUT2 #(
		.INIT('h2)
	) name4280 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w6425_,
		_w6426_
	);
	LUT2 #(
		.INIT('h1)
	) name4281 (
		\u8_wp_reg[1]/NET0131 ,
		_w6300_,
		_w6427_
	);
	LUT2 #(
		.INIT('h2)
	) name4282 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w6301_,
		_w6428_
	);
	LUT2 #(
		.INIT('h4)
	) name4283 (
		_w6427_,
		_w6428_,
		_w6429_
	);
	LUT2 #(
		.INIT('h1)
	) name4284 (
		\u4_wp_reg[1]/NET0131 ,
		_w6306_,
		_w6430_
	);
	LUT2 #(
		.INIT('h2)
	) name4285 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w6307_,
		_w6431_
	);
	LUT2 #(
		.INIT('h4)
	) name4286 (
		_w6430_,
		_w6431_,
		_w6432_
	);
	LUT2 #(
		.INIT('h1)
	) name4287 (
		\u5_wp_reg[1]/NET0131 ,
		_w6312_,
		_w6433_
	);
	LUT2 #(
		.INIT('h2)
	) name4288 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w6313_,
		_w6434_
	);
	LUT2 #(
		.INIT('h4)
	) name4289 (
		_w6433_,
		_w6434_,
		_w6435_
	);
	LUT2 #(
		.INIT('h1)
	) name4290 (
		\u3_wp_reg[1]/NET0131 ,
		_w6318_,
		_w6436_
	);
	LUT2 #(
		.INIT('h2)
	) name4291 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w6319_,
		_w6437_
	);
	LUT2 #(
		.INIT('h4)
	) name4292 (
		_w6436_,
		_w6437_,
		_w6438_
	);
	LUT2 #(
		.INIT('h1)
	) name4293 (
		\u6_wp_reg[1]/NET0131 ,
		_w6324_,
		_w6439_
	);
	LUT2 #(
		.INIT('h2)
	) name4294 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w6325_,
		_w6440_
	);
	LUT2 #(
		.INIT('h4)
	) name4295 (
		_w6439_,
		_w6440_,
		_w6441_
	);
	LUT2 #(
		.INIT('h1)
	) name4296 (
		\u7_wp_reg[1]/NET0131 ,
		_w6330_,
		_w6442_
	);
	LUT2 #(
		.INIT('h2)
	) name4297 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w6331_,
		_w6443_
	);
	LUT2 #(
		.INIT('h4)
	) name4298 (
		_w6442_,
		_w6443_,
		_w6444_
	);
	LUT2 #(
		.INIT('h1)
	) name4299 (
		\u15_rdd1_reg/NET0131 ,
		_w6135_,
		_w6445_
	);
	LUT2 #(
		.INIT('h2)
	) name4300 (
		\u15_crac_rd_reg/NET0131 ,
		_w6445_,
		_w6446_
	);
	LUT2 #(
		.INIT('h8)
	) name4301 (
		\u15_crac_rd_reg/NET0131 ,
		_w6135_,
		_w6447_
	);
	LUT2 #(
		.INIT('h8)
	) name4302 (
		\u15_crac_rd_done_reg/P0001 ,
		\u15_rdd3_reg/NET0131 ,
		_w6448_
	);
	LUT2 #(
		.INIT('h2)
	) name4303 (
		\u15_rdd2_reg/NET0131 ,
		_w6448_,
		_w6449_
	);
	LUT2 #(
		.INIT('h1)
	) name4304 (
		_w6447_,
		_w6449_,
		_w6450_
	);
	LUT2 #(
		.INIT('h8)
	) name4305 (
		\u15_rdd2_reg/NET0131 ,
		_w6215_,
		_w6451_
	);
	LUT2 #(
		.INIT('h4)
	) name4306 (
		\u15_crac_rd_done_reg/P0001 ,
		\u15_rdd3_reg/NET0131 ,
		_w6452_
	);
	LUT2 #(
		.INIT('h1)
	) name4307 (
		_w6451_,
		_w6452_,
		_w6453_
	);
	LUT2 #(
		.INIT('h8)
	) name4308 (
		\u2_res_cnt_reg[0]/P0001 ,
		_w5629_,
		_w6454_
	);
	LUT2 #(
		.INIT('h8)
	) name4309 (
		\u2_res_cnt_reg[1]/P0001 ,
		_w6454_,
		_w6455_
	);
	LUT2 #(
		.INIT('h8)
	) name4310 (
		\u2_res_cnt_reg[2]/P0001 ,
		_w6455_,
		_w6456_
	);
	LUT2 #(
		.INIT('h1)
	) name4311 (
		\u2_res_cnt_reg[3]/P0001 ,
		_w6456_,
		_w6457_
	);
	LUT2 #(
		.INIT('h8)
	) name4312 (
		\u2_res_cnt_reg[3]/P0001 ,
		_w6456_,
		_w6458_
	);
	LUT2 #(
		.INIT('h2)
	) name4313 (
		\u2_sync_resume_reg/NET0131 ,
		_w6457_,
		_w6459_
	);
	LUT2 #(
		.INIT('h4)
	) name4314 (
		_w6458_,
		_w6459_,
		_w6460_
	);
	LUT2 #(
		.INIT('h8)
	) name4315 (
		\u12_rf_we_reg/P0001 ,
		_w6143_,
		_w6461_
	);
	LUT2 #(
		.INIT('h8)
	) name4316 (
		\u12_dout_reg[0]/P0001 ,
		_w6461_,
		_w6462_
	);
	LUT2 #(
		.INIT('h8)
	) name4317 (
		\u12_dout_reg[1]/P0001 ,
		_w6461_,
		_w6463_
	);
	LUT2 #(
		.INIT('h1)
	) name4318 (
		\u14_crac_valid_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w6464_
	);
	LUT2 #(
		.INIT('h4)
	) name4319 (
		\u15_crac_wr_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w6465_
	);
	LUT2 #(
		.INIT('h4)
	) name4320 (
		\u15_crac_rd_reg/NET0131 ,
		_w6465_,
		_w6466_
	);
	LUT2 #(
		.INIT('h1)
	) name4321 (
		_w6464_,
		_w6466_,
		_w6467_
	);
	LUT2 #(
		.INIT('h8)
	) name4322 (
		\u15_rdd3_reg/NET0131 ,
		_w6215_,
		_w6468_
	);
	LUT2 #(
		.INIT('h8)
	) name4323 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[1]/NET0131 ,
		_w6469_
	);
	LUT2 #(
		.INIT('h8)
	) name4324 (
		\u2_cnt_reg[2]/NET0131 ,
		_w6469_,
		_w6470_
	);
	LUT2 #(
		.INIT('h8)
	) name4325 (
		\u2_cnt_reg[3]/NET0131 ,
		_w6470_,
		_w6471_
	);
	LUT2 #(
		.INIT('h8)
	) name4326 (
		\u2_cnt_reg[4]/NET0131 ,
		_w6471_,
		_w6472_
	);
	LUT2 #(
		.INIT('h8)
	) name4327 (
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		_w6473_
	);
	LUT2 #(
		.INIT('h8)
	) name4328 (
		_w6472_,
		_w6473_,
		_w6474_
	);
	LUT2 #(
		.INIT('h2)
	) name4329 (
		\u2_cnt_reg[7]/NET0131 ,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h4)
	) name4330 (
		\u2_cnt_reg[7]/NET0131 ,
		_w6474_,
		_w6476_
	);
	LUT2 #(
		.INIT('h1)
	) name4331 (
		suspended_o_pad,
		_w6475_,
		_w6477_
	);
	LUT2 #(
		.INIT('h4)
	) name4332 (
		_w6476_,
		_w6477_,
		_w6478_
	);
	LUT2 #(
		.INIT('h8)
	) name4333 (
		\u2_to_cnt_reg[0]/NET0131 ,
		\u2_to_cnt_reg[1]/NET0131 ,
		_w6479_
	);
	LUT2 #(
		.INIT('h8)
	) name4334 (
		\u2_to_cnt_reg[2]/NET0131 ,
		_w6479_,
		_w6480_
	);
	LUT2 #(
		.INIT('h8)
	) name4335 (
		\u2_to_cnt_reg[3]/NET0131 ,
		_w6480_,
		_w6481_
	);
	LUT2 #(
		.INIT('h1)
	) name4336 (
		\u2_to_cnt_reg[3]/NET0131 ,
		_w6480_,
		_w6482_
	);
	LUT2 #(
		.INIT('h1)
	) name4337 (
		\u2_bit_clk_e_reg/P0001 ,
		_w6481_,
		_w6483_
	);
	LUT2 #(
		.INIT('h4)
	) name4338 (
		_w6482_,
		_w6483_,
		_w6484_
	);
	LUT2 #(
		.INIT('h8)
	) name4339 (
		\u8_wp_reg[1]/NET0131 ,
		_w6403_,
		_w6485_
	);
	LUT2 #(
		.INIT('h2)
	) name4340 (
		\u8_mem_reg[2][5]/NET0131 ,
		_w6485_,
		_w6486_
	);
	LUT2 #(
		.INIT('h8)
	) name4341 (
		\u12_dout_reg[5]/P0001 ,
		_w6485_,
		_w6487_
	);
	LUT2 #(
		.INIT('h1)
	) name4342 (
		_w6486_,
		_w6487_,
		_w6488_
	);
	LUT2 #(
		.INIT('h4)
	) name4343 (
		\u3_wp_reg[1]/NET0131 ,
		_w6318_,
		_w6489_
	);
	LUT2 #(
		.INIT('h2)
	) name4344 (
		\u3_mem_reg[1][29]/NET0131 ,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('h8)
	) name4345 (
		\u12_dout_reg[29]/P0001 ,
		_w6489_,
		_w6491_
	);
	LUT2 #(
		.INIT('h1)
	) name4346 (
		_w6490_,
		_w6491_,
		_w6492_
	);
	LUT2 #(
		.INIT('h2)
	) name4347 (
		\u8_mem_reg[2][6]/NET0131 ,
		_w6485_,
		_w6493_
	);
	LUT2 #(
		.INIT('h8)
	) name4348 (
		\u12_dout_reg[6]/P0001 ,
		_w6485_,
		_w6494_
	);
	LUT2 #(
		.INIT('h1)
	) name4349 (
		_w6493_,
		_w6494_,
		_w6495_
	);
	LUT2 #(
		.INIT('h2)
	) name4350 (
		\u8_mem_reg[2][7]/NET0131 ,
		_w6485_,
		_w6496_
	);
	LUT2 #(
		.INIT('h8)
	) name4351 (
		\u12_dout_reg[7]/P0001 ,
		_w6485_,
		_w6497_
	);
	LUT2 #(
		.INIT('h1)
	) name4352 (
		_w6496_,
		_w6497_,
		_w6498_
	);
	LUT2 #(
		.INIT('h2)
	) name4353 (
		\u3_mem_reg[1][2]/NET0131 ,
		_w6489_,
		_w6499_
	);
	LUT2 #(
		.INIT('h8)
	) name4354 (
		\u12_dout_reg[2]/P0001 ,
		_w6489_,
		_w6500_
	);
	LUT2 #(
		.INIT('h1)
	) name4355 (
		_w6499_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h2)
	) name4356 (
		\u8_mem_reg[2][8]/NET0131 ,
		_w6485_,
		_w6502_
	);
	LUT2 #(
		.INIT('h8)
	) name4357 (
		\u12_dout_reg[8]/P0001 ,
		_w6485_,
		_w6503_
	);
	LUT2 #(
		.INIT('h1)
	) name4358 (
		_w6502_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h2)
	) name4359 (
		\u8_mem_reg[2][9]/NET0131 ,
		_w6485_,
		_w6505_
	);
	LUT2 #(
		.INIT('h8)
	) name4360 (
		\u12_dout_reg[9]/P0001 ,
		_w6485_,
		_w6506_
	);
	LUT2 #(
		.INIT('h1)
	) name4361 (
		_w6505_,
		_w6506_,
		_w6507_
	);
	LUT2 #(
		.INIT('h2)
	) name4362 (
		\u8_mem_reg[3][19]/NET0131 ,
		_w6301_,
		_w6508_
	);
	LUT2 #(
		.INIT('h8)
	) name4363 (
		\u12_dout_reg[19]/P0001 ,
		_w6301_,
		_w6509_
	);
	LUT2 #(
		.INIT('h1)
	) name4364 (
		_w6508_,
		_w6509_,
		_w6510_
	);
	LUT2 #(
		.INIT('h2)
	) name4365 (
		\u8_mem_reg[3][0]/NET0131 ,
		_w6301_,
		_w6511_
	);
	LUT2 #(
		.INIT('h8)
	) name4366 (
		\u12_dout_reg[0]/P0001 ,
		_w6301_,
		_w6512_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		_w6511_,
		_w6512_,
		_w6513_
	);
	LUT2 #(
		.INIT('h2)
	) name4368 (
		\u8_mem_reg[3][10]/NET0131 ,
		_w6301_,
		_w6514_
	);
	LUT2 #(
		.INIT('h8)
	) name4369 (
		\u12_dout_reg[10]/P0001 ,
		_w6301_,
		_w6515_
	);
	LUT2 #(
		.INIT('h1)
	) name4370 (
		_w6514_,
		_w6515_,
		_w6516_
	);
	LUT2 #(
		.INIT('h2)
	) name4371 (
		\u3_mem_reg[1][31]/NET0131 ,
		_w6489_,
		_w6517_
	);
	LUT2 #(
		.INIT('h8)
	) name4372 (
		\u12_dout_reg[31]/P0001 ,
		_w6489_,
		_w6518_
	);
	LUT2 #(
		.INIT('h1)
	) name4373 (
		_w6517_,
		_w6518_,
		_w6519_
	);
	LUT2 #(
		.INIT('h2)
	) name4374 (
		\u8_mem_reg[3][12]/NET0131 ,
		_w6301_,
		_w6520_
	);
	LUT2 #(
		.INIT('h8)
	) name4375 (
		\u12_dout_reg[12]/P0001 ,
		_w6301_,
		_w6521_
	);
	LUT2 #(
		.INIT('h1)
	) name4376 (
		_w6520_,
		_w6521_,
		_w6522_
	);
	LUT2 #(
		.INIT('h2)
	) name4377 (
		\u3_mem_reg[1][3]/NET0131 ,
		_w6489_,
		_w6523_
	);
	LUT2 #(
		.INIT('h8)
	) name4378 (
		\u12_dout_reg[3]/P0001 ,
		_w6489_,
		_w6524_
	);
	LUT2 #(
		.INIT('h1)
	) name4379 (
		_w6523_,
		_w6524_,
		_w6525_
	);
	LUT2 #(
		.INIT('h2)
	) name4380 (
		\u8_mem_reg[3][13]/NET0131 ,
		_w6301_,
		_w6526_
	);
	LUT2 #(
		.INIT('h8)
	) name4381 (
		\u12_dout_reg[13]/P0001 ,
		_w6301_,
		_w6527_
	);
	LUT2 #(
		.INIT('h1)
	) name4382 (
		_w6526_,
		_w6527_,
		_w6528_
	);
	LUT2 #(
		.INIT('h2)
	) name4383 (
		\u8_mem_reg[3][14]/NET0131 ,
		_w6301_,
		_w6529_
	);
	LUT2 #(
		.INIT('h8)
	) name4384 (
		\u12_dout_reg[14]/P0001 ,
		_w6301_,
		_w6530_
	);
	LUT2 #(
		.INIT('h1)
	) name4385 (
		_w6529_,
		_w6530_,
		_w6531_
	);
	LUT2 #(
		.INIT('h2)
	) name4386 (
		\u8_mem_reg[3][15]/NET0131 ,
		_w6301_,
		_w6532_
	);
	LUT2 #(
		.INIT('h8)
	) name4387 (
		\u12_dout_reg[15]/P0001 ,
		_w6301_,
		_w6533_
	);
	LUT2 #(
		.INIT('h1)
	) name4388 (
		_w6532_,
		_w6533_,
		_w6534_
	);
	LUT2 #(
		.INIT('h2)
	) name4389 (
		\u3_mem_reg[1][4]/NET0131 ,
		_w6489_,
		_w6535_
	);
	LUT2 #(
		.INIT('h8)
	) name4390 (
		\u12_dout_reg[4]/P0001 ,
		_w6489_,
		_w6536_
	);
	LUT2 #(
		.INIT('h1)
	) name4391 (
		_w6535_,
		_w6536_,
		_w6537_
	);
	LUT2 #(
		.INIT('h2)
	) name4392 (
		\u8_mem_reg[3][16]/NET0131 ,
		_w6301_,
		_w6538_
	);
	LUT2 #(
		.INIT('h8)
	) name4393 (
		\u12_dout_reg[16]/P0001 ,
		_w6301_,
		_w6539_
	);
	LUT2 #(
		.INIT('h1)
	) name4394 (
		_w6538_,
		_w6539_,
		_w6540_
	);
	LUT2 #(
		.INIT('h2)
	) name4395 (
		\u3_mem_reg[1][5]/NET0131 ,
		_w6489_,
		_w6541_
	);
	LUT2 #(
		.INIT('h8)
	) name4396 (
		\u12_dout_reg[5]/P0001 ,
		_w6489_,
		_w6542_
	);
	LUT2 #(
		.INIT('h1)
	) name4397 (
		_w6541_,
		_w6542_,
		_w6543_
	);
	LUT2 #(
		.INIT('h2)
	) name4398 (
		\u8_mem_reg[3][17]/NET0131 ,
		_w6301_,
		_w6544_
	);
	LUT2 #(
		.INIT('h8)
	) name4399 (
		\u12_dout_reg[17]/P0001 ,
		_w6301_,
		_w6545_
	);
	LUT2 #(
		.INIT('h1)
	) name4400 (
		_w6544_,
		_w6545_,
		_w6546_
	);
	LUT2 #(
		.INIT('h2)
	) name4401 (
		\u8_mem_reg[3][18]/NET0131 ,
		_w6301_,
		_w6547_
	);
	LUT2 #(
		.INIT('h8)
	) name4402 (
		\u12_dout_reg[18]/P0001 ,
		_w6301_,
		_w6548_
	);
	LUT2 #(
		.INIT('h1)
	) name4403 (
		_w6547_,
		_w6548_,
		_w6549_
	);
	LUT2 #(
		.INIT('h2)
	) name4404 (
		\u3_mem_reg[1][6]/NET0131 ,
		_w6489_,
		_w6550_
	);
	LUT2 #(
		.INIT('h8)
	) name4405 (
		\u12_dout_reg[6]/P0001 ,
		_w6489_,
		_w6551_
	);
	LUT2 #(
		.INIT('h1)
	) name4406 (
		_w6550_,
		_w6551_,
		_w6552_
	);
	LUT2 #(
		.INIT('h2)
	) name4407 (
		\u8_mem_reg[3][1]/NET0131 ,
		_w6301_,
		_w6553_
	);
	LUT2 #(
		.INIT('h8)
	) name4408 (
		\u12_dout_reg[1]/P0001 ,
		_w6301_,
		_w6554_
	);
	LUT2 #(
		.INIT('h1)
	) name4409 (
		_w6553_,
		_w6554_,
		_w6555_
	);
	LUT2 #(
		.INIT('h2)
	) name4410 (
		\u3_mem_reg[1][7]/NET0131 ,
		_w6489_,
		_w6556_
	);
	LUT2 #(
		.INIT('h8)
	) name4411 (
		\u12_dout_reg[7]/P0001 ,
		_w6489_,
		_w6557_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w6556_,
		_w6557_,
		_w6558_
	);
	LUT2 #(
		.INIT('h2)
	) name4413 (
		\u8_mem_reg[3][20]/NET0131 ,
		_w6301_,
		_w6559_
	);
	LUT2 #(
		.INIT('h8)
	) name4414 (
		\u12_dout_reg[20]/P0001 ,
		_w6301_,
		_w6560_
	);
	LUT2 #(
		.INIT('h1)
	) name4415 (
		_w6559_,
		_w6560_,
		_w6561_
	);
	LUT2 #(
		.INIT('h2)
	) name4416 (
		\u8_mem_reg[3][21]/NET0131 ,
		_w6301_,
		_w6562_
	);
	LUT2 #(
		.INIT('h8)
	) name4417 (
		\u12_dout_reg[21]/P0001 ,
		_w6301_,
		_w6563_
	);
	LUT2 #(
		.INIT('h1)
	) name4418 (
		_w6562_,
		_w6563_,
		_w6564_
	);
	LUT2 #(
		.INIT('h2)
	) name4419 (
		\u3_mem_reg[1][8]/NET0131 ,
		_w6489_,
		_w6565_
	);
	LUT2 #(
		.INIT('h8)
	) name4420 (
		\u12_dout_reg[8]/P0001 ,
		_w6489_,
		_w6566_
	);
	LUT2 #(
		.INIT('h1)
	) name4421 (
		_w6565_,
		_w6566_,
		_w6567_
	);
	LUT2 #(
		.INIT('h2)
	) name4422 (
		\u8_mem_reg[3][22]/NET0131 ,
		_w6301_,
		_w6568_
	);
	LUT2 #(
		.INIT('h8)
	) name4423 (
		\u12_dout_reg[22]/P0001 ,
		_w6301_,
		_w6569_
	);
	LUT2 #(
		.INIT('h1)
	) name4424 (
		_w6568_,
		_w6569_,
		_w6570_
	);
	LUT2 #(
		.INIT('h2)
	) name4425 (
		\u8_mem_reg[3][23]/NET0131 ,
		_w6301_,
		_w6571_
	);
	LUT2 #(
		.INIT('h8)
	) name4426 (
		\u12_dout_reg[23]/P0001 ,
		_w6301_,
		_w6572_
	);
	LUT2 #(
		.INIT('h1)
	) name4427 (
		_w6571_,
		_w6572_,
		_w6573_
	);
	LUT2 #(
		.INIT('h2)
	) name4428 (
		\u3_mem_reg[1][9]/NET0131 ,
		_w6489_,
		_w6574_
	);
	LUT2 #(
		.INIT('h8)
	) name4429 (
		\u12_dout_reg[9]/P0001 ,
		_w6489_,
		_w6575_
	);
	LUT2 #(
		.INIT('h1)
	) name4430 (
		_w6574_,
		_w6575_,
		_w6576_
	);
	LUT2 #(
		.INIT('h2)
	) name4431 (
		\u8_mem_reg[3][24]/NET0131 ,
		_w6301_,
		_w6577_
	);
	LUT2 #(
		.INIT('h8)
	) name4432 (
		\u12_dout_reg[24]/P0001 ,
		_w6301_,
		_w6578_
	);
	LUT2 #(
		.INIT('h1)
	) name4433 (
		_w6577_,
		_w6578_,
		_w6579_
	);
	LUT2 #(
		.INIT('h2)
	) name4434 (
		\u8_mem_reg[3][25]/NET0131 ,
		_w6301_,
		_w6580_
	);
	LUT2 #(
		.INIT('h8)
	) name4435 (
		\u12_dout_reg[25]/P0001 ,
		_w6301_,
		_w6581_
	);
	LUT2 #(
		.INIT('h1)
	) name4436 (
		_w6580_,
		_w6581_,
		_w6582_
	);
	LUT2 #(
		.INIT('h8)
	) name4437 (
		\u3_wp_reg[1]/NET0131 ,
		_w6407_,
		_w6583_
	);
	LUT2 #(
		.INIT('h2)
	) name4438 (
		\u3_mem_reg[2][0]/NET0131 ,
		_w6583_,
		_w6584_
	);
	LUT2 #(
		.INIT('h8)
	) name4439 (
		\u12_dout_reg[0]/P0001 ,
		_w6583_,
		_w6585_
	);
	LUT2 #(
		.INIT('h1)
	) name4440 (
		_w6584_,
		_w6585_,
		_w6586_
	);
	LUT2 #(
		.INIT('h2)
	) name4441 (
		\u8_mem_reg[3][27]/NET0131 ,
		_w6301_,
		_w6587_
	);
	LUT2 #(
		.INIT('h8)
	) name4442 (
		\u12_dout_reg[27]/P0001 ,
		_w6301_,
		_w6588_
	);
	LUT2 #(
		.INIT('h1)
	) name4443 (
		_w6587_,
		_w6588_,
		_w6589_
	);
	LUT2 #(
		.INIT('h2)
	) name4444 (
		\u3_mem_reg[2][10]/NET0131 ,
		_w6583_,
		_w6590_
	);
	LUT2 #(
		.INIT('h8)
	) name4445 (
		\u12_dout_reg[10]/P0001 ,
		_w6583_,
		_w6591_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		_w6590_,
		_w6591_,
		_w6592_
	);
	LUT2 #(
		.INIT('h2)
	) name4447 (
		\u8_mem_reg[3][29]/NET0131 ,
		_w6301_,
		_w6593_
	);
	LUT2 #(
		.INIT('h8)
	) name4448 (
		\u12_dout_reg[29]/P0001 ,
		_w6301_,
		_w6594_
	);
	LUT2 #(
		.INIT('h1)
	) name4449 (
		_w6593_,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h2)
	) name4450 (
		\u3_mem_reg[2][11]/NET0131 ,
		_w6583_,
		_w6596_
	);
	LUT2 #(
		.INIT('h8)
	) name4451 (
		\u12_dout_reg[11]/P0001 ,
		_w6583_,
		_w6597_
	);
	LUT2 #(
		.INIT('h1)
	) name4452 (
		_w6596_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h2)
	) name4453 (
		\u8_mem_reg[3][2]/NET0131 ,
		_w6301_,
		_w6599_
	);
	LUT2 #(
		.INIT('h8)
	) name4454 (
		\u12_dout_reg[2]/P0001 ,
		_w6301_,
		_w6600_
	);
	LUT2 #(
		.INIT('h1)
	) name4455 (
		_w6599_,
		_w6600_,
		_w6601_
	);
	LUT2 #(
		.INIT('h2)
	) name4456 (
		\u8_mem_reg[3][30]/NET0131 ,
		_w6301_,
		_w6602_
	);
	LUT2 #(
		.INIT('h8)
	) name4457 (
		\u12_dout_reg[30]/P0001 ,
		_w6301_,
		_w6603_
	);
	LUT2 #(
		.INIT('h1)
	) name4458 (
		_w6602_,
		_w6603_,
		_w6604_
	);
	LUT2 #(
		.INIT('h2)
	) name4459 (
		\u3_mem_reg[2][12]/NET0131 ,
		_w6583_,
		_w6605_
	);
	LUT2 #(
		.INIT('h8)
	) name4460 (
		\u12_dout_reg[12]/P0001 ,
		_w6583_,
		_w6606_
	);
	LUT2 #(
		.INIT('h1)
	) name4461 (
		_w6605_,
		_w6606_,
		_w6607_
	);
	LUT2 #(
		.INIT('h2)
	) name4462 (
		\u8_mem_reg[3][3]/NET0131 ,
		_w6301_,
		_w6608_
	);
	LUT2 #(
		.INIT('h8)
	) name4463 (
		\u12_dout_reg[3]/P0001 ,
		_w6301_,
		_w6609_
	);
	LUT2 #(
		.INIT('h1)
	) name4464 (
		_w6608_,
		_w6609_,
		_w6610_
	);
	LUT2 #(
		.INIT('h2)
	) name4465 (
		\u3_mem_reg[2][13]/NET0131 ,
		_w6583_,
		_w6611_
	);
	LUT2 #(
		.INIT('h8)
	) name4466 (
		\u12_dout_reg[13]/P0001 ,
		_w6583_,
		_w6612_
	);
	LUT2 #(
		.INIT('h1)
	) name4467 (
		_w6611_,
		_w6612_,
		_w6613_
	);
	LUT2 #(
		.INIT('h2)
	) name4468 (
		\u8_mem_reg[3][5]/NET0131 ,
		_w6301_,
		_w6614_
	);
	LUT2 #(
		.INIT('h8)
	) name4469 (
		\u12_dout_reg[5]/P0001 ,
		_w6301_,
		_w6615_
	);
	LUT2 #(
		.INIT('h1)
	) name4470 (
		_w6614_,
		_w6615_,
		_w6616_
	);
	LUT2 #(
		.INIT('h2)
	) name4471 (
		\u8_mem_reg[3][7]/NET0131 ,
		_w6301_,
		_w6617_
	);
	LUT2 #(
		.INIT('h8)
	) name4472 (
		\u12_dout_reg[7]/P0001 ,
		_w6301_,
		_w6618_
	);
	LUT2 #(
		.INIT('h1)
	) name4473 (
		_w6617_,
		_w6618_,
		_w6619_
	);
	LUT2 #(
		.INIT('h2)
	) name4474 (
		\u3_mem_reg[2][15]/NET0131 ,
		_w6583_,
		_w6620_
	);
	LUT2 #(
		.INIT('h8)
	) name4475 (
		\u12_dout_reg[15]/P0001 ,
		_w6583_,
		_w6621_
	);
	LUT2 #(
		.INIT('h1)
	) name4476 (
		_w6620_,
		_w6621_,
		_w6622_
	);
	LUT2 #(
		.INIT('h2)
	) name4477 (
		\u8_mem_reg[3][9]/NET0131 ,
		_w6301_,
		_w6623_
	);
	LUT2 #(
		.INIT('h8)
	) name4478 (
		\u12_dout_reg[9]/P0001 ,
		_w6301_,
		_w6624_
	);
	LUT2 #(
		.INIT('h1)
	) name4479 (
		_w6623_,
		_w6624_,
		_w6625_
	);
	LUT2 #(
		.INIT('h2)
	) name4480 (
		\u3_mem_reg[2][16]/NET0131 ,
		_w6583_,
		_w6626_
	);
	LUT2 #(
		.INIT('h8)
	) name4481 (
		\u12_dout_reg[16]/P0001 ,
		_w6583_,
		_w6627_
	);
	LUT2 #(
		.INIT('h1)
	) name4482 (
		_w6626_,
		_w6627_,
		_w6628_
	);
	LUT2 #(
		.INIT('h4)
	) name4483 (
		\u8_wp_reg[1]/NET0131 ,
		_w6300_,
		_w6629_
	);
	LUT2 #(
		.INIT('h2)
	) name4484 (
		\u8_mem_reg[1][4]/NET0131 ,
		_w6629_,
		_w6630_
	);
	LUT2 #(
		.INIT('h8)
	) name4485 (
		\u12_dout_reg[4]/P0001 ,
		_w6629_,
		_w6631_
	);
	LUT2 #(
		.INIT('h1)
	) name4486 (
		_w6630_,
		_w6631_,
		_w6632_
	);
	LUT2 #(
		.INIT('h2)
	) name4487 (
		\u3_mem_reg[2][18]/NET0131 ,
		_w6583_,
		_w6633_
	);
	LUT2 #(
		.INIT('h8)
	) name4488 (
		\u12_dout_reg[18]/P0001 ,
		_w6583_,
		_w6634_
	);
	LUT2 #(
		.INIT('h1)
	) name4489 (
		_w6633_,
		_w6634_,
		_w6635_
	);
	LUT2 #(
		.INIT('h2)
	) name4490 (
		\u3_mem_reg[2][19]/NET0131 ,
		_w6583_,
		_w6636_
	);
	LUT2 #(
		.INIT('h8)
	) name4491 (
		\u12_dout_reg[19]/P0001 ,
		_w6583_,
		_w6637_
	);
	LUT2 #(
		.INIT('h1)
	) name4492 (
		_w6636_,
		_w6637_,
		_w6638_
	);
	LUT2 #(
		.INIT('h2)
	) name4493 (
		\u3_mem_reg[2][1]/NET0131 ,
		_w6583_,
		_w6639_
	);
	LUT2 #(
		.INIT('h8)
	) name4494 (
		\u12_dout_reg[1]/P0001 ,
		_w6583_,
		_w6640_
	);
	LUT2 #(
		.INIT('h1)
	) name4495 (
		_w6639_,
		_w6640_,
		_w6641_
	);
	LUT2 #(
		.INIT('h2)
	) name4496 (
		\u3_mem_reg[1][30]/NET0131 ,
		_w6489_,
		_w6642_
	);
	LUT2 #(
		.INIT('h8)
	) name4497 (
		\u12_dout_reg[30]/P0001 ,
		_w6489_,
		_w6643_
	);
	LUT2 #(
		.INIT('h1)
	) name4498 (
		_w6642_,
		_w6643_,
		_w6644_
	);
	LUT2 #(
		.INIT('h2)
	) name4499 (
		\u3_mem_reg[2][21]/NET0131 ,
		_w6583_,
		_w6645_
	);
	LUT2 #(
		.INIT('h8)
	) name4500 (
		\u12_dout_reg[21]/P0001 ,
		_w6583_,
		_w6646_
	);
	LUT2 #(
		.INIT('h1)
	) name4501 (
		_w6645_,
		_w6646_,
		_w6647_
	);
	LUT2 #(
		.INIT('h2)
	) name4502 (
		\u3_mem_reg[2][22]/NET0131 ,
		_w6583_,
		_w6648_
	);
	LUT2 #(
		.INIT('h8)
	) name4503 (
		\u12_dout_reg[22]/P0001 ,
		_w6583_,
		_w6649_
	);
	LUT2 #(
		.INIT('h1)
	) name4504 (
		_w6648_,
		_w6649_,
		_w6650_
	);
	LUT2 #(
		.INIT('h2)
	) name4505 (
		\u3_mem_reg[2][24]/NET0131 ,
		_w6583_,
		_w6651_
	);
	LUT2 #(
		.INIT('h8)
	) name4506 (
		\u12_dout_reg[24]/P0001 ,
		_w6583_,
		_w6652_
	);
	LUT2 #(
		.INIT('h1)
	) name4507 (
		_w6651_,
		_w6652_,
		_w6653_
	);
	LUT2 #(
		.INIT('h2)
	) name4508 (
		\u3_mem_reg[2][26]/NET0131 ,
		_w6583_,
		_w6654_
	);
	LUT2 #(
		.INIT('h8)
	) name4509 (
		\u12_dout_reg[26]/P0001 ,
		_w6583_,
		_w6655_
	);
	LUT2 #(
		.INIT('h1)
	) name4510 (
		_w6654_,
		_w6655_,
		_w6656_
	);
	LUT2 #(
		.INIT('h2)
	) name4511 (
		\u3_mem_reg[2][27]/NET0131 ,
		_w6583_,
		_w6657_
	);
	LUT2 #(
		.INIT('h8)
	) name4512 (
		\u12_dout_reg[27]/P0001 ,
		_w6583_,
		_w6658_
	);
	LUT2 #(
		.INIT('h1)
	) name4513 (
		_w6657_,
		_w6658_,
		_w6659_
	);
	LUT2 #(
		.INIT('h2)
	) name4514 (
		\u3_mem_reg[2][28]/NET0131 ,
		_w6583_,
		_w6660_
	);
	LUT2 #(
		.INIT('h8)
	) name4515 (
		\u12_dout_reg[28]/P0001 ,
		_w6583_,
		_w6661_
	);
	LUT2 #(
		.INIT('h1)
	) name4516 (
		_w6660_,
		_w6661_,
		_w6662_
	);
	LUT2 #(
		.INIT('h2)
	) name4517 (
		\u3_mem_reg[2][29]/NET0131 ,
		_w6583_,
		_w6663_
	);
	LUT2 #(
		.INIT('h8)
	) name4518 (
		\u12_dout_reg[29]/P0001 ,
		_w6583_,
		_w6664_
	);
	LUT2 #(
		.INIT('h1)
	) name4519 (
		_w6663_,
		_w6664_,
		_w6665_
	);
	LUT2 #(
		.INIT('h2)
	) name4520 (
		\u3_mem_reg[2][2]/NET0131 ,
		_w6583_,
		_w6666_
	);
	LUT2 #(
		.INIT('h8)
	) name4521 (
		\u12_dout_reg[2]/P0001 ,
		_w6583_,
		_w6667_
	);
	LUT2 #(
		.INIT('h1)
	) name4522 (
		_w6666_,
		_w6667_,
		_w6668_
	);
	LUT2 #(
		.INIT('h2)
	) name4523 (
		\u3_mem_reg[2][30]/NET0131 ,
		_w6583_,
		_w6669_
	);
	LUT2 #(
		.INIT('h8)
	) name4524 (
		\u12_dout_reg[30]/P0001 ,
		_w6583_,
		_w6670_
	);
	LUT2 #(
		.INIT('h1)
	) name4525 (
		_w6669_,
		_w6670_,
		_w6671_
	);
	LUT2 #(
		.INIT('h2)
	) name4526 (
		\u3_mem_reg[2][31]/NET0131 ,
		_w6583_,
		_w6672_
	);
	LUT2 #(
		.INIT('h8)
	) name4527 (
		\u12_dout_reg[31]/P0001 ,
		_w6583_,
		_w6673_
	);
	LUT2 #(
		.INIT('h1)
	) name4528 (
		_w6672_,
		_w6673_,
		_w6674_
	);
	LUT2 #(
		.INIT('h2)
	) name4529 (
		\u3_mem_reg[2][3]/NET0131 ,
		_w6583_,
		_w6675_
	);
	LUT2 #(
		.INIT('h8)
	) name4530 (
		\u12_dout_reg[3]/P0001 ,
		_w6583_,
		_w6676_
	);
	LUT2 #(
		.INIT('h1)
	) name4531 (
		_w6675_,
		_w6676_,
		_w6677_
	);
	LUT2 #(
		.INIT('h2)
	) name4532 (
		\u3_mem_reg[2][4]/NET0131 ,
		_w6583_,
		_w6678_
	);
	LUT2 #(
		.INIT('h8)
	) name4533 (
		\u12_dout_reg[4]/P0001 ,
		_w6583_,
		_w6679_
	);
	LUT2 #(
		.INIT('h1)
	) name4534 (
		_w6678_,
		_w6679_,
		_w6680_
	);
	LUT2 #(
		.INIT('h2)
	) name4535 (
		\u3_mem_reg[2][5]/NET0131 ,
		_w6583_,
		_w6681_
	);
	LUT2 #(
		.INIT('h8)
	) name4536 (
		\u12_dout_reg[5]/P0001 ,
		_w6583_,
		_w6682_
	);
	LUT2 #(
		.INIT('h1)
	) name4537 (
		_w6681_,
		_w6682_,
		_w6683_
	);
	LUT2 #(
		.INIT('h2)
	) name4538 (
		\u3_mem_reg[2][6]/NET0131 ,
		_w6583_,
		_w6684_
	);
	LUT2 #(
		.INIT('h8)
	) name4539 (
		\u12_dout_reg[6]/P0001 ,
		_w6583_,
		_w6685_
	);
	LUT2 #(
		.INIT('h1)
	) name4540 (
		_w6684_,
		_w6685_,
		_w6686_
	);
	LUT2 #(
		.INIT('h2)
	) name4541 (
		\u3_mem_reg[2][7]/NET0131 ,
		_w6583_,
		_w6687_
	);
	LUT2 #(
		.INIT('h8)
	) name4542 (
		\u12_dout_reg[7]/P0001 ,
		_w6583_,
		_w6688_
	);
	LUT2 #(
		.INIT('h1)
	) name4543 (
		_w6687_,
		_w6688_,
		_w6689_
	);
	LUT2 #(
		.INIT('h2)
	) name4544 (
		\u3_mem_reg[2][8]/NET0131 ,
		_w6583_,
		_w6690_
	);
	LUT2 #(
		.INIT('h8)
	) name4545 (
		\u12_dout_reg[8]/P0001 ,
		_w6583_,
		_w6691_
	);
	LUT2 #(
		.INIT('h1)
	) name4546 (
		_w6690_,
		_w6691_,
		_w6692_
	);
	LUT2 #(
		.INIT('h2)
	) name4547 (
		\u3_mem_reg[2][9]/NET0131 ,
		_w6583_,
		_w6693_
	);
	LUT2 #(
		.INIT('h8)
	) name4548 (
		\u12_dout_reg[9]/P0001 ,
		_w6583_,
		_w6694_
	);
	LUT2 #(
		.INIT('h1)
	) name4549 (
		_w6693_,
		_w6694_,
		_w6695_
	);
	LUT2 #(
		.INIT('h2)
	) name4550 (
		\u3_mem_reg[3][0]/NET0131 ,
		_w6319_,
		_w6696_
	);
	LUT2 #(
		.INIT('h8)
	) name4551 (
		\u12_dout_reg[0]/P0001 ,
		_w6319_,
		_w6697_
	);
	LUT2 #(
		.INIT('h1)
	) name4552 (
		_w6696_,
		_w6697_,
		_w6698_
	);
	LUT2 #(
		.INIT('h2)
	) name4553 (
		\u3_mem_reg[3][10]/NET0131 ,
		_w6319_,
		_w6699_
	);
	LUT2 #(
		.INIT('h8)
	) name4554 (
		\u12_dout_reg[10]/P0001 ,
		_w6319_,
		_w6700_
	);
	LUT2 #(
		.INIT('h1)
	) name4555 (
		_w6699_,
		_w6700_,
		_w6701_
	);
	LUT2 #(
		.INIT('h2)
	) name4556 (
		\u3_mem_reg[3][11]/NET0131 ,
		_w6319_,
		_w6702_
	);
	LUT2 #(
		.INIT('h8)
	) name4557 (
		\u12_dout_reg[11]/P0001 ,
		_w6319_,
		_w6703_
	);
	LUT2 #(
		.INIT('h1)
	) name4558 (
		_w6702_,
		_w6703_,
		_w6704_
	);
	LUT2 #(
		.INIT('h2)
	) name4559 (
		\u3_mem_reg[3][12]/NET0131 ,
		_w6319_,
		_w6705_
	);
	LUT2 #(
		.INIT('h8)
	) name4560 (
		\u12_dout_reg[12]/P0001 ,
		_w6319_,
		_w6706_
	);
	LUT2 #(
		.INIT('h1)
	) name4561 (
		_w6705_,
		_w6706_,
		_w6707_
	);
	LUT2 #(
		.INIT('h2)
	) name4562 (
		\u3_mem_reg[3][13]/NET0131 ,
		_w6319_,
		_w6708_
	);
	LUT2 #(
		.INIT('h8)
	) name4563 (
		\u12_dout_reg[13]/P0001 ,
		_w6319_,
		_w6709_
	);
	LUT2 #(
		.INIT('h1)
	) name4564 (
		_w6708_,
		_w6709_,
		_w6710_
	);
	LUT2 #(
		.INIT('h2)
	) name4565 (
		\u3_mem_reg[3][14]/NET0131 ,
		_w6319_,
		_w6711_
	);
	LUT2 #(
		.INIT('h8)
	) name4566 (
		\u12_dout_reg[14]/P0001 ,
		_w6319_,
		_w6712_
	);
	LUT2 #(
		.INIT('h1)
	) name4567 (
		_w6711_,
		_w6712_,
		_w6713_
	);
	LUT2 #(
		.INIT('h2)
	) name4568 (
		\u3_mem_reg[3][15]/NET0131 ,
		_w6319_,
		_w6714_
	);
	LUT2 #(
		.INIT('h8)
	) name4569 (
		\u12_dout_reg[15]/P0001 ,
		_w6319_,
		_w6715_
	);
	LUT2 #(
		.INIT('h1)
	) name4570 (
		_w6714_,
		_w6715_,
		_w6716_
	);
	LUT2 #(
		.INIT('h2)
	) name4571 (
		\u3_mem_reg[3][16]/NET0131 ,
		_w6319_,
		_w6717_
	);
	LUT2 #(
		.INIT('h8)
	) name4572 (
		\u12_dout_reg[16]/P0001 ,
		_w6319_,
		_w6718_
	);
	LUT2 #(
		.INIT('h1)
	) name4573 (
		_w6717_,
		_w6718_,
		_w6719_
	);
	LUT2 #(
		.INIT('h2)
	) name4574 (
		\u3_mem_reg[3][17]/NET0131 ,
		_w6319_,
		_w6720_
	);
	LUT2 #(
		.INIT('h8)
	) name4575 (
		\u12_dout_reg[17]/P0001 ,
		_w6319_,
		_w6721_
	);
	LUT2 #(
		.INIT('h1)
	) name4576 (
		_w6720_,
		_w6721_,
		_w6722_
	);
	LUT2 #(
		.INIT('h2)
	) name4577 (
		\u3_mem_reg[3][18]/NET0131 ,
		_w6319_,
		_w6723_
	);
	LUT2 #(
		.INIT('h8)
	) name4578 (
		\u12_dout_reg[18]/P0001 ,
		_w6319_,
		_w6724_
	);
	LUT2 #(
		.INIT('h1)
	) name4579 (
		_w6723_,
		_w6724_,
		_w6725_
	);
	LUT2 #(
		.INIT('h2)
	) name4580 (
		\u3_mem_reg[3][19]/NET0131 ,
		_w6319_,
		_w6726_
	);
	LUT2 #(
		.INIT('h8)
	) name4581 (
		\u12_dout_reg[19]/P0001 ,
		_w6319_,
		_w6727_
	);
	LUT2 #(
		.INIT('h1)
	) name4582 (
		_w6726_,
		_w6727_,
		_w6728_
	);
	LUT2 #(
		.INIT('h2)
	) name4583 (
		\u3_mem_reg[3][1]/NET0131 ,
		_w6319_,
		_w6729_
	);
	LUT2 #(
		.INIT('h8)
	) name4584 (
		\u12_dout_reg[1]/P0001 ,
		_w6319_,
		_w6730_
	);
	LUT2 #(
		.INIT('h1)
	) name4585 (
		_w6729_,
		_w6730_,
		_w6731_
	);
	LUT2 #(
		.INIT('h2)
	) name4586 (
		\u3_mem_reg[3][21]/NET0131 ,
		_w6319_,
		_w6732_
	);
	LUT2 #(
		.INIT('h8)
	) name4587 (
		\u12_dout_reg[21]/P0001 ,
		_w6319_,
		_w6733_
	);
	LUT2 #(
		.INIT('h1)
	) name4588 (
		_w6732_,
		_w6733_,
		_w6734_
	);
	LUT2 #(
		.INIT('h2)
	) name4589 (
		\u3_mem_reg[3][22]/NET0131 ,
		_w6319_,
		_w6735_
	);
	LUT2 #(
		.INIT('h8)
	) name4590 (
		\u12_dout_reg[22]/P0001 ,
		_w6319_,
		_w6736_
	);
	LUT2 #(
		.INIT('h1)
	) name4591 (
		_w6735_,
		_w6736_,
		_w6737_
	);
	LUT2 #(
		.INIT('h2)
	) name4592 (
		\u3_mem_reg[3][23]/NET0131 ,
		_w6319_,
		_w6738_
	);
	LUT2 #(
		.INIT('h8)
	) name4593 (
		\u12_dout_reg[23]/P0001 ,
		_w6319_,
		_w6739_
	);
	LUT2 #(
		.INIT('h1)
	) name4594 (
		_w6738_,
		_w6739_,
		_w6740_
	);
	LUT2 #(
		.INIT('h2)
	) name4595 (
		\u3_mem_reg[3][24]/NET0131 ,
		_w6319_,
		_w6741_
	);
	LUT2 #(
		.INIT('h8)
	) name4596 (
		\u12_dout_reg[24]/P0001 ,
		_w6319_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name4597 (
		_w6741_,
		_w6742_,
		_w6743_
	);
	LUT2 #(
		.INIT('h2)
	) name4598 (
		\u3_mem_reg[3][26]/NET0131 ,
		_w6319_,
		_w6744_
	);
	LUT2 #(
		.INIT('h8)
	) name4599 (
		\u12_dout_reg[26]/P0001 ,
		_w6319_,
		_w6745_
	);
	LUT2 #(
		.INIT('h1)
	) name4600 (
		_w6744_,
		_w6745_,
		_w6746_
	);
	LUT2 #(
		.INIT('h2)
	) name4601 (
		\u3_mem_reg[3][27]/NET0131 ,
		_w6319_,
		_w6747_
	);
	LUT2 #(
		.INIT('h8)
	) name4602 (
		\u12_dout_reg[27]/P0001 ,
		_w6319_,
		_w6748_
	);
	LUT2 #(
		.INIT('h1)
	) name4603 (
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h2)
	) name4604 (
		\u8_mem_reg[3][28]/NET0131 ,
		_w6301_,
		_w6750_
	);
	LUT2 #(
		.INIT('h8)
	) name4605 (
		\u12_dout_reg[28]/P0001 ,
		_w6301_,
		_w6751_
	);
	LUT2 #(
		.INIT('h1)
	) name4606 (
		_w6750_,
		_w6751_,
		_w6752_
	);
	LUT2 #(
		.INIT('h2)
	) name4607 (
		\u3_mem_reg[3][28]/NET0131 ,
		_w6319_,
		_w6753_
	);
	LUT2 #(
		.INIT('h8)
	) name4608 (
		\u12_dout_reg[28]/P0001 ,
		_w6319_,
		_w6754_
	);
	LUT2 #(
		.INIT('h1)
	) name4609 (
		_w6753_,
		_w6754_,
		_w6755_
	);
	LUT2 #(
		.INIT('h2)
	) name4610 (
		\u3_mem_reg[3][29]/NET0131 ,
		_w6319_,
		_w6756_
	);
	LUT2 #(
		.INIT('h8)
	) name4611 (
		\u12_dout_reg[29]/P0001 ,
		_w6319_,
		_w6757_
	);
	LUT2 #(
		.INIT('h1)
	) name4612 (
		_w6756_,
		_w6757_,
		_w6758_
	);
	LUT2 #(
		.INIT('h2)
	) name4613 (
		\u3_mem_reg[3][2]/NET0131 ,
		_w6319_,
		_w6759_
	);
	LUT2 #(
		.INIT('h8)
	) name4614 (
		\u12_dout_reg[2]/P0001 ,
		_w6319_,
		_w6760_
	);
	LUT2 #(
		.INIT('h1)
	) name4615 (
		_w6759_,
		_w6760_,
		_w6761_
	);
	LUT2 #(
		.INIT('h2)
	) name4616 (
		\u3_mem_reg[3][30]/NET0131 ,
		_w6319_,
		_w6762_
	);
	LUT2 #(
		.INIT('h8)
	) name4617 (
		\u12_dout_reg[30]/P0001 ,
		_w6319_,
		_w6763_
	);
	LUT2 #(
		.INIT('h1)
	) name4618 (
		_w6762_,
		_w6763_,
		_w6764_
	);
	LUT2 #(
		.INIT('h2)
	) name4619 (
		\u3_mem_reg[3][31]/NET0131 ,
		_w6319_,
		_w6765_
	);
	LUT2 #(
		.INIT('h8)
	) name4620 (
		\u12_dout_reg[31]/P0001 ,
		_w6319_,
		_w6766_
	);
	LUT2 #(
		.INIT('h1)
	) name4621 (
		_w6765_,
		_w6766_,
		_w6767_
	);
	LUT2 #(
		.INIT('h2)
	) name4622 (
		\u3_mem_reg[3][4]/NET0131 ,
		_w6319_,
		_w6768_
	);
	LUT2 #(
		.INIT('h8)
	) name4623 (
		\u12_dout_reg[4]/P0001 ,
		_w6319_,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name4624 (
		_w6768_,
		_w6769_,
		_w6770_
	);
	LUT2 #(
		.INIT('h2)
	) name4625 (
		\u3_mem_reg[3][5]/NET0131 ,
		_w6319_,
		_w6771_
	);
	LUT2 #(
		.INIT('h8)
	) name4626 (
		\u12_dout_reg[5]/P0001 ,
		_w6319_,
		_w6772_
	);
	LUT2 #(
		.INIT('h1)
	) name4627 (
		_w6771_,
		_w6772_,
		_w6773_
	);
	LUT2 #(
		.INIT('h2)
	) name4628 (
		\u3_mem_reg[1][1]/NET0131 ,
		_w6489_,
		_w6774_
	);
	LUT2 #(
		.INIT('h8)
	) name4629 (
		\u12_dout_reg[1]/P0001 ,
		_w6489_,
		_w6775_
	);
	LUT2 #(
		.INIT('h1)
	) name4630 (
		_w6774_,
		_w6775_,
		_w6776_
	);
	LUT2 #(
		.INIT('h2)
	) name4631 (
		\u3_mem_reg[3][6]/NET0131 ,
		_w6319_,
		_w6777_
	);
	LUT2 #(
		.INIT('h8)
	) name4632 (
		\u12_dout_reg[6]/P0001 ,
		_w6319_,
		_w6778_
	);
	LUT2 #(
		.INIT('h1)
	) name4633 (
		_w6777_,
		_w6778_,
		_w6779_
	);
	LUT2 #(
		.INIT('h2)
	) name4634 (
		\u3_mem_reg[3][7]/NET0131 ,
		_w6319_,
		_w6780_
	);
	LUT2 #(
		.INIT('h8)
	) name4635 (
		\u12_dout_reg[7]/P0001 ,
		_w6319_,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name4636 (
		_w6780_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h2)
	) name4637 (
		\u3_mem_reg[3][8]/NET0131 ,
		_w6319_,
		_w6783_
	);
	LUT2 #(
		.INIT('h8)
	) name4638 (
		\u12_dout_reg[8]/P0001 ,
		_w6319_,
		_w6784_
	);
	LUT2 #(
		.INIT('h1)
	) name4639 (
		_w6783_,
		_w6784_,
		_w6785_
	);
	LUT2 #(
		.INIT('h2)
	) name4640 (
		\u3_mem_reg[3][9]/NET0131 ,
		_w6319_,
		_w6786_
	);
	LUT2 #(
		.INIT('h8)
	) name4641 (
		\u12_dout_reg[9]/P0001 ,
		_w6319_,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name4642 (
		_w6786_,
		_w6787_,
		_w6788_
	);
	LUT2 #(
		.INIT('h2)
	) name4643 (
		\u8_mem_reg[1][31]/NET0131 ,
		_w6629_,
		_w6789_
	);
	LUT2 #(
		.INIT('h8)
	) name4644 (
		\u12_dout_reg[31]/P0001 ,
		_w6629_,
		_w6790_
	);
	LUT2 #(
		.INIT('h1)
	) name4645 (
		_w6789_,
		_w6790_,
		_w6791_
	);
	LUT2 #(
		.INIT('h2)
	) name4646 (
		\u8_mem_reg[3][26]/NET0131 ,
		_w6301_,
		_w6792_
	);
	LUT2 #(
		.INIT('h8)
	) name4647 (
		\u12_dout_reg[26]/P0001 ,
		_w6301_,
		_w6793_
	);
	LUT2 #(
		.INIT('h1)
	) name4648 (
		_w6792_,
		_w6793_,
		_w6794_
	);
	LUT2 #(
		.INIT('h2)
	) name4649 (
		\u8_mem_reg[2][3]/NET0131 ,
		_w6485_,
		_w6795_
	);
	LUT2 #(
		.INIT('h8)
	) name4650 (
		\u12_dout_reg[3]/P0001 ,
		_w6485_,
		_w6796_
	);
	LUT2 #(
		.INIT('h1)
	) name4651 (
		_w6795_,
		_w6796_,
		_w6797_
	);
	LUT2 #(
		.INIT('h2)
	) name4652 (
		\u3_mem_reg[3][25]/NET0131 ,
		_w6319_,
		_w6798_
	);
	LUT2 #(
		.INIT('h8)
	) name4653 (
		\u12_dout_reg[25]/P0001 ,
		_w6319_,
		_w6799_
	);
	LUT2 #(
		.INIT('h1)
	) name4654 (
		_w6798_,
		_w6799_,
		_w6800_
	);
	LUT2 #(
		.INIT('h2)
	) name4655 (
		\u3_mem_reg[1][27]/NET0131 ,
		_w6489_,
		_w6801_
	);
	LUT2 #(
		.INIT('h8)
	) name4656 (
		\u12_dout_reg[27]/P0001 ,
		_w6489_,
		_w6802_
	);
	LUT2 #(
		.INIT('h1)
	) name4657 (
		_w6801_,
		_w6802_,
		_w6803_
	);
	LUT2 #(
		.INIT('h2)
	) name4658 (
		\u3_mem_reg[2][23]/NET0131 ,
		_w6583_,
		_w6804_
	);
	LUT2 #(
		.INIT('h8)
	) name4659 (
		\u12_dout_reg[23]/P0001 ,
		_w6583_,
		_w6805_
	);
	LUT2 #(
		.INIT('h1)
	) name4660 (
		_w6804_,
		_w6805_,
		_w6806_
	);
	LUT2 #(
		.INIT('h4)
	) name4661 (
		\u4_wp_reg[1]/NET0131 ,
		_w6306_,
		_w6807_
	);
	LUT2 #(
		.INIT('h2)
	) name4662 (
		\u4_mem_reg[1][0]/NET0131 ,
		_w6807_,
		_w6808_
	);
	LUT2 #(
		.INIT('h8)
	) name4663 (
		\u12_dout_reg[0]/P0001 ,
		_w6807_,
		_w6809_
	);
	LUT2 #(
		.INIT('h1)
	) name4664 (
		_w6808_,
		_w6809_,
		_w6810_
	);
	LUT2 #(
		.INIT('h2)
	) name4665 (
		\u4_mem_reg[1][10]/NET0131 ,
		_w6807_,
		_w6811_
	);
	LUT2 #(
		.INIT('h8)
	) name4666 (
		\u12_dout_reg[10]/P0001 ,
		_w6807_,
		_w6812_
	);
	LUT2 #(
		.INIT('h1)
	) name4667 (
		_w6811_,
		_w6812_,
		_w6813_
	);
	LUT2 #(
		.INIT('h2)
	) name4668 (
		\u4_mem_reg[1][11]/NET0131 ,
		_w6807_,
		_w6814_
	);
	LUT2 #(
		.INIT('h8)
	) name4669 (
		\u12_dout_reg[11]/P0001 ,
		_w6807_,
		_w6815_
	);
	LUT2 #(
		.INIT('h1)
	) name4670 (
		_w6814_,
		_w6815_,
		_w6816_
	);
	LUT2 #(
		.INIT('h2)
	) name4671 (
		\u4_mem_reg[1][12]/NET0131 ,
		_w6807_,
		_w6817_
	);
	LUT2 #(
		.INIT('h8)
	) name4672 (
		\u12_dout_reg[12]/P0001 ,
		_w6807_,
		_w6818_
	);
	LUT2 #(
		.INIT('h1)
	) name4673 (
		_w6817_,
		_w6818_,
		_w6819_
	);
	LUT2 #(
		.INIT('h2)
	) name4674 (
		\u4_mem_reg[1][13]/NET0131 ,
		_w6807_,
		_w6820_
	);
	LUT2 #(
		.INIT('h8)
	) name4675 (
		\u12_dout_reg[13]/P0001 ,
		_w6807_,
		_w6821_
	);
	LUT2 #(
		.INIT('h1)
	) name4676 (
		_w6820_,
		_w6821_,
		_w6822_
	);
	LUT2 #(
		.INIT('h2)
	) name4677 (
		\u4_mem_reg[1][14]/NET0131 ,
		_w6807_,
		_w6823_
	);
	LUT2 #(
		.INIT('h8)
	) name4678 (
		\u12_dout_reg[14]/P0001 ,
		_w6807_,
		_w6824_
	);
	LUT2 #(
		.INIT('h1)
	) name4679 (
		_w6823_,
		_w6824_,
		_w6825_
	);
	LUT2 #(
		.INIT('h2)
	) name4680 (
		\u4_mem_reg[1][15]/NET0131 ,
		_w6807_,
		_w6826_
	);
	LUT2 #(
		.INIT('h8)
	) name4681 (
		\u12_dout_reg[15]/P0001 ,
		_w6807_,
		_w6827_
	);
	LUT2 #(
		.INIT('h1)
	) name4682 (
		_w6826_,
		_w6827_,
		_w6828_
	);
	LUT2 #(
		.INIT('h2)
	) name4683 (
		\u4_mem_reg[1][16]/NET0131 ,
		_w6807_,
		_w6829_
	);
	LUT2 #(
		.INIT('h8)
	) name4684 (
		\u12_dout_reg[16]/P0001 ,
		_w6807_,
		_w6830_
	);
	LUT2 #(
		.INIT('h1)
	) name4685 (
		_w6829_,
		_w6830_,
		_w6831_
	);
	LUT2 #(
		.INIT('h2)
	) name4686 (
		\u4_mem_reg[1][17]/NET0131 ,
		_w6807_,
		_w6832_
	);
	LUT2 #(
		.INIT('h8)
	) name4687 (
		\u12_dout_reg[17]/P0001 ,
		_w6807_,
		_w6833_
	);
	LUT2 #(
		.INIT('h1)
	) name4688 (
		_w6832_,
		_w6833_,
		_w6834_
	);
	LUT2 #(
		.INIT('h2)
	) name4689 (
		\u4_mem_reg[1][18]/NET0131 ,
		_w6807_,
		_w6835_
	);
	LUT2 #(
		.INIT('h8)
	) name4690 (
		\u12_dout_reg[18]/P0001 ,
		_w6807_,
		_w6836_
	);
	LUT2 #(
		.INIT('h1)
	) name4691 (
		_w6835_,
		_w6836_,
		_w6837_
	);
	LUT2 #(
		.INIT('h2)
	) name4692 (
		\u4_mem_reg[1][19]/NET0131 ,
		_w6807_,
		_w6838_
	);
	LUT2 #(
		.INIT('h8)
	) name4693 (
		\u12_dout_reg[19]/P0001 ,
		_w6807_,
		_w6839_
	);
	LUT2 #(
		.INIT('h1)
	) name4694 (
		_w6838_,
		_w6839_,
		_w6840_
	);
	LUT2 #(
		.INIT('h2)
	) name4695 (
		\u4_mem_reg[1][1]/NET0131 ,
		_w6807_,
		_w6841_
	);
	LUT2 #(
		.INIT('h8)
	) name4696 (
		\u12_dout_reg[1]/P0001 ,
		_w6807_,
		_w6842_
	);
	LUT2 #(
		.INIT('h1)
	) name4697 (
		_w6841_,
		_w6842_,
		_w6843_
	);
	LUT2 #(
		.INIT('h2)
	) name4698 (
		\u4_mem_reg[1][20]/NET0131 ,
		_w6807_,
		_w6844_
	);
	LUT2 #(
		.INIT('h8)
	) name4699 (
		\u12_dout_reg[20]/P0001 ,
		_w6807_,
		_w6845_
	);
	LUT2 #(
		.INIT('h1)
	) name4700 (
		_w6844_,
		_w6845_,
		_w6846_
	);
	LUT2 #(
		.INIT('h2)
	) name4701 (
		\u4_mem_reg[1][21]/NET0131 ,
		_w6807_,
		_w6847_
	);
	LUT2 #(
		.INIT('h8)
	) name4702 (
		\u12_dout_reg[21]/P0001 ,
		_w6807_,
		_w6848_
	);
	LUT2 #(
		.INIT('h1)
	) name4703 (
		_w6847_,
		_w6848_,
		_w6849_
	);
	LUT2 #(
		.INIT('h2)
	) name4704 (
		\u4_mem_reg[1][22]/NET0131 ,
		_w6807_,
		_w6850_
	);
	LUT2 #(
		.INIT('h8)
	) name4705 (
		\u12_dout_reg[22]/P0001 ,
		_w6807_,
		_w6851_
	);
	LUT2 #(
		.INIT('h1)
	) name4706 (
		_w6850_,
		_w6851_,
		_w6852_
	);
	LUT2 #(
		.INIT('h2)
	) name4707 (
		\u4_mem_reg[1][23]/NET0131 ,
		_w6807_,
		_w6853_
	);
	LUT2 #(
		.INIT('h8)
	) name4708 (
		\u12_dout_reg[23]/P0001 ,
		_w6807_,
		_w6854_
	);
	LUT2 #(
		.INIT('h1)
	) name4709 (
		_w6853_,
		_w6854_,
		_w6855_
	);
	LUT2 #(
		.INIT('h2)
	) name4710 (
		\u4_mem_reg[1][24]/NET0131 ,
		_w6807_,
		_w6856_
	);
	LUT2 #(
		.INIT('h8)
	) name4711 (
		\u12_dout_reg[24]/P0001 ,
		_w6807_,
		_w6857_
	);
	LUT2 #(
		.INIT('h1)
	) name4712 (
		_w6856_,
		_w6857_,
		_w6858_
	);
	LUT2 #(
		.INIT('h2)
	) name4713 (
		\u4_mem_reg[1][25]/NET0131 ,
		_w6807_,
		_w6859_
	);
	LUT2 #(
		.INIT('h8)
	) name4714 (
		\u12_dout_reg[25]/P0001 ,
		_w6807_,
		_w6860_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w6859_,
		_w6860_,
		_w6861_
	);
	LUT2 #(
		.INIT('h2)
	) name4716 (
		\u4_mem_reg[1][26]/NET0131 ,
		_w6807_,
		_w6862_
	);
	LUT2 #(
		.INIT('h8)
	) name4717 (
		\u12_dout_reg[26]/P0001 ,
		_w6807_,
		_w6863_
	);
	LUT2 #(
		.INIT('h1)
	) name4718 (
		_w6862_,
		_w6863_,
		_w6864_
	);
	LUT2 #(
		.INIT('h2)
	) name4719 (
		\u4_mem_reg[1][27]/NET0131 ,
		_w6807_,
		_w6865_
	);
	LUT2 #(
		.INIT('h8)
	) name4720 (
		\u12_dout_reg[27]/P0001 ,
		_w6807_,
		_w6866_
	);
	LUT2 #(
		.INIT('h1)
	) name4721 (
		_w6865_,
		_w6866_,
		_w6867_
	);
	LUT2 #(
		.INIT('h2)
	) name4722 (
		\u4_mem_reg[1][28]/NET0131 ,
		_w6807_,
		_w6868_
	);
	LUT2 #(
		.INIT('h8)
	) name4723 (
		\u12_dout_reg[28]/P0001 ,
		_w6807_,
		_w6869_
	);
	LUT2 #(
		.INIT('h1)
	) name4724 (
		_w6868_,
		_w6869_,
		_w6870_
	);
	LUT2 #(
		.INIT('h2)
	) name4725 (
		\u4_mem_reg[1][29]/NET0131 ,
		_w6807_,
		_w6871_
	);
	LUT2 #(
		.INIT('h8)
	) name4726 (
		\u12_dout_reg[29]/P0001 ,
		_w6807_,
		_w6872_
	);
	LUT2 #(
		.INIT('h1)
	) name4727 (
		_w6871_,
		_w6872_,
		_w6873_
	);
	LUT2 #(
		.INIT('h2)
	) name4728 (
		\u4_mem_reg[1][2]/NET0131 ,
		_w6807_,
		_w6874_
	);
	LUT2 #(
		.INIT('h8)
	) name4729 (
		\u12_dout_reg[2]/P0001 ,
		_w6807_,
		_w6875_
	);
	LUT2 #(
		.INIT('h1)
	) name4730 (
		_w6874_,
		_w6875_,
		_w6876_
	);
	LUT2 #(
		.INIT('h2)
	) name4731 (
		\u4_mem_reg[1][30]/NET0131 ,
		_w6807_,
		_w6877_
	);
	LUT2 #(
		.INIT('h8)
	) name4732 (
		\u12_dout_reg[30]/P0001 ,
		_w6807_,
		_w6878_
	);
	LUT2 #(
		.INIT('h1)
	) name4733 (
		_w6877_,
		_w6878_,
		_w6879_
	);
	LUT2 #(
		.INIT('h2)
	) name4734 (
		\u4_mem_reg[1][31]/NET0131 ,
		_w6807_,
		_w6880_
	);
	LUT2 #(
		.INIT('h8)
	) name4735 (
		\u12_dout_reg[31]/P0001 ,
		_w6807_,
		_w6881_
	);
	LUT2 #(
		.INIT('h1)
	) name4736 (
		_w6880_,
		_w6881_,
		_w6882_
	);
	LUT2 #(
		.INIT('h2)
	) name4737 (
		\u4_mem_reg[1][3]/NET0131 ,
		_w6807_,
		_w6883_
	);
	LUT2 #(
		.INIT('h8)
	) name4738 (
		\u12_dout_reg[3]/P0001 ,
		_w6807_,
		_w6884_
	);
	LUT2 #(
		.INIT('h1)
	) name4739 (
		_w6883_,
		_w6884_,
		_w6885_
	);
	LUT2 #(
		.INIT('h2)
	) name4740 (
		\u4_mem_reg[1][4]/NET0131 ,
		_w6807_,
		_w6886_
	);
	LUT2 #(
		.INIT('h8)
	) name4741 (
		\u12_dout_reg[4]/P0001 ,
		_w6807_,
		_w6887_
	);
	LUT2 #(
		.INIT('h1)
	) name4742 (
		_w6886_,
		_w6887_,
		_w6888_
	);
	LUT2 #(
		.INIT('h2)
	) name4743 (
		\u4_mem_reg[1][5]/NET0131 ,
		_w6807_,
		_w6889_
	);
	LUT2 #(
		.INIT('h8)
	) name4744 (
		\u12_dout_reg[5]/P0001 ,
		_w6807_,
		_w6890_
	);
	LUT2 #(
		.INIT('h1)
	) name4745 (
		_w6889_,
		_w6890_,
		_w6891_
	);
	LUT2 #(
		.INIT('h2)
	) name4746 (
		\u4_mem_reg[1][6]/NET0131 ,
		_w6807_,
		_w6892_
	);
	LUT2 #(
		.INIT('h8)
	) name4747 (
		\u12_dout_reg[6]/P0001 ,
		_w6807_,
		_w6893_
	);
	LUT2 #(
		.INIT('h1)
	) name4748 (
		_w6892_,
		_w6893_,
		_w6894_
	);
	LUT2 #(
		.INIT('h2)
	) name4749 (
		\u4_mem_reg[1][7]/NET0131 ,
		_w6807_,
		_w6895_
	);
	LUT2 #(
		.INIT('h8)
	) name4750 (
		\u12_dout_reg[7]/P0001 ,
		_w6807_,
		_w6896_
	);
	LUT2 #(
		.INIT('h1)
	) name4751 (
		_w6895_,
		_w6896_,
		_w6897_
	);
	LUT2 #(
		.INIT('h2)
	) name4752 (
		\u4_mem_reg[1][8]/NET0131 ,
		_w6807_,
		_w6898_
	);
	LUT2 #(
		.INIT('h8)
	) name4753 (
		\u12_dout_reg[8]/P0001 ,
		_w6807_,
		_w6899_
	);
	LUT2 #(
		.INIT('h1)
	) name4754 (
		_w6898_,
		_w6899_,
		_w6900_
	);
	LUT2 #(
		.INIT('h2)
	) name4755 (
		\u4_mem_reg[1][9]/NET0131 ,
		_w6807_,
		_w6901_
	);
	LUT2 #(
		.INIT('h8)
	) name4756 (
		\u12_dout_reg[9]/P0001 ,
		_w6807_,
		_w6902_
	);
	LUT2 #(
		.INIT('h1)
	) name4757 (
		_w6901_,
		_w6902_,
		_w6903_
	);
	LUT2 #(
		.INIT('h8)
	) name4758 (
		\u4_wp_reg[1]/NET0131 ,
		_w6411_,
		_w6904_
	);
	LUT2 #(
		.INIT('h2)
	) name4759 (
		\u4_mem_reg[2][0]/NET0131 ,
		_w6904_,
		_w6905_
	);
	LUT2 #(
		.INIT('h8)
	) name4760 (
		\u12_dout_reg[0]/P0001 ,
		_w6904_,
		_w6906_
	);
	LUT2 #(
		.INIT('h1)
	) name4761 (
		_w6905_,
		_w6906_,
		_w6907_
	);
	LUT2 #(
		.INIT('h2)
	) name4762 (
		\u4_mem_reg[2][10]/NET0131 ,
		_w6904_,
		_w6908_
	);
	LUT2 #(
		.INIT('h8)
	) name4763 (
		\u12_dout_reg[10]/P0001 ,
		_w6904_,
		_w6909_
	);
	LUT2 #(
		.INIT('h1)
	) name4764 (
		_w6908_,
		_w6909_,
		_w6910_
	);
	LUT2 #(
		.INIT('h2)
	) name4765 (
		\u4_mem_reg[2][11]/NET0131 ,
		_w6904_,
		_w6911_
	);
	LUT2 #(
		.INIT('h8)
	) name4766 (
		\u12_dout_reg[11]/P0001 ,
		_w6904_,
		_w6912_
	);
	LUT2 #(
		.INIT('h1)
	) name4767 (
		_w6911_,
		_w6912_,
		_w6913_
	);
	LUT2 #(
		.INIT('h2)
	) name4768 (
		\u4_mem_reg[2][12]/NET0131 ,
		_w6904_,
		_w6914_
	);
	LUT2 #(
		.INIT('h8)
	) name4769 (
		\u12_dout_reg[12]/P0001 ,
		_w6904_,
		_w6915_
	);
	LUT2 #(
		.INIT('h1)
	) name4770 (
		_w6914_,
		_w6915_,
		_w6916_
	);
	LUT2 #(
		.INIT('h2)
	) name4771 (
		\u4_mem_reg[2][13]/NET0131 ,
		_w6904_,
		_w6917_
	);
	LUT2 #(
		.INIT('h8)
	) name4772 (
		\u12_dout_reg[13]/P0001 ,
		_w6904_,
		_w6918_
	);
	LUT2 #(
		.INIT('h1)
	) name4773 (
		_w6917_,
		_w6918_,
		_w6919_
	);
	LUT2 #(
		.INIT('h2)
	) name4774 (
		\u4_mem_reg[2][14]/NET0131 ,
		_w6904_,
		_w6920_
	);
	LUT2 #(
		.INIT('h8)
	) name4775 (
		\u12_dout_reg[14]/P0001 ,
		_w6904_,
		_w6921_
	);
	LUT2 #(
		.INIT('h1)
	) name4776 (
		_w6920_,
		_w6921_,
		_w6922_
	);
	LUT2 #(
		.INIT('h2)
	) name4777 (
		\u4_mem_reg[2][15]/NET0131 ,
		_w6904_,
		_w6923_
	);
	LUT2 #(
		.INIT('h8)
	) name4778 (
		\u12_dout_reg[15]/P0001 ,
		_w6904_,
		_w6924_
	);
	LUT2 #(
		.INIT('h1)
	) name4779 (
		_w6923_,
		_w6924_,
		_w6925_
	);
	LUT2 #(
		.INIT('h2)
	) name4780 (
		\u4_mem_reg[2][16]/NET0131 ,
		_w6904_,
		_w6926_
	);
	LUT2 #(
		.INIT('h8)
	) name4781 (
		\u12_dout_reg[16]/P0001 ,
		_w6904_,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name4782 (
		_w6926_,
		_w6927_,
		_w6928_
	);
	LUT2 #(
		.INIT('h2)
	) name4783 (
		\u4_mem_reg[2][17]/NET0131 ,
		_w6904_,
		_w6929_
	);
	LUT2 #(
		.INIT('h8)
	) name4784 (
		\u12_dout_reg[17]/P0001 ,
		_w6904_,
		_w6930_
	);
	LUT2 #(
		.INIT('h1)
	) name4785 (
		_w6929_,
		_w6930_,
		_w6931_
	);
	LUT2 #(
		.INIT('h2)
	) name4786 (
		\u4_mem_reg[2][18]/NET0131 ,
		_w6904_,
		_w6932_
	);
	LUT2 #(
		.INIT('h8)
	) name4787 (
		\u12_dout_reg[18]/P0001 ,
		_w6904_,
		_w6933_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		_w6932_,
		_w6933_,
		_w6934_
	);
	LUT2 #(
		.INIT('h2)
	) name4789 (
		\u4_mem_reg[2][19]/NET0131 ,
		_w6904_,
		_w6935_
	);
	LUT2 #(
		.INIT('h8)
	) name4790 (
		\u12_dout_reg[19]/P0001 ,
		_w6904_,
		_w6936_
	);
	LUT2 #(
		.INIT('h1)
	) name4791 (
		_w6935_,
		_w6936_,
		_w6937_
	);
	LUT2 #(
		.INIT('h2)
	) name4792 (
		\u4_mem_reg[2][1]/NET0131 ,
		_w6904_,
		_w6938_
	);
	LUT2 #(
		.INIT('h8)
	) name4793 (
		\u12_dout_reg[1]/P0001 ,
		_w6904_,
		_w6939_
	);
	LUT2 #(
		.INIT('h1)
	) name4794 (
		_w6938_,
		_w6939_,
		_w6940_
	);
	LUT2 #(
		.INIT('h2)
	) name4795 (
		\u4_mem_reg[2][20]/NET0131 ,
		_w6904_,
		_w6941_
	);
	LUT2 #(
		.INIT('h8)
	) name4796 (
		\u12_dout_reg[20]/P0001 ,
		_w6904_,
		_w6942_
	);
	LUT2 #(
		.INIT('h1)
	) name4797 (
		_w6941_,
		_w6942_,
		_w6943_
	);
	LUT2 #(
		.INIT('h2)
	) name4798 (
		\u4_mem_reg[2][21]/NET0131 ,
		_w6904_,
		_w6944_
	);
	LUT2 #(
		.INIT('h8)
	) name4799 (
		\u12_dout_reg[21]/P0001 ,
		_w6904_,
		_w6945_
	);
	LUT2 #(
		.INIT('h1)
	) name4800 (
		_w6944_,
		_w6945_,
		_w6946_
	);
	LUT2 #(
		.INIT('h2)
	) name4801 (
		\u4_mem_reg[2][22]/NET0131 ,
		_w6904_,
		_w6947_
	);
	LUT2 #(
		.INIT('h8)
	) name4802 (
		\u12_dout_reg[22]/P0001 ,
		_w6904_,
		_w6948_
	);
	LUT2 #(
		.INIT('h1)
	) name4803 (
		_w6947_,
		_w6948_,
		_w6949_
	);
	LUT2 #(
		.INIT('h2)
	) name4804 (
		\u4_mem_reg[2][23]/NET0131 ,
		_w6904_,
		_w6950_
	);
	LUT2 #(
		.INIT('h8)
	) name4805 (
		\u12_dout_reg[23]/P0001 ,
		_w6904_,
		_w6951_
	);
	LUT2 #(
		.INIT('h1)
	) name4806 (
		_w6950_,
		_w6951_,
		_w6952_
	);
	LUT2 #(
		.INIT('h2)
	) name4807 (
		\u4_mem_reg[2][24]/NET0131 ,
		_w6904_,
		_w6953_
	);
	LUT2 #(
		.INIT('h8)
	) name4808 (
		\u12_dout_reg[24]/P0001 ,
		_w6904_,
		_w6954_
	);
	LUT2 #(
		.INIT('h1)
	) name4809 (
		_w6953_,
		_w6954_,
		_w6955_
	);
	LUT2 #(
		.INIT('h2)
	) name4810 (
		\u4_mem_reg[2][25]/NET0131 ,
		_w6904_,
		_w6956_
	);
	LUT2 #(
		.INIT('h8)
	) name4811 (
		\u12_dout_reg[25]/P0001 ,
		_w6904_,
		_w6957_
	);
	LUT2 #(
		.INIT('h1)
	) name4812 (
		_w6956_,
		_w6957_,
		_w6958_
	);
	LUT2 #(
		.INIT('h2)
	) name4813 (
		\u4_mem_reg[2][26]/NET0131 ,
		_w6904_,
		_w6959_
	);
	LUT2 #(
		.INIT('h8)
	) name4814 (
		\u12_dout_reg[26]/P0001 ,
		_w6904_,
		_w6960_
	);
	LUT2 #(
		.INIT('h1)
	) name4815 (
		_w6959_,
		_w6960_,
		_w6961_
	);
	LUT2 #(
		.INIT('h2)
	) name4816 (
		\u4_mem_reg[2][27]/NET0131 ,
		_w6904_,
		_w6962_
	);
	LUT2 #(
		.INIT('h8)
	) name4817 (
		\u12_dout_reg[27]/P0001 ,
		_w6904_,
		_w6963_
	);
	LUT2 #(
		.INIT('h1)
	) name4818 (
		_w6962_,
		_w6963_,
		_w6964_
	);
	LUT2 #(
		.INIT('h2)
	) name4819 (
		\u4_mem_reg[2][28]/NET0131 ,
		_w6904_,
		_w6965_
	);
	LUT2 #(
		.INIT('h8)
	) name4820 (
		\u12_dout_reg[28]/P0001 ,
		_w6904_,
		_w6966_
	);
	LUT2 #(
		.INIT('h1)
	) name4821 (
		_w6965_,
		_w6966_,
		_w6967_
	);
	LUT2 #(
		.INIT('h2)
	) name4822 (
		\u4_mem_reg[2][29]/NET0131 ,
		_w6904_,
		_w6968_
	);
	LUT2 #(
		.INIT('h8)
	) name4823 (
		\u12_dout_reg[29]/P0001 ,
		_w6904_,
		_w6969_
	);
	LUT2 #(
		.INIT('h1)
	) name4824 (
		_w6968_,
		_w6969_,
		_w6970_
	);
	LUT2 #(
		.INIT('h2)
	) name4825 (
		\u4_mem_reg[2][2]/NET0131 ,
		_w6904_,
		_w6971_
	);
	LUT2 #(
		.INIT('h8)
	) name4826 (
		\u12_dout_reg[2]/P0001 ,
		_w6904_,
		_w6972_
	);
	LUT2 #(
		.INIT('h1)
	) name4827 (
		_w6971_,
		_w6972_,
		_w6973_
	);
	LUT2 #(
		.INIT('h2)
	) name4828 (
		\u4_mem_reg[2][30]/NET0131 ,
		_w6904_,
		_w6974_
	);
	LUT2 #(
		.INIT('h8)
	) name4829 (
		\u12_dout_reg[30]/P0001 ,
		_w6904_,
		_w6975_
	);
	LUT2 #(
		.INIT('h1)
	) name4830 (
		_w6974_,
		_w6975_,
		_w6976_
	);
	LUT2 #(
		.INIT('h2)
	) name4831 (
		\u4_mem_reg[2][31]/NET0131 ,
		_w6904_,
		_w6977_
	);
	LUT2 #(
		.INIT('h8)
	) name4832 (
		\u12_dout_reg[31]/P0001 ,
		_w6904_,
		_w6978_
	);
	LUT2 #(
		.INIT('h1)
	) name4833 (
		_w6977_,
		_w6978_,
		_w6979_
	);
	LUT2 #(
		.INIT('h2)
	) name4834 (
		\u4_mem_reg[2][3]/NET0131 ,
		_w6904_,
		_w6980_
	);
	LUT2 #(
		.INIT('h8)
	) name4835 (
		\u12_dout_reg[3]/P0001 ,
		_w6904_,
		_w6981_
	);
	LUT2 #(
		.INIT('h1)
	) name4836 (
		_w6980_,
		_w6981_,
		_w6982_
	);
	LUT2 #(
		.INIT('h2)
	) name4837 (
		\u4_mem_reg[2][4]/NET0131 ,
		_w6904_,
		_w6983_
	);
	LUT2 #(
		.INIT('h8)
	) name4838 (
		\u12_dout_reg[4]/P0001 ,
		_w6904_,
		_w6984_
	);
	LUT2 #(
		.INIT('h1)
	) name4839 (
		_w6983_,
		_w6984_,
		_w6985_
	);
	LUT2 #(
		.INIT('h2)
	) name4840 (
		\u4_mem_reg[2][5]/NET0131 ,
		_w6904_,
		_w6986_
	);
	LUT2 #(
		.INIT('h8)
	) name4841 (
		\u12_dout_reg[5]/P0001 ,
		_w6904_,
		_w6987_
	);
	LUT2 #(
		.INIT('h1)
	) name4842 (
		_w6986_,
		_w6987_,
		_w6988_
	);
	LUT2 #(
		.INIT('h2)
	) name4843 (
		\u4_mem_reg[2][6]/NET0131 ,
		_w6904_,
		_w6989_
	);
	LUT2 #(
		.INIT('h8)
	) name4844 (
		\u12_dout_reg[6]/P0001 ,
		_w6904_,
		_w6990_
	);
	LUT2 #(
		.INIT('h1)
	) name4845 (
		_w6989_,
		_w6990_,
		_w6991_
	);
	LUT2 #(
		.INIT('h2)
	) name4846 (
		\u4_mem_reg[2][7]/NET0131 ,
		_w6904_,
		_w6992_
	);
	LUT2 #(
		.INIT('h8)
	) name4847 (
		\u12_dout_reg[7]/P0001 ,
		_w6904_,
		_w6993_
	);
	LUT2 #(
		.INIT('h1)
	) name4848 (
		_w6992_,
		_w6993_,
		_w6994_
	);
	LUT2 #(
		.INIT('h2)
	) name4849 (
		\u4_mem_reg[2][8]/NET0131 ,
		_w6904_,
		_w6995_
	);
	LUT2 #(
		.INIT('h8)
	) name4850 (
		\u12_dout_reg[8]/P0001 ,
		_w6904_,
		_w6996_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		_w6995_,
		_w6996_,
		_w6997_
	);
	LUT2 #(
		.INIT('h2)
	) name4852 (
		\u4_mem_reg[2][9]/NET0131 ,
		_w6904_,
		_w6998_
	);
	LUT2 #(
		.INIT('h8)
	) name4853 (
		\u12_dout_reg[9]/P0001 ,
		_w6904_,
		_w6999_
	);
	LUT2 #(
		.INIT('h1)
	) name4854 (
		_w6998_,
		_w6999_,
		_w7000_
	);
	LUT2 #(
		.INIT('h2)
	) name4855 (
		\u4_mem_reg[3][0]/NET0131 ,
		_w6307_,
		_w7001_
	);
	LUT2 #(
		.INIT('h8)
	) name4856 (
		\u12_dout_reg[0]/P0001 ,
		_w6307_,
		_w7002_
	);
	LUT2 #(
		.INIT('h1)
	) name4857 (
		_w7001_,
		_w7002_,
		_w7003_
	);
	LUT2 #(
		.INIT('h2)
	) name4858 (
		\u4_mem_reg[3][10]/NET0131 ,
		_w6307_,
		_w7004_
	);
	LUT2 #(
		.INIT('h8)
	) name4859 (
		\u12_dout_reg[10]/P0001 ,
		_w6307_,
		_w7005_
	);
	LUT2 #(
		.INIT('h1)
	) name4860 (
		_w7004_,
		_w7005_,
		_w7006_
	);
	LUT2 #(
		.INIT('h2)
	) name4861 (
		\u4_mem_reg[3][11]/NET0131 ,
		_w6307_,
		_w7007_
	);
	LUT2 #(
		.INIT('h8)
	) name4862 (
		\u12_dout_reg[11]/P0001 ,
		_w6307_,
		_w7008_
	);
	LUT2 #(
		.INIT('h1)
	) name4863 (
		_w7007_,
		_w7008_,
		_w7009_
	);
	LUT2 #(
		.INIT('h2)
	) name4864 (
		\u4_mem_reg[3][12]/NET0131 ,
		_w6307_,
		_w7010_
	);
	LUT2 #(
		.INIT('h8)
	) name4865 (
		\u12_dout_reg[12]/P0001 ,
		_w6307_,
		_w7011_
	);
	LUT2 #(
		.INIT('h1)
	) name4866 (
		_w7010_,
		_w7011_,
		_w7012_
	);
	LUT2 #(
		.INIT('h2)
	) name4867 (
		\u4_mem_reg[3][13]/NET0131 ,
		_w6307_,
		_w7013_
	);
	LUT2 #(
		.INIT('h8)
	) name4868 (
		\u12_dout_reg[13]/P0001 ,
		_w6307_,
		_w7014_
	);
	LUT2 #(
		.INIT('h1)
	) name4869 (
		_w7013_,
		_w7014_,
		_w7015_
	);
	LUT2 #(
		.INIT('h2)
	) name4870 (
		\u4_mem_reg[3][14]/NET0131 ,
		_w6307_,
		_w7016_
	);
	LUT2 #(
		.INIT('h8)
	) name4871 (
		\u12_dout_reg[14]/P0001 ,
		_w6307_,
		_w7017_
	);
	LUT2 #(
		.INIT('h1)
	) name4872 (
		_w7016_,
		_w7017_,
		_w7018_
	);
	LUT2 #(
		.INIT('h2)
	) name4873 (
		\u4_mem_reg[3][15]/NET0131 ,
		_w6307_,
		_w7019_
	);
	LUT2 #(
		.INIT('h8)
	) name4874 (
		\u12_dout_reg[15]/P0001 ,
		_w6307_,
		_w7020_
	);
	LUT2 #(
		.INIT('h1)
	) name4875 (
		_w7019_,
		_w7020_,
		_w7021_
	);
	LUT2 #(
		.INIT('h2)
	) name4876 (
		\u4_mem_reg[3][16]/NET0131 ,
		_w6307_,
		_w7022_
	);
	LUT2 #(
		.INIT('h8)
	) name4877 (
		\u12_dout_reg[16]/P0001 ,
		_w6307_,
		_w7023_
	);
	LUT2 #(
		.INIT('h1)
	) name4878 (
		_w7022_,
		_w7023_,
		_w7024_
	);
	LUT2 #(
		.INIT('h2)
	) name4879 (
		\u4_mem_reg[3][17]/NET0131 ,
		_w6307_,
		_w7025_
	);
	LUT2 #(
		.INIT('h8)
	) name4880 (
		\u12_dout_reg[17]/P0001 ,
		_w6307_,
		_w7026_
	);
	LUT2 #(
		.INIT('h1)
	) name4881 (
		_w7025_,
		_w7026_,
		_w7027_
	);
	LUT2 #(
		.INIT('h2)
	) name4882 (
		\u4_mem_reg[3][18]/NET0131 ,
		_w6307_,
		_w7028_
	);
	LUT2 #(
		.INIT('h8)
	) name4883 (
		\u12_dout_reg[18]/P0001 ,
		_w6307_,
		_w7029_
	);
	LUT2 #(
		.INIT('h1)
	) name4884 (
		_w7028_,
		_w7029_,
		_w7030_
	);
	LUT2 #(
		.INIT('h2)
	) name4885 (
		\u4_mem_reg[3][19]/NET0131 ,
		_w6307_,
		_w7031_
	);
	LUT2 #(
		.INIT('h8)
	) name4886 (
		\u12_dout_reg[19]/P0001 ,
		_w6307_,
		_w7032_
	);
	LUT2 #(
		.INIT('h1)
	) name4887 (
		_w7031_,
		_w7032_,
		_w7033_
	);
	LUT2 #(
		.INIT('h2)
	) name4888 (
		\u4_mem_reg[3][1]/NET0131 ,
		_w6307_,
		_w7034_
	);
	LUT2 #(
		.INIT('h8)
	) name4889 (
		\u12_dout_reg[1]/P0001 ,
		_w6307_,
		_w7035_
	);
	LUT2 #(
		.INIT('h1)
	) name4890 (
		_w7034_,
		_w7035_,
		_w7036_
	);
	LUT2 #(
		.INIT('h2)
	) name4891 (
		\u4_mem_reg[3][20]/NET0131 ,
		_w6307_,
		_w7037_
	);
	LUT2 #(
		.INIT('h8)
	) name4892 (
		\u12_dout_reg[20]/P0001 ,
		_w6307_,
		_w7038_
	);
	LUT2 #(
		.INIT('h1)
	) name4893 (
		_w7037_,
		_w7038_,
		_w7039_
	);
	LUT2 #(
		.INIT('h2)
	) name4894 (
		\u4_mem_reg[3][21]/NET0131 ,
		_w6307_,
		_w7040_
	);
	LUT2 #(
		.INIT('h8)
	) name4895 (
		\u12_dout_reg[21]/P0001 ,
		_w6307_,
		_w7041_
	);
	LUT2 #(
		.INIT('h1)
	) name4896 (
		_w7040_,
		_w7041_,
		_w7042_
	);
	LUT2 #(
		.INIT('h2)
	) name4897 (
		\u4_mem_reg[3][22]/NET0131 ,
		_w6307_,
		_w7043_
	);
	LUT2 #(
		.INIT('h8)
	) name4898 (
		\u12_dout_reg[22]/P0001 ,
		_w6307_,
		_w7044_
	);
	LUT2 #(
		.INIT('h1)
	) name4899 (
		_w7043_,
		_w7044_,
		_w7045_
	);
	LUT2 #(
		.INIT('h2)
	) name4900 (
		\u4_mem_reg[3][23]/NET0131 ,
		_w6307_,
		_w7046_
	);
	LUT2 #(
		.INIT('h8)
	) name4901 (
		\u12_dout_reg[23]/P0001 ,
		_w6307_,
		_w7047_
	);
	LUT2 #(
		.INIT('h1)
	) name4902 (
		_w7046_,
		_w7047_,
		_w7048_
	);
	LUT2 #(
		.INIT('h2)
	) name4903 (
		\u4_mem_reg[3][24]/NET0131 ,
		_w6307_,
		_w7049_
	);
	LUT2 #(
		.INIT('h8)
	) name4904 (
		\u12_dout_reg[24]/P0001 ,
		_w6307_,
		_w7050_
	);
	LUT2 #(
		.INIT('h1)
	) name4905 (
		_w7049_,
		_w7050_,
		_w7051_
	);
	LUT2 #(
		.INIT('h2)
	) name4906 (
		\u4_mem_reg[3][25]/NET0131 ,
		_w6307_,
		_w7052_
	);
	LUT2 #(
		.INIT('h8)
	) name4907 (
		\u12_dout_reg[25]/P0001 ,
		_w6307_,
		_w7053_
	);
	LUT2 #(
		.INIT('h1)
	) name4908 (
		_w7052_,
		_w7053_,
		_w7054_
	);
	LUT2 #(
		.INIT('h2)
	) name4909 (
		\u4_mem_reg[3][26]/NET0131 ,
		_w6307_,
		_w7055_
	);
	LUT2 #(
		.INIT('h8)
	) name4910 (
		\u12_dout_reg[26]/P0001 ,
		_w6307_,
		_w7056_
	);
	LUT2 #(
		.INIT('h1)
	) name4911 (
		_w7055_,
		_w7056_,
		_w7057_
	);
	LUT2 #(
		.INIT('h2)
	) name4912 (
		\u4_mem_reg[3][27]/NET0131 ,
		_w6307_,
		_w7058_
	);
	LUT2 #(
		.INIT('h8)
	) name4913 (
		\u12_dout_reg[27]/P0001 ,
		_w6307_,
		_w7059_
	);
	LUT2 #(
		.INIT('h1)
	) name4914 (
		_w7058_,
		_w7059_,
		_w7060_
	);
	LUT2 #(
		.INIT('h2)
	) name4915 (
		\u4_mem_reg[3][28]/NET0131 ,
		_w6307_,
		_w7061_
	);
	LUT2 #(
		.INIT('h8)
	) name4916 (
		\u12_dout_reg[28]/P0001 ,
		_w6307_,
		_w7062_
	);
	LUT2 #(
		.INIT('h1)
	) name4917 (
		_w7061_,
		_w7062_,
		_w7063_
	);
	LUT2 #(
		.INIT('h2)
	) name4918 (
		\u4_mem_reg[3][29]/NET0131 ,
		_w6307_,
		_w7064_
	);
	LUT2 #(
		.INIT('h8)
	) name4919 (
		\u12_dout_reg[29]/P0001 ,
		_w6307_,
		_w7065_
	);
	LUT2 #(
		.INIT('h1)
	) name4920 (
		_w7064_,
		_w7065_,
		_w7066_
	);
	LUT2 #(
		.INIT('h2)
	) name4921 (
		\u4_mem_reg[3][2]/NET0131 ,
		_w6307_,
		_w7067_
	);
	LUT2 #(
		.INIT('h8)
	) name4922 (
		\u12_dout_reg[2]/P0001 ,
		_w6307_,
		_w7068_
	);
	LUT2 #(
		.INIT('h1)
	) name4923 (
		_w7067_,
		_w7068_,
		_w7069_
	);
	LUT2 #(
		.INIT('h2)
	) name4924 (
		\u4_mem_reg[3][30]/NET0131 ,
		_w6307_,
		_w7070_
	);
	LUT2 #(
		.INIT('h8)
	) name4925 (
		\u12_dout_reg[30]/P0001 ,
		_w6307_,
		_w7071_
	);
	LUT2 #(
		.INIT('h1)
	) name4926 (
		_w7070_,
		_w7071_,
		_w7072_
	);
	LUT2 #(
		.INIT('h2)
	) name4927 (
		\u4_mem_reg[3][31]/NET0131 ,
		_w6307_,
		_w7073_
	);
	LUT2 #(
		.INIT('h8)
	) name4928 (
		\u12_dout_reg[31]/P0001 ,
		_w6307_,
		_w7074_
	);
	LUT2 #(
		.INIT('h1)
	) name4929 (
		_w7073_,
		_w7074_,
		_w7075_
	);
	LUT2 #(
		.INIT('h2)
	) name4930 (
		\u4_mem_reg[3][3]/NET0131 ,
		_w6307_,
		_w7076_
	);
	LUT2 #(
		.INIT('h8)
	) name4931 (
		\u12_dout_reg[3]/P0001 ,
		_w6307_,
		_w7077_
	);
	LUT2 #(
		.INIT('h1)
	) name4932 (
		_w7076_,
		_w7077_,
		_w7078_
	);
	LUT2 #(
		.INIT('h2)
	) name4933 (
		\u4_mem_reg[3][4]/NET0131 ,
		_w6307_,
		_w7079_
	);
	LUT2 #(
		.INIT('h8)
	) name4934 (
		\u12_dout_reg[4]/P0001 ,
		_w6307_,
		_w7080_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		_w7079_,
		_w7080_,
		_w7081_
	);
	LUT2 #(
		.INIT('h2)
	) name4936 (
		\u4_mem_reg[3][5]/NET0131 ,
		_w6307_,
		_w7082_
	);
	LUT2 #(
		.INIT('h8)
	) name4937 (
		\u12_dout_reg[5]/P0001 ,
		_w6307_,
		_w7083_
	);
	LUT2 #(
		.INIT('h1)
	) name4938 (
		_w7082_,
		_w7083_,
		_w7084_
	);
	LUT2 #(
		.INIT('h2)
	) name4939 (
		\u4_mem_reg[3][6]/NET0131 ,
		_w6307_,
		_w7085_
	);
	LUT2 #(
		.INIT('h8)
	) name4940 (
		\u12_dout_reg[6]/P0001 ,
		_w6307_,
		_w7086_
	);
	LUT2 #(
		.INIT('h1)
	) name4941 (
		_w7085_,
		_w7086_,
		_w7087_
	);
	LUT2 #(
		.INIT('h2)
	) name4942 (
		\u4_mem_reg[3][7]/NET0131 ,
		_w6307_,
		_w7088_
	);
	LUT2 #(
		.INIT('h8)
	) name4943 (
		\u12_dout_reg[7]/P0001 ,
		_w6307_,
		_w7089_
	);
	LUT2 #(
		.INIT('h1)
	) name4944 (
		_w7088_,
		_w7089_,
		_w7090_
	);
	LUT2 #(
		.INIT('h2)
	) name4945 (
		\u4_mem_reg[3][8]/NET0131 ,
		_w6307_,
		_w7091_
	);
	LUT2 #(
		.INIT('h8)
	) name4946 (
		\u12_dout_reg[8]/P0001 ,
		_w6307_,
		_w7092_
	);
	LUT2 #(
		.INIT('h1)
	) name4947 (
		_w7091_,
		_w7092_,
		_w7093_
	);
	LUT2 #(
		.INIT('h2)
	) name4948 (
		\u4_mem_reg[3][9]/NET0131 ,
		_w6307_,
		_w7094_
	);
	LUT2 #(
		.INIT('h8)
	) name4949 (
		\u12_dout_reg[9]/P0001 ,
		_w6307_,
		_w7095_
	);
	LUT2 #(
		.INIT('h1)
	) name4950 (
		_w7094_,
		_w7095_,
		_w7096_
	);
	LUT2 #(
		.INIT('h2)
	) name4951 (
		\u3_mem_reg[2][14]/NET0131 ,
		_w6583_,
		_w7097_
	);
	LUT2 #(
		.INIT('h8)
	) name4952 (
		\u12_dout_reg[14]/P0001 ,
		_w6583_,
		_w7098_
	);
	LUT2 #(
		.INIT('h1)
	) name4953 (
		_w7097_,
		_w7098_,
		_w7099_
	);
	LUT2 #(
		.INIT('h4)
	) name4954 (
		\u5_wp_reg[1]/NET0131 ,
		_w6312_,
		_w7100_
	);
	LUT2 #(
		.INIT('h2)
	) name4955 (
		\u5_mem_reg[1][0]/NET0131 ,
		_w7100_,
		_w7101_
	);
	LUT2 #(
		.INIT('h8)
	) name4956 (
		\u12_dout_reg[0]/P0001 ,
		_w7100_,
		_w7102_
	);
	LUT2 #(
		.INIT('h1)
	) name4957 (
		_w7101_,
		_w7102_,
		_w7103_
	);
	LUT2 #(
		.INIT('h2)
	) name4958 (
		\u5_mem_reg[1][10]/NET0131 ,
		_w7100_,
		_w7104_
	);
	LUT2 #(
		.INIT('h8)
	) name4959 (
		\u12_dout_reg[10]/P0001 ,
		_w7100_,
		_w7105_
	);
	LUT2 #(
		.INIT('h1)
	) name4960 (
		_w7104_,
		_w7105_,
		_w7106_
	);
	LUT2 #(
		.INIT('h2)
	) name4961 (
		\u5_mem_reg[1][11]/NET0131 ,
		_w7100_,
		_w7107_
	);
	LUT2 #(
		.INIT('h8)
	) name4962 (
		\u12_dout_reg[11]/P0001 ,
		_w7100_,
		_w7108_
	);
	LUT2 #(
		.INIT('h1)
	) name4963 (
		_w7107_,
		_w7108_,
		_w7109_
	);
	LUT2 #(
		.INIT('h2)
	) name4964 (
		\u5_mem_reg[1][12]/NET0131 ,
		_w7100_,
		_w7110_
	);
	LUT2 #(
		.INIT('h8)
	) name4965 (
		\u12_dout_reg[12]/P0001 ,
		_w7100_,
		_w7111_
	);
	LUT2 #(
		.INIT('h1)
	) name4966 (
		_w7110_,
		_w7111_,
		_w7112_
	);
	LUT2 #(
		.INIT('h2)
	) name4967 (
		\u5_mem_reg[1][13]/NET0131 ,
		_w7100_,
		_w7113_
	);
	LUT2 #(
		.INIT('h8)
	) name4968 (
		\u12_dout_reg[13]/P0001 ,
		_w7100_,
		_w7114_
	);
	LUT2 #(
		.INIT('h1)
	) name4969 (
		_w7113_,
		_w7114_,
		_w7115_
	);
	LUT2 #(
		.INIT('h2)
	) name4970 (
		\u5_mem_reg[1][14]/NET0131 ,
		_w7100_,
		_w7116_
	);
	LUT2 #(
		.INIT('h8)
	) name4971 (
		\u12_dout_reg[14]/P0001 ,
		_w7100_,
		_w7117_
	);
	LUT2 #(
		.INIT('h1)
	) name4972 (
		_w7116_,
		_w7117_,
		_w7118_
	);
	LUT2 #(
		.INIT('h2)
	) name4973 (
		\u5_mem_reg[1][15]/NET0131 ,
		_w7100_,
		_w7119_
	);
	LUT2 #(
		.INIT('h8)
	) name4974 (
		\u12_dout_reg[15]/P0001 ,
		_w7100_,
		_w7120_
	);
	LUT2 #(
		.INIT('h1)
	) name4975 (
		_w7119_,
		_w7120_,
		_w7121_
	);
	LUT2 #(
		.INIT('h2)
	) name4976 (
		\u5_mem_reg[1][16]/NET0131 ,
		_w7100_,
		_w7122_
	);
	LUT2 #(
		.INIT('h8)
	) name4977 (
		\u12_dout_reg[16]/P0001 ,
		_w7100_,
		_w7123_
	);
	LUT2 #(
		.INIT('h1)
	) name4978 (
		_w7122_,
		_w7123_,
		_w7124_
	);
	LUT2 #(
		.INIT('h2)
	) name4979 (
		\u5_mem_reg[1][17]/NET0131 ,
		_w7100_,
		_w7125_
	);
	LUT2 #(
		.INIT('h8)
	) name4980 (
		\u12_dout_reg[17]/P0001 ,
		_w7100_,
		_w7126_
	);
	LUT2 #(
		.INIT('h1)
	) name4981 (
		_w7125_,
		_w7126_,
		_w7127_
	);
	LUT2 #(
		.INIT('h2)
	) name4982 (
		\u5_mem_reg[1][18]/NET0131 ,
		_w7100_,
		_w7128_
	);
	LUT2 #(
		.INIT('h8)
	) name4983 (
		\u12_dout_reg[18]/P0001 ,
		_w7100_,
		_w7129_
	);
	LUT2 #(
		.INIT('h1)
	) name4984 (
		_w7128_,
		_w7129_,
		_w7130_
	);
	LUT2 #(
		.INIT('h2)
	) name4985 (
		\u5_mem_reg[1][19]/NET0131 ,
		_w7100_,
		_w7131_
	);
	LUT2 #(
		.INIT('h8)
	) name4986 (
		\u12_dout_reg[19]/P0001 ,
		_w7100_,
		_w7132_
	);
	LUT2 #(
		.INIT('h1)
	) name4987 (
		_w7131_,
		_w7132_,
		_w7133_
	);
	LUT2 #(
		.INIT('h2)
	) name4988 (
		\u5_mem_reg[1][1]/NET0131 ,
		_w7100_,
		_w7134_
	);
	LUT2 #(
		.INIT('h8)
	) name4989 (
		\u12_dout_reg[1]/P0001 ,
		_w7100_,
		_w7135_
	);
	LUT2 #(
		.INIT('h1)
	) name4990 (
		_w7134_,
		_w7135_,
		_w7136_
	);
	LUT2 #(
		.INIT('h2)
	) name4991 (
		\u5_mem_reg[1][20]/NET0131 ,
		_w7100_,
		_w7137_
	);
	LUT2 #(
		.INIT('h8)
	) name4992 (
		\u12_dout_reg[20]/P0001 ,
		_w7100_,
		_w7138_
	);
	LUT2 #(
		.INIT('h1)
	) name4993 (
		_w7137_,
		_w7138_,
		_w7139_
	);
	LUT2 #(
		.INIT('h2)
	) name4994 (
		\u5_mem_reg[1][21]/NET0131 ,
		_w7100_,
		_w7140_
	);
	LUT2 #(
		.INIT('h8)
	) name4995 (
		\u12_dout_reg[21]/P0001 ,
		_w7100_,
		_w7141_
	);
	LUT2 #(
		.INIT('h1)
	) name4996 (
		_w7140_,
		_w7141_,
		_w7142_
	);
	LUT2 #(
		.INIT('h2)
	) name4997 (
		\u5_mem_reg[1][22]/NET0131 ,
		_w7100_,
		_w7143_
	);
	LUT2 #(
		.INIT('h8)
	) name4998 (
		\u12_dout_reg[22]/P0001 ,
		_w7100_,
		_w7144_
	);
	LUT2 #(
		.INIT('h1)
	) name4999 (
		_w7143_,
		_w7144_,
		_w7145_
	);
	LUT2 #(
		.INIT('h2)
	) name5000 (
		\u5_mem_reg[1][23]/NET0131 ,
		_w7100_,
		_w7146_
	);
	LUT2 #(
		.INIT('h8)
	) name5001 (
		\u12_dout_reg[23]/P0001 ,
		_w7100_,
		_w7147_
	);
	LUT2 #(
		.INIT('h1)
	) name5002 (
		_w7146_,
		_w7147_,
		_w7148_
	);
	LUT2 #(
		.INIT('h2)
	) name5003 (
		\u5_mem_reg[1][24]/NET0131 ,
		_w7100_,
		_w7149_
	);
	LUT2 #(
		.INIT('h8)
	) name5004 (
		\u12_dout_reg[24]/P0001 ,
		_w7100_,
		_w7150_
	);
	LUT2 #(
		.INIT('h1)
	) name5005 (
		_w7149_,
		_w7150_,
		_w7151_
	);
	LUT2 #(
		.INIT('h2)
	) name5006 (
		\u5_mem_reg[1][25]/NET0131 ,
		_w7100_,
		_w7152_
	);
	LUT2 #(
		.INIT('h8)
	) name5007 (
		\u12_dout_reg[25]/P0001 ,
		_w7100_,
		_w7153_
	);
	LUT2 #(
		.INIT('h1)
	) name5008 (
		_w7152_,
		_w7153_,
		_w7154_
	);
	LUT2 #(
		.INIT('h2)
	) name5009 (
		\u5_mem_reg[1][26]/NET0131 ,
		_w7100_,
		_w7155_
	);
	LUT2 #(
		.INIT('h8)
	) name5010 (
		\u12_dout_reg[26]/P0001 ,
		_w7100_,
		_w7156_
	);
	LUT2 #(
		.INIT('h1)
	) name5011 (
		_w7155_,
		_w7156_,
		_w7157_
	);
	LUT2 #(
		.INIT('h2)
	) name5012 (
		\u5_mem_reg[1][27]/NET0131 ,
		_w7100_,
		_w7158_
	);
	LUT2 #(
		.INIT('h8)
	) name5013 (
		\u12_dout_reg[27]/P0001 ,
		_w7100_,
		_w7159_
	);
	LUT2 #(
		.INIT('h1)
	) name5014 (
		_w7158_,
		_w7159_,
		_w7160_
	);
	LUT2 #(
		.INIT('h2)
	) name5015 (
		\u5_mem_reg[1][28]/NET0131 ,
		_w7100_,
		_w7161_
	);
	LUT2 #(
		.INIT('h8)
	) name5016 (
		\u12_dout_reg[28]/P0001 ,
		_w7100_,
		_w7162_
	);
	LUT2 #(
		.INIT('h1)
	) name5017 (
		_w7161_,
		_w7162_,
		_w7163_
	);
	LUT2 #(
		.INIT('h2)
	) name5018 (
		\u5_mem_reg[1][29]/NET0131 ,
		_w7100_,
		_w7164_
	);
	LUT2 #(
		.INIT('h8)
	) name5019 (
		\u12_dout_reg[29]/P0001 ,
		_w7100_,
		_w7165_
	);
	LUT2 #(
		.INIT('h1)
	) name5020 (
		_w7164_,
		_w7165_,
		_w7166_
	);
	LUT2 #(
		.INIT('h2)
	) name5021 (
		\u5_mem_reg[1][2]/NET0131 ,
		_w7100_,
		_w7167_
	);
	LUT2 #(
		.INIT('h8)
	) name5022 (
		\u12_dout_reg[2]/P0001 ,
		_w7100_,
		_w7168_
	);
	LUT2 #(
		.INIT('h1)
	) name5023 (
		_w7167_,
		_w7168_,
		_w7169_
	);
	LUT2 #(
		.INIT('h2)
	) name5024 (
		\u5_mem_reg[1][30]/NET0131 ,
		_w7100_,
		_w7170_
	);
	LUT2 #(
		.INIT('h8)
	) name5025 (
		\u12_dout_reg[30]/P0001 ,
		_w7100_,
		_w7171_
	);
	LUT2 #(
		.INIT('h1)
	) name5026 (
		_w7170_,
		_w7171_,
		_w7172_
	);
	LUT2 #(
		.INIT('h2)
	) name5027 (
		\u5_mem_reg[1][31]/NET0131 ,
		_w7100_,
		_w7173_
	);
	LUT2 #(
		.INIT('h8)
	) name5028 (
		\u12_dout_reg[31]/P0001 ,
		_w7100_,
		_w7174_
	);
	LUT2 #(
		.INIT('h1)
	) name5029 (
		_w7173_,
		_w7174_,
		_w7175_
	);
	LUT2 #(
		.INIT('h2)
	) name5030 (
		\u5_mem_reg[1][3]/NET0131 ,
		_w7100_,
		_w7176_
	);
	LUT2 #(
		.INIT('h8)
	) name5031 (
		\u12_dout_reg[3]/P0001 ,
		_w7100_,
		_w7177_
	);
	LUT2 #(
		.INIT('h1)
	) name5032 (
		_w7176_,
		_w7177_,
		_w7178_
	);
	LUT2 #(
		.INIT('h2)
	) name5033 (
		\u5_mem_reg[1][4]/NET0131 ,
		_w7100_,
		_w7179_
	);
	LUT2 #(
		.INIT('h8)
	) name5034 (
		\u12_dout_reg[4]/P0001 ,
		_w7100_,
		_w7180_
	);
	LUT2 #(
		.INIT('h1)
	) name5035 (
		_w7179_,
		_w7180_,
		_w7181_
	);
	LUT2 #(
		.INIT('h2)
	) name5036 (
		\u5_mem_reg[1][5]/NET0131 ,
		_w7100_,
		_w7182_
	);
	LUT2 #(
		.INIT('h8)
	) name5037 (
		\u12_dout_reg[5]/P0001 ,
		_w7100_,
		_w7183_
	);
	LUT2 #(
		.INIT('h1)
	) name5038 (
		_w7182_,
		_w7183_,
		_w7184_
	);
	LUT2 #(
		.INIT('h2)
	) name5039 (
		\u5_mem_reg[1][6]/NET0131 ,
		_w7100_,
		_w7185_
	);
	LUT2 #(
		.INIT('h8)
	) name5040 (
		\u12_dout_reg[6]/P0001 ,
		_w7100_,
		_w7186_
	);
	LUT2 #(
		.INIT('h1)
	) name5041 (
		_w7185_,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h2)
	) name5042 (
		\u5_mem_reg[1][7]/NET0131 ,
		_w7100_,
		_w7188_
	);
	LUT2 #(
		.INIT('h8)
	) name5043 (
		\u12_dout_reg[7]/P0001 ,
		_w7100_,
		_w7189_
	);
	LUT2 #(
		.INIT('h1)
	) name5044 (
		_w7188_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h2)
	) name5045 (
		\u5_mem_reg[1][8]/NET0131 ,
		_w7100_,
		_w7191_
	);
	LUT2 #(
		.INIT('h8)
	) name5046 (
		\u12_dout_reg[8]/P0001 ,
		_w7100_,
		_w7192_
	);
	LUT2 #(
		.INIT('h1)
	) name5047 (
		_w7191_,
		_w7192_,
		_w7193_
	);
	LUT2 #(
		.INIT('h2)
	) name5048 (
		\u5_mem_reg[1][9]/NET0131 ,
		_w7100_,
		_w7194_
	);
	LUT2 #(
		.INIT('h8)
	) name5049 (
		\u12_dout_reg[9]/P0001 ,
		_w7100_,
		_w7195_
	);
	LUT2 #(
		.INIT('h1)
	) name5050 (
		_w7194_,
		_w7195_,
		_w7196_
	);
	LUT2 #(
		.INIT('h8)
	) name5051 (
		\u5_wp_reg[1]/NET0131 ,
		_w6415_,
		_w7197_
	);
	LUT2 #(
		.INIT('h2)
	) name5052 (
		\u5_mem_reg[2][0]/NET0131 ,
		_w7197_,
		_w7198_
	);
	LUT2 #(
		.INIT('h8)
	) name5053 (
		\u12_dout_reg[0]/P0001 ,
		_w7197_,
		_w7199_
	);
	LUT2 #(
		.INIT('h1)
	) name5054 (
		_w7198_,
		_w7199_,
		_w7200_
	);
	LUT2 #(
		.INIT('h2)
	) name5055 (
		\u5_mem_reg[2][10]/NET0131 ,
		_w7197_,
		_w7201_
	);
	LUT2 #(
		.INIT('h8)
	) name5056 (
		\u12_dout_reg[10]/P0001 ,
		_w7197_,
		_w7202_
	);
	LUT2 #(
		.INIT('h1)
	) name5057 (
		_w7201_,
		_w7202_,
		_w7203_
	);
	LUT2 #(
		.INIT('h2)
	) name5058 (
		\u5_mem_reg[2][11]/NET0131 ,
		_w7197_,
		_w7204_
	);
	LUT2 #(
		.INIT('h8)
	) name5059 (
		\u12_dout_reg[11]/P0001 ,
		_w7197_,
		_w7205_
	);
	LUT2 #(
		.INIT('h1)
	) name5060 (
		_w7204_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('h2)
	) name5061 (
		\u5_mem_reg[2][12]/NET0131 ,
		_w7197_,
		_w7207_
	);
	LUT2 #(
		.INIT('h8)
	) name5062 (
		\u12_dout_reg[12]/P0001 ,
		_w7197_,
		_w7208_
	);
	LUT2 #(
		.INIT('h1)
	) name5063 (
		_w7207_,
		_w7208_,
		_w7209_
	);
	LUT2 #(
		.INIT('h2)
	) name5064 (
		\u5_mem_reg[2][13]/NET0131 ,
		_w7197_,
		_w7210_
	);
	LUT2 #(
		.INIT('h8)
	) name5065 (
		\u12_dout_reg[13]/P0001 ,
		_w7197_,
		_w7211_
	);
	LUT2 #(
		.INIT('h1)
	) name5066 (
		_w7210_,
		_w7211_,
		_w7212_
	);
	LUT2 #(
		.INIT('h2)
	) name5067 (
		\u5_mem_reg[2][14]/NET0131 ,
		_w7197_,
		_w7213_
	);
	LUT2 #(
		.INIT('h8)
	) name5068 (
		\u12_dout_reg[14]/P0001 ,
		_w7197_,
		_w7214_
	);
	LUT2 #(
		.INIT('h1)
	) name5069 (
		_w7213_,
		_w7214_,
		_w7215_
	);
	LUT2 #(
		.INIT('h2)
	) name5070 (
		\u5_mem_reg[2][15]/NET0131 ,
		_w7197_,
		_w7216_
	);
	LUT2 #(
		.INIT('h8)
	) name5071 (
		\u12_dout_reg[15]/P0001 ,
		_w7197_,
		_w7217_
	);
	LUT2 #(
		.INIT('h1)
	) name5072 (
		_w7216_,
		_w7217_,
		_w7218_
	);
	LUT2 #(
		.INIT('h2)
	) name5073 (
		\u5_mem_reg[2][16]/NET0131 ,
		_w7197_,
		_w7219_
	);
	LUT2 #(
		.INIT('h8)
	) name5074 (
		\u12_dout_reg[16]/P0001 ,
		_w7197_,
		_w7220_
	);
	LUT2 #(
		.INIT('h1)
	) name5075 (
		_w7219_,
		_w7220_,
		_w7221_
	);
	LUT2 #(
		.INIT('h2)
	) name5076 (
		\u5_mem_reg[2][17]/NET0131 ,
		_w7197_,
		_w7222_
	);
	LUT2 #(
		.INIT('h8)
	) name5077 (
		\u12_dout_reg[17]/P0001 ,
		_w7197_,
		_w7223_
	);
	LUT2 #(
		.INIT('h1)
	) name5078 (
		_w7222_,
		_w7223_,
		_w7224_
	);
	LUT2 #(
		.INIT('h2)
	) name5079 (
		\u5_mem_reg[2][18]/NET0131 ,
		_w7197_,
		_w7225_
	);
	LUT2 #(
		.INIT('h8)
	) name5080 (
		\u12_dout_reg[18]/P0001 ,
		_w7197_,
		_w7226_
	);
	LUT2 #(
		.INIT('h1)
	) name5081 (
		_w7225_,
		_w7226_,
		_w7227_
	);
	LUT2 #(
		.INIT('h2)
	) name5082 (
		\u5_mem_reg[2][19]/NET0131 ,
		_w7197_,
		_w7228_
	);
	LUT2 #(
		.INIT('h8)
	) name5083 (
		\u12_dout_reg[19]/P0001 ,
		_w7197_,
		_w7229_
	);
	LUT2 #(
		.INIT('h1)
	) name5084 (
		_w7228_,
		_w7229_,
		_w7230_
	);
	LUT2 #(
		.INIT('h2)
	) name5085 (
		\u5_mem_reg[2][1]/NET0131 ,
		_w7197_,
		_w7231_
	);
	LUT2 #(
		.INIT('h8)
	) name5086 (
		\u12_dout_reg[1]/P0001 ,
		_w7197_,
		_w7232_
	);
	LUT2 #(
		.INIT('h1)
	) name5087 (
		_w7231_,
		_w7232_,
		_w7233_
	);
	LUT2 #(
		.INIT('h2)
	) name5088 (
		\u5_mem_reg[2][20]/NET0131 ,
		_w7197_,
		_w7234_
	);
	LUT2 #(
		.INIT('h8)
	) name5089 (
		\u12_dout_reg[20]/P0001 ,
		_w7197_,
		_w7235_
	);
	LUT2 #(
		.INIT('h1)
	) name5090 (
		_w7234_,
		_w7235_,
		_w7236_
	);
	LUT2 #(
		.INIT('h2)
	) name5091 (
		\u5_mem_reg[2][21]/NET0131 ,
		_w7197_,
		_w7237_
	);
	LUT2 #(
		.INIT('h8)
	) name5092 (
		\u12_dout_reg[21]/P0001 ,
		_w7197_,
		_w7238_
	);
	LUT2 #(
		.INIT('h1)
	) name5093 (
		_w7237_,
		_w7238_,
		_w7239_
	);
	LUT2 #(
		.INIT('h2)
	) name5094 (
		\u5_mem_reg[2][22]/NET0131 ,
		_w7197_,
		_w7240_
	);
	LUT2 #(
		.INIT('h8)
	) name5095 (
		\u12_dout_reg[22]/P0001 ,
		_w7197_,
		_w7241_
	);
	LUT2 #(
		.INIT('h1)
	) name5096 (
		_w7240_,
		_w7241_,
		_w7242_
	);
	LUT2 #(
		.INIT('h2)
	) name5097 (
		\u5_mem_reg[2][23]/NET0131 ,
		_w7197_,
		_w7243_
	);
	LUT2 #(
		.INIT('h8)
	) name5098 (
		\u12_dout_reg[23]/P0001 ,
		_w7197_,
		_w7244_
	);
	LUT2 #(
		.INIT('h1)
	) name5099 (
		_w7243_,
		_w7244_,
		_w7245_
	);
	LUT2 #(
		.INIT('h2)
	) name5100 (
		\u5_mem_reg[2][24]/NET0131 ,
		_w7197_,
		_w7246_
	);
	LUT2 #(
		.INIT('h8)
	) name5101 (
		\u12_dout_reg[24]/P0001 ,
		_w7197_,
		_w7247_
	);
	LUT2 #(
		.INIT('h1)
	) name5102 (
		_w7246_,
		_w7247_,
		_w7248_
	);
	LUT2 #(
		.INIT('h2)
	) name5103 (
		\u5_mem_reg[2][25]/NET0131 ,
		_w7197_,
		_w7249_
	);
	LUT2 #(
		.INIT('h8)
	) name5104 (
		\u12_dout_reg[25]/P0001 ,
		_w7197_,
		_w7250_
	);
	LUT2 #(
		.INIT('h1)
	) name5105 (
		_w7249_,
		_w7250_,
		_w7251_
	);
	LUT2 #(
		.INIT('h2)
	) name5106 (
		\u5_mem_reg[2][26]/NET0131 ,
		_w7197_,
		_w7252_
	);
	LUT2 #(
		.INIT('h8)
	) name5107 (
		\u12_dout_reg[26]/P0001 ,
		_w7197_,
		_w7253_
	);
	LUT2 #(
		.INIT('h1)
	) name5108 (
		_w7252_,
		_w7253_,
		_w7254_
	);
	LUT2 #(
		.INIT('h2)
	) name5109 (
		\u5_mem_reg[2][27]/NET0131 ,
		_w7197_,
		_w7255_
	);
	LUT2 #(
		.INIT('h8)
	) name5110 (
		\u12_dout_reg[27]/P0001 ,
		_w7197_,
		_w7256_
	);
	LUT2 #(
		.INIT('h1)
	) name5111 (
		_w7255_,
		_w7256_,
		_w7257_
	);
	LUT2 #(
		.INIT('h2)
	) name5112 (
		\u5_mem_reg[2][28]/NET0131 ,
		_w7197_,
		_w7258_
	);
	LUT2 #(
		.INIT('h8)
	) name5113 (
		\u12_dout_reg[28]/P0001 ,
		_w7197_,
		_w7259_
	);
	LUT2 #(
		.INIT('h1)
	) name5114 (
		_w7258_,
		_w7259_,
		_w7260_
	);
	LUT2 #(
		.INIT('h2)
	) name5115 (
		\u5_mem_reg[2][29]/NET0131 ,
		_w7197_,
		_w7261_
	);
	LUT2 #(
		.INIT('h8)
	) name5116 (
		\u12_dout_reg[29]/P0001 ,
		_w7197_,
		_w7262_
	);
	LUT2 #(
		.INIT('h1)
	) name5117 (
		_w7261_,
		_w7262_,
		_w7263_
	);
	LUT2 #(
		.INIT('h2)
	) name5118 (
		\u5_mem_reg[2][2]/NET0131 ,
		_w7197_,
		_w7264_
	);
	LUT2 #(
		.INIT('h8)
	) name5119 (
		\u12_dout_reg[2]/P0001 ,
		_w7197_,
		_w7265_
	);
	LUT2 #(
		.INIT('h1)
	) name5120 (
		_w7264_,
		_w7265_,
		_w7266_
	);
	LUT2 #(
		.INIT('h2)
	) name5121 (
		\u5_mem_reg[2][30]/NET0131 ,
		_w7197_,
		_w7267_
	);
	LUT2 #(
		.INIT('h8)
	) name5122 (
		\u12_dout_reg[30]/P0001 ,
		_w7197_,
		_w7268_
	);
	LUT2 #(
		.INIT('h1)
	) name5123 (
		_w7267_,
		_w7268_,
		_w7269_
	);
	LUT2 #(
		.INIT('h2)
	) name5124 (
		\u5_mem_reg[2][31]/NET0131 ,
		_w7197_,
		_w7270_
	);
	LUT2 #(
		.INIT('h8)
	) name5125 (
		\u12_dout_reg[31]/P0001 ,
		_w7197_,
		_w7271_
	);
	LUT2 #(
		.INIT('h1)
	) name5126 (
		_w7270_,
		_w7271_,
		_w7272_
	);
	LUT2 #(
		.INIT('h2)
	) name5127 (
		\u5_mem_reg[2][3]/NET0131 ,
		_w7197_,
		_w7273_
	);
	LUT2 #(
		.INIT('h8)
	) name5128 (
		\u12_dout_reg[3]/P0001 ,
		_w7197_,
		_w7274_
	);
	LUT2 #(
		.INIT('h1)
	) name5129 (
		_w7273_,
		_w7274_,
		_w7275_
	);
	LUT2 #(
		.INIT('h2)
	) name5130 (
		\u5_mem_reg[2][4]/NET0131 ,
		_w7197_,
		_w7276_
	);
	LUT2 #(
		.INIT('h8)
	) name5131 (
		\u12_dout_reg[4]/P0001 ,
		_w7197_,
		_w7277_
	);
	LUT2 #(
		.INIT('h1)
	) name5132 (
		_w7276_,
		_w7277_,
		_w7278_
	);
	LUT2 #(
		.INIT('h2)
	) name5133 (
		\u5_mem_reg[2][5]/NET0131 ,
		_w7197_,
		_w7279_
	);
	LUT2 #(
		.INIT('h8)
	) name5134 (
		\u12_dout_reg[5]/P0001 ,
		_w7197_,
		_w7280_
	);
	LUT2 #(
		.INIT('h1)
	) name5135 (
		_w7279_,
		_w7280_,
		_w7281_
	);
	LUT2 #(
		.INIT('h2)
	) name5136 (
		\u5_mem_reg[2][6]/NET0131 ,
		_w7197_,
		_w7282_
	);
	LUT2 #(
		.INIT('h8)
	) name5137 (
		\u12_dout_reg[6]/P0001 ,
		_w7197_,
		_w7283_
	);
	LUT2 #(
		.INIT('h1)
	) name5138 (
		_w7282_,
		_w7283_,
		_w7284_
	);
	LUT2 #(
		.INIT('h2)
	) name5139 (
		\u5_mem_reg[2][7]/NET0131 ,
		_w7197_,
		_w7285_
	);
	LUT2 #(
		.INIT('h8)
	) name5140 (
		\u12_dout_reg[7]/P0001 ,
		_w7197_,
		_w7286_
	);
	LUT2 #(
		.INIT('h1)
	) name5141 (
		_w7285_,
		_w7286_,
		_w7287_
	);
	LUT2 #(
		.INIT('h2)
	) name5142 (
		\u5_mem_reg[2][8]/NET0131 ,
		_w7197_,
		_w7288_
	);
	LUT2 #(
		.INIT('h8)
	) name5143 (
		\u12_dout_reg[8]/P0001 ,
		_w7197_,
		_w7289_
	);
	LUT2 #(
		.INIT('h1)
	) name5144 (
		_w7288_,
		_w7289_,
		_w7290_
	);
	LUT2 #(
		.INIT('h2)
	) name5145 (
		\u5_mem_reg[2][9]/NET0131 ,
		_w7197_,
		_w7291_
	);
	LUT2 #(
		.INIT('h8)
	) name5146 (
		\u12_dout_reg[9]/P0001 ,
		_w7197_,
		_w7292_
	);
	LUT2 #(
		.INIT('h1)
	) name5147 (
		_w7291_,
		_w7292_,
		_w7293_
	);
	LUT2 #(
		.INIT('h2)
	) name5148 (
		\u5_mem_reg[3][0]/NET0131 ,
		_w6313_,
		_w7294_
	);
	LUT2 #(
		.INIT('h8)
	) name5149 (
		\u12_dout_reg[0]/P0001 ,
		_w6313_,
		_w7295_
	);
	LUT2 #(
		.INIT('h1)
	) name5150 (
		_w7294_,
		_w7295_,
		_w7296_
	);
	LUT2 #(
		.INIT('h2)
	) name5151 (
		\u5_mem_reg[3][10]/NET0131 ,
		_w6313_,
		_w7297_
	);
	LUT2 #(
		.INIT('h8)
	) name5152 (
		\u12_dout_reg[10]/P0001 ,
		_w6313_,
		_w7298_
	);
	LUT2 #(
		.INIT('h1)
	) name5153 (
		_w7297_,
		_w7298_,
		_w7299_
	);
	LUT2 #(
		.INIT('h2)
	) name5154 (
		\u5_mem_reg[3][11]/NET0131 ,
		_w6313_,
		_w7300_
	);
	LUT2 #(
		.INIT('h8)
	) name5155 (
		\u12_dout_reg[11]/P0001 ,
		_w6313_,
		_w7301_
	);
	LUT2 #(
		.INIT('h1)
	) name5156 (
		_w7300_,
		_w7301_,
		_w7302_
	);
	LUT2 #(
		.INIT('h2)
	) name5157 (
		\u5_mem_reg[3][12]/NET0131 ,
		_w6313_,
		_w7303_
	);
	LUT2 #(
		.INIT('h8)
	) name5158 (
		\u12_dout_reg[12]/P0001 ,
		_w6313_,
		_w7304_
	);
	LUT2 #(
		.INIT('h1)
	) name5159 (
		_w7303_,
		_w7304_,
		_w7305_
	);
	LUT2 #(
		.INIT('h2)
	) name5160 (
		\u5_mem_reg[3][13]/NET0131 ,
		_w6313_,
		_w7306_
	);
	LUT2 #(
		.INIT('h8)
	) name5161 (
		\u12_dout_reg[13]/P0001 ,
		_w6313_,
		_w7307_
	);
	LUT2 #(
		.INIT('h1)
	) name5162 (
		_w7306_,
		_w7307_,
		_w7308_
	);
	LUT2 #(
		.INIT('h2)
	) name5163 (
		\u5_mem_reg[3][14]/NET0131 ,
		_w6313_,
		_w7309_
	);
	LUT2 #(
		.INIT('h8)
	) name5164 (
		\u12_dout_reg[14]/P0001 ,
		_w6313_,
		_w7310_
	);
	LUT2 #(
		.INIT('h1)
	) name5165 (
		_w7309_,
		_w7310_,
		_w7311_
	);
	LUT2 #(
		.INIT('h2)
	) name5166 (
		\u5_mem_reg[3][15]/NET0131 ,
		_w6313_,
		_w7312_
	);
	LUT2 #(
		.INIT('h8)
	) name5167 (
		\u12_dout_reg[15]/P0001 ,
		_w6313_,
		_w7313_
	);
	LUT2 #(
		.INIT('h1)
	) name5168 (
		_w7312_,
		_w7313_,
		_w7314_
	);
	LUT2 #(
		.INIT('h2)
	) name5169 (
		\u5_mem_reg[3][16]/NET0131 ,
		_w6313_,
		_w7315_
	);
	LUT2 #(
		.INIT('h8)
	) name5170 (
		\u12_dout_reg[16]/P0001 ,
		_w6313_,
		_w7316_
	);
	LUT2 #(
		.INIT('h1)
	) name5171 (
		_w7315_,
		_w7316_,
		_w7317_
	);
	LUT2 #(
		.INIT('h2)
	) name5172 (
		\u5_mem_reg[3][17]/NET0131 ,
		_w6313_,
		_w7318_
	);
	LUT2 #(
		.INIT('h8)
	) name5173 (
		\u12_dout_reg[17]/P0001 ,
		_w6313_,
		_w7319_
	);
	LUT2 #(
		.INIT('h1)
	) name5174 (
		_w7318_,
		_w7319_,
		_w7320_
	);
	LUT2 #(
		.INIT('h2)
	) name5175 (
		\u5_mem_reg[3][18]/NET0131 ,
		_w6313_,
		_w7321_
	);
	LUT2 #(
		.INIT('h8)
	) name5176 (
		\u12_dout_reg[18]/P0001 ,
		_w6313_,
		_w7322_
	);
	LUT2 #(
		.INIT('h1)
	) name5177 (
		_w7321_,
		_w7322_,
		_w7323_
	);
	LUT2 #(
		.INIT('h2)
	) name5178 (
		\u5_mem_reg[3][19]/NET0131 ,
		_w6313_,
		_w7324_
	);
	LUT2 #(
		.INIT('h8)
	) name5179 (
		\u12_dout_reg[19]/P0001 ,
		_w6313_,
		_w7325_
	);
	LUT2 #(
		.INIT('h1)
	) name5180 (
		_w7324_,
		_w7325_,
		_w7326_
	);
	LUT2 #(
		.INIT('h2)
	) name5181 (
		\u5_mem_reg[3][1]/NET0131 ,
		_w6313_,
		_w7327_
	);
	LUT2 #(
		.INIT('h8)
	) name5182 (
		\u12_dout_reg[1]/P0001 ,
		_w6313_,
		_w7328_
	);
	LUT2 #(
		.INIT('h1)
	) name5183 (
		_w7327_,
		_w7328_,
		_w7329_
	);
	LUT2 #(
		.INIT('h2)
	) name5184 (
		\u5_mem_reg[3][20]/NET0131 ,
		_w6313_,
		_w7330_
	);
	LUT2 #(
		.INIT('h8)
	) name5185 (
		\u12_dout_reg[20]/P0001 ,
		_w6313_,
		_w7331_
	);
	LUT2 #(
		.INIT('h1)
	) name5186 (
		_w7330_,
		_w7331_,
		_w7332_
	);
	LUT2 #(
		.INIT('h2)
	) name5187 (
		\u5_mem_reg[3][21]/NET0131 ,
		_w6313_,
		_w7333_
	);
	LUT2 #(
		.INIT('h8)
	) name5188 (
		\u12_dout_reg[21]/P0001 ,
		_w6313_,
		_w7334_
	);
	LUT2 #(
		.INIT('h1)
	) name5189 (
		_w7333_,
		_w7334_,
		_w7335_
	);
	LUT2 #(
		.INIT('h2)
	) name5190 (
		\u5_mem_reg[3][22]/NET0131 ,
		_w6313_,
		_w7336_
	);
	LUT2 #(
		.INIT('h8)
	) name5191 (
		\u12_dout_reg[22]/P0001 ,
		_w6313_,
		_w7337_
	);
	LUT2 #(
		.INIT('h1)
	) name5192 (
		_w7336_,
		_w7337_,
		_w7338_
	);
	LUT2 #(
		.INIT('h2)
	) name5193 (
		\u5_mem_reg[3][23]/NET0131 ,
		_w6313_,
		_w7339_
	);
	LUT2 #(
		.INIT('h8)
	) name5194 (
		\u12_dout_reg[23]/P0001 ,
		_w6313_,
		_w7340_
	);
	LUT2 #(
		.INIT('h1)
	) name5195 (
		_w7339_,
		_w7340_,
		_w7341_
	);
	LUT2 #(
		.INIT('h2)
	) name5196 (
		\u5_mem_reg[3][24]/NET0131 ,
		_w6313_,
		_w7342_
	);
	LUT2 #(
		.INIT('h8)
	) name5197 (
		\u12_dout_reg[24]/P0001 ,
		_w6313_,
		_w7343_
	);
	LUT2 #(
		.INIT('h1)
	) name5198 (
		_w7342_,
		_w7343_,
		_w7344_
	);
	LUT2 #(
		.INIT('h2)
	) name5199 (
		\u5_mem_reg[3][25]/NET0131 ,
		_w6313_,
		_w7345_
	);
	LUT2 #(
		.INIT('h8)
	) name5200 (
		\u12_dout_reg[25]/P0001 ,
		_w6313_,
		_w7346_
	);
	LUT2 #(
		.INIT('h1)
	) name5201 (
		_w7345_,
		_w7346_,
		_w7347_
	);
	LUT2 #(
		.INIT('h2)
	) name5202 (
		\u5_mem_reg[3][26]/NET0131 ,
		_w6313_,
		_w7348_
	);
	LUT2 #(
		.INIT('h8)
	) name5203 (
		\u12_dout_reg[26]/P0001 ,
		_w6313_,
		_w7349_
	);
	LUT2 #(
		.INIT('h1)
	) name5204 (
		_w7348_,
		_w7349_,
		_w7350_
	);
	LUT2 #(
		.INIT('h2)
	) name5205 (
		\u5_mem_reg[3][27]/NET0131 ,
		_w6313_,
		_w7351_
	);
	LUT2 #(
		.INIT('h8)
	) name5206 (
		\u12_dout_reg[27]/P0001 ,
		_w6313_,
		_w7352_
	);
	LUT2 #(
		.INIT('h1)
	) name5207 (
		_w7351_,
		_w7352_,
		_w7353_
	);
	LUT2 #(
		.INIT('h2)
	) name5208 (
		\u5_mem_reg[3][28]/NET0131 ,
		_w6313_,
		_w7354_
	);
	LUT2 #(
		.INIT('h8)
	) name5209 (
		\u12_dout_reg[28]/P0001 ,
		_w6313_,
		_w7355_
	);
	LUT2 #(
		.INIT('h1)
	) name5210 (
		_w7354_,
		_w7355_,
		_w7356_
	);
	LUT2 #(
		.INIT('h2)
	) name5211 (
		\u5_mem_reg[3][29]/NET0131 ,
		_w6313_,
		_w7357_
	);
	LUT2 #(
		.INIT('h8)
	) name5212 (
		\u12_dout_reg[29]/P0001 ,
		_w6313_,
		_w7358_
	);
	LUT2 #(
		.INIT('h1)
	) name5213 (
		_w7357_,
		_w7358_,
		_w7359_
	);
	LUT2 #(
		.INIT('h2)
	) name5214 (
		\u5_mem_reg[3][2]/NET0131 ,
		_w6313_,
		_w7360_
	);
	LUT2 #(
		.INIT('h8)
	) name5215 (
		\u12_dout_reg[2]/P0001 ,
		_w6313_,
		_w7361_
	);
	LUT2 #(
		.INIT('h1)
	) name5216 (
		_w7360_,
		_w7361_,
		_w7362_
	);
	LUT2 #(
		.INIT('h2)
	) name5217 (
		\u5_mem_reg[3][30]/NET0131 ,
		_w6313_,
		_w7363_
	);
	LUT2 #(
		.INIT('h8)
	) name5218 (
		\u12_dout_reg[30]/P0001 ,
		_w6313_,
		_w7364_
	);
	LUT2 #(
		.INIT('h1)
	) name5219 (
		_w7363_,
		_w7364_,
		_w7365_
	);
	LUT2 #(
		.INIT('h2)
	) name5220 (
		\u5_mem_reg[3][31]/NET0131 ,
		_w6313_,
		_w7366_
	);
	LUT2 #(
		.INIT('h8)
	) name5221 (
		\u12_dout_reg[31]/P0001 ,
		_w6313_,
		_w7367_
	);
	LUT2 #(
		.INIT('h1)
	) name5222 (
		_w7366_,
		_w7367_,
		_w7368_
	);
	LUT2 #(
		.INIT('h2)
	) name5223 (
		\u5_mem_reg[3][3]/NET0131 ,
		_w6313_,
		_w7369_
	);
	LUT2 #(
		.INIT('h8)
	) name5224 (
		\u12_dout_reg[3]/P0001 ,
		_w6313_,
		_w7370_
	);
	LUT2 #(
		.INIT('h1)
	) name5225 (
		_w7369_,
		_w7370_,
		_w7371_
	);
	LUT2 #(
		.INIT('h2)
	) name5226 (
		\u5_mem_reg[3][4]/NET0131 ,
		_w6313_,
		_w7372_
	);
	LUT2 #(
		.INIT('h8)
	) name5227 (
		\u12_dout_reg[4]/P0001 ,
		_w6313_,
		_w7373_
	);
	LUT2 #(
		.INIT('h1)
	) name5228 (
		_w7372_,
		_w7373_,
		_w7374_
	);
	LUT2 #(
		.INIT('h2)
	) name5229 (
		\u5_mem_reg[3][5]/NET0131 ,
		_w6313_,
		_w7375_
	);
	LUT2 #(
		.INIT('h8)
	) name5230 (
		\u12_dout_reg[5]/P0001 ,
		_w6313_,
		_w7376_
	);
	LUT2 #(
		.INIT('h1)
	) name5231 (
		_w7375_,
		_w7376_,
		_w7377_
	);
	LUT2 #(
		.INIT('h2)
	) name5232 (
		\u5_mem_reg[3][6]/NET0131 ,
		_w6313_,
		_w7378_
	);
	LUT2 #(
		.INIT('h8)
	) name5233 (
		\u12_dout_reg[6]/P0001 ,
		_w6313_,
		_w7379_
	);
	LUT2 #(
		.INIT('h1)
	) name5234 (
		_w7378_,
		_w7379_,
		_w7380_
	);
	LUT2 #(
		.INIT('h2)
	) name5235 (
		\u5_mem_reg[3][7]/NET0131 ,
		_w6313_,
		_w7381_
	);
	LUT2 #(
		.INIT('h8)
	) name5236 (
		\u12_dout_reg[7]/P0001 ,
		_w6313_,
		_w7382_
	);
	LUT2 #(
		.INIT('h1)
	) name5237 (
		_w7381_,
		_w7382_,
		_w7383_
	);
	LUT2 #(
		.INIT('h2)
	) name5238 (
		\u5_mem_reg[3][8]/NET0131 ,
		_w6313_,
		_w7384_
	);
	LUT2 #(
		.INIT('h8)
	) name5239 (
		\u12_dout_reg[8]/P0001 ,
		_w6313_,
		_w7385_
	);
	LUT2 #(
		.INIT('h1)
	) name5240 (
		_w7384_,
		_w7385_,
		_w7386_
	);
	LUT2 #(
		.INIT('h2)
	) name5241 (
		\u5_mem_reg[3][9]/NET0131 ,
		_w6313_,
		_w7387_
	);
	LUT2 #(
		.INIT('h8)
	) name5242 (
		\u12_dout_reg[9]/P0001 ,
		_w6313_,
		_w7388_
	);
	LUT2 #(
		.INIT('h1)
	) name5243 (
		_w7387_,
		_w7388_,
		_w7389_
	);
	LUT2 #(
		.INIT('h2)
	) name5244 (
		\u8_mem_reg[3][6]/NET0131 ,
		_w6301_,
		_w7390_
	);
	LUT2 #(
		.INIT('h8)
	) name5245 (
		\u12_dout_reg[6]/P0001 ,
		_w6301_,
		_w7391_
	);
	LUT2 #(
		.INIT('h1)
	) name5246 (
		_w7390_,
		_w7391_,
		_w7392_
	);
	LUT2 #(
		.INIT('h2)
	) name5247 (
		\u8_mem_reg[1][28]/NET0131 ,
		_w6629_,
		_w7393_
	);
	LUT2 #(
		.INIT('h8)
	) name5248 (
		\u12_dout_reg[28]/P0001 ,
		_w6629_,
		_w7394_
	);
	LUT2 #(
		.INIT('h1)
	) name5249 (
		_w7393_,
		_w7394_,
		_w7395_
	);
	LUT2 #(
		.INIT('h2)
	) name5250 (
		\u3_mem_reg[2][20]/NET0131 ,
		_w6583_,
		_w7396_
	);
	LUT2 #(
		.INIT('h8)
	) name5251 (
		\u12_dout_reg[20]/P0001 ,
		_w6583_,
		_w7397_
	);
	LUT2 #(
		.INIT('h1)
	) name5252 (
		_w7396_,
		_w7397_,
		_w7398_
	);
	LUT2 #(
		.INIT('h2)
	) name5253 (
		\u8_mem_reg[3][31]/NET0131 ,
		_w6301_,
		_w7399_
	);
	LUT2 #(
		.INIT('h8)
	) name5254 (
		\u12_dout_reg[31]/P0001 ,
		_w6301_,
		_w7400_
	);
	LUT2 #(
		.INIT('h1)
	) name5255 (
		_w7399_,
		_w7400_,
		_w7401_
	);
	LUT2 #(
		.INIT('h4)
	) name5256 (
		\u6_wp_reg[1]/NET0131 ,
		_w6324_,
		_w7402_
	);
	LUT2 #(
		.INIT('h2)
	) name5257 (
		\u6_mem_reg[1][0]/NET0131 ,
		_w7402_,
		_w7403_
	);
	LUT2 #(
		.INIT('h8)
	) name5258 (
		\u12_dout_reg[0]/P0001 ,
		_w7402_,
		_w7404_
	);
	LUT2 #(
		.INIT('h1)
	) name5259 (
		_w7403_,
		_w7404_,
		_w7405_
	);
	LUT2 #(
		.INIT('h2)
	) name5260 (
		\u6_mem_reg[1][10]/NET0131 ,
		_w7402_,
		_w7406_
	);
	LUT2 #(
		.INIT('h8)
	) name5261 (
		\u12_dout_reg[10]/P0001 ,
		_w7402_,
		_w7407_
	);
	LUT2 #(
		.INIT('h1)
	) name5262 (
		_w7406_,
		_w7407_,
		_w7408_
	);
	LUT2 #(
		.INIT('h2)
	) name5263 (
		\u6_mem_reg[1][11]/NET0131 ,
		_w7402_,
		_w7409_
	);
	LUT2 #(
		.INIT('h8)
	) name5264 (
		\u12_dout_reg[11]/P0001 ,
		_w7402_,
		_w7410_
	);
	LUT2 #(
		.INIT('h1)
	) name5265 (
		_w7409_,
		_w7410_,
		_w7411_
	);
	LUT2 #(
		.INIT('h2)
	) name5266 (
		\u6_mem_reg[1][12]/NET0131 ,
		_w7402_,
		_w7412_
	);
	LUT2 #(
		.INIT('h8)
	) name5267 (
		\u12_dout_reg[12]/P0001 ,
		_w7402_,
		_w7413_
	);
	LUT2 #(
		.INIT('h1)
	) name5268 (
		_w7412_,
		_w7413_,
		_w7414_
	);
	LUT2 #(
		.INIT('h2)
	) name5269 (
		\u6_mem_reg[1][13]/NET0131 ,
		_w7402_,
		_w7415_
	);
	LUT2 #(
		.INIT('h8)
	) name5270 (
		\u12_dout_reg[13]/P0001 ,
		_w7402_,
		_w7416_
	);
	LUT2 #(
		.INIT('h1)
	) name5271 (
		_w7415_,
		_w7416_,
		_w7417_
	);
	LUT2 #(
		.INIT('h2)
	) name5272 (
		\u6_mem_reg[1][14]/NET0131 ,
		_w7402_,
		_w7418_
	);
	LUT2 #(
		.INIT('h8)
	) name5273 (
		\u12_dout_reg[14]/P0001 ,
		_w7402_,
		_w7419_
	);
	LUT2 #(
		.INIT('h1)
	) name5274 (
		_w7418_,
		_w7419_,
		_w7420_
	);
	LUT2 #(
		.INIT('h2)
	) name5275 (
		\u6_mem_reg[1][15]/NET0131 ,
		_w7402_,
		_w7421_
	);
	LUT2 #(
		.INIT('h8)
	) name5276 (
		\u12_dout_reg[15]/P0001 ,
		_w7402_,
		_w7422_
	);
	LUT2 #(
		.INIT('h1)
	) name5277 (
		_w7421_,
		_w7422_,
		_w7423_
	);
	LUT2 #(
		.INIT('h2)
	) name5278 (
		\u6_mem_reg[1][16]/NET0131 ,
		_w7402_,
		_w7424_
	);
	LUT2 #(
		.INIT('h8)
	) name5279 (
		\u12_dout_reg[16]/P0001 ,
		_w7402_,
		_w7425_
	);
	LUT2 #(
		.INIT('h1)
	) name5280 (
		_w7424_,
		_w7425_,
		_w7426_
	);
	LUT2 #(
		.INIT('h2)
	) name5281 (
		\u6_mem_reg[1][17]/NET0131 ,
		_w7402_,
		_w7427_
	);
	LUT2 #(
		.INIT('h8)
	) name5282 (
		\u12_dout_reg[17]/P0001 ,
		_w7402_,
		_w7428_
	);
	LUT2 #(
		.INIT('h1)
	) name5283 (
		_w7427_,
		_w7428_,
		_w7429_
	);
	LUT2 #(
		.INIT('h2)
	) name5284 (
		\u6_mem_reg[1][18]/NET0131 ,
		_w7402_,
		_w7430_
	);
	LUT2 #(
		.INIT('h8)
	) name5285 (
		\u12_dout_reg[18]/P0001 ,
		_w7402_,
		_w7431_
	);
	LUT2 #(
		.INIT('h1)
	) name5286 (
		_w7430_,
		_w7431_,
		_w7432_
	);
	LUT2 #(
		.INIT('h2)
	) name5287 (
		\u6_mem_reg[1][19]/NET0131 ,
		_w7402_,
		_w7433_
	);
	LUT2 #(
		.INIT('h8)
	) name5288 (
		\u12_dout_reg[19]/P0001 ,
		_w7402_,
		_w7434_
	);
	LUT2 #(
		.INIT('h1)
	) name5289 (
		_w7433_,
		_w7434_,
		_w7435_
	);
	LUT2 #(
		.INIT('h2)
	) name5290 (
		\u6_mem_reg[1][1]/NET0131 ,
		_w7402_,
		_w7436_
	);
	LUT2 #(
		.INIT('h8)
	) name5291 (
		\u12_dout_reg[1]/P0001 ,
		_w7402_,
		_w7437_
	);
	LUT2 #(
		.INIT('h1)
	) name5292 (
		_w7436_,
		_w7437_,
		_w7438_
	);
	LUT2 #(
		.INIT('h2)
	) name5293 (
		\u6_mem_reg[1][20]/NET0131 ,
		_w7402_,
		_w7439_
	);
	LUT2 #(
		.INIT('h8)
	) name5294 (
		\u12_dout_reg[20]/P0001 ,
		_w7402_,
		_w7440_
	);
	LUT2 #(
		.INIT('h1)
	) name5295 (
		_w7439_,
		_w7440_,
		_w7441_
	);
	LUT2 #(
		.INIT('h2)
	) name5296 (
		\u6_mem_reg[1][21]/NET0131 ,
		_w7402_,
		_w7442_
	);
	LUT2 #(
		.INIT('h8)
	) name5297 (
		\u12_dout_reg[21]/P0001 ,
		_w7402_,
		_w7443_
	);
	LUT2 #(
		.INIT('h1)
	) name5298 (
		_w7442_,
		_w7443_,
		_w7444_
	);
	LUT2 #(
		.INIT('h2)
	) name5299 (
		\u6_mem_reg[1][22]/NET0131 ,
		_w7402_,
		_w7445_
	);
	LUT2 #(
		.INIT('h8)
	) name5300 (
		\u12_dout_reg[22]/P0001 ,
		_w7402_,
		_w7446_
	);
	LUT2 #(
		.INIT('h1)
	) name5301 (
		_w7445_,
		_w7446_,
		_w7447_
	);
	LUT2 #(
		.INIT('h2)
	) name5302 (
		\u6_mem_reg[1][23]/NET0131 ,
		_w7402_,
		_w7448_
	);
	LUT2 #(
		.INIT('h8)
	) name5303 (
		\u12_dout_reg[23]/P0001 ,
		_w7402_,
		_w7449_
	);
	LUT2 #(
		.INIT('h1)
	) name5304 (
		_w7448_,
		_w7449_,
		_w7450_
	);
	LUT2 #(
		.INIT('h2)
	) name5305 (
		\u6_mem_reg[1][24]/NET0131 ,
		_w7402_,
		_w7451_
	);
	LUT2 #(
		.INIT('h8)
	) name5306 (
		\u12_dout_reg[24]/P0001 ,
		_w7402_,
		_w7452_
	);
	LUT2 #(
		.INIT('h1)
	) name5307 (
		_w7451_,
		_w7452_,
		_w7453_
	);
	LUT2 #(
		.INIT('h2)
	) name5308 (
		\u6_mem_reg[1][25]/NET0131 ,
		_w7402_,
		_w7454_
	);
	LUT2 #(
		.INIT('h8)
	) name5309 (
		\u12_dout_reg[25]/P0001 ,
		_w7402_,
		_w7455_
	);
	LUT2 #(
		.INIT('h1)
	) name5310 (
		_w7454_,
		_w7455_,
		_w7456_
	);
	LUT2 #(
		.INIT('h2)
	) name5311 (
		\u6_mem_reg[1][26]/NET0131 ,
		_w7402_,
		_w7457_
	);
	LUT2 #(
		.INIT('h8)
	) name5312 (
		\u12_dout_reg[26]/P0001 ,
		_w7402_,
		_w7458_
	);
	LUT2 #(
		.INIT('h1)
	) name5313 (
		_w7457_,
		_w7458_,
		_w7459_
	);
	LUT2 #(
		.INIT('h2)
	) name5314 (
		\u6_mem_reg[1][27]/NET0131 ,
		_w7402_,
		_w7460_
	);
	LUT2 #(
		.INIT('h8)
	) name5315 (
		\u12_dout_reg[27]/P0001 ,
		_w7402_,
		_w7461_
	);
	LUT2 #(
		.INIT('h1)
	) name5316 (
		_w7460_,
		_w7461_,
		_w7462_
	);
	LUT2 #(
		.INIT('h2)
	) name5317 (
		\u6_mem_reg[1][28]/NET0131 ,
		_w7402_,
		_w7463_
	);
	LUT2 #(
		.INIT('h8)
	) name5318 (
		\u12_dout_reg[28]/P0001 ,
		_w7402_,
		_w7464_
	);
	LUT2 #(
		.INIT('h1)
	) name5319 (
		_w7463_,
		_w7464_,
		_w7465_
	);
	LUT2 #(
		.INIT('h2)
	) name5320 (
		\u6_mem_reg[1][29]/NET0131 ,
		_w7402_,
		_w7466_
	);
	LUT2 #(
		.INIT('h8)
	) name5321 (
		\u12_dout_reg[29]/P0001 ,
		_w7402_,
		_w7467_
	);
	LUT2 #(
		.INIT('h1)
	) name5322 (
		_w7466_,
		_w7467_,
		_w7468_
	);
	LUT2 #(
		.INIT('h2)
	) name5323 (
		\u6_mem_reg[1][2]/NET0131 ,
		_w7402_,
		_w7469_
	);
	LUT2 #(
		.INIT('h8)
	) name5324 (
		\u12_dout_reg[2]/P0001 ,
		_w7402_,
		_w7470_
	);
	LUT2 #(
		.INIT('h1)
	) name5325 (
		_w7469_,
		_w7470_,
		_w7471_
	);
	LUT2 #(
		.INIT('h2)
	) name5326 (
		\u6_mem_reg[1][30]/NET0131 ,
		_w7402_,
		_w7472_
	);
	LUT2 #(
		.INIT('h8)
	) name5327 (
		\u12_dout_reg[30]/P0001 ,
		_w7402_,
		_w7473_
	);
	LUT2 #(
		.INIT('h1)
	) name5328 (
		_w7472_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h2)
	) name5329 (
		\u6_mem_reg[1][31]/NET0131 ,
		_w7402_,
		_w7475_
	);
	LUT2 #(
		.INIT('h8)
	) name5330 (
		\u12_dout_reg[31]/P0001 ,
		_w7402_,
		_w7476_
	);
	LUT2 #(
		.INIT('h1)
	) name5331 (
		_w7475_,
		_w7476_,
		_w7477_
	);
	LUT2 #(
		.INIT('h2)
	) name5332 (
		\u6_mem_reg[1][3]/NET0131 ,
		_w7402_,
		_w7478_
	);
	LUT2 #(
		.INIT('h8)
	) name5333 (
		\u12_dout_reg[3]/P0001 ,
		_w7402_,
		_w7479_
	);
	LUT2 #(
		.INIT('h1)
	) name5334 (
		_w7478_,
		_w7479_,
		_w7480_
	);
	LUT2 #(
		.INIT('h2)
	) name5335 (
		\u6_mem_reg[1][4]/NET0131 ,
		_w7402_,
		_w7481_
	);
	LUT2 #(
		.INIT('h8)
	) name5336 (
		\u12_dout_reg[4]/P0001 ,
		_w7402_,
		_w7482_
	);
	LUT2 #(
		.INIT('h1)
	) name5337 (
		_w7481_,
		_w7482_,
		_w7483_
	);
	LUT2 #(
		.INIT('h2)
	) name5338 (
		\u6_mem_reg[1][5]/NET0131 ,
		_w7402_,
		_w7484_
	);
	LUT2 #(
		.INIT('h8)
	) name5339 (
		\u12_dout_reg[5]/P0001 ,
		_w7402_,
		_w7485_
	);
	LUT2 #(
		.INIT('h1)
	) name5340 (
		_w7484_,
		_w7485_,
		_w7486_
	);
	LUT2 #(
		.INIT('h2)
	) name5341 (
		\u6_mem_reg[1][6]/NET0131 ,
		_w7402_,
		_w7487_
	);
	LUT2 #(
		.INIT('h8)
	) name5342 (
		\u12_dout_reg[6]/P0001 ,
		_w7402_,
		_w7488_
	);
	LUT2 #(
		.INIT('h1)
	) name5343 (
		_w7487_,
		_w7488_,
		_w7489_
	);
	LUT2 #(
		.INIT('h2)
	) name5344 (
		\u6_mem_reg[1][7]/NET0131 ,
		_w7402_,
		_w7490_
	);
	LUT2 #(
		.INIT('h8)
	) name5345 (
		\u12_dout_reg[7]/P0001 ,
		_w7402_,
		_w7491_
	);
	LUT2 #(
		.INIT('h1)
	) name5346 (
		_w7490_,
		_w7491_,
		_w7492_
	);
	LUT2 #(
		.INIT('h2)
	) name5347 (
		\u6_mem_reg[1][8]/NET0131 ,
		_w7402_,
		_w7493_
	);
	LUT2 #(
		.INIT('h8)
	) name5348 (
		\u12_dout_reg[8]/P0001 ,
		_w7402_,
		_w7494_
	);
	LUT2 #(
		.INIT('h1)
	) name5349 (
		_w7493_,
		_w7494_,
		_w7495_
	);
	LUT2 #(
		.INIT('h2)
	) name5350 (
		\u6_mem_reg[1][9]/NET0131 ,
		_w7402_,
		_w7496_
	);
	LUT2 #(
		.INIT('h8)
	) name5351 (
		\u12_dout_reg[9]/P0001 ,
		_w7402_,
		_w7497_
	);
	LUT2 #(
		.INIT('h1)
	) name5352 (
		_w7496_,
		_w7497_,
		_w7498_
	);
	LUT2 #(
		.INIT('h8)
	) name5353 (
		\u6_wp_reg[1]/NET0131 ,
		_w6419_,
		_w7499_
	);
	LUT2 #(
		.INIT('h2)
	) name5354 (
		\u6_mem_reg[2][0]/NET0131 ,
		_w7499_,
		_w7500_
	);
	LUT2 #(
		.INIT('h8)
	) name5355 (
		\u12_dout_reg[0]/P0001 ,
		_w7499_,
		_w7501_
	);
	LUT2 #(
		.INIT('h1)
	) name5356 (
		_w7500_,
		_w7501_,
		_w7502_
	);
	LUT2 #(
		.INIT('h2)
	) name5357 (
		\u6_mem_reg[2][10]/NET0131 ,
		_w7499_,
		_w7503_
	);
	LUT2 #(
		.INIT('h8)
	) name5358 (
		\u12_dout_reg[10]/P0001 ,
		_w7499_,
		_w7504_
	);
	LUT2 #(
		.INIT('h1)
	) name5359 (
		_w7503_,
		_w7504_,
		_w7505_
	);
	LUT2 #(
		.INIT('h2)
	) name5360 (
		\u6_mem_reg[2][11]/NET0131 ,
		_w7499_,
		_w7506_
	);
	LUT2 #(
		.INIT('h8)
	) name5361 (
		\u12_dout_reg[11]/P0001 ,
		_w7499_,
		_w7507_
	);
	LUT2 #(
		.INIT('h1)
	) name5362 (
		_w7506_,
		_w7507_,
		_w7508_
	);
	LUT2 #(
		.INIT('h2)
	) name5363 (
		\u6_mem_reg[2][12]/NET0131 ,
		_w7499_,
		_w7509_
	);
	LUT2 #(
		.INIT('h8)
	) name5364 (
		\u12_dout_reg[12]/P0001 ,
		_w7499_,
		_w7510_
	);
	LUT2 #(
		.INIT('h1)
	) name5365 (
		_w7509_,
		_w7510_,
		_w7511_
	);
	LUT2 #(
		.INIT('h2)
	) name5366 (
		\u6_mem_reg[2][13]/NET0131 ,
		_w7499_,
		_w7512_
	);
	LUT2 #(
		.INIT('h8)
	) name5367 (
		\u12_dout_reg[13]/P0001 ,
		_w7499_,
		_w7513_
	);
	LUT2 #(
		.INIT('h1)
	) name5368 (
		_w7512_,
		_w7513_,
		_w7514_
	);
	LUT2 #(
		.INIT('h2)
	) name5369 (
		\u6_mem_reg[2][14]/NET0131 ,
		_w7499_,
		_w7515_
	);
	LUT2 #(
		.INIT('h8)
	) name5370 (
		\u12_dout_reg[14]/P0001 ,
		_w7499_,
		_w7516_
	);
	LUT2 #(
		.INIT('h1)
	) name5371 (
		_w7515_,
		_w7516_,
		_w7517_
	);
	LUT2 #(
		.INIT('h2)
	) name5372 (
		\u6_mem_reg[2][15]/NET0131 ,
		_w7499_,
		_w7518_
	);
	LUT2 #(
		.INIT('h8)
	) name5373 (
		\u12_dout_reg[15]/P0001 ,
		_w7499_,
		_w7519_
	);
	LUT2 #(
		.INIT('h1)
	) name5374 (
		_w7518_,
		_w7519_,
		_w7520_
	);
	LUT2 #(
		.INIT('h2)
	) name5375 (
		\u6_mem_reg[2][16]/NET0131 ,
		_w7499_,
		_w7521_
	);
	LUT2 #(
		.INIT('h8)
	) name5376 (
		\u12_dout_reg[16]/P0001 ,
		_w7499_,
		_w7522_
	);
	LUT2 #(
		.INIT('h1)
	) name5377 (
		_w7521_,
		_w7522_,
		_w7523_
	);
	LUT2 #(
		.INIT('h2)
	) name5378 (
		\u6_mem_reg[2][17]/NET0131 ,
		_w7499_,
		_w7524_
	);
	LUT2 #(
		.INIT('h8)
	) name5379 (
		\u12_dout_reg[17]/P0001 ,
		_w7499_,
		_w7525_
	);
	LUT2 #(
		.INIT('h1)
	) name5380 (
		_w7524_,
		_w7525_,
		_w7526_
	);
	LUT2 #(
		.INIT('h2)
	) name5381 (
		\u6_mem_reg[2][18]/NET0131 ,
		_w7499_,
		_w7527_
	);
	LUT2 #(
		.INIT('h8)
	) name5382 (
		\u12_dout_reg[18]/P0001 ,
		_w7499_,
		_w7528_
	);
	LUT2 #(
		.INIT('h1)
	) name5383 (
		_w7527_,
		_w7528_,
		_w7529_
	);
	LUT2 #(
		.INIT('h2)
	) name5384 (
		\u6_mem_reg[2][19]/NET0131 ,
		_w7499_,
		_w7530_
	);
	LUT2 #(
		.INIT('h8)
	) name5385 (
		\u12_dout_reg[19]/P0001 ,
		_w7499_,
		_w7531_
	);
	LUT2 #(
		.INIT('h1)
	) name5386 (
		_w7530_,
		_w7531_,
		_w7532_
	);
	LUT2 #(
		.INIT('h2)
	) name5387 (
		\u6_mem_reg[2][1]/NET0131 ,
		_w7499_,
		_w7533_
	);
	LUT2 #(
		.INIT('h8)
	) name5388 (
		\u12_dout_reg[1]/P0001 ,
		_w7499_,
		_w7534_
	);
	LUT2 #(
		.INIT('h1)
	) name5389 (
		_w7533_,
		_w7534_,
		_w7535_
	);
	LUT2 #(
		.INIT('h2)
	) name5390 (
		\u6_mem_reg[2][20]/NET0131 ,
		_w7499_,
		_w7536_
	);
	LUT2 #(
		.INIT('h8)
	) name5391 (
		\u12_dout_reg[20]/P0001 ,
		_w7499_,
		_w7537_
	);
	LUT2 #(
		.INIT('h1)
	) name5392 (
		_w7536_,
		_w7537_,
		_w7538_
	);
	LUT2 #(
		.INIT('h2)
	) name5393 (
		\u6_mem_reg[2][21]/NET0131 ,
		_w7499_,
		_w7539_
	);
	LUT2 #(
		.INIT('h8)
	) name5394 (
		\u12_dout_reg[21]/P0001 ,
		_w7499_,
		_w7540_
	);
	LUT2 #(
		.INIT('h1)
	) name5395 (
		_w7539_,
		_w7540_,
		_w7541_
	);
	LUT2 #(
		.INIT('h2)
	) name5396 (
		\u6_mem_reg[2][22]/NET0131 ,
		_w7499_,
		_w7542_
	);
	LUT2 #(
		.INIT('h8)
	) name5397 (
		\u12_dout_reg[22]/P0001 ,
		_w7499_,
		_w7543_
	);
	LUT2 #(
		.INIT('h1)
	) name5398 (
		_w7542_,
		_w7543_,
		_w7544_
	);
	LUT2 #(
		.INIT('h2)
	) name5399 (
		\u6_mem_reg[2][23]/NET0131 ,
		_w7499_,
		_w7545_
	);
	LUT2 #(
		.INIT('h8)
	) name5400 (
		\u12_dout_reg[23]/P0001 ,
		_w7499_,
		_w7546_
	);
	LUT2 #(
		.INIT('h1)
	) name5401 (
		_w7545_,
		_w7546_,
		_w7547_
	);
	LUT2 #(
		.INIT('h2)
	) name5402 (
		\u6_mem_reg[2][24]/NET0131 ,
		_w7499_,
		_w7548_
	);
	LUT2 #(
		.INIT('h8)
	) name5403 (
		\u12_dout_reg[24]/P0001 ,
		_w7499_,
		_w7549_
	);
	LUT2 #(
		.INIT('h1)
	) name5404 (
		_w7548_,
		_w7549_,
		_w7550_
	);
	LUT2 #(
		.INIT('h2)
	) name5405 (
		\u6_mem_reg[2][25]/NET0131 ,
		_w7499_,
		_w7551_
	);
	LUT2 #(
		.INIT('h8)
	) name5406 (
		\u12_dout_reg[25]/P0001 ,
		_w7499_,
		_w7552_
	);
	LUT2 #(
		.INIT('h1)
	) name5407 (
		_w7551_,
		_w7552_,
		_w7553_
	);
	LUT2 #(
		.INIT('h2)
	) name5408 (
		\u6_mem_reg[2][26]/NET0131 ,
		_w7499_,
		_w7554_
	);
	LUT2 #(
		.INIT('h8)
	) name5409 (
		\u12_dout_reg[26]/P0001 ,
		_w7499_,
		_w7555_
	);
	LUT2 #(
		.INIT('h1)
	) name5410 (
		_w7554_,
		_w7555_,
		_w7556_
	);
	LUT2 #(
		.INIT('h2)
	) name5411 (
		\u6_mem_reg[2][27]/NET0131 ,
		_w7499_,
		_w7557_
	);
	LUT2 #(
		.INIT('h8)
	) name5412 (
		\u12_dout_reg[27]/P0001 ,
		_w7499_,
		_w7558_
	);
	LUT2 #(
		.INIT('h1)
	) name5413 (
		_w7557_,
		_w7558_,
		_w7559_
	);
	LUT2 #(
		.INIT('h2)
	) name5414 (
		\u6_mem_reg[2][28]/NET0131 ,
		_w7499_,
		_w7560_
	);
	LUT2 #(
		.INIT('h8)
	) name5415 (
		\u12_dout_reg[28]/P0001 ,
		_w7499_,
		_w7561_
	);
	LUT2 #(
		.INIT('h1)
	) name5416 (
		_w7560_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('h2)
	) name5417 (
		\u6_mem_reg[2][29]/NET0131 ,
		_w7499_,
		_w7563_
	);
	LUT2 #(
		.INIT('h8)
	) name5418 (
		\u12_dout_reg[29]/P0001 ,
		_w7499_,
		_w7564_
	);
	LUT2 #(
		.INIT('h1)
	) name5419 (
		_w7563_,
		_w7564_,
		_w7565_
	);
	LUT2 #(
		.INIT('h2)
	) name5420 (
		\u6_mem_reg[2][2]/NET0131 ,
		_w7499_,
		_w7566_
	);
	LUT2 #(
		.INIT('h8)
	) name5421 (
		\u12_dout_reg[2]/P0001 ,
		_w7499_,
		_w7567_
	);
	LUT2 #(
		.INIT('h1)
	) name5422 (
		_w7566_,
		_w7567_,
		_w7568_
	);
	LUT2 #(
		.INIT('h2)
	) name5423 (
		\u6_mem_reg[2][30]/NET0131 ,
		_w7499_,
		_w7569_
	);
	LUT2 #(
		.INIT('h8)
	) name5424 (
		\u12_dout_reg[30]/P0001 ,
		_w7499_,
		_w7570_
	);
	LUT2 #(
		.INIT('h1)
	) name5425 (
		_w7569_,
		_w7570_,
		_w7571_
	);
	LUT2 #(
		.INIT('h2)
	) name5426 (
		\u6_mem_reg[2][31]/NET0131 ,
		_w7499_,
		_w7572_
	);
	LUT2 #(
		.INIT('h8)
	) name5427 (
		\u12_dout_reg[31]/P0001 ,
		_w7499_,
		_w7573_
	);
	LUT2 #(
		.INIT('h1)
	) name5428 (
		_w7572_,
		_w7573_,
		_w7574_
	);
	LUT2 #(
		.INIT('h2)
	) name5429 (
		\u6_mem_reg[2][3]/NET0131 ,
		_w7499_,
		_w7575_
	);
	LUT2 #(
		.INIT('h8)
	) name5430 (
		\u12_dout_reg[3]/P0001 ,
		_w7499_,
		_w7576_
	);
	LUT2 #(
		.INIT('h1)
	) name5431 (
		_w7575_,
		_w7576_,
		_w7577_
	);
	LUT2 #(
		.INIT('h2)
	) name5432 (
		\u6_mem_reg[2][4]/NET0131 ,
		_w7499_,
		_w7578_
	);
	LUT2 #(
		.INIT('h8)
	) name5433 (
		\u12_dout_reg[4]/P0001 ,
		_w7499_,
		_w7579_
	);
	LUT2 #(
		.INIT('h1)
	) name5434 (
		_w7578_,
		_w7579_,
		_w7580_
	);
	LUT2 #(
		.INIT('h2)
	) name5435 (
		\u6_mem_reg[2][5]/NET0131 ,
		_w7499_,
		_w7581_
	);
	LUT2 #(
		.INIT('h8)
	) name5436 (
		\u12_dout_reg[5]/P0001 ,
		_w7499_,
		_w7582_
	);
	LUT2 #(
		.INIT('h1)
	) name5437 (
		_w7581_,
		_w7582_,
		_w7583_
	);
	LUT2 #(
		.INIT('h2)
	) name5438 (
		\u6_mem_reg[2][6]/NET0131 ,
		_w7499_,
		_w7584_
	);
	LUT2 #(
		.INIT('h8)
	) name5439 (
		\u12_dout_reg[6]/P0001 ,
		_w7499_,
		_w7585_
	);
	LUT2 #(
		.INIT('h1)
	) name5440 (
		_w7584_,
		_w7585_,
		_w7586_
	);
	LUT2 #(
		.INIT('h2)
	) name5441 (
		\u6_mem_reg[2][7]/NET0131 ,
		_w7499_,
		_w7587_
	);
	LUT2 #(
		.INIT('h8)
	) name5442 (
		\u12_dout_reg[7]/P0001 ,
		_w7499_,
		_w7588_
	);
	LUT2 #(
		.INIT('h1)
	) name5443 (
		_w7587_,
		_w7588_,
		_w7589_
	);
	LUT2 #(
		.INIT('h2)
	) name5444 (
		\u6_mem_reg[2][8]/NET0131 ,
		_w7499_,
		_w7590_
	);
	LUT2 #(
		.INIT('h8)
	) name5445 (
		\u12_dout_reg[8]/P0001 ,
		_w7499_,
		_w7591_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		_w7590_,
		_w7591_,
		_w7592_
	);
	LUT2 #(
		.INIT('h2)
	) name5447 (
		\u6_mem_reg[2][9]/NET0131 ,
		_w7499_,
		_w7593_
	);
	LUT2 #(
		.INIT('h8)
	) name5448 (
		\u12_dout_reg[9]/P0001 ,
		_w7499_,
		_w7594_
	);
	LUT2 #(
		.INIT('h1)
	) name5449 (
		_w7593_,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('h2)
	) name5450 (
		\u6_mem_reg[3][0]/NET0131 ,
		_w6325_,
		_w7596_
	);
	LUT2 #(
		.INIT('h8)
	) name5451 (
		\u12_dout_reg[0]/P0001 ,
		_w6325_,
		_w7597_
	);
	LUT2 #(
		.INIT('h1)
	) name5452 (
		_w7596_,
		_w7597_,
		_w7598_
	);
	LUT2 #(
		.INIT('h2)
	) name5453 (
		\u6_mem_reg[3][10]/NET0131 ,
		_w6325_,
		_w7599_
	);
	LUT2 #(
		.INIT('h8)
	) name5454 (
		\u12_dout_reg[10]/P0001 ,
		_w6325_,
		_w7600_
	);
	LUT2 #(
		.INIT('h1)
	) name5455 (
		_w7599_,
		_w7600_,
		_w7601_
	);
	LUT2 #(
		.INIT('h2)
	) name5456 (
		\u6_mem_reg[3][11]/NET0131 ,
		_w6325_,
		_w7602_
	);
	LUT2 #(
		.INIT('h8)
	) name5457 (
		\u12_dout_reg[11]/P0001 ,
		_w6325_,
		_w7603_
	);
	LUT2 #(
		.INIT('h1)
	) name5458 (
		_w7602_,
		_w7603_,
		_w7604_
	);
	LUT2 #(
		.INIT('h2)
	) name5459 (
		\u6_mem_reg[3][12]/NET0131 ,
		_w6325_,
		_w7605_
	);
	LUT2 #(
		.INIT('h8)
	) name5460 (
		\u12_dout_reg[12]/P0001 ,
		_w6325_,
		_w7606_
	);
	LUT2 #(
		.INIT('h1)
	) name5461 (
		_w7605_,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h2)
	) name5462 (
		\u6_mem_reg[3][13]/NET0131 ,
		_w6325_,
		_w7608_
	);
	LUT2 #(
		.INIT('h8)
	) name5463 (
		\u12_dout_reg[13]/P0001 ,
		_w6325_,
		_w7609_
	);
	LUT2 #(
		.INIT('h1)
	) name5464 (
		_w7608_,
		_w7609_,
		_w7610_
	);
	LUT2 #(
		.INIT('h2)
	) name5465 (
		\u6_mem_reg[3][14]/NET0131 ,
		_w6325_,
		_w7611_
	);
	LUT2 #(
		.INIT('h8)
	) name5466 (
		\u12_dout_reg[14]/P0001 ,
		_w6325_,
		_w7612_
	);
	LUT2 #(
		.INIT('h1)
	) name5467 (
		_w7611_,
		_w7612_,
		_w7613_
	);
	LUT2 #(
		.INIT('h2)
	) name5468 (
		\u6_mem_reg[3][15]/NET0131 ,
		_w6325_,
		_w7614_
	);
	LUT2 #(
		.INIT('h8)
	) name5469 (
		\u12_dout_reg[15]/P0001 ,
		_w6325_,
		_w7615_
	);
	LUT2 #(
		.INIT('h1)
	) name5470 (
		_w7614_,
		_w7615_,
		_w7616_
	);
	LUT2 #(
		.INIT('h2)
	) name5471 (
		\u6_mem_reg[3][16]/NET0131 ,
		_w6325_,
		_w7617_
	);
	LUT2 #(
		.INIT('h8)
	) name5472 (
		\u12_dout_reg[16]/P0001 ,
		_w6325_,
		_w7618_
	);
	LUT2 #(
		.INIT('h1)
	) name5473 (
		_w7617_,
		_w7618_,
		_w7619_
	);
	LUT2 #(
		.INIT('h2)
	) name5474 (
		\u6_mem_reg[3][17]/NET0131 ,
		_w6325_,
		_w7620_
	);
	LUT2 #(
		.INIT('h8)
	) name5475 (
		\u12_dout_reg[17]/P0001 ,
		_w6325_,
		_w7621_
	);
	LUT2 #(
		.INIT('h1)
	) name5476 (
		_w7620_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('h2)
	) name5477 (
		\u6_mem_reg[3][18]/NET0131 ,
		_w6325_,
		_w7623_
	);
	LUT2 #(
		.INIT('h8)
	) name5478 (
		\u12_dout_reg[18]/P0001 ,
		_w6325_,
		_w7624_
	);
	LUT2 #(
		.INIT('h1)
	) name5479 (
		_w7623_,
		_w7624_,
		_w7625_
	);
	LUT2 #(
		.INIT('h2)
	) name5480 (
		\u6_mem_reg[3][19]/NET0131 ,
		_w6325_,
		_w7626_
	);
	LUT2 #(
		.INIT('h8)
	) name5481 (
		\u12_dout_reg[19]/P0001 ,
		_w6325_,
		_w7627_
	);
	LUT2 #(
		.INIT('h1)
	) name5482 (
		_w7626_,
		_w7627_,
		_w7628_
	);
	LUT2 #(
		.INIT('h2)
	) name5483 (
		\u6_mem_reg[3][1]/NET0131 ,
		_w6325_,
		_w7629_
	);
	LUT2 #(
		.INIT('h8)
	) name5484 (
		\u12_dout_reg[1]/P0001 ,
		_w6325_,
		_w7630_
	);
	LUT2 #(
		.INIT('h1)
	) name5485 (
		_w7629_,
		_w7630_,
		_w7631_
	);
	LUT2 #(
		.INIT('h2)
	) name5486 (
		\u6_mem_reg[3][20]/NET0131 ,
		_w6325_,
		_w7632_
	);
	LUT2 #(
		.INIT('h8)
	) name5487 (
		\u12_dout_reg[20]/P0001 ,
		_w6325_,
		_w7633_
	);
	LUT2 #(
		.INIT('h1)
	) name5488 (
		_w7632_,
		_w7633_,
		_w7634_
	);
	LUT2 #(
		.INIT('h2)
	) name5489 (
		\u6_mem_reg[3][21]/NET0131 ,
		_w6325_,
		_w7635_
	);
	LUT2 #(
		.INIT('h8)
	) name5490 (
		\u12_dout_reg[21]/P0001 ,
		_w6325_,
		_w7636_
	);
	LUT2 #(
		.INIT('h1)
	) name5491 (
		_w7635_,
		_w7636_,
		_w7637_
	);
	LUT2 #(
		.INIT('h2)
	) name5492 (
		\u6_mem_reg[3][22]/NET0131 ,
		_w6325_,
		_w7638_
	);
	LUT2 #(
		.INIT('h8)
	) name5493 (
		\u12_dout_reg[22]/P0001 ,
		_w6325_,
		_w7639_
	);
	LUT2 #(
		.INIT('h1)
	) name5494 (
		_w7638_,
		_w7639_,
		_w7640_
	);
	LUT2 #(
		.INIT('h2)
	) name5495 (
		\u6_mem_reg[3][23]/NET0131 ,
		_w6325_,
		_w7641_
	);
	LUT2 #(
		.INIT('h8)
	) name5496 (
		\u12_dout_reg[23]/P0001 ,
		_w6325_,
		_w7642_
	);
	LUT2 #(
		.INIT('h1)
	) name5497 (
		_w7641_,
		_w7642_,
		_w7643_
	);
	LUT2 #(
		.INIT('h2)
	) name5498 (
		\u6_mem_reg[3][24]/NET0131 ,
		_w6325_,
		_w7644_
	);
	LUT2 #(
		.INIT('h8)
	) name5499 (
		\u12_dout_reg[24]/P0001 ,
		_w6325_,
		_w7645_
	);
	LUT2 #(
		.INIT('h1)
	) name5500 (
		_w7644_,
		_w7645_,
		_w7646_
	);
	LUT2 #(
		.INIT('h2)
	) name5501 (
		\u6_mem_reg[3][25]/NET0131 ,
		_w6325_,
		_w7647_
	);
	LUT2 #(
		.INIT('h8)
	) name5502 (
		\u12_dout_reg[25]/P0001 ,
		_w6325_,
		_w7648_
	);
	LUT2 #(
		.INIT('h1)
	) name5503 (
		_w7647_,
		_w7648_,
		_w7649_
	);
	LUT2 #(
		.INIT('h2)
	) name5504 (
		\u6_mem_reg[3][26]/NET0131 ,
		_w6325_,
		_w7650_
	);
	LUT2 #(
		.INIT('h8)
	) name5505 (
		\u12_dout_reg[26]/P0001 ,
		_w6325_,
		_w7651_
	);
	LUT2 #(
		.INIT('h1)
	) name5506 (
		_w7650_,
		_w7651_,
		_w7652_
	);
	LUT2 #(
		.INIT('h2)
	) name5507 (
		\u6_mem_reg[3][27]/NET0131 ,
		_w6325_,
		_w7653_
	);
	LUT2 #(
		.INIT('h8)
	) name5508 (
		\u12_dout_reg[27]/P0001 ,
		_w6325_,
		_w7654_
	);
	LUT2 #(
		.INIT('h1)
	) name5509 (
		_w7653_,
		_w7654_,
		_w7655_
	);
	LUT2 #(
		.INIT('h2)
	) name5510 (
		\u6_mem_reg[3][28]/NET0131 ,
		_w6325_,
		_w7656_
	);
	LUT2 #(
		.INIT('h8)
	) name5511 (
		\u12_dout_reg[28]/P0001 ,
		_w6325_,
		_w7657_
	);
	LUT2 #(
		.INIT('h1)
	) name5512 (
		_w7656_,
		_w7657_,
		_w7658_
	);
	LUT2 #(
		.INIT('h2)
	) name5513 (
		\u6_mem_reg[3][29]/NET0131 ,
		_w6325_,
		_w7659_
	);
	LUT2 #(
		.INIT('h8)
	) name5514 (
		\u12_dout_reg[29]/P0001 ,
		_w6325_,
		_w7660_
	);
	LUT2 #(
		.INIT('h1)
	) name5515 (
		_w7659_,
		_w7660_,
		_w7661_
	);
	LUT2 #(
		.INIT('h2)
	) name5516 (
		\u6_mem_reg[3][2]/NET0131 ,
		_w6325_,
		_w7662_
	);
	LUT2 #(
		.INIT('h8)
	) name5517 (
		\u12_dout_reg[2]/P0001 ,
		_w6325_,
		_w7663_
	);
	LUT2 #(
		.INIT('h1)
	) name5518 (
		_w7662_,
		_w7663_,
		_w7664_
	);
	LUT2 #(
		.INIT('h2)
	) name5519 (
		\u6_mem_reg[3][30]/NET0131 ,
		_w6325_,
		_w7665_
	);
	LUT2 #(
		.INIT('h8)
	) name5520 (
		\u12_dout_reg[30]/P0001 ,
		_w6325_,
		_w7666_
	);
	LUT2 #(
		.INIT('h1)
	) name5521 (
		_w7665_,
		_w7666_,
		_w7667_
	);
	LUT2 #(
		.INIT('h2)
	) name5522 (
		\u6_mem_reg[3][31]/NET0131 ,
		_w6325_,
		_w7668_
	);
	LUT2 #(
		.INIT('h8)
	) name5523 (
		\u12_dout_reg[31]/P0001 ,
		_w6325_,
		_w7669_
	);
	LUT2 #(
		.INIT('h1)
	) name5524 (
		_w7668_,
		_w7669_,
		_w7670_
	);
	LUT2 #(
		.INIT('h2)
	) name5525 (
		\u6_mem_reg[3][3]/NET0131 ,
		_w6325_,
		_w7671_
	);
	LUT2 #(
		.INIT('h8)
	) name5526 (
		\u12_dout_reg[3]/P0001 ,
		_w6325_,
		_w7672_
	);
	LUT2 #(
		.INIT('h1)
	) name5527 (
		_w7671_,
		_w7672_,
		_w7673_
	);
	LUT2 #(
		.INIT('h2)
	) name5528 (
		\u6_mem_reg[3][4]/NET0131 ,
		_w6325_,
		_w7674_
	);
	LUT2 #(
		.INIT('h8)
	) name5529 (
		\u12_dout_reg[4]/P0001 ,
		_w6325_,
		_w7675_
	);
	LUT2 #(
		.INIT('h1)
	) name5530 (
		_w7674_,
		_w7675_,
		_w7676_
	);
	LUT2 #(
		.INIT('h2)
	) name5531 (
		\u6_mem_reg[3][5]/NET0131 ,
		_w6325_,
		_w7677_
	);
	LUT2 #(
		.INIT('h8)
	) name5532 (
		\u12_dout_reg[5]/P0001 ,
		_w6325_,
		_w7678_
	);
	LUT2 #(
		.INIT('h1)
	) name5533 (
		_w7677_,
		_w7678_,
		_w7679_
	);
	LUT2 #(
		.INIT('h2)
	) name5534 (
		\u6_mem_reg[3][6]/NET0131 ,
		_w6325_,
		_w7680_
	);
	LUT2 #(
		.INIT('h8)
	) name5535 (
		\u12_dout_reg[6]/P0001 ,
		_w6325_,
		_w7681_
	);
	LUT2 #(
		.INIT('h1)
	) name5536 (
		_w7680_,
		_w7681_,
		_w7682_
	);
	LUT2 #(
		.INIT('h2)
	) name5537 (
		\u6_mem_reg[3][7]/NET0131 ,
		_w6325_,
		_w7683_
	);
	LUT2 #(
		.INIT('h8)
	) name5538 (
		\u12_dout_reg[7]/P0001 ,
		_w6325_,
		_w7684_
	);
	LUT2 #(
		.INIT('h1)
	) name5539 (
		_w7683_,
		_w7684_,
		_w7685_
	);
	LUT2 #(
		.INIT('h2)
	) name5540 (
		\u6_mem_reg[3][8]/NET0131 ,
		_w6325_,
		_w7686_
	);
	LUT2 #(
		.INIT('h8)
	) name5541 (
		\u12_dout_reg[8]/P0001 ,
		_w6325_,
		_w7687_
	);
	LUT2 #(
		.INIT('h1)
	) name5542 (
		_w7686_,
		_w7687_,
		_w7688_
	);
	LUT2 #(
		.INIT('h2)
	) name5543 (
		\u6_mem_reg[3][9]/NET0131 ,
		_w6325_,
		_w7689_
	);
	LUT2 #(
		.INIT('h8)
	) name5544 (
		\u12_dout_reg[9]/P0001 ,
		_w6325_,
		_w7690_
	);
	LUT2 #(
		.INIT('h1)
	) name5545 (
		_w7689_,
		_w7690_,
		_w7691_
	);
	LUT2 #(
		.INIT('h2)
	) name5546 (
		\u8_mem_reg[1][6]/NET0131 ,
		_w6629_,
		_w7692_
	);
	LUT2 #(
		.INIT('h8)
	) name5547 (
		\u12_dout_reg[6]/P0001 ,
		_w6629_,
		_w7693_
	);
	LUT2 #(
		.INIT('h1)
	) name5548 (
		_w7692_,
		_w7693_,
		_w7694_
	);
	LUT2 #(
		.INIT('h2)
	) name5549 (
		\u3_mem_reg[2][25]/NET0131 ,
		_w6583_,
		_w7695_
	);
	LUT2 #(
		.INIT('h8)
	) name5550 (
		\u12_dout_reg[25]/P0001 ,
		_w6583_,
		_w7696_
	);
	LUT2 #(
		.INIT('h1)
	) name5551 (
		_w7695_,
		_w7696_,
		_w7697_
	);
	LUT2 #(
		.INIT('h2)
	) name5552 (
		\u8_mem_reg[3][4]/NET0131 ,
		_w6301_,
		_w7698_
	);
	LUT2 #(
		.INIT('h8)
	) name5553 (
		\u12_dout_reg[4]/P0001 ,
		_w6301_,
		_w7699_
	);
	LUT2 #(
		.INIT('h1)
	) name5554 (
		_w7698_,
		_w7699_,
		_w7700_
	);
	LUT2 #(
		.INIT('h2)
	) name5555 (
		\u3_mem_reg[3][3]/NET0131 ,
		_w6319_,
		_w7701_
	);
	LUT2 #(
		.INIT('h8)
	) name5556 (
		\u12_dout_reg[3]/P0001 ,
		_w6319_,
		_w7702_
	);
	LUT2 #(
		.INIT('h1)
	) name5557 (
		_w7701_,
		_w7702_,
		_w7703_
	);
	LUT2 #(
		.INIT('h2)
	) name5558 (
		\u8_mem_reg[3][8]/NET0131 ,
		_w6301_,
		_w7704_
	);
	LUT2 #(
		.INIT('h8)
	) name5559 (
		\u12_dout_reg[8]/P0001 ,
		_w6301_,
		_w7705_
	);
	LUT2 #(
		.INIT('h1)
	) name5560 (
		_w7704_,
		_w7705_,
		_w7706_
	);
	LUT2 #(
		.INIT('h2)
	) name5561 (
		\u3_mem_reg[1][14]/NET0131 ,
		_w6489_,
		_w7707_
	);
	LUT2 #(
		.INIT('h8)
	) name5562 (
		\u12_dout_reg[14]/P0001 ,
		_w6489_,
		_w7708_
	);
	LUT2 #(
		.INIT('h1)
	) name5563 (
		_w7707_,
		_w7708_,
		_w7709_
	);
	LUT2 #(
		.INIT('h4)
	) name5564 (
		\u7_wp_reg[1]/NET0131 ,
		_w6330_,
		_w7710_
	);
	LUT2 #(
		.INIT('h2)
	) name5565 (
		\u7_mem_reg[1][0]/NET0131 ,
		_w7710_,
		_w7711_
	);
	LUT2 #(
		.INIT('h8)
	) name5566 (
		\u12_dout_reg[0]/P0001 ,
		_w7710_,
		_w7712_
	);
	LUT2 #(
		.INIT('h1)
	) name5567 (
		_w7711_,
		_w7712_,
		_w7713_
	);
	LUT2 #(
		.INIT('h2)
	) name5568 (
		\u7_mem_reg[1][10]/NET0131 ,
		_w7710_,
		_w7714_
	);
	LUT2 #(
		.INIT('h8)
	) name5569 (
		\u12_dout_reg[10]/P0001 ,
		_w7710_,
		_w7715_
	);
	LUT2 #(
		.INIT('h1)
	) name5570 (
		_w7714_,
		_w7715_,
		_w7716_
	);
	LUT2 #(
		.INIT('h2)
	) name5571 (
		\u7_mem_reg[1][11]/NET0131 ,
		_w7710_,
		_w7717_
	);
	LUT2 #(
		.INIT('h8)
	) name5572 (
		\u12_dout_reg[11]/P0001 ,
		_w7710_,
		_w7718_
	);
	LUT2 #(
		.INIT('h1)
	) name5573 (
		_w7717_,
		_w7718_,
		_w7719_
	);
	LUT2 #(
		.INIT('h2)
	) name5574 (
		\u3_mem_reg[1][23]/NET0131 ,
		_w6489_,
		_w7720_
	);
	LUT2 #(
		.INIT('h8)
	) name5575 (
		\u12_dout_reg[23]/P0001 ,
		_w6489_,
		_w7721_
	);
	LUT2 #(
		.INIT('h1)
	) name5576 (
		_w7720_,
		_w7721_,
		_w7722_
	);
	LUT2 #(
		.INIT('h2)
	) name5577 (
		\u7_mem_reg[1][12]/NET0131 ,
		_w7710_,
		_w7723_
	);
	LUT2 #(
		.INIT('h8)
	) name5578 (
		\u12_dout_reg[12]/P0001 ,
		_w7710_,
		_w7724_
	);
	LUT2 #(
		.INIT('h1)
	) name5579 (
		_w7723_,
		_w7724_,
		_w7725_
	);
	LUT2 #(
		.INIT('h2)
	) name5580 (
		\u7_mem_reg[1][13]/NET0131 ,
		_w7710_,
		_w7726_
	);
	LUT2 #(
		.INIT('h8)
	) name5581 (
		\u12_dout_reg[13]/P0001 ,
		_w7710_,
		_w7727_
	);
	LUT2 #(
		.INIT('h1)
	) name5582 (
		_w7726_,
		_w7727_,
		_w7728_
	);
	LUT2 #(
		.INIT('h2)
	) name5583 (
		\u7_mem_reg[1][14]/NET0131 ,
		_w7710_,
		_w7729_
	);
	LUT2 #(
		.INIT('h8)
	) name5584 (
		\u12_dout_reg[14]/P0001 ,
		_w7710_,
		_w7730_
	);
	LUT2 #(
		.INIT('h1)
	) name5585 (
		_w7729_,
		_w7730_,
		_w7731_
	);
	LUT2 #(
		.INIT('h2)
	) name5586 (
		\u7_mem_reg[1][15]/NET0131 ,
		_w7710_,
		_w7732_
	);
	LUT2 #(
		.INIT('h8)
	) name5587 (
		\u12_dout_reg[15]/P0001 ,
		_w7710_,
		_w7733_
	);
	LUT2 #(
		.INIT('h1)
	) name5588 (
		_w7732_,
		_w7733_,
		_w7734_
	);
	LUT2 #(
		.INIT('h2)
	) name5589 (
		\u7_mem_reg[1][16]/NET0131 ,
		_w7710_,
		_w7735_
	);
	LUT2 #(
		.INIT('h8)
	) name5590 (
		\u12_dout_reg[16]/P0001 ,
		_w7710_,
		_w7736_
	);
	LUT2 #(
		.INIT('h1)
	) name5591 (
		_w7735_,
		_w7736_,
		_w7737_
	);
	LUT2 #(
		.INIT('h2)
	) name5592 (
		\u7_mem_reg[1][17]/NET0131 ,
		_w7710_,
		_w7738_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		\u12_dout_reg[17]/P0001 ,
		_w7710_,
		_w7739_
	);
	LUT2 #(
		.INIT('h1)
	) name5594 (
		_w7738_,
		_w7739_,
		_w7740_
	);
	LUT2 #(
		.INIT('h2)
	) name5595 (
		\u7_mem_reg[1][18]/NET0131 ,
		_w7710_,
		_w7741_
	);
	LUT2 #(
		.INIT('h8)
	) name5596 (
		\u12_dout_reg[18]/P0001 ,
		_w7710_,
		_w7742_
	);
	LUT2 #(
		.INIT('h1)
	) name5597 (
		_w7741_,
		_w7742_,
		_w7743_
	);
	LUT2 #(
		.INIT('h2)
	) name5598 (
		\u7_mem_reg[1][19]/NET0131 ,
		_w7710_,
		_w7744_
	);
	LUT2 #(
		.INIT('h8)
	) name5599 (
		\u12_dout_reg[19]/P0001 ,
		_w7710_,
		_w7745_
	);
	LUT2 #(
		.INIT('h1)
	) name5600 (
		_w7744_,
		_w7745_,
		_w7746_
	);
	LUT2 #(
		.INIT('h2)
	) name5601 (
		\u7_mem_reg[1][1]/NET0131 ,
		_w7710_,
		_w7747_
	);
	LUT2 #(
		.INIT('h8)
	) name5602 (
		\u12_dout_reg[1]/P0001 ,
		_w7710_,
		_w7748_
	);
	LUT2 #(
		.INIT('h1)
	) name5603 (
		_w7747_,
		_w7748_,
		_w7749_
	);
	LUT2 #(
		.INIT('h2)
	) name5604 (
		\u7_mem_reg[1][20]/NET0131 ,
		_w7710_,
		_w7750_
	);
	LUT2 #(
		.INIT('h8)
	) name5605 (
		\u12_dout_reg[20]/P0001 ,
		_w7710_,
		_w7751_
	);
	LUT2 #(
		.INIT('h1)
	) name5606 (
		_w7750_,
		_w7751_,
		_w7752_
	);
	LUT2 #(
		.INIT('h2)
	) name5607 (
		\u7_mem_reg[1][21]/NET0131 ,
		_w7710_,
		_w7753_
	);
	LUT2 #(
		.INIT('h8)
	) name5608 (
		\u12_dout_reg[21]/P0001 ,
		_w7710_,
		_w7754_
	);
	LUT2 #(
		.INIT('h1)
	) name5609 (
		_w7753_,
		_w7754_,
		_w7755_
	);
	LUT2 #(
		.INIT('h2)
	) name5610 (
		\u7_mem_reg[1][22]/NET0131 ,
		_w7710_,
		_w7756_
	);
	LUT2 #(
		.INIT('h8)
	) name5611 (
		\u12_dout_reg[22]/P0001 ,
		_w7710_,
		_w7757_
	);
	LUT2 #(
		.INIT('h1)
	) name5612 (
		_w7756_,
		_w7757_,
		_w7758_
	);
	LUT2 #(
		.INIT('h2)
	) name5613 (
		\u7_mem_reg[1][23]/NET0131 ,
		_w7710_,
		_w7759_
	);
	LUT2 #(
		.INIT('h8)
	) name5614 (
		\u12_dout_reg[23]/P0001 ,
		_w7710_,
		_w7760_
	);
	LUT2 #(
		.INIT('h1)
	) name5615 (
		_w7759_,
		_w7760_,
		_w7761_
	);
	LUT2 #(
		.INIT('h2)
	) name5616 (
		\u7_mem_reg[1][24]/NET0131 ,
		_w7710_,
		_w7762_
	);
	LUT2 #(
		.INIT('h8)
	) name5617 (
		\u12_dout_reg[24]/P0001 ,
		_w7710_,
		_w7763_
	);
	LUT2 #(
		.INIT('h1)
	) name5618 (
		_w7762_,
		_w7763_,
		_w7764_
	);
	LUT2 #(
		.INIT('h2)
	) name5619 (
		\u7_mem_reg[1][25]/NET0131 ,
		_w7710_,
		_w7765_
	);
	LUT2 #(
		.INIT('h8)
	) name5620 (
		\u12_dout_reg[25]/P0001 ,
		_w7710_,
		_w7766_
	);
	LUT2 #(
		.INIT('h1)
	) name5621 (
		_w7765_,
		_w7766_,
		_w7767_
	);
	LUT2 #(
		.INIT('h2)
	) name5622 (
		\u7_mem_reg[1][26]/NET0131 ,
		_w7710_,
		_w7768_
	);
	LUT2 #(
		.INIT('h8)
	) name5623 (
		\u12_dout_reg[26]/P0001 ,
		_w7710_,
		_w7769_
	);
	LUT2 #(
		.INIT('h1)
	) name5624 (
		_w7768_,
		_w7769_,
		_w7770_
	);
	LUT2 #(
		.INIT('h2)
	) name5625 (
		\u7_mem_reg[1][27]/NET0131 ,
		_w7710_,
		_w7771_
	);
	LUT2 #(
		.INIT('h8)
	) name5626 (
		\u12_dout_reg[27]/P0001 ,
		_w7710_,
		_w7772_
	);
	LUT2 #(
		.INIT('h1)
	) name5627 (
		_w7771_,
		_w7772_,
		_w7773_
	);
	LUT2 #(
		.INIT('h2)
	) name5628 (
		\u7_mem_reg[1][28]/NET0131 ,
		_w7710_,
		_w7774_
	);
	LUT2 #(
		.INIT('h8)
	) name5629 (
		\u12_dout_reg[28]/P0001 ,
		_w7710_,
		_w7775_
	);
	LUT2 #(
		.INIT('h1)
	) name5630 (
		_w7774_,
		_w7775_,
		_w7776_
	);
	LUT2 #(
		.INIT('h2)
	) name5631 (
		\u7_mem_reg[1][29]/NET0131 ,
		_w7710_,
		_w7777_
	);
	LUT2 #(
		.INIT('h8)
	) name5632 (
		\u12_dout_reg[29]/P0001 ,
		_w7710_,
		_w7778_
	);
	LUT2 #(
		.INIT('h1)
	) name5633 (
		_w7777_,
		_w7778_,
		_w7779_
	);
	LUT2 #(
		.INIT('h2)
	) name5634 (
		\u7_mem_reg[1][2]/NET0131 ,
		_w7710_,
		_w7780_
	);
	LUT2 #(
		.INIT('h8)
	) name5635 (
		\u12_dout_reg[2]/P0001 ,
		_w7710_,
		_w7781_
	);
	LUT2 #(
		.INIT('h1)
	) name5636 (
		_w7780_,
		_w7781_,
		_w7782_
	);
	LUT2 #(
		.INIT('h2)
	) name5637 (
		\u7_mem_reg[1][30]/NET0131 ,
		_w7710_,
		_w7783_
	);
	LUT2 #(
		.INIT('h8)
	) name5638 (
		\u12_dout_reg[30]/P0001 ,
		_w7710_,
		_w7784_
	);
	LUT2 #(
		.INIT('h1)
	) name5639 (
		_w7783_,
		_w7784_,
		_w7785_
	);
	LUT2 #(
		.INIT('h2)
	) name5640 (
		\u7_mem_reg[1][31]/NET0131 ,
		_w7710_,
		_w7786_
	);
	LUT2 #(
		.INIT('h8)
	) name5641 (
		\u12_dout_reg[31]/P0001 ,
		_w7710_,
		_w7787_
	);
	LUT2 #(
		.INIT('h1)
	) name5642 (
		_w7786_,
		_w7787_,
		_w7788_
	);
	LUT2 #(
		.INIT('h2)
	) name5643 (
		\u7_mem_reg[1][3]/NET0131 ,
		_w7710_,
		_w7789_
	);
	LUT2 #(
		.INIT('h8)
	) name5644 (
		\u12_dout_reg[3]/P0001 ,
		_w7710_,
		_w7790_
	);
	LUT2 #(
		.INIT('h1)
	) name5645 (
		_w7789_,
		_w7790_,
		_w7791_
	);
	LUT2 #(
		.INIT('h2)
	) name5646 (
		\u7_mem_reg[1][4]/NET0131 ,
		_w7710_,
		_w7792_
	);
	LUT2 #(
		.INIT('h8)
	) name5647 (
		\u12_dout_reg[4]/P0001 ,
		_w7710_,
		_w7793_
	);
	LUT2 #(
		.INIT('h1)
	) name5648 (
		_w7792_,
		_w7793_,
		_w7794_
	);
	LUT2 #(
		.INIT('h2)
	) name5649 (
		\u7_mem_reg[1][5]/NET0131 ,
		_w7710_,
		_w7795_
	);
	LUT2 #(
		.INIT('h8)
	) name5650 (
		\u12_dout_reg[5]/P0001 ,
		_w7710_,
		_w7796_
	);
	LUT2 #(
		.INIT('h1)
	) name5651 (
		_w7795_,
		_w7796_,
		_w7797_
	);
	LUT2 #(
		.INIT('h2)
	) name5652 (
		\u7_mem_reg[1][6]/NET0131 ,
		_w7710_,
		_w7798_
	);
	LUT2 #(
		.INIT('h8)
	) name5653 (
		\u12_dout_reg[6]/P0001 ,
		_w7710_,
		_w7799_
	);
	LUT2 #(
		.INIT('h1)
	) name5654 (
		_w7798_,
		_w7799_,
		_w7800_
	);
	LUT2 #(
		.INIT('h2)
	) name5655 (
		\u7_mem_reg[1][7]/NET0131 ,
		_w7710_,
		_w7801_
	);
	LUT2 #(
		.INIT('h8)
	) name5656 (
		\u12_dout_reg[7]/P0001 ,
		_w7710_,
		_w7802_
	);
	LUT2 #(
		.INIT('h1)
	) name5657 (
		_w7801_,
		_w7802_,
		_w7803_
	);
	LUT2 #(
		.INIT('h2)
	) name5658 (
		\u7_mem_reg[1][8]/NET0131 ,
		_w7710_,
		_w7804_
	);
	LUT2 #(
		.INIT('h8)
	) name5659 (
		\u12_dout_reg[8]/P0001 ,
		_w7710_,
		_w7805_
	);
	LUT2 #(
		.INIT('h1)
	) name5660 (
		_w7804_,
		_w7805_,
		_w7806_
	);
	LUT2 #(
		.INIT('h2)
	) name5661 (
		\u3_mem_reg[3][20]/NET0131 ,
		_w6319_,
		_w7807_
	);
	LUT2 #(
		.INIT('h8)
	) name5662 (
		\u12_dout_reg[20]/P0001 ,
		_w6319_,
		_w7808_
	);
	LUT2 #(
		.INIT('h1)
	) name5663 (
		_w7807_,
		_w7808_,
		_w7809_
	);
	LUT2 #(
		.INIT('h2)
	) name5664 (
		\u7_mem_reg[1][9]/NET0131 ,
		_w7710_,
		_w7810_
	);
	LUT2 #(
		.INIT('h8)
	) name5665 (
		\u12_dout_reg[9]/P0001 ,
		_w7710_,
		_w7811_
	);
	LUT2 #(
		.INIT('h1)
	) name5666 (
		_w7810_,
		_w7811_,
		_w7812_
	);
	LUT2 #(
		.INIT('h8)
	) name5667 (
		\u7_wp_reg[1]/NET0131 ,
		_w6423_,
		_w7813_
	);
	LUT2 #(
		.INIT('h2)
	) name5668 (
		\u7_mem_reg[2][0]/NET0131 ,
		_w7813_,
		_w7814_
	);
	LUT2 #(
		.INIT('h8)
	) name5669 (
		\u12_dout_reg[0]/P0001 ,
		_w7813_,
		_w7815_
	);
	LUT2 #(
		.INIT('h1)
	) name5670 (
		_w7814_,
		_w7815_,
		_w7816_
	);
	LUT2 #(
		.INIT('h2)
	) name5671 (
		\u7_mem_reg[2][10]/NET0131 ,
		_w7813_,
		_w7817_
	);
	LUT2 #(
		.INIT('h8)
	) name5672 (
		\u12_dout_reg[10]/P0001 ,
		_w7813_,
		_w7818_
	);
	LUT2 #(
		.INIT('h1)
	) name5673 (
		_w7817_,
		_w7818_,
		_w7819_
	);
	LUT2 #(
		.INIT('h2)
	) name5674 (
		\u7_mem_reg[2][11]/NET0131 ,
		_w7813_,
		_w7820_
	);
	LUT2 #(
		.INIT('h8)
	) name5675 (
		\u12_dout_reg[11]/P0001 ,
		_w7813_,
		_w7821_
	);
	LUT2 #(
		.INIT('h1)
	) name5676 (
		_w7820_,
		_w7821_,
		_w7822_
	);
	LUT2 #(
		.INIT('h2)
	) name5677 (
		\u7_mem_reg[2][12]/NET0131 ,
		_w7813_,
		_w7823_
	);
	LUT2 #(
		.INIT('h8)
	) name5678 (
		\u12_dout_reg[12]/P0001 ,
		_w7813_,
		_w7824_
	);
	LUT2 #(
		.INIT('h1)
	) name5679 (
		_w7823_,
		_w7824_,
		_w7825_
	);
	LUT2 #(
		.INIT('h2)
	) name5680 (
		\u7_mem_reg[2][13]/NET0131 ,
		_w7813_,
		_w7826_
	);
	LUT2 #(
		.INIT('h8)
	) name5681 (
		\u12_dout_reg[13]/P0001 ,
		_w7813_,
		_w7827_
	);
	LUT2 #(
		.INIT('h1)
	) name5682 (
		_w7826_,
		_w7827_,
		_w7828_
	);
	LUT2 #(
		.INIT('h2)
	) name5683 (
		\u7_mem_reg[2][14]/NET0131 ,
		_w7813_,
		_w7829_
	);
	LUT2 #(
		.INIT('h8)
	) name5684 (
		\u12_dout_reg[14]/P0001 ,
		_w7813_,
		_w7830_
	);
	LUT2 #(
		.INIT('h1)
	) name5685 (
		_w7829_,
		_w7830_,
		_w7831_
	);
	LUT2 #(
		.INIT('h2)
	) name5686 (
		\u7_mem_reg[2][15]/NET0131 ,
		_w7813_,
		_w7832_
	);
	LUT2 #(
		.INIT('h8)
	) name5687 (
		\u12_dout_reg[15]/P0001 ,
		_w7813_,
		_w7833_
	);
	LUT2 #(
		.INIT('h1)
	) name5688 (
		_w7832_,
		_w7833_,
		_w7834_
	);
	LUT2 #(
		.INIT('h2)
	) name5689 (
		\u7_mem_reg[2][16]/NET0131 ,
		_w7813_,
		_w7835_
	);
	LUT2 #(
		.INIT('h8)
	) name5690 (
		\u12_dout_reg[16]/P0001 ,
		_w7813_,
		_w7836_
	);
	LUT2 #(
		.INIT('h1)
	) name5691 (
		_w7835_,
		_w7836_,
		_w7837_
	);
	LUT2 #(
		.INIT('h2)
	) name5692 (
		\u7_mem_reg[2][17]/NET0131 ,
		_w7813_,
		_w7838_
	);
	LUT2 #(
		.INIT('h8)
	) name5693 (
		\u12_dout_reg[17]/P0001 ,
		_w7813_,
		_w7839_
	);
	LUT2 #(
		.INIT('h1)
	) name5694 (
		_w7838_,
		_w7839_,
		_w7840_
	);
	LUT2 #(
		.INIT('h2)
	) name5695 (
		\u7_mem_reg[2][18]/NET0131 ,
		_w7813_,
		_w7841_
	);
	LUT2 #(
		.INIT('h8)
	) name5696 (
		\u12_dout_reg[18]/P0001 ,
		_w7813_,
		_w7842_
	);
	LUT2 #(
		.INIT('h1)
	) name5697 (
		_w7841_,
		_w7842_,
		_w7843_
	);
	LUT2 #(
		.INIT('h2)
	) name5698 (
		\u7_mem_reg[2][19]/NET0131 ,
		_w7813_,
		_w7844_
	);
	LUT2 #(
		.INIT('h8)
	) name5699 (
		\u12_dout_reg[19]/P0001 ,
		_w7813_,
		_w7845_
	);
	LUT2 #(
		.INIT('h1)
	) name5700 (
		_w7844_,
		_w7845_,
		_w7846_
	);
	LUT2 #(
		.INIT('h2)
	) name5701 (
		\u7_mem_reg[2][1]/NET0131 ,
		_w7813_,
		_w7847_
	);
	LUT2 #(
		.INIT('h8)
	) name5702 (
		\u12_dout_reg[1]/P0001 ,
		_w7813_,
		_w7848_
	);
	LUT2 #(
		.INIT('h1)
	) name5703 (
		_w7847_,
		_w7848_,
		_w7849_
	);
	LUT2 #(
		.INIT('h2)
	) name5704 (
		\u7_mem_reg[2][20]/NET0131 ,
		_w7813_,
		_w7850_
	);
	LUT2 #(
		.INIT('h8)
	) name5705 (
		\u12_dout_reg[20]/P0001 ,
		_w7813_,
		_w7851_
	);
	LUT2 #(
		.INIT('h1)
	) name5706 (
		_w7850_,
		_w7851_,
		_w7852_
	);
	LUT2 #(
		.INIT('h2)
	) name5707 (
		\u7_mem_reg[2][21]/NET0131 ,
		_w7813_,
		_w7853_
	);
	LUT2 #(
		.INIT('h8)
	) name5708 (
		\u12_dout_reg[21]/P0001 ,
		_w7813_,
		_w7854_
	);
	LUT2 #(
		.INIT('h1)
	) name5709 (
		_w7853_,
		_w7854_,
		_w7855_
	);
	LUT2 #(
		.INIT('h2)
	) name5710 (
		\u7_mem_reg[2][22]/NET0131 ,
		_w7813_,
		_w7856_
	);
	LUT2 #(
		.INIT('h8)
	) name5711 (
		\u12_dout_reg[22]/P0001 ,
		_w7813_,
		_w7857_
	);
	LUT2 #(
		.INIT('h1)
	) name5712 (
		_w7856_,
		_w7857_,
		_w7858_
	);
	LUT2 #(
		.INIT('h2)
	) name5713 (
		\u7_mem_reg[2][23]/NET0131 ,
		_w7813_,
		_w7859_
	);
	LUT2 #(
		.INIT('h8)
	) name5714 (
		\u12_dout_reg[23]/P0001 ,
		_w7813_,
		_w7860_
	);
	LUT2 #(
		.INIT('h1)
	) name5715 (
		_w7859_,
		_w7860_,
		_w7861_
	);
	LUT2 #(
		.INIT('h2)
	) name5716 (
		\u7_mem_reg[2][24]/NET0131 ,
		_w7813_,
		_w7862_
	);
	LUT2 #(
		.INIT('h8)
	) name5717 (
		\u12_dout_reg[24]/P0001 ,
		_w7813_,
		_w7863_
	);
	LUT2 #(
		.INIT('h1)
	) name5718 (
		_w7862_,
		_w7863_,
		_w7864_
	);
	LUT2 #(
		.INIT('h2)
	) name5719 (
		\u7_mem_reg[2][25]/NET0131 ,
		_w7813_,
		_w7865_
	);
	LUT2 #(
		.INIT('h8)
	) name5720 (
		\u12_dout_reg[25]/P0001 ,
		_w7813_,
		_w7866_
	);
	LUT2 #(
		.INIT('h1)
	) name5721 (
		_w7865_,
		_w7866_,
		_w7867_
	);
	LUT2 #(
		.INIT('h2)
	) name5722 (
		\u7_mem_reg[2][26]/NET0131 ,
		_w7813_,
		_w7868_
	);
	LUT2 #(
		.INIT('h8)
	) name5723 (
		\u12_dout_reg[26]/P0001 ,
		_w7813_,
		_w7869_
	);
	LUT2 #(
		.INIT('h1)
	) name5724 (
		_w7868_,
		_w7869_,
		_w7870_
	);
	LUT2 #(
		.INIT('h2)
	) name5725 (
		\u7_mem_reg[2][27]/NET0131 ,
		_w7813_,
		_w7871_
	);
	LUT2 #(
		.INIT('h8)
	) name5726 (
		\u12_dout_reg[27]/P0001 ,
		_w7813_,
		_w7872_
	);
	LUT2 #(
		.INIT('h1)
	) name5727 (
		_w7871_,
		_w7872_,
		_w7873_
	);
	LUT2 #(
		.INIT('h2)
	) name5728 (
		\u7_mem_reg[2][28]/NET0131 ,
		_w7813_,
		_w7874_
	);
	LUT2 #(
		.INIT('h8)
	) name5729 (
		\u12_dout_reg[28]/P0001 ,
		_w7813_,
		_w7875_
	);
	LUT2 #(
		.INIT('h1)
	) name5730 (
		_w7874_,
		_w7875_,
		_w7876_
	);
	LUT2 #(
		.INIT('h2)
	) name5731 (
		\u7_mem_reg[2][29]/NET0131 ,
		_w7813_,
		_w7877_
	);
	LUT2 #(
		.INIT('h8)
	) name5732 (
		\u12_dout_reg[29]/P0001 ,
		_w7813_,
		_w7878_
	);
	LUT2 #(
		.INIT('h1)
	) name5733 (
		_w7877_,
		_w7878_,
		_w7879_
	);
	LUT2 #(
		.INIT('h2)
	) name5734 (
		\u7_mem_reg[2][2]/NET0131 ,
		_w7813_,
		_w7880_
	);
	LUT2 #(
		.INIT('h8)
	) name5735 (
		\u12_dout_reg[2]/P0001 ,
		_w7813_,
		_w7881_
	);
	LUT2 #(
		.INIT('h1)
	) name5736 (
		_w7880_,
		_w7881_,
		_w7882_
	);
	LUT2 #(
		.INIT('h2)
	) name5737 (
		\u7_mem_reg[2][30]/NET0131 ,
		_w7813_,
		_w7883_
	);
	LUT2 #(
		.INIT('h8)
	) name5738 (
		\u12_dout_reg[30]/P0001 ,
		_w7813_,
		_w7884_
	);
	LUT2 #(
		.INIT('h1)
	) name5739 (
		_w7883_,
		_w7884_,
		_w7885_
	);
	LUT2 #(
		.INIT('h2)
	) name5740 (
		\u7_mem_reg[2][31]/NET0131 ,
		_w7813_,
		_w7886_
	);
	LUT2 #(
		.INIT('h8)
	) name5741 (
		\u12_dout_reg[31]/P0001 ,
		_w7813_,
		_w7887_
	);
	LUT2 #(
		.INIT('h1)
	) name5742 (
		_w7886_,
		_w7887_,
		_w7888_
	);
	LUT2 #(
		.INIT('h2)
	) name5743 (
		\u7_mem_reg[2][3]/NET0131 ,
		_w7813_,
		_w7889_
	);
	LUT2 #(
		.INIT('h8)
	) name5744 (
		\u12_dout_reg[3]/P0001 ,
		_w7813_,
		_w7890_
	);
	LUT2 #(
		.INIT('h1)
	) name5745 (
		_w7889_,
		_w7890_,
		_w7891_
	);
	LUT2 #(
		.INIT('h2)
	) name5746 (
		\u7_mem_reg[2][4]/NET0131 ,
		_w7813_,
		_w7892_
	);
	LUT2 #(
		.INIT('h8)
	) name5747 (
		\u12_dout_reg[4]/P0001 ,
		_w7813_,
		_w7893_
	);
	LUT2 #(
		.INIT('h1)
	) name5748 (
		_w7892_,
		_w7893_,
		_w7894_
	);
	LUT2 #(
		.INIT('h2)
	) name5749 (
		\u7_mem_reg[2][5]/NET0131 ,
		_w7813_,
		_w7895_
	);
	LUT2 #(
		.INIT('h8)
	) name5750 (
		\u12_dout_reg[5]/P0001 ,
		_w7813_,
		_w7896_
	);
	LUT2 #(
		.INIT('h1)
	) name5751 (
		_w7895_,
		_w7896_,
		_w7897_
	);
	LUT2 #(
		.INIT('h2)
	) name5752 (
		\u7_mem_reg[2][6]/NET0131 ,
		_w7813_,
		_w7898_
	);
	LUT2 #(
		.INIT('h8)
	) name5753 (
		\u12_dout_reg[6]/P0001 ,
		_w7813_,
		_w7899_
	);
	LUT2 #(
		.INIT('h1)
	) name5754 (
		_w7898_,
		_w7899_,
		_w7900_
	);
	LUT2 #(
		.INIT('h2)
	) name5755 (
		\u7_mem_reg[2][7]/NET0131 ,
		_w7813_,
		_w7901_
	);
	LUT2 #(
		.INIT('h8)
	) name5756 (
		\u12_dout_reg[7]/P0001 ,
		_w7813_,
		_w7902_
	);
	LUT2 #(
		.INIT('h1)
	) name5757 (
		_w7901_,
		_w7902_,
		_w7903_
	);
	LUT2 #(
		.INIT('h2)
	) name5758 (
		\u7_mem_reg[2][8]/NET0131 ,
		_w7813_,
		_w7904_
	);
	LUT2 #(
		.INIT('h8)
	) name5759 (
		\u12_dout_reg[8]/P0001 ,
		_w7813_,
		_w7905_
	);
	LUT2 #(
		.INIT('h1)
	) name5760 (
		_w7904_,
		_w7905_,
		_w7906_
	);
	LUT2 #(
		.INIT('h2)
	) name5761 (
		\u7_mem_reg[2][9]/NET0131 ,
		_w7813_,
		_w7907_
	);
	LUT2 #(
		.INIT('h8)
	) name5762 (
		\u12_dout_reg[9]/P0001 ,
		_w7813_,
		_w7908_
	);
	LUT2 #(
		.INIT('h1)
	) name5763 (
		_w7907_,
		_w7908_,
		_w7909_
	);
	LUT2 #(
		.INIT('h2)
	) name5764 (
		\u7_mem_reg[3][0]/NET0131 ,
		_w6331_,
		_w7910_
	);
	LUT2 #(
		.INIT('h8)
	) name5765 (
		\u12_dout_reg[0]/P0001 ,
		_w6331_,
		_w7911_
	);
	LUT2 #(
		.INIT('h1)
	) name5766 (
		_w7910_,
		_w7911_,
		_w7912_
	);
	LUT2 #(
		.INIT('h2)
	) name5767 (
		\u7_mem_reg[3][10]/NET0131 ,
		_w6331_,
		_w7913_
	);
	LUT2 #(
		.INIT('h8)
	) name5768 (
		\u12_dout_reg[10]/P0001 ,
		_w6331_,
		_w7914_
	);
	LUT2 #(
		.INIT('h1)
	) name5769 (
		_w7913_,
		_w7914_,
		_w7915_
	);
	LUT2 #(
		.INIT('h2)
	) name5770 (
		\u7_mem_reg[3][11]/NET0131 ,
		_w6331_,
		_w7916_
	);
	LUT2 #(
		.INIT('h8)
	) name5771 (
		\u12_dout_reg[11]/P0001 ,
		_w6331_,
		_w7917_
	);
	LUT2 #(
		.INIT('h1)
	) name5772 (
		_w7916_,
		_w7917_,
		_w7918_
	);
	LUT2 #(
		.INIT('h2)
	) name5773 (
		\u7_mem_reg[3][12]/NET0131 ,
		_w6331_,
		_w7919_
	);
	LUT2 #(
		.INIT('h8)
	) name5774 (
		\u12_dout_reg[12]/P0001 ,
		_w6331_,
		_w7920_
	);
	LUT2 #(
		.INIT('h1)
	) name5775 (
		_w7919_,
		_w7920_,
		_w7921_
	);
	LUT2 #(
		.INIT('h2)
	) name5776 (
		\u7_mem_reg[3][13]/NET0131 ,
		_w6331_,
		_w7922_
	);
	LUT2 #(
		.INIT('h8)
	) name5777 (
		\u12_dout_reg[13]/P0001 ,
		_w6331_,
		_w7923_
	);
	LUT2 #(
		.INIT('h1)
	) name5778 (
		_w7922_,
		_w7923_,
		_w7924_
	);
	LUT2 #(
		.INIT('h2)
	) name5779 (
		\u7_mem_reg[3][14]/NET0131 ,
		_w6331_,
		_w7925_
	);
	LUT2 #(
		.INIT('h8)
	) name5780 (
		\u12_dout_reg[14]/P0001 ,
		_w6331_,
		_w7926_
	);
	LUT2 #(
		.INIT('h1)
	) name5781 (
		_w7925_,
		_w7926_,
		_w7927_
	);
	LUT2 #(
		.INIT('h2)
	) name5782 (
		\u7_mem_reg[3][15]/NET0131 ,
		_w6331_,
		_w7928_
	);
	LUT2 #(
		.INIT('h8)
	) name5783 (
		\u12_dout_reg[15]/P0001 ,
		_w6331_,
		_w7929_
	);
	LUT2 #(
		.INIT('h1)
	) name5784 (
		_w7928_,
		_w7929_,
		_w7930_
	);
	LUT2 #(
		.INIT('h2)
	) name5785 (
		\u7_mem_reg[3][16]/NET0131 ,
		_w6331_,
		_w7931_
	);
	LUT2 #(
		.INIT('h8)
	) name5786 (
		\u12_dout_reg[16]/P0001 ,
		_w6331_,
		_w7932_
	);
	LUT2 #(
		.INIT('h1)
	) name5787 (
		_w7931_,
		_w7932_,
		_w7933_
	);
	LUT2 #(
		.INIT('h2)
	) name5788 (
		\u7_mem_reg[3][17]/NET0131 ,
		_w6331_,
		_w7934_
	);
	LUT2 #(
		.INIT('h8)
	) name5789 (
		\u12_dout_reg[17]/P0001 ,
		_w6331_,
		_w7935_
	);
	LUT2 #(
		.INIT('h1)
	) name5790 (
		_w7934_,
		_w7935_,
		_w7936_
	);
	LUT2 #(
		.INIT('h2)
	) name5791 (
		\u7_mem_reg[3][18]/NET0131 ,
		_w6331_,
		_w7937_
	);
	LUT2 #(
		.INIT('h8)
	) name5792 (
		\u12_dout_reg[18]/P0001 ,
		_w6331_,
		_w7938_
	);
	LUT2 #(
		.INIT('h1)
	) name5793 (
		_w7937_,
		_w7938_,
		_w7939_
	);
	LUT2 #(
		.INIT('h2)
	) name5794 (
		\u7_mem_reg[3][19]/NET0131 ,
		_w6331_,
		_w7940_
	);
	LUT2 #(
		.INIT('h8)
	) name5795 (
		\u12_dout_reg[19]/P0001 ,
		_w6331_,
		_w7941_
	);
	LUT2 #(
		.INIT('h1)
	) name5796 (
		_w7940_,
		_w7941_,
		_w7942_
	);
	LUT2 #(
		.INIT('h2)
	) name5797 (
		\u7_mem_reg[3][1]/NET0131 ,
		_w6331_,
		_w7943_
	);
	LUT2 #(
		.INIT('h8)
	) name5798 (
		\u12_dout_reg[1]/P0001 ,
		_w6331_,
		_w7944_
	);
	LUT2 #(
		.INIT('h1)
	) name5799 (
		_w7943_,
		_w7944_,
		_w7945_
	);
	LUT2 #(
		.INIT('h2)
	) name5800 (
		\u7_mem_reg[3][20]/NET0131 ,
		_w6331_,
		_w7946_
	);
	LUT2 #(
		.INIT('h8)
	) name5801 (
		\u12_dout_reg[20]/P0001 ,
		_w6331_,
		_w7947_
	);
	LUT2 #(
		.INIT('h1)
	) name5802 (
		_w7946_,
		_w7947_,
		_w7948_
	);
	LUT2 #(
		.INIT('h2)
	) name5803 (
		\u7_mem_reg[3][21]/NET0131 ,
		_w6331_,
		_w7949_
	);
	LUT2 #(
		.INIT('h8)
	) name5804 (
		\u12_dout_reg[21]/P0001 ,
		_w6331_,
		_w7950_
	);
	LUT2 #(
		.INIT('h1)
	) name5805 (
		_w7949_,
		_w7950_,
		_w7951_
	);
	LUT2 #(
		.INIT('h2)
	) name5806 (
		\u7_mem_reg[3][22]/NET0131 ,
		_w6331_,
		_w7952_
	);
	LUT2 #(
		.INIT('h8)
	) name5807 (
		\u12_dout_reg[22]/P0001 ,
		_w6331_,
		_w7953_
	);
	LUT2 #(
		.INIT('h1)
	) name5808 (
		_w7952_,
		_w7953_,
		_w7954_
	);
	LUT2 #(
		.INIT('h2)
	) name5809 (
		\u7_mem_reg[3][23]/NET0131 ,
		_w6331_,
		_w7955_
	);
	LUT2 #(
		.INIT('h8)
	) name5810 (
		\u12_dout_reg[23]/P0001 ,
		_w6331_,
		_w7956_
	);
	LUT2 #(
		.INIT('h1)
	) name5811 (
		_w7955_,
		_w7956_,
		_w7957_
	);
	LUT2 #(
		.INIT('h2)
	) name5812 (
		\u7_mem_reg[3][24]/NET0131 ,
		_w6331_,
		_w7958_
	);
	LUT2 #(
		.INIT('h8)
	) name5813 (
		\u12_dout_reg[24]/P0001 ,
		_w6331_,
		_w7959_
	);
	LUT2 #(
		.INIT('h1)
	) name5814 (
		_w7958_,
		_w7959_,
		_w7960_
	);
	LUT2 #(
		.INIT('h2)
	) name5815 (
		\u7_mem_reg[3][25]/NET0131 ,
		_w6331_,
		_w7961_
	);
	LUT2 #(
		.INIT('h8)
	) name5816 (
		\u12_dout_reg[25]/P0001 ,
		_w6331_,
		_w7962_
	);
	LUT2 #(
		.INIT('h1)
	) name5817 (
		_w7961_,
		_w7962_,
		_w7963_
	);
	LUT2 #(
		.INIT('h2)
	) name5818 (
		\u7_mem_reg[3][26]/NET0131 ,
		_w6331_,
		_w7964_
	);
	LUT2 #(
		.INIT('h8)
	) name5819 (
		\u12_dout_reg[26]/P0001 ,
		_w6331_,
		_w7965_
	);
	LUT2 #(
		.INIT('h1)
	) name5820 (
		_w7964_,
		_w7965_,
		_w7966_
	);
	LUT2 #(
		.INIT('h2)
	) name5821 (
		\u7_mem_reg[3][27]/NET0131 ,
		_w6331_,
		_w7967_
	);
	LUT2 #(
		.INIT('h8)
	) name5822 (
		\u12_dout_reg[27]/P0001 ,
		_w6331_,
		_w7968_
	);
	LUT2 #(
		.INIT('h1)
	) name5823 (
		_w7967_,
		_w7968_,
		_w7969_
	);
	LUT2 #(
		.INIT('h2)
	) name5824 (
		\u7_mem_reg[3][28]/NET0131 ,
		_w6331_,
		_w7970_
	);
	LUT2 #(
		.INIT('h8)
	) name5825 (
		\u12_dout_reg[28]/P0001 ,
		_w6331_,
		_w7971_
	);
	LUT2 #(
		.INIT('h1)
	) name5826 (
		_w7970_,
		_w7971_,
		_w7972_
	);
	LUT2 #(
		.INIT('h2)
	) name5827 (
		\u7_mem_reg[3][29]/NET0131 ,
		_w6331_,
		_w7973_
	);
	LUT2 #(
		.INIT('h8)
	) name5828 (
		\u12_dout_reg[29]/P0001 ,
		_w6331_,
		_w7974_
	);
	LUT2 #(
		.INIT('h1)
	) name5829 (
		_w7973_,
		_w7974_,
		_w7975_
	);
	LUT2 #(
		.INIT('h2)
	) name5830 (
		\u7_mem_reg[3][2]/NET0131 ,
		_w6331_,
		_w7976_
	);
	LUT2 #(
		.INIT('h8)
	) name5831 (
		\u12_dout_reg[2]/P0001 ,
		_w6331_,
		_w7977_
	);
	LUT2 #(
		.INIT('h1)
	) name5832 (
		_w7976_,
		_w7977_,
		_w7978_
	);
	LUT2 #(
		.INIT('h2)
	) name5833 (
		\u7_mem_reg[3][30]/NET0131 ,
		_w6331_,
		_w7979_
	);
	LUT2 #(
		.INIT('h8)
	) name5834 (
		\u12_dout_reg[30]/P0001 ,
		_w6331_,
		_w7980_
	);
	LUT2 #(
		.INIT('h1)
	) name5835 (
		_w7979_,
		_w7980_,
		_w7981_
	);
	LUT2 #(
		.INIT('h2)
	) name5836 (
		\u7_mem_reg[3][31]/NET0131 ,
		_w6331_,
		_w7982_
	);
	LUT2 #(
		.INIT('h8)
	) name5837 (
		\u12_dout_reg[31]/P0001 ,
		_w6331_,
		_w7983_
	);
	LUT2 #(
		.INIT('h1)
	) name5838 (
		_w7982_,
		_w7983_,
		_w7984_
	);
	LUT2 #(
		.INIT('h2)
	) name5839 (
		\u7_mem_reg[3][3]/NET0131 ,
		_w6331_,
		_w7985_
	);
	LUT2 #(
		.INIT('h8)
	) name5840 (
		\u12_dout_reg[3]/P0001 ,
		_w6331_,
		_w7986_
	);
	LUT2 #(
		.INIT('h1)
	) name5841 (
		_w7985_,
		_w7986_,
		_w7987_
	);
	LUT2 #(
		.INIT('h2)
	) name5842 (
		\u7_mem_reg[3][4]/NET0131 ,
		_w6331_,
		_w7988_
	);
	LUT2 #(
		.INIT('h8)
	) name5843 (
		\u12_dout_reg[4]/P0001 ,
		_w6331_,
		_w7989_
	);
	LUT2 #(
		.INIT('h1)
	) name5844 (
		_w7988_,
		_w7989_,
		_w7990_
	);
	LUT2 #(
		.INIT('h2)
	) name5845 (
		\u7_mem_reg[3][5]/NET0131 ,
		_w6331_,
		_w7991_
	);
	LUT2 #(
		.INIT('h8)
	) name5846 (
		\u12_dout_reg[5]/P0001 ,
		_w6331_,
		_w7992_
	);
	LUT2 #(
		.INIT('h1)
	) name5847 (
		_w7991_,
		_w7992_,
		_w7993_
	);
	LUT2 #(
		.INIT('h2)
	) name5848 (
		\u7_mem_reg[3][6]/NET0131 ,
		_w6331_,
		_w7994_
	);
	LUT2 #(
		.INIT('h8)
	) name5849 (
		\u12_dout_reg[6]/P0001 ,
		_w6331_,
		_w7995_
	);
	LUT2 #(
		.INIT('h1)
	) name5850 (
		_w7994_,
		_w7995_,
		_w7996_
	);
	LUT2 #(
		.INIT('h2)
	) name5851 (
		\u7_mem_reg[3][7]/NET0131 ,
		_w6331_,
		_w7997_
	);
	LUT2 #(
		.INIT('h8)
	) name5852 (
		\u12_dout_reg[7]/P0001 ,
		_w6331_,
		_w7998_
	);
	LUT2 #(
		.INIT('h1)
	) name5853 (
		_w7997_,
		_w7998_,
		_w7999_
	);
	LUT2 #(
		.INIT('h2)
	) name5854 (
		\u7_mem_reg[3][8]/NET0131 ,
		_w6331_,
		_w8000_
	);
	LUT2 #(
		.INIT('h8)
	) name5855 (
		\u12_dout_reg[8]/P0001 ,
		_w6331_,
		_w8001_
	);
	LUT2 #(
		.INIT('h1)
	) name5856 (
		_w8000_,
		_w8001_,
		_w8002_
	);
	LUT2 #(
		.INIT('h2)
	) name5857 (
		\u7_mem_reg[3][9]/NET0131 ,
		_w6331_,
		_w8003_
	);
	LUT2 #(
		.INIT('h8)
	) name5858 (
		\u12_dout_reg[9]/P0001 ,
		_w6331_,
		_w8004_
	);
	LUT2 #(
		.INIT('h1)
	) name5859 (
		_w8003_,
		_w8004_,
		_w8005_
	);
	LUT2 #(
		.INIT('h2)
	) name5860 (
		\u3_mem_reg[2][17]/NET0131 ,
		_w6583_,
		_w8006_
	);
	LUT2 #(
		.INIT('h8)
	) name5861 (
		\u12_dout_reg[17]/P0001 ,
		_w6583_,
		_w8007_
	);
	LUT2 #(
		.INIT('h1)
	) name5862 (
		_w8006_,
		_w8007_,
		_w8008_
	);
	LUT2 #(
		.INIT('h2)
	) name5863 (
		\u8_mem_reg[1][0]/NET0131 ,
		_w6629_,
		_w8009_
	);
	LUT2 #(
		.INIT('h8)
	) name5864 (
		\u12_dout_reg[0]/P0001 ,
		_w6629_,
		_w8010_
	);
	LUT2 #(
		.INIT('h1)
	) name5865 (
		_w8009_,
		_w8010_,
		_w8011_
	);
	LUT2 #(
		.INIT('h2)
	) name5866 (
		\u8_mem_reg[1][10]/NET0131 ,
		_w6629_,
		_w8012_
	);
	LUT2 #(
		.INIT('h8)
	) name5867 (
		\u12_dout_reg[10]/P0001 ,
		_w6629_,
		_w8013_
	);
	LUT2 #(
		.INIT('h1)
	) name5868 (
		_w8012_,
		_w8013_,
		_w8014_
	);
	LUT2 #(
		.INIT('h2)
	) name5869 (
		\u8_mem_reg[1][11]/NET0131 ,
		_w6629_,
		_w8015_
	);
	LUT2 #(
		.INIT('h8)
	) name5870 (
		\u12_dout_reg[11]/P0001 ,
		_w6629_,
		_w8016_
	);
	LUT2 #(
		.INIT('h1)
	) name5871 (
		_w8015_,
		_w8016_,
		_w8017_
	);
	LUT2 #(
		.INIT('h2)
	) name5872 (
		\u8_mem_reg[1][12]/NET0131 ,
		_w6629_,
		_w8018_
	);
	LUT2 #(
		.INIT('h8)
	) name5873 (
		\u12_dout_reg[12]/P0001 ,
		_w6629_,
		_w8019_
	);
	LUT2 #(
		.INIT('h1)
	) name5874 (
		_w8018_,
		_w8019_,
		_w8020_
	);
	LUT2 #(
		.INIT('h2)
	) name5875 (
		\u8_mem_reg[1][13]/NET0131 ,
		_w6629_,
		_w8021_
	);
	LUT2 #(
		.INIT('h8)
	) name5876 (
		\u12_dout_reg[13]/P0001 ,
		_w6629_,
		_w8022_
	);
	LUT2 #(
		.INIT('h1)
	) name5877 (
		_w8021_,
		_w8022_,
		_w8023_
	);
	LUT2 #(
		.INIT('h2)
	) name5878 (
		\u8_mem_reg[1][14]/NET0131 ,
		_w6629_,
		_w8024_
	);
	LUT2 #(
		.INIT('h8)
	) name5879 (
		\u12_dout_reg[14]/P0001 ,
		_w6629_,
		_w8025_
	);
	LUT2 #(
		.INIT('h1)
	) name5880 (
		_w8024_,
		_w8025_,
		_w8026_
	);
	LUT2 #(
		.INIT('h2)
	) name5881 (
		\u8_mem_reg[1][15]/NET0131 ,
		_w6629_,
		_w8027_
	);
	LUT2 #(
		.INIT('h8)
	) name5882 (
		\u12_dout_reg[15]/P0001 ,
		_w6629_,
		_w8028_
	);
	LUT2 #(
		.INIT('h1)
	) name5883 (
		_w8027_,
		_w8028_,
		_w8029_
	);
	LUT2 #(
		.INIT('h2)
	) name5884 (
		\u8_mem_reg[1][16]/NET0131 ,
		_w6629_,
		_w8030_
	);
	LUT2 #(
		.INIT('h8)
	) name5885 (
		\u12_dout_reg[16]/P0001 ,
		_w6629_,
		_w8031_
	);
	LUT2 #(
		.INIT('h1)
	) name5886 (
		_w8030_,
		_w8031_,
		_w8032_
	);
	LUT2 #(
		.INIT('h2)
	) name5887 (
		\u8_mem_reg[1][17]/NET0131 ,
		_w6629_,
		_w8033_
	);
	LUT2 #(
		.INIT('h8)
	) name5888 (
		\u12_dout_reg[17]/P0001 ,
		_w6629_,
		_w8034_
	);
	LUT2 #(
		.INIT('h1)
	) name5889 (
		_w8033_,
		_w8034_,
		_w8035_
	);
	LUT2 #(
		.INIT('h2)
	) name5890 (
		\u8_mem_reg[1][18]/NET0131 ,
		_w6629_,
		_w8036_
	);
	LUT2 #(
		.INIT('h8)
	) name5891 (
		\u12_dout_reg[18]/P0001 ,
		_w6629_,
		_w8037_
	);
	LUT2 #(
		.INIT('h1)
	) name5892 (
		_w8036_,
		_w8037_,
		_w8038_
	);
	LUT2 #(
		.INIT('h2)
	) name5893 (
		\u8_mem_reg[1][19]/NET0131 ,
		_w6629_,
		_w8039_
	);
	LUT2 #(
		.INIT('h8)
	) name5894 (
		\u12_dout_reg[19]/P0001 ,
		_w6629_,
		_w8040_
	);
	LUT2 #(
		.INIT('h1)
	) name5895 (
		_w8039_,
		_w8040_,
		_w8041_
	);
	LUT2 #(
		.INIT('h2)
	) name5896 (
		\u8_mem_reg[1][1]/NET0131 ,
		_w6629_,
		_w8042_
	);
	LUT2 #(
		.INIT('h8)
	) name5897 (
		\u12_dout_reg[1]/P0001 ,
		_w6629_,
		_w8043_
	);
	LUT2 #(
		.INIT('h1)
	) name5898 (
		_w8042_,
		_w8043_,
		_w8044_
	);
	LUT2 #(
		.INIT('h2)
	) name5899 (
		\u8_mem_reg[1][20]/NET0131 ,
		_w6629_,
		_w8045_
	);
	LUT2 #(
		.INIT('h8)
	) name5900 (
		\u12_dout_reg[20]/P0001 ,
		_w6629_,
		_w8046_
	);
	LUT2 #(
		.INIT('h1)
	) name5901 (
		_w8045_,
		_w8046_,
		_w8047_
	);
	LUT2 #(
		.INIT('h2)
	) name5902 (
		\u8_mem_reg[1][21]/NET0131 ,
		_w6629_,
		_w8048_
	);
	LUT2 #(
		.INIT('h8)
	) name5903 (
		\u12_dout_reg[21]/P0001 ,
		_w6629_,
		_w8049_
	);
	LUT2 #(
		.INIT('h1)
	) name5904 (
		_w8048_,
		_w8049_,
		_w8050_
	);
	LUT2 #(
		.INIT('h2)
	) name5905 (
		\u8_mem_reg[1][22]/NET0131 ,
		_w6629_,
		_w8051_
	);
	LUT2 #(
		.INIT('h8)
	) name5906 (
		\u12_dout_reg[22]/P0001 ,
		_w6629_,
		_w8052_
	);
	LUT2 #(
		.INIT('h1)
	) name5907 (
		_w8051_,
		_w8052_,
		_w8053_
	);
	LUT2 #(
		.INIT('h2)
	) name5908 (
		\u8_mem_reg[1][23]/NET0131 ,
		_w6629_,
		_w8054_
	);
	LUT2 #(
		.INIT('h8)
	) name5909 (
		\u12_dout_reg[23]/P0001 ,
		_w6629_,
		_w8055_
	);
	LUT2 #(
		.INIT('h1)
	) name5910 (
		_w8054_,
		_w8055_,
		_w8056_
	);
	LUT2 #(
		.INIT('h2)
	) name5911 (
		\u8_mem_reg[1][24]/NET0131 ,
		_w6629_,
		_w8057_
	);
	LUT2 #(
		.INIT('h8)
	) name5912 (
		\u12_dout_reg[24]/P0001 ,
		_w6629_,
		_w8058_
	);
	LUT2 #(
		.INIT('h1)
	) name5913 (
		_w8057_,
		_w8058_,
		_w8059_
	);
	LUT2 #(
		.INIT('h2)
	) name5914 (
		\u8_mem_reg[1][25]/NET0131 ,
		_w6629_,
		_w8060_
	);
	LUT2 #(
		.INIT('h8)
	) name5915 (
		\u12_dout_reg[25]/P0001 ,
		_w6629_,
		_w8061_
	);
	LUT2 #(
		.INIT('h1)
	) name5916 (
		_w8060_,
		_w8061_,
		_w8062_
	);
	LUT2 #(
		.INIT('h2)
	) name5917 (
		\u3_mem_reg[1][0]/NET0131 ,
		_w6489_,
		_w8063_
	);
	LUT2 #(
		.INIT('h8)
	) name5918 (
		\u12_dout_reg[0]/P0001 ,
		_w6489_,
		_w8064_
	);
	LUT2 #(
		.INIT('h1)
	) name5919 (
		_w8063_,
		_w8064_,
		_w8065_
	);
	LUT2 #(
		.INIT('h2)
	) name5920 (
		\u8_mem_reg[1][26]/NET0131 ,
		_w6629_,
		_w8066_
	);
	LUT2 #(
		.INIT('h8)
	) name5921 (
		\u12_dout_reg[26]/P0001 ,
		_w6629_,
		_w8067_
	);
	LUT2 #(
		.INIT('h1)
	) name5922 (
		_w8066_,
		_w8067_,
		_w8068_
	);
	LUT2 #(
		.INIT('h2)
	) name5923 (
		\u8_mem_reg[1][27]/NET0131 ,
		_w6629_,
		_w8069_
	);
	LUT2 #(
		.INIT('h8)
	) name5924 (
		\u12_dout_reg[27]/P0001 ,
		_w6629_,
		_w8070_
	);
	LUT2 #(
		.INIT('h1)
	) name5925 (
		_w8069_,
		_w8070_,
		_w8071_
	);
	LUT2 #(
		.INIT('h2)
	) name5926 (
		\u3_mem_reg[1][10]/NET0131 ,
		_w6489_,
		_w8072_
	);
	LUT2 #(
		.INIT('h8)
	) name5927 (
		\u12_dout_reg[10]/P0001 ,
		_w6489_,
		_w8073_
	);
	LUT2 #(
		.INIT('h1)
	) name5928 (
		_w8072_,
		_w8073_,
		_w8074_
	);
	LUT2 #(
		.INIT('h2)
	) name5929 (
		\u8_mem_reg[1][29]/NET0131 ,
		_w6629_,
		_w8075_
	);
	LUT2 #(
		.INIT('h8)
	) name5930 (
		\u12_dout_reg[29]/P0001 ,
		_w6629_,
		_w8076_
	);
	LUT2 #(
		.INIT('h1)
	) name5931 (
		_w8075_,
		_w8076_,
		_w8077_
	);
	LUT2 #(
		.INIT('h2)
	) name5932 (
		\u3_mem_reg[1][11]/NET0131 ,
		_w6489_,
		_w8078_
	);
	LUT2 #(
		.INIT('h8)
	) name5933 (
		\u12_dout_reg[11]/P0001 ,
		_w6489_,
		_w8079_
	);
	LUT2 #(
		.INIT('h1)
	) name5934 (
		_w8078_,
		_w8079_,
		_w8080_
	);
	LUT2 #(
		.INIT('h2)
	) name5935 (
		\u8_mem_reg[1][2]/NET0131 ,
		_w6629_,
		_w8081_
	);
	LUT2 #(
		.INIT('h8)
	) name5936 (
		\u12_dout_reg[2]/P0001 ,
		_w6629_,
		_w8082_
	);
	LUT2 #(
		.INIT('h1)
	) name5937 (
		_w8081_,
		_w8082_,
		_w8083_
	);
	LUT2 #(
		.INIT('h2)
	) name5938 (
		\u8_mem_reg[1][30]/NET0131 ,
		_w6629_,
		_w8084_
	);
	LUT2 #(
		.INIT('h8)
	) name5939 (
		\u12_dout_reg[30]/P0001 ,
		_w6629_,
		_w8085_
	);
	LUT2 #(
		.INIT('h1)
	) name5940 (
		_w8084_,
		_w8085_,
		_w8086_
	);
	LUT2 #(
		.INIT('h2)
	) name5941 (
		\u3_mem_reg[1][12]/NET0131 ,
		_w6489_,
		_w8087_
	);
	LUT2 #(
		.INIT('h8)
	) name5942 (
		\u12_dout_reg[12]/P0001 ,
		_w6489_,
		_w8088_
	);
	LUT2 #(
		.INIT('h1)
	) name5943 (
		_w8087_,
		_w8088_,
		_w8089_
	);
	LUT2 #(
		.INIT('h2)
	) name5944 (
		\u8_mem_reg[3][11]/NET0131 ,
		_w6301_,
		_w8090_
	);
	LUT2 #(
		.INIT('h8)
	) name5945 (
		\u12_dout_reg[11]/P0001 ,
		_w6301_,
		_w8091_
	);
	LUT2 #(
		.INIT('h1)
	) name5946 (
		_w8090_,
		_w8091_,
		_w8092_
	);
	LUT2 #(
		.INIT('h2)
	) name5947 (
		\u8_mem_reg[1][3]/NET0131 ,
		_w6629_,
		_w8093_
	);
	LUT2 #(
		.INIT('h8)
	) name5948 (
		\u12_dout_reg[3]/P0001 ,
		_w6629_,
		_w8094_
	);
	LUT2 #(
		.INIT('h1)
	) name5949 (
		_w8093_,
		_w8094_,
		_w8095_
	);
	LUT2 #(
		.INIT('h2)
	) name5950 (
		\u3_mem_reg[1][13]/NET0131 ,
		_w6489_,
		_w8096_
	);
	LUT2 #(
		.INIT('h8)
	) name5951 (
		\u12_dout_reg[13]/P0001 ,
		_w6489_,
		_w8097_
	);
	LUT2 #(
		.INIT('h1)
	) name5952 (
		_w8096_,
		_w8097_,
		_w8098_
	);
	LUT2 #(
		.INIT('h2)
	) name5953 (
		\u8_mem_reg[1][5]/NET0131 ,
		_w6629_,
		_w8099_
	);
	LUT2 #(
		.INIT('h8)
	) name5954 (
		\u12_dout_reg[5]/P0001 ,
		_w6629_,
		_w8100_
	);
	LUT2 #(
		.INIT('h1)
	) name5955 (
		_w8099_,
		_w8100_,
		_w8101_
	);
	LUT2 #(
		.INIT('h2)
	) name5956 (
		\u8_mem_reg[1][7]/NET0131 ,
		_w6629_,
		_w8102_
	);
	LUT2 #(
		.INIT('h8)
	) name5957 (
		\u12_dout_reg[7]/P0001 ,
		_w6629_,
		_w8103_
	);
	LUT2 #(
		.INIT('h1)
	) name5958 (
		_w8102_,
		_w8103_,
		_w8104_
	);
	LUT2 #(
		.INIT('h2)
	) name5959 (
		\u3_mem_reg[1][15]/NET0131 ,
		_w6489_,
		_w8105_
	);
	LUT2 #(
		.INIT('h8)
	) name5960 (
		\u12_dout_reg[15]/P0001 ,
		_w6489_,
		_w8106_
	);
	LUT2 #(
		.INIT('h1)
	) name5961 (
		_w8105_,
		_w8106_,
		_w8107_
	);
	LUT2 #(
		.INIT('h2)
	) name5962 (
		\u8_mem_reg[1][8]/NET0131 ,
		_w6629_,
		_w8108_
	);
	LUT2 #(
		.INIT('h8)
	) name5963 (
		\u12_dout_reg[8]/P0001 ,
		_w6629_,
		_w8109_
	);
	LUT2 #(
		.INIT('h1)
	) name5964 (
		_w8108_,
		_w8109_,
		_w8110_
	);
	LUT2 #(
		.INIT('h2)
	) name5965 (
		\u8_mem_reg[1][9]/NET0131 ,
		_w6629_,
		_w8111_
	);
	LUT2 #(
		.INIT('h8)
	) name5966 (
		\u12_dout_reg[9]/P0001 ,
		_w6629_,
		_w8112_
	);
	LUT2 #(
		.INIT('h1)
	) name5967 (
		_w8111_,
		_w8112_,
		_w8113_
	);
	LUT2 #(
		.INIT('h2)
	) name5968 (
		\u3_mem_reg[1][16]/NET0131 ,
		_w6489_,
		_w8114_
	);
	LUT2 #(
		.INIT('h8)
	) name5969 (
		\u12_dout_reg[16]/P0001 ,
		_w6489_,
		_w8115_
	);
	LUT2 #(
		.INIT('h1)
	) name5970 (
		_w8114_,
		_w8115_,
		_w8116_
	);
	LUT2 #(
		.INIT('h2)
	) name5971 (
		\u8_mem_reg[2][0]/NET0131 ,
		_w6485_,
		_w8117_
	);
	LUT2 #(
		.INIT('h8)
	) name5972 (
		\u12_dout_reg[0]/P0001 ,
		_w6485_,
		_w8118_
	);
	LUT2 #(
		.INIT('h1)
	) name5973 (
		_w8117_,
		_w8118_,
		_w8119_
	);
	LUT2 #(
		.INIT('h2)
	) name5974 (
		\u8_mem_reg[2][10]/NET0131 ,
		_w6485_,
		_w8120_
	);
	LUT2 #(
		.INIT('h8)
	) name5975 (
		\u12_dout_reg[10]/P0001 ,
		_w6485_,
		_w8121_
	);
	LUT2 #(
		.INIT('h1)
	) name5976 (
		_w8120_,
		_w8121_,
		_w8122_
	);
	LUT2 #(
		.INIT('h2)
	) name5977 (
		\u3_mem_reg[1][17]/NET0131 ,
		_w6489_,
		_w8123_
	);
	LUT2 #(
		.INIT('h8)
	) name5978 (
		\u12_dout_reg[17]/P0001 ,
		_w6489_,
		_w8124_
	);
	LUT2 #(
		.INIT('h1)
	) name5979 (
		_w8123_,
		_w8124_,
		_w8125_
	);
	LUT2 #(
		.INIT('h2)
	) name5980 (
		\u8_mem_reg[2][11]/NET0131 ,
		_w6485_,
		_w8126_
	);
	LUT2 #(
		.INIT('h8)
	) name5981 (
		\u12_dout_reg[11]/P0001 ,
		_w6485_,
		_w8127_
	);
	LUT2 #(
		.INIT('h1)
	) name5982 (
		_w8126_,
		_w8127_,
		_w8128_
	);
	LUT2 #(
		.INIT('h2)
	) name5983 (
		\u8_mem_reg[2][12]/NET0131 ,
		_w6485_,
		_w8129_
	);
	LUT2 #(
		.INIT('h8)
	) name5984 (
		\u12_dout_reg[12]/P0001 ,
		_w6485_,
		_w8130_
	);
	LUT2 #(
		.INIT('h1)
	) name5985 (
		_w8129_,
		_w8130_,
		_w8131_
	);
	LUT2 #(
		.INIT('h2)
	) name5986 (
		\u3_mem_reg[1][18]/NET0131 ,
		_w6489_,
		_w8132_
	);
	LUT2 #(
		.INIT('h8)
	) name5987 (
		\u12_dout_reg[18]/P0001 ,
		_w6489_,
		_w8133_
	);
	LUT2 #(
		.INIT('h1)
	) name5988 (
		_w8132_,
		_w8133_,
		_w8134_
	);
	LUT2 #(
		.INIT('h2)
	) name5989 (
		\u8_mem_reg[2][13]/NET0131 ,
		_w6485_,
		_w8135_
	);
	LUT2 #(
		.INIT('h8)
	) name5990 (
		\u12_dout_reg[13]/P0001 ,
		_w6485_,
		_w8136_
	);
	LUT2 #(
		.INIT('h1)
	) name5991 (
		_w8135_,
		_w8136_,
		_w8137_
	);
	LUT2 #(
		.INIT('h2)
	) name5992 (
		\u8_mem_reg[2][14]/NET0131 ,
		_w6485_,
		_w8138_
	);
	LUT2 #(
		.INIT('h8)
	) name5993 (
		\u12_dout_reg[14]/P0001 ,
		_w6485_,
		_w8139_
	);
	LUT2 #(
		.INIT('h1)
	) name5994 (
		_w8138_,
		_w8139_,
		_w8140_
	);
	LUT2 #(
		.INIT('h2)
	) name5995 (
		\u3_mem_reg[1][19]/NET0131 ,
		_w6489_,
		_w8141_
	);
	LUT2 #(
		.INIT('h8)
	) name5996 (
		\u12_dout_reg[19]/P0001 ,
		_w6489_,
		_w8142_
	);
	LUT2 #(
		.INIT('h1)
	) name5997 (
		_w8141_,
		_w8142_,
		_w8143_
	);
	LUT2 #(
		.INIT('h2)
	) name5998 (
		\u8_mem_reg[2][15]/NET0131 ,
		_w6485_,
		_w8144_
	);
	LUT2 #(
		.INIT('h8)
	) name5999 (
		\u12_dout_reg[15]/P0001 ,
		_w6485_,
		_w8145_
	);
	LUT2 #(
		.INIT('h1)
	) name6000 (
		_w8144_,
		_w8145_,
		_w8146_
	);
	LUT2 #(
		.INIT('h2)
	) name6001 (
		\u8_mem_reg[2][16]/NET0131 ,
		_w6485_,
		_w8147_
	);
	LUT2 #(
		.INIT('h8)
	) name6002 (
		\u12_dout_reg[16]/P0001 ,
		_w6485_,
		_w8148_
	);
	LUT2 #(
		.INIT('h1)
	) name6003 (
		_w8147_,
		_w8148_,
		_w8149_
	);
	LUT2 #(
		.INIT('h2)
	) name6004 (
		\u8_mem_reg[2][17]/NET0131 ,
		_w6485_,
		_w8150_
	);
	LUT2 #(
		.INIT('h8)
	) name6005 (
		\u12_dout_reg[17]/P0001 ,
		_w6485_,
		_w8151_
	);
	LUT2 #(
		.INIT('h1)
	) name6006 (
		_w8150_,
		_w8151_,
		_w8152_
	);
	LUT2 #(
		.INIT('h2)
	) name6007 (
		\u8_mem_reg[2][18]/NET0131 ,
		_w6485_,
		_w8153_
	);
	LUT2 #(
		.INIT('h8)
	) name6008 (
		\u12_dout_reg[18]/P0001 ,
		_w6485_,
		_w8154_
	);
	LUT2 #(
		.INIT('h1)
	) name6009 (
		_w8153_,
		_w8154_,
		_w8155_
	);
	LUT2 #(
		.INIT('h2)
	) name6010 (
		\u3_mem_reg[1][20]/NET0131 ,
		_w6489_,
		_w8156_
	);
	LUT2 #(
		.INIT('h8)
	) name6011 (
		\u12_dout_reg[20]/P0001 ,
		_w6489_,
		_w8157_
	);
	LUT2 #(
		.INIT('h1)
	) name6012 (
		_w8156_,
		_w8157_,
		_w8158_
	);
	LUT2 #(
		.INIT('h2)
	) name6013 (
		\u8_mem_reg[2][19]/NET0131 ,
		_w6485_,
		_w8159_
	);
	LUT2 #(
		.INIT('h8)
	) name6014 (
		\u12_dout_reg[19]/P0001 ,
		_w6485_,
		_w8160_
	);
	LUT2 #(
		.INIT('h1)
	) name6015 (
		_w8159_,
		_w8160_,
		_w8161_
	);
	LUT2 #(
		.INIT('h2)
	) name6016 (
		\u8_mem_reg[2][1]/NET0131 ,
		_w6485_,
		_w8162_
	);
	LUT2 #(
		.INIT('h8)
	) name6017 (
		\u12_dout_reg[1]/P0001 ,
		_w6485_,
		_w8163_
	);
	LUT2 #(
		.INIT('h1)
	) name6018 (
		_w8162_,
		_w8163_,
		_w8164_
	);
	LUT2 #(
		.INIT('h2)
	) name6019 (
		\u3_mem_reg[1][21]/NET0131 ,
		_w6489_,
		_w8165_
	);
	LUT2 #(
		.INIT('h8)
	) name6020 (
		\u12_dout_reg[21]/P0001 ,
		_w6489_,
		_w8166_
	);
	LUT2 #(
		.INIT('h1)
	) name6021 (
		_w8165_,
		_w8166_,
		_w8167_
	);
	LUT2 #(
		.INIT('h2)
	) name6022 (
		\u8_mem_reg[2][20]/NET0131 ,
		_w6485_,
		_w8168_
	);
	LUT2 #(
		.INIT('h8)
	) name6023 (
		\u12_dout_reg[20]/P0001 ,
		_w6485_,
		_w8169_
	);
	LUT2 #(
		.INIT('h1)
	) name6024 (
		_w8168_,
		_w8169_,
		_w8170_
	);
	LUT2 #(
		.INIT('h2)
	) name6025 (
		\u8_mem_reg[2][21]/NET0131 ,
		_w6485_,
		_w8171_
	);
	LUT2 #(
		.INIT('h8)
	) name6026 (
		\u12_dout_reg[21]/P0001 ,
		_w6485_,
		_w8172_
	);
	LUT2 #(
		.INIT('h1)
	) name6027 (
		_w8171_,
		_w8172_,
		_w8173_
	);
	LUT2 #(
		.INIT('h2)
	) name6028 (
		\u3_mem_reg[1][22]/NET0131 ,
		_w6489_,
		_w8174_
	);
	LUT2 #(
		.INIT('h8)
	) name6029 (
		\u12_dout_reg[22]/P0001 ,
		_w6489_,
		_w8175_
	);
	LUT2 #(
		.INIT('h1)
	) name6030 (
		_w8174_,
		_w8175_,
		_w8176_
	);
	LUT2 #(
		.INIT('h2)
	) name6031 (
		\u8_mem_reg[2][22]/NET0131 ,
		_w6485_,
		_w8177_
	);
	LUT2 #(
		.INIT('h8)
	) name6032 (
		\u12_dout_reg[22]/P0001 ,
		_w6485_,
		_w8178_
	);
	LUT2 #(
		.INIT('h1)
	) name6033 (
		_w8177_,
		_w8178_,
		_w8179_
	);
	LUT2 #(
		.INIT('h2)
	) name6034 (
		\u8_mem_reg[2][23]/NET0131 ,
		_w6485_,
		_w8180_
	);
	LUT2 #(
		.INIT('h8)
	) name6035 (
		\u12_dout_reg[23]/P0001 ,
		_w6485_,
		_w8181_
	);
	LUT2 #(
		.INIT('h1)
	) name6036 (
		_w8180_,
		_w8181_,
		_w8182_
	);
	LUT2 #(
		.INIT('h2)
	) name6037 (
		\u8_mem_reg[2][24]/NET0131 ,
		_w6485_,
		_w8183_
	);
	LUT2 #(
		.INIT('h8)
	) name6038 (
		\u12_dout_reg[24]/P0001 ,
		_w6485_,
		_w8184_
	);
	LUT2 #(
		.INIT('h1)
	) name6039 (
		_w8183_,
		_w8184_,
		_w8185_
	);
	LUT2 #(
		.INIT('h2)
	) name6040 (
		\u8_mem_reg[2][25]/NET0131 ,
		_w6485_,
		_w8186_
	);
	LUT2 #(
		.INIT('h8)
	) name6041 (
		\u12_dout_reg[25]/P0001 ,
		_w6485_,
		_w8187_
	);
	LUT2 #(
		.INIT('h1)
	) name6042 (
		_w8186_,
		_w8187_,
		_w8188_
	);
	LUT2 #(
		.INIT('h2)
	) name6043 (
		\u3_mem_reg[1][24]/NET0131 ,
		_w6489_,
		_w8189_
	);
	LUT2 #(
		.INIT('h8)
	) name6044 (
		\u12_dout_reg[24]/P0001 ,
		_w6489_,
		_w8190_
	);
	LUT2 #(
		.INIT('h1)
	) name6045 (
		_w8189_,
		_w8190_,
		_w8191_
	);
	LUT2 #(
		.INIT('h2)
	) name6046 (
		\u8_mem_reg[2][26]/NET0131 ,
		_w6485_,
		_w8192_
	);
	LUT2 #(
		.INIT('h8)
	) name6047 (
		\u12_dout_reg[26]/P0001 ,
		_w6485_,
		_w8193_
	);
	LUT2 #(
		.INIT('h1)
	) name6048 (
		_w8192_,
		_w8193_,
		_w8194_
	);
	LUT2 #(
		.INIT('h2)
	) name6049 (
		\u8_mem_reg[2][27]/NET0131 ,
		_w6485_,
		_w8195_
	);
	LUT2 #(
		.INIT('h8)
	) name6050 (
		\u12_dout_reg[27]/P0001 ,
		_w6485_,
		_w8196_
	);
	LUT2 #(
		.INIT('h1)
	) name6051 (
		_w8195_,
		_w8196_,
		_w8197_
	);
	LUT2 #(
		.INIT('h2)
	) name6052 (
		\u3_mem_reg[1][25]/NET0131 ,
		_w6489_,
		_w8198_
	);
	LUT2 #(
		.INIT('h8)
	) name6053 (
		\u12_dout_reg[25]/P0001 ,
		_w6489_,
		_w8199_
	);
	LUT2 #(
		.INIT('h1)
	) name6054 (
		_w8198_,
		_w8199_,
		_w8200_
	);
	LUT2 #(
		.INIT('h2)
	) name6055 (
		\u8_mem_reg[2][28]/NET0131 ,
		_w6485_,
		_w8201_
	);
	LUT2 #(
		.INIT('h8)
	) name6056 (
		\u12_dout_reg[28]/P0001 ,
		_w6485_,
		_w8202_
	);
	LUT2 #(
		.INIT('h1)
	) name6057 (
		_w8201_,
		_w8202_,
		_w8203_
	);
	LUT2 #(
		.INIT('h2)
	) name6058 (
		\u8_mem_reg[2][29]/NET0131 ,
		_w6485_,
		_w8204_
	);
	LUT2 #(
		.INIT('h8)
	) name6059 (
		\u12_dout_reg[29]/P0001 ,
		_w6485_,
		_w8205_
	);
	LUT2 #(
		.INIT('h1)
	) name6060 (
		_w8204_,
		_w8205_,
		_w8206_
	);
	LUT2 #(
		.INIT('h2)
	) name6061 (
		\u3_mem_reg[1][26]/NET0131 ,
		_w6489_,
		_w8207_
	);
	LUT2 #(
		.INIT('h8)
	) name6062 (
		\u12_dout_reg[26]/P0001 ,
		_w6489_,
		_w8208_
	);
	LUT2 #(
		.INIT('h1)
	) name6063 (
		_w8207_,
		_w8208_,
		_w8209_
	);
	LUT2 #(
		.INIT('h2)
	) name6064 (
		\u8_mem_reg[2][2]/NET0131 ,
		_w6485_,
		_w8210_
	);
	LUT2 #(
		.INIT('h8)
	) name6065 (
		\u12_dout_reg[2]/P0001 ,
		_w6485_,
		_w8211_
	);
	LUT2 #(
		.INIT('h1)
	) name6066 (
		_w8210_,
		_w8211_,
		_w8212_
	);
	LUT2 #(
		.INIT('h2)
	) name6067 (
		\u8_mem_reg[2][30]/NET0131 ,
		_w6485_,
		_w8213_
	);
	LUT2 #(
		.INIT('h8)
	) name6068 (
		\u12_dout_reg[30]/P0001 ,
		_w6485_,
		_w8214_
	);
	LUT2 #(
		.INIT('h1)
	) name6069 (
		_w8213_,
		_w8214_,
		_w8215_
	);
	LUT2 #(
		.INIT('h2)
	) name6070 (
		\u8_mem_reg[2][31]/NET0131 ,
		_w6485_,
		_w8216_
	);
	LUT2 #(
		.INIT('h8)
	) name6071 (
		\u12_dout_reg[31]/P0001 ,
		_w6485_,
		_w8217_
	);
	LUT2 #(
		.INIT('h1)
	) name6072 (
		_w8216_,
		_w8217_,
		_w8218_
	);
	LUT2 #(
		.INIT('h2)
	) name6073 (
		\u3_mem_reg[1][28]/NET0131 ,
		_w6489_,
		_w8219_
	);
	LUT2 #(
		.INIT('h8)
	) name6074 (
		\u12_dout_reg[28]/P0001 ,
		_w6489_,
		_w8220_
	);
	LUT2 #(
		.INIT('h1)
	) name6075 (
		_w8219_,
		_w8220_,
		_w8221_
	);
	LUT2 #(
		.INIT('h2)
	) name6076 (
		\u8_mem_reg[2][4]/NET0131 ,
		_w6485_,
		_w8222_
	);
	LUT2 #(
		.INIT('h8)
	) name6077 (
		\u12_dout_reg[4]/P0001 ,
		_w6485_,
		_w8223_
	);
	LUT2 #(
		.INIT('h1)
	) name6078 (
		_w8222_,
		_w8223_,
		_w8224_
	);
	LUT2 #(
		.INIT('h4)
	) name6079 (
		\u3_wp_reg[1]/NET0131 ,
		_w6407_,
		_w8225_
	);
	LUT2 #(
		.INIT('h4)
	) name6080 (
		\u4_wp_reg[1]/NET0131 ,
		_w6411_,
		_w8226_
	);
	LUT2 #(
		.INIT('h4)
	) name6081 (
		\u5_wp_reg[1]/NET0131 ,
		_w6415_,
		_w8227_
	);
	LUT2 #(
		.INIT('h4)
	) name6082 (
		\u6_wp_reg[1]/NET0131 ,
		_w6419_,
		_w8228_
	);
	LUT2 #(
		.INIT('h4)
	) name6083 (
		\u7_wp_reg[1]/NET0131 ,
		_w6423_,
		_w8229_
	);
	LUT2 #(
		.INIT('h4)
	) name6084 (
		\u8_wp_reg[1]/NET0131 ,
		_w6403_,
		_w8230_
	);
	LUT2 #(
		.INIT('h8)
	) name6085 (
		\u13_ints_r_reg[0]/NET0131 ,
		_w2741_,
		_w8231_
	);
	LUT2 #(
		.INIT('h8)
	) name6086 (
		\u13_occ0_r_reg[0]/NET0131 ,
		_w6151_,
		_w8232_
	);
	LUT2 #(
		.INIT('h8)
	) name6087 (
		\u13_intm_r_reg[0]/NET0131 ,
		_w6153_,
		_w8233_
	);
	LUT2 #(
		.INIT('h8)
	) name6088 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w6157_,
		_w8234_
	);
	LUT2 #(
		.INIT('h8)
	) name6089 (
		\u13_occ1_r_reg[0]/NET0131 ,
		_w6147_,
		_w8235_
	);
	LUT2 #(
		.INIT('h8)
	) name6090 (
		\u15_crac_din_reg[0]/NET0131 ,
		_w6159_,
		_w8236_
	);
	LUT2 #(
		.INIT('h1)
	) name6091 (
		_w8231_,
		_w8232_,
		_w8237_
	);
	LUT2 #(
		.INIT('h1)
	) name6092 (
		_w8233_,
		_w8234_,
		_w8238_
	);
	LUT2 #(
		.INIT('h1)
	) name6093 (
		_w8235_,
		_w8236_,
		_w8239_
	);
	LUT2 #(
		.INIT('h8)
	) name6094 (
		_w8238_,
		_w8239_,
		_w8240_
	);
	LUT2 #(
		.INIT('h8)
	) name6095 (
		_w8237_,
		_w8240_,
		_w8241_
	);
	LUT2 #(
		.INIT('h2)
	) name6096 (
		_w6146_,
		_w8241_,
		_w8242_
	);
	LUT2 #(
		.INIT('h8)
	) name6097 (
		\u9_dout_reg[0]/P0001 ,
		_w6168_,
		_w8243_
	);
	LUT2 #(
		.INIT('h8)
	) name6098 (
		\u10_dout_reg[0]/P0001 ,
		_w6170_,
		_w8244_
	);
	LUT2 #(
		.INIT('h8)
	) name6099 (
		\u11_dout_reg[0]/P0001 ,
		_w6145_,
		_w8245_
	);
	LUT2 #(
		.INIT('h1)
	) name6100 (
		_w8243_,
		_w8244_,
		_w8246_
	);
	LUT2 #(
		.INIT('h4)
	) name6101 (
		_w8245_,
		_w8246_,
		_w8247_
	);
	LUT2 #(
		.INIT('h4)
	) name6102 (
		_w8242_,
		_w8247_,
		_w8248_
	);
	LUT2 #(
		.INIT('h8)
	) name6103 (
		\u13_ints_r_reg[10]/NET0131 ,
		_w2741_,
		_w8249_
	);
	LUT2 #(
		.INIT('h8)
	) name6104 (
		\u13_occ0_r_reg[10]/NET0131 ,
		_w6151_,
		_w8250_
	);
	LUT2 #(
		.INIT('h8)
	) name6105 (
		\u13_intm_r_reg[10]/NET0131 ,
		_w6153_,
		_w8251_
	);
	LUT2 #(
		.INIT('h8)
	) name6106 (
		\u13_icc_r_reg[10]/NET0131 ,
		_w6157_,
		_w8252_
	);
	LUT2 #(
		.INIT('h8)
	) name6107 (
		\u13_occ1_r_reg[10]/NET0131 ,
		_w6147_,
		_w8253_
	);
	LUT2 #(
		.INIT('h8)
	) name6108 (
		\u15_crac_din_reg[10]/NET0131 ,
		_w6159_,
		_w8254_
	);
	LUT2 #(
		.INIT('h1)
	) name6109 (
		_w8249_,
		_w8250_,
		_w8255_
	);
	LUT2 #(
		.INIT('h1)
	) name6110 (
		_w8251_,
		_w8252_,
		_w8256_
	);
	LUT2 #(
		.INIT('h1)
	) name6111 (
		_w8253_,
		_w8254_,
		_w8257_
	);
	LUT2 #(
		.INIT('h8)
	) name6112 (
		_w8256_,
		_w8257_,
		_w8258_
	);
	LUT2 #(
		.INIT('h8)
	) name6113 (
		_w8255_,
		_w8258_,
		_w8259_
	);
	LUT2 #(
		.INIT('h2)
	) name6114 (
		_w6146_,
		_w8259_,
		_w8260_
	);
	LUT2 #(
		.INIT('h8)
	) name6115 (
		\u9_dout_reg[10]/P0001 ,
		_w6168_,
		_w8261_
	);
	LUT2 #(
		.INIT('h8)
	) name6116 (
		\u10_dout_reg[10]/P0001 ,
		_w6170_,
		_w8262_
	);
	LUT2 #(
		.INIT('h8)
	) name6117 (
		\u11_dout_reg[10]/P0001 ,
		_w6145_,
		_w8263_
	);
	LUT2 #(
		.INIT('h1)
	) name6118 (
		_w8261_,
		_w8262_,
		_w8264_
	);
	LUT2 #(
		.INIT('h4)
	) name6119 (
		_w8263_,
		_w8264_,
		_w8265_
	);
	LUT2 #(
		.INIT('h4)
	) name6120 (
		_w8260_,
		_w8265_,
		_w8266_
	);
	LUT2 #(
		.INIT('h8)
	) name6121 (
		\u13_ints_r_reg[11]/NET0131 ,
		_w2741_,
		_w8267_
	);
	LUT2 #(
		.INIT('h8)
	) name6122 (
		\u13_occ0_r_reg[11]/NET0131 ,
		_w6151_,
		_w8268_
	);
	LUT2 #(
		.INIT('h8)
	) name6123 (
		\u13_intm_r_reg[11]/NET0131 ,
		_w6153_,
		_w8269_
	);
	LUT2 #(
		.INIT('h8)
	) name6124 (
		\u13_icc_r_reg[11]/NET0131 ,
		_w6157_,
		_w8270_
	);
	LUT2 #(
		.INIT('h8)
	) name6125 (
		\u13_occ1_r_reg[11]/NET0131 ,
		_w6147_,
		_w8271_
	);
	LUT2 #(
		.INIT('h8)
	) name6126 (
		\u15_crac_din_reg[11]/NET0131 ,
		_w6159_,
		_w8272_
	);
	LUT2 #(
		.INIT('h1)
	) name6127 (
		_w8267_,
		_w8268_,
		_w8273_
	);
	LUT2 #(
		.INIT('h1)
	) name6128 (
		_w8269_,
		_w8270_,
		_w8274_
	);
	LUT2 #(
		.INIT('h1)
	) name6129 (
		_w8271_,
		_w8272_,
		_w8275_
	);
	LUT2 #(
		.INIT('h8)
	) name6130 (
		_w8274_,
		_w8275_,
		_w8276_
	);
	LUT2 #(
		.INIT('h8)
	) name6131 (
		_w8273_,
		_w8276_,
		_w8277_
	);
	LUT2 #(
		.INIT('h2)
	) name6132 (
		_w6146_,
		_w8277_,
		_w8278_
	);
	LUT2 #(
		.INIT('h8)
	) name6133 (
		\u9_dout_reg[11]/P0001 ,
		_w6168_,
		_w8279_
	);
	LUT2 #(
		.INIT('h8)
	) name6134 (
		\u10_dout_reg[11]/P0001 ,
		_w6170_,
		_w8280_
	);
	LUT2 #(
		.INIT('h8)
	) name6135 (
		\u11_dout_reg[11]/P0001 ,
		_w6145_,
		_w8281_
	);
	LUT2 #(
		.INIT('h1)
	) name6136 (
		_w8279_,
		_w8280_,
		_w8282_
	);
	LUT2 #(
		.INIT('h4)
	) name6137 (
		_w8281_,
		_w8282_,
		_w8283_
	);
	LUT2 #(
		.INIT('h4)
	) name6138 (
		_w8278_,
		_w8283_,
		_w8284_
	);
	LUT2 #(
		.INIT('h8)
	) name6139 (
		\u13_ints_r_reg[12]/NET0131 ,
		_w2741_,
		_w8285_
	);
	LUT2 #(
		.INIT('h8)
	) name6140 (
		\u13_occ0_r_reg[12]/NET0131 ,
		_w6151_,
		_w8286_
	);
	LUT2 #(
		.INIT('h8)
	) name6141 (
		\u13_intm_r_reg[12]/NET0131 ,
		_w6153_,
		_w8287_
	);
	LUT2 #(
		.INIT('h8)
	) name6142 (
		\u13_icc_r_reg[12]/NET0131 ,
		_w6157_,
		_w8288_
	);
	LUT2 #(
		.INIT('h8)
	) name6143 (
		\u13_occ1_r_reg[12]/NET0131 ,
		_w6147_,
		_w8289_
	);
	LUT2 #(
		.INIT('h8)
	) name6144 (
		\u15_crac_din_reg[12]/NET0131 ,
		_w6159_,
		_w8290_
	);
	LUT2 #(
		.INIT('h1)
	) name6145 (
		_w8285_,
		_w8286_,
		_w8291_
	);
	LUT2 #(
		.INIT('h1)
	) name6146 (
		_w8287_,
		_w8288_,
		_w8292_
	);
	LUT2 #(
		.INIT('h1)
	) name6147 (
		_w8289_,
		_w8290_,
		_w8293_
	);
	LUT2 #(
		.INIT('h8)
	) name6148 (
		_w8292_,
		_w8293_,
		_w8294_
	);
	LUT2 #(
		.INIT('h8)
	) name6149 (
		_w8291_,
		_w8294_,
		_w8295_
	);
	LUT2 #(
		.INIT('h2)
	) name6150 (
		_w6146_,
		_w8295_,
		_w8296_
	);
	LUT2 #(
		.INIT('h8)
	) name6151 (
		\u9_dout_reg[12]/P0001 ,
		_w6168_,
		_w8297_
	);
	LUT2 #(
		.INIT('h8)
	) name6152 (
		\u10_dout_reg[12]/P0001 ,
		_w6170_,
		_w8298_
	);
	LUT2 #(
		.INIT('h8)
	) name6153 (
		\u11_dout_reg[12]/P0001 ,
		_w6145_,
		_w8299_
	);
	LUT2 #(
		.INIT('h1)
	) name6154 (
		_w8297_,
		_w8298_,
		_w8300_
	);
	LUT2 #(
		.INIT('h4)
	) name6155 (
		_w8299_,
		_w8300_,
		_w8301_
	);
	LUT2 #(
		.INIT('h4)
	) name6156 (
		_w8296_,
		_w8301_,
		_w8302_
	);
	LUT2 #(
		.INIT('h8)
	) name6157 (
		\u13_ints_r_reg[13]/NET0131 ,
		_w2741_,
		_w8303_
	);
	LUT2 #(
		.INIT('h8)
	) name6158 (
		\u13_occ0_r_reg[13]/NET0131 ,
		_w6151_,
		_w8304_
	);
	LUT2 #(
		.INIT('h8)
	) name6159 (
		\u13_intm_r_reg[13]/NET0131 ,
		_w6153_,
		_w8305_
	);
	LUT2 #(
		.INIT('h8)
	) name6160 (
		\u13_icc_r_reg[13]/NET0131 ,
		_w6157_,
		_w8306_
	);
	LUT2 #(
		.INIT('h8)
	) name6161 (
		\u13_occ1_r_reg[13]/NET0131 ,
		_w6147_,
		_w8307_
	);
	LUT2 #(
		.INIT('h8)
	) name6162 (
		\u15_crac_din_reg[13]/NET0131 ,
		_w6159_,
		_w8308_
	);
	LUT2 #(
		.INIT('h1)
	) name6163 (
		_w8303_,
		_w8304_,
		_w8309_
	);
	LUT2 #(
		.INIT('h1)
	) name6164 (
		_w8305_,
		_w8306_,
		_w8310_
	);
	LUT2 #(
		.INIT('h1)
	) name6165 (
		_w8307_,
		_w8308_,
		_w8311_
	);
	LUT2 #(
		.INIT('h8)
	) name6166 (
		_w8310_,
		_w8311_,
		_w8312_
	);
	LUT2 #(
		.INIT('h8)
	) name6167 (
		_w8309_,
		_w8312_,
		_w8313_
	);
	LUT2 #(
		.INIT('h2)
	) name6168 (
		_w6146_,
		_w8313_,
		_w8314_
	);
	LUT2 #(
		.INIT('h8)
	) name6169 (
		\u9_dout_reg[13]/P0001 ,
		_w6168_,
		_w8315_
	);
	LUT2 #(
		.INIT('h8)
	) name6170 (
		\u10_dout_reg[13]/P0001 ,
		_w6170_,
		_w8316_
	);
	LUT2 #(
		.INIT('h8)
	) name6171 (
		\u11_dout_reg[13]/P0001 ,
		_w6145_,
		_w8317_
	);
	LUT2 #(
		.INIT('h1)
	) name6172 (
		_w8315_,
		_w8316_,
		_w8318_
	);
	LUT2 #(
		.INIT('h4)
	) name6173 (
		_w8317_,
		_w8318_,
		_w8319_
	);
	LUT2 #(
		.INIT('h4)
	) name6174 (
		_w8314_,
		_w8319_,
		_w8320_
	);
	LUT2 #(
		.INIT('h8)
	) name6175 (
		\u13_ints_r_reg[14]/NET0131 ,
		_w2741_,
		_w8321_
	);
	LUT2 #(
		.INIT('h8)
	) name6176 (
		\u13_occ0_r_reg[14]/NET0131 ,
		_w6151_,
		_w8322_
	);
	LUT2 #(
		.INIT('h8)
	) name6177 (
		\u13_intm_r_reg[14]/NET0131 ,
		_w6153_,
		_w8323_
	);
	LUT2 #(
		.INIT('h8)
	) name6178 (
		\u13_icc_r_reg[14]/NET0131 ,
		_w6157_,
		_w8324_
	);
	LUT2 #(
		.INIT('h8)
	) name6179 (
		\u13_occ1_r_reg[14]/NET0131 ,
		_w6147_,
		_w8325_
	);
	LUT2 #(
		.INIT('h8)
	) name6180 (
		\u15_crac_din_reg[14]/NET0131 ,
		_w6159_,
		_w8326_
	);
	LUT2 #(
		.INIT('h1)
	) name6181 (
		_w8321_,
		_w8322_,
		_w8327_
	);
	LUT2 #(
		.INIT('h1)
	) name6182 (
		_w8323_,
		_w8324_,
		_w8328_
	);
	LUT2 #(
		.INIT('h1)
	) name6183 (
		_w8325_,
		_w8326_,
		_w8329_
	);
	LUT2 #(
		.INIT('h8)
	) name6184 (
		_w8328_,
		_w8329_,
		_w8330_
	);
	LUT2 #(
		.INIT('h8)
	) name6185 (
		_w8327_,
		_w8330_,
		_w8331_
	);
	LUT2 #(
		.INIT('h2)
	) name6186 (
		_w6146_,
		_w8331_,
		_w8332_
	);
	LUT2 #(
		.INIT('h8)
	) name6187 (
		\u9_dout_reg[14]/P0001 ,
		_w6168_,
		_w8333_
	);
	LUT2 #(
		.INIT('h8)
	) name6188 (
		\u10_dout_reg[14]/P0001 ,
		_w6170_,
		_w8334_
	);
	LUT2 #(
		.INIT('h8)
	) name6189 (
		\u11_dout_reg[14]/P0001 ,
		_w6145_,
		_w8335_
	);
	LUT2 #(
		.INIT('h1)
	) name6190 (
		_w8333_,
		_w8334_,
		_w8336_
	);
	LUT2 #(
		.INIT('h4)
	) name6191 (
		_w8335_,
		_w8336_,
		_w8337_
	);
	LUT2 #(
		.INIT('h4)
	) name6192 (
		_w8332_,
		_w8337_,
		_w8338_
	);
	LUT2 #(
		.INIT('h8)
	) name6193 (
		\u13_intm_r_reg[15]/NET0131 ,
		_w6153_,
		_w8339_
	);
	LUT2 #(
		.INIT('h8)
	) name6194 (
		\u13_occ1_r_reg[15]/NET0131 ,
		_w6147_,
		_w8340_
	);
	LUT2 #(
		.INIT('h8)
	) name6195 (
		\u13_occ0_r_reg[15]/NET0131 ,
		_w6151_,
		_w8341_
	);
	LUT2 #(
		.INIT('h8)
	) name6196 (
		\u13_icc_r_reg[15]/NET0131 ,
		_w6157_,
		_w8342_
	);
	LUT2 #(
		.INIT('h8)
	) name6197 (
		\u13_ints_r_reg[15]/NET0131 ,
		_w2741_,
		_w8343_
	);
	LUT2 #(
		.INIT('h8)
	) name6198 (
		\u15_crac_din_reg[15]/NET0131 ,
		_w6159_,
		_w8344_
	);
	LUT2 #(
		.INIT('h1)
	) name6199 (
		_w8339_,
		_w8340_,
		_w8345_
	);
	LUT2 #(
		.INIT('h1)
	) name6200 (
		_w8341_,
		_w8342_,
		_w8346_
	);
	LUT2 #(
		.INIT('h1)
	) name6201 (
		_w8343_,
		_w8344_,
		_w8347_
	);
	LUT2 #(
		.INIT('h8)
	) name6202 (
		_w8346_,
		_w8347_,
		_w8348_
	);
	LUT2 #(
		.INIT('h8)
	) name6203 (
		_w8345_,
		_w8348_,
		_w8349_
	);
	LUT2 #(
		.INIT('h2)
	) name6204 (
		_w6146_,
		_w8349_,
		_w8350_
	);
	LUT2 #(
		.INIT('h8)
	) name6205 (
		\u9_dout_reg[15]/P0001 ,
		_w6168_,
		_w8351_
	);
	LUT2 #(
		.INIT('h8)
	) name6206 (
		\u10_dout_reg[15]/P0001 ,
		_w6170_,
		_w8352_
	);
	LUT2 #(
		.INIT('h8)
	) name6207 (
		\u11_dout_reg[15]/P0001 ,
		_w6145_,
		_w8353_
	);
	LUT2 #(
		.INIT('h1)
	) name6208 (
		_w8351_,
		_w8352_,
		_w8354_
	);
	LUT2 #(
		.INIT('h4)
	) name6209 (
		_w8353_,
		_w8354_,
		_w8355_
	);
	LUT2 #(
		.INIT('h4)
	) name6210 (
		_w8350_,
		_w8355_,
		_w8356_
	);
	LUT2 #(
		.INIT('h8)
	) name6211 (
		\u13_ints_r_reg[2]/NET0131 ,
		_w2741_,
		_w8357_
	);
	LUT2 #(
		.INIT('h8)
	) name6212 (
		\u13_occ0_r_reg[2]/NET0131 ,
		_w6151_,
		_w8358_
	);
	LUT2 #(
		.INIT('h8)
	) name6213 (
		\u13_intm_r_reg[2]/NET0131 ,
		_w6153_,
		_w8359_
	);
	LUT2 #(
		.INIT('h8)
	) name6214 (
		\u13_icc_r_reg[2]/NET0131 ,
		_w6157_,
		_w8360_
	);
	LUT2 #(
		.INIT('h8)
	) name6215 (
		\u13_occ1_r_reg[2]/NET0131 ,
		_w6147_,
		_w8361_
	);
	LUT2 #(
		.INIT('h8)
	) name6216 (
		\u15_crac_din_reg[2]/NET0131 ,
		_w6159_,
		_w8362_
	);
	LUT2 #(
		.INIT('h1)
	) name6217 (
		_w8357_,
		_w8358_,
		_w8363_
	);
	LUT2 #(
		.INIT('h1)
	) name6218 (
		_w8359_,
		_w8360_,
		_w8364_
	);
	LUT2 #(
		.INIT('h1)
	) name6219 (
		_w8361_,
		_w8362_,
		_w8365_
	);
	LUT2 #(
		.INIT('h8)
	) name6220 (
		_w8364_,
		_w8365_,
		_w8366_
	);
	LUT2 #(
		.INIT('h8)
	) name6221 (
		_w8363_,
		_w8366_,
		_w8367_
	);
	LUT2 #(
		.INIT('h2)
	) name6222 (
		_w6146_,
		_w8367_,
		_w8368_
	);
	LUT2 #(
		.INIT('h8)
	) name6223 (
		\u9_dout_reg[2]/P0001 ,
		_w6168_,
		_w8369_
	);
	LUT2 #(
		.INIT('h8)
	) name6224 (
		\u10_dout_reg[2]/P0001 ,
		_w6170_,
		_w8370_
	);
	LUT2 #(
		.INIT('h8)
	) name6225 (
		\u11_dout_reg[2]/P0001 ,
		_w6145_,
		_w8371_
	);
	LUT2 #(
		.INIT('h1)
	) name6226 (
		_w8369_,
		_w8370_,
		_w8372_
	);
	LUT2 #(
		.INIT('h4)
	) name6227 (
		_w8371_,
		_w8372_,
		_w8373_
	);
	LUT2 #(
		.INIT('h4)
	) name6228 (
		_w8368_,
		_w8373_,
		_w8374_
	);
	LUT2 #(
		.INIT('h8)
	) name6229 (
		\u13_ints_r_reg[3]/NET0131 ,
		_w2741_,
		_w8375_
	);
	LUT2 #(
		.INIT('h8)
	) name6230 (
		\u13_occ0_r_reg[3]/NET0131 ,
		_w6151_,
		_w8376_
	);
	LUT2 #(
		.INIT('h8)
	) name6231 (
		\u13_intm_r_reg[3]/NET0131 ,
		_w6153_,
		_w8377_
	);
	LUT2 #(
		.INIT('h8)
	) name6232 (
		\u13_icc_r_reg[3]/NET0131 ,
		_w6157_,
		_w8378_
	);
	LUT2 #(
		.INIT('h8)
	) name6233 (
		\u13_occ1_r_reg[3]/NET0131 ,
		_w6147_,
		_w8379_
	);
	LUT2 #(
		.INIT('h8)
	) name6234 (
		\u15_crac_din_reg[3]/NET0131 ,
		_w6159_,
		_w8380_
	);
	LUT2 #(
		.INIT('h1)
	) name6235 (
		_w8375_,
		_w8376_,
		_w8381_
	);
	LUT2 #(
		.INIT('h1)
	) name6236 (
		_w8377_,
		_w8378_,
		_w8382_
	);
	LUT2 #(
		.INIT('h1)
	) name6237 (
		_w8379_,
		_w8380_,
		_w8383_
	);
	LUT2 #(
		.INIT('h8)
	) name6238 (
		_w8382_,
		_w8383_,
		_w8384_
	);
	LUT2 #(
		.INIT('h8)
	) name6239 (
		_w8381_,
		_w8384_,
		_w8385_
	);
	LUT2 #(
		.INIT('h2)
	) name6240 (
		_w6146_,
		_w8385_,
		_w8386_
	);
	LUT2 #(
		.INIT('h8)
	) name6241 (
		\u9_dout_reg[3]/P0001 ,
		_w6168_,
		_w8387_
	);
	LUT2 #(
		.INIT('h8)
	) name6242 (
		\u10_dout_reg[3]/P0001 ,
		_w6170_,
		_w8388_
	);
	LUT2 #(
		.INIT('h8)
	) name6243 (
		\u11_dout_reg[3]/P0001 ,
		_w6145_,
		_w8389_
	);
	LUT2 #(
		.INIT('h1)
	) name6244 (
		_w8387_,
		_w8388_,
		_w8390_
	);
	LUT2 #(
		.INIT('h4)
	) name6245 (
		_w8389_,
		_w8390_,
		_w8391_
	);
	LUT2 #(
		.INIT('h4)
	) name6246 (
		_w8386_,
		_w8391_,
		_w8392_
	);
	LUT2 #(
		.INIT('h8)
	) name6247 (
		\u13_ints_r_reg[4]/NET0131 ,
		_w2741_,
		_w8393_
	);
	LUT2 #(
		.INIT('h8)
	) name6248 (
		\u13_occ0_r_reg[4]/NET0131 ,
		_w6151_,
		_w8394_
	);
	LUT2 #(
		.INIT('h8)
	) name6249 (
		\u13_intm_r_reg[4]/NET0131 ,
		_w6153_,
		_w8395_
	);
	LUT2 #(
		.INIT('h8)
	) name6250 (
		\u13_icc_r_reg[4]/NET0131 ,
		_w6157_,
		_w8396_
	);
	LUT2 #(
		.INIT('h8)
	) name6251 (
		\u13_occ1_r_reg[4]/NET0131 ,
		_w6147_,
		_w8397_
	);
	LUT2 #(
		.INIT('h8)
	) name6252 (
		\u15_crac_din_reg[4]/NET0131 ,
		_w6159_,
		_w8398_
	);
	LUT2 #(
		.INIT('h1)
	) name6253 (
		_w8393_,
		_w8394_,
		_w8399_
	);
	LUT2 #(
		.INIT('h1)
	) name6254 (
		_w8395_,
		_w8396_,
		_w8400_
	);
	LUT2 #(
		.INIT('h1)
	) name6255 (
		_w8397_,
		_w8398_,
		_w8401_
	);
	LUT2 #(
		.INIT('h8)
	) name6256 (
		_w8400_,
		_w8401_,
		_w8402_
	);
	LUT2 #(
		.INIT('h8)
	) name6257 (
		_w8399_,
		_w8402_,
		_w8403_
	);
	LUT2 #(
		.INIT('h2)
	) name6258 (
		_w6146_,
		_w8403_,
		_w8404_
	);
	LUT2 #(
		.INIT('h8)
	) name6259 (
		\u9_dout_reg[4]/P0001 ,
		_w6168_,
		_w8405_
	);
	LUT2 #(
		.INIT('h8)
	) name6260 (
		\u10_dout_reg[4]/P0001 ,
		_w6170_,
		_w8406_
	);
	LUT2 #(
		.INIT('h8)
	) name6261 (
		\u11_dout_reg[4]/P0001 ,
		_w6145_,
		_w8407_
	);
	LUT2 #(
		.INIT('h1)
	) name6262 (
		_w8405_,
		_w8406_,
		_w8408_
	);
	LUT2 #(
		.INIT('h4)
	) name6263 (
		_w8407_,
		_w8408_,
		_w8409_
	);
	LUT2 #(
		.INIT('h4)
	) name6264 (
		_w8404_,
		_w8409_,
		_w8410_
	);
	LUT2 #(
		.INIT('h8)
	) name6265 (
		\u13_ints_r_reg[5]/NET0131 ,
		_w2741_,
		_w8411_
	);
	LUT2 #(
		.INIT('h8)
	) name6266 (
		\u13_occ0_r_reg[5]/NET0131 ,
		_w6151_,
		_w8412_
	);
	LUT2 #(
		.INIT('h8)
	) name6267 (
		\u13_intm_r_reg[5]/NET0131 ,
		_w6153_,
		_w8413_
	);
	LUT2 #(
		.INIT('h8)
	) name6268 (
		\u13_icc_r_reg[5]/NET0131 ,
		_w6157_,
		_w8414_
	);
	LUT2 #(
		.INIT('h8)
	) name6269 (
		\u13_occ1_r_reg[5]/NET0131 ,
		_w6147_,
		_w8415_
	);
	LUT2 #(
		.INIT('h8)
	) name6270 (
		\u15_crac_din_reg[5]/NET0131 ,
		_w6159_,
		_w8416_
	);
	LUT2 #(
		.INIT('h1)
	) name6271 (
		_w8411_,
		_w8412_,
		_w8417_
	);
	LUT2 #(
		.INIT('h1)
	) name6272 (
		_w8413_,
		_w8414_,
		_w8418_
	);
	LUT2 #(
		.INIT('h1)
	) name6273 (
		_w8415_,
		_w8416_,
		_w8419_
	);
	LUT2 #(
		.INIT('h8)
	) name6274 (
		_w8418_,
		_w8419_,
		_w8420_
	);
	LUT2 #(
		.INIT('h8)
	) name6275 (
		_w8417_,
		_w8420_,
		_w8421_
	);
	LUT2 #(
		.INIT('h2)
	) name6276 (
		_w6146_,
		_w8421_,
		_w8422_
	);
	LUT2 #(
		.INIT('h8)
	) name6277 (
		\u9_dout_reg[5]/P0001 ,
		_w6168_,
		_w8423_
	);
	LUT2 #(
		.INIT('h8)
	) name6278 (
		\u10_dout_reg[5]/P0001 ,
		_w6170_,
		_w8424_
	);
	LUT2 #(
		.INIT('h8)
	) name6279 (
		\u11_dout_reg[5]/P0001 ,
		_w6145_,
		_w8425_
	);
	LUT2 #(
		.INIT('h1)
	) name6280 (
		_w8423_,
		_w8424_,
		_w8426_
	);
	LUT2 #(
		.INIT('h4)
	) name6281 (
		_w8425_,
		_w8426_,
		_w8427_
	);
	LUT2 #(
		.INIT('h4)
	) name6282 (
		_w8422_,
		_w8427_,
		_w8428_
	);
	LUT2 #(
		.INIT('h8)
	) name6283 (
		\u13_ints_r_reg[6]/NET0131 ,
		_w2741_,
		_w8429_
	);
	LUT2 #(
		.INIT('h8)
	) name6284 (
		\u13_occ0_r_reg[6]/NET0131 ,
		_w6151_,
		_w8430_
	);
	LUT2 #(
		.INIT('h8)
	) name6285 (
		\u13_intm_r_reg[6]/NET0131 ,
		_w6153_,
		_w8431_
	);
	LUT2 #(
		.INIT('h8)
	) name6286 (
		\u13_icc_r_reg[6]/NET0131 ,
		_w6157_,
		_w8432_
	);
	LUT2 #(
		.INIT('h8)
	) name6287 (
		\u13_occ1_r_reg[6]/NET0131 ,
		_w6147_,
		_w8433_
	);
	LUT2 #(
		.INIT('h8)
	) name6288 (
		\u15_crac_din_reg[6]/NET0131 ,
		_w6159_,
		_w8434_
	);
	LUT2 #(
		.INIT('h1)
	) name6289 (
		_w8429_,
		_w8430_,
		_w8435_
	);
	LUT2 #(
		.INIT('h1)
	) name6290 (
		_w8431_,
		_w8432_,
		_w8436_
	);
	LUT2 #(
		.INIT('h1)
	) name6291 (
		_w8433_,
		_w8434_,
		_w8437_
	);
	LUT2 #(
		.INIT('h8)
	) name6292 (
		_w8436_,
		_w8437_,
		_w8438_
	);
	LUT2 #(
		.INIT('h8)
	) name6293 (
		_w8435_,
		_w8438_,
		_w8439_
	);
	LUT2 #(
		.INIT('h2)
	) name6294 (
		_w6146_,
		_w8439_,
		_w8440_
	);
	LUT2 #(
		.INIT('h8)
	) name6295 (
		\u9_dout_reg[6]/P0001 ,
		_w6168_,
		_w8441_
	);
	LUT2 #(
		.INIT('h8)
	) name6296 (
		\u10_dout_reg[6]/P0001 ,
		_w6170_,
		_w8442_
	);
	LUT2 #(
		.INIT('h8)
	) name6297 (
		\u11_dout_reg[6]/P0001 ,
		_w6145_,
		_w8443_
	);
	LUT2 #(
		.INIT('h1)
	) name6298 (
		_w8441_,
		_w8442_,
		_w8444_
	);
	LUT2 #(
		.INIT('h4)
	) name6299 (
		_w8443_,
		_w8444_,
		_w8445_
	);
	LUT2 #(
		.INIT('h4)
	) name6300 (
		_w8440_,
		_w8445_,
		_w8446_
	);
	LUT2 #(
		.INIT('h8)
	) name6301 (
		\u13_intm_r_reg[7]/NET0131 ,
		_w6153_,
		_w8447_
	);
	LUT2 #(
		.INIT('h8)
	) name6302 (
		\u13_occ1_r_reg[7]/NET0131 ,
		_w6147_,
		_w8448_
	);
	LUT2 #(
		.INIT('h8)
	) name6303 (
		\u13_occ0_r_reg[7]/NET0131 ,
		_w6151_,
		_w8449_
	);
	LUT2 #(
		.INIT('h8)
	) name6304 (
		\u13_icc_r_reg[7]/NET0131 ,
		_w6157_,
		_w8450_
	);
	LUT2 #(
		.INIT('h8)
	) name6305 (
		\u13_ints_r_reg[7]/NET0131 ,
		_w2741_,
		_w8451_
	);
	LUT2 #(
		.INIT('h8)
	) name6306 (
		\u15_crac_din_reg[7]/NET0131 ,
		_w6159_,
		_w8452_
	);
	LUT2 #(
		.INIT('h1)
	) name6307 (
		_w8447_,
		_w8448_,
		_w8453_
	);
	LUT2 #(
		.INIT('h1)
	) name6308 (
		_w8449_,
		_w8450_,
		_w8454_
	);
	LUT2 #(
		.INIT('h1)
	) name6309 (
		_w8451_,
		_w8452_,
		_w8455_
	);
	LUT2 #(
		.INIT('h8)
	) name6310 (
		_w8454_,
		_w8455_,
		_w8456_
	);
	LUT2 #(
		.INIT('h8)
	) name6311 (
		_w8453_,
		_w8456_,
		_w8457_
	);
	LUT2 #(
		.INIT('h2)
	) name6312 (
		_w6146_,
		_w8457_,
		_w8458_
	);
	LUT2 #(
		.INIT('h8)
	) name6313 (
		\u9_dout_reg[7]/P0001 ,
		_w6168_,
		_w8459_
	);
	LUT2 #(
		.INIT('h8)
	) name6314 (
		\u10_dout_reg[7]/P0001 ,
		_w6170_,
		_w8460_
	);
	LUT2 #(
		.INIT('h8)
	) name6315 (
		\u11_dout_reg[7]/P0001 ,
		_w6145_,
		_w8461_
	);
	LUT2 #(
		.INIT('h1)
	) name6316 (
		_w8459_,
		_w8460_,
		_w8462_
	);
	LUT2 #(
		.INIT('h4)
	) name6317 (
		_w8461_,
		_w8462_,
		_w8463_
	);
	LUT2 #(
		.INIT('h4)
	) name6318 (
		_w8458_,
		_w8463_,
		_w8464_
	);
	LUT2 #(
		.INIT('h8)
	) name6319 (
		\u13_ints_r_reg[8]/NET0131 ,
		_w2741_,
		_w8465_
	);
	LUT2 #(
		.INIT('h8)
	) name6320 (
		\u13_occ0_r_reg[8]/NET0131 ,
		_w6151_,
		_w8466_
	);
	LUT2 #(
		.INIT('h8)
	) name6321 (
		\u13_intm_r_reg[8]/NET0131 ,
		_w6153_,
		_w8467_
	);
	LUT2 #(
		.INIT('h8)
	) name6322 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w6157_,
		_w8468_
	);
	LUT2 #(
		.INIT('h8)
	) name6323 (
		\u13_occ1_r_reg[8]/NET0131 ,
		_w6147_,
		_w8469_
	);
	LUT2 #(
		.INIT('h8)
	) name6324 (
		\u15_crac_din_reg[8]/NET0131 ,
		_w6159_,
		_w8470_
	);
	LUT2 #(
		.INIT('h1)
	) name6325 (
		_w8465_,
		_w8466_,
		_w8471_
	);
	LUT2 #(
		.INIT('h1)
	) name6326 (
		_w8467_,
		_w8468_,
		_w8472_
	);
	LUT2 #(
		.INIT('h1)
	) name6327 (
		_w8469_,
		_w8470_,
		_w8473_
	);
	LUT2 #(
		.INIT('h8)
	) name6328 (
		_w8472_,
		_w8473_,
		_w8474_
	);
	LUT2 #(
		.INIT('h8)
	) name6329 (
		_w8471_,
		_w8474_,
		_w8475_
	);
	LUT2 #(
		.INIT('h2)
	) name6330 (
		_w6146_,
		_w8475_,
		_w8476_
	);
	LUT2 #(
		.INIT('h8)
	) name6331 (
		\u9_dout_reg[8]/P0001 ,
		_w6168_,
		_w8477_
	);
	LUT2 #(
		.INIT('h8)
	) name6332 (
		\u10_dout_reg[8]/P0001 ,
		_w6170_,
		_w8478_
	);
	LUT2 #(
		.INIT('h8)
	) name6333 (
		\u11_dout_reg[8]/P0001 ,
		_w6145_,
		_w8479_
	);
	LUT2 #(
		.INIT('h1)
	) name6334 (
		_w8477_,
		_w8478_,
		_w8480_
	);
	LUT2 #(
		.INIT('h4)
	) name6335 (
		_w8479_,
		_w8480_,
		_w8481_
	);
	LUT2 #(
		.INIT('h4)
	) name6336 (
		_w8476_,
		_w8481_,
		_w8482_
	);
	LUT2 #(
		.INIT('h8)
	) name6337 (
		\u13_ints_r_reg[9]/NET0131 ,
		_w2741_,
		_w8483_
	);
	LUT2 #(
		.INIT('h8)
	) name6338 (
		\u13_occ0_r_reg[9]/NET0131 ,
		_w6151_,
		_w8484_
	);
	LUT2 #(
		.INIT('h8)
	) name6339 (
		\u13_intm_r_reg[9]/NET0131 ,
		_w6153_,
		_w8485_
	);
	LUT2 #(
		.INIT('h8)
	) name6340 (
		\u13_icc_r_reg[9]/NET0131 ,
		_w6157_,
		_w8486_
	);
	LUT2 #(
		.INIT('h8)
	) name6341 (
		\u13_occ1_r_reg[9]/NET0131 ,
		_w6147_,
		_w8487_
	);
	LUT2 #(
		.INIT('h8)
	) name6342 (
		\u15_crac_din_reg[9]/NET0131 ,
		_w6159_,
		_w8488_
	);
	LUT2 #(
		.INIT('h1)
	) name6343 (
		_w8483_,
		_w8484_,
		_w8489_
	);
	LUT2 #(
		.INIT('h1)
	) name6344 (
		_w8485_,
		_w8486_,
		_w8490_
	);
	LUT2 #(
		.INIT('h1)
	) name6345 (
		_w8487_,
		_w8488_,
		_w8491_
	);
	LUT2 #(
		.INIT('h8)
	) name6346 (
		_w8490_,
		_w8491_,
		_w8492_
	);
	LUT2 #(
		.INIT('h8)
	) name6347 (
		_w8489_,
		_w8492_,
		_w8493_
	);
	LUT2 #(
		.INIT('h2)
	) name6348 (
		_w6146_,
		_w8493_,
		_w8494_
	);
	LUT2 #(
		.INIT('h8)
	) name6349 (
		\u9_dout_reg[9]/P0001 ,
		_w6168_,
		_w8495_
	);
	LUT2 #(
		.INIT('h8)
	) name6350 (
		\u10_dout_reg[9]/P0001 ,
		_w6170_,
		_w8496_
	);
	LUT2 #(
		.INIT('h8)
	) name6351 (
		\u11_dout_reg[9]/P0001 ,
		_w6145_,
		_w8497_
	);
	LUT2 #(
		.INIT('h1)
	) name6352 (
		_w8495_,
		_w8496_,
		_w8498_
	);
	LUT2 #(
		.INIT('h4)
	) name6353 (
		_w8497_,
		_w8498_,
		_w8499_
	);
	LUT2 #(
		.INIT('h4)
	) name6354 (
		_w8494_,
		_w8499_,
		_w8500_
	);
	LUT2 #(
		.INIT('h8)
	) name6355 (
		\u12_rf_we_reg/P0001 ,
		_w6159_,
		_w8501_
	);
	LUT2 #(
		.INIT('h8)
	) name6356 (
		\u12_rf_we_reg/P0001 ,
		_w6157_,
		_w8502_
	);
	LUT2 #(
		.INIT('h8)
	) name6357 (
		\u12_rf_we_reg/P0001 ,
		_w6153_,
		_w8503_
	);
	LUT2 #(
		.INIT('h8)
	) name6358 (
		\u12_rf_we_reg/P0001 ,
		_w6151_,
		_w8504_
	);
	LUT2 #(
		.INIT('h8)
	) name6359 (
		\u12_rf_we_reg/P0001 ,
		_w6147_,
		_w8505_
	);
	LUT2 #(
		.INIT('h1)
	) name6360 (
		\u2_cnt_reg[4]/NET0131 ,
		_w6471_,
		_w8506_
	);
	LUT2 #(
		.INIT('h1)
	) name6361 (
		_w6472_,
		_w8506_,
		_w8507_
	);
	LUT2 #(
		.INIT('h1)
	) name6362 (
		suspended_o_pad,
		_w8507_,
		_w8508_
	);
	LUT2 #(
		.INIT('h1)
	) name6363 (
		_w6235_,
		_w6236_,
		_w8509_
	);
	LUT2 #(
		.INIT('h1)
	) name6364 (
		\u4_rp_reg[0]/P0001 ,
		_w8509_,
		_w8510_
	);
	LUT2 #(
		.INIT('h2)
	) name6365 (
		_w2765_,
		_w6243_,
		_w8511_
	);
	LUT2 #(
		.INIT('h1)
	) name6366 (
		_w2760_,
		_w6240_,
		_w8512_
	);
	LUT2 #(
		.INIT('h4)
	) name6367 (
		_w8511_,
		_w8512_,
		_w8513_
	);
	LUT2 #(
		.INIT('h2)
	) name6368 (
		\u4_rp_reg[0]/P0001 ,
		_w8513_,
		_w8514_
	);
	LUT2 #(
		.INIT('h8)
	) name6369 (
		\u4_rp_reg[0]/P0001 ,
		_w2765_,
		_w8515_
	);
	LUT2 #(
		.INIT('h2)
	) name6370 (
		_w6243_,
		_w8515_,
		_w8516_
	);
	LUT2 #(
		.INIT('h1)
	) name6371 (
		_w6235_,
		_w6239_,
		_w8517_
	);
	LUT2 #(
		.INIT('h1)
	) name6372 (
		_w8510_,
		_w8516_,
		_w8518_
	);
	LUT2 #(
		.INIT('h4)
	) name6373 (
		_w8517_,
		_w8518_,
		_w8519_
	);
	LUT2 #(
		.INIT('h4)
	) name6374 (
		_w8514_,
		_w8519_,
		_w8520_
	);
	LUT2 #(
		.INIT('h1)
	) name6375 (
		_w6248_,
		_w6249_,
		_w8521_
	);
	LUT2 #(
		.INIT('h1)
	) name6376 (
		\u5_rp_reg[0]/P0001 ,
		_w8521_,
		_w8522_
	);
	LUT2 #(
		.INIT('h2)
	) name6377 (
		_w2776_,
		_w6256_,
		_w8523_
	);
	LUT2 #(
		.INIT('h1)
	) name6378 (
		_w2771_,
		_w6253_,
		_w8524_
	);
	LUT2 #(
		.INIT('h4)
	) name6379 (
		_w8523_,
		_w8524_,
		_w8525_
	);
	LUT2 #(
		.INIT('h2)
	) name6380 (
		\u5_rp_reg[0]/P0001 ,
		_w8525_,
		_w8526_
	);
	LUT2 #(
		.INIT('h8)
	) name6381 (
		\u5_rp_reg[0]/P0001 ,
		_w2776_,
		_w8527_
	);
	LUT2 #(
		.INIT('h2)
	) name6382 (
		_w6256_,
		_w8527_,
		_w8528_
	);
	LUT2 #(
		.INIT('h1)
	) name6383 (
		_w6248_,
		_w6252_,
		_w8529_
	);
	LUT2 #(
		.INIT('h1)
	) name6384 (
		_w8522_,
		_w8528_,
		_w8530_
	);
	LUT2 #(
		.INIT('h4)
	) name6385 (
		_w8529_,
		_w8530_,
		_w8531_
	);
	LUT2 #(
		.INIT('h4)
	) name6386 (
		_w8526_,
		_w8531_,
		_w8532_
	);
	LUT2 #(
		.INIT('h1)
	) name6387 (
		\u14_crac_wr_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w8533_
	);
	LUT2 #(
		.INIT('h1)
	) name6388 (
		_w6465_,
		_w8533_,
		_w8534_
	);
	LUT2 #(
		.INIT('h8)
	) name6389 (
		\u6_rp_reg[0]/P0001 ,
		_w2801_,
		_w8535_
	);
	LUT2 #(
		.INIT('h4)
	) name6390 (
		_w6270_,
		_w8535_,
		_w8536_
	);
	LUT2 #(
		.INIT('h8)
	) name6391 (
		_w6261_,
		_w6266_,
		_w8537_
	);
	LUT2 #(
		.INIT('h2)
	) name6392 (
		_w6262_,
		_w6266_,
		_w8538_
	);
	LUT2 #(
		.INIT('h1)
	) name6393 (
		_w8537_,
		_w8538_,
		_w8539_
	);
	LUT2 #(
		.INIT('h1)
	) name6394 (
		_w2796_,
		_w8539_,
		_w8540_
	);
	LUT2 #(
		.INIT('h2)
	) name6395 (
		\u6_rp_reg[0]/P0001 ,
		_w8540_,
		_w8541_
	);
	LUT2 #(
		.INIT('h1)
	) name6396 (
		\u6_rp_reg[0]/P0001 ,
		_w6267_,
		_w8542_
	);
	LUT2 #(
		.INIT('h2)
	) name6397 (
		_w6270_,
		_w8535_,
		_w8543_
	);
	LUT2 #(
		.INIT('h1)
	) name6398 (
		_w8536_,
		_w8543_,
		_w8544_
	);
	LUT2 #(
		.INIT('h4)
	) name6399 (
		_w8542_,
		_w8544_,
		_w8545_
	);
	LUT2 #(
		.INIT('h4)
	) name6400 (
		_w8541_,
		_w8545_,
		_w8546_
	);
	LUT2 #(
		.INIT('h8)
	) name6401 (
		\u7_rp_reg[0]/P0001 ,
		_w2981_,
		_w8547_
	);
	LUT2 #(
		.INIT('h1)
	) name6402 (
		_w6276_,
		_w8547_,
		_w8548_
	);
	LUT2 #(
		.INIT('h8)
	) name6403 (
		_w6276_,
		_w8547_,
		_w8549_
	);
	LUT2 #(
		.INIT('h1)
	) name6404 (
		_w8548_,
		_w8549_,
		_w8550_
	);
	LUT2 #(
		.INIT('h1)
	) name6405 (
		_w6277_,
		_w6282_,
		_w8551_
	);
	LUT2 #(
		.INIT('h8)
	) name6406 (
		\u7_rp_reg[1]/NET0131 ,
		_w6280_,
		_w8552_
	);
	LUT2 #(
		.INIT('h2)
	) name6407 (
		\u7_rp_reg[0]/P0001 ,
		_w8552_,
		_w8553_
	);
	LUT2 #(
		.INIT('h1)
	) name6408 (
		_w8551_,
		_w8553_,
		_w8554_
	);
	LUT2 #(
		.INIT('h1)
	) name6409 (
		_w2805_,
		_w8551_,
		_w8555_
	);
	LUT2 #(
		.INIT('h2)
	) name6410 (
		\u7_rp_reg[0]/P0001 ,
		_w8555_,
		_w8556_
	);
	LUT2 #(
		.INIT('h8)
	) name6411 (
		\u7_rp_reg[0]/P0001 ,
		\u7_rp_reg[1]/NET0131 ,
		_w8557_
	);
	LUT2 #(
		.INIT('h1)
	) name6412 (
		_w6280_,
		_w8557_,
		_w8558_
	);
	LUT2 #(
		.INIT('h1)
	) name6413 (
		_w8550_,
		_w8558_,
		_w8559_
	);
	LUT2 #(
		.INIT('h4)
	) name6414 (
		_w8556_,
		_w8559_,
		_w8560_
	);
	LUT2 #(
		.INIT('h4)
	) name6415 (
		_w8554_,
		_w8560_,
		_w8561_
	);
	LUT2 #(
		.INIT('h8)
	) name6416 (
		\u3_rp_reg[0]/P0001 ,
		_w3009_,
		_w8562_
	);
	LUT2 #(
		.INIT('h1)
	) name6417 (
		_w6224_,
		_w8562_,
		_w8563_
	);
	LUT2 #(
		.INIT('h8)
	) name6418 (
		_w6224_,
		_w8562_,
		_w8564_
	);
	LUT2 #(
		.INIT('h1)
	) name6419 (
		_w8563_,
		_w8564_,
		_w8565_
	);
	LUT2 #(
		.INIT('h1)
	) name6420 (
		_w6225_,
		_w6230_,
		_w8566_
	);
	LUT2 #(
		.INIT('h8)
	) name6421 (
		\u3_rp_reg[1]/NET0131 ,
		_w6228_,
		_w8567_
	);
	LUT2 #(
		.INIT('h2)
	) name6422 (
		\u3_rp_reg[0]/P0001 ,
		_w8567_,
		_w8568_
	);
	LUT2 #(
		.INIT('h1)
	) name6423 (
		_w8566_,
		_w8568_,
		_w8569_
	);
	LUT2 #(
		.INIT('h1)
	) name6424 (
		_w2784_,
		_w8566_,
		_w8570_
	);
	LUT2 #(
		.INIT('h2)
	) name6425 (
		\u3_rp_reg[0]/P0001 ,
		_w8570_,
		_w8571_
	);
	LUT2 #(
		.INIT('h8)
	) name6426 (
		\u3_rp_reg[0]/P0001 ,
		\u3_rp_reg[1]/NET0131 ,
		_w8572_
	);
	LUT2 #(
		.INIT('h1)
	) name6427 (
		_w6228_,
		_w8572_,
		_w8573_
	);
	LUT2 #(
		.INIT('h1)
	) name6428 (
		_w8565_,
		_w8573_,
		_w8574_
	);
	LUT2 #(
		.INIT('h4)
	) name6429 (
		_w8571_,
		_w8574_,
		_w8575_
	);
	LUT2 #(
		.INIT('h4)
	) name6430 (
		_w8569_,
		_w8575_,
		_w8576_
	);
	LUT2 #(
		.INIT('h8)
	) name6431 (
		\u8_rp_reg[0]/P0001 ,
		_w2163_,
		_w8577_
	);
	LUT2 #(
		.INIT('h4)
	) name6432 (
		_w6296_,
		_w8577_,
		_w8578_
	);
	LUT2 #(
		.INIT('h8)
	) name6433 (
		_w6287_,
		_w6292_,
		_w8579_
	);
	LUT2 #(
		.INIT('h2)
	) name6434 (
		_w6288_,
		_w6292_,
		_w8580_
	);
	LUT2 #(
		.INIT('h1)
	) name6435 (
		_w8579_,
		_w8580_,
		_w8581_
	);
	LUT2 #(
		.INIT('h1)
	) name6436 (
		_w2160_,
		_w8581_,
		_w8582_
	);
	LUT2 #(
		.INIT('h2)
	) name6437 (
		\u8_rp_reg[0]/P0001 ,
		_w8582_,
		_w8583_
	);
	LUT2 #(
		.INIT('h1)
	) name6438 (
		\u8_rp_reg[0]/P0001 ,
		_w6293_,
		_w8584_
	);
	LUT2 #(
		.INIT('h2)
	) name6439 (
		_w6296_,
		_w8577_,
		_w8585_
	);
	LUT2 #(
		.INIT('h1)
	) name6440 (
		_w8578_,
		_w8585_,
		_w8586_
	);
	LUT2 #(
		.INIT('h4)
	) name6441 (
		_w8584_,
		_w8586_,
		_w8587_
	);
	LUT2 #(
		.INIT('h4)
	) name6442 (
		_w8583_,
		_w8587_,
		_w8588_
	);
	LUT2 #(
		.INIT('h8)
	) name6443 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[1]/P0001 ,
		_w8589_
	);
	LUT2 #(
		.INIT('h2)
	) name6444 (
		\u0_slt9_r_reg[0]/P0001 ,
		\u2_ld_reg/P0001 ,
		_w8590_
	);
	LUT2 #(
		.INIT('h1)
	) name6445 (
		_w8589_,
		_w8590_,
		_w8591_
	);
	LUT2 #(
		.INIT('h8)
	) name6446 (
		\u12_i3_re_reg/NET0131 ,
		\u9_rp_reg[0]/P0001 ,
		_w8592_
	);
	LUT2 #(
		.INIT('h1)
	) name6447 (
		\u9_rp_reg[1]/P0001 ,
		_w8592_,
		_w8593_
	);
	LUT2 #(
		.INIT('h8)
	) name6448 (
		\u9_rp_reg[1]/P0001 ,
		_w8592_,
		_w8594_
	);
	LUT2 #(
		.INIT('h2)
	) name6449 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w8593_,
		_w8595_
	);
	LUT2 #(
		.INIT('h4)
	) name6450 (
		_w8594_,
		_w8595_,
		_w8596_
	);
	LUT2 #(
		.INIT('h8)
	) name6451 (
		\u10_rp_reg[0]/P0001 ,
		\u12_i4_re_reg/P0001 ,
		_w8597_
	);
	LUT2 #(
		.INIT('h1)
	) name6452 (
		\u10_rp_reg[1]/P0001 ,
		_w8597_,
		_w8598_
	);
	LUT2 #(
		.INIT('h8)
	) name6453 (
		\u10_rp_reg[1]/P0001 ,
		_w8597_,
		_w8599_
	);
	LUT2 #(
		.INIT('h2)
	) name6454 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w8598_,
		_w8600_
	);
	LUT2 #(
		.INIT('h4)
	) name6455 (
		_w8599_,
		_w8600_,
		_w8601_
	);
	LUT2 #(
		.INIT('h8)
	) name6456 (
		\u11_rp_reg[0]/P0001 ,
		\u12_i6_re_reg/NET0131 ,
		_w8602_
	);
	LUT2 #(
		.INIT('h1)
	) name6457 (
		\u11_rp_reg[1]/P0001 ,
		_w8602_,
		_w8603_
	);
	LUT2 #(
		.INIT('h8)
	) name6458 (
		\u11_rp_reg[1]/P0001 ,
		_w8602_,
		_w8604_
	);
	LUT2 #(
		.INIT('h2)
	) name6459 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w8603_,
		_w8605_
	);
	LUT2 #(
		.INIT('h4)
	) name6460 (
		_w8604_,
		_w8605_,
		_w8606_
	);
	LUT2 #(
		.INIT('h1)
	) name6461 (
		\u9_rp_reg[2]/P0001 ,
		_w8594_,
		_w8607_
	);
	LUT2 #(
		.INIT('h8)
	) name6462 (
		\u9_rp_reg[2]/P0001 ,
		_w8594_,
		_w8608_
	);
	LUT2 #(
		.INIT('h2)
	) name6463 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w8607_,
		_w8609_
	);
	LUT2 #(
		.INIT('h4)
	) name6464 (
		_w8608_,
		_w8609_,
		_w8610_
	);
	LUT2 #(
		.INIT('h1)
	) name6465 (
		\u11_rp_reg[2]/P0001 ,
		_w8604_,
		_w8611_
	);
	LUT2 #(
		.INIT('h8)
	) name6466 (
		\u11_rp_reg[2]/P0001 ,
		_w8604_,
		_w8612_
	);
	LUT2 #(
		.INIT('h2)
	) name6467 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w8611_,
		_w8613_
	);
	LUT2 #(
		.INIT('h4)
	) name6468 (
		_w8612_,
		_w8613_,
		_w8614_
	);
	LUT2 #(
		.INIT('h1)
	) name6469 (
		\u10_rp_reg[2]/P0001 ,
		_w8599_,
		_w8615_
	);
	LUT2 #(
		.INIT('h8)
	) name6470 (
		\u10_rp_reg[2]/P0001 ,
		_w8599_,
		_w8616_
	);
	LUT2 #(
		.INIT('h2)
	) name6471 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w8615_,
		_w8617_
	);
	LUT2 #(
		.INIT('h4)
	) name6472 (
		_w8616_,
		_w8617_,
		_w8618_
	);
	LUT2 #(
		.INIT('h1)
	) name6473 (
		\u2_res_cnt_reg[2]/P0001 ,
		_w6455_,
		_w8619_
	);
	LUT2 #(
		.INIT('h2)
	) name6474 (
		\u2_sync_resume_reg/NET0131 ,
		_w6456_,
		_w8620_
	);
	LUT2 #(
		.INIT('h4)
	) name6475 (
		_w8619_,
		_w8620_,
		_w8621_
	);
	LUT2 #(
		.INIT('h1)
	) name6476 (
		\u11_rp_reg[0]/P0001 ,
		\u12_i6_re_reg/NET0131 ,
		_w8622_
	);
	LUT2 #(
		.INIT('h2)
	) name6477 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w8602_,
		_w8623_
	);
	LUT2 #(
		.INIT('h4)
	) name6478 (
		_w8622_,
		_w8623_,
		_w8624_
	);
	LUT2 #(
		.INIT('h8)
	) name6479 (
		\u13_crac_r_reg[0]/NET0131 ,
		_w6159_,
		_w8625_
	);
	LUT2 #(
		.INIT('h8)
	) name6480 (
		\u13_intm_r_reg[16]/NET0131 ,
		_w6153_,
		_w8626_
	);
	LUT2 #(
		.INIT('h8)
	) name6481 (
		\u13_icc_r_reg[16]/NET0131 ,
		_w6157_,
		_w8627_
	);
	LUT2 #(
		.INIT('h8)
	) name6482 (
		\u13_occ0_r_reg[16]/NET0131 ,
		_w6151_,
		_w8628_
	);
	LUT2 #(
		.INIT('h8)
	) name6483 (
		\u13_ints_r_reg[16]/NET0131 ,
		_w2741_,
		_w8629_
	);
	LUT2 #(
		.INIT('h1)
	) name6484 (
		_w8625_,
		_w8626_,
		_w8630_
	);
	LUT2 #(
		.INIT('h1)
	) name6485 (
		_w8627_,
		_w8628_,
		_w8631_
	);
	LUT2 #(
		.INIT('h4)
	) name6486 (
		_w8629_,
		_w8631_,
		_w8632_
	);
	LUT2 #(
		.INIT('h8)
	) name6487 (
		_w8630_,
		_w8632_,
		_w8633_
	);
	LUT2 #(
		.INIT('h2)
	) name6488 (
		_w6146_,
		_w8633_,
		_w8634_
	);
	LUT2 #(
		.INIT('h8)
	) name6489 (
		\u9_dout_reg[16]/P0001 ,
		_w6168_,
		_w8635_
	);
	LUT2 #(
		.INIT('h8)
	) name6490 (
		\u10_dout_reg[16]/P0001 ,
		_w6170_,
		_w8636_
	);
	LUT2 #(
		.INIT('h8)
	) name6491 (
		\u11_dout_reg[16]/P0001 ,
		_w6145_,
		_w8637_
	);
	LUT2 #(
		.INIT('h1)
	) name6492 (
		_w8635_,
		_w8636_,
		_w8638_
	);
	LUT2 #(
		.INIT('h4)
	) name6493 (
		_w8637_,
		_w8638_,
		_w8639_
	);
	LUT2 #(
		.INIT('h4)
	) name6494 (
		_w8634_,
		_w8639_,
		_w8640_
	);
	LUT2 #(
		.INIT('h8)
	) name6495 (
		\u13_icc_r_reg[17]/NET0131 ,
		_w6157_,
		_w8641_
	);
	LUT2 #(
		.INIT('h8)
	) name6496 (
		\u13_intm_r_reg[17]/NET0131 ,
		_w6153_,
		_w8642_
	);
	LUT2 #(
		.INIT('h8)
	) name6497 (
		\u13_crac_r_reg[1]/NET0131 ,
		_w6159_,
		_w8643_
	);
	LUT2 #(
		.INIT('h8)
	) name6498 (
		\u13_occ0_r_reg[17]/NET0131 ,
		_w6151_,
		_w8644_
	);
	LUT2 #(
		.INIT('h8)
	) name6499 (
		\u13_ints_r_reg[17]/NET0131 ,
		_w2741_,
		_w8645_
	);
	LUT2 #(
		.INIT('h1)
	) name6500 (
		_w8641_,
		_w8642_,
		_w8646_
	);
	LUT2 #(
		.INIT('h1)
	) name6501 (
		_w8643_,
		_w8644_,
		_w8647_
	);
	LUT2 #(
		.INIT('h4)
	) name6502 (
		_w8645_,
		_w8647_,
		_w8648_
	);
	LUT2 #(
		.INIT('h8)
	) name6503 (
		_w8646_,
		_w8648_,
		_w8649_
	);
	LUT2 #(
		.INIT('h2)
	) name6504 (
		_w6146_,
		_w8649_,
		_w8650_
	);
	LUT2 #(
		.INIT('h8)
	) name6505 (
		\u9_dout_reg[17]/P0001 ,
		_w6168_,
		_w8651_
	);
	LUT2 #(
		.INIT('h8)
	) name6506 (
		\u10_dout_reg[17]/P0001 ,
		_w6170_,
		_w8652_
	);
	LUT2 #(
		.INIT('h8)
	) name6507 (
		\u11_dout_reg[17]/P0001 ,
		_w6145_,
		_w8653_
	);
	LUT2 #(
		.INIT('h1)
	) name6508 (
		_w8651_,
		_w8652_,
		_w8654_
	);
	LUT2 #(
		.INIT('h4)
	) name6509 (
		_w8653_,
		_w8654_,
		_w8655_
	);
	LUT2 #(
		.INIT('h4)
	) name6510 (
		_w8650_,
		_w8655_,
		_w8656_
	);
	LUT2 #(
		.INIT('h8)
	) name6511 (
		\u13_crac_r_reg[3]/NET0131 ,
		_w6159_,
		_w8657_
	);
	LUT2 #(
		.INIT('h8)
	) name6512 (
		\u13_intm_r_reg[19]/NET0131 ,
		_w6153_,
		_w8658_
	);
	LUT2 #(
		.INIT('h8)
	) name6513 (
		\u13_icc_r_reg[19]/NET0131 ,
		_w6157_,
		_w8659_
	);
	LUT2 #(
		.INIT('h8)
	) name6514 (
		\u13_occ0_r_reg[19]/NET0131 ,
		_w6151_,
		_w8660_
	);
	LUT2 #(
		.INIT('h8)
	) name6515 (
		\u13_ints_r_reg[19]/NET0131 ,
		_w2741_,
		_w8661_
	);
	LUT2 #(
		.INIT('h1)
	) name6516 (
		_w8657_,
		_w8658_,
		_w8662_
	);
	LUT2 #(
		.INIT('h1)
	) name6517 (
		_w8659_,
		_w8660_,
		_w8663_
	);
	LUT2 #(
		.INIT('h4)
	) name6518 (
		_w8661_,
		_w8663_,
		_w8664_
	);
	LUT2 #(
		.INIT('h8)
	) name6519 (
		_w8662_,
		_w8664_,
		_w8665_
	);
	LUT2 #(
		.INIT('h2)
	) name6520 (
		_w6146_,
		_w8665_,
		_w8666_
	);
	LUT2 #(
		.INIT('h8)
	) name6521 (
		\u9_dout_reg[19]/P0001 ,
		_w6168_,
		_w8667_
	);
	LUT2 #(
		.INIT('h8)
	) name6522 (
		\u10_dout_reg[19]/P0001 ,
		_w6170_,
		_w8668_
	);
	LUT2 #(
		.INIT('h8)
	) name6523 (
		\u11_dout_reg[19]/P0001 ,
		_w6145_,
		_w8669_
	);
	LUT2 #(
		.INIT('h1)
	) name6524 (
		_w8667_,
		_w8668_,
		_w8670_
	);
	LUT2 #(
		.INIT('h4)
	) name6525 (
		_w8669_,
		_w8670_,
		_w8671_
	);
	LUT2 #(
		.INIT('h4)
	) name6526 (
		_w8666_,
		_w8671_,
		_w8672_
	);
	LUT2 #(
		.INIT('h1)
	) name6527 (
		\u12_i3_re_reg/NET0131 ,
		\u9_rp_reg[0]/P0001 ,
		_w8673_
	);
	LUT2 #(
		.INIT('h2)
	) name6528 (
		\u13_icc_r_reg[0]/NET0131 ,
		_w8592_,
		_w8674_
	);
	LUT2 #(
		.INIT('h4)
	) name6529 (
		_w8673_,
		_w8674_,
		_w8675_
	);
	LUT2 #(
		.INIT('h8)
	) name6530 (
		\u13_icc_r_reg[20]/NET0131 ,
		_w6157_,
		_w8676_
	);
	LUT2 #(
		.INIT('h8)
	) name6531 (
		\u13_intm_r_reg[20]/NET0131 ,
		_w6153_,
		_w8677_
	);
	LUT2 #(
		.INIT('h8)
	) name6532 (
		\u13_crac_r_reg[4]/NET0131 ,
		_w6159_,
		_w8678_
	);
	LUT2 #(
		.INIT('h8)
	) name6533 (
		\u13_occ0_r_reg[20]/NET0131 ,
		_w6151_,
		_w8679_
	);
	LUT2 #(
		.INIT('h8)
	) name6534 (
		\u13_ints_r_reg[20]/NET0131 ,
		_w2741_,
		_w8680_
	);
	LUT2 #(
		.INIT('h1)
	) name6535 (
		_w8676_,
		_w8677_,
		_w8681_
	);
	LUT2 #(
		.INIT('h1)
	) name6536 (
		_w8678_,
		_w8679_,
		_w8682_
	);
	LUT2 #(
		.INIT('h4)
	) name6537 (
		_w8680_,
		_w8682_,
		_w8683_
	);
	LUT2 #(
		.INIT('h8)
	) name6538 (
		_w8681_,
		_w8683_,
		_w8684_
	);
	LUT2 #(
		.INIT('h2)
	) name6539 (
		_w6146_,
		_w8684_,
		_w8685_
	);
	LUT2 #(
		.INIT('h8)
	) name6540 (
		\u9_dout_reg[20]/P0001 ,
		_w6168_,
		_w8686_
	);
	LUT2 #(
		.INIT('h8)
	) name6541 (
		\u10_dout_reg[20]/P0001 ,
		_w6170_,
		_w8687_
	);
	LUT2 #(
		.INIT('h8)
	) name6542 (
		\u11_dout_reg[20]/P0001 ,
		_w6145_,
		_w8688_
	);
	LUT2 #(
		.INIT('h1)
	) name6543 (
		_w8686_,
		_w8687_,
		_w8689_
	);
	LUT2 #(
		.INIT('h4)
	) name6544 (
		_w8688_,
		_w8689_,
		_w8690_
	);
	LUT2 #(
		.INIT('h4)
	) name6545 (
		_w8685_,
		_w8690_,
		_w8691_
	);
	LUT2 #(
		.INIT('h8)
	) name6546 (
		\u13_icc_r_reg[21]/NET0131 ,
		_w6157_,
		_w8692_
	);
	LUT2 #(
		.INIT('h8)
	) name6547 (
		\u13_intm_r_reg[21]/NET0131 ,
		_w6153_,
		_w8693_
	);
	LUT2 #(
		.INIT('h8)
	) name6548 (
		\u13_crac_r_reg[5]/NET0131 ,
		_w6159_,
		_w8694_
	);
	LUT2 #(
		.INIT('h8)
	) name6549 (
		\u13_occ0_r_reg[21]/NET0131 ,
		_w6151_,
		_w8695_
	);
	LUT2 #(
		.INIT('h8)
	) name6550 (
		\u13_ints_r_reg[21]/NET0131 ,
		_w2741_,
		_w8696_
	);
	LUT2 #(
		.INIT('h1)
	) name6551 (
		_w8692_,
		_w8693_,
		_w8697_
	);
	LUT2 #(
		.INIT('h1)
	) name6552 (
		_w8694_,
		_w8695_,
		_w8698_
	);
	LUT2 #(
		.INIT('h4)
	) name6553 (
		_w8696_,
		_w8698_,
		_w8699_
	);
	LUT2 #(
		.INIT('h8)
	) name6554 (
		_w8697_,
		_w8699_,
		_w8700_
	);
	LUT2 #(
		.INIT('h2)
	) name6555 (
		_w6146_,
		_w8700_,
		_w8701_
	);
	LUT2 #(
		.INIT('h8)
	) name6556 (
		\u9_dout_reg[21]/P0001 ,
		_w6168_,
		_w8702_
	);
	LUT2 #(
		.INIT('h8)
	) name6557 (
		\u10_dout_reg[21]/P0001 ,
		_w6170_,
		_w8703_
	);
	LUT2 #(
		.INIT('h8)
	) name6558 (
		\u11_dout_reg[21]/P0001 ,
		_w6145_,
		_w8704_
	);
	LUT2 #(
		.INIT('h1)
	) name6559 (
		_w8702_,
		_w8703_,
		_w8705_
	);
	LUT2 #(
		.INIT('h4)
	) name6560 (
		_w8704_,
		_w8705_,
		_w8706_
	);
	LUT2 #(
		.INIT('h4)
	) name6561 (
		_w8701_,
		_w8706_,
		_w8707_
	);
	LUT2 #(
		.INIT('h8)
	) name6562 (
		\u13_icc_r_reg[22]/NET0131 ,
		_w6157_,
		_w8708_
	);
	LUT2 #(
		.INIT('h8)
	) name6563 (
		\u13_intm_r_reg[22]/NET0131 ,
		_w6153_,
		_w8709_
	);
	LUT2 #(
		.INIT('h8)
	) name6564 (
		\u13_crac_r_reg[6]/NET0131 ,
		_w6159_,
		_w8710_
	);
	LUT2 #(
		.INIT('h8)
	) name6565 (
		\u13_occ0_r_reg[22]/NET0131 ,
		_w6151_,
		_w8711_
	);
	LUT2 #(
		.INIT('h8)
	) name6566 (
		\u13_ints_r_reg[22]/NET0131 ,
		_w2741_,
		_w8712_
	);
	LUT2 #(
		.INIT('h1)
	) name6567 (
		_w8708_,
		_w8709_,
		_w8713_
	);
	LUT2 #(
		.INIT('h1)
	) name6568 (
		_w8710_,
		_w8711_,
		_w8714_
	);
	LUT2 #(
		.INIT('h4)
	) name6569 (
		_w8712_,
		_w8714_,
		_w8715_
	);
	LUT2 #(
		.INIT('h8)
	) name6570 (
		_w8713_,
		_w8715_,
		_w8716_
	);
	LUT2 #(
		.INIT('h2)
	) name6571 (
		_w6146_,
		_w8716_,
		_w8717_
	);
	LUT2 #(
		.INIT('h8)
	) name6572 (
		\u9_dout_reg[22]/P0001 ,
		_w6168_,
		_w8718_
	);
	LUT2 #(
		.INIT('h8)
	) name6573 (
		\u10_dout_reg[22]/P0001 ,
		_w6170_,
		_w8719_
	);
	LUT2 #(
		.INIT('h8)
	) name6574 (
		\u11_dout_reg[22]/P0001 ,
		_w6145_,
		_w8720_
	);
	LUT2 #(
		.INIT('h1)
	) name6575 (
		_w8718_,
		_w8719_,
		_w8721_
	);
	LUT2 #(
		.INIT('h4)
	) name6576 (
		_w8720_,
		_w8721_,
		_w8722_
	);
	LUT2 #(
		.INIT('h4)
	) name6577 (
		_w8717_,
		_w8722_,
		_w8723_
	);
	LUT2 #(
		.INIT('h8)
	) name6578 (
		\u13_ints_r_reg[23]/NET0131 ,
		_w2741_,
		_w8724_
	);
	LUT2 #(
		.INIT('h8)
	) name6579 (
		\u13_intm_r_reg[23]/NET0131 ,
		_w6153_,
		_w8725_
	);
	LUT2 #(
		.INIT('h8)
	) name6580 (
		\u13_occ0_r_reg[23]/NET0131 ,
		_w6151_,
		_w8726_
	);
	LUT2 #(
		.INIT('h8)
	) name6581 (
		\u13_icc_r_reg[23]/NET0131 ,
		_w6157_,
		_w8727_
	);
	LUT2 #(
		.INIT('h1)
	) name6582 (
		_w8724_,
		_w8725_,
		_w8728_
	);
	LUT2 #(
		.INIT('h1)
	) name6583 (
		_w8726_,
		_w8727_,
		_w8729_
	);
	LUT2 #(
		.INIT('h8)
	) name6584 (
		_w8728_,
		_w8729_,
		_w8730_
	);
	LUT2 #(
		.INIT('h2)
	) name6585 (
		_w6146_,
		_w8730_,
		_w8731_
	);
	LUT2 #(
		.INIT('h8)
	) name6586 (
		\u9_dout_reg[23]/P0001 ,
		_w6168_,
		_w8732_
	);
	LUT2 #(
		.INIT('h8)
	) name6587 (
		\u11_dout_reg[23]/P0001 ,
		_w6145_,
		_w8733_
	);
	LUT2 #(
		.INIT('h8)
	) name6588 (
		\u10_dout_reg[23]/P0001 ,
		_w6170_,
		_w8734_
	);
	LUT2 #(
		.INIT('h1)
	) name6589 (
		_w8732_,
		_w8733_,
		_w8735_
	);
	LUT2 #(
		.INIT('h4)
	) name6590 (
		_w8734_,
		_w8735_,
		_w8736_
	);
	LUT2 #(
		.INIT('h4)
	) name6591 (
		_w8731_,
		_w8736_,
		_w8737_
	);
	LUT2 #(
		.INIT('h1)
	) name6592 (
		\u10_rp_reg[0]/P0001 ,
		\u12_i4_re_reg/P0001 ,
		_w8738_
	);
	LUT2 #(
		.INIT('h2)
	) name6593 (
		\u13_icc_r_reg[8]/NET0131 ,
		_w8597_,
		_w8739_
	);
	LUT2 #(
		.INIT('h4)
	) name6594 (
		_w8738_,
		_w8739_,
		_w8740_
	);
	LUT2 #(
		.INIT('h8)
	) name6595 (
		\u13_crac_r_reg[2]/NET0131 ,
		_w6159_,
		_w8741_
	);
	LUT2 #(
		.INIT('h8)
	) name6596 (
		\u13_intm_r_reg[18]/NET0131 ,
		_w6153_,
		_w8742_
	);
	LUT2 #(
		.INIT('h8)
	) name6597 (
		\u13_icc_r_reg[18]/NET0131 ,
		_w6157_,
		_w8743_
	);
	LUT2 #(
		.INIT('h8)
	) name6598 (
		\u13_occ0_r_reg[18]/NET0131 ,
		_w6151_,
		_w8744_
	);
	LUT2 #(
		.INIT('h8)
	) name6599 (
		\u13_ints_r_reg[18]/NET0131 ,
		_w2741_,
		_w8745_
	);
	LUT2 #(
		.INIT('h1)
	) name6600 (
		_w8741_,
		_w8742_,
		_w8746_
	);
	LUT2 #(
		.INIT('h1)
	) name6601 (
		_w8743_,
		_w8744_,
		_w8747_
	);
	LUT2 #(
		.INIT('h4)
	) name6602 (
		_w8745_,
		_w8747_,
		_w8748_
	);
	LUT2 #(
		.INIT('h8)
	) name6603 (
		_w8746_,
		_w8748_,
		_w8749_
	);
	LUT2 #(
		.INIT('h2)
	) name6604 (
		_w6146_,
		_w8749_,
		_w8750_
	);
	LUT2 #(
		.INIT('h8)
	) name6605 (
		\u9_dout_reg[18]/P0001 ,
		_w6168_,
		_w8751_
	);
	LUT2 #(
		.INIT('h8)
	) name6606 (
		\u10_dout_reg[18]/P0001 ,
		_w6170_,
		_w8752_
	);
	LUT2 #(
		.INIT('h8)
	) name6607 (
		\u11_dout_reg[18]/P0001 ,
		_w6145_,
		_w8753_
	);
	LUT2 #(
		.INIT('h1)
	) name6608 (
		_w8751_,
		_w8752_,
		_w8754_
	);
	LUT2 #(
		.INIT('h4)
	) name6609 (
		_w8753_,
		_w8754_,
		_w8755_
	);
	LUT2 #(
		.INIT('h4)
	) name6610 (
		_w8750_,
		_w8755_,
		_w8756_
	);
	LUT2 #(
		.INIT('h8)
	) name6611 (
		\u2_to_cnt_reg[4]/NET0131 ,
		_w6481_,
		_w8757_
	);
	LUT2 #(
		.INIT('h1)
	) name6612 (
		\u2_to_cnt_reg[4]/NET0131 ,
		_w6481_,
		_w8758_
	);
	LUT2 #(
		.INIT('h1)
	) name6613 (
		\u2_bit_clk_e_reg/P0001 ,
		_w8757_,
		_w8759_
	);
	LUT2 #(
		.INIT('h4)
	) name6614 (
		_w8758_,
		_w8759_,
		_w8760_
	);
	LUT2 #(
		.INIT('h1)
	) name6615 (
		\u2_to_cnt_reg[5]/NET0131 ,
		_w8757_,
		_w8761_
	);
	LUT2 #(
		.INIT('h8)
	) name6616 (
		\u2_to_cnt_reg[5]/NET0131 ,
		_w8757_,
		_w8762_
	);
	LUT2 #(
		.INIT('h1)
	) name6617 (
		\u2_bit_clk_e_reg/P0001 ,
		_w8761_,
		_w8763_
	);
	LUT2 #(
		.INIT('h4)
	) name6618 (
		_w8762_,
		_w8763_,
		_w8764_
	);
	LUT2 #(
		.INIT('h1)
	) name6619 (
		\u2_to_cnt_reg[2]/NET0131 ,
		_w6479_,
		_w8765_
	);
	LUT2 #(
		.INIT('h1)
	) name6620 (
		\u2_bit_clk_e_reg/P0001 ,
		_w6480_,
		_w8766_
	);
	LUT2 #(
		.INIT('h4)
	) name6621 (
		_w8765_,
		_w8766_,
		_w8767_
	);
	LUT2 #(
		.INIT('h8)
	) name6622 (
		\u12_i3_re_reg/NET0131 ,
		\u9_empty_reg/P0001 ,
		_w8768_
	);
	LUT2 #(
		.INIT('h1)
	) name6623 (
		\u23_int_set_reg[1]/NET0131 ,
		_w8768_,
		_w8769_
	);
	LUT2 #(
		.INIT('h8)
	) name6624 (
		\u10_empty_reg/P0001 ,
		\u12_i4_re_reg/P0001 ,
		_w8770_
	);
	LUT2 #(
		.INIT('h1)
	) name6625 (
		\u24_int_set_reg[1]/NET0131 ,
		_w8770_,
		_w8771_
	);
	LUT2 #(
		.INIT('h8)
	) name6626 (
		\u11_empty_reg/P0001 ,
		\u12_i6_re_reg/NET0131 ,
		_w8772_
	);
	LUT2 #(
		.INIT('h1)
	) name6627 (
		\u25_int_set_reg[1]/NET0131 ,
		_w8772_,
		_w8773_
	);
	LUT2 #(
		.INIT('h1)
	) name6628 (
		\u2_res_cnt_reg[0]/P0001 ,
		_w5629_,
		_w8774_
	);
	LUT2 #(
		.INIT('h2)
	) name6629 (
		\u2_sync_resume_reg/NET0131 ,
		_w6454_,
		_w8775_
	);
	LUT2 #(
		.INIT('h4)
	) name6630 (
		_w8774_,
		_w8775_,
		_w8776_
	);
	LUT2 #(
		.INIT('h8)
	) name6631 (
		wb_we_i_pad,
		_w2735_,
		_w8777_
	);
	LUT2 #(
		.INIT('h8)
	) name6632 (
		\u12_we1_reg/P0001 ,
		_w8777_,
		_w8778_
	);
	LUT2 #(
		.INIT('h4)
	) name6633 (
		\u12_we2_reg/P0001 ,
		_w8778_,
		_w8779_
	);
	LUT2 #(
		.INIT('h8)
	) name6634 (
		_w6139_,
		_w8779_,
		_w8780_
	);
	LUT2 #(
		.INIT('h8)
	) name6635 (
		_w6143_,
		_w8780_,
		_w8781_
	);
	LUT2 #(
		.INIT('h8)
	) name6636 (
		_w6151_,
		_w8780_,
		_w8782_
	);
	LUT2 #(
		.INIT('h8)
	) name6637 (
		_w6147_,
		_w8780_,
		_w8783_
	);
	LUT2 #(
		.INIT('h8)
	) name6638 (
		_w6159_,
		_w8780_,
		_w8784_
	);
	LUT2 #(
		.INIT('h8)
	) name6639 (
		_w6153_,
		_w8780_,
		_w8785_
	);
	LUT2 #(
		.INIT('h8)
	) name6640 (
		\u13_occ0_r_reg[24]/NET0131 ,
		_w6151_,
		_w8786_
	);
	LUT2 #(
		.INIT('h8)
	) name6641 (
		\u13_intm_r_reg[24]/NET0131 ,
		_w6153_,
		_w8787_
	);
	LUT2 #(
		.INIT('h8)
	) name6642 (
		\u13_ints_r_reg[24]/NET0131 ,
		_w2741_,
		_w8788_
	);
	LUT2 #(
		.INIT('h1)
	) name6643 (
		_w8786_,
		_w8787_,
		_w8789_
	);
	LUT2 #(
		.INIT('h4)
	) name6644 (
		_w8788_,
		_w8789_,
		_w8790_
	);
	LUT2 #(
		.INIT('h2)
	) name6645 (
		_w6146_,
		_w8790_,
		_w8791_
	);
	LUT2 #(
		.INIT('h8)
	) name6646 (
		\u9_dout_reg[24]/P0001 ,
		_w6168_,
		_w8792_
	);
	LUT2 #(
		.INIT('h8)
	) name6647 (
		\u11_dout_reg[24]/P0001 ,
		_w6145_,
		_w8793_
	);
	LUT2 #(
		.INIT('h8)
	) name6648 (
		\u10_dout_reg[24]/P0001 ,
		_w6170_,
		_w8794_
	);
	LUT2 #(
		.INIT('h1)
	) name6649 (
		_w8792_,
		_w8793_,
		_w8795_
	);
	LUT2 #(
		.INIT('h4)
	) name6650 (
		_w8794_,
		_w8795_,
		_w8796_
	);
	LUT2 #(
		.INIT('h4)
	) name6651 (
		_w8791_,
		_w8796_,
		_w8797_
	);
	LUT2 #(
		.INIT('h8)
	) name6652 (
		\u13_occ0_r_reg[25]/NET0131 ,
		_w6151_,
		_w8798_
	);
	LUT2 #(
		.INIT('h8)
	) name6653 (
		\u13_intm_r_reg[25]/NET0131 ,
		_w6153_,
		_w8799_
	);
	LUT2 #(
		.INIT('h8)
	) name6654 (
		\u13_ints_r_reg[25]/NET0131 ,
		_w2741_,
		_w8800_
	);
	LUT2 #(
		.INIT('h1)
	) name6655 (
		_w8798_,
		_w8799_,
		_w8801_
	);
	LUT2 #(
		.INIT('h4)
	) name6656 (
		_w8800_,
		_w8801_,
		_w8802_
	);
	LUT2 #(
		.INIT('h2)
	) name6657 (
		_w6146_,
		_w8802_,
		_w8803_
	);
	LUT2 #(
		.INIT('h8)
	) name6658 (
		\u9_dout_reg[25]/P0001 ,
		_w6168_,
		_w8804_
	);
	LUT2 #(
		.INIT('h8)
	) name6659 (
		\u11_dout_reg[25]/P0001 ,
		_w6145_,
		_w8805_
	);
	LUT2 #(
		.INIT('h8)
	) name6660 (
		\u10_dout_reg[25]/P0001 ,
		_w6170_,
		_w8806_
	);
	LUT2 #(
		.INIT('h1)
	) name6661 (
		_w8804_,
		_w8805_,
		_w8807_
	);
	LUT2 #(
		.INIT('h4)
	) name6662 (
		_w8806_,
		_w8807_,
		_w8808_
	);
	LUT2 #(
		.INIT('h4)
	) name6663 (
		_w8803_,
		_w8808_,
		_w8809_
	);
	LUT2 #(
		.INIT('h8)
	) name6664 (
		\u13_occ0_r_reg[26]/NET0131 ,
		_w6151_,
		_w8810_
	);
	LUT2 #(
		.INIT('h8)
	) name6665 (
		\u13_intm_r_reg[26]/NET0131 ,
		_w6153_,
		_w8811_
	);
	LUT2 #(
		.INIT('h8)
	) name6666 (
		\u13_ints_r_reg[26]/NET0131 ,
		_w2741_,
		_w8812_
	);
	LUT2 #(
		.INIT('h1)
	) name6667 (
		_w8810_,
		_w8811_,
		_w8813_
	);
	LUT2 #(
		.INIT('h4)
	) name6668 (
		_w8812_,
		_w8813_,
		_w8814_
	);
	LUT2 #(
		.INIT('h2)
	) name6669 (
		_w6146_,
		_w8814_,
		_w8815_
	);
	LUT2 #(
		.INIT('h8)
	) name6670 (
		\u9_dout_reg[26]/P0001 ,
		_w6168_,
		_w8816_
	);
	LUT2 #(
		.INIT('h8)
	) name6671 (
		\u11_dout_reg[26]/P0001 ,
		_w6145_,
		_w8817_
	);
	LUT2 #(
		.INIT('h8)
	) name6672 (
		\u10_dout_reg[26]/P0001 ,
		_w6170_,
		_w8818_
	);
	LUT2 #(
		.INIT('h1)
	) name6673 (
		_w8816_,
		_w8817_,
		_w8819_
	);
	LUT2 #(
		.INIT('h4)
	) name6674 (
		_w8818_,
		_w8819_,
		_w8820_
	);
	LUT2 #(
		.INIT('h4)
	) name6675 (
		_w8815_,
		_w8820_,
		_w8821_
	);
	LUT2 #(
		.INIT('h8)
	) name6676 (
		\u13_occ0_r_reg[27]/NET0131 ,
		_w6151_,
		_w8822_
	);
	LUT2 #(
		.INIT('h8)
	) name6677 (
		\u13_intm_r_reg[27]/NET0131 ,
		_w6153_,
		_w8823_
	);
	LUT2 #(
		.INIT('h8)
	) name6678 (
		\u13_ints_r_reg[27]/NET0131 ,
		_w2741_,
		_w8824_
	);
	LUT2 #(
		.INIT('h1)
	) name6679 (
		_w8822_,
		_w8823_,
		_w8825_
	);
	LUT2 #(
		.INIT('h4)
	) name6680 (
		_w8824_,
		_w8825_,
		_w8826_
	);
	LUT2 #(
		.INIT('h2)
	) name6681 (
		_w6146_,
		_w8826_,
		_w8827_
	);
	LUT2 #(
		.INIT('h8)
	) name6682 (
		\u9_dout_reg[27]/P0001 ,
		_w6168_,
		_w8828_
	);
	LUT2 #(
		.INIT('h8)
	) name6683 (
		\u11_dout_reg[27]/P0001 ,
		_w6145_,
		_w8829_
	);
	LUT2 #(
		.INIT('h8)
	) name6684 (
		\u10_dout_reg[27]/P0001 ,
		_w6170_,
		_w8830_
	);
	LUT2 #(
		.INIT('h1)
	) name6685 (
		_w8828_,
		_w8829_,
		_w8831_
	);
	LUT2 #(
		.INIT('h4)
	) name6686 (
		_w8830_,
		_w8831_,
		_w8832_
	);
	LUT2 #(
		.INIT('h4)
	) name6687 (
		_w8827_,
		_w8832_,
		_w8833_
	);
	LUT2 #(
		.INIT('h8)
	) name6688 (
		\u13_occ0_r_reg[28]/NET0131 ,
		_w6151_,
		_w8834_
	);
	LUT2 #(
		.INIT('h8)
	) name6689 (
		\u13_intm_r_reg[28]/NET0131 ,
		_w6153_,
		_w8835_
	);
	LUT2 #(
		.INIT('h8)
	) name6690 (
		\u13_ints_r_reg[28]/NET0131 ,
		_w2741_,
		_w8836_
	);
	LUT2 #(
		.INIT('h1)
	) name6691 (
		_w8834_,
		_w8835_,
		_w8837_
	);
	LUT2 #(
		.INIT('h4)
	) name6692 (
		_w8836_,
		_w8837_,
		_w8838_
	);
	LUT2 #(
		.INIT('h2)
	) name6693 (
		_w6146_,
		_w8838_,
		_w8839_
	);
	LUT2 #(
		.INIT('h8)
	) name6694 (
		\u9_dout_reg[28]/P0001 ,
		_w6168_,
		_w8840_
	);
	LUT2 #(
		.INIT('h8)
	) name6695 (
		\u11_dout_reg[28]/P0001 ,
		_w6145_,
		_w8841_
	);
	LUT2 #(
		.INIT('h8)
	) name6696 (
		\u10_dout_reg[28]/P0001 ,
		_w6170_,
		_w8842_
	);
	LUT2 #(
		.INIT('h1)
	) name6697 (
		_w8840_,
		_w8841_,
		_w8843_
	);
	LUT2 #(
		.INIT('h4)
	) name6698 (
		_w8842_,
		_w8843_,
		_w8844_
	);
	LUT2 #(
		.INIT('h4)
	) name6699 (
		_w8839_,
		_w8844_,
		_w8845_
	);
	LUT2 #(
		.INIT('h8)
	) name6700 (
		\u13_occ0_r_reg[29]/NET0131 ,
		_w6151_,
		_w8846_
	);
	LUT2 #(
		.INIT('h8)
	) name6701 (
		\u11_dout_reg[29]/P0001 ,
		_w6145_,
		_w8847_
	);
	LUT2 #(
		.INIT('h8)
	) name6702 (
		\u9_dout_reg[29]/P0001 ,
		_w6168_,
		_w8848_
	);
	LUT2 #(
		.INIT('h8)
	) name6703 (
		\u10_dout_reg[29]/P0001 ,
		_w6170_,
		_w8849_
	);
	LUT2 #(
		.INIT('h1)
	) name6704 (
		_w8846_,
		_w8847_,
		_w8850_
	);
	LUT2 #(
		.INIT('h1)
	) name6705 (
		_w8848_,
		_w8849_,
		_w8851_
	);
	LUT2 #(
		.INIT('h8)
	) name6706 (
		_w8850_,
		_w8851_,
		_w8852_
	);
	LUT2 #(
		.INIT('h8)
	) name6707 (
		\u13_occ0_r_reg[30]/NET0131 ,
		_w6151_,
		_w8853_
	);
	LUT2 #(
		.INIT('h8)
	) name6708 (
		\u11_dout_reg[30]/P0001 ,
		_w6145_,
		_w8854_
	);
	LUT2 #(
		.INIT('h8)
	) name6709 (
		\u9_dout_reg[30]/P0001 ,
		_w6168_,
		_w8855_
	);
	LUT2 #(
		.INIT('h8)
	) name6710 (
		\u10_dout_reg[30]/P0001 ,
		_w6170_,
		_w8856_
	);
	LUT2 #(
		.INIT('h1)
	) name6711 (
		_w8853_,
		_w8854_,
		_w8857_
	);
	LUT2 #(
		.INIT('h1)
	) name6712 (
		_w8855_,
		_w8856_,
		_w8858_
	);
	LUT2 #(
		.INIT('h8)
	) name6713 (
		_w8857_,
		_w8858_,
		_w8859_
	);
	LUT2 #(
		.INIT('h8)
	) name6714 (
		\u13_crac_r_reg[7]/NET0131 ,
		_w6159_,
		_w8860_
	);
	LUT2 #(
		.INIT('h8)
	) name6715 (
		\u13_occ0_r_reg[31]/NET0131 ,
		_w6151_,
		_w8861_
	);
	LUT2 #(
		.INIT('h8)
	) name6716 (
		\u10_dout_reg[31]/P0001 ,
		_w6170_,
		_w8862_
	);
	LUT2 #(
		.INIT('h8)
	) name6717 (
		\u11_dout_reg[31]/P0001 ,
		_w6145_,
		_w8863_
	);
	LUT2 #(
		.INIT('h8)
	) name6718 (
		\u9_dout_reg[31]/P0001 ,
		_w6168_,
		_w8864_
	);
	LUT2 #(
		.INIT('h1)
	) name6719 (
		_w8860_,
		_w8861_,
		_w8865_
	);
	LUT2 #(
		.INIT('h4)
	) name6720 (
		_w8862_,
		_w8865_,
		_w8866_
	);
	LUT2 #(
		.INIT('h1)
	) name6721 (
		_w8863_,
		_w8864_,
		_w8867_
	);
	LUT2 #(
		.INIT('h8)
	) name6722 (
		_w8866_,
		_w8867_,
		_w8868_
	);
	LUT2 #(
		.INIT('h1)
	) name6723 (
		\u2_res_cnt_reg[1]/P0001 ,
		_w6454_,
		_w8869_
	);
	LUT2 #(
		.INIT('h2)
	) name6724 (
		\u2_sync_resume_reg/NET0131 ,
		_w6455_,
		_w8870_
	);
	LUT2 #(
		.INIT('h4)
	) name6725 (
		_w8869_,
		_w8870_,
		_w8871_
	);
	LUT2 #(
		.INIT('h1)
	) name6726 (
		\u2_cnt_reg[3]/NET0131 ,
		_w6470_,
		_w8872_
	);
	LUT2 #(
		.INIT('h1)
	) name6727 (
		_w6471_,
		_w8872_,
		_w8873_
	);
	LUT2 #(
		.INIT('h1)
	) name6728 (
		suspended_o_pad,
		_w8873_,
		_w8874_
	);
	LUT2 #(
		.INIT('h8)
	) name6729 (
		\u13_intm_r_reg[26]/NET0131 ,
		\u13_ints_r_reg[26]/NET0131 ,
		_w8875_
	);
	LUT2 #(
		.INIT('h8)
	) name6730 (
		\u13_intm_r_reg[15]/NET0131 ,
		\u13_ints_r_reg[15]/NET0131 ,
		_w8876_
	);
	LUT2 #(
		.INIT('h8)
	) name6731 (
		\u13_intm_r_reg[0]/NET0131 ,
		\u13_ints_r_reg[0]/NET0131 ,
		_w8877_
	);
	LUT2 #(
		.INIT('h8)
	) name6732 (
		\u13_intm_r_reg[28]/NET0131 ,
		\u13_ints_r_reg[28]/NET0131 ,
		_w8878_
	);
	LUT2 #(
		.INIT('h8)
	) name6733 (
		\u13_intm_r_reg[1]/NET0131 ,
		\u13_ints_r_reg[1]/NET0131 ,
		_w8879_
	);
	LUT2 #(
		.INIT('h8)
	) name6734 (
		\u13_intm_r_reg[13]/NET0131 ,
		\u13_ints_r_reg[13]/NET0131 ,
		_w8880_
	);
	LUT2 #(
		.INIT('h8)
	) name6735 (
		\u13_intm_r_reg[11]/NET0131 ,
		\u13_ints_r_reg[11]/NET0131 ,
		_w8881_
	);
	LUT2 #(
		.INIT('h8)
	) name6736 (
		\u13_intm_r_reg[6]/NET0131 ,
		\u13_ints_r_reg[6]/NET0131 ,
		_w8882_
	);
	LUT2 #(
		.INIT('h8)
	) name6737 (
		\u13_intm_r_reg[5]/NET0131 ,
		\u13_ints_r_reg[5]/NET0131 ,
		_w8883_
	);
	LUT2 #(
		.INIT('h8)
	) name6738 (
		\u13_intm_r_reg[8]/NET0131 ,
		\u13_ints_r_reg[8]/NET0131 ,
		_w8884_
	);
	LUT2 #(
		.INIT('h8)
	) name6739 (
		\u13_intm_r_reg[7]/NET0131 ,
		\u13_ints_r_reg[7]/NET0131 ,
		_w8885_
	);
	LUT2 #(
		.INIT('h8)
	) name6740 (
		\u13_intm_r_reg[23]/NET0131 ,
		\u13_ints_r_reg[23]/NET0131 ,
		_w8886_
	);
	LUT2 #(
		.INIT('h8)
	) name6741 (
		\u13_intm_r_reg[24]/NET0131 ,
		\u13_ints_r_reg[24]/NET0131 ,
		_w8887_
	);
	LUT2 #(
		.INIT('h8)
	) name6742 (
		\u13_intm_r_reg[14]/NET0131 ,
		\u13_ints_r_reg[14]/NET0131 ,
		_w8888_
	);
	LUT2 #(
		.INIT('h8)
	) name6743 (
		\u13_intm_r_reg[22]/NET0131 ,
		\u13_ints_r_reg[22]/NET0131 ,
		_w8889_
	);
	LUT2 #(
		.INIT('h8)
	) name6744 (
		\u13_intm_r_reg[12]/NET0131 ,
		\u13_ints_r_reg[12]/NET0131 ,
		_w8890_
	);
	LUT2 #(
		.INIT('h8)
	) name6745 (
		\u13_intm_r_reg[19]/NET0131 ,
		\u13_ints_r_reg[19]/NET0131 ,
		_w8891_
	);
	LUT2 #(
		.INIT('h8)
	) name6746 (
		\u13_intm_r_reg[27]/NET0131 ,
		\u13_ints_r_reg[27]/NET0131 ,
		_w8892_
	);
	LUT2 #(
		.INIT('h8)
	) name6747 (
		\u13_intm_r_reg[9]/NET0131 ,
		\u13_ints_r_reg[9]/NET0131 ,
		_w8893_
	);
	LUT2 #(
		.INIT('h8)
	) name6748 (
		\u13_intm_r_reg[10]/NET0131 ,
		\u13_ints_r_reg[10]/NET0131 ,
		_w8894_
	);
	LUT2 #(
		.INIT('h8)
	) name6749 (
		\u13_intm_r_reg[4]/NET0131 ,
		\u13_ints_r_reg[4]/NET0131 ,
		_w8895_
	);
	LUT2 #(
		.INIT('h8)
	) name6750 (
		\u13_intm_r_reg[21]/NET0131 ,
		\u13_ints_r_reg[21]/NET0131 ,
		_w8896_
	);
	LUT2 #(
		.INIT('h8)
	) name6751 (
		\u13_intm_r_reg[17]/NET0131 ,
		\u13_ints_r_reg[17]/NET0131 ,
		_w8897_
	);
	LUT2 #(
		.INIT('h8)
	) name6752 (
		\u13_intm_r_reg[16]/NET0131 ,
		\u13_ints_r_reg[16]/NET0131 ,
		_w8898_
	);
	LUT2 #(
		.INIT('h8)
	) name6753 (
		\u13_intm_r_reg[20]/NET0131 ,
		\u13_ints_r_reg[20]/NET0131 ,
		_w8899_
	);
	LUT2 #(
		.INIT('h8)
	) name6754 (
		\u13_intm_r_reg[2]/NET0131 ,
		\u13_ints_r_reg[2]/NET0131 ,
		_w8900_
	);
	LUT2 #(
		.INIT('h8)
	) name6755 (
		\u13_intm_r_reg[25]/NET0131 ,
		\u13_ints_r_reg[25]/NET0131 ,
		_w8901_
	);
	LUT2 #(
		.INIT('h8)
	) name6756 (
		\u13_intm_r_reg[18]/NET0131 ,
		\u13_ints_r_reg[18]/NET0131 ,
		_w8902_
	);
	LUT2 #(
		.INIT('h8)
	) name6757 (
		\u13_intm_r_reg[3]/NET0131 ,
		\u13_ints_r_reg[3]/NET0131 ,
		_w8903_
	);
	LUT2 #(
		.INIT('h1)
	) name6758 (
		_w8875_,
		_w8876_,
		_w8904_
	);
	LUT2 #(
		.INIT('h1)
	) name6759 (
		_w8877_,
		_w8878_,
		_w8905_
	);
	LUT2 #(
		.INIT('h1)
	) name6760 (
		_w8879_,
		_w8880_,
		_w8906_
	);
	LUT2 #(
		.INIT('h1)
	) name6761 (
		_w8881_,
		_w8882_,
		_w8907_
	);
	LUT2 #(
		.INIT('h1)
	) name6762 (
		_w8883_,
		_w8884_,
		_w8908_
	);
	LUT2 #(
		.INIT('h1)
	) name6763 (
		_w8885_,
		_w8886_,
		_w8909_
	);
	LUT2 #(
		.INIT('h1)
	) name6764 (
		_w8887_,
		_w8888_,
		_w8910_
	);
	LUT2 #(
		.INIT('h1)
	) name6765 (
		_w8889_,
		_w8890_,
		_w8911_
	);
	LUT2 #(
		.INIT('h1)
	) name6766 (
		_w8891_,
		_w8892_,
		_w8912_
	);
	LUT2 #(
		.INIT('h1)
	) name6767 (
		_w8893_,
		_w8894_,
		_w8913_
	);
	LUT2 #(
		.INIT('h1)
	) name6768 (
		_w8895_,
		_w8896_,
		_w8914_
	);
	LUT2 #(
		.INIT('h1)
	) name6769 (
		_w8897_,
		_w8898_,
		_w8915_
	);
	LUT2 #(
		.INIT('h1)
	) name6770 (
		_w8899_,
		_w8900_,
		_w8916_
	);
	LUT2 #(
		.INIT('h1)
	) name6771 (
		_w8901_,
		_w8902_,
		_w8917_
	);
	LUT2 #(
		.INIT('h4)
	) name6772 (
		_w8903_,
		_w8917_,
		_w8918_
	);
	LUT2 #(
		.INIT('h8)
	) name6773 (
		_w8915_,
		_w8916_,
		_w8919_
	);
	LUT2 #(
		.INIT('h8)
	) name6774 (
		_w8913_,
		_w8914_,
		_w8920_
	);
	LUT2 #(
		.INIT('h8)
	) name6775 (
		_w8911_,
		_w8912_,
		_w8921_
	);
	LUT2 #(
		.INIT('h8)
	) name6776 (
		_w8909_,
		_w8910_,
		_w8922_
	);
	LUT2 #(
		.INIT('h8)
	) name6777 (
		_w8907_,
		_w8908_,
		_w8923_
	);
	LUT2 #(
		.INIT('h8)
	) name6778 (
		_w8905_,
		_w8906_,
		_w8924_
	);
	LUT2 #(
		.INIT('h8)
	) name6779 (
		_w8904_,
		_w8924_,
		_w8925_
	);
	LUT2 #(
		.INIT('h8)
	) name6780 (
		_w8922_,
		_w8923_,
		_w8926_
	);
	LUT2 #(
		.INIT('h8)
	) name6781 (
		_w8920_,
		_w8921_,
		_w8927_
	);
	LUT2 #(
		.INIT('h8)
	) name6782 (
		_w8918_,
		_w8919_,
		_w8928_
	);
	LUT2 #(
		.INIT('h8)
	) name6783 (
		_w8927_,
		_w8928_,
		_w8929_
	);
	LUT2 #(
		.INIT('h8)
	) name6784 (
		_w8925_,
		_w8926_,
		_w8930_
	);
	LUT2 #(
		.INIT('h8)
	) name6785 (
		_w8929_,
		_w8930_,
		_w8931_
	);
	LUT2 #(
		.INIT('h8)
	) name6786 (
		_w6157_,
		_w8780_,
		_w8932_
	);
	LUT2 #(
		.INIT('h1)
	) name6787 (
		_w2738_,
		_w8779_,
		_w8933_
	);
	LUT2 #(
		.INIT('h4)
	) name6788 (
		wb_ack_o_pad,
		wb_cyc_i_pad,
		_w8934_
	);
	LUT2 #(
		.INIT('h4)
	) name6789 (
		_w8933_,
		_w8934_,
		_w8935_
	);
	LUT2 #(
		.INIT('h1)
	) name6790 (
		_w6287_,
		_w6292_,
		_w8936_
	);
	LUT2 #(
		.INIT('h1)
	) name6791 (
		_w8579_,
		_w8936_,
		_w8937_
	);
	LUT2 #(
		.INIT('h2)
	) name6792 (
		_w6225_,
		_w6228_,
		_w8938_
	);
	LUT2 #(
		.INIT('h1)
	) name6793 (
		_w6229_,
		_w8938_,
		_w8939_
	);
	LUT2 #(
		.INIT('h2)
	) name6794 (
		_w6236_,
		_w6239_,
		_w8940_
	);
	LUT2 #(
		.INIT('h1)
	) name6795 (
		_w6240_,
		_w8940_,
		_w8941_
	);
	LUT2 #(
		.INIT('h2)
	) name6796 (
		_w6249_,
		_w6252_,
		_w8942_
	);
	LUT2 #(
		.INIT('h1)
	) name6797 (
		_w6253_,
		_w8942_,
		_w8943_
	);
	LUT2 #(
		.INIT('h1)
	) name6798 (
		_w6261_,
		_w6266_,
		_w8944_
	);
	LUT2 #(
		.INIT('h1)
	) name6799 (
		_w8537_,
		_w8944_,
		_w8945_
	);
	LUT2 #(
		.INIT('h2)
	) name6800 (
		_w6277_,
		_w6280_,
		_w8946_
	);
	LUT2 #(
		.INIT('h1)
	) name6801 (
		_w6281_,
		_w8946_,
		_w8947_
	);
	LUT2 #(
		.INIT('h8)
	) name6802 (
		_w2739_,
		_w8779_,
		_w8948_
	);
	LUT2 #(
		.INIT('h8)
	) name6803 (
		\u2_ld_reg/P0001 ,
		\u8_dout_reg[0]/P0001 ,
		_w8949_
	);
	LUT2 #(
		.INIT('h2)
	) name6804 (
		\u11_rp_reg[0]/P0001 ,
		\u11_wp_reg[1]/P0001 ,
		_w8950_
	);
	LUT2 #(
		.INIT('h2)
	) name6805 (
		\u11_rp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w8951_
	);
	LUT2 #(
		.INIT('h4)
	) name6806 (
		\u11_rp_reg[1]/P0001 ,
		\u11_wp_reg[2]/P0001 ,
		_w8952_
	);
	LUT2 #(
		.INIT('h1)
	) name6807 (
		_w8951_,
		_w8952_,
		_w8953_
	);
	LUT2 #(
		.INIT('h8)
	) name6808 (
		_w8950_,
		_w8953_,
		_w8954_
	);
	LUT2 #(
		.INIT('h1)
	) name6809 (
		_w8950_,
		_w8953_,
		_w8955_
	);
	LUT2 #(
		.INIT('h1)
	) name6810 (
		_w8954_,
		_w8955_,
		_w8956_
	);
	LUT2 #(
		.INIT('h2)
	) name6811 (
		\u9_rp_reg[0]/P0001 ,
		\u9_wp_reg[1]/P0001 ,
		_w8957_
	);
	LUT2 #(
		.INIT('h2)
	) name6812 (
		\u9_rp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w8958_
	);
	LUT2 #(
		.INIT('h4)
	) name6813 (
		\u9_rp_reg[1]/P0001 ,
		\u9_wp_reg[2]/P0001 ,
		_w8959_
	);
	LUT2 #(
		.INIT('h1)
	) name6814 (
		_w8958_,
		_w8959_,
		_w8960_
	);
	LUT2 #(
		.INIT('h8)
	) name6815 (
		_w8957_,
		_w8960_,
		_w8961_
	);
	LUT2 #(
		.INIT('h1)
	) name6816 (
		_w8957_,
		_w8960_,
		_w8962_
	);
	LUT2 #(
		.INIT('h1)
	) name6817 (
		_w8961_,
		_w8962_,
		_w8963_
	);
	LUT2 #(
		.INIT('h2)
	) name6818 (
		\u10_rp_reg[0]/P0001 ,
		\u10_wp_reg[1]/P0001 ,
		_w8964_
	);
	LUT2 #(
		.INIT('h2)
	) name6819 (
		\u10_rp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w8965_
	);
	LUT2 #(
		.INIT('h4)
	) name6820 (
		\u10_rp_reg[1]/P0001 ,
		\u10_wp_reg[2]/P0001 ,
		_w8966_
	);
	LUT2 #(
		.INIT('h1)
	) name6821 (
		_w8965_,
		_w8966_,
		_w8967_
	);
	LUT2 #(
		.INIT('h8)
	) name6822 (
		_w8964_,
		_w8967_,
		_w8968_
	);
	LUT2 #(
		.INIT('h1)
	) name6823 (
		_w8964_,
		_w8967_,
		_w8969_
	);
	LUT2 #(
		.INIT('h1)
	) name6824 (
		_w8968_,
		_w8969_,
		_w8970_
	);
	LUT2 #(
		.INIT('h1)
	) name6825 (
		\u13_ints_r_reg[0]/NET0131 ,
		\u15_crac_rd_done_reg/P0001 ,
		_w8971_
	);
	LUT2 #(
		.INIT('h1)
	) name6826 (
		_w2743_,
		_w8971_,
		_w8972_
	);
	LUT2 #(
		.INIT('h1)
	) name6827 (
		\u13_ints_r_reg[10]/NET0131 ,
		\u19_int_set_reg[2]/NET0131 ,
		_w8973_
	);
	LUT2 #(
		.INIT('h1)
	) name6828 (
		_w2743_,
		_w8973_,
		_w8974_
	);
	LUT2 #(
		.INIT('h1)
	) name6829 (
		\u13_ints_r_reg[12]/NET0131 ,
		\u20_int_set_reg[1]/NET0131 ,
		_w8975_
	);
	LUT2 #(
		.INIT('h1)
	) name6830 (
		_w2743_,
		_w8975_,
		_w8976_
	);
	LUT2 #(
		.INIT('h1)
	) name6831 (
		\u13_ints_r_reg[13]/NET0131 ,
		\u20_int_set_reg[2]/NET0131 ,
		_w8977_
	);
	LUT2 #(
		.INIT('h1)
	) name6832 (
		_w2743_,
		_w8977_,
		_w8978_
	);
	LUT2 #(
		.INIT('h1)
	) name6833 (
		\u13_ints_r_reg[15]/NET0131 ,
		\u21_int_set_reg[1]/NET0131 ,
		_w8979_
	);
	LUT2 #(
		.INIT('h1)
	) name6834 (
		_w2743_,
		_w8979_,
		_w8980_
	);
	LUT2 #(
		.INIT('h1)
	) name6835 (
		\u13_ints_r_reg[16]/NET0131 ,
		\u21_int_set_reg[2]/NET0131 ,
		_w8981_
	);
	LUT2 #(
		.INIT('h1)
	) name6836 (
		_w2743_,
		_w8981_,
		_w8982_
	);
	LUT2 #(
		.INIT('h1)
	) name6837 (
		\u13_ints_r_reg[18]/NET0131 ,
		\u22_int_set_reg[1]/NET0131 ,
		_w8983_
	);
	LUT2 #(
		.INIT('h1)
	) name6838 (
		_w2743_,
		_w8983_,
		_w8984_
	);
	LUT2 #(
		.INIT('h1)
	) name6839 (
		\u13_ints_r_reg[19]/NET0131 ,
		\u22_int_set_reg[2]/NET0131 ,
		_w8985_
	);
	LUT2 #(
		.INIT('h1)
	) name6840 (
		_w2743_,
		_w8985_,
		_w8986_
	);
	LUT2 #(
		.INIT('h1)
	) name6841 (
		\u13_ints_r_reg[21]/NET0131 ,
		\u23_int_set_reg[1]/NET0131 ,
		_w8987_
	);
	LUT2 #(
		.INIT('h1)
	) name6842 (
		_w2743_,
		_w8987_,
		_w8988_
	);
	LUT2 #(
		.INIT('h1)
	) name6843 (
		\u13_ints_r_reg[22]/NET0131 ,
		\u23_int_set_reg[2]/NET0131 ,
		_w8989_
	);
	LUT2 #(
		.INIT('h1)
	) name6844 (
		_w2743_,
		_w8989_,
		_w8990_
	);
	LUT2 #(
		.INIT('h1)
	) name6845 (
		\u13_ints_r_reg[24]/NET0131 ,
		\u24_int_set_reg[1]/NET0131 ,
		_w8991_
	);
	LUT2 #(
		.INIT('h1)
	) name6846 (
		_w2743_,
		_w8991_,
		_w8992_
	);
	LUT2 #(
		.INIT('h1)
	) name6847 (
		\u13_ints_r_reg[25]/NET0131 ,
		\u24_int_set_reg[2]/NET0131 ,
		_w8993_
	);
	LUT2 #(
		.INIT('h1)
	) name6848 (
		_w2743_,
		_w8993_,
		_w8994_
	);
	LUT2 #(
		.INIT('h1)
	) name6849 (
		\u13_ints_r_reg[27]/NET0131 ,
		\u25_int_set_reg[1]/NET0131 ,
		_w8995_
	);
	LUT2 #(
		.INIT('h1)
	) name6850 (
		_w2743_,
		_w8995_,
		_w8996_
	);
	LUT2 #(
		.INIT('h1)
	) name6851 (
		\u13_ints_r_reg[28]/NET0131 ,
		\u25_int_set_reg[2]/NET0131 ,
		_w8997_
	);
	LUT2 #(
		.INIT('h1)
	) name6852 (
		_w2743_,
		_w8997_,
		_w8998_
	);
	LUT2 #(
		.INIT('h1)
	) name6853 (
		\u13_ints_r_reg[3]/NET0131 ,
		\u17_int_set_reg[1]/NET0131 ,
		_w8999_
	);
	LUT2 #(
		.INIT('h1)
	) name6854 (
		_w2743_,
		_w8999_,
		_w9000_
	);
	LUT2 #(
		.INIT('h1)
	) name6855 (
		\u13_ints_r_reg[4]/NET0131 ,
		\u17_int_set_reg[2]/NET0131 ,
		_w9001_
	);
	LUT2 #(
		.INIT('h1)
	) name6856 (
		_w2743_,
		_w9001_,
		_w9002_
	);
	LUT2 #(
		.INIT('h1)
	) name6857 (
		\u13_ints_r_reg[6]/NET0131 ,
		\u18_int_set_reg[1]/NET0131 ,
		_w9003_
	);
	LUT2 #(
		.INIT('h1)
	) name6858 (
		_w2743_,
		_w9003_,
		_w9004_
	);
	LUT2 #(
		.INIT('h1)
	) name6859 (
		\u13_ints_r_reg[7]/NET0131 ,
		\u18_int_set_reg[2]/NET0131 ,
		_w9005_
	);
	LUT2 #(
		.INIT('h1)
	) name6860 (
		_w2743_,
		_w9005_,
		_w9006_
	);
	LUT2 #(
		.INIT('h1)
	) name6861 (
		\u13_ints_r_reg[9]/NET0131 ,
		\u19_int_set_reg[1]/NET0131 ,
		_w9007_
	);
	LUT2 #(
		.INIT('h1)
	) name6862 (
		_w2743_,
		_w9007_,
		_w9008_
	);
	LUT2 #(
		.INIT('h1)
	) name6863 (
		\u9_rp_reg[2]/P0001 ,
		\u9_wp_reg[3]/P0001 ,
		_w9009_
	);
	LUT2 #(
		.INIT('h8)
	) name6864 (
		\u9_rp_reg[2]/P0001 ,
		\u9_wp_reg[3]/P0001 ,
		_w9010_
	);
	LUT2 #(
		.INIT('h1)
	) name6865 (
		_w9009_,
		_w9010_,
		_w9011_
	);
	LUT2 #(
		.INIT('h4)
	) name6866 (
		\u9_rp_reg[0]/P0001 ,
		\u9_wp_reg[1]/P0001 ,
		_w9012_
	);
	LUT2 #(
		.INIT('h1)
	) name6867 (
		_w8957_,
		_w9012_,
		_w9013_
	);
	LUT2 #(
		.INIT('h8)
	) name6868 (
		_w8960_,
		_w9013_,
		_w9014_
	);
	LUT2 #(
		.INIT('h2)
	) name6869 (
		_w3312_,
		_w9011_,
		_w9015_
	);
	LUT2 #(
		.INIT('h8)
	) name6870 (
		_w9014_,
		_w9015_,
		_w9016_
	);
	LUT2 #(
		.INIT('h1)
	) name6871 (
		\wb_addr_i[29]_pad ,
		\wb_addr_i[30]_pad ,
		_w9017_
	);
	LUT2 #(
		.INIT('h4)
	) name6872 (
		\wb_addr_i[31]_pad ,
		_w9017_,
		_w9018_
	);
	LUT2 #(
		.INIT('h8)
	) name6873 (
		_w8777_,
		_w9018_,
		_w9019_
	);
	LUT2 #(
		.INIT('h4)
	) name6874 (
		_w8779_,
		_w9019_,
		_w9020_
	);
	LUT2 #(
		.INIT('h2)
	) name6875 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[4]/NET0131 ,
		_w9021_
	);
	LUT2 #(
		.INIT('h4)
	) name6876 (
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[6]/NET0131 ,
		_w9022_
	);
	LUT2 #(
		.INIT('h8)
	) name6877 (
		_w9021_,
		_w9022_,
		_w9023_
	);
	LUT2 #(
		.INIT('h1)
	) name6878 (
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w9024_
	);
	LUT2 #(
		.INIT('h2)
	) name6879 (
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w9025_
	);
	LUT2 #(
		.INIT('h8)
	) name6880 (
		_w9024_,
		_w9025_,
		_w9026_
	);
	LUT2 #(
		.INIT('h8)
	) name6881 (
		_w9023_,
		_w9026_,
		_w9027_
	);
	LUT2 #(
		.INIT('h1)
	) name6882 (
		\u10_rp_reg[2]/P0001 ,
		\u10_wp_reg[3]/P0001 ,
		_w9028_
	);
	LUT2 #(
		.INIT('h8)
	) name6883 (
		\u10_rp_reg[2]/P0001 ,
		\u10_wp_reg[3]/P0001 ,
		_w9029_
	);
	LUT2 #(
		.INIT('h1)
	) name6884 (
		_w9028_,
		_w9029_,
		_w9030_
	);
	LUT2 #(
		.INIT('h4)
	) name6885 (
		\u10_rp_reg[0]/P0001 ,
		\u10_wp_reg[1]/P0001 ,
		_w9031_
	);
	LUT2 #(
		.INIT('h1)
	) name6886 (
		_w8964_,
		_w9031_,
		_w9032_
	);
	LUT2 #(
		.INIT('h8)
	) name6887 (
		_w8967_,
		_w9032_,
		_w9033_
	);
	LUT2 #(
		.INIT('h2)
	) name6888 (
		_w3502_,
		_w9030_,
		_w9034_
	);
	LUT2 #(
		.INIT('h8)
	) name6889 (
		_w9033_,
		_w9034_,
		_w9035_
	);
	LUT2 #(
		.INIT('h1)
	) name6890 (
		\u11_rp_reg[2]/P0001 ,
		\u11_wp_reg[3]/P0001 ,
		_w9036_
	);
	LUT2 #(
		.INIT('h8)
	) name6891 (
		\u11_rp_reg[2]/P0001 ,
		\u11_wp_reg[3]/P0001 ,
		_w9037_
	);
	LUT2 #(
		.INIT('h1)
	) name6892 (
		_w9036_,
		_w9037_,
		_w9038_
	);
	LUT2 #(
		.INIT('h4)
	) name6893 (
		\u11_rp_reg[0]/P0001 ,
		\u11_wp_reg[1]/P0001 ,
		_w9039_
	);
	LUT2 #(
		.INIT('h1)
	) name6894 (
		_w8950_,
		_w9039_,
		_w9040_
	);
	LUT2 #(
		.INIT('h8)
	) name6895 (
		_w8953_,
		_w9040_,
		_w9041_
	);
	LUT2 #(
		.INIT('h2)
	) name6896 (
		_w3065_,
		_w9038_,
		_w9042_
	);
	LUT2 #(
		.INIT('h8)
	) name6897 (
		_w9041_,
		_w9042_,
		_w9043_
	);
	LUT2 #(
		.INIT('h1)
	) name6898 (
		\u2_cnt_reg[5]/NET0131 ,
		_w6472_,
		_w9044_
	);
	LUT2 #(
		.INIT('h8)
	) name6899 (
		\u2_cnt_reg[5]/NET0131 ,
		_w6472_,
		_w9045_
	);
	LUT2 #(
		.INIT('h1)
	) name6900 (
		_w9044_,
		_w9045_,
		_w9046_
	);
	LUT2 #(
		.INIT('h1)
	) name6901 (
		suspended_o_pad,
		_w9046_,
		_w9047_
	);
	LUT2 #(
		.INIT('h1)
	) name6902 (
		\u2_cnt_reg[6]/NET0131 ,
		_w9045_,
		_w9048_
	);
	LUT2 #(
		.INIT('h1)
	) name6903 (
		_w6474_,
		_w9048_,
		_w9049_
	);
	LUT2 #(
		.INIT('h1)
	) name6904 (
		suspended_o_pad,
		_w9049_,
		_w9050_
	);
	LUT2 #(
		.INIT('h1)
	) name6905 (
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[2]/NET0131 ,
		_w9051_
	);
	LUT2 #(
		.INIT('h8)
	) name6906 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w9052_
	);
	LUT2 #(
		.INIT('h8)
	) name6907 (
		_w9051_,
		_w9052_,
		_w9053_
	);
	LUT2 #(
		.INIT('h1)
	) name6908 (
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w9054_
	);
	LUT2 #(
		.INIT('h4)
	) name6909 (
		\u2_cnt_reg[6]/NET0131 ,
		_w9054_,
		_w9055_
	);
	LUT2 #(
		.INIT('h8)
	) name6910 (
		\u2_cnt_reg[7]/NET0131 ,
		_w9053_,
		_w9056_
	);
	LUT2 #(
		.INIT('h8)
	) name6911 (
		_w9055_,
		_w9056_,
		_w9057_
	);
	LUT2 #(
		.INIT('h1)
	) name6912 (
		\u2_cnt_reg[6]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w9058_
	);
	LUT2 #(
		.INIT('h8)
	) name6913 (
		_w9054_,
		_w9058_,
		_w9059_
	);
	LUT2 #(
		.INIT('h1)
	) name6914 (
		\u2_to_cnt_reg[2]/NET0131 ,
		\u2_to_cnt_reg[3]/NET0131 ,
		_w9060_
	);
	LUT2 #(
		.INIT('h4)
	) name6915 (
		\u2_to_cnt_reg[4]/NET0131 ,
		\u2_to_cnt_reg[5]/NET0131 ,
		_w9061_
	);
	LUT2 #(
		.INIT('h8)
	) name6916 (
		_w9060_,
		_w9061_,
		_w9062_
	);
	LUT2 #(
		.INIT('h2)
	) name6917 (
		\u2_to_cnt_reg[0]/NET0131 ,
		\u2_to_cnt_reg[1]/NET0131 ,
		_w9063_
	);
	LUT2 #(
		.INIT('h8)
	) name6918 (
		_w9062_,
		_w9063_,
		_w9064_
	);
	LUT2 #(
		.INIT('h2)
	) name6919 (
		\u2_to_cnt_reg[0]/NET0131 ,
		_w9064_,
		_w9065_
	);
	LUT2 #(
		.INIT('h1)
	) name6920 (
		\u2_bit_clk_e_reg/P0001 ,
		_w9065_,
		_w9066_
	);
	LUT2 #(
		.INIT('h2)
	) name6921 (
		\u2_to_cnt_reg[0]/NET0131 ,
		_w9062_,
		_w9067_
	);
	LUT2 #(
		.INIT('h1)
	) name6922 (
		\u2_to_cnt_reg[1]/NET0131 ,
		_w9067_,
		_w9068_
	);
	LUT2 #(
		.INIT('h1)
	) name6923 (
		\u2_bit_clk_e_reg/P0001 ,
		_w6479_,
		_w9069_
	);
	LUT2 #(
		.INIT('h4)
	) name6924 (
		_w9068_,
		_w9069_,
		_w9070_
	);
	LUT2 #(
		.INIT('h8)
	) name6925 (
		_w9030_,
		_w9033_,
		_w9071_
	);
	LUT2 #(
		.INIT('h8)
	) name6926 (
		_w9038_,
		_w9041_,
		_w9072_
	);
	LUT2 #(
		.INIT('h8)
	) name6927 (
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w9073_
	);
	LUT2 #(
		.INIT('h1)
	) name6928 (
		\u2_cnt_reg[5]/NET0131 ,
		\u2_cnt_reg[7]/NET0131 ,
		_w9074_
	);
	LUT2 #(
		.INIT('h8)
	) name6929 (
		_w9073_,
		_w9074_,
		_w9075_
	);
	LUT2 #(
		.INIT('h8)
	) name6930 (
		_w9023_,
		_w9075_,
		_w9076_
	);
	LUT2 #(
		.INIT('h8)
	) name6931 (
		_w9011_,
		_w9014_,
		_w9077_
	);
	LUT2 #(
		.INIT('h1)
	) name6932 (
		\u2_cnt_reg[1]/NET0131 ,
		\u2_cnt_reg[3]/NET0131 ,
		_w9078_
	);
	LUT2 #(
		.INIT('h4)
	) name6933 (
		\u2_cnt_reg[2]/NET0131 ,
		_w9078_,
		_w9079_
	);
	LUT2 #(
		.INIT('h4)
	) name6934 (
		\u2_cnt_reg[4]/NET0131 ,
		_w9079_,
		_w9080_
	);
	LUT2 #(
		.INIT('h2)
	) name6935 (
		_w6473_,
		_w9080_,
		_w9081_
	);
	LUT2 #(
		.INIT('h1)
	) name6936 (
		\u2_cnt_reg[7]/NET0131 ,
		_w9081_,
		_w9082_
	);
	LUT2 #(
		.INIT('h8)
	) name6937 (
		_w2738_,
		_w6168_,
		_w9083_
	);
	LUT2 #(
		.INIT('h8)
	) name6938 (
		_w2738_,
		_w6170_,
		_w9084_
	);
	LUT2 #(
		.INIT('h2)
	) name6939 (
		\u2_cnt_reg[3]/NET0131 ,
		_w9051_,
		_w9085_
	);
	LUT2 #(
		.INIT('h8)
	) name6940 (
		\u2_cnt_reg[4]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w9086_
	);
	LUT2 #(
		.INIT('h8)
	) name6941 (
		_w9085_,
		_w9086_,
		_w9087_
	);
	LUT2 #(
		.INIT('h2)
	) name6942 (
		_w9058_,
		_w9087_,
		_w9088_
	);
	LUT2 #(
		.INIT('h4)
	) name6943 (
		suspended_o_pad,
		\u2_cnt_reg[0]/NET0131 ,
		_w9089_
	);
	LUT2 #(
		.INIT('h1)
	) name6944 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[1]/NET0131 ,
		_w9090_
	);
	LUT2 #(
		.INIT('h1)
	) name6945 (
		_w6469_,
		_w9090_,
		_w9091_
	);
	LUT2 #(
		.INIT('h1)
	) name6946 (
		suspended_o_pad,
		_w9091_,
		_w9092_
	);
	LUT2 #(
		.INIT('h1)
	) name6947 (
		\u2_cnt_reg[2]/NET0131 ,
		_w6469_,
		_w9093_
	);
	LUT2 #(
		.INIT('h1)
	) name6948 (
		_w6470_,
		_w9093_,
		_w9094_
	);
	LUT2 #(
		.INIT('h1)
	) name6949 (
		suspended_o_pad,
		_w9094_,
		_w9095_
	);
	LUT2 #(
		.INIT('h2)
	) name6950 (
		_w9055_,
		_w9085_,
		_w9096_
	);
	LUT2 #(
		.INIT('h2)
	) name6951 (
		\u2_cnt_reg[7]/NET0131 ,
		_w9096_,
		_w9097_
	);
	LUT2 #(
		.INIT('h4)
	) name6952 (
		\u2_cnt_reg[0]/NET0131 ,
		_w9059_,
		_w9098_
	);
	LUT2 #(
		.INIT('h8)
	) name6953 (
		_w9079_,
		_w9098_,
		_w9099_
	);
	LUT2 #(
		.INIT('h8)
	) name6954 (
		\u2_cnt_reg[2]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w9100_
	);
	LUT2 #(
		.INIT('h8)
	) name6955 (
		_w9021_,
		_w9100_,
		_w9101_
	);
	LUT2 #(
		.INIT('h8)
	) name6956 (
		_w9058_,
		_w9078_,
		_w9102_
	);
	LUT2 #(
		.INIT('h8)
	) name6957 (
		_w9101_,
		_w9102_,
		_w9103_
	);
	LUT2 #(
		.INIT('h8)
	) name6958 (
		_w2738_,
		_w6145_,
		_w9104_
	);
	LUT2 #(
		.INIT('h8)
	) name6959 (
		\u2_cnt_reg[1]/NET0131 ,
		_w9073_,
		_w9105_
	);
	LUT2 #(
		.INIT('h2)
	) name6960 (
		_w9054_,
		_w9105_,
		_w9106_
	);
	LUT2 #(
		.INIT('h2)
	) name6961 (
		\u2_cnt_reg[6]/NET0131 ,
		_w9106_,
		_w9107_
	);
	LUT2 #(
		.INIT('h1)
	) name6962 (
		\u2_cnt_reg[7]/NET0131 ,
		_w9107_,
		_w9108_
	);
	LUT2 #(
		.INIT('h8)
	) name6963 (
		\u2_cnt_reg[4]/NET0131 ,
		_w9058_,
		_w9109_
	);
	LUT2 #(
		.INIT('h8)
	) name6964 (
		\u2_cnt_reg[5]/NET0131 ,
		_w9053_,
		_w9110_
	);
	LUT2 #(
		.INIT('h8)
	) name6965 (
		_w9109_,
		_w9110_,
		_w9111_
	);
	LUT2 #(
		.INIT('h2)
	) name6966 (
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w9112_
	);
	LUT2 #(
		.INIT('h8)
	) name6967 (
		\u9_mem_reg[1][0]/P0001 ,
		_w9112_,
		_w9113_
	);
	LUT2 #(
		.INIT('h1)
	) name6968 (
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w9114_
	);
	LUT2 #(
		.INIT('h8)
	) name6969 (
		\u9_mem_reg[0][0]/P0001 ,
		_w9114_,
		_w9115_
	);
	LUT2 #(
		.INIT('h8)
	) name6970 (
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w9116_
	);
	LUT2 #(
		.INIT('h8)
	) name6971 (
		\u9_mem_reg[3][0]/P0001 ,
		_w9116_,
		_w9117_
	);
	LUT2 #(
		.INIT('h4)
	) name6972 (
		\u9_rp_reg[0]/P0001 ,
		\u9_rp_reg[1]/P0001 ,
		_w9118_
	);
	LUT2 #(
		.INIT('h8)
	) name6973 (
		\u9_mem_reg[2][0]/P0001 ,
		_w9118_,
		_w9119_
	);
	LUT2 #(
		.INIT('h1)
	) name6974 (
		_w9113_,
		_w9115_,
		_w9120_
	);
	LUT2 #(
		.INIT('h1)
	) name6975 (
		_w9117_,
		_w9119_,
		_w9121_
	);
	LUT2 #(
		.INIT('h8)
	) name6976 (
		_w9120_,
		_w9121_,
		_w9122_
	);
	LUT2 #(
		.INIT('h8)
	) name6977 (
		\u9_mem_reg[2][10]/P0001 ,
		_w9118_,
		_w9123_
	);
	LUT2 #(
		.INIT('h8)
	) name6978 (
		\u9_mem_reg[0][10]/P0001 ,
		_w9114_,
		_w9124_
	);
	LUT2 #(
		.INIT('h8)
	) name6979 (
		\u9_mem_reg[3][10]/P0001 ,
		_w9116_,
		_w9125_
	);
	LUT2 #(
		.INIT('h8)
	) name6980 (
		\u9_mem_reg[1][10]/P0001 ,
		_w9112_,
		_w9126_
	);
	LUT2 #(
		.INIT('h1)
	) name6981 (
		_w9123_,
		_w9124_,
		_w9127_
	);
	LUT2 #(
		.INIT('h1)
	) name6982 (
		_w9125_,
		_w9126_,
		_w9128_
	);
	LUT2 #(
		.INIT('h8)
	) name6983 (
		_w9127_,
		_w9128_,
		_w9129_
	);
	LUT2 #(
		.INIT('h8)
	) name6984 (
		\u9_mem_reg[1][11]/P0001 ,
		_w9112_,
		_w9130_
	);
	LUT2 #(
		.INIT('h8)
	) name6985 (
		\u9_mem_reg[0][11]/P0001 ,
		_w9114_,
		_w9131_
	);
	LUT2 #(
		.INIT('h8)
	) name6986 (
		\u9_mem_reg[3][11]/P0001 ,
		_w9116_,
		_w9132_
	);
	LUT2 #(
		.INIT('h8)
	) name6987 (
		\u9_mem_reg[2][11]/P0001 ,
		_w9118_,
		_w9133_
	);
	LUT2 #(
		.INIT('h1)
	) name6988 (
		_w9130_,
		_w9131_,
		_w9134_
	);
	LUT2 #(
		.INIT('h1)
	) name6989 (
		_w9132_,
		_w9133_,
		_w9135_
	);
	LUT2 #(
		.INIT('h8)
	) name6990 (
		_w9134_,
		_w9135_,
		_w9136_
	);
	LUT2 #(
		.INIT('h8)
	) name6991 (
		\u9_mem_reg[1][12]/P0001 ,
		_w9112_,
		_w9137_
	);
	LUT2 #(
		.INIT('h8)
	) name6992 (
		\u9_mem_reg[0][12]/P0001 ,
		_w9114_,
		_w9138_
	);
	LUT2 #(
		.INIT('h8)
	) name6993 (
		\u9_mem_reg[3][12]/P0001 ,
		_w9116_,
		_w9139_
	);
	LUT2 #(
		.INIT('h8)
	) name6994 (
		\u9_mem_reg[2][12]/P0001 ,
		_w9118_,
		_w9140_
	);
	LUT2 #(
		.INIT('h1)
	) name6995 (
		_w9137_,
		_w9138_,
		_w9141_
	);
	LUT2 #(
		.INIT('h1)
	) name6996 (
		_w9139_,
		_w9140_,
		_w9142_
	);
	LUT2 #(
		.INIT('h8)
	) name6997 (
		_w9141_,
		_w9142_,
		_w9143_
	);
	LUT2 #(
		.INIT('h8)
	) name6998 (
		\u9_mem_reg[1][13]/P0001 ,
		_w9112_,
		_w9144_
	);
	LUT2 #(
		.INIT('h8)
	) name6999 (
		\u9_mem_reg[0][13]/P0001 ,
		_w9114_,
		_w9145_
	);
	LUT2 #(
		.INIT('h8)
	) name7000 (
		\u9_mem_reg[3][13]/P0001 ,
		_w9116_,
		_w9146_
	);
	LUT2 #(
		.INIT('h8)
	) name7001 (
		\u9_mem_reg[2][13]/P0001 ,
		_w9118_,
		_w9147_
	);
	LUT2 #(
		.INIT('h1)
	) name7002 (
		_w9144_,
		_w9145_,
		_w9148_
	);
	LUT2 #(
		.INIT('h1)
	) name7003 (
		_w9146_,
		_w9147_,
		_w9149_
	);
	LUT2 #(
		.INIT('h8)
	) name7004 (
		_w9148_,
		_w9149_,
		_w9150_
	);
	LUT2 #(
		.INIT('h8)
	) name7005 (
		\u9_mem_reg[1][14]/P0001 ,
		_w9112_,
		_w9151_
	);
	LUT2 #(
		.INIT('h8)
	) name7006 (
		\u9_mem_reg[0][14]/P0001 ,
		_w9114_,
		_w9152_
	);
	LUT2 #(
		.INIT('h8)
	) name7007 (
		\u9_mem_reg[3][14]/P0001 ,
		_w9116_,
		_w9153_
	);
	LUT2 #(
		.INIT('h8)
	) name7008 (
		\u9_mem_reg[2][14]/P0001 ,
		_w9118_,
		_w9154_
	);
	LUT2 #(
		.INIT('h1)
	) name7009 (
		_w9151_,
		_w9152_,
		_w9155_
	);
	LUT2 #(
		.INIT('h1)
	) name7010 (
		_w9153_,
		_w9154_,
		_w9156_
	);
	LUT2 #(
		.INIT('h8)
	) name7011 (
		_w9155_,
		_w9156_,
		_w9157_
	);
	LUT2 #(
		.INIT('h8)
	) name7012 (
		\u9_mem_reg[1][15]/P0001 ,
		_w9112_,
		_w9158_
	);
	LUT2 #(
		.INIT('h8)
	) name7013 (
		\u9_mem_reg[0][15]/P0001 ,
		_w9114_,
		_w9159_
	);
	LUT2 #(
		.INIT('h8)
	) name7014 (
		\u9_mem_reg[3][15]/P0001 ,
		_w9116_,
		_w9160_
	);
	LUT2 #(
		.INIT('h8)
	) name7015 (
		\u9_mem_reg[2][15]/P0001 ,
		_w9118_,
		_w9161_
	);
	LUT2 #(
		.INIT('h1)
	) name7016 (
		_w9158_,
		_w9159_,
		_w9162_
	);
	LUT2 #(
		.INIT('h1)
	) name7017 (
		_w9160_,
		_w9161_,
		_w9163_
	);
	LUT2 #(
		.INIT('h8)
	) name7018 (
		_w9162_,
		_w9163_,
		_w9164_
	);
	LUT2 #(
		.INIT('h8)
	) name7019 (
		\u9_mem_reg[2][16]/P0001 ,
		_w9118_,
		_w9165_
	);
	LUT2 #(
		.INIT('h8)
	) name7020 (
		\u9_mem_reg[1][16]/P0001 ,
		_w9112_,
		_w9166_
	);
	LUT2 #(
		.INIT('h8)
	) name7021 (
		\u9_mem_reg[3][16]/P0001 ,
		_w9116_,
		_w9167_
	);
	LUT2 #(
		.INIT('h8)
	) name7022 (
		\u9_mem_reg[0][16]/P0001 ,
		_w9114_,
		_w9168_
	);
	LUT2 #(
		.INIT('h1)
	) name7023 (
		_w9165_,
		_w9166_,
		_w9169_
	);
	LUT2 #(
		.INIT('h1)
	) name7024 (
		_w9167_,
		_w9168_,
		_w9170_
	);
	LUT2 #(
		.INIT('h8)
	) name7025 (
		_w9169_,
		_w9170_,
		_w9171_
	);
	LUT2 #(
		.INIT('h8)
	) name7026 (
		\u9_mem_reg[1][17]/P0001 ,
		_w9112_,
		_w9172_
	);
	LUT2 #(
		.INIT('h8)
	) name7027 (
		\u9_mem_reg[0][17]/P0001 ,
		_w9114_,
		_w9173_
	);
	LUT2 #(
		.INIT('h8)
	) name7028 (
		\u9_mem_reg[3][17]/P0001 ,
		_w9116_,
		_w9174_
	);
	LUT2 #(
		.INIT('h8)
	) name7029 (
		\u9_mem_reg[2][17]/P0001 ,
		_w9118_,
		_w9175_
	);
	LUT2 #(
		.INIT('h1)
	) name7030 (
		_w9172_,
		_w9173_,
		_w9176_
	);
	LUT2 #(
		.INIT('h1)
	) name7031 (
		_w9174_,
		_w9175_,
		_w9177_
	);
	LUT2 #(
		.INIT('h8)
	) name7032 (
		_w9176_,
		_w9177_,
		_w9178_
	);
	LUT2 #(
		.INIT('h8)
	) name7033 (
		\u9_mem_reg[1][18]/P0001 ,
		_w9112_,
		_w9179_
	);
	LUT2 #(
		.INIT('h8)
	) name7034 (
		\u9_mem_reg[2][18]/P0001 ,
		_w9118_,
		_w9180_
	);
	LUT2 #(
		.INIT('h8)
	) name7035 (
		\u9_mem_reg[3][18]/P0001 ,
		_w9116_,
		_w9181_
	);
	LUT2 #(
		.INIT('h8)
	) name7036 (
		\u9_mem_reg[0][18]/P0001 ,
		_w9114_,
		_w9182_
	);
	LUT2 #(
		.INIT('h1)
	) name7037 (
		_w9179_,
		_w9180_,
		_w9183_
	);
	LUT2 #(
		.INIT('h1)
	) name7038 (
		_w9181_,
		_w9182_,
		_w9184_
	);
	LUT2 #(
		.INIT('h8)
	) name7039 (
		_w9183_,
		_w9184_,
		_w9185_
	);
	LUT2 #(
		.INIT('h8)
	) name7040 (
		\u9_mem_reg[2][19]/P0001 ,
		_w9118_,
		_w9186_
	);
	LUT2 #(
		.INIT('h8)
	) name7041 (
		\u9_mem_reg[1][19]/P0001 ,
		_w9112_,
		_w9187_
	);
	LUT2 #(
		.INIT('h8)
	) name7042 (
		\u9_mem_reg[3][19]/P0001 ,
		_w9116_,
		_w9188_
	);
	LUT2 #(
		.INIT('h8)
	) name7043 (
		\u9_mem_reg[0][19]/P0001 ,
		_w9114_,
		_w9189_
	);
	LUT2 #(
		.INIT('h1)
	) name7044 (
		_w9186_,
		_w9187_,
		_w9190_
	);
	LUT2 #(
		.INIT('h1)
	) name7045 (
		_w9188_,
		_w9189_,
		_w9191_
	);
	LUT2 #(
		.INIT('h8)
	) name7046 (
		_w9190_,
		_w9191_,
		_w9192_
	);
	LUT2 #(
		.INIT('h8)
	) name7047 (
		\u9_mem_reg[1][1]/P0001 ,
		_w9112_,
		_w9193_
	);
	LUT2 #(
		.INIT('h8)
	) name7048 (
		\u9_mem_reg[0][1]/P0001 ,
		_w9114_,
		_w9194_
	);
	LUT2 #(
		.INIT('h8)
	) name7049 (
		\u9_mem_reg[3][1]/P0001 ,
		_w9116_,
		_w9195_
	);
	LUT2 #(
		.INIT('h8)
	) name7050 (
		\u9_mem_reg[2][1]/P0001 ,
		_w9118_,
		_w9196_
	);
	LUT2 #(
		.INIT('h1)
	) name7051 (
		_w9193_,
		_w9194_,
		_w9197_
	);
	LUT2 #(
		.INIT('h1)
	) name7052 (
		_w9195_,
		_w9196_,
		_w9198_
	);
	LUT2 #(
		.INIT('h8)
	) name7053 (
		_w9197_,
		_w9198_,
		_w9199_
	);
	LUT2 #(
		.INIT('h8)
	) name7054 (
		\u9_mem_reg[0][20]/P0001 ,
		_w9114_,
		_w9200_
	);
	LUT2 #(
		.INIT('h8)
	) name7055 (
		\u9_mem_reg[2][20]/P0001 ,
		_w9118_,
		_w9201_
	);
	LUT2 #(
		.INIT('h8)
	) name7056 (
		\u9_mem_reg[3][20]/P0001 ,
		_w9116_,
		_w9202_
	);
	LUT2 #(
		.INIT('h8)
	) name7057 (
		\u9_mem_reg[1][20]/P0001 ,
		_w9112_,
		_w9203_
	);
	LUT2 #(
		.INIT('h1)
	) name7058 (
		_w9200_,
		_w9201_,
		_w9204_
	);
	LUT2 #(
		.INIT('h1)
	) name7059 (
		_w9202_,
		_w9203_,
		_w9205_
	);
	LUT2 #(
		.INIT('h8)
	) name7060 (
		_w9204_,
		_w9205_,
		_w9206_
	);
	LUT2 #(
		.INIT('h8)
	) name7061 (
		\u9_mem_reg[2][21]/P0001 ,
		_w9118_,
		_w9207_
	);
	LUT2 #(
		.INIT('h8)
	) name7062 (
		\u9_mem_reg[1][21]/P0001 ,
		_w9112_,
		_w9208_
	);
	LUT2 #(
		.INIT('h8)
	) name7063 (
		\u9_mem_reg[3][21]/P0001 ,
		_w9116_,
		_w9209_
	);
	LUT2 #(
		.INIT('h8)
	) name7064 (
		\u9_mem_reg[0][21]/P0001 ,
		_w9114_,
		_w9210_
	);
	LUT2 #(
		.INIT('h1)
	) name7065 (
		_w9207_,
		_w9208_,
		_w9211_
	);
	LUT2 #(
		.INIT('h1)
	) name7066 (
		_w9209_,
		_w9210_,
		_w9212_
	);
	LUT2 #(
		.INIT('h8)
	) name7067 (
		_w9211_,
		_w9212_,
		_w9213_
	);
	LUT2 #(
		.INIT('h8)
	) name7068 (
		\u9_mem_reg[2][22]/P0001 ,
		_w9118_,
		_w9214_
	);
	LUT2 #(
		.INIT('h8)
	) name7069 (
		\u9_mem_reg[1][22]/P0001 ,
		_w9112_,
		_w9215_
	);
	LUT2 #(
		.INIT('h8)
	) name7070 (
		\u9_mem_reg[3][22]/P0001 ,
		_w9116_,
		_w9216_
	);
	LUT2 #(
		.INIT('h8)
	) name7071 (
		\u9_mem_reg[0][22]/P0001 ,
		_w9114_,
		_w9217_
	);
	LUT2 #(
		.INIT('h1)
	) name7072 (
		_w9214_,
		_w9215_,
		_w9218_
	);
	LUT2 #(
		.INIT('h1)
	) name7073 (
		_w9216_,
		_w9217_,
		_w9219_
	);
	LUT2 #(
		.INIT('h8)
	) name7074 (
		_w9218_,
		_w9219_,
		_w9220_
	);
	LUT2 #(
		.INIT('h8)
	) name7075 (
		\u9_mem_reg[1][23]/P0001 ,
		_w9112_,
		_w9221_
	);
	LUT2 #(
		.INIT('h8)
	) name7076 (
		\u9_mem_reg[2][23]/P0001 ,
		_w9118_,
		_w9222_
	);
	LUT2 #(
		.INIT('h8)
	) name7077 (
		\u9_mem_reg[3][23]/P0001 ,
		_w9116_,
		_w9223_
	);
	LUT2 #(
		.INIT('h8)
	) name7078 (
		\u9_mem_reg[0][23]/P0001 ,
		_w9114_,
		_w9224_
	);
	LUT2 #(
		.INIT('h1)
	) name7079 (
		_w9221_,
		_w9222_,
		_w9225_
	);
	LUT2 #(
		.INIT('h1)
	) name7080 (
		_w9223_,
		_w9224_,
		_w9226_
	);
	LUT2 #(
		.INIT('h8)
	) name7081 (
		_w9225_,
		_w9226_,
		_w9227_
	);
	LUT2 #(
		.INIT('h8)
	) name7082 (
		\u9_mem_reg[2][24]/P0001 ,
		_w9118_,
		_w9228_
	);
	LUT2 #(
		.INIT('h8)
	) name7083 (
		\u9_mem_reg[1][24]/P0001 ,
		_w9112_,
		_w9229_
	);
	LUT2 #(
		.INIT('h8)
	) name7084 (
		\u9_mem_reg[3][24]/P0001 ,
		_w9116_,
		_w9230_
	);
	LUT2 #(
		.INIT('h8)
	) name7085 (
		\u9_mem_reg[0][24]/P0001 ,
		_w9114_,
		_w9231_
	);
	LUT2 #(
		.INIT('h1)
	) name7086 (
		_w9228_,
		_w9229_,
		_w9232_
	);
	LUT2 #(
		.INIT('h1)
	) name7087 (
		_w9230_,
		_w9231_,
		_w9233_
	);
	LUT2 #(
		.INIT('h8)
	) name7088 (
		_w9232_,
		_w9233_,
		_w9234_
	);
	LUT2 #(
		.INIT('h8)
	) name7089 (
		\u9_mem_reg[2][26]/P0001 ,
		_w9118_,
		_w9235_
	);
	LUT2 #(
		.INIT('h8)
	) name7090 (
		\u9_mem_reg[1][26]/P0001 ,
		_w9112_,
		_w9236_
	);
	LUT2 #(
		.INIT('h8)
	) name7091 (
		\u9_mem_reg[3][26]/P0001 ,
		_w9116_,
		_w9237_
	);
	LUT2 #(
		.INIT('h8)
	) name7092 (
		\u9_mem_reg[0][26]/P0001 ,
		_w9114_,
		_w9238_
	);
	LUT2 #(
		.INIT('h1)
	) name7093 (
		_w9235_,
		_w9236_,
		_w9239_
	);
	LUT2 #(
		.INIT('h1)
	) name7094 (
		_w9237_,
		_w9238_,
		_w9240_
	);
	LUT2 #(
		.INIT('h8)
	) name7095 (
		_w9239_,
		_w9240_,
		_w9241_
	);
	LUT2 #(
		.INIT('h8)
	) name7096 (
		\u9_mem_reg[2][27]/P0001 ,
		_w9118_,
		_w9242_
	);
	LUT2 #(
		.INIT('h8)
	) name7097 (
		\u9_mem_reg[1][27]/P0001 ,
		_w9112_,
		_w9243_
	);
	LUT2 #(
		.INIT('h8)
	) name7098 (
		\u9_mem_reg[3][27]/P0001 ,
		_w9116_,
		_w9244_
	);
	LUT2 #(
		.INIT('h8)
	) name7099 (
		\u9_mem_reg[0][27]/P0001 ,
		_w9114_,
		_w9245_
	);
	LUT2 #(
		.INIT('h1)
	) name7100 (
		_w9242_,
		_w9243_,
		_w9246_
	);
	LUT2 #(
		.INIT('h1)
	) name7101 (
		_w9244_,
		_w9245_,
		_w9247_
	);
	LUT2 #(
		.INIT('h8)
	) name7102 (
		_w9246_,
		_w9247_,
		_w9248_
	);
	LUT2 #(
		.INIT('h8)
	) name7103 (
		\u9_mem_reg[2][28]/P0001 ,
		_w9118_,
		_w9249_
	);
	LUT2 #(
		.INIT('h8)
	) name7104 (
		\u9_mem_reg[1][28]/P0001 ,
		_w9112_,
		_w9250_
	);
	LUT2 #(
		.INIT('h8)
	) name7105 (
		\u9_mem_reg[3][28]/P0001 ,
		_w9116_,
		_w9251_
	);
	LUT2 #(
		.INIT('h8)
	) name7106 (
		\u9_mem_reg[0][28]/P0001 ,
		_w9114_,
		_w9252_
	);
	LUT2 #(
		.INIT('h1)
	) name7107 (
		_w9249_,
		_w9250_,
		_w9253_
	);
	LUT2 #(
		.INIT('h1)
	) name7108 (
		_w9251_,
		_w9252_,
		_w9254_
	);
	LUT2 #(
		.INIT('h8)
	) name7109 (
		_w9253_,
		_w9254_,
		_w9255_
	);
	LUT2 #(
		.INIT('h8)
	) name7110 (
		\u9_mem_reg[1][29]/P0001 ,
		_w9112_,
		_w9256_
	);
	LUT2 #(
		.INIT('h8)
	) name7111 (
		\u9_mem_reg[2][29]/P0001 ,
		_w9118_,
		_w9257_
	);
	LUT2 #(
		.INIT('h8)
	) name7112 (
		\u9_mem_reg[3][29]/P0001 ,
		_w9116_,
		_w9258_
	);
	LUT2 #(
		.INIT('h8)
	) name7113 (
		\u9_mem_reg[0][29]/P0001 ,
		_w9114_,
		_w9259_
	);
	LUT2 #(
		.INIT('h1)
	) name7114 (
		_w9256_,
		_w9257_,
		_w9260_
	);
	LUT2 #(
		.INIT('h1)
	) name7115 (
		_w9258_,
		_w9259_,
		_w9261_
	);
	LUT2 #(
		.INIT('h8)
	) name7116 (
		_w9260_,
		_w9261_,
		_w9262_
	);
	LUT2 #(
		.INIT('h8)
	) name7117 (
		\u9_mem_reg[1][2]/P0001 ,
		_w9112_,
		_w9263_
	);
	LUT2 #(
		.INIT('h8)
	) name7118 (
		\u9_mem_reg[0][2]/P0001 ,
		_w9114_,
		_w9264_
	);
	LUT2 #(
		.INIT('h8)
	) name7119 (
		\u9_mem_reg[3][2]/P0001 ,
		_w9116_,
		_w9265_
	);
	LUT2 #(
		.INIT('h8)
	) name7120 (
		\u9_mem_reg[2][2]/P0001 ,
		_w9118_,
		_w9266_
	);
	LUT2 #(
		.INIT('h1)
	) name7121 (
		_w9263_,
		_w9264_,
		_w9267_
	);
	LUT2 #(
		.INIT('h1)
	) name7122 (
		_w9265_,
		_w9266_,
		_w9268_
	);
	LUT2 #(
		.INIT('h8)
	) name7123 (
		_w9267_,
		_w9268_,
		_w9269_
	);
	LUT2 #(
		.INIT('h8)
	) name7124 (
		\u9_mem_reg[2][30]/P0001 ,
		_w9118_,
		_w9270_
	);
	LUT2 #(
		.INIT('h8)
	) name7125 (
		\u9_mem_reg[1][30]/P0001 ,
		_w9112_,
		_w9271_
	);
	LUT2 #(
		.INIT('h8)
	) name7126 (
		\u9_mem_reg[3][30]/P0001 ,
		_w9116_,
		_w9272_
	);
	LUT2 #(
		.INIT('h8)
	) name7127 (
		\u9_mem_reg[0][30]/P0001 ,
		_w9114_,
		_w9273_
	);
	LUT2 #(
		.INIT('h1)
	) name7128 (
		_w9270_,
		_w9271_,
		_w9274_
	);
	LUT2 #(
		.INIT('h1)
	) name7129 (
		_w9272_,
		_w9273_,
		_w9275_
	);
	LUT2 #(
		.INIT('h8)
	) name7130 (
		_w9274_,
		_w9275_,
		_w9276_
	);
	LUT2 #(
		.INIT('h8)
	) name7131 (
		\u9_mem_reg[2][31]/P0001 ,
		_w9118_,
		_w9277_
	);
	LUT2 #(
		.INIT('h8)
	) name7132 (
		\u9_mem_reg[1][31]/P0001 ,
		_w9112_,
		_w9278_
	);
	LUT2 #(
		.INIT('h8)
	) name7133 (
		\u9_mem_reg[3][31]/P0001 ,
		_w9116_,
		_w9279_
	);
	LUT2 #(
		.INIT('h8)
	) name7134 (
		\u9_mem_reg[0][31]/P0001 ,
		_w9114_,
		_w9280_
	);
	LUT2 #(
		.INIT('h1)
	) name7135 (
		_w9277_,
		_w9278_,
		_w9281_
	);
	LUT2 #(
		.INIT('h1)
	) name7136 (
		_w9279_,
		_w9280_,
		_w9282_
	);
	LUT2 #(
		.INIT('h8)
	) name7137 (
		_w9281_,
		_w9282_,
		_w9283_
	);
	LUT2 #(
		.INIT('h8)
	) name7138 (
		\u9_mem_reg[1][3]/P0001 ,
		_w9112_,
		_w9284_
	);
	LUT2 #(
		.INIT('h8)
	) name7139 (
		\u9_mem_reg[0][3]/P0001 ,
		_w9114_,
		_w9285_
	);
	LUT2 #(
		.INIT('h8)
	) name7140 (
		\u9_mem_reg[3][3]/P0001 ,
		_w9116_,
		_w9286_
	);
	LUT2 #(
		.INIT('h8)
	) name7141 (
		\u9_mem_reg[2][3]/P0001 ,
		_w9118_,
		_w9287_
	);
	LUT2 #(
		.INIT('h1)
	) name7142 (
		_w9284_,
		_w9285_,
		_w9288_
	);
	LUT2 #(
		.INIT('h1)
	) name7143 (
		_w9286_,
		_w9287_,
		_w9289_
	);
	LUT2 #(
		.INIT('h8)
	) name7144 (
		_w9288_,
		_w9289_,
		_w9290_
	);
	LUT2 #(
		.INIT('h8)
	) name7145 (
		\u9_mem_reg[1][5]/P0001 ,
		_w9112_,
		_w9291_
	);
	LUT2 #(
		.INIT('h8)
	) name7146 (
		\u9_mem_reg[0][5]/P0001 ,
		_w9114_,
		_w9292_
	);
	LUT2 #(
		.INIT('h8)
	) name7147 (
		\u9_mem_reg[3][5]/P0001 ,
		_w9116_,
		_w9293_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		\u9_mem_reg[2][5]/P0001 ,
		_w9118_,
		_w9294_
	);
	LUT2 #(
		.INIT('h1)
	) name7149 (
		_w9291_,
		_w9292_,
		_w9295_
	);
	LUT2 #(
		.INIT('h1)
	) name7150 (
		_w9293_,
		_w9294_,
		_w9296_
	);
	LUT2 #(
		.INIT('h8)
	) name7151 (
		_w9295_,
		_w9296_,
		_w9297_
	);
	LUT2 #(
		.INIT('h8)
	) name7152 (
		\u9_mem_reg[2][6]/P0001 ,
		_w9118_,
		_w9298_
	);
	LUT2 #(
		.INIT('h8)
	) name7153 (
		\u9_mem_reg[1][6]/P0001 ,
		_w9112_,
		_w9299_
	);
	LUT2 #(
		.INIT('h8)
	) name7154 (
		\u9_mem_reg[3][6]/P0001 ,
		_w9116_,
		_w9300_
	);
	LUT2 #(
		.INIT('h8)
	) name7155 (
		\u9_mem_reg[0][6]/P0001 ,
		_w9114_,
		_w9301_
	);
	LUT2 #(
		.INIT('h1)
	) name7156 (
		_w9298_,
		_w9299_,
		_w9302_
	);
	LUT2 #(
		.INIT('h1)
	) name7157 (
		_w9300_,
		_w9301_,
		_w9303_
	);
	LUT2 #(
		.INIT('h8)
	) name7158 (
		_w9302_,
		_w9303_,
		_w9304_
	);
	LUT2 #(
		.INIT('h8)
	) name7159 (
		\u9_mem_reg[2][7]/P0001 ,
		_w9118_,
		_w9305_
	);
	LUT2 #(
		.INIT('h8)
	) name7160 (
		\u9_mem_reg[0][7]/P0001 ,
		_w9114_,
		_w9306_
	);
	LUT2 #(
		.INIT('h8)
	) name7161 (
		\u9_mem_reg[3][7]/P0001 ,
		_w9116_,
		_w9307_
	);
	LUT2 #(
		.INIT('h8)
	) name7162 (
		\u9_mem_reg[1][7]/P0001 ,
		_w9112_,
		_w9308_
	);
	LUT2 #(
		.INIT('h1)
	) name7163 (
		_w9305_,
		_w9306_,
		_w9309_
	);
	LUT2 #(
		.INIT('h1)
	) name7164 (
		_w9307_,
		_w9308_,
		_w9310_
	);
	LUT2 #(
		.INIT('h8)
	) name7165 (
		_w9309_,
		_w9310_,
		_w9311_
	);
	LUT2 #(
		.INIT('h4)
	) name7166 (
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w9312_
	);
	LUT2 #(
		.INIT('h8)
	) name7167 (
		\u10_mem_reg[2][0]/P0001 ,
		_w9312_,
		_w9313_
	);
	LUT2 #(
		.INIT('h1)
	) name7168 (
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w9314_
	);
	LUT2 #(
		.INIT('h8)
	) name7169 (
		\u10_mem_reg[0][0]/P0001 ,
		_w9314_,
		_w9315_
	);
	LUT2 #(
		.INIT('h8)
	) name7170 (
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w9316_
	);
	LUT2 #(
		.INIT('h8)
	) name7171 (
		\u10_mem_reg[3][0]/P0001 ,
		_w9316_,
		_w9317_
	);
	LUT2 #(
		.INIT('h2)
	) name7172 (
		\u10_rp_reg[0]/P0001 ,
		\u10_rp_reg[1]/P0001 ,
		_w9318_
	);
	LUT2 #(
		.INIT('h8)
	) name7173 (
		\u10_mem_reg[1][0]/P0001 ,
		_w9318_,
		_w9319_
	);
	LUT2 #(
		.INIT('h1)
	) name7174 (
		_w9313_,
		_w9315_,
		_w9320_
	);
	LUT2 #(
		.INIT('h1)
	) name7175 (
		_w9317_,
		_w9319_,
		_w9321_
	);
	LUT2 #(
		.INIT('h8)
	) name7176 (
		_w9320_,
		_w9321_,
		_w9322_
	);
	LUT2 #(
		.INIT('h8)
	) name7177 (
		\u9_mem_reg[1][25]/P0001 ,
		_w9112_,
		_w9323_
	);
	LUT2 #(
		.INIT('h8)
	) name7178 (
		\u9_mem_reg[2][25]/P0001 ,
		_w9118_,
		_w9324_
	);
	LUT2 #(
		.INIT('h8)
	) name7179 (
		\u9_mem_reg[3][25]/P0001 ,
		_w9116_,
		_w9325_
	);
	LUT2 #(
		.INIT('h8)
	) name7180 (
		\u9_mem_reg[0][25]/P0001 ,
		_w9114_,
		_w9326_
	);
	LUT2 #(
		.INIT('h1)
	) name7181 (
		_w9323_,
		_w9324_,
		_w9327_
	);
	LUT2 #(
		.INIT('h1)
	) name7182 (
		_w9325_,
		_w9326_,
		_w9328_
	);
	LUT2 #(
		.INIT('h8)
	) name7183 (
		_w9327_,
		_w9328_,
		_w9329_
	);
	LUT2 #(
		.INIT('h8)
	) name7184 (
		\u10_mem_reg[1][11]/P0001 ,
		_w9318_,
		_w9330_
	);
	LUT2 #(
		.INIT('h8)
	) name7185 (
		\u10_mem_reg[0][11]/P0001 ,
		_w9314_,
		_w9331_
	);
	LUT2 #(
		.INIT('h8)
	) name7186 (
		\u10_mem_reg[3][11]/P0001 ,
		_w9316_,
		_w9332_
	);
	LUT2 #(
		.INIT('h8)
	) name7187 (
		\u10_mem_reg[2][11]/P0001 ,
		_w9312_,
		_w9333_
	);
	LUT2 #(
		.INIT('h1)
	) name7188 (
		_w9330_,
		_w9331_,
		_w9334_
	);
	LUT2 #(
		.INIT('h1)
	) name7189 (
		_w9332_,
		_w9333_,
		_w9335_
	);
	LUT2 #(
		.INIT('h8)
	) name7190 (
		_w9334_,
		_w9335_,
		_w9336_
	);
	LUT2 #(
		.INIT('h8)
	) name7191 (
		\u10_mem_reg[1][12]/P0001 ,
		_w9318_,
		_w9337_
	);
	LUT2 #(
		.INIT('h8)
	) name7192 (
		\u10_mem_reg[0][12]/P0001 ,
		_w9314_,
		_w9338_
	);
	LUT2 #(
		.INIT('h8)
	) name7193 (
		\u10_mem_reg[3][12]/P0001 ,
		_w9316_,
		_w9339_
	);
	LUT2 #(
		.INIT('h8)
	) name7194 (
		\u10_mem_reg[2][12]/P0001 ,
		_w9312_,
		_w9340_
	);
	LUT2 #(
		.INIT('h1)
	) name7195 (
		_w9337_,
		_w9338_,
		_w9341_
	);
	LUT2 #(
		.INIT('h1)
	) name7196 (
		_w9339_,
		_w9340_,
		_w9342_
	);
	LUT2 #(
		.INIT('h8)
	) name7197 (
		_w9341_,
		_w9342_,
		_w9343_
	);
	LUT2 #(
		.INIT('h8)
	) name7198 (
		\u10_mem_reg[2][13]/P0001 ,
		_w9312_,
		_w9344_
	);
	LUT2 #(
		.INIT('h8)
	) name7199 (
		\u10_mem_reg[0][13]/P0001 ,
		_w9314_,
		_w9345_
	);
	LUT2 #(
		.INIT('h8)
	) name7200 (
		\u10_mem_reg[3][13]/P0001 ,
		_w9316_,
		_w9346_
	);
	LUT2 #(
		.INIT('h8)
	) name7201 (
		\u10_mem_reg[1][13]/P0001 ,
		_w9318_,
		_w9347_
	);
	LUT2 #(
		.INIT('h1)
	) name7202 (
		_w9344_,
		_w9345_,
		_w9348_
	);
	LUT2 #(
		.INIT('h1)
	) name7203 (
		_w9346_,
		_w9347_,
		_w9349_
	);
	LUT2 #(
		.INIT('h8)
	) name7204 (
		_w9348_,
		_w9349_,
		_w9350_
	);
	LUT2 #(
		.INIT('h8)
	) name7205 (
		\u10_mem_reg[2][15]/P0001 ,
		_w9312_,
		_w9351_
	);
	LUT2 #(
		.INIT('h8)
	) name7206 (
		\u10_mem_reg[0][15]/P0001 ,
		_w9314_,
		_w9352_
	);
	LUT2 #(
		.INIT('h8)
	) name7207 (
		\u10_mem_reg[3][15]/P0001 ,
		_w9316_,
		_w9353_
	);
	LUT2 #(
		.INIT('h8)
	) name7208 (
		\u10_mem_reg[1][15]/P0001 ,
		_w9318_,
		_w9354_
	);
	LUT2 #(
		.INIT('h1)
	) name7209 (
		_w9351_,
		_w9352_,
		_w9355_
	);
	LUT2 #(
		.INIT('h1)
	) name7210 (
		_w9353_,
		_w9354_,
		_w9356_
	);
	LUT2 #(
		.INIT('h8)
	) name7211 (
		_w9355_,
		_w9356_,
		_w9357_
	);
	LUT2 #(
		.INIT('h8)
	) name7212 (
		\u10_mem_reg[1][16]/P0001 ,
		_w9318_,
		_w9358_
	);
	LUT2 #(
		.INIT('h8)
	) name7213 (
		\u10_mem_reg[0][16]/P0001 ,
		_w9314_,
		_w9359_
	);
	LUT2 #(
		.INIT('h8)
	) name7214 (
		\u10_mem_reg[3][16]/P0001 ,
		_w9316_,
		_w9360_
	);
	LUT2 #(
		.INIT('h8)
	) name7215 (
		\u10_mem_reg[2][16]/P0001 ,
		_w9312_,
		_w9361_
	);
	LUT2 #(
		.INIT('h1)
	) name7216 (
		_w9358_,
		_w9359_,
		_w9362_
	);
	LUT2 #(
		.INIT('h1)
	) name7217 (
		_w9360_,
		_w9361_,
		_w9363_
	);
	LUT2 #(
		.INIT('h8)
	) name7218 (
		_w9362_,
		_w9363_,
		_w9364_
	);
	LUT2 #(
		.INIT('h8)
	) name7219 (
		\u10_mem_reg[2][17]/P0001 ,
		_w9312_,
		_w9365_
	);
	LUT2 #(
		.INIT('h8)
	) name7220 (
		\u10_mem_reg[1][17]/P0001 ,
		_w9318_,
		_w9366_
	);
	LUT2 #(
		.INIT('h8)
	) name7221 (
		\u10_mem_reg[3][17]/P0001 ,
		_w9316_,
		_w9367_
	);
	LUT2 #(
		.INIT('h8)
	) name7222 (
		\u10_mem_reg[0][17]/P0001 ,
		_w9314_,
		_w9368_
	);
	LUT2 #(
		.INIT('h1)
	) name7223 (
		_w9365_,
		_w9366_,
		_w9369_
	);
	LUT2 #(
		.INIT('h1)
	) name7224 (
		_w9367_,
		_w9368_,
		_w9370_
	);
	LUT2 #(
		.INIT('h8)
	) name7225 (
		_w9369_,
		_w9370_,
		_w9371_
	);
	LUT2 #(
		.INIT('h8)
	) name7226 (
		\u10_mem_reg[1][18]/P0001 ,
		_w9318_,
		_w9372_
	);
	LUT2 #(
		.INIT('h8)
	) name7227 (
		\u10_mem_reg[2][18]/P0001 ,
		_w9312_,
		_w9373_
	);
	LUT2 #(
		.INIT('h8)
	) name7228 (
		\u10_mem_reg[3][18]/P0001 ,
		_w9316_,
		_w9374_
	);
	LUT2 #(
		.INIT('h8)
	) name7229 (
		\u10_mem_reg[0][18]/P0001 ,
		_w9314_,
		_w9375_
	);
	LUT2 #(
		.INIT('h1)
	) name7230 (
		_w9372_,
		_w9373_,
		_w9376_
	);
	LUT2 #(
		.INIT('h1)
	) name7231 (
		_w9374_,
		_w9375_,
		_w9377_
	);
	LUT2 #(
		.INIT('h8)
	) name7232 (
		_w9376_,
		_w9377_,
		_w9378_
	);
	LUT2 #(
		.INIT('h8)
	) name7233 (
		\u10_mem_reg[0][19]/P0001 ,
		_w9314_,
		_w9379_
	);
	LUT2 #(
		.INIT('h8)
	) name7234 (
		\u10_mem_reg[2][19]/P0001 ,
		_w9312_,
		_w9380_
	);
	LUT2 #(
		.INIT('h8)
	) name7235 (
		\u10_mem_reg[3][19]/P0001 ,
		_w9316_,
		_w9381_
	);
	LUT2 #(
		.INIT('h8)
	) name7236 (
		\u10_mem_reg[1][19]/P0001 ,
		_w9318_,
		_w9382_
	);
	LUT2 #(
		.INIT('h1)
	) name7237 (
		_w9379_,
		_w9380_,
		_w9383_
	);
	LUT2 #(
		.INIT('h1)
	) name7238 (
		_w9381_,
		_w9382_,
		_w9384_
	);
	LUT2 #(
		.INIT('h8)
	) name7239 (
		_w9383_,
		_w9384_,
		_w9385_
	);
	LUT2 #(
		.INIT('h8)
	) name7240 (
		\u10_mem_reg[2][1]/P0001 ,
		_w9312_,
		_w9386_
	);
	LUT2 #(
		.INIT('h8)
	) name7241 (
		\u10_mem_reg[0][1]/P0001 ,
		_w9314_,
		_w9387_
	);
	LUT2 #(
		.INIT('h8)
	) name7242 (
		\u10_mem_reg[3][1]/P0001 ,
		_w9316_,
		_w9388_
	);
	LUT2 #(
		.INIT('h8)
	) name7243 (
		\u10_mem_reg[1][1]/P0001 ,
		_w9318_,
		_w9389_
	);
	LUT2 #(
		.INIT('h1)
	) name7244 (
		_w9386_,
		_w9387_,
		_w9390_
	);
	LUT2 #(
		.INIT('h1)
	) name7245 (
		_w9388_,
		_w9389_,
		_w9391_
	);
	LUT2 #(
		.INIT('h8)
	) name7246 (
		_w9390_,
		_w9391_,
		_w9392_
	);
	LUT2 #(
		.INIT('h2)
	) name7247 (
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w9393_
	);
	LUT2 #(
		.INIT('h8)
	) name7248 (
		\u11_mem_reg[1][6]/P0001 ,
		_w9393_,
		_w9394_
	);
	LUT2 #(
		.INIT('h1)
	) name7249 (
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w9395_
	);
	LUT2 #(
		.INIT('h8)
	) name7250 (
		\u11_mem_reg[0][6]/P0001 ,
		_w9395_,
		_w9396_
	);
	LUT2 #(
		.INIT('h8)
	) name7251 (
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w9397_
	);
	LUT2 #(
		.INIT('h8)
	) name7252 (
		\u11_mem_reg[3][6]/P0001 ,
		_w9397_,
		_w9398_
	);
	LUT2 #(
		.INIT('h4)
	) name7253 (
		\u11_rp_reg[0]/P0001 ,
		\u11_rp_reg[1]/P0001 ,
		_w9399_
	);
	LUT2 #(
		.INIT('h8)
	) name7254 (
		\u11_mem_reg[2][6]/P0001 ,
		_w9399_,
		_w9400_
	);
	LUT2 #(
		.INIT('h1)
	) name7255 (
		_w9394_,
		_w9396_,
		_w9401_
	);
	LUT2 #(
		.INIT('h1)
	) name7256 (
		_w9398_,
		_w9400_,
		_w9402_
	);
	LUT2 #(
		.INIT('h8)
	) name7257 (
		_w9401_,
		_w9402_,
		_w9403_
	);
	LUT2 #(
		.INIT('h8)
	) name7258 (
		\u10_mem_reg[0][20]/P0001 ,
		_w9314_,
		_w9404_
	);
	LUT2 #(
		.INIT('h8)
	) name7259 (
		\u10_mem_reg[2][20]/P0001 ,
		_w9312_,
		_w9405_
	);
	LUT2 #(
		.INIT('h8)
	) name7260 (
		\u10_mem_reg[3][20]/P0001 ,
		_w9316_,
		_w9406_
	);
	LUT2 #(
		.INIT('h8)
	) name7261 (
		\u10_mem_reg[1][20]/P0001 ,
		_w9318_,
		_w9407_
	);
	LUT2 #(
		.INIT('h1)
	) name7262 (
		_w9404_,
		_w9405_,
		_w9408_
	);
	LUT2 #(
		.INIT('h1)
	) name7263 (
		_w9406_,
		_w9407_,
		_w9409_
	);
	LUT2 #(
		.INIT('h8)
	) name7264 (
		_w9408_,
		_w9409_,
		_w9410_
	);
	LUT2 #(
		.INIT('h8)
	) name7265 (
		\u10_mem_reg[0][21]/P0001 ,
		_w9314_,
		_w9411_
	);
	LUT2 #(
		.INIT('h8)
	) name7266 (
		\u10_mem_reg[2][21]/P0001 ,
		_w9312_,
		_w9412_
	);
	LUT2 #(
		.INIT('h8)
	) name7267 (
		\u10_mem_reg[3][21]/P0001 ,
		_w9316_,
		_w9413_
	);
	LUT2 #(
		.INIT('h8)
	) name7268 (
		\u10_mem_reg[1][21]/P0001 ,
		_w9318_,
		_w9414_
	);
	LUT2 #(
		.INIT('h1)
	) name7269 (
		_w9411_,
		_w9412_,
		_w9415_
	);
	LUT2 #(
		.INIT('h1)
	) name7270 (
		_w9413_,
		_w9414_,
		_w9416_
	);
	LUT2 #(
		.INIT('h8)
	) name7271 (
		_w9415_,
		_w9416_,
		_w9417_
	);
	LUT2 #(
		.INIT('h8)
	) name7272 (
		\u10_mem_reg[1][22]/P0001 ,
		_w9318_,
		_w9418_
	);
	LUT2 #(
		.INIT('h8)
	) name7273 (
		\u10_mem_reg[2][22]/P0001 ,
		_w9312_,
		_w9419_
	);
	LUT2 #(
		.INIT('h8)
	) name7274 (
		\u10_mem_reg[3][22]/P0001 ,
		_w9316_,
		_w9420_
	);
	LUT2 #(
		.INIT('h8)
	) name7275 (
		\u10_mem_reg[0][22]/P0001 ,
		_w9314_,
		_w9421_
	);
	LUT2 #(
		.INIT('h1)
	) name7276 (
		_w9418_,
		_w9419_,
		_w9422_
	);
	LUT2 #(
		.INIT('h1)
	) name7277 (
		_w9420_,
		_w9421_,
		_w9423_
	);
	LUT2 #(
		.INIT('h8)
	) name7278 (
		_w9422_,
		_w9423_,
		_w9424_
	);
	LUT2 #(
		.INIT('h8)
	) name7279 (
		\u10_mem_reg[0][23]/P0001 ,
		_w9314_,
		_w9425_
	);
	LUT2 #(
		.INIT('h8)
	) name7280 (
		\u10_mem_reg[2][23]/P0001 ,
		_w9312_,
		_w9426_
	);
	LUT2 #(
		.INIT('h8)
	) name7281 (
		\u10_mem_reg[3][23]/P0001 ,
		_w9316_,
		_w9427_
	);
	LUT2 #(
		.INIT('h8)
	) name7282 (
		\u10_mem_reg[1][23]/P0001 ,
		_w9318_,
		_w9428_
	);
	LUT2 #(
		.INIT('h1)
	) name7283 (
		_w9425_,
		_w9426_,
		_w9429_
	);
	LUT2 #(
		.INIT('h1)
	) name7284 (
		_w9427_,
		_w9428_,
		_w9430_
	);
	LUT2 #(
		.INIT('h8)
	) name7285 (
		_w9429_,
		_w9430_,
		_w9431_
	);
	LUT2 #(
		.INIT('h8)
	) name7286 (
		\u10_mem_reg[2][24]/P0001 ,
		_w9312_,
		_w9432_
	);
	LUT2 #(
		.INIT('h8)
	) name7287 (
		\u10_mem_reg[1][24]/P0001 ,
		_w9318_,
		_w9433_
	);
	LUT2 #(
		.INIT('h8)
	) name7288 (
		\u10_mem_reg[3][24]/P0001 ,
		_w9316_,
		_w9434_
	);
	LUT2 #(
		.INIT('h8)
	) name7289 (
		\u10_mem_reg[0][24]/P0001 ,
		_w9314_,
		_w9435_
	);
	LUT2 #(
		.INIT('h1)
	) name7290 (
		_w9432_,
		_w9433_,
		_w9436_
	);
	LUT2 #(
		.INIT('h1)
	) name7291 (
		_w9434_,
		_w9435_,
		_w9437_
	);
	LUT2 #(
		.INIT('h8)
	) name7292 (
		_w9436_,
		_w9437_,
		_w9438_
	);
	LUT2 #(
		.INIT('h8)
	) name7293 (
		\u10_mem_reg[1][25]/P0001 ,
		_w9318_,
		_w9439_
	);
	LUT2 #(
		.INIT('h8)
	) name7294 (
		\u10_mem_reg[2][25]/P0001 ,
		_w9312_,
		_w9440_
	);
	LUT2 #(
		.INIT('h8)
	) name7295 (
		\u10_mem_reg[3][25]/P0001 ,
		_w9316_,
		_w9441_
	);
	LUT2 #(
		.INIT('h8)
	) name7296 (
		\u10_mem_reg[0][25]/P0001 ,
		_w9314_,
		_w9442_
	);
	LUT2 #(
		.INIT('h1)
	) name7297 (
		_w9439_,
		_w9440_,
		_w9443_
	);
	LUT2 #(
		.INIT('h1)
	) name7298 (
		_w9441_,
		_w9442_,
		_w9444_
	);
	LUT2 #(
		.INIT('h8)
	) name7299 (
		_w9443_,
		_w9444_,
		_w9445_
	);
	LUT2 #(
		.INIT('h8)
	) name7300 (
		\u10_mem_reg[2][26]/P0001 ,
		_w9312_,
		_w9446_
	);
	LUT2 #(
		.INIT('h8)
	) name7301 (
		\u10_mem_reg[1][26]/P0001 ,
		_w9318_,
		_w9447_
	);
	LUT2 #(
		.INIT('h8)
	) name7302 (
		\u10_mem_reg[3][26]/P0001 ,
		_w9316_,
		_w9448_
	);
	LUT2 #(
		.INIT('h8)
	) name7303 (
		\u10_mem_reg[0][26]/P0001 ,
		_w9314_,
		_w9449_
	);
	LUT2 #(
		.INIT('h1)
	) name7304 (
		_w9446_,
		_w9447_,
		_w9450_
	);
	LUT2 #(
		.INIT('h1)
	) name7305 (
		_w9448_,
		_w9449_,
		_w9451_
	);
	LUT2 #(
		.INIT('h8)
	) name7306 (
		_w9450_,
		_w9451_,
		_w9452_
	);
	LUT2 #(
		.INIT('h8)
	) name7307 (
		\u10_mem_reg[0][27]/P0001 ,
		_w9314_,
		_w9453_
	);
	LUT2 #(
		.INIT('h8)
	) name7308 (
		\u10_mem_reg[2][27]/P0001 ,
		_w9312_,
		_w9454_
	);
	LUT2 #(
		.INIT('h8)
	) name7309 (
		\u10_mem_reg[3][27]/P0001 ,
		_w9316_,
		_w9455_
	);
	LUT2 #(
		.INIT('h8)
	) name7310 (
		\u10_mem_reg[1][27]/P0001 ,
		_w9318_,
		_w9456_
	);
	LUT2 #(
		.INIT('h1)
	) name7311 (
		_w9453_,
		_w9454_,
		_w9457_
	);
	LUT2 #(
		.INIT('h1)
	) name7312 (
		_w9455_,
		_w9456_,
		_w9458_
	);
	LUT2 #(
		.INIT('h8)
	) name7313 (
		_w9457_,
		_w9458_,
		_w9459_
	);
	LUT2 #(
		.INIT('h8)
	) name7314 (
		\u9_mem_reg[1][4]/P0001 ,
		_w9112_,
		_w9460_
	);
	LUT2 #(
		.INIT('h8)
	) name7315 (
		\u9_mem_reg[0][4]/P0001 ,
		_w9114_,
		_w9461_
	);
	LUT2 #(
		.INIT('h8)
	) name7316 (
		\u9_mem_reg[3][4]/P0001 ,
		_w9116_,
		_w9462_
	);
	LUT2 #(
		.INIT('h8)
	) name7317 (
		\u9_mem_reg[2][4]/P0001 ,
		_w9118_,
		_w9463_
	);
	LUT2 #(
		.INIT('h1)
	) name7318 (
		_w9460_,
		_w9461_,
		_w9464_
	);
	LUT2 #(
		.INIT('h1)
	) name7319 (
		_w9462_,
		_w9463_,
		_w9465_
	);
	LUT2 #(
		.INIT('h8)
	) name7320 (
		_w9464_,
		_w9465_,
		_w9466_
	);
	LUT2 #(
		.INIT('h8)
	) name7321 (
		\u10_mem_reg[0][28]/P0001 ,
		_w9314_,
		_w9467_
	);
	LUT2 #(
		.INIT('h8)
	) name7322 (
		\u10_mem_reg[2][28]/P0001 ,
		_w9312_,
		_w9468_
	);
	LUT2 #(
		.INIT('h8)
	) name7323 (
		\u10_mem_reg[3][28]/P0001 ,
		_w9316_,
		_w9469_
	);
	LUT2 #(
		.INIT('h8)
	) name7324 (
		\u10_mem_reg[1][28]/P0001 ,
		_w9318_,
		_w9470_
	);
	LUT2 #(
		.INIT('h1)
	) name7325 (
		_w9467_,
		_w9468_,
		_w9471_
	);
	LUT2 #(
		.INIT('h1)
	) name7326 (
		_w9469_,
		_w9470_,
		_w9472_
	);
	LUT2 #(
		.INIT('h8)
	) name7327 (
		_w9471_,
		_w9472_,
		_w9473_
	);
	LUT2 #(
		.INIT('h8)
	) name7328 (
		\u10_mem_reg[2][29]/P0001 ,
		_w9312_,
		_w9474_
	);
	LUT2 #(
		.INIT('h8)
	) name7329 (
		\u10_mem_reg[1][29]/P0001 ,
		_w9318_,
		_w9475_
	);
	LUT2 #(
		.INIT('h8)
	) name7330 (
		\u10_mem_reg[3][29]/P0001 ,
		_w9316_,
		_w9476_
	);
	LUT2 #(
		.INIT('h8)
	) name7331 (
		\u10_mem_reg[0][29]/P0001 ,
		_w9314_,
		_w9477_
	);
	LUT2 #(
		.INIT('h1)
	) name7332 (
		_w9474_,
		_w9475_,
		_w9478_
	);
	LUT2 #(
		.INIT('h1)
	) name7333 (
		_w9476_,
		_w9477_,
		_w9479_
	);
	LUT2 #(
		.INIT('h8)
	) name7334 (
		_w9478_,
		_w9479_,
		_w9480_
	);
	LUT2 #(
		.INIT('h8)
	) name7335 (
		\u11_mem_reg[1][0]/P0001 ,
		_w9393_,
		_w9481_
	);
	LUT2 #(
		.INIT('h8)
	) name7336 (
		\u11_mem_reg[0][0]/P0001 ,
		_w9395_,
		_w9482_
	);
	LUT2 #(
		.INIT('h8)
	) name7337 (
		\u11_mem_reg[3][0]/P0001 ,
		_w9397_,
		_w9483_
	);
	LUT2 #(
		.INIT('h8)
	) name7338 (
		\u11_mem_reg[2][0]/P0001 ,
		_w9399_,
		_w9484_
	);
	LUT2 #(
		.INIT('h1)
	) name7339 (
		_w9481_,
		_w9482_,
		_w9485_
	);
	LUT2 #(
		.INIT('h1)
	) name7340 (
		_w9483_,
		_w9484_,
		_w9486_
	);
	LUT2 #(
		.INIT('h8)
	) name7341 (
		_w9485_,
		_w9486_,
		_w9487_
	);
	LUT2 #(
		.INIT('h8)
	) name7342 (
		\u11_mem_reg[1][10]/P0001 ,
		_w9393_,
		_w9488_
	);
	LUT2 #(
		.INIT('h8)
	) name7343 (
		\u11_mem_reg[0][10]/P0001 ,
		_w9395_,
		_w9489_
	);
	LUT2 #(
		.INIT('h8)
	) name7344 (
		\u11_mem_reg[3][10]/P0001 ,
		_w9397_,
		_w9490_
	);
	LUT2 #(
		.INIT('h8)
	) name7345 (
		\u11_mem_reg[2][10]/P0001 ,
		_w9399_,
		_w9491_
	);
	LUT2 #(
		.INIT('h1)
	) name7346 (
		_w9488_,
		_w9489_,
		_w9492_
	);
	LUT2 #(
		.INIT('h1)
	) name7347 (
		_w9490_,
		_w9491_,
		_w9493_
	);
	LUT2 #(
		.INIT('h8)
	) name7348 (
		_w9492_,
		_w9493_,
		_w9494_
	);
	LUT2 #(
		.INIT('h8)
	) name7349 (
		\u10_mem_reg[0][30]/P0001 ,
		_w9314_,
		_w9495_
	);
	LUT2 #(
		.INIT('h8)
	) name7350 (
		\u10_mem_reg[2][30]/P0001 ,
		_w9312_,
		_w9496_
	);
	LUT2 #(
		.INIT('h8)
	) name7351 (
		\u10_mem_reg[3][30]/P0001 ,
		_w9316_,
		_w9497_
	);
	LUT2 #(
		.INIT('h8)
	) name7352 (
		\u10_mem_reg[1][30]/P0001 ,
		_w9318_,
		_w9498_
	);
	LUT2 #(
		.INIT('h1)
	) name7353 (
		_w9495_,
		_w9496_,
		_w9499_
	);
	LUT2 #(
		.INIT('h1)
	) name7354 (
		_w9497_,
		_w9498_,
		_w9500_
	);
	LUT2 #(
		.INIT('h8)
	) name7355 (
		_w9499_,
		_w9500_,
		_w9501_
	);
	LUT2 #(
		.INIT('h8)
	) name7356 (
		\u11_mem_reg[1][11]/P0001 ,
		_w9393_,
		_w9502_
	);
	LUT2 #(
		.INIT('h8)
	) name7357 (
		\u11_mem_reg[0][11]/P0001 ,
		_w9395_,
		_w9503_
	);
	LUT2 #(
		.INIT('h8)
	) name7358 (
		\u11_mem_reg[3][11]/P0001 ,
		_w9397_,
		_w9504_
	);
	LUT2 #(
		.INIT('h8)
	) name7359 (
		\u11_mem_reg[2][11]/P0001 ,
		_w9399_,
		_w9505_
	);
	LUT2 #(
		.INIT('h1)
	) name7360 (
		_w9502_,
		_w9503_,
		_w9506_
	);
	LUT2 #(
		.INIT('h1)
	) name7361 (
		_w9504_,
		_w9505_,
		_w9507_
	);
	LUT2 #(
		.INIT('h8)
	) name7362 (
		_w9506_,
		_w9507_,
		_w9508_
	);
	LUT2 #(
		.INIT('h8)
	) name7363 (
		\u11_mem_reg[1][12]/P0001 ,
		_w9393_,
		_w9509_
	);
	LUT2 #(
		.INIT('h8)
	) name7364 (
		\u11_mem_reg[0][12]/P0001 ,
		_w9395_,
		_w9510_
	);
	LUT2 #(
		.INIT('h8)
	) name7365 (
		\u11_mem_reg[3][12]/P0001 ,
		_w9397_,
		_w9511_
	);
	LUT2 #(
		.INIT('h8)
	) name7366 (
		\u11_mem_reg[2][12]/P0001 ,
		_w9399_,
		_w9512_
	);
	LUT2 #(
		.INIT('h1)
	) name7367 (
		_w9509_,
		_w9510_,
		_w9513_
	);
	LUT2 #(
		.INIT('h1)
	) name7368 (
		_w9511_,
		_w9512_,
		_w9514_
	);
	LUT2 #(
		.INIT('h8)
	) name7369 (
		_w9513_,
		_w9514_,
		_w9515_
	);
	LUT2 #(
		.INIT('h8)
	) name7370 (
		\u11_mem_reg[1][13]/P0001 ,
		_w9393_,
		_w9516_
	);
	LUT2 #(
		.INIT('h8)
	) name7371 (
		\u11_mem_reg[0][13]/P0001 ,
		_w9395_,
		_w9517_
	);
	LUT2 #(
		.INIT('h8)
	) name7372 (
		\u11_mem_reg[3][13]/P0001 ,
		_w9397_,
		_w9518_
	);
	LUT2 #(
		.INIT('h8)
	) name7373 (
		\u11_mem_reg[2][13]/P0001 ,
		_w9399_,
		_w9519_
	);
	LUT2 #(
		.INIT('h1)
	) name7374 (
		_w9516_,
		_w9517_,
		_w9520_
	);
	LUT2 #(
		.INIT('h1)
	) name7375 (
		_w9518_,
		_w9519_,
		_w9521_
	);
	LUT2 #(
		.INIT('h8)
	) name7376 (
		_w9520_,
		_w9521_,
		_w9522_
	);
	LUT2 #(
		.INIT('h8)
	) name7377 (
		\u11_mem_reg[2][14]/P0001 ,
		_w9399_,
		_w9523_
	);
	LUT2 #(
		.INIT('h8)
	) name7378 (
		\u11_mem_reg[0][14]/P0001 ,
		_w9395_,
		_w9524_
	);
	LUT2 #(
		.INIT('h8)
	) name7379 (
		\u11_mem_reg[3][14]/P0001 ,
		_w9397_,
		_w9525_
	);
	LUT2 #(
		.INIT('h8)
	) name7380 (
		\u11_mem_reg[1][14]/P0001 ,
		_w9393_,
		_w9526_
	);
	LUT2 #(
		.INIT('h1)
	) name7381 (
		_w9523_,
		_w9524_,
		_w9527_
	);
	LUT2 #(
		.INIT('h1)
	) name7382 (
		_w9525_,
		_w9526_,
		_w9528_
	);
	LUT2 #(
		.INIT('h8)
	) name7383 (
		_w9527_,
		_w9528_,
		_w9529_
	);
	LUT2 #(
		.INIT('h8)
	) name7384 (
		\u10_mem_reg[2][3]/P0001 ,
		_w9312_,
		_w9530_
	);
	LUT2 #(
		.INIT('h8)
	) name7385 (
		\u10_mem_reg[1][3]/P0001 ,
		_w9318_,
		_w9531_
	);
	LUT2 #(
		.INIT('h8)
	) name7386 (
		\u10_mem_reg[3][3]/P0001 ,
		_w9316_,
		_w9532_
	);
	LUT2 #(
		.INIT('h8)
	) name7387 (
		\u10_mem_reg[0][3]/P0001 ,
		_w9314_,
		_w9533_
	);
	LUT2 #(
		.INIT('h1)
	) name7388 (
		_w9530_,
		_w9531_,
		_w9534_
	);
	LUT2 #(
		.INIT('h1)
	) name7389 (
		_w9532_,
		_w9533_,
		_w9535_
	);
	LUT2 #(
		.INIT('h8)
	) name7390 (
		_w9534_,
		_w9535_,
		_w9536_
	);
	LUT2 #(
		.INIT('h8)
	) name7391 (
		\u11_mem_reg[1][15]/P0001 ,
		_w9393_,
		_w9537_
	);
	LUT2 #(
		.INIT('h8)
	) name7392 (
		\u11_mem_reg[0][15]/P0001 ,
		_w9395_,
		_w9538_
	);
	LUT2 #(
		.INIT('h8)
	) name7393 (
		\u11_mem_reg[3][15]/P0001 ,
		_w9397_,
		_w9539_
	);
	LUT2 #(
		.INIT('h8)
	) name7394 (
		\u11_mem_reg[2][15]/P0001 ,
		_w9399_,
		_w9540_
	);
	LUT2 #(
		.INIT('h1)
	) name7395 (
		_w9537_,
		_w9538_,
		_w9541_
	);
	LUT2 #(
		.INIT('h1)
	) name7396 (
		_w9539_,
		_w9540_,
		_w9542_
	);
	LUT2 #(
		.INIT('h8)
	) name7397 (
		_w9541_,
		_w9542_,
		_w9543_
	);
	LUT2 #(
		.INIT('h8)
	) name7398 (
		\u11_mem_reg[1][16]/P0001 ,
		_w9393_,
		_w9544_
	);
	LUT2 #(
		.INIT('h8)
	) name7399 (
		\u11_mem_reg[0][16]/P0001 ,
		_w9395_,
		_w9545_
	);
	LUT2 #(
		.INIT('h8)
	) name7400 (
		\u11_mem_reg[3][16]/P0001 ,
		_w9397_,
		_w9546_
	);
	LUT2 #(
		.INIT('h8)
	) name7401 (
		\u11_mem_reg[2][16]/P0001 ,
		_w9399_,
		_w9547_
	);
	LUT2 #(
		.INIT('h1)
	) name7402 (
		_w9544_,
		_w9545_,
		_w9548_
	);
	LUT2 #(
		.INIT('h1)
	) name7403 (
		_w9546_,
		_w9547_,
		_w9549_
	);
	LUT2 #(
		.INIT('h8)
	) name7404 (
		_w9548_,
		_w9549_,
		_w9550_
	);
	LUT2 #(
		.INIT('h8)
	) name7405 (
		\u10_mem_reg[2][4]/P0001 ,
		_w9312_,
		_w9551_
	);
	LUT2 #(
		.INIT('h8)
	) name7406 (
		\u10_mem_reg[1][4]/P0001 ,
		_w9318_,
		_w9552_
	);
	LUT2 #(
		.INIT('h8)
	) name7407 (
		\u10_mem_reg[3][4]/P0001 ,
		_w9316_,
		_w9553_
	);
	LUT2 #(
		.INIT('h8)
	) name7408 (
		\u10_mem_reg[0][4]/P0001 ,
		_w9314_,
		_w9554_
	);
	LUT2 #(
		.INIT('h1)
	) name7409 (
		_w9551_,
		_w9552_,
		_w9555_
	);
	LUT2 #(
		.INIT('h1)
	) name7410 (
		_w9553_,
		_w9554_,
		_w9556_
	);
	LUT2 #(
		.INIT('h8)
	) name7411 (
		_w9555_,
		_w9556_,
		_w9557_
	);
	LUT2 #(
		.INIT('h8)
	) name7412 (
		\u11_mem_reg[1][17]/P0001 ,
		_w9393_,
		_w9558_
	);
	LUT2 #(
		.INIT('h8)
	) name7413 (
		\u11_mem_reg[0][17]/P0001 ,
		_w9395_,
		_w9559_
	);
	LUT2 #(
		.INIT('h8)
	) name7414 (
		\u11_mem_reg[3][17]/P0001 ,
		_w9397_,
		_w9560_
	);
	LUT2 #(
		.INIT('h8)
	) name7415 (
		\u11_mem_reg[2][17]/P0001 ,
		_w9399_,
		_w9561_
	);
	LUT2 #(
		.INIT('h1)
	) name7416 (
		_w9558_,
		_w9559_,
		_w9562_
	);
	LUT2 #(
		.INIT('h1)
	) name7417 (
		_w9560_,
		_w9561_,
		_w9563_
	);
	LUT2 #(
		.INIT('h8)
	) name7418 (
		_w9562_,
		_w9563_,
		_w9564_
	);
	LUT2 #(
		.INIT('h8)
	) name7419 (
		\u11_mem_reg[2][18]/P0001 ,
		_w9399_,
		_w9565_
	);
	LUT2 #(
		.INIT('h8)
	) name7420 (
		\u11_mem_reg[1][18]/P0001 ,
		_w9393_,
		_w9566_
	);
	LUT2 #(
		.INIT('h8)
	) name7421 (
		\u11_mem_reg[3][18]/P0001 ,
		_w9397_,
		_w9567_
	);
	LUT2 #(
		.INIT('h8)
	) name7422 (
		\u11_mem_reg[0][18]/P0001 ,
		_w9395_,
		_w9568_
	);
	LUT2 #(
		.INIT('h1)
	) name7423 (
		_w9565_,
		_w9566_,
		_w9569_
	);
	LUT2 #(
		.INIT('h1)
	) name7424 (
		_w9567_,
		_w9568_,
		_w9570_
	);
	LUT2 #(
		.INIT('h8)
	) name7425 (
		_w9569_,
		_w9570_,
		_w9571_
	);
	LUT2 #(
		.INIT('h8)
	) name7426 (
		\u10_mem_reg[2][5]/P0001 ,
		_w9312_,
		_w9572_
	);
	LUT2 #(
		.INIT('h8)
	) name7427 (
		\u10_mem_reg[0][5]/P0001 ,
		_w9314_,
		_w9573_
	);
	LUT2 #(
		.INIT('h8)
	) name7428 (
		\u10_mem_reg[3][5]/P0001 ,
		_w9316_,
		_w9574_
	);
	LUT2 #(
		.INIT('h8)
	) name7429 (
		\u10_mem_reg[1][5]/P0001 ,
		_w9318_,
		_w9575_
	);
	LUT2 #(
		.INIT('h1)
	) name7430 (
		_w9572_,
		_w9573_,
		_w9576_
	);
	LUT2 #(
		.INIT('h1)
	) name7431 (
		_w9574_,
		_w9575_,
		_w9577_
	);
	LUT2 #(
		.INIT('h8)
	) name7432 (
		_w9576_,
		_w9577_,
		_w9578_
	);
	LUT2 #(
		.INIT('h8)
	) name7433 (
		\u11_mem_reg[2][19]/P0001 ,
		_w9399_,
		_w9579_
	);
	LUT2 #(
		.INIT('h8)
	) name7434 (
		\u11_mem_reg[1][19]/P0001 ,
		_w9393_,
		_w9580_
	);
	LUT2 #(
		.INIT('h8)
	) name7435 (
		\u11_mem_reg[3][19]/P0001 ,
		_w9397_,
		_w9581_
	);
	LUT2 #(
		.INIT('h8)
	) name7436 (
		\u11_mem_reg[0][19]/P0001 ,
		_w9395_,
		_w9582_
	);
	LUT2 #(
		.INIT('h1)
	) name7437 (
		_w9579_,
		_w9580_,
		_w9583_
	);
	LUT2 #(
		.INIT('h1)
	) name7438 (
		_w9581_,
		_w9582_,
		_w9584_
	);
	LUT2 #(
		.INIT('h8)
	) name7439 (
		_w9583_,
		_w9584_,
		_w9585_
	);
	LUT2 #(
		.INIT('h8)
	) name7440 (
		\u11_mem_reg[1][1]/P0001 ,
		_w9393_,
		_w9586_
	);
	LUT2 #(
		.INIT('h8)
	) name7441 (
		\u11_mem_reg[0][1]/P0001 ,
		_w9395_,
		_w9587_
	);
	LUT2 #(
		.INIT('h8)
	) name7442 (
		\u11_mem_reg[3][1]/P0001 ,
		_w9397_,
		_w9588_
	);
	LUT2 #(
		.INIT('h8)
	) name7443 (
		\u11_mem_reg[2][1]/P0001 ,
		_w9399_,
		_w9589_
	);
	LUT2 #(
		.INIT('h1)
	) name7444 (
		_w9586_,
		_w9587_,
		_w9590_
	);
	LUT2 #(
		.INIT('h1)
	) name7445 (
		_w9588_,
		_w9589_,
		_w9591_
	);
	LUT2 #(
		.INIT('h8)
	) name7446 (
		_w9590_,
		_w9591_,
		_w9592_
	);
	LUT2 #(
		.INIT('h8)
	) name7447 (
		\u10_mem_reg[2][6]/P0001 ,
		_w9312_,
		_w9593_
	);
	LUT2 #(
		.INIT('h8)
	) name7448 (
		\u10_mem_reg[1][6]/P0001 ,
		_w9318_,
		_w9594_
	);
	LUT2 #(
		.INIT('h8)
	) name7449 (
		\u10_mem_reg[3][6]/P0001 ,
		_w9316_,
		_w9595_
	);
	LUT2 #(
		.INIT('h8)
	) name7450 (
		\u10_mem_reg[0][6]/P0001 ,
		_w9314_,
		_w9596_
	);
	LUT2 #(
		.INIT('h1)
	) name7451 (
		_w9593_,
		_w9594_,
		_w9597_
	);
	LUT2 #(
		.INIT('h1)
	) name7452 (
		_w9595_,
		_w9596_,
		_w9598_
	);
	LUT2 #(
		.INIT('h8)
	) name7453 (
		_w9597_,
		_w9598_,
		_w9599_
	);
	LUT2 #(
		.INIT('h8)
	) name7454 (
		\u11_mem_reg[2][20]/P0001 ,
		_w9399_,
		_w9600_
	);
	LUT2 #(
		.INIT('h8)
	) name7455 (
		\u11_mem_reg[1][20]/P0001 ,
		_w9393_,
		_w9601_
	);
	LUT2 #(
		.INIT('h8)
	) name7456 (
		\u11_mem_reg[3][20]/P0001 ,
		_w9397_,
		_w9602_
	);
	LUT2 #(
		.INIT('h8)
	) name7457 (
		\u11_mem_reg[0][20]/P0001 ,
		_w9395_,
		_w9603_
	);
	LUT2 #(
		.INIT('h1)
	) name7458 (
		_w9600_,
		_w9601_,
		_w9604_
	);
	LUT2 #(
		.INIT('h1)
	) name7459 (
		_w9602_,
		_w9603_,
		_w9605_
	);
	LUT2 #(
		.INIT('h8)
	) name7460 (
		_w9604_,
		_w9605_,
		_w9606_
	);
	LUT2 #(
		.INIT('h8)
	) name7461 (
		\u11_mem_reg[1][21]/P0001 ,
		_w9393_,
		_w9607_
	);
	LUT2 #(
		.INIT('h8)
	) name7462 (
		\u11_mem_reg[2][21]/P0001 ,
		_w9399_,
		_w9608_
	);
	LUT2 #(
		.INIT('h8)
	) name7463 (
		\u11_mem_reg[3][21]/P0001 ,
		_w9397_,
		_w9609_
	);
	LUT2 #(
		.INIT('h8)
	) name7464 (
		\u11_mem_reg[0][21]/P0001 ,
		_w9395_,
		_w9610_
	);
	LUT2 #(
		.INIT('h1)
	) name7465 (
		_w9607_,
		_w9608_,
		_w9611_
	);
	LUT2 #(
		.INIT('h1)
	) name7466 (
		_w9609_,
		_w9610_,
		_w9612_
	);
	LUT2 #(
		.INIT('h8)
	) name7467 (
		_w9611_,
		_w9612_,
		_w9613_
	);
	LUT2 #(
		.INIT('h8)
	) name7468 (
		\u10_mem_reg[2][7]/P0001 ,
		_w9312_,
		_w9614_
	);
	LUT2 #(
		.INIT('h8)
	) name7469 (
		\u10_mem_reg[1][7]/P0001 ,
		_w9318_,
		_w9615_
	);
	LUT2 #(
		.INIT('h8)
	) name7470 (
		\u10_mem_reg[3][7]/P0001 ,
		_w9316_,
		_w9616_
	);
	LUT2 #(
		.INIT('h8)
	) name7471 (
		\u10_mem_reg[0][7]/P0001 ,
		_w9314_,
		_w9617_
	);
	LUT2 #(
		.INIT('h1)
	) name7472 (
		_w9614_,
		_w9615_,
		_w9618_
	);
	LUT2 #(
		.INIT('h1)
	) name7473 (
		_w9616_,
		_w9617_,
		_w9619_
	);
	LUT2 #(
		.INIT('h8)
	) name7474 (
		_w9618_,
		_w9619_,
		_w9620_
	);
	LUT2 #(
		.INIT('h8)
	) name7475 (
		\u11_mem_reg[2][22]/P0001 ,
		_w9399_,
		_w9621_
	);
	LUT2 #(
		.INIT('h8)
	) name7476 (
		\u11_mem_reg[1][22]/P0001 ,
		_w9393_,
		_w9622_
	);
	LUT2 #(
		.INIT('h8)
	) name7477 (
		\u11_mem_reg[3][22]/P0001 ,
		_w9397_,
		_w9623_
	);
	LUT2 #(
		.INIT('h8)
	) name7478 (
		\u11_mem_reg[0][22]/P0001 ,
		_w9395_,
		_w9624_
	);
	LUT2 #(
		.INIT('h1)
	) name7479 (
		_w9621_,
		_w9622_,
		_w9625_
	);
	LUT2 #(
		.INIT('h1)
	) name7480 (
		_w9623_,
		_w9624_,
		_w9626_
	);
	LUT2 #(
		.INIT('h8)
	) name7481 (
		_w9625_,
		_w9626_,
		_w9627_
	);
	LUT2 #(
		.INIT('h8)
	) name7482 (
		\u11_mem_reg[2][23]/P0001 ,
		_w9399_,
		_w9628_
	);
	LUT2 #(
		.INIT('h8)
	) name7483 (
		\u11_mem_reg[1][23]/P0001 ,
		_w9393_,
		_w9629_
	);
	LUT2 #(
		.INIT('h8)
	) name7484 (
		\u11_mem_reg[3][23]/P0001 ,
		_w9397_,
		_w9630_
	);
	LUT2 #(
		.INIT('h8)
	) name7485 (
		\u11_mem_reg[0][23]/P0001 ,
		_w9395_,
		_w9631_
	);
	LUT2 #(
		.INIT('h1)
	) name7486 (
		_w9628_,
		_w9629_,
		_w9632_
	);
	LUT2 #(
		.INIT('h1)
	) name7487 (
		_w9630_,
		_w9631_,
		_w9633_
	);
	LUT2 #(
		.INIT('h8)
	) name7488 (
		_w9632_,
		_w9633_,
		_w9634_
	);
	LUT2 #(
		.INIT('h8)
	) name7489 (
		\u10_mem_reg[2][8]/P0001 ,
		_w9312_,
		_w9635_
	);
	LUT2 #(
		.INIT('h8)
	) name7490 (
		\u10_mem_reg[0][8]/P0001 ,
		_w9314_,
		_w9636_
	);
	LUT2 #(
		.INIT('h8)
	) name7491 (
		\u10_mem_reg[3][8]/P0001 ,
		_w9316_,
		_w9637_
	);
	LUT2 #(
		.INIT('h8)
	) name7492 (
		\u10_mem_reg[1][8]/P0001 ,
		_w9318_,
		_w9638_
	);
	LUT2 #(
		.INIT('h1)
	) name7493 (
		_w9635_,
		_w9636_,
		_w9639_
	);
	LUT2 #(
		.INIT('h1)
	) name7494 (
		_w9637_,
		_w9638_,
		_w9640_
	);
	LUT2 #(
		.INIT('h8)
	) name7495 (
		_w9639_,
		_w9640_,
		_w9641_
	);
	LUT2 #(
		.INIT('h8)
	) name7496 (
		\u11_mem_reg[2][24]/P0001 ,
		_w9399_,
		_w9642_
	);
	LUT2 #(
		.INIT('h8)
	) name7497 (
		\u11_mem_reg[1][24]/P0001 ,
		_w9393_,
		_w9643_
	);
	LUT2 #(
		.INIT('h8)
	) name7498 (
		\u11_mem_reg[3][24]/P0001 ,
		_w9397_,
		_w9644_
	);
	LUT2 #(
		.INIT('h8)
	) name7499 (
		\u11_mem_reg[0][24]/P0001 ,
		_w9395_,
		_w9645_
	);
	LUT2 #(
		.INIT('h1)
	) name7500 (
		_w9642_,
		_w9643_,
		_w9646_
	);
	LUT2 #(
		.INIT('h1)
	) name7501 (
		_w9644_,
		_w9645_,
		_w9647_
	);
	LUT2 #(
		.INIT('h8)
	) name7502 (
		_w9646_,
		_w9647_,
		_w9648_
	);
	LUT2 #(
		.INIT('h8)
	) name7503 (
		\u11_mem_reg[2][25]/P0001 ,
		_w9399_,
		_w9649_
	);
	LUT2 #(
		.INIT('h8)
	) name7504 (
		\u11_mem_reg[1][25]/P0001 ,
		_w9393_,
		_w9650_
	);
	LUT2 #(
		.INIT('h8)
	) name7505 (
		\u11_mem_reg[3][25]/P0001 ,
		_w9397_,
		_w9651_
	);
	LUT2 #(
		.INIT('h8)
	) name7506 (
		\u11_mem_reg[0][25]/P0001 ,
		_w9395_,
		_w9652_
	);
	LUT2 #(
		.INIT('h1)
	) name7507 (
		_w9649_,
		_w9650_,
		_w9653_
	);
	LUT2 #(
		.INIT('h1)
	) name7508 (
		_w9651_,
		_w9652_,
		_w9654_
	);
	LUT2 #(
		.INIT('h8)
	) name7509 (
		_w9653_,
		_w9654_,
		_w9655_
	);
	LUT2 #(
		.INIT('h8)
	) name7510 (
		\u10_mem_reg[1][9]/P0001 ,
		_w9318_,
		_w9656_
	);
	LUT2 #(
		.INIT('h8)
	) name7511 (
		\u10_mem_reg[0][9]/P0001 ,
		_w9314_,
		_w9657_
	);
	LUT2 #(
		.INIT('h8)
	) name7512 (
		\u10_mem_reg[3][9]/P0001 ,
		_w9316_,
		_w9658_
	);
	LUT2 #(
		.INIT('h8)
	) name7513 (
		\u10_mem_reg[2][9]/P0001 ,
		_w9312_,
		_w9659_
	);
	LUT2 #(
		.INIT('h1)
	) name7514 (
		_w9656_,
		_w9657_,
		_w9660_
	);
	LUT2 #(
		.INIT('h1)
	) name7515 (
		_w9658_,
		_w9659_,
		_w9661_
	);
	LUT2 #(
		.INIT('h8)
	) name7516 (
		_w9660_,
		_w9661_,
		_w9662_
	);
	LUT2 #(
		.INIT('h8)
	) name7517 (
		\u11_mem_reg[2][26]/P0001 ,
		_w9399_,
		_w9663_
	);
	LUT2 #(
		.INIT('h8)
	) name7518 (
		\u11_mem_reg[1][26]/P0001 ,
		_w9393_,
		_w9664_
	);
	LUT2 #(
		.INIT('h8)
	) name7519 (
		\u11_mem_reg[3][26]/P0001 ,
		_w9397_,
		_w9665_
	);
	LUT2 #(
		.INIT('h8)
	) name7520 (
		\u11_mem_reg[0][26]/P0001 ,
		_w9395_,
		_w9666_
	);
	LUT2 #(
		.INIT('h1)
	) name7521 (
		_w9663_,
		_w9664_,
		_w9667_
	);
	LUT2 #(
		.INIT('h1)
	) name7522 (
		_w9665_,
		_w9666_,
		_w9668_
	);
	LUT2 #(
		.INIT('h8)
	) name7523 (
		_w9667_,
		_w9668_,
		_w9669_
	);
	LUT2 #(
		.INIT('h8)
	) name7524 (
		\u11_mem_reg[2][27]/P0001 ,
		_w9399_,
		_w9670_
	);
	LUT2 #(
		.INIT('h8)
	) name7525 (
		\u11_mem_reg[1][27]/P0001 ,
		_w9393_,
		_w9671_
	);
	LUT2 #(
		.INIT('h8)
	) name7526 (
		\u11_mem_reg[3][27]/P0001 ,
		_w9397_,
		_w9672_
	);
	LUT2 #(
		.INIT('h8)
	) name7527 (
		\u11_mem_reg[0][27]/P0001 ,
		_w9395_,
		_w9673_
	);
	LUT2 #(
		.INIT('h1)
	) name7528 (
		_w9670_,
		_w9671_,
		_w9674_
	);
	LUT2 #(
		.INIT('h1)
	) name7529 (
		_w9672_,
		_w9673_,
		_w9675_
	);
	LUT2 #(
		.INIT('h8)
	) name7530 (
		_w9674_,
		_w9675_,
		_w9676_
	);
	LUT2 #(
		.INIT('h8)
	) name7531 (
		\u11_mem_reg[2][28]/P0001 ,
		_w9399_,
		_w9677_
	);
	LUT2 #(
		.INIT('h8)
	) name7532 (
		\u11_mem_reg[1][28]/P0001 ,
		_w9393_,
		_w9678_
	);
	LUT2 #(
		.INIT('h8)
	) name7533 (
		\u11_mem_reg[3][28]/P0001 ,
		_w9397_,
		_w9679_
	);
	LUT2 #(
		.INIT('h8)
	) name7534 (
		\u11_mem_reg[0][28]/P0001 ,
		_w9395_,
		_w9680_
	);
	LUT2 #(
		.INIT('h1)
	) name7535 (
		_w9677_,
		_w9678_,
		_w9681_
	);
	LUT2 #(
		.INIT('h1)
	) name7536 (
		_w9679_,
		_w9680_,
		_w9682_
	);
	LUT2 #(
		.INIT('h8)
	) name7537 (
		_w9681_,
		_w9682_,
		_w9683_
	);
	LUT2 #(
		.INIT('h8)
	) name7538 (
		\u10_mem_reg[3][14]/P0001 ,
		_w9316_,
		_w9684_
	);
	LUT2 #(
		.INIT('h8)
	) name7539 (
		\u10_mem_reg[2][14]/P0001 ,
		_w9312_,
		_w9685_
	);
	LUT2 #(
		.INIT('h8)
	) name7540 (
		\u10_mem_reg[0][14]/P0001 ,
		_w9314_,
		_w9686_
	);
	LUT2 #(
		.INIT('h8)
	) name7541 (
		\u10_mem_reg[1][14]/P0001 ,
		_w9318_,
		_w9687_
	);
	LUT2 #(
		.INIT('h1)
	) name7542 (
		_w9684_,
		_w9685_,
		_w9688_
	);
	LUT2 #(
		.INIT('h1)
	) name7543 (
		_w9686_,
		_w9687_,
		_w9689_
	);
	LUT2 #(
		.INIT('h8)
	) name7544 (
		_w9688_,
		_w9689_,
		_w9690_
	);
	LUT2 #(
		.INIT('h8)
	) name7545 (
		\u11_mem_reg[2][29]/P0001 ,
		_w9399_,
		_w9691_
	);
	LUT2 #(
		.INIT('h8)
	) name7546 (
		\u11_mem_reg[1][29]/P0001 ,
		_w9393_,
		_w9692_
	);
	LUT2 #(
		.INIT('h8)
	) name7547 (
		\u11_mem_reg[3][29]/P0001 ,
		_w9397_,
		_w9693_
	);
	LUT2 #(
		.INIT('h8)
	) name7548 (
		\u11_mem_reg[0][29]/P0001 ,
		_w9395_,
		_w9694_
	);
	LUT2 #(
		.INIT('h1)
	) name7549 (
		_w9691_,
		_w9692_,
		_w9695_
	);
	LUT2 #(
		.INIT('h1)
	) name7550 (
		_w9693_,
		_w9694_,
		_w9696_
	);
	LUT2 #(
		.INIT('h8)
	) name7551 (
		_w9695_,
		_w9696_,
		_w9697_
	);
	LUT2 #(
		.INIT('h8)
	) name7552 (
		\u11_mem_reg[1][2]/P0001 ,
		_w9393_,
		_w9698_
	);
	LUT2 #(
		.INIT('h8)
	) name7553 (
		\u11_mem_reg[0][2]/P0001 ,
		_w9395_,
		_w9699_
	);
	LUT2 #(
		.INIT('h8)
	) name7554 (
		\u11_mem_reg[3][2]/P0001 ,
		_w9397_,
		_w9700_
	);
	LUT2 #(
		.INIT('h8)
	) name7555 (
		\u11_mem_reg[2][2]/P0001 ,
		_w9399_,
		_w9701_
	);
	LUT2 #(
		.INIT('h1)
	) name7556 (
		_w9698_,
		_w9699_,
		_w9702_
	);
	LUT2 #(
		.INIT('h1)
	) name7557 (
		_w9700_,
		_w9701_,
		_w9703_
	);
	LUT2 #(
		.INIT('h8)
	) name7558 (
		_w9702_,
		_w9703_,
		_w9704_
	);
	LUT2 #(
		.INIT('h8)
	) name7559 (
		\u11_mem_reg[2][30]/P0001 ,
		_w9399_,
		_w9705_
	);
	LUT2 #(
		.INIT('h8)
	) name7560 (
		\u11_mem_reg[1][30]/P0001 ,
		_w9393_,
		_w9706_
	);
	LUT2 #(
		.INIT('h8)
	) name7561 (
		\u11_mem_reg[3][30]/P0001 ,
		_w9397_,
		_w9707_
	);
	LUT2 #(
		.INIT('h8)
	) name7562 (
		\u11_mem_reg[0][30]/P0001 ,
		_w9395_,
		_w9708_
	);
	LUT2 #(
		.INIT('h1)
	) name7563 (
		_w9705_,
		_w9706_,
		_w9709_
	);
	LUT2 #(
		.INIT('h1)
	) name7564 (
		_w9707_,
		_w9708_,
		_w9710_
	);
	LUT2 #(
		.INIT('h8)
	) name7565 (
		_w9709_,
		_w9710_,
		_w9711_
	);
	LUT2 #(
		.INIT('h8)
	) name7566 (
		\u11_mem_reg[2][31]/P0001 ,
		_w9399_,
		_w9712_
	);
	LUT2 #(
		.INIT('h8)
	) name7567 (
		\u11_mem_reg[1][31]/P0001 ,
		_w9393_,
		_w9713_
	);
	LUT2 #(
		.INIT('h8)
	) name7568 (
		\u11_mem_reg[3][31]/P0001 ,
		_w9397_,
		_w9714_
	);
	LUT2 #(
		.INIT('h8)
	) name7569 (
		\u11_mem_reg[0][31]/P0001 ,
		_w9395_,
		_w9715_
	);
	LUT2 #(
		.INIT('h1)
	) name7570 (
		_w9712_,
		_w9713_,
		_w9716_
	);
	LUT2 #(
		.INIT('h1)
	) name7571 (
		_w9714_,
		_w9715_,
		_w9717_
	);
	LUT2 #(
		.INIT('h8)
	) name7572 (
		_w9716_,
		_w9717_,
		_w9718_
	);
	LUT2 #(
		.INIT('h8)
	) name7573 (
		\u11_mem_reg[1][3]/P0001 ,
		_w9393_,
		_w9719_
	);
	LUT2 #(
		.INIT('h8)
	) name7574 (
		\u11_mem_reg[0][3]/P0001 ,
		_w9395_,
		_w9720_
	);
	LUT2 #(
		.INIT('h8)
	) name7575 (
		\u11_mem_reg[3][3]/P0001 ,
		_w9397_,
		_w9721_
	);
	LUT2 #(
		.INIT('h8)
	) name7576 (
		\u11_mem_reg[2][3]/P0001 ,
		_w9399_,
		_w9722_
	);
	LUT2 #(
		.INIT('h1)
	) name7577 (
		_w9719_,
		_w9720_,
		_w9723_
	);
	LUT2 #(
		.INIT('h1)
	) name7578 (
		_w9721_,
		_w9722_,
		_w9724_
	);
	LUT2 #(
		.INIT('h8)
	) name7579 (
		_w9723_,
		_w9724_,
		_w9725_
	);
	LUT2 #(
		.INIT('h8)
	) name7580 (
		\u11_mem_reg[1][4]/P0001 ,
		_w9393_,
		_w9726_
	);
	LUT2 #(
		.INIT('h8)
	) name7581 (
		\u11_mem_reg[0][4]/P0001 ,
		_w9395_,
		_w9727_
	);
	LUT2 #(
		.INIT('h8)
	) name7582 (
		\u11_mem_reg[3][4]/P0001 ,
		_w9397_,
		_w9728_
	);
	LUT2 #(
		.INIT('h8)
	) name7583 (
		\u11_mem_reg[2][4]/P0001 ,
		_w9399_,
		_w9729_
	);
	LUT2 #(
		.INIT('h1)
	) name7584 (
		_w9726_,
		_w9727_,
		_w9730_
	);
	LUT2 #(
		.INIT('h1)
	) name7585 (
		_w9728_,
		_w9729_,
		_w9731_
	);
	LUT2 #(
		.INIT('h8)
	) name7586 (
		_w9730_,
		_w9731_,
		_w9732_
	);
	LUT2 #(
		.INIT('h8)
	) name7587 (
		\u11_mem_reg[1][5]/P0001 ,
		_w9393_,
		_w9733_
	);
	LUT2 #(
		.INIT('h8)
	) name7588 (
		\u11_mem_reg[0][5]/P0001 ,
		_w9395_,
		_w9734_
	);
	LUT2 #(
		.INIT('h8)
	) name7589 (
		\u11_mem_reg[3][5]/P0001 ,
		_w9397_,
		_w9735_
	);
	LUT2 #(
		.INIT('h8)
	) name7590 (
		\u11_mem_reg[2][5]/P0001 ,
		_w9399_,
		_w9736_
	);
	LUT2 #(
		.INIT('h1)
	) name7591 (
		_w9733_,
		_w9734_,
		_w9737_
	);
	LUT2 #(
		.INIT('h1)
	) name7592 (
		_w9735_,
		_w9736_,
		_w9738_
	);
	LUT2 #(
		.INIT('h8)
	) name7593 (
		_w9737_,
		_w9738_,
		_w9739_
	);
	LUT2 #(
		.INIT('h8)
	) name7594 (
		\u11_mem_reg[2][7]/P0001 ,
		_w9399_,
		_w9740_
	);
	LUT2 #(
		.INIT('h8)
	) name7595 (
		\u11_mem_reg[0][7]/P0001 ,
		_w9395_,
		_w9741_
	);
	LUT2 #(
		.INIT('h8)
	) name7596 (
		\u11_mem_reg[3][7]/P0001 ,
		_w9397_,
		_w9742_
	);
	LUT2 #(
		.INIT('h8)
	) name7597 (
		\u11_mem_reg[1][7]/P0001 ,
		_w9393_,
		_w9743_
	);
	LUT2 #(
		.INIT('h1)
	) name7598 (
		_w9740_,
		_w9741_,
		_w9744_
	);
	LUT2 #(
		.INIT('h1)
	) name7599 (
		_w9742_,
		_w9743_,
		_w9745_
	);
	LUT2 #(
		.INIT('h8)
	) name7600 (
		_w9744_,
		_w9745_,
		_w9746_
	);
	LUT2 #(
		.INIT('h8)
	) name7601 (
		\u11_mem_reg[1][8]/P0001 ,
		_w9393_,
		_w9747_
	);
	LUT2 #(
		.INIT('h8)
	) name7602 (
		\u11_mem_reg[0][8]/P0001 ,
		_w9395_,
		_w9748_
	);
	LUT2 #(
		.INIT('h8)
	) name7603 (
		\u11_mem_reg[3][8]/P0001 ,
		_w9397_,
		_w9749_
	);
	LUT2 #(
		.INIT('h8)
	) name7604 (
		\u11_mem_reg[2][8]/P0001 ,
		_w9399_,
		_w9750_
	);
	LUT2 #(
		.INIT('h1)
	) name7605 (
		_w9747_,
		_w9748_,
		_w9751_
	);
	LUT2 #(
		.INIT('h1)
	) name7606 (
		_w9749_,
		_w9750_,
		_w9752_
	);
	LUT2 #(
		.INIT('h8)
	) name7607 (
		_w9751_,
		_w9752_,
		_w9753_
	);
	LUT2 #(
		.INIT('h8)
	) name7608 (
		\u11_mem_reg[1][9]/P0001 ,
		_w9393_,
		_w9754_
	);
	LUT2 #(
		.INIT('h8)
	) name7609 (
		\u11_mem_reg[0][9]/P0001 ,
		_w9395_,
		_w9755_
	);
	LUT2 #(
		.INIT('h8)
	) name7610 (
		\u11_mem_reg[3][9]/P0001 ,
		_w9397_,
		_w9756_
	);
	LUT2 #(
		.INIT('h8)
	) name7611 (
		\u11_mem_reg[2][9]/P0001 ,
		_w9399_,
		_w9757_
	);
	LUT2 #(
		.INIT('h1)
	) name7612 (
		_w9754_,
		_w9755_,
		_w9758_
	);
	LUT2 #(
		.INIT('h1)
	) name7613 (
		_w9756_,
		_w9757_,
		_w9759_
	);
	LUT2 #(
		.INIT('h8)
	) name7614 (
		_w9758_,
		_w9759_,
		_w9760_
	);
	LUT2 #(
		.INIT('h8)
	) name7615 (
		\u10_mem_reg[2][10]/P0001 ,
		_w9312_,
		_w9761_
	);
	LUT2 #(
		.INIT('h8)
	) name7616 (
		\u10_mem_reg[0][10]/P0001 ,
		_w9314_,
		_w9762_
	);
	LUT2 #(
		.INIT('h8)
	) name7617 (
		\u10_mem_reg[3][10]/P0001 ,
		_w9316_,
		_w9763_
	);
	LUT2 #(
		.INIT('h8)
	) name7618 (
		\u10_mem_reg[1][10]/P0001 ,
		_w9318_,
		_w9764_
	);
	LUT2 #(
		.INIT('h1)
	) name7619 (
		_w9761_,
		_w9762_,
		_w9765_
	);
	LUT2 #(
		.INIT('h1)
	) name7620 (
		_w9763_,
		_w9764_,
		_w9766_
	);
	LUT2 #(
		.INIT('h8)
	) name7621 (
		_w9765_,
		_w9766_,
		_w9767_
	);
	LUT2 #(
		.INIT('h8)
	) name7622 (
		\u10_mem_reg[2][2]/P0001 ,
		_w9312_,
		_w9768_
	);
	LUT2 #(
		.INIT('h8)
	) name7623 (
		\u10_mem_reg[1][2]/P0001 ,
		_w9318_,
		_w9769_
	);
	LUT2 #(
		.INIT('h8)
	) name7624 (
		\u10_mem_reg[3][2]/P0001 ,
		_w9316_,
		_w9770_
	);
	LUT2 #(
		.INIT('h8)
	) name7625 (
		\u10_mem_reg[0][2]/P0001 ,
		_w9314_,
		_w9771_
	);
	LUT2 #(
		.INIT('h1)
	) name7626 (
		_w9768_,
		_w9769_,
		_w9772_
	);
	LUT2 #(
		.INIT('h1)
	) name7627 (
		_w9770_,
		_w9771_,
		_w9773_
	);
	LUT2 #(
		.INIT('h8)
	) name7628 (
		_w9772_,
		_w9773_,
		_w9774_
	);
	LUT2 #(
		.INIT('h8)
	) name7629 (
		\u9_mem_reg[1][8]/P0001 ,
		_w9112_,
		_w9775_
	);
	LUT2 #(
		.INIT('h8)
	) name7630 (
		\u9_mem_reg[0][8]/P0001 ,
		_w9114_,
		_w9776_
	);
	LUT2 #(
		.INIT('h8)
	) name7631 (
		\u9_mem_reg[3][8]/P0001 ,
		_w9116_,
		_w9777_
	);
	LUT2 #(
		.INIT('h8)
	) name7632 (
		\u9_mem_reg[2][8]/P0001 ,
		_w9118_,
		_w9778_
	);
	LUT2 #(
		.INIT('h1)
	) name7633 (
		_w9775_,
		_w9776_,
		_w9779_
	);
	LUT2 #(
		.INIT('h1)
	) name7634 (
		_w9777_,
		_w9778_,
		_w9780_
	);
	LUT2 #(
		.INIT('h8)
	) name7635 (
		_w9779_,
		_w9780_,
		_w9781_
	);
	LUT2 #(
		.INIT('h8)
	) name7636 (
		\u10_mem_reg[1][31]/P0001 ,
		_w9318_,
		_w9782_
	);
	LUT2 #(
		.INIT('h8)
	) name7637 (
		\u10_mem_reg[2][31]/P0001 ,
		_w9312_,
		_w9783_
	);
	LUT2 #(
		.INIT('h8)
	) name7638 (
		\u10_mem_reg[3][31]/P0001 ,
		_w9316_,
		_w9784_
	);
	LUT2 #(
		.INIT('h8)
	) name7639 (
		\u10_mem_reg[0][31]/P0001 ,
		_w9314_,
		_w9785_
	);
	LUT2 #(
		.INIT('h1)
	) name7640 (
		_w9782_,
		_w9783_,
		_w9786_
	);
	LUT2 #(
		.INIT('h1)
	) name7641 (
		_w9784_,
		_w9785_,
		_w9787_
	);
	LUT2 #(
		.INIT('h8)
	) name7642 (
		_w9786_,
		_w9787_,
		_w9788_
	);
	LUT2 #(
		.INIT('h8)
	) name7643 (
		\u9_mem_reg[1][9]/P0001 ,
		_w9112_,
		_w9789_
	);
	LUT2 #(
		.INIT('h8)
	) name7644 (
		\u9_mem_reg[0][9]/P0001 ,
		_w9114_,
		_w9790_
	);
	LUT2 #(
		.INIT('h8)
	) name7645 (
		\u9_mem_reg[3][9]/P0001 ,
		_w9116_,
		_w9791_
	);
	LUT2 #(
		.INIT('h8)
	) name7646 (
		\u9_mem_reg[2][9]/P0001 ,
		_w9118_,
		_w9792_
	);
	LUT2 #(
		.INIT('h1)
	) name7647 (
		_w9789_,
		_w9790_,
		_w9793_
	);
	LUT2 #(
		.INIT('h1)
	) name7648 (
		_w9791_,
		_w9792_,
		_w9794_
	);
	LUT2 #(
		.INIT('h8)
	) name7649 (
		_w9793_,
		_w9794_,
		_w9795_
	);
	LUT2 #(
		.INIT('h2)
	) name7650 (
		\u13_icc_r_reg[10]/NET0131 ,
		\u13_icc_r_reg[11]/NET0131 ,
		_w9796_
	);
	LUT2 #(
		.INIT('h8)
	) name7651 (
		\u1_slt4_reg[5]/P0001 ,
		_w9796_,
		_w9797_
	);
	LUT2 #(
		.INIT('h8)
	) name7652 (
		\u1_slt4_reg[3]/P0001 ,
		_w5671_,
		_w9798_
	);
	LUT2 #(
		.INIT('h8)
	) name7653 (
		\u10_din_tmp1_reg[3]/P0001 ,
		_w3501_,
		_w9799_
	);
	LUT2 #(
		.INIT('h1)
	) name7654 (
		_w9797_,
		_w9798_,
		_w9800_
	);
	LUT2 #(
		.INIT('h4)
	) name7655 (
		_w9799_,
		_w9800_,
		_w9801_
	);
	LUT2 #(
		.INIT('h8)
	) name7656 (
		_w2737_,
		_w9018_,
		_w9802_
	);
	LUT2 #(
		.INIT('h8)
	) name7657 (
		\u1_slt3_reg[1]/P0001 ,
		_w5701_,
		_w9803_
	);
	LUT2 #(
		.INIT('h2)
	) name7658 (
		\u13_icc_r_reg[2]/NET0131 ,
		\u13_icc_r_reg[3]/NET0131 ,
		_w9804_
	);
	LUT2 #(
		.INIT('h8)
	) name7659 (
		\u1_slt3_reg[3]/P0001 ,
		_w9804_,
		_w9805_
	);
	LUT2 #(
		.INIT('h8)
	) name7660 (
		\u9_din_tmp1_reg[1]/P0001 ,
		_w3311_,
		_w9806_
	);
	LUT2 #(
		.INIT('h1)
	) name7661 (
		_w9803_,
		_w9805_,
		_w9807_
	);
	LUT2 #(
		.INIT('h4)
	) name7662 (
		_w9806_,
		_w9807_,
		_w9808_
	);
	LUT2 #(
		.INIT('h8)
	) name7663 (
		\u1_slt3_reg[2]/P0001 ,
		_w5701_,
		_w9809_
	);
	LUT2 #(
		.INIT('h8)
	) name7664 (
		\u1_slt3_reg[4]/P0001 ,
		_w9804_,
		_w9810_
	);
	LUT2 #(
		.INIT('h8)
	) name7665 (
		\u9_din_tmp1_reg[2]/P0001 ,
		_w3311_,
		_w9811_
	);
	LUT2 #(
		.INIT('h1)
	) name7666 (
		_w9809_,
		_w9810_,
		_w9812_
	);
	LUT2 #(
		.INIT('h4)
	) name7667 (
		_w9811_,
		_w9812_,
		_w9813_
	);
	LUT2 #(
		.INIT('h8)
	) name7668 (
		\u1_slt3_reg[8]/P0001 ,
		_w5701_,
		_w9814_
	);
	LUT2 #(
		.INIT('h8)
	) name7669 (
		\u1_slt3_reg[10]/P0001 ,
		_w9804_,
		_w9815_
	);
	LUT2 #(
		.INIT('h8)
	) name7670 (
		\u9_din_tmp1_reg[8]/P0001 ,
		_w3311_,
		_w9816_
	);
	LUT2 #(
		.INIT('h1)
	) name7671 (
		_w9814_,
		_w9815_,
		_w9817_
	);
	LUT2 #(
		.INIT('h4)
	) name7672 (
		_w9816_,
		_w9817_,
		_w9818_
	);
	LUT2 #(
		.INIT('h8)
	) name7673 (
		\u1_slt3_reg[17]/P0001 ,
		_w5701_,
		_w9819_
	);
	LUT2 #(
		.INIT('h8)
	) name7674 (
		\u1_slt3_reg[5]/P0001 ,
		_w3311_,
		_w9820_
	);
	LUT2 #(
		.INIT('h8)
	) name7675 (
		\u1_slt3_reg[19]/P0001 ,
		_w9804_,
		_w9821_
	);
	LUT2 #(
		.INIT('h1)
	) name7676 (
		_w9819_,
		_w9820_,
		_w9822_
	);
	LUT2 #(
		.INIT('h4)
	) name7677 (
		_w9821_,
		_w9822_,
		_w9823_
	);
	LUT2 #(
		.INIT('h8)
	) name7678 (
		\u1_slt3_reg[16]/P0001 ,
		_w5701_,
		_w9824_
	);
	LUT2 #(
		.INIT('h8)
	) name7679 (
		\u1_slt3_reg[4]/P0001 ,
		_w3311_,
		_w9825_
	);
	LUT2 #(
		.INIT('h8)
	) name7680 (
		\u1_slt3_reg[18]/P0001 ,
		_w9804_,
		_w9826_
	);
	LUT2 #(
		.INIT('h1)
	) name7681 (
		_w9824_,
		_w9825_,
		_w9827_
	);
	LUT2 #(
		.INIT('h4)
	) name7682 (
		_w9826_,
		_w9827_,
		_w9828_
	);
	LUT2 #(
		.INIT('h8)
	) name7683 (
		\u1_slt3_reg[15]/P0001 ,
		_w5701_,
		_w9829_
	);
	LUT2 #(
		.INIT('h8)
	) name7684 (
		\u1_slt3_reg[17]/P0001 ,
		_w9804_,
		_w9830_
	);
	LUT2 #(
		.INIT('h8)
	) name7685 (
		\u9_din_tmp1_reg[15]/P0001 ,
		_w3311_,
		_w9831_
	);
	LUT2 #(
		.INIT('h1)
	) name7686 (
		_w9829_,
		_w9830_,
		_w9832_
	);
	LUT2 #(
		.INIT('h4)
	) name7687 (
		_w9831_,
		_w9832_,
		_w9833_
	);
	LUT2 #(
		.INIT('h8)
	) name7688 (
		\u1_slt3_reg[14]/P0001 ,
		_w5701_,
		_w9834_
	);
	LUT2 #(
		.INIT('h8)
	) name7689 (
		\u1_slt3_reg[16]/P0001 ,
		_w9804_,
		_w9835_
	);
	LUT2 #(
		.INIT('h8)
	) name7690 (
		\u9_din_tmp1_reg[14]/P0001 ,
		_w3311_,
		_w9836_
	);
	LUT2 #(
		.INIT('h1)
	) name7691 (
		_w9834_,
		_w9835_,
		_w9837_
	);
	LUT2 #(
		.INIT('h4)
	) name7692 (
		_w9836_,
		_w9837_,
		_w9838_
	);
	LUT2 #(
		.INIT('h8)
	) name7693 (
		\u1_slt3_reg[13]/P0001 ,
		_w5701_,
		_w9839_
	);
	LUT2 #(
		.INIT('h8)
	) name7694 (
		\u1_slt3_reg[15]/P0001 ,
		_w9804_,
		_w9840_
	);
	LUT2 #(
		.INIT('h8)
	) name7695 (
		\u9_din_tmp1_reg[13]/P0001 ,
		_w3311_,
		_w9841_
	);
	LUT2 #(
		.INIT('h1)
	) name7696 (
		_w9839_,
		_w9840_,
		_w9842_
	);
	LUT2 #(
		.INIT('h4)
	) name7697 (
		_w9841_,
		_w9842_,
		_w9843_
	);
	LUT2 #(
		.INIT('h8)
	) name7698 (
		\u1_slt3_reg[12]/P0001 ,
		_w5701_,
		_w9844_
	);
	LUT2 #(
		.INIT('h8)
	) name7699 (
		\u1_slt3_reg[14]/P0001 ,
		_w9804_,
		_w9845_
	);
	LUT2 #(
		.INIT('h8)
	) name7700 (
		\u9_din_tmp1_reg[12]/P0001 ,
		_w3311_,
		_w9846_
	);
	LUT2 #(
		.INIT('h1)
	) name7701 (
		_w9844_,
		_w9845_,
		_w9847_
	);
	LUT2 #(
		.INIT('h4)
	) name7702 (
		_w9846_,
		_w9847_,
		_w9848_
	);
	LUT2 #(
		.INIT('h8)
	) name7703 (
		\u1_slt3_reg[13]/P0001 ,
		_w9804_,
		_w9849_
	);
	LUT2 #(
		.INIT('h8)
	) name7704 (
		\u1_slt3_reg[11]/P0001 ,
		_w5701_,
		_w9850_
	);
	LUT2 #(
		.INIT('h8)
	) name7705 (
		\u9_din_tmp1_reg[11]/P0001 ,
		_w3311_,
		_w9851_
	);
	LUT2 #(
		.INIT('h1)
	) name7706 (
		_w9849_,
		_w9850_,
		_w9852_
	);
	LUT2 #(
		.INIT('h4)
	) name7707 (
		_w9851_,
		_w9852_,
		_w9853_
	);
	LUT2 #(
		.INIT('h8)
	) name7708 (
		\u1_slt3_reg[9]/P0001 ,
		_w5701_,
		_w9854_
	);
	LUT2 #(
		.INIT('h8)
	) name7709 (
		\u1_slt3_reg[11]/P0001 ,
		_w9804_,
		_w9855_
	);
	LUT2 #(
		.INIT('h8)
	) name7710 (
		\u9_din_tmp1_reg[9]/P0001 ,
		_w3311_,
		_w9856_
	);
	LUT2 #(
		.INIT('h1)
	) name7711 (
		_w9854_,
		_w9855_,
		_w9857_
	);
	LUT2 #(
		.INIT('h4)
	) name7712 (
		_w9856_,
		_w9857_,
		_w9858_
	);
	LUT2 #(
		.INIT('h8)
	) name7713 (
		\u1_slt3_reg[3]/P0001 ,
		_w5701_,
		_w9859_
	);
	LUT2 #(
		.INIT('h8)
	) name7714 (
		\u1_slt3_reg[5]/P0001 ,
		_w9804_,
		_w9860_
	);
	LUT2 #(
		.INIT('h8)
	) name7715 (
		\u9_din_tmp1_reg[3]/P0001 ,
		_w3311_,
		_w9861_
	);
	LUT2 #(
		.INIT('h1)
	) name7716 (
		_w9859_,
		_w9860_,
		_w9862_
	);
	LUT2 #(
		.INIT('h4)
	) name7717 (
		_w9861_,
		_w9862_,
		_w9863_
	);
	LUT2 #(
		.INIT('h8)
	) name7718 (
		\u1_slt3_reg[12]/P0001 ,
		_w9804_,
		_w9864_
	);
	LUT2 #(
		.INIT('h8)
	) name7719 (
		\u1_slt3_reg[10]/P0001 ,
		_w5701_,
		_w9865_
	);
	LUT2 #(
		.INIT('h8)
	) name7720 (
		\u9_din_tmp1_reg[10]/P0001 ,
		_w3311_,
		_w9866_
	);
	LUT2 #(
		.INIT('h1)
	) name7721 (
		_w9864_,
		_w9865_,
		_w9867_
	);
	LUT2 #(
		.INIT('h4)
	) name7722 (
		_w9866_,
		_w9867_,
		_w9868_
	);
	LUT2 #(
		.INIT('h2)
	) name7723 (
		\u13_icc_r_reg[18]/NET0131 ,
		\u13_icc_r_reg[19]/NET0131 ,
		_w9869_
	);
	LUT2 #(
		.INIT('h8)
	) name7724 (
		\u1_slt6_reg[13]/P0001 ,
		_w9869_,
		_w9870_
	);
	LUT2 #(
		.INIT('h8)
	) name7725 (
		\u1_slt6_reg[11]/P0001 ,
		_w5936_,
		_w9871_
	);
	LUT2 #(
		.INIT('h8)
	) name7726 (
		\u11_din_tmp1_reg[11]/P0001 ,
		_w3064_,
		_w9872_
	);
	LUT2 #(
		.INIT('h1)
	) name7727 (
		_w9870_,
		_w9871_,
		_w9873_
	);
	LUT2 #(
		.INIT('h4)
	) name7728 (
		_w9872_,
		_w9873_,
		_w9874_
	);
	LUT2 #(
		.INIT('h8)
	) name7729 (
		\u1_slt4_reg[9]/P0001 ,
		_w5671_,
		_w9875_
	);
	LUT2 #(
		.INIT('h8)
	) name7730 (
		\u1_slt4_reg[11]/P0001 ,
		_w9796_,
		_w9876_
	);
	LUT2 #(
		.INIT('h8)
	) name7731 (
		\u10_din_tmp1_reg[9]/P0001 ,
		_w3501_,
		_w9877_
	);
	LUT2 #(
		.INIT('h1)
	) name7732 (
		_w9875_,
		_w9876_,
		_w9878_
	);
	LUT2 #(
		.INIT('h4)
	) name7733 (
		_w9877_,
		_w9878_,
		_w9879_
	);
	LUT2 #(
		.INIT('h8)
	) name7734 (
		\u1_slt3_reg[6]/P0001 ,
		_w5701_,
		_w9880_
	);
	LUT2 #(
		.INIT('h8)
	) name7735 (
		\u1_slt3_reg[8]/P0001 ,
		_w9804_,
		_w9881_
	);
	LUT2 #(
		.INIT('h8)
	) name7736 (
		\u9_din_tmp1_reg[6]/P0001 ,
		_w3311_,
		_w9882_
	);
	LUT2 #(
		.INIT('h1)
	) name7737 (
		_w9880_,
		_w9881_,
		_w9883_
	);
	LUT2 #(
		.INIT('h4)
	) name7738 (
		_w9882_,
		_w9883_,
		_w9884_
	);
	LUT2 #(
		.INIT('h8)
	) name7739 (
		\u1_slt4_reg[0]/P0001 ,
		_w5671_,
		_w9885_
	);
	LUT2 #(
		.INIT('h8)
	) name7740 (
		\u1_slt4_reg[2]/P0001 ,
		_w9796_,
		_w9886_
	);
	LUT2 #(
		.INIT('h8)
	) name7741 (
		\u10_din_tmp1_reg[0]/P0001 ,
		_w3501_,
		_w9887_
	);
	LUT2 #(
		.INIT('h1)
	) name7742 (
		_w9885_,
		_w9886_,
		_w9888_
	);
	LUT2 #(
		.INIT('h4)
	) name7743 (
		_w9887_,
		_w9888_,
		_w9889_
	);
	LUT2 #(
		.INIT('h8)
	) name7744 (
		\u1_slt4_reg[12]/P0001 ,
		_w9796_,
		_w9890_
	);
	LUT2 #(
		.INIT('h8)
	) name7745 (
		\u1_slt4_reg[10]/P0001 ,
		_w5671_,
		_w9891_
	);
	LUT2 #(
		.INIT('h8)
	) name7746 (
		\u10_din_tmp1_reg[10]/P0001 ,
		_w3501_,
		_w9892_
	);
	LUT2 #(
		.INIT('h1)
	) name7747 (
		_w9890_,
		_w9891_,
		_w9893_
	);
	LUT2 #(
		.INIT('h4)
	) name7748 (
		_w9892_,
		_w9893_,
		_w9894_
	);
	LUT2 #(
		.INIT('h8)
	) name7749 (
		\u1_slt4_reg[13]/P0001 ,
		_w9796_,
		_w9895_
	);
	LUT2 #(
		.INIT('h8)
	) name7750 (
		\u1_slt4_reg[11]/P0001 ,
		_w5671_,
		_w9896_
	);
	LUT2 #(
		.INIT('h8)
	) name7751 (
		\u10_din_tmp1_reg[11]/P0001 ,
		_w3501_,
		_w9897_
	);
	LUT2 #(
		.INIT('h1)
	) name7752 (
		_w9895_,
		_w9896_,
		_w9898_
	);
	LUT2 #(
		.INIT('h4)
	) name7753 (
		_w9897_,
		_w9898_,
		_w9899_
	);
	LUT2 #(
		.INIT('h8)
	) name7754 (
		\u1_slt4_reg[14]/P0001 ,
		_w9796_,
		_w9900_
	);
	LUT2 #(
		.INIT('h8)
	) name7755 (
		\u1_slt4_reg[12]/P0001 ,
		_w5671_,
		_w9901_
	);
	LUT2 #(
		.INIT('h8)
	) name7756 (
		\u10_din_tmp1_reg[12]/P0001 ,
		_w3501_,
		_w9902_
	);
	LUT2 #(
		.INIT('h1)
	) name7757 (
		_w9900_,
		_w9901_,
		_w9903_
	);
	LUT2 #(
		.INIT('h4)
	) name7758 (
		_w9902_,
		_w9903_,
		_w9904_
	);
	LUT2 #(
		.INIT('h8)
	) name7759 (
		\u1_slt3_reg[7]/P0001 ,
		_w5701_,
		_w9905_
	);
	LUT2 #(
		.INIT('h8)
	) name7760 (
		\u1_slt3_reg[9]/P0001 ,
		_w9804_,
		_w9906_
	);
	LUT2 #(
		.INIT('h8)
	) name7761 (
		\u9_din_tmp1_reg[7]/P0001 ,
		_w3311_,
		_w9907_
	);
	LUT2 #(
		.INIT('h1)
	) name7762 (
		_w9905_,
		_w9906_,
		_w9908_
	);
	LUT2 #(
		.INIT('h4)
	) name7763 (
		_w9907_,
		_w9908_,
		_w9909_
	);
	LUT2 #(
		.INIT('h8)
	) name7764 (
		\u1_slt4_reg[15]/P0001 ,
		_w9796_,
		_w9910_
	);
	LUT2 #(
		.INIT('h8)
	) name7765 (
		\u1_slt4_reg[13]/P0001 ,
		_w5671_,
		_w9911_
	);
	LUT2 #(
		.INIT('h8)
	) name7766 (
		\u10_din_tmp1_reg[13]/P0001 ,
		_w3501_,
		_w9912_
	);
	LUT2 #(
		.INIT('h1)
	) name7767 (
		_w9910_,
		_w9911_,
		_w9913_
	);
	LUT2 #(
		.INIT('h4)
	) name7768 (
		_w9912_,
		_w9913_,
		_w9914_
	);
	LUT2 #(
		.INIT('h8)
	) name7769 (
		\u1_slt3_reg[5]/P0001 ,
		_w5701_,
		_w9915_
	);
	LUT2 #(
		.INIT('h8)
	) name7770 (
		\u1_slt3_reg[7]/P0001 ,
		_w9804_,
		_w9916_
	);
	LUT2 #(
		.INIT('h8)
	) name7771 (
		\u9_din_tmp1_reg[5]/P0001 ,
		_w3311_,
		_w9917_
	);
	LUT2 #(
		.INIT('h1)
	) name7772 (
		_w9915_,
		_w9916_,
		_w9918_
	);
	LUT2 #(
		.INIT('h4)
	) name7773 (
		_w9917_,
		_w9918_,
		_w9919_
	);
	LUT2 #(
		.INIT('h8)
	) name7774 (
		\u1_slt6_reg[0]/P0001 ,
		_w5936_,
		_w9920_
	);
	LUT2 #(
		.INIT('h8)
	) name7775 (
		\u1_slt6_reg[2]/P0001 ,
		_w9869_,
		_w9921_
	);
	LUT2 #(
		.INIT('h8)
	) name7776 (
		\u11_din_tmp1_reg[0]/P0001 ,
		_w3064_,
		_w9922_
	);
	LUT2 #(
		.INIT('h1)
	) name7777 (
		_w9920_,
		_w9921_,
		_w9923_
	);
	LUT2 #(
		.INIT('h4)
	) name7778 (
		_w9922_,
		_w9923_,
		_w9924_
	);
	LUT2 #(
		.INIT('h8)
	) name7779 (
		\u1_slt6_reg[12]/P0001 ,
		_w9869_,
		_w9925_
	);
	LUT2 #(
		.INIT('h8)
	) name7780 (
		\u1_slt6_reg[10]/P0001 ,
		_w5936_,
		_w9926_
	);
	LUT2 #(
		.INIT('h8)
	) name7781 (
		\u11_din_tmp1_reg[10]/P0001 ,
		_w3064_,
		_w9927_
	);
	LUT2 #(
		.INIT('h1)
	) name7782 (
		_w9925_,
		_w9926_,
		_w9928_
	);
	LUT2 #(
		.INIT('h4)
	) name7783 (
		_w9927_,
		_w9928_,
		_w9929_
	);
	LUT2 #(
		.INIT('h8)
	) name7784 (
		\u1_slt4_reg[17]/P0001 ,
		_w9796_,
		_w9930_
	);
	LUT2 #(
		.INIT('h8)
	) name7785 (
		\u1_slt4_reg[15]/P0001 ,
		_w5671_,
		_w9931_
	);
	LUT2 #(
		.INIT('h8)
	) name7786 (
		\u10_din_tmp1_reg[15]/P0001 ,
		_w3501_,
		_w9932_
	);
	LUT2 #(
		.INIT('h1)
	) name7787 (
		_w9930_,
		_w9931_,
		_w9933_
	);
	LUT2 #(
		.INIT('h4)
	) name7788 (
		_w9932_,
		_w9933_,
		_w9934_
	);
	LUT2 #(
		.INIT('h8)
	) name7789 (
		\u1_slt6_reg[14]/P0001 ,
		_w9869_,
		_w9935_
	);
	LUT2 #(
		.INIT('h8)
	) name7790 (
		\u1_slt6_reg[12]/P0001 ,
		_w5936_,
		_w9936_
	);
	LUT2 #(
		.INIT('h8)
	) name7791 (
		\u11_din_tmp1_reg[12]/P0001 ,
		_w3064_,
		_w9937_
	);
	LUT2 #(
		.INIT('h1)
	) name7792 (
		_w9935_,
		_w9936_,
		_w9938_
	);
	LUT2 #(
		.INIT('h4)
	) name7793 (
		_w9937_,
		_w9938_,
		_w9939_
	);
	LUT2 #(
		.INIT('h8)
	) name7794 (
		\u1_slt6_reg[15]/P0001 ,
		_w9869_,
		_w9940_
	);
	LUT2 #(
		.INIT('h8)
	) name7795 (
		\u1_slt6_reg[13]/P0001 ,
		_w5936_,
		_w9941_
	);
	LUT2 #(
		.INIT('h8)
	) name7796 (
		\u11_din_tmp1_reg[13]/P0001 ,
		_w3064_,
		_w9942_
	);
	LUT2 #(
		.INIT('h1)
	) name7797 (
		_w9940_,
		_w9941_,
		_w9943_
	);
	LUT2 #(
		.INIT('h4)
	) name7798 (
		_w9942_,
		_w9943_,
		_w9944_
	);
	LUT2 #(
		.INIT('h8)
	) name7799 (
		\u1_slt4_reg[18]/P0001 ,
		_w9796_,
		_w9945_
	);
	LUT2 #(
		.INIT('h8)
	) name7800 (
		\u1_slt4_reg[4]/P0001 ,
		_w3501_,
		_w9946_
	);
	LUT2 #(
		.INIT('h8)
	) name7801 (
		\u1_slt4_reg[16]/P0001 ,
		_w5671_,
		_w9947_
	);
	LUT2 #(
		.INIT('h1)
	) name7802 (
		_w9945_,
		_w9946_,
		_w9948_
	);
	LUT2 #(
		.INIT('h4)
	) name7803 (
		_w9947_,
		_w9948_,
		_w9949_
	);
	LUT2 #(
		.INIT('h8)
	) name7804 (
		\u1_slt6_reg[16]/P0001 ,
		_w9869_,
		_w9950_
	);
	LUT2 #(
		.INIT('h8)
	) name7805 (
		\u1_slt6_reg[14]/P0001 ,
		_w5936_,
		_w9951_
	);
	LUT2 #(
		.INIT('h8)
	) name7806 (
		\u11_din_tmp1_reg[14]/P0001 ,
		_w3064_,
		_w9952_
	);
	LUT2 #(
		.INIT('h1)
	) name7807 (
		_w9950_,
		_w9951_,
		_w9953_
	);
	LUT2 #(
		.INIT('h4)
	) name7808 (
		_w9952_,
		_w9953_,
		_w9954_
	);
	LUT2 #(
		.INIT('h8)
	) name7809 (
		\u1_slt4_reg[19]/P0001 ,
		_w9796_,
		_w9955_
	);
	LUT2 #(
		.INIT('h8)
	) name7810 (
		\u1_slt4_reg[5]/P0001 ,
		_w3501_,
		_w9956_
	);
	LUT2 #(
		.INIT('h8)
	) name7811 (
		\u1_slt4_reg[17]/P0001 ,
		_w5671_,
		_w9957_
	);
	LUT2 #(
		.INIT('h1)
	) name7812 (
		_w9955_,
		_w9956_,
		_w9958_
	);
	LUT2 #(
		.INIT('h4)
	) name7813 (
		_w9957_,
		_w9958_,
		_w9959_
	);
	LUT2 #(
		.INIT('h8)
	) name7814 (
		\u1_slt6_reg[19]/P0001 ,
		_w9869_,
		_w9960_
	);
	LUT2 #(
		.INIT('h8)
	) name7815 (
		\u1_slt6_reg[5]/P0001 ,
		_w3064_,
		_w9961_
	);
	LUT2 #(
		.INIT('h8)
	) name7816 (
		\u1_slt6_reg[17]/P0001 ,
		_w5936_,
		_w9962_
	);
	LUT2 #(
		.INIT('h1)
	) name7817 (
		_w9960_,
		_w9961_,
		_w9963_
	);
	LUT2 #(
		.INIT('h4)
	) name7818 (
		_w9962_,
		_w9963_,
		_w9964_
	);
	LUT2 #(
		.INIT('h8)
	) name7819 (
		\u1_slt6_reg[1]/P0001 ,
		_w5936_,
		_w9965_
	);
	LUT2 #(
		.INIT('h8)
	) name7820 (
		\u1_slt6_reg[3]/P0001 ,
		_w9869_,
		_w9966_
	);
	LUT2 #(
		.INIT('h8)
	) name7821 (
		\u11_din_tmp1_reg[1]/P0001 ,
		_w3064_,
		_w9967_
	);
	LUT2 #(
		.INIT('h1)
	) name7822 (
		_w9965_,
		_w9966_,
		_w9968_
	);
	LUT2 #(
		.INIT('h4)
	) name7823 (
		_w9967_,
		_w9968_,
		_w9969_
	);
	LUT2 #(
		.INIT('h8)
	) name7824 (
		\u1_slt4_reg[1]/P0001 ,
		_w5671_,
		_w9970_
	);
	LUT2 #(
		.INIT('h8)
	) name7825 (
		\u1_slt4_reg[3]/P0001 ,
		_w9796_,
		_w9971_
	);
	LUT2 #(
		.INIT('h8)
	) name7826 (
		\u10_din_tmp1_reg[1]/P0001 ,
		_w3501_,
		_w9972_
	);
	LUT2 #(
		.INIT('h1)
	) name7827 (
		_w9970_,
		_w9971_,
		_w9973_
	);
	LUT2 #(
		.INIT('h4)
	) name7828 (
		_w9972_,
		_w9973_,
		_w9974_
	);
	LUT2 #(
		.INIT('h8)
	) name7829 (
		\u1_slt4_reg[16]/P0001 ,
		_w9796_,
		_w9975_
	);
	LUT2 #(
		.INIT('h8)
	) name7830 (
		\u1_slt4_reg[14]/P0001 ,
		_w5671_,
		_w9976_
	);
	LUT2 #(
		.INIT('h8)
	) name7831 (
		\u10_din_tmp1_reg[14]/P0001 ,
		_w3501_,
		_w9977_
	);
	LUT2 #(
		.INIT('h1)
	) name7832 (
		_w9975_,
		_w9976_,
		_w9978_
	);
	LUT2 #(
		.INIT('h4)
	) name7833 (
		_w9977_,
		_w9978_,
		_w9979_
	);
	LUT2 #(
		.INIT('h8)
	) name7834 (
		\u1_slt6_reg[4]/P0001 ,
		_w9869_,
		_w9980_
	);
	LUT2 #(
		.INIT('h8)
	) name7835 (
		\u1_slt6_reg[2]/P0001 ,
		_w5936_,
		_w9981_
	);
	LUT2 #(
		.INIT('h8)
	) name7836 (
		\u11_din_tmp1_reg[2]/P0001 ,
		_w3064_,
		_w9982_
	);
	LUT2 #(
		.INIT('h1)
	) name7837 (
		_w9980_,
		_w9981_,
		_w9983_
	);
	LUT2 #(
		.INIT('h4)
	) name7838 (
		_w9982_,
		_w9983_,
		_w9984_
	);
	LUT2 #(
		.INIT('h8)
	) name7839 (
		\u1_slt6_reg[18]/P0001 ,
		_w9869_,
		_w9985_
	);
	LUT2 #(
		.INIT('h8)
	) name7840 (
		\u1_slt6_reg[4]/P0001 ,
		_w3064_,
		_w9986_
	);
	LUT2 #(
		.INIT('h8)
	) name7841 (
		\u1_slt6_reg[16]/P0001 ,
		_w5936_,
		_w9987_
	);
	LUT2 #(
		.INIT('h1)
	) name7842 (
		_w9985_,
		_w9986_,
		_w9988_
	);
	LUT2 #(
		.INIT('h4)
	) name7843 (
		_w9987_,
		_w9988_,
		_w9989_
	);
	LUT2 #(
		.INIT('h8)
	) name7844 (
		\u1_slt6_reg[5]/P0001 ,
		_w9869_,
		_w9990_
	);
	LUT2 #(
		.INIT('h8)
	) name7845 (
		\u1_slt6_reg[3]/P0001 ,
		_w5936_,
		_w9991_
	);
	LUT2 #(
		.INIT('h8)
	) name7846 (
		\u11_din_tmp1_reg[3]/P0001 ,
		_w3064_,
		_w9992_
	);
	LUT2 #(
		.INIT('h1)
	) name7847 (
		_w9990_,
		_w9991_,
		_w9993_
	);
	LUT2 #(
		.INIT('h4)
	) name7848 (
		_w9992_,
		_w9993_,
		_w9994_
	);
	LUT2 #(
		.INIT('h8)
	) name7849 (
		\u1_slt6_reg[6]/P0001 ,
		_w9869_,
		_w9995_
	);
	LUT2 #(
		.INIT('h8)
	) name7850 (
		\u1_slt6_reg[4]/P0001 ,
		_w5936_,
		_w9996_
	);
	LUT2 #(
		.INIT('h8)
	) name7851 (
		\u11_din_tmp1_reg[4]/P0001 ,
		_w3064_,
		_w9997_
	);
	LUT2 #(
		.INIT('h1)
	) name7852 (
		_w9995_,
		_w9996_,
		_w9998_
	);
	LUT2 #(
		.INIT('h4)
	) name7853 (
		_w9997_,
		_w9998_,
		_w9999_
	);
	LUT2 #(
		.INIT('h8)
	) name7854 (
		\u1_slt6_reg[7]/P0001 ,
		_w9869_,
		_w10000_
	);
	LUT2 #(
		.INIT('h8)
	) name7855 (
		\u1_slt6_reg[5]/P0001 ,
		_w5936_,
		_w10001_
	);
	LUT2 #(
		.INIT('h8)
	) name7856 (
		\u11_din_tmp1_reg[5]/P0001 ,
		_w3064_,
		_w10002_
	);
	LUT2 #(
		.INIT('h1)
	) name7857 (
		_w10000_,
		_w10001_,
		_w10003_
	);
	LUT2 #(
		.INIT('h4)
	) name7858 (
		_w10002_,
		_w10003_,
		_w10004_
	);
	LUT2 #(
		.INIT('h8)
	) name7859 (
		\u1_slt6_reg[8]/P0001 ,
		_w9869_,
		_w10005_
	);
	LUT2 #(
		.INIT('h8)
	) name7860 (
		\u1_slt6_reg[6]/P0001 ,
		_w5936_,
		_w10006_
	);
	LUT2 #(
		.INIT('h8)
	) name7861 (
		\u11_din_tmp1_reg[6]/P0001 ,
		_w3064_,
		_w10007_
	);
	LUT2 #(
		.INIT('h1)
	) name7862 (
		_w10005_,
		_w10006_,
		_w10008_
	);
	LUT2 #(
		.INIT('h4)
	) name7863 (
		_w10007_,
		_w10008_,
		_w10009_
	);
	LUT2 #(
		.INIT('h8)
	) name7864 (
		\u1_slt6_reg[9]/P0001 ,
		_w9869_,
		_w10010_
	);
	LUT2 #(
		.INIT('h8)
	) name7865 (
		\u1_slt6_reg[7]/P0001 ,
		_w5936_,
		_w10011_
	);
	LUT2 #(
		.INIT('h8)
	) name7866 (
		\u11_din_tmp1_reg[7]/P0001 ,
		_w3064_,
		_w10012_
	);
	LUT2 #(
		.INIT('h1)
	) name7867 (
		_w10010_,
		_w10011_,
		_w10013_
	);
	LUT2 #(
		.INIT('h4)
	) name7868 (
		_w10012_,
		_w10013_,
		_w10014_
	);
	LUT2 #(
		.INIT('h8)
	) name7869 (
		\u1_slt6_reg[10]/P0001 ,
		_w9869_,
		_w10015_
	);
	LUT2 #(
		.INIT('h8)
	) name7870 (
		\u1_slt6_reg[8]/P0001 ,
		_w5936_,
		_w10016_
	);
	LUT2 #(
		.INIT('h8)
	) name7871 (
		\u11_din_tmp1_reg[8]/P0001 ,
		_w3064_,
		_w10017_
	);
	LUT2 #(
		.INIT('h1)
	) name7872 (
		_w10015_,
		_w10016_,
		_w10018_
	);
	LUT2 #(
		.INIT('h4)
	) name7873 (
		_w10017_,
		_w10018_,
		_w10019_
	);
	LUT2 #(
		.INIT('h8)
	) name7874 (
		\u1_slt6_reg[9]/P0001 ,
		_w5936_,
		_w10020_
	);
	LUT2 #(
		.INIT('h8)
	) name7875 (
		\u1_slt6_reg[11]/P0001 ,
		_w9869_,
		_w10021_
	);
	LUT2 #(
		.INIT('h8)
	) name7876 (
		\u11_din_tmp1_reg[9]/P0001 ,
		_w3064_,
		_w10022_
	);
	LUT2 #(
		.INIT('h1)
	) name7877 (
		_w10020_,
		_w10021_,
		_w10023_
	);
	LUT2 #(
		.INIT('h4)
	) name7878 (
		_w10022_,
		_w10023_,
		_w10024_
	);
	LUT2 #(
		.INIT('h8)
	) name7879 (
		\u1_slt4_reg[4]/P0001 ,
		_w9796_,
		_w10025_
	);
	LUT2 #(
		.INIT('h8)
	) name7880 (
		\u1_slt4_reg[2]/P0001 ,
		_w5671_,
		_w10026_
	);
	LUT2 #(
		.INIT('h8)
	) name7881 (
		\u10_din_tmp1_reg[2]/P0001 ,
		_w3501_,
		_w10027_
	);
	LUT2 #(
		.INIT('h1)
	) name7882 (
		_w10025_,
		_w10026_,
		_w10028_
	);
	LUT2 #(
		.INIT('h4)
	) name7883 (
		_w10027_,
		_w10028_,
		_w10029_
	);
	LUT2 #(
		.INIT('h8)
	) name7884 (
		\u1_slt4_reg[6]/P0001 ,
		_w9796_,
		_w10030_
	);
	LUT2 #(
		.INIT('h8)
	) name7885 (
		\u1_slt4_reg[4]/P0001 ,
		_w5671_,
		_w10031_
	);
	LUT2 #(
		.INIT('h8)
	) name7886 (
		\u10_din_tmp1_reg[4]/P0001 ,
		_w3501_,
		_w10032_
	);
	LUT2 #(
		.INIT('h1)
	) name7887 (
		_w10030_,
		_w10031_,
		_w10033_
	);
	LUT2 #(
		.INIT('h4)
	) name7888 (
		_w10032_,
		_w10033_,
		_w10034_
	);
	LUT2 #(
		.INIT('h8)
	) name7889 (
		\u1_slt4_reg[7]/P0001 ,
		_w9796_,
		_w10035_
	);
	LUT2 #(
		.INIT('h8)
	) name7890 (
		\u1_slt4_reg[5]/P0001 ,
		_w5671_,
		_w10036_
	);
	LUT2 #(
		.INIT('h8)
	) name7891 (
		\u10_din_tmp1_reg[5]/P0001 ,
		_w3501_,
		_w10037_
	);
	LUT2 #(
		.INIT('h1)
	) name7892 (
		_w10035_,
		_w10036_,
		_w10038_
	);
	LUT2 #(
		.INIT('h4)
	) name7893 (
		_w10037_,
		_w10038_,
		_w10039_
	);
	LUT2 #(
		.INIT('h8)
	) name7894 (
		\u1_slt4_reg[8]/P0001 ,
		_w9796_,
		_w10040_
	);
	LUT2 #(
		.INIT('h8)
	) name7895 (
		\u1_slt4_reg[6]/P0001 ,
		_w5671_,
		_w10041_
	);
	LUT2 #(
		.INIT('h8)
	) name7896 (
		\u10_din_tmp1_reg[6]/P0001 ,
		_w3501_,
		_w10042_
	);
	LUT2 #(
		.INIT('h1)
	) name7897 (
		_w10040_,
		_w10041_,
		_w10043_
	);
	LUT2 #(
		.INIT('h4)
	) name7898 (
		_w10042_,
		_w10043_,
		_w10044_
	);
	LUT2 #(
		.INIT('h8)
	) name7899 (
		\u1_slt4_reg[9]/P0001 ,
		_w9796_,
		_w10045_
	);
	LUT2 #(
		.INIT('h8)
	) name7900 (
		\u1_slt4_reg[7]/P0001 ,
		_w5671_,
		_w10046_
	);
	LUT2 #(
		.INIT('h8)
	) name7901 (
		\u10_din_tmp1_reg[7]/P0001 ,
		_w3501_,
		_w10047_
	);
	LUT2 #(
		.INIT('h1)
	) name7902 (
		_w10045_,
		_w10046_,
		_w10048_
	);
	LUT2 #(
		.INIT('h4)
	) name7903 (
		_w10047_,
		_w10048_,
		_w10049_
	);
	LUT2 #(
		.INIT('h8)
	) name7904 (
		\u1_slt4_reg[10]/P0001 ,
		_w9796_,
		_w10050_
	);
	LUT2 #(
		.INIT('h8)
	) name7905 (
		\u1_slt4_reg[8]/P0001 ,
		_w5671_,
		_w10051_
	);
	LUT2 #(
		.INIT('h8)
	) name7906 (
		\u10_din_tmp1_reg[8]/P0001 ,
		_w3501_,
		_w10052_
	);
	LUT2 #(
		.INIT('h1)
	) name7907 (
		_w10050_,
		_w10051_,
		_w10053_
	);
	LUT2 #(
		.INIT('h4)
	) name7908 (
		_w10052_,
		_w10053_,
		_w10054_
	);
	LUT2 #(
		.INIT('h8)
	) name7909 (
		\u1_slt6_reg[17]/P0001 ,
		_w9869_,
		_w10055_
	);
	LUT2 #(
		.INIT('h8)
	) name7910 (
		\u1_slt6_reg[15]/P0001 ,
		_w5936_,
		_w10056_
	);
	LUT2 #(
		.INIT('h8)
	) name7911 (
		\u11_din_tmp1_reg[15]/P0001 ,
		_w3064_,
		_w10057_
	);
	LUT2 #(
		.INIT('h1)
	) name7912 (
		_w10055_,
		_w10056_,
		_w10058_
	);
	LUT2 #(
		.INIT('h4)
	) name7913 (
		_w10057_,
		_w10058_,
		_w10059_
	);
	LUT2 #(
		.INIT('h8)
	) name7914 (
		\u1_slt3_reg[0]/P0001 ,
		_w5701_,
		_w10060_
	);
	LUT2 #(
		.INIT('h8)
	) name7915 (
		\u1_slt3_reg[2]/P0001 ,
		_w9804_,
		_w10061_
	);
	LUT2 #(
		.INIT('h8)
	) name7916 (
		\u9_din_tmp1_reg[0]/P0001 ,
		_w3311_,
		_w10062_
	);
	LUT2 #(
		.INIT('h1)
	) name7917 (
		_w10060_,
		_w10061_,
		_w10063_
	);
	LUT2 #(
		.INIT('h4)
	) name7918 (
		_w10062_,
		_w10063_,
		_w10064_
	);
	LUT2 #(
		.INIT('h8)
	) name7919 (
		\u1_slt3_reg[4]/P0001 ,
		_w5701_,
		_w10065_
	);
	LUT2 #(
		.INIT('h8)
	) name7920 (
		\u1_slt3_reg[6]/P0001 ,
		_w9804_,
		_w10066_
	);
	LUT2 #(
		.INIT('h8)
	) name7921 (
		\u9_din_tmp1_reg[4]/P0001 ,
		_w3311_,
		_w10067_
	);
	LUT2 #(
		.INIT('h1)
	) name7922 (
		_w10065_,
		_w10066_,
		_w10068_
	);
	LUT2 #(
		.INIT('h4)
	) name7923 (
		_w10067_,
		_w10068_,
		_w10069_
	);
	LUT2 #(
		.INIT('h2)
	) name7924 (
		\u2_cnt_reg[0]/NET0131 ,
		\u2_cnt_reg[5]/NET0131 ,
		_w10070_
	);
	LUT2 #(
		.INIT('h8)
	) name7925 (
		_w9079_,
		_w10070_,
		_w10071_
	);
	LUT2 #(
		.INIT('h8)
	) name7926 (
		_w9109_,
		_w10071_,
		_w10072_
	);
	LUT2 #(
		.INIT('h2)
	) name7927 (
		\u11_mem_reg[0][24]/P0001 ,
		_w5933_,
		_w10073_
	);
	LUT2 #(
		.INIT('h8)
	) name7928 (
		_w5933_,
		_w5975_,
		_w10074_
	);
	LUT2 #(
		.INIT('h1)
	) name7929 (
		_w10073_,
		_w10074_,
		_w10075_
	);
	LUT2 #(
		.INIT('h2)
	) name7930 (
		\u10_mem_reg[0][20]/P0001 ,
		_w5928_,
		_w10076_
	);
	LUT2 #(
		.INIT('h8)
	) name7931 (
		_w5683_,
		_w5928_,
		_w10077_
	);
	LUT2 #(
		.INIT('h1)
	) name7932 (
		_w10076_,
		_w10077_,
		_w10078_
	);
	LUT2 #(
		.INIT('h2)
	) name7933 (
		\u9_mem_reg[0][31]/P0001 ,
		_w5698_,
		_w10079_
	);
	LUT2 #(
		.INIT('h8)
	) name7934 (
		_w5698_,
		_w5789_,
		_w10080_
	);
	LUT2 #(
		.INIT('h1)
	) name7935 (
		_w10079_,
		_w10080_,
		_w10081_
	);
	LUT2 #(
		.INIT('h2)
	) name7936 (
		\u9_mem_reg[0][20]/P0001 ,
		_w5698_,
		_w10082_
	);
	LUT2 #(
		.INIT('h8)
	) name7937 (
		_w5698_,
		_w5741_,
		_w10083_
	);
	LUT2 #(
		.INIT('h1)
	) name7938 (
		_w10082_,
		_w10083_,
		_w10084_
	);
	LUT2 #(
		.INIT('h2)
	) name7939 (
		\u9_mem_reg[0][21]/P0001 ,
		_w5698_,
		_w10085_
	);
	LUT2 #(
		.INIT('h8)
	) name7940 (
		_w5698_,
		_w5745_,
		_w10086_
	);
	LUT2 #(
		.INIT('h1)
	) name7941 (
		_w10085_,
		_w10086_,
		_w10087_
	);
	LUT2 #(
		.INIT('h2)
	) name7942 (
		\u9_mem_reg[0][23]/P0001 ,
		_w5698_,
		_w10088_
	);
	LUT2 #(
		.INIT('h8)
	) name7943 (
		_w5698_,
		_w5757_,
		_w10089_
	);
	LUT2 #(
		.INIT('h1)
	) name7944 (
		_w10088_,
		_w10089_,
		_w10090_
	);
	LUT2 #(
		.INIT('h2)
	) name7945 (
		\u9_mem_reg[0][24]/P0001 ,
		_w5698_,
		_w10091_
	);
	LUT2 #(
		.INIT('h8)
	) name7946 (
		_w5698_,
		_w5761_,
		_w10092_
	);
	LUT2 #(
		.INIT('h1)
	) name7947 (
		_w10091_,
		_w10092_,
		_w10093_
	);
	LUT2 #(
		.INIT('h2)
	) name7948 (
		\u9_mem_reg[0][25]/P0001 ,
		_w5698_,
		_w10094_
	);
	LUT2 #(
		.INIT('h8)
	) name7949 (
		_w5698_,
		_w5765_,
		_w10095_
	);
	LUT2 #(
		.INIT('h1)
	) name7950 (
		_w10094_,
		_w10095_,
		_w10096_
	);
	LUT2 #(
		.INIT('h2)
	) name7951 (
		\u9_mem_reg[0][26]/P0001 ,
		_w5698_,
		_w10097_
	);
	LUT2 #(
		.INIT('h8)
	) name7952 (
		_w5698_,
		_w5769_,
		_w10098_
	);
	LUT2 #(
		.INIT('h1)
	) name7953 (
		_w10097_,
		_w10098_,
		_w10099_
	);
	LUT2 #(
		.INIT('h2)
	) name7954 (
		\u9_mem_reg[0][27]/P0001 ,
		_w5698_,
		_w10100_
	);
	LUT2 #(
		.INIT('h8)
	) name7955 (
		_w5698_,
		_w5773_,
		_w10101_
	);
	LUT2 #(
		.INIT('h1)
	) name7956 (
		_w10100_,
		_w10101_,
		_w10102_
	);
	LUT2 #(
		.INIT('h2)
	) name7957 (
		\u9_mem_reg[0][28]/P0001 ,
		_w5698_,
		_w10103_
	);
	LUT2 #(
		.INIT('h8)
	) name7958 (
		_w5698_,
		_w5777_,
		_w10104_
	);
	LUT2 #(
		.INIT('h1)
	) name7959 (
		_w10103_,
		_w10104_,
		_w10105_
	);
	LUT2 #(
		.INIT('h2)
	) name7960 (
		\u9_mem_reg[0][29]/P0001 ,
		_w5698_,
		_w10106_
	);
	LUT2 #(
		.INIT('h8)
	) name7961 (
		_w5698_,
		_w5781_,
		_w10107_
	);
	LUT2 #(
		.INIT('h1)
	) name7962 (
		_w10106_,
		_w10107_,
		_w10108_
	);
	LUT2 #(
		.INIT('h2)
	) name7963 (
		\u9_mem_reg[0][30]/P0001 ,
		_w5698_,
		_w10109_
	);
	LUT2 #(
		.INIT('h8)
	) name7964 (
		_w5698_,
		_w5785_,
		_w10110_
	);
	LUT2 #(
		.INIT('h1)
	) name7965 (
		_w10109_,
		_w10110_,
		_w10111_
	);
	LUT2 #(
		.INIT('h2)
	) name7966 (
		\u11_mem_reg[0][21]/P0001 ,
		_w5933_,
		_w10112_
	);
	LUT2 #(
		.INIT('h8)
	) name7967 (
		_w5933_,
		_w5963_,
		_w10113_
	);
	LUT2 #(
		.INIT('h1)
	) name7968 (
		_w10112_,
		_w10113_,
		_w10114_
	);
	LUT2 #(
		.INIT('h2)
	) name7969 (
		\u10_mem_reg[0][22]/P0001 ,
		_w5928_,
		_w10115_
	);
	LUT2 #(
		.INIT('h8)
	) name7970 (
		_w5691_,
		_w5928_,
		_w10116_
	);
	LUT2 #(
		.INIT('h1)
	) name7971 (
		_w10115_,
		_w10116_,
		_w10117_
	);
	LUT2 #(
		.INIT('h2)
	) name7972 (
		\u11_mem_reg[0][27]/P0001 ,
		_w5933_,
		_w10118_
	);
	LUT2 #(
		.INIT('h8)
	) name7973 (
		_w5933_,
		_w5987_,
		_w10119_
	);
	LUT2 #(
		.INIT('h1)
	) name7974 (
		_w10118_,
		_w10119_,
		_w10120_
	);
	LUT2 #(
		.INIT('h2)
	) name7975 (
		\u11_mem_reg[0][31]/P0001 ,
		_w5933_,
		_w10121_
	);
	LUT2 #(
		.INIT('h8)
	) name7976 (
		_w5933_,
		_w6003_,
		_w10122_
	);
	LUT2 #(
		.INIT('h1)
	) name7977 (
		_w10121_,
		_w10122_,
		_w10123_
	);
	LUT2 #(
		.INIT('h2)
	) name7978 (
		\u11_mem_reg[0][29]/P0001 ,
		_w5933_,
		_w10124_
	);
	LUT2 #(
		.INIT('h8)
	) name7979 (
		_w5933_,
		_w5995_,
		_w10125_
	);
	LUT2 #(
		.INIT('h1)
	) name7980 (
		_w10124_,
		_w10125_,
		_w10126_
	);
	LUT2 #(
		.INIT('h2)
	) name7981 (
		\u11_mem_reg[0][20]/P0001 ,
		_w5933_,
		_w10127_
	);
	LUT2 #(
		.INIT('h8)
	) name7982 (
		_w5933_,
		_w5959_,
		_w10128_
	);
	LUT2 #(
		.INIT('h1)
	) name7983 (
		_w10127_,
		_w10128_,
		_w10129_
	);
	LUT2 #(
		.INIT('h2)
	) name7984 (
		\u11_mem_reg[0][22]/P0001 ,
		_w5933_,
		_w10130_
	);
	LUT2 #(
		.INIT('h8)
	) name7985 (
		_w5933_,
		_w5967_,
		_w10131_
	);
	LUT2 #(
		.INIT('h1)
	) name7986 (
		_w10130_,
		_w10131_,
		_w10132_
	);
	LUT2 #(
		.INIT('h2)
	) name7987 (
		\u11_mem_reg[0][23]/P0001 ,
		_w5933_,
		_w10133_
	);
	LUT2 #(
		.INIT('h8)
	) name7988 (
		_w5933_,
		_w5971_,
		_w10134_
	);
	LUT2 #(
		.INIT('h1)
	) name7989 (
		_w10133_,
		_w10134_,
		_w10135_
	);
	LUT2 #(
		.INIT('h2)
	) name7990 (
		\u11_mem_reg[0][25]/P0001 ,
		_w5933_,
		_w10136_
	);
	LUT2 #(
		.INIT('h8)
	) name7991 (
		_w5933_,
		_w5979_,
		_w10137_
	);
	LUT2 #(
		.INIT('h1)
	) name7992 (
		_w10136_,
		_w10137_,
		_w10138_
	);
	LUT2 #(
		.INIT('h2)
	) name7993 (
		\u10_mem_reg[0][21]/P0001 ,
		_w5928_,
		_w10139_
	);
	LUT2 #(
		.INIT('h8)
	) name7994 (
		_w5687_,
		_w5928_,
		_w10140_
	);
	LUT2 #(
		.INIT('h1)
	) name7995 (
		_w10139_,
		_w10140_,
		_w10141_
	);
	LUT2 #(
		.INIT('h2)
	) name7996 (
		\u11_mem_reg[0][26]/P0001 ,
		_w5933_,
		_w10142_
	);
	LUT2 #(
		.INIT('h8)
	) name7997 (
		_w5933_,
		_w5983_,
		_w10143_
	);
	LUT2 #(
		.INIT('h1)
	) name7998 (
		_w10142_,
		_w10143_,
		_w10144_
	);
	LUT2 #(
		.INIT('h2)
	) name7999 (
		\u10_mem_reg[0][23]/P0001 ,
		_w5928_,
		_w10145_
	);
	LUT2 #(
		.INIT('h8)
	) name8000 (
		_w5695_,
		_w5928_,
		_w10146_
	);
	LUT2 #(
		.INIT('h1)
	) name8001 (
		_w10145_,
		_w10146_,
		_w10147_
	);
	LUT2 #(
		.INIT('h2)
	) name8002 (
		\u11_mem_reg[0][30]/P0001 ,
		_w5933_,
		_w10148_
	);
	LUT2 #(
		.INIT('h8)
	) name8003 (
		_w5933_,
		_w5999_,
		_w10149_
	);
	LUT2 #(
		.INIT('h1)
	) name8004 (
		_w10148_,
		_w10149_,
		_w10150_
	);
	LUT2 #(
		.INIT('h2)
	) name8005 (
		\u10_mem_reg[0][24]/P0001 ,
		_w5928_,
		_w10151_
	);
	LUT2 #(
		.INIT('h8)
	) name8006 (
		_w5714_,
		_w5928_,
		_w10152_
	);
	LUT2 #(
		.INIT('h1)
	) name8007 (
		_w10151_,
		_w10152_,
		_w10153_
	);
	LUT2 #(
		.INIT('h2)
	) name8008 (
		\u10_mem_reg[0][25]/P0001 ,
		_w5928_,
		_w10154_
	);
	LUT2 #(
		.INIT('h8)
	) name8009 (
		_w5718_,
		_w5928_,
		_w10155_
	);
	LUT2 #(
		.INIT('h1)
	) name8010 (
		_w10154_,
		_w10155_,
		_w10156_
	);
	LUT2 #(
		.INIT('h2)
	) name8011 (
		\u10_mem_reg[0][26]/P0001 ,
		_w5928_,
		_w10157_
	);
	LUT2 #(
		.INIT('h8)
	) name8012 (
		_w5722_,
		_w5928_,
		_w10158_
	);
	LUT2 #(
		.INIT('h1)
	) name8013 (
		_w10157_,
		_w10158_,
		_w10159_
	);
	LUT2 #(
		.INIT('h2)
	) name8014 (
		\u10_mem_reg[0][27]/P0001 ,
		_w5928_,
		_w10160_
	);
	LUT2 #(
		.INIT('h8)
	) name8015 (
		_w5726_,
		_w5928_,
		_w10161_
	);
	LUT2 #(
		.INIT('h1)
	) name8016 (
		_w10160_,
		_w10161_,
		_w10162_
	);
	LUT2 #(
		.INIT('h2)
	) name8017 (
		\u10_mem_reg[0][28]/P0001 ,
		_w5928_,
		_w10163_
	);
	LUT2 #(
		.INIT('h8)
	) name8018 (
		_w5730_,
		_w5928_,
		_w10164_
	);
	LUT2 #(
		.INIT('h1)
	) name8019 (
		_w10163_,
		_w10164_,
		_w10165_
	);
	LUT2 #(
		.INIT('h2)
	) name8020 (
		\u11_mem_reg[0][28]/P0001 ,
		_w5933_,
		_w10166_
	);
	LUT2 #(
		.INIT('h8)
	) name8021 (
		_w5933_,
		_w5991_,
		_w10167_
	);
	LUT2 #(
		.INIT('h1)
	) name8022 (
		_w10166_,
		_w10167_,
		_w10168_
	);
	LUT2 #(
		.INIT('h2)
	) name8023 (
		\u10_mem_reg[0][30]/P0001 ,
		_w5928_,
		_w10169_
	);
	LUT2 #(
		.INIT('h8)
	) name8024 (
		_w5793_,
		_w5928_,
		_w10170_
	);
	LUT2 #(
		.INIT('h1)
	) name8025 (
		_w10169_,
		_w10170_,
		_w10171_
	);
	LUT2 #(
		.INIT('h2)
	) name8026 (
		\u10_mem_reg[0][31]/P0001 ,
		_w5928_,
		_w10172_
	);
	LUT2 #(
		.INIT('h8)
	) name8027 (
		_w5797_,
		_w5928_,
		_w10173_
	);
	LUT2 #(
		.INIT('h1)
	) name8028 (
		_w10172_,
		_w10173_,
		_w10174_
	);
	LUT2 #(
		.INIT('h2)
	) name8029 (
		\u10_mem_reg[0][29]/P0001 ,
		_w5928_,
		_w10175_
	);
	LUT2 #(
		.INIT('h8)
	) name8030 (
		_w5749_,
		_w5928_,
		_w10176_
	);
	LUT2 #(
		.INIT('h1)
	) name8031 (
		_w10175_,
		_w10176_,
		_w10177_
	);
	LUT2 #(
		.INIT('h2)
	) name8032 (
		\u9_mem_reg[0][22]/P0001 ,
		_w5698_,
		_w10178_
	);
	LUT2 #(
		.INIT('h8)
	) name8033 (
		_w5698_,
		_w5753_,
		_w10179_
	);
	LUT2 #(
		.INIT('h1)
	) name8034 (
		_w10178_,
		_w10179_,
		_w10180_
	);
	LUT2 #(
		.INIT('h2)
	) name8035 (
		\u2_bit_clk_r1_reg/P0001 ,
		\u2_bit_clk_r_reg/P0001 ,
		_w10181_
	);
	LUT2 #(
		.INIT('h4)
	) name8036 (
		\u2_bit_clk_r1_reg/P0001 ,
		\u2_bit_clk_r_reg/P0001 ,
		_w10182_
	);
	LUT2 #(
		.INIT('h1)
	) name8037 (
		_w10181_,
		_w10182_,
		_w10183_
	);
	LUT2 #(
		.INIT('h4)
	) name8038 (
		\dma_ack_i[6]_pad ,
		\dma_req_o[6]_pad ,
		_w10184_
	);
	LUT2 #(
		.INIT('h4)
	) name8039 (
		\dma_ack_i[6]_pad ,
		\u13_icc_r_reg[6]/NET0131 ,
		_w10185_
	);
	LUT2 #(
		.INIT('h8)
	) name8040 (
		_w4429_,
		_w10185_,
		_w10186_
	);
	LUT2 #(
		.INIT('h8)
	) name8041 (
		\u16_u6_dma_req_r1_reg/P0001 ,
		_w10186_,
		_w10187_
	);
	LUT2 #(
		.INIT('h1)
	) name8042 (
		_w10184_,
		_w10187_,
		_w10188_
	);
	LUT2 #(
		.INIT('h4)
	) name8043 (
		\dma_ack_i[7]_pad ,
		\dma_req_o[7]_pad ,
		_w10189_
	);
	LUT2 #(
		.INIT('h4)
	) name8044 (
		\dma_ack_i[7]_pad ,
		\u13_icc_r_reg[14]/NET0131 ,
		_w10190_
	);
	LUT2 #(
		.INIT('h8)
	) name8045 (
		_w4462_,
		_w10190_,
		_w10191_
	);
	LUT2 #(
		.INIT('h8)
	) name8046 (
		\u16_u7_dma_req_r1_reg/P0001 ,
		_w10191_,
		_w10192_
	);
	LUT2 #(
		.INIT('h1)
	) name8047 (
		_w10189_,
		_w10192_,
		_w10193_
	);
	LUT2 #(
		.INIT('h1)
	) name8048 (
		\u2_sync_beat_reg/P0001 ,
		\u2_sync_resume_reg/NET0131 ,
		_w10194_
	);
	LUT2 #(
		.INIT('h2)
	) name8049 (
		\u3_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w10195_
	);
	LUT2 #(
		.INIT('h8)
	) name8050 (
		\u14_u0_full_empty_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w10196_
	);
	LUT2 #(
		.INIT('h1)
	) name8051 (
		_w10195_,
		_w10196_,
		_w10197_
	);
	LUT2 #(
		.INIT('h2)
	) name8052 (
		\u4_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w10198_
	);
	LUT2 #(
		.INIT('h8)
	) name8053 (
		\u14_u1_full_empty_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w10199_
	);
	LUT2 #(
		.INIT('h1)
	) name8054 (
		_w10198_,
		_w10199_,
		_w10200_
	);
	LUT2 #(
		.INIT('h2)
	) name8055 (
		\u5_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w10201_
	);
	LUT2 #(
		.INIT('h8)
	) name8056 (
		\u14_u2_full_empty_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w10202_
	);
	LUT2 #(
		.INIT('h1)
	) name8057 (
		_w10201_,
		_w10202_,
		_w10203_
	);
	LUT2 #(
		.INIT('h2)
	) name8058 (
		\u6_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w10204_
	);
	LUT2 #(
		.INIT('h8)
	) name8059 (
		\u14_u3_full_empty_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w10205_
	);
	LUT2 #(
		.INIT('h1)
	) name8060 (
		_w10204_,
		_w10205_,
		_w10206_
	);
	LUT2 #(
		.INIT('h2)
	) name8061 (
		\u7_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w10207_
	);
	LUT2 #(
		.INIT('h8)
	) name8062 (
		\u14_u4_full_empty_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w10208_
	);
	LUT2 #(
		.INIT('h1)
	) name8063 (
		_w10207_,
		_w10208_,
		_w10209_
	);
	LUT2 #(
		.INIT('h2)
	) name8064 (
		\u8_empty_reg/NET0131 ,
		\valid_s_reg/NET0131 ,
		_w10210_
	);
	LUT2 #(
		.INIT('h8)
	) name8065 (
		\u14_u5_full_empty_r_reg/P0001 ,
		\valid_s_reg/NET0131 ,
		_w10211_
	);
	LUT2 #(
		.INIT('h1)
	) name8066 (
		_w10210_,
		_w10211_,
		_w10212_
	);
	LUT2 #(
		.INIT('h4)
	) name8067 (
		\in_valid_s_reg[0]/NET0131 ,
		\u9_full_reg/NET0131 ,
		_w10213_
	);
	LUT2 #(
		.INIT('h8)
	) name8068 (
		\in_valid_s_reg[0]/NET0131 ,
		\u14_u6_full_empty_r_reg/P0001 ,
		_w10214_
	);
	LUT2 #(
		.INIT('h1)
	) name8069 (
		_w10213_,
		_w10214_,
		_w10215_
	);
	LUT2 #(
		.INIT('h4)
	) name8070 (
		\in_valid_s_reg[1]/NET0131 ,
		\u10_full_reg/NET0131 ,
		_w10216_
	);
	LUT2 #(
		.INIT('h8)
	) name8071 (
		\in_valid_s_reg[1]/NET0131 ,
		\u14_u7_full_empty_r_reg/P0001 ,
		_w10217_
	);
	LUT2 #(
		.INIT('h1)
	) name8072 (
		_w10216_,
		_w10217_,
		_w10218_
	);
	LUT2 #(
		.INIT('h4)
	) name8073 (
		\in_valid_s_reg[2]/NET0131 ,
		\u11_full_reg/NET0131 ,
		_w10219_
	);
	LUT2 #(
		.INIT('h8)
	) name8074 (
		\in_valid_s_reg[2]/NET0131 ,
		\u14_u8_full_empty_r_reg/P0001 ,
		_w10220_
	);
	LUT2 #(
		.INIT('h1)
	) name8075 (
		_w10219_,
		_w10220_,
		_w10221_
	);
	LUT2 #(
		.INIT('h8)
	) name8076 (
		\u1_sr_reg[11]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w10222_
	);
	LUT2 #(
		.INIT('h2)
	) name8077 (
		\u1_slt0_reg[11]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w10223_
	);
	LUT2 #(
		.INIT('h1)
	) name8078 (
		_w10222_,
		_w10223_,
		_w10224_
	);
	LUT2 #(
		.INIT('h8)
	) name8079 (
		\u1_sr_reg[12]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w10225_
	);
	LUT2 #(
		.INIT('h2)
	) name8080 (
		\u1_slt0_reg[12]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w10226_
	);
	LUT2 #(
		.INIT('h1)
	) name8081 (
		_w10225_,
		_w10226_,
		_w10227_
	);
	LUT2 #(
		.INIT('h8)
	) name8082 (
		\u1_sr_reg[15]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w10228_
	);
	LUT2 #(
		.INIT('h2)
	) name8083 (
		\u1_slt0_reg[15]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w10229_
	);
	LUT2 #(
		.INIT('h1)
	) name8084 (
		_w10228_,
		_w10229_,
		_w10230_
	);
	LUT2 #(
		.INIT('h8)
	) name8085 (
		\u1_sr_reg[9]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w10231_
	);
	LUT2 #(
		.INIT('h2)
	) name8086 (
		\u1_slt0_reg[9]/P0001 ,
		\u2_out_le_reg[0]/P0001 ,
		_w10232_
	);
	LUT2 #(
		.INIT('h1)
	) name8087 (
		_w10231_,
		_w10232_,
		_w10233_
	);
	LUT2 #(
		.INIT('h8)
	) name8088 (
		\u1_sr_reg[10]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10234_
	);
	LUT2 #(
		.INIT('h2)
	) name8089 (
		\u1_slt1_reg[10]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10235_
	);
	LUT2 #(
		.INIT('h1)
	) name8090 (
		_w10234_,
		_w10235_,
		_w10236_
	);
	LUT2 #(
		.INIT('h8)
	) name8091 (
		\u1_sr_reg[11]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10237_
	);
	LUT2 #(
		.INIT('h2)
	) name8092 (
		\u1_slt1_reg[11]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10238_
	);
	LUT2 #(
		.INIT('h1)
	) name8093 (
		_w10237_,
		_w10238_,
		_w10239_
	);
	LUT2 #(
		.INIT('h8)
	) name8094 (
		\u1_sr_reg[5]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10240_
	);
	LUT2 #(
		.INIT('h2)
	) name8095 (
		\u1_slt1_reg[5]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10241_
	);
	LUT2 #(
		.INIT('h1)
	) name8096 (
		_w10240_,
		_w10241_,
		_w10242_
	);
	LUT2 #(
		.INIT('h8)
	) name8097 (
		\u1_sr_reg[6]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10243_
	);
	LUT2 #(
		.INIT('h2)
	) name8098 (
		\u1_slt1_reg[6]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10244_
	);
	LUT2 #(
		.INIT('h1)
	) name8099 (
		_w10243_,
		_w10244_,
		_w10245_
	);
	LUT2 #(
		.INIT('h8)
	) name8100 (
		\u1_sr_reg[7]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10246_
	);
	LUT2 #(
		.INIT('h2)
	) name8101 (
		\u1_slt1_reg[7]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10247_
	);
	LUT2 #(
		.INIT('h1)
	) name8102 (
		_w10246_,
		_w10247_,
		_w10248_
	);
	LUT2 #(
		.INIT('h8)
	) name8103 (
		\u1_sr_reg[8]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10249_
	);
	LUT2 #(
		.INIT('h2)
	) name8104 (
		\u1_slt1_reg[8]/P0001 ,
		\u2_out_le_reg[1]/P0001 ,
		_w10250_
	);
	LUT2 #(
		.INIT('h1)
	) name8105 (
		_w10249_,
		_w10250_,
		_w10251_
	);
	assign \_al_n1  = 1'b0;
	assign \g16/_0_  = _w2157_ ;
	assign \g23/_0_  = _w2168_ ;
	assign \g29500/_0_  = _w2178_ ;
	assign \g29503/_3_  = _w2181_ ;
	assign \g29505/_3_  = _w2183_ ;
	assign \g29507/_3_  = _w2186_ ;
	assign \g29509/_3_  = _w2189_ ;
	assign \g29511/_0_  = _w2190_ ;
	assign \g29513/_3_  = _w2193_ ;
	assign \g29515/_3_  = _w2196_ ;
	assign \g29517/_3_  = _w2199_ ;
	assign \g29519/_0_  = _w2202_ ;
	assign \g29522/_0_  = _w2203_ ;
	assign \g29524/_0_  = _w2204_ ;
	assign \g29526/_0_  = _w2205_ ;
	assign \g29528/_0_  = _w2206_ ;
	assign \g29530/_0_  = _w2207_ ;
	assign \g29532/_0_  = _w2208_ ;
	assign \g29534/_3_  = _w2211_ ;
	assign \g29536/_3_  = _w2214_ ;
	assign \g29538/_3_  = _w2217_ ;
	assign \g29540/_3_  = _w2220_ ;
	assign \g29542/_3_  = _w2223_ ;
	assign \g29544/_3_  = _w2226_ ;
	assign \g29546/_3_  = _w2229_ ;
	assign \g29548/_3_  = _w2232_ ;
	assign \g29550/_0_  = _w2233_ ;
	assign \g29552/_0_  = _w2234_ ;
	assign \g29554/_0_  = _w2235_ ;
	assign \g29556/_0_  = _w2236_ ;
	assign \g29558/_0_  = _w2237_ ;
	assign \g29560/_0_  = _w2238_ ;
	assign \g29562/_0_  = _w2239_ ;
	assign \g29564/_0_  = _w2240_ ;
	assign \g29566/_0_  = _w2241_ ;
	assign \g29568/_0_  = _w2242_ ;
	assign \g29570/_0_  = _w2243_ ;
	assign \g29572/_0_  = _w2244_ ;
	assign \g29574/_3_  = _w2247_ ;
	assign \g29576/_3_  = _w2250_ ;
	assign \g29578/_3_  = _w2253_ ;
	assign \g29580/_3_  = _w2256_ ;
	assign \g29582/_3_  = _w2259_ ;
	assign \g29584/_3_  = _w2262_ ;
	assign \g29586/_3_  = _w2265_ ;
	assign \g29588/_3_  = _w2268_ ;
	assign \g29590/_3_  = _w2271_ ;
	assign \g29592/_3_  = _w2274_ ;
	assign \g29594/_3_  = _w2277_ ;
	assign \g29596/_3_  = _w2280_ ;
	assign \g29598/_3_  = _w2283_ ;
	assign \g29600/_3_  = _w2286_ ;
	assign \g29602/_3_  = _w2289_ ;
	assign \g29604/_3_  = _w2292_ ;
	assign \g29606/_0_  = _w2293_ ;
	assign \g29608/_0_  = _w2294_ ;
	assign \g29610/_0_  = _w2295_ ;
	assign \g29612/_0_  = _w2296_ ;
	assign \g29614/_3_  = _w2299_ ;
	assign \g29616/_3_  = _w2302_ ;
	assign \g29618/_3_  = _w2305_ ;
	assign \g29620/_3_  = _w2308_ ;
	assign \g29622/_3_  = _w2311_ ;
	assign \g29624/_3_  = _w2314_ ;
	assign \g29626/_3_  = _w2317_ ;
	assign \g29628/_3_  = _w2320_ ;
	assign \g29630/_3_  = _w2323_ ;
	assign \g29632/_3_  = _w2326_ ;
	assign \g29634/_3_  = _w2329_ ;
	assign \g29636/_3_  = _w2332_ ;
	assign \g29638/_3_  = _w2335_ ;
	assign \g29640/_3_  = _w2338_ ;
	assign \g29642/_3_  = _w2341_ ;
	assign \g29644/_3_  = _w2344_ ;
	assign \g29646/_3_  = _w2347_ ;
	assign \g29648/_3_  = _w2350_ ;
	assign \g29650/_3_  = _w2353_ ;
	assign \g29652/_3_  = _w2356_ ;
	assign \g29654/_3_  = _w2359_ ;
	assign \g29656/_3_  = _w2362_ ;
	assign \g29658/_3_  = _w2365_ ;
	assign \g29660/_3_  = _w2368_ ;
	assign \g29662/_3_  = _w2371_ ;
	assign \g29664/_3_  = _w2374_ ;
	assign \g29666/_3_  = _w2377_ ;
	assign \g29668/_3_  = _w2380_ ;
	assign \g29670/_3_  = _w2383_ ;
	assign \g29672/_3_  = _w2386_ ;
	assign \g29674/_3_  = _w2389_ ;
	assign \g29676/_3_  = _w2392_ ;
	assign \g29678/_3_  = _w2395_ ;
	assign \g29680/_3_  = _w2398_ ;
	assign \g29682/_3_  = _w2401_ ;
	assign \g29684/_3_  = _w2404_ ;
	assign \g29686/_3_  = _w2407_ ;
	assign \g29688/_3_  = _w2410_ ;
	assign \g29690/_3_  = _w2413_ ;
	assign \g29692/_3_  = _w2416_ ;
	assign \g29694/_0_  = _w2417_ ;
	assign \g29696/_0_  = _w2418_ ;
	assign \g29698/_0_  = _w2419_ ;
	assign \g29700/_0_  = _w2420_ ;
	assign \g29702/_0_  = _w2421_ ;
	assign \g29704/_0_  = _w2422_ ;
	assign \g29706/_0_  = _w2423_ ;
	assign \g29708/_0_  = _w2424_ ;
	assign \g29710/_0_  = _w2425_ ;
	assign \g29712/_0_  = _w2426_ ;
	assign \g29714/_0_  = _w2427_ ;
	assign \g29716/_0_  = _w2428_ ;
	assign \g29718/_0_  = _w2429_ ;
	assign \g29720/_0_  = _w2430_ ;
	assign \g29722/_0_  = _w2431_ ;
	assign \g29724/_0_  = _w2432_ ;
	assign \g29726/_0_  = _w2433_ ;
	assign \g29728/_0_  = _w2434_ ;
	assign \g29730/_0_  = _w2435_ ;
	assign \g29732/_0_  = _w2436_ ;
	assign \g29734/_3_  = _w2439_ ;
	assign \g29736/_3_  = _w2442_ ;
	assign \g29738/_3_  = _w2445_ ;
	assign \g29740/_3_  = _w2448_ ;
	assign \g29742/_3_  = _w2451_ ;
	assign \g29744/_3_  = _w2454_ ;
	assign \g29746/_3_  = _w2457_ ;
	assign \g29748/_3_  = _w2460_ ;
	assign \g29750/_3_  = _w2463_ ;
	assign \g29752/_3_  = _w2466_ ;
	assign \g29754/_3_  = _w2469_ ;
	assign \g29756/_3_  = _w2472_ ;
	assign \g29758/_3_  = _w2475_ ;
	assign \g29760/_3_  = _w2478_ ;
	assign \g29762/_3_  = _w2481_ ;
	assign \g29764/_3_  = _w2484_ ;
	assign \g29766/_3_  = _w2487_ ;
	assign \g29768/_3_  = _w2490_ ;
	assign \g29770/_3_  = _w2493_ ;
	assign \g29772/_3_  = _w2496_ ;
	assign \g29774/_3_  = _w2499_ ;
	assign \g29776/_3_  = _w2502_ ;
	assign \g29778/_3_  = _w2505_ ;
	assign \g29780/_3_  = _w2508_ ;
	assign \g29782/_3_  = _w2511_ ;
	assign \g29784/_3_  = _w2514_ ;
	assign \g29786/_3_  = _w2517_ ;
	assign \g29788/_3_  = _w2520_ ;
	assign \g29790/_3_  = _w2523_ ;
	assign \g29792/_3_  = _w2526_ ;
	assign \g29794/_3_  = _w2529_ ;
	assign \g29796/_3_  = _w2532_ ;
	assign \g29798/_3_  = _w2535_ ;
	assign \g29800/_3_  = _w2538_ ;
	assign \g29802/_3_  = _w2541_ ;
	assign \g29804/_3_  = _w2544_ ;
	assign \g29806/_3_  = _w2547_ ;
	assign \g29808/_3_  = _w2550_ ;
	assign \g29810/_3_  = _w2553_ ;
	assign \g29812/_3_  = _w2556_ ;
	assign \g29814/_3_  = _w2559_ ;
	assign \g29816/_3_  = _w2562_ ;
	assign \g29818/_3_  = _w2565_ ;
	assign \g29820/_3_  = _w2568_ ;
	assign \g29822/_3_  = _w2571_ ;
	assign \g29824/_3_  = _w2574_ ;
	assign \g29826/_3_  = _w2577_ ;
	assign \g29828/_3_  = _w2580_ ;
	assign \g29830/_3_  = _w2583_ ;
	assign \g29832/_3_  = _w2586_ ;
	assign \g29834/_3_  = _w2589_ ;
	assign \g29836/_3_  = _w2592_ ;
	assign \g29838/_3_  = _w2595_ ;
	assign \g29840/_3_  = _w2598_ ;
	assign \g29842/_3_  = _w2601_ ;
	assign \g29844/_3_  = _w2604_ ;
	assign \g29846/_3_  = _w2607_ ;
	assign \g29848/_3_  = _w2610_ ;
	assign \g29850/_3_  = _w2613_ ;
	assign \g29852/_3_  = _w2616_ ;
	assign \g29854/_3_  = _w2619_ ;
	assign \g29856/_3_  = _w2622_ ;
	assign \g29858/_3_  = _w2625_ ;
	assign \g29860/_3_  = _w2628_ ;
	assign \g29862/_3_  = _w2631_ ;
	assign \g29864/_3_  = _w2634_ ;
	assign \g29866/_3_  = _w2637_ ;
	assign \g29868/_3_  = _w2640_ ;
	assign \g29870/_3_  = _w2643_ ;
	assign \g29872/_3_  = _w2646_ ;
	assign \g29874/_3_  = _w2649_ ;
	assign \g29876/_3_  = _w2652_ ;
	assign \g29878/_3_  = _w2655_ ;
	assign \g29880/_3_  = _w2658_ ;
	assign \g29904/_0_  = _w2670_ ;
	assign \g29905/_0_  = _w2682_ ;
	assign \g29906/_0_  = _w2694_ ;
	assign \g29907/_0_  = _w2706_ ;
	assign \g29908/_0_  = _w2718_ ;
	assign \g29909/_0_  = _w2730_ ;
	assign \g29914/_3_  = _w2733_ ;
	assign \g29952/_0_  = _w2744_ ;
	assign \g29953/_0_  = _w2746_ ;
	assign \g29954/_0_  = _w2748_ ;
	assign \g29955/_0_  = _w2750_ ;
	assign \g29956/_0_  = _w2752_ ;
	assign \g29957/_0_  = _w2754_ ;
	assign \g29975/_0_  = _w2668_ ;
	assign \g29976/_0_  = _w2680_ ;
	assign \g29977/_0_  = _w2692_ ;
	assign \g29978/_0_  = _w2704_ ;
	assign \g29979/_0_  = _w2716_ ;
	assign \g29980/_0_  = _w2728_ ;
	assign \g29989/_3_  = _w2757_ ;
	assign \g30020/_0_  = _w2768_ ;
	assign \g30021/_0_  = _w2779_ ;
	assign \g30045/_0_  = _w2783_ ;
	assign \g30046/_0_  = _w2793_ ;
	assign \g30047/_0_  = _w2804_ ;
	assign \g30048/_0_  = _w2814_ ;
	assign \g30049/_0_  = _w2666_ ;
	assign \g30050/_0_  = _w2678_ ;
	assign \g30051/_0_  = _w2690_ ;
	assign \g30052/_0_  = _w2702_ ;
	assign \g30053/_0_  = _w2714_ ;
	assign \g30054/_0_  = _w2726_ ;
	assign \g30062/_0_  = _w2818_ ;
	assign \g30063/_0_  = _w2822_ ;
	assign \g30064/_0_  = _w2824_ ;
	assign \g30065/_0_  = _w2826_ ;
	assign \g30066/_0_  = _w2828_ ;
	assign \g30067/_0_  = _w2832_ ;
	assign \g30068/_0_  = _w2836_ ;
	assign \g30069/_0_  = _w2840_ ;
	assign \g30070/_0_  = _w2843_ ;
	assign \g30071/_0_  = _w2846_ ;
	assign \g30072/_0_  = _w2849_ ;
	assign \g30073/_0_  = _w2852_ ;
	assign \g30074/_0_  = _w2855_ ;
	assign \g30075/_0_  = _w2858_ ;
	assign \g30136/_3_  = _w2861_ ;
	assign \g30707/_0_  = _w2867_ ;
	assign \g30708/_0_  = _w2872_ ;
	assign \g30711/_0_  = _w2877_ ;
	assign \g30714/_0_  = _w2882_ ;
	assign \g30715/_0_  = _w2887_ ;
	assign \g30720/_0_  = _w2892_ ;
	assign \g30725/_0_  = _w2897_ ;
	assign \g30741/_0_  = _w2914_ ;
	assign \g30742/_0_  = _w2924_ ;
	assign \g30743/_0_  = _w2941_ ;
	assign \g30744/_0_  = _w2951_ ;
	assign \g30745/_0_  = _w2968_ ;
	assign \g30746/_0_  = _w2978_ ;
	assign \g30747/_0_  = _w2996_ ;
	assign \g30748/_0_  = _w3006_ ;
	assign \g30749/_0_  = _w3024_ ;
	assign \g30750/_0_  = _w3041_ ;
	assign \g30751/_0_  = _w3051_ ;
	assign \g30752/_0_  = _w3061_ ;
	assign \g30789/_0_  = _w3071_ ;
	assign \g30790/_0_  = _w3112_ ;
	assign \g30791/_0_  = _w3152_ ;
	assign \g30792/_0_  = _w3178_ ;
	assign \g30793/_0_  = _w3204_ ;
	assign \g30794/_0_  = _w3230_ ;
	assign \g30795/_0_  = _w3256_ ;
	assign \g30796/_0_  = _w3282_ ;
	assign \g30797/_0_  = _w3308_ ;
	assign \g30798/_0_  = _w3318_ ;
	assign \g30799/_0_  = _w3344_ ;
	assign \g30800/_0_  = _w3370_ ;
	assign \g30801/_0_  = _w3384_ ;
	assign \g30802/_0_  = _w3398_ ;
	assign \g30803/_0_  = _w3417_ ;
	assign \g30804/_0_  = _w3436_ ;
	assign \g30805/_0_  = _w3448_ ;
	assign \g30806/_0_  = _w3460_ ;
	assign \g30807/_0_  = _w3479_ ;
	assign \g30808/_0_  = _w3498_ ;
	assign \g30809/_0_  = _w3508_ ;
	assign \g30810/_0_  = _w3549_ ;
	assign \g30811/_0_  = _w3589_ ;
	assign \g30812/_0_  = _w3615_ ;
	assign \g30813/_0_  = _w3641_ ;
	assign \g30814/_0_  = _w3667_ ;
	assign \g30815/_0_  = _w3693_ ;
	assign \g30816/_0_  = _w3719_ ;
	assign \g30817/_0_  = _w3745_ ;
	assign \g30818/_0_  = _w3771_ ;
	assign \g30819/_0_  = _w3797_ ;
	assign \g30820/_0_  = _w3811_ ;
	assign \g30821/_0_  = _w3825_ ;
	assign \g30822/_0_  = _w3844_ ;
	assign \g30823/_0_  = _w3863_ ;
	assign \g30824/_0_  = _w3875_ ;
	assign \g30825/_0_  = _w3887_ ;
	assign \g30826/_0_  = _w3906_ ;
	assign \g30827/_0_  = _w3925_ ;
	assign \g30828/_0_  = _w3966_ ;
	assign \g30829/_0_  = _w4006_ ;
	assign \g30830/_0_  = _w4032_ ;
	assign \g30831/_0_  = _w4058_ ;
	assign \g30832/_0_  = _w4084_ ;
	assign \g30833/_0_  = _w4110_ ;
	assign \g30834/_0_  = _w4136_ ;
	assign \g30835/_0_  = _w4162_ ;
	assign \g30836/_0_  = _w4188_ ;
	assign \g30837/_0_  = _w4214_ ;
	assign \g30838/_0_  = _w4228_ ;
	assign \g30839/_0_  = _w4242_ ;
	assign \g30840/_0_  = _w4261_ ;
	assign \g30841/_0_  = _w4280_ ;
	assign \g30842/_0_  = _w4292_ ;
	assign \g30843/_0_  = _w4304_ ;
	assign \g30844/_0_  = _w4323_ ;
	assign \g30845/_0_  = _w4342_ ;
	assign \g30846/_0_  = _w4383_ ;
	assign \g30847/_0_  = _w4422_ ;
	assign \g30848/_0_  = _w4429_ ;
	assign \g30849/_0_  = _w4455_ ;
	assign \g30850/_0_  = _w4462_ ;
	assign \g30851/_0_  = _w4488_ ;
	assign \g30852/_0_  = _w4514_ ;
	assign \g30853/_0_  = _w2153_ ;
	assign \g30854/_0_  = _w4539_ ;
	assign \g30855/_0_  = _w4565_ ;
	assign \g30856/_0_  = _w4591_ ;
	assign \g30857/_0_  = _w4617_ ;
	assign \g30858/_0_  = _w4643_ ;
	assign \g30859/_0_  = _w4657_ ;
	assign \g30860/_0_  = _w4671_ ;
	assign \g30861/_0_  = _w4690_ ;
	assign \g30862/_0_  = _w4709_ ;
	assign \g30863/_0_  = _w4721_ ;
	assign \g30864/_0_  = _w4733_ ;
	assign \g30865/_0_  = _w4752_ ;
	assign \g30866/_0_  = _w4771_ ;
	assign \g30867/_0_  = _w4812_ ;
	assign \g30868/_0_  = _w4852_ ;
	assign \g30869/_0_  = _w4878_ ;
	assign \g30870/_0_  = _w4903_ ;
	assign \g30871/_0_  = _w4929_ ;
	assign \g30872/_0_  = _w4955_ ;
	assign \g30873/_0_  = _w4981_ ;
	assign \g30874/_0_  = _w5006_ ;
	assign \g30875/_0_  = _w5032_ ;
	assign \g30876/_0_  = _w5073_ ;
	assign \g30877/_0_  = _w5099_ ;
	assign \g30878/_0_  = _w5139_ ;
	assign \g30879/_0_  = _w5165_ ;
	assign \g30880/_0_  = _w5179_ ;
	assign \g30881/_0_  = _w5205_ ;
	assign \g30882/_0_  = _w5219_ ;
	assign \g30883/_0_  = _w5245_ ;
	assign \g30884/_0_  = _w5264_ ;
	assign \g30885/_0_  = _w5290_ ;
	assign \g30886/_0_  = _w5309_ ;
	assign \g30887/_0_  = _w5335_ ;
	assign \g30888/_0_  = _w5361_ ;
	assign \g30889/_0_  = _w5373_ ;
	assign \g30890/_0_  = _w5385_ ;
	assign \g30891/_0_  = _w5411_ ;
	assign \g30892/_0_  = _w5430_ ;
	assign \g30893/_0_  = _w5456_ ;
	assign \g30894/_0_  = _w5475_ ;
	assign \g30895/_0_  = _w5489_ ;
	assign \g30896/_0_  = _w5503_ ;
	assign \g30897/_0_  = _w5522_ ;
	assign \g30898/_0_  = _w5541_ ;
	assign \g30899/_0_  = _w5553_ ;
	assign \g30900/_0_  = _w5565_ ;
	assign \g30901/_0_  = _w5584_ ;
	assign \g30902/_0_  = _w5603_ ;
	assign \g30906/_0_  = _w5606_ ;
	assign \g30907/_0_  = _w5609_ ;
	assign \g30908/_0_  = _w5612_ ;
	assign \g30909/_0_  = _w5616_ ;
	assign \g30910/_0_  = _w5620_ ;
	assign \g30911/_0_  = _w5624_ ;
	assign \g30918/_0_  = _w5631_ ;
	assign \g30919/_0_  = _w5634_ ;
	assign \g30920/_0_  = _w5639_ ;
	assign \g30921/_0_  = _w5643_ ;
	assign \g30922/_0_  = _w5647_ ;
	assign \g30923/_0_  = _w5651_ ;
	assign \g30924/_0_  = _w5656_ ;
	assign \g30925/_0_  = _w5661_ ;
	assign \g30926/_0_  = _w5666_ ;
	assign \g30946/_0_  = _w5675_ ;
	assign \g30947/_0_  = _w5681_ ;
	assign \g30948/_0_  = _w5685_ ;
	assign \g30949/_0_  = _w5689_ ;
	assign \g30950/_0_  = _w5693_ ;
	assign \g30951/_0_  = _w5697_ ;
	assign \g30952/_0_  = _w5706_ ;
	assign \g30953/_0_  = _w5712_ ;
	assign \g30954/_0_  = _w5716_ ;
	assign \g30955/_0_  = _w5720_ ;
	assign \g30956/_0_  = _w5724_ ;
	assign \g30957/_0_  = _w5728_ ;
	assign \g30958/_0_  = _w5732_ ;
	assign \g30959/_0_  = _w5736_ ;
	assign \g30960/_0_  = _w5739_ ;
	assign \g30961/_0_  = _w5743_ ;
	assign \g30962/_0_  = _w5747_ ;
	assign \g30963/_0_  = _w5751_ ;
	assign \g30964/_0_  = _w5755_ ;
	assign \g30965/_0_  = _w5759_ ;
	assign \g30966/_0_  = _w5763_ ;
	assign \g30967/_0_  = _w5767_ ;
	assign \g30968/_0_  = _w5771_ ;
	assign \g30969/_0_  = _w5775_ ;
	assign \g30970/_0_  = _w5779_ ;
	assign \g30971/_0_  = _w5783_ ;
	assign \g30972/_0_  = _w5787_ ;
	assign \g30973/_0_  = _w5791_ ;
	assign \g30974/_0_  = _w5795_ ;
	assign \g30975/_0_  = _w5799_ ;
	assign \g30976/_0_  = _w5804_ ;
	assign \g30977/_0_  = _w5807_ ;
	assign \g30978/_0_  = _w5810_ ;
	assign \g30979/_0_  = _w5813_ ;
	assign \g30980/_0_  = _w5816_ ;
	assign \g30981/_0_  = _w5819_ ;
	assign \g30982/_0_  = _w5822_ ;
	assign \g30983/_0_  = _w5825_ ;
	assign \g30984/_0_  = _w5828_ ;
	assign \g30985/_0_  = _w5831_ ;
	assign \g30986/_0_  = _w5834_ ;
	assign \g30987/_0_  = _w5837_ ;
	assign \g30988/_0_  = _w5840_ ;
	assign \g30989/_0_  = _w5843_ ;
	assign \g30990/_0_  = _w5846_ ;
	assign \g30991/_0_  = _w5849_ ;
	assign \g30992/_0_  = _w5852_ ;
	assign \g30993/_0_  = _w5855_ ;
	assign \g30994/_0_  = _w5858_ ;
	assign \g30995/_0_  = _w5861_ ;
	assign \g30996/_0_  = _w5864_ ;
	assign \g30997/_0_  = _w5867_ ;
	assign \g30998/_0_  = _w5870_ ;
	assign \g30999/_0_  = _w5873_ ;
	assign \g31000/_0_  = _w5876_ ;
	assign \g31001/_0_  = _w5879_ ;
	assign \g31002/_0_  = _w5882_ ;
	assign \g31003/_0_  = _w5885_ ;
	assign \g31004/_0_  = _w5888_ ;
	assign \g31005/_0_  = _w5891_ ;
	assign \g31006/_0_  = _w5894_ ;
	assign \g31007/_0_  = _w5897_ ;
	assign \g31008/_0_  = _w5900_ ;
	assign \g31009/_0_  = _w5903_ ;
	assign \g31010/_0_  = _w5906_ ;
	assign \g31011/_0_  = _w5909_ ;
	assign \g31012/_0_  = _w5912_ ;
	assign \g31013/_0_  = _w5915_ ;
	assign \g31014/_0_  = _w5918_ ;
	assign \g31015/_0_  = _w5921_ ;
	assign \g31016/_0_  = _w5924_ ;
	assign \g31017/_0_  = _w5927_ ;
	assign \g31018/_0_  = _w5932_ ;
	assign \g31019/_0_  = _w5941_ ;
	assign \g31020/_0_  = _w5947_ ;
	assign \g31021/_0_  = _w5950_ ;
	assign \g31022/_0_  = _w5954_ ;
	assign \g31023/_0_  = _w5957_ ;
	assign \g31024/_0_  = _w5961_ ;
	assign \g31025/_0_  = _w5965_ ;
	assign \g31026/_0_  = _w5969_ ;
	assign \g31027/_0_  = _w5973_ ;
	assign \g31028/_0_  = _w5977_ ;
	assign \g31029/_0_  = _w5981_ ;
	assign \g31030/_0_  = _w5985_ ;
	assign \g31031/_0_  = _w5989_ ;
	assign \g31032/_0_  = _w5993_ ;
	assign \g31033/_0_  = _w5997_ ;
	assign \g31034/_0_  = _w6001_ ;
	assign \g31035/_0_  = _w6005_ ;
	assign \g31036/_0_  = _w6010_ ;
	assign \g31037/_0_  = _w6013_ ;
	assign \g31038/_0_  = _w6016_ ;
	assign \g31039/_0_  = _w6019_ ;
	assign \g31040/_0_  = _w6022_ ;
	assign \g31041/_0_  = _w6025_ ;
	assign \g31042/_0_  = _w6028_ ;
	assign \g31043/_0_  = _w6031_ ;
	assign \g31044/_0_  = _w6035_ ;
	assign \g31045/_0_  = _w6038_ ;
	assign \g31046/_0_  = _w6041_ ;
	assign \g31047/_0_  = _w6044_ ;
	assign \g31048/_0_  = _w6047_ ;
	assign \g31049/_0_  = _w6050_ ;
	assign \g31050/_0_  = _w6053_ ;
	assign \g31051/_0_  = _w6056_ ;
	assign \g31052/_0_  = _w6059_ ;
	assign \g31053/_0_  = _w6062_ ;
	assign \g31054/_0_  = _w6065_ ;
	assign \g31055/_0_  = _w6068_ ;
	assign \g31056/_0_  = _w6071_ ;
	assign \g31057/_0_  = _w6074_ ;
	assign \g31058/_0_  = _w6077_ ;
	assign \g31059/_0_  = _w6080_ ;
	assign \g31060/_0_  = _w6083_ ;
	assign \g31061/_0_  = _w6086_ ;
	assign \g31062/_0_  = _w6089_ ;
	assign \g31063/_0_  = _w6092_ ;
	assign \g31064/_0_  = _w6095_ ;
	assign \g31065/_0_  = _w6098_ ;
	assign \g31066/_0_  = _w6101_ ;
	assign \g31067/_0_  = _w6104_ ;
	assign \g31068/_0_  = _w6107_ ;
	assign \g31069/_0_  = _w6110_ ;
	assign \g31070/_0_  = _w6113_ ;
	assign \g31071/_0_  = _w6116_ ;
	assign \g31072/_0_  = _w6119_ ;
	assign \g31073/_0_  = _w6122_ ;
	assign \g31074/_0_  = _w6125_ ;
	assign \g31075/_0_  = _w6128_ ;
	assign \g31076/_0_  = _w6131_ ;
	assign \g31077/_0_  = _w6134_ ;
	assign \g31084/u3_syn_4  = _w3068_ ;
	assign \g31085/u3_syn_4  = _w5668_ ;
	assign \g31096/u3_syn_4  = _w5733_ ;
	assign \g31115/u3_syn_4  = _w5801_ ;
	assign \g31136/u3_syn_4  = _w3315_ ;
	assign \g31158/u3_syn_4  = _w3505_ ;
	assign \g31176/u3_syn_4  = _w5951_ ;
	assign \g31193/u3_syn_4  = _w6032_ ;
	assign \g31195/u3_syn_4  = _w6007_ ;
	assign \g31247/u3_syn_4  = _w5699_ ;
	assign \g31280/u3_syn_4  = _w5929_ ;
	assign \g31285/u3_syn_4  = _w5934_ ;
	assign \g31568/_0_  = _w6138_ ;
	assign \g31631/_0_  = _w6175_ ;
	assign \g31672/_0_  = _w6182_ ;
	assign \g31731/_0_  = _w6186_ ;
	assign \g31732/_0_  = _w6190_ ;
	assign \g31742/_2_  = _w6192_ ;
	assign \g31744/_2_  = _w6194_ ;
	assign \g31746/_2_  = _w6196_ ;
	assign \g31748/_2_  = _w6198_ ;
	assign \g31751/_2_  = _w6200_ ;
	assign \g31754/_2_  = _w6202_ ;
	assign \g31756/_2_  = _w6204_ ;
	assign \g31758/_2_  = _w6206_ ;
	assign \g31760/_2_  = _w6208_ ;
	assign \g31761/_0_  = _w6210_ ;
	assign \g31789/_0_  = _w6213_ ;
	assign \g31807/_3_  = _w6218_ ;
	assign \g31825/_3_  = _w6221_ ;
	assign \g32607/_0_  = _w6234_ ;
	assign \g32608/_0_  = _w6247_ ;
	assign \g32609/_0_  = _w6260_ ;
	assign \g32610/_0_  = _w6273_ ;
	assign \g32611/_0_  = _w6286_ ;
	assign \g32612/_0_  = _w6299_ ;
	assign \g32613/_0_  = _w6305_ ;
	assign \g32614/_0_  = _w6311_ ;
	assign \g32615/_0_  = _w6317_ ;
	assign \g32616/_0_  = _w6323_ ;
	assign \g32617/_0_  = _w6329_ ;
	assign \g32618/_0_  = _w6335_ ;
	assign \g32645/_0__syn_2  = _w6336_ ;
	assign \g32687/_0__syn_2  = _w6337_ ;
	assign \g32749/_0__syn_2  = _w6338_ ;
	assign \g32757/_0_  = _w6346_ ;
	assign \g32758/_0_  = _w6353_ ;
	assign \g32759/_0_  = _w6360_ ;
	assign \g32760/_0_  = _w6367_ ;
	assign \g32761/_0_  = _w6374_ ;
	assign \g32762/_0_  = _w6381_ ;
	assign \g32763/_0_  = _w6388_ ;
	assign \g32764/_0_  = _w6395_ ;
	assign \g32765/_0_  = _w6402_ ;
	assign \g32769/_0_  = _w6406_ ;
	assign \g32835/_1_  = _w3313_ ;
	assign \g32839/_0_  = _w6410_ ;
	assign \g32844/_0_  = _w6414_ ;
	assign \g32901/_1_  = _w3503_ ;
	assign \g32902/_0_  = _w6418_ ;
	assign \g32963/_1_  = _w3066_ ;
	assign \g32972/_0_  = _w6422_ ;
	assign \g32977/_0_  = _w6426_ ;
	assign \g32979/_0_  = _w6429_ ;
	assign \g32980/_0_  = _w6432_ ;
	assign \g32981/_0_  = _w6435_ ;
	assign \g32982/_0_  = _w6438_ ;
	assign \g32983/_0_  = _w6441_ ;
	assign \g32987/_0_  = _w6444_ ;
	assign \g33018/_0_  = _w6446_ ;
	assign \g33019/_0_  = _w6450_ ;
	assign \g33088/_0_  = _w6453_ ;
	assign \g33261/_0_  = _w6460_ ;
	assign \g33264/_0_  = _w6462_ ;
	assign \g33275/_0_  = _w6463_ ;
	assign \g33276/_0_  = _w6467_ ;
	assign \g33277/_0_  = _w6468_ ;
	assign \g33371/_0_  = _w6478_ ;
	assign \g33382/_0_  = _w6484_ ;
	assign \g33401/_0_  = _w6488_ ;
	assign \g33402/_0_  = _w6492_ ;
	assign \g33403/_0_  = _w6495_ ;
	assign \g33404/_0_  = _w6498_ ;
	assign \g33405/_0_  = _w6501_ ;
	assign \g33406/_0_  = _w6504_ ;
	assign \g33407/_0_  = _w6507_ ;
	assign \g33408/_0_  = _w6510_ ;
	assign \g33409/_0_  = _w6513_ ;
	assign \g33410/_0_  = _w6516_ ;
	assign \g33411/_0_  = _w6519_ ;
	assign \g33412/_0_  = _w6522_ ;
	assign \g33413/_0_  = _w6525_ ;
	assign \g33414/_0_  = _w6528_ ;
	assign \g33415/_0_  = _w6531_ ;
	assign \g33416/_0_  = _w6534_ ;
	assign \g33417/_0_  = _w6537_ ;
	assign \g33418/_0_  = _w6540_ ;
	assign \g33419/_0_  = _w6543_ ;
	assign \g33420/_0_  = _w6546_ ;
	assign \g33421/_0_  = _w6549_ ;
	assign \g33422/_0_  = _w6552_ ;
	assign \g33423/_0_  = _w6555_ ;
	assign \g33424/_0_  = _w6558_ ;
	assign \g33425/_0_  = _w6561_ ;
	assign \g33426/_0_  = _w6564_ ;
	assign \g33427/_0_  = _w6567_ ;
	assign \g33428/_0_  = _w6570_ ;
	assign \g33429/_0_  = _w6573_ ;
	assign \g33430/_0_  = _w6576_ ;
	assign \g33431/_0_  = _w6579_ ;
	assign \g33432/_0_  = _w6582_ ;
	assign \g33433/_0_  = _w6586_ ;
	assign \g33434/_0_  = _w6589_ ;
	assign \g33435/_0_  = _w6592_ ;
	assign \g33436/_0_  = _w6595_ ;
	assign \g33437/_0_  = _w6598_ ;
	assign \g33438/_0_  = _w6601_ ;
	assign \g33439/_0_  = _w6604_ ;
	assign \g33440/_0_  = _w6607_ ;
	assign \g33441/_0_  = _w6610_ ;
	assign \g33442/_0_  = _w6613_ ;
	assign \g33443/_0_  = _w6616_ ;
	assign \g33444/_0_  = _w6619_ ;
	assign \g33445/_0_  = _w6622_ ;
	assign \g33446/_0_  = _w6625_ ;
	assign \g33447/_0_  = _w6628_ ;
	assign \g33448/_0_  = _w6632_ ;
	assign \g33449/_0_  = _w6635_ ;
	assign \g33450/_0_  = _w6638_ ;
	assign \g33451/_0_  = _w6641_ ;
	assign \g33452/_0_  = _w6644_ ;
	assign \g33453/_0_  = _w6647_ ;
	assign \g33454/_0_  = _w6650_ ;
	assign \g33455/_0_  = _w6653_ ;
	assign \g33456/_0_  = _w6656_ ;
	assign \g33457/_0_  = _w6659_ ;
	assign \g33458/_0_  = _w6662_ ;
	assign \g33459/_0_  = _w6665_ ;
	assign \g33460/_0_  = _w6668_ ;
	assign \g33461/_0_  = _w6671_ ;
	assign \g33462/_0_  = _w6674_ ;
	assign \g33463/_0_  = _w6677_ ;
	assign \g33464/_0_  = _w6680_ ;
	assign \g33465/_0_  = _w6683_ ;
	assign \g33466/_0_  = _w6686_ ;
	assign \g33467/_0_  = _w6689_ ;
	assign \g33468/_0_  = _w6692_ ;
	assign \g33469/_0_  = _w6695_ ;
	assign \g33470/_0_  = _w6698_ ;
	assign \g33471/_0_  = _w6701_ ;
	assign \g33472/_0_  = _w6704_ ;
	assign \g33473/_0_  = _w6707_ ;
	assign \g33474/_0_  = _w6710_ ;
	assign \g33475/_0_  = _w6713_ ;
	assign \g33476/_0_  = _w6716_ ;
	assign \g33477/_0_  = _w6719_ ;
	assign \g33478/_0_  = _w6722_ ;
	assign \g33479/_0_  = _w6725_ ;
	assign \g33480/_0_  = _w6728_ ;
	assign \g33481/_0_  = _w6731_ ;
	assign \g33482/_0_  = _w6734_ ;
	assign \g33483/_0_  = _w6737_ ;
	assign \g33484/_0_  = _w6740_ ;
	assign \g33485/_0_  = _w6743_ ;
	assign \g33486/_0_  = _w6746_ ;
	assign \g33487/_0_  = _w6749_ ;
	assign \g33488/_0_  = _w6752_ ;
	assign \g33489/_0_  = _w6755_ ;
	assign \g33490/_0_  = _w6758_ ;
	assign \g33491/_0_  = _w6761_ ;
	assign \g33492/_0_  = _w6764_ ;
	assign \g33493/_0_  = _w6767_ ;
	assign \g33494/_0_  = _w6770_ ;
	assign \g33495/_0_  = _w6773_ ;
	assign \g33496/_0_  = _w6776_ ;
	assign \g33497/_0_  = _w6779_ ;
	assign \g33498/_0_  = _w6782_ ;
	assign \g33499/_0_  = _w6785_ ;
	assign \g33500/_0_  = _w6788_ ;
	assign \g33501/_0_  = _w6791_ ;
	assign \g33502/_0_  = _w6794_ ;
	assign \g33503/_0_  = _w6797_ ;
	assign \g33504/_0_  = _w6800_ ;
	assign \g33505/_0_  = _w6803_ ;
	assign \g33506/_0_  = _w6806_ ;
	assign \g33507/_0_  = _w6810_ ;
	assign \g33508/_0_  = _w6813_ ;
	assign \g33509/_0_  = _w6816_ ;
	assign \g33510/_0_  = _w6819_ ;
	assign \g33511/_0_  = _w6822_ ;
	assign \g33512/_0_  = _w6825_ ;
	assign \g33513/_0_  = _w6828_ ;
	assign \g33514/_0_  = _w6831_ ;
	assign \g33515/_0_  = _w6834_ ;
	assign \g33516/_0_  = _w6837_ ;
	assign \g33517/_0_  = _w6840_ ;
	assign \g33518/_0_  = _w6843_ ;
	assign \g33519/_0_  = _w6846_ ;
	assign \g33520/_0_  = _w6849_ ;
	assign \g33521/_0_  = _w6852_ ;
	assign \g33522/_0_  = _w6855_ ;
	assign \g33523/_0_  = _w6858_ ;
	assign \g33524/_0_  = _w6861_ ;
	assign \g33525/_0_  = _w6864_ ;
	assign \g33526/_0_  = _w6867_ ;
	assign \g33527/_0_  = _w6870_ ;
	assign \g33528/_0_  = _w6873_ ;
	assign \g33529/_0_  = _w6876_ ;
	assign \g33530/_0_  = _w6879_ ;
	assign \g33531/_0_  = _w6882_ ;
	assign \g33532/_0_  = _w6885_ ;
	assign \g33533/_0_  = _w6888_ ;
	assign \g33534/_0_  = _w6891_ ;
	assign \g33535/_0_  = _w6894_ ;
	assign \g33536/_0_  = _w6897_ ;
	assign \g33537/_0_  = _w6900_ ;
	assign \g33538/_0_  = _w6903_ ;
	assign \g33539/_0_  = _w6907_ ;
	assign \g33540/_0_  = _w6910_ ;
	assign \g33541/_0_  = _w6913_ ;
	assign \g33542/_0_  = _w6916_ ;
	assign \g33543/_0_  = _w6919_ ;
	assign \g33544/_0_  = _w6922_ ;
	assign \g33545/_0_  = _w6925_ ;
	assign \g33546/_0_  = _w6928_ ;
	assign \g33547/_0_  = _w6931_ ;
	assign \g33548/_0_  = _w6934_ ;
	assign \g33549/_0_  = _w6937_ ;
	assign \g33550/_0_  = _w6940_ ;
	assign \g33551/_0_  = _w6943_ ;
	assign \g33552/_0_  = _w6946_ ;
	assign \g33553/_0_  = _w6949_ ;
	assign \g33554/_0_  = _w6952_ ;
	assign \g33555/_0_  = _w6955_ ;
	assign \g33556/_0_  = _w6958_ ;
	assign \g33557/_0_  = _w6961_ ;
	assign \g33558/_0_  = _w6964_ ;
	assign \g33559/_0_  = _w6967_ ;
	assign \g33560/_0_  = _w6970_ ;
	assign \g33561/_0_  = _w6973_ ;
	assign \g33562/_0_  = _w6976_ ;
	assign \g33563/_0_  = _w6979_ ;
	assign \g33564/_0_  = _w6982_ ;
	assign \g33565/_0_  = _w6985_ ;
	assign \g33566/_0_  = _w6988_ ;
	assign \g33567/_0_  = _w6991_ ;
	assign \g33568/_0_  = _w6994_ ;
	assign \g33569/_0_  = _w6997_ ;
	assign \g33570/_0_  = _w7000_ ;
	assign \g33571/_0_  = _w7003_ ;
	assign \g33572/_0_  = _w7006_ ;
	assign \g33573/_0_  = _w7009_ ;
	assign \g33574/_0_  = _w7012_ ;
	assign \g33575/_0_  = _w7015_ ;
	assign \g33576/_0_  = _w7018_ ;
	assign \g33577/_0_  = _w7021_ ;
	assign \g33578/_0_  = _w7024_ ;
	assign \g33579/_0_  = _w7027_ ;
	assign \g33580/_0_  = _w7030_ ;
	assign \g33581/_0_  = _w7033_ ;
	assign \g33582/_0_  = _w7036_ ;
	assign \g33583/_0_  = _w7039_ ;
	assign \g33584/_0_  = _w7042_ ;
	assign \g33585/_0_  = _w7045_ ;
	assign \g33586/_0_  = _w7048_ ;
	assign \g33587/_0_  = _w7051_ ;
	assign \g33588/_0_  = _w7054_ ;
	assign \g33589/_0_  = _w7057_ ;
	assign \g33590/_0_  = _w7060_ ;
	assign \g33591/_0_  = _w7063_ ;
	assign \g33592/_0_  = _w7066_ ;
	assign \g33593/_0_  = _w7069_ ;
	assign \g33594/_0_  = _w7072_ ;
	assign \g33595/_0_  = _w7075_ ;
	assign \g33596/_0_  = _w7078_ ;
	assign \g33597/_0_  = _w7081_ ;
	assign \g33598/_0_  = _w7084_ ;
	assign \g33599/_0_  = _w7087_ ;
	assign \g33600/_0_  = _w7090_ ;
	assign \g33601/_0_  = _w7093_ ;
	assign \g33602/_0_  = _w7096_ ;
	assign \g33603/_0_  = _w7099_ ;
	assign \g33604/_0_  = _w7103_ ;
	assign \g33605/_0_  = _w7106_ ;
	assign \g33606/_0_  = _w7109_ ;
	assign \g33607/_0_  = _w7112_ ;
	assign \g33608/_0_  = _w7115_ ;
	assign \g33609/_0_  = _w7118_ ;
	assign \g33610/_0_  = _w7121_ ;
	assign \g33611/_0_  = _w7124_ ;
	assign \g33612/_0_  = _w7127_ ;
	assign \g33613/_0_  = _w7130_ ;
	assign \g33614/_0_  = _w7133_ ;
	assign \g33615/_0_  = _w7136_ ;
	assign \g33616/_0_  = _w7139_ ;
	assign \g33617/_0_  = _w7142_ ;
	assign \g33618/_0_  = _w7145_ ;
	assign \g33619/_0_  = _w7148_ ;
	assign \g33620/_0_  = _w7151_ ;
	assign \g33621/_0_  = _w7154_ ;
	assign \g33622/_0_  = _w7157_ ;
	assign \g33623/_0_  = _w7160_ ;
	assign \g33624/_0_  = _w7163_ ;
	assign \g33625/_0_  = _w7166_ ;
	assign \g33626/_0_  = _w7169_ ;
	assign \g33627/_0_  = _w7172_ ;
	assign \g33628/_0_  = _w7175_ ;
	assign \g33629/_0_  = _w7178_ ;
	assign \g33630/_0_  = _w7181_ ;
	assign \g33631/_0_  = _w7184_ ;
	assign \g33632/_0_  = _w7187_ ;
	assign \g33633/_0_  = _w7190_ ;
	assign \g33634/_0_  = _w7193_ ;
	assign \g33635/_0_  = _w7196_ ;
	assign \g33636/_0_  = _w7200_ ;
	assign \g33637/_0_  = _w7203_ ;
	assign \g33638/_0_  = _w7206_ ;
	assign \g33639/_0_  = _w7209_ ;
	assign \g33640/_0_  = _w7212_ ;
	assign \g33641/_0_  = _w7215_ ;
	assign \g33642/_0_  = _w7218_ ;
	assign \g33643/_0_  = _w7221_ ;
	assign \g33644/_0_  = _w7224_ ;
	assign \g33645/_0_  = _w7227_ ;
	assign \g33646/_0_  = _w7230_ ;
	assign \g33647/_0_  = _w7233_ ;
	assign \g33648/_0_  = _w7236_ ;
	assign \g33649/_0_  = _w7239_ ;
	assign \g33650/_0_  = _w7242_ ;
	assign \g33651/_0_  = _w7245_ ;
	assign \g33652/_0_  = _w7248_ ;
	assign \g33653/_0_  = _w7251_ ;
	assign \g33654/_0_  = _w7254_ ;
	assign \g33655/_0_  = _w7257_ ;
	assign \g33656/_0_  = _w7260_ ;
	assign \g33657/_0_  = _w7263_ ;
	assign \g33658/_0_  = _w7266_ ;
	assign \g33659/_0_  = _w7269_ ;
	assign \g33660/_0_  = _w7272_ ;
	assign \g33661/_0_  = _w7275_ ;
	assign \g33662/_0_  = _w7278_ ;
	assign \g33663/_0_  = _w7281_ ;
	assign \g33664/_0_  = _w7284_ ;
	assign \g33665/_0_  = _w7287_ ;
	assign \g33666/_0_  = _w7290_ ;
	assign \g33667/_0_  = _w7293_ ;
	assign \g33668/_0_  = _w7296_ ;
	assign \g33669/_0_  = _w7299_ ;
	assign \g33670/_0_  = _w7302_ ;
	assign \g33671/_0_  = _w7305_ ;
	assign \g33672/_0_  = _w7308_ ;
	assign \g33673/_0_  = _w7311_ ;
	assign \g33674/_0_  = _w7314_ ;
	assign \g33675/_0_  = _w7317_ ;
	assign \g33676/_0_  = _w7320_ ;
	assign \g33677/_0_  = _w7323_ ;
	assign \g33678/_0_  = _w7326_ ;
	assign \g33679/_0_  = _w7329_ ;
	assign \g33680/_0_  = _w7332_ ;
	assign \g33681/_0_  = _w7335_ ;
	assign \g33682/_0_  = _w7338_ ;
	assign \g33683/_0_  = _w7341_ ;
	assign \g33684/_0_  = _w7344_ ;
	assign \g33685/_0_  = _w7347_ ;
	assign \g33686/_0_  = _w7350_ ;
	assign \g33687/_0_  = _w7353_ ;
	assign \g33688/_0_  = _w7356_ ;
	assign \g33689/_0_  = _w7359_ ;
	assign \g33690/_0_  = _w7362_ ;
	assign \g33691/_0_  = _w7365_ ;
	assign \g33692/_0_  = _w7368_ ;
	assign \g33693/_0_  = _w7371_ ;
	assign \g33694/_0_  = _w7374_ ;
	assign \g33695/_0_  = _w7377_ ;
	assign \g33696/_0_  = _w7380_ ;
	assign \g33697/_0_  = _w7383_ ;
	assign \g33698/_0_  = _w7386_ ;
	assign \g33699/_0_  = _w7389_ ;
	assign \g33700/_0_  = _w7392_ ;
	assign \g33701/_0_  = _w7395_ ;
	assign \g33702/_0_  = _w7398_ ;
	assign \g33703/_0_  = _w7401_ ;
	assign \g33704/_0_  = _w7405_ ;
	assign \g33705/_0_  = _w7408_ ;
	assign \g33706/_0_  = _w7411_ ;
	assign \g33707/_0_  = _w7414_ ;
	assign \g33708/_0_  = _w7417_ ;
	assign \g33709/_0_  = _w7420_ ;
	assign \g33710/_0_  = _w7423_ ;
	assign \g33711/_0_  = _w7426_ ;
	assign \g33712/_0_  = _w7429_ ;
	assign \g33713/_0_  = _w7432_ ;
	assign \g33714/_0_  = _w7435_ ;
	assign \g33715/_0_  = _w7438_ ;
	assign \g33716/_0_  = _w7441_ ;
	assign \g33717/_0_  = _w7444_ ;
	assign \g33718/_0_  = _w7447_ ;
	assign \g33719/_0_  = _w7450_ ;
	assign \g33720/_0_  = _w7453_ ;
	assign \g33721/_0_  = _w7456_ ;
	assign \g33722/_0_  = _w7459_ ;
	assign \g33723/_0_  = _w7462_ ;
	assign \g33724/_0_  = _w7465_ ;
	assign \g33725/_0_  = _w7468_ ;
	assign \g33726/_0_  = _w7471_ ;
	assign \g33727/_0_  = _w7474_ ;
	assign \g33728/_0_  = _w7477_ ;
	assign \g33729/_0_  = _w7480_ ;
	assign \g33730/_0_  = _w7483_ ;
	assign \g33731/_0_  = _w7486_ ;
	assign \g33732/_0_  = _w7489_ ;
	assign \g33733/_0_  = _w7492_ ;
	assign \g33734/_0_  = _w7495_ ;
	assign \g33735/_0_  = _w7498_ ;
	assign \g33736/_0_  = _w7502_ ;
	assign \g33737/_0_  = _w7505_ ;
	assign \g33738/_0_  = _w7508_ ;
	assign \g33739/_0_  = _w7511_ ;
	assign \g33740/_0_  = _w7514_ ;
	assign \g33741/_0_  = _w7517_ ;
	assign \g33742/_0_  = _w7520_ ;
	assign \g33743/_0_  = _w7523_ ;
	assign \g33744/_0_  = _w7526_ ;
	assign \g33745/_0_  = _w7529_ ;
	assign \g33746/_0_  = _w7532_ ;
	assign \g33747/_0_  = _w7535_ ;
	assign \g33748/_0_  = _w7538_ ;
	assign \g33749/_0_  = _w7541_ ;
	assign \g33750/_0_  = _w7544_ ;
	assign \g33751/_0_  = _w7547_ ;
	assign \g33752/_0_  = _w7550_ ;
	assign \g33753/_0_  = _w7553_ ;
	assign \g33754/_0_  = _w7556_ ;
	assign \g33755/_0_  = _w7559_ ;
	assign \g33756/_0_  = _w7562_ ;
	assign \g33757/_0_  = _w7565_ ;
	assign \g33758/_0_  = _w7568_ ;
	assign \g33759/_0_  = _w7571_ ;
	assign \g33760/_0_  = _w7574_ ;
	assign \g33761/_0_  = _w7577_ ;
	assign \g33762/_0_  = _w7580_ ;
	assign \g33763/_0_  = _w7583_ ;
	assign \g33764/_0_  = _w7586_ ;
	assign \g33765/_0_  = _w7589_ ;
	assign \g33766/_0_  = _w7592_ ;
	assign \g33767/_0_  = _w7595_ ;
	assign \g33768/_0_  = _w7598_ ;
	assign \g33769/_0_  = _w7601_ ;
	assign \g33770/_0_  = _w7604_ ;
	assign \g33771/_0_  = _w7607_ ;
	assign \g33772/_0_  = _w7610_ ;
	assign \g33773/_0_  = _w7613_ ;
	assign \g33774/_0_  = _w7616_ ;
	assign \g33775/_0_  = _w7619_ ;
	assign \g33776/_0_  = _w7622_ ;
	assign \g33777/_0_  = _w7625_ ;
	assign \g33778/_0_  = _w7628_ ;
	assign \g33779/_0_  = _w7631_ ;
	assign \g33780/_0_  = _w7634_ ;
	assign \g33781/_0_  = _w7637_ ;
	assign \g33782/_0_  = _w7640_ ;
	assign \g33783/_0_  = _w7643_ ;
	assign \g33784/_0_  = _w7646_ ;
	assign \g33785/_0_  = _w7649_ ;
	assign \g33786/_0_  = _w7652_ ;
	assign \g33787/_0_  = _w7655_ ;
	assign \g33788/_0_  = _w7658_ ;
	assign \g33789/_0_  = _w7661_ ;
	assign \g33790/_0_  = _w7664_ ;
	assign \g33791/_0_  = _w7667_ ;
	assign \g33792/_0_  = _w7670_ ;
	assign \g33793/_0_  = _w7673_ ;
	assign \g33794/_0_  = _w7676_ ;
	assign \g33795/_0_  = _w7679_ ;
	assign \g33796/_0_  = _w7682_ ;
	assign \g33797/_0_  = _w7685_ ;
	assign \g33798/_0_  = _w7688_ ;
	assign \g33799/_0_  = _w7691_ ;
	assign \g33800/_0_  = _w7694_ ;
	assign \g33801/_0_  = _w7697_ ;
	assign \g33802/_0_  = _w7700_ ;
	assign \g33803/_0_  = _w7703_ ;
	assign \g33804/_0_  = _w7706_ ;
	assign \g33805/_0_  = _w7709_ ;
	assign \g33806/_0_  = _w7713_ ;
	assign \g33807/_0_  = _w7716_ ;
	assign \g33808/_0_  = _w7719_ ;
	assign \g33809/_0_  = _w7722_ ;
	assign \g33810/_0_  = _w7725_ ;
	assign \g33811/_0_  = _w7728_ ;
	assign \g33812/_0_  = _w7731_ ;
	assign \g33813/_0_  = _w7734_ ;
	assign \g33814/_0_  = _w7737_ ;
	assign \g33815/_0_  = _w7740_ ;
	assign \g33816/_0_  = _w7743_ ;
	assign \g33817/_0_  = _w7746_ ;
	assign \g33818/_0_  = _w7749_ ;
	assign \g33819/_0_  = _w7752_ ;
	assign \g33820/_0_  = _w7755_ ;
	assign \g33821/_0_  = _w7758_ ;
	assign \g33822/_0_  = _w7761_ ;
	assign \g33823/_0_  = _w7764_ ;
	assign \g33824/_0_  = _w7767_ ;
	assign \g33825/_0_  = _w7770_ ;
	assign \g33826/_0_  = _w7773_ ;
	assign \g33827/_0_  = _w7776_ ;
	assign \g33828/_0_  = _w7779_ ;
	assign \g33829/_0_  = _w7782_ ;
	assign \g33830/_0_  = _w7785_ ;
	assign \g33831/_0_  = _w7788_ ;
	assign \g33832/_0_  = _w7791_ ;
	assign \g33833/_0_  = _w7794_ ;
	assign \g33834/_0_  = _w7797_ ;
	assign \g33835/_0_  = _w7800_ ;
	assign \g33836/_0_  = _w7803_ ;
	assign \g33837/_0_  = _w7806_ ;
	assign \g33838/_0_  = _w7809_ ;
	assign \g33839/_0_  = _w7812_ ;
	assign \g33840/_0_  = _w7816_ ;
	assign \g33841/_0_  = _w7819_ ;
	assign \g33842/_0_  = _w7822_ ;
	assign \g33843/_0_  = _w7825_ ;
	assign \g33844/_0_  = _w7828_ ;
	assign \g33845/_0_  = _w7831_ ;
	assign \g33846/_0_  = _w7834_ ;
	assign \g33847/_0_  = _w7837_ ;
	assign \g33848/_0_  = _w7840_ ;
	assign \g33849/_0_  = _w7843_ ;
	assign \g33850/_0_  = _w7846_ ;
	assign \g33851/_0_  = _w7849_ ;
	assign \g33852/_0_  = _w7852_ ;
	assign \g33853/_0_  = _w7855_ ;
	assign \g33854/_0_  = _w7858_ ;
	assign \g33855/_0_  = _w7861_ ;
	assign \g33856/_0_  = _w7864_ ;
	assign \g33857/_0_  = _w7867_ ;
	assign \g33858/_0_  = _w7870_ ;
	assign \g33859/_0_  = _w7873_ ;
	assign \g33860/_0_  = _w7876_ ;
	assign \g33861/_0_  = _w7879_ ;
	assign \g33862/_0_  = _w7882_ ;
	assign \g33863/_0_  = _w7885_ ;
	assign \g33864/_0_  = _w7888_ ;
	assign \g33865/_0_  = _w7891_ ;
	assign \g33866/_0_  = _w7894_ ;
	assign \g33867/_0_  = _w7897_ ;
	assign \g33868/_0_  = _w7900_ ;
	assign \g33869/_0_  = _w7903_ ;
	assign \g33870/_0_  = _w7906_ ;
	assign \g33871/_0_  = _w7909_ ;
	assign \g33872/_0_  = _w7912_ ;
	assign \g33873/_0_  = _w7915_ ;
	assign \g33874/_0_  = _w7918_ ;
	assign \g33875/_0_  = _w7921_ ;
	assign \g33876/_0_  = _w7924_ ;
	assign \g33877/_0_  = _w7927_ ;
	assign \g33878/_0_  = _w7930_ ;
	assign \g33879/_0_  = _w7933_ ;
	assign \g33880/_0_  = _w7936_ ;
	assign \g33881/_0_  = _w7939_ ;
	assign \g33882/_0_  = _w7942_ ;
	assign \g33883/_0_  = _w7945_ ;
	assign \g33884/_0_  = _w7948_ ;
	assign \g33885/_0_  = _w7951_ ;
	assign \g33886/_0_  = _w7954_ ;
	assign \g33887/_0_  = _w7957_ ;
	assign \g33888/_0_  = _w7960_ ;
	assign \g33889/_0_  = _w7963_ ;
	assign \g33890/_0_  = _w7966_ ;
	assign \g33891/_0_  = _w7969_ ;
	assign \g33892/_0_  = _w7972_ ;
	assign \g33893/_0_  = _w7975_ ;
	assign \g33894/_0_  = _w7978_ ;
	assign \g33895/_0_  = _w7981_ ;
	assign \g33896/_0_  = _w7984_ ;
	assign \g33897/_0_  = _w7987_ ;
	assign \g33898/_0_  = _w7990_ ;
	assign \g33899/_0_  = _w7993_ ;
	assign \g33900/_0_  = _w7996_ ;
	assign \g33901/_0_  = _w7999_ ;
	assign \g33902/_0_  = _w8002_ ;
	assign \g33903/_0_  = _w8005_ ;
	assign \g33904/_0_  = _w8008_ ;
	assign \g33905/_0_  = _w8011_ ;
	assign \g33906/_0_  = _w8014_ ;
	assign \g33907/_0_  = _w8017_ ;
	assign \g33908/_0_  = _w8020_ ;
	assign \g33909/_0_  = _w8023_ ;
	assign \g33910/_0_  = _w8026_ ;
	assign \g33911/_0_  = _w8029_ ;
	assign \g33912/_0_  = _w8032_ ;
	assign \g33913/_0_  = _w8035_ ;
	assign \g33914/_0_  = _w8038_ ;
	assign \g33915/_0_  = _w8041_ ;
	assign \g33916/_0_  = _w8044_ ;
	assign \g33917/_0_  = _w8047_ ;
	assign \g33918/_0_  = _w8050_ ;
	assign \g33919/_0_  = _w8053_ ;
	assign \g33920/_0_  = _w8056_ ;
	assign \g33921/_0_  = _w8059_ ;
	assign \g33922/_0_  = _w8062_ ;
	assign \g33923/_0_  = _w8065_ ;
	assign \g33924/_0_  = _w8068_ ;
	assign \g33925/_0_  = _w8071_ ;
	assign \g33926/_0_  = _w8074_ ;
	assign \g33927/_0_  = _w8077_ ;
	assign \g33928/_0_  = _w8080_ ;
	assign \g33929/_0_  = _w8083_ ;
	assign \g33930/_0_  = _w8086_ ;
	assign \g33931/_0_  = _w8089_ ;
	assign \g33932/_0_  = _w8092_ ;
	assign \g33933/_0_  = _w8095_ ;
	assign \g33934/_0_  = _w8098_ ;
	assign \g33935/_0_  = _w8101_ ;
	assign \g33936/_0_  = _w8104_ ;
	assign \g33937/_0_  = _w8107_ ;
	assign \g33938/_0_  = _w8110_ ;
	assign \g33939/_0_  = _w8113_ ;
	assign \g33940/_0_  = _w8116_ ;
	assign \g33941/_0_  = _w8119_ ;
	assign \g33942/_0_  = _w8122_ ;
	assign \g33943/_0_  = _w8125_ ;
	assign \g33944/_0_  = _w8128_ ;
	assign \g33945/_0_  = _w8131_ ;
	assign \g33946/_0_  = _w8134_ ;
	assign \g33947/_0_  = _w8137_ ;
	assign \g33948/_0_  = _w8140_ ;
	assign \g33949/_0_  = _w8143_ ;
	assign \g33950/_0_  = _w8146_ ;
	assign \g33951/_0_  = _w8149_ ;
	assign \g33952/_0_  = _w8152_ ;
	assign \g33953/_0_  = _w8155_ ;
	assign \g33954/_0_  = _w8158_ ;
	assign \g33955/_0_  = _w8161_ ;
	assign \g33956/_0_  = _w8164_ ;
	assign \g33957/_0_  = _w8167_ ;
	assign \g33958/_0_  = _w8170_ ;
	assign \g33959/_0_  = _w8173_ ;
	assign \g33960/_0_  = _w8176_ ;
	assign \g33961/_0_  = _w8179_ ;
	assign \g33962/_0_  = _w8182_ ;
	assign \g33963/_0_  = _w8185_ ;
	assign \g33964/_0_  = _w8188_ ;
	assign \g33965/_0_  = _w8191_ ;
	assign \g33966/_0_  = _w8194_ ;
	assign \g33967/_0_  = _w8197_ ;
	assign \g33968/_0_  = _w8200_ ;
	assign \g33969/_0_  = _w8203_ ;
	assign \g33970/_0_  = _w8206_ ;
	assign \g33971/_0_  = _w8209_ ;
	assign \g33972/_0_  = _w8212_ ;
	assign \g33973/_0_  = _w8215_ ;
	assign \g33974/_0_  = _w8218_ ;
	assign \g33975/_0_  = _w8221_ ;
	assign \g33976/_0_  = _w8224_ ;
	assign \g33977/u3_syn_4  = _w8225_ ;
	assign \g33981/u3_syn_4  = _w8226_ ;
	assign \g34014/u3_syn_4  = _w8227_ ;
	assign \g34047/u3_syn_4  = _w8228_ ;
	assign \g34084/u3_syn_4  = _w8229_ ;
	assign \g34123/u3_syn_4  = _w8230_ ;
	assign \g34306/_0_  = _w8248_ ;
	assign \g34316/_0_  = _w8266_ ;
	assign \g34324/_0_  = _w8284_ ;
	assign \g34326/_0_  = _w8302_ ;
	assign \g34328/_0_  = _w8320_ ;
	assign \g34331/_0_  = _w8338_ ;
	assign \g34333/_0_  = _w8356_ ;
	assign \g34344/_0_  = _w8374_ ;
	assign \g34347/_0_  = _w8392_ ;
	assign \g34351/_0_  = _w8410_ ;
	assign \g34361/_0_  = _w8428_ ;
	assign \g34368/_0_  = _w8446_ ;
	assign \g34377/_0_  = _w8464_ ;
	assign \g34385/_0_  = _w8482_ ;
	assign \g34393/_0_  = _w8500_ ;
	assign \g34414/_1_  = _w8501_ ;
	assign \g34451/_1_  = _w8502_ ;
	assign \g34476/_1_  = _w8503_ ;
	assign \g34487/_0_  = _w8504_ ;
	assign \g34490/_1_  = _w8505_ ;
	assign \g34715/_0_  = _w8508_ ;
	assign \g34878/_0_  = _w8520_ ;
	assign \g34882/_0_  = _w8532_ ;
	assign \g34883/_0_  = _w8534_ ;
	assign \g34893/_0_  = _w8546_ ;
	assign \g34896/_0_  = _w8561_ ;
	assign \g34898/_0_  = _w8576_ ;
	assign \g34899/_0_  = _w8588_ ;
	assign \g34916/_3_  = _w8591_ ;
	assign \g35264/_0_  = _w8596_ ;
	assign \g35265/_0_  = _w8601_ ;
	assign \g35266/_0_  = _w8606_ ;
	assign \g35267/_0_  = _w8610_ ;
	assign \g35268/_0_  = _w8614_ ;
	assign \g35269/_0_  = _w8618_ ;
	assign \g35270/_0_  = _w8621_ ;
	assign \g35271/_0_  = _w8624_ ;
	assign \g35272/_0_  = _w8640_ ;
	assign \g35273/_0_  = _w8656_ ;
	assign \g35274/_0_  = _w8672_ ;
	assign \g35275/_0_  = _w8675_ ;
	assign \g35276/_0_  = _w8691_ ;
	assign \g35277/_0_  = _w8707_ ;
	assign \g35278/_0_  = _w8723_ ;
	assign \g35279/_0_  = _w8737_ ;
	assign \g35283/_0_  = _w8740_ ;
	assign \g35287/_0_  = _w3062_ ;
	assign \g35294/_0_  = _w6339_ ;
	assign \g35300/_0_  = _w2758_ ;
	assign \g35304/_0_  = _w2769_ ;
	assign \g35308/_0_  = _w2794_ ;
	assign \g35312/_0_  = _w2807_ ;
	assign \g35316/_0_  = _w2158_ ;
	assign \g35318/_0_  = _w3309_ ;
	assign \g35326/_0_  = _w8756_ ;
	assign \g35334/_0_  = _w3499_ ;
	assign \g35336/_0_  = _w8760_ ;
	assign \g35337/_0_  = _w8764_ ;
	assign \g35338/_0_  = _w8767_ ;
	assign \g35357/_0_  = _w8769_ ;
	assign \g35358/_0_  = _w8771_ ;
	assign \g35359/_0_  = _w8773_ ;
	assign \g35419/_0_  = _w8776_ ;
	assign \g35438/_0_  = _w8781_ ;
	assign \g35439/_0_  = _w8782_ ;
	assign \g35440/_0_  = _w8783_ ;
	assign \g35441/_0_  = _w8784_ ;
	assign \g35442/_0_  = _w8785_ ;
	assign \g35444/_0_  = _w8797_ ;
	assign \g35445/_0_  = _w8809_ ;
	assign \g35446/_0_  = _w8821_ ;
	assign \g35447/_0_  = _w8833_ ;
	assign \g35448/_0_  = _w8845_ ;
	assign \g35449/_0_  = _w8852_ ;
	assign \g35450/_0_  = _w8859_ ;
	assign \g35451/_0_  = _w8868_ ;
	assign \g35452/_0_  = _w8871_ ;
	assign \g35463/_0_  = _w8874_ ;
	assign \g35464/_0_  = _w8931_ ;
	assign \g35466/_0_  = _w8932_ ;
	assign \g35485/_2_  = _w8935_ ;
	assign \g35495/_0_  = _w8937_ ;
	assign \g35496/_0_  = _w8939_ ;
	assign \g35499/_0_  = _w8941_ ;
	assign \g35500/_0_  = _w8943_ ;
	assign \g35501/_0_  = _w8945_ ;
	assign \g35502/_0_  = _w8947_ ;
	assign \g35563/_0_  = _w8948_ ;
	assign \g35633/_0_  = _w8949_ ;
	assign \g35717/_0_  = _w8956_ ;
	assign \g35718/_0_  = _w8963_ ;
	assign \g35719/_0_  = _w8970_ ;
	assign \g35809/_0_  = _w8972_ ;
	assign \g35810/_0_  = _w8974_ ;
	assign \g35811/_0_  = _w8976_ ;
	assign \g35812/_0_  = _w8978_ ;
	assign \g35813/_0_  = _w8980_ ;
	assign \g35814/_0_  = _w8982_ ;
	assign \g35815/_0_  = _w8984_ ;
	assign \g35816/_0_  = _w8986_ ;
	assign \g35817/_0_  = _w8988_ ;
	assign \g35818/_0_  = _w8990_ ;
	assign \g35819/_0_  = _w8992_ ;
	assign \g35820/_0_  = _w8994_ ;
	assign \g35821/_0_  = _w8996_ ;
	assign \g35822/_0_  = _w8998_ ;
	assign \g35823/_0_  = _w9000_ ;
	assign \g35824/_0_  = _w9002_ ;
	assign \g35825/_0_  = _w9004_ ;
	assign \g35826/_0_  = _w9006_ ;
	assign \g35827/_0_  = _w9008_ ;
	assign \g35830/_0_  = _w9016_ ;
	assign \g35833/_0_  = _w9020_ ;
	assign \g35835/_0_  = _w9027_ ;
	assign \g35836/_0_  = _w9035_ ;
	assign \g35837/_0_  = _w9043_ ;
	assign \g35839/_0_  = _w9047_ ;
	assign \g35840/_0_  = _w9050_ ;
	assign \g35841/_0_  = _w9057_ ;
	assign \g35843/_0_  = _w9059_ ;
	assign \g35844/_0_  = _w9066_ ;
	assign \g35845/_0_  = _w9070_ ;
	assign \g35853/_0_  = _w9071_ ;
	assign \g35854/_0_  = _w9072_ ;
	assign \g35855/_0_  = _w9076_ ;
	assign \g35856/_0_  = _w9077_ ;
	assign \g36306/_0_  = _w9082_ ;
	assign \g36414/_0_  = _w9083_ ;
	assign \g36415/_0_  = _w9084_ ;
	assign \g36449/_0_  = _w9088_ ;
	assign \g36550/_0_  = _w9089_ ;
	assign \g36551/_0_  = _w9092_ ;
	assign \g36553/_0_  = _w9095_ ;
	assign \g36560/_0_  = _w9097_ ;
	assign \g36562/_3_  = _w9099_ ;
	assign \g36563/_0_  = _w9103_ ;
	assign \g36612/_0_  = _w9104_ ;
	assign \g36614/_2_  = _w9108_ ;
	assign \g36695/_0_  = _w9111_ ;
	assign \g36784/_0_  = _w9122_ ;
	assign \g36785/_0_  = _w9129_ ;
	assign \g36786/_0_  = _w9136_ ;
	assign \g36787/_0_  = _w9143_ ;
	assign \g36788/_0_  = _w9150_ ;
	assign \g36789/_0_  = _w9157_ ;
	assign \g36790/_0_  = _w9164_ ;
	assign \g36791/_0_  = _w9171_ ;
	assign \g36792/_0_  = _w9178_ ;
	assign \g36793/_0_  = _w9185_ ;
	assign \g36794/_0_  = _w9192_ ;
	assign \g36796/_0_  = _w9199_ ;
	assign \g36797/_0_  = _w9206_ ;
	assign \g36798/_0_  = _w9213_ ;
	assign \g36799/_0_  = _w9220_ ;
	assign \g36800/_0_  = _w9227_ ;
	assign \g36801/_0_  = _w9234_ ;
	assign \g36802/_0_  = _w9241_ ;
	assign \g36803/_0_  = _w9248_ ;
	assign \g36804/_0_  = _w9255_ ;
	assign \g36805/_0_  = _w9262_ ;
	assign \g36806/_0_  = _w9269_ ;
	assign \g36807/_0_  = _w9276_ ;
	assign \g36808/_0_  = _w9283_ ;
	assign \g36809/_0_  = _w9290_ ;
	assign \g36810/_0_  = _w9297_ ;
	assign \g36811/_0_  = _w9304_ ;
	assign \g36813/_0_  = _w9311_ ;
	assign \g36814/_0_  = _w9322_ ;
	assign \g36815/_0_  = _w9329_ ;
	assign \g36820/_0_  = _w9336_ ;
	assign \g36825/_0_  = _w9343_ ;
	assign \g36832/_0_  = _w9350_ ;
	assign \g36846/_0_  = _w9357_ ;
	assign \g36855/_0_  = _w9364_ ;
	assign \g36857/_0_  = _w9371_ ;
	assign \g36859/_0_  = _w9378_ ;
	assign \g36860/_0_  = _w9385_ ;
	assign \g36861/_0_  = _w9392_ ;
	assign \g36862/_0_  = _w9403_ ;
	assign \g36863/_0_  = _w9410_ ;
	assign \g36864/_0_  = _w9417_ ;
	assign \g36867/_0_  = _w9424_ ;
	assign \g36870/_0_  = _w9431_ ;
	assign \g36871/_0_  = _w9438_ ;
	assign \g36877/_0_  = _w9445_ ;
	assign \g36879/_0_  = _w9452_ ;
	assign \g36892/_0_  = _w9459_ ;
	assign \g36893/_0_  = _w9466_ ;
	assign \g36901/_0_  = _w9473_ ;
	assign \g36909/_0_  = _w9480_ ;
	assign \g36914/_0_  = _w9487_ ;
	assign \g36919/_0_  = _w9494_ ;
	assign \g36922/_0_  = _w9501_ ;
	assign \g36923/_0_  = _w9508_ ;
	assign \g36927/_0_  = _w9515_ ;
	assign \g36930/_0_  = _w9522_ ;
	assign \g36931/_0_  = _w9529_ ;
	assign \g36933/_0_  = _w9536_ ;
	assign \g36934/_0_  = _w9543_ ;
	assign \g36935/_0_  = _w9550_ ;
	assign \g36936/_0_  = _w9557_ ;
	assign \g36937/_0_  = _w9564_ ;
	assign \g36938/_0_  = _w9571_ ;
	assign \g36939/_0_  = _w9578_ ;
	assign \g36940/_0_  = _w9585_ ;
	assign \g36941/_0_  = _w9592_ ;
	assign \g36943/_0_  = _w9599_ ;
	assign \g36944/_0_  = _w9606_ ;
	assign \g36945/_0_  = _w9613_ ;
	assign \g36946/_0_  = _w9620_ ;
	assign \g36947/_0_  = _w9627_ ;
	assign \g36948/_0_  = _w9634_ ;
	assign \g36949/_0_  = _w9641_ ;
	assign \g36950/_0_  = _w9648_ ;
	assign \g36951/_0_  = _w9655_ ;
	assign \g36952/_0_  = _w9662_ ;
	assign \g36953/_0_  = _w9669_ ;
	assign \g36954/_0_  = _w9676_ ;
	assign \g36957/_0_  = _w9683_ ;
	assign \g36958/_0_  = _w9690_ ;
	assign \g36959/_0_  = _w9697_ ;
	assign \g36960/_0_  = _w9704_ ;
	assign \g36961/_0_  = _w9711_ ;
	assign \g36962/_0_  = _w9718_ ;
	assign \g36963/_0_  = _w9725_ ;
	assign \g36970/_0_  = _w9732_ ;
	assign \g36977/_0_  = _w9739_ ;
	assign \g36986/_0_  = _w9746_ ;
	assign \g36991/_0_  = _w9753_ ;
	assign \g36994/_0_  = _w9760_ ;
	assign \g37015/_0_  = _w9767_ ;
	assign \g37057/_0_  = _w9774_ ;
	assign \g37073/_0_  = _w9781_ ;
	assign \g37128/_0_  = _w9788_ ;
	assign \g37129/_0_  = _w9795_ ;
	assign \g37138/_0_  = _w9801_ ;
	assign \g37139/_0_  = _w9802_ ;
	assign \g37140/_0_  = _w9808_ ;
	assign \g37141/_0_  = _w9813_ ;
	assign \g37142/_0_  = _w9818_ ;
	assign \g37143/_0_  = _w9823_ ;
	assign \g37144/_0_  = _w9828_ ;
	assign \g37145/_0_  = _w9833_ ;
	assign \g37146/_0_  = _w9838_ ;
	assign \g37147/_0_  = _w9843_ ;
	assign \g37148/_0_  = _w9848_ ;
	assign \g37149/_0_  = _w9853_ ;
	assign \g37150/_0_  = _w9858_ ;
	assign \g37151/_0_  = _w9863_ ;
	assign \g37152/_0_  = _w9868_ ;
	assign \g37153/_0_  = _w9874_ ;
	assign \g37154/_0_  = _w9879_ ;
	assign \g37155/_0_  = _w9884_ ;
	assign \g37156/_0_  = _w9889_ ;
	assign \g37157/_0_  = _w9894_ ;
	assign \g37158/_0_  = _w9899_ ;
	assign \g37159/_0_  = _w9904_ ;
	assign \g37160/_0_  = _w9909_ ;
	assign \g37161/_0_  = _w9914_ ;
	assign \g37162/_0_  = _w9919_ ;
	assign \g37163/_0_  = _w9924_ ;
	assign \g37164/_0_  = _w9929_ ;
	assign \g37165/_0_  = _w9934_ ;
	assign \g37166/_0_  = _w9939_ ;
	assign \g37167/_0_  = _w9944_ ;
	assign \g37168/_0_  = _w9949_ ;
	assign \g37169/_0_  = _w9954_ ;
	assign \g37170/_0_  = _w9959_ ;
	assign \g37171/_0_  = _w9964_ ;
	assign \g37172/_0_  = _w9969_ ;
	assign \g37173/_0_  = _w9974_ ;
	assign \g37174/_0_  = _w9979_ ;
	assign \g37175/_0_  = _w9984_ ;
	assign \g37176/_0_  = _w9989_ ;
	assign \g37177/_0_  = _w9994_ ;
	assign \g37178/_0_  = _w9999_ ;
	assign \g37179/_0_  = _w10004_ ;
	assign \g37180/_0_  = _w10009_ ;
	assign \g37181/_0_  = _w10014_ ;
	assign \g37182/_0_  = _w10019_ ;
	assign \g37183/_0_  = _w10024_ ;
	assign \g37184/_0_  = _w10029_ ;
	assign \g37185/_0_  = _w10034_ ;
	assign \g37187/_0_  = _w10039_ ;
	assign \g37188/_0_  = _w10044_ ;
	assign \g37190/_0_  = _w10049_ ;
	assign \g37191/_0_  = _w10054_ ;
	assign \g37192/_0_  = _w10059_ ;
	assign \g37193/_0_  = _w10064_ ;
	assign \g37194/_0_  = _w10069_ ;
	assign \g37372/_3_  = _w10072_ ;
	assign \g37377/_0_  = _w10075_ ;
	assign \g37378/_0_  = _w10078_ ;
	assign \g37379/_0_  = _w10081_ ;
	assign \g37380/_0_  = _w10084_ ;
	assign \g37381/_0_  = _w10087_ ;
	assign \g37382/_0_  = _w10090_ ;
	assign \g37383/_0_  = _w10093_ ;
	assign \g37384/_0_  = _w10096_ ;
	assign \g37385/_0_  = _w10099_ ;
	assign \g37386/_0_  = _w10102_ ;
	assign \g37387/_0_  = _w10105_ ;
	assign \g37388/_0_  = _w10108_ ;
	assign \g37389/_0_  = _w10111_ ;
	assign \g37390/_0_  = _w10114_ ;
	assign \g37391/_0_  = _w10117_ ;
	assign \g37392/_0_  = _w10120_ ;
	assign \g37393/_0_  = _w10123_ ;
	assign \g37394/_0_  = _w10126_ ;
	assign \g37395/_0_  = _w10129_ ;
	assign \g37396/_0_  = _w10132_ ;
	assign \g37397/_0_  = _w10135_ ;
	assign \g37398/_0_  = _w10138_ ;
	assign \g37399/_0_  = _w10141_ ;
	assign \g37400/_0_  = _w10144_ ;
	assign \g37401/_0_  = _w10147_ ;
	assign \g37402/_0_  = _w10150_ ;
	assign \g37403/_0_  = _w10153_ ;
	assign \g37404/_0_  = _w10156_ ;
	assign \g37405/_0_  = _w10159_ ;
	assign \g37406/_0_  = _w10162_ ;
	assign \g37407/_0_  = _w10165_ ;
	assign \g37408/_0_  = _w10168_ ;
	assign \g37409/_0_  = _w10171_ ;
	assign \g37410/_0_  = _w10174_ ;
	assign \g37411/_0_  = _w10177_ ;
	assign \g37412/_0_  = _w10180_ ;
	assign \g37413/_0_  = _w10183_ ;
	assign \g37576/_3_  = _w9064_ ;
	assign \g37590/_2_  = _w2738_ ;
	assign \g40278/_0_  = _w8778_ ;
	assign \g40379/_0_  = _w8521_ ;
	assign \g40389/_2_  = _w9013_ ;
	assign \g40390/_2_  = _w9032_ ;
	assign \g40391/_0_  = _w6289_ ;
	assign \g40393/_2_  = _w9040_ ;
	assign \g40395/_0_  = _w8551_ ;
	assign \g40397/_0_  = _w8509_ ;
	assign \g40400/_0_  = _w6263_ ;
	assign \g40402/_0_  = _w8566_ ;
	assign \g45458/_0_  = _w2155_ ;
	assign \g45675/_0_  = _w10188_ ;
	assign \g45677/_0_  = _w10186_ ;
	assign \g45678/_0_  = _w10193_ ;
	assign \g45682/_0_  = _w10191_ ;
	assign sync_pad_o_pad = _w10194_ ;
	assign \u14_u0_full_empty_r_reg/P0001_reg_syn_3  = _w10197_ ;
	assign \u14_u1_full_empty_r_reg/P0001_reg_syn_3  = _w10200_ ;
	assign \u14_u2_full_empty_r_reg/P0001_reg_syn_3  = _w10203_ ;
	assign \u14_u3_full_empty_r_reg/P0001_reg_syn_3  = _w10206_ ;
	assign \u14_u4_full_empty_r_reg/P0001_reg_syn_3  = _w10209_ ;
	assign \u14_u5_full_empty_r_reg/P0001_reg_syn_3  = _w10212_ ;
	assign \u14_u6_full_empty_r_reg/P0001_reg_syn_3  = _w10215_ ;
	assign \u14_u7_full_empty_r_reg/P0001_reg_syn_3  = _w10218_ ;
	assign \u14_u8_full_empty_r_reg/P0001_reg_syn_3  = _w10221_ ;
	assign \u1_slt0_reg[11]/P0001_reg_syn_3  = _w10224_ ;
	assign \u1_slt0_reg[12]/P0001_reg_syn_3  = _w10227_ ;
	assign \u1_slt0_reg[15]/P0001_reg_syn_3  = _w10230_ ;
	assign \u1_slt0_reg[9]/P0001_reg_syn_3  = _w10233_ ;
	assign \u1_slt1_reg[10]/P0001_reg_syn_3  = _w10236_ ;
	assign \u1_slt1_reg[11]/P0001_reg_syn_3  = _w10239_ ;
	assign \u1_slt1_reg[5]/P0001_reg_syn_3  = _w10242_ ;
	assign \u1_slt1_reg[6]/P0001_reg_syn_3  = _w10245_ ;
	assign \u1_slt1_reg[7]/P0001_reg_syn_3  = _w10248_ ;
	assign \u1_slt1_reg[8]/P0001_reg_syn_3  = _w10251_ ;
	assign wb_err_o_pad = 1'b0;
endmodule;