module top( \EN_DISP_reg/NET0131  , \FLAG_reg/NET0131  , \MAR_reg[0]/NET0131  , \MAR_reg[1]/NET0131  , \MAR_reg[2]/NET0131  , \MAR_reg[3]/NET0131  , \MAR_reg[4]/NET0131  , \MAX_reg[0]/NET0131  , \MAX_reg[1]/NET0131  , \MAX_reg[2]/NET0131  , \MAX_reg[3]/NET0131  , \MAX_reg[4]/NET0131  , \MAX_reg[5]/NET0131  , \MAX_reg[6]/NET0131  , \MAX_reg[7]/NET0131  , \MAX_reg[8]/NET0131  , \NUM_reg[0]/NET0131  , \NUM_reg[1]/NET0131  , \NUM_reg[2]/NET0131  , \NUM_reg[3]/NET0131  , \NUM_reg[4]/NET0131  , \RES_DISP_reg/NET0131  , START_pad , \STATO_reg[0]/NET0131  , \STATO_reg[1]/NET0131  , \STATO_reg[2]/NET0131  , \TEMP_reg[0]/NET0131  , \TEMP_reg[1]/NET0131  , \TEMP_reg[2]/NET0131  , \TEMP_reg[3]/NET0131  , \TEMP_reg[4]/NET0131  , \TEMP_reg[5]/NET0131  , \TEMP_reg[6]/NET0131  , \TEMP_reg[7]/NET0131  , \TEMP_reg[8]/NET0131  , \DISPMAX2[0]_pad  , \DISPMAX2[1]_pad  , \DISPMAX2[2]_pad  , \DISPMAX2[4]_pad  , \DISPMAX2[5]_pad  , \DISPMAX2[6]_pad  , \DISPMAX3[0]_pad  , \DISPMAX3[1]_pad  , \DISPMAX3[2]_pad  , \DISPMAX3[3]_pad  , \DISPMAX3[4]_pad  , \DISPMAX3[5]_pad  , \DISPMAX3[6]_pad  , \DISPNUM1[0]_pad  , \DISPNUM1[6]_pad  , \DISPNUM2[0]_pad  , \DISPNUM2[1]_pad  , \DISPNUM2[2]_pad  , \DISPNUM2[3]_pad  , \DISPNUM2[4]_pad  , \DISPNUM2[5]_pad  , \DISPNUM2[6]_pad  , SIGN_pad , \_al_n0  , \_al_n1  , \g2955/_2_  , \g2956/_2_  , \g2957/_2_  , \g2958/_2_  , \g2959/_2_  , \g2960/_2_  , \g2961/_2_  , \g2962/_2_  , \g2963/_2_  , \g2985/_0_  , \g3032/_0_  , \g3033/_0_  , \g3034/_0_  , \g3038/_0_  , \g3247/_0_  , \g3279/_0_  , \g3309/_0_  , \g3335/_0_  , \g3336/_0_  , \g3337/_0_  , \g3338/_0_  , \g3339/_0_  , \g3340/_0_  , \g3341/_0_  , \g3360/_0_  , \g3361/_0_  , \g3369/_0_  , \g3373/_0_  , \g3382/_0_  , \g3451/_0_  , \g3475/_0_  , \g3490/_0_  , \g3514/_0_  , \g3774/_1_  , \g4511/_0_  );
  input \EN_DISP_reg/NET0131  ;
  input \FLAG_reg/NET0131  ;
  input \MAR_reg[0]/NET0131  ;
  input \MAR_reg[1]/NET0131  ;
  input \MAR_reg[2]/NET0131  ;
  input \MAR_reg[3]/NET0131  ;
  input \MAR_reg[4]/NET0131  ;
  input \MAX_reg[0]/NET0131  ;
  input \MAX_reg[1]/NET0131  ;
  input \MAX_reg[2]/NET0131  ;
  input \MAX_reg[3]/NET0131  ;
  input \MAX_reg[4]/NET0131  ;
  input \MAX_reg[5]/NET0131  ;
  input \MAX_reg[6]/NET0131  ;
  input \MAX_reg[7]/NET0131  ;
  input \MAX_reg[8]/NET0131  ;
  input \NUM_reg[0]/NET0131  ;
  input \NUM_reg[1]/NET0131  ;
  input \NUM_reg[2]/NET0131  ;
  input \NUM_reg[3]/NET0131  ;
  input \NUM_reg[4]/NET0131  ;
  input \RES_DISP_reg/NET0131  ;
  input START_pad ;
  input \STATO_reg[0]/NET0131  ;
  input \STATO_reg[1]/NET0131  ;
  input \STATO_reg[2]/NET0131  ;
  input \TEMP_reg[0]/NET0131  ;
  input \TEMP_reg[1]/NET0131  ;
  input \TEMP_reg[2]/NET0131  ;
  input \TEMP_reg[3]/NET0131  ;
  input \TEMP_reg[4]/NET0131  ;
  input \TEMP_reg[5]/NET0131  ;
  input \TEMP_reg[6]/NET0131  ;
  input \TEMP_reg[7]/NET0131  ;
  input \TEMP_reg[8]/NET0131  ;
  output \DISPMAX2[0]_pad  ;
  output \DISPMAX2[1]_pad  ;
  output \DISPMAX2[2]_pad  ;
  output \DISPMAX2[4]_pad  ;
  output \DISPMAX2[5]_pad  ;
  output \DISPMAX2[6]_pad  ;
  output \DISPMAX3[0]_pad  ;
  output \DISPMAX3[1]_pad  ;
  output \DISPMAX3[2]_pad  ;
  output \DISPMAX3[3]_pad  ;
  output \DISPMAX3[4]_pad  ;
  output \DISPMAX3[5]_pad  ;
  output \DISPMAX3[6]_pad  ;
  output \DISPNUM1[0]_pad  ;
  output \DISPNUM1[6]_pad  ;
  output \DISPNUM2[0]_pad  ;
  output \DISPNUM2[1]_pad  ;
  output \DISPNUM2[2]_pad  ;
  output \DISPNUM2[3]_pad  ;
  output \DISPNUM2[4]_pad  ;
  output \DISPNUM2[5]_pad  ;
  output \DISPNUM2[6]_pad  ;
  output SIGN_pad ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g2955/_2_  ;
  output \g2956/_2_  ;
  output \g2957/_2_  ;
  output \g2958/_2_  ;
  output \g2959/_2_  ;
  output \g2960/_2_  ;
  output \g2961/_2_  ;
  output \g2962/_2_  ;
  output \g2963/_2_  ;
  output \g2985/_0_  ;
  output \g3032/_0_  ;
  output \g3033/_0_  ;
  output \g3034/_0_  ;
  output \g3038/_0_  ;
  output \g3247/_0_  ;
  output \g3279/_0_  ;
  output \g3309/_0_  ;
  output \g3335/_0_  ;
  output \g3336/_0_  ;
  output \g3337/_0_  ;
  output \g3338/_0_  ;
  output \g3339/_0_  ;
  output \g3340/_0_  ;
  output \g3341/_0_  ;
  output \g3360/_0_  ;
  output \g3361/_0_  ;
  output \g3369/_0_  ;
  output \g3373/_0_  ;
  output \g3382/_0_  ;
  output \g3451/_0_  ;
  output \g3475/_0_  ;
  output \g3490/_0_  ;
  output \g3514/_0_  ;
  output \g3774/_1_  ;
  output \g4511/_0_  ;
  wire n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 ;
  assign n36 = \MAX_reg[4]/NET0131  & ~\MAX_reg[8]/NET0131  ;
  assign n37 = ~\MAX_reg[0]/NET0131  & ~\MAX_reg[1]/NET0131  ;
  assign n38 = \MAX_reg[8]/NET0131  & ~n37 ;
  assign n39 = \MAX_reg[0]/NET0131  & \MAX_reg[1]/NET0131  ;
  assign n40 = n38 & ~n39 ;
  assign n41 = \MAX_reg[1]/NET0131  & ~\MAX_reg[8]/NET0131  ;
  assign n42 = ~n40 & ~n41 ;
  assign n43 = \MAX_reg[2]/NET0131  & ~n38 ;
  assign n44 = ~\MAX_reg[2]/NET0131  & n38 ;
  assign n45 = ~n43 & ~n44 ;
  assign n46 = \MAX_reg[3]/NET0131  & ~\MAX_reg[8]/NET0131  ;
  assign n47 = ~\MAX_reg[2]/NET0131  & n37 ;
  assign n49 = \MAX_reg[3]/NET0131  & ~n47 ;
  assign n48 = ~\MAX_reg[3]/NET0131  & n47 ;
  assign n50 = \MAX_reg[8]/NET0131  & ~n48 ;
  assign n51 = ~n49 & n50 ;
  assign n52 = ~n46 & ~n51 ;
  assign n53 = ~n45 & ~n52 ;
  assign n54 = ~n42 & n53 ;
  assign n55 = n36 & n54 ;
  assign n56 = ~\MAX_reg[4]/NET0131  & n48 ;
  assign n57 = \MAX_reg[8]/NET0131  & ~n56 ;
  assign n58 = n42 & n45 ;
  assign n59 = ~n57 & ~n58 ;
  assign n60 = ~n52 & n59 ;
  assign n61 = ~n36 & ~n60 ;
  assign n62 = ~n55 & ~n61 ;
  assign n63 = ~\EN_DISP_reg/NET0131  & \RES_DISP_reg/NET0131  ;
  assign n64 = ~n62 & n63 ;
  assign n65 = n61 & n63 ;
  assign n66 = n45 & n52 ;
  assign n67 = n36 & ~n66 ;
  assign n68 = ~n61 & ~n67 ;
  assign n69 = ~n55 & n63 ;
  assign n70 = ~n68 & n69 ;
  assign n71 = ~n54 & n67 ;
  assign n72 = n63 & ~n71 ;
  assign n73 = ~n55 & n68 ;
  assign n74 = n63 & ~n73 ;
  assign n75 = \RES_DISP_reg/NET0131  & ~n67 ;
  assign n76 = ~n55 & n75 ;
  assign n77 = ~\EN_DISP_reg/NET0131  & ~n76 ;
  assign n89 = ~n53 & n67 ;
  assign n90 = n36 & ~n58 ;
  assign n91 = ~n52 & ~n59 ;
  assign n92 = ~n90 & ~n91 ;
  assign n93 = ~n55 & ~n92 ;
  assign n94 = ~n89 & n93 ;
  assign n95 = ~\MAX_reg[0]/NET0131  & ~n94 ;
  assign n78 = n42 & ~n61 ;
  assign n79 = ~n67 & ~n78 ;
  assign n80 = n45 & n79 ;
  assign n81 = ~n45 & ~n79 ;
  assign n82 = ~n80 & ~n81 ;
  assign n96 = ~n82 & ~n94 ;
  assign n97 = ~n95 & ~n96 ;
  assign n83 = ~\MAX_reg[0]/NET0131  & ~n82 ;
  assign n85 = n42 & ~n68 ;
  assign n84 = ~n42 & n68 ;
  assign n86 = ~n55 & ~n84 ;
  assign n87 = ~n85 & n86 ;
  assign n98 = ~n83 & n87 ;
  assign n99 = ~n97 & n98 ;
  assign n88 = n83 & ~n87 ;
  assign n100 = ~n57 & ~n88 ;
  assign n101 = ~n99 & n100 ;
  assign n102 = n63 & ~n101 ;
  assign n103 = ~n57 & n94 ;
  assign n104 = ~n57 & ~n82 ;
  assign n105 = ~n87 & n95 ;
  assign n106 = n104 & ~n105 ;
  assign n107 = ~n87 & ~n94 ;
  assign n108 = ~n57 & ~n107 ;
  assign n109 = n97 & n108 ;
  assign n110 = ~n106 & ~n109 ;
  assign n111 = ~n103 & ~n110 ;
  assign n112 = n63 & ~n111 ;
  assign n113 = ~n57 & ~n109 ;
  assign n114 = ~n57 & ~n96 ;
  assign n115 = ~n105 & n114 ;
  assign n116 = ~n83 & ~n94 ;
  assign n117 = ~n115 & n116 ;
  assign n118 = n113 & n117 ;
  assign n119 = n63 & ~n118 ;
  assign n120 = ~n103 & ~n109 ;
  assign n121 = n115 & n120 ;
  assign n122 = n63 & ~n121 ;
  assign n123 = n87 & n95 ;
  assign n124 = n104 & n123 ;
  assign n125 = n63 & ~n124 ;
  assign n126 = n104 & n107 ;
  assign n127 = \MAX_reg[0]/NET0131  & n126 ;
  assign n128 = ~n114 & ~n127 ;
  assign n129 = ~n115 & ~n128 ;
  assign n130 = ~n109 & ~n129 ;
  assign n131 = ~n103 & ~n130 ;
  assign n132 = n63 & ~n131 ;
  assign n133 = n113 & ~n126 ;
  assign n134 = \RES_DISP_reg/NET0131  & ~n103 ;
  assign n135 = ~n133 & n134 ;
  assign n136 = ~\EN_DISP_reg/NET0131  & ~n135 ;
  assign n137 = ~\NUM_reg[1]/NET0131  & ~\NUM_reg[2]/NET0131  ;
  assign n138 = \NUM_reg[3]/NET0131  & ~n137 ;
  assign n139 = ~\NUM_reg[4]/NET0131  & ~n138 ;
  assign n140 = n63 & n139 ;
  assign n141 = ~\EN_DISP_reg/NET0131  & ~\RES_DISP_reg/NET0131  ;
  assign n142 = \NUM_reg[4]/NET0131  & ~n137 ;
  assign n143 = \NUM_reg[3]/NET0131  & n137 ;
  assign n144 = ~n142 & ~n143 ;
  assign n145 = ~\NUM_reg[1]/NET0131  & ~n139 ;
  assign n146 = \NUM_reg[1]/NET0131  & n139 ;
  assign n147 = ~n145 & ~n146 ;
  assign n152 = \NUM_reg[2]/NET0131  & ~n145 ;
  assign n153 = \NUM_reg[4]/NET0131  & n137 ;
  assign n154 = ~n152 & ~n153 ;
  assign n155 = ~n147 & ~n154 ;
  assign n156 = n144 & ~n155 ;
  assign n157 = ~\NUM_reg[0]/NET0131  & n144 ;
  assign n158 = ~n156 & ~n157 ;
  assign n159 = n144 & n154 ;
  assign n148 = ~\NUM_reg[2]/NET0131  & n147 ;
  assign n160 = \NUM_reg[0]/NET0131  & n148 ;
  assign n161 = n159 & ~n160 ;
  assign n162 = ~\NUM_reg[0]/NET0131  & ~n148 ;
  assign n163 = n161 & ~n162 ;
  assign n164 = ~n155 & ~n163 ;
  assign n165 = ~n158 & ~n164 ;
  assign n166 = n144 & ~n165 ;
  assign n149 = ~\NUM_reg[0]/NET0131  & n148 ;
  assign n150 = ~n138 & n149 ;
  assign n151 = ~n144 & ~n150 ;
  assign n167 = n63 & ~n151 ;
  assign n168 = ~n166 & n167 ;
  assign n169 = ~n149 & n154 ;
  assign n170 = ~n158 & ~n169 ;
  assign n171 = n144 & ~n170 ;
  assign n172 = n63 & ~n171 ;
  assign n173 = n147 & n157 ;
  assign n174 = ~n159 & ~n173 ;
  assign n175 = n156 & ~n174 ;
  assign n176 = ~\NUM_reg[0]/NET0131  & n159 ;
  assign n177 = n175 & ~n176 ;
  assign n178 = n63 & ~n177 ;
  assign n179 = ~n158 & n174 ;
  assign n180 = n63 & ~n179 ;
  assign n181 = ~n147 & n176 ;
  assign n182 = n63 & ~n181 ;
  assign n183 = ~n161 & n175 ;
  assign n184 = ~n158 & ~n183 ;
  assign n185 = n144 & ~n184 ;
  assign n186 = n63 & ~n185 ;
  assign n187 = ~n148 & ~n158 ;
  assign n188 = \RES_DISP_reg/NET0131  & n144 ;
  assign n189 = ~n187 & n188 ;
  assign n190 = ~\EN_DISP_reg/NET0131  & ~n189 ;
  assign n191 = ~\MAX_reg[8]/NET0131  & \RES_DISP_reg/NET0131  ;
  assign n192 = ~\EN_DISP_reg/NET0131  & ~n191 ;
  assign n204 = \MAR_reg[0]/NET0131  & ~\MAR_reg[2]/NET0131  ;
  assign n205 = \MAR_reg[3]/NET0131  & n204 ;
  assign n193 = ~\MAR_reg[1]/NET0131  & ~\MAR_reg[2]/NET0131  ;
  assign n194 = \MAR_reg[4]/NET0131  & n193 ;
  assign n202 = ~\MAR_reg[1]/NET0131  & \MAR_reg[2]/NET0131  ;
  assign n203 = ~\MAR_reg[3]/NET0131  & n202 ;
  assign n206 = ~n194 & ~n203 ;
  assign n207 = ~n205 & n206 ;
  assign n195 = \MAR_reg[2]/NET0131  & ~\MAR_reg[3]/NET0131  ;
  assign n196 = ~\MAR_reg[3]/NET0131  & \MAR_reg[4]/NET0131  ;
  assign n197 = ~n195 & ~n196 ;
  assign n198 = ~\MAR_reg[0]/NET0131  & ~n197 ;
  assign n199 = \MAR_reg[1]/NET0131  & ~\MAR_reg[4]/NET0131  ;
  assign n200 = \MAR_reg[0]/NET0131  & ~n195 ;
  assign n201 = n199 & n200 ;
  assign n208 = ~n198 & ~n201 ;
  assign n209 = n207 & n208 ;
  assign n210 = \TEMP_reg[6]/NET0131  & n209 ;
  assign n215 = ~\MAR_reg[3]/NET0131  & ~\MAR_reg[4]/NET0131  ;
  assign n216 = \MAR_reg[2]/NET0131  & n215 ;
  assign n217 = ~\MAR_reg[1]/NET0131  & n196 ;
  assign n218 = ~n216 & ~n217 ;
  assign n219 = ~\MAR_reg[0]/NET0131  & ~n218 ;
  assign n211 = ~\MAR_reg[2]/NET0131  & \MAR_reg[4]/NET0131  ;
  assign n212 = ~n199 & ~n211 ;
  assign n213 = \MAR_reg[0]/NET0131  & ~n212 ;
  assign n214 = ~\MAR_reg[2]/NET0131  & n196 ;
  assign n220 = \MAR_reg[3]/NET0131  & ~\MAR_reg[4]/NET0131  ;
  assign n221 = ~\MAR_reg[2]/NET0131  & n220 ;
  assign n222 = ~n214 & ~n221 ;
  assign n223 = ~n213 & n222 ;
  assign n224 = ~n219 & n223 ;
  assign n225 = \TEMP_reg[7]/NET0131  & n224 ;
  assign n226 = ~n210 & ~n225 ;
  assign n239 = ~n214 & ~n216 ;
  assign n254 = ~n199 & ~n221 ;
  assign n255 = n239 & n254 ;
  assign n256 = \MAR_reg[0]/NET0131  & ~n255 ;
  assign n257 = \MAR_reg[1]/NET0131  & ~n239 ;
  assign n258 = \MAR_reg[3]/NET0131  & \MAR_reg[4]/NET0131  ;
  assign n259 = n193 & n258 ;
  assign n260 = \MAR_reg[4]/NET0131  & n195 ;
  assign n261 = ~n259 & ~n260 ;
  assign n262 = ~\MAR_reg[0]/NET0131  & ~n261 ;
  assign n263 = ~n257 & ~n262 ;
  assign n264 = ~n256 & n263 ;
  assign n265 = \TEMP_reg[0]/NET0131  & n264 ;
  assign n266 = ~n193 & ~n221 ;
  assign n267 = ~\MAR_reg[0]/NET0131  & ~n266 ;
  assign n227 = \MAR_reg[1]/NET0131  & \MAR_reg[2]/NET0131  ;
  assign n228 = \MAR_reg[3]/NET0131  & n227 ;
  assign n270 = ~n228 & ~n259 ;
  assign n240 = \MAR_reg[0]/NET0131  & \MAR_reg[1]/NET0131  ;
  assign n268 = \MAR_reg[4]/NET0131  & n240 ;
  assign n269 = n202 & n215 ;
  assign n271 = ~n268 & ~n269 ;
  assign n272 = n270 & n271 ;
  assign n273 = ~n267 & n272 ;
  assign n274 = \TEMP_reg[1]/NET0131  & n273 ;
  assign n275 = ~n265 & ~n274 ;
  assign n276 = ~\TEMP_reg[1]/NET0131  & ~n273 ;
  assign n277 = ~n275 & ~n276 ;
  assign n278 = n196 & ~n227 ;
  assign n279 = \MAR_reg[0]/NET0131  & ~\MAR_reg[1]/NET0131  ;
  assign n280 = ~n221 & n279 ;
  assign n281 = ~n196 & ~n280 ;
  assign n282 = ~n278 & ~n281 ;
  assign n283 = ~n194 & ~n221 ;
  assign n284 = ~\MAR_reg[0]/NET0131  & ~n283 ;
  assign n285 = \MAR_reg[4]/NET0131  & n205 ;
  assign n286 = ~n284 & ~n285 ;
  assign n287 = ~n282 & n286 ;
  assign n288 = \TEMP_reg[3]/NET0131  & n287 ;
  assign n290 = \MAR_reg[0]/NET0131  & ~n283 ;
  assign n291 = ~\MAR_reg[0]/NET0131  & n195 ;
  assign n289 = n215 & n240 ;
  assign n292 = ~n278 & ~n289 ;
  assign n293 = ~n291 & n292 ;
  assign n294 = ~n290 & n293 ;
  assign n295 = \TEMP_reg[2]/NET0131  & n294 ;
  assign n296 = ~n288 & ~n295 ;
  assign n297 = ~n277 & n296 ;
  assign n298 = ~\TEMP_reg[3]/NET0131  & ~n287 ;
  assign n299 = ~\TEMP_reg[2]/NET0131  & ~n294 ;
  assign n300 = ~n288 & n299 ;
  assign n301 = ~n298 & ~n300 ;
  assign n302 = ~n297 & n301 ;
  assign n231 = \MAR_reg[0]/NET0131  & ~n194 ;
  assign n232 = n197 & n231 ;
  assign n233 = ~n217 & ~n221 ;
  assign n234 = ~n228 & n233 ;
  assign n229 = ~n193 & ~n227 ;
  assign n230 = ~\MAR_reg[4]/NET0131  & ~n229 ;
  assign n235 = ~n198 & ~n230 ;
  assign n236 = n234 & n235 ;
  assign n237 = ~n232 & n236 ;
  assign n238 = \TEMP_reg[5]/NET0131  & n237 ;
  assign n242 = ~n215 & ~n227 ;
  assign n243 = ~n199 & ~n242 ;
  assign n244 = ~n202 & n220 ;
  assign n245 = ~n243 & ~n244 ;
  assign n246 = ~\MAR_reg[0]/NET0131  & ~n245 ;
  assign n241 = ~n239 & n240 ;
  assign n247 = \MAR_reg[2]/NET0131  & ~\MAR_reg[4]/NET0131  ;
  assign n248 = \MAR_reg[1]/NET0131  & \MAR_reg[3]/NET0131  ;
  assign n249 = ~n211 & n248 ;
  assign n250 = ~n247 & n249 ;
  assign n251 = ~n241 & ~n250 ;
  assign n252 = ~n246 & n251 ;
  assign n253 = \TEMP_reg[4]/NET0131  & n252 ;
  assign n303 = ~n238 & ~n253 ;
  assign n304 = ~n302 & n303 ;
  assign n305 = n226 & n304 ;
  assign n306 = ~\TEMP_reg[7]/NET0131  & ~n224 ;
  assign n307 = ~\TEMP_reg[6]/NET0131  & ~n209 ;
  assign n308 = ~\TEMP_reg[5]/NET0131  & ~n237 ;
  assign n309 = ~\TEMP_reg[4]/NET0131  & ~n252 ;
  assign n310 = ~n308 & ~n309 ;
  assign n311 = ~n238 & ~n310 ;
  assign n312 = ~n307 & ~n311 ;
  assign n313 = n226 & ~n312 ;
  assign n314 = ~n306 & ~n313 ;
  assign n315 = ~n305 & n314 ;
  assign n316 = ~\MAR_reg[0]/NET0131  & ~\MAR_reg[1]/NET0131  ;
  assign n317 = ~n239 & n316 ;
  assign n318 = n220 & n240 ;
  assign n319 = ~n285 & ~n318 ;
  assign n320 = ~n317 & n319 ;
  assign n321 = \TEMP_reg[8]/NET0131  & ~n320 ;
  assign n322 = ~\TEMP_reg[8]/NET0131  & n320 ;
  assign n323 = ~n321 & ~n322 ;
  assign n324 = n315 & n323 ;
  assign n325 = ~n315 & ~n323 ;
  assign n326 = ~n324 & ~n325 ;
  assign n327 = ~n210 & ~n307 ;
  assign n328 = ~n304 & ~n311 ;
  assign n329 = n327 & ~n328 ;
  assign n330 = ~n327 & n328 ;
  assign n331 = ~n329 & ~n330 ;
  assign n332 = ~\TEMP_reg[0]/NET0131  & ~n264 ;
  assign n371 = ~n276 & ~n332 ;
  assign n372 = n275 & n371 ;
  assign n373 = ~n331 & n372 ;
  assign n333 = ~n225 & ~n306 ;
  assign n334 = n277 & ~n299 ;
  assign n335 = ~n253 & n296 ;
  assign n336 = ~n334 & n335 ;
  assign n337 = ~n253 & n298 ;
  assign n338 = ~n309 & ~n337 ;
  assign n339 = ~n308 & n338 ;
  assign n340 = ~n336 & n339 ;
  assign n341 = ~n210 & ~n238 ;
  assign n342 = ~n340 & n341 ;
  assign n343 = ~n307 & ~n342 ;
  assign n344 = ~n333 & ~n343 ;
  assign n345 = n333 & n343 ;
  assign n374 = ~n344 & ~n345 ;
  assign n375 = n373 & n374 ;
  assign n346 = ~n265 & ~n332 ;
  assign n347 = ~n288 & ~n298 ;
  assign n348 = ~n295 & ~n334 ;
  assign n349 = n347 & ~n348 ;
  assign n351 = ~n295 & ~n299 ;
  assign n352 = ~n277 & ~n351 ;
  assign n353 = n277 & n351 ;
  assign n357 = ~n352 & ~n353 ;
  assign n358 = ~n349 & n357 ;
  assign n354 = ~n253 & ~n309 ;
  assign n356 = n302 & n354 ;
  assign n350 = ~n347 & n348 ;
  assign n355 = ~n302 & ~n354 ;
  assign n359 = ~n350 & ~n355 ;
  assign n360 = ~n356 & n359 ;
  assign n361 = n358 & n360 ;
  assign n362 = n346 & ~n361 ;
  assign n363 = ~n238 & ~n308 ;
  assign n364 = ~n336 & n338 ;
  assign n365 = n346 & ~n364 ;
  assign n366 = ~n346 & n364 ;
  assign n367 = ~n365 & ~n366 ;
  assign n368 = n363 & ~n367 ;
  assign n369 = ~n363 & n367 ;
  assign n370 = ~n368 & ~n369 ;
  assign n376 = ~n362 & ~n370 ;
  assign n377 = n375 & n376 ;
  assign n378 = ~n326 & ~n377 ;
  assign n382 = \MAX_reg[7]/NET0131  & n224 ;
  assign n391 = ~\MAX_reg[1]/NET0131  & ~n273 ;
  assign n392 = \MAX_reg[0]/NET0131  & n264 ;
  assign n393 = ~n391 & n392 ;
  assign n389 = \MAX_reg[2]/NET0131  & n294 ;
  assign n390 = \MAX_reg[1]/NET0131  & n273 ;
  assign n394 = ~n389 & ~n390 ;
  assign n395 = ~n393 & n394 ;
  assign n387 = ~\MAX_reg[3]/NET0131  & ~n287 ;
  assign n388 = ~\MAX_reg[2]/NET0131  & ~n294 ;
  assign n396 = ~n387 & ~n388 ;
  assign n397 = ~n395 & n396 ;
  assign n385 = \MAX_reg[3]/NET0131  & n287 ;
  assign n386 = \MAX_reg[4]/NET0131  & n252 ;
  assign n398 = ~n385 & ~n386 ;
  assign n399 = ~n397 & n398 ;
  assign n383 = ~\MAX_reg[4]/NET0131  & ~n252 ;
  assign n384 = ~\MAX_reg[5]/NET0131  & ~n237 ;
  assign n400 = ~n383 & ~n384 ;
  assign n401 = ~n399 & n400 ;
  assign n402 = \MAX_reg[6]/NET0131  & n209 ;
  assign n403 = \MAX_reg[5]/NET0131  & n237 ;
  assign n404 = ~n402 & ~n403 ;
  assign n405 = ~n401 & n404 ;
  assign n406 = ~\MAX_reg[7]/NET0131  & ~n224 ;
  assign n407 = ~\MAX_reg[6]/NET0131  & ~n209 ;
  assign n408 = ~n406 & ~n407 ;
  assign n409 = ~n405 & n408 ;
  assign n410 = ~n382 & ~n409 ;
  assign n411 = \MAX_reg[8]/NET0131  & ~n320 ;
  assign n412 = ~\MAX_reg[8]/NET0131  & n320 ;
  assign n413 = ~n411 & ~n412 ;
  assign n414 = n410 & n413 ;
  assign n415 = ~n410 & ~n413 ;
  assign n416 = ~n414 & ~n415 ;
  assign n417 = \MAX_reg[0]/NET0131  & n416 ;
  assign n418 = ~n264 & ~n416 ;
  assign n419 = ~n417 & ~n418 ;
  assign n420 = n378 & n419 ;
  assign n379 = ~\MAX_reg[0]/NET0131  & ~n378 ;
  assign n380 = \STATO_reg[1]/NET0131  & ~\STATO_reg[2]/NET0131  ;
  assign n381 = \STATO_reg[0]/NET0131  & n380 ;
  assign n421 = ~n379 & n381 ;
  assign n422 = ~n420 & n421 ;
  assign n423 = ~\STATO_reg[0]/NET0131  & ~\STATO_reg[1]/NET0131  ;
  assign n424 = \STATO_reg[2]/NET0131  & n423 ;
  assign n425 = ~\STATO_reg[1]/NET0131  & ~\STATO_reg[2]/NET0131  ;
  assign n426 = ~n424 & ~n425 ;
  assign n427 = \MAX_reg[0]/NET0131  & ~n426 ;
  assign n428 = ~\STATO_reg[0]/NET0131  & n380 ;
  assign n429 = ~n264 & n428 ;
  assign n430 = ~n427 & ~n429 ;
  assign n431 = ~n422 & n430 ;
  assign n433 = \MAX_reg[1]/NET0131  & n416 ;
  assign n434 = ~n273 & ~n416 ;
  assign n435 = ~n433 & ~n434 ;
  assign n436 = n378 & n435 ;
  assign n432 = ~\MAX_reg[1]/NET0131  & ~n378 ;
  assign n437 = n381 & ~n432 ;
  assign n438 = ~n436 & n437 ;
  assign n439 = \MAX_reg[1]/NET0131  & ~n426 ;
  assign n440 = ~n273 & n428 ;
  assign n441 = ~n439 & ~n440 ;
  assign n442 = ~n438 & n441 ;
  assign n444 = \MAX_reg[2]/NET0131  & n416 ;
  assign n445 = ~n294 & ~n416 ;
  assign n446 = ~n444 & ~n445 ;
  assign n447 = n378 & n446 ;
  assign n443 = ~\MAX_reg[2]/NET0131  & ~n378 ;
  assign n448 = n381 & ~n443 ;
  assign n449 = ~n447 & n448 ;
  assign n450 = \MAX_reg[2]/NET0131  & ~n426 ;
  assign n451 = ~n294 & n428 ;
  assign n452 = ~n450 & ~n451 ;
  assign n453 = ~n449 & n452 ;
  assign n455 = \MAX_reg[3]/NET0131  & n416 ;
  assign n456 = ~n287 & ~n416 ;
  assign n457 = ~n455 & ~n456 ;
  assign n458 = n378 & n457 ;
  assign n454 = ~\MAX_reg[3]/NET0131  & ~n378 ;
  assign n459 = n381 & ~n454 ;
  assign n460 = ~n458 & n459 ;
  assign n461 = \MAX_reg[3]/NET0131  & ~n426 ;
  assign n462 = ~n287 & n428 ;
  assign n463 = ~n461 & ~n462 ;
  assign n464 = ~n460 & n463 ;
  assign n466 = \MAX_reg[4]/NET0131  & n416 ;
  assign n467 = ~n252 & ~n416 ;
  assign n468 = ~n466 & ~n467 ;
  assign n469 = n378 & n468 ;
  assign n465 = ~\MAX_reg[4]/NET0131  & ~n378 ;
  assign n470 = n381 & ~n465 ;
  assign n471 = ~n469 & n470 ;
  assign n472 = \MAX_reg[4]/NET0131  & ~n426 ;
  assign n473 = ~n252 & n428 ;
  assign n474 = ~n472 & ~n473 ;
  assign n475 = ~n471 & n474 ;
  assign n477 = \MAX_reg[5]/NET0131  & n416 ;
  assign n478 = ~n237 & ~n416 ;
  assign n479 = ~n477 & ~n478 ;
  assign n480 = n378 & n479 ;
  assign n476 = ~\MAX_reg[5]/NET0131  & ~n378 ;
  assign n481 = n381 & ~n476 ;
  assign n482 = ~n480 & n481 ;
  assign n483 = \MAX_reg[5]/NET0131  & ~n426 ;
  assign n484 = ~n237 & n428 ;
  assign n485 = ~n483 & ~n484 ;
  assign n486 = ~n482 & n485 ;
  assign n488 = \MAX_reg[6]/NET0131  & n416 ;
  assign n489 = ~n209 & ~n416 ;
  assign n490 = ~n488 & ~n489 ;
  assign n491 = n378 & n490 ;
  assign n487 = ~\MAX_reg[6]/NET0131  & ~n378 ;
  assign n492 = n381 & ~n487 ;
  assign n493 = ~n491 & n492 ;
  assign n494 = \MAX_reg[6]/NET0131  & ~n426 ;
  assign n495 = ~n209 & n428 ;
  assign n496 = ~n494 & ~n495 ;
  assign n497 = ~n493 & n496 ;
  assign n499 = \MAX_reg[7]/NET0131  & n416 ;
  assign n500 = ~n224 & ~n416 ;
  assign n501 = ~n499 & ~n500 ;
  assign n502 = n378 & n501 ;
  assign n498 = ~\MAX_reg[7]/NET0131  & ~n378 ;
  assign n503 = n381 & ~n498 ;
  assign n504 = ~n502 & n503 ;
  assign n505 = \MAX_reg[7]/NET0131  & ~n426 ;
  assign n506 = ~n224 & n428 ;
  assign n507 = ~n505 & ~n506 ;
  assign n508 = ~n504 & n507 ;
  assign n513 = ~\MAX_reg[8]/NET0131  & ~n378 ;
  assign n509 = ~\MAX_reg[8]/NET0131  & ~n410 ;
  assign n510 = n320 & n410 ;
  assign n511 = ~n509 & ~n510 ;
  assign n512 = n378 & ~n511 ;
  assign n514 = n381 & ~n512 ;
  assign n515 = ~n513 & n514 ;
  assign n516 = \MAX_reg[8]/NET0131  & ~n426 ;
  assign n517 = ~n320 & n428 ;
  assign n518 = ~n516 & ~n517 ;
  assign n519 = ~n515 & n518 ;
  assign n520 = \STATO_reg[0]/NET0131  & n425 ;
  assign n521 = ~START_pad & n520 ;
  assign n522 = ~n428 & ~n521 ;
  assign n523 = ~n423 & n522 ;
  assign n524 = \FLAG_reg/NET0131  & ~n523 ;
  assign n525 = ~\FLAG_reg/NET0131  & ~n378 ;
  assign n526 = ~n326 & n381 ;
  assign n527 = ~n525 & n526 ;
  assign n528 = ~n524 & ~n527 ;
  assign n529 = \FLAG_reg/NET0131  & n326 ;
  assign n530 = \NUM_reg[0]/NET0131  & n529 ;
  assign n531 = n381 & ~n530 ;
  assign n532 = n523 & ~n531 ;
  assign n533 = \NUM_reg[1]/NET0131  & ~n532 ;
  assign n534 = ~\NUM_reg[1]/NET0131  & n381 ;
  assign n535 = n530 & n534 ;
  assign n536 = ~n533 & ~n535 ;
  assign n537 = \NUM_reg[2]/NET0131  & ~n523 ;
  assign n538 = \NUM_reg[0]/NET0131  & \NUM_reg[1]/NET0131  ;
  assign n541 = n529 & n538 ;
  assign n542 = ~\NUM_reg[2]/NET0131  & ~n541 ;
  assign n539 = \NUM_reg[2]/NET0131  & n538 ;
  assign n540 = n529 & n539 ;
  assign n543 = n381 & ~n540 ;
  assign n544 = ~n542 & n543 ;
  assign n545 = ~n537 & ~n544 ;
  assign n546 = \NUM_reg[3]/NET0131  & n540 ;
  assign n547 = n381 & ~n546 ;
  assign n548 = n523 & ~n547 ;
  assign n549 = \NUM_reg[4]/NET0131  & ~n548 ;
  assign n550 = ~\NUM_reg[4]/NET0131  & n381 ;
  assign n551 = n546 & n550 ;
  assign n552 = ~n549 & ~n551 ;
  assign n553 = \NUM_reg[3]/NET0131  & ~n548 ;
  assign n554 = n540 & n547 ;
  assign n555 = ~n553 & ~n554 ;
  assign n556 = ~n381 & n523 ;
  assign n557 = \MAR_reg[4]/NET0131  & ~n556 ;
  assign n558 = \MAR_reg[2]/NET0131  & n240 ;
  assign n559 = \MAR_reg[3]/NET0131  & n424 ;
  assign n560 = n558 & n559 ;
  assign n561 = ~n557 & ~n560 ;
  assign n562 = \TEMP_reg[5]/NET0131  & ~n426 ;
  assign n563 = ~n237 & n380 ;
  assign n564 = ~n562 & ~n563 ;
  assign n565 = ~\STATO_reg[2]/NET0131  & n423 ;
  assign n566 = n522 & ~n565 ;
  assign n567 = ~n381 & n566 ;
  assign n568 = \MAR_reg[3]/NET0131  & ~n567 ;
  assign n570 = \MAR_reg[2]/NET0131  & n318 ;
  assign n569 = ~\MAR_reg[3]/NET0131  & ~n558 ;
  assign n571 = n424 & ~n569 ;
  assign n572 = ~n570 & n571 ;
  assign n573 = ~n568 & ~n572 ;
  assign n574 = \TEMP_reg[0]/NET0131  & ~n426 ;
  assign n575 = ~n264 & n380 ;
  assign n576 = ~n574 & ~n575 ;
  assign n577 = \TEMP_reg[8]/NET0131  & ~n426 ;
  assign n578 = ~n320 & n380 ;
  assign n579 = ~n577 & ~n578 ;
  assign n580 = \TEMP_reg[1]/NET0131  & ~n426 ;
  assign n581 = ~n273 & n380 ;
  assign n582 = ~n580 & ~n581 ;
  assign n583 = \TEMP_reg[2]/NET0131  & ~n426 ;
  assign n584 = ~n294 & n380 ;
  assign n585 = ~n583 & ~n584 ;
  assign n586 = \TEMP_reg[3]/NET0131  & ~n426 ;
  assign n587 = ~n287 & n380 ;
  assign n588 = ~n586 & ~n587 ;
  assign n589 = \TEMP_reg[4]/NET0131  & ~n426 ;
  assign n590 = ~n252 & n380 ;
  assign n591 = ~n589 & ~n590 ;
  assign n592 = \TEMP_reg[6]/NET0131  & ~n426 ;
  assign n593 = ~n209 & n380 ;
  assign n594 = ~n592 & ~n593 ;
  assign n595 = ~n240 & ~n316 ;
  assign n596 = n258 & n558 ;
  assign n597 = ~n595 & ~n596 ;
  assign n598 = n424 & ~n597 ;
  assign n599 = \MAR_reg[1]/NET0131  & ~n567 ;
  assign n600 = ~n598 & ~n599 ;
  assign n601 = START_pad & n520 ;
  assign n602 = n424 & ~n596 ;
  assign n603 = ~n380 & ~n520 ;
  assign n604 = ~n602 & n603 ;
  assign n605 = \EN_DISP_reg/NET0131  & ~n604 ;
  assign n606 = ~n601 & ~n605 ;
  assign n607 = ~n258 & n558 ;
  assign n608 = ~\MAR_reg[2]/NET0131  & ~n240 ;
  assign n609 = n424 & ~n608 ;
  assign n610 = ~n607 & n609 ;
  assign n611 = \MAR_reg[2]/NET0131  & ~n567 ;
  assign n612 = ~n610 & ~n611 ;
  assign n613 = \MAR_reg[0]/NET0131  & ~n596 ;
  assign n614 = n424 & ~n613 ;
  assign n615 = \MAR_reg[0]/NET0131  & ~n567 ;
  assign n616 = ~n614 & ~n615 ;
  assign n617 = \TEMP_reg[7]/NET0131  & ~n426 ;
  assign n618 = ~n224 & n380 ;
  assign n619 = ~n617 & ~n618 ;
  assign n620 = START_pad & n596 ;
  assign n621 = n424 & n620 ;
  assign n622 = ~n381 & ~n621 ;
  assign n623 = n424 & ~n620 ;
  assign n624 = n566 & ~n623 ;
  assign n625 = ~n424 & n603 ;
  assign n626 = ~\RES_DISP_reg/NET0131  & ~n601 ;
  assign n627 = ~n625 & ~n626 ;
  assign n628 = ~n428 & ~n601 ;
  assign n629 = ~n602 & n628 ;
  assign n630 = \NUM_reg[0]/NET0131  & ~n532 ;
  assign n631 = n529 & n531 ;
  assign n632 = ~n630 & ~n631 ;
  assign \DISPMAX2[0]_pad  = n64 ;
  assign \DISPMAX2[1]_pad  = n65 ;
  assign \DISPMAX2[2]_pad  = n70 ;
  assign \DISPMAX2[4]_pad  = n72 ;
  assign \DISPMAX2[5]_pad  = n74 ;
  assign \DISPMAX2[6]_pad  = n77 ;
  assign \DISPMAX3[0]_pad  = n102 ;
  assign \DISPMAX3[1]_pad  = n112 ;
  assign \DISPMAX3[2]_pad  = n119 ;
  assign \DISPMAX3[3]_pad  = n122 ;
  assign \DISPMAX3[4]_pad  = n125 ;
  assign \DISPMAX3[5]_pad  = n132 ;
  assign \DISPMAX3[6]_pad  = n136 ;
  assign \DISPNUM1[0]_pad  = n140 ;
  assign \DISPNUM1[6]_pad  = n141 ;
  assign \DISPNUM2[0]_pad  = n168 ;
  assign \DISPNUM2[1]_pad  = n172 ;
  assign \DISPNUM2[2]_pad  = n178 ;
  assign \DISPNUM2[3]_pad  = n180 ;
  assign \DISPNUM2[4]_pad  = n182 ;
  assign \DISPNUM2[5]_pad  = n186 ;
  assign \DISPNUM2[6]_pad  = n190 ;
  assign SIGN_pad = n192 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g2955/_2_  = ~n431 ;
  assign \g2956/_2_  = ~n442 ;
  assign \g2957/_2_  = ~n453 ;
  assign \g2958/_2_  = ~n464 ;
  assign \g2959/_2_  = ~n475 ;
  assign \g2960/_2_  = ~n486 ;
  assign \g2961/_2_  = ~n497 ;
  assign \g2962/_2_  = ~n508 ;
  assign \g2963/_2_  = ~n519 ;
  assign \g2985/_0_  = ~n528 ;
  assign \g3032/_0_  = ~n536 ;
  assign \g3033/_0_  = ~n545 ;
  assign \g3034/_0_  = ~n552 ;
  assign \g3038/_0_  = ~n555 ;
  assign \g3247/_0_  = ~n561 ;
  assign \g3279/_0_  = ~n564 ;
  assign \g3309/_0_  = ~n573 ;
  assign \g3335/_0_  = ~n576 ;
  assign \g3336/_0_  = ~n579 ;
  assign \g3337/_0_  = ~n582 ;
  assign \g3338/_0_  = ~n585 ;
  assign \g3339/_0_  = ~n588 ;
  assign \g3340/_0_  = ~n591 ;
  assign \g3341/_0_  = ~n594 ;
  assign \g3360/_0_  = ~n600 ;
  assign \g3361/_0_  = ~n606 ;
  assign \g3369/_0_  = ~n612 ;
  assign \g3373/_0_  = ~n616 ;
  assign \g3382/_0_  = ~n619 ;
  assign \g3451/_0_  = ~n622 ;
  assign \g3475/_0_  = ~n624 ;
  assign \g3490/_0_  = n627 ;
  assign \g3514/_0_  = ~n629 ;
  assign \g3774/_1_  = n63 ;
  assign \g4511/_0_  = ~n632 ;
endmodule
