module top (ACCRPY_pad, \BULL0_pad , \BULL1_pad , \BULL2_pad , \BULL3_pad , \BULL4_pad , \BULL5_pad , \BULL6_pad , CAPSD_pad, \CAT0_pad , \CAT1_pad , \CAT2_pad , \CAT3_pad , \CAT4_pad , \CAT5_pad , COMPPAR_pad, \DEL1_pad , END_pad, FBI_pad, \IBT0_pad , \IBT1_pad , \IBT2_pad , ICLR_pad, KBG_N_pad, LSD_pad, MARSSR_pad, MMERR_pad, ORWD_N_pad, OVACC_pad, OWL_N_pad, \PLUTO0_pad , \PLUTO1_pad , \PLUTO2_pad , \PLUTO3_pad , \PLUTO4_pad , \PLUTO5_pad , PY_pad, RATR_pad, SDO_pad, \STAR0_pad , \STAR1_pad , \STAR2_pad , \STAR3_pad , VACC_pad, VERR_N_pad, VLENESR_pad, \VST1_pad , VSUMESR_pad, WATCH_pad, ACCRPY_P_pad, \BULL0_P_pad , \BULL1_P_pad , \BULL2_P_pad , \BULL3_P_pad , \BULL4_P_pad , \BULL5_P_pad , \BULL6_P_pad , COMPPAR_P_pad, \DEL1_P_pad , END_P_pad, KBG_F_pad, LSD_P_pad, MARSSR_P_pad, ORWD_F_pad, OVACC_P_pad, OWL_F_pad, \PLUTO0_P_pad , \PLUTO1_P_pad , \PLUTO2_P_pad , \PLUTO3_P_pad , \PLUTO4_P_pad , \PLUTO5_P_pad , PY_P_pad, RATR_P_pad, \STAR0_P_pad , \STAR1_P_pad , \STAR2_P_pad , \STAR3_P_pad , VERR_F_pad, VLENESR_P_pad, \VST0_P_pad , \VST1_P_pad , VSUMESR_P_pad, WATCH_P_pad, \n1022 );
	input ACCRPY_pad ;
	input \BULL0_pad  ;
	input \BULL1_pad  ;
	input \BULL2_pad  ;
	input \BULL3_pad  ;
	input \BULL4_pad  ;
	input \BULL5_pad  ;
	input \BULL6_pad  ;
	input CAPSD_pad ;
	input \CAT0_pad  ;
	input \CAT1_pad  ;
	input \CAT2_pad  ;
	input \CAT3_pad  ;
	input \CAT4_pad  ;
	input \CAT5_pad  ;
	input COMPPAR_pad ;
	input \DEL1_pad  ;
	input END_pad ;
	input FBI_pad ;
	input \IBT0_pad  ;
	input \IBT1_pad  ;
	input \IBT2_pad  ;
	input ICLR_pad ;
	input KBG_N_pad ;
	input LSD_pad ;
	input MARSSR_pad ;
	input MMERR_pad ;
	input ORWD_N_pad ;
	input OVACC_pad ;
	input OWL_N_pad ;
	input \PLUTO0_pad  ;
	input \PLUTO1_pad  ;
	input \PLUTO2_pad  ;
	input \PLUTO3_pad  ;
	input \PLUTO4_pad  ;
	input \PLUTO5_pad  ;
	input PY_pad ;
	input RATR_pad ;
	input SDO_pad ;
	input \STAR0_pad  ;
	input \STAR1_pad  ;
	input \STAR2_pad  ;
	input \STAR3_pad  ;
	input VACC_pad ;
	input VERR_N_pad ;
	input VLENESR_pad ;
	input \VST1_pad  ;
	input VSUMESR_pad ;
	input WATCH_pad ;
	output ACCRPY_P_pad ;
	output \BULL0_P_pad  ;
	output \BULL1_P_pad  ;
	output \BULL2_P_pad  ;
	output \BULL3_P_pad  ;
	output \BULL4_P_pad  ;
	output \BULL5_P_pad  ;
	output \BULL6_P_pad  ;
	output COMPPAR_P_pad ;
	output \DEL1_P_pad  ;
	output END_P_pad ;
	output KBG_F_pad ;
	output LSD_P_pad ;
	output MARSSR_P_pad ;
	output ORWD_F_pad ;
	output OVACC_P_pad ;
	output OWL_F_pad ;
	output \PLUTO0_P_pad  ;
	output \PLUTO1_P_pad  ;
	output \PLUTO2_P_pad  ;
	output \PLUTO3_P_pad  ;
	output \PLUTO4_P_pad  ;
	output \PLUTO5_P_pad  ;
	output PY_P_pad ;
	output RATR_P_pad ;
	output \STAR0_P_pad  ;
	output \STAR1_P_pad  ;
	output \STAR2_P_pad  ;
	output \STAR3_P_pad  ;
	output VERR_F_pad ;
	output VLENESR_P_pad ;
	output \VST0_P_pad  ;
	output \VST1_P_pad  ;
	output VSUMESR_P_pad ;
	output WATCH_P_pad ;
	output \n1022  ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w149_ ;
	wire _w148_ ;
	wire _w147_ ;
	wire _w146_ ;
	wire _w145_ ;
	wire _w144_ ;
	wire _w143_ ;
	wire _w142_ ;
	wire _w141_ ;
	wire _w140_ ;
	wire _w139_ ;
	wire _w138_ ;
	wire _w137_ ;
	wire _w136_ ;
	wire _w135_ ;
	wire _w134_ ;
	wire _w133_ ;
	wire _w132_ ;
	wire _w131_ ;
	wire _w130_ ;
	wire _w129_ ;
	wire _w128_ ;
	wire _w127_ ;
	wire _w126_ ;
	wire _w125_ ;
	wire _w124_ ;
	wire _w123_ ;
	wire _w122_ ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w58_ ;
	wire _w59_ ;
	wire _w60_ ;
	wire _w61_ ;
	wire _w62_ ;
	wire _w63_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	LUT3 #(
		.INIT('h35)
	) name0 (
		\CAT2_pad ,
		\CAT3_pad ,
		\IBT0_pad ,
		_w51_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		\IBT2_pad ,
		WATCH_pad,
		_w52_
	);
	LUT3 #(
		.INIT('h35)
	) name2 (
		\CAT4_pad ,
		\CAT5_pad ,
		\IBT0_pad ,
		_w53_
	);
	LUT4 #(
		.INIT('h1fbf)
	) name3 (
		\IBT1_pad ,
		_w51_,
		_w52_,
		_w53_,
		_w54_
	);
	LUT4 #(
		.INIT('h0070)
	) name4 (
		\CAT1_pad ,
		\IBT0_pad ,
		\IBT1_pad ,
		\IBT2_pad ,
		_w55_
	);
	LUT2 #(
		.INIT('h2)
	) name5 (
		\CAT0_pad ,
		\IBT0_pad ,
		_w56_
	);
	LUT3 #(
		.INIT('hd0)
	) name6 (
		\CAT0_pad ,
		\IBT0_pad ,
		WATCH_pad,
		_w57_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w55_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\STAR0_pad ,
		\STAR1_pad ,
		_w59_
	);
	LUT4 #(
		.INIT('h0080)
	) name9 (
		FBI_pad,
		\STAR0_pad ,
		\STAR1_pad ,
		\STAR2_pad ,
		_w60_
	);
	LUT3 #(
		.INIT('h70)
	) name10 (
		_w55_,
		_w57_,
		_w60_,
		_w61_
	);
	LUT4 #(
		.INIT('hc888)
	) name11 (
		ACCRPY_pad,
		OWL_N_pad,
		_w54_,
		_w61_,
		_w62_
	);
	LUT3 #(
		.INIT('h48)
	) name12 (
		\BULL0_pad ,
		OWL_N_pad,
		WATCH_pad,
		_w63_
	);
	LUT3 #(
		.INIT('h80)
	) name13 (
		\BULL0_pad ,
		\BULL1_pad ,
		WATCH_pad,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		OWL_N_pad,
		WATCH_pad,
		_w65_
	);
	LUT4 #(
		.INIT('h60c0)
	) name15 (
		\BULL0_pad ,
		\BULL1_pad ,
		OWL_N_pad,
		WATCH_pad,
		_w66_
	);
	LUT4 #(
		.INIT('h070f)
	) name16 (
		\BULL0_pad ,
		\BULL1_pad ,
		\BULL2_pad ,
		WATCH_pad,
		_w67_
	);
	LUT4 #(
		.INIT('h8000)
	) name17 (
		\BULL0_pad ,
		\BULL1_pad ,
		\BULL2_pad ,
		WATCH_pad,
		_w68_
	);
	LUT3 #(
		.INIT('h02)
	) name18 (
		OWL_N_pad,
		_w67_,
		_w68_,
		_w69_
	);
	LUT3 #(
		.INIT('h48)
	) name19 (
		\BULL3_pad ,
		OWL_N_pad,
		_w68_,
		_w70_
	);
	LUT4 #(
		.INIT('h60c0)
	) name20 (
		\BULL3_pad ,
		\BULL4_pad ,
		OWL_N_pad,
		_w68_,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\BULL5_pad ,
		OWL_N_pad,
		_w72_
	);
	LUT4 #(
		.INIT('h2800)
	) name22 (
		\BULL3_pad ,
		\BULL4_pad ,
		\BULL5_pad ,
		OWL_N_pad,
		_w73_
	);
	LUT4 #(
		.INIT('hfc70)
	) name23 (
		\BULL3_pad ,
		_w68_,
		_w72_,
		_w73_,
		_w74_
	);
	LUT4 #(
		.INIT('h8000)
	) name24 (
		\BULL2_pad ,
		\BULL3_pad ,
		\BULL4_pad ,
		\BULL5_pad ,
		_w75_
	);
	LUT4 #(
		.INIT('hf755)
	) name25 (
		\BULL6_pad ,
		OWL_N_pad,
		_w64_,
		_w75_,
		_w76_
	);
	LUT4 #(
		.INIT('h0080)
	) name26 (
		\BULL3_pad ,
		\BULL4_pad ,
		\BULL5_pad ,
		\BULL6_pad ,
		_w77_
	);
	LUT2 #(
		.INIT('h8)
	) name27 (
		_w68_,
		_w77_,
		_w78_
	);
	LUT3 #(
		.INIT('ha2)
	) name28 (
		OWL_N_pad,
		_w76_,
		_w78_,
		_w79_
	);
	LUT4 #(
		.INIT('h6a00)
	) name29 (
		COMPPAR_pad,
		\DEL1_pad ,
		FBI_pad,
		OWL_N_pad,
		_w80_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		CAPSD_pad,
		ICLR_pad,
		_w81_
	);
	LUT4 #(
		.INIT('hc888)
	) name31 (
		END_pad,
		OWL_N_pad,
		_w54_,
		_w61_,
		_w82_
	);
	LUT2 #(
		.INIT('h2)
	) name32 (
		_w54_,
		_w58_,
		_w83_
	);
	LUT3 #(
		.INIT('h20)
	) name33 (
		FBI_pad,
		\STAR2_pad ,
		\STAR3_pad ,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w59_,
		_w84_,
		_w85_
	);
	LUT3 #(
		.INIT('hd0)
	) name35 (
		_w54_,
		_w58_,
		_w85_,
		_w86_
	);
	LUT3 #(
		.INIT('h08)
	) name36 (
		\STAR0_pad ,
		\STAR1_pad ,
		\STAR2_pad ,
		_w87_
	);
	LUT4 #(
		.INIT('haa2a)
	) name37 (
		FBI_pad,
		\STAR0_pad ,
		\STAR1_pad ,
		\STAR2_pad ,
		_w88_
	);
	LUT3 #(
		.INIT('h70)
	) name38 (
		_w55_,
		_w57_,
		_w88_,
		_w89_
	);
	LUT3 #(
		.INIT('h2a)
	) name39 (
		KBG_N_pad,
		_w54_,
		_w89_,
		_w90_
	);
	LUT3 #(
		.INIT('h75)
	) name40 (
		OWL_N_pad,
		_w86_,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		LSD_pad,
		OWL_N_pad,
		_w92_
	);
	LUT3 #(
		.INIT('h70)
	) name42 (
		_w59_,
		_w84_,
		_w92_,
		_w93_
	);
	LUT4 #(
		.INIT('h002a)
	) name43 (
		FBI_pad,
		LSD_pad,
		OWL_N_pad,
		\STAR3_pad ,
		_w94_
	);
	LUT3 #(
		.INIT('h80)
	) name44 (
		_w65_,
		_w87_,
		_w94_,
		_w95_
	);
	LUT4 #(
		.INIT('h37bf)
	) name45 (
		\IBT1_pad ,
		\IBT2_pad ,
		_w51_,
		_w53_,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name46 (
		_w55_,
		_w56_,
		_w97_
	);
	LUT4 #(
		.INIT('heeae)
	) name47 (
		_w93_,
		_w95_,
		_w96_,
		_w97_,
		_w98_
	);
	LUT4 #(
		.INIT('h0400)
	) name48 (
		\BULL3_pad ,
		\BULL4_pad ,
		\BULL5_pad ,
		\BULL6_pad ,
		_w99_
	);
	LUT4 #(
		.INIT('h0400)
	) name49 (
		\BULL0_pad ,
		\BULL1_pad ,
		\BULL2_pad ,
		WATCH_pad,
		_w100_
	);
	LUT4 #(
		.INIT('hc888)
	) name50 (
		MARSSR_pad,
		OWL_N_pad,
		_w99_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		ICLR_pad,
		VACC_pad,
		_w102_
	);
	LUT3 #(
		.INIT('h10)
	) name52 (
		END_pad,
		ICLR_pad,
		KBG_N_pad,
		_w103_
	);
	LUT3 #(
		.INIT('h70)
	) name53 (
		_w99_,
		_w100_,
		_w103_,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name54 (
		OWL_N_pad,
		\PLUTO0_pad ,
		_w105_
	);
	LUT4 #(
		.INIT('h0400)
	) name55 (
		\IBT0_pad ,
		\IBT1_pad ,
		\IBT2_pad ,
		OWL_N_pad,
		_w106_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w105_,
		_w106_,
		_w107_
	);
	LUT3 #(
		.INIT('h2a)
	) name57 (
		KBG_N_pad,
		_w99_,
		_w100_,
		_w108_
	);
	LUT4 #(
		.INIT('h00a8)
	) name58 (
		COMPPAR_pad,
		MMERR_pad,
		SDO_pad,
		\VST1_pad ,
		_w109_
	);
	LUT2 #(
		.INIT('h2)
	) name59 (
		END_pad,
		_w109_,
		_w110_
	);
	LUT3 #(
		.INIT('h31)
	) name60 (
		END_pad,
		_w105_,
		_w109_,
		_w111_
	);
	LUT3 #(
		.INIT('h15)
	) name61 (
		_w107_,
		_w108_,
		_w111_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		OWL_N_pad,
		\PLUTO1_pad ,
		_w113_
	);
	LUT4 #(
		.INIT('h0800)
	) name63 (
		\IBT0_pad ,
		\IBT1_pad ,
		\IBT2_pad ,
		OWL_N_pad,
		_w114_
	);
	LUT4 #(
		.INIT('hfdf0)
	) name64 (
		_w108_,
		_w110_,
		_w113_,
		_w114_,
		_w115_
	);
	LUT2 #(
		.INIT('h8)
	) name65 (
		OWL_N_pad,
		\PLUTO2_pad ,
		_w116_
	);
	LUT4 #(
		.INIT('h1000)
	) name66 (
		\IBT0_pad ,
		\IBT1_pad ,
		\IBT2_pad ,
		OWL_N_pad,
		_w117_
	);
	LUT4 #(
		.INIT('hfdf0)
	) name67 (
		_w108_,
		_w110_,
		_w116_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		OWL_N_pad,
		\PLUTO3_pad ,
		_w119_
	);
	LUT4 #(
		.INIT('h2000)
	) name69 (
		\IBT0_pad ,
		\IBT1_pad ,
		\IBT2_pad ,
		OWL_N_pad,
		_w120_
	);
	LUT4 #(
		.INIT('hfdf0)
	) name70 (
		_w108_,
		_w110_,
		_w119_,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h8)
	) name71 (
		OWL_N_pad,
		\PLUTO4_pad ,
		_w122_
	);
	LUT4 #(
		.INIT('h4000)
	) name72 (
		\IBT0_pad ,
		\IBT1_pad ,
		\IBT2_pad ,
		OWL_N_pad,
		_w123_
	);
	LUT4 #(
		.INIT('hfdf0)
	) name73 (
		_w108_,
		_w110_,
		_w122_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		OWL_N_pad,
		\PLUTO5_pad ,
		_w125_
	);
	LUT4 #(
		.INIT('h8000)
	) name75 (
		\IBT0_pad ,
		\IBT1_pad ,
		\IBT2_pad ,
		OWL_N_pad,
		_w126_
	);
	LUT4 #(
		.INIT('hfdf0)
	) name76 (
		_w108_,
		_w110_,
		_w125_,
		_w126_,
		_w127_
	);
	LUT4 #(
		.INIT('h0b08)
	) name77 (
		\DEL1_pad ,
		FBI_pad,
		ICLR_pad,
		PY_pad,
		_w128_
	);
	LUT4 #(
		.INIT('h0a08)
	) name78 (
		COMPPAR_pad,
		MMERR_pad,
		RATR_pad,
		SDO_pad,
		_w129_
	);
	LUT3 #(
		.INIT('hc8)
	) name79 (
		END_pad,
		OWL_N_pad,
		RATR_pad,
		_w130_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		_w129_,
		_w130_,
		_w131_
	);
	LUT3 #(
		.INIT('hb0)
	) name81 (
		FBI_pad,
		OWL_N_pad,
		\STAR0_pad ,
		_w132_
	);
	LUT4 #(
		.INIT('h40ff)
	) name82 (
		FBI_pad,
		ORWD_N_pad,
		OWL_N_pad,
		\STAR0_pad ,
		_w133_
	);
	LUT3 #(
		.INIT('h07)
	) name83 (
		_w55_,
		_w57_,
		_w132_,
		_w134_
	);
	LUT3 #(
		.INIT('h13)
	) name84 (
		_w54_,
		_w133_,
		_w134_,
		_w135_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		FBI_pad,
		OWL_N_pad,
		_w136_
	);
	LUT3 #(
		.INIT('h4f)
	) name86 (
		FBI_pad,
		ORWD_N_pad,
		OWL_N_pad,
		_w137_
	);
	LUT3 #(
		.INIT('h07)
	) name87 (
		_w55_,
		_w57_,
		_w136_,
		_w138_
	);
	LUT4 #(
		.INIT('h5450)
	) name88 (
		\STAR0_pad ,
		_w54_,
		_w137_,
		_w138_,
		_w139_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w135_,
		_w139_,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		FBI_pad,
		ORWD_N_pad,
		_w141_
	);
	LUT3 #(
		.INIT('h15)
	) name91 (
		FBI_pad,
		_w55_,
		_w57_,
		_w142_
	);
	LUT4 #(
		.INIT('h040c)
	) name92 (
		_w54_,
		_w59_,
		_w141_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		OWL_N_pad,
		\STAR1_pad ,
		_w144_
	);
	LUT4 #(
		.INIT('hec00)
	) name94 (
		_w54_,
		_w133_,
		_w134_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		\STAR0_pad ,
		\STAR1_pad ,
		_w146_
	);
	LUT4 #(
		.INIT('h1300)
	) name96 (
		_w54_,
		_w137_,
		_w138_,
		_w146_,
		_w147_
	);
	LUT3 #(
		.INIT('hf4)
	) name97 (
		_w143_,
		_w145_,
		_w147_,
		_w148_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		OWL_N_pad,
		\STAR2_pad ,
		_w149_
	);
	LUT4 #(
		.INIT('h040c)
	) name99 (
		_w54_,
		_w87_,
		_w137_,
		_w138_,
		_w150_
	);
	LUT3 #(
		.INIT('hf4)
	) name100 (
		_w143_,
		_w149_,
		_w150_,
		_w151_
	);
	LUT3 #(
		.INIT('h80)
	) name101 (
		\STAR0_pad ,
		\STAR1_pad ,
		\STAR2_pad ,
		_w152_
	);
	LUT4 #(
		.INIT('h1300)
	) name102 (
		_w54_,
		_w141_,
		_w142_,
		_w152_,
		_w153_
	);
	LUT4 #(
		.INIT('h8000)
	) name103 (
		FBI_pad,
		\STAR0_pad ,
		\STAR1_pad ,
		\STAR2_pad ,
		_w154_
	);
	LUT4 #(
		.INIT('h4000)
	) name104 (
		ORWD_N_pad,
		\STAR0_pad ,
		\STAR1_pad ,
		\STAR2_pad ,
		_w155_
	);
	LUT4 #(
		.INIT('h020f)
	) name105 (
		_w54_,
		_w58_,
		_w154_,
		_w155_,
		_w156_
	);
	LUT4 #(
		.INIT('h082a)
	) name106 (
		OWL_N_pad,
		\STAR3_pad ,
		_w153_,
		_w156_,
		_w157_
	);
	LUT3 #(
		.INIT('h2a)
	) name107 (
		VERR_N_pad,
		_w99_,
		_w100_,
		_w158_
	);
	LUT3 #(
		.INIT('h70)
	) name108 (
		_w54_,
		_w89_,
		_w158_,
		_w159_
	);
	LUT3 #(
		.INIT('h75)
	) name109 (
		OWL_N_pad,
		_w86_,
		_w159_,
		_w160_
	);
	LUT3 #(
		.INIT('hc4)
	) name110 (
		KBG_N_pad,
		OWL_N_pad,
		VLENESR_pad,
		_w161_
	);
	LUT4 #(
		.INIT('h3210)
	) name111 (
		FBI_pad,
		ICLR_pad,
		SDO_pad,
		\VST1_pad ,
		_w162_
	);
	LUT4 #(
		.INIT('h3120)
	) name112 (
		FBI_pad,
		ICLR_pad,
		PY_pad,
		\VST1_pad ,
		_w163_
	);
	LUT4 #(
		.INIT('hcc80)
	) name113 (
		END_pad,
		OWL_N_pad,
		\VST1_pad ,
		VSUMESR_pad,
		_w164_
	);
	LUT4 #(
		.INIT('hcc08)
	) name114 (
		OVACC_pad,
		OWL_N_pad,
		VACC_pad,
		WATCH_pad,
		_w165_
	);
	LUT3 #(
		.INIT('h70)
	) name115 (
		_w55_,
		_w57_,
		_w87_,
		_w166_
	);
	LUT4 #(
		.INIT('h1113)
	) name116 (
		_w54_,
		_w137_,
		_w138_,
		_w166_,
		_w167_
	);
	assign ACCRPY_P_pad = _w62_ ;
	assign \BULL0_P_pad  = _w63_ ;
	assign \BULL1_P_pad  = _w66_ ;
	assign \BULL2_P_pad  = _w69_ ;
	assign \BULL3_P_pad  = _w70_ ;
	assign \BULL4_P_pad  = _w71_ ;
	assign \BULL5_P_pad  = _w74_ ;
	assign \BULL6_P_pad  = _w79_ ;
	assign COMPPAR_P_pad = _w80_ ;
	assign \DEL1_P_pad  = _w81_ ;
	assign END_P_pad = _w82_ ;
	assign KBG_F_pad = _w91_ ;
	assign LSD_P_pad = _w98_ ;
	assign MARSSR_P_pad = _w101_ ;
	assign ORWD_F_pad = _w83_ ;
	assign OVACC_P_pad = _w102_ ;
	assign OWL_F_pad = _w104_ ;
	assign \PLUTO0_P_pad  = _w112_ ;
	assign \PLUTO1_P_pad  = _w115_ ;
	assign \PLUTO2_P_pad  = _w118_ ;
	assign \PLUTO3_P_pad  = _w121_ ;
	assign \PLUTO4_P_pad  = _w124_ ;
	assign \PLUTO5_P_pad  = _w127_ ;
	assign PY_P_pad = _w128_ ;
	assign RATR_P_pad = _w131_ ;
	assign \STAR0_P_pad  = _w140_ ;
	assign \STAR1_P_pad  = _w148_ ;
	assign \STAR2_P_pad  = _w151_ ;
	assign \STAR3_P_pad  = _w157_ ;
	assign VERR_F_pad = _w160_ ;
	assign VLENESR_P_pad = _w161_ ;
	assign \VST0_P_pad  = _w162_ ;
	assign \VST1_P_pad  = _w163_ ;
	assign VSUMESR_P_pad = _w164_ ;
	assign WATCH_P_pad = _w165_ ;
	assign \n1022  = _w167_ ;
endmodule;