module top (\G0_pad , \G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G18_pad , \G1_pad , \G2_pad , \G38_reg/NET0131 , \G39_reg/NET0131 , \G3_pad , \G40_reg/NET0131 , \G41_reg/NET0131 , \G42_reg/NET0131 , \G4_pad , \G5_pad , \G6_pad , \G7_pad , \G8_pad , \G9_pad , \G288_pad , \G290_pad , \G296_pad , \G302_pad , \G315_pad , \G325_pad , \G327_pad , \G45_pad , \G47_pad , \G49_pad , \G53_pad , \G55_pad , \_al_n0 , \_al_n1 , \g1404/_0_ , \g1412/_0_ , \g1416/_0_ , \g1451/_2_ , \g1459/_3_ , \g1511/_3_ , \g1527/_3_ , \g1529/_3_ , \g31/_0_ , \g33/_1_ , \g56/_3_ );
	input \G0_pad  ;
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G18_pad  ;
	input \G1_pad  ;
	input \G2_pad  ;
	input \G38_reg/NET0131  ;
	input \G39_reg/NET0131  ;
	input \G3_pad  ;
	input \G40_reg/NET0131  ;
	input \G41_reg/NET0131  ;
	input \G42_reg/NET0131  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G6_pad  ;
	input \G7_pad  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G288_pad  ;
	output \G290_pad  ;
	output \G296_pad  ;
	output \G302_pad  ;
	output \G315_pad  ;
	output \G325_pad  ;
	output \G327_pad  ;
	output \G45_pad  ;
	output \G47_pad  ;
	output \G49_pad  ;
	output \G53_pad  ;
	output \G55_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1404/_0_  ;
	output \g1412/_0_  ;
	output \g1416/_0_  ;
	output \g1451/_2_  ;
	output \g1459/_3_  ;
	output \g1511/_3_  ;
	output \g1527/_3_  ;
	output \g1529/_3_  ;
	output \g31/_0_  ;
	output \g33/_1_  ;
	output \g56/_3_  ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w195_ ;
	wire _w194_ ;
	wire _w193_ ;
	wire _w192_ ;
	wire _w191_ ;
	wire _w190_ ;
	wire _w189_ ;
	wire _w188_ ;
	wire _w187_ ;
	wire _w186_ ;
	wire _w185_ ;
	wire _w184_ ;
	wire _w183_ ;
	wire _w182_ ;
	wire _w181_ ;
	wire _w180_ ;
	wire _w179_ ;
	wire _w178_ ;
	wire _w177_ ;
	wire _w176_ ;
	wire _w175_ ;
	wire _w174_ ;
	wire _w173_ ;
	wire _w172_ ;
	wire _w171_ ;
	wire _w170_ ;
	wire _w169_ ;
	wire _w168_ ;
	wire _w167_ ;
	wire _w166_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w82_ ;
	wire _w81_ ;
	wire _w80_ ;
	wire _w79_ ;
	wire _w78_ ;
	wire _w77_ ;
	wire _w76_ ;
	wire _w75_ ;
	wire _w74_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w36_ ;
	wire _w35_ ;
	wire _w34_ ;
	wire _w33_ ;
	wire _w32_ ;
	wire _w31_ ;
	wire _w30_ ;
	wire _w29_ ;
	wire _w28_ ;
	wire _w27_ ;
	wire _w26_ ;
	wire _w25_ ;
	wire _w24_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w42_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	wire _w104_ ;
	wire _w105_ ;
	wire _w106_ ;
	wire _w107_ ;
	wire _w108_ ;
	wire _w109_ ;
	wire _w110_ ;
	wire _w111_ ;
	wire _w112_ ;
	wire _w113_ ;
	wire _w114_ ;
	wire _w115_ ;
	wire _w116_ ;
	wire _w117_ ;
	wire _w118_ ;
	wire _w119_ ;
	wire _w120_ ;
	wire _w121_ ;
	wire _w122_ ;
	wire _w123_ ;
	wire _w124_ ;
	wire _w125_ ;
	wire _w126_ ;
	wire _w127_ ;
	wire _w128_ ;
	wire _w129_ ;
	wire _w130_ ;
	wire _w131_ ;
	wire _w132_ ;
	wire _w133_ ;
	wire _w134_ ;
	wire _w135_ ;
	wire _w136_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w150_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w24_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w25_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\G42_reg/NET0131 ,
		_w25_,
		_w26_
	);
	LUT2 #(
		.INIT('h8)
	) name3 (
		_w24_,
		_w26_,
		_w27_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w28_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\G15_pad ,
		\G39_reg/NET0131 ,
		_w29_
	);
	LUT2 #(
		.INIT('h4)
	) name6 (
		\G42_reg/NET0131 ,
		_w28_,
		_w30_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w29_,
		_w30_,
		_w31_
	);
	LUT2 #(
		.INIT('h8)
	) name8 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w32_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		\G42_reg/NET0131 ,
		_w32_,
		_w33_
	);
	LUT2 #(
		.INIT('h4)
	) name10 (
		\G38_reg/NET0131 ,
		_w33_,
		_w34_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\G39_reg/NET0131 ,
		_w34_,
		_w35_
	);
	LUT2 #(
		.INIT('h2)
	) name12 (
		\G16_pad ,
		\G4_pad ,
		_w36_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w37_
	);
	LUT2 #(
		.INIT('h8)
	) name14 (
		\G40_reg/NET0131 ,
		_w37_,
		_w38_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		\G38_reg/NET0131 ,
		_w38_,
		_w39_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		\G40_reg/NET0131 ,
		_w37_,
		_w40_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\G39_reg/NET0131 ,
		_w40_,
		_w41_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		_w39_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h4)
	) name19 (
		_w36_,
		_w42_,
		_w43_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w44_
	);
	LUT2 #(
		.INIT('h8)
	) name21 (
		\G38_reg/NET0131 ,
		_w44_,
		_w45_
	);
	LUT2 #(
		.INIT('h2)
	) name22 (
		\G40_reg/NET0131 ,
		_w45_,
		_w46_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		\G4_pad ,
		_w46_,
		_w47_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\G16_pad ,
		_w37_,
		_w48_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		\G40_reg/NET0131 ,
		_w48_,
		_w49_
	);
	LUT2 #(
		.INIT('h1)
	) name26 (
		_w47_,
		_w49_,
		_w50_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\G39_reg/NET0131 ,
		_w50_,
		_w51_
	);
	LUT2 #(
		.INIT('h2)
	) name28 (
		\G16_pad ,
		\G38_reg/NET0131 ,
		_w52_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		\G39_reg/NET0131 ,
		\G40_reg/NET0131 ,
		_w53_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w44_,
		_w53_,
		_w54_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\G1_pad ,
		_w52_,
		_w55_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		_w43_,
		_w56_,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name34 (
		_w51_,
		_w57_,
		_w58_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w24_,
		_w37_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w54_,
		_w59_,
		_w60_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		\G38_reg/NET0131 ,
		_w60_,
		_w61_
	);
	LUT2 #(
		.INIT('h8)
	) name38 (
		\G42_reg/NET0131 ,
		_w24_,
		_w62_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w25_,
		_w62_,
		_w63_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\G42_reg/NET0131 ,
		_w29_,
		_w64_
	);
	LUT2 #(
		.INIT('h8)
	) name41 (
		_w28_,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		\G10_pad ,
		\G11_pad ,
		_w66_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\G10_pad ,
		\G11_pad ,
		_w67_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\G12_pad ,
		_w67_,
		_w68_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w69_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		\G15_pad ,
		_w52_,
		_w70_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w66_,
		_w69_,
		_w71_
	);
	LUT2 #(
		.INIT('h8)
	) name48 (
		_w70_,
		_w71_,
		_w72_
	);
	LUT2 #(
		.INIT('h2)
	) name49 (
		_w33_,
		_w68_,
		_w73_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		_w72_,
		_w73_,
		_w74_
	);
	LUT2 #(
		.INIT('h4)
	) name51 (
		\G5_pad ,
		_w27_,
		_w75_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\G39_reg/NET0131 ,
		_w46_,
		_w76_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w42_,
		_w76_,
		_w77_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\G40_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w78_
	);
	LUT2 #(
		.INIT('h4)
	) name55 (
		\G42_reg/NET0131 ,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w80_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w79_,
		_w80_,
		_w81_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\G5_pad ,
		_w27_,
		_w82_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		\G6_pad ,
		\G7_pad ,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name60 (
		\G8_pad ,
		\G9_pad ,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name61 (
		_w83_,
		_w84_,
		_w85_
	);
	LUT2 #(
		.INIT('h1)
	) name62 (
		\G40_reg/NET0131 ,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h8)
	) name63 (
		\G38_reg/NET0131 ,
		\G39_reg/NET0131 ,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w86_,
		_w87_,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		_w89_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\G38_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w90_
	);
	LUT2 #(
		.INIT('h2)
	) name67 (
		\G40_reg/NET0131 ,
		_w90_,
		_w91_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		\G13_pad ,
		\G15_pad ,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name69 (
		\G42_reg/NET0131 ,
		_w92_,
		_w93_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		\G15_pad ,
		\G42_reg/NET0131 ,
		_w94_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		_w91_,
		_w94_,
		_w95_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w93_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\G39_reg/NET0131 ,
		_w96_,
		_w97_
	);
	LUT2 #(
		.INIT('h2)
	) name74 (
		\G41_reg/NET0131 ,
		_w89_,
		_w98_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		_w88_,
		_w98_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w97_,
		_w99_,
		_w100_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		\G1_pad ,
		_w28_,
		_w101_
	);
	LUT2 #(
		.INIT('h8)
	) name78 (
		\G15_pad ,
		\G40_reg/NET0131 ,
		_w102_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		\G42_reg/NET0131 ,
		\G6_pad ,
		_w103_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		\G7_pad ,
		\G8_pad ,
		_w104_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		\G9_pad ,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		_w102_,
		_w103_,
		_w106_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		_w105_,
		_w106_,
		_w107_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w101_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h2)
	) name85 (
		_w80_,
		_w108_,
		_w109_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		\G41_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w110_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		\G39_reg/NET0131 ,
		_w110_,
		_w111_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		\G40_reg/NET0131 ,
		_w94_,
		_w112_
	);
	LUT2 #(
		.INIT('h4)
	) name89 (
		_w64_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name90 (
		_w111_,
		_w113_,
		_w114_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		_w115_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\G39_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w116_
	);
	LUT2 #(
		.INIT('h8)
	) name93 (
		_w115_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('h1)
	) name94 (
		_w114_,
		_w117_,
		_w118_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		_w109_,
		_w118_,
		_w119_
	);
	LUT2 #(
		.INIT('h4)
	) name96 (
		_w100_,
		_w119_,
		_w120_
	);
	LUT2 #(
		.INIT('h2)
	) name97 (
		\G16_pad ,
		_w120_,
		_w121_
	);
	LUT2 #(
		.INIT('h2)
	) name98 (
		\G15_pad ,
		\G39_reg/NET0131 ,
		_w122_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\G14_pad ,
		_w122_,
		_w123_
	);
	LUT2 #(
		.INIT('h8)
	) name100 (
		_w79_,
		_w123_,
		_w124_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		\G4_pad ,
		_w40_,
		_w125_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		\G39_reg/NET0131 ,
		_w125_,
		_w126_
	);
	LUT2 #(
		.INIT('h4)
	) name103 (
		\G41_reg/NET0131 ,
		\G5_pad ,
		_w127_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		\G42_reg/NET0131 ,
		_w127_,
		_w128_
	);
	LUT2 #(
		.INIT('h2)
	) name105 (
		\G2_pad ,
		_w128_,
		_w129_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		\G1_pad ,
		\G3_pad ,
		_w130_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		_w110_,
		_w130_,
		_w131_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w128_,
		_w131_,
		_w132_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		_w24_,
		_w129_,
		_w133_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w132_,
		_w133_,
		_w134_
	);
	LUT2 #(
		.INIT('h1)
	) name111 (
		_w124_,
		_w126_,
		_w135_
	);
	LUT2 #(
		.INIT('h4)
	) name112 (
		_w134_,
		_w135_,
		_w136_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\G38_reg/NET0131 ,
		_w136_,
		_w137_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\G4_pad ,
		_w76_,
		_w138_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\G0_pad ,
		\G39_reg/NET0131 ,
		_w139_
	);
	LUT2 #(
		.INIT('h2)
	) name116 (
		\G38_reg/NET0131 ,
		_w69_,
		_w140_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w139_,
		_w140_,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name118 (
		_w38_,
		_w141_,
		_w142_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w138_,
		_w142_,
		_w143_
	);
	LUT2 #(
		.INIT('h4)
	) name120 (
		_w137_,
		_w143_,
		_w144_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		_w121_,
		_w144_,
		_w145_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		\G18_pad ,
		_w145_,
		_w146_
	);
	LUT2 #(
		.INIT('h4)
	) name123 (
		\G38_reg/NET0131 ,
		_w132_,
		_w147_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		\G0_pad ,
		_w37_,
		_w148_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		\G4_pad ,
		_w44_,
		_w149_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\G38_reg/NET0131 ,
		_w148_,
		_w150_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		_w149_,
		_w150_,
		_w151_
	);
	LUT2 #(
		.INIT('h2)
	) name128 (
		_w24_,
		_w147_,
		_w152_
	);
	LUT2 #(
		.INIT('h4)
	) name129 (
		_w151_,
		_w152_,
		_w153_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\G42_reg/NET0131 ,
		_w66_,
		_w154_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\G15_pad ,
		_w32_,
		_w155_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w154_,
		_w155_,
		_w156_
	);
	LUT2 #(
		.INIT('h8)
	) name133 (
		\G16_pad ,
		_w69_,
		_w157_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w89_,
		_w157_,
		_w158_
	);
	LUT2 #(
		.INIT('h4)
	) name135 (
		_w40_,
		_w158_,
		_w159_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w39_,
		_w156_,
		_w160_
	);
	LUT2 #(
		.INIT('h8)
	) name137 (
		_w159_,
		_w160_,
		_w161_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w162_
	);
	LUT2 #(
		.INIT('h4)
	) name139 (
		\G14_pad ,
		\G15_pad ,
		_w163_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\G41_reg/NET0131 ,
		_w163_,
		_w164_
	);
	LUT2 #(
		.INIT('h2)
	) name141 (
		_w162_,
		_w164_,
		_w165_
	);
	LUT2 #(
		.INIT('h8)
	) name142 (
		\G2_pad ,
		_w130_,
		_w166_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		\G16_pad ,
		_w166_,
		_w167_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		\G41_reg/NET0131 ,
		_w167_,
		_w168_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		_w80_,
		_w165_,
		_w169_
	);
	LUT2 #(
		.INIT('h4)
	) name146 (
		_w168_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\G39_reg/NET0131 ,
		\G4_pad ,
		_w171_
	);
	LUT2 #(
		.INIT('h4)
	) name148 (
		\G40_reg/NET0131 ,
		_w171_,
		_w172_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		\G15_pad ,
		\G38_reg/NET0131 ,
		_w173_
	);
	LUT2 #(
		.INIT('h8)
	) name150 (
		_w85_,
		_w173_,
		_w174_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		\G16_pad ,
		_w174_,
		_w175_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w37_,
		_w172_,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name153 (
		_w175_,
		_w176_,
		_w177_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w161_,
		_w170_,
		_w178_
	);
	LUT2 #(
		.INIT('h4)
	) name155 (
		_w177_,
		_w178_,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		_w153_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\G18_pad ,
		_w180_,
		_w181_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		\G39_reg/NET0131 ,
		_w32_,
		_w182_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		\G38_reg/NET0131 ,
		_w33_,
		_w183_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w62_,
		_w182_,
		_w184_
	);
	LUT2 #(
		.INIT('h8)
	) name161 (
		_w183_,
		_w184_,
		_w185_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		\G10_pad ,
		\G12_pad ,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		\G11_pad ,
		_w186_,
		_w187_
	);
	LUT2 #(
		.INIT('h2)
	) name164 (
		_w122_,
		_w187_,
		_w188_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w34_,
		_w188_,
		_w189_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w185_,
		_w189_,
		_w190_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		_w36_,
		_w190_,
		_w191_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		\G0_pad ,
		_w90_,
		_w192_
	);
	LUT2 #(
		.INIT('h8)
	) name169 (
		\G16_pad ,
		\G38_reg/NET0131 ,
		_w193_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		\G16_pad ,
		\G1_pad ,
		_w194_
	);
	LUT2 #(
		.INIT('h4)
	) name171 (
		\G38_reg/NET0131 ,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		\G42_reg/NET0131 ,
		_w195_,
		_w196_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w193_,
		_w196_,
		_w197_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		\G39_reg/NET0131 ,
		_w28_,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w192_,
		_w198_,
		_w199_
	);
	LUT2 #(
		.INIT('h4)
	) name176 (
		_w197_,
		_w199_,
		_w200_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		\G0_pad ,
		_w87_,
		_w201_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\G1_pad ,
		\G39_reg/NET0131 ,
		_w202_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		\G41_reg/NET0131 ,
		_w202_,
		_w203_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w201_,
		_w203_,
		_w204_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\G38_reg/NET0131 ,
		\G41_reg/NET0131 ,
		_w205_
	);
	LUT2 #(
		.INIT('h8)
	) name182 (
		\G40_reg/NET0131 ,
		\G42_reg/NET0131 ,
		_w206_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w205_,
		_w206_,
		_w207_
	);
	LUT2 #(
		.INIT('h4)
	) name184 (
		_w204_,
		_w207_,
		_w208_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		_w200_,
		_w208_,
		_w209_
	);
	LUT2 #(
		.INIT('h4)
	) name186 (
		_w191_,
		_w209_,
		_w210_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		\G18_pad ,
		_w210_,
		_w211_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		\G42_reg/NET0131 ,
		_w53_,
		_w212_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w62_,
		_w212_,
		_w213_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\G1_pad ,
		_w25_,
		_w214_
	);
	LUT2 #(
		.INIT('h4)
	) name191 (
		_w213_,
		_w214_,
		_w215_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\G3_pad ,
		_w54_,
		_w216_
	);
	LUT2 #(
		.INIT('h8)
	) name193 (
		_w195_,
		_w216_,
		_w217_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		_w52_,
		_w59_,
		_w218_
	);
	LUT2 #(
		.INIT('h8)
	) name195 (
		\G15_pad ,
		_w81_,
		_w219_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		\G38_reg/NET0131 ,
		_w124_,
		_w220_
	);
	LUT2 #(
		.INIT('h4)
	) name197 (
		\G16_pad ,
		\G41_reg/NET0131 ,
		_w221_
	);
	LUT2 #(
		.INIT('h2)
	) name198 (
		\G42_reg/NET0131 ,
		_w221_,
		_w222_
	);
	LUT2 #(
		.INIT('h2)
	) name199 (
		\G41_reg/NET0131 ,
		\G4_pad ,
		_w223_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		\G41_reg/NET0131 ,
		\G5_pad ,
		_w224_
	);
	LUT2 #(
		.INIT('h2)
	) name201 (
		\G39_reg/NET0131 ,
		_w224_,
		_w225_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w223_,
		_w225_,
		_w226_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\G40_reg/NET0131 ,
		_w222_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		_w226_,
		_w227_,
		_w228_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		\G16_pad ,
		_w53_,
		_w229_
	);
	LUT2 #(
		.INIT('h1)
	) name206 (
		_w62_,
		_w229_,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name207 (
		\G41_reg/NET0131 ,
		_w166_,
		_w231_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w230_,
		_w231_,
		_w232_
	);
	LUT2 #(
		.INIT('h8)
	) name209 (
		_w102_,
		_w110_,
		_w233_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		\G16_pad ,
		_w162_,
		_w234_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		_w233_,
		_w234_,
		_w235_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		\G39_reg/NET0131 ,
		_w125_,
		_w236_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w165_,
		_w235_,
		_w237_
	);
	LUT2 #(
		.INIT('h8)
	) name214 (
		_w236_,
		_w237_,
		_w238_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w228_,
		_w232_,
		_w239_
	);
	LUT2 #(
		.INIT('h4)
	) name216 (
		_w238_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		\G38_reg/NET0131 ,
		_w240_,
		_w241_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\G16_pad ,
		_w92_,
		_w242_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		_w69_,
		_w242_,
		_w243_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w201_,
		_w243_,
		_w244_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		_w38_,
		_w244_,
		_w245_
	);
	LUT2 #(
		.INIT('h2)
	) name222 (
		\G15_pad ,
		_w44_,
		_w246_
	);
	LUT2 #(
		.INIT('h2)
	) name223 (
		\G16_pad ,
		_w246_,
		_w247_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		_w40_,
		_w171_,
		_w248_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w247_,
		_w248_,
		_w249_
	);
	LUT2 #(
		.INIT('h1)
	) name226 (
		\G39_reg/NET0131 ,
		_w115_,
		_w250_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		\G40_reg/NET0131 ,
		_w223_,
		_w251_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w250_,
		_w251_,
		_w252_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w175_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w245_,
		_w249_,
		_w254_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		_w253_,
		_w254_,
		_w255_
	);
	LUT2 #(
		.INIT('h4)
	) name232 (
		_w241_,
		_w255_,
		_w256_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\G18_pad ,
		_w256_,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name234 (
		_w48_,
		_w172_,
		_w258_
	);
	LUT2 #(
		.INIT('h8)
	) name235 (
		_w68_,
		_w154_,
		_w259_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		\G16_pad ,
		_w122_,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name237 (
		_w223_,
		_w260_,
		_w261_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		_w91_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w259_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		_w26_,
		_w53_,
		_w264_
	);
	LUT2 #(
		.INIT('h8)
	) name241 (
		_w167_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name242 (
		_w258_,
		_w265_,
		_w266_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w263_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w153_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		\G18_pad ,
		_w268_,
		_w269_
	);
	assign \G288_pad  = _w27_ ;
	assign \G290_pad  = _w31_ ;
	assign \G296_pad  = _w35_ ;
	assign \G302_pad  = _w58_ ;
	assign \G315_pad  = _w61_ ;
	assign \G325_pad  = _w63_ ;
	assign \G327_pad  = _w65_ ;
	assign \G45_pad  = _w74_ ;
	assign \G47_pad  = _w75_ ;
	assign \G49_pad  = _w77_ ;
	assign \G53_pad  = _w81_ ;
	assign \G55_pad  = _w82_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g1404/_0_  = _w146_ ;
	assign \g1412/_0_  = _w181_ ;
	assign \g1416/_0_  = _w211_ ;
	assign \g1451/_2_  = _w215_ ;
	assign \g1459/_3_  = _w217_ ;
	assign \g1511/_3_  = _w218_ ;
	assign \g1527/_3_  = _w219_ ;
	assign \g1529/_3_  = _w220_ ;
	assign \g31/_0_  = _w257_ ;
	assign \g33/_1_  = _w269_ ;
	assign \g56/_3_  = _w177_ ;
endmodule;