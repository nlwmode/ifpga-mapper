module top (\a0_pad , \a1_pad , \a2_pad , \a3_pad , \a4_pad , \b0_pad , \b1_pad , \b2_pad , \b3_pad , \b4_pad , b_pad, \c0_pad , \c1_pad , \c2_pad , \c3_pad , \c4_pad , c_pad, \d0_pad , \d1_pad , \d2_pad , \d3_pad , \d4_pad , d_pad, \e0_pad , \e1_pad , \e2_pad , \e3_pad , \e4_pad , e_pad, \f0_pad , \f1_pad , \f2_pad , \f3_pad , \f4_pad , f_pad, \g0_pad , \g1_pad , \g2_pad , \g3_pad , \g4_pad , g_pad, \h0_pad , \h1_pad , \h2_pad , \h3_pad , \h4_pad , h_pad, \i0_pad , \i1_pad , \i2_pad , \i3_pad , i_pad, \j0_pad , \j1_pad , \j2_pad , \j3_pad , j_pad, \k0_pad , \k1_pad , \k2_pad , \k3_pad , k_pad, \l0_pad , \l1_pad , \l2_pad , \l3_pad , l_pad, \m0_pad , \m1_pad , \m2_pad , \m3_pad , m_pad, \n0_pad , \n1_pad , \n2_pad , \n3_pad , n_pad, \o0_pad , \o1_pad , \o2_pad , \o3_pad , o_pad, \p1_pad , \p2_pad , \p3_pad , p_pad, \q1_pad , \q2_pad , \q3_pad , q_pad, \r0_pad , \r1_pad , \r2_pad , \r3_pad , r_pad, \s0_pad , \s1_pad , \s2_pad , \s3_pad , s_pad, \t0_pad , \t1_pad , \t2_pad , \t3_pad , t_pad, \u0_pad , \u1_pad , \u2_pad , \u3_pad , u_pad, \v0_pad , \v1_pad , \v2_pad , \v3_pad , v_pad, \w0_pad , \w1_pad , \w2_pad , \w3_pad , w_pad, \x0_pad , \x1_pad , \x2_pad , \x3_pad , x_pad, \y0_pad , \y1_pad , \y2_pad , \y3_pad , y_pad, \z0_pad , \z1_pad , \z2_pad , \z3_pad , z_pad, \a5_pad , \a6_pad , \a7_pad , \a8_pad , \b5_pad , \b6_pad , \b7_pad , \b8_pad , \c5_pad , \c6_pad , \c7_pad , \c8_pad , \d5_pad , \d6_pad , \d7_pad , \e5_pad , \e6_pad , \e7_pad , \f5_pad , \f6_pad , \f7_pad , \g5_pad , \g6_pad , \g7_pad , \h5_pad , \h6_pad , \h7_pad , \i4_pad , \i5_pad , \i6_pad , \i7_pad , \j4_pad , \j5_pad , \j6_pad , \j7_pad , \k4_pad , \k5_pad , \k6_pad , \k7_pad , \l4_pad , \l5_pad , \l6_pad , \l7_pad , \m4_pad , \m5_pad , \m6_pad , \m7_pad , \n4_pad , \n5_pad , \n6_pad , \n7_pad , \o4_pad , \o5_pad , \o6_pad , \o7_pad , \p4_pad , \p5_pad , \p6_pad , \p7_pad , \q4_pad , \q5_pad , \q6_pad , \q7_pad , \r4_pad , \r5_pad , \r6_pad , \r7_pad , \s4_pad , \s5_pad , \s6_pad , \s7_pad , \t4_pad , \t5_pad , \t6_pad , \t7_pad , \u4_pad , \u5_pad , \u6_pad , \u7_pad , \v4_pad , \v5_pad , \v6_pad , \v7_pad , \w4_pad , \w5_pad , \w6_pad , \w7_pad , \x4_pad , \x5_pad , \x6_pad , \x7_pad , \y4_pad , \y5_pad , \y6_pad , \y7_pad , \z4_pad , \z5_pad , \z6_pad , \z7_pad );
	input \a0_pad  ;
	input \a1_pad  ;
	input \a2_pad  ;
	input \a3_pad  ;
	input \a4_pad  ;
	input \b0_pad  ;
	input \b1_pad  ;
	input \b2_pad  ;
	input \b3_pad  ;
	input \b4_pad  ;
	input b_pad ;
	input \c0_pad  ;
	input \c1_pad  ;
	input \c2_pad  ;
	input \c3_pad  ;
	input \c4_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input \d1_pad  ;
	input \d2_pad  ;
	input \d3_pad  ;
	input \d4_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input \e1_pad  ;
	input \e2_pad  ;
	input \e3_pad  ;
	input \e4_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input \f1_pad  ;
	input \f2_pad  ;
	input \f3_pad  ;
	input \f4_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input \g1_pad  ;
	input \g2_pad  ;
	input \g3_pad  ;
	input \g4_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input \h1_pad  ;
	input \h2_pad  ;
	input \h3_pad  ;
	input \h4_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input \i1_pad  ;
	input \i2_pad  ;
	input \i3_pad  ;
	input i_pad ;
	input \j0_pad  ;
	input \j1_pad  ;
	input \j2_pad  ;
	input \j3_pad  ;
	input j_pad ;
	input \k0_pad  ;
	input \k1_pad  ;
	input \k2_pad  ;
	input \k3_pad  ;
	input k_pad ;
	input \l0_pad  ;
	input \l1_pad  ;
	input \l2_pad  ;
	input \l3_pad  ;
	input l_pad ;
	input \m0_pad  ;
	input \m1_pad  ;
	input \m2_pad  ;
	input \m3_pad  ;
	input m_pad ;
	input \n0_pad  ;
	input \n1_pad  ;
	input \n2_pad  ;
	input \n3_pad  ;
	input n_pad ;
	input \o0_pad  ;
	input \o1_pad  ;
	input \o2_pad  ;
	input \o3_pad  ;
	input o_pad ;
	input \p1_pad  ;
	input \p2_pad  ;
	input \p3_pad  ;
	input p_pad ;
	input \q1_pad  ;
	input \q2_pad  ;
	input \q3_pad  ;
	input q_pad ;
	input \r0_pad  ;
	input \r1_pad  ;
	input \r2_pad  ;
	input \r3_pad  ;
	input r_pad ;
	input \s0_pad  ;
	input \s1_pad  ;
	input \s2_pad  ;
	input \s3_pad  ;
	input s_pad ;
	input \t0_pad  ;
	input \t1_pad  ;
	input \t2_pad  ;
	input \t3_pad  ;
	input t_pad ;
	input \u0_pad  ;
	input \u1_pad  ;
	input \u2_pad  ;
	input \u3_pad  ;
	input u_pad ;
	input \v0_pad  ;
	input \v1_pad  ;
	input \v2_pad  ;
	input \v3_pad  ;
	input v_pad ;
	input \w0_pad  ;
	input \w1_pad  ;
	input \w2_pad  ;
	input \w3_pad  ;
	input w_pad ;
	input \x0_pad  ;
	input \x1_pad  ;
	input \x2_pad  ;
	input \x3_pad  ;
	input x_pad ;
	input \y0_pad  ;
	input \y1_pad  ;
	input \y2_pad  ;
	input \y3_pad  ;
	input y_pad ;
	input \z0_pad  ;
	input \z1_pad  ;
	input \z2_pad  ;
	input \z3_pad  ;
	input z_pad ;
	output \a5_pad  ;
	output \a6_pad  ;
	output \a7_pad  ;
	output \a8_pad  ;
	output \b5_pad  ;
	output \b6_pad  ;
	output \b7_pad  ;
	output \b8_pad  ;
	output \c5_pad  ;
	output \c6_pad  ;
	output \c7_pad  ;
	output \c8_pad  ;
	output \d5_pad  ;
	output \d6_pad  ;
	output \d7_pad  ;
	output \e5_pad  ;
	output \e6_pad  ;
	output \e7_pad  ;
	output \f5_pad  ;
	output \f6_pad  ;
	output \f7_pad  ;
	output \g5_pad  ;
	output \g6_pad  ;
	output \g7_pad  ;
	output \h5_pad  ;
	output \h6_pad  ;
	output \h7_pad  ;
	output \i4_pad  ;
	output \i5_pad  ;
	output \i6_pad  ;
	output \i7_pad  ;
	output \j4_pad  ;
	output \j5_pad  ;
	output \j6_pad  ;
	output \j7_pad  ;
	output \k4_pad  ;
	output \k5_pad  ;
	output \k6_pad  ;
	output \k7_pad  ;
	output \l4_pad  ;
	output \l5_pad  ;
	output \l6_pad  ;
	output \l7_pad  ;
	output \m4_pad  ;
	output \m5_pad  ;
	output \m6_pad  ;
	output \m7_pad  ;
	output \n4_pad  ;
	output \n5_pad  ;
	output \n6_pad  ;
	output \n7_pad  ;
	output \o4_pad  ;
	output \o5_pad  ;
	output \o6_pad  ;
	output \o7_pad  ;
	output \p4_pad  ;
	output \p5_pad  ;
	output \p6_pad  ;
	output \p7_pad  ;
	output \q4_pad  ;
	output \q5_pad  ;
	output \q6_pad  ;
	output \q7_pad  ;
	output \r4_pad  ;
	output \r5_pad  ;
	output \r6_pad  ;
	output \r7_pad  ;
	output \s4_pad  ;
	output \s5_pad  ;
	output \s6_pad  ;
	output \s7_pad  ;
	output \t4_pad  ;
	output \t5_pad  ;
	output \t6_pad  ;
	output \t7_pad  ;
	output \u4_pad  ;
	output \u5_pad  ;
	output \u6_pad  ;
	output \u7_pad  ;
	output \v4_pad  ;
	output \v5_pad  ;
	output \v6_pad  ;
	output \v7_pad  ;
	output \w4_pad  ;
	output \w5_pad  ;
	output \w6_pad  ;
	output \w7_pad  ;
	output \x4_pad  ;
	output \x5_pad  ;
	output \x6_pad  ;
	output \x7_pad  ;
	output \y4_pad  ;
	output \y5_pad  ;
	output \y6_pad  ;
	output \y7_pad  ;
	output \z4_pad  ;
	output \z5_pad  ;
	output \z6_pad  ;
	output \z7_pad  ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w256_ ;
	wire _w255_ ;
	wire _w254_ ;
	wire _w253_ ;
	wire _w252_ ;
	wire _w251_ ;
	wire _w250_ ;
	wire _w249_ ;
	wire _w248_ ;
	wire _w247_ ;
	wire _w246_ ;
	wire _w245_ ;
	wire _w244_ ;
	wire _w243_ ;
	wire _w242_ ;
	wire _w241_ ;
	wire _w240_ ;
	wire _w239_ ;
	wire _w238_ ;
	wire _w237_ ;
	wire _w236_ ;
	wire _w235_ ;
	wire _w234_ ;
	wire _w233_ ;
	wire _w232_ ;
	wire _w231_ ;
	wire _w230_ ;
	wire _w229_ ;
	wire _w228_ ;
	wire _w227_ ;
	wire _w226_ ;
	wire _w225_ ;
	wire _w224_ ;
	wire _w223_ ;
	wire _w222_ ;
	wire _w221_ ;
	wire _w220_ ;
	wire _w219_ ;
	wire _w218_ ;
	wire _w217_ ;
	wire _w216_ ;
	wire _w215_ ;
	wire _w214_ ;
	wire _w213_ ;
	wire _w212_ ;
	wire _w211_ ;
	wire _w210_ ;
	wire _w209_ ;
	wire _w208_ ;
	wire _w207_ ;
	wire _w206_ ;
	wire _w205_ ;
	wire _w204_ ;
	wire _w203_ ;
	wire _w202_ ;
	wire _w201_ ;
	wire _w200_ ;
	wire _w199_ ;
	wire _w198_ ;
	wire _w197_ ;
	wire _w196_ ;
	wire _w165_ ;
	wire _w164_ ;
	wire _w163_ ;
	wire _w162_ ;
	wire _w161_ ;
	wire _w160_ ;
	wire _w159_ ;
	wire _w158_ ;
	wire _w157_ ;
	wire _w156_ ;
	wire _w155_ ;
	wire _w154_ ;
	wire _w153_ ;
	wire _w152_ ;
	wire _w151_ ;
	wire _w150_ ;
	wire _w137_ ;
	wire _w138_ ;
	wire _w139_ ;
	wire _w140_ ;
	wire _w141_ ;
	wire _w142_ ;
	wire _w143_ ;
	wire _w144_ ;
	wire _w145_ ;
	wire _w146_ ;
	wire _w147_ ;
	wire _w148_ ;
	wire _w149_ ;
	wire _w166_ ;
	wire _w167_ ;
	wire _w168_ ;
	wire _w169_ ;
	wire _w170_ ;
	wire _w171_ ;
	wire _w172_ ;
	wire _w173_ ;
	wire _w174_ ;
	wire _w175_ ;
	wire _w176_ ;
	wire _w177_ ;
	wire _w178_ ;
	wire _w179_ ;
	wire _w180_ ;
	wire _w181_ ;
	wire _w182_ ;
	wire _w183_ ;
	wire _w184_ ;
	wire _w185_ ;
	wire _w186_ ;
	wire _w187_ ;
	wire _w188_ ;
	wire _w189_ ;
	wire _w190_ ;
	wire _w191_ ;
	wire _w192_ ;
	wire _w193_ ;
	wire _w194_ ;
	wire _w195_ ;
	wire _w264_ ;
	wire _w265_ ;
	wire _w266_ ;
	wire _w267_ ;
	wire _w268_ ;
	wire _w269_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w286_ ;
	wire _w287_ ;
	wire _w288_ ;
	wire _w289_ ;
	wire _w290_ ;
	wire _w291_ ;
	wire _w292_ ;
	wire _w293_ ;
	wire _w294_ ;
	wire _w295_ ;
	wire _w296_ ;
	wire _w297_ ;
	wire _w298_ ;
	wire _w299_ ;
	wire _w300_ ;
	wire _w301_ ;
	wire _w302_ ;
	wire _w303_ ;
	wire _w304_ ;
	wire _w305_ ;
	wire _w306_ ;
	wire _w307_ ;
	wire _w308_ ;
	wire _w309_ ;
	wire _w310_ ;
	wire _w311_ ;
	wire _w312_ ;
	wire _w313_ ;
	wire _w314_ ;
	wire _w315_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w384_ ;
	wire _w385_ ;
	wire _w386_ ;
	wire _w387_ ;
	wire _w388_ ;
	wire _w389_ ;
	wire _w390_ ;
	wire _w391_ ;
	wire _w392_ ;
	wire _w393_ ;
	LUT3 #(
		.INIT('h20)
	) name0 (
		i_pad,
		p_pad,
		r_pad,
		_w137_
	);
	LUT4 #(
		.INIT('h00ea)
	) name1 (
		\f1_pad ,
		i_pad,
		r_pad,
		\y1_pad ,
		_w138_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		_w137_,
		_w138_,
		_w139_
	);
	LUT3 #(
		.INIT('h80)
	) name3 (
		\a4_pad ,
		\y3_pad ,
		\z3_pad ,
		_w140_
	);
	LUT4 #(
		.INIT('h8000)
	) name4 (
		\a4_pad ,
		\b4_pad ,
		\y3_pad ,
		\z3_pad ,
		_w141_
	);
	LUT2 #(
		.INIT('h8)
	) name5 (
		\c4_pad ,
		_w141_,
		_w142_
	);
	LUT4 #(
		.INIT('h485a)
	) name6 (
		\d4_pad ,
		\f4_pad ,
		\h0_pad ,
		\j0_pad ,
		_w143_
	);
	LUT2 #(
		.INIT('h6)
	) name7 (
		\g4_pad ,
		\k0_pad ,
		_w144_
	);
	LUT2 #(
		.INIT('h6)
	) name8 (
		\e4_pad ,
		\i0_pad ,
		_w145_
	);
	LUT3 #(
		.INIT('hc4)
	) name9 (
		\f4_pad ,
		\h4_pad ,
		\j0_pad ,
		_w146_
	);
	LUT4 #(
		.INIT('h1000)
	) name10 (
		_w145_,
		_w144_,
		_w146_,
		_w143_,
		_w147_
	);
	LUT2 #(
		.INIT('h8)
	) name11 (
		\d2_pad ,
		\l0_pad ,
		_w148_
	);
	LUT4 #(
		.INIT('h0001)
	) name12 (
		\h0_pad ,
		\i0_pad ,
		\j0_pad ,
		\k0_pad ,
		_w149_
	);
	LUT2 #(
		.INIT('h8)
	) name13 (
		_w148_,
		_w149_,
		_w150_
	);
	LUT4 #(
		.INIT('h0015)
	) name14 (
		\a2_pad ,
		_w142_,
		_w147_,
		_w150_,
		_w151_
	);
	LUT4 #(
		.INIT('h0c06)
	) name15 (
		\e2_pad ,
		\f2_pad ,
		\n0_pad ,
		_w151_,
		_w152_
	);
	LUT3 #(
		.INIT('h20)
	) name16 (
		f_pad,
		\g3_pad ,
		h_pad,
		_w153_
	);
	LUT4 #(
		.INIT('h00ea)
	) name17 (
		\f3_pad ,
		f_pad,
		h_pad,
		\y1_pad ,
		_w154_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		_w153_,
		_w154_,
		_w155_
	);
	LUT3 #(
		.INIT('h20)
	) name19 (
		\c4_pad ,
		\d4_pad ,
		_w141_,
		_w156_
	);
	LUT4 #(
		.INIT('h2000)
	) name20 (
		\c4_pad ,
		\d4_pad ,
		\e4_pad ,
		_w141_,
		_w157_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		\l0_pad ,
		\n0_pad ,
		_w158_
	);
	LUT3 #(
		.INIT('h48)
	) name22 (
		\f4_pad ,
		_w158_,
		_w157_,
		_w159_
	);
	LUT3 #(
		.INIT('h20)
	) name23 (
		i_pad,
		q_pad,
		r_pad,
		_w160_
	);
	LUT4 #(
		.INIT('h00ea)
	) name24 (
		\g1_pad ,
		i_pad,
		r_pad,
		\y1_pad ,
		_w161_
	);
	LUT2 #(
		.INIT('h4)
	) name25 (
		_w160_,
		_w161_,
		_w162_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\h2_pad ,
		\n0_pad ,
		_w163_
	);
	LUT3 #(
		.INIT('h20)
	) name27 (
		f_pad,
		\h3_pad ,
		h_pad,
		_w164_
	);
	LUT4 #(
		.INIT('h00ec)
	) name28 (
		f_pad,
		\g3_pad ,
		h_pad,
		\y1_pad ,
		_w165_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		_w164_,
		_w165_,
		_w166_
	);
	LUT4 #(
		.INIT('h60c0)
	) name30 (
		\f4_pad ,
		\g4_pad ,
		_w158_,
		_w157_,
		_w167_
	);
	LUT3 #(
		.INIT('h04)
	) name31 (
		\b0_pad ,
		s_pad,
		t_pad,
		_w168_
	);
	LUT4 #(
		.INIT('h00dc)
	) name32 (
		\b0_pad ,
		\h1_pad ,
		s_pad,
		\y1_pad ,
		_w169_
	);
	LUT2 #(
		.INIT('h4)
	) name33 (
		_w168_,
		_w169_,
		_w170_
	);
	LUT2 #(
		.INIT('h2)
	) name34 (
		\l0_pad ,
		\n0_pad ,
		_w171_
	);
	LUT3 #(
		.INIT('h20)
	) name35 (
		f_pad,
		g_pad,
		h_pad,
		_w172_
	);
	LUT4 #(
		.INIT('h00ec)
	) name36 (
		f_pad,
		\h3_pad ,
		h_pad,
		\y1_pad ,
		_w173_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		_w172_,
		_w173_,
		_w174_
	);
	LUT3 #(
		.INIT('h13)
	) name38 (
		\d2_pad ,
		\h4_pad ,
		\l0_pad ,
		_w175_
	);
	LUT4 #(
		.INIT('h002a)
	) name39 (
		b_pad,
		\g2_pad ,
		\h2_pad ,
		\n0_pad ,
		_w176_
	);
	LUT2 #(
		.INIT('h4)
	) name40 (
		_w175_,
		_w176_,
		_w177_
	);
	LUT3 #(
		.INIT('h04)
	) name41 (
		\b0_pad ,
		s_pad,
		u_pad,
		_w178_
	);
	LUT4 #(
		.INIT('h00dc)
	) name42 (
		\b0_pad ,
		\i1_pad ,
		s_pad,
		\y1_pad ,
		_w179_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w178_,
		_w179_,
		_w180_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		\o2_pad ,
		\p2_pad ,
		_w181_
	);
	LUT3 #(
		.INIT('h02)
	) name45 (
		\g0_pad ,
		\o2_pad ,
		\p2_pad ,
		_w182_
	);
	LUT3 #(
		.INIT('hc4)
	) name46 (
		\j2_pad ,
		\o2_pad ,
		\p2_pad ,
		_w183_
	);
	LUT3 #(
		.INIT('h20)
	) name47 (
		\l2_pad ,
		\m2_pad ,
		\n2_pad ,
		_w184_
	);
	LUT4 #(
		.INIT('h0010)
	) name48 (
		\x1_pad ,
		_w183_,
		_w184_,
		_w182_,
		_w185_
	);
	LUT3 #(
		.INIT('h32)
	) name49 (
		\i2_pad ,
		\y1_pad ,
		_w185_,
		_w186_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		\j2_pad ,
		\k2_pad ,
		_w187_
	);
	LUT4 #(
		.INIT('haa02)
	) name51 (
		\i3_pad ,
		\j2_pad ,
		\k2_pad ,
		\x1_pad ,
		_w188_
	);
	LUT4 #(
		.INIT('h00c8)
	) name52 (
		\j2_pad ,
		\j3_pad ,
		\k2_pad ,
		\x1_pad ,
		_w189_
	);
	LUT3 #(
		.INIT('h01)
	) name53 (
		c_pad,
		d_pad,
		e_pad,
		_w190_
	);
	LUT3 #(
		.INIT('h04)
	) name54 (
		_w189_,
		_w190_,
		_w188_,
		_w191_
	);
	LUT4 #(
		.INIT('h0002)
	) name55 (
		c_pad,
		d_pad,
		e_pad,
		\s2_pad ,
		_w192_
	);
	LUT3 #(
		.INIT('h02)
	) name56 (
		d_pad,
		e_pad,
		\r0_pad ,
		_w193_
	);
	LUT3 #(
		.INIT('h0d)
	) name57 (
		e_pad,
		\h1_pad ,
		\y1_pad ,
		_w194_
	);
	LUT3 #(
		.INIT('h10)
	) name58 (
		_w193_,
		_w192_,
		_w194_,
		_w195_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		_w191_,
		_w195_,
		_w196_
	);
	LUT3 #(
		.INIT('h04)
	) name60 (
		\b0_pad ,
		s_pad,
		v_pad,
		_w197_
	);
	LUT4 #(
		.INIT('h00dc)
	) name61 (
		\b0_pad ,
		\j1_pad ,
		s_pad,
		\y1_pad ,
		_w198_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w197_,
		_w198_,
		_w199_
	);
	LUT4 #(
		.INIT('h001f)
	) name63 (
		\e0_pad ,
		\f0_pad ,
		\g0_pad ,
		\o2_pad ,
		_w200_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		\p2_pad ,
		\x1_pad ,
		_w201_
	);
	LUT4 #(
		.INIT('h5155)
	) name65 (
		\j2_pad ,
		_w184_,
		_w200_,
		_w201_,
		_w202_
	);
	LUT2 #(
		.INIT('h1)
	) name66 (
		\j2_pad ,
		\o2_pad ,
		_w203_
	);
	LUT4 #(
		.INIT('h0200)
	) name67 (
		_w184_,
		_w203_,
		_w200_,
		_w201_,
		_w204_
	);
	LUT3 #(
		.INIT('h01)
	) name68 (
		\y1_pad ,
		_w204_,
		_w202_,
		_w205_
	);
	LUT4 #(
		.INIT('hcc04)
	) name69 (
		\j2_pad ,
		\j3_pad ,
		\k2_pad ,
		\x1_pad ,
		_w206_
	);
	LUT4 #(
		.INIT('h00e0)
	) name70 (
		\j2_pad ,
		\k2_pad ,
		\k3_pad ,
		\x1_pad ,
		_w207_
	);
	LUT3 #(
		.INIT('h02)
	) name71 (
		_w190_,
		_w207_,
		_w206_,
		_w208_
	);
	LUT4 #(
		.INIT('h0002)
	) name72 (
		c_pad,
		d_pad,
		e_pad,
		\t2_pad ,
		_w209_
	);
	LUT3 #(
		.INIT('h02)
	) name73 (
		d_pad,
		e_pad,
		\s0_pad ,
		_w210_
	);
	LUT3 #(
		.INIT('h0d)
	) name74 (
		e_pad,
		\i1_pad ,
		\y1_pad ,
		_w211_
	);
	LUT3 #(
		.INIT('h10)
	) name75 (
		_w210_,
		_w209_,
		_w211_,
		_w212_
	);
	LUT2 #(
		.INIT('h4)
	) name76 (
		_w208_,
		_w212_,
		_w213_
	);
	LUT3 #(
		.INIT('h04)
	) name77 (
		\b0_pad ,
		s_pad,
		w_pad,
		_w214_
	);
	LUT4 #(
		.INIT('h00dc)
	) name78 (
		\b0_pad ,
		\k1_pad ,
		s_pad,
		\y1_pad ,
		_w215_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		_w214_,
		_w215_,
		_w216_
	);
	LUT4 #(
		.INIT('h00ef)
	) name80 (
		\e0_pad ,
		\f0_pad ,
		\g0_pad ,
		\p2_pad ,
		_w217_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\o2_pad ,
		\x1_pad ,
		_w218_
	);
	LUT3 #(
		.INIT('h20)
	) name82 (
		_w184_,
		_w217_,
		_w218_,
		_w219_
	);
	LUT3 #(
		.INIT('h12)
	) name83 (
		\k2_pad ,
		\y1_pad ,
		_w219_,
		_w220_
	);
	LUT4 #(
		.INIT('hf010)
	) name84 (
		\j2_pad ,
		\k2_pad ,
		\k3_pad ,
		\x1_pad ,
		_w221_
	);
	LUT4 #(
		.INIT('h00e0)
	) name85 (
		\j2_pad ,
		\k2_pad ,
		\l3_pad ,
		\x1_pad ,
		_w222_
	);
	LUT3 #(
		.INIT('h02)
	) name86 (
		_w190_,
		_w222_,
		_w221_,
		_w223_
	);
	LUT4 #(
		.INIT('h0002)
	) name87 (
		c_pad,
		d_pad,
		e_pad,
		\u2_pad ,
		_w224_
	);
	LUT3 #(
		.INIT('h02)
	) name88 (
		d_pad,
		e_pad,
		\t0_pad ,
		_w225_
	);
	LUT3 #(
		.INIT('h0d)
	) name89 (
		e_pad,
		\j1_pad ,
		\y1_pad ,
		_w226_
	);
	LUT3 #(
		.INIT('h10)
	) name90 (
		_w225_,
		_w224_,
		_w226_,
		_w227_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w223_,
		_w227_,
		_w228_
	);
	LUT3 #(
		.INIT('h04)
	) name92 (
		\b0_pad ,
		s_pad,
		x_pad,
		_w229_
	);
	LUT4 #(
		.INIT('h00dc)
	) name93 (
		\b0_pad ,
		\l1_pad ,
		s_pad,
		\y1_pad ,
		_w230_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w229_,
		_w230_,
		_w231_
	);
	LUT4 #(
		.INIT('h0100)
	) name95 (
		c_pad,
		d_pad,
		e_pad,
		\x1_pad ,
		_w232_
	);
	LUT3 #(
		.INIT('h21)
	) name96 (
		\l2_pad ,
		\y1_pad ,
		_w232_,
		_w233_
	);
	LUT4 #(
		.INIT('hf010)
	) name97 (
		\j2_pad ,
		\k2_pad ,
		\l3_pad ,
		\x1_pad ,
		_w234_
	);
	LUT4 #(
		.INIT('h00e0)
	) name98 (
		\j2_pad ,
		\k2_pad ,
		\m3_pad ,
		\x1_pad ,
		_w235_
	);
	LUT3 #(
		.INIT('h02)
	) name99 (
		_w190_,
		_w235_,
		_w234_,
		_w236_
	);
	LUT4 #(
		.INIT('h0002)
	) name100 (
		c_pad,
		d_pad,
		e_pad,
		\v2_pad ,
		_w237_
	);
	LUT3 #(
		.INIT('h02)
	) name101 (
		d_pad,
		e_pad,
		\u0_pad ,
		_w238_
	);
	LUT3 #(
		.INIT('h0d)
	) name102 (
		e_pad,
		\k1_pad ,
		\y1_pad ,
		_w239_
	);
	LUT3 #(
		.INIT('h10)
	) name103 (
		_w238_,
		_w237_,
		_w239_,
		_w240_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w236_,
		_w240_,
		_w241_
	);
	LUT3 #(
		.INIT('h04)
	) name105 (
		\b0_pad ,
		s_pad,
		y_pad,
		_w242_
	);
	LUT4 #(
		.INIT('h00dc)
	) name106 (
		\b0_pad ,
		\m1_pad ,
		s_pad,
		\y1_pad ,
		_w243_
	);
	LUT2 #(
		.INIT('h4)
	) name107 (
		_w242_,
		_w243_,
		_w244_
	);
	LUT3 #(
		.INIT('h08)
	) name108 (
		\l2_pad ,
		\m2_pad ,
		_w232_,
		_w245_
	);
	LUT4 #(
		.INIT('h0c06)
	) name109 (
		\l2_pad ,
		\m2_pad ,
		\y1_pad ,
		_w232_,
		_w246_
	);
	LUT4 #(
		.INIT('hf010)
	) name110 (
		\j2_pad ,
		\k2_pad ,
		\m3_pad ,
		\x1_pad ,
		_w247_
	);
	LUT4 #(
		.INIT('h00e0)
	) name111 (
		\j2_pad ,
		\k2_pad ,
		\n3_pad ,
		\x1_pad ,
		_w248_
	);
	LUT3 #(
		.INIT('h02)
	) name112 (
		_w190_,
		_w248_,
		_w247_,
		_w249_
	);
	LUT4 #(
		.INIT('h0002)
	) name113 (
		c_pad,
		d_pad,
		e_pad,
		\w2_pad ,
		_w250_
	);
	LUT3 #(
		.INIT('h02)
	) name114 (
		d_pad,
		e_pad,
		\v0_pad ,
		_w251_
	);
	LUT3 #(
		.INIT('h0d)
	) name115 (
		e_pad,
		\l1_pad ,
		\y1_pad ,
		_w252_
	);
	LUT3 #(
		.INIT('h10)
	) name116 (
		_w251_,
		_w250_,
		_w252_,
		_w253_
	);
	LUT2 #(
		.INIT('h4)
	) name117 (
		_w249_,
		_w253_,
		_w254_
	);
	LUT2 #(
		.INIT('hb)
	) name118 (
		\a2_pad ,
		\x1_pad ,
		_w255_
	);
	LUT3 #(
		.INIT('h04)
	) name119 (
		\b0_pad ,
		s_pad,
		z_pad,
		_w256_
	);
	LUT4 #(
		.INIT('h00dc)
	) name120 (
		\b0_pad ,
		\n1_pad ,
		s_pad,
		\y1_pad ,
		_w257_
	);
	LUT2 #(
		.INIT('h4)
	) name121 (
		_w256_,
		_w257_,
		_w258_
	);
	LUT4 #(
		.INIT('h0080)
	) name122 (
		\l2_pad ,
		\m2_pad ,
		\n2_pad ,
		_w232_,
		_w259_
	);
	LUT3 #(
		.INIT('h12)
	) name123 (
		\n2_pad ,
		\y1_pad ,
		_w245_,
		_w260_
	);
	LUT4 #(
		.INIT('hf010)
	) name124 (
		\j2_pad ,
		\k2_pad ,
		\n3_pad ,
		\x1_pad ,
		_w261_
	);
	LUT4 #(
		.INIT('h00e0)
	) name125 (
		\j2_pad ,
		\k2_pad ,
		\o3_pad ,
		\x1_pad ,
		_w262_
	);
	LUT3 #(
		.INIT('h02)
	) name126 (
		_w190_,
		_w262_,
		_w261_,
		_w263_
	);
	LUT4 #(
		.INIT('h0002)
	) name127 (
		c_pad,
		d_pad,
		e_pad,
		\x2_pad ,
		_w264_
	);
	LUT3 #(
		.INIT('h02)
	) name128 (
		d_pad,
		e_pad,
		\w0_pad ,
		_w265_
	);
	LUT3 #(
		.INIT('h0d)
	) name129 (
		e_pad,
		\m1_pad ,
		\y1_pad ,
		_w266_
	);
	LUT3 #(
		.INIT('h10)
	) name130 (
		_w265_,
		_w264_,
		_w266_,
		_w267_
	);
	LUT2 #(
		.INIT('h4)
	) name131 (
		_w263_,
		_w267_,
		_w268_
	);
	LUT4 #(
		.INIT('h0080)
	) name132 (
		\i2_pad ,
		\q2_pad ,
		\r2_pad ,
		\x1_pad ,
		_w269_
	);
	LUT4 #(
		.INIT('hfcec)
	) name133 (
		\o0_pad ,
		\y1_pad ,
		_w190_,
		_w269_,
		_w270_
	);
	LUT3 #(
		.INIT('h10)
	) name134 (
		\a0_pad ,
		\b0_pad ,
		s_pad,
		_w271_
	);
	LUT4 #(
		.INIT('h00dc)
	) name135 (
		\b0_pad ,
		\o1_pad ,
		s_pad,
		\y1_pad ,
		_w272_
	);
	LUT2 #(
		.INIT('h4)
	) name136 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT3 #(
		.INIT('h12)
	) name137 (
		\o2_pad ,
		\y1_pad ,
		_w259_,
		_w274_
	);
	LUT4 #(
		.INIT('hf010)
	) name138 (
		\j2_pad ,
		\k2_pad ,
		\o3_pad ,
		\x1_pad ,
		_w275_
	);
	LUT4 #(
		.INIT('h00e0)
	) name139 (
		\j2_pad ,
		\k2_pad ,
		\p3_pad ,
		\x1_pad ,
		_w276_
	);
	LUT3 #(
		.INIT('h02)
	) name140 (
		_w190_,
		_w276_,
		_w275_,
		_w277_
	);
	LUT4 #(
		.INIT('h0002)
	) name141 (
		c_pad,
		d_pad,
		e_pad,
		\y2_pad ,
		_w278_
	);
	LUT3 #(
		.INIT('h02)
	) name142 (
		d_pad,
		e_pad,
		\x0_pad ,
		_w279_
	);
	LUT3 #(
		.INIT('h0d)
	) name143 (
		e_pad,
		\n1_pad ,
		\y1_pad ,
		_w280_
	);
	LUT3 #(
		.INIT('h10)
	) name144 (
		_w279_,
		_w278_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h4)
	) name145 (
		_w277_,
		_w281_,
		_w282_
	);
	LUT3 #(
		.INIT('ha8)
	) name146 (
		\i2_pad ,
		\q2_pad ,
		\r2_pad ,
		_w283_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		_w187_,
		_w283_,
		_w284_
	);
	LUT3 #(
		.INIT('h51)
	) name148 (
		\x1_pad ,
		_w187_,
		_w283_,
		_w285_
	);
	LUT4 #(
		.INIT('h00ac)
	) name149 (
		\j0_pad ,
		\k0_pad ,
		\l2_pad ,
		\n2_pad ,
		_w286_
	);
	LUT4 #(
		.INIT('hac00)
	) name150 (
		\h0_pad ,
		\i0_pad ,
		\l2_pad ,
		\n2_pad ,
		_w287_
	);
	LUT4 #(
		.INIT('hc840)
	) name151 (
		\m2_pad ,
		_w181_,
		_w287_,
		_w286_,
		_w288_
	);
	LUT4 #(
		.INIT('hc8c0)
	) name152 (
		\d0_pad ,
		\i2_pad ,
		\q2_pad ,
		\r2_pad ,
		_w289_
	);
	LUT3 #(
		.INIT('h4c)
	) name153 (
		\i2_pad ,
		\i3_pad ,
		\r2_pad ,
		_w290_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		\c0_pad ,
		\r2_pad ,
		_w291_
	);
	LUT4 #(
		.INIT('h8808)
	) name155 (
		\i2_pad ,
		\q2_pad ,
		\r2_pad ,
		\z1_pad ,
		_w292_
	);
	LUT4 #(
		.INIT('he0ee)
	) name156 (
		_w289_,
		_w290_,
		_w291_,
		_w292_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		\a2_pad ,
		\y1_pad ,
		_w294_
	);
	LUT4 #(
		.INIT('hd800)
	) name158 (
		_w285_,
		_w293_,
		_w288_,
		_w294_,
		_w295_
	);
	LUT3 #(
		.INIT('h2a)
	) name159 (
		\a2_pad ,
		\e2_pad ,
		\f2_pad ,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		\d0_pad ,
		\e2_pad ,
		_w297_
	);
	LUT4 #(
		.INIT('h00d0)
	) name161 (
		\d0_pad ,
		\f2_pad ,
		\m0_pad ,
		\y1_pad ,
		_w298_
	);
	LUT3 #(
		.INIT('h20)
	) name162 (
		_w296_,
		_w297_,
		_w298_,
		_w299_
	);
	LUT2 #(
		.INIT('he)
	) name163 (
		_w295_,
		_w299_,
		_w300_
	);
	LUT3 #(
		.INIT('h08)
	) name164 (
		\b0_pad ,
		s_pad,
		t_pad,
		_w301_
	);
	LUT4 #(
		.INIT('h00ec)
	) name165 (
		\b0_pad ,
		\p1_pad ,
		s_pad,
		\y1_pad ,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		_w301_,
		_w302_,
		_w303_
	);
	LUT4 #(
		.INIT('h060c)
	) name167 (
		\o2_pad ,
		\p2_pad ,
		\y1_pad ,
		_w259_,
		_w304_
	);
	LUT4 #(
		.INIT('hf010)
	) name168 (
		\j2_pad ,
		\k2_pad ,
		\p3_pad ,
		\x1_pad ,
		_w305_
	);
	LUT4 #(
		.INIT('h00e0)
	) name169 (
		\j2_pad ,
		\k2_pad ,
		\q3_pad ,
		\x1_pad ,
		_w306_
	);
	LUT3 #(
		.INIT('h02)
	) name170 (
		_w190_,
		_w306_,
		_w305_,
		_w307_
	);
	LUT4 #(
		.INIT('h0002)
	) name171 (
		c_pad,
		d_pad,
		e_pad,
		\z2_pad ,
		_w308_
	);
	LUT3 #(
		.INIT('h02)
	) name172 (
		d_pad,
		e_pad,
		\y0_pad ,
		_w309_
	);
	LUT3 #(
		.INIT('h0d)
	) name173 (
		e_pad,
		\o1_pad ,
		\y1_pad ,
		_w310_
	);
	LUT3 #(
		.INIT('h10)
	) name174 (
		_w309_,
		_w308_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h4)
	) name175 (
		_w307_,
		_w311_,
		_w312_
	);
	LUT4 #(
		.INIT('h00ea)
	) name176 (
		\c2_pad ,
		\g2_pad ,
		\h2_pad ,
		\n0_pad ,
		_w313_
	);
	LUT3 #(
		.INIT('h08)
	) name177 (
		\b0_pad ,
		s_pad,
		u_pad,
		_w314_
	);
	LUT4 #(
		.INIT('h00ec)
	) name178 (
		\b0_pad ,
		\q1_pad ,
		s_pad,
		\y1_pad ,
		_w315_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT4 #(
		.INIT('h5545)
	) name180 (
		\i2_pad ,
		_w183_,
		_w184_,
		_w182_,
		_w317_
	);
	LUT3 #(
		.INIT('h02)
	) name181 (
		\q2_pad ,
		\x1_pad ,
		_w317_,
		_w318_
	);
	LUT4 #(
		.INIT('h0a09)
	) name182 (
		\q2_pad ,
		\x1_pad ,
		\y1_pad ,
		_w317_,
		_w319_
	);
	LUT4 #(
		.INIT('hf010)
	) name183 (
		\j2_pad ,
		\k2_pad ,
		\q3_pad ,
		\x1_pad ,
		_w320_
	);
	LUT4 #(
		.INIT('h00e0)
	) name184 (
		\j2_pad ,
		\k2_pad ,
		\r3_pad ,
		\x1_pad ,
		_w321_
	);
	LUT3 #(
		.INIT('h02)
	) name185 (
		_w190_,
		_w321_,
		_w320_,
		_w322_
	);
	LUT4 #(
		.INIT('h0004)
	) name186 (
		\a3_pad ,
		c_pad,
		d_pad,
		e_pad,
		_w323_
	);
	LUT3 #(
		.INIT('h02)
	) name187 (
		d_pad,
		e_pad,
		\z0_pad ,
		_w324_
	);
	LUT3 #(
		.INIT('h0d)
	) name188 (
		e_pad,
		\p1_pad ,
		\y1_pad ,
		_w325_
	);
	LUT3 #(
		.INIT('h10)
	) name189 (
		_w324_,
		_w323_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w322_,
		_w326_,
		_w327_
	);
	LUT3 #(
		.INIT('h02)
	) name191 (
		i_pad,
		j_pad,
		r_pad,
		_w328_
	);
	LUT4 #(
		.INIT('h00ce)
	) name192 (
		i_pad,
		\r0_pad ,
		r_pad,
		\y1_pad ,
		_w329_
	);
	LUT2 #(
		.INIT('h4)
	) name193 (
		_w328_,
		_w329_,
		_w330_
	);
	LUT3 #(
		.INIT('h08)
	) name194 (
		\b0_pad ,
		s_pad,
		v_pad,
		_w331_
	);
	LUT4 #(
		.INIT('h00ec)
	) name195 (
		\b0_pad ,
		\r1_pad ,
		s_pad,
		\y1_pad ,
		_w332_
	);
	LUT2 #(
		.INIT('h4)
	) name196 (
		_w331_,
		_w332_,
		_w333_
	);
	LUT3 #(
		.INIT('h12)
	) name197 (
		\r2_pad ,
		\y1_pad ,
		_w318_,
		_w334_
	);
	LUT4 #(
		.INIT('hf010)
	) name198 (
		\j2_pad ,
		\k2_pad ,
		\r3_pad ,
		\x1_pad ,
		_w335_
	);
	LUT4 #(
		.INIT('h00e0)
	) name199 (
		\j2_pad ,
		\k2_pad ,
		\s3_pad ,
		\x1_pad ,
		_w336_
	);
	LUT3 #(
		.INIT('h02)
	) name200 (
		_w190_,
		_w336_,
		_w335_,
		_w337_
	);
	LUT4 #(
		.INIT('h0004)
	) name201 (
		\b3_pad ,
		c_pad,
		d_pad,
		e_pad,
		_w338_
	);
	LUT3 #(
		.INIT('h04)
	) name202 (
		\a1_pad ,
		d_pad,
		e_pad,
		_w339_
	);
	LUT3 #(
		.INIT('h0d)
	) name203 (
		e_pad,
		\q1_pad ,
		\y1_pad ,
		_w340_
	);
	LUT3 #(
		.INIT('h10)
	) name204 (
		_w339_,
		_w338_,
		_w340_,
		_w341_
	);
	LUT2 #(
		.INIT('h4)
	) name205 (
		_w337_,
		_w341_,
		_w342_
	);
	LUT3 #(
		.INIT('h02)
	) name206 (
		i_pad,
		k_pad,
		r_pad,
		_w343_
	);
	LUT4 #(
		.INIT('h00f2)
	) name207 (
		i_pad,
		r_pad,
		\s0_pad ,
		\y1_pad ,
		_w344_
	);
	LUT2 #(
		.INIT('h4)
	) name208 (
		_w343_,
		_w344_,
		_w345_
	);
	LUT3 #(
		.INIT('h08)
	) name209 (
		\b0_pad ,
		s_pad,
		w_pad,
		_w346_
	);
	LUT4 #(
		.INIT('h00ec)
	) name210 (
		\b0_pad ,
		\s1_pad ,
		s_pad,
		\y1_pad ,
		_w347_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT3 #(
		.INIT('h02)
	) name212 (
		f_pad,
		h_pad,
		\t2_pad ,
		_w349_
	);
	LUT4 #(
		.INIT('h00f2)
	) name213 (
		f_pad,
		h_pad,
		\s2_pad ,
		\y1_pad ,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w349_,
		_w350_,
		_w351_
	);
	LUT4 #(
		.INIT('hf010)
	) name215 (
		\j2_pad ,
		\k2_pad ,
		\s3_pad ,
		\x1_pad ,
		_w352_
	);
	LUT4 #(
		.INIT('h00e0)
	) name216 (
		\j2_pad ,
		\k2_pad ,
		\t3_pad ,
		\x1_pad ,
		_w353_
	);
	LUT3 #(
		.INIT('h02)
	) name217 (
		_w190_,
		_w353_,
		_w352_,
		_w354_
	);
	LUT4 #(
		.INIT('h0004)
	) name218 (
		\c3_pad ,
		c_pad,
		d_pad,
		e_pad,
		_w355_
	);
	LUT3 #(
		.INIT('h04)
	) name219 (
		\b1_pad ,
		d_pad,
		e_pad,
		_w356_
	);
	LUT3 #(
		.INIT('h0d)
	) name220 (
		e_pad,
		\r1_pad ,
		\y1_pad ,
		_w357_
	);
	LUT3 #(
		.INIT('h10)
	) name221 (
		_w356_,
		_w355_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w354_,
		_w358_,
		_w359_
	);
	LUT3 #(
		.INIT('h02)
	) name223 (
		i_pad,
		l_pad,
		r_pad,
		_w360_
	);
	LUT4 #(
		.INIT('h00f2)
	) name224 (
		i_pad,
		r_pad,
		\t0_pad ,
		\y1_pad ,
		_w361_
	);
	LUT2 #(
		.INIT('h4)
	) name225 (
		_w360_,
		_w361_,
		_w362_
	);
	LUT3 #(
		.INIT('h08)
	) name226 (
		\b0_pad ,
		s_pad,
		x_pad,
		_w363_
	);
	LUT4 #(
		.INIT('h00f8)
	) name227 (
		\b0_pad ,
		s_pad,
		\t1_pad ,
		\y1_pad ,
		_w364_
	);
	LUT2 #(
		.INIT('h4)
	) name228 (
		_w363_,
		_w364_,
		_w365_
	);
	LUT3 #(
		.INIT('h02)
	) name229 (
		f_pad,
		h_pad,
		\u2_pad ,
		_w366_
	);
	LUT4 #(
		.INIT('h00f2)
	) name230 (
		f_pad,
		h_pad,
		\t2_pad ,
		\y1_pad ,
		_w367_
	);
	LUT2 #(
		.INIT('h4)
	) name231 (
		_w366_,
		_w367_,
		_w368_
	);
	LUT4 #(
		.INIT('hf010)
	) name232 (
		\j2_pad ,
		\k2_pad ,
		\t3_pad ,
		\x1_pad ,
		_w369_
	);
	LUT4 #(
		.INIT('h00e0)
	) name233 (
		\j2_pad ,
		\k2_pad ,
		\u3_pad ,
		\x1_pad ,
		_w370_
	);
	LUT3 #(
		.INIT('h02)
	) name234 (
		_w190_,
		_w370_,
		_w369_,
		_w371_
	);
	LUT4 #(
		.INIT('h0002)
	) name235 (
		c_pad,
		\d3_pad ,
		d_pad,
		e_pad,
		_w372_
	);
	LUT3 #(
		.INIT('h04)
	) name236 (
		\c1_pad ,
		d_pad,
		e_pad,
		_w373_
	);
	LUT3 #(
		.INIT('h0d)
	) name237 (
		e_pad,
		\s1_pad ,
		\y1_pad ,
		_w374_
	);
	LUT3 #(
		.INIT('h10)
	) name238 (
		_w373_,
		_w372_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		_w371_,
		_w375_,
		_w376_
	);
	LUT3 #(
		.INIT('h02)
	) name240 (
		i_pad,
		m_pad,
		r_pad,
		_w377_
	);
	LUT4 #(
		.INIT('h00f2)
	) name241 (
		i_pad,
		r_pad,
		\u0_pad ,
		\y1_pad ,
		_w378_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		_w377_,
		_w378_,
		_w379_
	);
	LUT3 #(
		.INIT('h08)
	) name243 (
		\b0_pad ,
		s_pad,
		y_pad,
		_w380_
	);
	LUT4 #(
		.INIT('h00f8)
	) name244 (
		\b0_pad ,
		s_pad,
		\u1_pad ,
		\y1_pad ,
		_w381_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		_w380_,
		_w381_,
		_w382_
	);
	LUT3 #(
		.INIT('h02)
	) name246 (
		f_pad,
		h_pad,
		\v2_pad ,
		_w383_
	);
	LUT4 #(
		.INIT('h00f2)
	) name247 (
		f_pad,
		h_pad,
		\u2_pad ,
		\y1_pad ,
		_w384_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT4 #(
		.INIT('hf010)
	) name249 (
		\j2_pad ,
		\k2_pad ,
		\u3_pad ,
		\x1_pad ,
		_w386_
	);
	LUT4 #(
		.INIT('h00e0)
	) name250 (
		\j2_pad ,
		\k2_pad ,
		\v3_pad ,
		\x1_pad ,
		_w387_
	);
	LUT3 #(
		.INIT('h02)
	) name251 (
		_w190_,
		_w387_,
		_w386_,
		_w388_
	);
	LUT4 #(
		.INIT('h0002)
	) name252 (
		c_pad,
		d_pad,
		\e3_pad ,
		e_pad,
		_w389_
	);
	LUT3 #(
		.INIT('h04)
	) name253 (
		\d1_pad ,
		d_pad,
		e_pad,
		_w390_
	);
	LUT3 #(
		.INIT('h0d)
	) name254 (
		e_pad,
		\t1_pad ,
		\y1_pad ,
		_w391_
	);
	LUT3 #(
		.INIT('h10)
	) name255 (
		_w390_,
		_w389_,
		_w391_,
		_w392_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		_w388_,
		_w392_,
		_w393_
	);
	LUT3 #(
		.INIT('h02)
	) name257 (
		i_pad,
		n_pad,
		r_pad,
		_w394_
	);
	LUT4 #(
		.INIT('h00f2)
	) name258 (
		i_pad,
		r_pad,
		\v0_pad ,
		\y1_pad ,
		_w395_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w394_,
		_w395_,
		_w396_
	);
	LUT3 #(
		.INIT('h08)
	) name260 (
		\b0_pad ,
		s_pad,
		z_pad,
		_w397_
	);
	LUT4 #(
		.INIT('h00f8)
	) name261 (
		\b0_pad ,
		s_pad,
		\v1_pad ,
		\y1_pad ,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		_w397_,
		_w398_,
		_w399_
	);
	LUT3 #(
		.INIT('h02)
	) name263 (
		f_pad,
		h_pad,
		\w2_pad ,
		_w400_
	);
	LUT4 #(
		.INIT('h00f2)
	) name264 (
		f_pad,
		h_pad,
		\v2_pad ,
		\y1_pad ,
		_w401_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		_w400_,
		_w401_,
		_w402_
	);
	LUT4 #(
		.INIT('hf010)
	) name266 (
		\j2_pad ,
		\k2_pad ,
		\v3_pad ,
		\x1_pad ,
		_w403_
	);
	LUT4 #(
		.INIT('h00e0)
	) name267 (
		\j2_pad ,
		\k2_pad ,
		\w3_pad ,
		\x1_pad ,
		_w404_
	);
	LUT3 #(
		.INIT('h02)
	) name268 (
		_w190_,
		_w404_,
		_w403_,
		_w405_
	);
	LUT4 #(
		.INIT('h0002)
	) name269 (
		c_pad,
		d_pad,
		e_pad,
		\f3_pad ,
		_w406_
	);
	LUT3 #(
		.INIT('h02)
	) name270 (
		d_pad,
		\e1_pad ,
		e_pad,
		_w407_
	);
	LUT3 #(
		.INIT('h0d)
	) name271 (
		e_pad,
		\u1_pad ,
		\y1_pad ,
		_w408_
	);
	LUT3 #(
		.INIT('h10)
	) name272 (
		_w407_,
		_w406_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h4)
	) name273 (
		_w405_,
		_w409_,
		_w410_
	);
	LUT3 #(
		.INIT('h02)
	) name274 (
		i_pad,
		o_pad,
		r_pad,
		_w411_
	);
	LUT4 #(
		.INIT('h00f2)
	) name275 (
		i_pad,
		r_pad,
		\w0_pad ,
		\y1_pad ,
		_w412_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		_w411_,
		_w412_,
		_w413_
	);
	LUT3 #(
		.INIT('h40)
	) name277 (
		\a0_pad ,
		\b0_pad ,
		s_pad,
		_w414_
	);
	LUT4 #(
		.INIT('h00f8)
	) name278 (
		\b0_pad ,
		s_pad,
		\w1_pad ,
		\y1_pad ,
		_w415_
	);
	LUT2 #(
		.INIT('h4)
	) name279 (
		_w414_,
		_w415_,
		_w416_
	);
	LUT3 #(
		.INIT('h02)
	) name280 (
		f_pad,
		h_pad,
		\x2_pad ,
		_w417_
	);
	LUT4 #(
		.INIT('h00f2)
	) name281 (
		f_pad,
		h_pad,
		\w2_pad ,
		\y1_pad ,
		_w418_
	);
	LUT2 #(
		.INIT('h4)
	) name282 (
		_w417_,
		_w418_,
		_w419_
	);
	LUT4 #(
		.INIT('hf010)
	) name283 (
		\j2_pad ,
		\k2_pad ,
		\w3_pad ,
		\x1_pad ,
		_w420_
	);
	LUT4 #(
		.INIT('h0e00)
	) name284 (
		\j2_pad ,
		\k2_pad ,
		\x1_pad ,
		\x3_pad ,
		_w421_
	);
	LUT3 #(
		.INIT('h02)
	) name285 (
		_w190_,
		_w421_,
		_w420_,
		_w422_
	);
	LUT4 #(
		.INIT('h0002)
	) name286 (
		c_pad,
		d_pad,
		e_pad,
		\g3_pad ,
		_w423_
	);
	LUT3 #(
		.INIT('h02)
	) name287 (
		d_pad,
		e_pad,
		\f1_pad ,
		_w424_
	);
	LUT3 #(
		.INIT('h0d)
	) name288 (
		e_pad,
		\v1_pad ,
		\y1_pad ,
		_w425_
	);
	LUT3 #(
		.INIT('h10)
	) name289 (
		_w424_,
		_w423_,
		_w425_,
		_w426_
	);
	LUT2 #(
		.INIT('h4)
	) name290 (
		_w422_,
		_w426_,
		_w427_
	);
	LUT3 #(
		.INIT('h02)
	) name291 (
		i_pad,
		p_pad,
		r_pad,
		_w428_
	);
	LUT4 #(
		.INIT('h00f2)
	) name292 (
		i_pad,
		r_pad,
		\x0_pad ,
		\y1_pad ,
		_w429_
	);
	LUT2 #(
		.INIT('h4)
	) name293 (
		_w428_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('he)
	) name294 (
		\y1_pad ,
		_w232_,
		_w431_
	);
	LUT3 #(
		.INIT('h02)
	) name295 (
		f_pad,
		h_pad,
		\y2_pad ,
		_w432_
	);
	LUT4 #(
		.INIT('h00f2)
	) name296 (
		f_pad,
		h_pad,
		\x2_pad ,
		\y1_pad ,
		_w433_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		_w432_,
		_w433_,
		_w434_
	);
	LUT4 #(
		.INIT('hf100)
	) name298 (
		\j2_pad ,
		\k2_pad ,
		\x1_pad ,
		\x3_pad ,
		_w435_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		_w190_,
		_w435_,
		_w436_
	);
	LUT4 #(
		.INIT('h0002)
	) name300 (
		c_pad,
		d_pad,
		e_pad,
		\h3_pad ,
		_w437_
	);
	LUT3 #(
		.INIT('h02)
	) name301 (
		d_pad,
		e_pad,
		\g1_pad ,
		_w438_
	);
	LUT3 #(
		.INIT('h0d)
	) name302 (
		e_pad,
		\w1_pad ,
		\y1_pad ,
		_w439_
	);
	LUT3 #(
		.INIT('h10)
	) name303 (
		_w437_,
		_w438_,
		_w439_,
		_w440_
	);
	LUT2 #(
		.INIT('h4)
	) name304 (
		_w436_,
		_w440_,
		_w441_
	);
	LUT3 #(
		.INIT('h02)
	) name305 (
		i_pad,
		q_pad,
		r_pad,
		_w442_
	);
	LUT4 #(
		.INIT('h00f2)
	) name306 (
		i_pad,
		r_pad,
		\y0_pad ,
		\y1_pad ,
		_w443_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w442_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('he)
	) name308 (
		\n0_pad ,
		_w269_,
		_w445_
	);
	LUT3 #(
		.INIT('h02)
	) name309 (
		f_pad,
		h_pad,
		\z2_pad ,
		_w446_
	);
	LUT4 #(
		.INIT('h0f02)
	) name310 (
		f_pad,
		h_pad,
		\y1_pad ,
		\y2_pad ,
		_w447_
	);
	LUT2 #(
		.INIT('h4)
	) name311 (
		_w446_,
		_w447_,
		_w448_
	);
	LUT3 #(
		.INIT('h01)
	) name312 (
		\l0_pad ,
		\n0_pad ,
		\y3_pad ,
		_w449_
	);
	LUT3 #(
		.INIT('h20)
	) name313 (
		i_pad,
		j_pad,
		r_pad,
		_w450_
	);
	LUT4 #(
		.INIT('h0f08)
	) name314 (
		i_pad,
		r_pad,
		\y1_pad ,
		\z0_pad ,
		_w451_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		_w450_,
		_w451_,
		_w452_
	);
	LUT3 #(
		.INIT('h01)
	) name316 (
		\i3_pad ,
		_w187_,
		_w283_,
		_w453_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name317 (
		\c0_pad ,
		\d0_pad ,
		\q2_pad ,
		\r2_pad ,
		_w454_
	);
	LUT3 #(
		.INIT('h31)
	) name318 (
		\i2_pad ,
		\x1_pad ,
		_w454_,
		_w455_
	);
	LUT4 #(
		.INIT('h0d00)
	) name319 (
		_w284_,
		_w288_,
		_w453_,
		_w455_,
		_w456_
	);
	LUT4 #(
		.INIT('h5054)
	) name320 (
		\y1_pad ,
		\z1_pad ,
		_w269_,
		_w456_,
		_w457_
	);
	LUT3 #(
		.INIT('h02)
	) name321 (
		\i3_pad ,
		_w187_,
		_w283_,
		_w458_
	);
	LUT3 #(
		.INIT('h2a)
	) name322 (
		\c0_pad ,
		\d0_pad ,
		\r2_pad ,
		_w459_
	);
	LUT2 #(
		.INIT('h2)
	) name323 (
		_w289_,
		_w459_,
		_w460_
	);
	LUT4 #(
		.INIT('h0007)
	) name324 (
		_w284_,
		_w288_,
		_w458_,
		_w460_,
		_w461_
	);
	LUT3 #(
		.INIT('h01)
	) name325 (
		\x1_pad ,
		\y1_pad ,
		\z1_pad ,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w461_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('he)
	) name327 (
		_w457_,
		_w463_,
		_w464_
	);
	LUT3 #(
		.INIT('h02)
	) name328 (
		f_pad,
		g_pad,
		h_pad,
		_w465_
	);
	LUT4 #(
		.INIT('h0f02)
	) name329 (
		f_pad,
		h_pad,
		\y1_pad ,
		\z2_pad ,
		_w466_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		_w465_,
		_w466_,
		_w467_
	);
	LUT4 #(
		.INIT('h0110)
	) name331 (
		\l0_pad ,
		\n0_pad ,
		\y3_pad ,
		\z3_pad ,
		_w468_
	);
	LUT3 #(
		.INIT('h20)
	) name332 (
		i_pad,
		k_pad,
		r_pad,
		_w469_
	);
	LUT4 #(
		.INIT('h00ea)
	) name333 (
		\a1_pad ,
		i_pad,
		r_pad,
		\y1_pad ,
		_w470_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w469_,
		_w470_,
		_w471_
	);
	LUT4 #(
		.INIT('h0007)
	) name335 (
		_w142_,
		_w147_,
		_w150_,
		_w296_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		\y1_pad ,
		_w472_,
		_w473_
	);
	LUT3 #(
		.INIT('h40)
	) name337 (
		\b3_pad ,
		f_pad,
		h_pad,
		_w474_
	);
	LUT4 #(
		.INIT('h00ea)
	) name338 (
		\a3_pad ,
		f_pad,
		h_pad,
		\y1_pad ,
		_w475_
	);
	LUT2 #(
		.INIT('h4)
	) name339 (
		_w474_,
		_w475_,
		_w476_
	);
	LUT3 #(
		.INIT('h15)
	) name340 (
		\a4_pad ,
		\y3_pad ,
		\z3_pad ,
		_w477_
	);
	LUT3 #(
		.INIT('h04)
	) name341 (
		_w140_,
		_w158_,
		_w477_,
		_w478_
	);
	LUT3 #(
		.INIT('h20)
	) name342 (
		i_pad,
		l_pad,
		r_pad,
		_w479_
	);
	LUT4 #(
		.INIT('h00ea)
	) name343 (
		\b1_pad ,
		i_pad,
		r_pad,
		\y1_pad ,
		_w480_
	);
	LUT2 #(
		.INIT('h4)
	) name344 (
		_w479_,
		_w480_,
		_w481_
	);
	LUT3 #(
		.INIT('h01)
	) name345 (
		\e4_pad ,
		\f4_pad ,
		\g4_pad ,
		_w482_
	);
	LUT4 #(
		.INIT('h8000)
	) name346 (
		\c4_pad ,
		\d4_pad ,
		_w141_,
		_w482_,
		_w483_
	);
	LUT3 #(
		.INIT('h48)
	) name347 (
		\b2_pad ,
		_w158_,
		_w483_,
		_w484_
	);
	LUT3 #(
		.INIT('h40)
	) name348 (
		\c3_pad ,
		f_pad,
		h_pad,
		_w485_
	);
	LUT4 #(
		.INIT('h00ea)
	) name349 (
		\b3_pad ,
		f_pad,
		h_pad,
		\y1_pad ,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w485_,
		_w486_,
		_w487_
	);
	LUT3 #(
		.INIT('h60)
	) name351 (
		\b4_pad ,
		_w140_,
		_w158_,
		_w488_
	);
	LUT3 #(
		.INIT('h20)
	) name352 (
		i_pad,
		m_pad,
		r_pad,
		_w489_
	);
	LUT4 #(
		.INIT('h00ea)
	) name353 (
		\c1_pad ,
		i_pad,
		r_pad,
		\y1_pad ,
		_w490_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		_w489_,
		_w490_,
		_w491_
	);
	LUT4 #(
		.INIT('h60c0)
	) name355 (
		\b2_pad ,
		\c2_pad ,
		_w158_,
		_w483_,
		_w492_
	);
	LUT3 #(
		.INIT('h40)
	) name356 (
		\d3_pad ,
		f_pad,
		h_pad,
		_w493_
	);
	LUT4 #(
		.INIT('h00ea)
	) name357 (
		\c3_pad ,
		f_pad,
		h_pad,
		\y1_pad ,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		_w493_,
		_w494_,
		_w495_
	);
	LUT3 #(
		.INIT('h60)
	) name359 (
		\c4_pad ,
		_w141_,
		_w158_,
		_w496_
	);
	LUT3 #(
		.INIT('h20)
	) name360 (
		i_pad,
		n_pad,
		r_pad,
		_w497_
	);
	LUT4 #(
		.INIT('h00ea)
	) name361 (
		\d1_pad ,
		i_pad,
		r_pad,
		\y1_pad ,
		_w498_
	);
	LUT2 #(
		.INIT('h4)
	) name362 (
		_w497_,
		_w498_,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		\d2_pad ,
		\l0_pad ,
		_w500_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		_w176_,
		_w500_,
		_w501_
	);
	LUT3 #(
		.INIT('h40)
	) name365 (
		\e3_pad ,
		f_pad,
		h_pad,
		_w502_
	);
	LUT4 #(
		.INIT('h00ea)
	) name366 (
		\d3_pad ,
		f_pad,
		h_pad,
		\y1_pad ,
		_w503_
	);
	LUT2 #(
		.INIT('h4)
	) name367 (
		_w502_,
		_w503_,
		_w504_
	);
	LUT4 #(
		.INIT('h6c00)
	) name368 (
		\c4_pad ,
		\d4_pad ,
		_w141_,
		_w158_,
		_w505_
	);
	LUT3 #(
		.INIT('h20)
	) name369 (
		i_pad,
		o_pad,
		r_pad,
		_w506_
	);
	LUT4 #(
		.INIT('h00ea)
	) name370 (
		\e1_pad ,
		i_pad,
		r_pad,
		\y1_pad ,
		_w507_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		_w506_,
		_w507_,
		_w508_
	);
	LUT3 #(
		.INIT('h21)
	) name372 (
		\e2_pad ,
		\n0_pad ,
		_w151_,
		_w509_
	);
	LUT3 #(
		.INIT('h40)
	) name373 (
		\f3_pad ,
		f_pad,
		h_pad,
		_w510_
	);
	LUT4 #(
		.INIT('h00ea)
	) name374 (
		\e3_pad ,
		f_pad,
		h_pad,
		\y1_pad ,
		_w511_
	);
	LUT2 #(
		.INIT('h4)
	) name375 (
		_w510_,
		_w511_,
		_w512_
	);
	LUT3 #(
		.INIT('h48)
	) name376 (
		\e4_pad ,
		_w158_,
		_w156_,
		_w513_
	);
	assign \a5_pad  = _w139_ ;
	assign \a6_pad  = _w152_ ;
	assign \a7_pad  = _w155_ ;
	assign \a8_pad  = _w159_ ;
	assign \b5_pad  = _w162_ ;
	assign \b6_pad  = _w163_ ;
	assign \b7_pad  = _w166_ ;
	assign \b8_pad  = _w167_ ;
	assign \c5_pad  = _w170_ ;
	assign \c6_pad  = _w171_ ;
	assign \c7_pad  = _w174_ ;
	assign \c8_pad  = _w177_ ;
	assign \d5_pad  = _w180_ ;
	assign \d6_pad  = _w186_ ;
	assign \d7_pad  = _w196_ ;
	assign \e5_pad  = _w199_ ;
	assign \e6_pad  = _w205_ ;
	assign \e7_pad  = _w213_ ;
	assign \f5_pad  = _w216_ ;
	assign \f6_pad  = _w220_ ;
	assign \f7_pad  = _w228_ ;
	assign \g5_pad  = _w231_ ;
	assign \g6_pad  = _w233_ ;
	assign \g7_pad  = _w241_ ;
	assign \h5_pad  = _w244_ ;
	assign \h6_pad  = _w246_ ;
	assign \h7_pad  = _w254_ ;
	assign \i4_pad  = _w255_ ;
	assign \i5_pad  = _w258_ ;
	assign \i6_pad  = _w260_ ;
	assign \i7_pad  = _w268_ ;
	assign \j4_pad  = _w270_ ;
	assign \j5_pad  = _w273_ ;
	assign \j6_pad  = _w274_ ;
	assign \j7_pad  = _w282_ ;
	assign \k4_pad  = _w300_ ;
	assign \k5_pad  = _w303_ ;
	assign \k6_pad  = _w304_ ;
	assign \k7_pad  = _w312_ ;
	assign \l4_pad  = _w313_ ;
	assign \l5_pad  = _w316_ ;
	assign \l6_pad  = _w319_ ;
	assign \l7_pad  = _w327_ ;
	assign \m4_pad  = _w330_ ;
	assign \m5_pad  = _w333_ ;
	assign \m6_pad  = _w334_ ;
	assign \m7_pad  = _w342_ ;
	assign \n4_pad  = _w345_ ;
	assign \n5_pad  = _w348_ ;
	assign \n6_pad  = _w351_ ;
	assign \n7_pad  = _w359_ ;
	assign \o4_pad  = _w362_ ;
	assign \o5_pad  = _w365_ ;
	assign \o6_pad  = _w368_ ;
	assign \o7_pad  = _w376_ ;
	assign \p4_pad  = _w379_ ;
	assign \p5_pad  = _w382_ ;
	assign \p6_pad  = _w385_ ;
	assign \p7_pad  = _w393_ ;
	assign \q4_pad  = _w396_ ;
	assign \q5_pad  = _w399_ ;
	assign \q6_pad  = _w402_ ;
	assign \q7_pad  = _w410_ ;
	assign \r4_pad  = _w413_ ;
	assign \r5_pad  = _w416_ ;
	assign \r6_pad  = _w419_ ;
	assign \r7_pad  = _w427_ ;
	assign \s4_pad  = _w430_ ;
	assign \s5_pad  = _w431_ ;
	assign \s6_pad  = _w434_ ;
	assign \s7_pad  = _w441_ ;
	assign \t4_pad  = _w444_ ;
	assign \t5_pad  = _w445_ ;
	assign \t6_pad  = _w448_ ;
	assign \t7_pad  = _w449_ ;
	assign \u4_pad  = _w452_ ;
	assign \u5_pad  = _w464_ ;
	assign \u6_pad  = _w467_ ;
	assign \u7_pad  = _w468_ ;
	assign \v4_pad  = _w471_ ;
	assign \v5_pad  = _w473_ ;
	assign \v6_pad  = _w476_ ;
	assign \v7_pad  = _w478_ ;
	assign \w4_pad  = _w481_ ;
	assign \w5_pad  = _w484_ ;
	assign \w6_pad  = _w487_ ;
	assign \w7_pad  = _w488_ ;
	assign \x4_pad  = _w491_ ;
	assign \x5_pad  = _w492_ ;
	assign \x6_pad  = _w495_ ;
	assign \x7_pad  = _w496_ ;
	assign \y4_pad  = _w499_ ;
	assign \y5_pad  = _w501_ ;
	assign \y6_pad  = _w504_ ;
	assign \y7_pad  = _w505_ ;
	assign \z4_pad  = _w508_ ;
	assign \z5_pad  = _w509_ ;
	assign \z6_pad  = _w512_ ;
	assign \z7_pad  = _w513_ ;
endmodule;