module top (\in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] , \result[0] , \result[1] , \result[2] , \result[3] , \result[4] , \result[5] , \result[6] , \result[7] , \result[8] , \result[9] , \result[10] , \result[11] , \result[12] , \result[13] , \result[14] , \result[15] , \result[16] , \result[17] , \result[18] , \result[19] , \result[20] , \result[21] , \result[22] , \result[23] , \result[24] , \result[25] , \result[26] , \result[27] , \result[28] , \result[29] , \result[30] , \result[31] , \result[32] , \result[33] , \result[34] , \result[35] , \result[36] , \result[37] , \result[38] , \result[39] , \result[40] , \result[41] , \result[42] , \result[43] , \result[44] , \result[45] , \result[46] , \result[47] , \result[48] , \result[49] , \result[50] , \result[51] , \result[52] , \result[53] , \result[54] , \result[55] , \result[56] , \result[57] , \result[58] , \result[59] , \result[60] , \result[61] , \result[62] , \result[63] , \result[64] , \result[65] , \result[66] , \result[67] , \result[68] , \result[69] , \result[70] , \result[71] , \result[72] , \result[73] , \result[74] , \result[75] , \result[76] , \result[77] , \result[78] , \result[79] , \result[80] , \result[81] , \result[82] , \result[83] , \result[84] , \result[85] , \result[86] , \result[87] , \result[88] , \result[89] , \result[90] , \result[91] , \result[92] , \result[93] , \result[94] , \result[95] , \result[96] , \result[97] , \result[98] , \result[99] , \result[100] , \result[101] , \result[102] , \result[103] , \result[104] , \result[105] , \result[106] , \result[107] , \result[108] , \result[109] , \result[110] , \result[111] , \result[112] , \result[113] , \result[114] , \result[115] , \result[116] , \result[117] , \result[118] , \result[119] , \result[120] , \result[121] , \result[122] , \result[123] , \result[124] , \result[125] , \result[126] , \result[127] , \address[0] , \address[1] );
	input \in0[0]  ;
	input \in0[1]  ;
	input \in0[2]  ;
	input \in0[3]  ;
	input \in0[4]  ;
	input \in0[5]  ;
	input \in0[6]  ;
	input \in0[7]  ;
	input \in0[8]  ;
	input \in0[9]  ;
	input \in0[10]  ;
	input \in0[11]  ;
	input \in0[12]  ;
	input \in0[13]  ;
	input \in0[14]  ;
	input \in0[15]  ;
	input \in0[16]  ;
	input \in0[17]  ;
	input \in0[18]  ;
	input \in0[19]  ;
	input \in0[20]  ;
	input \in0[21]  ;
	input \in0[22]  ;
	input \in0[23]  ;
	input \in0[24]  ;
	input \in0[25]  ;
	input \in0[26]  ;
	input \in0[27]  ;
	input \in0[28]  ;
	input \in0[29]  ;
	input \in0[30]  ;
	input \in0[31]  ;
	input \in0[32]  ;
	input \in0[33]  ;
	input \in0[34]  ;
	input \in0[35]  ;
	input \in0[36]  ;
	input \in0[37]  ;
	input \in0[38]  ;
	input \in0[39]  ;
	input \in0[40]  ;
	input \in0[41]  ;
	input \in0[42]  ;
	input \in0[43]  ;
	input \in0[44]  ;
	input \in0[45]  ;
	input \in0[46]  ;
	input \in0[47]  ;
	input \in0[48]  ;
	input \in0[49]  ;
	input \in0[50]  ;
	input \in0[51]  ;
	input \in0[52]  ;
	input \in0[53]  ;
	input \in0[54]  ;
	input \in0[55]  ;
	input \in0[56]  ;
	input \in0[57]  ;
	input \in0[58]  ;
	input \in0[59]  ;
	input \in0[60]  ;
	input \in0[61]  ;
	input \in0[62]  ;
	input \in0[63]  ;
	input \in0[64]  ;
	input \in0[65]  ;
	input \in0[66]  ;
	input \in0[67]  ;
	input \in0[68]  ;
	input \in0[69]  ;
	input \in0[70]  ;
	input \in0[71]  ;
	input \in0[72]  ;
	input \in0[73]  ;
	input \in0[74]  ;
	input \in0[75]  ;
	input \in0[76]  ;
	input \in0[77]  ;
	input \in0[78]  ;
	input \in0[79]  ;
	input \in0[80]  ;
	input \in0[81]  ;
	input \in0[82]  ;
	input \in0[83]  ;
	input \in0[84]  ;
	input \in0[85]  ;
	input \in0[86]  ;
	input \in0[87]  ;
	input \in0[88]  ;
	input \in0[89]  ;
	input \in0[90]  ;
	input \in0[91]  ;
	input \in0[92]  ;
	input \in0[93]  ;
	input \in0[94]  ;
	input \in0[95]  ;
	input \in0[96]  ;
	input \in0[97]  ;
	input \in0[98]  ;
	input \in0[99]  ;
	input \in0[100]  ;
	input \in0[101]  ;
	input \in0[102]  ;
	input \in0[103]  ;
	input \in0[104]  ;
	input \in0[105]  ;
	input \in0[106]  ;
	input \in0[107]  ;
	input \in0[108]  ;
	input \in0[109]  ;
	input \in0[110]  ;
	input \in0[111]  ;
	input \in0[112]  ;
	input \in0[113]  ;
	input \in0[114]  ;
	input \in0[115]  ;
	input \in0[116]  ;
	input \in0[117]  ;
	input \in0[118]  ;
	input \in0[119]  ;
	input \in0[120]  ;
	input \in0[121]  ;
	input \in0[122]  ;
	input \in0[123]  ;
	input \in0[124]  ;
	input \in0[125]  ;
	input \in0[126]  ;
	input \in0[127]  ;
	input \in1[0]  ;
	input \in1[1]  ;
	input \in1[2]  ;
	input \in1[3]  ;
	input \in1[4]  ;
	input \in1[5]  ;
	input \in1[6]  ;
	input \in1[7]  ;
	input \in1[8]  ;
	input \in1[9]  ;
	input \in1[10]  ;
	input \in1[11]  ;
	input \in1[12]  ;
	input \in1[13]  ;
	input \in1[14]  ;
	input \in1[15]  ;
	input \in1[16]  ;
	input \in1[17]  ;
	input \in1[18]  ;
	input \in1[19]  ;
	input \in1[20]  ;
	input \in1[21]  ;
	input \in1[22]  ;
	input \in1[23]  ;
	input \in1[24]  ;
	input \in1[25]  ;
	input \in1[26]  ;
	input \in1[27]  ;
	input \in1[28]  ;
	input \in1[29]  ;
	input \in1[30]  ;
	input \in1[31]  ;
	input \in1[32]  ;
	input \in1[33]  ;
	input \in1[34]  ;
	input \in1[35]  ;
	input \in1[36]  ;
	input \in1[37]  ;
	input \in1[38]  ;
	input \in1[39]  ;
	input \in1[40]  ;
	input \in1[41]  ;
	input \in1[42]  ;
	input \in1[43]  ;
	input \in1[44]  ;
	input \in1[45]  ;
	input \in1[46]  ;
	input \in1[47]  ;
	input \in1[48]  ;
	input \in1[49]  ;
	input \in1[50]  ;
	input \in1[51]  ;
	input \in1[52]  ;
	input \in1[53]  ;
	input \in1[54]  ;
	input \in1[55]  ;
	input \in1[56]  ;
	input \in1[57]  ;
	input \in1[58]  ;
	input \in1[59]  ;
	input \in1[60]  ;
	input \in1[61]  ;
	input \in1[62]  ;
	input \in1[63]  ;
	input \in1[64]  ;
	input \in1[65]  ;
	input \in1[66]  ;
	input \in1[67]  ;
	input \in1[68]  ;
	input \in1[69]  ;
	input \in1[70]  ;
	input \in1[71]  ;
	input \in1[72]  ;
	input \in1[73]  ;
	input \in1[74]  ;
	input \in1[75]  ;
	input \in1[76]  ;
	input \in1[77]  ;
	input \in1[78]  ;
	input \in1[79]  ;
	input \in1[80]  ;
	input \in1[81]  ;
	input \in1[82]  ;
	input \in1[83]  ;
	input \in1[84]  ;
	input \in1[85]  ;
	input \in1[86]  ;
	input \in1[87]  ;
	input \in1[88]  ;
	input \in1[89]  ;
	input \in1[90]  ;
	input \in1[91]  ;
	input \in1[92]  ;
	input \in1[93]  ;
	input \in1[94]  ;
	input \in1[95]  ;
	input \in1[96]  ;
	input \in1[97]  ;
	input \in1[98]  ;
	input \in1[99]  ;
	input \in1[100]  ;
	input \in1[101]  ;
	input \in1[102]  ;
	input \in1[103]  ;
	input \in1[104]  ;
	input \in1[105]  ;
	input \in1[106]  ;
	input \in1[107]  ;
	input \in1[108]  ;
	input \in1[109]  ;
	input \in1[110]  ;
	input \in1[111]  ;
	input \in1[112]  ;
	input \in1[113]  ;
	input \in1[114]  ;
	input \in1[115]  ;
	input \in1[116]  ;
	input \in1[117]  ;
	input \in1[118]  ;
	input \in1[119]  ;
	input \in1[120]  ;
	input \in1[121]  ;
	input \in1[122]  ;
	input \in1[123]  ;
	input \in1[124]  ;
	input \in1[125]  ;
	input \in1[126]  ;
	input \in1[127]  ;
	input \in2[0]  ;
	input \in2[1]  ;
	input \in2[2]  ;
	input \in2[3]  ;
	input \in2[4]  ;
	input \in2[5]  ;
	input \in2[6]  ;
	input \in2[7]  ;
	input \in2[8]  ;
	input \in2[9]  ;
	input \in2[10]  ;
	input \in2[11]  ;
	input \in2[12]  ;
	input \in2[13]  ;
	input \in2[14]  ;
	input \in2[15]  ;
	input \in2[16]  ;
	input \in2[17]  ;
	input \in2[18]  ;
	input \in2[19]  ;
	input \in2[20]  ;
	input \in2[21]  ;
	input \in2[22]  ;
	input \in2[23]  ;
	input \in2[24]  ;
	input \in2[25]  ;
	input \in2[26]  ;
	input \in2[27]  ;
	input \in2[28]  ;
	input \in2[29]  ;
	input \in2[30]  ;
	input \in2[31]  ;
	input \in2[32]  ;
	input \in2[33]  ;
	input \in2[34]  ;
	input \in2[35]  ;
	input \in2[36]  ;
	input \in2[37]  ;
	input \in2[38]  ;
	input \in2[39]  ;
	input \in2[40]  ;
	input \in2[41]  ;
	input \in2[42]  ;
	input \in2[43]  ;
	input \in2[44]  ;
	input \in2[45]  ;
	input \in2[46]  ;
	input \in2[47]  ;
	input \in2[48]  ;
	input \in2[49]  ;
	input \in2[50]  ;
	input \in2[51]  ;
	input \in2[52]  ;
	input \in2[53]  ;
	input \in2[54]  ;
	input \in2[55]  ;
	input \in2[56]  ;
	input \in2[57]  ;
	input \in2[58]  ;
	input \in2[59]  ;
	input \in2[60]  ;
	input \in2[61]  ;
	input \in2[62]  ;
	input \in2[63]  ;
	input \in2[64]  ;
	input \in2[65]  ;
	input \in2[66]  ;
	input \in2[67]  ;
	input \in2[68]  ;
	input \in2[69]  ;
	input \in2[70]  ;
	input \in2[71]  ;
	input \in2[72]  ;
	input \in2[73]  ;
	input \in2[74]  ;
	input \in2[75]  ;
	input \in2[76]  ;
	input \in2[77]  ;
	input \in2[78]  ;
	input \in2[79]  ;
	input \in2[80]  ;
	input \in2[81]  ;
	input \in2[82]  ;
	input \in2[83]  ;
	input \in2[84]  ;
	input \in2[85]  ;
	input \in2[86]  ;
	input \in2[87]  ;
	input \in2[88]  ;
	input \in2[89]  ;
	input \in2[90]  ;
	input \in2[91]  ;
	input \in2[92]  ;
	input \in2[93]  ;
	input \in2[94]  ;
	input \in2[95]  ;
	input \in2[96]  ;
	input \in2[97]  ;
	input \in2[98]  ;
	input \in2[99]  ;
	input \in2[100]  ;
	input \in2[101]  ;
	input \in2[102]  ;
	input \in2[103]  ;
	input \in2[104]  ;
	input \in2[105]  ;
	input \in2[106]  ;
	input \in2[107]  ;
	input \in2[108]  ;
	input \in2[109]  ;
	input \in2[110]  ;
	input \in2[111]  ;
	input \in2[112]  ;
	input \in2[113]  ;
	input \in2[114]  ;
	input \in2[115]  ;
	input \in2[116]  ;
	input \in2[117]  ;
	input \in2[118]  ;
	input \in2[119]  ;
	input \in2[120]  ;
	input \in2[121]  ;
	input \in2[122]  ;
	input \in2[123]  ;
	input \in2[124]  ;
	input \in2[125]  ;
	input \in2[126]  ;
	input \in2[127]  ;
	input \in3[0]  ;
	input \in3[1]  ;
	input \in3[2]  ;
	input \in3[3]  ;
	input \in3[4]  ;
	input \in3[5]  ;
	input \in3[6]  ;
	input \in3[7]  ;
	input \in3[8]  ;
	input \in3[9]  ;
	input \in3[10]  ;
	input \in3[11]  ;
	input \in3[12]  ;
	input \in3[13]  ;
	input \in3[14]  ;
	input \in3[15]  ;
	input \in3[16]  ;
	input \in3[17]  ;
	input \in3[18]  ;
	input \in3[19]  ;
	input \in3[20]  ;
	input \in3[21]  ;
	input \in3[22]  ;
	input \in3[23]  ;
	input \in3[24]  ;
	input \in3[25]  ;
	input \in3[26]  ;
	input \in3[27]  ;
	input \in3[28]  ;
	input \in3[29]  ;
	input \in3[30]  ;
	input \in3[31]  ;
	input \in3[32]  ;
	input \in3[33]  ;
	input \in3[34]  ;
	input \in3[35]  ;
	input \in3[36]  ;
	input \in3[37]  ;
	input \in3[38]  ;
	input \in3[39]  ;
	input \in3[40]  ;
	input \in3[41]  ;
	input \in3[42]  ;
	input \in3[43]  ;
	input \in3[44]  ;
	input \in3[45]  ;
	input \in3[46]  ;
	input \in3[47]  ;
	input \in3[48]  ;
	input \in3[49]  ;
	input \in3[50]  ;
	input \in3[51]  ;
	input \in3[52]  ;
	input \in3[53]  ;
	input \in3[54]  ;
	input \in3[55]  ;
	input \in3[56]  ;
	input \in3[57]  ;
	input \in3[58]  ;
	input \in3[59]  ;
	input \in3[60]  ;
	input \in3[61]  ;
	input \in3[62]  ;
	input \in3[63]  ;
	input \in3[64]  ;
	input \in3[65]  ;
	input \in3[66]  ;
	input \in3[67]  ;
	input \in3[68]  ;
	input \in3[69]  ;
	input \in3[70]  ;
	input \in3[71]  ;
	input \in3[72]  ;
	input \in3[73]  ;
	input \in3[74]  ;
	input \in3[75]  ;
	input \in3[76]  ;
	input \in3[77]  ;
	input \in3[78]  ;
	input \in3[79]  ;
	input \in3[80]  ;
	input \in3[81]  ;
	input \in3[82]  ;
	input \in3[83]  ;
	input \in3[84]  ;
	input \in3[85]  ;
	input \in3[86]  ;
	input \in3[87]  ;
	input \in3[88]  ;
	input \in3[89]  ;
	input \in3[90]  ;
	input \in3[91]  ;
	input \in3[92]  ;
	input \in3[93]  ;
	input \in3[94]  ;
	input \in3[95]  ;
	input \in3[96]  ;
	input \in3[97]  ;
	input \in3[98]  ;
	input \in3[99]  ;
	input \in3[100]  ;
	input \in3[101]  ;
	input \in3[102]  ;
	input \in3[103]  ;
	input \in3[104]  ;
	input \in3[105]  ;
	input \in3[106]  ;
	input \in3[107]  ;
	input \in3[108]  ;
	input \in3[109]  ;
	input \in3[110]  ;
	input \in3[111]  ;
	input \in3[112]  ;
	input \in3[113]  ;
	input \in3[114]  ;
	input \in3[115]  ;
	input \in3[116]  ;
	input \in3[117]  ;
	input \in3[118]  ;
	input \in3[119]  ;
	input \in3[120]  ;
	input \in3[121]  ;
	input \in3[122]  ;
	input \in3[123]  ;
	input \in3[124]  ;
	input \in3[125]  ;
	input \in3[126]  ;
	input \in3[127]  ;
	output \result[0]  ;
	output \result[1]  ;
	output \result[2]  ;
	output \result[3]  ;
	output \result[4]  ;
	output \result[5]  ;
	output \result[6]  ;
	output \result[7]  ;
	output \result[8]  ;
	output \result[9]  ;
	output \result[10]  ;
	output \result[11]  ;
	output \result[12]  ;
	output \result[13]  ;
	output \result[14]  ;
	output \result[15]  ;
	output \result[16]  ;
	output \result[17]  ;
	output \result[18]  ;
	output \result[19]  ;
	output \result[20]  ;
	output \result[21]  ;
	output \result[22]  ;
	output \result[23]  ;
	output \result[24]  ;
	output \result[25]  ;
	output \result[26]  ;
	output \result[27]  ;
	output \result[28]  ;
	output \result[29]  ;
	output \result[30]  ;
	output \result[31]  ;
	output \result[32]  ;
	output \result[33]  ;
	output \result[34]  ;
	output \result[35]  ;
	output \result[36]  ;
	output \result[37]  ;
	output \result[38]  ;
	output \result[39]  ;
	output \result[40]  ;
	output \result[41]  ;
	output \result[42]  ;
	output \result[43]  ;
	output \result[44]  ;
	output \result[45]  ;
	output \result[46]  ;
	output \result[47]  ;
	output \result[48]  ;
	output \result[49]  ;
	output \result[50]  ;
	output \result[51]  ;
	output \result[52]  ;
	output \result[53]  ;
	output \result[54]  ;
	output \result[55]  ;
	output \result[56]  ;
	output \result[57]  ;
	output \result[58]  ;
	output \result[59]  ;
	output \result[60]  ;
	output \result[61]  ;
	output \result[62]  ;
	output \result[63]  ;
	output \result[64]  ;
	output \result[65]  ;
	output \result[66]  ;
	output \result[67]  ;
	output \result[68]  ;
	output \result[69]  ;
	output \result[70]  ;
	output \result[71]  ;
	output \result[72]  ;
	output \result[73]  ;
	output \result[74]  ;
	output \result[75]  ;
	output \result[76]  ;
	output \result[77]  ;
	output \result[78]  ;
	output \result[79]  ;
	output \result[80]  ;
	output \result[81]  ;
	output \result[82]  ;
	output \result[83]  ;
	output \result[84]  ;
	output \result[85]  ;
	output \result[86]  ;
	output \result[87]  ;
	output \result[88]  ;
	output \result[89]  ;
	output \result[90]  ;
	output \result[91]  ;
	output \result[92]  ;
	output \result[93]  ;
	output \result[94]  ;
	output \result[95]  ;
	output \result[96]  ;
	output \result[97]  ;
	output \result[98]  ;
	output \result[99]  ;
	output \result[100]  ;
	output \result[101]  ;
	output \result[102]  ;
	output \result[103]  ;
	output \result[104]  ;
	output \result[105]  ;
	output \result[106]  ;
	output \result[107]  ;
	output \result[108]  ;
	output \result[109]  ;
	output \result[110]  ;
	output \result[111]  ;
	output \result[112]  ;
	output \result[113]  ;
	output \result[114]  ;
	output \result[115]  ;
	output \result[116]  ;
	output \result[117]  ;
	output \result[118]  ;
	output \result[119]  ;
	output \result[120]  ;
	output \result[121]  ;
	output \result[122]  ;
	output \result[123]  ;
	output \result[124]  ;
	output \result[125]  ;
	output \result[126]  ;
	output \result[127]  ;
	output \address[0]  ;
	output \address[1]  ;
	wire _w2574_ ;
	wire _w2573_ ;
	wire _w2572_ ;
	wire _w2571_ ;
	wire _w2570_ ;
	wire _w2569_ ;
	wire _w2568_ ;
	wire _w2567_ ;
	wire _w2566_ ;
	wire _w2565_ ;
	wire _w2564_ ;
	wire _w2563_ ;
	wire _w2562_ ;
	wire _w2561_ ;
	wire _w2560_ ;
	wire _w2559_ ;
	wire _w2558_ ;
	wire _w2557_ ;
	wire _w2556_ ;
	wire _w2555_ ;
	wire _w2554_ ;
	wire _w2553_ ;
	wire _w2552_ ;
	wire _w2551_ ;
	wire _w2550_ ;
	wire _w2549_ ;
	wire _w2548_ ;
	wire _w2547_ ;
	wire _w2546_ ;
	wire _w2545_ ;
	wire _w2544_ ;
	wire _w2543_ ;
	wire _w2542_ ;
	wire _w2541_ ;
	wire _w2540_ ;
	wire _w2539_ ;
	wire _w2538_ ;
	wire _w2537_ ;
	wire _w2536_ ;
	wire _w2535_ ;
	wire _w2534_ ;
	wire _w2533_ ;
	wire _w2532_ ;
	wire _w2531_ ;
	wire _w2530_ ;
	wire _w2529_ ;
	wire _w2528_ ;
	wire _w2527_ ;
	wire _w2526_ ;
	wire _w2525_ ;
	wire _w2524_ ;
	wire _w2523_ ;
	wire _w2522_ ;
	wire _w2521_ ;
	wire _w2520_ ;
	wire _w2519_ ;
	wire _w2518_ ;
	wire _w2517_ ;
	wire _w2516_ ;
	wire _w2515_ ;
	wire _w2514_ ;
	wire _w2513_ ;
	wire _w2512_ ;
	wire _w2511_ ;
	wire _w2510_ ;
	wire _w2509_ ;
	wire _w2508_ ;
	wire _w2507_ ;
	wire _w2506_ ;
	wire _w2505_ ;
	wire _w2504_ ;
	wire _w2503_ ;
	wire _w2502_ ;
	wire _w2501_ ;
	wire _w2500_ ;
	wire _w2499_ ;
	wire _w2498_ ;
	wire _w2497_ ;
	wire _w2496_ ;
	wire _w2495_ ;
	wire _w2494_ ;
	wire _w2493_ ;
	wire _w2492_ ;
	wire _w2491_ ;
	wire _w2490_ ;
	wire _w2489_ ;
	wire _w2488_ ;
	wire _w2487_ ;
	wire _w2486_ ;
	wire _w2485_ ;
	wire _w2484_ ;
	wire _w2483_ ;
	wire _w2482_ ;
	wire _w2481_ ;
	wire _w2480_ ;
	wire _w2479_ ;
	wire _w2478_ ;
	wire _w2477_ ;
	wire _w2476_ ;
	wire _w2475_ ;
	wire _w2474_ ;
	wire _w2473_ ;
	wire _w2472_ ;
	wire _w2471_ ;
	wire _w2470_ ;
	wire _w2469_ ;
	wire _w2468_ ;
	wire _w2467_ ;
	wire _w2466_ ;
	wire _w2465_ ;
	wire _w2464_ ;
	wire _w2463_ ;
	wire _w2462_ ;
	wire _w2461_ ;
	wire _w2460_ ;
	wire _w2459_ ;
	wire _w2458_ ;
	wire _w2457_ ;
	wire _w2456_ ;
	wire _w2455_ ;
	wire _w2454_ ;
	wire _w2453_ ;
	wire _w2452_ ;
	wire _w2451_ ;
	wire _w2450_ ;
	wire _w2449_ ;
	wire _w2448_ ;
	wire _w2447_ ;
	wire _w2446_ ;
	wire _w2445_ ;
	wire _w2444_ ;
	wire _w2443_ ;
	wire _w2442_ ;
	wire _w2441_ ;
	wire _w2440_ ;
	wire _w2439_ ;
	wire _w2438_ ;
	wire _w2437_ ;
	wire _w2436_ ;
	wire _w2435_ ;
	wire _w2434_ ;
	wire _w2433_ ;
	wire _w2432_ ;
	wire _w2431_ ;
	wire _w2430_ ;
	wire _w2429_ ;
	wire _w2428_ ;
	wire _w2427_ ;
	wire _w2426_ ;
	wire _w2425_ ;
	wire _w2424_ ;
	wire _w2423_ ;
	wire _w2422_ ;
	wire _w2421_ ;
	wire _w2420_ ;
	wire _w2419_ ;
	wire _w2418_ ;
	wire _w2417_ ;
	wire _w2416_ ;
	wire _w2415_ ;
	wire _w2414_ ;
	wire _w2413_ ;
	wire _w2412_ ;
	wire _w2411_ ;
	wire _w2410_ ;
	wire _w2409_ ;
	wire _w2408_ ;
	wire _w2407_ ;
	wire _w2406_ ;
	wire _w2405_ ;
	wire _w2404_ ;
	wire _w2403_ ;
	wire _w2402_ ;
	wire _w2401_ ;
	wire _w2400_ ;
	wire _w2399_ ;
	wire _w2398_ ;
	wire _w2397_ ;
	wire _w2396_ ;
	wire _w2395_ ;
	wire _w2394_ ;
	wire _w2393_ ;
	wire _w2392_ ;
	wire _w2391_ ;
	wire _w2390_ ;
	wire _w2389_ ;
	wire _w2388_ ;
	wire _w2387_ ;
	wire _w2386_ ;
	wire _w2385_ ;
	wire _w2384_ ;
	wire _w2383_ ;
	wire _w2382_ ;
	wire _w2381_ ;
	wire _w2380_ ;
	wire _w2379_ ;
	wire _w2378_ ;
	wire _w2377_ ;
	wire _w2376_ ;
	wire _w2375_ ;
	wire _w2374_ ;
	wire _w2373_ ;
	wire _w2372_ ;
	wire _w2371_ ;
	wire _w2370_ ;
	wire _w2369_ ;
	wire _w2368_ ;
	wire _w2367_ ;
	wire _w2366_ ;
	wire _w2365_ ;
	wire _w2364_ ;
	wire _w2363_ ;
	wire _w2362_ ;
	wire _w2361_ ;
	wire _w2360_ ;
	wire _w2359_ ;
	wire _w2358_ ;
	wire _w2357_ ;
	wire _w2356_ ;
	wire _w2355_ ;
	wire _w2354_ ;
	wire _w2353_ ;
	wire _w2352_ ;
	wire _w2351_ ;
	wire _w2350_ ;
	wire _w2349_ ;
	wire _w2348_ ;
	wire _w2347_ ;
	wire _w2346_ ;
	wire _w2345_ ;
	wire _w2344_ ;
	wire _w2343_ ;
	wire _w2342_ ;
	wire _w2341_ ;
	wire _w2340_ ;
	wire _w2339_ ;
	wire _w2338_ ;
	wire _w2337_ ;
	wire _w2336_ ;
	wire _w2335_ ;
	wire _w2334_ ;
	wire _w2333_ ;
	wire _w2332_ ;
	wire _w2331_ ;
	wire _w2330_ ;
	wire _w2329_ ;
	wire _w2328_ ;
	wire _w2327_ ;
	wire _w2326_ ;
	wire _w2325_ ;
	wire _w2324_ ;
	wire _w2323_ ;
	wire _w2322_ ;
	wire _w2321_ ;
	wire _w2320_ ;
	wire _w2319_ ;
	wire _w2318_ ;
	wire _w2317_ ;
	wire _w2316_ ;
	wire _w2315_ ;
	wire _w2314_ ;
	wire _w2313_ ;
	wire _w2312_ ;
	wire _w2311_ ;
	wire _w2310_ ;
	wire _w2309_ ;
	wire _w2308_ ;
	wire _w2307_ ;
	wire _w2306_ ;
	wire _w2305_ ;
	wire _w2304_ ;
	wire _w2303_ ;
	wire _w2302_ ;
	wire _w2301_ ;
	wire _w2300_ ;
	wire _w2299_ ;
	wire _w2298_ ;
	wire _w2297_ ;
	wire _w2296_ ;
	wire _w2295_ ;
	wire _w2294_ ;
	wire _w2293_ ;
	wire _w2292_ ;
	wire _w2291_ ;
	wire _w2290_ ;
	wire _w2289_ ;
	wire _w2288_ ;
	wire _w2287_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2269_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2250_ ;
	wire _w2249_ ;
	wire _w2248_ ;
	wire _w2247_ ;
	wire _w2246_ ;
	wire _w2245_ ;
	wire _w2244_ ;
	wire _w2243_ ;
	wire _w2242_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2239_ ;
	wire _w2238_ ;
	wire _w2237_ ;
	wire _w2236_ ;
	wire _w2235_ ;
	wire _w2234_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2123_ ;
	wire _w2122_ ;
	wire _w2121_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1757_ ;
	wire _w1756_ ;
	wire _w1755_ ;
	wire _w1754_ ;
	wire _w1753_ ;
	wire _w1752_ ;
	wire _w1751_ ;
	wire _w1750_ ;
	wire _w1749_ ;
	wire _w1748_ ;
	wire _w1747_ ;
	wire _w1746_ ;
	wire _w1745_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1721_ ;
	wire _w1720_ ;
	wire _w1719_ ;
	wire _w1718_ ;
	wire _w1717_ ;
	wire _w1716_ ;
	wire _w1715_ ;
	wire _w1714_ ;
	wire _w1713_ ;
	wire _w1712_ ;
	wire _w1711_ ;
	wire _w1710_ ;
	wire _w1709_ ;
	wire _w1708_ ;
	wire _w1707_ ;
	wire _w1706_ ;
	wire _w1705_ ;
	wire _w1704_ ;
	wire _w1703_ ;
	wire _w1702_ ;
	wire _w1701_ ;
	wire _w1700_ ;
	wire _w1699_ ;
	wire _w1698_ ;
	wire _w1697_ ;
	wire _w1696_ ;
	wire _w1695_ ;
	wire _w1694_ ;
	wire _w1693_ ;
	wire _w1692_ ;
	wire _w1691_ ;
	wire _w1690_ ;
	wire _w1689_ ;
	wire _w1688_ ;
	wire _w1687_ ;
	wire _w1686_ ;
	wire _w1685_ ;
	wire _w1684_ ;
	wire _w1683_ ;
	wire _w1682_ ;
	wire _w1681_ ;
	wire _w1680_ ;
	wire _w1679_ ;
	wire _w1678_ ;
	wire _w1677_ ;
	wire _w1676_ ;
	wire _w1675_ ;
	wire _w1674_ ;
	wire _w1673_ ;
	wire _w1672_ ;
	wire _w1671_ ;
	wire _w1670_ ;
	wire _w1669_ ;
	wire _w1668_ ;
	wire _w1667_ ;
	wire _w1666_ ;
	wire _w1665_ ;
	wire _w1664_ ;
	wire _w1663_ ;
	wire _w1662_ ;
	wire _w1661_ ;
	wire _w1660_ ;
	wire _w1659_ ;
	wire _w1658_ ;
	wire _w1657_ ;
	wire _w1656_ ;
	wire _w1655_ ;
	wire _w1654_ ;
	wire _w1653_ ;
	wire _w1652_ ;
	wire _w1651_ ;
	wire _w1650_ ;
	wire _w1649_ ;
	wire _w1648_ ;
	wire _w1647_ ;
	wire _w1646_ ;
	wire _w1645_ ;
	wire _w1644_ ;
	wire _w1643_ ;
	wire _w1642_ ;
	wire _w1641_ ;
	wire _w1640_ ;
	wire _w1639_ ;
	wire _w1638_ ;
	wire _w1637_ ;
	wire _w1636_ ;
	wire _w1635_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w797_ ;
	wire _w796_ ;
	wire _w795_ ;
	wire _w794_ ;
	wire _w793_ ;
	wire _w792_ ;
	wire _w791_ ;
	wire _w790_ ;
	wire _w789_ ;
	wire _w788_ ;
	wire _w787_ ;
	wire _w786_ ;
	wire _w785_ ;
	wire _w784_ ;
	wire _w783_ ;
	wire _w782_ ;
	wire _w781_ ;
	wire _w780_ ;
	wire _w779_ ;
	wire _w778_ ;
	wire _w777_ ;
	wire _w776_ ;
	wire _w775_ ;
	wire _w774_ ;
	wire _w773_ ;
	wire _w772_ ;
	wire _w771_ ;
	wire _w640_ ;
	wire _w639_ ;
	wire _w638_ ;
	wire _w637_ ;
	wire _w636_ ;
	wire _w635_ ;
	wire _w634_ ;
	wire _w633_ ;
	wire _w632_ ;
	wire _w631_ ;
	wire _w630_ ;
	wire _w629_ ;
	wire _w628_ ;
	wire _w627_ ;
	wire _w626_ ;
	wire _w625_ ;
	wire _w624_ ;
	wire _w623_ ;
	wire _w622_ ;
	wire _w621_ ;
	wire _w620_ ;
	wire _w619_ ;
	wire _w618_ ;
	wire _w617_ ;
	wire _w616_ ;
	wire _w615_ ;
	wire _w614_ ;
	wire _w613_ ;
	wire _w612_ ;
	wire _w611_ ;
	wire _w610_ ;
	wire _w609_ ;
	wire _w608_ ;
	wire _w607_ ;
	wire _w606_ ;
	wire _w605_ ;
	wire _w604_ ;
	wire _w603_ ;
	wire _w602_ ;
	wire _w601_ ;
	wire _w600_ ;
	wire _w599_ ;
	wire _w598_ ;
	wire _w597_ ;
	wire _w596_ ;
	wire _w595_ ;
	wire _w594_ ;
	wire _w593_ ;
	wire _w592_ ;
	wire _w591_ ;
	wire _w590_ ;
	wire _w589_ ;
	wire _w588_ ;
	wire _w587_ ;
	wire _w586_ ;
	wire _w585_ ;
	wire _w584_ ;
	wire _w583_ ;
	wire _w582_ ;
	wire _w581_ ;
	wire _w580_ ;
	wire _w579_ ;
	wire _w578_ ;
	wire _w577_ ;
	wire _w576_ ;
	wire _w575_ ;
	wire _w574_ ;
	wire _w573_ ;
	wire _w542_ ;
	wire _w541_ ;
	wire _w540_ ;
	wire _w539_ ;
	wire _w538_ ;
	wire _w537_ ;
	wire _w536_ ;
	wire _w535_ ;
	wire _w534_ ;
	wire _w533_ ;
	wire _w532_ ;
	wire _w531_ ;
	wire _w530_ ;
	wire _w529_ ;
	wire _w528_ ;
	wire _w527_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w1055_ ;
	wire _w1056_ ;
	wire _w1057_ ;
	wire _w1058_ ;
	wire _w1059_ ;
	wire _w1060_ ;
	wire _w1061_ ;
	wire _w1062_ ;
	wire _w1063_ ;
	wire _w1064_ ;
	wire _w1065_ ;
	wire _w1066_ ;
	wire _w1067_ ;
	wire _w1068_ ;
	wire _w1069_ ;
	wire _w1070_ ;
	wire _w1071_ ;
	wire _w1072_ ;
	wire _w1073_ ;
	wire _w1074_ ;
	wire _w1075_ ;
	wire _w1076_ ;
	wire _w1077_ ;
	wire _w1078_ ;
	wire _w1079_ ;
	wire _w1080_ ;
	wire _w1081_ ;
	wire _w1082_ ;
	wire _w1083_ ;
	wire _w1084_ ;
	wire _w1085_ ;
	wire _w1086_ ;
	wire _w1087_ ;
	wire _w1088_ ;
	wire _w1089_ ;
	wire _w1090_ ;
	wire _w1091_ ;
	wire _w1092_ ;
	wire _w1093_ ;
	wire _w1094_ ;
	wire _w1095_ ;
	wire _w1096_ ;
	wire _w1097_ ;
	wire _w1098_ ;
	wire _w1099_ ;
	wire _w1100_ ;
	wire _w1101_ ;
	wire _w1102_ ;
	wire _w1103_ ;
	wire _w1104_ ;
	wire _w1105_ ;
	wire _w1106_ ;
	wire _w1107_ ;
	wire _w1108_ ;
	wire _w1109_ ;
	wire _w1110_ ;
	wire _w1111_ ;
	wire _w1112_ ;
	wire _w1113_ ;
	wire _w1114_ ;
	wire _w1115_ ;
	wire _w1116_ ;
	wire _w1117_ ;
	wire _w1118_ ;
	wire _w1119_ ;
	wire _w1120_ ;
	wire _w1121_ ;
	wire _w1122_ ;
	wire _w1123_ ;
	wire _w1124_ ;
	wire _w1125_ ;
	wire _w1126_ ;
	wire _w1127_ ;
	wire _w1128_ ;
	wire _w1129_ ;
	wire _w1130_ ;
	wire _w1131_ ;
	wire _w1132_ ;
	wire _w1133_ ;
	wire _w1134_ ;
	wire _w1135_ ;
	wire _w1136_ ;
	wire _w1137_ ;
	wire _w1138_ ;
	wire _w1139_ ;
	wire _w1140_ ;
	wire _w1141_ ;
	wire _w1142_ ;
	wire _w1143_ ;
	wire _w1144_ ;
	wire _w1145_ ;
	wire _w1146_ ;
	wire _w1147_ ;
	wire _w1148_ ;
	wire _w1149_ ;
	wire _w1150_ ;
	wire _w1151_ ;
	wire _w1152_ ;
	wire _w1153_ ;
	wire _w1154_ ;
	wire _w1155_ ;
	wire _w1156_ ;
	wire _w1157_ ;
	wire _w1158_ ;
	wire _w1159_ ;
	wire _w1160_ ;
	wire _w1161_ ;
	wire _w1162_ ;
	wire _w1163_ ;
	wire _w1164_ ;
	wire _w1165_ ;
	wire _w1166_ ;
	wire _w1167_ ;
	wire _w1168_ ;
	wire _w1169_ ;
	wire _w1170_ ;
	wire _w1171_ ;
	wire _w1172_ ;
	wire _w1173_ ;
	wire _w1174_ ;
	wire _w1175_ ;
	wire _w1176_ ;
	wire _w1177_ ;
	wire _w1178_ ;
	wire _w1179_ ;
	wire _w1180_ ;
	wire _w1181_ ;
	wire _w1182_ ;
	wire _w1183_ ;
	wire _w1184_ ;
	wire _w1185_ ;
	wire _w1186_ ;
	wire _w1187_ ;
	wire _w1188_ ;
	wire _w1189_ ;
	wire _w1190_ ;
	wire _w1191_ ;
	wire _w1192_ ;
	wire _w1193_ ;
	wire _w1194_ ;
	wire _w1195_ ;
	wire _w1196_ ;
	wire _w1197_ ;
	wire _w1198_ ;
	wire _w1199_ ;
	wire _w1200_ ;
	wire _w1201_ ;
	wire _w1202_ ;
	wire _w1203_ ;
	wire _w1204_ ;
	wire _w1205_ ;
	wire _w1206_ ;
	wire _w1207_ ;
	wire _w1208_ ;
	wire _w1209_ ;
	wire _w1210_ ;
	wire _w1211_ ;
	wire _w1212_ ;
	wire _w1213_ ;
	wire _w1214_ ;
	wire _w1215_ ;
	wire _w1216_ ;
	wire _w1217_ ;
	wire _w1218_ ;
	wire _w1219_ ;
	wire _w1220_ ;
	wire _w1221_ ;
	wire _w1222_ ;
	wire _w1223_ ;
	wire _w1224_ ;
	wire _w1225_ ;
	wire _w1226_ ;
	wire _w1227_ ;
	wire _w1228_ ;
	wire _w1229_ ;
	wire _w1230_ ;
	wire _w1231_ ;
	wire _w1232_ ;
	wire _w1233_ ;
	wire _w1234_ ;
	wire _w1235_ ;
	wire _w1236_ ;
	wire _w1237_ ;
	wire _w1238_ ;
	wire _w1239_ ;
	wire _w1240_ ;
	wire _w1241_ ;
	wire _w1242_ ;
	wire _w1243_ ;
	wire _w1244_ ;
	wire _w1245_ ;
	wire _w1246_ ;
	wire _w1247_ ;
	wire _w1248_ ;
	wire _w1249_ ;
	wire _w1250_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1253_ ;
	wire _w1254_ ;
	wire _w1255_ ;
	wire _w1256_ ;
	wire _w1257_ ;
	wire _w1258_ ;
	wire _w1259_ ;
	wire _w1260_ ;
	wire _w1261_ ;
	wire _w1262_ ;
	wire _w1263_ ;
	wire _w1264_ ;
	wire _w1265_ ;
	wire _w1266_ ;
	wire _w1267_ ;
	wire _w1268_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1271_ ;
	wire _w1272_ ;
	wire _w1273_ ;
	wire _w1274_ ;
	wire _w1275_ ;
	wire _w1276_ ;
	wire _w1277_ ;
	wire _w1278_ ;
	wire _w1279_ ;
	wire _w1280_ ;
	wire _w1281_ ;
	wire _w1282_ ;
	wire _w1283_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1286_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1301_ ;
	wire _w1302_ ;
	wire _w1303_ ;
	wire _w1304_ ;
	wire _w1305_ ;
	wire _w1306_ ;
	wire _w1307_ ;
	wire _w1308_ ;
	wire _w1309_ ;
	wire _w1310_ ;
	wire _w1311_ ;
	wire _w1312_ ;
	wire _w1313_ ;
	wire _w1314_ ;
	wire _w1315_ ;
	wire _w1316_ ;
	wire _w1317_ ;
	wire _w1318_ ;
	wire _w1319_ ;
	wire _w1320_ ;
	wire _w1321_ ;
	wire _w1322_ ;
	wire _w1323_ ;
	wire _w1324_ ;
	wire _w1325_ ;
	wire _w1326_ ;
	wire _w1327_ ;
	wire _w1328_ ;
	wire _w1329_ ;
	wire _w1330_ ;
	wire _w1331_ ;
	wire _w1332_ ;
	wire _w1333_ ;
	wire _w1334_ ;
	wire _w1335_ ;
	wire _w1336_ ;
	wire _w1337_ ;
	wire _w1338_ ;
	wire _w1339_ ;
	wire _w1340_ ;
	wire _w1341_ ;
	wire _w1342_ ;
	wire _w1343_ ;
	wire _w1344_ ;
	wire _w1345_ ;
	wire _w1346_ ;
	wire _w1347_ ;
	wire _w1348_ ;
	wire _w1349_ ;
	wire _w1350_ ;
	wire _w1351_ ;
	wire _w1352_ ;
	wire _w1353_ ;
	wire _w1354_ ;
	wire _w1355_ ;
	wire _w1356_ ;
	wire _w1357_ ;
	wire _w1358_ ;
	wire _w1359_ ;
	wire _w1360_ ;
	wire _w1361_ ;
	wire _w1362_ ;
	wire _w1363_ ;
	wire _w1364_ ;
	wire _w1365_ ;
	wire _w1366_ ;
	wire _w1367_ ;
	wire _w1368_ ;
	wire _w1369_ ;
	wire _w1370_ ;
	wire _w1371_ ;
	wire _w1372_ ;
	wire _w1373_ ;
	wire _w1374_ ;
	wire _w1375_ ;
	wire _w1376_ ;
	wire _w1377_ ;
	wire _w1378_ ;
	wire _w1379_ ;
	wire _w1380_ ;
	wire _w1381_ ;
	wire _w1382_ ;
	wire _w1383_ ;
	wire _w1384_ ;
	wire _w1385_ ;
	wire _w1386_ ;
	wire _w1387_ ;
	wire _w1388_ ;
	wire _w1389_ ;
	wire _w1390_ ;
	wire _w1391_ ;
	wire _w1392_ ;
	wire _w1393_ ;
	wire _w1394_ ;
	wire _w1395_ ;
	wire _w1396_ ;
	wire _w1397_ ;
	wire _w1398_ ;
	wire _w1399_ ;
	wire _w1400_ ;
	wire _w1401_ ;
	wire _w1402_ ;
	wire _w1403_ ;
	wire _w1404_ ;
	wire _w1405_ ;
	wire _w1406_ ;
	wire _w1407_ ;
	wire _w1408_ ;
	wire _w1409_ ;
	wire _w1410_ ;
	wire _w1411_ ;
	wire _w1412_ ;
	wire _w1413_ ;
	wire _w1414_ ;
	wire _w1415_ ;
	wire _w1416_ ;
	wire _w1417_ ;
	wire _w1418_ ;
	wire _w1419_ ;
	wire _w1420_ ;
	wire _w1421_ ;
	wire _w1422_ ;
	wire _w1423_ ;
	wire _w1424_ ;
	wire _w1425_ ;
	wire _w1426_ ;
	wire _w1427_ ;
	wire _w1428_ ;
	wire _w1429_ ;
	wire _w1430_ ;
	wire _w1431_ ;
	wire _w1432_ ;
	wire _w1433_ ;
	wire _w1434_ ;
	wire _w1435_ ;
	wire _w1436_ ;
	wire _w1437_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1501_ ;
	wire _w1502_ ;
	wire _w1503_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	LUT4 #(
		.INIT('h8caf)
	) name0 (
		\in2[122] ,
		\in2[123] ,
		\in3[122] ,
		\in3[123] ,
		_w514_
	);
	LUT4 #(
		.INIT('h8caf)
	) name1 (
		\in2[120] ,
		\in2[121] ,
		\in3[120] ,
		\in3[121] ,
		_w515_
	);
	LUT2 #(
		.INIT('h8)
	) name2 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h2)
	) name3 (
		\in2[127] ,
		\in3[127] ,
		_w517_
	);
	LUT4 #(
		.INIT('h8caf)
	) name4 (
		\in2[125] ,
		\in2[126] ,
		\in3[125] ,
		\in3[126] ,
		_w518_
	);
	LUT4 #(
		.INIT('hf531)
	) name5 (
		\in2[124] ,
		\in2[125] ,
		\in3[124] ,
		\in3[125] ,
		_w519_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name6 (
		\in2[126] ,
		\in2[127] ,
		\in3[126] ,
		\in3[127] ,
		_w520_
	);
	LUT4 #(
		.INIT('h0455)
	) name7 (
		_w517_,
		_w518_,
		_w519_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\in2[123] ,
		\in3[123] ,
		_w522_
	);
	LUT4 #(
		.INIT('h080a)
	) name9 (
		\in2[120] ,
		\in2[121] ,
		\in3[120] ,
		\in3[121] ,
		_w523_
	);
	LUT4 #(
		.INIT('hf531)
	) name10 (
		\in2[121] ,
		\in2[122] ,
		\in3[121] ,
		\in3[122] ,
		_w524_
	);
	LUT4 #(
		.INIT('h1311)
	) name11 (
		_w514_,
		_w522_,
		_w523_,
		_w524_,
		_w525_
	);
	LUT3 #(
		.INIT('h10)
	) name12 (
		_w516_,
		_w521_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\in2[115] ,
		\in3[115] ,
		_w527_
	);
	LUT4 #(
		.INIT('h8caf)
	) name14 (
		\in2[114] ,
		\in2[115] ,
		\in3[114] ,
		\in3[115] ,
		_w528_
	);
	LUT4 #(
		.INIT('h080a)
	) name15 (
		\in2[112] ,
		\in2[113] ,
		\in3[112] ,
		\in3[113] ,
		_w529_
	);
	LUT4 #(
		.INIT('hf531)
	) name16 (
		\in2[113] ,
		\in2[114] ,
		\in3[113] ,
		\in3[114] ,
		_w530_
	);
	LUT4 #(
		.INIT('h1511)
	) name17 (
		_w527_,
		_w528_,
		_w529_,
		_w530_,
		_w531_
	);
	LUT4 #(
		.INIT('h8caf)
	) name18 (
		\in2[118] ,
		\in2[119] ,
		\in3[118] ,
		\in3[119] ,
		_w532_
	);
	LUT4 #(
		.INIT('h8caf)
	) name19 (
		\in2[116] ,
		\in2[117] ,
		\in3[116] ,
		\in3[117] ,
		_w533_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w532_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h4)
	) name21 (
		_w531_,
		_w534_,
		_w535_
	);
	LUT4 #(
		.INIT('h8caf)
	) name22 (
		\in2[110] ,
		\in2[111] ,
		\in3[110] ,
		\in3[111] ,
		_w536_
	);
	LUT4 #(
		.INIT('h8caf)
	) name23 (
		\in2[108] ,
		\in2[109] ,
		\in3[108] ,
		\in3[109] ,
		_w537_
	);
	LUT2 #(
		.INIT('h8)
	) name24 (
		_w536_,
		_w537_,
		_w538_
	);
	LUT2 #(
		.INIT('h2)
	) name25 (
		\in2[111] ,
		\in3[111] ,
		_w539_
	);
	LUT4 #(
		.INIT('h080a)
	) name26 (
		\in2[108] ,
		\in2[109] ,
		\in3[108] ,
		\in3[109] ,
		_w540_
	);
	LUT4 #(
		.INIT('hf531)
	) name27 (
		\in2[109] ,
		\in2[110] ,
		\in3[109] ,
		\in3[110] ,
		_w541_
	);
	LUT4 #(
		.INIT('h1311)
	) name28 (
		_w536_,
		_w539_,
		_w540_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		_w538_,
		_w542_,
		_w543_
	);
	LUT4 #(
		.INIT('h8caf)
	) name30 (
		\in2[98] ,
		\in2[99] ,
		\in3[98] ,
		\in3[99] ,
		_w544_
	);
	LUT4 #(
		.INIT('h8caf)
	) name31 (
		\in2[96] ,
		\in2[97] ,
		\in3[96] ,
		\in3[97] ,
		_w545_
	);
	LUT2 #(
		.INIT('h8)
	) name32 (
		_w544_,
		_w545_,
		_w546_
	);
	LUT2 #(
		.INIT('h2)
	) name33 (
		\in2[103] ,
		\in3[103] ,
		_w547_
	);
	LUT4 #(
		.INIT('h8caf)
	) name34 (
		\in2[102] ,
		\in2[103] ,
		\in3[102] ,
		\in3[103] ,
		_w548_
	);
	LUT4 #(
		.INIT('h080a)
	) name35 (
		\in2[100] ,
		\in2[101] ,
		\in3[100] ,
		\in3[101] ,
		_w549_
	);
	LUT4 #(
		.INIT('hf531)
	) name36 (
		\in2[101] ,
		\in2[102] ,
		\in3[101] ,
		\in3[102] ,
		_w550_
	);
	LUT3 #(
		.INIT('h8a)
	) name37 (
		_w548_,
		_w549_,
		_w550_,
		_w551_
	);
	LUT4 #(
		.INIT('h1511)
	) name38 (
		_w547_,
		_w548_,
		_w549_,
		_w550_,
		_w552_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\in2[99] ,
		\in3[99] ,
		_w553_
	);
	LUT4 #(
		.INIT('h080a)
	) name40 (
		\in2[96] ,
		\in2[97] ,
		\in3[96] ,
		\in3[97] ,
		_w554_
	);
	LUT4 #(
		.INIT('hf531)
	) name41 (
		\in2[97] ,
		\in2[98] ,
		\in3[97] ,
		\in3[98] ,
		_w555_
	);
	LUT4 #(
		.INIT('h1311)
	) name42 (
		_w544_,
		_w553_,
		_w554_,
		_w555_,
		_w556_
	);
	LUT3 #(
		.INIT('h40)
	) name43 (
		_w546_,
		_w552_,
		_w556_,
		_w557_
	);
	LUT2 #(
		.INIT('h2)
	) name44 (
		\in2[91] ,
		\in3[91] ,
		_w558_
	);
	LUT4 #(
		.INIT('h8caf)
	) name45 (
		\in2[90] ,
		\in2[91] ,
		\in3[90] ,
		\in3[91] ,
		_w559_
	);
	LUT4 #(
		.INIT('h080a)
	) name46 (
		\in2[88] ,
		\in2[89] ,
		\in3[88] ,
		\in3[89] ,
		_w560_
	);
	LUT4 #(
		.INIT('hf531)
	) name47 (
		\in2[89] ,
		\in2[90] ,
		\in3[89] ,
		\in3[90] ,
		_w561_
	);
	LUT4 #(
		.INIT('h1511)
	) name48 (
		_w558_,
		_w559_,
		_w560_,
		_w561_,
		_w562_
	);
	LUT4 #(
		.INIT('h8caf)
	) name49 (
		\in2[94] ,
		\in2[95] ,
		\in3[94] ,
		\in3[95] ,
		_w563_
	);
	LUT4 #(
		.INIT('h8caf)
	) name50 (
		\in2[92] ,
		\in2[93] ,
		\in3[92] ,
		\in3[93] ,
		_w564_
	);
	LUT2 #(
		.INIT('h8)
	) name51 (
		_w563_,
		_w564_,
		_w565_
	);
	LUT2 #(
		.INIT('h4)
	) name52 (
		_w562_,
		_w565_,
		_w566_
	);
	LUT4 #(
		.INIT('h8caf)
	) name53 (
		\in2[86] ,
		\in2[87] ,
		\in3[86] ,
		\in3[87] ,
		_w567_
	);
	LUT4 #(
		.INIT('h8caf)
	) name54 (
		\in2[84] ,
		\in2[85] ,
		\in3[84] ,
		\in3[85] ,
		_w568_
	);
	LUT2 #(
		.INIT('h8)
	) name55 (
		_w567_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\in2[87] ,
		\in3[87] ,
		_w570_
	);
	LUT4 #(
		.INIT('h080a)
	) name57 (
		\in2[84] ,
		\in2[85] ,
		\in3[84] ,
		\in3[85] ,
		_w571_
	);
	LUT4 #(
		.INIT('hf531)
	) name58 (
		\in2[85] ,
		\in2[86] ,
		\in3[85] ,
		\in3[86] ,
		_w572_
	);
	LUT4 #(
		.INIT('h1311)
	) name59 (
		_w567_,
		_w570_,
		_w571_,
		_w572_,
		_w573_
	);
	LUT2 #(
		.INIT('h4)
	) name60 (
		_w569_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h2)
	) name61 (
		\in2[79] ,
		\in3[79] ,
		_w575_
	);
	LUT4 #(
		.INIT('h8caf)
	) name62 (
		\in2[78] ,
		\in2[79] ,
		\in3[78] ,
		\in3[79] ,
		_w576_
	);
	LUT4 #(
		.INIT('h080a)
	) name63 (
		\in2[76] ,
		\in2[77] ,
		\in3[76] ,
		\in3[77] ,
		_w577_
	);
	LUT4 #(
		.INIT('hf531)
	) name64 (
		\in2[77] ,
		\in2[78] ,
		\in3[77] ,
		\in3[78] ,
		_w578_
	);
	LUT4 #(
		.INIT('h1511)
	) name65 (
		_w575_,
		_w576_,
		_w577_,
		_w578_,
		_w579_
	);
	LUT4 #(
		.INIT('h8caf)
	) name66 (
		\in2[82] ,
		\in2[83] ,
		\in3[82] ,
		\in3[83] ,
		_w580_
	);
	LUT4 #(
		.INIT('h8caf)
	) name67 (
		\in2[80] ,
		\in2[81] ,
		\in3[80] ,
		\in3[81] ,
		_w581_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w580_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name69 (
		_w579_,
		_w582_,
		_w583_
	);
	LUT4 #(
		.INIT('h8caf)
	) name70 (
		\in2[74] ,
		\in2[75] ,
		\in3[74] ,
		\in3[75] ,
		_w584_
	);
	LUT4 #(
		.INIT('h8caf)
	) name71 (
		\in2[72] ,
		\in2[73] ,
		\in3[72] ,
		\in3[73] ,
		_w585_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w584_,
		_w585_,
		_w586_
	);
	LUT2 #(
		.INIT('h2)
	) name73 (
		\in2[75] ,
		\in3[75] ,
		_w587_
	);
	LUT4 #(
		.INIT('h080a)
	) name74 (
		\in2[72] ,
		\in2[73] ,
		\in3[72] ,
		\in3[73] ,
		_w588_
	);
	LUT4 #(
		.INIT('hf531)
	) name75 (
		\in2[73] ,
		\in2[74] ,
		\in3[73] ,
		\in3[74] ,
		_w589_
	);
	LUT4 #(
		.INIT('h1311)
	) name76 (
		_w584_,
		_w587_,
		_w588_,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name77 (
		_w586_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\in2[67] ,
		\in3[67] ,
		_w592_
	);
	LUT4 #(
		.INIT('h8caf)
	) name79 (
		\in2[66] ,
		\in2[67] ,
		\in3[66] ,
		\in3[67] ,
		_w593_
	);
	LUT4 #(
		.INIT('h080a)
	) name80 (
		\in2[64] ,
		\in2[65] ,
		\in3[64] ,
		\in3[65] ,
		_w594_
	);
	LUT4 #(
		.INIT('hf531)
	) name81 (
		\in2[65] ,
		\in2[66] ,
		\in3[65] ,
		\in3[66] ,
		_w595_
	);
	LUT4 #(
		.INIT('h1511)
	) name82 (
		_w592_,
		_w593_,
		_w594_,
		_w595_,
		_w596_
	);
	LUT4 #(
		.INIT('h8caf)
	) name83 (
		\in2[70] ,
		\in2[71] ,
		\in3[70] ,
		\in3[71] ,
		_w597_
	);
	LUT4 #(
		.INIT('h8caf)
	) name84 (
		\in2[68] ,
		\in2[69] ,
		\in3[68] ,
		\in3[69] ,
		_w598_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w597_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w596_,
		_w599_,
		_w600_
	);
	LUT4 #(
		.INIT('h8caf)
	) name87 (
		\in2[58] ,
		\in2[59] ,
		\in3[58] ,
		\in3[59] ,
		_w601_
	);
	LUT4 #(
		.INIT('h8caf)
	) name88 (
		\in2[60] ,
		\in2[61] ,
		\in3[60] ,
		\in3[61] ,
		_w602_
	);
	LUT4 #(
		.INIT('h8caf)
	) name89 (
		\in2[62] ,
		\in2[63] ,
		\in3[62] ,
		\in3[63] ,
		_w603_
	);
	LUT4 #(
		.INIT('h8caf)
	) name90 (
		\in2[56] ,
		\in2[57] ,
		\in3[56] ,
		\in3[57] ,
		_w604_
	);
	LUT4 #(
		.INIT('h8000)
	) name91 (
		_w601_,
		_w602_,
		_w603_,
		_w604_,
		_w605_
	);
	LUT2 #(
		.INIT('h2)
	) name92 (
		\in2[63] ,
		\in3[63] ,
		_w606_
	);
	LUT4 #(
		.INIT('h7310)
	) name93 (
		\in2[62] ,
		\in2[63] ,
		\in3[62] ,
		\in3[63] ,
		_w607_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		\in2[59] ,
		\in3[59] ,
		_w608_
	);
	LUT2 #(
		.INIT('h8)
	) name95 (
		_w602_,
		_w608_,
		_w609_
	);
	LUT4 #(
		.INIT('h080a)
	) name96 (
		\in2[56] ,
		\in2[57] ,
		\in3[56] ,
		\in3[57] ,
		_w610_
	);
	LUT4 #(
		.INIT('hf531)
	) name97 (
		\in2[57] ,
		\in2[58] ,
		\in3[57] ,
		\in3[58] ,
		_w611_
	);
	LUT4 #(
		.INIT('h8088)
	) name98 (
		_w601_,
		_w602_,
		_w610_,
		_w611_,
		_w612_
	);
	LUT4 #(
		.INIT('h080a)
	) name99 (
		\in2[60] ,
		\in2[61] ,
		\in3[60] ,
		\in3[61] ,
		_w613_
	);
	LUT4 #(
		.INIT('hf531)
	) name100 (
		\in2[61] ,
		\in2[62] ,
		\in3[61] ,
		\in3[62] ,
		_w614_
	);
	LUT3 #(
		.INIT('h10)
	) name101 (
		_w606_,
		_w613_,
		_w614_,
		_w615_
	);
	LUT4 #(
		.INIT('h5455)
	) name102 (
		_w607_,
		_w609_,
		_w612_,
		_w615_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w605_,
		_w616_,
		_w617_
	);
	LUT4 #(
		.INIT('hf531)
	) name104 (
		\in2[28] ,
		\in2[29] ,
		\in3[28] ,
		\in3[29] ,
		_w618_
	);
	LUT4 #(
		.INIT('h8caf)
	) name105 (
		\in2[27] ,
		\in2[28] ,
		\in3[27] ,
		\in3[28] ,
		_w619_
	);
	LUT2 #(
		.INIT('h2)
	) name106 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT4 #(
		.INIT('h8caf)
	) name107 (
		\in2[25] ,
		\in2[26] ,
		\in3[25] ,
		\in3[26] ,
		_w621_
	);
	LUT4 #(
		.INIT('hf531)
	) name108 (
		\in2[24] ,
		\in2[25] ,
		\in3[24] ,
		\in3[25] ,
		_w622_
	);
	LUT2 #(
		.INIT('h2)
	) name109 (
		_w621_,
		_w622_,
		_w623_
	);
	LUT4 #(
		.INIT('hf531)
	) name110 (
		\in2[22] ,
		\in2[23] ,
		\in3[22] ,
		\in3[23] ,
		_w624_
	);
	LUT4 #(
		.INIT('h8caf)
	) name111 (
		\in2[21] ,
		\in2[22] ,
		\in3[21] ,
		\in3[22] ,
		_w625_
	);
	LUT2 #(
		.INIT('h2)
	) name112 (
		_w624_,
		_w625_,
		_w626_
	);
	LUT4 #(
		.INIT('h8caf)
	) name113 (
		\in2[19] ,
		\in2[20] ,
		\in3[19] ,
		\in3[20] ,
		_w627_
	);
	LUT4 #(
		.INIT('hf531)
	) name114 (
		\in2[18] ,
		\in2[19] ,
		\in3[18] ,
		\in3[19] ,
		_w628_
	);
	LUT2 #(
		.INIT('h2)
	) name115 (
		_w627_,
		_w628_,
		_w629_
	);
	LUT4 #(
		.INIT('hf531)
	) name116 (
		\in2[16] ,
		\in2[17] ,
		\in3[16] ,
		\in3[17] ,
		_w630_
	);
	LUT4 #(
		.INIT('h8caf)
	) name117 (
		\in2[15] ,
		\in2[16] ,
		\in3[15] ,
		\in3[16] ,
		_w631_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		_w630_,
		_w631_,
		_w632_
	);
	LUT4 #(
		.INIT('h8caf)
	) name119 (
		\in2[13] ,
		\in2[14] ,
		\in3[13] ,
		\in3[14] ,
		_w633_
	);
	LUT4 #(
		.INIT('hf531)
	) name120 (
		\in2[12] ,
		\in2[13] ,
		\in3[12] ,
		\in3[13] ,
		_w634_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		_w633_,
		_w634_,
		_w635_
	);
	LUT4 #(
		.INIT('hf531)
	) name122 (
		\in2[10] ,
		\in2[11] ,
		\in3[10] ,
		\in3[11] ,
		_w636_
	);
	LUT4 #(
		.INIT('h8caf)
	) name123 (
		\in2[9] ,
		\in2[10] ,
		\in3[9] ,
		\in3[10] ,
		_w637_
	);
	LUT2 #(
		.INIT('h2)
	) name124 (
		_w636_,
		_w637_,
		_w638_
	);
	LUT4 #(
		.INIT('h8caf)
	) name125 (
		\in2[7] ,
		\in2[8] ,
		\in3[7] ,
		\in3[8] ,
		_w639_
	);
	LUT4 #(
		.INIT('hf531)
	) name126 (
		\in2[6] ,
		\in2[7] ,
		\in3[6] ,
		\in3[7] ,
		_w640_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT4 #(
		.INIT('hf531)
	) name128 (
		\in2[4] ,
		\in2[5] ,
		\in3[4] ,
		\in3[5] ,
		_w642_
	);
	LUT4 #(
		.INIT('h8caf)
	) name129 (
		\in2[3] ,
		\in2[4] ,
		\in3[3] ,
		\in3[4] ,
		_w643_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		_w642_,
		_w643_,
		_w644_
	);
	LUT4 #(
		.INIT('hf531)
	) name131 (
		\in2[0] ,
		\in2[1] ,
		\in3[0] ,
		\in3[1] ,
		_w645_
	);
	LUT4 #(
		.INIT('h8caf)
	) name132 (
		\in2[1] ,
		\in2[2] ,
		\in3[1] ,
		\in3[2] ,
		_w646_
	);
	LUT4 #(
		.INIT('hf531)
	) name133 (
		\in2[2] ,
		\in2[3] ,
		\in3[2] ,
		\in3[3] ,
		_w647_
	);
	LUT4 #(
		.INIT('h8a00)
	) name134 (
		_w642_,
		_w645_,
		_w646_,
		_w647_,
		_w648_
	);
	LUT4 #(
		.INIT('h8caf)
	) name135 (
		\in2[5] ,
		\in2[6] ,
		\in3[5] ,
		\in3[6] ,
		_w649_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w639_,
		_w649_,
		_w650_
	);
	LUT4 #(
		.INIT('h5455)
	) name137 (
		_w641_,
		_w644_,
		_w648_,
		_w650_,
		_w651_
	);
	LUT4 #(
		.INIT('hf531)
	) name138 (
		\in2[8] ,
		\in2[9] ,
		\in3[8] ,
		\in3[9] ,
		_w652_
	);
	LUT2 #(
		.INIT('h8)
	) name139 (
		_w636_,
		_w652_,
		_w653_
	);
	LUT4 #(
		.INIT('h8caf)
	) name140 (
		\in2[11] ,
		\in2[12] ,
		\in3[11] ,
		\in3[12] ,
		_w654_
	);
	LUT2 #(
		.INIT('h8)
	) name141 (
		_w633_,
		_w654_,
		_w655_
	);
	LUT4 #(
		.INIT('h1500)
	) name142 (
		_w638_,
		_w651_,
		_w653_,
		_w655_,
		_w656_
	);
	LUT4 #(
		.INIT('hf531)
	) name143 (
		\in2[14] ,
		\in2[15] ,
		\in3[14] ,
		\in3[15] ,
		_w657_
	);
	LUT2 #(
		.INIT('h8)
	) name144 (
		_w630_,
		_w657_,
		_w658_
	);
	LUT4 #(
		.INIT('h5455)
	) name145 (
		_w632_,
		_w635_,
		_w656_,
		_w658_,
		_w659_
	);
	LUT4 #(
		.INIT('h8caf)
	) name146 (
		\in2[17] ,
		\in2[18] ,
		\in3[17] ,
		\in3[18] ,
		_w660_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		_w627_,
		_w660_,
		_w661_
	);
	LUT4 #(
		.INIT('hf531)
	) name148 (
		\in2[20] ,
		\in2[21] ,
		\in3[20] ,
		\in3[21] ,
		_w662_
	);
	LUT2 #(
		.INIT('h8)
	) name149 (
		_w624_,
		_w662_,
		_w663_
	);
	LUT4 #(
		.INIT('h1500)
	) name150 (
		_w629_,
		_w659_,
		_w661_,
		_w663_,
		_w664_
	);
	LUT4 #(
		.INIT('h8caf)
	) name151 (
		\in2[23] ,
		\in2[24] ,
		\in3[23] ,
		\in3[24] ,
		_w665_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w621_,
		_w665_,
		_w666_
	);
	LUT4 #(
		.INIT('h5455)
	) name153 (
		_w623_,
		_w626_,
		_w664_,
		_w666_,
		_w667_
	);
	LUT4 #(
		.INIT('hf531)
	) name154 (
		\in2[26] ,
		\in2[27] ,
		\in3[26] ,
		\in3[27] ,
		_w668_
	);
	LUT2 #(
		.INIT('h8)
	) name155 (
		_w618_,
		_w668_,
		_w669_
	);
	LUT2 #(
		.INIT('h4)
	) name156 (
		\in2[31] ,
		\in3[31] ,
		_w670_
	);
	LUT4 #(
		.INIT('h8caf)
	) name157 (
		\in2[32] ,
		\in2[33] ,
		\in3[32] ,
		\in3[33] ,
		_w671_
	);
	LUT4 #(
		.INIT('h8caf)
	) name158 (
		\in2[34] ,
		\in2[35] ,
		\in3[34] ,
		\in3[35] ,
		_w672_
	);
	LUT4 #(
		.INIT('h8caf)
	) name159 (
		\in2[38] ,
		\in2[39] ,
		\in3[38] ,
		\in3[39] ,
		_w673_
	);
	LUT4 #(
		.INIT('h4000)
	) name160 (
		_w670_,
		_w671_,
		_w672_,
		_w673_,
		_w674_
	);
	LUT4 #(
		.INIT('h8caf)
	) name161 (
		\in2[36] ,
		\in2[37] ,
		\in3[36] ,
		\in3[37] ,
		_w675_
	);
	LUT4 #(
		.INIT('h8caf)
	) name162 (
		\in2[29] ,
		\in2[30] ,
		\in3[29] ,
		\in3[30] ,
		_w676_
	);
	LUT2 #(
		.INIT('h8)
	) name163 (
		_w675_,
		_w676_,
		_w677_
	);
	LUT2 #(
		.INIT('h8)
	) name164 (
		_w674_,
		_w677_,
		_w678_
	);
	LUT4 #(
		.INIT('h1500)
	) name165 (
		_w620_,
		_w667_,
		_w669_,
		_w678_,
		_w679_
	);
	LUT4 #(
		.INIT('hf531)
	) name166 (
		\in2[30] ,
		\in2[31] ,
		\in3[30] ,
		\in3[31] ,
		_w680_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		_w675_,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h8)
	) name168 (
		_w674_,
		_w681_,
		_w682_
	);
	LUT4 #(
		.INIT('h8caf)
	) name169 (
		\in2[46] ,
		\in2[47] ,
		\in3[46] ,
		\in3[47] ,
		_w683_
	);
	LUT2 #(
		.INIT('h2)
	) name170 (
		\in2[47] ,
		\in3[47] ,
		_w684_
	);
	LUT4 #(
		.INIT('h7310)
	) name171 (
		\in2[46] ,
		\in2[47] ,
		\in3[46] ,
		\in3[47] ,
		_w685_
	);
	LUT4 #(
		.INIT('h8caf)
	) name172 (
		\in2[44] ,
		\in2[45] ,
		\in3[44] ,
		\in3[45] ,
		_w686_
	);
	LUT2 #(
		.INIT('h2)
	) name173 (
		\in2[43] ,
		\in3[43] ,
		_w687_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		_w686_,
		_w687_,
		_w688_
	);
	LUT4 #(
		.INIT('h8caf)
	) name175 (
		\in2[42] ,
		\in2[43] ,
		\in3[42] ,
		\in3[43] ,
		_w689_
	);
	LUT4 #(
		.INIT('h080a)
	) name176 (
		\in2[40] ,
		\in2[41] ,
		\in3[40] ,
		\in3[41] ,
		_w690_
	);
	LUT4 #(
		.INIT('hf531)
	) name177 (
		\in2[41] ,
		\in2[42] ,
		\in3[41] ,
		\in3[42] ,
		_w691_
	);
	LUT4 #(
		.INIT('h8088)
	) name178 (
		_w686_,
		_w689_,
		_w690_,
		_w691_,
		_w692_
	);
	LUT4 #(
		.INIT('h080a)
	) name179 (
		\in2[44] ,
		\in2[45] ,
		\in3[44] ,
		\in3[45] ,
		_w693_
	);
	LUT4 #(
		.INIT('hf531)
	) name180 (
		\in2[45] ,
		\in2[46] ,
		\in3[45] ,
		\in3[46] ,
		_w694_
	);
	LUT3 #(
		.INIT('h10)
	) name181 (
		_w684_,
		_w693_,
		_w694_,
		_w695_
	);
	LUT4 #(
		.INIT('h5455)
	) name182 (
		_w685_,
		_w688_,
		_w692_,
		_w695_,
		_w696_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		\in2[39] ,
		\in3[39] ,
		_w697_
	);
	LUT4 #(
		.INIT('h7310)
	) name184 (
		\in2[38] ,
		\in2[39] ,
		\in3[38] ,
		\in3[39] ,
		_w698_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\in2[35] ,
		\in3[35] ,
		_w699_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		_w675_,
		_w699_,
		_w700_
	);
	LUT4 #(
		.INIT('h080a)
	) name187 (
		\in2[32] ,
		\in2[33] ,
		\in3[32] ,
		\in3[33] ,
		_w701_
	);
	LUT4 #(
		.INIT('hf531)
	) name188 (
		\in2[33] ,
		\in2[34] ,
		\in3[33] ,
		\in3[34] ,
		_w702_
	);
	LUT4 #(
		.INIT('h8088)
	) name189 (
		_w672_,
		_w675_,
		_w701_,
		_w702_,
		_w703_
	);
	LUT4 #(
		.INIT('h080a)
	) name190 (
		\in2[36] ,
		\in2[37] ,
		\in3[36] ,
		\in3[37] ,
		_w704_
	);
	LUT4 #(
		.INIT('hf531)
	) name191 (
		\in2[37] ,
		\in2[38] ,
		\in3[37] ,
		\in3[38] ,
		_w705_
	);
	LUT3 #(
		.INIT('h10)
	) name192 (
		_w697_,
		_w704_,
		_w705_,
		_w706_
	);
	LUT4 #(
		.INIT('h5455)
	) name193 (
		_w698_,
		_w700_,
		_w703_,
		_w706_,
		_w707_
	);
	LUT3 #(
		.INIT('h01)
	) name194 (
		_w682_,
		_w696_,
		_w707_,
		_w708_
	);
	LUT4 #(
		.INIT('h8caf)
	) name195 (
		\in2[40] ,
		\in2[41] ,
		\in3[40] ,
		\in3[41] ,
		_w709_
	);
	LUT4 #(
		.INIT('h8000)
	) name196 (
		_w683_,
		_w686_,
		_w689_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h2)
	) name197 (
		_w685_,
		_w710_,
		_w711_
	);
	LUT4 #(
		.INIT('h0010)
	) name198 (
		_w688_,
		_w692_,
		_w695_,
		_w710_,
		_w712_
	);
	LUT4 #(
		.INIT('h8caf)
	) name199 (
		\in2[52] ,
		\in2[53] ,
		\in3[52] ,
		\in3[53] ,
		_w713_
	);
	LUT4 #(
		.INIT('h8caf)
	) name200 (
		\in2[50] ,
		\in2[51] ,
		\in3[50] ,
		\in3[51] ,
		_w714_
	);
	LUT4 #(
		.INIT('h8caf)
	) name201 (
		\in2[54] ,
		\in2[55] ,
		\in3[54] ,
		\in3[55] ,
		_w715_
	);
	LUT4 #(
		.INIT('h8caf)
	) name202 (
		\in2[48] ,
		\in2[49] ,
		\in3[48] ,
		\in3[49] ,
		_w716_
	);
	LUT4 #(
		.INIT('h8000)
	) name203 (
		_w713_,
		_w714_,
		_w715_,
		_w716_,
		_w717_
	);
	LUT3 #(
		.INIT('h10)
	) name204 (
		_w711_,
		_w712_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h2)
	) name205 (
		\in2[55] ,
		\in3[55] ,
		_w719_
	);
	LUT4 #(
		.INIT('h7310)
	) name206 (
		\in2[54] ,
		\in2[55] ,
		\in3[54] ,
		\in3[55] ,
		_w720_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		\in2[51] ,
		\in3[51] ,
		_w721_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		_w713_,
		_w721_,
		_w722_
	);
	LUT4 #(
		.INIT('h080a)
	) name209 (
		\in2[48] ,
		\in2[49] ,
		\in3[48] ,
		\in3[49] ,
		_w723_
	);
	LUT4 #(
		.INIT('hf531)
	) name210 (
		\in2[49] ,
		\in2[50] ,
		\in3[49] ,
		\in3[50] ,
		_w724_
	);
	LUT4 #(
		.INIT('h8088)
	) name211 (
		_w713_,
		_w714_,
		_w723_,
		_w724_,
		_w725_
	);
	LUT4 #(
		.INIT('h080a)
	) name212 (
		\in2[52] ,
		\in2[53] ,
		\in3[52] ,
		\in3[53] ,
		_w726_
	);
	LUT4 #(
		.INIT('hf531)
	) name213 (
		\in2[53] ,
		\in2[54] ,
		\in3[53] ,
		\in3[54] ,
		_w727_
	);
	LUT3 #(
		.INIT('h10)
	) name214 (
		_w719_,
		_w726_,
		_w727_,
		_w728_
	);
	LUT4 #(
		.INIT('h5455)
	) name215 (
		_w720_,
		_w722_,
		_w725_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w616_,
		_w729_,
		_w730_
	);
	LUT4 #(
		.INIT('h4f00)
	) name217 (
		_w679_,
		_w708_,
		_w718_,
		_w730_,
		_w731_
	);
	LUT4 #(
		.INIT('h8caf)
	) name218 (
		\in2[64] ,
		\in2[65] ,
		\in3[64] ,
		\in3[65] ,
		_w732_
	);
	LUT4 #(
		.INIT('h8000)
	) name219 (
		_w593_,
		_w597_,
		_w598_,
		_w732_,
		_w733_
	);
	LUT4 #(
		.INIT('h5455)
	) name220 (
		_w600_,
		_w617_,
		_w731_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h2)
	) name221 (
		\in2[71] ,
		\in3[71] ,
		_w735_
	);
	LUT4 #(
		.INIT('h080a)
	) name222 (
		\in2[68] ,
		\in2[69] ,
		\in3[68] ,
		\in3[69] ,
		_w736_
	);
	LUT4 #(
		.INIT('hf531)
	) name223 (
		\in2[69] ,
		\in2[70] ,
		\in3[69] ,
		\in3[70] ,
		_w737_
	);
	LUT4 #(
		.INIT('h1311)
	) name224 (
		_w597_,
		_w735_,
		_w736_,
		_w737_,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name225 (
		_w590_,
		_w738_,
		_w739_
	);
	LUT4 #(
		.INIT('h8caf)
	) name226 (
		\in2[76] ,
		\in2[77] ,
		\in3[76] ,
		\in3[77] ,
		_w740_
	);
	LUT4 #(
		.INIT('h8000)
	) name227 (
		_w576_,
		_w580_,
		_w581_,
		_w740_,
		_w741_
	);
	LUT4 #(
		.INIT('h1500)
	) name228 (
		_w591_,
		_w734_,
		_w739_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h2)
	) name229 (
		\in2[83] ,
		\in3[83] ,
		_w743_
	);
	LUT4 #(
		.INIT('h080a)
	) name230 (
		\in2[80] ,
		\in2[81] ,
		\in3[80] ,
		\in3[81] ,
		_w744_
	);
	LUT4 #(
		.INIT('hf531)
	) name231 (
		\in2[81] ,
		\in2[82] ,
		\in3[81] ,
		\in3[82] ,
		_w745_
	);
	LUT4 #(
		.INIT('h1311)
	) name232 (
		_w580_,
		_w743_,
		_w744_,
		_w745_,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name233 (
		_w573_,
		_w746_,
		_w747_
	);
	LUT4 #(
		.INIT('h5455)
	) name234 (
		_w574_,
		_w583_,
		_w742_,
		_w747_,
		_w748_
	);
	LUT4 #(
		.INIT('h8caf)
	) name235 (
		\in2[88] ,
		\in2[89] ,
		\in3[88] ,
		\in3[89] ,
		_w749_
	);
	LUT4 #(
		.INIT('h8000)
	) name236 (
		_w559_,
		_w563_,
		_w564_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h2)
	) name237 (
		\in2[95] ,
		\in3[95] ,
		_w751_
	);
	LUT4 #(
		.INIT('h080a)
	) name238 (
		\in2[92] ,
		\in2[93] ,
		\in3[92] ,
		\in3[93] ,
		_w752_
	);
	LUT4 #(
		.INIT('hf531)
	) name239 (
		\in2[93] ,
		\in2[94] ,
		\in3[93] ,
		\in3[94] ,
		_w753_
	);
	LUT4 #(
		.INIT('h1311)
	) name240 (
		_w563_,
		_w751_,
		_w752_,
		_w753_,
		_w754_
	);
	LUT3 #(
		.INIT('h80)
	) name241 (
		_w552_,
		_w556_,
		_w754_,
		_w755_
	);
	LUT4 #(
		.INIT('h1500)
	) name242 (
		_w566_,
		_w748_,
		_w750_,
		_w755_,
		_w756_
	);
	LUT4 #(
		.INIT('h8caf)
	) name243 (
		\in2[100] ,
		\in2[101] ,
		\in3[100] ,
		\in3[101] ,
		_w757_
	);
	LUT3 #(
		.INIT('h15)
	) name244 (
		_w547_,
		_w548_,
		_w757_,
		_w758_
	);
	LUT4 #(
		.INIT('h8caf)
	) name245 (
		\in2[106] ,
		\in2[107] ,
		\in3[106] ,
		\in3[107] ,
		_w759_
	);
	LUT4 #(
		.INIT('h8caf)
	) name246 (
		\in2[104] ,
		\in2[105] ,
		\in3[104] ,
		\in3[105] ,
		_w760_
	);
	LUT2 #(
		.INIT('h8)
	) name247 (
		_w759_,
		_w760_,
		_w761_
	);
	LUT3 #(
		.INIT('hb0)
	) name248 (
		_w551_,
		_w758_,
		_w761_,
		_w762_
	);
	LUT2 #(
		.INIT('h2)
	) name249 (
		\in2[107] ,
		\in3[107] ,
		_w763_
	);
	LUT4 #(
		.INIT('h080a)
	) name250 (
		\in2[104] ,
		\in2[105] ,
		\in3[104] ,
		\in3[105] ,
		_w764_
	);
	LUT4 #(
		.INIT('hf531)
	) name251 (
		\in2[105] ,
		\in2[106] ,
		\in3[105] ,
		\in3[106] ,
		_w765_
	);
	LUT4 #(
		.INIT('h1311)
	) name252 (
		_w759_,
		_w763_,
		_w764_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h8)
	) name253 (
		_w542_,
		_w766_,
		_w767_
	);
	LUT4 #(
		.INIT('hef00)
	) name254 (
		_w557_,
		_w756_,
		_w762_,
		_w767_,
		_w768_
	);
	LUT4 #(
		.INIT('h8caf)
	) name255 (
		\in2[112] ,
		\in2[113] ,
		\in3[112] ,
		\in3[113] ,
		_w769_
	);
	LUT4 #(
		.INIT('h8000)
	) name256 (
		_w528_,
		_w532_,
		_w533_,
		_w769_,
		_w770_
	);
	LUT4 #(
		.INIT('h5455)
	) name257 (
		_w535_,
		_w543_,
		_w768_,
		_w770_,
		_w771_
	);
	LUT2 #(
		.INIT('h2)
	) name258 (
		\in2[119] ,
		\in3[119] ,
		_w772_
	);
	LUT4 #(
		.INIT('h080a)
	) name259 (
		\in2[116] ,
		\in2[117] ,
		\in3[116] ,
		\in3[117] ,
		_w773_
	);
	LUT4 #(
		.INIT('hf531)
	) name260 (
		\in2[117] ,
		\in2[118] ,
		\in3[117] ,
		\in3[118] ,
		_w774_
	);
	LUT4 #(
		.INIT('h1311)
	) name261 (
		_w532_,
		_w772_,
		_w773_,
		_w774_,
		_w775_
	);
	LUT3 #(
		.INIT('h40)
	) name262 (
		_w521_,
		_w525_,
		_w775_,
		_w776_
	);
	LUT4 #(
		.INIT('haf23)
	) name263 (
		\in2[124] ,
		\in2[127] ,
		\in3[124] ,
		\in3[127] ,
		_w777_
	);
	LUT2 #(
		.INIT('h8)
	) name264 (
		_w518_,
		_w777_,
		_w778_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		_w521_,
		_w778_,
		_w779_
	);
	LUT3 #(
		.INIT('ha8)
	) name266 (
		\in2[0] ,
		_w521_,
		_w778_,
		_w780_
	);
	LUT4 #(
		.INIT('h1500)
	) name267 (
		_w526_,
		_w771_,
		_w776_,
		_w780_,
		_w781_
	);
	LUT4 #(
		.INIT('h0015)
	) name268 (
		_w526_,
		_w771_,
		_w776_,
		_w779_,
		_w782_
	);
	LUT3 #(
		.INIT('h31)
	) name269 (
		\in3[0] ,
		_w781_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h2)
	) name270 (
		\in0[115] ,
		\in1[115] ,
		_w784_
	);
	LUT4 #(
		.INIT('h8caf)
	) name271 (
		\in0[114] ,
		\in0[115] ,
		\in1[114] ,
		\in1[115] ,
		_w785_
	);
	LUT4 #(
		.INIT('h080a)
	) name272 (
		\in0[112] ,
		\in0[113] ,
		\in1[112] ,
		\in1[113] ,
		_w786_
	);
	LUT4 #(
		.INIT('hf531)
	) name273 (
		\in0[113] ,
		\in0[114] ,
		\in1[113] ,
		\in1[114] ,
		_w787_
	);
	LUT4 #(
		.INIT('h1511)
	) name274 (
		_w784_,
		_w785_,
		_w786_,
		_w787_,
		_w788_
	);
	LUT4 #(
		.INIT('h8caf)
	) name275 (
		\in0[116] ,
		\in0[117] ,
		\in1[116] ,
		\in1[117] ,
		_w789_
	);
	LUT2 #(
		.INIT('h4)
	) name276 (
		_w788_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h2)
	) name277 (
		\in0[79] ,
		\in1[79] ,
		_w791_
	);
	LUT4 #(
		.INIT('h8caf)
	) name278 (
		\in0[78] ,
		\in0[79] ,
		\in1[78] ,
		\in1[79] ,
		_w792_
	);
	LUT4 #(
		.INIT('h080a)
	) name279 (
		\in0[76] ,
		\in0[77] ,
		\in1[76] ,
		\in1[77] ,
		_w793_
	);
	LUT4 #(
		.INIT('hf531)
	) name280 (
		\in0[77] ,
		\in0[78] ,
		\in1[77] ,
		\in1[78] ,
		_w794_
	);
	LUT4 #(
		.INIT('h1511)
	) name281 (
		_w791_,
		_w792_,
		_w793_,
		_w794_,
		_w795_
	);
	LUT4 #(
		.INIT('h8caf)
	) name282 (
		\in0[80] ,
		\in0[81] ,
		\in1[80] ,
		\in1[81] ,
		_w796_
	);
	LUT2 #(
		.INIT('h4)
	) name283 (
		_w795_,
		_w796_,
		_w797_
	);
	LUT4 #(
		.INIT('h8caf)
	) name284 (
		\in0[74] ,
		\in0[75] ,
		\in1[74] ,
		\in1[75] ,
		_w798_
	);
	LUT4 #(
		.INIT('h8caf)
	) name285 (
		\in0[72] ,
		\in0[73] ,
		\in1[72] ,
		\in1[73] ,
		_w799_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		_w798_,
		_w799_,
		_w800_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		\in0[75] ,
		\in1[75] ,
		_w801_
	);
	LUT4 #(
		.INIT('h080a)
	) name288 (
		\in0[72] ,
		\in0[73] ,
		\in1[72] ,
		\in1[73] ,
		_w802_
	);
	LUT4 #(
		.INIT('hf531)
	) name289 (
		\in0[73] ,
		\in0[74] ,
		\in1[73] ,
		\in1[74] ,
		_w803_
	);
	LUT4 #(
		.INIT('h1311)
	) name290 (
		_w798_,
		_w801_,
		_w802_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		_w800_,
		_w804_,
		_w805_
	);
	LUT2 #(
		.INIT('h2)
	) name292 (
		\in0[67] ,
		\in1[67] ,
		_w806_
	);
	LUT4 #(
		.INIT('h8caf)
	) name293 (
		\in0[66] ,
		\in0[67] ,
		\in1[66] ,
		\in1[67] ,
		_w807_
	);
	LUT4 #(
		.INIT('h080a)
	) name294 (
		\in0[64] ,
		\in0[65] ,
		\in1[64] ,
		\in1[65] ,
		_w808_
	);
	LUT4 #(
		.INIT('hf531)
	) name295 (
		\in0[65] ,
		\in0[66] ,
		\in1[65] ,
		\in1[66] ,
		_w809_
	);
	LUT4 #(
		.INIT('h1511)
	) name296 (
		_w806_,
		_w807_,
		_w808_,
		_w809_,
		_w810_
	);
	LUT4 #(
		.INIT('h8caf)
	) name297 (
		\in0[70] ,
		\in0[71] ,
		\in1[70] ,
		\in1[71] ,
		_w811_
	);
	LUT4 #(
		.INIT('h8caf)
	) name298 (
		\in0[68] ,
		\in0[69] ,
		\in1[68] ,
		\in1[69] ,
		_w812_
	);
	LUT2 #(
		.INIT('h8)
	) name299 (
		_w811_,
		_w812_,
		_w813_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		_w810_,
		_w813_,
		_w814_
	);
	LUT4 #(
		.INIT('hf531)
	) name301 (
		\in0[28] ,
		\in0[29] ,
		\in1[28] ,
		\in1[29] ,
		_w815_
	);
	LUT4 #(
		.INIT('h8caf)
	) name302 (
		\in0[27] ,
		\in0[28] ,
		\in1[27] ,
		\in1[28] ,
		_w816_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		_w815_,
		_w816_,
		_w817_
	);
	LUT4 #(
		.INIT('h8caf)
	) name304 (
		\in0[25] ,
		\in0[26] ,
		\in1[25] ,
		\in1[26] ,
		_w818_
	);
	LUT4 #(
		.INIT('hf531)
	) name305 (
		\in0[24] ,
		\in0[25] ,
		\in1[24] ,
		\in1[25] ,
		_w819_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		_w818_,
		_w819_,
		_w820_
	);
	LUT4 #(
		.INIT('hf531)
	) name307 (
		\in0[22] ,
		\in0[23] ,
		\in1[22] ,
		\in1[23] ,
		_w821_
	);
	LUT4 #(
		.INIT('h8caf)
	) name308 (
		\in0[21] ,
		\in0[22] ,
		\in1[21] ,
		\in1[22] ,
		_w822_
	);
	LUT2 #(
		.INIT('h2)
	) name309 (
		_w821_,
		_w822_,
		_w823_
	);
	LUT4 #(
		.INIT('h8caf)
	) name310 (
		\in0[19] ,
		\in0[20] ,
		\in1[19] ,
		\in1[20] ,
		_w824_
	);
	LUT4 #(
		.INIT('hf531)
	) name311 (
		\in0[18] ,
		\in0[19] ,
		\in1[18] ,
		\in1[19] ,
		_w825_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		_w824_,
		_w825_,
		_w826_
	);
	LUT4 #(
		.INIT('hf531)
	) name313 (
		\in0[16] ,
		\in0[17] ,
		\in1[16] ,
		\in1[17] ,
		_w827_
	);
	LUT4 #(
		.INIT('h8caf)
	) name314 (
		\in0[15] ,
		\in0[16] ,
		\in1[15] ,
		\in1[16] ,
		_w828_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		_w827_,
		_w828_,
		_w829_
	);
	LUT4 #(
		.INIT('h8caf)
	) name316 (
		\in0[13] ,
		\in0[14] ,
		\in1[13] ,
		\in1[14] ,
		_w830_
	);
	LUT4 #(
		.INIT('hf531)
	) name317 (
		\in0[12] ,
		\in0[13] ,
		\in1[12] ,
		\in1[13] ,
		_w831_
	);
	LUT2 #(
		.INIT('h2)
	) name318 (
		_w830_,
		_w831_,
		_w832_
	);
	LUT4 #(
		.INIT('hf531)
	) name319 (
		\in0[10] ,
		\in0[11] ,
		\in1[10] ,
		\in1[11] ,
		_w833_
	);
	LUT4 #(
		.INIT('h8caf)
	) name320 (
		\in0[9] ,
		\in0[10] ,
		\in1[9] ,
		\in1[10] ,
		_w834_
	);
	LUT2 #(
		.INIT('h2)
	) name321 (
		_w833_,
		_w834_,
		_w835_
	);
	LUT4 #(
		.INIT('h8caf)
	) name322 (
		\in0[7] ,
		\in0[8] ,
		\in1[7] ,
		\in1[8] ,
		_w836_
	);
	LUT4 #(
		.INIT('hf531)
	) name323 (
		\in0[6] ,
		\in0[7] ,
		\in1[6] ,
		\in1[7] ,
		_w837_
	);
	LUT2 #(
		.INIT('h2)
	) name324 (
		_w836_,
		_w837_,
		_w838_
	);
	LUT4 #(
		.INIT('hf531)
	) name325 (
		\in0[4] ,
		\in0[5] ,
		\in1[4] ,
		\in1[5] ,
		_w839_
	);
	LUT4 #(
		.INIT('h8caf)
	) name326 (
		\in0[3] ,
		\in0[4] ,
		\in1[3] ,
		\in1[4] ,
		_w840_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		_w839_,
		_w840_,
		_w841_
	);
	LUT4 #(
		.INIT('hf531)
	) name328 (
		\in0[0] ,
		\in0[1] ,
		\in1[0] ,
		\in1[1] ,
		_w842_
	);
	LUT4 #(
		.INIT('h8caf)
	) name329 (
		\in0[1] ,
		\in0[2] ,
		\in1[1] ,
		\in1[2] ,
		_w843_
	);
	LUT4 #(
		.INIT('hf531)
	) name330 (
		\in0[2] ,
		\in0[3] ,
		\in1[2] ,
		\in1[3] ,
		_w844_
	);
	LUT4 #(
		.INIT('h8a00)
	) name331 (
		_w839_,
		_w842_,
		_w843_,
		_w844_,
		_w845_
	);
	LUT4 #(
		.INIT('h8caf)
	) name332 (
		\in0[5] ,
		\in0[6] ,
		\in1[5] ,
		\in1[6] ,
		_w846_
	);
	LUT2 #(
		.INIT('h8)
	) name333 (
		_w836_,
		_w846_,
		_w847_
	);
	LUT4 #(
		.INIT('h5455)
	) name334 (
		_w838_,
		_w841_,
		_w845_,
		_w847_,
		_w848_
	);
	LUT4 #(
		.INIT('hf531)
	) name335 (
		\in0[8] ,
		\in0[9] ,
		\in1[8] ,
		\in1[9] ,
		_w849_
	);
	LUT2 #(
		.INIT('h8)
	) name336 (
		_w833_,
		_w849_,
		_w850_
	);
	LUT4 #(
		.INIT('h8caf)
	) name337 (
		\in0[11] ,
		\in0[12] ,
		\in1[11] ,
		\in1[12] ,
		_w851_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w830_,
		_w851_,
		_w852_
	);
	LUT4 #(
		.INIT('h1500)
	) name339 (
		_w835_,
		_w848_,
		_w850_,
		_w852_,
		_w853_
	);
	LUT4 #(
		.INIT('hf531)
	) name340 (
		\in0[14] ,
		\in0[15] ,
		\in1[14] ,
		\in1[15] ,
		_w854_
	);
	LUT2 #(
		.INIT('h8)
	) name341 (
		_w827_,
		_w854_,
		_w855_
	);
	LUT4 #(
		.INIT('h5455)
	) name342 (
		_w829_,
		_w832_,
		_w853_,
		_w855_,
		_w856_
	);
	LUT4 #(
		.INIT('h8caf)
	) name343 (
		\in0[17] ,
		\in0[18] ,
		\in1[17] ,
		\in1[18] ,
		_w857_
	);
	LUT2 #(
		.INIT('h8)
	) name344 (
		_w824_,
		_w857_,
		_w858_
	);
	LUT4 #(
		.INIT('hf531)
	) name345 (
		\in0[20] ,
		\in0[21] ,
		\in1[20] ,
		\in1[21] ,
		_w859_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		_w821_,
		_w859_,
		_w860_
	);
	LUT4 #(
		.INIT('h1500)
	) name347 (
		_w826_,
		_w856_,
		_w858_,
		_w860_,
		_w861_
	);
	LUT4 #(
		.INIT('h8caf)
	) name348 (
		\in0[23] ,
		\in0[24] ,
		\in1[23] ,
		\in1[24] ,
		_w862_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		_w818_,
		_w862_,
		_w863_
	);
	LUT4 #(
		.INIT('h5455)
	) name350 (
		_w820_,
		_w823_,
		_w861_,
		_w863_,
		_w864_
	);
	LUT4 #(
		.INIT('hf531)
	) name351 (
		\in0[26] ,
		\in0[27] ,
		\in1[26] ,
		\in1[27] ,
		_w865_
	);
	LUT2 #(
		.INIT('h8)
	) name352 (
		_w815_,
		_w865_,
		_w866_
	);
	LUT2 #(
		.INIT('h4)
	) name353 (
		\in0[31] ,
		\in1[31] ,
		_w867_
	);
	LUT4 #(
		.INIT('h8caf)
	) name354 (
		\in0[32] ,
		\in0[33] ,
		\in1[32] ,
		\in1[33] ,
		_w868_
	);
	LUT4 #(
		.INIT('h8caf)
	) name355 (
		\in0[34] ,
		\in0[35] ,
		\in1[34] ,
		\in1[35] ,
		_w869_
	);
	LUT4 #(
		.INIT('h8caf)
	) name356 (
		\in0[38] ,
		\in0[39] ,
		\in1[38] ,
		\in1[39] ,
		_w870_
	);
	LUT4 #(
		.INIT('h4000)
	) name357 (
		_w867_,
		_w868_,
		_w869_,
		_w870_,
		_w871_
	);
	LUT4 #(
		.INIT('h8caf)
	) name358 (
		\in0[36] ,
		\in0[37] ,
		\in1[36] ,
		\in1[37] ,
		_w872_
	);
	LUT4 #(
		.INIT('h8caf)
	) name359 (
		\in0[29] ,
		\in0[30] ,
		\in1[29] ,
		\in1[30] ,
		_w873_
	);
	LUT2 #(
		.INIT('h8)
	) name360 (
		_w872_,
		_w873_,
		_w874_
	);
	LUT2 #(
		.INIT('h8)
	) name361 (
		_w871_,
		_w874_,
		_w875_
	);
	LUT4 #(
		.INIT('h1500)
	) name362 (
		_w817_,
		_w864_,
		_w866_,
		_w875_,
		_w876_
	);
	LUT4 #(
		.INIT('hf531)
	) name363 (
		\in0[30] ,
		\in0[31] ,
		\in1[30] ,
		\in1[31] ,
		_w877_
	);
	LUT2 #(
		.INIT('h2)
	) name364 (
		_w872_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		_w871_,
		_w878_,
		_w879_
	);
	LUT4 #(
		.INIT('h8caf)
	) name366 (
		\in0[46] ,
		\in0[47] ,
		\in1[46] ,
		\in1[47] ,
		_w880_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		\in0[47] ,
		\in1[47] ,
		_w881_
	);
	LUT4 #(
		.INIT('h7310)
	) name368 (
		\in0[46] ,
		\in0[47] ,
		\in1[46] ,
		\in1[47] ,
		_w882_
	);
	LUT4 #(
		.INIT('h8caf)
	) name369 (
		\in0[44] ,
		\in0[45] ,
		\in1[44] ,
		\in1[45] ,
		_w883_
	);
	LUT2 #(
		.INIT('h2)
	) name370 (
		\in0[43] ,
		\in1[43] ,
		_w884_
	);
	LUT2 #(
		.INIT('h8)
	) name371 (
		_w883_,
		_w884_,
		_w885_
	);
	LUT4 #(
		.INIT('h8caf)
	) name372 (
		\in0[42] ,
		\in0[43] ,
		\in1[42] ,
		\in1[43] ,
		_w886_
	);
	LUT4 #(
		.INIT('h080a)
	) name373 (
		\in0[40] ,
		\in0[41] ,
		\in1[40] ,
		\in1[41] ,
		_w887_
	);
	LUT4 #(
		.INIT('hf531)
	) name374 (
		\in0[41] ,
		\in0[42] ,
		\in1[41] ,
		\in1[42] ,
		_w888_
	);
	LUT4 #(
		.INIT('h8088)
	) name375 (
		_w883_,
		_w886_,
		_w887_,
		_w888_,
		_w889_
	);
	LUT4 #(
		.INIT('h080a)
	) name376 (
		\in0[44] ,
		\in0[45] ,
		\in1[44] ,
		\in1[45] ,
		_w890_
	);
	LUT4 #(
		.INIT('hf531)
	) name377 (
		\in0[45] ,
		\in0[46] ,
		\in1[45] ,
		\in1[46] ,
		_w891_
	);
	LUT3 #(
		.INIT('h10)
	) name378 (
		_w881_,
		_w890_,
		_w891_,
		_w892_
	);
	LUT4 #(
		.INIT('h5455)
	) name379 (
		_w882_,
		_w885_,
		_w889_,
		_w892_,
		_w893_
	);
	LUT2 #(
		.INIT('h2)
	) name380 (
		\in0[39] ,
		\in1[39] ,
		_w894_
	);
	LUT4 #(
		.INIT('h7310)
	) name381 (
		\in0[38] ,
		\in0[39] ,
		\in1[38] ,
		\in1[39] ,
		_w895_
	);
	LUT2 #(
		.INIT('h2)
	) name382 (
		\in0[35] ,
		\in1[35] ,
		_w896_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		_w872_,
		_w896_,
		_w897_
	);
	LUT4 #(
		.INIT('h080a)
	) name384 (
		\in0[32] ,
		\in0[33] ,
		\in1[32] ,
		\in1[33] ,
		_w898_
	);
	LUT4 #(
		.INIT('hf531)
	) name385 (
		\in0[33] ,
		\in0[34] ,
		\in1[33] ,
		\in1[34] ,
		_w899_
	);
	LUT4 #(
		.INIT('h8088)
	) name386 (
		_w869_,
		_w872_,
		_w898_,
		_w899_,
		_w900_
	);
	LUT4 #(
		.INIT('h080a)
	) name387 (
		\in0[36] ,
		\in0[37] ,
		\in1[36] ,
		\in1[37] ,
		_w901_
	);
	LUT4 #(
		.INIT('hf531)
	) name388 (
		\in0[37] ,
		\in0[38] ,
		\in1[37] ,
		\in1[38] ,
		_w902_
	);
	LUT3 #(
		.INIT('h10)
	) name389 (
		_w894_,
		_w901_,
		_w902_,
		_w903_
	);
	LUT4 #(
		.INIT('h5455)
	) name390 (
		_w895_,
		_w897_,
		_w900_,
		_w903_,
		_w904_
	);
	LUT3 #(
		.INIT('h01)
	) name391 (
		_w879_,
		_w893_,
		_w904_,
		_w905_
	);
	LUT4 #(
		.INIT('h8caf)
	) name392 (
		\in0[40] ,
		\in0[41] ,
		\in1[40] ,
		\in1[41] ,
		_w906_
	);
	LUT4 #(
		.INIT('h8000)
	) name393 (
		_w880_,
		_w883_,
		_w886_,
		_w906_,
		_w907_
	);
	LUT2 #(
		.INIT('h2)
	) name394 (
		_w882_,
		_w907_,
		_w908_
	);
	LUT4 #(
		.INIT('h0010)
	) name395 (
		_w885_,
		_w889_,
		_w892_,
		_w907_,
		_w909_
	);
	LUT4 #(
		.INIT('h8caf)
	) name396 (
		\in0[58] ,
		\in0[59] ,
		\in1[58] ,
		\in1[59] ,
		_w910_
	);
	LUT4 #(
		.INIT('h8caf)
	) name397 (
		\in0[60] ,
		\in0[61] ,
		\in1[60] ,
		\in1[61] ,
		_w911_
	);
	LUT4 #(
		.INIT('h8caf)
	) name398 (
		\in0[62] ,
		\in0[63] ,
		\in1[62] ,
		\in1[63] ,
		_w912_
	);
	LUT4 #(
		.INIT('h8caf)
	) name399 (
		\in0[56] ,
		\in0[57] ,
		\in1[56] ,
		\in1[57] ,
		_w913_
	);
	LUT4 #(
		.INIT('h8000)
	) name400 (
		_w910_,
		_w911_,
		_w912_,
		_w913_,
		_w914_
	);
	LUT4 #(
		.INIT('h8caf)
	) name401 (
		\in0[52] ,
		\in0[53] ,
		\in1[52] ,
		\in1[53] ,
		_w915_
	);
	LUT4 #(
		.INIT('h8caf)
	) name402 (
		\in0[50] ,
		\in0[51] ,
		\in1[50] ,
		\in1[51] ,
		_w916_
	);
	LUT4 #(
		.INIT('h8caf)
	) name403 (
		\in0[54] ,
		\in0[55] ,
		\in1[54] ,
		\in1[55] ,
		_w917_
	);
	LUT4 #(
		.INIT('h8caf)
	) name404 (
		\in0[48] ,
		\in0[49] ,
		\in1[48] ,
		\in1[49] ,
		_w918_
	);
	LUT4 #(
		.INIT('h8000)
	) name405 (
		_w915_,
		_w916_,
		_w917_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w914_,
		_w919_,
		_w920_
	);
	LUT3 #(
		.INIT('h10)
	) name407 (
		_w908_,
		_w909_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h2)
	) name408 (
		\in0[51] ,
		\in1[51] ,
		_w922_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w915_,
		_w922_,
		_w923_
	);
	LUT4 #(
		.INIT('h080a)
	) name410 (
		\in0[48] ,
		\in0[49] ,
		\in1[48] ,
		\in1[49] ,
		_w924_
	);
	LUT4 #(
		.INIT('hf531)
	) name411 (
		\in0[49] ,
		\in0[50] ,
		\in1[49] ,
		\in1[50] ,
		_w925_
	);
	LUT4 #(
		.INIT('h8088)
	) name412 (
		_w915_,
		_w916_,
		_w924_,
		_w925_,
		_w926_
	);
	LUT4 #(
		.INIT('h080a)
	) name413 (
		\in0[52] ,
		\in0[53] ,
		\in1[52] ,
		\in1[53] ,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name414 (
		\in0[55] ,
		\in1[55] ,
		_w928_
	);
	LUT4 #(
		.INIT('hf531)
	) name415 (
		\in0[53] ,
		\in0[54] ,
		\in1[53] ,
		\in1[54] ,
		_w929_
	);
	LUT3 #(
		.INIT('h10)
	) name416 (
		_w927_,
		_w928_,
		_w929_,
		_w930_
	);
	LUT3 #(
		.INIT('h10)
	) name417 (
		_w923_,
		_w926_,
		_w930_,
		_w931_
	);
	LUT4 #(
		.INIT('h7310)
	) name418 (
		\in0[54] ,
		\in0[55] ,
		\in1[54] ,
		\in1[55] ,
		_w932_
	);
	LUT2 #(
		.INIT('h2)
	) name419 (
		_w914_,
		_w932_,
		_w933_
	);
	LUT2 #(
		.INIT('h2)
	) name420 (
		\in0[63] ,
		\in1[63] ,
		_w934_
	);
	LUT4 #(
		.INIT('h7310)
	) name421 (
		\in0[62] ,
		\in0[63] ,
		\in1[62] ,
		\in1[63] ,
		_w935_
	);
	LUT2 #(
		.INIT('h2)
	) name422 (
		\in0[59] ,
		\in1[59] ,
		_w936_
	);
	LUT2 #(
		.INIT('h8)
	) name423 (
		_w911_,
		_w936_,
		_w937_
	);
	LUT4 #(
		.INIT('h080a)
	) name424 (
		\in0[56] ,
		\in0[57] ,
		\in1[56] ,
		\in1[57] ,
		_w938_
	);
	LUT4 #(
		.INIT('hf531)
	) name425 (
		\in0[57] ,
		\in0[58] ,
		\in1[57] ,
		\in1[58] ,
		_w939_
	);
	LUT4 #(
		.INIT('h8088)
	) name426 (
		_w910_,
		_w911_,
		_w938_,
		_w939_,
		_w940_
	);
	LUT4 #(
		.INIT('h080a)
	) name427 (
		\in0[60] ,
		\in0[61] ,
		\in1[60] ,
		\in1[61] ,
		_w941_
	);
	LUT4 #(
		.INIT('hf531)
	) name428 (
		\in0[61] ,
		\in0[62] ,
		\in1[61] ,
		\in1[62] ,
		_w942_
	);
	LUT3 #(
		.INIT('h10)
	) name429 (
		_w934_,
		_w941_,
		_w942_,
		_w943_
	);
	LUT4 #(
		.INIT('h5455)
	) name430 (
		_w935_,
		_w937_,
		_w940_,
		_w943_,
		_w944_
	);
	LUT3 #(
		.INIT('h0b)
	) name431 (
		_w931_,
		_w933_,
		_w944_,
		_w945_
	);
	LUT4 #(
		.INIT('h4f00)
	) name432 (
		_w876_,
		_w905_,
		_w921_,
		_w945_,
		_w946_
	);
	LUT4 #(
		.INIT('h8caf)
	) name433 (
		\in0[64] ,
		\in0[65] ,
		\in1[64] ,
		\in1[65] ,
		_w947_
	);
	LUT4 #(
		.INIT('h8000)
	) name434 (
		_w807_,
		_w811_,
		_w812_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h2)
	) name435 (
		\in0[71] ,
		\in1[71] ,
		_w949_
	);
	LUT4 #(
		.INIT('h080a)
	) name436 (
		\in0[68] ,
		\in0[69] ,
		\in1[68] ,
		\in1[69] ,
		_w950_
	);
	LUT4 #(
		.INIT('hf531)
	) name437 (
		\in0[69] ,
		\in0[70] ,
		\in1[69] ,
		\in1[70] ,
		_w951_
	);
	LUT4 #(
		.INIT('h1311)
	) name438 (
		_w811_,
		_w949_,
		_w950_,
		_w951_,
		_w952_
	);
	LUT2 #(
		.INIT('h8)
	) name439 (
		_w804_,
		_w952_,
		_w953_
	);
	LUT4 #(
		.INIT('h4500)
	) name440 (
		_w814_,
		_w946_,
		_w948_,
		_w953_,
		_w954_
	);
	LUT4 #(
		.INIT('h8caf)
	) name441 (
		\in0[76] ,
		\in0[77] ,
		\in1[76] ,
		\in1[77] ,
		_w955_
	);
	LUT3 #(
		.INIT('h80)
	) name442 (
		_w792_,
		_w796_,
		_w955_,
		_w956_
	);
	LUT4 #(
		.INIT('h5455)
	) name443 (
		_w797_,
		_w805_,
		_w954_,
		_w956_,
		_w957_
	);
	LUT4 #(
		.INIT('h8caf)
	) name444 (
		\in0[86] ,
		\in0[87] ,
		\in1[86] ,
		\in1[87] ,
		_w958_
	);
	LUT4 #(
		.INIT('h8caf)
	) name445 (
		\in0[84] ,
		\in0[85] ,
		\in1[84] ,
		\in1[85] ,
		_w959_
	);
	LUT2 #(
		.INIT('h8)
	) name446 (
		_w958_,
		_w959_,
		_w960_
	);
	LUT4 #(
		.INIT('h8caf)
	) name447 (
		\in0[82] ,
		\in0[83] ,
		\in1[82] ,
		\in1[83] ,
		_w961_
	);
	LUT3 #(
		.INIT('h80)
	) name448 (
		_w958_,
		_w959_,
		_w961_,
		_w962_
	);
	LUT2 #(
		.INIT('h2)
	) name449 (
		\in0[83] ,
		\in1[83] ,
		_w963_
	);
	LUT4 #(
		.INIT('h080a)
	) name450 (
		\in0[80] ,
		\in0[81] ,
		\in1[80] ,
		\in1[81] ,
		_w964_
	);
	LUT4 #(
		.INIT('hf531)
	) name451 (
		\in0[81] ,
		\in0[82] ,
		\in1[81] ,
		\in1[82] ,
		_w965_
	);
	LUT4 #(
		.INIT('h1311)
	) name452 (
		_w961_,
		_w963_,
		_w964_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h2)
	) name453 (
		\in0[91] ,
		\in1[91] ,
		_w967_
	);
	LUT4 #(
		.INIT('h8caf)
	) name454 (
		\in0[90] ,
		\in0[91] ,
		\in1[90] ,
		\in1[91] ,
		_w968_
	);
	LUT4 #(
		.INIT('h080a)
	) name455 (
		\in0[88] ,
		\in0[89] ,
		\in1[88] ,
		\in1[89] ,
		_w969_
	);
	LUT4 #(
		.INIT('hf531)
	) name456 (
		\in0[89] ,
		\in0[90] ,
		\in1[89] ,
		\in1[90] ,
		_w970_
	);
	LUT3 #(
		.INIT('h8a)
	) name457 (
		_w968_,
		_w969_,
		_w970_,
		_w971_
	);
	LUT4 #(
		.INIT('h1511)
	) name458 (
		_w967_,
		_w968_,
		_w969_,
		_w970_,
		_w972_
	);
	LUT2 #(
		.INIT('h2)
	) name459 (
		\in0[87] ,
		\in1[87] ,
		_w973_
	);
	LUT4 #(
		.INIT('h080a)
	) name460 (
		\in0[84] ,
		\in0[85] ,
		\in1[84] ,
		\in1[85] ,
		_w974_
	);
	LUT4 #(
		.INIT('hf531)
	) name461 (
		\in0[85] ,
		\in0[86] ,
		\in1[85] ,
		\in1[86] ,
		_w975_
	);
	LUT4 #(
		.INIT('h1311)
	) name462 (
		_w958_,
		_w973_,
		_w974_,
		_w975_,
		_w976_
	);
	LUT4 #(
		.INIT('hd000)
	) name463 (
		_w960_,
		_w966_,
		_w972_,
		_w976_,
		_w977_
	);
	LUT4 #(
		.INIT('h8caf)
	) name464 (
		\in0[88] ,
		\in0[89] ,
		\in1[88] ,
		\in1[89] ,
		_w978_
	);
	LUT3 #(
		.INIT('h15)
	) name465 (
		_w967_,
		_w968_,
		_w978_,
		_w979_
	);
	LUT4 #(
		.INIT('h8caf)
	) name466 (
		\in0[98] ,
		\in0[99] ,
		\in1[98] ,
		\in1[99] ,
		_w980_
	);
	LUT4 #(
		.INIT('h8caf)
	) name467 (
		\in0[96] ,
		\in0[97] ,
		\in1[96] ,
		\in1[97] ,
		_w981_
	);
	LUT2 #(
		.INIT('h8)
	) name468 (
		_w980_,
		_w981_,
		_w982_
	);
	LUT4 #(
		.INIT('h8caf)
	) name469 (
		\in0[94] ,
		\in0[95] ,
		\in1[94] ,
		\in1[95] ,
		_w983_
	);
	LUT4 #(
		.INIT('h8caf)
	) name470 (
		\in0[92] ,
		\in0[93] ,
		\in1[92] ,
		\in1[93] ,
		_w984_
	);
	LUT4 #(
		.INIT('h8000)
	) name471 (
		_w980_,
		_w981_,
		_w983_,
		_w984_,
		_w985_
	);
	LUT3 #(
		.INIT('hb0)
	) name472 (
		_w971_,
		_w979_,
		_w985_,
		_w986_
	);
	LUT4 #(
		.INIT('h4f00)
	) name473 (
		_w957_,
		_w962_,
		_w977_,
		_w986_,
		_w987_
	);
	LUT2 #(
		.INIT('h2)
	) name474 (
		\in0[95] ,
		\in1[95] ,
		_w988_
	);
	LUT4 #(
		.INIT('h080a)
	) name475 (
		\in0[92] ,
		\in0[93] ,
		\in1[92] ,
		\in1[93] ,
		_w989_
	);
	LUT4 #(
		.INIT('hf531)
	) name476 (
		\in0[93] ,
		\in0[94] ,
		\in1[93] ,
		\in1[94] ,
		_w990_
	);
	LUT4 #(
		.INIT('h1311)
	) name477 (
		_w983_,
		_w988_,
		_w989_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		\in0[103] ,
		\in1[103] ,
		_w992_
	);
	LUT4 #(
		.INIT('h8caf)
	) name479 (
		\in0[102] ,
		\in0[103] ,
		\in1[102] ,
		\in1[103] ,
		_w993_
	);
	LUT4 #(
		.INIT('h080a)
	) name480 (
		\in0[100] ,
		\in0[101] ,
		\in1[100] ,
		\in1[101] ,
		_w994_
	);
	LUT4 #(
		.INIT('hf531)
	) name481 (
		\in0[101] ,
		\in0[102] ,
		\in1[101] ,
		\in1[102] ,
		_w995_
	);
	LUT3 #(
		.INIT('h8a)
	) name482 (
		_w993_,
		_w994_,
		_w995_,
		_w996_
	);
	LUT4 #(
		.INIT('h1511)
	) name483 (
		_w992_,
		_w993_,
		_w994_,
		_w995_,
		_w997_
	);
	LUT2 #(
		.INIT('h2)
	) name484 (
		\in0[99] ,
		\in1[99] ,
		_w998_
	);
	LUT4 #(
		.INIT('h080a)
	) name485 (
		\in0[96] ,
		\in0[97] ,
		\in1[96] ,
		\in1[97] ,
		_w999_
	);
	LUT4 #(
		.INIT('hf531)
	) name486 (
		\in0[97] ,
		\in0[98] ,
		\in1[97] ,
		\in1[98] ,
		_w1000_
	);
	LUT4 #(
		.INIT('h1311)
	) name487 (
		_w980_,
		_w998_,
		_w999_,
		_w1000_,
		_w1001_
	);
	LUT4 #(
		.INIT('hd000)
	) name488 (
		_w982_,
		_w991_,
		_w997_,
		_w1001_,
		_w1002_
	);
	LUT4 #(
		.INIT('h8caf)
	) name489 (
		\in0[100] ,
		\in0[101] ,
		\in1[100] ,
		\in1[101] ,
		_w1003_
	);
	LUT3 #(
		.INIT('h15)
	) name490 (
		_w992_,
		_w993_,
		_w1003_,
		_w1004_
	);
	LUT4 #(
		.INIT('h8caf)
	) name491 (
		\in0[110] ,
		\in0[111] ,
		\in1[110] ,
		\in1[111] ,
		_w1005_
	);
	LUT4 #(
		.INIT('h8caf)
	) name492 (
		\in0[108] ,
		\in0[109] ,
		\in1[108] ,
		\in1[109] ,
		_w1006_
	);
	LUT4 #(
		.INIT('h8caf)
	) name493 (
		\in0[106] ,
		\in0[107] ,
		\in1[106] ,
		\in1[107] ,
		_w1007_
	);
	LUT4 #(
		.INIT('h8caf)
	) name494 (
		\in0[104] ,
		\in0[105] ,
		\in1[104] ,
		\in1[105] ,
		_w1008_
	);
	LUT4 #(
		.INIT('h8000)
	) name495 (
		_w1005_,
		_w1006_,
		_w1007_,
		_w1008_,
		_w1009_
	);
	LUT3 #(
		.INIT('hb0)
	) name496 (
		_w996_,
		_w1004_,
		_w1009_,
		_w1010_
	);
	LUT2 #(
		.INIT('h2)
	) name497 (
		\in0[107] ,
		\in1[107] ,
		_w1011_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		_w1006_,
		_w1011_,
		_w1012_
	);
	LUT4 #(
		.INIT('h080a)
	) name499 (
		\in0[104] ,
		\in0[105] ,
		\in1[104] ,
		\in1[105] ,
		_w1013_
	);
	LUT4 #(
		.INIT('hf531)
	) name500 (
		\in0[105] ,
		\in0[106] ,
		\in1[105] ,
		\in1[106] ,
		_w1014_
	);
	LUT4 #(
		.INIT('h8088)
	) name501 (
		_w1006_,
		_w1007_,
		_w1013_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		\in0[111] ,
		\in1[111] ,
		_w1016_
	);
	LUT4 #(
		.INIT('h080a)
	) name503 (
		\in0[108] ,
		\in0[109] ,
		\in1[108] ,
		\in1[109] ,
		_w1017_
	);
	LUT4 #(
		.INIT('hf531)
	) name504 (
		\in0[109] ,
		\in0[110] ,
		\in1[109] ,
		\in1[110] ,
		_w1018_
	);
	LUT4 #(
		.INIT('h1311)
	) name505 (
		_w1005_,
		_w1016_,
		_w1017_,
		_w1018_,
		_w1019_
	);
	LUT4 #(
		.INIT('h5700)
	) name506 (
		_w1005_,
		_w1012_,
		_w1015_,
		_w1019_,
		_w1020_
	);
	LUT4 #(
		.INIT('h4f00)
	) name507 (
		_w987_,
		_w1002_,
		_w1010_,
		_w1020_,
		_w1021_
	);
	LUT4 #(
		.INIT('h8caf)
	) name508 (
		\in0[112] ,
		\in0[113] ,
		\in1[112] ,
		\in1[113] ,
		_w1022_
	);
	LUT3 #(
		.INIT('h80)
	) name509 (
		_w785_,
		_w789_,
		_w1022_,
		_w1023_
	);
	LUT4 #(
		.INIT('h8caf)
	) name510 (
		\in0[122] ,
		\in0[123] ,
		\in1[122] ,
		\in1[123] ,
		_w1024_
	);
	LUT4 #(
		.INIT('h8caf)
	) name511 (
		\in0[120] ,
		\in0[121] ,
		\in1[120] ,
		\in1[121] ,
		_w1025_
	);
	LUT2 #(
		.INIT('h8)
	) name512 (
		_w1024_,
		_w1025_,
		_w1026_
	);
	LUT4 #(
		.INIT('h8caf)
	) name513 (
		\in0[118] ,
		\in0[119] ,
		\in1[118] ,
		\in1[119] ,
		_w1027_
	);
	LUT3 #(
		.INIT('h80)
	) name514 (
		_w1024_,
		_w1025_,
		_w1027_,
		_w1028_
	);
	LUT4 #(
		.INIT('hba00)
	) name515 (
		_w790_,
		_w1021_,
		_w1023_,
		_w1028_,
		_w1029_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\in0[119] ,
		\in1[119] ,
		_w1030_
	);
	LUT4 #(
		.INIT('h080a)
	) name517 (
		\in0[116] ,
		\in0[117] ,
		\in1[116] ,
		\in1[117] ,
		_w1031_
	);
	LUT4 #(
		.INIT('hf531)
	) name518 (
		\in0[117] ,
		\in0[118] ,
		\in1[117] ,
		\in1[118] ,
		_w1032_
	);
	LUT4 #(
		.INIT('h1311)
	) name519 (
		_w1027_,
		_w1030_,
		_w1031_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h2)
	) name520 (
		\in0[127] ,
		\in1[127] ,
		_w1034_
	);
	LUT4 #(
		.INIT('h8caf)
	) name521 (
		\in0[125] ,
		\in0[126] ,
		\in1[125] ,
		\in1[126] ,
		_w1035_
	);
	LUT4 #(
		.INIT('hf531)
	) name522 (
		\in0[124] ,
		\in0[125] ,
		\in1[124] ,
		\in1[125] ,
		_w1036_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name523 (
		\in0[126] ,
		\in0[127] ,
		\in1[126] ,
		\in1[127] ,
		_w1037_
	);
	LUT4 #(
		.INIT('h0455)
	) name524 (
		_w1034_,
		_w1035_,
		_w1036_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		\in0[123] ,
		\in1[123] ,
		_w1039_
	);
	LUT4 #(
		.INIT('h080a)
	) name526 (
		\in0[120] ,
		\in0[121] ,
		\in1[120] ,
		\in1[121] ,
		_w1040_
	);
	LUT4 #(
		.INIT('hf531)
	) name527 (
		\in0[121] ,
		\in0[122] ,
		\in1[121] ,
		\in1[122] ,
		_w1041_
	);
	LUT4 #(
		.INIT('h1311)
	) name528 (
		_w1024_,
		_w1039_,
		_w1040_,
		_w1041_,
		_w1042_
	);
	LUT4 #(
		.INIT('h0d00)
	) name529 (
		_w1026_,
		_w1033_,
		_w1038_,
		_w1042_,
		_w1043_
	);
	LUT4 #(
		.INIT('haf23)
	) name530 (
		\in0[124] ,
		\in0[127] ,
		\in1[124] ,
		\in1[127] ,
		_w1044_
	);
	LUT2 #(
		.INIT('h8)
	) name531 (
		_w1035_,
		_w1044_,
		_w1045_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w1038_,
		_w1045_,
		_w1046_
	);
	LUT3 #(
		.INIT('ha8)
	) name533 (
		\in0[126] ,
		_w1038_,
		_w1045_,
		_w1047_
	);
	LUT3 #(
		.INIT('hb0)
	) name534 (
		_w1029_,
		_w1043_,
		_w1047_,
		_w1048_
	);
	LUT3 #(
		.INIT('h0b)
	) name535 (
		_w1029_,
		_w1043_,
		_w1046_,
		_w1049_
	);
	LUT4 #(
		.INIT('haa20)
	) name536 (
		\in1[126] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1050_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		_w1048_,
		_w1050_,
		_w1051_
	);
	LUT3 #(
		.INIT('ha8)
	) name538 (
		\in2[126] ,
		_w521_,
		_w778_,
		_w1052_
	);
	LUT4 #(
		.INIT('h1500)
	) name539 (
		_w526_,
		_w771_,
		_w776_,
		_w1052_,
		_w1053_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name540 (
		\in3[126] ,
		_w782_,
		_w1051_,
		_w1053_,
		_w1054_
	);
	LUT3 #(
		.INIT('ha8)
	) name541 (
		\in0[125] ,
		_w1038_,
		_w1045_,
		_w1055_
	);
	LUT3 #(
		.INIT('hb0)
	) name542 (
		_w1029_,
		_w1043_,
		_w1055_,
		_w1056_
	);
	LUT4 #(
		.INIT('haa20)
	) name543 (
		\in1[125] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w1056_,
		_w1057_,
		_w1058_
	);
	LUT3 #(
		.INIT('ha8)
	) name545 (
		\in2[125] ,
		_w521_,
		_w778_,
		_w1059_
	);
	LUT4 #(
		.INIT('h1500)
	) name546 (
		_w526_,
		_w771_,
		_w776_,
		_w1059_,
		_w1060_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name547 (
		\in3[125] ,
		_w782_,
		_w1058_,
		_w1060_,
		_w1061_
	);
	LUT4 #(
		.INIT('h0888)
	) name548 (
		\in0[127] ,
		\in1[127] ,
		\in2[127] ,
		\in3[127] ,
		_w1062_
	);
	LUT3 #(
		.INIT('ha8)
	) name549 (
		\in0[124] ,
		_w1038_,
		_w1045_,
		_w1063_
	);
	LUT3 #(
		.INIT('hb0)
	) name550 (
		_w1029_,
		_w1043_,
		_w1063_,
		_w1064_
	);
	LUT4 #(
		.INIT('haa20)
	) name551 (
		\in1[124] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w1064_,
		_w1065_,
		_w1066_
	);
	LUT3 #(
		.INIT('ha8)
	) name553 (
		\in2[124] ,
		_w521_,
		_w778_,
		_w1067_
	);
	LUT4 #(
		.INIT('h1500)
	) name554 (
		_w526_,
		_w771_,
		_w776_,
		_w1067_,
		_w1068_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name555 (
		\in3[124] ,
		_w782_,
		_w1066_,
		_w1068_,
		_w1069_
	);
	LUT4 #(
		.INIT('h0800)
	) name556 (
		_w1054_,
		_w1061_,
		_w1062_,
		_w1069_,
		_w1070_
	);
	LUT4 #(
		.INIT('h000d)
	) name557 (
		\in3[124] ,
		_w782_,
		_w1066_,
		_w1068_,
		_w1071_
	);
	LUT4 #(
		.INIT('h000d)
	) name558 (
		\in3[125] ,
		_w782_,
		_w1058_,
		_w1060_,
		_w1072_
	);
	LUT4 #(
		.INIT('h8880)
	) name559 (
		_w1054_,
		_w1061_,
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT4 #(
		.INIT('h7000)
	) name560 (
		\in0[127] ,
		\in1[127] ,
		\in2[127] ,
		\in3[127] ,
		_w1074_
	);
	LUT4 #(
		.INIT('h000d)
	) name561 (
		\in3[126] ,
		_w782_,
		_w1051_,
		_w1053_,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name562 (
		_w1074_,
		_w1075_,
		_w1076_
	);
	LUT3 #(
		.INIT('h45)
	) name563 (
		_w1062_,
		_w1073_,
		_w1076_,
		_w1077_
	);
	LUT4 #(
		.INIT('h2322)
	) name564 (
		_w1062_,
		_w1070_,
		_w1073_,
		_w1076_,
		_w1078_
	);
	LUT3 #(
		.INIT('ha8)
	) name565 (
		\in0[123] ,
		_w1038_,
		_w1045_,
		_w1079_
	);
	LUT3 #(
		.INIT('hb0)
	) name566 (
		_w1029_,
		_w1043_,
		_w1079_,
		_w1080_
	);
	LUT4 #(
		.INIT('haa20)
	) name567 (
		\in1[123] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w1080_,
		_w1081_,
		_w1082_
	);
	LUT3 #(
		.INIT('ha8)
	) name569 (
		\in2[123] ,
		_w521_,
		_w778_,
		_w1083_
	);
	LUT4 #(
		.INIT('h1500)
	) name570 (
		_w526_,
		_w771_,
		_w776_,
		_w1083_,
		_w1084_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name571 (
		\in3[123] ,
		_w782_,
		_w1082_,
		_w1084_,
		_w1085_
	);
	LUT3 #(
		.INIT('ha8)
	) name572 (
		\in0[122] ,
		_w1038_,
		_w1045_,
		_w1086_
	);
	LUT3 #(
		.INIT('hb0)
	) name573 (
		_w1029_,
		_w1043_,
		_w1086_,
		_w1087_
	);
	LUT4 #(
		.INIT('haa20)
	) name574 (
		\in1[122] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1088_
	);
	LUT2 #(
		.INIT('h1)
	) name575 (
		_w1087_,
		_w1088_,
		_w1089_
	);
	LUT3 #(
		.INIT('h02)
	) name576 (
		\in3[122] ,
		_w1087_,
		_w1088_,
		_w1090_
	);
	LUT3 #(
		.INIT('h02)
	) name577 (
		\in2[122] ,
		_w1087_,
		_w1088_,
		_w1091_
	);
	LUT3 #(
		.INIT('h1b)
	) name578 (
		_w782_,
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h8)
	) name579 (
		_w1085_,
		_w1092_,
		_w1093_
	);
	LUT3 #(
		.INIT('ha8)
	) name580 (
		\in0[120] ,
		_w1038_,
		_w1045_,
		_w1094_
	);
	LUT3 #(
		.INIT('hb0)
	) name581 (
		_w1029_,
		_w1043_,
		_w1094_,
		_w1095_
	);
	LUT4 #(
		.INIT('haa20)
	) name582 (
		\in1[120] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1096_
	);
	LUT2 #(
		.INIT('h1)
	) name583 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT3 #(
		.INIT('h02)
	) name584 (
		\in3[120] ,
		_w1095_,
		_w1096_,
		_w1098_
	);
	LUT3 #(
		.INIT('h02)
	) name585 (
		\in2[120] ,
		_w1095_,
		_w1096_,
		_w1099_
	);
	LUT3 #(
		.INIT('h1b)
	) name586 (
		_w782_,
		_w1098_,
		_w1099_,
		_w1100_
	);
	LUT3 #(
		.INIT('ha8)
	) name587 (
		\in0[121] ,
		_w1038_,
		_w1045_,
		_w1101_
	);
	LUT3 #(
		.INIT('hb0)
	) name588 (
		_w1029_,
		_w1043_,
		_w1101_,
		_w1102_
	);
	LUT4 #(
		.INIT('haa20)
	) name589 (
		\in1[121] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1103_
	);
	LUT2 #(
		.INIT('h1)
	) name590 (
		_w1102_,
		_w1103_,
		_w1104_
	);
	LUT3 #(
		.INIT('ha8)
	) name591 (
		\in2[121] ,
		_w521_,
		_w778_,
		_w1105_
	);
	LUT4 #(
		.INIT('h1500)
	) name592 (
		_w526_,
		_w771_,
		_w776_,
		_w1105_,
		_w1106_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name593 (
		\in3[121] ,
		_w782_,
		_w1104_,
		_w1106_,
		_w1107_
	);
	LUT4 #(
		.INIT('h8000)
	) name594 (
		_w1085_,
		_w1092_,
		_w1100_,
		_w1107_,
		_w1108_
	);
	LUT4 #(
		.INIT('h000d)
	) name595 (
		\in3[123] ,
		_w782_,
		_w1082_,
		_w1084_,
		_w1109_
	);
	LUT3 #(
		.INIT('ha8)
	) name596 (
		\in2[120] ,
		_w521_,
		_w778_,
		_w1110_
	);
	LUT4 #(
		.INIT('h1500)
	) name597 (
		_w526_,
		_w771_,
		_w776_,
		_w1110_,
		_w1111_
	);
	LUT4 #(
		.INIT('h000d)
	) name598 (
		\in3[120] ,
		_w782_,
		_w1097_,
		_w1111_,
		_w1112_
	);
	LUT4 #(
		.INIT('h000d)
	) name599 (
		\in3[121] ,
		_w782_,
		_w1104_,
		_w1106_,
		_w1113_
	);
	LUT3 #(
		.INIT('ha8)
	) name600 (
		\in2[122] ,
		_w521_,
		_w778_,
		_w1114_
	);
	LUT4 #(
		.INIT('h1500)
	) name601 (
		_w526_,
		_w771_,
		_w776_,
		_w1114_,
		_w1115_
	);
	LUT4 #(
		.INIT('h000d)
	) name602 (
		\in3[122] ,
		_w782_,
		_w1089_,
		_w1115_,
		_w1116_
	);
	LUT4 #(
		.INIT('h0007)
	) name603 (
		_w1107_,
		_w1112_,
		_w1113_,
		_w1116_,
		_w1117_
	);
	LUT3 #(
		.INIT('h31)
	) name604 (
		_w1093_,
		_w1109_,
		_w1117_,
		_w1118_
	);
	LUT3 #(
		.INIT('h10)
	) name605 (
		_w1077_,
		_w1108_,
		_w1118_,
		_w1119_
	);
	LUT3 #(
		.INIT('ha8)
	) name606 (
		\in0[111] ,
		_w1038_,
		_w1045_,
		_w1120_
	);
	LUT3 #(
		.INIT('hb0)
	) name607 (
		_w1029_,
		_w1043_,
		_w1120_,
		_w1121_
	);
	LUT4 #(
		.INIT('haa20)
	) name608 (
		\in1[111] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1122_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		_w1121_,
		_w1122_,
		_w1123_
	);
	LUT3 #(
		.INIT('ha8)
	) name610 (
		\in2[111] ,
		_w521_,
		_w778_,
		_w1124_
	);
	LUT4 #(
		.INIT('h1500)
	) name611 (
		_w526_,
		_w771_,
		_w776_,
		_w1124_,
		_w1125_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name612 (
		\in3[111] ,
		_w782_,
		_w1123_,
		_w1125_,
		_w1126_
	);
	LUT3 #(
		.INIT('ha8)
	) name613 (
		\in0[110] ,
		_w1038_,
		_w1045_,
		_w1127_
	);
	LUT3 #(
		.INIT('hb0)
	) name614 (
		_w1029_,
		_w1043_,
		_w1127_,
		_w1128_
	);
	LUT4 #(
		.INIT('haa20)
	) name615 (
		\in1[110] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1129_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		_w1128_,
		_w1129_,
		_w1130_
	);
	LUT3 #(
		.INIT('h02)
	) name617 (
		\in3[110] ,
		_w1128_,
		_w1129_,
		_w1131_
	);
	LUT3 #(
		.INIT('h02)
	) name618 (
		\in2[110] ,
		_w1128_,
		_w1129_,
		_w1132_
	);
	LUT3 #(
		.INIT('h1b)
	) name619 (
		_w782_,
		_w1131_,
		_w1132_,
		_w1133_
	);
	LUT2 #(
		.INIT('h8)
	) name620 (
		_w1126_,
		_w1133_,
		_w1134_
	);
	LUT3 #(
		.INIT('ha8)
	) name621 (
		\in0[108] ,
		_w1038_,
		_w1045_,
		_w1135_
	);
	LUT3 #(
		.INIT('hb0)
	) name622 (
		_w1029_,
		_w1043_,
		_w1135_,
		_w1136_
	);
	LUT4 #(
		.INIT('haa20)
	) name623 (
		\in1[108] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1137_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w1136_,
		_w1137_,
		_w1138_
	);
	LUT3 #(
		.INIT('h02)
	) name625 (
		\in3[108] ,
		_w1136_,
		_w1137_,
		_w1139_
	);
	LUT3 #(
		.INIT('h02)
	) name626 (
		\in2[108] ,
		_w1136_,
		_w1137_,
		_w1140_
	);
	LUT3 #(
		.INIT('h1b)
	) name627 (
		_w782_,
		_w1139_,
		_w1140_,
		_w1141_
	);
	LUT3 #(
		.INIT('ha8)
	) name628 (
		\in0[109] ,
		_w1038_,
		_w1045_,
		_w1142_
	);
	LUT3 #(
		.INIT('hb0)
	) name629 (
		_w1029_,
		_w1043_,
		_w1142_,
		_w1143_
	);
	LUT4 #(
		.INIT('haa20)
	) name630 (
		\in1[109] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name631 (
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT3 #(
		.INIT('ha8)
	) name632 (
		\in2[109] ,
		_w521_,
		_w778_,
		_w1146_
	);
	LUT4 #(
		.INIT('h1500)
	) name633 (
		_w526_,
		_w771_,
		_w776_,
		_w1146_,
		_w1147_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name634 (
		\in3[109] ,
		_w782_,
		_w1145_,
		_w1147_,
		_w1148_
	);
	LUT4 #(
		.INIT('h8000)
	) name635 (
		_w1126_,
		_w1133_,
		_w1141_,
		_w1148_,
		_w1149_
	);
	LUT3 #(
		.INIT('ha8)
	) name636 (
		\in0[115] ,
		_w1038_,
		_w1045_,
		_w1150_
	);
	LUT3 #(
		.INIT('hb0)
	) name637 (
		_w1029_,
		_w1043_,
		_w1150_,
		_w1151_
	);
	LUT4 #(
		.INIT('haa20)
	) name638 (
		\in1[115] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w1151_,
		_w1152_,
		_w1153_
	);
	LUT3 #(
		.INIT('ha8)
	) name640 (
		\in2[115] ,
		_w521_,
		_w778_,
		_w1154_
	);
	LUT4 #(
		.INIT('h1500)
	) name641 (
		_w526_,
		_w771_,
		_w776_,
		_w1154_,
		_w1155_
	);
	LUT4 #(
		.INIT('h000d)
	) name642 (
		\in3[115] ,
		_w782_,
		_w1153_,
		_w1155_,
		_w1156_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name643 (
		\in3[115] ,
		_w782_,
		_w1153_,
		_w1155_,
		_w1157_
	);
	LUT3 #(
		.INIT('ha8)
	) name644 (
		\in0[114] ,
		_w1038_,
		_w1045_,
		_w1158_
	);
	LUT3 #(
		.INIT('hb0)
	) name645 (
		_w1029_,
		_w1043_,
		_w1158_,
		_w1159_
	);
	LUT4 #(
		.INIT('haa20)
	) name646 (
		\in1[114] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w1159_,
		_w1160_,
		_w1161_
	);
	LUT3 #(
		.INIT('h02)
	) name648 (
		\in3[114] ,
		_w1159_,
		_w1160_,
		_w1162_
	);
	LUT3 #(
		.INIT('h02)
	) name649 (
		\in2[114] ,
		_w1159_,
		_w1160_,
		_w1163_
	);
	LUT3 #(
		.INIT('h1b)
	) name650 (
		_w782_,
		_w1162_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h8)
	) name651 (
		_w1157_,
		_w1164_,
		_w1165_
	);
	LUT3 #(
		.INIT('ha8)
	) name652 (
		\in0[113] ,
		_w1038_,
		_w1045_,
		_w1166_
	);
	LUT3 #(
		.INIT('hb0)
	) name653 (
		_w1029_,
		_w1043_,
		_w1166_,
		_w1167_
	);
	LUT4 #(
		.INIT('haa20)
	) name654 (
		\in1[113] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1168_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		_w1167_,
		_w1168_,
		_w1169_
	);
	LUT3 #(
		.INIT('ha8)
	) name656 (
		\in2[113] ,
		_w521_,
		_w778_,
		_w1170_
	);
	LUT4 #(
		.INIT('h1500)
	) name657 (
		_w526_,
		_w771_,
		_w776_,
		_w1170_,
		_w1171_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name658 (
		\in3[113] ,
		_w782_,
		_w1169_,
		_w1171_,
		_w1172_
	);
	LUT3 #(
		.INIT('ha8)
	) name659 (
		\in2[112] ,
		_w521_,
		_w778_,
		_w1173_
	);
	LUT4 #(
		.INIT('h1500)
	) name660 (
		_w526_,
		_w771_,
		_w776_,
		_w1173_,
		_w1174_
	);
	LUT3 #(
		.INIT('ha8)
	) name661 (
		\in0[112] ,
		_w1038_,
		_w1045_,
		_w1175_
	);
	LUT3 #(
		.INIT('hb0)
	) name662 (
		_w1029_,
		_w1043_,
		_w1175_,
		_w1176_
	);
	LUT4 #(
		.INIT('haa20)
	) name663 (
		\in1[112] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1177_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w1176_,
		_w1177_,
		_w1178_
	);
	LUT4 #(
		.INIT('h000d)
	) name665 (
		\in3[112] ,
		_w782_,
		_w1174_,
		_w1178_,
		_w1179_
	);
	LUT4 #(
		.INIT('h000d)
	) name666 (
		\in3[113] ,
		_w782_,
		_w1169_,
		_w1171_,
		_w1180_
	);
	LUT3 #(
		.INIT('ha8)
	) name667 (
		\in2[114] ,
		_w521_,
		_w778_,
		_w1181_
	);
	LUT4 #(
		.INIT('h1500)
	) name668 (
		_w526_,
		_w771_,
		_w776_,
		_w1181_,
		_w1182_
	);
	LUT4 #(
		.INIT('h000d)
	) name669 (
		\in3[114] ,
		_w782_,
		_w1161_,
		_w1182_,
		_w1183_
	);
	LUT4 #(
		.INIT('h0007)
	) name670 (
		_w1172_,
		_w1179_,
		_w1180_,
		_w1183_,
		_w1184_
	);
	LUT3 #(
		.INIT('h51)
	) name671 (
		_w1156_,
		_w1165_,
		_w1184_,
		_w1185_
	);
	LUT4 #(
		.INIT('h000d)
	) name672 (
		\in3[111] ,
		_w782_,
		_w1123_,
		_w1125_,
		_w1186_
	);
	LUT3 #(
		.INIT('ha8)
	) name673 (
		\in2[108] ,
		_w521_,
		_w778_,
		_w1187_
	);
	LUT4 #(
		.INIT('h1500)
	) name674 (
		_w526_,
		_w771_,
		_w776_,
		_w1187_,
		_w1188_
	);
	LUT4 #(
		.INIT('h000d)
	) name675 (
		\in3[108] ,
		_w782_,
		_w1138_,
		_w1188_,
		_w1189_
	);
	LUT3 #(
		.INIT('ha8)
	) name676 (
		\in2[110] ,
		_w521_,
		_w778_,
		_w1190_
	);
	LUT4 #(
		.INIT('h1500)
	) name677 (
		_w526_,
		_w771_,
		_w776_,
		_w1190_,
		_w1191_
	);
	LUT4 #(
		.INIT('h000d)
	) name678 (
		\in3[110] ,
		_w782_,
		_w1130_,
		_w1191_,
		_w1192_
	);
	LUT4 #(
		.INIT('h000d)
	) name679 (
		\in3[109] ,
		_w782_,
		_w1145_,
		_w1147_,
		_w1193_
	);
	LUT4 #(
		.INIT('h0007)
	) name680 (
		_w1148_,
		_w1189_,
		_w1192_,
		_w1193_,
		_w1194_
	);
	LUT3 #(
		.INIT('h31)
	) name681 (
		_w1134_,
		_w1186_,
		_w1194_,
		_w1195_
	);
	LUT3 #(
		.INIT('h40)
	) name682 (
		_w1149_,
		_w1185_,
		_w1195_,
		_w1196_
	);
	LUT3 #(
		.INIT('ha8)
	) name683 (
		\in0[103] ,
		_w1038_,
		_w1045_,
		_w1197_
	);
	LUT3 #(
		.INIT('hb0)
	) name684 (
		_w1029_,
		_w1043_,
		_w1197_,
		_w1198_
	);
	LUT4 #(
		.INIT('haa20)
	) name685 (
		\in1[103] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1199_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		_w1198_,
		_w1199_,
		_w1200_
	);
	LUT3 #(
		.INIT('ha8)
	) name687 (
		\in2[103] ,
		_w521_,
		_w778_,
		_w1201_
	);
	LUT4 #(
		.INIT('h1500)
	) name688 (
		_w526_,
		_w771_,
		_w776_,
		_w1201_,
		_w1202_
	);
	LUT4 #(
		.INIT('h000d)
	) name689 (
		\in3[103] ,
		_w782_,
		_w1200_,
		_w1202_,
		_w1203_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name690 (
		\in3[103] ,
		_w782_,
		_w1200_,
		_w1202_,
		_w1204_
	);
	LUT3 #(
		.INIT('ha8)
	) name691 (
		\in0[102] ,
		_w1038_,
		_w1045_,
		_w1205_
	);
	LUT3 #(
		.INIT('hb0)
	) name692 (
		_w1029_,
		_w1043_,
		_w1205_,
		_w1206_
	);
	LUT4 #(
		.INIT('haa20)
	) name693 (
		\in1[102] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1207_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w1206_,
		_w1207_,
		_w1208_
	);
	LUT3 #(
		.INIT('h02)
	) name695 (
		\in3[102] ,
		_w1206_,
		_w1207_,
		_w1209_
	);
	LUT3 #(
		.INIT('h02)
	) name696 (
		\in2[102] ,
		_w1206_,
		_w1207_,
		_w1210_
	);
	LUT3 #(
		.INIT('h1b)
	) name697 (
		_w782_,
		_w1209_,
		_w1210_,
		_w1211_
	);
	LUT2 #(
		.INIT('h8)
	) name698 (
		_w1204_,
		_w1211_,
		_w1212_
	);
	LUT3 #(
		.INIT('ha8)
	) name699 (
		\in0[101] ,
		_w1038_,
		_w1045_,
		_w1213_
	);
	LUT3 #(
		.INIT('hb0)
	) name700 (
		_w1029_,
		_w1043_,
		_w1213_,
		_w1214_
	);
	LUT4 #(
		.INIT('haa20)
	) name701 (
		\in1[101] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1215_
	);
	LUT2 #(
		.INIT('h1)
	) name702 (
		_w1214_,
		_w1215_,
		_w1216_
	);
	LUT3 #(
		.INIT('ha8)
	) name703 (
		\in2[101] ,
		_w521_,
		_w778_,
		_w1217_
	);
	LUT4 #(
		.INIT('h1500)
	) name704 (
		_w526_,
		_w771_,
		_w776_,
		_w1217_,
		_w1218_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name705 (
		\in3[101] ,
		_w782_,
		_w1216_,
		_w1218_,
		_w1219_
	);
	LUT3 #(
		.INIT('ha8)
	) name706 (
		\in2[100] ,
		_w521_,
		_w778_,
		_w1220_
	);
	LUT4 #(
		.INIT('h1500)
	) name707 (
		_w526_,
		_w771_,
		_w776_,
		_w1220_,
		_w1221_
	);
	LUT3 #(
		.INIT('ha8)
	) name708 (
		\in0[100] ,
		_w1038_,
		_w1045_,
		_w1222_
	);
	LUT3 #(
		.INIT('hb0)
	) name709 (
		_w1029_,
		_w1043_,
		_w1222_,
		_w1223_
	);
	LUT4 #(
		.INIT('haa20)
	) name710 (
		\in1[100] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1224_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w1223_,
		_w1224_,
		_w1225_
	);
	LUT4 #(
		.INIT('h000d)
	) name712 (
		\in3[100] ,
		_w782_,
		_w1221_,
		_w1225_,
		_w1226_
	);
	LUT3 #(
		.INIT('ha8)
	) name713 (
		\in2[102] ,
		_w521_,
		_w778_,
		_w1227_
	);
	LUT4 #(
		.INIT('h1500)
	) name714 (
		_w526_,
		_w771_,
		_w776_,
		_w1227_,
		_w1228_
	);
	LUT4 #(
		.INIT('h000d)
	) name715 (
		\in3[102] ,
		_w782_,
		_w1208_,
		_w1228_,
		_w1229_
	);
	LUT4 #(
		.INIT('h000d)
	) name716 (
		\in3[101] ,
		_w782_,
		_w1216_,
		_w1218_,
		_w1230_
	);
	LUT4 #(
		.INIT('h0007)
	) name717 (
		_w1219_,
		_w1226_,
		_w1229_,
		_w1230_,
		_w1231_
	);
	LUT3 #(
		.INIT('ha8)
	) name718 (
		\in0[107] ,
		_w1038_,
		_w1045_,
		_w1232_
	);
	LUT3 #(
		.INIT('hb0)
	) name719 (
		_w1029_,
		_w1043_,
		_w1232_,
		_w1233_
	);
	LUT4 #(
		.INIT('haa20)
	) name720 (
		\in1[107] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1234_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		_w1233_,
		_w1234_,
		_w1235_
	);
	LUT3 #(
		.INIT('ha8)
	) name722 (
		\in2[107] ,
		_w521_,
		_w778_,
		_w1236_
	);
	LUT4 #(
		.INIT('h1500)
	) name723 (
		_w526_,
		_w771_,
		_w776_,
		_w1236_,
		_w1237_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name724 (
		\in3[107] ,
		_w782_,
		_w1235_,
		_w1237_,
		_w1238_
	);
	LUT3 #(
		.INIT('ha8)
	) name725 (
		\in0[106] ,
		_w1038_,
		_w1045_,
		_w1239_
	);
	LUT3 #(
		.INIT('hb0)
	) name726 (
		_w1029_,
		_w1043_,
		_w1239_,
		_w1240_
	);
	LUT4 #(
		.INIT('haa20)
	) name727 (
		\in1[106] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1241_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		_w1240_,
		_w1241_,
		_w1242_
	);
	LUT3 #(
		.INIT('h02)
	) name729 (
		\in3[106] ,
		_w1240_,
		_w1241_,
		_w1243_
	);
	LUT3 #(
		.INIT('h02)
	) name730 (
		\in2[106] ,
		_w1240_,
		_w1241_,
		_w1244_
	);
	LUT3 #(
		.INIT('h1b)
	) name731 (
		_w782_,
		_w1243_,
		_w1244_,
		_w1245_
	);
	LUT2 #(
		.INIT('h8)
	) name732 (
		_w1238_,
		_w1245_,
		_w1246_
	);
	LUT3 #(
		.INIT('ha8)
	) name733 (
		\in0[105] ,
		_w1038_,
		_w1045_,
		_w1247_
	);
	LUT3 #(
		.INIT('hb0)
	) name734 (
		_w1029_,
		_w1043_,
		_w1247_,
		_w1248_
	);
	LUT4 #(
		.INIT('haa20)
	) name735 (
		\in1[105] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w1248_,
		_w1249_,
		_w1250_
	);
	LUT3 #(
		.INIT('ha8)
	) name737 (
		\in2[105] ,
		_w521_,
		_w778_,
		_w1251_
	);
	LUT4 #(
		.INIT('h1500)
	) name738 (
		_w526_,
		_w771_,
		_w776_,
		_w1251_,
		_w1252_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name739 (
		\in3[105] ,
		_w782_,
		_w1250_,
		_w1252_,
		_w1253_
	);
	LUT3 #(
		.INIT('ha8)
	) name740 (
		\in0[104] ,
		_w1038_,
		_w1045_,
		_w1254_
	);
	LUT3 #(
		.INIT('hb0)
	) name741 (
		_w1029_,
		_w1043_,
		_w1254_,
		_w1255_
	);
	LUT4 #(
		.INIT('haa20)
	) name742 (
		\in1[104] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w1255_,
		_w1256_,
		_w1257_
	);
	LUT3 #(
		.INIT('h02)
	) name744 (
		\in3[104] ,
		_w1255_,
		_w1256_,
		_w1258_
	);
	LUT3 #(
		.INIT('h02)
	) name745 (
		\in2[104] ,
		_w1255_,
		_w1256_,
		_w1259_
	);
	LUT3 #(
		.INIT('h1b)
	) name746 (
		_w782_,
		_w1258_,
		_w1259_,
		_w1260_
	);
	LUT4 #(
		.INIT('h8000)
	) name747 (
		_w1238_,
		_w1245_,
		_w1253_,
		_w1260_,
		_w1261_
	);
	LUT4 #(
		.INIT('hae00)
	) name748 (
		_w1203_,
		_w1212_,
		_w1231_,
		_w1261_,
		_w1262_
	);
	LUT3 #(
		.INIT('ha8)
	) name749 (
		\in0[99] ,
		_w1038_,
		_w1045_,
		_w1263_
	);
	LUT3 #(
		.INIT('hb0)
	) name750 (
		_w1029_,
		_w1043_,
		_w1263_,
		_w1264_
	);
	LUT4 #(
		.INIT('haa20)
	) name751 (
		\in1[99] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w1264_,
		_w1265_,
		_w1266_
	);
	LUT3 #(
		.INIT('ha8)
	) name753 (
		\in2[99] ,
		_w521_,
		_w778_,
		_w1267_
	);
	LUT4 #(
		.INIT('h1500)
	) name754 (
		_w526_,
		_w771_,
		_w776_,
		_w1267_,
		_w1268_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name755 (
		\in3[99] ,
		_w782_,
		_w1266_,
		_w1268_,
		_w1269_
	);
	LUT3 #(
		.INIT('ha8)
	) name756 (
		\in0[98] ,
		_w1038_,
		_w1045_,
		_w1270_
	);
	LUT3 #(
		.INIT('hb0)
	) name757 (
		_w1029_,
		_w1043_,
		_w1270_,
		_w1271_
	);
	LUT4 #(
		.INIT('haa20)
	) name758 (
		\in1[98] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name759 (
		_w1271_,
		_w1272_,
		_w1273_
	);
	LUT3 #(
		.INIT('h02)
	) name760 (
		\in3[98] ,
		_w1271_,
		_w1272_,
		_w1274_
	);
	LUT3 #(
		.INIT('h02)
	) name761 (
		\in2[98] ,
		_w1271_,
		_w1272_,
		_w1275_
	);
	LUT3 #(
		.INIT('h1b)
	) name762 (
		_w782_,
		_w1274_,
		_w1275_,
		_w1276_
	);
	LUT2 #(
		.INIT('h8)
	) name763 (
		_w1269_,
		_w1276_,
		_w1277_
	);
	LUT3 #(
		.INIT('ha8)
	) name764 (
		\in0[96] ,
		_w1038_,
		_w1045_,
		_w1278_
	);
	LUT3 #(
		.INIT('hb0)
	) name765 (
		_w1029_,
		_w1043_,
		_w1278_,
		_w1279_
	);
	LUT4 #(
		.INIT('haa20)
	) name766 (
		\in1[96] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1280_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w1279_,
		_w1280_,
		_w1281_
	);
	LUT3 #(
		.INIT('h02)
	) name768 (
		\in3[96] ,
		_w1279_,
		_w1280_,
		_w1282_
	);
	LUT3 #(
		.INIT('h02)
	) name769 (
		\in2[96] ,
		_w1279_,
		_w1280_,
		_w1283_
	);
	LUT3 #(
		.INIT('h1b)
	) name770 (
		_w782_,
		_w1282_,
		_w1283_,
		_w1284_
	);
	LUT3 #(
		.INIT('ha8)
	) name771 (
		\in0[97] ,
		_w1038_,
		_w1045_,
		_w1285_
	);
	LUT3 #(
		.INIT('hb0)
	) name772 (
		_w1029_,
		_w1043_,
		_w1285_,
		_w1286_
	);
	LUT4 #(
		.INIT('haa20)
	) name773 (
		\in1[97] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1287_
	);
	LUT2 #(
		.INIT('h1)
	) name774 (
		_w1286_,
		_w1287_,
		_w1288_
	);
	LUT3 #(
		.INIT('ha8)
	) name775 (
		\in2[97] ,
		_w521_,
		_w778_,
		_w1289_
	);
	LUT4 #(
		.INIT('h1500)
	) name776 (
		_w526_,
		_w771_,
		_w776_,
		_w1289_,
		_w1290_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name777 (
		\in3[97] ,
		_w782_,
		_w1288_,
		_w1290_,
		_w1291_
	);
	LUT4 #(
		.INIT('h8000)
	) name778 (
		_w1269_,
		_w1276_,
		_w1284_,
		_w1291_,
		_w1292_
	);
	LUT4 #(
		.INIT('h000d)
	) name779 (
		\in3[99] ,
		_w782_,
		_w1266_,
		_w1268_,
		_w1293_
	);
	LUT3 #(
		.INIT('ha8)
	) name780 (
		\in2[96] ,
		_w521_,
		_w778_,
		_w1294_
	);
	LUT4 #(
		.INIT('h1500)
	) name781 (
		_w526_,
		_w771_,
		_w776_,
		_w1294_,
		_w1295_
	);
	LUT4 #(
		.INIT('h000d)
	) name782 (
		\in3[96] ,
		_w782_,
		_w1281_,
		_w1295_,
		_w1296_
	);
	LUT4 #(
		.INIT('h000d)
	) name783 (
		\in3[97] ,
		_w782_,
		_w1288_,
		_w1290_,
		_w1297_
	);
	LUT3 #(
		.INIT('ha8)
	) name784 (
		\in2[98] ,
		_w521_,
		_w778_,
		_w1298_
	);
	LUT4 #(
		.INIT('h1500)
	) name785 (
		_w526_,
		_w771_,
		_w776_,
		_w1298_,
		_w1299_
	);
	LUT4 #(
		.INIT('h000d)
	) name786 (
		\in3[98] ,
		_w782_,
		_w1273_,
		_w1299_,
		_w1300_
	);
	LUT4 #(
		.INIT('h0007)
	) name787 (
		_w1291_,
		_w1296_,
		_w1297_,
		_w1300_,
		_w1301_
	);
	LUT3 #(
		.INIT('h31)
	) name788 (
		_w1277_,
		_w1293_,
		_w1301_,
		_w1302_
	);
	LUT4 #(
		.INIT('h0301)
	) name789 (
		_w1277_,
		_w1292_,
		_w1293_,
		_w1301_,
		_w1303_
	);
	LUT3 #(
		.INIT('ha8)
	) name790 (
		\in0[87] ,
		_w1038_,
		_w1045_,
		_w1304_
	);
	LUT3 #(
		.INIT('hb0)
	) name791 (
		_w1029_,
		_w1043_,
		_w1304_,
		_w1305_
	);
	LUT4 #(
		.INIT('haa20)
	) name792 (
		\in1[87] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1306_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		_w1305_,
		_w1306_,
		_w1307_
	);
	LUT3 #(
		.INIT('ha8)
	) name794 (
		\in2[87] ,
		_w521_,
		_w778_,
		_w1308_
	);
	LUT4 #(
		.INIT('h1500)
	) name795 (
		_w526_,
		_w771_,
		_w776_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name796 (
		\in3[87] ,
		_w782_,
		_w1307_,
		_w1309_,
		_w1310_
	);
	LUT3 #(
		.INIT('ha8)
	) name797 (
		\in0[86] ,
		_w1038_,
		_w1045_,
		_w1311_
	);
	LUT3 #(
		.INIT('hb0)
	) name798 (
		_w1029_,
		_w1043_,
		_w1311_,
		_w1312_
	);
	LUT4 #(
		.INIT('haa20)
	) name799 (
		\in1[86] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1313_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w1312_,
		_w1313_,
		_w1314_
	);
	LUT3 #(
		.INIT('h02)
	) name801 (
		\in3[86] ,
		_w1312_,
		_w1313_,
		_w1315_
	);
	LUT3 #(
		.INIT('h02)
	) name802 (
		\in2[86] ,
		_w1312_,
		_w1313_,
		_w1316_
	);
	LUT3 #(
		.INIT('h1b)
	) name803 (
		_w782_,
		_w1315_,
		_w1316_,
		_w1317_
	);
	LUT2 #(
		.INIT('h8)
	) name804 (
		_w1310_,
		_w1317_,
		_w1318_
	);
	LUT3 #(
		.INIT('ha8)
	) name805 (
		\in0[84] ,
		_w1038_,
		_w1045_,
		_w1319_
	);
	LUT3 #(
		.INIT('hb0)
	) name806 (
		_w1029_,
		_w1043_,
		_w1319_,
		_w1320_
	);
	LUT4 #(
		.INIT('haa20)
	) name807 (
		\in1[84] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1321_
	);
	LUT2 #(
		.INIT('h1)
	) name808 (
		_w1320_,
		_w1321_,
		_w1322_
	);
	LUT3 #(
		.INIT('h02)
	) name809 (
		\in3[84] ,
		_w1320_,
		_w1321_,
		_w1323_
	);
	LUT3 #(
		.INIT('h02)
	) name810 (
		\in2[84] ,
		_w1320_,
		_w1321_,
		_w1324_
	);
	LUT3 #(
		.INIT('h1b)
	) name811 (
		_w782_,
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT3 #(
		.INIT('ha8)
	) name812 (
		\in0[85] ,
		_w1038_,
		_w1045_,
		_w1326_
	);
	LUT3 #(
		.INIT('hb0)
	) name813 (
		_w1029_,
		_w1043_,
		_w1326_,
		_w1327_
	);
	LUT4 #(
		.INIT('haa20)
	) name814 (
		\in1[85] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1328_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w1327_,
		_w1328_,
		_w1329_
	);
	LUT3 #(
		.INIT('ha8)
	) name816 (
		\in2[85] ,
		_w521_,
		_w778_,
		_w1330_
	);
	LUT4 #(
		.INIT('h1500)
	) name817 (
		_w526_,
		_w771_,
		_w776_,
		_w1330_,
		_w1331_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name818 (
		\in3[85] ,
		_w782_,
		_w1329_,
		_w1331_,
		_w1332_
	);
	LUT4 #(
		.INIT('h8000)
	) name819 (
		_w1310_,
		_w1317_,
		_w1325_,
		_w1332_,
		_w1333_
	);
	LUT3 #(
		.INIT('ha8)
	) name820 (
		\in0[91] ,
		_w1038_,
		_w1045_,
		_w1334_
	);
	LUT3 #(
		.INIT('hb0)
	) name821 (
		_w1029_,
		_w1043_,
		_w1334_,
		_w1335_
	);
	LUT4 #(
		.INIT('haa20)
	) name822 (
		\in1[91] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1336_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		_w1335_,
		_w1336_,
		_w1337_
	);
	LUT3 #(
		.INIT('ha8)
	) name824 (
		\in2[91] ,
		_w521_,
		_w778_,
		_w1338_
	);
	LUT4 #(
		.INIT('h1500)
	) name825 (
		_w526_,
		_w771_,
		_w776_,
		_w1338_,
		_w1339_
	);
	LUT4 #(
		.INIT('h000d)
	) name826 (
		\in3[91] ,
		_w782_,
		_w1337_,
		_w1339_,
		_w1340_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name827 (
		\in3[91] ,
		_w782_,
		_w1337_,
		_w1339_,
		_w1341_
	);
	LUT3 #(
		.INIT('ha8)
	) name828 (
		\in0[90] ,
		_w1038_,
		_w1045_,
		_w1342_
	);
	LUT3 #(
		.INIT('hb0)
	) name829 (
		_w1029_,
		_w1043_,
		_w1342_,
		_w1343_
	);
	LUT4 #(
		.INIT('haa20)
	) name830 (
		\in1[90] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1344_
	);
	LUT2 #(
		.INIT('h1)
	) name831 (
		_w1343_,
		_w1344_,
		_w1345_
	);
	LUT3 #(
		.INIT('h02)
	) name832 (
		\in3[90] ,
		_w1343_,
		_w1344_,
		_w1346_
	);
	LUT3 #(
		.INIT('h02)
	) name833 (
		\in2[90] ,
		_w1343_,
		_w1344_,
		_w1347_
	);
	LUT3 #(
		.INIT('h1b)
	) name834 (
		_w782_,
		_w1346_,
		_w1347_,
		_w1348_
	);
	LUT2 #(
		.INIT('h8)
	) name835 (
		_w1341_,
		_w1348_,
		_w1349_
	);
	LUT3 #(
		.INIT('ha8)
	) name836 (
		\in0[89] ,
		_w1038_,
		_w1045_,
		_w1350_
	);
	LUT3 #(
		.INIT('hb0)
	) name837 (
		_w1029_,
		_w1043_,
		_w1350_,
		_w1351_
	);
	LUT4 #(
		.INIT('haa20)
	) name838 (
		\in1[89] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1352_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w1351_,
		_w1352_,
		_w1353_
	);
	LUT3 #(
		.INIT('ha8)
	) name840 (
		\in2[89] ,
		_w521_,
		_w778_,
		_w1354_
	);
	LUT4 #(
		.INIT('h1500)
	) name841 (
		_w526_,
		_w771_,
		_w776_,
		_w1354_,
		_w1355_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name842 (
		\in3[89] ,
		_w782_,
		_w1353_,
		_w1355_,
		_w1356_
	);
	LUT3 #(
		.INIT('ha8)
	) name843 (
		\in2[88] ,
		_w521_,
		_w778_,
		_w1357_
	);
	LUT4 #(
		.INIT('h1500)
	) name844 (
		_w526_,
		_w771_,
		_w776_,
		_w1357_,
		_w1358_
	);
	LUT3 #(
		.INIT('ha8)
	) name845 (
		\in0[88] ,
		_w1038_,
		_w1045_,
		_w1359_
	);
	LUT3 #(
		.INIT('hb0)
	) name846 (
		_w1029_,
		_w1043_,
		_w1359_,
		_w1360_
	);
	LUT4 #(
		.INIT('haa20)
	) name847 (
		\in1[88] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1361_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w1360_,
		_w1361_,
		_w1362_
	);
	LUT4 #(
		.INIT('h000d)
	) name849 (
		\in3[88] ,
		_w782_,
		_w1358_,
		_w1362_,
		_w1363_
	);
	LUT4 #(
		.INIT('h000d)
	) name850 (
		\in3[89] ,
		_w782_,
		_w1353_,
		_w1355_,
		_w1364_
	);
	LUT3 #(
		.INIT('ha8)
	) name851 (
		\in2[90] ,
		_w521_,
		_w778_,
		_w1365_
	);
	LUT4 #(
		.INIT('h1500)
	) name852 (
		_w526_,
		_w771_,
		_w776_,
		_w1365_,
		_w1366_
	);
	LUT4 #(
		.INIT('h000d)
	) name853 (
		\in3[90] ,
		_w782_,
		_w1345_,
		_w1366_,
		_w1367_
	);
	LUT4 #(
		.INIT('h0007)
	) name854 (
		_w1356_,
		_w1363_,
		_w1364_,
		_w1367_,
		_w1368_
	);
	LUT3 #(
		.INIT('h51)
	) name855 (
		_w1340_,
		_w1349_,
		_w1368_,
		_w1369_
	);
	LUT4 #(
		.INIT('h000d)
	) name856 (
		\in3[87] ,
		_w782_,
		_w1307_,
		_w1309_,
		_w1370_
	);
	LUT3 #(
		.INIT('ha8)
	) name857 (
		\in2[84] ,
		_w521_,
		_w778_,
		_w1371_
	);
	LUT4 #(
		.INIT('h1500)
	) name858 (
		_w526_,
		_w771_,
		_w776_,
		_w1371_,
		_w1372_
	);
	LUT4 #(
		.INIT('h000d)
	) name859 (
		\in3[84] ,
		_w782_,
		_w1322_,
		_w1372_,
		_w1373_
	);
	LUT3 #(
		.INIT('ha8)
	) name860 (
		\in2[86] ,
		_w521_,
		_w778_,
		_w1374_
	);
	LUT4 #(
		.INIT('h1500)
	) name861 (
		_w526_,
		_w771_,
		_w776_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('h000d)
	) name862 (
		\in3[86] ,
		_w782_,
		_w1314_,
		_w1375_,
		_w1376_
	);
	LUT4 #(
		.INIT('h000d)
	) name863 (
		\in3[85] ,
		_w782_,
		_w1329_,
		_w1331_,
		_w1377_
	);
	LUT4 #(
		.INIT('h0007)
	) name864 (
		_w1332_,
		_w1373_,
		_w1376_,
		_w1377_,
		_w1378_
	);
	LUT3 #(
		.INIT('h31)
	) name865 (
		_w1318_,
		_w1370_,
		_w1378_,
		_w1379_
	);
	LUT3 #(
		.INIT('h40)
	) name866 (
		_w1333_,
		_w1369_,
		_w1379_,
		_w1380_
	);
	LUT3 #(
		.INIT('ha8)
	) name867 (
		\in0[79] ,
		_w1038_,
		_w1045_,
		_w1381_
	);
	LUT3 #(
		.INIT('hb0)
	) name868 (
		_w1029_,
		_w1043_,
		_w1381_,
		_w1382_
	);
	LUT4 #(
		.INIT('haa20)
	) name869 (
		\in1[79] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1383_
	);
	LUT2 #(
		.INIT('h1)
	) name870 (
		_w1382_,
		_w1383_,
		_w1384_
	);
	LUT3 #(
		.INIT('ha8)
	) name871 (
		\in2[79] ,
		_w521_,
		_w778_,
		_w1385_
	);
	LUT4 #(
		.INIT('h1500)
	) name872 (
		_w526_,
		_w771_,
		_w776_,
		_w1385_,
		_w1386_
	);
	LUT4 #(
		.INIT('h000d)
	) name873 (
		\in3[79] ,
		_w782_,
		_w1384_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name874 (
		\in3[79] ,
		_w782_,
		_w1384_,
		_w1386_,
		_w1388_
	);
	LUT3 #(
		.INIT('ha8)
	) name875 (
		\in0[78] ,
		_w1038_,
		_w1045_,
		_w1389_
	);
	LUT3 #(
		.INIT('hb0)
	) name876 (
		_w1029_,
		_w1043_,
		_w1389_,
		_w1390_
	);
	LUT4 #(
		.INIT('haa20)
	) name877 (
		\in1[78] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1391_
	);
	LUT2 #(
		.INIT('h1)
	) name878 (
		_w1390_,
		_w1391_,
		_w1392_
	);
	LUT3 #(
		.INIT('h02)
	) name879 (
		\in3[78] ,
		_w1390_,
		_w1391_,
		_w1393_
	);
	LUT3 #(
		.INIT('h02)
	) name880 (
		\in2[78] ,
		_w1390_,
		_w1391_,
		_w1394_
	);
	LUT3 #(
		.INIT('h1b)
	) name881 (
		_w782_,
		_w1393_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		_w1388_,
		_w1395_,
		_w1396_
	);
	LUT3 #(
		.INIT('ha8)
	) name883 (
		\in0[77] ,
		_w1038_,
		_w1045_,
		_w1397_
	);
	LUT3 #(
		.INIT('hb0)
	) name884 (
		_w1029_,
		_w1043_,
		_w1397_,
		_w1398_
	);
	LUT4 #(
		.INIT('haa20)
	) name885 (
		\in1[77] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1399_
	);
	LUT2 #(
		.INIT('h1)
	) name886 (
		_w1398_,
		_w1399_,
		_w1400_
	);
	LUT3 #(
		.INIT('ha8)
	) name887 (
		\in2[77] ,
		_w521_,
		_w778_,
		_w1401_
	);
	LUT4 #(
		.INIT('h1500)
	) name888 (
		_w526_,
		_w771_,
		_w776_,
		_w1401_,
		_w1402_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name889 (
		\in3[77] ,
		_w782_,
		_w1400_,
		_w1402_,
		_w1403_
	);
	LUT3 #(
		.INIT('ha8)
	) name890 (
		\in2[76] ,
		_w521_,
		_w778_,
		_w1404_
	);
	LUT4 #(
		.INIT('h1500)
	) name891 (
		_w526_,
		_w771_,
		_w776_,
		_w1404_,
		_w1405_
	);
	LUT3 #(
		.INIT('ha8)
	) name892 (
		\in0[76] ,
		_w1038_,
		_w1045_,
		_w1406_
	);
	LUT3 #(
		.INIT('hb0)
	) name893 (
		_w1029_,
		_w1043_,
		_w1406_,
		_w1407_
	);
	LUT4 #(
		.INIT('haa20)
	) name894 (
		\in1[76] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1408_
	);
	LUT2 #(
		.INIT('h1)
	) name895 (
		_w1407_,
		_w1408_,
		_w1409_
	);
	LUT4 #(
		.INIT('h000d)
	) name896 (
		\in3[76] ,
		_w782_,
		_w1405_,
		_w1409_,
		_w1410_
	);
	LUT3 #(
		.INIT('ha8)
	) name897 (
		\in2[78] ,
		_w521_,
		_w778_,
		_w1411_
	);
	LUT4 #(
		.INIT('h1500)
	) name898 (
		_w526_,
		_w771_,
		_w776_,
		_w1411_,
		_w1412_
	);
	LUT4 #(
		.INIT('h000d)
	) name899 (
		\in3[78] ,
		_w782_,
		_w1392_,
		_w1412_,
		_w1413_
	);
	LUT4 #(
		.INIT('h000d)
	) name900 (
		\in3[77] ,
		_w782_,
		_w1400_,
		_w1402_,
		_w1414_
	);
	LUT4 #(
		.INIT('h0007)
	) name901 (
		_w1403_,
		_w1410_,
		_w1413_,
		_w1414_,
		_w1415_
	);
	LUT3 #(
		.INIT('ha8)
	) name902 (
		\in0[83] ,
		_w1038_,
		_w1045_,
		_w1416_
	);
	LUT3 #(
		.INIT('hb0)
	) name903 (
		_w1029_,
		_w1043_,
		_w1416_,
		_w1417_
	);
	LUT4 #(
		.INIT('haa20)
	) name904 (
		\in1[83] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1418_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT3 #(
		.INIT('ha8)
	) name906 (
		\in2[83] ,
		_w521_,
		_w778_,
		_w1420_
	);
	LUT4 #(
		.INIT('h1500)
	) name907 (
		_w526_,
		_w771_,
		_w776_,
		_w1420_,
		_w1421_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name908 (
		\in3[83] ,
		_w782_,
		_w1419_,
		_w1421_,
		_w1422_
	);
	LUT3 #(
		.INIT('ha8)
	) name909 (
		\in0[82] ,
		_w1038_,
		_w1045_,
		_w1423_
	);
	LUT3 #(
		.INIT('hb0)
	) name910 (
		_w1029_,
		_w1043_,
		_w1423_,
		_w1424_
	);
	LUT4 #(
		.INIT('haa20)
	) name911 (
		\in1[82] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1425_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1424_,
		_w1425_,
		_w1426_
	);
	LUT3 #(
		.INIT('h02)
	) name913 (
		\in3[82] ,
		_w1424_,
		_w1425_,
		_w1427_
	);
	LUT3 #(
		.INIT('h02)
	) name914 (
		\in2[82] ,
		_w1424_,
		_w1425_,
		_w1428_
	);
	LUT3 #(
		.INIT('h1b)
	) name915 (
		_w782_,
		_w1427_,
		_w1428_,
		_w1429_
	);
	LUT2 #(
		.INIT('h8)
	) name916 (
		_w1422_,
		_w1429_,
		_w1430_
	);
	LUT3 #(
		.INIT('ha8)
	) name917 (
		\in0[81] ,
		_w1038_,
		_w1045_,
		_w1431_
	);
	LUT3 #(
		.INIT('hb0)
	) name918 (
		_w1029_,
		_w1043_,
		_w1431_,
		_w1432_
	);
	LUT4 #(
		.INIT('haa20)
	) name919 (
		\in1[81] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1433_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1432_,
		_w1433_,
		_w1434_
	);
	LUT3 #(
		.INIT('ha8)
	) name921 (
		\in2[81] ,
		_w521_,
		_w778_,
		_w1435_
	);
	LUT4 #(
		.INIT('h1500)
	) name922 (
		_w526_,
		_w771_,
		_w776_,
		_w1435_,
		_w1436_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name923 (
		\in3[81] ,
		_w782_,
		_w1434_,
		_w1436_,
		_w1437_
	);
	LUT3 #(
		.INIT('ha8)
	) name924 (
		\in0[80] ,
		_w1038_,
		_w1045_,
		_w1438_
	);
	LUT3 #(
		.INIT('hb0)
	) name925 (
		_w1029_,
		_w1043_,
		_w1438_,
		_w1439_
	);
	LUT4 #(
		.INIT('haa20)
	) name926 (
		\in1[80] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1440_
	);
	LUT2 #(
		.INIT('h1)
	) name927 (
		_w1439_,
		_w1440_,
		_w1441_
	);
	LUT3 #(
		.INIT('h02)
	) name928 (
		\in3[80] ,
		_w1439_,
		_w1440_,
		_w1442_
	);
	LUT3 #(
		.INIT('h02)
	) name929 (
		\in2[80] ,
		_w1439_,
		_w1440_,
		_w1443_
	);
	LUT3 #(
		.INIT('h1b)
	) name930 (
		_w782_,
		_w1442_,
		_w1443_,
		_w1444_
	);
	LUT4 #(
		.INIT('h8000)
	) name931 (
		_w1422_,
		_w1429_,
		_w1437_,
		_w1444_,
		_w1445_
	);
	LUT4 #(
		.INIT('hae00)
	) name932 (
		_w1387_,
		_w1396_,
		_w1415_,
		_w1445_,
		_w1446_
	);
	LUT3 #(
		.INIT('ha8)
	) name933 (
		\in0[75] ,
		_w1038_,
		_w1045_,
		_w1447_
	);
	LUT3 #(
		.INIT('hb0)
	) name934 (
		_w1029_,
		_w1043_,
		_w1447_,
		_w1448_
	);
	LUT4 #(
		.INIT('haa20)
	) name935 (
		\in1[75] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1449_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1448_,
		_w1449_,
		_w1450_
	);
	LUT3 #(
		.INIT('ha8)
	) name937 (
		\in2[75] ,
		_w521_,
		_w778_,
		_w1451_
	);
	LUT4 #(
		.INIT('h1500)
	) name938 (
		_w526_,
		_w771_,
		_w776_,
		_w1451_,
		_w1452_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name939 (
		\in3[75] ,
		_w782_,
		_w1450_,
		_w1452_,
		_w1453_
	);
	LUT3 #(
		.INIT('ha8)
	) name940 (
		\in0[74] ,
		_w1038_,
		_w1045_,
		_w1454_
	);
	LUT3 #(
		.INIT('hb0)
	) name941 (
		_w1029_,
		_w1043_,
		_w1454_,
		_w1455_
	);
	LUT4 #(
		.INIT('haa20)
	) name942 (
		\in1[74] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1456_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		_w1455_,
		_w1456_,
		_w1457_
	);
	LUT3 #(
		.INIT('h02)
	) name944 (
		\in3[74] ,
		_w1455_,
		_w1456_,
		_w1458_
	);
	LUT3 #(
		.INIT('h02)
	) name945 (
		\in2[74] ,
		_w1455_,
		_w1456_,
		_w1459_
	);
	LUT3 #(
		.INIT('h1b)
	) name946 (
		_w782_,
		_w1458_,
		_w1459_,
		_w1460_
	);
	LUT2 #(
		.INIT('h8)
	) name947 (
		_w1453_,
		_w1460_,
		_w1461_
	);
	LUT3 #(
		.INIT('ha8)
	) name948 (
		\in0[72] ,
		_w1038_,
		_w1045_,
		_w1462_
	);
	LUT3 #(
		.INIT('hb0)
	) name949 (
		_w1029_,
		_w1043_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('haa20)
	) name950 (
		\in1[72] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1464_
	);
	LUT2 #(
		.INIT('h1)
	) name951 (
		_w1463_,
		_w1464_,
		_w1465_
	);
	LUT3 #(
		.INIT('h02)
	) name952 (
		\in3[72] ,
		_w1463_,
		_w1464_,
		_w1466_
	);
	LUT3 #(
		.INIT('h02)
	) name953 (
		\in2[72] ,
		_w1463_,
		_w1464_,
		_w1467_
	);
	LUT3 #(
		.INIT('h1b)
	) name954 (
		_w782_,
		_w1466_,
		_w1467_,
		_w1468_
	);
	LUT3 #(
		.INIT('ha8)
	) name955 (
		\in0[73] ,
		_w1038_,
		_w1045_,
		_w1469_
	);
	LUT3 #(
		.INIT('hb0)
	) name956 (
		_w1029_,
		_w1043_,
		_w1469_,
		_w1470_
	);
	LUT4 #(
		.INIT('haa20)
	) name957 (
		\in1[73] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1471_
	);
	LUT2 #(
		.INIT('h1)
	) name958 (
		_w1470_,
		_w1471_,
		_w1472_
	);
	LUT3 #(
		.INIT('ha8)
	) name959 (
		\in2[73] ,
		_w521_,
		_w778_,
		_w1473_
	);
	LUT4 #(
		.INIT('h1500)
	) name960 (
		_w526_,
		_w771_,
		_w776_,
		_w1473_,
		_w1474_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name961 (
		\in3[73] ,
		_w782_,
		_w1472_,
		_w1474_,
		_w1475_
	);
	LUT4 #(
		.INIT('h8000)
	) name962 (
		_w1453_,
		_w1460_,
		_w1468_,
		_w1475_,
		_w1476_
	);
	LUT4 #(
		.INIT('h000d)
	) name963 (
		\in3[75] ,
		_w782_,
		_w1450_,
		_w1452_,
		_w1477_
	);
	LUT3 #(
		.INIT('ha8)
	) name964 (
		\in2[72] ,
		_w521_,
		_w778_,
		_w1478_
	);
	LUT4 #(
		.INIT('h1500)
	) name965 (
		_w526_,
		_w771_,
		_w776_,
		_w1478_,
		_w1479_
	);
	LUT4 #(
		.INIT('h000d)
	) name966 (
		\in3[72] ,
		_w782_,
		_w1465_,
		_w1479_,
		_w1480_
	);
	LUT4 #(
		.INIT('h000d)
	) name967 (
		\in3[73] ,
		_w782_,
		_w1472_,
		_w1474_,
		_w1481_
	);
	LUT3 #(
		.INIT('ha8)
	) name968 (
		\in2[74] ,
		_w521_,
		_w778_,
		_w1482_
	);
	LUT4 #(
		.INIT('h1500)
	) name969 (
		_w526_,
		_w771_,
		_w776_,
		_w1482_,
		_w1483_
	);
	LUT4 #(
		.INIT('h000d)
	) name970 (
		\in3[74] ,
		_w782_,
		_w1457_,
		_w1483_,
		_w1484_
	);
	LUT4 #(
		.INIT('h0007)
	) name971 (
		_w1475_,
		_w1480_,
		_w1481_,
		_w1484_,
		_w1485_
	);
	LUT3 #(
		.INIT('h31)
	) name972 (
		_w1461_,
		_w1477_,
		_w1485_,
		_w1486_
	);
	LUT4 #(
		.INIT('h0301)
	) name973 (
		_w1461_,
		_w1476_,
		_w1477_,
		_w1485_,
		_w1487_
	);
	LUT3 #(
		.INIT('ha8)
	) name974 (
		\in0[67] ,
		_w1038_,
		_w1045_,
		_w1488_
	);
	LUT3 #(
		.INIT('hb0)
	) name975 (
		_w1029_,
		_w1043_,
		_w1488_,
		_w1489_
	);
	LUT4 #(
		.INIT('haa20)
	) name976 (
		\in1[67] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1490_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		_w1489_,
		_w1490_,
		_w1491_
	);
	LUT3 #(
		.INIT('ha8)
	) name978 (
		\in2[67] ,
		_w521_,
		_w778_,
		_w1492_
	);
	LUT4 #(
		.INIT('h1500)
	) name979 (
		_w526_,
		_w771_,
		_w776_,
		_w1492_,
		_w1493_
	);
	LUT4 #(
		.INIT('h000d)
	) name980 (
		\in3[67] ,
		_w782_,
		_w1491_,
		_w1493_,
		_w1494_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name981 (
		\in3[67] ,
		_w782_,
		_w1491_,
		_w1493_,
		_w1495_
	);
	LUT3 #(
		.INIT('ha8)
	) name982 (
		\in0[66] ,
		_w1038_,
		_w1045_,
		_w1496_
	);
	LUT3 #(
		.INIT('hb0)
	) name983 (
		_w1029_,
		_w1043_,
		_w1496_,
		_w1497_
	);
	LUT4 #(
		.INIT('haa20)
	) name984 (
		\in1[66] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1498_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		_w1497_,
		_w1498_,
		_w1499_
	);
	LUT3 #(
		.INIT('h02)
	) name986 (
		\in3[66] ,
		_w1497_,
		_w1498_,
		_w1500_
	);
	LUT3 #(
		.INIT('h02)
	) name987 (
		\in2[66] ,
		_w1497_,
		_w1498_,
		_w1501_
	);
	LUT3 #(
		.INIT('h1b)
	) name988 (
		_w782_,
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT2 #(
		.INIT('h8)
	) name989 (
		_w1495_,
		_w1502_,
		_w1503_
	);
	LUT3 #(
		.INIT('ha8)
	) name990 (
		\in0[65] ,
		_w1038_,
		_w1045_,
		_w1504_
	);
	LUT3 #(
		.INIT('hb0)
	) name991 (
		_w1029_,
		_w1043_,
		_w1504_,
		_w1505_
	);
	LUT4 #(
		.INIT('haa20)
	) name992 (
		\in1[65] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1506_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		_w1505_,
		_w1506_,
		_w1507_
	);
	LUT3 #(
		.INIT('ha8)
	) name994 (
		\in2[65] ,
		_w521_,
		_w778_,
		_w1508_
	);
	LUT4 #(
		.INIT('h1500)
	) name995 (
		_w526_,
		_w771_,
		_w776_,
		_w1508_,
		_w1509_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name996 (
		\in3[65] ,
		_w782_,
		_w1507_,
		_w1509_,
		_w1510_
	);
	LUT3 #(
		.INIT('ha8)
	) name997 (
		\in2[64] ,
		_w521_,
		_w778_,
		_w1511_
	);
	LUT4 #(
		.INIT('h1500)
	) name998 (
		_w526_,
		_w771_,
		_w776_,
		_w1511_,
		_w1512_
	);
	LUT3 #(
		.INIT('ha8)
	) name999 (
		\in0[64] ,
		_w1038_,
		_w1045_,
		_w1513_
	);
	LUT3 #(
		.INIT('hb0)
	) name1000 (
		_w1029_,
		_w1043_,
		_w1513_,
		_w1514_
	);
	LUT4 #(
		.INIT('haa20)
	) name1001 (
		\in1[64] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1515_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1514_,
		_w1515_,
		_w1516_
	);
	LUT4 #(
		.INIT('h000d)
	) name1003 (
		\in3[64] ,
		_w782_,
		_w1512_,
		_w1516_,
		_w1517_
	);
	LUT4 #(
		.INIT('h000d)
	) name1004 (
		\in3[65] ,
		_w782_,
		_w1507_,
		_w1509_,
		_w1518_
	);
	LUT3 #(
		.INIT('ha8)
	) name1005 (
		\in2[66] ,
		_w521_,
		_w778_,
		_w1519_
	);
	LUT4 #(
		.INIT('h1500)
	) name1006 (
		_w526_,
		_w771_,
		_w776_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h000d)
	) name1007 (
		\in3[66] ,
		_w782_,
		_w1499_,
		_w1520_,
		_w1521_
	);
	LUT4 #(
		.INIT('h0007)
	) name1008 (
		_w1510_,
		_w1517_,
		_w1518_,
		_w1521_,
		_w1522_
	);
	LUT3 #(
		.INIT('ha8)
	) name1009 (
		\in0[71] ,
		_w1038_,
		_w1045_,
		_w1523_
	);
	LUT3 #(
		.INIT('hb0)
	) name1010 (
		_w1029_,
		_w1043_,
		_w1523_,
		_w1524_
	);
	LUT4 #(
		.INIT('haa20)
	) name1011 (
		\in1[71] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1525_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w1524_,
		_w1525_,
		_w1526_
	);
	LUT3 #(
		.INIT('ha8)
	) name1013 (
		\in2[71] ,
		_w521_,
		_w778_,
		_w1527_
	);
	LUT4 #(
		.INIT('h1500)
	) name1014 (
		_w526_,
		_w771_,
		_w776_,
		_w1527_,
		_w1528_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1015 (
		\in3[71] ,
		_w782_,
		_w1526_,
		_w1528_,
		_w1529_
	);
	LUT3 #(
		.INIT('ha8)
	) name1016 (
		\in0[70] ,
		_w1038_,
		_w1045_,
		_w1530_
	);
	LUT3 #(
		.INIT('hb0)
	) name1017 (
		_w1029_,
		_w1043_,
		_w1530_,
		_w1531_
	);
	LUT4 #(
		.INIT('haa20)
	) name1018 (
		\in1[70] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1532_
	);
	LUT2 #(
		.INIT('h1)
	) name1019 (
		_w1531_,
		_w1532_,
		_w1533_
	);
	LUT3 #(
		.INIT('h02)
	) name1020 (
		\in3[70] ,
		_w1531_,
		_w1532_,
		_w1534_
	);
	LUT3 #(
		.INIT('h02)
	) name1021 (
		\in2[70] ,
		_w1531_,
		_w1532_,
		_w1535_
	);
	LUT3 #(
		.INIT('h1b)
	) name1022 (
		_w782_,
		_w1534_,
		_w1535_,
		_w1536_
	);
	LUT2 #(
		.INIT('h8)
	) name1023 (
		_w1529_,
		_w1536_,
		_w1537_
	);
	LUT3 #(
		.INIT('ha8)
	) name1024 (
		\in0[69] ,
		_w1038_,
		_w1045_,
		_w1538_
	);
	LUT3 #(
		.INIT('hb0)
	) name1025 (
		_w1029_,
		_w1043_,
		_w1538_,
		_w1539_
	);
	LUT4 #(
		.INIT('haa20)
	) name1026 (
		\in1[69] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1540_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		_w1539_,
		_w1540_,
		_w1541_
	);
	LUT3 #(
		.INIT('ha8)
	) name1028 (
		\in2[69] ,
		_w521_,
		_w778_,
		_w1542_
	);
	LUT4 #(
		.INIT('h1500)
	) name1029 (
		_w526_,
		_w771_,
		_w776_,
		_w1542_,
		_w1543_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1030 (
		\in3[69] ,
		_w782_,
		_w1541_,
		_w1543_,
		_w1544_
	);
	LUT3 #(
		.INIT('ha8)
	) name1031 (
		\in0[68] ,
		_w1038_,
		_w1045_,
		_w1545_
	);
	LUT3 #(
		.INIT('hb0)
	) name1032 (
		_w1029_,
		_w1043_,
		_w1545_,
		_w1546_
	);
	LUT4 #(
		.INIT('haa20)
	) name1033 (
		\in1[68] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1547_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w1546_,
		_w1547_,
		_w1548_
	);
	LUT3 #(
		.INIT('h02)
	) name1035 (
		\in3[68] ,
		_w1546_,
		_w1547_,
		_w1549_
	);
	LUT3 #(
		.INIT('h02)
	) name1036 (
		\in2[68] ,
		_w1546_,
		_w1547_,
		_w1550_
	);
	LUT3 #(
		.INIT('h1b)
	) name1037 (
		_w782_,
		_w1549_,
		_w1550_,
		_w1551_
	);
	LUT4 #(
		.INIT('h8000)
	) name1038 (
		_w1529_,
		_w1536_,
		_w1544_,
		_w1551_,
		_w1552_
	);
	LUT4 #(
		.INIT('hae00)
	) name1039 (
		_w1494_,
		_w1503_,
		_w1522_,
		_w1552_,
		_w1553_
	);
	LUT3 #(
		.INIT('ha8)
	) name1040 (
		\in0[63] ,
		_w1038_,
		_w1045_,
		_w1554_
	);
	LUT3 #(
		.INIT('hb0)
	) name1041 (
		_w1029_,
		_w1043_,
		_w1554_,
		_w1555_
	);
	LUT4 #(
		.INIT('haa20)
	) name1042 (
		\in1[63] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1556_
	);
	LUT2 #(
		.INIT('h1)
	) name1043 (
		_w1555_,
		_w1556_,
		_w1557_
	);
	LUT3 #(
		.INIT('ha8)
	) name1044 (
		\in2[63] ,
		_w521_,
		_w778_,
		_w1558_
	);
	LUT4 #(
		.INIT('h1500)
	) name1045 (
		_w526_,
		_w771_,
		_w776_,
		_w1558_,
		_w1559_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1046 (
		\in3[63] ,
		_w782_,
		_w1557_,
		_w1559_,
		_w1560_
	);
	LUT3 #(
		.INIT('ha8)
	) name1047 (
		\in0[61] ,
		_w1038_,
		_w1045_,
		_w1561_
	);
	LUT3 #(
		.INIT('hb0)
	) name1048 (
		_w1029_,
		_w1043_,
		_w1561_,
		_w1562_
	);
	LUT4 #(
		.INIT('haa20)
	) name1049 (
		\in1[61] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1563_
	);
	LUT2 #(
		.INIT('h1)
	) name1050 (
		_w1562_,
		_w1563_,
		_w1564_
	);
	LUT3 #(
		.INIT('ha8)
	) name1051 (
		\in2[61] ,
		_w521_,
		_w778_,
		_w1565_
	);
	LUT4 #(
		.INIT('h1500)
	) name1052 (
		_w526_,
		_w771_,
		_w776_,
		_w1565_,
		_w1566_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1053 (
		\in3[61] ,
		_w782_,
		_w1564_,
		_w1566_,
		_w1567_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		_w1560_,
		_w1567_,
		_w1568_
	);
	LUT3 #(
		.INIT('ha8)
	) name1055 (
		\in0[59] ,
		_w1038_,
		_w1045_,
		_w1569_
	);
	LUT3 #(
		.INIT('hb0)
	) name1056 (
		_w1029_,
		_w1043_,
		_w1569_,
		_w1570_
	);
	LUT4 #(
		.INIT('haa20)
	) name1057 (
		\in1[59] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1571_
	);
	LUT2 #(
		.INIT('h1)
	) name1058 (
		_w1570_,
		_w1571_,
		_w1572_
	);
	LUT3 #(
		.INIT('ha8)
	) name1059 (
		\in2[59] ,
		_w521_,
		_w778_,
		_w1573_
	);
	LUT4 #(
		.INIT('h1500)
	) name1060 (
		_w526_,
		_w771_,
		_w776_,
		_w1573_,
		_w1574_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1061 (
		\in3[59] ,
		_w782_,
		_w1572_,
		_w1574_,
		_w1575_
	);
	LUT3 #(
		.INIT('ha8)
	) name1062 (
		\in0[58] ,
		_w1038_,
		_w1045_,
		_w1576_
	);
	LUT3 #(
		.INIT('hb0)
	) name1063 (
		_w1029_,
		_w1043_,
		_w1576_,
		_w1577_
	);
	LUT4 #(
		.INIT('haa20)
	) name1064 (
		\in1[58] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name1065 (
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT3 #(
		.INIT('ha8)
	) name1066 (
		\in2[58] ,
		_w521_,
		_w778_,
		_w1580_
	);
	LUT4 #(
		.INIT('h1500)
	) name1067 (
		_w526_,
		_w771_,
		_w776_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1068 (
		\in3[58] ,
		_w782_,
		_w1579_,
		_w1581_,
		_w1582_
	);
	LUT3 #(
		.INIT('ha8)
	) name1069 (
		\in0[60] ,
		_w1038_,
		_w1045_,
		_w1583_
	);
	LUT3 #(
		.INIT('hb0)
	) name1070 (
		_w1029_,
		_w1043_,
		_w1583_,
		_w1584_
	);
	LUT4 #(
		.INIT('haa20)
	) name1071 (
		\in1[60] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1585_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w1584_,
		_w1585_,
		_w1586_
	);
	LUT3 #(
		.INIT('ha8)
	) name1073 (
		\in2[60] ,
		_w521_,
		_w778_,
		_w1587_
	);
	LUT4 #(
		.INIT('h1500)
	) name1074 (
		_w526_,
		_w771_,
		_w776_,
		_w1587_,
		_w1588_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1075 (
		\in3[60] ,
		_w782_,
		_w1586_,
		_w1588_,
		_w1589_
	);
	LUT3 #(
		.INIT('h80)
	) name1076 (
		_w1575_,
		_w1582_,
		_w1589_,
		_w1590_
	);
	LUT3 #(
		.INIT('ha8)
	) name1077 (
		\in0[62] ,
		_w1038_,
		_w1045_,
		_w1591_
	);
	LUT3 #(
		.INIT('hb0)
	) name1078 (
		_w1029_,
		_w1043_,
		_w1591_,
		_w1592_
	);
	LUT4 #(
		.INIT('haa20)
	) name1079 (
		\in1[62] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name1080 (
		_w1592_,
		_w1593_,
		_w1594_
	);
	LUT3 #(
		.INIT('h02)
	) name1081 (
		\in3[62] ,
		_w1592_,
		_w1593_,
		_w1595_
	);
	LUT3 #(
		.INIT('h02)
	) name1082 (
		\in2[62] ,
		_w1592_,
		_w1593_,
		_w1596_
	);
	LUT3 #(
		.INIT('h1b)
	) name1083 (
		_w782_,
		_w1595_,
		_w1596_,
		_w1597_
	);
	LUT3 #(
		.INIT('ha8)
	) name1084 (
		\in0[57] ,
		_w1038_,
		_w1045_,
		_w1598_
	);
	LUT3 #(
		.INIT('hb0)
	) name1085 (
		_w1029_,
		_w1043_,
		_w1598_,
		_w1599_
	);
	LUT4 #(
		.INIT('haa20)
	) name1086 (
		\in1[57] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1600_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT3 #(
		.INIT('ha8)
	) name1088 (
		\in2[57] ,
		_w521_,
		_w778_,
		_w1602_
	);
	LUT4 #(
		.INIT('h1500)
	) name1089 (
		_w526_,
		_w771_,
		_w776_,
		_w1602_,
		_w1603_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1090 (
		\in3[57] ,
		_w782_,
		_w1601_,
		_w1603_,
		_w1604_
	);
	LUT3 #(
		.INIT('ha8)
	) name1091 (
		\in0[56] ,
		_w1038_,
		_w1045_,
		_w1605_
	);
	LUT3 #(
		.INIT('hb0)
	) name1092 (
		_w1029_,
		_w1043_,
		_w1605_,
		_w1606_
	);
	LUT4 #(
		.INIT('haa20)
	) name1093 (
		\in1[56] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1607_
	);
	LUT2 #(
		.INIT('h1)
	) name1094 (
		_w1606_,
		_w1607_,
		_w1608_
	);
	LUT3 #(
		.INIT('ha8)
	) name1095 (
		\in2[56] ,
		_w521_,
		_w778_,
		_w1609_
	);
	LUT4 #(
		.INIT('h1500)
	) name1096 (
		_w526_,
		_w771_,
		_w776_,
		_w1609_,
		_w1610_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1097 (
		\in3[56] ,
		_w782_,
		_w1608_,
		_w1610_,
		_w1611_
	);
	LUT3 #(
		.INIT('h80)
	) name1098 (
		_w1597_,
		_w1604_,
		_w1611_,
		_w1612_
	);
	LUT3 #(
		.INIT('h80)
	) name1099 (
		_w1568_,
		_w1590_,
		_w1612_,
		_w1613_
	);
	LUT3 #(
		.INIT('ha8)
	) name1100 (
		\in2[62] ,
		_w521_,
		_w778_,
		_w1614_
	);
	LUT4 #(
		.INIT('h1500)
	) name1101 (
		_w526_,
		_w771_,
		_w776_,
		_w1614_,
		_w1615_
	);
	LUT4 #(
		.INIT('h000d)
	) name1102 (
		\in3[62] ,
		_w782_,
		_w1594_,
		_w1615_,
		_w1616_
	);
	LUT4 #(
		.INIT('h000d)
	) name1103 (
		\in3[63] ,
		_w782_,
		_w1557_,
		_w1559_,
		_w1617_
	);
	LUT3 #(
		.INIT('h07)
	) name1104 (
		_w1560_,
		_w1616_,
		_w1617_,
		_w1618_
	);
	LUT3 #(
		.INIT('h80)
	) name1105 (
		_w1560_,
		_w1567_,
		_w1597_,
		_w1619_
	);
	LUT4 #(
		.INIT('h000d)
	) name1106 (
		\in3[56] ,
		_w782_,
		_w1608_,
		_w1610_,
		_w1620_
	);
	LUT4 #(
		.INIT('h000d)
	) name1107 (
		\in3[58] ,
		_w782_,
		_w1579_,
		_w1581_,
		_w1621_
	);
	LUT4 #(
		.INIT('h000d)
	) name1108 (
		\in3[57] ,
		_w782_,
		_w1601_,
		_w1603_,
		_w1622_
	);
	LUT4 #(
		.INIT('h0007)
	) name1109 (
		_w1604_,
		_w1620_,
		_w1621_,
		_w1622_,
		_w1623_
	);
	LUT4 #(
		.INIT('h000d)
	) name1110 (
		\in3[59] ,
		_w782_,
		_w1572_,
		_w1574_,
		_w1624_
	);
	LUT4 #(
		.INIT('h000d)
	) name1111 (
		\in3[60] ,
		_w782_,
		_w1586_,
		_w1588_,
		_w1625_
	);
	LUT4 #(
		.INIT('h000d)
	) name1112 (
		\in3[61] ,
		_w782_,
		_w1564_,
		_w1566_,
		_w1626_
	);
	LUT4 #(
		.INIT('h0007)
	) name1113 (
		_w1589_,
		_w1624_,
		_w1625_,
		_w1626_,
		_w1627_
	);
	LUT4 #(
		.INIT('h08cc)
	) name1114 (
		_w1590_,
		_w1619_,
		_w1623_,
		_w1627_,
		_w1628_
	);
	LUT3 #(
		.INIT('h04)
	) name1115 (
		_w1613_,
		_w1618_,
		_w1628_,
		_w1629_
	);
	LUT3 #(
		.INIT('ha8)
	) name1116 (
		\in0[28] ,
		_w1038_,
		_w1045_,
		_w1630_
	);
	LUT3 #(
		.INIT('hb0)
	) name1117 (
		_w1029_,
		_w1043_,
		_w1630_,
		_w1631_
	);
	LUT4 #(
		.INIT('haa20)
	) name1118 (
		\in1[28] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name1119 (
		_w1631_,
		_w1632_,
		_w1633_
	);
	LUT3 #(
		.INIT('ha8)
	) name1120 (
		\in2[28] ,
		_w521_,
		_w778_,
		_w1634_
	);
	LUT4 #(
		.INIT('h1500)
	) name1121 (
		_w526_,
		_w771_,
		_w776_,
		_w1634_,
		_w1635_
	);
	LUT4 #(
		.INIT('h000d)
	) name1122 (
		\in3[28] ,
		_w782_,
		_w1633_,
		_w1635_,
		_w1636_
	);
	LUT3 #(
		.INIT('ha8)
	) name1123 (
		\in0[29] ,
		_w1038_,
		_w1045_,
		_w1637_
	);
	LUT3 #(
		.INIT('hb0)
	) name1124 (
		_w1029_,
		_w1043_,
		_w1637_,
		_w1638_
	);
	LUT4 #(
		.INIT('haa20)
	) name1125 (
		\in1[29] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name1126 (
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT3 #(
		.INIT('ha8)
	) name1127 (
		\in2[29] ,
		_w521_,
		_w778_,
		_w1641_
	);
	LUT4 #(
		.INIT('h1500)
	) name1128 (
		_w526_,
		_w771_,
		_w776_,
		_w1641_,
		_w1642_
	);
	LUT4 #(
		.INIT('h000d)
	) name1129 (
		\in3[29] ,
		_w782_,
		_w1640_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h1)
	) name1130 (
		_w1636_,
		_w1643_,
		_w1644_
	);
	LUT3 #(
		.INIT('ha8)
	) name1131 (
		\in0[34] ,
		_w1038_,
		_w1045_,
		_w1645_
	);
	LUT3 #(
		.INIT('hb0)
	) name1132 (
		_w1029_,
		_w1043_,
		_w1645_,
		_w1646_
	);
	LUT4 #(
		.INIT('haa20)
	) name1133 (
		\in1[34] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1647_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		_w1646_,
		_w1647_,
		_w1648_
	);
	LUT3 #(
		.INIT('h02)
	) name1135 (
		\in3[34] ,
		_w1646_,
		_w1647_,
		_w1649_
	);
	LUT3 #(
		.INIT('h02)
	) name1136 (
		\in2[34] ,
		_w1646_,
		_w1647_,
		_w1650_
	);
	LUT3 #(
		.INIT('h1b)
	) name1137 (
		_w782_,
		_w1649_,
		_w1650_,
		_w1651_
	);
	LUT3 #(
		.INIT('ha8)
	) name1138 (
		\in0[33] ,
		_w1038_,
		_w1045_,
		_w1652_
	);
	LUT3 #(
		.INIT('hb0)
	) name1139 (
		_w1029_,
		_w1043_,
		_w1652_,
		_w1653_
	);
	LUT4 #(
		.INIT('haa20)
	) name1140 (
		\in1[33] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1654_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		_w1653_,
		_w1654_,
		_w1655_
	);
	LUT3 #(
		.INIT('ha8)
	) name1142 (
		\in2[33] ,
		_w521_,
		_w778_,
		_w1656_
	);
	LUT4 #(
		.INIT('h1500)
	) name1143 (
		_w526_,
		_w771_,
		_w776_,
		_w1656_,
		_w1657_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1144 (
		\in3[33] ,
		_w782_,
		_w1655_,
		_w1657_,
		_w1658_
	);
	LUT3 #(
		.INIT('ha8)
	) name1145 (
		\in0[35] ,
		_w1038_,
		_w1045_,
		_w1659_
	);
	LUT3 #(
		.INIT('hb0)
	) name1146 (
		_w1029_,
		_w1043_,
		_w1659_,
		_w1660_
	);
	LUT4 #(
		.INIT('haa20)
	) name1147 (
		\in1[35] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1661_
	);
	LUT2 #(
		.INIT('h1)
	) name1148 (
		_w1660_,
		_w1661_,
		_w1662_
	);
	LUT3 #(
		.INIT('ha8)
	) name1149 (
		\in2[35] ,
		_w521_,
		_w778_,
		_w1663_
	);
	LUT4 #(
		.INIT('h1500)
	) name1150 (
		_w526_,
		_w771_,
		_w776_,
		_w1663_,
		_w1664_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1151 (
		\in3[35] ,
		_w782_,
		_w1662_,
		_w1664_,
		_w1665_
	);
	LUT3 #(
		.INIT('h80)
	) name1152 (
		_w1651_,
		_w1658_,
		_w1665_,
		_w1666_
	);
	LUT3 #(
		.INIT('ha8)
	) name1153 (
		\in0[32] ,
		_w1038_,
		_w1045_,
		_w1667_
	);
	LUT3 #(
		.INIT('hb0)
	) name1154 (
		_w1029_,
		_w1043_,
		_w1667_,
		_w1668_
	);
	LUT4 #(
		.INIT('haa20)
	) name1155 (
		\in1[32] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1669_
	);
	LUT2 #(
		.INIT('h1)
	) name1156 (
		_w1668_,
		_w1669_,
		_w1670_
	);
	LUT3 #(
		.INIT('h02)
	) name1157 (
		\in3[32] ,
		_w1668_,
		_w1669_,
		_w1671_
	);
	LUT3 #(
		.INIT('h02)
	) name1158 (
		\in2[32] ,
		_w1668_,
		_w1669_,
		_w1672_
	);
	LUT3 #(
		.INIT('h1b)
	) name1159 (
		_w782_,
		_w1671_,
		_w1672_,
		_w1673_
	);
	LUT3 #(
		.INIT('ha8)
	) name1160 (
		\in0[31] ,
		_w1038_,
		_w1045_,
		_w1674_
	);
	LUT3 #(
		.INIT('hb0)
	) name1161 (
		_w1029_,
		_w1043_,
		_w1674_,
		_w1675_
	);
	LUT4 #(
		.INIT('haa20)
	) name1162 (
		\in1[31] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1676_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		_w1675_,
		_w1676_,
		_w1677_
	);
	LUT3 #(
		.INIT('ha8)
	) name1164 (
		\in2[31] ,
		_w521_,
		_w778_,
		_w1678_
	);
	LUT4 #(
		.INIT('h1500)
	) name1165 (
		_w526_,
		_w771_,
		_w776_,
		_w1678_,
		_w1679_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1166 (
		\in3[31] ,
		_w782_,
		_w1677_,
		_w1679_,
		_w1680_
	);
	LUT3 #(
		.INIT('ha8)
	) name1167 (
		\in0[36] ,
		_w1038_,
		_w1045_,
		_w1681_
	);
	LUT3 #(
		.INIT('hb0)
	) name1168 (
		_w1029_,
		_w1043_,
		_w1681_,
		_w1682_
	);
	LUT4 #(
		.INIT('haa20)
	) name1169 (
		\in1[36] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name1170 (
		_w1682_,
		_w1683_,
		_w1684_
	);
	LUT3 #(
		.INIT('ha8)
	) name1171 (
		\in2[36] ,
		_w521_,
		_w778_,
		_w1685_
	);
	LUT4 #(
		.INIT('h1500)
	) name1172 (
		_w526_,
		_w771_,
		_w776_,
		_w1685_,
		_w1686_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1173 (
		\in3[36] ,
		_w782_,
		_w1684_,
		_w1686_,
		_w1687_
	);
	LUT3 #(
		.INIT('h80)
	) name1174 (
		_w1673_,
		_w1680_,
		_w1687_,
		_w1688_
	);
	LUT3 #(
		.INIT('ha8)
	) name1175 (
		\in0[38] ,
		_w1038_,
		_w1045_,
		_w1689_
	);
	LUT3 #(
		.INIT('hb0)
	) name1176 (
		_w1029_,
		_w1043_,
		_w1689_,
		_w1690_
	);
	LUT4 #(
		.INIT('haa20)
	) name1177 (
		\in1[38] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1691_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		_w1690_,
		_w1691_,
		_w1692_
	);
	LUT3 #(
		.INIT('h02)
	) name1179 (
		\in3[38] ,
		_w1690_,
		_w1691_,
		_w1693_
	);
	LUT3 #(
		.INIT('h02)
	) name1180 (
		\in2[38] ,
		_w1690_,
		_w1691_,
		_w1694_
	);
	LUT3 #(
		.INIT('h1b)
	) name1181 (
		_w782_,
		_w1693_,
		_w1694_,
		_w1695_
	);
	LUT3 #(
		.INIT('ha8)
	) name1182 (
		\in0[39] ,
		_w1038_,
		_w1045_,
		_w1696_
	);
	LUT3 #(
		.INIT('hb0)
	) name1183 (
		_w1029_,
		_w1043_,
		_w1696_,
		_w1697_
	);
	LUT4 #(
		.INIT('haa20)
	) name1184 (
		\in1[39] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1698_
	);
	LUT2 #(
		.INIT('h1)
	) name1185 (
		_w1697_,
		_w1698_,
		_w1699_
	);
	LUT3 #(
		.INIT('ha8)
	) name1186 (
		\in2[39] ,
		_w521_,
		_w778_,
		_w1700_
	);
	LUT4 #(
		.INIT('h1500)
	) name1187 (
		_w526_,
		_w771_,
		_w776_,
		_w1700_,
		_w1701_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1188 (
		\in3[39] ,
		_w782_,
		_w1699_,
		_w1701_,
		_w1702_
	);
	LUT3 #(
		.INIT('ha8)
	) name1189 (
		\in0[37] ,
		_w1038_,
		_w1045_,
		_w1703_
	);
	LUT3 #(
		.INIT('hb0)
	) name1190 (
		_w1029_,
		_w1043_,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('haa20)
	) name1191 (
		\in1[37] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1705_
	);
	LUT2 #(
		.INIT('h1)
	) name1192 (
		_w1704_,
		_w1705_,
		_w1706_
	);
	LUT3 #(
		.INIT('ha8)
	) name1193 (
		\in2[37] ,
		_w521_,
		_w778_,
		_w1707_
	);
	LUT4 #(
		.INIT('h1500)
	) name1194 (
		_w526_,
		_w771_,
		_w776_,
		_w1707_,
		_w1708_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1195 (
		\in3[37] ,
		_w782_,
		_w1706_,
		_w1708_,
		_w1709_
	);
	LUT3 #(
		.INIT('h80)
	) name1196 (
		_w1695_,
		_w1702_,
		_w1709_,
		_w1710_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1197 (
		\in3[29] ,
		_w782_,
		_w1640_,
		_w1642_,
		_w1711_
	);
	LUT3 #(
		.INIT('ha8)
	) name1198 (
		\in0[30] ,
		_w1038_,
		_w1045_,
		_w1712_
	);
	LUT3 #(
		.INIT('hb0)
	) name1199 (
		_w1029_,
		_w1043_,
		_w1712_,
		_w1713_
	);
	LUT4 #(
		.INIT('haa20)
	) name1200 (
		\in1[30] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1714_
	);
	LUT2 #(
		.INIT('h1)
	) name1201 (
		_w1713_,
		_w1714_,
		_w1715_
	);
	LUT3 #(
		.INIT('ha8)
	) name1202 (
		\in2[30] ,
		_w521_,
		_w778_,
		_w1716_
	);
	LUT4 #(
		.INIT('h1500)
	) name1203 (
		_w526_,
		_w771_,
		_w776_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1204 (
		\in3[30] ,
		_w782_,
		_w1715_,
		_w1717_,
		_w1718_
	);
	LUT2 #(
		.INIT('h8)
	) name1205 (
		_w1711_,
		_w1718_,
		_w1719_
	);
	LUT4 #(
		.INIT('h8000)
	) name1206 (
		_w1666_,
		_w1688_,
		_w1710_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h4)
	) name1207 (
		_w1644_,
		_w1720_,
		_w1721_
	);
	LUT3 #(
		.INIT('ha8)
	) name1208 (
		\in0[21] ,
		_w1038_,
		_w1045_,
		_w1722_
	);
	LUT3 #(
		.INIT('hb0)
	) name1209 (
		_w1029_,
		_w1043_,
		_w1722_,
		_w1723_
	);
	LUT4 #(
		.INIT('haa20)
	) name1210 (
		\in1[21] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1724_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w1723_,
		_w1724_,
		_w1725_
	);
	LUT3 #(
		.INIT('ha8)
	) name1212 (
		\in2[21] ,
		_w521_,
		_w778_,
		_w1726_
	);
	LUT4 #(
		.INIT('h1500)
	) name1213 (
		_w526_,
		_w771_,
		_w776_,
		_w1726_,
		_w1727_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1214 (
		\in3[21] ,
		_w782_,
		_w1725_,
		_w1727_,
		_w1728_
	);
	LUT3 #(
		.INIT('ha8)
	) name1215 (
		\in0[20] ,
		_w1038_,
		_w1045_,
		_w1729_
	);
	LUT3 #(
		.INIT('hb0)
	) name1216 (
		_w1029_,
		_w1043_,
		_w1729_,
		_w1730_
	);
	LUT4 #(
		.INIT('haa20)
	) name1217 (
		\in1[20] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1731_
	);
	LUT2 #(
		.INIT('h1)
	) name1218 (
		_w1730_,
		_w1731_,
		_w1732_
	);
	LUT3 #(
		.INIT('ha8)
	) name1219 (
		\in2[20] ,
		_w521_,
		_w778_,
		_w1733_
	);
	LUT4 #(
		.INIT('h1500)
	) name1220 (
		_w526_,
		_w771_,
		_w776_,
		_w1733_,
		_w1734_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1221 (
		\in3[20] ,
		_w782_,
		_w1732_,
		_w1734_,
		_w1735_
	);
	LUT4 #(
		.INIT('h000d)
	) name1222 (
		\in3[20] ,
		_w782_,
		_w1732_,
		_w1734_,
		_w1736_
	);
	LUT3 #(
		.INIT('ha8)
	) name1223 (
		\in2[19] ,
		_w521_,
		_w778_,
		_w1737_
	);
	LUT4 #(
		.INIT('h1500)
	) name1224 (
		_w526_,
		_w771_,
		_w776_,
		_w1737_,
		_w1738_
	);
	LUT3 #(
		.INIT('ha8)
	) name1225 (
		\in0[19] ,
		_w1038_,
		_w1045_,
		_w1739_
	);
	LUT3 #(
		.INIT('hb0)
	) name1226 (
		_w1029_,
		_w1043_,
		_w1739_,
		_w1740_
	);
	LUT4 #(
		.INIT('haa20)
	) name1227 (
		\in1[19] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1741_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w1740_,
		_w1741_,
		_w1742_
	);
	LUT4 #(
		.INIT('h000d)
	) name1229 (
		\in3[19] ,
		_w782_,
		_w1738_,
		_w1742_,
		_w1743_
	);
	LUT4 #(
		.INIT('h8880)
	) name1230 (
		_w1728_,
		_w1735_,
		_w1736_,
		_w1743_,
		_w1744_
	);
	LUT3 #(
		.INIT('ha8)
	) name1231 (
		\in0[23] ,
		_w1038_,
		_w1045_,
		_w1745_
	);
	LUT3 #(
		.INIT('hb0)
	) name1232 (
		_w1029_,
		_w1043_,
		_w1745_,
		_w1746_
	);
	LUT4 #(
		.INIT('haa20)
	) name1233 (
		\in1[23] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1747_
	);
	LUT2 #(
		.INIT('h1)
	) name1234 (
		_w1746_,
		_w1747_,
		_w1748_
	);
	LUT3 #(
		.INIT('ha8)
	) name1235 (
		\in2[23] ,
		_w521_,
		_w778_,
		_w1749_
	);
	LUT4 #(
		.INIT('h1500)
	) name1236 (
		_w526_,
		_w771_,
		_w776_,
		_w1749_,
		_w1750_
	);
	LUT4 #(
		.INIT('h000d)
	) name1237 (
		\in3[23] ,
		_w782_,
		_w1748_,
		_w1750_,
		_w1751_
	);
	LUT3 #(
		.INIT('ha8)
	) name1238 (
		\in0[24] ,
		_w1038_,
		_w1045_,
		_w1752_
	);
	LUT3 #(
		.INIT('hb0)
	) name1239 (
		_w1029_,
		_w1043_,
		_w1752_,
		_w1753_
	);
	LUT4 #(
		.INIT('haa20)
	) name1240 (
		\in1[24] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1754_
	);
	LUT2 #(
		.INIT('h1)
	) name1241 (
		_w1753_,
		_w1754_,
		_w1755_
	);
	LUT3 #(
		.INIT('ha8)
	) name1242 (
		\in2[24] ,
		_w521_,
		_w778_,
		_w1756_
	);
	LUT4 #(
		.INIT('h1500)
	) name1243 (
		_w526_,
		_w771_,
		_w776_,
		_w1756_,
		_w1757_
	);
	LUT4 #(
		.INIT('h000d)
	) name1244 (
		\in3[24] ,
		_w782_,
		_w1755_,
		_w1757_,
		_w1758_
	);
	LUT3 #(
		.INIT('ha8)
	) name1245 (
		\in0[22] ,
		_w1038_,
		_w1045_,
		_w1759_
	);
	LUT3 #(
		.INIT('hb0)
	) name1246 (
		_w1029_,
		_w1043_,
		_w1759_,
		_w1760_
	);
	LUT4 #(
		.INIT('haa20)
	) name1247 (
		\in1[22] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1761_
	);
	LUT2 #(
		.INIT('h1)
	) name1248 (
		_w1760_,
		_w1761_,
		_w1762_
	);
	LUT3 #(
		.INIT('ha8)
	) name1249 (
		\in2[22] ,
		_w521_,
		_w778_,
		_w1763_
	);
	LUT4 #(
		.INIT('h1500)
	) name1250 (
		_w526_,
		_w771_,
		_w776_,
		_w1763_,
		_w1764_
	);
	LUT4 #(
		.INIT('h000d)
	) name1251 (
		\in3[22] ,
		_w782_,
		_w1762_,
		_w1764_,
		_w1765_
	);
	LUT4 #(
		.INIT('h000d)
	) name1252 (
		\in3[21] ,
		_w782_,
		_w1725_,
		_w1727_,
		_w1766_
	);
	LUT4 #(
		.INIT('h0001)
	) name1253 (
		_w1751_,
		_w1758_,
		_w1765_,
		_w1766_,
		_w1767_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1254 (
		\in3[22] ,
		_w782_,
		_w1762_,
		_w1764_,
		_w1768_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1255 (
		\in3[23] ,
		_w782_,
		_w1748_,
		_w1750_,
		_w1769_
	);
	LUT4 #(
		.INIT('h0111)
	) name1256 (
		_w1751_,
		_w1758_,
		_w1768_,
		_w1769_,
		_w1770_
	);
	LUT3 #(
		.INIT('ha8)
	) name1257 (
		\in0[25] ,
		_w1038_,
		_w1045_,
		_w1771_
	);
	LUT3 #(
		.INIT('hb0)
	) name1258 (
		_w1029_,
		_w1043_,
		_w1771_,
		_w1772_
	);
	LUT4 #(
		.INIT('haa20)
	) name1259 (
		\in1[25] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name1260 (
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT3 #(
		.INIT('ha8)
	) name1261 (
		\in2[25] ,
		_w521_,
		_w778_,
		_w1775_
	);
	LUT4 #(
		.INIT('h1500)
	) name1262 (
		_w526_,
		_w771_,
		_w776_,
		_w1775_,
		_w1776_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1263 (
		\in3[25] ,
		_w782_,
		_w1774_,
		_w1776_,
		_w1777_
	);
	LUT3 #(
		.INIT('ha8)
	) name1264 (
		\in0[26] ,
		_w1038_,
		_w1045_,
		_w1778_
	);
	LUT3 #(
		.INIT('hb0)
	) name1265 (
		_w1029_,
		_w1043_,
		_w1778_,
		_w1779_
	);
	LUT4 #(
		.INIT('haa20)
	) name1266 (
		\in1[26] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1780_
	);
	LUT2 #(
		.INIT('h1)
	) name1267 (
		_w1779_,
		_w1780_,
		_w1781_
	);
	LUT3 #(
		.INIT('ha8)
	) name1268 (
		\in2[26] ,
		_w521_,
		_w778_,
		_w1782_
	);
	LUT4 #(
		.INIT('h1500)
	) name1269 (
		_w526_,
		_w771_,
		_w776_,
		_w1782_,
		_w1783_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1270 (
		\in3[26] ,
		_w782_,
		_w1781_,
		_w1783_,
		_w1784_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1271 (
		\in3[24] ,
		_w782_,
		_w1755_,
		_w1757_,
		_w1785_
	);
	LUT3 #(
		.INIT('h80)
	) name1272 (
		_w1777_,
		_w1784_,
		_w1785_,
		_w1786_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1273 (
		_w1744_,
		_w1767_,
		_w1770_,
		_w1786_,
		_w1787_
	);
	LUT3 #(
		.INIT('ha8)
	) name1274 (
		\in0[12] ,
		_w1038_,
		_w1045_,
		_w1788_
	);
	LUT3 #(
		.INIT('hb0)
	) name1275 (
		_w1029_,
		_w1043_,
		_w1788_,
		_w1789_
	);
	LUT4 #(
		.INIT('haa20)
	) name1276 (
		\in1[12] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1790_
	);
	LUT2 #(
		.INIT('h1)
	) name1277 (
		_w1789_,
		_w1790_,
		_w1791_
	);
	LUT3 #(
		.INIT('ha8)
	) name1278 (
		\in2[12] ,
		_w521_,
		_w778_,
		_w1792_
	);
	LUT4 #(
		.INIT('h1500)
	) name1279 (
		_w526_,
		_w771_,
		_w776_,
		_w1792_,
		_w1793_
	);
	LUT4 #(
		.INIT('h000d)
	) name1280 (
		\in3[12] ,
		_w782_,
		_w1791_,
		_w1793_,
		_w1794_
	);
	LUT3 #(
		.INIT('ha8)
	) name1281 (
		\in0[11] ,
		_w1038_,
		_w1045_,
		_w1795_
	);
	LUT3 #(
		.INIT('hb0)
	) name1282 (
		_w1029_,
		_w1043_,
		_w1795_,
		_w1796_
	);
	LUT4 #(
		.INIT('haa20)
	) name1283 (
		\in1[11] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1797_
	);
	LUT2 #(
		.INIT('h1)
	) name1284 (
		_w1796_,
		_w1797_,
		_w1798_
	);
	LUT3 #(
		.INIT('ha8)
	) name1285 (
		\in2[11] ,
		_w521_,
		_w778_,
		_w1799_
	);
	LUT4 #(
		.INIT('h1500)
	) name1286 (
		_w526_,
		_w771_,
		_w776_,
		_w1799_,
		_w1800_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1287 (
		\in3[11] ,
		_w782_,
		_w1798_,
		_w1800_,
		_w1801_
	);
	LUT2 #(
		.INIT('h1)
	) name1288 (
		_w1794_,
		_w1801_,
		_w1802_
	);
	LUT3 #(
		.INIT('ha8)
	) name1289 (
		\in0[14] ,
		_w1038_,
		_w1045_,
		_w1803_
	);
	LUT3 #(
		.INIT('hb0)
	) name1290 (
		_w1029_,
		_w1043_,
		_w1803_,
		_w1804_
	);
	LUT4 #(
		.INIT('haa20)
	) name1291 (
		\in1[14] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name1292 (
		_w1804_,
		_w1805_,
		_w1806_
	);
	LUT3 #(
		.INIT('ha8)
	) name1293 (
		\in2[14] ,
		_w521_,
		_w778_,
		_w1807_
	);
	LUT4 #(
		.INIT('h1500)
	) name1294 (
		_w526_,
		_w771_,
		_w776_,
		_w1807_,
		_w1808_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1295 (
		\in3[14] ,
		_w782_,
		_w1806_,
		_w1808_,
		_w1809_
	);
	LUT3 #(
		.INIT('ha8)
	) name1296 (
		\in0[15] ,
		_w1038_,
		_w1045_,
		_w1810_
	);
	LUT3 #(
		.INIT('hb0)
	) name1297 (
		_w1029_,
		_w1043_,
		_w1810_,
		_w1811_
	);
	LUT4 #(
		.INIT('haa20)
	) name1298 (
		\in1[15] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1812_
	);
	LUT2 #(
		.INIT('h1)
	) name1299 (
		_w1811_,
		_w1812_,
		_w1813_
	);
	LUT3 #(
		.INIT('ha8)
	) name1300 (
		\in2[15] ,
		_w521_,
		_w778_,
		_w1814_
	);
	LUT4 #(
		.INIT('h1500)
	) name1301 (
		_w526_,
		_w771_,
		_w776_,
		_w1814_,
		_w1815_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1302 (
		\in3[15] ,
		_w782_,
		_w1813_,
		_w1815_,
		_w1816_
	);
	LUT3 #(
		.INIT('ha8)
	) name1303 (
		\in0[13] ,
		_w1038_,
		_w1045_,
		_w1817_
	);
	LUT3 #(
		.INIT('hb0)
	) name1304 (
		_w1029_,
		_w1043_,
		_w1817_,
		_w1818_
	);
	LUT4 #(
		.INIT('haa20)
	) name1305 (
		\in1[13] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1819_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		_w1818_,
		_w1819_,
		_w1820_
	);
	LUT3 #(
		.INIT('ha8)
	) name1307 (
		\in2[13] ,
		_w521_,
		_w778_,
		_w1821_
	);
	LUT4 #(
		.INIT('h1500)
	) name1308 (
		_w526_,
		_w771_,
		_w776_,
		_w1821_,
		_w1822_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1309 (
		\in3[13] ,
		_w782_,
		_w1820_,
		_w1822_,
		_w1823_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1310 (
		\in3[12] ,
		_w782_,
		_w1791_,
		_w1793_,
		_w1824_
	);
	LUT4 #(
		.INIT('h8000)
	) name1311 (
		_w1809_,
		_w1816_,
		_w1823_,
		_w1824_,
		_w1825_
	);
	LUT4 #(
		.INIT('h000d)
	) name1312 (
		\in3[13] ,
		_w782_,
		_w1820_,
		_w1822_,
		_w1826_
	);
	LUT4 #(
		.INIT('h000d)
	) name1313 (
		\in3[14] ,
		_w782_,
		_w1806_,
		_w1808_,
		_w1827_
	);
	LUT4 #(
		.INIT('h8880)
	) name1314 (
		_w1809_,
		_w1816_,
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT3 #(
		.INIT('ha8)
	) name1315 (
		\in0[17] ,
		_w1038_,
		_w1045_,
		_w1829_
	);
	LUT3 #(
		.INIT('hb0)
	) name1316 (
		_w1029_,
		_w1043_,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('haa20)
	) name1317 (
		\in1[17] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1831_
	);
	LUT2 #(
		.INIT('h1)
	) name1318 (
		_w1830_,
		_w1831_,
		_w1832_
	);
	LUT3 #(
		.INIT('ha8)
	) name1319 (
		\in2[17] ,
		_w521_,
		_w778_,
		_w1833_
	);
	LUT4 #(
		.INIT('h1500)
	) name1320 (
		_w526_,
		_w771_,
		_w776_,
		_w1833_,
		_w1834_
	);
	LUT4 #(
		.INIT('h000d)
	) name1321 (
		\in3[17] ,
		_w782_,
		_w1832_,
		_w1834_,
		_w1835_
	);
	LUT3 #(
		.INIT('ha8)
	) name1322 (
		\in0[18] ,
		_w1038_,
		_w1045_,
		_w1836_
	);
	LUT3 #(
		.INIT('hb0)
	) name1323 (
		_w1029_,
		_w1043_,
		_w1836_,
		_w1837_
	);
	LUT4 #(
		.INIT('haa20)
	) name1324 (
		\in1[18] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1838_
	);
	LUT2 #(
		.INIT('h1)
	) name1325 (
		_w1837_,
		_w1838_,
		_w1839_
	);
	LUT3 #(
		.INIT('ha8)
	) name1326 (
		\in2[18] ,
		_w521_,
		_w778_,
		_w1840_
	);
	LUT4 #(
		.INIT('h1500)
	) name1327 (
		_w526_,
		_w771_,
		_w776_,
		_w1840_,
		_w1841_
	);
	LUT4 #(
		.INIT('h000d)
	) name1328 (
		\in3[18] ,
		_w782_,
		_w1839_,
		_w1841_,
		_w1842_
	);
	LUT3 #(
		.INIT('ha8)
	) name1329 (
		\in0[16] ,
		_w1038_,
		_w1045_,
		_w1843_
	);
	LUT3 #(
		.INIT('hb0)
	) name1330 (
		_w1029_,
		_w1043_,
		_w1843_,
		_w1844_
	);
	LUT4 #(
		.INIT('haa20)
	) name1331 (
		\in1[16] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1845_
	);
	LUT2 #(
		.INIT('h1)
	) name1332 (
		_w1844_,
		_w1845_,
		_w1846_
	);
	LUT3 #(
		.INIT('ha8)
	) name1333 (
		\in2[16] ,
		_w521_,
		_w778_,
		_w1847_
	);
	LUT4 #(
		.INIT('h1500)
	) name1334 (
		_w526_,
		_w771_,
		_w776_,
		_w1847_,
		_w1848_
	);
	LUT4 #(
		.INIT('h000d)
	) name1335 (
		\in3[16] ,
		_w782_,
		_w1846_,
		_w1848_,
		_w1849_
	);
	LUT4 #(
		.INIT('h000d)
	) name1336 (
		\in3[15] ,
		_w782_,
		_w1813_,
		_w1815_,
		_w1850_
	);
	LUT4 #(
		.INIT('h0001)
	) name1337 (
		_w1835_,
		_w1842_,
		_w1849_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1338 (
		_w1802_,
		_w1825_,
		_w1828_,
		_w1851_,
		_w1852_
	);
	LUT3 #(
		.INIT('ha8)
	) name1339 (
		\in0[4] ,
		_w1038_,
		_w1045_,
		_w1853_
	);
	LUT3 #(
		.INIT('hb0)
	) name1340 (
		_w1029_,
		_w1043_,
		_w1853_,
		_w1854_
	);
	LUT4 #(
		.INIT('haa20)
	) name1341 (
		\in1[4] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name1342 (
		_w1854_,
		_w1855_,
		_w1856_
	);
	LUT3 #(
		.INIT('ha8)
	) name1343 (
		\in2[4] ,
		_w521_,
		_w778_,
		_w1857_
	);
	LUT4 #(
		.INIT('h1500)
	) name1344 (
		_w526_,
		_w771_,
		_w776_,
		_w1857_,
		_w1858_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1345 (
		\in3[4] ,
		_w782_,
		_w1856_,
		_w1858_,
		_w1859_
	);
	LUT3 #(
		.INIT('ha8)
	) name1346 (
		\in0[5] ,
		_w1038_,
		_w1045_,
		_w1860_
	);
	LUT3 #(
		.INIT('hb0)
	) name1347 (
		_w1029_,
		_w1043_,
		_w1860_,
		_w1861_
	);
	LUT4 #(
		.INIT('haa20)
	) name1348 (
		\in1[5] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name1349 (
		_w1861_,
		_w1862_,
		_w1863_
	);
	LUT3 #(
		.INIT('h02)
	) name1350 (
		\in3[5] ,
		_w1861_,
		_w1862_,
		_w1864_
	);
	LUT3 #(
		.INIT('h02)
	) name1351 (
		\in2[5] ,
		_w1861_,
		_w1862_,
		_w1865_
	);
	LUT3 #(
		.INIT('h1b)
	) name1352 (
		_w782_,
		_w1864_,
		_w1865_,
		_w1866_
	);
	LUT3 #(
		.INIT('ha8)
	) name1353 (
		\in0[3] ,
		_w1038_,
		_w1045_,
		_w1867_
	);
	LUT3 #(
		.INIT('hb0)
	) name1354 (
		_w1029_,
		_w1043_,
		_w1867_,
		_w1868_
	);
	LUT4 #(
		.INIT('haa20)
	) name1355 (
		\in1[3] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1869_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT3 #(
		.INIT('ha8)
	) name1357 (
		\in2[3] ,
		_w521_,
		_w778_,
		_w1871_
	);
	LUT4 #(
		.INIT('h1500)
	) name1358 (
		_w526_,
		_w771_,
		_w776_,
		_w1871_,
		_w1872_
	);
	LUT4 #(
		.INIT('h000d)
	) name1359 (
		\in3[3] ,
		_w782_,
		_w1870_,
		_w1872_,
		_w1873_
	);
	LUT4 #(
		.INIT('h000d)
	) name1360 (
		\in3[4] ,
		_w782_,
		_w1856_,
		_w1858_,
		_w1874_
	);
	LUT4 #(
		.INIT('h8880)
	) name1361 (
		_w1859_,
		_w1866_,
		_w1873_,
		_w1874_,
		_w1875_
	);
	LUT3 #(
		.INIT('ha8)
	) name1362 (
		\in0[1] ,
		_w1038_,
		_w1045_,
		_w1876_
	);
	LUT3 #(
		.INIT('hb0)
	) name1363 (
		_w1029_,
		_w1043_,
		_w1876_,
		_w1877_
	);
	LUT4 #(
		.INIT('haa20)
	) name1364 (
		\in1[1] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1878_
	);
	LUT2 #(
		.INIT('h1)
	) name1365 (
		_w1877_,
		_w1878_,
		_w1879_
	);
	LUT3 #(
		.INIT('h02)
	) name1366 (
		\in3[1] ,
		_w1877_,
		_w1878_,
		_w1880_
	);
	LUT3 #(
		.INIT('h02)
	) name1367 (
		\in2[1] ,
		_w1877_,
		_w1878_,
		_w1881_
	);
	LUT3 #(
		.INIT('h1b)
	) name1368 (
		_w782_,
		_w1880_,
		_w1881_,
		_w1882_
	);
	LUT3 #(
		.INIT('ha8)
	) name1369 (
		\in0[0] ,
		_w1038_,
		_w1045_,
		_w1883_
	);
	LUT3 #(
		.INIT('hb0)
	) name1370 (
		_w1029_,
		_w1043_,
		_w1883_,
		_w1884_
	);
	LUT4 #(
		.INIT('haa20)
	) name1371 (
		\in1[0] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1885_
	);
	LUT2 #(
		.INIT('h1)
	) name1372 (
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT4 #(
		.INIT('h0031)
	) name1373 (
		\in3[0] ,
		_w781_,
		_w782_,
		_w1886_,
		_w1887_
	);
	LUT3 #(
		.INIT('ha8)
	) name1374 (
		\in2[1] ,
		_w521_,
		_w778_,
		_w1888_
	);
	LUT4 #(
		.INIT('h1500)
	) name1375 (
		_w526_,
		_w771_,
		_w776_,
		_w1888_,
		_w1889_
	);
	LUT4 #(
		.INIT('h000d)
	) name1376 (
		\in3[1] ,
		_w782_,
		_w1879_,
		_w1889_,
		_w1890_
	);
	LUT3 #(
		.INIT('ha8)
	) name1377 (
		\in0[2] ,
		_w1038_,
		_w1045_,
		_w1891_
	);
	LUT3 #(
		.INIT('hb0)
	) name1378 (
		_w1029_,
		_w1043_,
		_w1891_,
		_w1892_
	);
	LUT4 #(
		.INIT('haa20)
	) name1379 (
		\in1[2] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1893_
	);
	LUT2 #(
		.INIT('h1)
	) name1380 (
		_w1892_,
		_w1893_,
		_w1894_
	);
	LUT3 #(
		.INIT('ha8)
	) name1381 (
		\in2[2] ,
		_w521_,
		_w778_,
		_w1895_
	);
	LUT4 #(
		.INIT('h1500)
	) name1382 (
		_w526_,
		_w771_,
		_w776_,
		_w1895_,
		_w1896_
	);
	LUT4 #(
		.INIT('h000d)
	) name1383 (
		\in3[2] ,
		_w782_,
		_w1894_,
		_w1896_,
		_w1897_
	);
	LUT4 #(
		.INIT('h0007)
	) name1384 (
		_w1882_,
		_w1887_,
		_w1890_,
		_w1897_,
		_w1898_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1385 (
		\in3[3] ,
		_w782_,
		_w1870_,
		_w1872_,
		_w1899_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1386 (
		\in3[2] ,
		_w782_,
		_w1894_,
		_w1896_,
		_w1900_
	);
	LUT4 #(
		.INIT('h8000)
	) name1387 (
		_w1859_,
		_w1866_,
		_w1899_,
		_w1900_,
		_w1901_
	);
	LUT3 #(
		.INIT('ha8)
	) name1388 (
		\in0[7] ,
		_w1038_,
		_w1045_,
		_w1902_
	);
	LUT3 #(
		.INIT('hb0)
	) name1389 (
		_w1029_,
		_w1043_,
		_w1902_,
		_w1903_
	);
	LUT4 #(
		.INIT('haa20)
	) name1390 (
		\in1[7] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1904_
	);
	LUT2 #(
		.INIT('h1)
	) name1391 (
		_w1903_,
		_w1904_,
		_w1905_
	);
	LUT3 #(
		.INIT('ha8)
	) name1392 (
		\in2[7] ,
		_w521_,
		_w778_,
		_w1906_
	);
	LUT4 #(
		.INIT('h1500)
	) name1393 (
		_w526_,
		_w771_,
		_w776_,
		_w1906_,
		_w1907_
	);
	LUT4 #(
		.INIT('h000d)
	) name1394 (
		\in3[7] ,
		_w782_,
		_w1905_,
		_w1907_,
		_w1908_
	);
	LUT3 #(
		.INIT('ha8)
	) name1395 (
		\in0[6] ,
		_w1038_,
		_w1045_,
		_w1909_
	);
	LUT3 #(
		.INIT('hb0)
	) name1396 (
		_w1029_,
		_w1043_,
		_w1909_,
		_w1910_
	);
	LUT4 #(
		.INIT('haa20)
	) name1397 (
		\in1[6] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1911_
	);
	LUT2 #(
		.INIT('h1)
	) name1398 (
		_w1910_,
		_w1911_,
		_w1912_
	);
	LUT3 #(
		.INIT('ha8)
	) name1399 (
		\in2[6] ,
		_w521_,
		_w778_,
		_w1913_
	);
	LUT4 #(
		.INIT('h1500)
	) name1400 (
		_w526_,
		_w771_,
		_w776_,
		_w1913_,
		_w1914_
	);
	LUT4 #(
		.INIT('h000d)
	) name1401 (
		\in3[6] ,
		_w782_,
		_w1912_,
		_w1914_,
		_w1915_
	);
	LUT3 #(
		.INIT('ha8)
	) name1402 (
		\in2[5] ,
		_w521_,
		_w778_,
		_w1916_
	);
	LUT4 #(
		.INIT('h1500)
	) name1403 (
		_w526_,
		_w771_,
		_w776_,
		_w1916_,
		_w1917_
	);
	LUT4 #(
		.INIT('h000d)
	) name1404 (
		\in3[5] ,
		_w782_,
		_w1863_,
		_w1917_,
		_w1918_
	);
	LUT3 #(
		.INIT('h01)
	) name1405 (
		_w1908_,
		_w1915_,
		_w1918_,
		_w1919_
	);
	LUT4 #(
		.INIT('h4500)
	) name1406 (
		_w1875_,
		_w1898_,
		_w1901_,
		_w1919_,
		_w1920_
	);
	LUT3 #(
		.INIT('h0d)
	) name1407 (
		\in3[6] ,
		_w782_,
		_w1914_,
		_w1921_
	);
	LUT3 #(
		.INIT('h04)
	) name1408 (
		_w1908_,
		_w1912_,
		_w1921_,
		_w1922_
	);
	LUT3 #(
		.INIT('ha8)
	) name1409 (
		\in0[10] ,
		_w1038_,
		_w1045_,
		_w1923_
	);
	LUT3 #(
		.INIT('hb0)
	) name1410 (
		_w1029_,
		_w1043_,
		_w1923_,
		_w1924_
	);
	LUT4 #(
		.INIT('haa20)
	) name1411 (
		\in1[10] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1925_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		_w1924_,
		_w1925_,
		_w1926_
	);
	LUT3 #(
		.INIT('ha8)
	) name1413 (
		\in2[10] ,
		_w521_,
		_w778_,
		_w1927_
	);
	LUT4 #(
		.INIT('h1500)
	) name1414 (
		_w526_,
		_w771_,
		_w776_,
		_w1927_,
		_w1928_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1415 (
		\in3[10] ,
		_w782_,
		_w1926_,
		_w1928_,
		_w1929_
	);
	LUT3 #(
		.INIT('ha8)
	) name1416 (
		\in0[9] ,
		_w1038_,
		_w1045_,
		_w1930_
	);
	LUT3 #(
		.INIT('hb0)
	) name1417 (
		_w1029_,
		_w1043_,
		_w1930_,
		_w1931_
	);
	LUT4 #(
		.INIT('haa20)
	) name1418 (
		\in1[9] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1932_
	);
	LUT2 #(
		.INIT('h1)
	) name1419 (
		_w1931_,
		_w1932_,
		_w1933_
	);
	LUT3 #(
		.INIT('ha8)
	) name1420 (
		\in2[9] ,
		_w521_,
		_w778_,
		_w1934_
	);
	LUT4 #(
		.INIT('h1500)
	) name1421 (
		_w526_,
		_w771_,
		_w776_,
		_w1934_,
		_w1935_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1422 (
		\in3[9] ,
		_w782_,
		_w1933_,
		_w1935_,
		_w1936_
	);
	LUT3 #(
		.INIT('ha8)
	) name1423 (
		\in0[8] ,
		_w1038_,
		_w1045_,
		_w1937_
	);
	LUT3 #(
		.INIT('hb0)
	) name1424 (
		_w1029_,
		_w1043_,
		_w1937_,
		_w1938_
	);
	LUT4 #(
		.INIT('haa20)
	) name1425 (
		\in1[8] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1939_
	);
	LUT2 #(
		.INIT('h1)
	) name1426 (
		_w1938_,
		_w1939_,
		_w1940_
	);
	LUT3 #(
		.INIT('ha8)
	) name1427 (
		\in2[8] ,
		_w521_,
		_w778_,
		_w1941_
	);
	LUT4 #(
		.INIT('h1500)
	) name1428 (
		_w526_,
		_w771_,
		_w776_,
		_w1941_,
		_w1942_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1429 (
		\in3[8] ,
		_w782_,
		_w1940_,
		_w1942_,
		_w1943_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1430 (
		\in3[7] ,
		_w782_,
		_w1905_,
		_w1907_,
		_w1944_
	);
	LUT4 #(
		.INIT('h8000)
	) name1431 (
		_w1929_,
		_w1936_,
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h4)
	) name1432 (
		_w1922_,
		_w1945_,
		_w1946_
	);
	LUT4 #(
		.INIT('h000d)
	) name1433 (
		\in3[8] ,
		_w782_,
		_w1940_,
		_w1942_,
		_w1947_
	);
	LUT4 #(
		.INIT('h000d)
	) name1434 (
		\in3[9] ,
		_w782_,
		_w1933_,
		_w1935_,
		_w1948_
	);
	LUT4 #(
		.INIT('h8880)
	) name1435 (
		_w1929_,
		_w1936_,
		_w1947_,
		_w1948_,
		_w1949_
	);
	LUT4 #(
		.INIT('h000d)
	) name1436 (
		\in3[11] ,
		_w782_,
		_w1798_,
		_w1800_,
		_w1950_
	);
	LUT4 #(
		.INIT('h000d)
	) name1437 (
		\in3[10] ,
		_w782_,
		_w1926_,
		_w1928_,
		_w1951_
	);
	LUT3 #(
		.INIT('h01)
	) name1438 (
		_w1794_,
		_w1950_,
		_w1951_,
		_w1952_
	);
	LUT4 #(
		.INIT('h0400)
	) name1439 (
		_w1828_,
		_w1851_,
		_w1949_,
		_w1952_,
		_w1953_
	);
	LUT4 #(
		.INIT('h1055)
	) name1440 (
		_w1852_,
		_w1920_,
		_w1946_,
		_w1953_,
		_w1954_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1441 (
		\in3[16] ,
		_w782_,
		_w1846_,
		_w1848_,
		_w1955_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1442 (
		\in3[17] ,
		_w782_,
		_w1832_,
		_w1834_,
		_w1956_
	);
	LUT4 #(
		.INIT('h0111)
	) name1443 (
		_w1835_,
		_w1842_,
		_w1955_,
		_w1956_,
		_w1957_
	);
	LUT3 #(
		.INIT('h02)
	) name1444 (
		\in3[19] ,
		_w1740_,
		_w1741_,
		_w1958_
	);
	LUT3 #(
		.INIT('h02)
	) name1445 (
		\in2[19] ,
		_w1740_,
		_w1741_,
		_w1959_
	);
	LUT3 #(
		.INIT('h1b)
	) name1446 (
		_w782_,
		_w1958_,
		_w1959_,
		_w1960_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1447 (
		\in3[18] ,
		_w782_,
		_w1839_,
		_w1841_,
		_w1961_
	);
	LUT4 #(
		.INIT('h8000)
	) name1448 (
		_w1728_,
		_w1735_,
		_w1960_,
		_w1961_,
		_w1962_
	);
	LUT4 #(
		.INIT('h0400)
	) name1449 (
		_w1770_,
		_w1786_,
		_w1957_,
		_w1962_,
		_w1963_
	);
	LUT4 #(
		.INIT('h000d)
	) name1450 (
		\in3[25] ,
		_w782_,
		_w1774_,
		_w1776_,
		_w1964_
	);
	LUT4 #(
		.INIT('h000d)
	) name1451 (
		\in3[26] ,
		_w782_,
		_w1781_,
		_w1783_,
		_w1965_
	);
	LUT3 #(
		.INIT('ha8)
	) name1452 (
		\in0[27] ,
		_w1038_,
		_w1045_,
		_w1966_
	);
	LUT3 #(
		.INIT('hb0)
	) name1453 (
		_w1029_,
		_w1043_,
		_w1966_,
		_w1967_
	);
	LUT4 #(
		.INIT('haa20)
	) name1454 (
		\in1[27] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w1968_
	);
	LUT2 #(
		.INIT('h1)
	) name1455 (
		_w1967_,
		_w1968_,
		_w1969_
	);
	LUT3 #(
		.INIT('ha8)
	) name1456 (
		\in2[27] ,
		_w521_,
		_w778_,
		_w1970_
	);
	LUT4 #(
		.INIT('h1500)
	) name1457 (
		_w526_,
		_w771_,
		_w776_,
		_w1970_,
		_w1971_
	);
	LUT4 #(
		.INIT('h000d)
	) name1458 (
		\in3[27] ,
		_w782_,
		_w1969_,
		_w1971_,
		_w1972_
	);
	LUT4 #(
		.INIT('h0057)
	) name1459 (
		_w1784_,
		_w1964_,
		_w1965_,
		_w1972_,
		_w1973_
	);
	LUT4 #(
		.INIT('h1500)
	) name1460 (
		_w1787_,
		_w1954_,
		_w1963_,
		_w1973_,
		_w1974_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1461 (
		\in3[27] ,
		_w782_,
		_w1969_,
		_w1971_,
		_w1975_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1462 (
		\in3[28] ,
		_w782_,
		_w1633_,
		_w1635_,
		_w1976_
	);
	LUT2 #(
		.INIT('h8)
	) name1463 (
		_w1975_,
		_w1976_,
		_w1977_
	);
	LUT2 #(
		.INIT('h8)
	) name1464 (
		_w1720_,
		_w1977_,
		_w1978_
	);
	LUT3 #(
		.INIT('ha8)
	) name1465 (
		\in2[38] ,
		_w521_,
		_w778_,
		_w1979_
	);
	LUT4 #(
		.INIT('h1500)
	) name1466 (
		_w526_,
		_w771_,
		_w776_,
		_w1979_,
		_w1980_
	);
	LUT4 #(
		.INIT('h000d)
	) name1467 (
		\in3[38] ,
		_w782_,
		_w1692_,
		_w1980_,
		_w1981_
	);
	LUT4 #(
		.INIT('h000d)
	) name1468 (
		\in3[39] ,
		_w782_,
		_w1699_,
		_w1701_,
		_w1982_
	);
	LUT3 #(
		.INIT('h07)
	) name1469 (
		_w1702_,
		_w1981_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h4)
	) name1470 (
		_w1710_,
		_w1983_,
		_w1984_
	);
	LUT3 #(
		.INIT('ha8)
	) name1471 (
		\in2[34] ,
		_w521_,
		_w778_,
		_w1985_
	);
	LUT4 #(
		.INIT('h1500)
	) name1472 (
		_w526_,
		_w771_,
		_w776_,
		_w1985_,
		_w1986_
	);
	LUT4 #(
		.INIT('h000d)
	) name1473 (
		\in3[34] ,
		_w782_,
		_w1648_,
		_w1986_,
		_w1987_
	);
	LUT4 #(
		.INIT('h000d)
	) name1474 (
		\in3[35] ,
		_w782_,
		_w1662_,
		_w1664_,
		_w1988_
	);
	LUT4 #(
		.INIT('hcc80)
	) name1475 (
		_w1665_,
		_w1687_,
		_w1987_,
		_w1988_,
		_w1989_
	);
	LUT3 #(
		.INIT('ha8)
	) name1476 (
		\in2[32] ,
		_w521_,
		_w778_,
		_w1990_
	);
	LUT4 #(
		.INIT('h1500)
	) name1477 (
		_w526_,
		_w771_,
		_w776_,
		_w1990_,
		_w1991_
	);
	LUT4 #(
		.INIT('h000d)
	) name1478 (
		\in3[32] ,
		_w782_,
		_w1670_,
		_w1991_,
		_w1992_
	);
	LUT4 #(
		.INIT('h000d)
	) name1479 (
		\in3[33] ,
		_w782_,
		_w1655_,
		_w1657_,
		_w1993_
	);
	LUT2 #(
		.INIT('h1)
	) name1480 (
		_w1992_,
		_w1993_,
		_w1994_
	);
	LUT4 #(
		.INIT('h8000)
	) name1481 (
		_w1651_,
		_w1658_,
		_w1665_,
		_w1687_,
		_w1995_
	);
	LUT3 #(
		.INIT('h45)
	) name1482 (
		_w1989_,
		_w1994_,
		_w1995_,
		_w1996_
	);
	LUT4 #(
		.INIT('h000d)
	) name1483 (
		\in3[36] ,
		_w782_,
		_w1684_,
		_w1686_,
		_w1997_
	);
	LUT4 #(
		.INIT('h000d)
	) name1484 (
		\in3[37] ,
		_w782_,
		_w1706_,
		_w1708_,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name1485 (
		_w1997_,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('h8)
	) name1486 (
		_w1983_,
		_w1999_,
		_w2000_
	);
	LUT3 #(
		.INIT('h15)
	) name1487 (
		_w1984_,
		_w1996_,
		_w2000_,
		_w2001_
	);
	LUT3 #(
		.INIT('ha8)
	) name1488 (
		\in0[46] ,
		_w1038_,
		_w1045_,
		_w2002_
	);
	LUT3 #(
		.INIT('hb0)
	) name1489 (
		_w1029_,
		_w1043_,
		_w2002_,
		_w2003_
	);
	LUT4 #(
		.INIT('haa20)
	) name1490 (
		\in1[46] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2004_
	);
	LUT2 #(
		.INIT('h1)
	) name1491 (
		_w2003_,
		_w2004_,
		_w2005_
	);
	LUT3 #(
		.INIT('h02)
	) name1492 (
		\in3[46] ,
		_w2003_,
		_w2004_,
		_w2006_
	);
	LUT3 #(
		.INIT('h02)
	) name1493 (
		\in2[46] ,
		_w2003_,
		_w2004_,
		_w2007_
	);
	LUT3 #(
		.INIT('h1b)
	) name1494 (
		_w782_,
		_w2006_,
		_w2007_,
		_w2008_
	);
	LUT3 #(
		.INIT('ha8)
	) name1495 (
		\in0[47] ,
		_w1038_,
		_w1045_,
		_w2009_
	);
	LUT3 #(
		.INIT('hb0)
	) name1496 (
		_w1029_,
		_w1043_,
		_w2009_,
		_w2010_
	);
	LUT4 #(
		.INIT('haa20)
	) name1497 (
		\in1[47] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2011_
	);
	LUT2 #(
		.INIT('h1)
	) name1498 (
		_w2010_,
		_w2011_,
		_w2012_
	);
	LUT3 #(
		.INIT('ha8)
	) name1499 (
		\in2[47] ,
		_w521_,
		_w778_,
		_w2013_
	);
	LUT4 #(
		.INIT('h1500)
	) name1500 (
		_w526_,
		_w771_,
		_w776_,
		_w2013_,
		_w2014_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1501 (
		\in3[47] ,
		_w782_,
		_w2012_,
		_w2014_,
		_w2015_
	);
	LUT3 #(
		.INIT('ha8)
	) name1502 (
		\in0[45] ,
		_w1038_,
		_w1045_,
		_w2016_
	);
	LUT3 #(
		.INIT('hb0)
	) name1503 (
		_w1029_,
		_w1043_,
		_w2016_,
		_w2017_
	);
	LUT4 #(
		.INIT('haa20)
	) name1504 (
		\in1[45] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2018_
	);
	LUT2 #(
		.INIT('h1)
	) name1505 (
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT3 #(
		.INIT('ha8)
	) name1506 (
		\in2[45] ,
		_w521_,
		_w778_,
		_w2020_
	);
	LUT4 #(
		.INIT('h1500)
	) name1507 (
		_w526_,
		_w771_,
		_w776_,
		_w2020_,
		_w2021_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1508 (
		\in3[45] ,
		_w782_,
		_w2019_,
		_w2021_,
		_w2022_
	);
	LUT3 #(
		.INIT('h80)
	) name1509 (
		_w2008_,
		_w2015_,
		_w2022_,
		_w2023_
	);
	LUT3 #(
		.INIT('ha8)
	) name1510 (
		\in0[44] ,
		_w1038_,
		_w1045_,
		_w2024_
	);
	LUT3 #(
		.INIT('hb0)
	) name1511 (
		_w1029_,
		_w1043_,
		_w2024_,
		_w2025_
	);
	LUT4 #(
		.INIT('haa20)
	) name1512 (
		\in1[44] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2026_
	);
	LUT2 #(
		.INIT('h1)
	) name1513 (
		_w2025_,
		_w2026_,
		_w2027_
	);
	LUT3 #(
		.INIT('ha8)
	) name1514 (
		\in2[44] ,
		_w521_,
		_w778_,
		_w2028_
	);
	LUT4 #(
		.INIT('h1500)
	) name1515 (
		_w526_,
		_w771_,
		_w776_,
		_w2028_,
		_w2029_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1516 (
		\in3[44] ,
		_w782_,
		_w2027_,
		_w2029_,
		_w2030_
	);
	LUT3 #(
		.INIT('ha8)
	) name1517 (
		\in0[43] ,
		_w1038_,
		_w1045_,
		_w2031_
	);
	LUT3 #(
		.INIT('hb0)
	) name1518 (
		_w1029_,
		_w1043_,
		_w2031_,
		_w2032_
	);
	LUT4 #(
		.INIT('haa20)
	) name1519 (
		\in1[43] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2033_
	);
	LUT2 #(
		.INIT('h1)
	) name1520 (
		_w2032_,
		_w2033_,
		_w2034_
	);
	LUT3 #(
		.INIT('h02)
	) name1521 (
		\in3[43] ,
		_w2032_,
		_w2033_,
		_w2035_
	);
	LUT3 #(
		.INIT('h02)
	) name1522 (
		\in2[43] ,
		_w2032_,
		_w2033_,
		_w2036_
	);
	LUT3 #(
		.INIT('h1b)
	) name1523 (
		_w782_,
		_w2035_,
		_w2036_,
		_w2037_
	);
	LUT3 #(
		.INIT('ha8)
	) name1524 (
		\in0[42] ,
		_w1038_,
		_w1045_,
		_w2038_
	);
	LUT3 #(
		.INIT('hb0)
	) name1525 (
		_w1029_,
		_w1043_,
		_w2038_,
		_w2039_
	);
	LUT4 #(
		.INIT('haa20)
	) name1526 (
		\in1[42] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2040_
	);
	LUT2 #(
		.INIT('h1)
	) name1527 (
		_w2039_,
		_w2040_,
		_w2041_
	);
	LUT3 #(
		.INIT('ha8)
	) name1528 (
		\in2[42] ,
		_w521_,
		_w778_,
		_w2042_
	);
	LUT4 #(
		.INIT('h1500)
	) name1529 (
		_w526_,
		_w771_,
		_w776_,
		_w2042_,
		_w2043_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1530 (
		\in3[42] ,
		_w782_,
		_w2041_,
		_w2043_,
		_w2044_
	);
	LUT3 #(
		.INIT('h80)
	) name1531 (
		_w2030_,
		_w2037_,
		_w2044_,
		_w2045_
	);
	LUT3 #(
		.INIT('ha8)
	) name1532 (
		\in0[41] ,
		_w1038_,
		_w1045_,
		_w2046_
	);
	LUT3 #(
		.INIT('hb0)
	) name1533 (
		_w1029_,
		_w1043_,
		_w2046_,
		_w2047_
	);
	LUT4 #(
		.INIT('haa20)
	) name1534 (
		\in1[41] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2048_
	);
	LUT2 #(
		.INIT('h1)
	) name1535 (
		_w2047_,
		_w2048_,
		_w2049_
	);
	LUT3 #(
		.INIT('ha8)
	) name1536 (
		\in2[41] ,
		_w521_,
		_w778_,
		_w2050_
	);
	LUT4 #(
		.INIT('h1500)
	) name1537 (
		_w526_,
		_w771_,
		_w776_,
		_w2050_,
		_w2051_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1538 (
		\in3[41] ,
		_w782_,
		_w2049_,
		_w2051_,
		_w2052_
	);
	LUT3 #(
		.INIT('ha8)
	) name1539 (
		\in2[40] ,
		_w521_,
		_w778_,
		_w2053_
	);
	LUT4 #(
		.INIT('h1500)
	) name1540 (
		_w526_,
		_w771_,
		_w776_,
		_w2053_,
		_w2054_
	);
	LUT3 #(
		.INIT('ha8)
	) name1541 (
		\in0[40] ,
		_w1038_,
		_w1045_,
		_w2055_
	);
	LUT3 #(
		.INIT('hb0)
	) name1542 (
		_w1029_,
		_w1043_,
		_w2055_,
		_w2056_
	);
	LUT4 #(
		.INIT('haa20)
	) name1543 (
		\in1[40] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name1544 (
		_w2056_,
		_w2057_,
		_w2058_
	);
	LUT4 #(
		.INIT('h000d)
	) name1545 (
		\in3[40] ,
		_w782_,
		_w2054_,
		_w2058_,
		_w2059_
	);
	LUT4 #(
		.INIT('h000d)
	) name1546 (
		\in3[42] ,
		_w782_,
		_w2041_,
		_w2043_,
		_w2060_
	);
	LUT4 #(
		.INIT('h000d)
	) name1547 (
		\in3[41] ,
		_w782_,
		_w2049_,
		_w2051_,
		_w2061_
	);
	LUT4 #(
		.INIT('h0007)
	) name1548 (
		_w2052_,
		_w2059_,
		_w2060_,
		_w2061_,
		_w2062_
	);
	LUT3 #(
		.INIT('ha8)
	) name1549 (
		\in2[43] ,
		_w521_,
		_w778_,
		_w2063_
	);
	LUT4 #(
		.INIT('h1500)
	) name1550 (
		_w526_,
		_w771_,
		_w776_,
		_w2063_,
		_w2064_
	);
	LUT4 #(
		.INIT('h000d)
	) name1551 (
		\in3[43] ,
		_w782_,
		_w2034_,
		_w2064_,
		_w2065_
	);
	LUT4 #(
		.INIT('h000d)
	) name1552 (
		\in3[44] ,
		_w782_,
		_w2027_,
		_w2029_,
		_w2066_
	);
	LUT4 #(
		.INIT('h000d)
	) name1553 (
		\in3[45] ,
		_w782_,
		_w2019_,
		_w2021_,
		_w2067_
	);
	LUT4 #(
		.INIT('h0007)
	) name1554 (
		_w2030_,
		_w2065_,
		_w2066_,
		_w2067_,
		_w2068_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1555 (
		_w2023_,
		_w2045_,
		_w2062_,
		_w2068_,
		_w2069_
	);
	LUT4 #(
		.INIT('h000d)
	) name1556 (
		\in3[30] ,
		_w782_,
		_w1715_,
		_w1717_,
		_w2070_
	);
	LUT4 #(
		.INIT('h000d)
	) name1557 (
		\in3[31] ,
		_w782_,
		_w1677_,
		_w1679_,
		_w2071_
	);
	LUT2 #(
		.INIT('h1)
	) name1558 (
		_w2070_,
		_w2071_,
		_w2072_
	);
	LUT4 #(
		.INIT('h0080)
	) name1559 (
		_w1666_,
		_w1688_,
		_w1710_,
		_w2072_,
		_w2073_
	);
	LUT3 #(
		.INIT('ha8)
	) name1560 (
		\in2[46] ,
		_w521_,
		_w778_,
		_w2074_
	);
	LUT4 #(
		.INIT('h1500)
	) name1561 (
		_w526_,
		_w771_,
		_w776_,
		_w2074_,
		_w2075_
	);
	LUT4 #(
		.INIT('h000d)
	) name1562 (
		\in3[46] ,
		_w782_,
		_w2005_,
		_w2075_,
		_w2076_
	);
	LUT4 #(
		.INIT('h000d)
	) name1563 (
		\in3[47] ,
		_w782_,
		_w2012_,
		_w2014_,
		_w2077_
	);
	LUT3 #(
		.INIT('h07)
	) name1564 (
		_w2015_,
		_w2076_,
		_w2077_,
		_w2078_
	);
	LUT3 #(
		.INIT('h10)
	) name1565 (
		_w2069_,
		_w2073_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h4)
	) name1566 (
		_w2001_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('h4500)
	) name1567 (
		_w1721_,
		_w1974_,
		_w1978_,
		_w2080_,
		_w2081_
	);
	LUT3 #(
		.INIT('h02)
	) name1568 (
		\in3[40] ,
		_w2056_,
		_w2057_,
		_w2082_
	);
	LUT3 #(
		.INIT('h02)
	) name1569 (
		\in2[40] ,
		_w2056_,
		_w2057_,
		_w2083_
	);
	LUT3 #(
		.INIT('h1b)
	) name1570 (
		_w782_,
		_w2082_,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h8)
	) name1571 (
		_w2052_,
		_w2084_,
		_w2085_
	);
	LUT4 #(
		.INIT('h70f0)
	) name1572 (
		_w2023_,
		_w2045_,
		_w2078_,
		_w2085_,
		_w2086_
	);
	LUT3 #(
		.INIT('ha8)
	) name1573 (
		\in0[55] ,
		_w1038_,
		_w1045_,
		_w2087_
	);
	LUT3 #(
		.INIT('hb0)
	) name1574 (
		_w1029_,
		_w1043_,
		_w2087_,
		_w2088_
	);
	LUT4 #(
		.INIT('haa20)
	) name1575 (
		\in1[55] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2089_
	);
	LUT2 #(
		.INIT('h1)
	) name1576 (
		_w2088_,
		_w2089_,
		_w2090_
	);
	LUT3 #(
		.INIT('ha8)
	) name1577 (
		\in2[55] ,
		_w521_,
		_w778_,
		_w2091_
	);
	LUT4 #(
		.INIT('h1500)
	) name1578 (
		_w526_,
		_w771_,
		_w776_,
		_w2091_,
		_w2092_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1579 (
		\in3[55] ,
		_w782_,
		_w2090_,
		_w2092_,
		_w2093_
	);
	LUT3 #(
		.INIT('ha8)
	) name1580 (
		\in0[54] ,
		_w1038_,
		_w1045_,
		_w2094_
	);
	LUT3 #(
		.INIT('hb0)
	) name1581 (
		_w1029_,
		_w1043_,
		_w2094_,
		_w2095_
	);
	LUT4 #(
		.INIT('haa20)
	) name1582 (
		\in1[54] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2096_
	);
	LUT2 #(
		.INIT('h1)
	) name1583 (
		_w2095_,
		_w2096_,
		_w2097_
	);
	LUT3 #(
		.INIT('h02)
	) name1584 (
		\in3[54] ,
		_w2095_,
		_w2096_,
		_w2098_
	);
	LUT3 #(
		.INIT('h02)
	) name1585 (
		\in2[54] ,
		_w2095_,
		_w2096_,
		_w2099_
	);
	LUT3 #(
		.INIT('h1b)
	) name1586 (
		_w782_,
		_w2098_,
		_w2099_,
		_w2100_
	);
	LUT2 #(
		.INIT('h8)
	) name1587 (
		_w2093_,
		_w2100_,
		_w2101_
	);
	LUT3 #(
		.INIT('ha8)
	) name1588 (
		\in0[52] ,
		_w1038_,
		_w1045_,
		_w2102_
	);
	LUT3 #(
		.INIT('hb0)
	) name1589 (
		_w1029_,
		_w1043_,
		_w2102_,
		_w2103_
	);
	LUT4 #(
		.INIT('haa20)
	) name1590 (
		\in1[52] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2104_
	);
	LUT2 #(
		.INIT('h1)
	) name1591 (
		_w2103_,
		_w2104_,
		_w2105_
	);
	LUT3 #(
		.INIT('h02)
	) name1592 (
		\in3[52] ,
		_w2103_,
		_w2104_,
		_w2106_
	);
	LUT3 #(
		.INIT('h02)
	) name1593 (
		\in2[52] ,
		_w2103_,
		_w2104_,
		_w2107_
	);
	LUT3 #(
		.INIT('h1b)
	) name1594 (
		_w782_,
		_w2106_,
		_w2107_,
		_w2108_
	);
	LUT3 #(
		.INIT('ha8)
	) name1595 (
		\in0[53] ,
		_w1038_,
		_w1045_,
		_w2109_
	);
	LUT3 #(
		.INIT('hb0)
	) name1596 (
		_w1029_,
		_w1043_,
		_w2109_,
		_w2110_
	);
	LUT4 #(
		.INIT('haa20)
	) name1597 (
		\in1[53] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2111_
	);
	LUT2 #(
		.INIT('h1)
	) name1598 (
		_w2110_,
		_w2111_,
		_w2112_
	);
	LUT3 #(
		.INIT('ha8)
	) name1599 (
		\in2[53] ,
		_w521_,
		_w778_,
		_w2113_
	);
	LUT4 #(
		.INIT('h1500)
	) name1600 (
		_w526_,
		_w771_,
		_w776_,
		_w2113_,
		_w2114_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1601 (
		\in3[53] ,
		_w782_,
		_w2112_,
		_w2114_,
		_w2115_
	);
	LUT4 #(
		.INIT('h8000)
	) name1602 (
		_w2093_,
		_w2100_,
		_w2108_,
		_w2115_,
		_w2116_
	);
	LUT3 #(
		.INIT('ha8)
	) name1603 (
		\in0[51] ,
		_w1038_,
		_w1045_,
		_w2117_
	);
	LUT3 #(
		.INIT('hb0)
	) name1604 (
		_w1029_,
		_w1043_,
		_w2117_,
		_w2118_
	);
	LUT4 #(
		.INIT('haa20)
	) name1605 (
		\in1[51] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2119_
	);
	LUT2 #(
		.INIT('h1)
	) name1606 (
		_w2118_,
		_w2119_,
		_w2120_
	);
	LUT3 #(
		.INIT('ha8)
	) name1607 (
		\in2[51] ,
		_w521_,
		_w778_,
		_w2121_
	);
	LUT4 #(
		.INIT('h1500)
	) name1608 (
		_w526_,
		_w771_,
		_w776_,
		_w2121_,
		_w2122_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1609 (
		\in3[51] ,
		_w782_,
		_w2120_,
		_w2122_,
		_w2123_
	);
	LUT3 #(
		.INIT('ha8)
	) name1610 (
		\in0[50] ,
		_w1038_,
		_w1045_,
		_w2124_
	);
	LUT3 #(
		.INIT('hb0)
	) name1611 (
		_w1029_,
		_w1043_,
		_w2124_,
		_w2125_
	);
	LUT4 #(
		.INIT('haa20)
	) name1612 (
		\in1[50] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2126_
	);
	LUT2 #(
		.INIT('h1)
	) name1613 (
		_w2125_,
		_w2126_,
		_w2127_
	);
	LUT3 #(
		.INIT('h02)
	) name1614 (
		\in3[50] ,
		_w2125_,
		_w2126_,
		_w2128_
	);
	LUT3 #(
		.INIT('h02)
	) name1615 (
		\in2[50] ,
		_w2125_,
		_w2126_,
		_w2129_
	);
	LUT3 #(
		.INIT('h1b)
	) name1616 (
		_w782_,
		_w2128_,
		_w2129_,
		_w2130_
	);
	LUT3 #(
		.INIT('ha8)
	) name1617 (
		\in0[49] ,
		_w1038_,
		_w1045_,
		_w2131_
	);
	LUT3 #(
		.INIT('hb0)
	) name1618 (
		_w1029_,
		_w1043_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('haa20)
	) name1619 (
		\in1[49] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name1620 (
		_w2132_,
		_w2133_,
		_w2134_
	);
	LUT3 #(
		.INIT('ha8)
	) name1621 (
		\in2[49] ,
		_w521_,
		_w778_,
		_w2135_
	);
	LUT4 #(
		.INIT('h1500)
	) name1622 (
		_w526_,
		_w771_,
		_w776_,
		_w2135_,
		_w2136_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1623 (
		\in3[49] ,
		_w782_,
		_w2134_,
		_w2136_,
		_w2137_
	);
	LUT3 #(
		.INIT('ha8)
	) name1624 (
		\in0[48] ,
		_w1038_,
		_w1045_,
		_w2138_
	);
	LUT3 #(
		.INIT('hb0)
	) name1625 (
		_w1029_,
		_w1043_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('haa20)
	) name1626 (
		\in1[48] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2140_
	);
	LUT2 #(
		.INIT('h1)
	) name1627 (
		_w2139_,
		_w2140_,
		_w2141_
	);
	LUT3 #(
		.INIT('h02)
	) name1628 (
		\in3[48] ,
		_w2139_,
		_w2140_,
		_w2142_
	);
	LUT3 #(
		.INIT('h02)
	) name1629 (
		\in2[48] ,
		_w2139_,
		_w2140_,
		_w2143_
	);
	LUT3 #(
		.INIT('h1b)
	) name1630 (
		_w782_,
		_w2142_,
		_w2143_,
		_w2144_
	);
	LUT4 #(
		.INIT('h8000)
	) name1631 (
		_w2123_,
		_w2130_,
		_w2137_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h8)
	) name1632 (
		_w2116_,
		_w2145_,
		_w2146_
	);
	LUT3 #(
		.INIT('hb0)
	) name1633 (
		_w2069_,
		_w2086_,
		_w2146_,
		_w2147_
	);
	LUT3 #(
		.INIT('h80)
	) name1634 (
		_w2123_,
		_w2130_,
		_w2137_,
		_w2148_
	);
	LUT3 #(
		.INIT('ha8)
	) name1635 (
		\in2[48] ,
		_w521_,
		_w778_,
		_w2149_
	);
	LUT4 #(
		.INIT('h1500)
	) name1636 (
		_w526_,
		_w771_,
		_w776_,
		_w2149_,
		_w2150_
	);
	LUT4 #(
		.INIT('h000d)
	) name1637 (
		\in3[48] ,
		_w782_,
		_w2141_,
		_w2150_,
		_w2151_
	);
	LUT4 #(
		.INIT('h000d)
	) name1638 (
		\in3[49] ,
		_w782_,
		_w2134_,
		_w2136_,
		_w2152_
	);
	LUT2 #(
		.INIT('h1)
	) name1639 (
		_w2151_,
		_w2152_,
		_w2153_
	);
	LUT4 #(
		.INIT('h000d)
	) name1640 (
		\in3[51] ,
		_w782_,
		_w2120_,
		_w2122_,
		_w2154_
	);
	LUT3 #(
		.INIT('ha8)
	) name1641 (
		\in2[50] ,
		_w521_,
		_w778_,
		_w2155_
	);
	LUT4 #(
		.INIT('h1500)
	) name1642 (
		_w526_,
		_w771_,
		_w776_,
		_w2155_,
		_w2156_
	);
	LUT4 #(
		.INIT('h000d)
	) name1643 (
		\in3[50] ,
		_w782_,
		_w2127_,
		_w2156_,
		_w2157_
	);
	LUT3 #(
		.INIT('h13)
	) name1644 (
		_w2123_,
		_w2154_,
		_w2157_,
		_w2158_
	);
	LUT4 #(
		.INIT('h08aa)
	) name1645 (
		_w2116_,
		_w2148_,
		_w2153_,
		_w2158_,
		_w2159_
	);
	LUT4 #(
		.INIT('h000d)
	) name1646 (
		\in3[55] ,
		_w782_,
		_w2090_,
		_w2092_,
		_w2160_
	);
	LUT3 #(
		.INIT('ha8)
	) name1647 (
		\in2[52] ,
		_w521_,
		_w778_,
		_w2161_
	);
	LUT4 #(
		.INIT('h1500)
	) name1648 (
		_w526_,
		_w771_,
		_w776_,
		_w2161_,
		_w2162_
	);
	LUT4 #(
		.INIT('h000d)
	) name1649 (
		\in3[52] ,
		_w782_,
		_w2105_,
		_w2162_,
		_w2163_
	);
	LUT4 #(
		.INIT('h000d)
	) name1650 (
		\in3[53] ,
		_w782_,
		_w2112_,
		_w2114_,
		_w2164_
	);
	LUT3 #(
		.INIT('ha8)
	) name1651 (
		\in2[54] ,
		_w521_,
		_w778_,
		_w2165_
	);
	LUT4 #(
		.INIT('h1500)
	) name1652 (
		_w526_,
		_w771_,
		_w776_,
		_w2165_,
		_w2166_
	);
	LUT4 #(
		.INIT('h000d)
	) name1653 (
		\in3[54] ,
		_w782_,
		_w2097_,
		_w2166_,
		_w2167_
	);
	LUT4 #(
		.INIT('h0007)
	) name1654 (
		_w2115_,
		_w2163_,
		_w2164_,
		_w2167_,
		_w2168_
	);
	LUT3 #(
		.INIT('h31)
	) name1655 (
		_w2101_,
		_w2160_,
		_w2168_,
		_w2169_
	);
	LUT4 #(
		.INIT('h0200)
	) name1656 (
		_w1618_,
		_w1628_,
		_w2159_,
		_w2169_,
		_w2170_
	);
	LUT4 #(
		.INIT('h1055)
	) name1657 (
		_w1629_,
		_w2081_,
		_w2147_,
		_w2170_,
		_w2171_
	);
	LUT3 #(
		.INIT('h02)
	) name1658 (
		\in3[64] ,
		_w1514_,
		_w1515_,
		_w2172_
	);
	LUT3 #(
		.INIT('h02)
	) name1659 (
		\in2[64] ,
		_w1514_,
		_w1515_,
		_w2173_
	);
	LUT3 #(
		.INIT('h1b)
	) name1660 (
		_w782_,
		_w2172_,
		_w2173_,
		_w2174_
	);
	LUT4 #(
		.INIT('h8000)
	) name1661 (
		_w1495_,
		_w1502_,
		_w1510_,
		_w2174_,
		_w2175_
	);
	LUT2 #(
		.INIT('h8)
	) name1662 (
		_w1552_,
		_w2175_,
		_w2176_
	);
	LUT4 #(
		.INIT('h000d)
	) name1663 (
		\in3[71] ,
		_w782_,
		_w1526_,
		_w1528_,
		_w2177_
	);
	LUT3 #(
		.INIT('ha8)
	) name1664 (
		\in2[68] ,
		_w521_,
		_w778_,
		_w2178_
	);
	LUT4 #(
		.INIT('h1500)
	) name1665 (
		_w526_,
		_w771_,
		_w776_,
		_w2178_,
		_w2179_
	);
	LUT4 #(
		.INIT('h000d)
	) name1666 (
		\in3[68] ,
		_w782_,
		_w1548_,
		_w2179_,
		_w2180_
	);
	LUT3 #(
		.INIT('ha8)
	) name1667 (
		\in2[70] ,
		_w521_,
		_w778_,
		_w2181_
	);
	LUT4 #(
		.INIT('h1500)
	) name1668 (
		_w526_,
		_w771_,
		_w776_,
		_w2181_,
		_w2182_
	);
	LUT4 #(
		.INIT('h000d)
	) name1669 (
		\in3[70] ,
		_w782_,
		_w1533_,
		_w2182_,
		_w2183_
	);
	LUT4 #(
		.INIT('h000d)
	) name1670 (
		\in3[69] ,
		_w782_,
		_w1541_,
		_w1543_,
		_w2184_
	);
	LUT4 #(
		.INIT('h0007)
	) name1671 (
		_w1544_,
		_w2180_,
		_w2183_,
		_w2184_,
		_w2185_
	);
	LUT3 #(
		.INIT('h31)
	) name1672 (
		_w1537_,
		_w2177_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h8)
	) name1673 (
		_w1486_,
		_w2186_,
		_w2187_
	);
	LUT4 #(
		.INIT('h1500)
	) name1674 (
		_w1553_,
		_w2171_,
		_w2176_,
		_w2187_,
		_w2188_
	);
	LUT3 #(
		.INIT('h02)
	) name1675 (
		\in3[76] ,
		_w1407_,
		_w1408_,
		_w2189_
	);
	LUT3 #(
		.INIT('h02)
	) name1676 (
		\in2[76] ,
		_w1407_,
		_w1408_,
		_w2190_
	);
	LUT3 #(
		.INIT('h1b)
	) name1677 (
		_w782_,
		_w2189_,
		_w2190_,
		_w2191_
	);
	LUT4 #(
		.INIT('h8000)
	) name1678 (
		_w1388_,
		_w1395_,
		_w1403_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h8)
	) name1679 (
		_w1445_,
		_w2192_,
		_w2193_
	);
	LUT4 #(
		.INIT('h5455)
	) name1680 (
		_w1446_,
		_w1487_,
		_w2188_,
		_w2193_,
		_w2194_
	);
	LUT4 #(
		.INIT('h000d)
	) name1681 (
		\in3[83] ,
		_w782_,
		_w1419_,
		_w1421_,
		_w2195_
	);
	LUT3 #(
		.INIT('ha8)
	) name1682 (
		\in2[80] ,
		_w521_,
		_w778_,
		_w2196_
	);
	LUT4 #(
		.INIT('h1500)
	) name1683 (
		_w526_,
		_w771_,
		_w776_,
		_w2196_,
		_w2197_
	);
	LUT4 #(
		.INIT('h000d)
	) name1684 (
		\in3[80] ,
		_w782_,
		_w1441_,
		_w2197_,
		_w2198_
	);
	LUT4 #(
		.INIT('h000d)
	) name1685 (
		\in3[81] ,
		_w782_,
		_w1434_,
		_w1436_,
		_w2199_
	);
	LUT3 #(
		.INIT('ha8)
	) name1686 (
		\in2[82] ,
		_w521_,
		_w778_,
		_w2200_
	);
	LUT4 #(
		.INIT('h1500)
	) name1687 (
		_w526_,
		_w771_,
		_w776_,
		_w2200_,
		_w2201_
	);
	LUT4 #(
		.INIT('h000d)
	) name1688 (
		\in3[82] ,
		_w782_,
		_w1426_,
		_w2201_,
		_w2202_
	);
	LUT4 #(
		.INIT('h0007)
	) name1689 (
		_w1437_,
		_w2198_,
		_w2199_,
		_w2202_,
		_w2203_
	);
	LUT3 #(
		.INIT('h31)
	) name1690 (
		_w1430_,
		_w2195_,
		_w2203_,
		_w2204_
	);
	LUT3 #(
		.INIT('h80)
	) name1691 (
		_w1369_,
		_w1379_,
		_w2204_,
		_w2205_
	);
	LUT3 #(
		.INIT('h02)
	) name1692 (
		\in3[88] ,
		_w1360_,
		_w1361_,
		_w2206_
	);
	LUT3 #(
		.INIT('h02)
	) name1693 (
		\in2[88] ,
		_w1360_,
		_w1361_,
		_w2207_
	);
	LUT3 #(
		.INIT('h1b)
	) name1694 (
		_w782_,
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h8)
	) name1695 (
		_w1356_,
		_w2208_,
		_w2209_
	);
	LUT4 #(
		.INIT('h1151)
	) name1696 (
		_w1340_,
		_w1349_,
		_w1368_,
		_w2209_,
		_w2210_
	);
	LUT3 #(
		.INIT('ha8)
	) name1697 (
		\in0[95] ,
		_w1038_,
		_w1045_,
		_w2211_
	);
	LUT3 #(
		.INIT('hb0)
	) name1698 (
		_w1029_,
		_w1043_,
		_w2211_,
		_w2212_
	);
	LUT4 #(
		.INIT('haa20)
	) name1699 (
		\in1[95] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2213_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		_w2212_,
		_w2213_,
		_w2214_
	);
	LUT3 #(
		.INIT('ha8)
	) name1701 (
		\in2[95] ,
		_w521_,
		_w778_,
		_w2215_
	);
	LUT4 #(
		.INIT('h1500)
	) name1702 (
		_w526_,
		_w771_,
		_w776_,
		_w2215_,
		_w2216_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1703 (
		\in3[95] ,
		_w782_,
		_w2214_,
		_w2216_,
		_w2217_
	);
	LUT3 #(
		.INIT('ha8)
	) name1704 (
		\in0[94] ,
		_w1038_,
		_w1045_,
		_w2218_
	);
	LUT3 #(
		.INIT('hb0)
	) name1705 (
		_w1029_,
		_w1043_,
		_w2218_,
		_w2219_
	);
	LUT4 #(
		.INIT('haa20)
	) name1706 (
		\in1[94] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2220_
	);
	LUT2 #(
		.INIT('h1)
	) name1707 (
		_w2219_,
		_w2220_,
		_w2221_
	);
	LUT3 #(
		.INIT('h02)
	) name1708 (
		\in3[94] ,
		_w2219_,
		_w2220_,
		_w2222_
	);
	LUT3 #(
		.INIT('h02)
	) name1709 (
		\in2[94] ,
		_w2219_,
		_w2220_,
		_w2223_
	);
	LUT3 #(
		.INIT('h1b)
	) name1710 (
		_w782_,
		_w2222_,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('h8)
	) name1711 (
		_w2217_,
		_w2224_,
		_w2225_
	);
	LUT3 #(
		.INIT('ha8)
	) name1712 (
		\in0[93] ,
		_w1038_,
		_w1045_,
		_w2226_
	);
	LUT3 #(
		.INIT('hb0)
	) name1713 (
		_w1029_,
		_w1043_,
		_w2226_,
		_w2227_
	);
	LUT4 #(
		.INIT('haa20)
	) name1714 (
		\in1[93] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2228_
	);
	LUT2 #(
		.INIT('h1)
	) name1715 (
		_w2227_,
		_w2228_,
		_w2229_
	);
	LUT3 #(
		.INIT('ha8)
	) name1716 (
		\in2[93] ,
		_w521_,
		_w778_,
		_w2230_
	);
	LUT4 #(
		.INIT('h1500)
	) name1717 (
		_w526_,
		_w771_,
		_w776_,
		_w2230_,
		_w2231_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1718 (
		\in3[93] ,
		_w782_,
		_w2229_,
		_w2231_,
		_w2232_
	);
	LUT3 #(
		.INIT('ha8)
	) name1719 (
		\in0[92] ,
		_w1038_,
		_w1045_,
		_w2233_
	);
	LUT3 #(
		.INIT('hb0)
	) name1720 (
		_w1029_,
		_w1043_,
		_w2233_,
		_w2234_
	);
	LUT4 #(
		.INIT('haa20)
	) name1721 (
		\in1[92] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2235_
	);
	LUT2 #(
		.INIT('h1)
	) name1722 (
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT3 #(
		.INIT('h02)
	) name1723 (
		\in3[92] ,
		_w2234_,
		_w2235_,
		_w2237_
	);
	LUT3 #(
		.INIT('h02)
	) name1724 (
		\in2[92] ,
		_w2234_,
		_w2235_,
		_w2238_
	);
	LUT3 #(
		.INIT('h1b)
	) name1725 (
		_w782_,
		_w2237_,
		_w2238_,
		_w2239_
	);
	LUT4 #(
		.INIT('h8000)
	) name1726 (
		_w2217_,
		_w2224_,
		_w2232_,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h4)
	) name1727 (
		_w2210_,
		_w2240_,
		_w2241_
	);
	LUT4 #(
		.INIT('h1500)
	) name1728 (
		_w1380_,
		_w2194_,
		_w2205_,
		_w2241_,
		_w2242_
	);
	LUT4 #(
		.INIT('h000d)
	) name1729 (
		\in3[95] ,
		_w782_,
		_w2214_,
		_w2216_,
		_w2243_
	);
	LUT3 #(
		.INIT('ha8)
	) name1730 (
		\in2[92] ,
		_w521_,
		_w778_,
		_w2244_
	);
	LUT4 #(
		.INIT('h1500)
	) name1731 (
		_w526_,
		_w771_,
		_w776_,
		_w2244_,
		_w2245_
	);
	LUT4 #(
		.INIT('h000d)
	) name1732 (
		\in3[92] ,
		_w782_,
		_w2236_,
		_w2245_,
		_w2246_
	);
	LUT3 #(
		.INIT('ha8)
	) name1733 (
		\in2[94] ,
		_w521_,
		_w778_,
		_w2247_
	);
	LUT4 #(
		.INIT('h1500)
	) name1734 (
		_w526_,
		_w771_,
		_w776_,
		_w2247_,
		_w2248_
	);
	LUT4 #(
		.INIT('h000d)
	) name1735 (
		\in3[94] ,
		_w782_,
		_w2221_,
		_w2248_,
		_w2249_
	);
	LUT4 #(
		.INIT('h000d)
	) name1736 (
		\in3[93] ,
		_w782_,
		_w2229_,
		_w2231_,
		_w2250_
	);
	LUT4 #(
		.INIT('h0007)
	) name1737 (
		_w2232_,
		_w2246_,
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT3 #(
		.INIT('h31)
	) name1738 (
		_w2225_,
		_w2243_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h8)
	) name1739 (
		_w1302_,
		_w2252_,
		_w2253_
	);
	LUT3 #(
		.INIT('h02)
	) name1740 (
		\in3[100] ,
		_w1223_,
		_w1224_,
		_w2254_
	);
	LUT3 #(
		.INIT('h02)
	) name1741 (
		\in2[100] ,
		_w1223_,
		_w1224_,
		_w2255_
	);
	LUT3 #(
		.INIT('h1b)
	) name1742 (
		_w782_,
		_w2254_,
		_w2255_,
		_w2256_
	);
	LUT4 #(
		.INIT('h8000)
	) name1743 (
		_w1204_,
		_w1211_,
		_w1219_,
		_w2256_,
		_w2257_
	);
	LUT2 #(
		.INIT('h8)
	) name1744 (
		_w1261_,
		_w2257_,
		_w2258_
	);
	LUT4 #(
		.INIT('h4500)
	) name1745 (
		_w1303_,
		_w2242_,
		_w2253_,
		_w2258_,
		_w2259_
	);
	LUT4 #(
		.INIT('h000d)
	) name1746 (
		\in3[107] ,
		_w782_,
		_w1235_,
		_w1237_,
		_w2260_
	);
	LUT3 #(
		.INIT('ha8)
	) name1747 (
		\in2[104] ,
		_w521_,
		_w778_,
		_w2261_
	);
	LUT4 #(
		.INIT('h1500)
	) name1748 (
		_w526_,
		_w771_,
		_w776_,
		_w2261_,
		_w2262_
	);
	LUT4 #(
		.INIT('h000d)
	) name1749 (
		\in3[104] ,
		_w782_,
		_w1257_,
		_w2262_,
		_w2263_
	);
	LUT4 #(
		.INIT('h000d)
	) name1750 (
		\in3[105] ,
		_w782_,
		_w1250_,
		_w1252_,
		_w2264_
	);
	LUT3 #(
		.INIT('ha8)
	) name1751 (
		\in2[106] ,
		_w521_,
		_w778_,
		_w2265_
	);
	LUT4 #(
		.INIT('h1500)
	) name1752 (
		_w526_,
		_w771_,
		_w776_,
		_w2265_,
		_w2266_
	);
	LUT4 #(
		.INIT('h000d)
	) name1753 (
		\in3[106] ,
		_w782_,
		_w1242_,
		_w2266_,
		_w2267_
	);
	LUT4 #(
		.INIT('h0007)
	) name1754 (
		_w1253_,
		_w2263_,
		_w2264_,
		_w2267_,
		_w2268_
	);
	LUT3 #(
		.INIT('h31)
	) name1755 (
		_w1246_,
		_w2260_,
		_w2268_,
		_w2269_
	);
	LUT3 #(
		.INIT('h80)
	) name1756 (
		_w1185_,
		_w1195_,
		_w2269_,
		_w2270_
	);
	LUT4 #(
		.INIT('h5455)
	) name1757 (
		_w1196_,
		_w1262_,
		_w2259_,
		_w2270_,
		_w2271_
	);
	LUT3 #(
		.INIT('h02)
	) name1758 (
		\in3[112] ,
		_w1176_,
		_w1177_,
		_w2272_
	);
	LUT3 #(
		.INIT('h02)
	) name1759 (
		\in2[112] ,
		_w1176_,
		_w1177_,
		_w2273_
	);
	LUT3 #(
		.INIT('h1b)
	) name1760 (
		_w782_,
		_w2272_,
		_w2273_,
		_w2274_
	);
	LUT2 #(
		.INIT('h8)
	) name1761 (
		_w1172_,
		_w2274_,
		_w2275_
	);
	LUT4 #(
		.INIT('h1151)
	) name1762 (
		_w1156_,
		_w1165_,
		_w1184_,
		_w2275_,
		_w2276_
	);
	LUT3 #(
		.INIT('ha8)
	) name1763 (
		\in0[119] ,
		_w1038_,
		_w1045_,
		_w2277_
	);
	LUT3 #(
		.INIT('hb0)
	) name1764 (
		_w1029_,
		_w1043_,
		_w2277_,
		_w2278_
	);
	LUT4 #(
		.INIT('haa20)
	) name1765 (
		\in1[119] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2279_
	);
	LUT2 #(
		.INIT('h1)
	) name1766 (
		_w2278_,
		_w2279_,
		_w2280_
	);
	LUT3 #(
		.INIT('ha8)
	) name1767 (
		\in2[119] ,
		_w521_,
		_w778_,
		_w2281_
	);
	LUT4 #(
		.INIT('h1500)
	) name1768 (
		_w526_,
		_w771_,
		_w776_,
		_w2281_,
		_w2282_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1769 (
		\in3[119] ,
		_w782_,
		_w2280_,
		_w2282_,
		_w2283_
	);
	LUT3 #(
		.INIT('ha8)
	) name1770 (
		\in0[118] ,
		_w1038_,
		_w1045_,
		_w2284_
	);
	LUT3 #(
		.INIT('hb0)
	) name1771 (
		_w1029_,
		_w1043_,
		_w2284_,
		_w2285_
	);
	LUT4 #(
		.INIT('haa20)
	) name1772 (
		\in1[118] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2286_
	);
	LUT2 #(
		.INIT('h1)
	) name1773 (
		_w2285_,
		_w2286_,
		_w2287_
	);
	LUT3 #(
		.INIT('h02)
	) name1774 (
		\in3[118] ,
		_w2285_,
		_w2286_,
		_w2288_
	);
	LUT3 #(
		.INIT('h02)
	) name1775 (
		\in2[118] ,
		_w2285_,
		_w2286_,
		_w2289_
	);
	LUT3 #(
		.INIT('h1b)
	) name1776 (
		_w782_,
		_w2288_,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h8)
	) name1777 (
		_w2283_,
		_w2290_,
		_w2291_
	);
	LUT3 #(
		.INIT('ha8)
	) name1778 (
		\in0[117] ,
		_w1038_,
		_w1045_,
		_w2292_
	);
	LUT3 #(
		.INIT('hb0)
	) name1779 (
		_w1029_,
		_w1043_,
		_w2292_,
		_w2293_
	);
	LUT4 #(
		.INIT('haa20)
	) name1780 (
		\in1[117] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2294_
	);
	LUT2 #(
		.INIT('h1)
	) name1781 (
		_w2293_,
		_w2294_,
		_w2295_
	);
	LUT3 #(
		.INIT('ha8)
	) name1782 (
		\in2[117] ,
		_w521_,
		_w778_,
		_w2296_
	);
	LUT4 #(
		.INIT('h1500)
	) name1783 (
		_w526_,
		_w771_,
		_w776_,
		_w2296_,
		_w2297_
	);
	LUT4 #(
		.INIT('h0fdf)
	) name1784 (
		\in3[117] ,
		_w782_,
		_w2295_,
		_w2297_,
		_w2298_
	);
	LUT3 #(
		.INIT('ha8)
	) name1785 (
		\in0[116] ,
		_w1038_,
		_w1045_,
		_w2299_
	);
	LUT3 #(
		.INIT('hb0)
	) name1786 (
		_w1029_,
		_w1043_,
		_w2299_,
		_w2300_
	);
	LUT4 #(
		.INIT('haa20)
	) name1787 (
		\in1[116] ,
		_w1029_,
		_w1043_,
		_w1046_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name1788 (
		_w2300_,
		_w2301_,
		_w2302_
	);
	LUT3 #(
		.INIT('h02)
	) name1789 (
		\in3[116] ,
		_w2300_,
		_w2301_,
		_w2303_
	);
	LUT3 #(
		.INIT('h02)
	) name1790 (
		\in2[116] ,
		_w2300_,
		_w2301_,
		_w2304_
	);
	LUT3 #(
		.INIT('h1b)
	) name1791 (
		_w782_,
		_w2303_,
		_w2304_,
		_w2305_
	);
	LUT4 #(
		.INIT('h8000)
	) name1792 (
		_w2283_,
		_w2290_,
		_w2298_,
		_w2305_,
		_w2306_
	);
	LUT2 #(
		.INIT('h4)
	) name1793 (
		_w2276_,
		_w2306_,
		_w2307_
	);
	LUT4 #(
		.INIT('h000d)
	) name1794 (
		\in3[119] ,
		_w782_,
		_w2280_,
		_w2282_,
		_w2308_
	);
	LUT3 #(
		.INIT('ha8)
	) name1795 (
		\in2[116] ,
		_w521_,
		_w778_,
		_w2309_
	);
	LUT4 #(
		.INIT('h1500)
	) name1796 (
		_w526_,
		_w771_,
		_w776_,
		_w2309_,
		_w2310_
	);
	LUT4 #(
		.INIT('h000d)
	) name1797 (
		\in3[116] ,
		_w782_,
		_w2302_,
		_w2310_,
		_w2311_
	);
	LUT3 #(
		.INIT('ha8)
	) name1798 (
		\in2[118] ,
		_w521_,
		_w778_,
		_w2312_
	);
	LUT4 #(
		.INIT('h1500)
	) name1799 (
		_w526_,
		_w771_,
		_w776_,
		_w2312_,
		_w2313_
	);
	LUT4 #(
		.INIT('h000d)
	) name1800 (
		\in3[118] ,
		_w782_,
		_w2287_,
		_w2313_,
		_w2314_
	);
	LUT4 #(
		.INIT('h000d)
	) name1801 (
		\in3[117] ,
		_w782_,
		_w2295_,
		_w2297_,
		_w2315_
	);
	LUT4 #(
		.INIT('h0007)
	) name1802 (
		_w2298_,
		_w2311_,
		_w2314_,
		_w2315_,
		_w2316_
	);
	LUT3 #(
		.INIT('h31)
	) name1803 (
		_w2291_,
		_w2308_,
		_w2316_,
		_w2317_
	);
	LUT3 #(
		.INIT('h40)
	) name1804 (
		_w1077_,
		_w1118_,
		_w2317_,
		_w2318_
	);
	LUT4 #(
		.INIT('h4055)
	) name1805 (
		_w1119_,
		_w2271_,
		_w2307_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('hb)
	) name1806 (
		_w1078_,
		_w2319_,
		_w2320_
	);
	LUT4 #(
		.INIT('h4755)
	) name1807 (
		_w783_,
		_w1078_,
		_w1886_,
		_w2319_,
		_w2321_
	);
	LUT3 #(
		.INIT('h0d)
	) name1808 (
		\in3[1] ,
		_w782_,
		_w1889_,
		_w2322_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1809 (
		_w1078_,
		_w1879_,
		_w2319_,
		_w2322_,
		_w2323_
	);
	LUT3 #(
		.INIT('h0d)
	) name1810 (
		\in3[2] ,
		_w782_,
		_w1896_,
		_w2324_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1811 (
		_w1078_,
		_w1894_,
		_w2319_,
		_w2324_,
		_w2325_
	);
	LUT3 #(
		.INIT('h0d)
	) name1812 (
		\in3[3] ,
		_w782_,
		_w1872_,
		_w2326_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1813 (
		_w1078_,
		_w1870_,
		_w2319_,
		_w2326_,
		_w2327_
	);
	LUT3 #(
		.INIT('h0d)
	) name1814 (
		\in3[4] ,
		_w782_,
		_w1858_,
		_w2328_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1815 (
		_w1078_,
		_w1856_,
		_w2319_,
		_w2328_,
		_w2329_
	);
	LUT3 #(
		.INIT('h0d)
	) name1816 (
		\in3[5] ,
		_w782_,
		_w1917_,
		_w2330_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1817 (
		_w1078_,
		_w1863_,
		_w2319_,
		_w2330_,
		_w2331_
	);
	LUT4 #(
		.INIT('h1b0f)
	) name1818 (
		_w1078_,
		_w1912_,
		_w1921_,
		_w2319_,
		_w2332_
	);
	LUT3 #(
		.INIT('h0d)
	) name1819 (
		\in3[7] ,
		_w782_,
		_w1907_,
		_w2333_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1820 (
		_w1078_,
		_w1905_,
		_w2319_,
		_w2333_,
		_w2334_
	);
	LUT3 #(
		.INIT('h0d)
	) name1821 (
		\in3[8] ,
		_w782_,
		_w1942_,
		_w2335_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1822 (
		_w1078_,
		_w1940_,
		_w2319_,
		_w2335_,
		_w2336_
	);
	LUT3 #(
		.INIT('h0d)
	) name1823 (
		\in3[9] ,
		_w782_,
		_w1935_,
		_w2337_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1824 (
		_w1078_,
		_w1933_,
		_w2319_,
		_w2337_,
		_w2338_
	);
	LUT3 #(
		.INIT('h0d)
	) name1825 (
		\in3[10] ,
		_w782_,
		_w1928_,
		_w2339_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1826 (
		_w1078_,
		_w1926_,
		_w2319_,
		_w2339_,
		_w2340_
	);
	LUT3 #(
		.INIT('h0d)
	) name1827 (
		\in3[11] ,
		_w782_,
		_w1800_,
		_w2341_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1828 (
		_w1078_,
		_w1798_,
		_w2319_,
		_w2341_,
		_w2342_
	);
	LUT3 #(
		.INIT('h0d)
	) name1829 (
		\in3[12] ,
		_w782_,
		_w1793_,
		_w2343_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1830 (
		_w1078_,
		_w1791_,
		_w2319_,
		_w2343_,
		_w2344_
	);
	LUT3 #(
		.INIT('h0d)
	) name1831 (
		\in3[13] ,
		_w782_,
		_w1822_,
		_w2345_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1832 (
		_w1078_,
		_w1820_,
		_w2319_,
		_w2345_,
		_w2346_
	);
	LUT3 #(
		.INIT('h0d)
	) name1833 (
		\in3[14] ,
		_w782_,
		_w1808_,
		_w2347_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1834 (
		_w1078_,
		_w1806_,
		_w2319_,
		_w2347_,
		_w2348_
	);
	LUT3 #(
		.INIT('h0d)
	) name1835 (
		\in3[15] ,
		_w782_,
		_w1815_,
		_w2349_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1836 (
		_w1078_,
		_w1813_,
		_w2319_,
		_w2349_,
		_w2350_
	);
	LUT3 #(
		.INIT('h0d)
	) name1837 (
		\in3[16] ,
		_w782_,
		_w1848_,
		_w2351_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1838 (
		_w1078_,
		_w1846_,
		_w2319_,
		_w2351_,
		_w2352_
	);
	LUT3 #(
		.INIT('h0d)
	) name1839 (
		\in3[17] ,
		_w782_,
		_w1834_,
		_w2353_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1840 (
		_w1078_,
		_w1832_,
		_w2319_,
		_w2353_,
		_w2354_
	);
	LUT3 #(
		.INIT('h0d)
	) name1841 (
		\in3[18] ,
		_w782_,
		_w1841_,
		_w2355_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1842 (
		_w1078_,
		_w1839_,
		_w2319_,
		_w2355_,
		_w2356_
	);
	LUT3 #(
		.INIT('h0d)
	) name1843 (
		\in3[19] ,
		_w782_,
		_w1738_,
		_w2357_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1844 (
		_w1078_,
		_w1742_,
		_w2319_,
		_w2357_,
		_w2358_
	);
	LUT3 #(
		.INIT('h0d)
	) name1845 (
		\in3[20] ,
		_w782_,
		_w1734_,
		_w2359_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1846 (
		_w1078_,
		_w1732_,
		_w2319_,
		_w2359_,
		_w2360_
	);
	LUT3 #(
		.INIT('h0d)
	) name1847 (
		\in3[21] ,
		_w782_,
		_w1727_,
		_w2361_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1848 (
		_w1078_,
		_w1725_,
		_w2319_,
		_w2361_,
		_w2362_
	);
	LUT3 #(
		.INIT('h0d)
	) name1849 (
		\in3[22] ,
		_w782_,
		_w1764_,
		_w2363_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1850 (
		_w1078_,
		_w1762_,
		_w2319_,
		_w2363_,
		_w2364_
	);
	LUT3 #(
		.INIT('h0d)
	) name1851 (
		\in3[23] ,
		_w782_,
		_w1750_,
		_w2365_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1852 (
		_w1078_,
		_w1748_,
		_w2319_,
		_w2365_,
		_w2366_
	);
	LUT3 #(
		.INIT('h0d)
	) name1853 (
		\in3[24] ,
		_w782_,
		_w1757_,
		_w2367_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1854 (
		_w1078_,
		_w1755_,
		_w2319_,
		_w2367_,
		_w2368_
	);
	LUT3 #(
		.INIT('h0d)
	) name1855 (
		\in3[25] ,
		_w782_,
		_w1776_,
		_w2369_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1856 (
		_w1078_,
		_w1774_,
		_w2319_,
		_w2369_,
		_w2370_
	);
	LUT3 #(
		.INIT('h0d)
	) name1857 (
		\in3[26] ,
		_w782_,
		_w1783_,
		_w2371_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1858 (
		_w1078_,
		_w1781_,
		_w2319_,
		_w2371_,
		_w2372_
	);
	LUT3 #(
		.INIT('h0d)
	) name1859 (
		\in3[27] ,
		_w782_,
		_w1971_,
		_w2373_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1860 (
		_w1078_,
		_w1969_,
		_w2319_,
		_w2373_,
		_w2374_
	);
	LUT3 #(
		.INIT('h0d)
	) name1861 (
		\in3[28] ,
		_w782_,
		_w1635_,
		_w2375_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1862 (
		_w1078_,
		_w1633_,
		_w2319_,
		_w2375_,
		_w2376_
	);
	LUT3 #(
		.INIT('h0d)
	) name1863 (
		\in3[29] ,
		_w782_,
		_w1642_,
		_w2377_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1864 (
		_w1078_,
		_w1640_,
		_w2319_,
		_w2377_,
		_w2378_
	);
	LUT3 #(
		.INIT('h0d)
	) name1865 (
		\in3[30] ,
		_w782_,
		_w1717_,
		_w2379_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1866 (
		_w1078_,
		_w1715_,
		_w2319_,
		_w2379_,
		_w2380_
	);
	LUT3 #(
		.INIT('h0d)
	) name1867 (
		\in3[31] ,
		_w782_,
		_w1679_,
		_w2381_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1868 (
		_w1078_,
		_w1677_,
		_w2319_,
		_w2381_,
		_w2382_
	);
	LUT3 #(
		.INIT('h0d)
	) name1869 (
		\in3[32] ,
		_w782_,
		_w1991_,
		_w2383_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1870 (
		_w1078_,
		_w1670_,
		_w2319_,
		_w2383_,
		_w2384_
	);
	LUT3 #(
		.INIT('h0d)
	) name1871 (
		\in3[33] ,
		_w782_,
		_w1657_,
		_w2385_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1872 (
		_w1078_,
		_w1655_,
		_w2319_,
		_w2385_,
		_w2386_
	);
	LUT3 #(
		.INIT('h0d)
	) name1873 (
		\in3[34] ,
		_w782_,
		_w1986_,
		_w2387_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1874 (
		_w1078_,
		_w1648_,
		_w2319_,
		_w2387_,
		_w2388_
	);
	LUT3 #(
		.INIT('h0d)
	) name1875 (
		\in3[35] ,
		_w782_,
		_w1664_,
		_w2389_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1876 (
		_w1078_,
		_w1662_,
		_w2319_,
		_w2389_,
		_w2390_
	);
	LUT3 #(
		.INIT('h0d)
	) name1877 (
		\in3[36] ,
		_w782_,
		_w1686_,
		_w2391_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1878 (
		_w1078_,
		_w1684_,
		_w2319_,
		_w2391_,
		_w2392_
	);
	LUT3 #(
		.INIT('h0d)
	) name1879 (
		\in3[37] ,
		_w782_,
		_w1708_,
		_w2393_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1880 (
		_w1078_,
		_w1706_,
		_w2319_,
		_w2393_,
		_w2394_
	);
	LUT3 #(
		.INIT('h0d)
	) name1881 (
		\in3[38] ,
		_w782_,
		_w1980_,
		_w2395_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1882 (
		_w1078_,
		_w1692_,
		_w2319_,
		_w2395_,
		_w2396_
	);
	LUT3 #(
		.INIT('h0d)
	) name1883 (
		\in3[39] ,
		_w782_,
		_w1701_,
		_w2397_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1884 (
		_w1078_,
		_w1699_,
		_w2319_,
		_w2397_,
		_w2398_
	);
	LUT3 #(
		.INIT('h0d)
	) name1885 (
		\in3[40] ,
		_w782_,
		_w2054_,
		_w2399_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1886 (
		_w1078_,
		_w2058_,
		_w2319_,
		_w2399_,
		_w2400_
	);
	LUT3 #(
		.INIT('h0d)
	) name1887 (
		\in3[41] ,
		_w782_,
		_w2051_,
		_w2401_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1888 (
		_w1078_,
		_w2049_,
		_w2319_,
		_w2401_,
		_w2402_
	);
	LUT3 #(
		.INIT('h0d)
	) name1889 (
		\in3[42] ,
		_w782_,
		_w2043_,
		_w2403_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1890 (
		_w1078_,
		_w2041_,
		_w2319_,
		_w2403_,
		_w2404_
	);
	LUT3 #(
		.INIT('h0d)
	) name1891 (
		\in3[43] ,
		_w782_,
		_w2064_,
		_w2405_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1892 (
		_w1078_,
		_w2034_,
		_w2319_,
		_w2405_,
		_w2406_
	);
	LUT3 #(
		.INIT('h0d)
	) name1893 (
		\in3[44] ,
		_w782_,
		_w2029_,
		_w2407_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1894 (
		_w1078_,
		_w2027_,
		_w2319_,
		_w2407_,
		_w2408_
	);
	LUT3 #(
		.INIT('h0d)
	) name1895 (
		\in3[45] ,
		_w782_,
		_w2021_,
		_w2409_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1896 (
		_w1078_,
		_w2019_,
		_w2319_,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('h0d)
	) name1897 (
		\in3[46] ,
		_w782_,
		_w2075_,
		_w2411_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1898 (
		_w1078_,
		_w2005_,
		_w2319_,
		_w2411_,
		_w2412_
	);
	LUT3 #(
		.INIT('h0d)
	) name1899 (
		\in3[47] ,
		_w782_,
		_w2014_,
		_w2413_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1900 (
		_w1078_,
		_w2012_,
		_w2319_,
		_w2413_,
		_w2414_
	);
	LUT3 #(
		.INIT('h0d)
	) name1901 (
		\in3[48] ,
		_w782_,
		_w2150_,
		_w2415_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1902 (
		_w1078_,
		_w2141_,
		_w2319_,
		_w2415_,
		_w2416_
	);
	LUT3 #(
		.INIT('h0d)
	) name1903 (
		\in3[49] ,
		_w782_,
		_w2136_,
		_w2417_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1904 (
		_w1078_,
		_w2134_,
		_w2319_,
		_w2417_,
		_w2418_
	);
	LUT3 #(
		.INIT('h0d)
	) name1905 (
		\in3[50] ,
		_w782_,
		_w2156_,
		_w2419_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1906 (
		_w1078_,
		_w2127_,
		_w2319_,
		_w2419_,
		_w2420_
	);
	LUT3 #(
		.INIT('h0d)
	) name1907 (
		\in3[51] ,
		_w782_,
		_w2122_,
		_w2421_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1908 (
		_w1078_,
		_w2120_,
		_w2319_,
		_w2421_,
		_w2422_
	);
	LUT3 #(
		.INIT('h0d)
	) name1909 (
		\in3[52] ,
		_w782_,
		_w2162_,
		_w2423_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1910 (
		_w1078_,
		_w2105_,
		_w2319_,
		_w2423_,
		_w2424_
	);
	LUT3 #(
		.INIT('h0d)
	) name1911 (
		\in3[53] ,
		_w782_,
		_w2114_,
		_w2425_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1912 (
		_w1078_,
		_w2112_,
		_w2319_,
		_w2425_,
		_w2426_
	);
	LUT3 #(
		.INIT('h0d)
	) name1913 (
		\in3[54] ,
		_w782_,
		_w2166_,
		_w2427_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1914 (
		_w1078_,
		_w2097_,
		_w2319_,
		_w2427_,
		_w2428_
	);
	LUT3 #(
		.INIT('h0d)
	) name1915 (
		\in3[55] ,
		_w782_,
		_w2092_,
		_w2429_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1916 (
		_w1078_,
		_w2090_,
		_w2319_,
		_w2429_,
		_w2430_
	);
	LUT3 #(
		.INIT('h0d)
	) name1917 (
		\in3[56] ,
		_w782_,
		_w1610_,
		_w2431_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1918 (
		_w1078_,
		_w1608_,
		_w2319_,
		_w2431_,
		_w2432_
	);
	LUT3 #(
		.INIT('h0d)
	) name1919 (
		\in3[57] ,
		_w782_,
		_w1603_,
		_w2433_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1920 (
		_w1078_,
		_w1601_,
		_w2319_,
		_w2433_,
		_w2434_
	);
	LUT3 #(
		.INIT('h0d)
	) name1921 (
		\in3[58] ,
		_w782_,
		_w1581_,
		_w2435_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1922 (
		_w1078_,
		_w1579_,
		_w2319_,
		_w2435_,
		_w2436_
	);
	LUT3 #(
		.INIT('h0d)
	) name1923 (
		\in3[59] ,
		_w782_,
		_w1574_,
		_w2437_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1924 (
		_w1078_,
		_w1572_,
		_w2319_,
		_w2437_,
		_w2438_
	);
	LUT3 #(
		.INIT('h0d)
	) name1925 (
		\in3[60] ,
		_w782_,
		_w1588_,
		_w2439_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1926 (
		_w1078_,
		_w1586_,
		_w2319_,
		_w2439_,
		_w2440_
	);
	LUT3 #(
		.INIT('h0d)
	) name1927 (
		\in3[61] ,
		_w782_,
		_w1566_,
		_w2441_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1928 (
		_w1078_,
		_w1564_,
		_w2319_,
		_w2441_,
		_w2442_
	);
	LUT3 #(
		.INIT('h0d)
	) name1929 (
		\in3[62] ,
		_w782_,
		_w1615_,
		_w2443_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1930 (
		_w1078_,
		_w1594_,
		_w2319_,
		_w2443_,
		_w2444_
	);
	LUT3 #(
		.INIT('h0d)
	) name1931 (
		\in3[63] ,
		_w782_,
		_w1559_,
		_w2445_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1932 (
		_w1078_,
		_w1557_,
		_w2319_,
		_w2445_,
		_w2446_
	);
	LUT3 #(
		.INIT('h0d)
	) name1933 (
		\in3[64] ,
		_w782_,
		_w1512_,
		_w2447_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1934 (
		_w1078_,
		_w1516_,
		_w2319_,
		_w2447_,
		_w2448_
	);
	LUT3 #(
		.INIT('h0d)
	) name1935 (
		\in3[65] ,
		_w782_,
		_w1509_,
		_w2449_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1936 (
		_w1078_,
		_w1507_,
		_w2319_,
		_w2449_,
		_w2450_
	);
	LUT3 #(
		.INIT('h0d)
	) name1937 (
		\in3[66] ,
		_w782_,
		_w1520_,
		_w2451_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1938 (
		_w1078_,
		_w1499_,
		_w2319_,
		_w2451_,
		_w2452_
	);
	LUT3 #(
		.INIT('h0d)
	) name1939 (
		\in3[67] ,
		_w782_,
		_w1493_,
		_w2453_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1940 (
		_w1078_,
		_w1491_,
		_w2319_,
		_w2453_,
		_w2454_
	);
	LUT3 #(
		.INIT('h0d)
	) name1941 (
		\in3[68] ,
		_w782_,
		_w2179_,
		_w2455_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1942 (
		_w1078_,
		_w1548_,
		_w2319_,
		_w2455_,
		_w2456_
	);
	LUT3 #(
		.INIT('h0d)
	) name1943 (
		\in3[69] ,
		_w782_,
		_w1543_,
		_w2457_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1944 (
		_w1078_,
		_w1541_,
		_w2319_,
		_w2457_,
		_w2458_
	);
	LUT3 #(
		.INIT('h0d)
	) name1945 (
		\in3[70] ,
		_w782_,
		_w2182_,
		_w2459_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1946 (
		_w1078_,
		_w1533_,
		_w2319_,
		_w2459_,
		_w2460_
	);
	LUT3 #(
		.INIT('h0d)
	) name1947 (
		\in3[71] ,
		_w782_,
		_w1528_,
		_w2461_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1948 (
		_w1078_,
		_w1526_,
		_w2319_,
		_w2461_,
		_w2462_
	);
	LUT3 #(
		.INIT('h0d)
	) name1949 (
		\in3[72] ,
		_w782_,
		_w1479_,
		_w2463_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1950 (
		_w1078_,
		_w1465_,
		_w2319_,
		_w2463_,
		_w2464_
	);
	LUT3 #(
		.INIT('h0d)
	) name1951 (
		\in3[73] ,
		_w782_,
		_w1474_,
		_w2465_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1952 (
		_w1078_,
		_w1472_,
		_w2319_,
		_w2465_,
		_w2466_
	);
	LUT3 #(
		.INIT('h0d)
	) name1953 (
		\in3[74] ,
		_w782_,
		_w1483_,
		_w2467_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1954 (
		_w1078_,
		_w1457_,
		_w2319_,
		_w2467_,
		_w2468_
	);
	LUT3 #(
		.INIT('h0d)
	) name1955 (
		\in3[75] ,
		_w782_,
		_w1452_,
		_w2469_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1956 (
		_w1078_,
		_w1450_,
		_w2319_,
		_w2469_,
		_w2470_
	);
	LUT3 #(
		.INIT('h0d)
	) name1957 (
		\in3[76] ,
		_w782_,
		_w1405_,
		_w2471_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1958 (
		_w1078_,
		_w1409_,
		_w2319_,
		_w2471_,
		_w2472_
	);
	LUT3 #(
		.INIT('h0d)
	) name1959 (
		\in3[77] ,
		_w782_,
		_w1402_,
		_w2473_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1960 (
		_w1078_,
		_w1400_,
		_w2319_,
		_w2473_,
		_w2474_
	);
	LUT3 #(
		.INIT('h0d)
	) name1961 (
		\in3[78] ,
		_w782_,
		_w1412_,
		_w2475_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1962 (
		_w1078_,
		_w1392_,
		_w2319_,
		_w2475_,
		_w2476_
	);
	LUT3 #(
		.INIT('h0d)
	) name1963 (
		\in3[79] ,
		_w782_,
		_w1386_,
		_w2477_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1964 (
		_w1078_,
		_w1384_,
		_w2319_,
		_w2477_,
		_w2478_
	);
	LUT3 #(
		.INIT('h0d)
	) name1965 (
		\in3[80] ,
		_w782_,
		_w2197_,
		_w2479_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1966 (
		_w1078_,
		_w1441_,
		_w2319_,
		_w2479_,
		_w2480_
	);
	LUT3 #(
		.INIT('h0d)
	) name1967 (
		\in3[81] ,
		_w782_,
		_w1436_,
		_w2481_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1968 (
		_w1078_,
		_w1434_,
		_w2319_,
		_w2481_,
		_w2482_
	);
	LUT3 #(
		.INIT('h0d)
	) name1969 (
		\in3[82] ,
		_w782_,
		_w2201_,
		_w2483_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1970 (
		_w1078_,
		_w1426_,
		_w2319_,
		_w2483_,
		_w2484_
	);
	LUT3 #(
		.INIT('h0d)
	) name1971 (
		\in3[83] ,
		_w782_,
		_w1421_,
		_w2485_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1972 (
		_w1078_,
		_w1419_,
		_w2319_,
		_w2485_,
		_w2486_
	);
	LUT3 #(
		.INIT('h0d)
	) name1973 (
		\in3[84] ,
		_w782_,
		_w1372_,
		_w2487_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1974 (
		_w1078_,
		_w1322_,
		_w2319_,
		_w2487_,
		_w2488_
	);
	LUT3 #(
		.INIT('h0d)
	) name1975 (
		\in3[85] ,
		_w782_,
		_w1331_,
		_w2489_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1976 (
		_w1078_,
		_w1329_,
		_w2319_,
		_w2489_,
		_w2490_
	);
	LUT3 #(
		.INIT('h0d)
	) name1977 (
		\in3[86] ,
		_w782_,
		_w1375_,
		_w2491_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1978 (
		_w1078_,
		_w1314_,
		_w2319_,
		_w2491_,
		_w2492_
	);
	LUT3 #(
		.INIT('h0d)
	) name1979 (
		\in3[87] ,
		_w782_,
		_w1309_,
		_w2493_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1980 (
		_w1078_,
		_w1307_,
		_w2319_,
		_w2493_,
		_w2494_
	);
	LUT3 #(
		.INIT('h0d)
	) name1981 (
		\in3[88] ,
		_w782_,
		_w1358_,
		_w2495_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1982 (
		_w1078_,
		_w1362_,
		_w2319_,
		_w2495_,
		_w2496_
	);
	LUT3 #(
		.INIT('h0d)
	) name1983 (
		\in3[89] ,
		_w782_,
		_w1355_,
		_w2497_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1984 (
		_w1078_,
		_w1353_,
		_w2319_,
		_w2497_,
		_w2498_
	);
	LUT3 #(
		.INIT('h0d)
	) name1985 (
		\in3[90] ,
		_w782_,
		_w1366_,
		_w2499_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1986 (
		_w1078_,
		_w1345_,
		_w2319_,
		_w2499_,
		_w2500_
	);
	LUT3 #(
		.INIT('h0d)
	) name1987 (
		\in3[91] ,
		_w782_,
		_w1339_,
		_w2501_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1988 (
		_w1078_,
		_w1337_,
		_w2319_,
		_w2501_,
		_w2502_
	);
	LUT3 #(
		.INIT('h0d)
	) name1989 (
		\in3[92] ,
		_w782_,
		_w2245_,
		_w2503_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1990 (
		_w1078_,
		_w2236_,
		_w2319_,
		_w2503_,
		_w2504_
	);
	LUT3 #(
		.INIT('h0d)
	) name1991 (
		\in3[93] ,
		_w782_,
		_w2231_,
		_w2505_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1992 (
		_w1078_,
		_w2229_,
		_w2319_,
		_w2505_,
		_w2506_
	);
	LUT3 #(
		.INIT('h0d)
	) name1993 (
		\in3[94] ,
		_w782_,
		_w2248_,
		_w2507_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1994 (
		_w1078_,
		_w2221_,
		_w2319_,
		_w2507_,
		_w2508_
	);
	LUT3 #(
		.INIT('h0d)
	) name1995 (
		\in3[95] ,
		_w782_,
		_w2216_,
		_w2509_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1996 (
		_w1078_,
		_w2214_,
		_w2319_,
		_w2509_,
		_w2510_
	);
	LUT3 #(
		.INIT('h0d)
	) name1997 (
		\in3[96] ,
		_w782_,
		_w1295_,
		_w2511_
	);
	LUT4 #(
		.INIT('h10bf)
	) name1998 (
		_w1078_,
		_w1281_,
		_w2319_,
		_w2511_,
		_w2512_
	);
	LUT3 #(
		.INIT('h0d)
	) name1999 (
		\in3[97] ,
		_w782_,
		_w1290_,
		_w2513_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2000 (
		_w1078_,
		_w1288_,
		_w2319_,
		_w2513_,
		_w2514_
	);
	LUT3 #(
		.INIT('h0d)
	) name2001 (
		\in3[98] ,
		_w782_,
		_w1299_,
		_w2515_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2002 (
		_w1078_,
		_w1273_,
		_w2319_,
		_w2515_,
		_w2516_
	);
	LUT3 #(
		.INIT('h0d)
	) name2003 (
		\in3[99] ,
		_w782_,
		_w1268_,
		_w2517_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2004 (
		_w1078_,
		_w1266_,
		_w2319_,
		_w2517_,
		_w2518_
	);
	LUT3 #(
		.INIT('h0d)
	) name2005 (
		\in3[100] ,
		_w782_,
		_w1221_,
		_w2519_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2006 (
		_w1078_,
		_w1225_,
		_w2319_,
		_w2519_,
		_w2520_
	);
	LUT3 #(
		.INIT('h0d)
	) name2007 (
		\in3[101] ,
		_w782_,
		_w1218_,
		_w2521_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2008 (
		_w1078_,
		_w1216_,
		_w2319_,
		_w2521_,
		_w2522_
	);
	LUT3 #(
		.INIT('h0d)
	) name2009 (
		\in3[102] ,
		_w782_,
		_w1228_,
		_w2523_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2010 (
		_w1078_,
		_w1208_,
		_w2319_,
		_w2523_,
		_w2524_
	);
	LUT3 #(
		.INIT('h0d)
	) name2011 (
		\in3[103] ,
		_w782_,
		_w1202_,
		_w2525_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2012 (
		_w1078_,
		_w1200_,
		_w2319_,
		_w2525_,
		_w2526_
	);
	LUT3 #(
		.INIT('h0d)
	) name2013 (
		\in3[104] ,
		_w782_,
		_w2262_,
		_w2527_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2014 (
		_w1078_,
		_w1257_,
		_w2319_,
		_w2527_,
		_w2528_
	);
	LUT3 #(
		.INIT('h0d)
	) name2015 (
		\in3[105] ,
		_w782_,
		_w1252_,
		_w2529_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2016 (
		_w1078_,
		_w1250_,
		_w2319_,
		_w2529_,
		_w2530_
	);
	LUT3 #(
		.INIT('h0d)
	) name2017 (
		\in3[106] ,
		_w782_,
		_w2266_,
		_w2531_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2018 (
		_w1078_,
		_w1242_,
		_w2319_,
		_w2531_,
		_w2532_
	);
	LUT3 #(
		.INIT('h0d)
	) name2019 (
		\in3[107] ,
		_w782_,
		_w1237_,
		_w2533_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2020 (
		_w1078_,
		_w1235_,
		_w2319_,
		_w2533_,
		_w2534_
	);
	LUT3 #(
		.INIT('h0d)
	) name2021 (
		\in3[108] ,
		_w782_,
		_w1188_,
		_w2535_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2022 (
		_w1078_,
		_w1138_,
		_w2319_,
		_w2535_,
		_w2536_
	);
	LUT3 #(
		.INIT('h0d)
	) name2023 (
		\in3[109] ,
		_w782_,
		_w1147_,
		_w2537_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2024 (
		_w1078_,
		_w1145_,
		_w2319_,
		_w2537_,
		_w2538_
	);
	LUT3 #(
		.INIT('h0d)
	) name2025 (
		\in3[110] ,
		_w782_,
		_w1191_,
		_w2539_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2026 (
		_w1078_,
		_w1130_,
		_w2319_,
		_w2539_,
		_w2540_
	);
	LUT3 #(
		.INIT('h0d)
	) name2027 (
		\in3[111] ,
		_w782_,
		_w1125_,
		_w2541_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2028 (
		_w1078_,
		_w1123_,
		_w2319_,
		_w2541_,
		_w2542_
	);
	LUT3 #(
		.INIT('h0d)
	) name2029 (
		\in3[112] ,
		_w782_,
		_w1174_,
		_w2543_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2030 (
		_w1078_,
		_w1178_,
		_w2319_,
		_w2543_,
		_w2544_
	);
	LUT3 #(
		.INIT('h0d)
	) name2031 (
		\in3[113] ,
		_w782_,
		_w1171_,
		_w2545_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2032 (
		_w1078_,
		_w1169_,
		_w2319_,
		_w2545_,
		_w2546_
	);
	LUT3 #(
		.INIT('h0d)
	) name2033 (
		\in3[114] ,
		_w782_,
		_w1182_,
		_w2547_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2034 (
		_w1078_,
		_w1161_,
		_w2319_,
		_w2547_,
		_w2548_
	);
	LUT3 #(
		.INIT('h0d)
	) name2035 (
		\in3[115] ,
		_w782_,
		_w1155_,
		_w2549_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2036 (
		_w1078_,
		_w1153_,
		_w2319_,
		_w2549_,
		_w2550_
	);
	LUT3 #(
		.INIT('h0d)
	) name2037 (
		\in3[116] ,
		_w782_,
		_w2310_,
		_w2551_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2038 (
		_w1078_,
		_w2302_,
		_w2319_,
		_w2551_,
		_w2552_
	);
	LUT3 #(
		.INIT('h0d)
	) name2039 (
		\in3[117] ,
		_w782_,
		_w2297_,
		_w2553_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2040 (
		_w1078_,
		_w2295_,
		_w2319_,
		_w2553_,
		_w2554_
	);
	LUT3 #(
		.INIT('h0d)
	) name2041 (
		\in3[118] ,
		_w782_,
		_w2313_,
		_w2555_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2042 (
		_w1078_,
		_w2287_,
		_w2319_,
		_w2555_,
		_w2556_
	);
	LUT3 #(
		.INIT('h0d)
	) name2043 (
		\in3[119] ,
		_w782_,
		_w2282_,
		_w2557_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2044 (
		_w1078_,
		_w2280_,
		_w2319_,
		_w2557_,
		_w2558_
	);
	LUT3 #(
		.INIT('h0d)
	) name2045 (
		\in3[120] ,
		_w782_,
		_w1111_,
		_w2559_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2046 (
		_w1078_,
		_w1097_,
		_w2319_,
		_w2559_,
		_w2560_
	);
	LUT3 #(
		.INIT('h0d)
	) name2047 (
		\in3[121] ,
		_w782_,
		_w1106_,
		_w2561_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2048 (
		_w1078_,
		_w1104_,
		_w2319_,
		_w2561_,
		_w2562_
	);
	LUT3 #(
		.INIT('h0d)
	) name2049 (
		\in3[122] ,
		_w782_,
		_w1115_,
		_w2563_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2050 (
		_w1078_,
		_w1089_,
		_w2319_,
		_w2563_,
		_w2564_
	);
	LUT3 #(
		.INIT('h0d)
	) name2051 (
		\in3[123] ,
		_w782_,
		_w1084_,
		_w2565_
	);
	LUT4 #(
		.INIT('h10bf)
	) name2052 (
		_w1078_,
		_w1082_,
		_w2319_,
		_w2565_,
		_w2566_
	);
	LUT3 #(
		.INIT('h0d)
	) name2053 (
		\in3[124] ,
		_w782_,
		_w1068_,
		_w2567_
	);
	LUT4 #(
		.INIT('h10df)
	) name2054 (
		_w1066_,
		_w1078_,
		_w2319_,
		_w2567_,
		_w2568_
	);
	LUT3 #(
		.INIT('h0d)
	) name2055 (
		\in3[125] ,
		_w782_,
		_w1060_,
		_w2569_
	);
	LUT4 #(
		.INIT('h10df)
	) name2056 (
		_w1058_,
		_w1078_,
		_w2319_,
		_w2569_,
		_w2570_
	);
	LUT3 #(
		.INIT('h0d)
	) name2057 (
		\in3[126] ,
		_w782_,
		_w1053_,
		_w2571_
	);
	LUT4 #(
		.INIT('h10df)
	) name2058 (
		_w1051_,
		_w1078_,
		_w2319_,
		_w2571_,
		_w2572_
	);
	LUT4 #(
		.INIT('h8000)
	) name2059 (
		\in0[127] ,
		\in1[127] ,
		\in2[127] ,
		\in3[127] ,
		_w2573_
	);
	LUT4 #(
		.INIT('h5355)
	) name2060 (
		_w782_,
		_w1049_,
		_w1078_,
		_w2319_,
		_w2574_
	);
	assign \result[0]  = _w2321_ ;
	assign \result[1]  = _w2323_ ;
	assign \result[2]  = _w2325_ ;
	assign \result[3]  = _w2327_ ;
	assign \result[4]  = _w2329_ ;
	assign \result[5]  = _w2331_ ;
	assign \result[6]  = _w2332_ ;
	assign \result[7]  = _w2334_ ;
	assign \result[8]  = _w2336_ ;
	assign \result[9]  = _w2338_ ;
	assign \result[10]  = _w2340_ ;
	assign \result[11]  = _w2342_ ;
	assign \result[12]  = _w2344_ ;
	assign \result[13]  = _w2346_ ;
	assign \result[14]  = _w2348_ ;
	assign \result[15]  = _w2350_ ;
	assign \result[16]  = _w2352_ ;
	assign \result[17]  = _w2354_ ;
	assign \result[18]  = _w2356_ ;
	assign \result[19]  = _w2358_ ;
	assign \result[20]  = _w2360_ ;
	assign \result[21]  = _w2362_ ;
	assign \result[22]  = _w2364_ ;
	assign \result[23]  = _w2366_ ;
	assign \result[24]  = _w2368_ ;
	assign \result[25]  = _w2370_ ;
	assign \result[26]  = _w2372_ ;
	assign \result[27]  = _w2374_ ;
	assign \result[28]  = _w2376_ ;
	assign \result[29]  = _w2378_ ;
	assign \result[30]  = _w2380_ ;
	assign \result[31]  = _w2382_ ;
	assign \result[32]  = _w2384_ ;
	assign \result[33]  = _w2386_ ;
	assign \result[34]  = _w2388_ ;
	assign \result[35]  = _w2390_ ;
	assign \result[36]  = _w2392_ ;
	assign \result[37]  = _w2394_ ;
	assign \result[38]  = _w2396_ ;
	assign \result[39]  = _w2398_ ;
	assign \result[40]  = _w2400_ ;
	assign \result[41]  = _w2402_ ;
	assign \result[42]  = _w2404_ ;
	assign \result[43]  = _w2406_ ;
	assign \result[44]  = _w2408_ ;
	assign \result[45]  = _w2410_ ;
	assign \result[46]  = _w2412_ ;
	assign \result[47]  = _w2414_ ;
	assign \result[48]  = _w2416_ ;
	assign \result[49]  = _w2418_ ;
	assign \result[50]  = _w2420_ ;
	assign \result[51]  = _w2422_ ;
	assign \result[52]  = _w2424_ ;
	assign \result[53]  = _w2426_ ;
	assign \result[54]  = _w2428_ ;
	assign \result[55]  = _w2430_ ;
	assign \result[56]  = _w2432_ ;
	assign \result[57]  = _w2434_ ;
	assign \result[58]  = _w2436_ ;
	assign \result[59]  = _w2438_ ;
	assign \result[60]  = _w2440_ ;
	assign \result[61]  = _w2442_ ;
	assign \result[62]  = _w2444_ ;
	assign \result[63]  = _w2446_ ;
	assign \result[64]  = _w2448_ ;
	assign \result[65]  = _w2450_ ;
	assign \result[66]  = _w2452_ ;
	assign \result[67]  = _w2454_ ;
	assign \result[68]  = _w2456_ ;
	assign \result[69]  = _w2458_ ;
	assign \result[70]  = _w2460_ ;
	assign \result[71]  = _w2462_ ;
	assign \result[72]  = _w2464_ ;
	assign \result[73]  = _w2466_ ;
	assign \result[74]  = _w2468_ ;
	assign \result[75]  = _w2470_ ;
	assign \result[76]  = _w2472_ ;
	assign \result[77]  = _w2474_ ;
	assign \result[78]  = _w2476_ ;
	assign \result[79]  = _w2478_ ;
	assign \result[80]  = _w2480_ ;
	assign \result[81]  = _w2482_ ;
	assign \result[82]  = _w2484_ ;
	assign \result[83]  = _w2486_ ;
	assign \result[84]  = _w2488_ ;
	assign \result[85]  = _w2490_ ;
	assign \result[86]  = _w2492_ ;
	assign \result[87]  = _w2494_ ;
	assign \result[88]  = _w2496_ ;
	assign \result[89]  = _w2498_ ;
	assign \result[90]  = _w2500_ ;
	assign \result[91]  = _w2502_ ;
	assign \result[92]  = _w2504_ ;
	assign \result[93]  = _w2506_ ;
	assign \result[94]  = _w2508_ ;
	assign \result[95]  = _w2510_ ;
	assign \result[96]  = _w2512_ ;
	assign \result[97]  = _w2514_ ;
	assign \result[98]  = _w2516_ ;
	assign \result[99]  = _w2518_ ;
	assign \result[100]  = _w2520_ ;
	assign \result[101]  = _w2522_ ;
	assign \result[102]  = _w2524_ ;
	assign \result[103]  = _w2526_ ;
	assign \result[104]  = _w2528_ ;
	assign \result[105]  = _w2530_ ;
	assign \result[106]  = _w2532_ ;
	assign \result[107]  = _w2534_ ;
	assign \result[108]  = _w2536_ ;
	assign \result[109]  = _w2538_ ;
	assign \result[110]  = _w2540_ ;
	assign \result[111]  = _w2542_ ;
	assign \result[112]  = _w2544_ ;
	assign \result[113]  = _w2546_ ;
	assign \result[114]  = _w2548_ ;
	assign \result[115]  = _w2550_ ;
	assign \result[116]  = _w2552_ ;
	assign \result[117]  = _w2554_ ;
	assign \result[118]  = _w2556_ ;
	assign \result[119]  = _w2558_ ;
	assign \result[120]  = _w2560_ ;
	assign \result[121]  = _w2562_ ;
	assign \result[122]  = _w2564_ ;
	assign \result[123]  = _w2566_ ;
	assign \result[124]  = _w2568_ ;
	assign \result[125]  = _w2570_ ;
	assign \result[126]  = _w2572_ ;
	assign \result[127]  = _w2573_ ;
	assign \address[0]  = _w2574_ ;
	assign \address[1]  = _w2320_ ;
endmodule;