module top (\a0_pad , a_pad, b_pad, \c0_pad , c_pad, \d0_pad , d_pad, \e0_pad , e_pad, \f0_pad , f_pad, \g0_pad , g_pad, \h0_pad , h_pad, \i0_pad , i_pad, j_pad, k_pad, l_pad, m_pad, n_pad, o_pad, p_pad, q_pad, r_pad, s_pad, t_pad, u_pad, v_pad, w_pad, x_pad, y_pad, z_pad, \j0_pad , \k0_pad , \l0_pad , \m0_pad , \n0_pad , \o0_pad , \p0_pad , \q0_pad , \r0_pad , \s0_pad );
	input \a0_pad  ;
	input a_pad ;
	input b_pad ;
	input \c0_pad  ;
	input c_pad ;
	input \d0_pad  ;
	input d_pad ;
	input \e0_pad  ;
	input e_pad ;
	input \f0_pad  ;
	input f_pad ;
	input \g0_pad  ;
	input g_pad ;
	input \h0_pad  ;
	input h_pad ;
	input \i0_pad  ;
	input i_pad ;
	input j_pad ;
	input k_pad ;
	input l_pad ;
	input m_pad ;
	input n_pad ;
	input o_pad ;
	input p_pad ;
	input q_pad ;
	input r_pad ;
	input s_pad ;
	input t_pad ;
	input u_pad ;
	input v_pad ;
	input w_pad ;
	input x_pad ;
	input y_pad ;
	input z_pad ;
	output \j0_pad  ;
	output \k0_pad  ;
	output \l0_pad  ;
	output \m0_pad  ;
	output \n0_pad  ;
	output \o0_pad  ;
	output \p0_pad  ;
	output \q0_pad  ;
	output \r0_pad  ;
	output \s0_pad  ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w103_ ;
	wire _w102_ ;
	wire _w101_ ;
	wire _w100_ ;
	wire _w99_ ;
	wire _w98_ ;
	wire _w97_ ;
	wire _w96_ ;
	wire _w95_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w57_ ;
	wire _w56_ ;
	wire _w55_ ;
	wire _w54_ ;
	wire _w53_ ;
	wire _w52_ ;
	wire _w51_ ;
	wire _w50_ ;
	wire _w49_ ;
	wire _w42_ ;
	wire _w37_ ;
	wire _w38_ ;
	wire _w39_ ;
	wire _w40_ ;
	wire _w41_ ;
	wire _w43_ ;
	wire _w44_ ;
	wire _w16_ ;
	wire _w75_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w65_ ;
	wire _w66_ ;
	wire _w67_ ;
	wire _w68_ ;
	wire _w69_ ;
	wire _w70_ ;
	wire _w71_ ;
	wire _w72_ ;
	wire _w73_ ;
	wire _w74_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\h0_pad ,
		_w16_
	);
	LUT2 #(
		.INIT('h8)
	) name1 (
		c_pad,
		d_pad,
		_w37_
	);
	LUT2 #(
		.INIT('h6)
	) name2 (
		c_pad,
		d_pad,
		_w38_
	);
	LUT4 #(
		.INIT('h069f)
	) name3 (
		c_pad,
		d_pad,
		\h0_pad ,
		\i0_pad ,
		_w39_
	);
	LUT2 #(
		.INIT('h9)
	) name4 (
		e_pad,
		h_pad,
		_w40_
	);
	LUT4 #(
		.INIT('h9acf)
	) name5 (
		c_pad,
		d_pad,
		f_pad,
		g_pad,
		_w41_
	);
	LUT3 #(
		.INIT('h41)
	) name6 (
		b_pad,
		_w40_,
		_w41_,
		_w42_
	);
	LUT2 #(
		.INIT('h2)
	) name7 (
		i_pad,
		j_pad,
		_w43_
	);
	LUT4 #(
		.INIT('h7d00)
	) name8 (
		b_pad,
		_w38_,
		_w40_,
		_w43_,
		_w44_
	);
	LUT2 #(
		.INIT('h4)
	) name9 (
		_w42_,
		_w44_,
		_w45_
	);
	LUT4 #(
		.INIT('hfac8)
	) name10 (
		p_pad,
		q_pad,
		u_pad,
		v_pad,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		s_pad,
		x_pad,
		_w47_
	);
	LUT4 #(
		.INIT('hfac8)
	) name12 (
		r_pad,
		t_pad,
		w_pad,
		y_pad,
		_w48_
	);
	LUT3 #(
		.INIT('h40)
	) name13 (
		_w47_,
		_w46_,
		_w48_,
		_w49_
	);
	LUT3 #(
		.INIT('h40)
	) name14 (
		\a0_pad ,
		b_pad,
		z_pad,
		_w50_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		_w37_,
		_w50_,
		_w51_
	);
	LUT3 #(
		.INIT('h10)
	) name16 (
		\c0_pad ,
		_w49_,
		_w51_,
		_w52_
	);
	LUT2 #(
		.INIT('h6)
	) name17 (
		\c0_pad ,
		\d0_pad ,
		_w53_
	);
	LUT3 #(
		.INIT('h40)
	) name18 (
		_w49_,
		_w51_,
		_w53_,
		_w54_
	);
	LUT3 #(
		.INIT('h80)
	) name19 (
		\c0_pad ,
		\d0_pad ,
		\e0_pad ,
		_w55_
	);
	LUT3 #(
		.INIT('h78)
	) name20 (
		\c0_pad ,
		\d0_pad ,
		\e0_pad ,
		_w56_
	);
	LUT3 #(
		.INIT('h40)
	) name21 (
		_w49_,
		_w51_,
		_w56_,
		_w57_
	);
	LUT4 #(
		.INIT('h7f80)
	) name22 (
		\c0_pad ,
		\d0_pad ,
		\e0_pad ,
		\f0_pad ,
		_w58_
	);
	LUT3 #(
		.INIT('h40)
	) name23 (
		_w49_,
		_w51_,
		_w58_,
		_w59_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		\f0_pad ,
		\g0_pad ,
		_w60_
	);
	LUT2 #(
		.INIT('h8)
	) name25 (
		\f0_pad ,
		\g0_pad ,
		_w61_
	);
	LUT2 #(
		.INIT('h6)
	) name26 (
		\f0_pad ,
		\g0_pad ,
		_w62_
	);
	LUT3 #(
		.INIT('h93)
	) name27 (
		\f0_pad ,
		\g0_pad ,
		_w55_,
		_w63_
	);
	LUT3 #(
		.INIT('hbf)
	) name28 (
		_w49_,
		_w51_,
		_w63_,
		_w64_
	);
	LUT3 #(
		.INIT('h80)
	) name29 (
		r_pad,
		s_pad,
		t_pad,
		_w65_
	);
	LUT4 #(
		.INIT('h4000)
	) name30 (
		l_pad,
		r_pad,
		s_pad,
		t_pad,
		_w66_
	);
	LUT2 #(
		.INIT('h1)
	) name31 (
		q_pad,
		_w66_,
		_w67_
	);
	LUT3 #(
		.INIT('h40)
	) name32 (
		m_pad,
		s_pad,
		t_pad,
		_w68_
	);
	LUT4 #(
		.INIT('h0acf)
	) name33 (
		n_pad,
		o_pad,
		s_pad,
		t_pad,
		_w69_
	);
	LUT3 #(
		.INIT('h31)
	) name34 (
		r_pad,
		_w68_,
		_w69_,
		_w70_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		q_pad,
		r_pad,
		_w71_
	);
	LUT3 #(
		.INIT('h40)
	) name36 (
		p_pad,
		s_pad,
		t_pad,
		_w72_
	);
	LUT2 #(
		.INIT('h8)
	) name37 (
		_w71_,
		_w72_,
		_w73_
	);
	LUT4 #(
		.INIT('h0057)
	) name38 (
		p_pad,
		_w67_,
		_w70_,
		_w73_,
		_w74_
	);
	LUT3 #(
		.INIT('he8)
	) name39 (
		r_pad,
		s_pad,
		t_pad,
		_w75_
	);
	LUT4 #(
		.INIT('h177f)
	) name40 (
		q_pad,
		r_pad,
		s_pad,
		t_pad,
		_w76_
	);
	LUT3 #(
		.INIT('he0)
	) name41 (
		\c0_pad ,
		\d0_pad ,
		\e0_pad ,
		_w77_
	);
	LUT4 #(
		.INIT('h1fe0)
	) name42 (
		\c0_pad ,
		\d0_pad ,
		\e0_pad ,
		\f0_pad ,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name43 (
		\g0_pad ,
		_w78_,
		_w79_
	);
	LUT3 #(
		.INIT('h40)
	) name44 (
		k_pad,
		s_pad,
		t_pad,
		_w80_
	);
	LUT3 #(
		.INIT('h2a)
	) name45 (
		\h0_pad ,
		_w71_,
		_w80_,
		_w81_
	);
	LUT3 #(
		.INIT('h20)
	) name46 (
		_w79_,
		_w76_,
		_w81_,
		_w82_
	);
	LUT2 #(
		.INIT('h4)
	) name47 (
		_w74_,
		_w82_,
		_w83_
	);
	LUT4 #(
		.INIT('hf53f)
	) name48 (
		m_pad,
		n_pad,
		r_pad,
		s_pad,
		_w84_
	);
	LUT3 #(
		.INIT('h80)
	) name49 (
		p_pad,
		q_pad,
		t_pad,
		_w85_
	);
	LUT2 #(
		.INIT('h4)
	) name50 (
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		l_pad,
		q_pad,
		_w87_
	);
	LUT4 #(
		.INIT('hf531)
	) name52 (
		k_pad,
		l_pad,
		p_pad,
		q_pad,
		_w88_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		p_pad,
		q_pad,
		_w89_
	);
	LUT3 #(
		.INIT('h04)
	) name54 (
		_w89_,
		_w65_,
		_w88_,
		_w90_
	);
	LUT3 #(
		.INIT('h80)
	) name55 (
		q_pad,
		r_pad,
		s_pad,
		_w91_
	);
	LUT3 #(
		.INIT('h08)
	) name56 (
		o_pad,
		p_pad,
		t_pad,
		_w92_
	);
	LUT2 #(
		.INIT('h8)
	) name57 (
		_w91_,
		_w92_,
		_w93_
	);
	LUT4 #(
		.INIT('haaa8)
	) name58 (
		_w79_,
		_w90_,
		_w93_,
		_w86_,
		_w94_
	);
	LUT2 #(
		.INIT('h4)
	) name59 (
		\a0_pad ,
		a_pad,
		_w95_
	);
	LUT3 #(
		.INIT('he0)
	) name60 (
		\h0_pad ,
		_w94_,
		_w95_,
		_w96_
	);
	LUT2 #(
		.INIT('h4)
	) name61 (
		_w83_,
		_w96_,
		_w97_
	);
	LUT4 #(
		.INIT('ha0a8)
	) name62 (
		q_pad,
		r_pad,
		_w68_,
		_w69_,
		_w98_
	);
	LUT4 #(
		.INIT('h0008)
	) name63 (
		_w61_,
		_w77_,
		_w76_,
		_w66_,
		_w99_
	);
	LUT2 #(
		.INIT('h4)
	) name64 (
		_w98_,
		_w99_,
		_w100_
	);
	LUT4 #(
		.INIT('h8ccc)
	) name65 (
		m_pad,
		q_pad,
		s_pad,
		t_pad,
		_w101_
	);
	LUT4 #(
		.INIT('hc400)
	) name66 (
		r_pad,
		_w75_,
		_w69_,
		_w101_,
		_w102_
	);
	LUT2 #(
		.INIT('h8)
	) name67 (
		_w65_,
		_w87_,
		_w103_
	);
	LUT2 #(
		.INIT('h2)
	) name68 (
		_w60_,
		_w77_,
		_w104_
	);
	LUT3 #(
		.INIT('he0)
	) name69 (
		_w102_,
		_w103_,
		_w104_,
		_w105_
	);
	LUT2 #(
		.INIT('h1)
	) name70 (
		_w62_,
		_w78_,
		_w106_
	);
	LUT3 #(
		.INIT('h20)
	) name71 (
		k_pad,
		p_pad,
		t_pad,
		_w107_
	);
	LUT4 #(
		.INIT('h1000)
	) name72 (
		_w62_,
		_w78_,
		_w91_,
		_w107_,
		_w108_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\i0_pad ,
		_w108_,
		_w109_
	);
	LUT4 #(
		.INIT('h5700)
	) name74 (
		p_pad,
		_w100_,
		_w105_,
		_w109_,
		_w110_
	);
	LUT4 #(
		.INIT('h020a)
	) name75 (
		\i0_pad ,
		_w71_,
		_w76_,
		_w80_,
		_w111_
	);
	LUT2 #(
		.INIT('h8)
	) name76 (
		_w106_,
		_w111_,
		_w112_
	);
	LUT3 #(
		.INIT('h8a)
	) name77 (
		_w95_,
		_w74_,
		_w112_,
		_w113_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w110_,
		_w113_,
		_w114_
	);
	assign \j0_pad  = _w16_ ;
	assign \k0_pad  = _w39_ ;
	assign \l0_pad  = _w45_ ;
	assign \m0_pad  = _w52_ ;
	assign \n0_pad  = _w54_ ;
	assign \o0_pad  = _w57_ ;
	assign \p0_pad  = _w59_ ;
	assign \q0_pad  = _w64_ ;
	assign \r0_pad  = _w97_ ;
	assign \s0_pad  = _w114_ ;
endmodule;