module top (\g1000_reg/NET0131 , \g1001_reg/NET0131 , \g1002_reg/NET0131 , \g1003_reg/NET0131 , \g1004_reg/NET0131 , \g1005_reg/NET0131 , \g1006_reg/NET0131 , \g1007_reg/NET0131 , \g1008_reg/NET0131 , \g1009_reg/NET0131 , \g1010_reg/NET0131 , \g1011_reg/NET0131 , \g1018_reg/NET0131 , \g101_reg/NET0131 , \g1024_reg/NET0131 , \g1030_reg/NET0131 , \g1033_reg/NET0131 , \g1036_reg/NET0131 , \g1038_reg/NET0131 , \g1040_reg/NET0131 , \g1041_reg/NET0131 , \g1045_reg/NET0131 , \g1048_reg/NET0131 , \g1051_reg/NET0131 , \g1053_reg/NET0131 , \g1055_reg/NET0131 , \g1056_reg/NET0131 , \g105_reg/NET0131 , \g1060_reg/NET0131 , \g1063_reg/NET0131 , \g1066_reg/NET0131 , \g1068_reg/NET0131 , \g1070_reg/NET0131 , \g1071_reg/NET0131 , \g1075_reg/NET0131 , \g1078_reg/NET0131 , \g1081_reg/NET0131 , \g1083_reg/NET0131 , \g1085_reg/NET0131 , \g1088_reg/NET0131 , \g1089_reg/NET0131 , \g1090_reg/NET0131 , \g1091_reg/NET0131 , \g1092_reg/NET0131 , \g1095_reg/NET0131 , \g1098_reg/NET0131 , \g109_reg/NET0131 , \g1101_reg/NET0131 , \g1104_reg/NET0131 , \g1107_reg/NET0131 , \g1110_reg/NET0131 , \g1113_reg/NET0131 , \g1114_reg/NET0131 , \g1115_reg/NET0131 , \g1116_reg/NET0131 , \g1119_reg/NET0131 , \g1122_reg/NET0131 , \g1125_reg/NET0131 , \g1128_reg/NET0131 , \g1131_reg/NET0131 , \g1134_reg/NET0131 , \g1135_reg/NET0131 , \g1136_reg/NET0131 , \g1138_reg/NET0131 , \g113_reg/NET0131 , \g1140_reg/NET0131 , \g1151_reg/NET0131 , \g1164_reg/NET0131 , \g1165_reg/NET0131 , \g1166_reg/NET0131 , \g1167_reg/NET0131 , \g1171_reg/NET0131 , \g1173_reg/NET0131 , \g1174_reg/NET0131 , \g1175_reg/NET0131 , \g1176_reg/NET0131 , \g1177_reg/NET0131 , \g117_reg/NET0131 , \g1180_reg/NET0131 , \g1183_reg/NET0131 , \g1186_reg/NET0131 , \g1192_reg/NET0131 , \g1193_reg/NET0131 , \g1196_reg/NET0131 , \g1210_reg/NET0131 , \g1211_reg/NET0131 , \g1215_reg/NET0131 , \g1216_reg/NET0131 , \g1217_reg/NET0131 , \g1218_reg/NET0131 , \g1219_reg/NET0131 , \g121_reg/NET0131 , \g1220_reg/NET0131 , \g1222_reg/NET0131 , \g1223_reg/NET0131 , \g1224_reg/NET0131 , \g1227_reg/NET0131 , \g1228_reg/NET0131 , \g1230_reg/NET0131 , \g1234_reg/NET0131 , \g1240_reg/NET0131 , \g1243_reg/NET0131 , \g1245_reg/NET0131 , \g1249_pad , \g1251_reg/NET0131 , \g1253_reg/NET0131 , \g1255_reg/NET0131 , \g1257_reg/NET0131 , \g1259_reg/NET0131 , \g125_reg/NET0131 , \g1261_reg/NET0131 , \g1262_reg/NET0131 , \g1263_reg/NET0131 , \g1264_reg/NET0131 , \g1265_reg/NET0131 , \g1266_reg/NET0131 , \g1267_reg/NET0131 , \g1268_reg/NET0131 , \g1269_reg/NET0131 , \g1270_reg/NET0131 , \g1271_reg/NET0131 , \g1272_reg/NET0131 , \g1273_reg/NET0131 , \g1276_reg/NET0131 , \g1279_reg/NET0131 , \g1282_reg/NET0131 , \g1285_reg/NET0131 , \g1288_reg/NET0131 , \g1291_reg/NET0131 , \g1294_reg/NET0131 , \g1297_reg/NET0131 , \g129_reg/NET0131 , \g1300_reg/NET0131 , \g1303_reg/NET0131 , \g1306_reg/NET0131 , \g130_reg/NET0131 , \g1316_reg/NET0131 , \g1319_reg/NET0131 , \g131_reg/NET0131 , \g1326_reg/NET0131 , \g132_reg/NET0131 , \g1332_reg/NET0131 , \g1339_reg/NET0131 , \g133_reg/NET0131 , \g1345_reg/NET0131 , \g1346_reg/NET0131 , \g134_reg/NET0131 , \g1352_reg/NET0131 , \g1358_reg/NET0131 , \g1365_reg/NET0131 , \g1372_reg/NET0131 , \g1378_reg/NET0131 , \g1384_reg/NET0131 , \g1385_reg/NET0131 , \g1386_reg/NET0131 , \g1387_reg/NET0131 , \g1388_reg/NET0131 , \g1389_reg/NET0131 , \g1390_reg/NET0131 , \g1391_reg/NET0131 , \g1392_reg/NET0131 , \g1393_reg/NET0131 , \g1394_reg/NET0131 , \g1395_reg/NET0131 , \g1396_reg/NET0131 , \g1397_reg/NET0131 , \g1398_reg/NET0131 , \g1399_reg/NET0131 , \g1400_reg/NET0131 , \g1401_reg/NET0131 , \g1402_reg/NET0131 , \g1403_reg/NET0131 , \g1404_reg/NET0131 , \g1405_reg/NET0131 , \g1406_reg/NET0131 , \g1407_reg/NET0131 , \g1408_reg/NET0131 , \g1409_reg/NET0131 , \g1410_reg/NET0131 , \g1411_reg/NET0131 , \g1412_reg/NET0131 , \g1413_reg/NET0131 , \g1414_reg/NET0131 , \g1415_reg/NET0131 , \g1416_reg/NET0131 , \g1417_reg/NET0131 , \g1418_reg/NET0131 , \g1419_reg/NET0131 , \g141_reg/NET0131 , \g1420_reg/NET0131 , \g1421_reg/NET0131 , \g1422_reg/NET0131 , \g1423_reg/NET0131 , \g1424_reg/NET0131 , \g1425_reg/NET0131 , \g1426_reg/NET0131 , \g142_reg/NET0131 , \g1430_reg/NET0131 , \g1435_reg/NET0131 , \g1439_reg/NET0131 , \g143_reg/NET0131 , \g1444_reg/NET0131 , \g1448_reg/NET0131 , \g144_reg/NET0131 , \g1453_reg/NET0131 , \g1457_reg/NET0131 , \g145_reg/NET0131 , \g1462_reg/NET0131 , \g1466_reg/NET0131 , \g146_reg/NET0131 , \g1471_reg/NET0131 , \g1476_reg/NET0131 , \g147_reg/NET0131 , \g1481_reg/NET0131 , \g1486_reg/NET0131 , \g148_reg/NET0131 , \g1491_reg/NET0131 , \g1496_reg/NET0131 , \g149_reg/NET0131 , \g1501_reg/NET0131 , \g1506_reg/NET0131 , \g150_reg/NET0131 , \g1511_reg/NET0131 , \g1512_reg/NET0131 , \g1513_reg/NET0131 , \g1514_reg/NET0131 , \g1515_reg/NET0131 , \g1516_reg/NET0131 , \g151_reg/NET0131 , \g1523_reg/NET0131 , \g1524_reg/NET0131 , \g1525_reg/NET0131 , \g1526_reg/NET0131 , \g1527_reg/NET0131 , \g1528_reg/NET0131 , \g1529_reg/NET0131 , \g152_reg/NET0131 , \g1530_reg/NET0131 , \g1531_reg/NET0131 , \g1532_reg/NET0131 , \g1533_reg/NET0131 , \g1534_reg/NET0131 , \g1535_reg/NET0131 , \g1536_reg/NET0131 , \g1537_reg/NET0131 , \g1538_reg/NET0131 , \g1539_reg/NET0131 , \g153_reg/NET0131 , \g1540_reg/NET0131 , \g1541_reg/NET0131 , \g1542_reg/NET0131 , \g1543_reg/NET0131 , \g1544_reg/NET0131 , \g1545_reg/NET0131 , \g1546_reg/NET0131 , \g154_reg/NET0131 , \g1550_reg/NET0131 , \g1551_reg/NET0131 , \g1552_reg/NET0131 , \g1553_reg/NET0131 , \g1554_reg/NET0131 , \g1555_reg/NET0131 , \g1556_reg/NET0131 , \g1557_reg/NET0131 , \g1558_reg/NET0131 , \g1559_reg/NET0131 , \g155_reg/NET0131 , \g1560_reg/NET0131 , \g1561_reg/NET0131 , \g1563_reg/NET0131 , \g1567_reg/NET0131 , \g156_reg/NET0131 , \g1570_reg/NET0131 , \g1573_reg/NET0131 , \g1576_reg/NET0131 , \g1579_reg/NET0131 , \g157_reg/NET0131 , \g1582_reg/NET0131 , \g1585_reg/NET0131 , \g1588_reg/NET0131 , \g158_reg/NET0131 , \g1591_reg/NET0131 , \g1594_reg/NET0131 , \g1597_reg/NET0131 , \g159_reg/NET0131 , \g1600_reg/NET0131 , \g1603_reg/NET0131 , \g1606_reg/NET0131 , \g1609_reg/NET0131 , \g160_reg/NET0131 , \g1612_reg/NET0131 , \g1615_reg/NET0131 , \g1618_reg/NET0131 , \g161_reg/NET0131 , \g1621_reg/NET0131 , \g1624_reg/NET0131 , \g1627_reg/NET0131 , \g16297_pad , \g162_reg/NET0131 , \g1630_reg/NET0131 , \g1633_reg/NET0131 , \g16355_pad , \g1636_reg/NET0131 , \g16399_pad , \g1639_reg/NET0131 , \g163_reg/NET0131 , \g1642_reg/NET0131 , \g16437_pad , \g1645_reg/NET0131 , \g1648_reg/NET0131 , \g164_reg/NET0131 , \g1651_reg/NET0131 , \g1654_reg/NET0131 , \g1660_reg/NET0131 , \g1662_reg/NET0131 , \g1664_reg/NET0131 , \g1666_reg/NET0131 , \g1668_reg/NET0131 , \g1670_reg/NET0131 , \g1672_reg/NET0131 , \g1679_reg/NET0131 , \g1680_reg/NET0131 , \g1686_reg/NET0131 , \g168_reg/NET0131 , \g1693_reg/NET0131 , \g1694_reg/NET0131 , \g1695_reg/NET0131 , \g1696_reg/NET0131 , \g1697_reg/NET0131 , \g1698_reg/NET0131 , \g1699_reg/NET0131 , \g169_reg/NET0131 , \g1700_reg/NET0131 , \g1701_reg/NET0131 , \g1702_reg/NET0131 , \g1703_reg/NET0131 , \g1704_reg/NET0131 , \g1705_reg/NET0131 , \g170_reg/NET0131 , \g171_reg/NET0131 , \g1724_reg/NET0131 , \g1727_reg/NET0131 , \g172_reg/NET0131 , \g1730_reg/NET0131 , \g1732_reg/NET0131 , \g1734_reg/NET0131 , \g1735_reg/NET0131 , \g1739_reg/NET0131 , \g173_reg/NET0131 , \g1742_reg/NET0131 , \g1745_reg/NET0131 , \g1747_reg/NET0131 , \g1749_reg/NET0131 , \g174_reg/NET0131 , \g1750_reg/NET0131 , \g1754_reg/NET0131 , \g1757_reg/NET0131 , \g175_reg/NET0131 , \g1760_reg/NET0131 , \g1762_reg/NET0131 , \g1764_reg/NET0131 , \g1765_reg/NET0131 , \g1769_reg/NET0131 , \g176_reg/NET0131 , \g1772_reg/NET0131 , \g1775_reg/NET0131 , \g1777_reg/NET0131 , \g1779_reg/NET0131 , \g177_reg/NET0131 , \g1783_reg/NET0131 , \g1784_reg/NET0131 , \g1785_reg/NET0131 , \g1789_reg/NET0131 , \g178_reg/NET0131 , \g1792_reg/NET0131 , \g1795_reg/NET0131 , \g1798_reg/NET0131 , \g179_reg/NET0131 , \g1801_reg/NET0131 , \g1804_reg/NET0131 , \g1807_reg/NET0131 , \g1808_reg/NET0131 , \g1809_reg/NET0131 , \g1810_reg/NET0131 , \g1813_reg/NET0131 , \g1816_reg/NET0131 , \g1819_reg/NET0131 , \g1822_reg/NET0131 , \g1825_reg/NET0131 , \g1828_reg/NET0131 , \g1829_reg/NET0131 , \g1830_reg/NET0131 , \g1832_reg/NET0131 , \g1834_reg/NET0131 , \g1845_reg/NET0131 , \g1846_reg/NET0131 , \g1849_reg/NET0131 , \g1852_reg/NET0131 , \g1858_reg/NET0131 , \g1859_reg/NET0131 , \g185_reg/NET0131 , \g1860_reg/NET0131 , \g1861_reg/NET0131 , \g1865_reg/NET0131 , \g1867_reg/NET0131 , \g1868_reg/NET0131 , \g1869_reg/NET0131 , \g186_reg/NET0131 , \g1870_reg/NET0131 , \g1871_reg/NET0131 , \g1874_reg/NET0131 , \g1877_reg/NET0131 , \g1880_reg/NET0131 , \g1886_reg/NET0131 , \g1887_reg/NET0131 , \g189_reg/NET0131 , \g1904_reg/NET0131 , \g1905_reg/NET0131 , \g1909_reg/NET0131 , \g1910_reg/NET0131 , \g1911_reg/NET0131 , \g1912_reg/NET0131 , \g1913_reg/NET0131 , \g1914_reg/NET0131 , \g1916_reg/NET0131 , \g1917_reg/NET0131 , \g1918_reg/NET0131 , \g1921_reg/NET0131 , \g1922_reg/NET0131 , \g1924_reg/NET0131 , \g1928_reg/NET0131 , \g192_reg/NET0131 , \g1939_reg/NET0131 , \g1943_pad , \g1945_reg/NET0131 , \g1947_reg/NET0131 , \g1949_reg/NET0131 , \g1951_reg/NET0131 , \g1953_reg/NET0131 , \g1955_reg/NET0131 , \g1956_reg/NET0131 , \g1957_reg/NET0131 , \g1958_reg/NET0131 , \g1959_reg/NET0131 , \g195_reg/NET0131 , \g1960_reg/NET0131 , \g1961_reg/NET0131 , \g1962_reg/NET0131 , \g1963_reg/NET0131 , \g1964_reg/NET0131 , \g1965_reg/NET0131 , \g1966_reg/NET0131 , \g1967_reg/NET0131 , \g1970_reg/NET0131 , \g1973_reg/NET0131 , \g1976_reg/NET0131 , \g1979_reg/NET0131 , \g1982_reg/NET0131 , \g1985_reg/NET0131 , \g1988_reg/NET0131 , \g198_reg/NET0131 , \g1991_reg/NET0131 , \g1994_reg/NET0131 , \g1997_reg/NET0131 , \g2000_reg/NET0131 , \g201_reg/NET0131 , \g204_reg/NET0131 , \g2078_reg/NET0131 , \g2079_reg/NET0131 , \g207_reg/NET0131 , \g2080_reg/NET0131 , \g2081_reg/NET0131 , \g2082_reg/NET0131 , \g2083_reg/NET0131 , \g2084_reg/NET0131 , \g2085_reg/NET0131 , \g2086_reg/NET0131 , \g2087_reg/NET0131 , \g2088_reg/NET0131 , \g2089_reg/NET0131 , \g2090_reg/NET0131 , \g2091_reg/NET0131 , \g2092_reg/NET0131 , \g2093_reg/NET0131 , \g2094_reg/NET0131 , \g2095_reg/NET0131 , \g2096_reg/NET0131 , \g2097_reg/NET0131 , \g2098_reg/NET0131 , \g2099_reg/NET0131 , \g2100_reg/NET0131 , \g2101_reg/NET0131 , \g2102_reg/NET0131 , \g2103_reg/NET0131 , \g2104_reg/NET0131 , \g2105_reg/NET0131 , \g2106_reg/NET0131 , \g2107_reg/NET0131 , \g2108_reg/NET0131 , \g2109_reg/NET0131 , \g210_reg/NET0131 , \g2110_reg/NET0131 , \g2111_reg/NET0131 , \g2112_reg/NET0131 , \g2113_reg/NET0131 , \g2114_reg/NET0131 , \g2115_reg/NET0131 , \g2116_reg/NET0131 , \g2117_reg/NET0131 , \g2118_reg/NET0131 , \g2119_reg/NET0131 , \g213_reg/NET0131 , \g2165_reg/NET0131 , \g216_reg/NET0131 , \g2170_reg/NET0131 , \g2175_reg/NET0131 , \g2180_reg/NET0131 , \g2185_reg/NET0131 , \g2190_reg/NET0131 , \g2195_reg/NET0131 , \g219_reg/NET0131 , \g2200_reg/NET0131 , \g2205_reg/NET0131 , \g2206_reg/NET0131 , \g2207_reg/NET0131 , \g2208_reg/NET0131 , \g2209_reg/NET0131 , \g2210_reg/NET0131 , \g2217_reg/NET0131 , \g2218_reg/NET0131 , \g2219_reg/NET0131 , \g2220_reg/NET0131 , \g2221_reg/NET0131 , \g2222_reg/NET0131 , \g2223_reg/NET0131 , \g2224_reg/NET0131 , \g2225_reg/NET0131 , \g2226_reg/NET0131 , \g2227_reg/NET0131 , \g2228_reg/NET0131 , \g2229_reg/NET0131 , \g222_reg/NET0131 , \g2230_reg/NET0131 , \g2231_reg/NET0131 , \g2232_reg/NET0131 , \g2233_reg/NET0131 , \g2234_reg/NET0131 , \g2235_reg/NET0131 , \g2236_reg/NET0131 , \g2237_reg/NET0131 , \g2238_reg/NET0131 , \g2239_reg/NET0131 , \g2240_reg/NET0131 , \g2244_reg/NET0131 , \g2245_reg/NET0131 , \g2246_reg/NET0131 , \g2247_reg/NET0131 , \g2248_reg/NET0131 , \g2249_reg/NET0131 , \g2250_reg/NET0131 , \g2251_reg/NET0131 , \g2252_reg/NET0131 , \g2253_reg/NET0131 , \g2254_reg/NET0131 , \g2255_reg/NET0131 , \g225_reg/NET0131 , \g2261_reg/NET0131 , \g2264_reg/NET0131 , \g2267_reg/NET0131 , \g2270_reg/NET0131 , \g2273_reg/NET0131 , \g2276_reg/NET0131 , \g2279_reg/NET0131 , \g2282_reg/NET0131 , \g2285_reg/NET0131 , \g2288_reg/NET0131 , \g228_reg/NET0131 , \g2291_reg/NET0131 , \g2294_reg/NET0131 , \g2297_reg/NET0131 , \g2300_reg/NET0131 , \g2303_reg/NET0131 , \g2306_reg/NET0131 , \g2309_reg/NET0131 , \g2312_reg/NET0131 , \g2315_reg/NET0131 , \g2318_reg/NET0131 , \g231_reg/NET0131 , \g2321_reg/NET0131 , \g2324_reg/NET0131 , \g2327_reg/NET0131 , \g2330_reg/NET0131 , \g2333_reg/NET0131 , \g2336_reg/NET0131 , \g2339_reg/NET0131 , \g2342_reg/NET0131 , \g2345_reg/NET0131 , \g2348_reg/NET0131 , \g234_reg/NET0131 , \g2354_reg/NET0131 , \g2356_reg/NET0131 , \g2358_reg/NET0131 , \g2360_reg/NET0131 , \g2362_reg/NET0131 , \g2364_reg/NET0131 , \g2366_reg/NET0131 , \g2373_reg/NET0131 , \g2374_reg/NET0131 , \g237_reg/NET0131 , \g2380_reg/NET0131 , \g2387_reg/NET0131 , \g2388_reg/NET0131 , \g2389_reg/NET0131 , \g2390_reg/NET0131 , \g2391_reg/NET0131 , \g2392_reg/NET0131 , \g2393_reg/NET0131 , \g2394_reg/NET0131 , \g2395_reg/NET0131 , \g2396_reg/NET0131 , \g2397_reg/NET0131 , \g2398_reg/NET0131 , \g2399_reg/NET0131 , \g240_reg/NET0131 , \g2418_reg/NET0131 , \g2421_reg/NET0131 , \g2424_reg/NET0131 , \g2426_reg/NET0131 , \g2428_reg/NET0131 , \g2429_reg/NET0131 , \g2433_reg/NET0131 , \g2436_reg/NET0131 , \g2439_reg/NET0131 , \g243_reg/NET0131 , \g2441_reg/NET0131 , \g2443_reg/NET0131 , \g2444_reg/NET0131 , \g2448_reg/NET0131 , \g2451_reg/NET0131 , \g2454_reg/NET0131 , \g2456_reg/NET0131 , \g2458_reg/NET0131 , \g2459_reg/NET0131 , \g2463_reg/NET0131 , \g2466_reg/NET0131 , \g2469_reg/NET0131 , \g246_reg/NET0131 , \g2471_reg/NET0131 , \g2473_reg/NET0131 , \g2477_reg/NET0131 , \g2478_reg/NET0131 , \g2479_reg/NET0131 , \g2483_reg/NET0131 , \g2486_reg/NET0131 , \g2489_reg/NET0131 , \g2492_reg/NET0131 , \g2495_reg/NET0131 , \g2498_reg/NET0131 , \g249_reg/NET0131 , \g2501_reg/NET0131 , \g2502_reg/NET0131 , \g2503_reg/NET0131 , \g2504_reg/NET0131 , \g2507_reg/NET0131 , \g2510_reg/NET0131 , \g2513_reg/NET0131 , \g2516_reg/NET0131 , \g2519_reg/NET0131 , \g2522_reg/NET0131 , \g2523_reg/NET0131 , \g2524_reg/NET0131 , \g2526_reg/NET0131 , \g2528_reg/NET0131 , \g252_reg/NET0131 , \g2539_reg/NET0131 , \g2540_reg/NET0131 , \g2543_reg/NET0131 , \g2546_reg/NET0131 , \g2552_reg/NET0131 , \g2553_reg/NET0131 , \g2554_reg/NET0131 , \g2555_reg/NET0131 , \g2559_reg/NET0131 , \g255_reg/NET0131 , \g2561_reg/NET0131 , \g2562_reg/NET0131 , \g2563_reg/NET0131 , \g2564_reg/NET0131 , \g2565_reg/NET0131 , \g2568_reg/NET0131 , \g2571_reg/NET0131 , \g2574_reg/NET0131 , \g2580_reg/NET0131 , \g2581_reg/NET0131 , \g258_reg/NET0131 , \g2598_reg/NET0131 , \g2599_reg/NET0131 , \g2603_reg/NET0131 , \g2604_reg/NET0131 , \g2605_reg/NET0131 , \g2606_reg/NET0131 , \g2607_reg/NET0131 , \g2608_reg/NET0131 , \g2610_reg/NET0131 , \g2611_reg/NET0131 , \g2612_reg/NET0131 , \g2615_reg/NET0131 , \g2616_reg/NET0131 , \g2618_reg/NET0131 , \g261_reg/NET0131 , \g2622_reg/NET0131 , \g2633_reg/NET0131 , \g2637_pad , \g2639_reg/NET0131 , \g2641_reg/NET0131 , \g2643_reg/NET0131 , \g2645_reg/NET0131 , \g2647_reg/NET0131 , \g2649_reg/NET0131 , \g264_reg/NET0131 , \g2650_reg/NET0131 , \g2651_reg/NET0131 , \g2652_reg/NET0131 , \g2653_reg/NET0131 , \g2654_reg/NET0131 , \g2655_reg/NET0131 , \g2656_reg/NET0131 , \g2657_reg/NET0131 , \g2658_reg/NET0131 , \g2659_reg/NET0131 , \g2660_reg/NET0131 , \g2661_reg/NET0131 , \g2664_reg/NET0131 , \g2667_reg/NET0131 , \g2670_reg/NET0131 , \g2673_reg/NET0131 , \g2676_reg/NET0131 , \g2679_reg/NET0131 , \g267_reg/NET0131 , \g2682_reg/NET0131 , \g2685_reg/NET0131 , \g2688_reg/NET0131 , \g2691_reg/NET0131 , \g2694_reg/NET0131 , \g270_reg/NET0131 , \g273_reg/NET0131 , \g2772_reg/NET0131 , \g2773_reg/NET0131 , \g2774_reg/NET0131 , \g2775_reg/NET0131 , \g2776_reg/NET0131 , \g2777_reg/NET0131 , \g2778_reg/NET0131 , \g2779_reg/NET0131 , \g2780_reg/NET0131 , \g2781_reg/NET0131 , \g2782_reg/NET0131 , \g2783_reg/NET0131 , \g2784_reg/NET0131 , \g2785_reg/NET0131 , \g2786_reg/NET0131 , \g2787_reg/NET0131 , \g2788_reg/NET0131 , \g2789_reg/NET0131 , \g2790_reg/NET0131 , \g2791_reg/NET0131 , \g2792_reg/NET0131 , \g2793_reg/NET0131 , \g2794_reg/NET0131 , \g2795_reg/NET0131 , \g2796_reg/NET0131 , \g2797_reg/NET0131 , \g2798_reg/NET0131 , \g2799_reg/NET0131 , \g279_reg/NET0131 , \g2800_reg/NET0131 , \g2801_reg/NET0131 , \g2802_reg/NET0131 , \g2803_reg/NET0131 , \g2804_reg/NET0131 , \g2805_reg/NET0131 , \g2806_reg/NET0131 , \g2807_reg/NET0131 , \g2808_reg/NET0131 , \g2809_reg/NET0131 , \g2810_reg/NET0131 , \g2811_reg/NET0131 , \g2812_reg/NET0131 , \g2813_reg/NET0131 , \g2814_reg/NET0131 , \g2817_reg/NET0131 , \g281_reg/NET0131 , \g283_reg/NET0131 , \g285_reg/NET0131 , \g2874_reg/NET0131 , \g2879_reg/NET0131 , \g287_reg/NET0131 , \g2883_reg/NET0131 , \g2888_reg/NET0131 , \g2892_reg/NET0131 , \g2896_reg/NET0131 , \g289_reg/NET0131 , \g2900_reg/NET0131 , \g2903_reg/NET0131 , \g2908_reg/NET0131 , \g2912_reg/NET0131 , \g2917_reg/NET0131 , \g291_reg/NET0131 , \g2920_reg/NET0131 , \g2924_reg/NET0131 , \g2929_reg/NET0131 , \g2933_reg/NET0131 , \g2934_reg/NET0131 , \g2935_reg/NET0131 , \g2938_reg/NET0131 , \g2941_reg/NET0131 , \g2944_reg/NET0131 , \g2947_reg/NET0131 , \g2950_reg/NET0131 , \g2953_reg/NET0131 , \g2956_reg/NET0131 , \g2959_reg/NET0131 , \g2962_reg/NET0131 , \g2963_reg/NET0131 , \g2966_reg/NET0131 , \g2969_reg/NET0131 , \g2972_reg/NET0131 , \g2975_reg/NET0131 , \g2978_reg/NET0131 , \g2981_reg/NET0131 , \g2984_reg/NET0131 , \g2985_reg/NET0131 , \g2986_reg/NET0131 , \g2987_reg/NET0131 , \g298_reg/NET0131 , \g2990_reg/NET0131 , \g2991_reg/NET0131 , \g2992_reg/NET0131 , \g2993_reg/NET0131 , \g2997_reg/NET0131 , \g2998_reg/NET0131 , \g299_reg/NET0131 , \g3002_reg/NET0131 , \g3006_reg/NET0131 , \g3010_reg/NET0131 , \g3013_reg/NET0131 , \g3018_reg/NET0131 , \g3024_reg/NET0131 , \g3028_reg/NET0131 , \g3032_reg/NET0131 , \g3036_reg/NET0131 , \g3043_reg/NET0131 , \g3044_reg/NET0131 , \g3045_reg/NET0131 , \g3046_reg/NET0131 , \g3047_reg/NET0131 , \g3048_reg/NET0131 , \g3049_reg/NET0131 , \g3050_reg/NET0131 , \g3051_reg/NET0131 , \g3052_reg/NET0131 , \g3053_reg/NET0131 , \g3054_reg/NET0131 , \g3055_reg/NET0131 , \g3056_reg/NET0131 , \g3057_reg/NET0131 , \g3058_reg/NET0131 , \g3059_reg/NET0131 , \g305_reg/NET0131 , \g3060_reg/NET0131 , \g3061_reg/NET0131 , \g3062_reg/NET0131 , \g3063_reg/NET0131 , \g3064_reg/NET0131 , \g3065_reg/NET0131 , \g3066_reg/NET0131 , \g3067_reg/NET0131 , \g3068_reg/NET0131 , \g3069_reg/NET0131 , \g3070_reg/NET0131 , \g3071_reg/NET0131 , \g3072_reg/NET0131 , \g3073_reg/NET0131 , \g3074_reg/NET0131 , \g3075_reg/NET0131 , \g3076_reg/NET0131 , \g3077_reg/NET0131 , \g3078_reg/NET0131 , \g3079_reg/NET0131 , \g3080_reg/NET0131 , \g3083_reg/NET0131 , \g3097_reg/NET0131 , \g3110_reg/NET0131 , \g3114_reg/NET0131 , \g3120_reg/NET0131 , \g312_reg/NET0131 , \g3139_reg/NET0131 , \g313_reg/NET0131 , \g314_reg/NET0131 , \g315_reg/NET0131 , \g316_reg/NET0131 , \g317_reg/NET0131 , \g318_reg/NET0131 , \g319_reg/NET0131 , \g320_reg/NET0131 , \g321_reg/NET0131 , \g3229_pad , \g322_reg/NET0131 , \g3230_pad , \g3231_pad , \g3233_pad , \g3234_pad , \g323_reg/NET0131 , \g324_reg/NET0131 , \g343_reg/NET0131 , \g346_reg/NET0131 , \g349_reg/NET0131 , \g351_reg/NET0131 , \g353_reg/NET0131 , \g354_reg/NET0131 , \g358_reg/NET0131 , \g361_reg/NET0131 , \g364_reg/NET0131 , \g366_reg/NET0131 , \g368_reg/NET0131 , \g369_reg/NET0131 , \g373_reg/NET0131 , \g376_reg/NET0131 , \g379_reg/NET0131 , \g381_reg/NET0131 , \g383_reg/NET0131 , \g384_reg/NET0131 , \g388_reg/NET0131 , \g391_reg/NET0131 , \g394_reg/NET0131 , \g396_reg/NET0131 , \g398_reg/NET0131 , \g402_reg/NET0131 , \g403_reg/NET0131 , \g404_reg/NET0131 , \g408_reg/NET0131 , \g411_reg/NET0131 , \g414_reg/NET0131 , \g417_reg/NET0131 , \g420_reg/NET0131 , \g423_reg/NET0131 , \g426_reg/NET0131 , \g427_reg/NET0131 , \g428_reg/NET0131 , \g429_reg/NET0131 , \g432_reg/NET0131 , \g435_reg/NET0131 , \g438_reg/NET0131 , \g441_reg/NET0131 , \g444_reg/NET0131 , \g447_reg/NET0131 , \g448_reg/NET0131 , \g449_reg/NET0131 , \g451_reg/NET0131 , \g453_reg/NET0131 , \g464_reg/NET0131 , \g465_reg/NET0131 , \g468_reg/NET0131 , \g471_reg/NET0131 , \g477_reg/NET0131 , \g478_reg/NET0131 , \g479_reg/NET0131 , \g480_reg/NET0131 , \g484_reg/NET0131 , \g486_reg/NET0131 , \g487_reg/NET0131 , \g488_reg/NET0131 , \g489_reg/NET0131 , \g490_reg/NET0131 , \g493_reg/NET0131 , \g496_reg/NET0131 , \g499_reg/NET0131 , \g506_reg/NET0131 , \g507_reg/NET0131 , \g51_pad , \g524_reg/NET0131 , \g525_reg/NET0131 , \g529_reg/NET0131 , \g530_reg/NET0131 , \g531_reg/NET0131 , \g532_reg/NET0131 , \g533_reg/NET0131 , \g534_reg/NET0131 , \g536_reg/NET0131 , \g537_reg/NET0131 , \g5388_pad , \g538_reg/NET0131 , \g541_reg/NET0131 , \g542_reg/NET0131 , \g544_reg/NET0131 , \g548_reg/NET0131 , \g559_reg/NET0131 , \g563_pad , \g5657_pad , \g565_reg/NET0131 , \g567_reg/NET0131 , \g569_reg/NET0131 , \g571_reg/NET0131 , \g573_reg/NET0131 , \g575_reg/NET0131 , \g576_reg/NET0131 , \g577_reg/NET0131 , \g578_reg/NET0131 , \g579_reg/NET0131 , \g580_reg/NET0131 , \g581_reg/NET0131 , \g582_reg/NET0131 , \g583_reg/NET0131 , \g584_reg/NET0131 , \g585_reg/NET0131 , \g586_reg/NET0131 , \g587_reg/NET0131 , \g590_reg/NET0131 , \g593_reg/NET0131 , \g596_reg/NET0131 , \g599_reg/NET0131 , \g602_reg/NET0131 , \g605_reg/NET0131 , \g608_reg/NET0131 , \g611_reg/NET0131 , \g614_reg/NET0131 , \g617_reg/NET0131 , \g620_reg/NET0131 , \g698_reg/NET0131 , \g699_reg/NET0131 , \g700_reg/NET0131 , \g701_reg/NET0131 , \g702_reg/NET0131 , \g703_reg/NET0131 , \g704_reg/NET0131 , \g705_reg/NET0131 , \g706_reg/NET0131 , \g707_reg/NET0131 , \g708_reg/NET0131 , \g709_reg/NET0131 , \g710_reg/NET0131 , \g711_reg/NET0131 , \g712_reg/NET0131 , \g713_reg/NET0131 , \g714_reg/NET0131 , \g715_reg/NET0131 , \g716_reg/NET0131 , \g717_reg/NET0131 , \g718_reg/NET0131 , \g719_reg/NET0131 , \g720_reg/NET0131 , \g721_reg/NET0131 , \g722_reg/NET0131 , \g723_reg/NET0131 , \g724_reg/NET0131 , \g725_reg/NET0131 , \g726_reg/NET0131 , \g727_reg/NET0131 , \g728_reg/NET0131 , \g729_reg/NET0131 , \g730_reg/NET0131 , \g731_reg/NET0131 , \g732_reg/NET0131 , \g733_reg/NET0131 , \g734_reg/NET0131 , \g735_reg/NET0131 , \g736_reg/NET0131 , \g737_reg/NET0131 , \g738_reg/NET0131 , \g739_reg/NET0131 , \g785_reg/NET0131 , \g789_reg/NET0131 , \g793_reg/NET0131 , \g7961_pad , \g797_reg/NET0131 , \g801_reg/NET0131 , \g805_reg/NET0131 , \g809_reg/NET0131 , \g813_reg/NET0131 , \g817_reg/NET0131 , \g818_reg/NET0131 , \g819_reg/NET0131 , \g820_reg/NET0131 , \g821_reg/NET0131 , \g822_reg/NET0131 , \g8259_pad , \g8260_pad , \g8261_pad , \g8262_pad , \g8263_pad , \g8264_pad , \g8265_pad , \g8266_pad , \g8268_pad , \g8269_pad , \g8270_pad , \g8271_pad , \g8272_pad , \g8273_pad , \g8274_pad , \g8275_pad , \g829_reg/NET0131 , \g830_reg/NET0131 , \g831_reg/NET0131 , \g832_reg/NET0131 , \g833_reg/NET0131 , \g834_reg/NET0131 , \g835_reg/NET0131 , \g836_reg/NET0131 , \g837_reg/NET0131 , \g838_reg/NET0131 , \g839_reg/NET0131 , \g840_reg/NET0131 , \g841_reg/NET0131 , \g842_reg/NET0131 , \g843_reg/NET0131 , \g844_reg/NET0131 , \g845_reg/NET0131 , \g846_reg/NET0131 , \g847_reg/NET0131 , \g848_reg/NET0131 , \g849_reg/NET0131 , \g850_reg/NET0131 , \g851_reg/NET0131 , \g852_reg/NET0131 , \g856_reg/NET0131 , \g857_reg/NET0131 , \g858_reg/NET0131 , \g859_reg/NET0131 , \g860_reg/NET0131 , \g861_reg/NET0131 , \g862_reg/NET0131 , \g863_reg/NET0131 , \g864_reg/NET0131 , \g865_reg/NET0131 , \g866_reg/NET0131 , \g867_reg/NET0131 , \g873_reg/NET0131 , \g876_reg/NET0131 , \g879_reg/NET0131 , \g882_reg/NET0131 , \g885_reg/NET0131 , \g888_reg/NET0131 , \g891_reg/NET0131 , \g894_reg/NET0131 , \g897_reg/NET0131 , \g900_reg/NET0131 , \g903_reg/NET0131 , \g906_reg/NET0131 , \g909_reg/NET0131 , \g912_reg/NET0131 , \g915_reg/NET0131 , \g918_reg/NET0131 , \g921_reg/NET0131 , \g924_reg/NET0131 , \g927_reg/NET0131 , \g930_reg/NET0131 , \g933_reg/NET0131 , \g936_reg/NET0131 , \g939_reg/NET0131 , \g942_reg/NET0131 , \g945_reg/NET0131 , \g948_reg/NET0131 , \g951_reg/NET0131 , \g954_reg/NET0131 , \g957_reg/NET0131 , \g960_reg/NET0131 , \g966_reg/NET0131 , \g968_reg/NET0131 , \g970_reg/NET0131 , \g972_reg/NET0131 , \g974_reg/NET0131 , \g976_reg/NET0131 , \g978_reg/NET0131 , \g97_reg/NET0131 , \g985_reg/NET0131 , \g986_reg/NET0131 , \g992_reg/NET0131 , \g999_reg/NET0131 , \_al_n0 , \_al_n1 , \g101_reg/P0001 , \g105_reg/P0001 , \g109_reg/P0001 , \g1138_reg/P0001 , \g113_reg/P0001 , \g1140_reg/P0001 , \g117_reg/P0001 , \g121_reg/P0001 , \g125_reg/P0001 , \g1471_reg/P0001 , \g1476_reg/P0001 , \g1481_reg/P0001 , \g1486_reg/P0001 , \g1491_reg/P0001 , \g1496_reg/P0001 , \g1501_reg/P0001 , \g1506_reg/P0001 , \g16496_pad , \g1660_reg/P0001 , \g1662_reg/P0001 , \g1664_reg/P0001 , \g1666_reg/P0001 , \g1668_reg/P0001 , \g1670_reg/P0001 , \g1672_reg/P0001 , \g18/_0_ , \g1832_reg/P0001 , \g1834_reg/P0001 , \g2165_reg/P0001 , \g2170_reg/P0001 , \g2175_reg/P0001 , \g2180_reg/P0001 , \g2185_reg/P0001 , \g2190_reg/P0001 , \g2195_reg/P0001 , \g2200_reg/P0001 , \g2354_reg/P0001 , \g2356_reg/P0001 , \g2358_reg/P0001 , \g2360_reg/P0001 , \g2362_reg/P0001 , \g2364_reg/P0001 , \g2366_reg/P0001 , \g2526_reg/P0001 , \g2528_reg/P0001 , \g25489_pad , \g279_reg/P0001 , \g281_reg/P0001 , \g283_reg/P0001 , \g285_reg/P0001 , \g2879_reg/NET0131_syn_2 , \g287_reg/P0001 , \g289_reg/P0001 , \g291_reg/P0001 , \g451_reg/P0001 , \g453_reg/P0001 , \g59421/_3_ , \g59425/_1_ , \g59435/_0_ , \g59436/_0_ , \g59441/_3_ , \g59442/_0_ , \g59445/_0_ , \g59453/_0_ , \g59462/_3_ , \g59466/_3_ , \g59467/_3_ , \g59468/_3_ , \g59469/_3_ , \g59470/_3_ , \g59471/_3_ , \g59472/_3_ , \g59473/_3_ , \g59489/_0_ , \g59498/_0_ , \g59499/_0_ , \g59500/_0_ , \g59502/_2_ , \g59503/_0_ , \g59505/_2_ , \g59507/_0_ , \g59508/_0_ , \g59533/_3_ , \g59534/_3_ , \g59535/_3_ , \g59536/_3_ , \g59537/_3_ , \g59538/_3_ , \g59539/_3_ , \g59540/_3_ , \g59548/_0_ , \g59550/_0_ , \g59551/_0_ , \g59552/_0_ , \g59554/_0_ , \g59555/_0_ , \g59556/_0_ , \g59557/_0_ , \g59558/_0_ , \g59559/_0_ , \g59560/_0_ , \g59561/_0_ , \g59639/_0_ , \g59694/_2_ , \g59695/_0_ , \g59697/_2_ , \g59698/_0_ , \g59699/_0_ , \g59700/_0_ , \g59705/_0_ , \g59706/_0_ , \g59707/_0_ , \g59708/_0_ , \g59709/_0_ , \g59710/_0_ , \g59711/_0_ , \g59712/_0_ , \g59713/_0_ , \g59714/_0_ , \g59715/_0_ , \g59716/_0_ , \g59717/_0_ , \g59718/_0_ , \g59719/_0_ , \g59720/_0_ , \g59721/_0_ , \g59722/_0_ , \g59723/_0_ , \g59724/_0_ , \g59725/_0_ , \g59726/_0_ , \g59727/_0_ , \g59728/_0_ , \g59729/_0_ , \g59730/_0_ , \g59731/_0_ , \g59732/_0_ , \g59733/_0_ , \g59734/_0_ , \g59735/_0_ , \g59736/_0_ , \g59737/_0_ , \g59738/_0_ , \g59739/_0_ , \g59740/_0_ , \g59741/_0_ , \g59742/_0_ , \g59743/_0_ , \g59744/_0_ , \g59745/_0_ , \g59747/_0_ , \g59748/_0_ , \g59749/_0_ , \g59750/_0_ , \g59751/_0_ , \g59752/_0_ , \g59753/_0_ , \g59754/_0_ , \g59755/_0_ , \g59756/_0_ , \g59757/_0_ , \g59758/_0_ , \g59759/_0_ , \g59760/_0_ , \g59761/_0_ , \g59762/_0_ , \g59763/_0_ , \g59764/_0_ , \g59765/_0_ , \g59766/_0_ , \g59915/_0_ , \g59952/_2_ , \g60046/_0_ , \g60048/_0_ , \g60049/_0_ , \g60051/_0_ , \g60063/_0_ , \g60103/_0_ , \g60104/_0_ , \g60105/_0_ , \g60107/_2_ , \g60108/_0_ , \g60109/_0_ , \g60110/_0_ , \g60112/_2_ , \g60119/_0_ , \g60120/_0_ , \g60121/_0_ , \g60122/_0_ , \g60123/_0_ , \g60124/_0_ , \g60126/_0_ , \g60127/_0_ , \g60128/_0_ , \g60129/_0_ , \g60130/_0_ , \g60135/_0_ , \g60136/_0_ , \g60137/_0_ , \g60138/_0_ , \g60139/_0_ , \g60143/_3_ , \g60144/_0_ , \g60145/_0_ , \g60339/_0_ , \g60404/_0_ , \g60427/_0_ , \g60428/_0_ , \g60429/_0_ , \g60434/_0_ , \g60435/_0_ , \g60437/_0_ , \g60438/_0_ , \g60439/_0_ , \g60440/_0_ , \g60441/_0_ , \g60448/_0_ , \g60451/_0_ , \g60452/_0_ , \g60453/_0_ , \g60459/_0_ , \g60460/_0_ , \g60523/_0_ , \g60534/_0_ , \g60535/_0_ , \g60536/_0_ , \g60585/_0_ , \g60586/_0_ , \g60587/_0_ , \g60588/_0_ , \g60591/_0_ , \g60592/_0_ , \g60599/_0_ , \g60601/_0_ , \g60602/_0_ , \g60603/_0_ , \g60604/_0_ , \g60605/_0_ , \g60606/_0_ , \g60607/_0_ , \g60608/_0_ , \g60609/_0_ , \g60613/_0_ , \g60614/_0_ , \g60615/_0_ , \g60694/_0_ , \g60708/_0_ , \g60709/_0_ , \g60710/_0_ , \g60785/_0_ , \g60787/_0_ , \g60788/_0_ , \g60799/_0_ , \g60801/_0_ , \g60802/_0_ , \g60803/_1__syn_2 , \g60805/_1__syn_2 , \g60806/_1__syn_2 , \g60808/_0_ , \g60810/_0_ , \g60811/_0_ , \g60825/_3_ , \g60896/_0_ , \g60980/_0_ , \g60981/_0_ , \g60985/_0_ , \g60986/_0_ , \g61012/_0_ , \g61013/_0_ , \g61015/_0_ , \g61017/_0_ , \g61122/_0_ , \g61123/_0_ , \g61124/_0_ , \g61125/_0_ , \g61222/_0_ , \g61223/_0_ , \g61224/_0_ , \g61225/_0_ , \g61228/_0_ , \g61229/_0_ , \g61230/_0_ , \g61231/_0_ , \g61281/_0_ , \g61293/_1_ , \g61307/_0__syn_2 , \g61309/_0__syn_2 , \g61310/_0__syn_2 , \g61311/_1_ , \g61312/_1_ , \g61313/_1_ , \g61324/_1_ , \g61325/_1_ , \g61326/_1_ , \g61328/_1_ , \g61329/_1_ , \g61330/_1_ , \g61332/_1_ , \g61333/_1_ , \g61334/_1_ , \g61335/_1_ , \g61336/_0_ , \g61338/_0_ , \g61339/_0_ , \g61340/_0_ , \g61377/_1_ , \g61378/_1_ , \g61379/_1_ , \g61388/_1_ , \g61391/_0_ , \g61394/_1_ , \g61395/_1_ , \g61396/_1_ , \g61398/_1_ , \g61399/_1_ , \g61421/_1_ , \g61422/_1_ , \g61423/_1_ , \g61524/_0_ , \g61525/_0_ , \g61526/_0_ , \g61527/_0_ , \g61528/_0_ , \g61529/_0_ , \g61530/_0_ , \g61531/_0_ , \g61532/_0_ , \g61533/_0_ , \g61534/_0_ , \g61535/_0_ , \g61536/_0_ , \g61537/_0_ , \g61538/_0_ , \g61539/_0_ , \g61540/_0_ , \g61541/_0_ , \g61542/_0_ , \g61543/_0_ , \g61544/_0_ , \g61545/_0_ , \g61546/_0_ , \g61547/_0_ , \g61548/_0_ , \g61549/_0_ , \g61550/_0_ , \g61551/_0_ , \g61552/_0_ , \g61553/_0_ , \g61554/_0_ , \g61555/_0_ , \g61556/_0_ , \g61557/_0_ , \g61558/_0_ , \g61559/_0_ , \g61560/_0_ , \g61561/_0_ , \g61562/_0_ , \g61563/_0_ , \g61564/_0_ , \g61565/_0_ , \g61566/_0_ , \g61620/_0_ , \g61621/_0_ , \g61622/_0_ , \g61623/_0_ , \g61753/_0_ , \g61764/_0_ , \g61786/_0_ , \g61795/_0_ , \g61801/_0_ , \g61803/_0_ , \g61808/_0_ , \g61848/_0_ , \g61850/_0_ , \g61851/_0_ , \g62097/_0_ , \g62102/_0_ , \g62115/_0_ , \g62119/_0_ , \g62130/_1_ , \g62131/_0_ , \g62132/_0_ , \g62139/_1_ , \g62140/_1_ , \g62141/_1_ , \g62144/_0_ , \g62145/_0_ , \g62146/_0_ , \g62147/_0_ , \g62150/_0_ , \g62151/_1_ , \g62152/_0_ , \g62153/_1_ , \g62156/_1_ , \g62157/_0_ , \g62159/_0_ , \g62161/_0_ , \g62187/_1_ , \g62190/_1_ , \g62191/_1_ , \g62192/_1_ , \g62194/_1_ , \g62195/_1_ , \g62196/_1_ , \g62203/_0_ , \g62204/_1_ , \g62207/_0__syn_2 , \g62208/_1_ , \g62209/_1_ , \g62210/_1_ , \g62211/_1_ , \g62212/_1_ , \g62217/_0_ , \g62286/_0_ , \g62287/_0_ , \g62288/_0_ , \g62289/_0_ , \g62290/_0_ , \g62291/_0_ , \g62292/_0_ , \g62435/_0_ , \g62436/_0_ , \g62439/_0_ , \g62456/_0_ , \g62486/_1_ , \g62492/_1_ , \g62494/_0_ , \g62495/_1_ , \g62497/_0_ , \g62537/_0_ , \g62544/_0_ , \g62546/_0_ , \g62547/_0_ , \g62549/_3_ , \g62552/_0_ , \g62554/_0_ , \g62555/_0_ , \g62556/_0_ , \g62558/_0_ , \g62559/_0_ , \g62561/_0_ , \g62562/_0_ , \g62566/_0_ , \g62567/_0_ , \g62568/_0_ , \g62569/_0_ , \g62570/_0_ , \g62571/_0_ , \g62572/_0_ , \g62573/_0_ , \g62574/_0_ , \g62575/_0_ , \g62576/_0_ , \g62577/_0_ , \g62578/_0_ , \g62579/_0_ , \g62580/_0_ , \g62581/_0_ , \g62582/_0_ , \g62583/_0_ , \g62584/_0_ , \g62585/_0_ , \g62586/_0_ , \g62587/_0_ , \g62588/_0_ , \g62589/_0_ , \g62590/_0_ , \g62591/_0_ , \g62592/_0_ , \g62593/_0_ , \g62594/_0_ , \g62595/_0_ , \g62596/_0_ , \g62597/_0_ , \g62602/_0_ , \g62607/_0_ , \g62608/_0_ , \g62609/_0_ , \g62619/_0_ , \g62620/_0_ , \g62621/_0_ , \g62622/_0_ , \g62623/_0_ , \g62624/_0_ , \g62626/_0_ , \g62627/_0_ , \g62628/_0_ , \g62629/_0_ , \g62630/_0_ , \g62631/_0_ , \g62632/_0_ , \g62633/_0_ , \g62634/_0_ , \g62635/_0_ , \g62636/_0_ , \g62637/_0_ , \g62638/_0_ , \g62639/_0_ , \g62640/_0_ , \g62641/_0_ , \g62642/_0_ , \g62643/_0_ , \g62644/_0_ , \g62645/_0_ , \g62646/_0_ , \g62647/_0_ , \g62648/_0_ , \g62649/_0_ , \g62650/_0_ , \g62651/_0_ , \g62652/_0_ , \g62653/_0_ , \g62654/_0_ , \g62655/_0_ , \g62656/_0_ , \g62657/_0_ , \g62658/_0_ , \g62659/_0_ , \g62660/_0_ , \g62661/_0_ , \g62674/_0_ , \g62682/_0_ , \g62683/_0_ , \g62689/_0_ , \g62690/_0_ , \g62691/_0_ , \g62694/_0_ , \g62695/_0_ , \g62696/_0_ , \g62698/_0_ , \g62699/_0_ , \g62700/_0_ , \g62723/_0_ , \g62724/_0_ , \g62725/_0_ , \g62726/_0_ , \g62727/_0_ , \g62728/_0_ , \g62735/_0_ , \g62736/_0_ , \g62737/_0_ , \g62738/_0_ , \g62739/_0_ , \g62740/_0_ , \g62754/_0_ , \g62762/_0_ , \g62763/_0_ , \g62764/_0_ , \g62780/_0_ , \g62781/_0_ , \g62785/_0_ , \g62786/_0_ , \g62787/_0_ , \g62791/_0_ , \g62792/_0_ , \g62794/_0_ , \g62804/_0_ , \g62806/_0_ , \g62807/_0_ , \g62811/_0_ , \g62968/_0_ , \g63005/_0_ , \g63041/_0_ , \g63116/_0_ , \g63157/_0_ , \g63164/_0_ , \g63170/_0_ , \g63189/_0_ , \g63202/_0_ , \g63206/_0_ , \g63207/_0_ , \g63265/_0_ , \g63266/_0_ , \g63269/_0_ , \g63271/_0_ , \g63272/_0_ , \g63273/_0_ , \g63274/_0_ , \g63275/_0_ , \g63276/_0_ , \g63277/_0_ , \g63278/_0_ , \g63280/_0_ , \g63281/_0_ , \g63282/_0_ , \g63283/_0_ , \g63284/_0_ , \g63285/_0_ , \g63286/_0_ , \g63287/_0_ , \g63288/_0_ , \g63289/_0_ , \g63290/_0_ , \g63292/_0_ , \g63293/_0_ , \g63294/_0_ , \g63295/_0_ , \g63296/_0_ , \g63297/_0_ , \g63298/_0_ , \g63299/_0_ , \g63302/_0_ , \g63303/_0_ , \g63304/_0_ , \g63305/_0_ , \g63306/_0_ , \g63307/_0_ , \g63308/_0_ , \g63309/_0_ , \g63310/_0_ , \g63311/_0_ , \g63312/_0_ , \g63313/_0_ , \g63314/_0_ , \g63315/_0_ , \g63316/_0_ , \g63317/_0_ , \g63318/_0_ , \g63319/_0_ , \g63320/_0_ , \g63321/_0_ , \g63322/_0_ , \g63323/_0_ , \g63324/_0_ , \g63325/_0_ , \g63326/_0_ , \g63327/_0_ , \g63328/_0_ , \g63329/_0_ , \g63330/_0_ , \g63331/_0_ , \g63339/_0_ , \g63505/_0_ , \g63525/_0_ , \g63543/_1_ , \g63602/_0_ , \g63653/_0_ , \g63663/_1_ , \g63677/_0_ , \g63694/_0_ , \g63729/_0_ , \g63766/_0_ , \g63771/_1_ , \g63773/_1_ , \g63784/_1_ , \g63964/_0_ , \g63965/_0_ , \g63966/_0_ , \g63967/_0_ , \g64257/_1_ , \g64266/_0_ , \g64275/_0_ , \g64400/_0_ , \g64416/_0_ , \g64470/_3_ , \g64473/_0_ , \g64474/_0_ , \g64475/_0_ , \g64479/_0_ , \g64480/_0_ , \g64481/_0_ , \g64483/_0_ , \g64484/_0_ , \g64485/_0_ , \g64486/_0_ , \g64493/_0_ , \g64494/_0_ , \g64495/_0_ , \g64496/_0_ , \g64505/_3_ , \g64507/_0_ , \g64508/_0_ , \g64510/_0_ , \g64511/_0_ , \g64544/_0_ , \g64545/_0_ , \g64546/_0_ , \g64639/_0_ , \g64641/_0_ , \g64642/_0_ , \g64645/_0_ , \g64650/_0_ , \g64737/_0_ , \g64738/_0_ , \g65066/_0_ , \g65070/_0_ , \g65090/_0_ , \g65102/_0_ , \g65102/_3_ , \g65126/_3_ , \g65147/_3_ , \g65163/_0_ , \g65176/_3_ , \g65178/_0_ , \g65182/_0_ , \g65190/_1_ , \g65191/_0_ , \g65196/_0_ , \g65268/_0_ , \g65275/_0_ , \g65290/_0_ , \g65290/_3_ , \g65291/_0_ , \g65292/_0_ , \g65298/_0_ , \g65298/_3_ , \g65314/_0_ , \g65314/_3_ , \g65319/_3_ , \g65335/_0_ , \g65342/_0_ , \g65348/_0_ , \g65422/_0_ , \g65465/_1_ , \g65469/_1_ , \g65478/_1_ , \g65507/_0_ , \g65548/_0_ , \g65699/_1_ , \g65713/_1_ , \g65835/_0_ , \g65860/_0_ , \g65863/_0_ , \g66094/_1_ , \g66102/_0_ , \g66107/_0_ , \g66130/_3_ , \g66131/_3_ , \g66228/_1_ , \g66348/_1_ , \g66543/_0_ , \g66549/_1_ , \g66640/_3_ , \g66641/_3_ , \g66950/_1_ , \g67111/_0_ , \g67219/_0_ , \g67263/_0_ , \g67909/_1_ , \g68049/_0_ , \g68220/_0_ , \g68413/_0_ , \g68511/_0_ , \g68536/_0_ , \g68543/_1_ , \g68554/_0_ , \g68559/_0_ , \g70915/_0_ , \g71108/_1_ , \g71115/_2_ , \g71244_dup/_0_ , \g71368/_0_ , \g71581/_0_ , \g71720/_0_ , \g785_reg/P0001 , \g789_reg/P0001 , \g797_reg/P0001 , \g809_reg/P0001 , \g813_reg/P0001 , \g966_reg/P0001 , \g968_reg/P0001 , \g970_reg/P0001 , \g972_reg/P0001 , \g974_reg/P0001 , \g976_reg/P0001 , \g978_reg/P0001 );
	input \g1000_reg/NET0131  ;
	input \g1001_reg/NET0131  ;
	input \g1002_reg/NET0131  ;
	input \g1003_reg/NET0131  ;
	input \g1004_reg/NET0131  ;
	input \g1005_reg/NET0131  ;
	input \g1006_reg/NET0131  ;
	input \g1007_reg/NET0131  ;
	input \g1008_reg/NET0131  ;
	input \g1009_reg/NET0131  ;
	input \g1010_reg/NET0131  ;
	input \g1011_reg/NET0131  ;
	input \g1018_reg/NET0131  ;
	input \g101_reg/NET0131  ;
	input \g1024_reg/NET0131  ;
	input \g1030_reg/NET0131  ;
	input \g1033_reg/NET0131  ;
	input \g1036_reg/NET0131  ;
	input \g1038_reg/NET0131  ;
	input \g1040_reg/NET0131  ;
	input \g1041_reg/NET0131  ;
	input \g1045_reg/NET0131  ;
	input \g1048_reg/NET0131  ;
	input \g1051_reg/NET0131  ;
	input \g1053_reg/NET0131  ;
	input \g1055_reg/NET0131  ;
	input \g1056_reg/NET0131  ;
	input \g105_reg/NET0131  ;
	input \g1060_reg/NET0131  ;
	input \g1063_reg/NET0131  ;
	input \g1066_reg/NET0131  ;
	input \g1068_reg/NET0131  ;
	input \g1070_reg/NET0131  ;
	input \g1071_reg/NET0131  ;
	input \g1075_reg/NET0131  ;
	input \g1078_reg/NET0131  ;
	input \g1081_reg/NET0131  ;
	input \g1083_reg/NET0131  ;
	input \g1085_reg/NET0131  ;
	input \g1088_reg/NET0131  ;
	input \g1089_reg/NET0131  ;
	input \g1090_reg/NET0131  ;
	input \g1091_reg/NET0131  ;
	input \g1092_reg/NET0131  ;
	input \g1095_reg/NET0131  ;
	input \g1098_reg/NET0131  ;
	input \g109_reg/NET0131  ;
	input \g1101_reg/NET0131  ;
	input \g1104_reg/NET0131  ;
	input \g1107_reg/NET0131  ;
	input \g1110_reg/NET0131  ;
	input \g1113_reg/NET0131  ;
	input \g1114_reg/NET0131  ;
	input \g1115_reg/NET0131  ;
	input \g1116_reg/NET0131  ;
	input \g1119_reg/NET0131  ;
	input \g1122_reg/NET0131  ;
	input \g1125_reg/NET0131  ;
	input \g1128_reg/NET0131  ;
	input \g1131_reg/NET0131  ;
	input \g1134_reg/NET0131  ;
	input \g1135_reg/NET0131  ;
	input \g1136_reg/NET0131  ;
	input \g1138_reg/NET0131  ;
	input \g113_reg/NET0131  ;
	input \g1140_reg/NET0131  ;
	input \g1151_reg/NET0131  ;
	input \g1164_reg/NET0131  ;
	input \g1165_reg/NET0131  ;
	input \g1166_reg/NET0131  ;
	input \g1167_reg/NET0131  ;
	input \g1171_reg/NET0131  ;
	input \g1173_reg/NET0131  ;
	input \g1174_reg/NET0131  ;
	input \g1175_reg/NET0131  ;
	input \g1176_reg/NET0131  ;
	input \g1177_reg/NET0131  ;
	input \g117_reg/NET0131  ;
	input \g1180_reg/NET0131  ;
	input \g1183_reg/NET0131  ;
	input \g1186_reg/NET0131  ;
	input \g1192_reg/NET0131  ;
	input \g1193_reg/NET0131  ;
	input \g1196_reg/NET0131  ;
	input \g1210_reg/NET0131  ;
	input \g1211_reg/NET0131  ;
	input \g1215_reg/NET0131  ;
	input \g1216_reg/NET0131  ;
	input \g1217_reg/NET0131  ;
	input \g1218_reg/NET0131  ;
	input \g1219_reg/NET0131  ;
	input \g121_reg/NET0131  ;
	input \g1220_reg/NET0131  ;
	input \g1222_reg/NET0131  ;
	input \g1223_reg/NET0131  ;
	input \g1224_reg/NET0131  ;
	input \g1227_reg/NET0131  ;
	input \g1228_reg/NET0131  ;
	input \g1230_reg/NET0131  ;
	input \g1234_reg/NET0131  ;
	input \g1240_reg/NET0131  ;
	input \g1243_reg/NET0131  ;
	input \g1245_reg/NET0131  ;
	input \g1249_pad  ;
	input \g1251_reg/NET0131  ;
	input \g1253_reg/NET0131  ;
	input \g1255_reg/NET0131  ;
	input \g1257_reg/NET0131  ;
	input \g1259_reg/NET0131  ;
	input \g125_reg/NET0131  ;
	input \g1261_reg/NET0131  ;
	input \g1262_reg/NET0131  ;
	input \g1263_reg/NET0131  ;
	input \g1264_reg/NET0131  ;
	input \g1265_reg/NET0131  ;
	input \g1266_reg/NET0131  ;
	input \g1267_reg/NET0131  ;
	input \g1268_reg/NET0131  ;
	input \g1269_reg/NET0131  ;
	input \g1270_reg/NET0131  ;
	input \g1271_reg/NET0131  ;
	input \g1272_reg/NET0131  ;
	input \g1273_reg/NET0131  ;
	input \g1276_reg/NET0131  ;
	input \g1279_reg/NET0131  ;
	input \g1282_reg/NET0131  ;
	input \g1285_reg/NET0131  ;
	input \g1288_reg/NET0131  ;
	input \g1291_reg/NET0131  ;
	input \g1294_reg/NET0131  ;
	input \g1297_reg/NET0131  ;
	input \g129_reg/NET0131  ;
	input \g1300_reg/NET0131  ;
	input \g1303_reg/NET0131  ;
	input \g1306_reg/NET0131  ;
	input \g130_reg/NET0131  ;
	input \g1316_reg/NET0131  ;
	input \g1319_reg/NET0131  ;
	input \g131_reg/NET0131  ;
	input \g1326_reg/NET0131  ;
	input \g132_reg/NET0131  ;
	input \g1332_reg/NET0131  ;
	input \g1339_reg/NET0131  ;
	input \g133_reg/NET0131  ;
	input \g1345_reg/NET0131  ;
	input \g1346_reg/NET0131  ;
	input \g134_reg/NET0131  ;
	input \g1352_reg/NET0131  ;
	input \g1358_reg/NET0131  ;
	input \g1365_reg/NET0131  ;
	input \g1372_reg/NET0131  ;
	input \g1378_reg/NET0131  ;
	input \g1384_reg/NET0131  ;
	input \g1385_reg/NET0131  ;
	input \g1386_reg/NET0131  ;
	input \g1387_reg/NET0131  ;
	input \g1388_reg/NET0131  ;
	input \g1389_reg/NET0131  ;
	input \g1390_reg/NET0131  ;
	input \g1391_reg/NET0131  ;
	input \g1392_reg/NET0131  ;
	input \g1393_reg/NET0131  ;
	input \g1394_reg/NET0131  ;
	input \g1395_reg/NET0131  ;
	input \g1396_reg/NET0131  ;
	input \g1397_reg/NET0131  ;
	input \g1398_reg/NET0131  ;
	input \g1399_reg/NET0131  ;
	input \g1400_reg/NET0131  ;
	input \g1401_reg/NET0131  ;
	input \g1402_reg/NET0131  ;
	input \g1403_reg/NET0131  ;
	input \g1404_reg/NET0131  ;
	input \g1405_reg/NET0131  ;
	input \g1406_reg/NET0131  ;
	input \g1407_reg/NET0131  ;
	input \g1408_reg/NET0131  ;
	input \g1409_reg/NET0131  ;
	input \g1410_reg/NET0131  ;
	input \g1411_reg/NET0131  ;
	input \g1412_reg/NET0131  ;
	input \g1413_reg/NET0131  ;
	input \g1414_reg/NET0131  ;
	input \g1415_reg/NET0131  ;
	input \g1416_reg/NET0131  ;
	input \g1417_reg/NET0131  ;
	input \g1418_reg/NET0131  ;
	input \g1419_reg/NET0131  ;
	input \g141_reg/NET0131  ;
	input \g1420_reg/NET0131  ;
	input \g1421_reg/NET0131  ;
	input \g1422_reg/NET0131  ;
	input \g1423_reg/NET0131  ;
	input \g1424_reg/NET0131  ;
	input \g1425_reg/NET0131  ;
	input \g1426_reg/NET0131  ;
	input \g142_reg/NET0131  ;
	input \g1430_reg/NET0131  ;
	input \g1435_reg/NET0131  ;
	input \g1439_reg/NET0131  ;
	input \g143_reg/NET0131  ;
	input \g1444_reg/NET0131  ;
	input \g1448_reg/NET0131  ;
	input \g144_reg/NET0131  ;
	input \g1453_reg/NET0131  ;
	input \g1457_reg/NET0131  ;
	input \g145_reg/NET0131  ;
	input \g1462_reg/NET0131  ;
	input \g1466_reg/NET0131  ;
	input \g146_reg/NET0131  ;
	input \g1471_reg/NET0131  ;
	input \g1476_reg/NET0131  ;
	input \g147_reg/NET0131  ;
	input \g1481_reg/NET0131  ;
	input \g1486_reg/NET0131  ;
	input \g148_reg/NET0131  ;
	input \g1491_reg/NET0131  ;
	input \g1496_reg/NET0131  ;
	input \g149_reg/NET0131  ;
	input \g1501_reg/NET0131  ;
	input \g1506_reg/NET0131  ;
	input \g150_reg/NET0131  ;
	input \g1511_reg/NET0131  ;
	input \g1512_reg/NET0131  ;
	input \g1513_reg/NET0131  ;
	input \g1514_reg/NET0131  ;
	input \g1515_reg/NET0131  ;
	input \g1516_reg/NET0131  ;
	input \g151_reg/NET0131  ;
	input \g1523_reg/NET0131  ;
	input \g1524_reg/NET0131  ;
	input \g1525_reg/NET0131  ;
	input \g1526_reg/NET0131  ;
	input \g1527_reg/NET0131  ;
	input \g1528_reg/NET0131  ;
	input \g1529_reg/NET0131  ;
	input \g152_reg/NET0131  ;
	input \g1530_reg/NET0131  ;
	input \g1531_reg/NET0131  ;
	input \g1532_reg/NET0131  ;
	input \g1533_reg/NET0131  ;
	input \g1534_reg/NET0131  ;
	input \g1535_reg/NET0131  ;
	input \g1536_reg/NET0131  ;
	input \g1537_reg/NET0131  ;
	input \g1538_reg/NET0131  ;
	input \g1539_reg/NET0131  ;
	input \g153_reg/NET0131  ;
	input \g1540_reg/NET0131  ;
	input \g1541_reg/NET0131  ;
	input \g1542_reg/NET0131  ;
	input \g1543_reg/NET0131  ;
	input \g1544_reg/NET0131  ;
	input \g1545_reg/NET0131  ;
	input \g1546_reg/NET0131  ;
	input \g154_reg/NET0131  ;
	input \g1550_reg/NET0131  ;
	input \g1551_reg/NET0131  ;
	input \g1552_reg/NET0131  ;
	input \g1553_reg/NET0131  ;
	input \g1554_reg/NET0131  ;
	input \g1555_reg/NET0131  ;
	input \g1556_reg/NET0131  ;
	input \g1557_reg/NET0131  ;
	input \g1558_reg/NET0131  ;
	input \g1559_reg/NET0131  ;
	input \g155_reg/NET0131  ;
	input \g1560_reg/NET0131  ;
	input \g1561_reg/NET0131  ;
	input \g1563_reg/NET0131  ;
	input \g1567_reg/NET0131  ;
	input \g156_reg/NET0131  ;
	input \g1570_reg/NET0131  ;
	input \g1573_reg/NET0131  ;
	input \g1576_reg/NET0131  ;
	input \g1579_reg/NET0131  ;
	input \g157_reg/NET0131  ;
	input \g1582_reg/NET0131  ;
	input \g1585_reg/NET0131  ;
	input \g1588_reg/NET0131  ;
	input \g158_reg/NET0131  ;
	input \g1591_reg/NET0131  ;
	input \g1594_reg/NET0131  ;
	input \g1597_reg/NET0131  ;
	input \g159_reg/NET0131  ;
	input \g1600_reg/NET0131  ;
	input \g1603_reg/NET0131  ;
	input \g1606_reg/NET0131  ;
	input \g1609_reg/NET0131  ;
	input \g160_reg/NET0131  ;
	input \g1612_reg/NET0131  ;
	input \g1615_reg/NET0131  ;
	input \g1618_reg/NET0131  ;
	input \g161_reg/NET0131  ;
	input \g1621_reg/NET0131  ;
	input \g1624_reg/NET0131  ;
	input \g1627_reg/NET0131  ;
	input \g16297_pad  ;
	input \g162_reg/NET0131  ;
	input \g1630_reg/NET0131  ;
	input \g1633_reg/NET0131  ;
	input \g16355_pad  ;
	input \g1636_reg/NET0131  ;
	input \g16399_pad  ;
	input \g1639_reg/NET0131  ;
	input \g163_reg/NET0131  ;
	input \g1642_reg/NET0131  ;
	input \g16437_pad  ;
	input \g1645_reg/NET0131  ;
	input \g1648_reg/NET0131  ;
	input \g164_reg/NET0131  ;
	input \g1651_reg/NET0131  ;
	input \g1654_reg/NET0131  ;
	input \g1660_reg/NET0131  ;
	input \g1662_reg/NET0131  ;
	input \g1664_reg/NET0131  ;
	input \g1666_reg/NET0131  ;
	input \g1668_reg/NET0131  ;
	input \g1670_reg/NET0131  ;
	input \g1672_reg/NET0131  ;
	input \g1679_reg/NET0131  ;
	input \g1680_reg/NET0131  ;
	input \g1686_reg/NET0131  ;
	input \g168_reg/NET0131  ;
	input \g1693_reg/NET0131  ;
	input \g1694_reg/NET0131  ;
	input \g1695_reg/NET0131  ;
	input \g1696_reg/NET0131  ;
	input \g1697_reg/NET0131  ;
	input \g1698_reg/NET0131  ;
	input \g1699_reg/NET0131  ;
	input \g169_reg/NET0131  ;
	input \g1700_reg/NET0131  ;
	input \g1701_reg/NET0131  ;
	input \g1702_reg/NET0131  ;
	input \g1703_reg/NET0131  ;
	input \g1704_reg/NET0131  ;
	input \g1705_reg/NET0131  ;
	input \g170_reg/NET0131  ;
	input \g171_reg/NET0131  ;
	input \g1724_reg/NET0131  ;
	input \g1727_reg/NET0131  ;
	input \g172_reg/NET0131  ;
	input \g1730_reg/NET0131  ;
	input \g1732_reg/NET0131  ;
	input \g1734_reg/NET0131  ;
	input \g1735_reg/NET0131  ;
	input \g1739_reg/NET0131  ;
	input \g173_reg/NET0131  ;
	input \g1742_reg/NET0131  ;
	input \g1745_reg/NET0131  ;
	input \g1747_reg/NET0131  ;
	input \g1749_reg/NET0131  ;
	input \g174_reg/NET0131  ;
	input \g1750_reg/NET0131  ;
	input \g1754_reg/NET0131  ;
	input \g1757_reg/NET0131  ;
	input \g175_reg/NET0131  ;
	input \g1760_reg/NET0131  ;
	input \g1762_reg/NET0131  ;
	input \g1764_reg/NET0131  ;
	input \g1765_reg/NET0131  ;
	input \g1769_reg/NET0131  ;
	input \g176_reg/NET0131  ;
	input \g1772_reg/NET0131  ;
	input \g1775_reg/NET0131  ;
	input \g1777_reg/NET0131  ;
	input \g1779_reg/NET0131  ;
	input \g177_reg/NET0131  ;
	input \g1783_reg/NET0131  ;
	input \g1784_reg/NET0131  ;
	input \g1785_reg/NET0131  ;
	input \g1789_reg/NET0131  ;
	input \g178_reg/NET0131  ;
	input \g1792_reg/NET0131  ;
	input \g1795_reg/NET0131  ;
	input \g1798_reg/NET0131  ;
	input \g179_reg/NET0131  ;
	input \g1801_reg/NET0131  ;
	input \g1804_reg/NET0131  ;
	input \g1807_reg/NET0131  ;
	input \g1808_reg/NET0131  ;
	input \g1809_reg/NET0131  ;
	input \g1810_reg/NET0131  ;
	input \g1813_reg/NET0131  ;
	input \g1816_reg/NET0131  ;
	input \g1819_reg/NET0131  ;
	input \g1822_reg/NET0131  ;
	input \g1825_reg/NET0131  ;
	input \g1828_reg/NET0131  ;
	input \g1829_reg/NET0131  ;
	input \g1830_reg/NET0131  ;
	input \g1832_reg/NET0131  ;
	input \g1834_reg/NET0131  ;
	input \g1845_reg/NET0131  ;
	input \g1846_reg/NET0131  ;
	input \g1849_reg/NET0131  ;
	input \g1852_reg/NET0131  ;
	input \g1858_reg/NET0131  ;
	input \g1859_reg/NET0131  ;
	input \g185_reg/NET0131  ;
	input \g1860_reg/NET0131  ;
	input \g1861_reg/NET0131  ;
	input \g1865_reg/NET0131  ;
	input \g1867_reg/NET0131  ;
	input \g1868_reg/NET0131  ;
	input \g1869_reg/NET0131  ;
	input \g186_reg/NET0131  ;
	input \g1870_reg/NET0131  ;
	input \g1871_reg/NET0131  ;
	input \g1874_reg/NET0131  ;
	input \g1877_reg/NET0131  ;
	input \g1880_reg/NET0131  ;
	input \g1886_reg/NET0131  ;
	input \g1887_reg/NET0131  ;
	input \g189_reg/NET0131  ;
	input \g1904_reg/NET0131  ;
	input \g1905_reg/NET0131  ;
	input \g1909_reg/NET0131  ;
	input \g1910_reg/NET0131  ;
	input \g1911_reg/NET0131  ;
	input \g1912_reg/NET0131  ;
	input \g1913_reg/NET0131  ;
	input \g1914_reg/NET0131  ;
	input \g1916_reg/NET0131  ;
	input \g1917_reg/NET0131  ;
	input \g1918_reg/NET0131  ;
	input \g1921_reg/NET0131  ;
	input \g1922_reg/NET0131  ;
	input \g1924_reg/NET0131  ;
	input \g1928_reg/NET0131  ;
	input \g192_reg/NET0131  ;
	input \g1939_reg/NET0131  ;
	input \g1943_pad  ;
	input \g1945_reg/NET0131  ;
	input \g1947_reg/NET0131  ;
	input \g1949_reg/NET0131  ;
	input \g1951_reg/NET0131  ;
	input \g1953_reg/NET0131  ;
	input \g1955_reg/NET0131  ;
	input \g1956_reg/NET0131  ;
	input \g1957_reg/NET0131  ;
	input \g1958_reg/NET0131  ;
	input \g1959_reg/NET0131  ;
	input \g195_reg/NET0131  ;
	input \g1960_reg/NET0131  ;
	input \g1961_reg/NET0131  ;
	input \g1962_reg/NET0131  ;
	input \g1963_reg/NET0131  ;
	input \g1964_reg/NET0131  ;
	input \g1965_reg/NET0131  ;
	input \g1966_reg/NET0131  ;
	input \g1967_reg/NET0131  ;
	input \g1970_reg/NET0131  ;
	input \g1973_reg/NET0131  ;
	input \g1976_reg/NET0131  ;
	input \g1979_reg/NET0131  ;
	input \g1982_reg/NET0131  ;
	input \g1985_reg/NET0131  ;
	input \g1988_reg/NET0131  ;
	input \g198_reg/NET0131  ;
	input \g1991_reg/NET0131  ;
	input \g1994_reg/NET0131  ;
	input \g1997_reg/NET0131  ;
	input \g2000_reg/NET0131  ;
	input \g201_reg/NET0131  ;
	input \g204_reg/NET0131  ;
	input \g2078_reg/NET0131  ;
	input \g2079_reg/NET0131  ;
	input \g207_reg/NET0131  ;
	input \g2080_reg/NET0131  ;
	input \g2081_reg/NET0131  ;
	input \g2082_reg/NET0131  ;
	input \g2083_reg/NET0131  ;
	input \g2084_reg/NET0131  ;
	input \g2085_reg/NET0131  ;
	input \g2086_reg/NET0131  ;
	input \g2087_reg/NET0131  ;
	input \g2088_reg/NET0131  ;
	input \g2089_reg/NET0131  ;
	input \g2090_reg/NET0131  ;
	input \g2091_reg/NET0131  ;
	input \g2092_reg/NET0131  ;
	input \g2093_reg/NET0131  ;
	input \g2094_reg/NET0131  ;
	input \g2095_reg/NET0131  ;
	input \g2096_reg/NET0131  ;
	input \g2097_reg/NET0131  ;
	input \g2098_reg/NET0131  ;
	input \g2099_reg/NET0131  ;
	input \g2100_reg/NET0131  ;
	input \g2101_reg/NET0131  ;
	input \g2102_reg/NET0131  ;
	input \g2103_reg/NET0131  ;
	input \g2104_reg/NET0131  ;
	input \g2105_reg/NET0131  ;
	input \g2106_reg/NET0131  ;
	input \g2107_reg/NET0131  ;
	input \g2108_reg/NET0131  ;
	input \g2109_reg/NET0131  ;
	input \g210_reg/NET0131  ;
	input \g2110_reg/NET0131  ;
	input \g2111_reg/NET0131  ;
	input \g2112_reg/NET0131  ;
	input \g2113_reg/NET0131  ;
	input \g2114_reg/NET0131  ;
	input \g2115_reg/NET0131  ;
	input \g2116_reg/NET0131  ;
	input \g2117_reg/NET0131  ;
	input \g2118_reg/NET0131  ;
	input \g2119_reg/NET0131  ;
	input \g213_reg/NET0131  ;
	input \g2165_reg/NET0131  ;
	input \g216_reg/NET0131  ;
	input \g2170_reg/NET0131  ;
	input \g2175_reg/NET0131  ;
	input \g2180_reg/NET0131  ;
	input \g2185_reg/NET0131  ;
	input \g2190_reg/NET0131  ;
	input \g2195_reg/NET0131  ;
	input \g219_reg/NET0131  ;
	input \g2200_reg/NET0131  ;
	input \g2205_reg/NET0131  ;
	input \g2206_reg/NET0131  ;
	input \g2207_reg/NET0131  ;
	input \g2208_reg/NET0131  ;
	input \g2209_reg/NET0131  ;
	input \g2210_reg/NET0131  ;
	input \g2217_reg/NET0131  ;
	input \g2218_reg/NET0131  ;
	input \g2219_reg/NET0131  ;
	input \g2220_reg/NET0131  ;
	input \g2221_reg/NET0131  ;
	input \g2222_reg/NET0131  ;
	input \g2223_reg/NET0131  ;
	input \g2224_reg/NET0131  ;
	input \g2225_reg/NET0131  ;
	input \g2226_reg/NET0131  ;
	input \g2227_reg/NET0131  ;
	input \g2228_reg/NET0131  ;
	input \g2229_reg/NET0131  ;
	input \g222_reg/NET0131  ;
	input \g2230_reg/NET0131  ;
	input \g2231_reg/NET0131  ;
	input \g2232_reg/NET0131  ;
	input \g2233_reg/NET0131  ;
	input \g2234_reg/NET0131  ;
	input \g2235_reg/NET0131  ;
	input \g2236_reg/NET0131  ;
	input \g2237_reg/NET0131  ;
	input \g2238_reg/NET0131  ;
	input \g2239_reg/NET0131  ;
	input \g2240_reg/NET0131  ;
	input \g2244_reg/NET0131  ;
	input \g2245_reg/NET0131  ;
	input \g2246_reg/NET0131  ;
	input \g2247_reg/NET0131  ;
	input \g2248_reg/NET0131  ;
	input \g2249_reg/NET0131  ;
	input \g2250_reg/NET0131  ;
	input \g2251_reg/NET0131  ;
	input \g2252_reg/NET0131  ;
	input \g2253_reg/NET0131  ;
	input \g2254_reg/NET0131  ;
	input \g2255_reg/NET0131  ;
	input \g225_reg/NET0131  ;
	input \g2261_reg/NET0131  ;
	input \g2264_reg/NET0131  ;
	input \g2267_reg/NET0131  ;
	input \g2270_reg/NET0131  ;
	input \g2273_reg/NET0131  ;
	input \g2276_reg/NET0131  ;
	input \g2279_reg/NET0131  ;
	input \g2282_reg/NET0131  ;
	input \g2285_reg/NET0131  ;
	input \g2288_reg/NET0131  ;
	input \g228_reg/NET0131  ;
	input \g2291_reg/NET0131  ;
	input \g2294_reg/NET0131  ;
	input \g2297_reg/NET0131  ;
	input \g2300_reg/NET0131  ;
	input \g2303_reg/NET0131  ;
	input \g2306_reg/NET0131  ;
	input \g2309_reg/NET0131  ;
	input \g2312_reg/NET0131  ;
	input \g2315_reg/NET0131  ;
	input \g2318_reg/NET0131  ;
	input \g231_reg/NET0131  ;
	input \g2321_reg/NET0131  ;
	input \g2324_reg/NET0131  ;
	input \g2327_reg/NET0131  ;
	input \g2330_reg/NET0131  ;
	input \g2333_reg/NET0131  ;
	input \g2336_reg/NET0131  ;
	input \g2339_reg/NET0131  ;
	input \g2342_reg/NET0131  ;
	input \g2345_reg/NET0131  ;
	input \g2348_reg/NET0131  ;
	input \g234_reg/NET0131  ;
	input \g2354_reg/NET0131  ;
	input \g2356_reg/NET0131  ;
	input \g2358_reg/NET0131  ;
	input \g2360_reg/NET0131  ;
	input \g2362_reg/NET0131  ;
	input \g2364_reg/NET0131  ;
	input \g2366_reg/NET0131  ;
	input \g2373_reg/NET0131  ;
	input \g2374_reg/NET0131  ;
	input \g237_reg/NET0131  ;
	input \g2380_reg/NET0131  ;
	input \g2387_reg/NET0131  ;
	input \g2388_reg/NET0131  ;
	input \g2389_reg/NET0131  ;
	input \g2390_reg/NET0131  ;
	input \g2391_reg/NET0131  ;
	input \g2392_reg/NET0131  ;
	input \g2393_reg/NET0131  ;
	input \g2394_reg/NET0131  ;
	input \g2395_reg/NET0131  ;
	input \g2396_reg/NET0131  ;
	input \g2397_reg/NET0131  ;
	input \g2398_reg/NET0131  ;
	input \g2399_reg/NET0131  ;
	input \g240_reg/NET0131  ;
	input \g2418_reg/NET0131  ;
	input \g2421_reg/NET0131  ;
	input \g2424_reg/NET0131  ;
	input \g2426_reg/NET0131  ;
	input \g2428_reg/NET0131  ;
	input \g2429_reg/NET0131  ;
	input \g2433_reg/NET0131  ;
	input \g2436_reg/NET0131  ;
	input \g2439_reg/NET0131  ;
	input \g243_reg/NET0131  ;
	input \g2441_reg/NET0131  ;
	input \g2443_reg/NET0131  ;
	input \g2444_reg/NET0131  ;
	input \g2448_reg/NET0131  ;
	input \g2451_reg/NET0131  ;
	input \g2454_reg/NET0131  ;
	input \g2456_reg/NET0131  ;
	input \g2458_reg/NET0131  ;
	input \g2459_reg/NET0131  ;
	input \g2463_reg/NET0131  ;
	input \g2466_reg/NET0131  ;
	input \g2469_reg/NET0131  ;
	input \g246_reg/NET0131  ;
	input \g2471_reg/NET0131  ;
	input \g2473_reg/NET0131  ;
	input \g2477_reg/NET0131  ;
	input \g2478_reg/NET0131  ;
	input \g2479_reg/NET0131  ;
	input \g2483_reg/NET0131  ;
	input \g2486_reg/NET0131  ;
	input \g2489_reg/NET0131  ;
	input \g2492_reg/NET0131  ;
	input \g2495_reg/NET0131  ;
	input \g2498_reg/NET0131  ;
	input \g249_reg/NET0131  ;
	input \g2501_reg/NET0131  ;
	input \g2502_reg/NET0131  ;
	input \g2503_reg/NET0131  ;
	input \g2504_reg/NET0131  ;
	input \g2507_reg/NET0131  ;
	input \g2510_reg/NET0131  ;
	input \g2513_reg/NET0131  ;
	input \g2516_reg/NET0131  ;
	input \g2519_reg/NET0131  ;
	input \g2522_reg/NET0131  ;
	input \g2523_reg/NET0131  ;
	input \g2524_reg/NET0131  ;
	input \g2526_reg/NET0131  ;
	input \g2528_reg/NET0131  ;
	input \g252_reg/NET0131  ;
	input \g2539_reg/NET0131  ;
	input \g2540_reg/NET0131  ;
	input \g2543_reg/NET0131  ;
	input \g2546_reg/NET0131  ;
	input \g2552_reg/NET0131  ;
	input \g2553_reg/NET0131  ;
	input \g2554_reg/NET0131  ;
	input \g2555_reg/NET0131  ;
	input \g2559_reg/NET0131  ;
	input \g255_reg/NET0131  ;
	input \g2561_reg/NET0131  ;
	input \g2562_reg/NET0131  ;
	input \g2563_reg/NET0131  ;
	input \g2564_reg/NET0131  ;
	input \g2565_reg/NET0131  ;
	input \g2568_reg/NET0131  ;
	input \g2571_reg/NET0131  ;
	input \g2574_reg/NET0131  ;
	input \g2580_reg/NET0131  ;
	input \g2581_reg/NET0131  ;
	input \g258_reg/NET0131  ;
	input \g2598_reg/NET0131  ;
	input \g2599_reg/NET0131  ;
	input \g2603_reg/NET0131  ;
	input \g2604_reg/NET0131  ;
	input \g2605_reg/NET0131  ;
	input \g2606_reg/NET0131  ;
	input \g2607_reg/NET0131  ;
	input \g2608_reg/NET0131  ;
	input \g2610_reg/NET0131  ;
	input \g2611_reg/NET0131  ;
	input \g2612_reg/NET0131  ;
	input \g2615_reg/NET0131  ;
	input \g2616_reg/NET0131  ;
	input \g2618_reg/NET0131  ;
	input \g261_reg/NET0131  ;
	input \g2622_reg/NET0131  ;
	input \g2633_reg/NET0131  ;
	input \g2637_pad  ;
	input \g2639_reg/NET0131  ;
	input \g2641_reg/NET0131  ;
	input \g2643_reg/NET0131  ;
	input \g2645_reg/NET0131  ;
	input \g2647_reg/NET0131  ;
	input \g2649_reg/NET0131  ;
	input \g264_reg/NET0131  ;
	input \g2650_reg/NET0131  ;
	input \g2651_reg/NET0131  ;
	input \g2652_reg/NET0131  ;
	input \g2653_reg/NET0131  ;
	input \g2654_reg/NET0131  ;
	input \g2655_reg/NET0131  ;
	input \g2656_reg/NET0131  ;
	input \g2657_reg/NET0131  ;
	input \g2658_reg/NET0131  ;
	input \g2659_reg/NET0131  ;
	input \g2660_reg/NET0131  ;
	input \g2661_reg/NET0131  ;
	input \g2664_reg/NET0131  ;
	input \g2667_reg/NET0131  ;
	input \g2670_reg/NET0131  ;
	input \g2673_reg/NET0131  ;
	input \g2676_reg/NET0131  ;
	input \g2679_reg/NET0131  ;
	input \g267_reg/NET0131  ;
	input \g2682_reg/NET0131  ;
	input \g2685_reg/NET0131  ;
	input \g2688_reg/NET0131  ;
	input \g2691_reg/NET0131  ;
	input \g2694_reg/NET0131  ;
	input \g270_reg/NET0131  ;
	input \g273_reg/NET0131  ;
	input \g2772_reg/NET0131  ;
	input \g2773_reg/NET0131  ;
	input \g2774_reg/NET0131  ;
	input \g2775_reg/NET0131  ;
	input \g2776_reg/NET0131  ;
	input \g2777_reg/NET0131  ;
	input \g2778_reg/NET0131  ;
	input \g2779_reg/NET0131  ;
	input \g2780_reg/NET0131  ;
	input \g2781_reg/NET0131  ;
	input \g2782_reg/NET0131  ;
	input \g2783_reg/NET0131  ;
	input \g2784_reg/NET0131  ;
	input \g2785_reg/NET0131  ;
	input \g2786_reg/NET0131  ;
	input \g2787_reg/NET0131  ;
	input \g2788_reg/NET0131  ;
	input \g2789_reg/NET0131  ;
	input \g2790_reg/NET0131  ;
	input \g2791_reg/NET0131  ;
	input \g2792_reg/NET0131  ;
	input \g2793_reg/NET0131  ;
	input \g2794_reg/NET0131  ;
	input \g2795_reg/NET0131  ;
	input \g2796_reg/NET0131  ;
	input \g2797_reg/NET0131  ;
	input \g2798_reg/NET0131  ;
	input \g2799_reg/NET0131  ;
	input \g279_reg/NET0131  ;
	input \g2800_reg/NET0131  ;
	input \g2801_reg/NET0131  ;
	input \g2802_reg/NET0131  ;
	input \g2803_reg/NET0131  ;
	input \g2804_reg/NET0131  ;
	input \g2805_reg/NET0131  ;
	input \g2806_reg/NET0131  ;
	input \g2807_reg/NET0131  ;
	input \g2808_reg/NET0131  ;
	input \g2809_reg/NET0131  ;
	input \g2810_reg/NET0131  ;
	input \g2811_reg/NET0131  ;
	input \g2812_reg/NET0131  ;
	input \g2813_reg/NET0131  ;
	input \g2814_reg/NET0131  ;
	input \g2817_reg/NET0131  ;
	input \g281_reg/NET0131  ;
	input \g283_reg/NET0131  ;
	input \g285_reg/NET0131  ;
	input \g2874_reg/NET0131  ;
	input \g2879_reg/NET0131  ;
	input \g287_reg/NET0131  ;
	input \g2883_reg/NET0131  ;
	input \g2888_reg/NET0131  ;
	input \g2892_reg/NET0131  ;
	input \g2896_reg/NET0131  ;
	input \g289_reg/NET0131  ;
	input \g2900_reg/NET0131  ;
	input \g2903_reg/NET0131  ;
	input \g2908_reg/NET0131  ;
	input \g2912_reg/NET0131  ;
	input \g2917_reg/NET0131  ;
	input \g291_reg/NET0131  ;
	input \g2920_reg/NET0131  ;
	input \g2924_reg/NET0131  ;
	input \g2929_reg/NET0131  ;
	input \g2933_reg/NET0131  ;
	input \g2934_reg/NET0131  ;
	input \g2935_reg/NET0131  ;
	input \g2938_reg/NET0131  ;
	input \g2941_reg/NET0131  ;
	input \g2944_reg/NET0131  ;
	input \g2947_reg/NET0131  ;
	input \g2950_reg/NET0131  ;
	input \g2953_reg/NET0131  ;
	input \g2956_reg/NET0131  ;
	input \g2959_reg/NET0131  ;
	input \g2962_reg/NET0131  ;
	input \g2963_reg/NET0131  ;
	input \g2966_reg/NET0131  ;
	input \g2969_reg/NET0131  ;
	input \g2972_reg/NET0131  ;
	input \g2975_reg/NET0131  ;
	input \g2978_reg/NET0131  ;
	input \g2981_reg/NET0131  ;
	input \g2984_reg/NET0131  ;
	input \g2985_reg/NET0131  ;
	input \g2986_reg/NET0131  ;
	input \g2987_reg/NET0131  ;
	input \g298_reg/NET0131  ;
	input \g2990_reg/NET0131  ;
	input \g2991_reg/NET0131  ;
	input \g2992_reg/NET0131  ;
	input \g2993_reg/NET0131  ;
	input \g2997_reg/NET0131  ;
	input \g2998_reg/NET0131  ;
	input \g299_reg/NET0131  ;
	input \g3002_reg/NET0131  ;
	input \g3006_reg/NET0131  ;
	input \g3010_reg/NET0131  ;
	input \g3013_reg/NET0131  ;
	input \g3018_reg/NET0131  ;
	input \g3024_reg/NET0131  ;
	input \g3028_reg/NET0131  ;
	input \g3032_reg/NET0131  ;
	input \g3036_reg/NET0131  ;
	input \g3043_reg/NET0131  ;
	input \g3044_reg/NET0131  ;
	input \g3045_reg/NET0131  ;
	input \g3046_reg/NET0131  ;
	input \g3047_reg/NET0131  ;
	input \g3048_reg/NET0131  ;
	input \g3049_reg/NET0131  ;
	input \g3050_reg/NET0131  ;
	input \g3051_reg/NET0131  ;
	input \g3052_reg/NET0131  ;
	input \g3053_reg/NET0131  ;
	input \g3054_reg/NET0131  ;
	input \g3055_reg/NET0131  ;
	input \g3056_reg/NET0131  ;
	input \g3057_reg/NET0131  ;
	input \g3058_reg/NET0131  ;
	input \g3059_reg/NET0131  ;
	input \g305_reg/NET0131  ;
	input \g3060_reg/NET0131  ;
	input \g3061_reg/NET0131  ;
	input \g3062_reg/NET0131  ;
	input \g3063_reg/NET0131  ;
	input \g3064_reg/NET0131  ;
	input \g3065_reg/NET0131  ;
	input \g3066_reg/NET0131  ;
	input \g3067_reg/NET0131  ;
	input \g3068_reg/NET0131  ;
	input \g3069_reg/NET0131  ;
	input \g3070_reg/NET0131  ;
	input \g3071_reg/NET0131  ;
	input \g3072_reg/NET0131  ;
	input \g3073_reg/NET0131  ;
	input \g3074_reg/NET0131  ;
	input \g3075_reg/NET0131  ;
	input \g3076_reg/NET0131  ;
	input \g3077_reg/NET0131  ;
	input \g3078_reg/NET0131  ;
	input \g3079_reg/NET0131  ;
	input \g3080_reg/NET0131  ;
	input \g3083_reg/NET0131  ;
	input \g3097_reg/NET0131  ;
	input \g3110_reg/NET0131  ;
	input \g3114_reg/NET0131  ;
	input \g3120_reg/NET0131  ;
	input \g312_reg/NET0131  ;
	input \g3139_reg/NET0131  ;
	input \g313_reg/NET0131  ;
	input \g314_reg/NET0131  ;
	input \g315_reg/NET0131  ;
	input \g316_reg/NET0131  ;
	input \g317_reg/NET0131  ;
	input \g318_reg/NET0131  ;
	input \g319_reg/NET0131  ;
	input \g320_reg/NET0131  ;
	input \g321_reg/NET0131  ;
	input \g3229_pad  ;
	input \g322_reg/NET0131  ;
	input \g3230_pad  ;
	input \g3231_pad  ;
	input \g3233_pad  ;
	input \g3234_pad  ;
	input \g323_reg/NET0131  ;
	input \g324_reg/NET0131  ;
	input \g343_reg/NET0131  ;
	input \g346_reg/NET0131  ;
	input \g349_reg/NET0131  ;
	input \g351_reg/NET0131  ;
	input \g353_reg/NET0131  ;
	input \g354_reg/NET0131  ;
	input \g358_reg/NET0131  ;
	input \g361_reg/NET0131  ;
	input \g364_reg/NET0131  ;
	input \g366_reg/NET0131  ;
	input \g368_reg/NET0131  ;
	input \g369_reg/NET0131  ;
	input \g373_reg/NET0131  ;
	input \g376_reg/NET0131  ;
	input \g379_reg/NET0131  ;
	input \g381_reg/NET0131  ;
	input \g383_reg/NET0131  ;
	input \g384_reg/NET0131  ;
	input \g388_reg/NET0131  ;
	input \g391_reg/NET0131  ;
	input \g394_reg/NET0131  ;
	input \g396_reg/NET0131  ;
	input \g398_reg/NET0131  ;
	input \g402_reg/NET0131  ;
	input \g403_reg/NET0131  ;
	input \g404_reg/NET0131  ;
	input \g408_reg/NET0131  ;
	input \g411_reg/NET0131  ;
	input \g414_reg/NET0131  ;
	input \g417_reg/NET0131  ;
	input \g420_reg/NET0131  ;
	input \g423_reg/NET0131  ;
	input \g426_reg/NET0131  ;
	input \g427_reg/NET0131  ;
	input \g428_reg/NET0131  ;
	input \g429_reg/NET0131  ;
	input \g432_reg/NET0131  ;
	input \g435_reg/NET0131  ;
	input \g438_reg/NET0131  ;
	input \g441_reg/NET0131  ;
	input \g444_reg/NET0131  ;
	input \g447_reg/NET0131  ;
	input \g448_reg/NET0131  ;
	input \g449_reg/NET0131  ;
	input \g451_reg/NET0131  ;
	input \g453_reg/NET0131  ;
	input \g464_reg/NET0131  ;
	input \g465_reg/NET0131  ;
	input \g468_reg/NET0131  ;
	input \g471_reg/NET0131  ;
	input \g477_reg/NET0131  ;
	input \g478_reg/NET0131  ;
	input \g479_reg/NET0131  ;
	input \g480_reg/NET0131  ;
	input \g484_reg/NET0131  ;
	input \g486_reg/NET0131  ;
	input \g487_reg/NET0131  ;
	input \g488_reg/NET0131  ;
	input \g489_reg/NET0131  ;
	input \g490_reg/NET0131  ;
	input \g493_reg/NET0131  ;
	input \g496_reg/NET0131  ;
	input \g499_reg/NET0131  ;
	input \g506_reg/NET0131  ;
	input \g507_reg/NET0131  ;
	input \g51_pad  ;
	input \g524_reg/NET0131  ;
	input \g525_reg/NET0131  ;
	input \g529_reg/NET0131  ;
	input \g530_reg/NET0131  ;
	input \g531_reg/NET0131  ;
	input \g532_reg/NET0131  ;
	input \g533_reg/NET0131  ;
	input \g534_reg/NET0131  ;
	input \g536_reg/NET0131  ;
	input \g537_reg/NET0131  ;
	input \g5388_pad  ;
	input \g538_reg/NET0131  ;
	input \g541_reg/NET0131  ;
	input \g542_reg/NET0131  ;
	input \g544_reg/NET0131  ;
	input \g548_reg/NET0131  ;
	input \g559_reg/NET0131  ;
	input \g563_pad  ;
	input \g5657_pad  ;
	input \g565_reg/NET0131  ;
	input \g567_reg/NET0131  ;
	input \g569_reg/NET0131  ;
	input \g571_reg/NET0131  ;
	input \g573_reg/NET0131  ;
	input \g575_reg/NET0131  ;
	input \g576_reg/NET0131  ;
	input \g577_reg/NET0131  ;
	input \g578_reg/NET0131  ;
	input \g579_reg/NET0131  ;
	input \g580_reg/NET0131  ;
	input \g581_reg/NET0131  ;
	input \g582_reg/NET0131  ;
	input \g583_reg/NET0131  ;
	input \g584_reg/NET0131  ;
	input \g585_reg/NET0131  ;
	input \g586_reg/NET0131  ;
	input \g587_reg/NET0131  ;
	input \g590_reg/NET0131  ;
	input \g593_reg/NET0131  ;
	input \g596_reg/NET0131  ;
	input \g599_reg/NET0131  ;
	input \g602_reg/NET0131  ;
	input \g605_reg/NET0131  ;
	input \g608_reg/NET0131  ;
	input \g611_reg/NET0131  ;
	input \g614_reg/NET0131  ;
	input \g617_reg/NET0131  ;
	input \g620_reg/NET0131  ;
	input \g698_reg/NET0131  ;
	input \g699_reg/NET0131  ;
	input \g700_reg/NET0131  ;
	input \g701_reg/NET0131  ;
	input \g702_reg/NET0131  ;
	input \g703_reg/NET0131  ;
	input \g704_reg/NET0131  ;
	input \g705_reg/NET0131  ;
	input \g706_reg/NET0131  ;
	input \g707_reg/NET0131  ;
	input \g708_reg/NET0131  ;
	input \g709_reg/NET0131  ;
	input \g710_reg/NET0131  ;
	input \g711_reg/NET0131  ;
	input \g712_reg/NET0131  ;
	input \g713_reg/NET0131  ;
	input \g714_reg/NET0131  ;
	input \g715_reg/NET0131  ;
	input \g716_reg/NET0131  ;
	input \g717_reg/NET0131  ;
	input \g718_reg/NET0131  ;
	input \g719_reg/NET0131  ;
	input \g720_reg/NET0131  ;
	input \g721_reg/NET0131  ;
	input \g722_reg/NET0131  ;
	input \g723_reg/NET0131  ;
	input \g724_reg/NET0131  ;
	input \g725_reg/NET0131  ;
	input \g726_reg/NET0131  ;
	input \g727_reg/NET0131  ;
	input \g728_reg/NET0131  ;
	input \g729_reg/NET0131  ;
	input \g730_reg/NET0131  ;
	input \g731_reg/NET0131  ;
	input \g732_reg/NET0131  ;
	input \g733_reg/NET0131  ;
	input \g734_reg/NET0131  ;
	input \g735_reg/NET0131  ;
	input \g736_reg/NET0131  ;
	input \g737_reg/NET0131  ;
	input \g738_reg/NET0131  ;
	input \g739_reg/NET0131  ;
	input \g785_reg/NET0131  ;
	input \g789_reg/NET0131  ;
	input \g793_reg/NET0131  ;
	input \g7961_pad  ;
	input \g797_reg/NET0131  ;
	input \g801_reg/NET0131  ;
	input \g805_reg/NET0131  ;
	input \g809_reg/NET0131  ;
	input \g813_reg/NET0131  ;
	input \g817_reg/NET0131  ;
	input \g818_reg/NET0131  ;
	input \g819_reg/NET0131  ;
	input \g820_reg/NET0131  ;
	input \g821_reg/NET0131  ;
	input \g822_reg/NET0131  ;
	input \g8259_pad  ;
	input \g8260_pad  ;
	input \g8261_pad  ;
	input \g8262_pad  ;
	input \g8263_pad  ;
	input \g8264_pad  ;
	input \g8265_pad  ;
	input \g8266_pad  ;
	input \g8268_pad  ;
	input \g8269_pad  ;
	input \g8270_pad  ;
	input \g8271_pad  ;
	input \g8272_pad  ;
	input \g8273_pad  ;
	input \g8274_pad  ;
	input \g8275_pad  ;
	input \g829_reg/NET0131  ;
	input \g830_reg/NET0131  ;
	input \g831_reg/NET0131  ;
	input \g832_reg/NET0131  ;
	input \g833_reg/NET0131  ;
	input \g834_reg/NET0131  ;
	input \g835_reg/NET0131  ;
	input \g836_reg/NET0131  ;
	input \g837_reg/NET0131  ;
	input \g838_reg/NET0131  ;
	input \g839_reg/NET0131  ;
	input \g840_reg/NET0131  ;
	input \g841_reg/NET0131  ;
	input \g842_reg/NET0131  ;
	input \g843_reg/NET0131  ;
	input \g844_reg/NET0131  ;
	input \g845_reg/NET0131  ;
	input \g846_reg/NET0131  ;
	input \g847_reg/NET0131  ;
	input \g848_reg/NET0131  ;
	input \g849_reg/NET0131  ;
	input \g850_reg/NET0131  ;
	input \g851_reg/NET0131  ;
	input \g852_reg/NET0131  ;
	input \g856_reg/NET0131  ;
	input \g857_reg/NET0131  ;
	input \g858_reg/NET0131  ;
	input \g859_reg/NET0131  ;
	input \g860_reg/NET0131  ;
	input \g861_reg/NET0131  ;
	input \g862_reg/NET0131  ;
	input \g863_reg/NET0131  ;
	input \g864_reg/NET0131  ;
	input \g865_reg/NET0131  ;
	input \g866_reg/NET0131  ;
	input \g867_reg/NET0131  ;
	input \g873_reg/NET0131  ;
	input \g876_reg/NET0131  ;
	input \g879_reg/NET0131  ;
	input \g882_reg/NET0131  ;
	input \g885_reg/NET0131  ;
	input \g888_reg/NET0131  ;
	input \g891_reg/NET0131  ;
	input \g894_reg/NET0131  ;
	input \g897_reg/NET0131  ;
	input \g900_reg/NET0131  ;
	input \g903_reg/NET0131  ;
	input \g906_reg/NET0131  ;
	input \g909_reg/NET0131  ;
	input \g912_reg/NET0131  ;
	input \g915_reg/NET0131  ;
	input \g918_reg/NET0131  ;
	input \g921_reg/NET0131  ;
	input \g924_reg/NET0131  ;
	input \g927_reg/NET0131  ;
	input \g930_reg/NET0131  ;
	input \g933_reg/NET0131  ;
	input \g936_reg/NET0131  ;
	input \g939_reg/NET0131  ;
	input \g942_reg/NET0131  ;
	input \g945_reg/NET0131  ;
	input \g948_reg/NET0131  ;
	input \g951_reg/NET0131  ;
	input \g954_reg/NET0131  ;
	input \g957_reg/NET0131  ;
	input \g960_reg/NET0131  ;
	input \g966_reg/NET0131  ;
	input \g968_reg/NET0131  ;
	input \g970_reg/NET0131  ;
	input \g972_reg/NET0131  ;
	input \g974_reg/NET0131  ;
	input \g976_reg/NET0131  ;
	input \g978_reg/NET0131  ;
	input \g97_reg/NET0131  ;
	input \g985_reg/NET0131  ;
	input \g986_reg/NET0131  ;
	input \g992_reg/NET0131  ;
	input \g999_reg/NET0131  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g101_reg/P0001  ;
	output \g105_reg/P0001  ;
	output \g109_reg/P0001  ;
	output \g1138_reg/P0001  ;
	output \g113_reg/P0001  ;
	output \g1140_reg/P0001  ;
	output \g117_reg/P0001  ;
	output \g121_reg/P0001  ;
	output \g125_reg/P0001  ;
	output \g1471_reg/P0001  ;
	output \g1476_reg/P0001  ;
	output \g1481_reg/P0001  ;
	output \g1486_reg/P0001  ;
	output \g1491_reg/P0001  ;
	output \g1496_reg/P0001  ;
	output \g1501_reg/P0001  ;
	output \g1506_reg/P0001  ;
	output \g16496_pad  ;
	output \g1660_reg/P0001  ;
	output \g1662_reg/P0001  ;
	output \g1664_reg/P0001  ;
	output \g1666_reg/P0001  ;
	output \g1668_reg/P0001  ;
	output \g1670_reg/P0001  ;
	output \g1672_reg/P0001  ;
	output \g18/_0_  ;
	output \g1832_reg/P0001  ;
	output \g1834_reg/P0001  ;
	output \g2165_reg/P0001  ;
	output \g2170_reg/P0001  ;
	output \g2175_reg/P0001  ;
	output \g2180_reg/P0001  ;
	output \g2185_reg/P0001  ;
	output \g2190_reg/P0001  ;
	output \g2195_reg/P0001  ;
	output \g2200_reg/P0001  ;
	output \g2354_reg/P0001  ;
	output \g2356_reg/P0001  ;
	output \g2358_reg/P0001  ;
	output \g2360_reg/P0001  ;
	output \g2362_reg/P0001  ;
	output \g2364_reg/P0001  ;
	output \g2366_reg/P0001  ;
	output \g2526_reg/P0001  ;
	output \g2528_reg/P0001  ;
	output \g25489_pad  ;
	output \g279_reg/P0001  ;
	output \g281_reg/P0001  ;
	output \g283_reg/P0001  ;
	output \g285_reg/P0001  ;
	output \g2879_reg/NET0131_syn_2  ;
	output \g287_reg/P0001  ;
	output \g289_reg/P0001  ;
	output \g291_reg/P0001  ;
	output \g451_reg/P0001  ;
	output \g453_reg/P0001  ;
	output \g59421/_3_  ;
	output \g59425/_1_  ;
	output \g59435/_0_  ;
	output \g59436/_0_  ;
	output \g59441/_3_  ;
	output \g59442/_0_  ;
	output \g59445/_0_  ;
	output \g59453/_0_  ;
	output \g59462/_3_  ;
	output \g59466/_3_  ;
	output \g59467/_3_  ;
	output \g59468/_3_  ;
	output \g59469/_3_  ;
	output \g59470/_3_  ;
	output \g59471/_3_  ;
	output \g59472/_3_  ;
	output \g59473/_3_  ;
	output \g59489/_0_  ;
	output \g59498/_0_  ;
	output \g59499/_0_  ;
	output \g59500/_0_  ;
	output \g59502/_2_  ;
	output \g59503/_0_  ;
	output \g59505/_2_  ;
	output \g59507/_0_  ;
	output \g59508/_0_  ;
	output \g59533/_3_  ;
	output \g59534/_3_  ;
	output \g59535/_3_  ;
	output \g59536/_3_  ;
	output \g59537/_3_  ;
	output \g59538/_3_  ;
	output \g59539/_3_  ;
	output \g59540/_3_  ;
	output \g59548/_0_  ;
	output \g59550/_0_  ;
	output \g59551/_0_  ;
	output \g59552/_0_  ;
	output \g59554/_0_  ;
	output \g59555/_0_  ;
	output \g59556/_0_  ;
	output \g59557/_0_  ;
	output \g59558/_0_  ;
	output \g59559/_0_  ;
	output \g59560/_0_  ;
	output \g59561/_0_  ;
	output \g59639/_0_  ;
	output \g59694/_2_  ;
	output \g59695/_0_  ;
	output \g59697/_2_  ;
	output \g59698/_0_  ;
	output \g59699/_0_  ;
	output \g59700/_0_  ;
	output \g59705/_0_  ;
	output \g59706/_0_  ;
	output \g59707/_0_  ;
	output \g59708/_0_  ;
	output \g59709/_0_  ;
	output \g59710/_0_  ;
	output \g59711/_0_  ;
	output \g59712/_0_  ;
	output \g59713/_0_  ;
	output \g59714/_0_  ;
	output \g59715/_0_  ;
	output \g59716/_0_  ;
	output \g59717/_0_  ;
	output \g59718/_0_  ;
	output \g59719/_0_  ;
	output \g59720/_0_  ;
	output \g59721/_0_  ;
	output \g59722/_0_  ;
	output \g59723/_0_  ;
	output \g59724/_0_  ;
	output \g59725/_0_  ;
	output \g59726/_0_  ;
	output \g59727/_0_  ;
	output \g59728/_0_  ;
	output \g59729/_0_  ;
	output \g59730/_0_  ;
	output \g59731/_0_  ;
	output \g59732/_0_  ;
	output \g59733/_0_  ;
	output \g59734/_0_  ;
	output \g59735/_0_  ;
	output \g59736/_0_  ;
	output \g59737/_0_  ;
	output \g59738/_0_  ;
	output \g59739/_0_  ;
	output \g59740/_0_  ;
	output \g59741/_0_  ;
	output \g59742/_0_  ;
	output \g59743/_0_  ;
	output \g59744/_0_  ;
	output \g59745/_0_  ;
	output \g59747/_0_  ;
	output \g59748/_0_  ;
	output \g59749/_0_  ;
	output \g59750/_0_  ;
	output \g59751/_0_  ;
	output \g59752/_0_  ;
	output \g59753/_0_  ;
	output \g59754/_0_  ;
	output \g59755/_0_  ;
	output \g59756/_0_  ;
	output \g59757/_0_  ;
	output \g59758/_0_  ;
	output \g59759/_0_  ;
	output \g59760/_0_  ;
	output \g59761/_0_  ;
	output \g59762/_0_  ;
	output \g59763/_0_  ;
	output \g59764/_0_  ;
	output \g59765/_0_  ;
	output \g59766/_0_  ;
	output \g59915/_0_  ;
	output \g59952/_2_  ;
	output \g60046/_0_  ;
	output \g60048/_0_  ;
	output \g60049/_0_  ;
	output \g60051/_0_  ;
	output \g60063/_0_  ;
	output \g60103/_0_  ;
	output \g60104/_0_  ;
	output \g60105/_0_  ;
	output \g60107/_2_  ;
	output \g60108/_0_  ;
	output \g60109/_0_  ;
	output \g60110/_0_  ;
	output \g60112/_2_  ;
	output \g60119/_0_  ;
	output \g60120/_0_  ;
	output \g60121/_0_  ;
	output \g60122/_0_  ;
	output \g60123/_0_  ;
	output \g60124/_0_  ;
	output \g60126/_0_  ;
	output \g60127/_0_  ;
	output \g60128/_0_  ;
	output \g60129/_0_  ;
	output \g60130/_0_  ;
	output \g60135/_0_  ;
	output \g60136/_0_  ;
	output \g60137/_0_  ;
	output \g60138/_0_  ;
	output \g60139/_0_  ;
	output \g60143/_3_  ;
	output \g60144/_0_  ;
	output \g60145/_0_  ;
	output \g60339/_0_  ;
	output \g60404/_0_  ;
	output \g60427/_0_  ;
	output \g60428/_0_  ;
	output \g60429/_0_  ;
	output \g60434/_0_  ;
	output \g60435/_0_  ;
	output \g60437/_0_  ;
	output \g60438/_0_  ;
	output \g60439/_0_  ;
	output \g60440/_0_  ;
	output \g60441/_0_  ;
	output \g60448/_0_  ;
	output \g60451/_0_  ;
	output \g60452/_0_  ;
	output \g60453/_0_  ;
	output \g60459/_0_  ;
	output \g60460/_0_  ;
	output \g60523/_0_  ;
	output \g60534/_0_  ;
	output \g60535/_0_  ;
	output \g60536/_0_  ;
	output \g60585/_0_  ;
	output \g60586/_0_  ;
	output \g60587/_0_  ;
	output \g60588/_0_  ;
	output \g60591/_0_  ;
	output \g60592/_0_  ;
	output \g60599/_0_  ;
	output \g60601/_0_  ;
	output \g60602/_0_  ;
	output \g60603/_0_  ;
	output \g60604/_0_  ;
	output \g60605/_0_  ;
	output \g60606/_0_  ;
	output \g60607/_0_  ;
	output \g60608/_0_  ;
	output \g60609/_0_  ;
	output \g60613/_0_  ;
	output \g60614/_0_  ;
	output \g60615/_0_  ;
	output \g60694/_0_  ;
	output \g60708/_0_  ;
	output \g60709/_0_  ;
	output \g60710/_0_  ;
	output \g60785/_0_  ;
	output \g60787/_0_  ;
	output \g60788/_0_  ;
	output \g60799/_0_  ;
	output \g60801/_0_  ;
	output \g60802/_0_  ;
	output \g60803/_1__syn_2  ;
	output \g60805/_1__syn_2  ;
	output \g60806/_1__syn_2  ;
	output \g60808/_0_  ;
	output \g60810/_0_  ;
	output \g60811/_0_  ;
	output \g60825/_3_  ;
	output \g60896/_0_  ;
	output \g60980/_0_  ;
	output \g60981/_0_  ;
	output \g60985/_0_  ;
	output \g60986/_0_  ;
	output \g61012/_0_  ;
	output \g61013/_0_  ;
	output \g61015/_0_  ;
	output \g61017/_0_  ;
	output \g61122/_0_  ;
	output \g61123/_0_  ;
	output \g61124/_0_  ;
	output \g61125/_0_  ;
	output \g61222/_0_  ;
	output \g61223/_0_  ;
	output \g61224/_0_  ;
	output \g61225/_0_  ;
	output \g61228/_0_  ;
	output \g61229/_0_  ;
	output \g61230/_0_  ;
	output \g61231/_0_  ;
	output \g61281/_0_  ;
	output \g61293/_1_  ;
	output \g61307/_0__syn_2  ;
	output \g61309/_0__syn_2  ;
	output \g61310/_0__syn_2  ;
	output \g61311/_1_  ;
	output \g61312/_1_  ;
	output \g61313/_1_  ;
	output \g61324/_1_  ;
	output \g61325/_1_  ;
	output \g61326/_1_  ;
	output \g61328/_1_  ;
	output \g61329/_1_  ;
	output \g61330/_1_  ;
	output \g61332/_1_  ;
	output \g61333/_1_  ;
	output \g61334/_1_  ;
	output \g61335/_1_  ;
	output \g61336/_0_  ;
	output \g61338/_0_  ;
	output \g61339/_0_  ;
	output \g61340/_0_  ;
	output \g61377/_1_  ;
	output \g61378/_1_  ;
	output \g61379/_1_  ;
	output \g61388/_1_  ;
	output \g61391/_0_  ;
	output \g61394/_1_  ;
	output \g61395/_1_  ;
	output \g61396/_1_  ;
	output \g61398/_1_  ;
	output \g61399/_1_  ;
	output \g61421/_1_  ;
	output \g61422/_1_  ;
	output \g61423/_1_  ;
	output \g61524/_0_  ;
	output \g61525/_0_  ;
	output \g61526/_0_  ;
	output \g61527/_0_  ;
	output \g61528/_0_  ;
	output \g61529/_0_  ;
	output \g61530/_0_  ;
	output \g61531/_0_  ;
	output \g61532/_0_  ;
	output \g61533/_0_  ;
	output \g61534/_0_  ;
	output \g61535/_0_  ;
	output \g61536/_0_  ;
	output \g61537/_0_  ;
	output \g61538/_0_  ;
	output \g61539/_0_  ;
	output \g61540/_0_  ;
	output \g61541/_0_  ;
	output \g61542/_0_  ;
	output \g61543/_0_  ;
	output \g61544/_0_  ;
	output \g61545/_0_  ;
	output \g61546/_0_  ;
	output \g61547/_0_  ;
	output \g61548/_0_  ;
	output \g61549/_0_  ;
	output \g61550/_0_  ;
	output \g61551/_0_  ;
	output \g61552/_0_  ;
	output \g61553/_0_  ;
	output \g61554/_0_  ;
	output \g61555/_0_  ;
	output \g61556/_0_  ;
	output \g61557/_0_  ;
	output \g61558/_0_  ;
	output \g61559/_0_  ;
	output \g61560/_0_  ;
	output \g61561/_0_  ;
	output \g61562/_0_  ;
	output \g61563/_0_  ;
	output \g61564/_0_  ;
	output \g61565/_0_  ;
	output \g61566/_0_  ;
	output \g61620/_0_  ;
	output \g61621/_0_  ;
	output \g61622/_0_  ;
	output \g61623/_0_  ;
	output \g61753/_0_  ;
	output \g61764/_0_  ;
	output \g61786/_0_  ;
	output \g61795/_0_  ;
	output \g61801/_0_  ;
	output \g61803/_0_  ;
	output \g61808/_0_  ;
	output \g61848/_0_  ;
	output \g61850/_0_  ;
	output \g61851/_0_  ;
	output \g62097/_0_  ;
	output \g62102/_0_  ;
	output \g62115/_0_  ;
	output \g62119/_0_  ;
	output \g62130/_1_  ;
	output \g62131/_0_  ;
	output \g62132/_0_  ;
	output \g62139/_1_  ;
	output \g62140/_1_  ;
	output \g62141/_1_  ;
	output \g62144/_0_  ;
	output \g62145/_0_  ;
	output \g62146/_0_  ;
	output \g62147/_0_  ;
	output \g62150/_0_  ;
	output \g62151/_1_  ;
	output \g62152/_0_  ;
	output \g62153/_1_  ;
	output \g62156/_1_  ;
	output \g62157/_0_  ;
	output \g62159/_0_  ;
	output \g62161/_0_  ;
	output \g62187/_1_  ;
	output \g62190/_1_  ;
	output \g62191/_1_  ;
	output \g62192/_1_  ;
	output \g62194/_1_  ;
	output \g62195/_1_  ;
	output \g62196/_1_  ;
	output \g62203/_0_  ;
	output \g62204/_1_  ;
	output \g62207/_0__syn_2  ;
	output \g62208/_1_  ;
	output \g62209/_1_  ;
	output \g62210/_1_  ;
	output \g62211/_1_  ;
	output \g62212/_1_  ;
	output \g62217/_0_  ;
	output \g62286/_0_  ;
	output \g62287/_0_  ;
	output \g62288/_0_  ;
	output \g62289/_0_  ;
	output \g62290/_0_  ;
	output \g62291/_0_  ;
	output \g62292/_0_  ;
	output \g62435/_0_  ;
	output \g62436/_0_  ;
	output \g62439/_0_  ;
	output \g62456/_0_  ;
	output \g62486/_1_  ;
	output \g62492/_1_  ;
	output \g62494/_0_  ;
	output \g62495/_1_  ;
	output \g62497/_0_  ;
	output \g62537/_0_  ;
	output \g62544/_0_  ;
	output \g62546/_0_  ;
	output \g62547/_0_  ;
	output \g62549/_3_  ;
	output \g62552/_0_  ;
	output \g62554/_0_  ;
	output \g62555/_0_  ;
	output \g62556/_0_  ;
	output \g62558/_0_  ;
	output \g62559/_0_  ;
	output \g62561/_0_  ;
	output \g62562/_0_  ;
	output \g62566/_0_  ;
	output \g62567/_0_  ;
	output \g62568/_0_  ;
	output \g62569/_0_  ;
	output \g62570/_0_  ;
	output \g62571/_0_  ;
	output \g62572/_0_  ;
	output \g62573/_0_  ;
	output \g62574/_0_  ;
	output \g62575/_0_  ;
	output \g62576/_0_  ;
	output \g62577/_0_  ;
	output \g62578/_0_  ;
	output \g62579/_0_  ;
	output \g62580/_0_  ;
	output \g62581/_0_  ;
	output \g62582/_0_  ;
	output \g62583/_0_  ;
	output \g62584/_0_  ;
	output \g62585/_0_  ;
	output \g62586/_0_  ;
	output \g62587/_0_  ;
	output \g62588/_0_  ;
	output \g62589/_0_  ;
	output \g62590/_0_  ;
	output \g62591/_0_  ;
	output \g62592/_0_  ;
	output \g62593/_0_  ;
	output \g62594/_0_  ;
	output \g62595/_0_  ;
	output \g62596/_0_  ;
	output \g62597/_0_  ;
	output \g62602/_0_  ;
	output \g62607/_0_  ;
	output \g62608/_0_  ;
	output \g62609/_0_  ;
	output \g62619/_0_  ;
	output \g62620/_0_  ;
	output \g62621/_0_  ;
	output \g62622/_0_  ;
	output \g62623/_0_  ;
	output \g62624/_0_  ;
	output \g62626/_0_  ;
	output \g62627/_0_  ;
	output \g62628/_0_  ;
	output \g62629/_0_  ;
	output \g62630/_0_  ;
	output \g62631/_0_  ;
	output \g62632/_0_  ;
	output \g62633/_0_  ;
	output \g62634/_0_  ;
	output \g62635/_0_  ;
	output \g62636/_0_  ;
	output \g62637/_0_  ;
	output \g62638/_0_  ;
	output \g62639/_0_  ;
	output \g62640/_0_  ;
	output \g62641/_0_  ;
	output \g62642/_0_  ;
	output \g62643/_0_  ;
	output \g62644/_0_  ;
	output \g62645/_0_  ;
	output \g62646/_0_  ;
	output \g62647/_0_  ;
	output \g62648/_0_  ;
	output \g62649/_0_  ;
	output \g62650/_0_  ;
	output \g62651/_0_  ;
	output \g62652/_0_  ;
	output \g62653/_0_  ;
	output \g62654/_0_  ;
	output \g62655/_0_  ;
	output \g62656/_0_  ;
	output \g62657/_0_  ;
	output \g62658/_0_  ;
	output \g62659/_0_  ;
	output \g62660/_0_  ;
	output \g62661/_0_  ;
	output \g62674/_0_  ;
	output \g62682/_0_  ;
	output \g62683/_0_  ;
	output \g62689/_0_  ;
	output \g62690/_0_  ;
	output \g62691/_0_  ;
	output \g62694/_0_  ;
	output \g62695/_0_  ;
	output \g62696/_0_  ;
	output \g62698/_0_  ;
	output \g62699/_0_  ;
	output \g62700/_0_  ;
	output \g62723/_0_  ;
	output \g62724/_0_  ;
	output \g62725/_0_  ;
	output \g62726/_0_  ;
	output \g62727/_0_  ;
	output \g62728/_0_  ;
	output \g62735/_0_  ;
	output \g62736/_0_  ;
	output \g62737/_0_  ;
	output \g62738/_0_  ;
	output \g62739/_0_  ;
	output \g62740/_0_  ;
	output \g62754/_0_  ;
	output \g62762/_0_  ;
	output \g62763/_0_  ;
	output \g62764/_0_  ;
	output \g62780/_0_  ;
	output \g62781/_0_  ;
	output \g62785/_0_  ;
	output \g62786/_0_  ;
	output \g62787/_0_  ;
	output \g62791/_0_  ;
	output \g62792/_0_  ;
	output \g62794/_0_  ;
	output \g62804/_0_  ;
	output \g62806/_0_  ;
	output \g62807/_0_  ;
	output \g62811/_0_  ;
	output \g62968/_0_  ;
	output \g63005/_0_  ;
	output \g63041/_0_  ;
	output \g63116/_0_  ;
	output \g63157/_0_  ;
	output \g63164/_0_  ;
	output \g63170/_0_  ;
	output \g63189/_0_  ;
	output \g63202/_0_  ;
	output \g63206/_0_  ;
	output \g63207/_0_  ;
	output \g63265/_0_  ;
	output \g63266/_0_  ;
	output \g63269/_0_  ;
	output \g63271/_0_  ;
	output \g63272/_0_  ;
	output \g63273/_0_  ;
	output \g63274/_0_  ;
	output \g63275/_0_  ;
	output \g63276/_0_  ;
	output \g63277/_0_  ;
	output \g63278/_0_  ;
	output \g63280/_0_  ;
	output \g63281/_0_  ;
	output \g63282/_0_  ;
	output \g63283/_0_  ;
	output \g63284/_0_  ;
	output \g63285/_0_  ;
	output \g63286/_0_  ;
	output \g63287/_0_  ;
	output \g63288/_0_  ;
	output \g63289/_0_  ;
	output \g63290/_0_  ;
	output \g63292/_0_  ;
	output \g63293/_0_  ;
	output \g63294/_0_  ;
	output \g63295/_0_  ;
	output \g63296/_0_  ;
	output \g63297/_0_  ;
	output \g63298/_0_  ;
	output \g63299/_0_  ;
	output \g63302/_0_  ;
	output \g63303/_0_  ;
	output \g63304/_0_  ;
	output \g63305/_0_  ;
	output \g63306/_0_  ;
	output \g63307/_0_  ;
	output \g63308/_0_  ;
	output \g63309/_0_  ;
	output \g63310/_0_  ;
	output \g63311/_0_  ;
	output \g63312/_0_  ;
	output \g63313/_0_  ;
	output \g63314/_0_  ;
	output \g63315/_0_  ;
	output \g63316/_0_  ;
	output \g63317/_0_  ;
	output \g63318/_0_  ;
	output \g63319/_0_  ;
	output \g63320/_0_  ;
	output \g63321/_0_  ;
	output \g63322/_0_  ;
	output \g63323/_0_  ;
	output \g63324/_0_  ;
	output \g63325/_0_  ;
	output \g63326/_0_  ;
	output \g63327/_0_  ;
	output \g63328/_0_  ;
	output \g63329/_0_  ;
	output \g63330/_0_  ;
	output \g63331/_0_  ;
	output \g63339/_0_  ;
	output \g63505/_0_  ;
	output \g63525/_0_  ;
	output \g63543/_1_  ;
	output \g63602/_0_  ;
	output \g63653/_0_  ;
	output \g63663/_1_  ;
	output \g63677/_0_  ;
	output \g63694/_0_  ;
	output \g63729/_0_  ;
	output \g63766/_0_  ;
	output \g63771/_1_  ;
	output \g63773/_1_  ;
	output \g63784/_1_  ;
	output \g63964/_0_  ;
	output \g63965/_0_  ;
	output \g63966/_0_  ;
	output \g63967/_0_  ;
	output \g64257/_1_  ;
	output \g64266/_0_  ;
	output \g64275/_0_  ;
	output \g64400/_0_  ;
	output \g64416/_0_  ;
	output \g64470/_3_  ;
	output \g64473/_0_  ;
	output \g64474/_0_  ;
	output \g64475/_0_  ;
	output \g64479/_0_  ;
	output \g64480/_0_  ;
	output \g64481/_0_  ;
	output \g64483/_0_  ;
	output \g64484/_0_  ;
	output \g64485/_0_  ;
	output \g64486/_0_  ;
	output \g64493/_0_  ;
	output \g64494/_0_  ;
	output \g64495/_0_  ;
	output \g64496/_0_  ;
	output \g64505/_3_  ;
	output \g64507/_0_  ;
	output \g64508/_0_  ;
	output \g64510/_0_  ;
	output \g64511/_0_  ;
	output \g64544/_0_  ;
	output \g64545/_0_  ;
	output \g64546/_0_  ;
	output \g64639/_0_  ;
	output \g64641/_0_  ;
	output \g64642/_0_  ;
	output \g64645/_0_  ;
	output \g64650/_0_  ;
	output \g64737/_0_  ;
	output \g64738/_0_  ;
	output \g65066/_0_  ;
	output \g65070/_0_  ;
	output \g65090/_0_  ;
	output \g65102/_0_  ;
	output \g65102/_3_  ;
	output \g65126/_3_  ;
	output \g65147/_3_  ;
	output \g65163/_0_  ;
	output \g65176/_3_  ;
	output \g65178/_0_  ;
	output \g65182/_0_  ;
	output \g65190/_1_  ;
	output \g65191/_0_  ;
	output \g65196/_0_  ;
	output \g65268/_0_  ;
	output \g65275/_0_  ;
	output \g65290/_0_  ;
	output \g65290/_3_  ;
	output \g65291/_0_  ;
	output \g65292/_0_  ;
	output \g65298/_0_  ;
	output \g65298/_3_  ;
	output \g65314/_0_  ;
	output \g65314/_3_  ;
	output \g65319/_3_  ;
	output \g65335/_0_  ;
	output \g65342/_0_  ;
	output \g65348/_0_  ;
	output \g65422/_0_  ;
	output \g65465/_1_  ;
	output \g65469/_1_  ;
	output \g65478/_1_  ;
	output \g65507/_0_  ;
	output \g65548/_0_  ;
	output \g65699/_1_  ;
	output \g65713/_1_  ;
	output \g65835/_0_  ;
	output \g65860/_0_  ;
	output \g65863/_0_  ;
	output \g66094/_1_  ;
	output \g66102/_0_  ;
	output \g66107/_0_  ;
	output \g66130/_3_  ;
	output \g66131/_3_  ;
	output \g66228/_1_  ;
	output \g66348/_1_  ;
	output \g66543/_0_  ;
	output \g66549/_1_  ;
	output \g66640/_3_  ;
	output \g66641/_3_  ;
	output \g66950/_1_  ;
	output \g67111/_0_  ;
	output \g67219/_0_  ;
	output \g67263/_0_  ;
	output \g67909/_1_  ;
	output \g68049/_0_  ;
	output \g68220/_0_  ;
	output \g68413/_0_  ;
	output \g68511/_0_  ;
	output \g68536/_0_  ;
	output \g68543/_1_  ;
	output \g68554/_0_  ;
	output \g68559/_0_  ;
	output \g70915/_0_  ;
	output \g71108/_1_  ;
	output \g71115/_2_  ;
	output \g71244_dup/_0_  ;
	output \g71368/_0_  ;
	output \g71581/_0_  ;
	output \g71720/_0_  ;
	output \g785_reg/P0001  ;
	output \g789_reg/P0001  ;
	output \g797_reg/P0001  ;
	output \g809_reg/P0001  ;
	output \g813_reg/P0001  ;
	output \g966_reg/P0001  ;
	output \g968_reg/P0001  ;
	output \g970_reg/P0001  ;
	output \g972_reg/P0001  ;
	output \g974_reg/P0001  ;
	output \g976_reg/P0001  ;
	output \g978_reg/P0001  ;
	wire _w5127_ ;
	wire _w5126_ ;
	wire _w5125_ ;
	wire _w5124_ ;
	wire _w5123_ ;
	wire _w5122_ ;
	wire _w5121_ ;
	wire _w5120_ ;
	wire _w5119_ ;
	wire _w5117_ ;
	wire _w5116_ ;
	wire _w5115_ ;
	wire _w5114_ ;
	wire _w5113_ ;
	wire _w5112_ ;
	wire _w5111_ ;
	wire _w5110_ ;
	wire _w5109_ ;
	wire _w5108_ ;
	wire _w5107_ ;
	wire _w5106_ ;
	wire _w5105_ ;
	wire _w5104_ ;
	wire _w5102_ ;
	wire _w5101_ ;
	wire _w5100_ ;
	wire _w5099_ ;
	wire _w5098_ ;
	wire _w5097_ ;
	wire _w5096_ ;
	wire _w5095_ ;
	wire _w5094_ ;
	wire _w5093_ ;
	wire _w5092_ ;
	wire _w5091_ ;
	wire _w5090_ ;
	wire _w5089_ ;
	wire _w5088_ ;
	wire _w5087_ ;
	wire _w5086_ ;
	wire _w5085_ ;
	wire _w5084_ ;
	wire _w5083_ ;
	wire _w5082_ ;
	wire _w5081_ ;
	wire _w5080_ ;
	wire _w5079_ ;
	wire _w5078_ ;
	wire _w5077_ ;
	wire _w5076_ ;
	wire _w5075_ ;
	wire _w5074_ ;
	wire _w5073_ ;
	wire _w5072_ ;
	wire _w5071_ ;
	wire _w5070_ ;
	wire _w5069_ ;
	wire _w5068_ ;
	wire _w5067_ ;
	wire _w5066_ ;
	wire _w5065_ ;
	wire _w5064_ ;
	wire _w5063_ ;
	wire _w5062_ ;
	wire _w5061_ ;
	wire _w5060_ ;
	wire _w5059_ ;
	wire _w5058_ ;
	wire _w5057_ ;
	wire _w5056_ ;
	wire _w5055_ ;
	wire _w5054_ ;
	wire _w5053_ ;
	wire _w5052_ ;
	wire _w5051_ ;
	wire _w5050_ ;
	wire _w5049_ ;
	wire _w5048_ ;
	wire _w5047_ ;
	wire _w5046_ ;
	wire _w5045_ ;
	wire _w5044_ ;
	wire _w5043_ ;
	wire _w5042_ ;
	wire _w5041_ ;
	wire _w5040_ ;
	wire _w5039_ ;
	wire _w5038_ ;
	wire _w5037_ ;
	wire _w5036_ ;
	wire _w5035_ ;
	wire _w5034_ ;
	wire _w5033_ ;
	wire _w5032_ ;
	wire _w5031_ ;
	wire _w5030_ ;
	wire _w5029_ ;
	wire _w5028_ ;
	wire _w5027_ ;
	wire _w5026_ ;
	wire _w5025_ ;
	wire _w5024_ ;
	wire _w5023_ ;
	wire _w5022_ ;
	wire _w5021_ ;
	wire _w5020_ ;
	wire _w5019_ ;
	wire _w5018_ ;
	wire _w5017_ ;
	wire _w5016_ ;
	wire _w5015_ ;
	wire _w5014_ ;
	wire _w5013_ ;
	wire _w5012_ ;
	wire _w5011_ ;
	wire _w5010_ ;
	wire _w5009_ ;
	wire _w5008_ ;
	wire _w5007_ ;
	wire _w5006_ ;
	wire _w5005_ ;
	wire _w5004_ ;
	wire _w5003_ ;
	wire _w5002_ ;
	wire _w5001_ ;
	wire _w5000_ ;
	wire _w4999_ ;
	wire _w4998_ ;
	wire _w4997_ ;
	wire _w4996_ ;
	wire _w4995_ ;
	wire _w4994_ ;
	wire _w4993_ ;
	wire _w4992_ ;
	wire _w4991_ ;
	wire _w4990_ ;
	wire _w4989_ ;
	wire _w4988_ ;
	wire _w4987_ ;
	wire _w4986_ ;
	wire _w4985_ ;
	wire _w4984_ ;
	wire _w4983_ ;
	wire _w4982_ ;
	wire _w4981_ ;
	wire _w4980_ ;
	wire _w4979_ ;
	wire _w4978_ ;
	wire _w4977_ ;
	wire _w4976_ ;
	wire _w4975_ ;
	wire _w4974_ ;
	wire _w4973_ ;
	wire _w4972_ ;
	wire _w4971_ ;
	wire _w4970_ ;
	wire _w4969_ ;
	wire _w4968_ ;
	wire _w4967_ ;
	wire _w4966_ ;
	wire _w4965_ ;
	wire _w4964_ ;
	wire _w4963_ ;
	wire _w4962_ ;
	wire _w4961_ ;
	wire _w4960_ ;
	wire _w4959_ ;
	wire _w4958_ ;
	wire _w4957_ ;
	wire _w4956_ ;
	wire _w4955_ ;
	wire _w4954_ ;
	wire _w4953_ ;
	wire _w4952_ ;
	wire _w4951_ ;
	wire _w4950_ ;
	wire _w4949_ ;
	wire _w4948_ ;
	wire _w4947_ ;
	wire _w4946_ ;
	wire _w4945_ ;
	wire _w4944_ ;
	wire _w4943_ ;
	wire _w4942_ ;
	wire _w4941_ ;
	wire _w4940_ ;
	wire _w4939_ ;
	wire _w4938_ ;
	wire _w4937_ ;
	wire _w4936_ ;
	wire _w4935_ ;
	wire _w4934_ ;
	wire _w4933_ ;
	wire _w4932_ ;
	wire _w4931_ ;
	wire _w4930_ ;
	wire _w4929_ ;
	wire _w4928_ ;
	wire _w4927_ ;
	wire _w4926_ ;
	wire _w4925_ ;
	wire _w4924_ ;
	wire _w4923_ ;
	wire _w4922_ ;
	wire _w4921_ ;
	wire _w4920_ ;
	wire _w4919_ ;
	wire _w4918_ ;
	wire _w4917_ ;
	wire _w4916_ ;
	wire _w4915_ ;
	wire _w4914_ ;
	wire _w4913_ ;
	wire _w4912_ ;
	wire _w4911_ ;
	wire _w4910_ ;
	wire _w4909_ ;
	wire _w4908_ ;
	wire _w4907_ ;
	wire _w4906_ ;
	wire _w4905_ ;
	wire _w4904_ ;
	wire _w4903_ ;
	wire _w4902_ ;
	wire _w4901_ ;
	wire _w4900_ ;
	wire _w4899_ ;
	wire _w4898_ ;
	wire _w4897_ ;
	wire _w4896_ ;
	wire _w4895_ ;
	wire _w4894_ ;
	wire _w4893_ ;
	wire _w4892_ ;
	wire _w4891_ ;
	wire _w4890_ ;
	wire _w4889_ ;
	wire _w4888_ ;
	wire _w4887_ ;
	wire _w4886_ ;
	wire _w4885_ ;
	wire _w4884_ ;
	wire _w4883_ ;
	wire _w4882_ ;
	wire _w4881_ ;
	wire _w4880_ ;
	wire _w4879_ ;
	wire _w4878_ ;
	wire _w4877_ ;
	wire _w4876_ ;
	wire _w4875_ ;
	wire _w4874_ ;
	wire _w4873_ ;
	wire _w4872_ ;
	wire _w4871_ ;
	wire _w4870_ ;
	wire _w4869_ ;
	wire _w4868_ ;
	wire _w4867_ ;
	wire _w4866_ ;
	wire _w4865_ ;
	wire _w4864_ ;
	wire _w4863_ ;
	wire _w4862_ ;
	wire _w4861_ ;
	wire _w4860_ ;
	wire _w4859_ ;
	wire _w4858_ ;
	wire _w4857_ ;
	wire _w4856_ ;
	wire _w4855_ ;
	wire _w4854_ ;
	wire _w4853_ ;
	wire _w4852_ ;
	wire _w4851_ ;
	wire _w4850_ ;
	wire _w4849_ ;
	wire _w4848_ ;
	wire _w4847_ ;
	wire _w4846_ ;
	wire _w4845_ ;
	wire _w4844_ ;
	wire _w4843_ ;
	wire _w4842_ ;
	wire _w4841_ ;
	wire _w4840_ ;
	wire _w4839_ ;
	wire _w4838_ ;
	wire _w4837_ ;
	wire _w4836_ ;
	wire _w4835_ ;
	wire _w4834_ ;
	wire _w4833_ ;
	wire _w4832_ ;
	wire _w4831_ ;
	wire _w4830_ ;
	wire _w4829_ ;
	wire _w4828_ ;
	wire _w4827_ ;
	wire _w4826_ ;
	wire _w4825_ ;
	wire _w4824_ ;
	wire _w4823_ ;
	wire _w4822_ ;
	wire _w4821_ ;
	wire _w4820_ ;
	wire _w4819_ ;
	wire _w4818_ ;
	wire _w4817_ ;
	wire _w4816_ ;
	wire _w4815_ ;
	wire _w4814_ ;
	wire _w4813_ ;
	wire _w4812_ ;
	wire _w4811_ ;
	wire _w4810_ ;
	wire _w4809_ ;
	wire _w4808_ ;
	wire _w4807_ ;
	wire _w4806_ ;
	wire _w4805_ ;
	wire _w4804_ ;
	wire _w4803_ ;
	wire _w4802_ ;
	wire _w4801_ ;
	wire _w4800_ ;
	wire _w4799_ ;
	wire _w4798_ ;
	wire _w4797_ ;
	wire _w4796_ ;
	wire _w4795_ ;
	wire _w4794_ ;
	wire _w4793_ ;
	wire _w4792_ ;
	wire _w4791_ ;
	wire _w4790_ ;
	wire _w4789_ ;
	wire _w4788_ ;
	wire _w4787_ ;
	wire _w4786_ ;
	wire _w4785_ ;
	wire _w4784_ ;
	wire _w4783_ ;
	wire _w4782_ ;
	wire _w4781_ ;
	wire _w4780_ ;
	wire _w4779_ ;
	wire _w4778_ ;
	wire _w4777_ ;
	wire _w4776_ ;
	wire _w4775_ ;
	wire _w4774_ ;
	wire _w4773_ ;
	wire _w4772_ ;
	wire _w4771_ ;
	wire _w4770_ ;
	wire _w4769_ ;
	wire _w4768_ ;
	wire _w4767_ ;
	wire _w4766_ ;
	wire _w4765_ ;
	wire _w4764_ ;
	wire _w4763_ ;
	wire _w4762_ ;
	wire _w4761_ ;
	wire _w4760_ ;
	wire _w4759_ ;
	wire _w4758_ ;
	wire _w4757_ ;
	wire _w4756_ ;
	wire _w4755_ ;
	wire _w4754_ ;
	wire _w4753_ ;
	wire _w4752_ ;
	wire _w4751_ ;
	wire _w4750_ ;
	wire _w4749_ ;
	wire _w4748_ ;
	wire _w4747_ ;
	wire _w4746_ ;
	wire _w4745_ ;
	wire _w4744_ ;
	wire _w4743_ ;
	wire _w4742_ ;
	wire _w4741_ ;
	wire _w4740_ ;
	wire _w4739_ ;
	wire _w4738_ ;
	wire _w4737_ ;
	wire _w4736_ ;
	wire _w4735_ ;
	wire _w4734_ ;
	wire _w4733_ ;
	wire _w4732_ ;
	wire _w4731_ ;
	wire _w4730_ ;
	wire _w4729_ ;
	wire _w4728_ ;
	wire _w4727_ ;
	wire _w4726_ ;
	wire _w4725_ ;
	wire _w4724_ ;
	wire _w4723_ ;
	wire _w4722_ ;
	wire _w4721_ ;
	wire _w4720_ ;
	wire _w4719_ ;
	wire _w4718_ ;
	wire _w4717_ ;
	wire _w4716_ ;
	wire _w4715_ ;
	wire _w4714_ ;
	wire _w4713_ ;
	wire _w4712_ ;
	wire _w4711_ ;
	wire _w4710_ ;
	wire _w4709_ ;
	wire _w4708_ ;
	wire _w4707_ ;
	wire _w4706_ ;
	wire _w4705_ ;
	wire _w4704_ ;
	wire _w4703_ ;
	wire _w4702_ ;
	wire _w4701_ ;
	wire _w4700_ ;
	wire _w4699_ ;
	wire _w4698_ ;
	wire _w4697_ ;
	wire _w4696_ ;
	wire _w4695_ ;
	wire _w4694_ ;
	wire _w4693_ ;
	wire _w4692_ ;
	wire _w4691_ ;
	wire _w4690_ ;
	wire _w4689_ ;
	wire _w4688_ ;
	wire _w4687_ ;
	wire _w4686_ ;
	wire _w4685_ ;
	wire _w4684_ ;
	wire _w4683_ ;
	wire _w4682_ ;
	wire _w4681_ ;
	wire _w4680_ ;
	wire _w4679_ ;
	wire _w4678_ ;
	wire _w4677_ ;
	wire _w4676_ ;
	wire _w4675_ ;
	wire _w4674_ ;
	wire _w4673_ ;
	wire _w4672_ ;
	wire _w4671_ ;
	wire _w4670_ ;
	wire _w4669_ ;
	wire _w4668_ ;
	wire _w4667_ ;
	wire _w4666_ ;
	wire _w4665_ ;
	wire _w4664_ ;
	wire _w4663_ ;
	wire _w4662_ ;
	wire _w4661_ ;
	wire _w4660_ ;
	wire _w4659_ ;
	wire _w4658_ ;
	wire _w4657_ ;
	wire _w4656_ ;
	wire _w4655_ ;
	wire _w4654_ ;
	wire _w4653_ ;
	wire _w4652_ ;
	wire _w4651_ ;
	wire _w4650_ ;
	wire _w4649_ ;
	wire _w4648_ ;
	wire _w4647_ ;
	wire _w4646_ ;
	wire _w4645_ ;
	wire _w4644_ ;
	wire _w4643_ ;
	wire _w4642_ ;
	wire _w4641_ ;
	wire _w4640_ ;
	wire _w4639_ ;
	wire _w4638_ ;
	wire _w4637_ ;
	wire _w4636_ ;
	wire _w4635_ ;
	wire _w4634_ ;
	wire _w4633_ ;
	wire _w4632_ ;
	wire _w4631_ ;
	wire _w4630_ ;
	wire _w4629_ ;
	wire _w4628_ ;
	wire _w4627_ ;
	wire _w4626_ ;
	wire _w4625_ ;
	wire _w4624_ ;
	wire _w4623_ ;
	wire _w4622_ ;
	wire _w4621_ ;
	wire _w4620_ ;
	wire _w4619_ ;
	wire _w4618_ ;
	wire _w4617_ ;
	wire _w4616_ ;
	wire _w4615_ ;
	wire _w4614_ ;
	wire _w4613_ ;
	wire _w4612_ ;
	wire _w4611_ ;
	wire _w4610_ ;
	wire _w4609_ ;
	wire _w4608_ ;
	wire _w4607_ ;
	wire _w4606_ ;
	wire _w4605_ ;
	wire _w4604_ ;
	wire _w4603_ ;
	wire _w4602_ ;
	wire _w4601_ ;
	wire _w4600_ ;
	wire _w4599_ ;
	wire _w4598_ ;
	wire _w4597_ ;
	wire _w4596_ ;
	wire _w4595_ ;
	wire _w4594_ ;
	wire _w4593_ ;
	wire _w4592_ ;
	wire _w4591_ ;
	wire _w4590_ ;
	wire _w4589_ ;
	wire _w4588_ ;
	wire _w4587_ ;
	wire _w4586_ ;
	wire _w4585_ ;
	wire _w4584_ ;
	wire _w4583_ ;
	wire _w4582_ ;
	wire _w4581_ ;
	wire _w4580_ ;
	wire _w4579_ ;
	wire _w4578_ ;
	wire _w4577_ ;
	wire _w4576_ ;
	wire _w4575_ ;
	wire _w4574_ ;
	wire _w4573_ ;
	wire _w4572_ ;
	wire _w4571_ ;
	wire _w4570_ ;
	wire _w4569_ ;
	wire _w4568_ ;
	wire _w4567_ ;
	wire _w4566_ ;
	wire _w4565_ ;
	wire _w4564_ ;
	wire _w4563_ ;
	wire _w4562_ ;
	wire _w4561_ ;
	wire _w4560_ ;
	wire _w4559_ ;
	wire _w4558_ ;
	wire _w4557_ ;
	wire _w4556_ ;
	wire _w4555_ ;
	wire _w4554_ ;
	wire _w4553_ ;
	wire _w4552_ ;
	wire _w4551_ ;
	wire _w4550_ ;
	wire _w4549_ ;
	wire _w4548_ ;
	wire _w4547_ ;
	wire _w4546_ ;
	wire _w4545_ ;
	wire _w4544_ ;
	wire _w4543_ ;
	wire _w4542_ ;
	wire _w4541_ ;
	wire _w4540_ ;
	wire _w4539_ ;
	wire _w4538_ ;
	wire _w4537_ ;
	wire _w4536_ ;
	wire _w4535_ ;
	wire _w4534_ ;
	wire _w4533_ ;
	wire _w4532_ ;
	wire _w4531_ ;
	wire _w4530_ ;
	wire _w4529_ ;
	wire _w4528_ ;
	wire _w4527_ ;
	wire _w4526_ ;
	wire _w4525_ ;
	wire _w4524_ ;
	wire _w4523_ ;
	wire _w4522_ ;
	wire _w4521_ ;
	wire _w4520_ ;
	wire _w4519_ ;
	wire _w4518_ ;
	wire _w4517_ ;
	wire _w4516_ ;
	wire _w4515_ ;
	wire _w4514_ ;
	wire _w4513_ ;
	wire _w4512_ ;
	wire _w4511_ ;
	wire _w4510_ ;
	wire _w4509_ ;
	wire _w4508_ ;
	wire _w4507_ ;
	wire _w4506_ ;
	wire _w4505_ ;
	wire _w4504_ ;
	wire _w4503_ ;
	wire _w4502_ ;
	wire _w4501_ ;
	wire _w4500_ ;
	wire _w4499_ ;
	wire _w4498_ ;
	wire _w4497_ ;
	wire _w4496_ ;
	wire _w4495_ ;
	wire _w4494_ ;
	wire _w4493_ ;
	wire _w4492_ ;
	wire _w4491_ ;
	wire _w4490_ ;
	wire _w4489_ ;
	wire _w4488_ ;
	wire _w4487_ ;
	wire _w4486_ ;
	wire _w4485_ ;
	wire _w4484_ ;
	wire _w4483_ ;
	wire _w4482_ ;
	wire _w4481_ ;
	wire _w4480_ ;
	wire _w4479_ ;
	wire _w4478_ ;
	wire _w4477_ ;
	wire _w4476_ ;
	wire _w4475_ ;
	wire _w4474_ ;
	wire _w4473_ ;
	wire _w4472_ ;
	wire _w4471_ ;
	wire _w4470_ ;
	wire _w4469_ ;
	wire _w4468_ ;
	wire _w4467_ ;
	wire _w4466_ ;
	wire _w4465_ ;
	wire _w4464_ ;
	wire _w4463_ ;
	wire _w4462_ ;
	wire _w4461_ ;
	wire _w4460_ ;
	wire _w4459_ ;
	wire _w4458_ ;
	wire _w4457_ ;
	wire _w4456_ ;
	wire _w4455_ ;
	wire _w4454_ ;
	wire _w4453_ ;
	wire _w4452_ ;
	wire _w4451_ ;
	wire _w4450_ ;
	wire _w4449_ ;
	wire _w4448_ ;
	wire _w4447_ ;
	wire _w4446_ ;
	wire _w4445_ ;
	wire _w4444_ ;
	wire _w4443_ ;
	wire _w4442_ ;
	wire _w4441_ ;
	wire _w4440_ ;
	wire _w4439_ ;
	wire _w4438_ ;
	wire _w4437_ ;
	wire _w4436_ ;
	wire _w4435_ ;
	wire _w4434_ ;
	wire _w4433_ ;
	wire _w4432_ ;
	wire _w4431_ ;
	wire _w4430_ ;
	wire _w4429_ ;
	wire _w4428_ ;
	wire _w4427_ ;
	wire _w4426_ ;
	wire _w4425_ ;
	wire _w4424_ ;
	wire _w4423_ ;
	wire _w4422_ ;
	wire _w4421_ ;
	wire _w4420_ ;
	wire _w4419_ ;
	wire _w4418_ ;
	wire _w4417_ ;
	wire _w4416_ ;
	wire _w4415_ ;
	wire _w4414_ ;
	wire _w4413_ ;
	wire _w4412_ ;
	wire _w4411_ ;
	wire _w4410_ ;
	wire _w4409_ ;
	wire _w4408_ ;
	wire _w4407_ ;
	wire _w4406_ ;
	wire _w4405_ ;
	wire _w4404_ ;
	wire _w4403_ ;
	wire _w4402_ ;
	wire _w4401_ ;
	wire _w4400_ ;
	wire _w4399_ ;
	wire _w4398_ ;
	wire _w4397_ ;
	wire _w4396_ ;
	wire _w4395_ ;
	wire _w4394_ ;
	wire _w4393_ ;
	wire _w4392_ ;
	wire _w4391_ ;
	wire _w4390_ ;
	wire _w4389_ ;
	wire _w4388_ ;
	wire _w4387_ ;
	wire _w4386_ ;
	wire _w4385_ ;
	wire _w4384_ ;
	wire _w4383_ ;
	wire _w4382_ ;
	wire _w4381_ ;
	wire _w4380_ ;
	wire _w4379_ ;
	wire _w4378_ ;
	wire _w4377_ ;
	wire _w4376_ ;
	wire _w4375_ ;
	wire _w4374_ ;
	wire _w4373_ ;
	wire _w4372_ ;
	wire _w4371_ ;
	wire _w4370_ ;
	wire _w4369_ ;
	wire _w4368_ ;
	wire _w4367_ ;
	wire _w4366_ ;
	wire _w4365_ ;
	wire _w4364_ ;
	wire _w4363_ ;
	wire _w4362_ ;
	wire _w4361_ ;
	wire _w4360_ ;
	wire _w4359_ ;
	wire _w4358_ ;
	wire _w4357_ ;
	wire _w4356_ ;
	wire _w4355_ ;
	wire _w4354_ ;
	wire _w4353_ ;
	wire _w4352_ ;
	wire _w4351_ ;
	wire _w4350_ ;
	wire _w4349_ ;
	wire _w4348_ ;
	wire _w4347_ ;
	wire _w4346_ ;
	wire _w4345_ ;
	wire _w4344_ ;
	wire _w4343_ ;
	wire _w4342_ ;
	wire _w4341_ ;
	wire _w4340_ ;
	wire _w4339_ ;
	wire _w4338_ ;
	wire _w4337_ ;
	wire _w4336_ ;
	wire _w4335_ ;
	wire _w4334_ ;
	wire _w4333_ ;
	wire _w4332_ ;
	wire _w4331_ ;
	wire _w4330_ ;
	wire _w4329_ ;
	wire _w4328_ ;
	wire _w4327_ ;
	wire _w4326_ ;
	wire _w4325_ ;
	wire _w4324_ ;
	wire _w4323_ ;
	wire _w4322_ ;
	wire _w4321_ ;
	wire _w4320_ ;
	wire _w4319_ ;
	wire _w4318_ ;
	wire _w4317_ ;
	wire _w4316_ ;
	wire _w4315_ ;
	wire _w4314_ ;
	wire _w4313_ ;
	wire _w4312_ ;
	wire _w4311_ ;
	wire _w4310_ ;
	wire _w4309_ ;
	wire _w4308_ ;
	wire _w4307_ ;
	wire _w4306_ ;
	wire _w4305_ ;
	wire _w4304_ ;
	wire _w4303_ ;
	wire _w4302_ ;
	wire _w4301_ ;
	wire _w4300_ ;
	wire _w4299_ ;
	wire _w4298_ ;
	wire _w4297_ ;
	wire _w4296_ ;
	wire _w4295_ ;
	wire _w4294_ ;
	wire _w4293_ ;
	wire _w4292_ ;
	wire _w4291_ ;
	wire _w4290_ ;
	wire _w4289_ ;
	wire _w4288_ ;
	wire _w4287_ ;
	wire _w4286_ ;
	wire _w4285_ ;
	wire _w4284_ ;
	wire _w4283_ ;
	wire _w4282_ ;
	wire _w4281_ ;
	wire _w4280_ ;
	wire _w4279_ ;
	wire _w4278_ ;
	wire _w4277_ ;
	wire _w4276_ ;
	wire _w4275_ ;
	wire _w4274_ ;
	wire _w4273_ ;
	wire _w4272_ ;
	wire _w4271_ ;
	wire _w4270_ ;
	wire _w4269_ ;
	wire _w4268_ ;
	wire _w4267_ ;
	wire _w4266_ ;
	wire _w4265_ ;
	wire _w4264_ ;
	wire _w4263_ ;
	wire _w4262_ ;
	wire _w4261_ ;
	wire _w4260_ ;
	wire _w4259_ ;
	wire _w4258_ ;
	wire _w4257_ ;
	wire _w4256_ ;
	wire _w4255_ ;
	wire _w4254_ ;
	wire _w4253_ ;
	wire _w4252_ ;
	wire _w4251_ ;
	wire _w4250_ ;
	wire _w4249_ ;
	wire _w4248_ ;
	wire _w4247_ ;
	wire _w4246_ ;
	wire _w4245_ ;
	wire _w4244_ ;
	wire _w4243_ ;
	wire _w4242_ ;
	wire _w4241_ ;
	wire _w4240_ ;
	wire _w4239_ ;
	wire _w4238_ ;
	wire _w4237_ ;
	wire _w4236_ ;
	wire _w4235_ ;
	wire _w4234_ ;
	wire _w4233_ ;
	wire _w4232_ ;
	wire _w4231_ ;
	wire _w4230_ ;
	wire _w4229_ ;
	wire _w4228_ ;
	wire _w4227_ ;
	wire _w4226_ ;
	wire _w4225_ ;
	wire _w4224_ ;
	wire _w4223_ ;
	wire _w4222_ ;
	wire _w4221_ ;
	wire _w4220_ ;
	wire _w4219_ ;
	wire _w4218_ ;
	wire _w4217_ ;
	wire _w4216_ ;
	wire _w4215_ ;
	wire _w4214_ ;
	wire _w4213_ ;
	wire _w4212_ ;
	wire _w4211_ ;
	wire _w4210_ ;
	wire _w4209_ ;
	wire _w4208_ ;
	wire _w4207_ ;
	wire _w4206_ ;
	wire _w4205_ ;
	wire _w4204_ ;
	wire _w4203_ ;
	wire _w4202_ ;
	wire _w4201_ ;
	wire _w4200_ ;
	wire _w4199_ ;
	wire _w4198_ ;
	wire _w4197_ ;
	wire _w4196_ ;
	wire _w4195_ ;
	wire _w4194_ ;
	wire _w4193_ ;
	wire _w4192_ ;
	wire _w4191_ ;
	wire _w4190_ ;
	wire _w4189_ ;
	wire _w4188_ ;
	wire _w4187_ ;
	wire _w4186_ ;
	wire _w4185_ ;
	wire _w4184_ ;
	wire _w4183_ ;
	wire _w4182_ ;
	wire _w4181_ ;
	wire _w4180_ ;
	wire _w4179_ ;
	wire _w4178_ ;
	wire _w4177_ ;
	wire _w4176_ ;
	wire _w4175_ ;
	wire _w4174_ ;
	wire _w4173_ ;
	wire _w4172_ ;
	wire _w4171_ ;
	wire _w4170_ ;
	wire _w4169_ ;
	wire _w4168_ ;
	wire _w4167_ ;
	wire _w4166_ ;
	wire _w4165_ ;
	wire _w4164_ ;
	wire _w4163_ ;
	wire _w4162_ ;
	wire _w4161_ ;
	wire _w4160_ ;
	wire _w4159_ ;
	wire _w4158_ ;
	wire _w4157_ ;
	wire _w4156_ ;
	wire _w4155_ ;
	wire _w4154_ ;
	wire _w4153_ ;
	wire _w4152_ ;
	wire _w4151_ ;
	wire _w4150_ ;
	wire _w4149_ ;
	wire _w4148_ ;
	wire _w4147_ ;
	wire _w4146_ ;
	wire _w4145_ ;
	wire _w4144_ ;
	wire _w4143_ ;
	wire _w4142_ ;
	wire _w4141_ ;
	wire _w4140_ ;
	wire _w4139_ ;
	wire _w4138_ ;
	wire _w4137_ ;
	wire _w4136_ ;
	wire _w4135_ ;
	wire _w4134_ ;
	wire _w4133_ ;
	wire _w4132_ ;
	wire _w4131_ ;
	wire _w4130_ ;
	wire _w4129_ ;
	wire _w4128_ ;
	wire _w4127_ ;
	wire _w4126_ ;
	wire _w4125_ ;
	wire _w4124_ ;
	wire _w4123_ ;
	wire _w4122_ ;
	wire _w4121_ ;
	wire _w4120_ ;
	wire _w4119_ ;
	wire _w4118_ ;
	wire _w4117_ ;
	wire _w4116_ ;
	wire _w4115_ ;
	wire _w4114_ ;
	wire _w4113_ ;
	wire _w4112_ ;
	wire _w4111_ ;
	wire _w4110_ ;
	wire _w4109_ ;
	wire _w4108_ ;
	wire _w4107_ ;
	wire _w4106_ ;
	wire _w4105_ ;
	wire _w4104_ ;
	wire _w4103_ ;
	wire _w4102_ ;
	wire _w4101_ ;
	wire _w4100_ ;
	wire _w4099_ ;
	wire _w4098_ ;
	wire _w4097_ ;
	wire _w4096_ ;
	wire _w4095_ ;
	wire _w4094_ ;
	wire _w4093_ ;
	wire _w4092_ ;
	wire _w4091_ ;
	wire _w4090_ ;
	wire _w4089_ ;
	wire _w4088_ ;
	wire _w4087_ ;
	wire _w4086_ ;
	wire _w4085_ ;
	wire _w4084_ ;
	wire _w4083_ ;
	wire _w4082_ ;
	wire _w4081_ ;
	wire _w4080_ ;
	wire _w4079_ ;
	wire _w4078_ ;
	wire _w4077_ ;
	wire _w4076_ ;
	wire _w4075_ ;
	wire _w4074_ ;
	wire _w4073_ ;
	wire _w4072_ ;
	wire _w4071_ ;
	wire _w4070_ ;
	wire _w4069_ ;
	wire _w4068_ ;
	wire _w4067_ ;
	wire _w4066_ ;
	wire _w4065_ ;
	wire _w4064_ ;
	wire _w4063_ ;
	wire _w4062_ ;
	wire _w4061_ ;
	wire _w4060_ ;
	wire _w4059_ ;
	wire _w4058_ ;
	wire _w4057_ ;
	wire _w4056_ ;
	wire _w4055_ ;
	wire _w4054_ ;
	wire _w4053_ ;
	wire _w4052_ ;
	wire _w4051_ ;
	wire _w4050_ ;
	wire _w4049_ ;
	wire _w4048_ ;
	wire _w4047_ ;
	wire _w4046_ ;
	wire _w4045_ ;
	wire _w4044_ ;
	wire _w4043_ ;
	wire _w4042_ ;
	wire _w4041_ ;
	wire _w4040_ ;
	wire _w4039_ ;
	wire _w4038_ ;
	wire _w4037_ ;
	wire _w4036_ ;
	wire _w4035_ ;
	wire _w4034_ ;
	wire _w4033_ ;
	wire _w4032_ ;
	wire _w4031_ ;
	wire _w4030_ ;
	wire _w4029_ ;
	wire _w4028_ ;
	wire _w4027_ ;
	wire _w4026_ ;
	wire _w4025_ ;
	wire _w4024_ ;
	wire _w4023_ ;
	wire _w4022_ ;
	wire _w4021_ ;
	wire _w4020_ ;
	wire _w4019_ ;
	wire _w4018_ ;
	wire _w4017_ ;
	wire _w4016_ ;
	wire _w4015_ ;
	wire _w4014_ ;
	wire _w4013_ ;
	wire _w4012_ ;
	wire _w4011_ ;
	wire _w4010_ ;
	wire _w4009_ ;
	wire _w4008_ ;
	wire _w4007_ ;
	wire _w4006_ ;
	wire _w4005_ ;
	wire _w4004_ ;
	wire _w4003_ ;
	wire _w4002_ ;
	wire _w4001_ ;
	wire _w4000_ ;
	wire _w3999_ ;
	wire _w3998_ ;
	wire _w3997_ ;
	wire _w3996_ ;
	wire _w3995_ ;
	wire _w3994_ ;
	wire _w3993_ ;
	wire _w3992_ ;
	wire _w3991_ ;
	wire _w3990_ ;
	wire _w3989_ ;
	wire _w3988_ ;
	wire _w3987_ ;
	wire _w3986_ ;
	wire _w3985_ ;
	wire _w3984_ ;
	wire _w3983_ ;
	wire _w3982_ ;
	wire _w3981_ ;
	wire _w3980_ ;
	wire _w3979_ ;
	wire _w3978_ ;
	wire _w3977_ ;
	wire _w3976_ ;
	wire _w3975_ ;
	wire _w3974_ ;
	wire _w3973_ ;
	wire _w3972_ ;
	wire _w3971_ ;
	wire _w3970_ ;
	wire _w3969_ ;
	wire _w3968_ ;
	wire _w3967_ ;
	wire _w3966_ ;
	wire _w3965_ ;
	wire _w3964_ ;
	wire _w3963_ ;
	wire _w3962_ ;
	wire _w3961_ ;
	wire _w3960_ ;
	wire _w3959_ ;
	wire _w3958_ ;
	wire _w3957_ ;
	wire _w3956_ ;
	wire _w3955_ ;
	wire _w3954_ ;
	wire _w3953_ ;
	wire _w3952_ ;
	wire _w3951_ ;
	wire _w3950_ ;
	wire _w3949_ ;
	wire _w3948_ ;
	wire _w3947_ ;
	wire _w3946_ ;
	wire _w3945_ ;
	wire _w3944_ ;
	wire _w3943_ ;
	wire _w3942_ ;
	wire _w3941_ ;
	wire _w3940_ ;
	wire _w3939_ ;
	wire _w3938_ ;
	wire _w3937_ ;
	wire _w3936_ ;
	wire _w3935_ ;
	wire _w3934_ ;
	wire _w3933_ ;
	wire _w3932_ ;
	wire _w3931_ ;
	wire _w3930_ ;
	wire _w3929_ ;
	wire _w3928_ ;
	wire _w3927_ ;
	wire _w3926_ ;
	wire _w3925_ ;
	wire _w3924_ ;
	wire _w3923_ ;
	wire _w3922_ ;
	wire _w3921_ ;
	wire _w3920_ ;
	wire _w3919_ ;
	wire _w3918_ ;
	wire _w3917_ ;
	wire _w3916_ ;
	wire _w3915_ ;
	wire _w3914_ ;
	wire _w3913_ ;
	wire _w3912_ ;
	wire _w3911_ ;
	wire _w3910_ ;
	wire _w3909_ ;
	wire _w3908_ ;
	wire _w3907_ ;
	wire _w3906_ ;
	wire _w3905_ ;
	wire _w3904_ ;
	wire _w3903_ ;
	wire _w3902_ ;
	wire _w3901_ ;
	wire _w3900_ ;
	wire _w3899_ ;
	wire _w3898_ ;
	wire _w3897_ ;
	wire _w3896_ ;
	wire _w3895_ ;
	wire _w3894_ ;
	wire _w3893_ ;
	wire _w3892_ ;
	wire _w3891_ ;
	wire _w3890_ ;
	wire _w3889_ ;
	wire _w3888_ ;
	wire _w3887_ ;
	wire _w3886_ ;
	wire _w3885_ ;
	wire _w3884_ ;
	wire _w3883_ ;
	wire _w3882_ ;
	wire _w3881_ ;
	wire _w3880_ ;
	wire _w3879_ ;
	wire _w3878_ ;
	wire _w3877_ ;
	wire _w3876_ ;
	wire _w3875_ ;
	wire _w3874_ ;
	wire _w3873_ ;
	wire _w3872_ ;
	wire _w3871_ ;
	wire _w3870_ ;
	wire _w3869_ ;
	wire _w3868_ ;
	wire _w3867_ ;
	wire _w3866_ ;
	wire _w3865_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w2288_ ;
	wire _w2286_ ;
	wire _w2285_ ;
	wire _w2284_ ;
	wire _w2283_ ;
	wire _w2282_ ;
	wire _w2281_ ;
	wire _w2280_ ;
	wire _w2279_ ;
	wire _w2278_ ;
	wire _w2277_ ;
	wire _w2276_ ;
	wire _w2275_ ;
	wire _w2274_ ;
	wire _w2273_ ;
	wire _w2272_ ;
	wire _w2271_ ;
	wire _w2270_ ;
	wire _w2268_ ;
	wire _w2267_ ;
	wire _w2266_ ;
	wire _w2265_ ;
	wire _w2264_ ;
	wire _w2263_ ;
	wire _w2262_ ;
	wire _w2261_ ;
	wire _w2260_ ;
	wire _w2259_ ;
	wire _w2258_ ;
	wire _w2257_ ;
	wire _w2256_ ;
	wire _w2255_ ;
	wire _w2254_ ;
	wire _w2253_ ;
	wire _w2252_ ;
	wire _w2251_ ;
	wire _w2247_ ;
	wire _w2245_ ;
	wire _w2243_ ;
	wire _w2241_ ;
	wire _w2240_ ;
	wire _w2238_ ;
	wire _w2236_ ;
	wire _w2233_ ;
	wire _w2232_ ;
	wire _w2231_ ;
	wire _w2230_ ;
	wire _w2229_ ;
	wire _w2228_ ;
	wire _w2227_ ;
	wire _w2226_ ;
	wire _w2225_ ;
	wire _w2224_ ;
	wire _w2223_ ;
	wire _w2222_ ;
	wire _w2221_ ;
	wire _w2220_ ;
	wire _w2219_ ;
	wire _w2218_ ;
	wire _w2217_ ;
	wire _w2216_ ;
	wire _w2215_ ;
	wire _w2214_ ;
	wire _w2213_ ;
	wire _w2212_ ;
	wire _w2211_ ;
	wire _w2210_ ;
	wire _w2209_ ;
	wire _w2208_ ;
	wire _w2207_ ;
	wire _w2206_ ;
	wire _w2205_ ;
	wire _w2204_ ;
	wire _w2203_ ;
	wire _w2202_ ;
	wire _w2201_ ;
	wire _w2200_ ;
	wire _w2199_ ;
	wire _w2198_ ;
	wire _w2197_ ;
	wire _w2196_ ;
	wire _w2195_ ;
	wire _w2194_ ;
	wire _w2193_ ;
	wire _w2192_ ;
	wire _w2191_ ;
	wire _w2190_ ;
	wire _w2189_ ;
	wire _w2188_ ;
	wire _w2187_ ;
	wire _w2186_ ;
	wire _w2185_ ;
	wire _w2184_ ;
	wire _w2183_ ;
	wire _w2182_ ;
	wire _w2181_ ;
	wire _w2180_ ;
	wire _w2179_ ;
	wire _w2178_ ;
	wire _w2177_ ;
	wire _w2176_ ;
	wire _w2175_ ;
	wire _w2174_ ;
	wire _w2173_ ;
	wire _w2172_ ;
	wire _w2171_ ;
	wire _w2170_ ;
	wire _w2169_ ;
	wire _w2168_ ;
	wire _w2167_ ;
	wire _w2166_ ;
	wire _w2165_ ;
	wire _w2164_ ;
	wire _w2163_ ;
	wire _w2162_ ;
	wire _w2161_ ;
	wire _w2160_ ;
	wire _w2159_ ;
	wire _w2158_ ;
	wire _w2157_ ;
	wire _w2156_ ;
	wire _w2155_ ;
	wire _w2154_ ;
	wire _w2153_ ;
	wire _w2152_ ;
	wire _w2151_ ;
	wire _w2150_ ;
	wire _w2149_ ;
	wire _w2148_ ;
	wire _w2147_ ;
	wire _w2146_ ;
	wire _w2145_ ;
	wire _w2144_ ;
	wire _w2143_ ;
	wire _w2142_ ;
	wire _w2141_ ;
	wire _w2140_ ;
	wire _w2139_ ;
	wire _w2138_ ;
	wire _w2137_ ;
	wire _w2136_ ;
	wire _w2135_ ;
	wire _w2134_ ;
	wire _w2133_ ;
	wire _w2132_ ;
	wire _w2131_ ;
	wire _w2130_ ;
	wire _w2129_ ;
	wire _w2128_ ;
	wire _w2127_ ;
	wire _w2126_ ;
	wire _w2125_ ;
	wire _w2124_ ;
	wire _w2122_ ;
	wire _w2120_ ;
	wire _w2119_ ;
	wire _w2118_ ;
	wire _w2117_ ;
	wire _w2116_ ;
	wire _w2115_ ;
	wire _w2114_ ;
	wire _w2113_ ;
	wire _w2112_ ;
	wire _w2111_ ;
	wire _w2110_ ;
	wire _w2109_ ;
	wire _w2108_ ;
	wire _w2107_ ;
	wire _w2106_ ;
	wire _w2105_ ;
	wire _w2104_ ;
	wire _w2103_ ;
	wire _w2102_ ;
	wire _w2101_ ;
	wire _w2100_ ;
	wire _w2099_ ;
	wire _w2098_ ;
	wire _w2097_ ;
	wire _w2096_ ;
	wire _w2095_ ;
	wire _w2094_ ;
	wire _w2093_ ;
	wire _w2092_ ;
	wire _w2091_ ;
	wire _w2090_ ;
	wire _w2089_ ;
	wire _w2088_ ;
	wire _w2087_ ;
	wire _w2086_ ;
	wire _w2085_ ;
	wire _w2084_ ;
	wire _w2083_ ;
	wire _w2082_ ;
	wire _w2081_ ;
	wire _w2080_ ;
	wire _w2079_ ;
	wire _w2078_ ;
	wire _w2077_ ;
	wire _w2076_ ;
	wire _w2075_ ;
	wire _w2074_ ;
	wire _w2073_ ;
	wire _w2072_ ;
	wire _w2071_ ;
	wire _w2070_ ;
	wire _w2069_ ;
	wire _w2068_ ;
	wire _w2067_ ;
	wire _w2066_ ;
	wire _w2065_ ;
	wire _w2064_ ;
	wire _w2063_ ;
	wire _w2062_ ;
	wire _w2061_ ;
	wire _w2060_ ;
	wire _w2059_ ;
	wire _w2058_ ;
	wire _w2057_ ;
	wire _w2056_ ;
	wire _w2055_ ;
	wire _w2054_ ;
	wire _w2053_ ;
	wire _w2052_ ;
	wire _w2051_ ;
	wire _w2050_ ;
	wire _w2049_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1955_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1950_ ;
	wire _w1948_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1825_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1764_ ;
	wire _w1763_ ;
	wire _w1762_ ;
	wire _w1761_ ;
	wire _w1760_ ;
	wire _w1759_ ;
	wire _w1758_ ;
	wire _w1756_ ;
	wire _w1754_ ;
	wire _w1752_ ;
	wire _w1750_ ;
	wire _w1748_ ;
	wire _w1746_ ;
	wire _w1744_ ;
	wire _w1743_ ;
	wire _w1742_ ;
	wire _w1741_ ;
	wire _w1740_ ;
	wire _w1739_ ;
	wire _w1738_ ;
	wire _w1737_ ;
	wire _w1736_ ;
	wire _w1735_ ;
	wire _w1734_ ;
	wire _w1733_ ;
	wire _w1732_ ;
	wire _w1731_ ;
	wire _w1730_ ;
	wire _w1729_ ;
	wire _w1728_ ;
	wire _w1727_ ;
	wire _w1726_ ;
	wire _w1725_ ;
	wire _w1724_ ;
	wire _w1723_ ;
	wire _w1722_ ;
	wire _w1437_ ;
	wire _w1436_ ;
	wire _w1435_ ;
	wire _w1434_ ;
	wire _w1433_ ;
	wire _w1432_ ;
	wire _w1431_ ;
	wire _w1430_ ;
	wire _w1429_ ;
	wire _w1428_ ;
	wire _w1427_ ;
	wire _w1426_ ;
	wire _w1425_ ;
	wire _w1424_ ;
	wire _w1423_ ;
	wire _w1422_ ;
	wire _w1421_ ;
	wire _w1420_ ;
	wire _w1418_ ;
	wire _w1416_ ;
	wire _w1414_ ;
	wire _w1412_ ;
	wire _w1410_ ;
	wire _w1408_ ;
	wire _w1406_ ;
	wire _w1404_ ;
	wire _w1403_ ;
	wire _w1402_ ;
	wire _w1401_ ;
	wire _w1969_ ;
	wire _w860_ ;
	wire _w3217_ ;
	wire _w1400_ ;
	wire _w1399_ ;
	wire _w1397_ ;
	wire _w1395_ ;
	wire _w1393_ ;
	wire _w1391_ ;
	wire _w1389_ ;
	wire _w1388_ ;
	wire _w1956_ ;
	wire _w847_ ;
	wire _w3204_ ;
	wire _w1384_ ;
	wire _w1382_ ;
	wire _w1381_ ;
	wire _w1949_ ;
	wire _w840_ ;
	wire _w3197_ ;
	wire _w1380_ ;
	wire _w1379_ ;
	wire _w1947_ ;
	wire _w838_ ;
	wire _w3195_ ;
	wire _w1378_ ;
	wire _w1377_ ;
	wire _w1376_ ;
	wire _w1375_ ;
	wire _w1372_ ;
	wire _w1370_ ;
	wire _w1368_ ;
	wire _w1366_ ;
	wire _w1364_ ;
	wire _w1362_ ;
	wire _w1360_ ;
	wire _w1357_ ;
	wire _w1355_ ;
	wire _w1353_ ;
	wire _w1351_ ;
	wire _w1350_ ;
	wire _w1349_ ;
	wire _w1347_ ;
	wire _w1345_ ;
	wire _w1344_ ;
	wire _w1342_ ;
	wire _w1340_ ;
	wire _w1339_ ;
	wire _w1337_ ;
	wire _w1335_ ;
	wire _w1332_ ;
	wire _w1330_ ;
	wire _w1329_ ;
	wire _w1327_ ;
	wire _w1326_ ;
	wire _w1324_ ;
	wire _w1322_ ;
	wire _w1320_ ;
	wire _w1318_ ;
	wire _w1314_ ;
	wire _w1341_ ;
	wire _w232_ ;
	wire _w2589_ ;
	wire _w1313_ ;
	wire _w1311_ ;
	wire _w1338_ ;
	wire _w229_ ;
	wire _w2586_ ;
	wire _w1310_ ;
	wire _w1309_ ;
	wire _w1308_ ;
	wire _w1383_ ;
	wire _w1951_ ;
	wire _w842_ ;
	wire _w3199_ ;
	wire _w2235_ ;
	wire _w1126_ ;
	wire _w3483_ ;
	wire _w1667_ ;
	wire _w1253_ ;
	wire _w1398_ ;
	wire _w2250_ ;
	wire _w1141_ ;
	wire _w3498_ ;
	wire _w1682_ ;
	wire _w1268_ ;
	wire _w1374_ ;
	wire _w1241_ ;
	wire _w1334_ ;
	wire _w1929_ ;
	wire _w820_ ;
	wire _w3177_ ;
	wire _w1361_ ;
	wire _w1387_ ;
	wire _w2239_ ;
	wire _w1130_ ;
	wire _w3487_ ;
	wire _w1671_ ;
	wire _w1396_ ;
	wire _w2248_ ;
	wire _w1139_ ;
	wire _w3496_ ;
	wire _w1680_ ;
	wire _w1266_ ;
	wire _w1385_ ;
	wire _w2237_ ;
	wire _w1128_ ;
	wire _w3485_ ;
	wire _w1669_ ;
	wire _w1824_ ;
	wire _w715_ ;
	wire _w3072_ ;
	wire _w1256_ ;
	wire _w1419_ ;
	wire _w1757_ ;
	wire _w648_ ;
	wire _w3005_ ;
	wire _w1283_ ;
	wire _w1417_ ;
	wire _w1755_ ;
	wire _w646_ ;
	wire _w3003_ ;
	wire _w1281_ ;
	wire _w1415_ ;
	wire _w1753_ ;
	wire _w644_ ;
	wire _w3001_ ;
	wire _w1279_ ;
	wire _w1328_ ;
	wire _w2234_ ;
	wire _w5103_ ;
	wire _w16_ ;
	wire _w2373_ ;
	wire _w1639_ ;
	wire _w1325_ ;
	wire _w1636_ ;
	wire _w1323_ ;
	wire _w1634_ ;
	wire _w1359_ ;
	wire _w1954_ ;
	wire _w845_ ;
	wire _w3202_ ;
	wire _w1386_ ;
	wire _w1365_ ;
	wire _w1321_ ;
	wire _w1348_ ;
	wire _w239_ ;
	wire _w2596_ ;
	wire _w1632_ ;
	wire _w1319_ ;
	wire _w1346_ ;
	wire _w237_ ;
	wire _w2594_ ;
	wire _w1630_ ;
	wire _w1503_ ;
	wire _w1413_ ;
	wire _w1751_ ;
	wire _w642_ ;
	wire _w2999_ ;
	wire _w101_ ;
	wire _w2458_ ;
	wire _w1277_ ;
	wire _w1257_ ;
	wire _w1245_ ;
	wire _w1367_ ;
	wire _w1962_ ;
	wire _w853_ ;
	wire _w3210_ ;
	wire _w1394_ ;
	wire _w1373_ ;
	wire _w1392_ ;
	wire _w2244_ ;
	wire _w1135_ ;
	wire _w3492_ ;
	wire _w1676_ ;
	wire _w1358_ ;
	wire _w73_ ;
	wire _w2430_ ;
	wire _w1696_ ;
	wire _w1411_ ;
	wire _w1749_ ;
	wire _w640_ ;
	wire _w2997_ ;
	wire _w1275_ ;
	wire _w1255_ ;
	wire _w1243_ ;
	wire _w1409_ ;
	wire _w1747_ ;
	wire _w638_ ;
	wire _w2995_ ;
	wire _w1720_ ;
	wire _w1273_ ;
	wire _w1371_ ;
	wire _w86_ ;
	wire _w2443_ ;
	wire _w1709_ ;
	wire _w1317_ ;
	wire _w1628_ ;
	wire _w1501_ ;
	wire _w1390_ ;
	wire _w2242_ ;
	wire _w1133_ ;
	wire _w3490_ ;
	wire _w2269_ ;
	wire _w51_ ;
	wire _w2408_ ;
	wire _w1674_ ;
	wire _w1352_ ;
	wire _w1356_ ;
	wire _w2289_ ;
	wire _w71_ ;
	wire _w2428_ ;
	wire _w1694_ ;
	wire _w1312_ ;
	wire _w1623_ ;
	wire _w1303_ ;
	wire _w1354_ ;
	wire _w2287_ ;
	wire _w69_ ;
	wire _w2426_ ;
	wire _w1692_ ;
	wire _w227_ ;
	wire _w2584_ ;
	wire _w1336_ ;
	wire _w1407_ ;
	wire _w1745_ ;
	wire _w636_ ;
	wire _w2993_ ;
	wire _w1718_ ;
	wire _w2123_ ;
	wire _w1014_ ;
	wire _w3371_ ;
	wire _w1555_ ;
	wire _w1271_ ;
	wire _w1369_ ;
	wire _w1315_ ;
	wire _w1626_ ;
	wire _w1306_ ;
	wire _w1333_ ;
	wire _w224_ ;
	wire _w2581_ ;
	wire _w1316_ ;
	wire _w1343_ ;
	wire _w234_ ;
	wire _w2591_ ;
	wire _w2249_ ;
	wire _w5118_ ;
	wire _w31_ ;
	wire _w2388_ ;
	wire _w1654_ ;
	wire _w1262_ ;
	wire _w1331_ ;
	wire _w222_ ;
	wire _w2579_ ;
	wire _w1304_ ;
	wire _w1250_ ;
	wire _w1405_ ;
	wire _w120_ ;
	wire _w2477_ ;
	wire _w1263_ ;
	wire _w2246_ ;
	wire _w1137_ ;
	wire _w3494_ ;
	wire _w1678_ ;
	wire _w1264_ ;
	wire _w1301_ ;
	wire _w1286_ ;
	wire _w1363_ ;
	wire _w1260_ ;
	wire _w1826_ ;
	wire _w717_ ;
	wire _w3074_ ;
	wire _w1258_ ;
	wire _w1231_ ;
	wire _w1233_ ;
	wire _w1235_ ;
	wire _w1237_ ;
	wire _w1239_ ;
	wire _w1251_ ;
	wire _w1252_ ;
	wire _w1254_ ;
	wire _w1259_ ;
	wire _w1261_ ;
	wire _w1265_ ;
	wire _w1267_ ;
	wire _w2121_ ;
	wire _w1012_ ;
	wire _w3369_ ;
	wire _w1553_ ;
	wire _w1269_ ;
	wire _w1270_ ;
	wire _w1272_ ;
	wire _w1274_ ;
	wire _w1276_ ;
	wire _w1278_ ;
	wire _w1280_ ;
	wire _w1282_ ;
	wire _w1284_ ;
	wire _w1285_ ;
	wire _w1287_ ;
	wire _w1288_ ;
	wire _w1289_ ;
	wire _w1290_ ;
	wire _w1291_ ;
	wire _w1292_ ;
	wire _w1293_ ;
	wire _w1294_ ;
	wire _w1295_ ;
	wire _w1296_ ;
	wire _w1297_ ;
	wire _w1298_ ;
	wire _w1299_ ;
	wire _w1300_ ;
	wire _w1302_ ;
	wire _w1305_ ;
	wire _w1307_ ;
	wire _w1438_ ;
	wire _w1439_ ;
	wire _w1440_ ;
	wire _w1441_ ;
	wire _w333_ ;
	wire _w2690_ ;
	wire _w1442_ ;
	wire _w1443_ ;
	wire _w335_ ;
	wire _w2692_ ;
	wire _w1444_ ;
	wire _w1445_ ;
	wire _w337_ ;
	wire _w2694_ ;
	wire _w1446_ ;
	wire _w1447_ ;
	wire _w339_ ;
	wire _w2696_ ;
	wire _w1448_ ;
	wire _w1449_ ;
	wire _w341_ ;
	wire _w2698_ ;
	wire _w1450_ ;
	wire _w1451_ ;
	wire _w343_ ;
	wire _w2700_ ;
	wire _w1452_ ;
	wire _w1453_ ;
	wire _w345_ ;
	wire _w2702_ ;
	wire _w1454_ ;
	wire _w1455_ ;
	wire _w1456_ ;
	wire _w1457_ ;
	wire _w1458_ ;
	wire _w1459_ ;
	wire _w1460_ ;
	wire _w1461_ ;
	wire _w1462_ ;
	wire _w1463_ ;
	wire _w1464_ ;
	wire _w1465_ ;
	wire _w1466_ ;
	wire _w1467_ ;
	wire _w1468_ ;
	wire _w1469_ ;
	wire _w1470_ ;
	wire _w1471_ ;
	wire _w1472_ ;
	wire _w1473_ ;
	wire _w1474_ ;
	wire _w1475_ ;
	wire _w1476_ ;
	wire _w1477_ ;
	wire _w1478_ ;
	wire _w1479_ ;
	wire _w1480_ ;
	wire _w1481_ ;
	wire _w1482_ ;
	wire _w1483_ ;
	wire _w1484_ ;
	wire _w1485_ ;
	wire _w1486_ ;
	wire _w1487_ ;
	wire _w1488_ ;
	wire _w1489_ ;
	wire _w1490_ ;
	wire _w1491_ ;
	wire _w1492_ ;
	wire _w1493_ ;
	wire _w1494_ ;
	wire _w1495_ ;
	wire _w1496_ ;
	wire _w1497_ ;
	wire _w1498_ ;
	wire _w1499_ ;
	wire _w1500_ ;
	wire _w1502_ ;
	wire _w1504_ ;
	wire _w1505_ ;
	wire _w1506_ ;
	wire _w1507_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1521_ ;
	wire _w1522_ ;
	wire _w1523_ ;
	wire _w1524_ ;
	wire _w1525_ ;
	wire _w1526_ ;
	wire _w1527_ ;
	wire _w419_ ;
	wire _w2776_ ;
	wire _w1528_ ;
	wire _w1529_ ;
	wire _w421_ ;
	wire _w2778_ ;
	wire _w1530_ ;
	wire _w1531_ ;
	wire _w1532_ ;
	wire _w1533_ ;
	wire _w1534_ ;
	wire _w1535_ ;
	wire _w1536_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1554_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1567_ ;
	wire _w1568_ ;
	wire _w1569_ ;
	wire _w1570_ ;
	wire _w1571_ ;
	wire _w1572_ ;
	wire _w1573_ ;
	wire _w1574_ ;
	wire _w1575_ ;
	wire _w1576_ ;
	wire _w1577_ ;
	wire _w1578_ ;
	wire _w1579_ ;
	wire _w1580_ ;
	wire _w1581_ ;
	wire _w1582_ ;
	wire _w1583_ ;
	wire _w1584_ ;
	wire _w1585_ ;
	wire _w1586_ ;
	wire _w1587_ ;
	wire _w1588_ ;
	wire _w1589_ ;
	wire _w1590_ ;
	wire _w1591_ ;
	wire _w1592_ ;
	wire _w1593_ ;
	wire _w1594_ ;
	wire _w1595_ ;
	wire _w1596_ ;
	wire _w1597_ ;
	wire _w1598_ ;
	wire _w1599_ ;
	wire _w1600_ ;
	wire _w1601_ ;
	wire _w1602_ ;
	wire _w1603_ ;
	wire _w1604_ ;
	wire _w1605_ ;
	wire _w1606_ ;
	wire _w1607_ ;
	wire _w1608_ ;
	wire _w1609_ ;
	wire _w1610_ ;
	wire _w1611_ ;
	wire _w1612_ ;
	wire _w1613_ ;
	wire _w1614_ ;
	wire _w1615_ ;
	wire _w1616_ ;
	wire _w1617_ ;
	wire _w1618_ ;
	wire _w1619_ ;
	wire _w1620_ ;
	wire _w1621_ ;
	wire _w1622_ ;
	wire _w1624_ ;
	wire _w1625_ ;
	wire _w1627_ ;
	wire _w1629_ ;
	wire _w1631_ ;
	wire _w1633_ ;
	wire _w1635_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w541_ ;
	wire _w2898_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w544_ ;
	wire _w2901_ ;
	wire _w1653_ ;
	wire _w546_ ;
	wire _w2903_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w548_ ;
	wire _w2905_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w550_ ;
	wire _w2907_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w552_ ;
	wire _w2909_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w554_ ;
	wire _w2911_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w557_ ;
	wire _w2914_ ;
	wire _w1666_ ;
	wire _w1668_ ;
	wire _w1670_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1675_ ;
	wire _w1677_ ;
	wire _w1679_ ;
	wire _w1681_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1693_ ;
	wire _w1695_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1719_ ;
	wire _w1721_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2427_ ;
	wire _w2429_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2580_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2585_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2590_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2595_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w2617_ ;
	wire _w2618_ ;
	wire _w2619_ ;
	wire _w2620_ ;
	wire _w2621_ ;
	wire _w2622_ ;
	wire _w2623_ ;
	wire _w2624_ ;
	wire _w2625_ ;
	wire _w2626_ ;
	wire _w2627_ ;
	wire _w2628_ ;
	wire _w2629_ ;
	wire _w2630_ ;
	wire _w2631_ ;
	wire _w2632_ ;
	wire _w2633_ ;
	wire _w2634_ ;
	wire _w2635_ ;
	wire _w2636_ ;
	wire _w2637_ ;
	wire _w2638_ ;
	wire _w2639_ ;
	wire _w2640_ ;
	wire _w2641_ ;
	wire _w2642_ ;
	wire _w2643_ ;
	wire _w2644_ ;
	wire _w2645_ ;
	wire _w2646_ ;
	wire _w2647_ ;
	wire _w2648_ ;
	wire _w2649_ ;
	wire _w2650_ ;
	wire _w2651_ ;
	wire _w2652_ ;
	wire _w2653_ ;
	wire _w2654_ ;
	wire _w2655_ ;
	wire _w2656_ ;
	wire _w2657_ ;
	wire _w2658_ ;
	wire _w2659_ ;
	wire _w2660_ ;
	wire _w2661_ ;
	wire _w2662_ ;
	wire _w2663_ ;
	wire _w2664_ ;
	wire _w2665_ ;
	wire _w2666_ ;
	wire _w2667_ ;
	wire _w2668_ ;
	wire _w2669_ ;
	wire _w2670_ ;
	wire _w2671_ ;
	wire _w2672_ ;
	wire _w2673_ ;
	wire _w2674_ ;
	wire _w2675_ ;
	wire _w2676_ ;
	wire _w2677_ ;
	wire _w2678_ ;
	wire _w2679_ ;
	wire _w2680_ ;
	wire _w2681_ ;
	wire _w2682_ ;
	wire _w2683_ ;
	wire _w2684_ ;
	wire _w2685_ ;
	wire _w2686_ ;
	wire _w2687_ ;
	wire _w2688_ ;
	wire _w2689_ ;
	wire _w2691_ ;
	wire _w2693_ ;
	wire _w2695_ ;
	wire _w2697_ ;
	wire _w2699_ ;
	wire _w2701_ ;
	wire _w2703_ ;
	wire _w2704_ ;
	wire _w2705_ ;
	wire _w2706_ ;
	wire _w2707_ ;
	wire _w2708_ ;
	wire _w2709_ ;
	wire _w2710_ ;
	wire _w2711_ ;
	wire _w2712_ ;
	wire _w2713_ ;
	wire _w2714_ ;
	wire _w2715_ ;
	wire _w2716_ ;
	wire _w2717_ ;
	wire _w2718_ ;
	wire _w2719_ ;
	wire _w2720_ ;
	wire _w2721_ ;
	wire _w2722_ ;
	wire _w2723_ ;
	wire _w2724_ ;
	wire _w2725_ ;
	wire _w2726_ ;
	wire _w2727_ ;
	wire _w2728_ ;
	wire _w2729_ ;
	wire _w2730_ ;
	wire _w2731_ ;
	wire _w2732_ ;
	wire _w2733_ ;
	wire _w2734_ ;
	wire _w2735_ ;
	wire _w2736_ ;
	wire _w2737_ ;
	wire _w2738_ ;
	wire _w2739_ ;
	wire _w2740_ ;
	wire _w2741_ ;
	wire _w2742_ ;
	wire _w2743_ ;
	wire _w2744_ ;
	wire _w2745_ ;
	wire _w2746_ ;
	wire _w2747_ ;
	wire _w2748_ ;
	wire _w2749_ ;
	wire _w2750_ ;
	wire _w2751_ ;
	wire _w2752_ ;
	wire _w2753_ ;
	wire _w2754_ ;
	wire _w2755_ ;
	wire _w2756_ ;
	wire _w2757_ ;
	wire _w2758_ ;
	wire _w2759_ ;
	wire _w2760_ ;
	wire _w2761_ ;
	wire _w2762_ ;
	wire _w2763_ ;
	wire _w2764_ ;
	wire _w2765_ ;
	wire _w2766_ ;
	wire _w2767_ ;
	wire _w2768_ ;
	wire _w2769_ ;
	wire _w2770_ ;
	wire _w2771_ ;
	wire _w2772_ ;
	wire _w2773_ ;
	wire _w2774_ ;
	wire _w2775_ ;
	wire _w2777_ ;
	wire _w2779_ ;
	wire _w2780_ ;
	wire _w2781_ ;
	wire _w2782_ ;
	wire _w2783_ ;
	wire _w2784_ ;
	wire _w2785_ ;
	wire _w2786_ ;
	wire _w2787_ ;
	wire _w2788_ ;
	wire _w2789_ ;
	wire _w2790_ ;
	wire _w2791_ ;
	wire _w2792_ ;
	wire _w2793_ ;
	wire _w2794_ ;
	wire _w2795_ ;
	wire _w2796_ ;
	wire _w2797_ ;
	wire _w2798_ ;
	wire _w2799_ ;
	wire _w2800_ ;
	wire _w2801_ ;
	wire _w2802_ ;
	wire _w2803_ ;
	wire _w2804_ ;
	wire _w2805_ ;
	wire _w2806_ ;
	wire _w2807_ ;
	wire _w2808_ ;
	wire _w2809_ ;
	wire _w2810_ ;
	wire _w2811_ ;
	wire _w2812_ ;
	wire _w2813_ ;
	wire _w2814_ ;
	wire _w2815_ ;
	wire _w2816_ ;
	wire _w2817_ ;
	wire _w2818_ ;
	wire _w2819_ ;
	wire _w2820_ ;
	wire _w2821_ ;
	wire _w2822_ ;
	wire _w2823_ ;
	wire _w2824_ ;
	wire _w2825_ ;
	wire _w2826_ ;
	wire _w2827_ ;
	wire _w2828_ ;
	wire _w2829_ ;
	wire _w2830_ ;
	wire _w2831_ ;
	wire _w2832_ ;
	wire _w2833_ ;
	wire _w2834_ ;
	wire _w2835_ ;
	wire _w2836_ ;
	wire _w2837_ ;
	wire _w2838_ ;
	wire _w2839_ ;
	wire _w2840_ ;
	wire _w2841_ ;
	wire _w2842_ ;
	wire _w2843_ ;
	wire _w2844_ ;
	wire _w2845_ ;
	wire _w2846_ ;
	wire _w2847_ ;
	wire _w2848_ ;
	wire _w2849_ ;
	wire _w2850_ ;
	wire _w2851_ ;
	wire _w2852_ ;
	wire _w2853_ ;
	wire _w2854_ ;
	wire _w2855_ ;
	wire _w2856_ ;
	wire _w2857_ ;
	wire _w2858_ ;
	wire _w2859_ ;
	wire _w2860_ ;
	wire _w2861_ ;
	wire _w2862_ ;
	wire _w2863_ ;
	wire _w2864_ ;
	wire _w2865_ ;
	wire _w2866_ ;
	wire _w2867_ ;
	wire _w2868_ ;
	wire _w2869_ ;
	wire _w2870_ ;
	wire _w2871_ ;
	wire _w2872_ ;
	wire _w2873_ ;
	wire _w2874_ ;
	wire _w2875_ ;
	wire _w2876_ ;
	wire _w2877_ ;
	wire _w2878_ ;
	wire _w2879_ ;
	wire _w2880_ ;
	wire _w2881_ ;
	wire _w2882_ ;
	wire _w2883_ ;
	wire _w2884_ ;
	wire _w2885_ ;
	wire _w2886_ ;
	wire _w2887_ ;
	wire _w2888_ ;
	wire _w2889_ ;
	wire _w2890_ ;
	wire _w2891_ ;
	wire _w2892_ ;
	wire _w2893_ ;
	wire _w2894_ ;
	wire _w2895_ ;
	wire _w2896_ ;
	wire _w2897_ ;
	wire _w2899_ ;
	wire _w2900_ ;
	wire _w2902_ ;
	wire _w2904_ ;
	wire _w2906_ ;
	wire _w2908_ ;
	wire _w2910_ ;
	wire _w2912_ ;
	wire _w2913_ ;
	wire _w2915_ ;
	wire _w2916_ ;
	wire _w2917_ ;
	wire _w2918_ ;
	wire _w2919_ ;
	wire _w2920_ ;
	wire _w2921_ ;
	wire _w2922_ ;
	wire _w2923_ ;
	wire _w2924_ ;
	wire _w2925_ ;
	wire _w2926_ ;
	wire _w2927_ ;
	wire _w2928_ ;
	wire _w2929_ ;
	wire _w2930_ ;
	wire _w2931_ ;
	wire _w2932_ ;
	wire _w2933_ ;
	wire _w2934_ ;
	wire _w2935_ ;
	wire _w2936_ ;
	wire _w2937_ ;
	wire _w2938_ ;
	wire _w2939_ ;
	wire _w2940_ ;
	wire _w2941_ ;
	wire _w2942_ ;
	wire _w2943_ ;
	wire _w2944_ ;
	wire _w2945_ ;
	wire _w2946_ ;
	wire _w2947_ ;
	wire _w2948_ ;
	wire _w2949_ ;
	wire _w2950_ ;
	wire _w2951_ ;
	wire _w2952_ ;
	wire _w2953_ ;
	wire _w2954_ ;
	wire _w2955_ ;
	wire _w2956_ ;
	wire _w2957_ ;
	wire _w2958_ ;
	wire _w2959_ ;
	wire _w2960_ ;
	wire _w2961_ ;
	wire _w2962_ ;
	wire _w2963_ ;
	wire _w2964_ ;
	wire _w2965_ ;
	wire _w2966_ ;
	wire _w2967_ ;
	wire _w2968_ ;
	wire _w2969_ ;
	wire _w2970_ ;
	wire _w2971_ ;
	wire _w2972_ ;
	wire _w2973_ ;
	wire _w2974_ ;
	wire _w2975_ ;
	wire _w2976_ ;
	wire _w2977_ ;
	wire _w2978_ ;
	wire _w2979_ ;
	wire _w2980_ ;
	wire _w2981_ ;
	wire _w2982_ ;
	wire _w2983_ ;
	wire _w2984_ ;
	wire _w2985_ ;
	wire _w2986_ ;
	wire _w2987_ ;
	wire _w2988_ ;
	wire _w2989_ ;
	wire _w2990_ ;
	wire _w2991_ ;
	wire _w2992_ ;
	wire _w2994_ ;
	wire _w2996_ ;
	wire _w2998_ ;
	wire _w3000_ ;
	wire _w3002_ ;
	wire _w3004_ ;
	wire _w3006_ ;
	wire _w3007_ ;
	wire _w3008_ ;
	wire _w3009_ ;
	wire _w3010_ ;
	wire _w3011_ ;
	wire _w3012_ ;
	wire _w3013_ ;
	wire _w3014_ ;
	wire _w3015_ ;
	wire _w3016_ ;
	wire _w3017_ ;
	wire _w3018_ ;
	wire _w3019_ ;
	wire _w3020_ ;
	wire _w3021_ ;
	wire _w3022_ ;
	wire _w3023_ ;
	wire _w3024_ ;
	wire _w3025_ ;
	wire _w3026_ ;
	wire _w3027_ ;
	wire _w3028_ ;
	wire _w3029_ ;
	wire _w3030_ ;
	wire _w3031_ ;
	wire _w3032_ ;
	wire _w3033_ ;
	wire _w3034_ ;
	wire _w3035_ ;
	wire _w3036_ ;
	wire _w3037_ ;
	wire _w3038_ ;
	wire _w3039_ ;
	wire _w3040_ ;
	wire _w3041_ ;
	wire _w3042_ ;
	wire _w3043_ ;
	wire _w3044_ ;
	wire _w3045_ ;
	wire _w3046_ ;
	wire _w3047_ ;
	wire _w3048_ ;
	wire _w3049_ ;
	wire _w3050_ ;
	wire _w3051_ ;
	wire _w3052_ ;
	wire _w3053_ ;
	wire _w3054_ ;
	wire _w3055_ ;
	wire _w3056_ ;
	wire _w3057_ ;
	wire _w3058_ ;
	wire _w3059_ ;
	wire _w3060_ ;
	wire _w3061_ ;
	wire _w3062_ ;
	wire _w3063_ ;
	wire _w3064_ ;
	wire _w3065_ ;
	wire _w3066_ ;
	wire _w3067_ ;
	wire _w3068_ ;
	wire _w3069_ ;
	wire _w3070_ ;
	wire _w3071_ ;
	wire _w3073_ ;
	wire _w3075_ ;
	wire _w3076_ ;
	wire _w3077_ ;
	wire _w3078_ ;
	wire _w3079_ ;
	wire _w3080_ ;
	wire _w3081_ ;
	wire _w3082_ ;
	wire _w3083_ ;
	wire _w3084_ ;
	wire _w3085_ ;
	wire _w3086_ ;
	wire _w3087_ ;
	wire _w3088_ ;
	wire _w3089_ ;
	wire _w3090_ ;
	wire _w3091_ ;
	wire _w3092_ ;
	wire _w3093_ ;
	wire _w3094_ ;
	wire _w3095_ ;
	wire _w3096_ ;
	wire _w3097_ ;
	wire _w3098_ ;
	wire _w3099_ ;
	wire _w3100_ ;
	wire _w3101_ ;
	wire _w3102_ ;
	wire _w3103_ ;
	wire _w3104_ ;
	wire _w3105_ ;
	wire _w3106_ ;
	wire _w3107_ ;
	wire _w3108_ ;
	wire _w3109_ ;
	wire _w3110_ ;
	wire _w3111_ ;
	wire _w3112_ ;
	wire _w3113_ ;
	wire _w3114_ ;
	wire _w3115_ ;
	wire _w3116_ ;
	wire _w3117_ ;
	wire _w3118_ ;
	wire _w3119_ ;
	wire _w3120_ ;
	wire _w3121_ ;
	wire _w3122_ ;
	wire _w3123_ ;
	wire _w3124_ ;
	wire _w3125_ ;
	wire _w3126_ ;
	wire _w3127_ ;
	wire _w3128_ ;
	wire _w3129_ ;
	wire _w3130_ ;
	wire _w3131_ ;
	wire _w3132_ ;
	wire _w3133_ ;
	wire _w3134_ ;
	wire _w3135_ ;
	wire _w3136_ ;
	wire _w3137_ ;
	wire _w3138_ ;
	wire _w3139_ ;
	wire _w3140_ ;
	wire _w3141_ ;
	wire _w3142_ ;
	wire _w3143_ ;
	wire _w3144_ ;
	wire _w3145_ ;
	wire _w3146_ ;
	wire _w3147_ ;
	wire _w3148_ ;
	wire _w3149_ ;
	wire _w3150_ ;
	wire _w3151_ ;
	wire _w3152_ ;
	wire _w3153_ ;
	wire _w3154_ ;
	wire _w3155_ ;
	wire _w3156_ ;
	wire _w3157_ ;
	wire _w3158_ ;
	wire _w3159_ ;
	wire _w3160_ ;
	wire _w3161_ ;
	wire _w3162_ ;
	wire _w3163_ ;
	wire _w3164_ ;
	wire _w3165_ ;
	wire _w3166_ ;
	wire _w3167_ ;
	wire _w3168_ ;
	wire _w3169_ ;
	wire _w3170_ ;
	wire _w3171_ ;
	wire _w3172_ ;
	wire _w3173_ ;
	wire _w3174_ ;
	wire _w3175_ ;
	wire _w3176_ ;
	wire _w3178_ ;
	wire _w3179_ ;
	wire _w3180_ ;
	wire _w3181_ ;
	wire _w3182_ ;
	wire _w3183_ ;
	wire _w3184_ ;
	wire _w3185_ ;
	wire _w3186_ ;
	wire _w3187_ ;
	wire _w3188_ ;
	wire _w3189_ ;
	wire _w3190_ ;
	wire _w3191_ ;
	wire _w3192_ ;
	wire _w3193_ ;
	wire _w3194_ ;
	wire _w3196_ ;
	wire _w3198_ ;
	wire _w3200_ ;
	wire _w3201_ ;
	wire _w3203_ ;
	wire _w3205_ ;
	wire _w3206_ ;
	wire _w3207_ ;
	wire _w3208_ ;
	wire _w3209_ ;
	wire _w3211_ ;
	wire _w3212_ ;
	wire _w3213_ ;
	wire _w3214_ ;
	wire _w3215_ ;
	wire _w3216_ ;
	wire _w3218_ ;
	wire _w3219_ ;
	wire _w3220_ ;
	wire _w3221_ ;
	wire _w3222_ ;
	wire _w3223_ ;
	wire _w3224_ ;
	wire _w3225_ ;
	wire _w3226_ ;
	wire _w3227_ ;
	wire _w3228_ ;
	wire _w3229_ ;
	wire _w3230_ ;
	wire _w3231_ ;
	wire _w3232_ ;
	wire _w3233_ ;
	wire _w3234_ ;
	wire _w3235_ ;
	wire _w3236_ ;
	wire _w3237_ ;
	wire _w3238_ ;
	wire _w3239_ ;
	wire _w3240_ ;
	wire _w3241_ ;
	wire _w3242_ ;
	wire _w3243_ ;
	wire _w3244_ ;
	wire _w3245_ ;
	wire _w3246_ ;
	wire _w3247_ ;
	wire _w3248_ ;
	wire _w3249_ ;
	wire _w3250_ ;
	wire _w3251_ ;
	wire _w3252_ ;
	wire _w3253_ ;
	wire _w3254_ ;
	wire _w3255_ ;
	wire _w3256_ ;
	wire _w3257_ ;
	wire _w3258_ ;
	wire _w3259_ ;
	wire _w3260_ ;
	wire _w3261_ ;
	wire _w3262_ ;
	wire _w3263_ ;
	wire _w3264_ ;
	wire _w3265_ ;
	wire _w3266_ ;
	wire _w3267_ ;
	wire _w3268_ ;
	wire _w3269_ ;
	wire _w3270_ ;
	wire _w3271_ ;
	wire _w3272_ ;
	wire _w3273_ ;
	wire _w3274_ ;
	wire _w3275_ ;
	wire _w3276_ ;
	wire _w3277_ ;
	wire _w3278_ ;
	wire _w3279_ ;
	wire _w3280_ ;
	wire _w3281_ ;
	wire _w3282_ ;
	wire _w3283_ ;
	wire _w3284_ ;
	wire _w3285_ ;
	wire _w3286_ ;
	wire _w3287_ ;
	wire _w3288_ ;
	wire _w3289_ ;
	wire _w3290_ ;
	wire _w3291_ ;
	wire _w3292_ ;
	wire _w3293_ ;
	wire _w3294_ ;
	wire _w3295_ ;
	wire _w3296_ ;
	wire _w3297_ ;
	wire _w3298_ ;
	wire _w3299_ ;
	wire _w3300_ ;
	wire _w3301_ ;
	wire _w3302_ ;
	wire _w3303_ ;
	wire _w3304_ ;
	wire _w3305_ ;
	wire _w3306_ ;
	wire _w3307_ ;
	wire _w3308_ ;
	wire _w3309_ ;
	wire _w3310_ ;
	wire _w3311_ ;
	wire _w3312_ ;
	wire _w3313_ ;
	wire _w3314_ ;
	wire _w3315_ ;
	wire _w3316_ ;
	wire _w3317_ ;
	wire _w3318_ ;
	wire _w3319_ ;
	wire _w3320_ ;
	wire _w3321_ ;
	wire _w3322_ ;
	wire _w3323_ ;
	wire _w3324_ ;
	wire _w3325_ ;
	wire _w3326_ ;
	wire _w3327_ ;
	wire _w3328_ ;
	wire _w3329_ ;
	wire _w3330_ ;
	wire _w3331_ ;
	wire _w3332_ ;
	wire _w3333_ ;
	wire _w3334_ ;
	wire _w3335_ ;
	wire _w3336_ ;
	wire _w3337_ ;
	wire _w3338_ ;
	wire _w3339_ ;
	wire _w3340_ ;
	wire _w3341_ ;
	wire _w3342_ ;
	wire _w3343_ ;
	wire _w3344_ ;
	wire _w3345_ ;
	wire _w3346_ ;
	wire _w3347_ ;
	wire _w3348_ ;
	wire _w3349_ ;
	wire _w3350_ ;
	wire _w3351_ ;
	wire _w3352_ ;
	wire _w3353_ ;
	wire _w3354_ ;
	wire _w3355_ ;
	wire _w3356_ ;
	wire _w3357_ ;
	wire _w3358_ ;
	wire _w3359_ ;
	wire _w3360_ ;
	wire _w3361_ ;
	wire _w3362_ ;
	wire _w3363_ ;
	wire _w3364_ ;
	wire _w3365_ ;
	wire _w3366_ ;
	wire _w3367_ ;
	wire _w3368_ ;
	wire _w3370_ ;
	wire _w3372_ ;
	wire _w3373_ ;
	wire _w3374_ ;
	wire _w3375_ ;
	wire _w3376_ ;
	wire _w3377_ ;
	wire _w3378_ ;
	wire _w3379_ ;
	wire _w3380_ ;
	wire _w3381_ ;
	wire _w3382_ ;
	wire _w3383_ ;
	wire _w3384_ ;
	wire _w3385_ ;
	wire _w3386_ ;
	wire _w3387_ ;
	wire _w3388_ ;
	wire _w3389_ ;
	wire _w3390_ ;
	wire _w3391_ ;
	wire _w3392_ ;
	wire _w3393_ ;
	wire _w3394_ ;
	wire _w3395_ ;
	wire _w3396_ ;
	wire _w3397_ ;
	wire _w3398_ ;
	wire _w3399_ ;
	wire _w3400_ ;
	wire _w3401_ ;
	wire _w3402_ ;
	wire _w3403_ ;
	wire _w3404_ ;
	wire _w3405_ ;
	wire _w3406_ ;
	wire _w3407_ ;
	wire _w3408_ ;
	wire _w3409_ ;
	wire _w3410_ ;
	wire _w3411_ ;
	wire _w3412_ ;
	wire _w3413_ ;
	wire _w3414_ ;
	wire _w3415_ ;
	wire _w3416_ ;
	wire _w3417_ ;
	wire _w3418_ ;
	wire _w3419_ ;
	wire _w3420_ ;
	wire _w3421_ ;
	wire _w3422_ ;
	wire _w3423_ ;
	wire _w3424_ ;
	wire _w3425_ ;
	wire _w3426_ ;
	wire _w3427_ ;
	wire _w3428_ ;
	wire _w3429_ ;
	wire _w3430_ ;
	wire _w3431_ ;
	wire _w3432_ ;
	wire _w3433_ ;
	wire _w3434_ ;
	wire _w3435_ ;
	wire _w3436_ ;
	wire _w3437_ ;
	wire _w3438_ ;
	wire _w3439_ ;
	wire _w3440_ ;
	wire _w3441_ ;
	wire _w3442_ ;
	wire _w3443_ ;
	wire _w3444_ ;
	wire _w3445_ ;
	wire _w3446_ ;
	wire _w3447_ ;
	wire _w3448_ ;
	wire _w3449_ ;
	wire _w3450_ ;
	wire _w3451_ ;
	wire _w3452_ ;
	wire _w3453_ ;
	wire _w3454_ ;
	wire _w3455_ ;
	wire _w3456_ ;
	wire _w3457_ ;
	wire _w3458_ ;
	wire _w3459_ ;
	wire _w3460_ ;
	wire _w3461_ ;
	wire _w3462_ ;
	wire _w3463_ ;
	wire _w3464_ ;
	wire _w3465_ ;
	wire _w3466_ ;
	wire _w3467_ ;
	wire _w3468_ ;
	wire _w3469_ ;
	wire _w3470_ ;
	wire _w3471_ ;
	wire _w3472_ ;
	wire _w3473_ ;
	wire _w3474_ ;
	wire _w3475_ ;
	wire _w3476_ ;
	wire _w3477_ ;
	wire _w3478_ ;
	wire _w3479_ ;
	wire _w3480_ ;
	wire _w3481_ ;
	wire _w3482_ ;
	wire _w3484_ ;
	wire _w3486_ ;
	wire _w3488_ ;
	wire _w3489_ ;
	wire _w3491_ ;
	wire _w3493_ ;
	wire _w3495_ ;
	wire _w3497_ ;
	wire _w3499_ ;
	wire _w3500_ ;
	wire _w3501_ ;
	wire _w3502_ ;
	wire _w3503_ ;
	wire _w3504_ ;
	wire _w3505_ ;
	wire _w3506_ ;
	wire _w3507_ ;
	wire _w3508_ ;
	wire _w3509_ ;
	wire _w3510_ ;
	wire _w3511_ ;
	wire _w3512_ ;
	wire _w3513_ ;
	wire _w3514_ ;
	wire _w3515_ ;
	wire _w3516_ ;
	wire _w3517_ ;
	wire _w3518_ ;
	wire _w3519_ ;
	wire _w3520_ ;
	wire _w3521_ ;
	wire _w3522_ ;
	wire _w3523_ ;
	wire _w3524_ ;
	wire _w3525_ ;
	wire _w3526_ ;
	wire _w3527_ ;
	wire _w3528_ ;
	wire _w3529_ ;
	wire _w3530_ ;
	wire _w3531_ ;
	wire _w3532_ ;
	wire _w3533_ ;
	wire _w3534_ ;
	wire _w3535_ ;
	wire _w3536_ ;
	wire _w3537_ ;
	LUT1 #(
		.INIT('h1)
	) name0 (
		\g101_reg/NET0131 ,
		_w16_
	);
	LUT1 #(
		.INIT('h1)
	) name1 (
		\g105_reg/NET0131 ,
		_w31_
	);
	LUT1 #(
		.INIT('h1)
	) name2 (
		\g109_reg/NET0131 ,
		_w51_
	);
	LUT1 #(
		.INIT('h1)
	) name3 (
		\g1138_reg/NET0131 ,
		_w69_
	);
	LUT1 #(
		.INIT('h1)
	) name4 (
		\g113_reg/NET0131 ,
		_w71_
	);
	LUT1 #(
		.INIT('h1)
	) name5 (
		\g1140_reg/NET0131 ,
		_w73_
	);
	LUT1 #(
		.INIT('h1)
	) name6 (
		\g117_reg/NET0131 ,
		_w86_
	);
	LUT1 #(
		.INIT('h1)
	) name7 (
		\g121_reg/NET0131 ,
		_w101_
	);
	LUT1 #(
		.INIT('h1)
	) name8 (
		\g125_reg/NET0131 ,
		_w120_
	);
	LUT1 #(
		.INIT('h1)
	) name9 (
		\g1471_reg/NET0131 ,
		_w222_
	);
	LUT1 #(
		.INIT('h1)
	) name10 (
		\g1476_reg/NET0131 ,
		_w224_
	);
	LUT1 #(
		.INIT('h1)
	) name11 (
		\g1481_reg/NET0131 ,
		_w227_
	);
	LUT1 #(
		.INIT('h1)
	) name12 (
		\g1486_reg/NET0131 ,
		_w229_
	);
	LUT1 #(
		.INIT('h1)
	) name13 (
		\g1491_reg/NET0131 ,
		_w232_
	);
	LUT1 #(
		.INIT('h1)
	) name14 (
		\g1496_reg/NET0131 ,
		_w234_
	);
	LUT1 #(
		.INIT('h1)
	) name15 (
		\g1501_reg/NET0131 ,
		_w237_
	);
	LUT1 #(
		.INIT('h1)
	) name16 (
		\g1506_reg/NET0131 ,
		_w239_
	);
	LUT1 #(
		.INIT('h1)
	) name17 (
		\g1660_reg/NET0131 ,
		_w333_
	);
	LUT1 #(
		.INIT('h1)
	) name18 (
		\g1662_reg/NET0131 ,
		_w335_
	);
	LUT1 #(
		.INIT('h1)
	) name19 (
		\g1664_reg/NET0131 ,
		_w337_
	);
	LUT1 #(
		.INIT('h1)
	) name20 (
		\g1666_reg/NET0131 ,
		_w339_
	);
	LUT1 #(
		.INIT('h1)
	) name21 (
		\g1668_reg/NET0131 ,
		_w341_
	);
	LUT1 #(
		.INIT('h1)
	) name22 (
		\g1670_reg/NET0131 ,
		_w343_
	);
	LUT1 #(
		.INIT('h1)
	) name23 (
		\g1672_reg/NET0131 ,
		_w345_
	);
	LUT1 #(
		.INIT('h1)
	) name24 (
		\g1832_reg/NET0131 ,
		_w419_
	);
	LUT1 #(
		.INIT('h1)
	) name25 (
		\g1834_reg/NET0131 ,
		_w421_
	);
	LUT1 #(
		.INIT('h1)
	) name26 (
		\g2165_reg/NET0131 ,
		_w541_
	);
	LUT1 #(
		.INIT('h1)
	) name27 (
		\g2170_reg/NET0131 ,
		_w544_
	);
	LUT1 #(
		.INIT('h1)
	) name28 (
		\g2175_reg/NET0131 ,
		_w546_
	);
	LUT1 #(
		.INIT('h1)
	) name29 (
		\g2180_reg/NET0131 ,
		_w548_
	);
	LUT1 #(
		.INIT('h1)
	) name30 (
		\g2185_reg/NET0131 ,
		_w550_
	);
	LUT1 #(
		.INIT('h1)
	) name31 (
		\g2190_reg/NET0131 ,
		_w552_
	);
	LUT1 #(
		.INIT('h1)
	) name32 (
		\g2195_reg/NET0131 ,
		_w554_
	);
	LUT1 #(
		.INIT('h1)
	) name33 (
		\g2200_reg/NET0131 ,
		_w557_
	);
	LUT1 #(
		.INIT('h1)
	) name34 (
		\g2354_reg/NET0131 ,
		_w636_
	);
	LUT1 #(
		.INIT('h1)
	) name35 (
		\g2356_reg/NET0131 ,
		_w638_
	);
	LUT1 #(
		.INIT('h1)
	) name36 (
		\g2358_reg/NET0131 ,
		_w640_
	);
	LUT1 #(
		.INIT('h1)
	) name37 (
		\g2360_reg/NET0131 ,
		_w642_
	);
	LUT1 #(
		.INIT('h1)
	) name38 (
		\g2362_reg/NET0131 ,
		_w644_
	);
	LUT1 #(
		.INIT('h1)
	) name39 (
		\g2364_reg/NET0131 ,
		_w646_
	);
	LUT1 #(
		.INIT('h1)
	) name40 (
		\g2366_reg/NET0131 ,
		_w648_
	);
	LUT1 #(
		.INIT('h1)
	) name41 (
		\g2526_reg/NET0131 ,
		_w715_
	);
	LUT1 #(
		.INIT('h1)
	) name42 (
		\g2528_reg/NET0131 ,
		_w717_
	);
	LUT1 #(
		.INIT('h1)
	) name43 (
		\g279_reg/NET0131 ,
		_w820_
	);
	LUT1 #(
		.INIT('h1)
	) name44 (
		\g281_reg/NET0131 ,
		_w838_
	);
	LUT1 #(
		.INIT('h1)
	) name45 (
		\g283_reg/NET0131 ,
		_w840_
	);
	LUT1 #(
		.INIT('h1)
	) name46 (
		\g285_reg/NET0131 ,
		_w842_
	);
	LUT1 #(
		.INIT('h1)
	) name47 (
		\g2879_reg/NET0131 ,
		_w845_
	);
	LUT1 #(
		.INIT('h1)
	) name48 (
		\g287_reg/NET0131 ,
		_w847_
	);
	LUT1 #(
		.INIT('h1)
	) name49 (
		\g289_reg/NET0131 ,
		_w853_
	);
	LUT1 #(
		.INIT('h1)
	) name50 (
		\g291_reg/NET0131 ,
		_w860_
	);
	LUT1 #(
		.INIT('h1)
	) name51 (
		\g451_reg/NET0131 ,
		_w1012_
	);
	LUT1 #(
		.INIT('h1)
	) name52 (
		\g453_reg/NET0131 ,
		_w1014_
	);
	LUT1 #(
		.INIT('h1)
	) name53 (
		\g785_reg/NET0131 ,
		_w1126_
	);
	LUT1 #(
		.INIT('h1)
	) name54 (
		\g789_reg/NET0131 ,
		_w1128_
	);
	LUT1 #(
		.INIT('h1)
	) name55 (
		\g793_reg/NET0131 ,
		_w1130_
	);
	LUT1 #(
		.INIT('h1)
	) name56 (
		\g797_reg/NET0131 ,
		_w1133_
	);
	LUT1 #(
		.INIT('h1)
	) name57 (
		\g801_reg/NET0131 ,
		_w1135_
	);
	LUT1 #(
		.INIT('h1)
	) name58 (
		\g805_reg/NET0131 ,
		_w1137_
	);
	LUT1 #(
		.INIT('h1)
	) name59 (
		\g809_reg/NET0131 ,
		_w1139_
	);
	LUT1 #(
		.INIT('h1)
	) name60 (
		\g813_reg/NET0131 ,
		_w1141_
	);
	LUT1 #(
		.INIT('h1)
	) name61 (
		\g966_reg/NET0131 ,
		_w1231_
	);
	LUT1 #(
		.INIT('h1)
	) name62 (
		\g968_reg/NET0131 ,
		_w1233_
	);
	LUT1 #(
		.INIT('h1)
	) name63 (
		\g970_reg/NET0131 ,
		_w1235_
	);
	LUT1 #(
		.INIT('h1)
	) name64 (
		\g972_reg/NET0131 ,
		_w1237_
	);
	LUT1 #(
		.INIT('h1)
	) name65 (
		\g974_reg/NET0131 ,
		_w1239_
	);
	LUT1 #(
		.INIT('h1)
	) name66 (
		\g976_reg/NET0131 ,
		_w1241_
	);
	LUT1 #(
		.INIT('h1)
	) name67 (
		\g978_reg/NET0131 ,
		_w1243_
	);
	LUT1 #(
		.INIT('h1)
	) name68 (
		\g97_reg/NET0131 ,
		_w1245_
	);
	LUT3 #(
		.INIT('h73)
	) name69 (
		\g2986_reg/NET0131 ,
		\g2987_reg/NET0131 ,
		\g5388_pad ,
		_w1250_
	);
	LUT2 #(
		.INIT('h2)
	) name70 (
		\g1092_reg/NET0131 ,
		\g2394_reg/NET0131 ,
		_w1251_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name71 (
		\g1088_reg/NET0131 ,
		\g2393_reg/NET0131 ,
		\g2395_reg/NET0131 ,
		\g7961_pad ,
		_w1252_
	);
	LUT2 #(
		.INIT('h4)
	) name72 (
		_w1251_,
		_w1252_,
		_w1253_
	);
	LUT2 #(
		.INIT('h8)
	) name73 (
		\g1092_reg/NET0131 ,
		\g2336_reg/NET0131 ,
		_w1254_
	);
	LUT4 #(
		.INIT('h135f)
	) name74 (
		\g1088_reg/NET0131 ,
		\g2333_reg/NET0131 ,
		\g2339_reg/NET0131 ,
		\g7961_pad ,
		_w1255_
	);
	LUT2 #(
		.INIT('h4)
	) name75 (
		_w1254_,
		_w1255_,
		_w1256_
	);
	LUT3 #(
		.INIT('h9a)
	) name76 (
		\g2200_reg/NET0131 ,
		_w1254_,
		_w1255_,
		_w1257_
	);
	LUT2 #(
		.INIT('h8)
	) name77 (
		\g2306_reg/NET0131 ,
		\g7961_pad ,
		_w1258_
	);
	LUT4 #(
		.INIT('h153f)
	) name78 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2309_reg/NET0131 ,
		\g2312_reg/NET0131 ,
		_w1259_
	);
	LUT2 #(
		.INIT('h4)
	) name79 (
		_w1258_,
		_w1259_,
		_w1260_
	);
	LUT3 #(
		.INIT('h9a)
	) name80 (
		\g2170_reg/NET0131 ,
		_w1258_,
		_w1259_,
		_w1261_
	);
	LUT2 #(
		.INIT('h8)
	) name81 (
		_w1257_,
		_w1261_,
		_w1262_
	);
	LUT4 #(
		.INIT('h135f)
	) name82 (
		\g1088_reg/NET0131 ,
		\g2324_reg/NET0131 ,
		\g2330_reg/NET0131 ,
		\g7961_pad ,
		_w1263_
	);
	LUT2 #(
		.INIT('h8)
	) name83 (
		\g1092_reg/NET0131 ,
		\g2327_reg/NET0131 ,
		_w1264_
	);
	LUT2 #(
		.INIT('h2)
	) name84 (
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT3 #(
		.INIT('ha6)
	) name85 (
		\g2190_reg/NET0131 ,
		_w1263_,
		_w1264_,
		_w1266_
	);
	LUT2 #(
		.INIT('h2)
	) name86 (
		\g1088_reg/NET0131 ,
		\g2247_reg/NET0131 ,
		_w1267_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name87 (
		\g1092_reg/NET0131 ,
		\g2248_reg/NET0131 ,
		\g2249_reg/NET0131 ,
		\g7961_pad ,
		_w1268_
	);
	LUT2 #(
		.INIT('h4)
	) name88 (
		_w1267_,
		_w1268_,
		_w1269_
	);
	LUT2 #(
		.INIT('h8)
	) name89 (
		\g2342_reg/NET0131 ,
		\g7961_pad ,
		_w1270_
	);
	LUT4 #(
		.INIT('h153f)
	) name90 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2345_reg/NET0131 ,
		\g2348_reg/NET0131 ,
		_w1271_
	);
	LUT2 #(
		.INIT('h4)
	) name91 (
		_w1270_,
		_w1271_,
		_w1272_
	);
	LUT4 #(
		.INIT('h4b44)
	) name92 (
		_w1267_,
		_w1268_,
		_w1270_,
		_w1271_,
		_w1273_
	);
	LUT4 #(
		.INIT('h153f)
	) name93 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2318_reg/NET0131 ,
		\g2321_reg/NET0131 ,
		_w1274_
	);
	LUT2 #(
		.INIT('h8)
	) name94 (
		\g2315_reg/NET0131 ,
		\g7961_pad ,
		_w1275_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w1274_,
		_w1275_,
		_w1276_
	);
	LUT3 #(
		.INIT('ha6)
	) name96 (
		\g2180_reg/NET0131 ,
		_w1274_,
		_w1275_,
		_w1277_
	);
	LUT3 #(
		.INIT('h45)
	) name97 (
		_w1266_,
		_w1273_,
		_w1277_,
		_w1278_
	);
	LUT2 #(
		.INIT('h4)
	) name98 (
		_w1262_,
		_w1278_,
		_w1279_
	);
	LUT4 #(
		.INIT('h135f)
	) name99 (
		_w1257_,
		_w1261_,
		_w1266_,
		_w1277_,
		_w1280_
	);
	LUT3 #(
		.INIT('h15)
	) name100 (
		_w1261_,
		_w1266_,
		_w1277_,
		_w1281_
	);
	LUT4 #(
		.INIT('h223f)
	) name101 (
		_w1257_,
		_w1273_,
		_w1280_,
		_w1281_,
		_w1282_
	);
	LUT2 #(
		.INIT('h8)
	) name102 (
		\g1088_reg/NET0131 ,
		\g2285_reg/NET0131 ,
		_w1283_
	);
	LUT4 #(
		.INIT('h135f)
	) name103 (
		\g1092_reg/NET0131 ,
		\g2279_reg/NET0131 ,
		\g2282_reg/NET0131 ,
		\g7961_pad ,
		_w1284_
	);
	LUT2 #(
		.INIT('h4)
	) name104 (
		_w1283_,
		_w1284_,
		_w1285_
	);
	LUT3 #(
		.INIT('h9a)
	) name105 (
		\g2185_reg/NET0131 ,
		_w1283_,
		_w1284_,
		_w1286_
	);
	LUT4 #(
		.INIT('h2000)
	) name106 (
		_w1266_,
		_w1273_,
		_w1277_,
		_w1286_,
		_w1287_
	);
	LUT2 #(
		.INIT('h8)
	) name107 (
		\g1092_reg/NET0131 ,
		\g2291_reg/NET0131 ,
		_w1288_
	);
	LUT4 #(
		.INIT('h135f)
	) name108 (
		\g1088_reg/NET0131 ,
		\g2288_reg/NET0131 ,
		\g2294_reg/NET0131 ,
		\g7961_pad ,
		_w1289_
	);
	LUT2 #(
		.INIT('h4)
	) name109 (
		_w1288_,
		_w1289_,
		_w1290_
	);
	LUT3 #(
		.INIT('h9a)
	) name110 (
		\g2195_reg/NET0131 ,
		_w1288_,
		_w1289_,
		_w1291_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		\g1088_reg/NET0131 ,
		\g2250_reg/NET0131 ,
		_w1292_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name112 (
		\g1092_reg/NET0131 ,
		\g2251_reg/NET0131 ,
		\g2252_reg/NET0131 ,
		\g7961_pad ,
		_w1293_
	);
	LUT2 #(
		.INIT('h4)
	) name113 (
		_w1292_,
		_w1293_,
		_w1294_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\g2297_reg/NET0131 ,
		\g7961_pad ,
		_w1295_
	);
	LUT4 #(
		.INIT('h153f)
	) name115 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2300_reg/NET0131 ,
		\g2303_reg/NET0131 ,
		_w1296_
	);
	LUT2 #(
		.INIT('h4)
	) name116 (
		_w1295_,
		_w1296_,
		_w1297_
	);
	LUT4 #(
		.INIT('h4b44)
	) name117 (
		_w1292_,
		_w1293_,
		_w1295_,
		_w1296_,
		_w1298_
	);
	LUT2 #(
		.INIT('h2)
	) name118 (
		_w1291_,
		_w1298_,
		_w1299_
	);
	LUT4 #(
		.INIT('h135f)
	) name119 (
		\g1088_reg/NET0131 ,
		\g2261_reg/NET0131 ,
		\g2267_reg/NET0131 ,
		\g7961_pad ,
		_w1300_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		\g1092_reg/NET0131 ,
		\g2264_reg/NET0131 ,
		_w1301_
	);
	LUT2 #(
		.INIT('h2)
	) name121 (
		_w1300_,
		_w1301_,
		_w1302_
	);
	LUT3 #(
		.INIT('ha6)
	) name122 (
		\g2165_reg/NET0131 ,
		_w1300_,
		_w1301_,
		_w1303_
	);
	LUT2 #(
		.INIT('h8)
	) name123 (
		\g2270_reg/NET0131 ,
		\g7961_pad ,
		_w1304_
	);
	LUT4 #(
		.INIT('h153f)
	) name124 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2273_reg/NET0131 ,
		\g2276_reg/NET0131 ,
		_w1305_
	);
	LUT2 #(
		.INIT('h4)
	) name125 (
		_w1304_,
		_w1305_,
		_w1306_
	);
	LUT3 #(
		.INIT('h9a)
	) name126 (
		\g2175_reg/NET0131 ,
		_w1304_,
		_w1305_,
		_w1307_
	);
	LUT4 #(
		.INIT('h8000)
	) name127 (
		_w1257_,
		_w1261_,
		_w1303_,
		_w1307_,
		_w1308_
	);
	LUT3 #(
		.INIT('h80)
	) name128 (
		_w1287_,
		_w1299_,
		_w1308_,
		_w1309_
	);
	LUT4 #(
		.INIT('haa8a)
	) name129 (
		_w1253_,
		_w1279_,
		_w1282_,
		_w1309_,
		_w1310_
	);
	LUT2 #(
		.INIT('h2)
	) name130 (
		\g1092_reg/NET0131 ,
		\g2246_reg/NET0131 ,
		_w1311_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name131 (
		\g1088_reg/NET0131 ,
		\g2244_reg/NET0131 ,
		\g2245_reg/NET0131 ,
		\g7961_pad ,
		_w1312_
	);
	LUT2 #(
		.INIT('h4)
	) name132 (
		_w1311_,
		_w1312_,
		_w1313_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name133 (
		\g1088_reg/NET0131 ,
		\g2229_reg/NET0131 ,
		\g2230_reg/NET0131 ,
		\g7961_pad ,
		_w1314_
	);
	LUT2 #(
		.INIT('h2)
	) name134 (
		\g1092_reg/NET0131 ,
		\g2231_reg/NET0131 ,
		_w1315_
	);
	LUT3 #(
		.INIT('ha6)
	) name135 (
		\g2195_reg/NET0131 ,
		_w1314_,
		_w1315_,
		_w1316_
	);
	LUT2 #(
		.INIT('h2)
	) name136 (
		\g1092_reg/NET0131 ,
		\g2237_reg/NET0131 ,
		_w1317_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name137 (
		\g1088_reg/NET0131 ,
		\g2235_reg/NET0131 ,
		\g2236_reg/NET0131 ,
		\g7961_pad ,
		_w1318_
	);
	LUT4 #(
		.INIT('h4b44)
	) name138 (
		_w1292_,
		_w1293_,
		_w1317_,
		_w1318_,
		_w1319_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name139 (
		\g1088_reg/NET0131 ,
		\g2223_reg/NET0131 ,
		\g2224_reg/NET0131 ,
		\g7961_pad ,
		_w1320_
	);
	LUT2 #(
		.INIT('h2)
	) name140 (
		\g1092_reg/NET0131 ,
		\g2225_reg/NET0131 ,
		_w1321_
	);
	LUT3 #(
		.INIT('ha6)
	) name141 (
		\g2185_reg/NET0131 ,
		_w1320_,
		_w1321_,
		_w1322_
	);
	LUT4 #(
		.INIT('hf531)
	) name142 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2205_reg/NET0131 ,
		\g2207_reg/NET0131 ,
		_w1323_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		\g2206_reg/NET0131 ,
		\g7961_pad ,
		_w1324_
	);
	LUT3 #(
		.INIT('ha6)
	) name144 (
		\g2165_reg/NET0131 ,
		_w1323_,
		_w1324_,
		_w1325_
	);
	LUT4 #(
		.INIT('h2000)
	) name145 (
		_w1316_,
		_w1319_,
		_w1322_,
		_w1325_,
		_w1326_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name146 (
		\g1088_reg/NET0131 ,
		\g2232_reg/NET0131 ,
		\g2233_reg/NET0131 ,
		\g7961_pad ,
		_w1327_
	);
	LUT2 #(
		.INIT('h2)
	) name147 (
		\g1092_reg/NET0131 ,
		\g2234_reg/NET0131 ,
		_w1328_
	);
	LUT3 #(
		.INIT('ha6)
	) name148 (
		\g2200_reg/NET0131 ,
		_w1327_,
		_w1328_,
		_w1329_
	);
	LUT4 #(
		.INIT('hf531)
	) name149 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2208_reg/NET0131 ,
		\g2210_reg/NET0131 ,
		_w1330_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		\g2209_reg/NET0131 ,
		\g7961_pad ,
		_w1331_
	);
	LUT3 #(
		.INIT('ha6)
	) name151 (
		\g2170_reg/NET0131 ,
		_w1330_,
		_w1331_,
		_w1332_
	);
	LUT3 #(
		.INIT('h8a)
	) name152 (
		\g1563_reg/NET0131 ,
		_w1311_,
		_w1312_,
		_w1333_
	);
	LUT4 #(
		.INIT('hf531)
	) name153 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2220_reg/NET0131 ,
		\g2222_reg/NET0131 ,
		_w1334_
	);
	LUT2 #(
		.INIT('h4)
	) name154 (
		\g2221_reg/NET0131 ,
		\g7961_pad ,
		_w1335_
	);
	LUT3 #(
		.INIT('ha6)
	) name155 (
		\g2180_reg/NET0131 ,
		_w1334_,
		_w1335_,
		_w1336_
	);
	LUT4 #(
		.INIT('h8000)
	) name156 (
		_w1329_,
		_w1332_,
		_w1333_,
		_w1336_,
		_w1337_
	);
	LUT2 #(
		.INIT('h8)
	) name157 (
		_w1326_,
		_w1337_,
		_w1338_
	);
	LUT2 #(
		.INIT('h8)
	) name158 (
		_w1286_,
		_w1291_,
		_w1339_
	);
	LUT3 #(
		.INIT('h2a)
	) name159 (
		_w1298_,
		_w1303_,
		_w1307_,
		_w1340_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		_w1298_,
		_w1307_,
		_w1341_
	);
	LUT3 #(
		.INIT('h15)
	) name161 (
		_w1286_,
		_w1291_,
		_w1303_,
		_w1342_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name162 (
		_w1339_,
		_w1340_,
		_w1341_,
		_w1342_,
		_w1343_
	);
	LUT4 #(
		.INIT('h51f3)
	) name163 (
		_w1286_,
		_w1291_,
		_w1298_,
		_w1307_,
		_w1344_
	);
	LUT2 #(
		.INIT('h4)
	) name164 (
		_w1303_,
		_w1344_,
		_w1345_
	);
	LUT4 #(
		.INIT('hf531)
	) name165 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2217_reg/NET0131 ,
		\g2219_reg/NET0131 ,
		_w1346_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		\g2218_reg/NET0131 ,
		\g7961_pad ,
		_w1347_
	);
	LUT3 #(
		.INIT('ha6)
	) name167 (
		\g2175_reg/NET0131 ,
		_w1346_,
		_w1347_,
		_w1348_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name168 (
		\g1088_reg/NET0131 ,
		\g2226_reg/NET0131 ,
		\g2227_reg/NET0131 ,
		\g7961_pad ,
		_w1349_
	);
	LUT2 #(
		.INIT('h2)
	) name169 (
		\g1092_reg/NET0131 ,
		\g2228_reg/NET0131 ,
		_w1350_
	);
	LUT3 #(
		.INIT('ha6)
	) name170 (
		\g2190_reg/NET0131 ,
		_w1349_,
		_w1350_,
		_w1351_
	);
	LUT2 #(
		.INIT('h8)
	) name171 (
		_w1348_,
		_w1351_,
		_w1352_
	);
	LUT2 #(
		.INIT('h2)
	) name172 (
		\g1092_reg/NET0131 ,
		\g2240_reg/NET0131 ,
		_w1353_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name173 (
		\g1088_reg/NET0131 ,
		\g2238_reg/NET0131 ,
		\g2239_reg/NET0131 ,
		\g7961_pad ,
		_w1354_
	);
	LUT4 #(
		.INIT('hb4bb)
	) name174 (
		_w1267_,
		_w1268_,
		_w1353_,
		_w1354_,
		_w1355_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		\g1092_reg/NET0131 ,
		\g2398_reg/NET0131 ,
		_w1356_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name176 (
		\g1088_reg/NET0131 ,
		\g2396_reg/NET0131 ,
		\g2397_reg/NET0131 ,
		\g7961_pad ,
		_w1357_
	);
	LUT2 #(
		.INIT('h4)
	) name177 (
		_w1356_,
		_w1357_,
		_w1358_
	);
	LUT4 #(
		.INIT('h0080)
	) name178 (
		_w1348_,
		_w1351_,
		_w1355_,
		_w1358_,
		_w1359_
	);
	LUT3 #(
		.INIT('hb0)
	) name179 (
		_w1303_,
		_w1344_,
		_w1359_,
		_w1360_
	);
	LUT4 #(
		.INIT('h1555)
	) name180 (
		_w1313_,
		_w1338_,
		_w1343_,
		_w1360_,
		_w1361_
	);
	LUT2 #(
		.INIT('h2)
	) name181 (
		\g1088_reg/NET0131 ,
		\g2389_reg/NET0131 ,
		_w1362_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name182 (
		\g1092_reg/NET0131 ,
		\g2387_reg/NET0131 ,
		\g2388_reg/NET0131 ,
		\g7961_pad ,
		_w1363_
	);
	LUT2 #(
		.INIT('h4)
	) name183 (
		_w1362_,
		_w1363_,
		_w1364_
	);
	LUT3 #(
		.INIT('h8a)
	) name184 (
		\g1563_reg/NET0131 ,
		_w1362_,
		_w1363_,
		_w1365_
	);
	LUT2 #(
		.INIT('h2)
	) name185 (
		\g1092_reg/NET0131 ,
		\g2391_reg/NET0131 ,
		_w1366_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name186 (
		\g1088_reg/NET0131 ,
		\g2390_reg/NET0131 ,
		\g2392_reg/NET0131 ,
		\g7961_pad ,
		_w1367_
	);
	LUT2 #(
		.INIT('h4)
	) name187 (
		_w1366_,
		_w1367_,
		_w1368_
	);
	LUT4 #(
		.INIT('h0400)
	) name188 (
		_w1251_,
		_w1252_,
		_w1362_,
		_w1363_,
		_w1369_
	);
	LUT2 #(
		.INIT('h8)
	) name189 (
		_w1368_,
		_w1369_,
		_w1370_
	);
	LUT2 #(
		.INIT('h2)
	) name190 (
		\g1088_reg/NET0131 ,
		\g2477_reg/NET0131 ,
		_w1371_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name191 (
		\g1092_reg/NET0131 ,
		\g2478_reg/NET0131 ,
		\g2479_reg/NET0131 ,
		\g7961_pad ,
		_w1372_
	);
	LUT2 #(
		.INIT('h4)
	) name192 (
		_w1371_,
		_w1372_,
		_w1373_
	);
	LUT4 #(
		.INIT('h0080)
	) name193 (
		_w1348_,
		_w1351_,
		_w1355_,
		_w1373_,
		_w1374_
	);
	LUT3 #(
		.INIT('h80)
	) name194 (
		_w1326_,
		_w1337_,
		_w1374_,
		_w1375_
	);
	LUT4 #(
		.INIT('h070f)
	) name195 (
		_w1326_,
		_w1337_,
		_w1370_,
		_w1374_,
		_w1376_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name196 (
		_w1251_,
		_w1252_,
		_w1356_,
		_w1357_,
		_w1377_
	);
	LUT3 #(
		.INIT('h20)
	) name197 (
		_w1355_,
		_w1364_,
		_w1377_,
		_w1378_
	);
	LUT4 #(
		.INIT('h8000)
	) name198 (
		_w1326_,
		_w1337_,
		_w1352_,
		_w1378_,
		_w1379_
	);
	LUT3 #(
		.INIT('h08)
	) name199 (
		_w1368_,
		_w1376_,
		_w1379_,
		_w1380_
	);
	LUT4 #(
		.INIT('h4f00)
	) name200 (
		_w1310_,
		_w1361_,
		_w1365_,
		_w1380_,
		_w1381_
	);
	LUT2 #(
		.INIT('h2)
	) name201 (
		_w1343_,
		_w1345_,
		_w1382_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name202 (
		_w1253_,
		_w1287_,
		_w1299_,
		_w1308_,
		_w1383_
	);
	LUT3 #(
		.INIT('h40)
	) name203 (
		_w1279_,
		_w1282_,
		_w1383_,
		_w1384_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name204 (
		_w1362_,
		_w1363_,
		_w1366_,
		_w1367_,
		_w1385_
	);
	LUT2 #(
		.INIT('h8)
	) name205 (
		_w1333_,
		_w1385_,
		_w1386_
	);
	LUT4 #(
		.INIT('h7f00)
	) name206 (
		_w1326_,
		_w1337_,
		_w1374_,
		_w1386_,
		_w1387_
	);
	LUT4 #(
		.INIT('h5100)
	) name207 (
		_w1370_,
		_w1382_,
		_w1384_,
		_w1387_,
		_w1388_
	);
	LUT4 #(
		.INIT('heee2)
	) name208 (
		\g2390_reg/NET0131 ,
		\g7961_pad ,
		_w1381_,
		_w1388_,
		_w1389_
	);
	LUT4 #(
		.INIT('h0100)
	) name209 (
		\g2991_reg/NET0131 ,
		\g2992_reg/NET0131 ,
		\g3114_reg/NET0131 ,
		\g3120_reg/NET0131 ,
		_w1390_
	);
	LUT2 #(
		.INIT('h1)
	) name210 (
		\g2984_reg/NET0131 ,
		\g2985_reg/NET0131 ,
		_w1391_
	);
	LUT3 #(
		.INIT('h0e)
	) name211 (
		\g2984_reg/NET0131 ,
		\g2985_reg/NET0131 ,
		\g3120_reg/NET0131 ,
		_w1392_
	);
	LUT2 #(
		.INIT('h4)
	) name212 (
		\g3114_reg/NET0131 ,
		\g3139_reg/NET0131 ,
		_w1393_
	);
	LUT4 #(
		.INIT('h4ccc)
	) name213 (
		\g3097_reg/NET0131 ,
		\g3114_reg/NET0131 ,
		\g3120_reg/NET0131 ,
		\g3139_reg/NET0131 ,
		_w1394_
	);
	LUT4 #(
		.INIT('h0045)
	) name214 (
		_w1390_,
		_w1392_,
		_w1393_,
		_w1394_,
		_w1395_
	);
	LUT2 #(
		.INIT('h4)
	) name215 (
		\g3230_pad ,
		\g3233_pad ,
		_w1396_
	);
	LUT2 #(
		.INIT('hb)
	) name216 (
		\g3230_pad ,
		\g3233_pad ,
		_w1397_
	);
	LUT4 #(
		.INIT('h0001)
	) name217 (
		\g3110_reg/NET0131 ,
		\g3114_reg/NET0131 ,
		\g3120_reg/NET0131 ,
		\g3139_reg/NET0131 ,
		_w1398_
	);
	LUT2 #(
		.INIT('h2)
	) name218 (
		_w1396_,
		_w1398_,
		_w1399_
	);
	LUT2 #(
		.INIT('hd)
	) name219 (
		_w1396_,
		_w1398_,
		_w1400_
	);
	LUT3 #(
		.INIT('h01)
	) name220 (
		\g3110_reg/NET0131 ,
		\g3120_reg/NET0131 ,
		\g3139_reg/NET0131 ,
		_w1401_
	);
	LUT3 #(
		.INIT('h01)
	) name221 (
		\g2991_reg/NET0131 ,
		\g2992_reg/NET0131 ,
		\g3114_reg/NET0131 ,
		_w1402_
	);
	LUT3 #(
		.INIT('h5d)
	) name222 (
		_w1396_,
		_w1401_,
		_w1402_,
		_w1403_
	);
	LUT3 #(
		.INIT('h96)
	) name223 (
		\g8260_pad ,
		\g8263_pad ,
		\g8266_pad ,
		_w1404_
	);
	LUT3 #(
		.INIT('h69)
	) name224 (
		\g8259_pad ,
		\g8261_pad ,
		\g8265_pad ,
		_w1405_
	);
	LUT2 #(
		.INIT('h9)
	) name225 (
		\g8262_pad ,
		\g8264_pad ,
		_w1406_
	);
	LUT4 #(
		.INIT('h6996)
	) name226 (
		\g2990_reg/NET0131 ,
		_w1404_,
		_w1405_,
		_w1406_,
		_w1407_
	);
	LUT2 #(
		.INIT('h2)
	) name227 (
		\g3120_reg/NET0131 ,
		\g3231_pad ,
		_w1408_
	);
	LUT4 #(
		.INIT('h6996)
	) name228 (
		_w1404_,
		_w1405_,
		_w1406_,
		_w1408_,
		_w1409_
	);
	LUT3 #(
		.INIT('hd8)
	) name229 (
		\g2987_reg/NET0131 ,
		\g2997_reg/NET0131 ,
		\g3061_reg/NET0131 ,
		_w1410_
	);
	LUT3 #(
		.INIT('h96)
	) name230 (
		\g8270_pad ,
		\g8271_pad ,
		\g8273_pad ,
		_w1411_
	);
	LUT3 #(
		.INIT('h69)
	) name231 (
		\g8268_pad ,
		\g8269_pad ,
		\g8272_pad ,
		_w1412_
	);
	LUT2 #(
		.INIT('h9)
	) name232 (
		\g8274_pad ,
		\g8275_pad ,
		_w1413_
	);
	LUT4 #(
		.INIT('h6996)
	) name233 (
		\g3083_reg/NET0131 ,
		_w1411_,
		_w1412_,
		_w1413_,
		_w1414_
	);
	LUT4 #(
		.INIT('h6996)
	) name234 (
		_w1408_,
		_w1411_,
		_w1412_,
		_w1413_,
		_w1415_
	);
	LUT4 #(
		.INIT('h0002)
	) name235 (
		\g2574_reg/NET0131 ,
		\g2618_reg/NET0131 ,
		\g2633_reg/NET0131 ,
		\g2637_pad ,
		_w1416_
	);
	LUT2 #(
		.INIT('h8)
	) name236 (
		\g2688_reg/NET0131 ,
		\g5657_pad ,
		_w1417_
	);
	LUT4 #(
		.INIT('h135f)
	) name237 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2691_reg/NET0131 ,
		\g2694_reg/NET0131 ,
		_w1418_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w1417_,
		_w1418_,
		_w1419_
	);
	LUT2 #(
		.INIT('h4)
	) name239 (
		\g2797_reg/NET0131 ,
		\g5657_pad ,
		_w1420_
	);
	LUT4 #(
		.INIT('hf351)
	) name240 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2796_reg/NET0131 ,
		\g2798_reg/NET0131 ,
		_w1421_
	);
	LUT2 #(
		.INIT('h4)
	) name241 (
		_w1420_,
		_w1421_,
		_w1422_
	);
	LUT2 #(
		.INIT('h4)
	) name242 (
		\g2779_reg/NET0131 ,
		\g5657_pad ,
		_w1423_
	);
	LUT4 #(
		.INIT('hf351)
	) name243 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2778_reg/NET0131 ,
		\g2780_reg/NET0131 ,
		_w1424_
	);
	LUT2 #(
		.INIT('h4)
	) name244 (
		_w1423_,
		_w1424_,
		_w1425_
	);
	LUT2 #(
		.INIT('h4)
	) name245 (
		\g2791_reg/NET0131 ,
		\g5657_pad ,
		_w1426_
	);
	LUT4 #(
		.INIT('hf351)
	) name246 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2790_reg/NET0131 ,
		\g2792_reg/NET0131 ,
		_w1427_
	);
	LUT4 #(
		.INIT('h0b00)
	) name247 (
		_w1423_,
		_w1424_,
		_w1426_,
		_w1427_,
		_w1428_
	);
	LUT2 #(
		.INIT('h4)
	) name248 (
		\g2788_reg/NET0131 ,
		\g5657_pad ,
		_w1429_
	);
	LUT4 #(
		.INIT('hf351)
	) name249 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2787_reg/NET0131 ,
		\g2789_reg/NET0131 ,
		_w1430_
	);
	LUT2 #(
		.INIT('h4)
	) name250 (
		\g2785_reg/NET0131 ,
		\g5657_pad ,
		_w1431_
	);
	LUT4 #(
		.INIT('hf351)
	) name251 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2784_reg/NET0131 ,
		\g2786_reg/NET0131 ,
		_w1432_
	);
	LUT4 #(
		.INIT('h0400)
	) name252 (
		_w1429_,
		_w1430_,
		_w1431_,
		_w1432_,
		_w1433_
	);
	LUT2 #(
		.INIT('h4)
	) name253 (
		\g2794_reg/NET0131 ,
		\g5657_pad ,
		_w1434_
	);
	LUT4 #(
		.INIT('hf351)
	) name254 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2793_reg/NET0131 ,
		\g2795_reg/NET0131 ,
		_w1435_
	);
	LUT4 #(
		.INIT('h0b00)
	) name255 (
		_w1420_,
		_w1421_,
		_w1434_,
		_w1435_,
		_w1436_
	);
	LUT2 #(
		.INIT('h4)
	) name256 (
		\g2782_reg/NET0131 ,
		\g5657_pad ,
		_w1437_
	);
	LUT4 #(
		.INIT('hf351)
	) name257 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2781_reg/NET0131 ,
		\g2783_reg/NET0131 ,
		_w1438_
	);
	LUT2 #(
		.INIT('h4)
	) name258 (
		_w1437_,
		_w1438_,
		_w1439_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		\g2773_reg/NET0131 ,
		\g5657_pad ,
		_w1440_
	);
	LUT4 #(
		.INIT('hf351)
	) name260 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2772_reg/NET0131 ,
		\g2774_reg/NET0131 ,
		_w1441_
	);
	LUT4 #(
		.INIT('h0b00)
	) name261 (
		_w1437_,
		_w1438_,
		_w1440_,
		_w1441_,
		_w1442_
	);
	LUT4 #(
		.INIT('h8000)
	) name262 (
		_w1428_,
		_w1433_,
		_w1436_,
		_w1442_,
		_w1443_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		\g1018_reg/NET0131 ,
		\g2813_reg/NET0131 ,
		_w1444_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name264 (
		\g1024_reg/NET0131 ,
		\g2811_reg/NET0131 ,
		\g2812_reg/NET0131 ,
		\g5657_pad ,
		_w1445_
	);
	LUT2 #(
		.INIT('h2)
	) name265 (
		\g1024_reg/NET0131 ,
		\g2805_reg/NET0131 ,
		_w1446_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name266 (
		\g1018_reg/NET0131 ,
		\g2806_reg/NET0131 ,
		\g2807_reg/NET0131 ,
		\g5657_pad ,
		_w1447_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name267 (
		_w1444_,
		_w1445_,
		_w1446_,
		_w1447_,
		_w1448_
	);
	LUT2 #(
		.INIT('h4)
	) name268 (
		\g2776_reg/NET0131 ,
		\g5657_pad ,
		_w1449_
	);
	LUT4 #(
		.INIT('hf351)
	) name269 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2775_reg/NET0131 ,
		\g2777_reg/NET0131 ,
		_w1450_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		\g2800_reg/NET0131 ,
		\g5657_pad ,
		_w1451_
	);
	LUT4 #(
		.INIT('hf351)
	) name271 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2799_reg/NET0131 ,
		\g2801_reg/NET0131 ,
		_w1452_
	);
	LUT2 #(
		.INIT('h4)
	) name272 (
		_w1451_,
		_w1452_,
		_w1453_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name273 (
		_w1449_,
		_w1450_,
		_w1451_,
		_w1452_,
		_w1454_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		_w1448_,
		_w1454_,
		_w1455_
	);
	LUT4 #(
		.INIT('ha999)
	) name275 (
		_w1419_,
		_w1422_,
		_w1443_,
		_w1455_,
		_w1456_
	);
	LUT2 #(
		.INIT('h8)
	) name276 (
		\g2679_reg/NET0131 ,
		\g5657_pad ,
		_w1457_
	);
	LUT4 #(
		.INIT('h135f)
	) name277 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2682_reg/NET0131 ,
		\g2685_reg/NET0131 ,
		_w1458_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		_w1457_,
		_w1458_,
		_w1459_
	);
	LUT3 #(
		.INIT('h08)
	) name279 (
		_w1448_,
		_w1454_,
		_w1459_,
		_w1460_
	);
	LUT4 #(
		.INIT('h4044)
	) name280 (
		_w1451_,
		_w1452_,
		_w1457_,
		_w1458_,
		_w1461_
	);
	LUT4 #(
		.INIT('h0b00)
	) name281 (
		_w1451_,
		_w1452_,
		_w1457_,
		_w1458_,
		_w1462_
	);
	LUT3 #(
		.INIT('h70)
	) name282 (
		_w1443_,
		_w1455_,
		_w1462_,
		_w1463_
	);
	LUT4 #(
		.INIT('hec13)
	) name283 (
		_w1443_,
		_w1453_,
		_w1455_,
		_w1459_,
		_w1464_
	);
	LUT3 #(
		.INIT('h80)
	) name284 (
		_w1416_,
		_w1456_,
		_w1464_,
		_w1465_
	);
	LUT2 #(
		.INIT('h8)
	) name285 (
		\g1243_reg/NET0131 ,
		_w1416_,
		_w1466_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w1461_,
		_w1466_,
		_w1467_
	);
	LUT3 #(
		.INIT('h70)
	) name287 (
		_w1443_,
		_w1460_,
		_w1467_,
		_w1468_
	);
	LUT4 #(
		.INIT('h4c5f)
	) name288 (
		_w1456_,
		_w1463_,
		_w1466_,
		_w1468_,
		_w1469_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w1465_,
		_w1469_,
		_w1470_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name290 (
		_w1417_,
		_w1418_,
		_w1423_,
		_w1424_,
		_w1471_
	);
	LUT3 #(
		.INIT('h70)
	) name291 (
		_w1443_,
		_w1455_,
		_w1471_,
		_w1472_
	);
	LUT4 #(
		.INIT('h0400)
	) name292 (
		_w1417_,
		_w1418_,
		_w1423_,
		_w1424_,
		_w1473_
	);
	LUT3 #(
		.INIT('h80)
	) name293 (
		_w1419_,
		_w1448_,
		_w1454_,
		_w1474_
	);
	LUT4 #(
		.INIT('h5666)
	) name294 (
		_w1419_,
		_w1425_,
		_w1443_,
		_w1455_,
		_w1475_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name295 (
		_w1437_,
		_w1438_,
		_w1457_,
		_w1458_,
		_w1476_
	);
	LUT3 #(
		.INIT('h70)
	) name296 (
		_w1443_,
		_w1455_,
		_w1476_,
		_w1477_
	);
	LUT4 #(
		.INIT('h0400)
	) name297 (
		_w1437_,
		_w1438_,
		_w1457_,
		_w1458_,
		_w1478_
	);
	LUT3 #(
		.INIT('h80)
	) name298 (
		_w1448_,
		_w1454_,
		_w1459_,
		_w1479_
	);
	LUT4 #(
		.INIT('h15ea)
	) name299 (
		_w1439_,
		_w1443_,
		_w1455_,
		_w1459_,
		_w1480_
	);
	LUT3 #(
		.INIT('hd7)
	) name300 (
		_w1416_,
		_w1475_,
		_w1480_,
		_w1481_
	);
	LUT4 #(
		.INIT('h4b44)
	) name301 (
		_w1417_,
		_w1418_,
		_w1440_,
		_w1441_,
		_w1482_
	);
	LUT2 #(
		.INIT('h2)
	) name302 (
		_w1416_,
		_w1482_,
		_w1483_
	);
	LUT4 #(
		.INIT('h00d7)
	) name303 (
		_w1416_,
		_w1475_,
		_w1480_,
		_w1483_,
		_w1484_
	);
	LUT3 #(
		.INIT('h02)
	) name304 (
		_w1416_,
		_w1473_,
		_w1482_,
		_w1485_
	);
	LUT3 #(
		.INIT('h70)
	) name305 (
		_w1443_,
		_w1474_,
		_w1485_,
		_w1486_
	);
	LUT4 #(
		.INIT('h0200)
	) name306 (
		_w1416_,
		_w1472_,
		_w1480_,
		_w1486_,
		_w1487_
	);
	LUT3 #(
		.INIT('h02)
	) name307 (
		_w1416_,
		_w1478_,
		_w1482_,
		_w1488_
	);
	LUT3 #(
		.INIT('h70)
	) name308 (
		_w1443_,
		_w1479_,
		_w1488_,
		_w1489_
	);
	LUT3 #(
		.INIT('h10)
	) name309 (
		_w1475_,
		_w1477_,
		_w1489_,
		_w1490_
	);
	LUT4 #(
		.INIT('h4044)
	) name310 (
		_w1449_,
		_w1450_,
		_w1457_,
		_w1458_,
		_w1491_
	);
	LUT4 #(
		.INIT('hb4bb)
	) name311 (
		_w1449_,
		_w1450_,
		_w1457_,
		_w1458_,
		_w1492_
	);
	LUT3 #(
		.INIT('h08)
	) name312 (
		_w1448_,
		_w1454_,
		_w1491_,
		_w1493_
	);
	LUT3 #(
		.INIT('h13)
	) name313 (
		_w1443_,
		_w1492_,
		_w1493_,
		_w1494_
	);
	LUT3 #(
		.INIT('h2a)
	) name314 (
		_w1416_,
		_w1443_,
		_w1460_,
		_w1495_
	);
	LUT2 #(
		.INIT('h4)
	) name315 (
		_w1494_,
		_w1495_,
		_w1496_
	);
	LUT4 #(
		.INIT('h0100)
	) name316 (
		_w1484_,
		_w1487_,
		_w1490_,
		_w1496_,
		_w1497_
	);
	LUT3 #(
		.INIT('hf9)
	) name317 (
		_w1481_,
		_w1483_,
		_w1496_,
		_w1498_
	);
	LUT4 #(
		.INIT('h4b44)
	) name318 (
		_w1434_,
		_w1435_,
		_w1457_,
		_w1458_,
		_w1499_
	);
	LUT4 #(
		.INIT('h4b44)
	) name319 (
		_w1417_,
		_w1418_,
		_w1431_,
		_w1432_,
		_w1500_
	);
	LUT4 #(
		.INIT('h4b44)
	) name320 (
		_w1429_,
		_w1430_,
		_w1457_,
		_w1458_,
		_w1501_
	);
	LUT4 #(
		.INIT('hd77d)
	) name321 (
		_w1416_,
		_w1499_,
		_w1500_,
		_w1501_,
		_w1502_
	);
	LUT4 #(
		.INIT('h4b44)
	) name322 (
		_w1417_,
		_w1418_,
		_w1426_,
		_w1427_,
		_w1503_
	);
	LUT2 #(
		.INIT('h8)
	) name323 (
		\g1880_reg/NET0131 ,
		\g1924_reg/NET0131 ,
		_w1504_
	);
	LUT3 #(
		.INIT('h70)
	) name324 (
		\g1880_reg/NET0131 ,
		\g1924_reg/NET0131 ,
		\g5657_pad ,
		_w1505_
	);
	LUT3 #(
		.INIT('h54)
	) name325 (
		\g2574_reg/NET0131 ,
		\g2622_reg/NET0131 ,
		\g5657_pad ,
		_w1506_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w1505_,
		_w1506_,
		_w1507_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		\g1186_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w1508_
	);
	LUT3 #(
		.INIT('h20)
	) name328 (
		\g1186_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		\g5657_pad ,
		_w1509_
	);
	LUT4 #(
		.INIT('h1500)
	) name329 (
		\g1186_reg/NET0131 ,
		\g499_reg/NET0131 ,
		\g544_reg/NET0131 ,
		\g5657_pad ,
		_w1510_
	);
	LUT3 #(
		.INIT('h54)
	) name330 (
		\g1880_reg/NET0131 ,
		\g1928_reg/NET0131 ,
		\g5657_pad ,
		_w1511_
	);
	LUT4 #(
		.INIT('h0200)
	) name331 (
		_w1506_,
		_w1509_,
		_w1510_,
		_w1511_,
		_w1512_
	);
	LUT4 #(
		.INIT('h0002)
	) name332 (
		_w1416_,
		_w1503_,
		_w1507_,
		_w1512_,
		_w1513_
	);
	LUT3 #(
		.INIT('h10)
	) name333 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		_w1514_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		\g2612_reg/NET0131 ,
		\g3229_pad ,
		_w1515_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		\g2574_reg/NET0131 ,
		\g2618_reg/NET0131 ,
		_w1516_
	);
	LUT4 #(
		.INIT('h0007)
	) name336 (
		\g2574_reg/NET0131 ,
		\g2618_reg/NET0131 ,
		\g2633_reg/NET0131 ,
		\g2637_pad ,
		_w1517_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\g2615_reg/NET0131 ,
		\g3229_pad ,
		_w1518_
	);
	LUT4 #(
		.INIT('h0020)
	) name338 (
		_w1514_,
		_w1515_,
		_w1517_,
		_w1518_,
		_w1519_
	);
	LUT3 #(
		.INIT('h10)
	) name339 (
		_w1507_,
		_w1512_,
		_w1519_,
		_w1520_
	);
	LUT4 #(
		.INIT('h00d7)
	) name340 (
		\g1196_reg/NET0131 ,
		_w1502_,
		_w1513_,
		_w1520_,
		_w1521_
	);
	LUT4 #(
		.INIT('h007d)
	) name341 (
		\g1196_reg/NET0131 ,
		_w1502_,
		_w1513_,
		_w1520_,
		_w1522_
	);
	LUT4 #(
		.INIT('h04bf)
	) name342 (
		_w1497_,
		_w1498_,
		_w1521_,
		_w1522_,
		_w1523_
	);
	LUT2 #(
		.INIT('he)
	) name343 (
		_w1470_,
		_w1523_,
		_w1524_
	);
	LUT3 #(
		.INIT('he4)
	) name344 (
		\g2987_reg/NET0131 ,
		\g3051_reg/NET0131 ,
		\g3070_reg/NET0131 ,
		_w1525_
	);
	LUT3 #(
		.INIT('he4)
	) name345 (
		\g2987_reg/NET0131 ,
		\g3060_reg/NET0131 ,
		\g3078_reg/NET0131 ,
		_w1526_
	);
	LUT3 #(
		.INIT('he4)
	) name346 (
		\g2987_reg/NET0131 ,
		\g3057_reg/NET0131 ,
		\g3075_reg/NET0131 ,
		_w1527_
	);
	LUT3 #(
		.INIT('he4)
	) name347 (
		\g2987_reg/NET0131 ,
		\g3058_reg/NET0131 ,
		\g3076_reg/NET0131 ,
		_w1528_
	);
	LUT3 #(
		.INIT('he4)
	) name348 (
		\g2987_reg/NET0131 ,
		\g3053_reg/NET0131 ,
		\g3072_reg/NET0131 ,
		_w1529_
	);
	LUT3 #(
		.INIT('he4)
	) name349 (
		\g2987_reg/NET0131 ,
		\g3059_reg/NET0131 ,
		\g3077_reg/NET0131 ,
		_w1530_
	);
	LUT3 #(
		.INIT('he4)
	) name350 (
		\g2987_reg/NET0131 ,
		\g3056_reg/NET0131 ,
		\g3074_reg/NET0131 ,
		_w1531_
	);
	LUT3 #(
		.INIT('he4)
	) name351 (
		\g2987_reg/NET0131 ,
		\g3052_reg/NET0131 ,
		\g3071_reg/NET0131 ,
		_w1532_
	);
	LUT3 #(
		.INIT('he4)
	) name352 (
		\g2987_reg/NET0131 ,
		\g3055_reg/NET0131 ,
		\g3073_reg/NET0131 ,
		_w1533_
	);
	LUT4 #(
		.INIT('h0002)
	) name353 (
		\g1880_reg/NET0131 ,
		\g1924_reg/NET0131 ,
		\g1939_reg/NET0131 ,
		\g1943_pad ,
		_w1534_
	);
	LUT2 #(
		.INIT('h4)
	) name354 (
		\g2100_reg/NET0131 ,
		\g5657_pad ,
		_w1535_
	);
	LUT4 #(
		.INIT('hf351)
	) name355 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2099_reg/NET0131 ,
		\g2101_reg/NET0131 ,
		_w1536_
	);
	LUT2 #(
		.INIT('h2)
	) name356 (
		\g1024_reg/NET0131 ,
		\g2111_reg/NET0131 ,
		_w1537_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name357 (
		\g1018_reg/NET0131 ,
		\g2112_reg/NET0131 ,
		\g2113_reg/NET0131 ,
		\g5657_pad ,
		_w1538_
	);
	LUT4 #(
		.INIT('h4044)
	) name358 (
		_w1535_,
		_w1536_,
		_w1537_,
		_w1538_,
		_w1539_
	);
	LUT2 #(
		.INIT('h4)
	) name359 (
		\g2097_reg/NET0131 ,
		\g5657_pad ,
		_w1540_
	);
	LUT4 #(
		.INIT('hf351)
	) name360 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2096_reg/NET0131 ,
		\g2098_reg/NET0131 ,
		_w1541_
	);
	LUT2 #(
		.INIT('h2)
	) name361 (
		\g1018_reg/NET0131 ,
		\g2119_reg/NET0131 ,
		_w1542_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name362 (
		\g1024_reg/NET0131 ,
		\g2117_reg/NET0131 ,
		\g2118_reg/NET0131 ,
		\g5657_pad ,
		_w1543_
	);
	LUT4 #(
		.INIT('h4044)
	) name363 (
		_w1540_,
		_w1541_,
		_w1542_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h8)
	) name364 (
		_w1539_,
		_w1544_,
		_w1545_
	);
	LUT2 #(
		.INIT('h4)
	) name365 (
		\g2103_reg/NET0131 ,
		\g5657_pad ,
		_w1546_
	);
	LUT4 #(
		.INIT('hf351)
	) name366 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2102_reg/NET0131 ,
		\g2104_reg/NET0131 ,
		_w1547_
	);
	LUT2 #(
		.INIT('h4)
	) name367 (
		_w1546_,
		_w1547_,
		_w1548_
	);
	LUT2 #(
		.INIT('h4)
	) name368 (
		\g2094_reg/NET0131 ,
		\g5657_pad ,
		_w1549_
	);
	LUT4 #(
		.INIT('hf351)
	) name369 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2093_reg/NET0131 ,
		\g2095_reg/NET0131 ,
		_w1550_
	);
	LUT4 #(
		.INIT('h0b00)
	) name370 (
		_w1546_,
		_w1547_,
		_w1549_,
		_w1550_,
		_w1551_
	);
	LUT2 #(
		.INIT('h4)
	) name371 (
		\g2079_reg/NET0131 ,
		\g5657_pad ,
		_w1552_
	);
	LUT4 #(
		.INIT('hf351)
	) name372 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2078_reg/NET0131 ,
		\g2080_reg/NET0131 ,
		_w1553_
	);
	LUT2 #(
		.INIT('h4)
	) name373 (
		\g2091_reg/NET0131 ,
		\g5657_pad ,
		_w1554_
	);
	LUT4 #(
		.INIT('hf351)
	) name374 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2090_reg/NET0131 ,
		\g2092_reg/NET0131 ,
		_w1555_
	);
	LUT4 #(
		.INIT('h0400)
	) name375 (
		_w1552_,
		_w1553_,
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h4)
	) name376 (
		\g2088_reg/NET0131 ,
		\g5657_pad ,
		_w1557_
	);
	LUT4 #(
		.INIT('hf351)
	) name377 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2087_reg/NET0131 ,
		\g2089_reg/NET0131 ,
		_w1558_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		_w1557_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h4)
	) name379 (
		\g2082_reg/NET0131 ,
		\g5657_pad ,
		_w1560_
	);
	LUT4 #(
		.INIT('hf351)
	) name380 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2081_reg/NET0131 ,
		\g2083_reg/NET0131 ,
		_w1561_
	);
	LUT2 #(
		.INIT('h4)
	) name381 (
		_w1560_,
		_w1561_,
		_w1562_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name382 (
		_w1557_,
		_w1558_,
		_w1560_,
		_w1561_,
		_w1563_
	);
	LUT2 #(
		.INIT('h4)
	) name383 (
		\g2085_reg/NET0131 ,
		\g5657_pad ,
		_w1564_
	);
	LUT4 #(
		.INIT('hf351)
	) name384 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2084_reg/NET0131 ,
		\g2086_reg/NET0131 ,
		_w1565_
	);
	LUT2 #(
		.INIT('h4)
	) name385 (
		_w1564_,
		_w1565_,
		_w1566_
	);
	LUT2 #(
		.INIT('h4)
	) name386 (
		\g2106_reg/NET0131 ,
		\g5657_pad ,
		_w1567_
	);
	LUT4 #(
		.INIT('hf351)
	) name387 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2105_reg/NET0131 ,
		\g2107_reg/NET0131 ,
		_w1568_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name389 (
		_w1564_,
		_w1565_,
		_w1567_,
		_w1568_,
		_w1570_
	);
	LUT4 #(
		.INIT('h8000)
	) name390 (
		_w1551_,
		_w1556_,
		_w1563_,
		_w1570_,
		_w1571_
	);
	LUT2 #(
		.INIT('h8)
	) name391 (
		\g1018_reg/NET0131 ,
		\g1988_reg/NET0131 ,
		_w1572_
	);
	LUT4 #(
		.INIT('h135f)
	) name392 (
		\g1024_reg/NET0131 ,
		\g1985_reg/NET0131 ,
		\g1991_reg/NET0131 ,
		\g5657_pad ,
		_w1573_
	);
	LUT2 #(
		.INIT('h4)
	) name393 (
		_w1572_,
		_w1573_,
		_w1574_
	);
	LUT4 #(
		.INIT('hec13)
	) name394 (
		_w1545_,
		_w1559_,
		_w1571_,
		_w1574_,
		_w1575_
	);
	LUT2 #(
		.INIT('h8)
	) name395 (
		\g1024_reg/NET0131 ,
		\g2000_reg/NET0131 ,
		_w1576_
	);
	LUT4 #(
		.INIT('h135f)
	) name396 (
		\g1018_reg/NET0131 ,
		\g1994_reg/NET0131 ,
		\g1997_reg/NET0131 ,
		\g5657_pad ,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name397 (
		_w1576_,
		_w1577_,
		_w1578_
	);
	LUT4 #(
		.INIT('hec13)
	) name398 (
		_w1545_,
		_w1566_,
		_w1571_,
		_w1578_,
		_w1579_
	);
	LUT4 #(
		.INIT('h4b44)
	) name399 (
		_w1552_,
		_w1553_,
		_w1576_,
		_w1577_,
		_w1580_
	);
	LUT4 #(
		.INIT('h2882)
	) name400 (
		_w1534_,
		_w1575_,
		_w1579_,
		_w1580_,
		_w1581_
	);
	LUT4 #(
		.INIT('hec13)
	) name401 (
		_w1545_,
		_w1562_,
		_w1571_,
		_w1574_,
		_w1582_
	);
	LUT4 #(
		.INIT('h4b44)
	) name402 (
		_w1540_,
		_w1541_,
		_w1576_,
		_w1577_,
		_w1583_
	);
	LUT2 #(
		.INIT('h8)
	) name403 (
		_w1534_,
		_w1583_,
		_w1584_
	);
	LUT2 #(
		.INIT('h2)
	) name404 (
		_w1534_,
		_w1583_,
		_w1585_
	);
	LUT4 #(
		.INIT('h4b44)
	) name405 (
		_w1554_,
		_w1555_,
		_w1576_,
		_w1577_,
		_w1586_
	);
	LUT4 #(
		.INIT('h4b44)
	) name406 (
		_w1549_,
		_w1550_,
		_w1572_,
		_w1573_,
		_w1587_
	);
	LUT4 #(
		.INIT('h4b44)
	) name407 (
		_w1535_,
		_w1536_,
		_w1572_,
		_w1573_,
		_w1588_
	);
	LUT4 #(
		.INIT('hd77d)
	) name408 (
		_w1534_,
		_w1586_,
		_w1587_,
		_w1588_,
		_w1589_
	);
	LUT4 #(
		.INIT('h7d82)
	) name409 (
		_w1534_,
		_w1582_,
		_w1583_,
		_w1589_,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name410 (
		_w1581_,
		_w1590_,
		_w1591_
	);
	LUT2 #(
		.INIT('h8)
	) name411 (
		\g1196_reg/NET0131 ,
		_w1589_,
		_w1592_
	);
	LUT4 #(
		.INIT('h2700)
	) name412 (
		_w1582_,
		_w1584_,
		_w1585_,
		_w1592_,
		_w1593_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\g1196_reg/NET0131 ,
		_w1589_,
		_w1594_
	);
	LUT4 #(
		.INIT('hd800)
	) name414 (
		_w1582_,
		_w1584_,
		_w1585_,
		_w1594_,
		_w1595_
	);
	LUT3 #(
		.INIT('ha2)
	) name415 (
		\g1196_reg/NET0131 ,
		_w1534_,
		_w1580_,
		_w1596_
	);
	LUT4 #(
		.INIT('hd700)
	) name416 (
		_w1534_,
		_w1575_,
		_w1579_,
		_w1596_,
		_w1597_
	);
	LUT3 #(
		.INIT('h08)
	) name417 (
		\g1196_reg/NET0131 ,
		_w1534_,
		_w1580_,
		_w1598_
	);
	LUT3 #(
		.INIT('h9f)
	) name418 (
		_w1575_,
		_w1579_,
		_w1598_,
		_w1599_
	);
	LUT4 #(
		.INIT('h0100)
	) name419 (
		_w1593_,
		_w1595_,
		_w1597_,
		_w1599_,
		_w1600_
	);
	LUT4 #(
		.INIT('hec13)
	) name420 (
		_w1545_,
		_w1569_,
		_w1571_,
		_w1574_,
		_w1601_
	);
	LUT4 #(
		.INIT('hec13)
	) name421 (
		_w1545_,
		_w1548_,
		_w1571_,
		_w1578_,
		_w1602_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		\g1243_reg/NET0131 ,
		_w1534_,
		_w1603_
	);
	LUT3 #(
		.INIT('h10)
	) name423 (
		_w1509_,
		_w1510_,
		_w1511_,
		_w1604_
	);
	LUT3 #(
		.INIT('h10)
	) name424 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		_w1605_
	);
	LUT2 #(
		.INIT('h4)
	) name425 (
		\g1918_reg/NET0131 ,
		\g3229_pad ,
		_w1606_
	);
	LUT4 #(
		.INIT('h0007)
	) name426 (
		\g1880_reg/NET0131 ,
		\g1924_reg/NET0131 ,
		\g1939_reg/NET0131 ,
		\g1943_pad ,
		_w1607_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		\g1921_reg/NET0131 ,
		\g3229_pad ,
		_w1608_
	);
	LUT4 #(
		.INIT('h0020)
	) name428 (
		_w1605_,
		_w1606_,
		_w1607_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h4)
	) name429 (
		_w1604_,
		_w1609_,
		_w1610_
	);
	LUT4 #(
		.INIT('h009f)
	) name430 (
		_w1601_,
		_w1602_,
		_w1603_,
		_w1610_,
		_w1611_
	);
	LUT3 #(
		.INIT('h1f)
	) name431 (
		_w1591_,
		_w1600_,
		_w1611_,
		_w1612_
	);
	LUT2 #(
		.INIT('h4)
	) name432 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w1613_
	);
	LUT4 #(
		.INIT('hef00)
	) name433 (
		_w1507_,
		_w1512_,
		_w1517_,
		_w1613_,
		_w1614_
	);
	LUT3 #(
		.INIT('h80)
	) name434 (
		\g2574_reg/NET0131 ,
		_w1448_,
		_w1454_,
		_w1615_
	);
	LUT2 #(
		.INIT('h4)
	) name435 (
		\g2809_reg/NET0131 ,
		\g5657_pad ,
		_w1616_
	);
	LUT4 #(
		.INIT('hf351)
	) name436 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2808_reg/NET0131 ,
		\g2810_reg/NET0131 ,
		_w1617_
	);
	LUT3 #(
		.INIT('h8a)
	) name437 (
		\g2574_reg/NET0131 ,
		_w1616_,
		_w1617_,
		_w1618_
	);
	LUT4 #(
		.INIT('h4c44)
	) name438 (
		\g2574_reg/NET0131 ,
		_w1613_,
		_w1616_,
		_w1617_,
		_w1619_
	);
	LUT4 #(
		.INIT('h2033)
	) name439 (
		_w1443_,
		_w1614_,
		_w1615_,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h2)
	) name440 (
		_w1416_,
		_w1514_,
		_w1621_
	);
	LUT2 #(
		.INIT('h4)
	) name441 (
		_w1499_,
		_w1621_,
		_w1622_
	);
	LUT3 #(
		.INIT('h32)
	) name442 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		_w1623_
	);
	LUT4 #(
		.INIT('h0054)
	) name443 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2603_reg/NET0131 ,
		_w1624_
	);
	LUT2 #(
		.INIT('h8)
	) name444 (
		_w1517_,
		_w1624_,
		_w1625_
	);
	LUT4 #(
		.INIT('he0f0)
	) name445 (
		_w1507_,
		_w1512_,
		_w1623_,
		_w1625_,
		_w1626_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w1622_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('hd)
	) name447 (
		_w1620_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h4)
	) name448 (
		_w1500_,
		_w1621_,
		_w1629_
	);
	LUT4 #(
		.INIT('h0054)
	) name449 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2606_reg/NET0131 ,
		_w1630_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		_w1517_,
		_w1630_,
		_w1631_
	);
	LUT3 #(
		.INIT('h10)
	) name451 (
		_w1507_,
		_w1512_,
		_w1631_,
		_w1632_
	);
	LUT3 #(
		.INIT('h02)
	) name452 (
		_w1623_,
		_w1629_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('hd)
	) name453 (
		_w1620_,
		_w1633_,
		_w1634_
	);
	LUT3 #(
		.INIT('h54)
	) name454 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		_w1635_
	);
	LUT2 #(
		.INIT('h2)
	) name455 (
		_w1416_,
		_w1635_,
		_w1636_
	);
	LUT4 #(
		.INIT('h0054)
	) name456 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2607_reg/NET0131 ,
		_w1637_
	);
	LUT2 #(
		.INIT('h8)
	) name457 (
		_w1517_,
		_w1637_,
		_w1638_
	);
	LUT4 #(
		.INIT('he0f0)
	) name458 (
		_w1507_,
		_w1512_,
		_w1623_,
		_w1638_,
		_w1639_
	);
	LUT4 #(
		.INIT('hefcc)
	) name459 (
		_w1480_,
		_w1614_,
		_w1636_,
		_w1639_,
		_w1640_
	);
	LUT4 #(
		.INIT('h0010)
	) name460 (
		_w1507_,
		_w1512_,
		_w1517_,
		_w1618_,
		_w1641_
	);
	LUT4 #(
		.INIT('h80cc)
	) name461 (
		_w1443_,
		_w1613_,
		_w1615_,
		_w1641_,
		_w1642_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w1501_,
		_w1621_,
		_w1643_
	);
	LUT4 #(
		.INIT('h0054)
	) name463 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2605_reg/NET0131 ,
		_w1644_
	);
	LUT2 #(
		.INIT('h8)
	) name464 (
		_w1517_,
		_w1644_,
		_w1645_
	);
	LUT3 #(
		.INIT('h10)
	) name465 (
		_w1507_,
		_w1512_,
		_w1645_,
		_w1646_
	);
	LUT3 #(
		.INIT('h02)
	) name466 (
		_w1623_,
		_w1643_,
		_w1646_,
		_w1647_
	);
	LUT2 #(
		.INIT('he)
	) name467 (
		_w1642_,
		_w1647_,
		_w1648_
	);
	LUT4 #(
		.INIT('h0054)
	) name468 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2608_reg/NET0131 ,
		_w1649_
	);
	LUT2 #(
		.INIT('h8)
	) name469 (
		_w1517_,
		_w1649_,
		_w1650_
	);
	LUT4 #(
		.INIT('he0f0)
	) name470 (
		_w1507_,
		_w1512_,
		_w1623_,
		_w1650_,
		_w1651_
	);
	LUT4 #(
		.INIT('hefcc)
	) name471 (
		_w1475_,
		_w1614_,
		_w1636_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h4)
	) name472 (
		_w1503_,
		_w1621_,
		_w1653_
	);
	LUT4 #(
		.INIT('h0054)
	) name473 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2604_reg/NET0131 ,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		_w1517_,
		_w1654_,
		_w1655_
	);
	LUT3 #(
		.INIT('h10)
	) name475 (
		_w1507_,
		_w1512_,
		_w1655_,
		_w1656_
	);
	LUT3 #(
		.INIT('h02)
	) name476 (
		_w1623_,
		_w1653_,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('he)
	) name477 (
		_w1642_,
		_w1657_,
		_w1658_
	);
	LUT2 #(
		.INIT('h2)
	) name478 (
		_w1416_,
		_w1461_,
		_w1659_
	);
	LUT3 #(
		.INIT('h70)
	) name479 (
		_w1443_,
		_w1460_,
		_w1659_,
		_w1660_
	);
	LUT3 #(
		.INIT('h8c)
	) name480 (
		_w1463_,
		_w1613_,
		_w1660_,
		_w1661_
	);
	LUT3 #(
		.INIT('h70)
	) name481 (
		_w1443_,
		_w1460_,
		_w1621_,
		_w1662_
	);
	LUT4 #(
		.INIT('h0054)
	) name482 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2610_reg/NET0131 ,
		_w1663_
	);
	LUT2 #(
		.INIT('h8)
	) name483 (
		_w1517_,
		_w1663_,
		_w1664_
	);
	LUT4 #(
		.INIT('he0f0)
	) name484 (
		_w1507_,
		_w1512_,
		_w1623_,
		_w1664_,
		_w1665_
	);
	LUT3 #(
		.INIT('hb0)
	) name485 (
		_w1494_,
		_w1662_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('he)
	) name486 (
		_w1661_,
		_w1666_,
		_w1667_
	);
	LUT2 #(
		.INIT('h4)
	) name487 (
		_w1482_,
		_w1621_,
		_w1668_
	);
	LUT4 #(
		.INIT('h0054)
	) name488 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2611_reg/NET0131 ,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name489 (
		_w1517_,
		_w1669_,
		_w1670_
	);
	LUT3 #(
		.INIT('h10)
	) name490 (
		_w1507_,
		_w1512_,
		_w1670_,
		_w1671_
	);
	LUT4 #(
		.INIT('h5551)
	) name491 (
		_w1613_,
		_w1623_,
		_w1668_,
		_w1671_,
		_w1672_
	);
	LUT4 #(
		.INIT('haaa2)
	) name492 (
		_w1416_,
		_w1623_,
		_w1668_,
		_w1671_,
		_w1673_
	);
	LUT3 #(
		.INIT('h13)
	) name493 (
		_w1456_,
		_w1672_,
		_w1673_,
		_w1674_
	);
	LUT3 #(
		.INIT('he4)
	) name494 (
		\g2987_reg/NET0131 ,
		\g3048_reg/NET0131 ,
		\g3067_reg/NET0131 ,
		_w1675_
	);
	LUT3 #(
		.INIT('he4)
	) name495 (
		\g2987_reg/NET0131 ,
		\g3049_reg/NET0131 ,
		\g3068_reg/NET0131 ,
		_w1676_
	);
	LUT3 #(
		.INIT('he4)
	) name496 (
		\g2987_reg/NET0131 ,
		\g3050_reg/NET0131 ,
		\g3069_reg/NET0131 ,
		_w1677_
	);
	LUT3 #(
		.INIT('he4)
	) name497 (
		\g2987_reg/NET0131 ,
		\g3046_reg/NET0131 ,
		\g3065_reg/NET0131 ,
		_w1678_
	);
	LUT3 #(
		.INIT('he4)
	) name498 (
		\g2987_reg/NET0131 ,
		\g3045_reg/NET0131 ,
		\g3064_reg/NET0131 ,
		_w1679_
	);
	LUT3 #(
		.INIT('he4)
	) name499 (
		\g2987_reg/NET0131 ,
		\g3044_reg/NET0131 ,
		\g3063_reg/NET0131 ,
		_w1680_
	);
	LUT3 #(
		.INIT('he4)
	) name500 (
		\g2987_reg/NET0131 ,
		\g3043_reg/NET0131 ,
		\g3062_reg/NET0131 ,
		_w1681_
	);
	LUT3 #(
		.INIT('he4)
	) name501 (
		\g2987_reg/NET0131 ,
		\g3047_reg/NET0131 ,
		\g3066_reg/NET0131 ,
		_w1682_
	);
	LUT2 #(
		.INIT('h1)
	) name502 (
		\g2373_reg/NET0131 ,
		\g2374_reg/NET0131 ,
		_w1683_
	);
	LUT2 #(
		.INIT('h1)
	) name503 (
		\g1679_reg/NET0131 ,
		\g1680_reg/NET0131 ,
		_w1684_
	);
	LUT3 #(
		.INIT('ha8)
	) name504 (
		\g1092_reg/NET0131 ,
		\g1679_reg/NET0131 ,
		\g1680_reg/NET0131 ,
		_w1685_
	);
	LUT4 #(
		.INIT('h0808)
	) name505 (
		\g1092_reg/NET0131 ,
		\g1679_reg/NET0131 ,
		\g1680_reg/NET0131 ,
		\g1686_reg/NET0131 ,
		_w1686_
	);
	LUT3 #(
		.INIT('ha8)
	) name506 (
		\g1092_reg/NET0131 ,
		\g298_reg/NET0131 ,
		\g299_reg/NET0131 ,
		_w1687_
	);
	LUT3 #(
		.INIT('hc8)
	) name507 (
		\g1092_reg/NET0131 ,
		\g986_reg/NET0131 ,
		\g992_reg/NET0131 ,
		_w1688_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		\g985_reg/NET0131 ,
		\g986_reg/NET0131 ,
		_w1689_
	);
	LUT3 #(
		.INIT('ha8)
	) name509 (
		\g1092_reg/NET0131 ,
		\g985_reg/NET0131 ,
		\g986_reg/NET0131 ,
		_w1690_
	);
	LUT4 #(
		.INIT('h8a00)
	) name510 (
		_w1685_,
		_w1687_,
		_w1688_,
		_w1690_,
		_w1691_
	);
	LUT3 #(
		.INIT('hc8)
	) name511 (
		\g1092_reg/NET0131 ,
		\g2374_reg/NET0131 ,
		\g2380_reg/NET0131 ,
		_w1692_
	);
	LUT4 #(
		.INIT('habaa)
	) name512 (
		_w1683_,
		_w1686_,
		_w1691_,
		_w1692_,
		_w1693_
	);
	LUT2 #(
		.INIT('h2)
	) name513 (
		\g315_reg/NET0131 ,
		\g7961_pad ,
		_w1694_
	);
	LUT2 #(
		.INIT('h4)
	) name514 (
		\g315_reg/NET0131 ,
		\g7961_pad ,
		_w1695_
	);
	LUT4 #(
		.INIT('hf351)
	) name515 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g316_reg/NET0131 ,
		\g317_reg/NET0131 ,
		_w1696_
	);
	LUT2 #(
		.INIT('h4)
	) name516 (
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h2)
	) name517 (
		\g1088_reg/NET0131 ,
		\g314_reg/NET0131 ,
		_w1698_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name518 (
		\g1092_reg/NET0131 ,
		\g312_reg/NET0131 ,
		\g313_reg/NET0131 ,
		\g7961_pad ,
		_w1699_
	);
	LUT2 #(
		.INIT('h4)
	) name519 (
		_w1698_,
		_w1699_,
		_w1700_
	);
	LUT4 #(
		.INIT('h4044)
	) name520 (
		_w1695_,
		_w1696_,
		_w1698_,
		_w1699_,
		_w1701_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name521 (
		\g1092_reg/NET0131 ,
		\g145_reg/NET0131 ,
		\g146_reg/NET0131 ,
		\g7961_pad ,
		_w1702_
	);
	LUT2 #(
		.INIT('h2)
	) name522 (
		\g1088_reg/NET0131 ,
		\g144_reg/NET0131 ,
		_w1703_
	);
	LUT3 #(
		.INIT('ha6)
	) name523 (
		\g109_reg/NET0131 ,
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name524 (
		\g1092_reg/NET0131 ,
		\g157_reg/NET0131 ,
		\g158_reg/NET0131 ,
		\g7961_pad ,
		_w1705_
	);
	LUT2 #(
		.INIT('h2)
	) name525 (
		\g1088_reg/NET0131 ,
		\g156_reg/NET0131 ,
		_w1706_
	);
	LUT3 #(
		.INIT('ha6)
	) name526 (
		\g125_reg/NET0131 ,
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT4 #(
		.INIT('hf531)
	) name527 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g132_reg/NET0131 ,
		\g134_reg/NET0131 ,
		_w1708_
	);
	LUT2 #(
		.INIT('h4)
	) name528 (
		\g133_reg/NET0131 ,
		\g7961_pad ,
		_w1709_
	);
	LUT3 #(
		.INIT('ha6)
	) name529 (
		\g101_reg/NET0131 ,
		_w1708_,
		_w1709_,
		_w1710_
	);
	LUT3 #(
		.INIT('h80)
	) name530 (
		_w1704_,
		_w1707_,
		_w1710_,
		_w1711_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name531 (
		\g1088_reg/NET0131 ,
		\g150_reg/NET0131 ,
		\g151_reg/NET0131 ,
		\g7961_pad ,
		_w1712_
	);
	LUT2 #(
		.INIT('h2)
	) name532 (
		\g1092_reg/NET0131 ,
		\g152_reg/NET0131 ,
		_w1713_
	);
	LUT3 #(
		.INIT('ha6)
	) name533 (
		\g117_reg/NET0131 ,
		_w1712_,
		_w1713_,
		_w1714_
	);
	LUT4 #(
		.INIT('hf531)
	) name534 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g141_reg/NET0131 ,
		\g143_reg/NET0131 ,
		_w1715_
	);
	LUT2 #(
		.INIT('h4)
	) name535 (
		\g142_reg/NET0131 ,
		\g7961_pad ,
		_w1716_
	);
	LUT3 #(
		.INIT('ha6)
	) name536 (
		\g105_reg/NET0131 ,
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT4 #(
		.INIT('hf531)
	) name537 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g147_reg/NET0131 ,
		\g149_reg/NET0131 ,
		_w1718_
	);
	LUT2 #(
		.INIT('h4)
	) name538 (
		\g148_reg/NET0131 ,
		\g7961_pad ,
		_w1719_
	);
	LUT3 #(
		.INIT('ha6)
	) name539 (
		\g113_reg/NET0131 ,
		_w1718_,
		_w1719_,
		_w1720_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name540 (
		\g1088_reg/NET0131 ,
		\g153_reg/NET0131 ,
		\g154_reg/NET0131 ,
		\g7961_pad ,
		_w1721_
	);
	LUT2 #(
		.INIT('h2)
	) name541 (
		\g1092_reg/NET0131 ,
		\g155_reg/NET0131 ,
		_w1722_
	);
	LUT3 #(
		.INIT('ha6)
	) name542 (
		\g121_reg/NET0131 ,
		_w1721_,
		_w1722_,
		_w1723_
	);
	LUT4 #(
		.INIT('h8000)
	) name543 (
		_w1714_,
		_w1717_,
		_w1720_,
		_w1723_,
		_w1724_
	);
	LUT4 #(
		.INIT('hf531)
	) name544 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g129_reg/NET0131 ,
		\g131_reg/NET0131 ,
		_w1725_
	);
	LUT2 #(
		.INIT('h4)
	) name545 (
		\g130_reg/NET0131 ,
		\g7961_pad ,
		_w1726_
	);
	LUT3 #(
		.INIT('ha6)
	) name546 (
		\g97_reg/NET0131 ,
		_w1725_,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h2)
	) name547 (
		\g1088_reg/NET0131 ,
		\g171_reg/NET0131 ,
		_w1728_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name548 (
		\g1092_reg/NET0131 ,
		\g172_reg/NET0131 ,
		\g173_reg/NET0131 ,
		\g7961_pad ,
		_w1729_
	);
	LUT2 #(
		.INIT('h4)
	) name549 (
		_w1728_,
		_w1729_,
		_w1730_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		\g163_reg/NET0131 ,
		\g7961_pad ,
		_w1731_
	);
	LUT4 #(
		.INIT('hf531)
	) name551 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g162_reg/NET0131 ,
		\g164_reg/NET0131 ,
		_w1732_
	);
	LUT4 #(
		.INIT('h4b44)
	) name552 (
		_w1728_,
		_w1729_,
		_w1731_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		\g1088_reg/NET0131 ,
		\g168_reg/NET0131 ,
		_w1734_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name554 (
		\g1092_reg/NET0131 ,
		\g169_reg/NET0131 ,
		\g170_reg/NET0131 ,
		\g7961_pad ,
		_w1735_
	);
	LUT2 #(
		.INIT('h4)
	) name555 (
		_w1734_,
		_w1735_,
		_w1736_
	);
	LUT3 #(
		.INIT('h8a)
	) name556 (
		\g1563_reg/NET0131 ,
		_w1734_,
		_w1735_,
		_w1737_
	);
	LUT2 #(
		.INIT('h2)
	) name557 (
		\g1088_reg/NET0131 ,
		\g174_reg/NET0131 ,
		_w1738_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name558 (
		\g1092_reg/NET0131 ,
		\g175_reg/NET0131 ,
		\g176_reg/NET0131 ,
		\g7961_pad ,
		_w1739_
	);
	LUT2 #(
		.INIT('h4)
	) name559 (
		_w1738_,
		_w1739_,
		_w1740_
	);
	LUT2 #(
		.INIT('h2)
	) name560 (
		\g1092_reg/NET0131 ,
		\g161_reg/NET0131 ,
		_w1741_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name561 (
		\g1088_reg/NET0131 ,
		\g159_reg/NET0131 ,
		\g160_reg/NET0131 ,
		\g7961_pad ,
		_w1742_
	);
	LUT4 #(
		.INIT('h4b44)
	) name562 (
		_w1738_,
		_w1739_,
		_w1741_,
		_w1742_,
		_w1743_
	);
	LUT3 #(
		.INIT('h04)
	) name563 (
		_w1733_,
		_w1737_,
		_w1743_,
		_w1744_
	);
	LUT2 #(
		.INIT('h2)
	) name564 (
		\g1088_reg/NET0131 ,
		\g320_reg/NET0131 ,
		_w1745_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name565 (
		\g1092_reg/NET0131 ,
		\g318_reg/NET0131 ,
		\g319_reg/NET0131 ,
		\g7961_pad ,
		_w1746_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		_w1745_,
		_w1746_,
		_w1747_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		\g1088_reg/NET0131 ,
		\g321_reg/NET0131 ,
		_w1748_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name568 (
		\g1092_reg/NET0131 ,
		\g322_reg/NET0131 ,
		\g323_reg/NET0131 ,
		\g7961_pad ,
		_w1749_
	);
	LUT2 #(
		.INIT('h4)
	) name569 (
		_w1748_,
		_w1749_,
		_w1750_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name570 (
		_w1745_,
		_w1746_,
		_w1748_,
		_w1749_,
		_w1751_
	);
	LUT4 #(
		.INIT('h0400)
	) name571 (
		_w1733_,
		_w1737_,
		_w1743_,
		_w1751_,
		_w1752_
	);
	LUT4 #(
		.INIT('h8000)
	) name572 (
		_w1711_,
		_w1724_,
		_w1727_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h8)
	) name573 (
		_w1701_,
		_w1753_,
		_w1754_
	);
	LUT2 #(
		.INIT('h8)
	) name574 (
		\g267_reg/NET0131 ,
		\g7961_pad ,
		_w1755_
	);
	LUT4 #(
		.INIT('h153f)
	) name575 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g270_reg/NET0131 ,
		\g273_reg/NET0131 ,
		_w1756_
	);
	LUT2 #(
		.INIT('h4)
	) name576 (
		_w1755_,
		_w1756_,
		_w1757_
	);
	LUT4 #(
		.INIT('h4b44)
	) name577 (
		_w1728_,
		_w1729_,
		_w1755_,
		_w1756_,
		_w1758_
	);
	LUT4 #(
		.INIT('h153f)
	) name578 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g261_reg/NET0131 ,
		\g264_reg/NET0131 ,
		_w1759_
	);
	LUT2 #(
		.INIT('h8)
	) name579 (
		\g258_reg/NET0131 ,
		\g7961_pad ,
		_w1760_
	);
	LUT2 #(
		.INIT('h2)
	) name580 (
		_w1759_,
		_w1760_,
		_w1761_
	);
	LUT3 #(
		.INIT('ha6)
	) name581 (
		\g125_reg/NET0131 ,
		_w1759_,
		_w1760_,
		_w1762_
	);
	LUT2 #(
		.INIT('h8)
	) name582 (
		\g222_reg/NET0131 ,
		\g7961_pad ,
		_w1763_
	);
	LUT4 #(
		.INIT('h153f)
	) name583 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g225_reg/NET0131 ,
		\g228_reg/NET0131 ,
		_w1764_
	);
	LUT2 #(
		.INIT('h4)
	) name584 (
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT4 #(
		.INIT('h4b44)
	) name585 (
		_w1738_,
		_w1739_,
		_w1763_,
		_w1764_,
		_w1766_
	);
	LUT4 #(
		.INIT('h135f)
	) name586 (
		\g1088_reg/NET0131 ,
		\g231_reg/NET0131 ,
		\g237_reg/NET0131 ,
		\g7961_pad ,
		_w1767_
	);
	LUT2 #(
		.INIT('h8)
	) name587 (
		\g1092_reg/NET0131 ,
		\g234_reg/NET0131 ,
		_w1768_
	);
	LUT2 #(
		.INIT('h2)
	) name588 (
		_w1767_,
		_w1768_,
		_w1769_
	);
	LUT3 #(
		.INIT('ha6)
	) name589 (
		\g101_reg/NET0131 ,
		_w1767_,
		_w1768_,
		_w1770_
	);
	LUT4 #(
		.INIT('h0400)
	) name590 (
		_w1758_,
		_w1762_,
		_w1766_,
		_w1770_,
		_w1771_
	);
	LUT4 #(
		.INIT('h135f)
	) name591 (
		\g1088_reg/NET0131 ,
		\g249_reg/NET0131 ,
		\g255_reg/NET0131 ,
		\g7961_pad ,
		_w1772_
	);
	LUT2 #(
		.INIT('h8)
	) name592 (
		\g1092_reg/NET0131 ,
		\g252_reg/NET0131 ,
		_w1773_
	);
	LUT2 #(
		.INIT('h2)
	) name593 (
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT3 #(
		.INIT('ha6)
	) name594 (
		\g117_reg/NET0131 ,
		_w1772_,
		_w1773_,
		_w1775_
	);
	LUT4 #(
		.INIT('h153f)
	) name595 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g243_reg/NET0131 ,
		\g246_reg/NET0131 ,
		_w1776_
	);
	LUT2 #(
		.INIT('h8)
	) name596 (
		\g240_reg/NET0131 ,
		\g7961_pad ,
		_w1777_
	);
	LUT2 #(
		.INIT('h2)
	) name597 (
		_w1776_,
		_w1777_,
		_w1778_
	);
	LUT3 #(
		.INIT('ha6)
	) name598 (
		\g109_reg/NET0131 ,
		_w1776_,
		_w1777_,
		_w1779_
	);
	LUT2 #(
		.INIT('h8)
	) name599 (
		_w1775_,
		_w1779_,
		_w1780_
	);
	LUT4 #(
		.INIT('h135f)
	) name600 (
		\g1092_reg/NET0131 ,
		\g186_reg/NET0131 ,
		\g189_reg/NET0131 ,
		\g7961_pad ,
		_w1781_
	);
	LUT2 #(
		.INIT('h8)
	) name601 (
		\g1088_reg/NET0131 ,
		\g192_reg/NET0131 ,
		_w1782_
	);
	LUT2 #(
		.INIT('h2)
	) name602 (
		_w1781_,
		_w1782_,
		_w1783_
	);
	LUT3 #(
		.INIT('ha6)
	) name603 (
		\g97_reg/NET0131 ,
		_w1781_,
		_w1782_,
		_w1784_
	);
	LUT2 #(
		.INIT('h8)
	) name604 (
		\g213_reg/NET0131 ,
		\g7961_pad ,
		_w1785_
	);
	LUT4 #(
		.INIT('h153f)
	) name605 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g216_reg/NET0131 ,
		\g219_reg/NET0131 ,
		_w1786_
	);
	LUT2 #(
		.INIT('h4)
	) name606 (
		_w1785_,
		_w1786_,
		_w1787_
	);
	LUT3 #(
		.INIT('h9a)
	) name607 (
		\g121_reg/NET0131 ,
		_w1785_,
		_w1786_,
		_w1788_
	);
	LUT4 #(
		.INIT('h153f)
	) name608 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g198_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w1789_
	);
	LUT2 #(
		.INIT('h8)
	) name609 (
		\g195_reg/NET0131 ,
		\g7961_pad ,
		_w1790_
	);
	LUT2 #(
		.INIT('h2)
	) name610 (
		_w1789_,
		_w1790_,
		_w1791_
	);
	LUT3 #(
		.INIT('ha6)
	) name611 (
		\g105_reg/NET0131 ,
		_w1789_,
		_w1790_,
		_w1792_
	);
	LUT2 #(
		.INIT('h8)
	) name612 (
		\g1088_reg/NET0131 ,
		\g210_reg/NET0131 ,
		_w1793_
	);
	LUT4 #(
		.INIT('h135f)
	) name613 (
		\g1092_reg/NET0131 ,
		\g204_reg/NET0131 ,
		\g207_reg/NET0131 ,
		\g7961_pad ,
		_w1794_
	);
	LUT2 #(
		.INIT('h4)
	) name614 (
		_w1793_,
		_w1794_,
		_w1795_
	);
	LUT3 #(
		.INIT('h9a)
	) name615 (
		\g113_reg/NET0131 ,
		_w1793_,
		_w1794_,
		_w1796_
	);
	LUT4 #(
		.INIT('h8000)
	) name616 (
		_w1784_,
		_w1788_,
		_w1792_,
		_w1796_,
		_w1797_
	);
	LUT3 #(
		.INIT('h80)
	) name617 (
		_w1771_,
		_w1780_,
		_w1797_,
		_w1798_
	);
	LUT4 #(
		.INIT('hc800)
	) name618 (
		_w1762_,
		_w1770_,
		_w1775_,
		_w1779_,
		_w1799_
	);
	LUT3 #(
		.INIT('h2a)
	) name619 (
		_w1758_,
		_w1762_,
		_w1775_,
		_w1800_
	);
	LUT2 #(
		.INIT('h4)
	) name620 (
		_w1799_,
		_w1800_,
		_w1801_
	);
	LUT4 #(
		.INIT('h0007)
	) name621 (
		_w1762_,
		_w1770_,
		_w1775_,
		_w1779_,
		_w1802_
	);
	LUT3 #(
		.INIT('h0b)
	) name622 (
		_w1758_,
		_w1762_,
		_w1770_,
		_w1803_
	);
	LUT3 #(
		.INIT('h23)
	) name623 (
		_w1780_,
		_w1802_,
		_w1803_,
		_w1804_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name624 (
		_w1747_,
		_w1798_,
		_w1801_,
		_w1804_,
		_w1805_
	);
	LUT4 #(
		.INIT('h2a3f)
	) name625 (
		_w1766_,
		_w1784_,
		_w1788_,
		_w1792_,
		_w1806_
	);
	LUT2 #(
		.INIT('h4)
	) name626 (
		_w1766_,
		_w1788_,
		_w1807_
	);
	LUT3 #(
		.INIT('h15)
	) name627 (
		_w1784_,
		_w1792_,
		_w1796_,
		_w1808_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name628 (
		_w1796_,
		_w1806_,
		_w1807_,
		_w1808_,
		_w1809_
	);
	LUT4 #(
		.INIT('h0004)
	) name629 (
		_w1733_,
		_w1737_,
		_w1743_,
		_w1750_,
		_w1810_
	);
	LUT3 #(
		.INIT('h80)
	) name630 (
		_w1724_,
		_w1727_,
		_w1810_,
		_w1811_
	);
	LUT2 #(
		.INIT('h8)
	) name631 (
		_w1784_,
		_w1792_,
		_w1812_
	);
	LUT3 #(
		.INIT('h2a)
	) name632 (
		_w1766_,
		_w1788_,
		_w1796_,
		_w1813_
	);
	LUT2 #(
		.INIT('h4)
	) name633 (
		_w1812_,
		_w1813_,
		_w1814_
	);
	LUT3 #(
		.INIT('h8a)
	) name634 (
		_w1711_,
		_w1812_,
		_w1813_,
		_w1815_
	);
	LUT4 #(
		.INIT('h1555)
	) name635 (
		_w1736_,
		_w1809_,
		_w1811_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h8)
	) name636 (
		\g1563_reg/NET0131 ,
		_w1701_,
		_w1817_
	);
	LUT4 #(
		.INIT('h1055)
	) name637 (
		_w1754_,
		_w1805_,
		_w1816_,
		_w1817_,
		_w1818_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name638 (
		_w1747_,
		_w1771_,
		_w1780_,
		_w1797_,
		_w1819_
	);
	LUT3 #(
		.INIT('h40)
	) name639 (
		_w1801_,
		_w1804_,
		_w1819_,
		_w1820_
	);
	LUT4 #(
		.INIT('h0400)
	) name640 (
		_w1698_,
		_w1699_,
		_w1745_,
		_w1746_,
		_w1821_
	);
	LUT2 #(
		.INIT('h2)
	) name641 (
		_w1697_,
		_w1821_,
		_w1822_
	);
	LUT3 #(
		.INIT('h0b)
	) name642 (
		_w1812_,
		_w1813_,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h8)
	) name643 (
		_w1809_,
		_w1823_,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		\g315_reg/NET0131 ,
		\g7961_pad ,
		_w1825_
	);
	LUT2 #(
		.INIT('h2)
	) name645 (
		\g1092_reg/NET0131 ,
		\g404_reg/NET0131 ,
		_w1826_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name646 (
		\g1088_reg/NET0131 ,
		\g402_reg/NET0131 ,
		\g403_reg/NET0131 ,
		\g7961_pad ,
		_w1827_
	);
	LUT2 #(
		.INIT('h4)
	) name647 (
		_w1826_,
		_w1827_,
		_w1828_
	);
	LUT4 #(
		.INIT('h0004)
	) name648 (
		_w1733_,
		_w1737_,
		_w1743_,
		_w1828_,
		_w1829_
	);
	LUT4 #(
		.INIT('h8000)
	) name649 (
		_w1711_,
		_w1724_,
		_w1727_,
		_w1829_,
		_w1830_
	);
	LUT4 #(
		.INIT('hcd45)
	) name650 (
		_w1697_,
		_w1700_,
		_w1737_,
		_w1747_,
		_w1831_
	);
	LUT3 #(
		.INIT('h01)
	) name651 (
		_w1825_,
		_w1830_,
		_w1831_,
		_w1832_
	);
	LUT3 #(
		.INIT('hb0)
	) name652 (
		_w1820_,
		_w1824_,
		_w1832_,
		_w1833_
	);
	LUT3 #(
		.INIT('hea)
	) name653 (
		_w1694_,
		_w1818_,
		_w1833_,
		_w1834_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		\g1092_reg/NET0131 ,
		\g316_reg/NET0131 ,
		_w1835_
	);
	LUT2 #(
		.INIT('h1)
	) name655 (
		\g1092_reg/NET0131 ,
		\g316_reg/NET0131 ,
		_w1836_
	);
	LUT3 #(
		.INIT('h01)
	) name656 (
		_w1830_,
		_w1831_,
		_w1836_,
		_w1837_
	);
	LUT3 #(
		.INIT('hb0)
	) name657 (
		_w1820_,
		_w1824_,
		_w1837_,
		_w1838_
	);
	LUT3 #(
		.INIT('hec)
	) name658 (
		_w1818_,
		_w1835_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h4)
	) name659 (
		\g1088_reg/NET0131 ,
		\g317_reg/NET0131 ,
		_w1840_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		\g1088_reg/NET0131 ,
		\g317_reg/NET0131 ,
		_w1841_
	);
	LUT3 #(
		.INIT('h01)
	) name661 (
		_w1830_,
		_w1831_,
		_w1841_,
		_w1842_
	);
	LUT3 #(
		.INIT('hb0)
	) name662 (
		_w1820_,
		_w1824_,
		_w1842_,
		_w1843_
	);
	LUT3 #(
		.INIT('hec)
	) name663 (
		_w1818_,
		_w1840_,
		_w1843_,
		_w1844_
	);
	LUT2 #(
		.INIT('h2)
	) name664 (
		\g1003_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w1845_
	);
	LUT2 #(
		.INIT('h4)
	) name665 (
		\g1003_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w1846_
	);
	LUT4 #(
		.INIT('h8acf)
	) name666 (
		\g1002_reg/NET0131 ,
		\g1004_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		\g7961_pad ,
		_w1847_
	);
	LUT2 #(
		.INIT('h4)
	) name667 (
		_w1846_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h4)
	) name668 (
		\g1007_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w1849_
	);
	LUT4 #(
		.INIT('h8acf)
	) name669 (
		\g1005_reg/NET0131 ,
		\g1006_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		_w1850_
	);
	LUT2 #(
		.INIT('h4)
	) name670 (
		_w1849_,
		_w1850_,
		_w1851_
	);
	LUT4 #(
		.INIT('hf531)
	) name671 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g856_reg/NET0131 ,
		\g858_reg/NET0131 ,
		_w1852_
	);
	LUT2 #(
		.INIT('h2)
	) name672 (
		\g7961_pad ,
		\g857_reg/NET0131 ,
		_w1853_
	);
	LUT3 #(
		.INIT('ha2)
	) name673 (
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		\g857_reg/NET0131 ,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		_w1852_,
		_w1854_,
		_w1855_
	);
	LUT4 #(
		.INIT('h0bbb)
	) name675 (
		_w1849_,
		_w1850_,
		_w1852_,
		_w1854_,
		_w1856_
	);
	LUT2 #(
		.INIT('h4)
	) name676 (
		\g1001_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w1857_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name677 (
		\g1000_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g999_reg/NET0131 ,
		_w1858_
	);
	LUT2 #(
		.INIT('h4)
	) name678 (
		_w1857_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w1856_,
		_w1859_,
		_w1860_
	);
	LUT4 #(
		.INIT('hf351)
	) name680 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g830_reg/NET0131 ,
		\g831_reg/NET0131 ,
		_w1861_
	);
	LUT2 #(
		.INIT('h2)
	) name681 (
		\g1088_reg/NET0131 ,
		\g829_reg/NET0131 ,
		_w1862_
	);
	LUT3 #(
		.INIT('ha6)
	) name682 (
		\g793_reg/NET0131 ,
		_w1861_,
		_w1862_,
		_w1863_
	);
	LUT4 #(
		.INIT('hf531)
	) name683 (
		\g1088_reg/NET0131 ,
		\g7961_pad ,
		\g832_reg/NET0131 ,
		\g833_reg/NET0131 ,
		_w1864_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		\g1092_reg/NET0131 ,
		\g834_reg/NET0131 ,
		_w1865_
	);
	LUT3 #(
		.INIT('ha6)
	) name685 (
		\g797_reg/NET0131 ,
		_w1864_,
		_w1865_,
		_w1866_
	);
	LUT4 #(
		.INIT('hf531)
	) name686 (
		\g1088_reg/NET0131 ,
		\g7961_pad ,
		\g817_reg/NET0131 ,
		\g818_reg/NET0131 ,
		_w1867_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		\g1092_reg/NET0131 ,
		\g819_reg/NET0131 ,
		_w1868_
	);
	LUT3 #(
		.INIT('ha6)
	) name688 (
		\g785_reg/NET0131 ,
		_w1867_,
		_w1868_,
		_w1869_
	);
	LUT4 #(
		.INIT('hf351)
	) name689 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g842_reg/NET0131 ,
		\g843_reg/NET0131 ,
		_w1870_
	);
	LUT2 #(
		.INIT('h2)
	) name690 (
		\g1088_reg/NET0131 ,
		\g841_reg/NET0131 ,
		_w1871_
	);
	LUT3 #(
		.INIT('ha6)
	) name691 (
		\g809_reg/NET0131 ,
		_w1870_,
		_w1871_,
		_w1872_
	);
	LUT4 #(
		.INIT('h8000)
	) name692 (
		_w1863_,
		_w1866_,
		_w1869_,
		_w1872_,
		_w1873_
	);
	LUT2 #(
		.INIT('h2)
	) name693 (
		\g1088_reg/NET0131 ,
		\g859_reg/NET0131 ,
		_w1874_
	);
	LUT4 #(
		.INIT('hf351)
	) name694 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g860_reg/NET0131 ,
		\g861_reg/NET0131 ,
		_w1875_
	);
	LUT2 #(
		.INIT('h4)
	) name695 (
		_w1874_,
		_w1875_,
		_w1876_
	);
	LUT2 #(
		.INIT('h2)
	) name696 (
		\g7961_pad ,
		\g851_reg/NET0131 ,
		_w1877_
	);
	LUT4 #(
		.INIT('hf531)
	) name697 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g850_reg/NET0131 ,
		\g852_reg/NET0131 ,
		_w1878_
	);
	LUT4 #(
		.INIT('h4b44)
	) name698 (
		_w1874_,
		_w1875_,
		_w1877_,
		_w1878_,
		_w1879_
	);
	LUT4 #(
		.INIT('hf531)
	) name699 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g838_reg/NET0131 ,
		\g840_reg/NET0131 ,
		_w1880_
	);
	LUT2 #(
		.INIT('h2)
	) name700 (
		\g7961_pad ,
		\g839_reg/NET0131 ,
		_w1881_
	);
	LUT3 #(
		.INIT('hc4)
	) name701 (
		\g7961_pad ,
		\g805_reg/NET0131 ,
		\g839_reg/NET0131 ,
		_w1882_
	);
	LUT2 #(
		.INIT('h8)
	) name702 (
		_w1880_,
		_w1882_,
		_w1883_
	);
	LUT4 #(
		.INIT('hf351)
	) name703 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g821_reg/NET0131 ,
		\g822_reg/NET0131 ,
		_w1884_
	);
	LUT2 #(
		.INIT('h2)
	) name704 (
		\g1088_reg/NET0131 ,
		\g820_reg/NET0131 ,
		_w1885_
	);
	LUT3 #(
		.INIT('h51)
	) name705 (
		\g789_reg/NET0131 ,
		_w1884_,
		_w1885_,
		_w1886_
	);
	LUT3 #(
		.INIT('h01)
	) name706 (
		_w1879_,
		_w1883_,
		_w1886_,
		_w1887_
	);
	LUT3 #(
		.INIT('hc4)
	) name707 (
		\g1088_reg/NET0131 ,
		\g789_reg/NET0131 ,
		\g820_reg/NET0131 ,
		_w1888_
	);
	LUT2 #(
		.INIT('h8)
	) name708 (
		_w1884_,
		_w1888_,
		_w1889_
	);
	LUT2 #(
		.INIT('h2)
	) name709 (
		_w1852_,
		_w1853_,
		_w1890_
	);
	LUT3 #(
		.INIT('ha2)
	) name710 (
		\g1563_reg/NET0131 ,
		_w1852_,
		_w1853_,
		_w1891_
	);
	LUT3 #(
		.INIT('h51)
	) name711 (
		\g805_reg/NET0131 ,
		_w1880_,
		_w1881_,
		_w1892_
	);
	LUT3 #(
		.INIT('h04)
	) name712 (
		_w1889_,
		_w1891_,
		_w1892_,
		_w1893_
	);
	LUT3 #(
		.INIT('h80)
	) name713 (
		_w1873_,
		_w1887_,
		_w1893_,
		_w1894_
	);
	LUT4 #(
		.INIT('hf351)
	) name714 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g836_reg/NET0131 ,
		\g837_reg/NET0131 ,
		_w1895_
	);
	LUT2 #(
		.INIT('h2)
	) name715 (
		\g1088_reg/NET0131 ,
		\g835_reg/NET0131 ,
		_w1896_
	);
	LUT3 #(
		.INIT('ha6)
	) name716 (
		\g801_reg/NET0131 ,
		_w1895_,
		_w1896_,
		_w1897_
	);
	LUT2 #(
		.INIT('h2)
	) name717 (
		\g1088_reg/NET0131 ,
		\g862_reg/NET0131 ,
		_w1898_
	);
	LUT4 #(
		.INIT('hf351)
	) name718 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g863_reg/NET0131 ,
		\g864_reg/NET0131 ,
		_w1899_
	);
	LUT2 #(
		.INIT('h4)
	) name719 (
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h2)
	) name720 (
		\g7961_pad ,
		\g848_reg/NET0131 ,
		_w1901_
	);
	LUT4 #(
		.INIT('hf531)
	) name721 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g847_reg/NET0131 ,
		\g849_reg/NET0131 ,
		_w1902_
	);
	LUT4 #(
		.INIT('h4b44)
	) name722 (
		_w1898_,
		_w1899_,
		_w1901_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h2)
	) name723 (
		_w1897_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h4)
	) name724 (
		\g1009_reg/NET0131 ,
		\g7961_pad ,
		_w1905_
	);
	LUT4 #(
		.INIT('h8caf)
	) name725 (
		\g1008_reg/NET0131 ,
		\g1010_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w1906_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		_w1905_,
		_w1906_,
		_w1907_
	);
	LUT4 #(
		.INIT('hf531)
	) name727 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g844_reg/NET0131 ,
		\g846_reg/NET0131 ,
		_w1908_
	);
	LUT2 #(
		.INIT('h2)
	) name728 (
		\g7961_pad ,
		\g845_reg/NET0131 ,
		_w1909_
	);
	LUT3 #(
		.INIT('ha6)
	) name729 (
		\g813_reg/NET0131 ,
		_w1908_,
		_w1909_,
		_w1910_
	);
	LUT4 #(
		.INIT('h0200)
	) name730 (
		_w1897_,
		_w1903_,
		_w1907_,
		_w1910_,
		_w1911_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		_w1859_,
		_w1911_,
		_w1912_
	);
	LUT4 #(
		.INIT('ha888)
	) name732 (
		_w1848_,
		_w1860_,
		_w1894_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h4)
	) name733 (
		\g1090_reg/NET0131 ,
		\g7961_pad ,
		_w1914_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name734 (
		\g1088_reg/NET0131 ,
		\g1089_reg/NET0131 ,
		\g1091_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w1915_
	);
	LUT2 #(
		.INIT('h4)
	) name735 (
		_w1914_,
		_w1915_,
		_w1916_
	);
	LUT4 #(
		.INIT('h0020)
	) name736 (
		_w1897_,
		_w1903_,
		_w1910_,
		_w1916_,
		_w1917_
	);
	LUT4 #(
		.INIT('h8000)
	) name737 (
		_w1873_,
		_w1887_,
		_w1893_,
		_w1917_,
		_w1918_
	);
	LUT4 #(
		.INIT('h0400)
	) name738 (
		_w1849_,
		_w1850_,
		_w1857_,
		_w1858_,
		_w1919_
	);
	LUT2 #(
		.INIT('h8)
	) name739 (
		_w1848_,
		_w1919_,
		_w1920_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		_w1918_,
		_w1920_,
		_w1921_
	);
	LUT2 #(
		.INIT('h4)
	) name741 (
		_w1913_,
		_w1921_,
		_w1922_
	);
	LUT2 #(
		.INIT('h8)
	) name742 (
		\g1088_reg/NET0131 ,
		\g897_reg/NET0131 ,
		_w1923_
	);
	LUT4 #(
		.INIT('h153f)
	) name743 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g891_reg/NET0131 ,
		\g894_reg/NET0131 ,
		_w1924_
	);
	LUT2 #(
		.INIT('h4)
	) name744 (
		_w1923_,
		_w1924_,
		_w1925_
	);
	LUT3 #(
		.INIT('h9a)
	) name745 (
		\g801_reg/NET0131 ,
		_w1923_,
		_w1924_,
		_w1926_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		\g7961_pad ,
		\g909_reg/NET0131 ,
		_w1927_
	);
	LUT4 #(
		.INIT('h153f)
	) name747 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g912_reg/NET0131 ,
		\g915_reg/NET0131 ,
		_w1928_
	);
	LUT2 #(
		.INIT('h4)
	) name748 (
		_w1927_,
		_w1928_,
		_w1929_
	);
	LUT4 #(
		.INIT('h4b44)
	) name749 (
		_w1898_,
		_w1899_,
		_w1927_,
		_w1928_,
		_w1930_
	);
	LUT2 #(
		.INIT('h8)
	) name750 (
		\g7961_pad ,
		\g882_reg/NET0131 ,
		_w1931_
	);
	LUT4 #(
		.INIT('h153f)
	) name751 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g885_reg/NET0131 ,
		\g888_reg/NET0131 ,
		_w1932_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		_w1931_,
		_w1932_,
		_w1933_
	);
	LUT3 #(
		.INIT('h9a)
	) name753 (
		\g793_reg/NET0131 ,
		_w1931_,
		_w1932_,
		_w1934_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		\g7961_pad ,
		\g900_reg/NET0131 ,
		_w1935_
	);
	LUT4 #(
		.INIT('h153f)
	) name755 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g903_reg/NET0131 ,
		\g906_reg/NET0131 ,
		_w1936_
	);
	LUT2 #(
		.INIT('h4)
	) name756 (
		_w1935_,
		_w1936_,
		_w1937_
	);
	LUT3 #(
		.INIT('h9a)
	) name757 (
		\g809_reg/NET0131 ,
		_w1935_,
		_w1936_,
		_w1938_
	);
	LUT4 #(
		.INIT('h3200)
	) name758 (
		_w1926_,
		_w1930_,
		_w1934_,
		_w1938_,
		_w1939_
	);
	LUT4 #(
		.INIT('h153f)
	) name759 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g873_reg/NET0131 ,
		\g876_reg/NET0131 ,
		_w1940_
	);
	LUT2 #(
		.INIT('h8)
	) name760 (
		\g1088_reg/NET0131 ,
		\g879_reg/NET0131 ,
		_w1941_
	);
	LUT2 #(
		.INIT('h2)
	) name761 (
		_w1940_,
		_w1941_,
		_w1942_
	);
	LUT3 #(
		.INIT('ha6)
	) name762 (
		\g785_reg/NET0131 ,
		_w1940_,
		_w1941_,
		_w1943_
	);
	LUT3 #(
		.INIT('h07)
	) name763 (
		_w1926_,
		_w1934_,
		_w1943_,
		_w1944_
	);
	LUT2 #(
		.INIT('h4)
	) name764 (
		_w1939_,
		_w1944_,
		_w1945_
	);
	LUT4 #(
		.INIT('h0045)
	) name765 (
		_w1926_,
		_w1930_,
		_w1934_,
		_w1938_,
		_w1946_
	);
	LUT2 #(
		.INIT('h8)
	) name766 (
		_w1926_,
		_w1938_,
		_w1947_
	);
	LUT4 #(
		.INIT('h135f)
	) name767 (
		_w1926_,
		_w1934_,
		_w1938_,
		_w1943_,
		_w1948_
	);
	LUT3 #(
		.INIT('h13)
	) name768 (
		_w1930_,
		_w1946_,
		_w1948_,
		_w1949_
	);
	LUT3 #(
		.INIT('h8a)
	) name769 (
		_w1891_,
		_w1945_,
		_w1949_,
		_w1950_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		\g1563_reg/NET0131 ,
		_w1911_,
		_w1951_
	);
	LUT2 #(
		.INIT('h8)
	) name771 (
		_w1894_,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h8)
	) name772 (
		\g7961_pad ,
		\g927_reg/NET0131 ,
		_w1953_
	);
	LUT4 #(
		.INIT('h153f)
	) name773 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g930_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w1954_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		_w1953_,
		_w1954_,
		_w1955_
	);
	LUT3 #(
		.INIT('h9a)
	) name775 (
		\g797_reg/NET0131 ,
		_w1953_,
		_w1954_,
		_w1956_
	);
	LUT2 #(
		.INIT('h8)
	) name776 (
		\g7961_pad ,
		\g954_reg/NET0131 ,
		_w1957_
	);
	LUT4 #(
		.INIT('h153f)
	) name777 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g957_reg/NET0131 ,
		\g960_reg/NET0131 ,
		_w1958_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		_w1957_,
		_w1958_,
		_w1959_
	);
	LUT4 #(
		.INIT('h4b44)
	) name779 (
		_w1874_,
		_w1875_,
		_w1957_,
		_w1958_,
		_w1960_
	);
	LUT2 #(
		.INIT('h8)
	) name780 (
		\g7961_pad ,
		\g918_reg/NET0131 ,
		_w1961_
	);
	LUT4 #(
		.INIT('h153f)
	) name781 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g921_reg/NET0131 ,
		\g924_reg/NET0131 ,
		_w1962_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w1961_,
		_w1962_,
		_w1963_
	);
	LUT3 #(
		.INIT('h9a)
	) name783 (
		\g789_reg/NET0131 ,
		_w1961_,
		_w1962_,
		_w1964_
	);
	LUT2 #(
		.INIT('h8)
	) name784 (
		\g1092_reg/NET0131 ,
		\g948_reg/NET0131 ,
		_w1965_
	);
	LUT4 #(
		.INIT('h153f)
	) name785 (
		\g1088_reg/NET0131 ,
		\g7961_pad ,
		\g945_reg/NET0131 ,
		\g951_reg/NET0131 ,
		_w1966_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		_w1965_,
		_w1966_,
		_w1967_
	);
	LUT3 #(
		.INIT('h9a)
	) name787 (
		\g813_reg/NET0131 ,
		_w1965_,
		_w1966_,
		_w1968_
	);
	LUT4 #(
		.INIT('h4ddd)
	) name788 (
		_w1956_,
		_w1960_,
		_w1964_,
		_w1968_,
		_w1969_
	);
	LUT2 #(
		.INIT('h8)
	) name789 (
		\g1088_reg/NET0131 ,
		\g942_reg/NET0131 ,
		_w1970_
	);
	LUT4 #(
		.INIT('h153f)
	) name790 (
		\g1092_reg/NET0131 ,
		\g7961_pad ,
		\g936_reg/NET0131 ,
		\g939_reg/NET0131 ,
		_w1971_
	);
	LUT2 #(
		.INIT('h4)
	) name791 (
		_w1970_,
		_w1971_,
		_w1972_
	);
	LUT3 #(
		.INIT('h9a)
	) name792 (
		\g805_reg/NET0131 ,
		_w1970_,
		_w1971_,
		_w1973_
	);
	LUT4 #(
		.INIT('h004c)
	) name793 (
		_w1956_,
		_w1960_,
		_w1964_,
		_w1968_,
		_w1974_
	);
	LUT4 #(
		.INIT('h8808)
	) name794 (
		_w1891_,
		_w1969_,
		_w1973_,
		_w1974_,
		_w1975_
	);
	LUT4 #(
		.INIT('h45cf)
	) name795 (
		_w1956_,
		_w1960_,
		_w1968_,
		_w1973_,
		_w1976_
	);
	LUT2 #(
		.INIT('h2)
	) name796 (
		_w1891_,
		_w1964_,
		_w1977_
	);
	LUT2 #(
		.INIT('h8)
	) name797 (
		_w1976_,
		_w1977_,
		_w1978_
	);
	LUT3 #(
		.INIT('h15)
	) name798 (
		_w1920_,
		_w1976_,
		_w1977_,
		_w1979_
	);
	LUT3 #(
		.INIT('h10)
	) name799 (
		_w1918_,
		_w1975_,
		_w1979_,
		_w1980_
	);
	LUT3 #(
		.INIT('h08)
	) name800 (
		\g1563_reg/NET0131 ,
		_w1852_,
		_w1853_,
		_w1981_
	);
	LUT4 #(
		.INIT('h0800)
	) name801 (
		_w1934_,
		_w1943_,
		_w1960_,
		_w1968_,
		_w1982_
	);
	LUT4 #(
		.INIT('h4000)
	) name802 (
		_w1930_,
		_w1956_,
		_w1964_,
		_w1973_,
		_w1983_
	);
	LUT4 #(
		.INIT('h8000)
	) name803 (
		\g1563_reg/NET0131 ,
		_w1947_,
		_w1982_,
		_w1983_,
		_w1984_
	);
	LUT3 #(
		.INIT('h02)
	) name804 (
		_w1851_,
		_w1981_,
		_w1984_,
		_w1985_
	);
	LUT4 #(
		.INIT('hb000)
	) name805 (
		_w1950_,
		_w1952_,
		_w1980_,
		_w1985_,
		_w1986_
	);
	LUT2 #(
		.INIT('h1)
	) name806 (
		\g1003_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w1987_
	);
	LUT4 #(
		.INIT('h1555)
	) name807 (
		_w1859_,
		_w1947_,
		_w1982_,
		_w1983_,
		_w1988_
	);
	LUT3 #(
		.INIT('ha2)
	) name808 (
		_w1969_,
		_w1973_,
		_w1974_,
		_w1989_
	);
	LUT2 #(
		.INIT('h8)
	) name809 (
		_w1851_,
		_w1891_,
		_w1990_
	);
	LUT3 #(
		.INIT('hb0)
	) name810 (
		_w1964_,
		_w1976_,
		_w1990_,
		_w1991_
	);
	LUT3 #(
		.INIT('h20)
	) name811 (
		_w1988_,
		_w1989_,
		_w1991_,
		_w1992_
	);
	LUT2 #(
		.INIT('h4)
	) name812 (
		_w1859_,
		_w1891_,
		_w1993_
	);
	LUT4 #(
		.INIT('h1055)
	) name813 (
		_w1848_,
		_w1945_,
		_w1949_,
		_w1993_,
		_w1994_
	);
	LUT3 #(
		.INIT('h45)
	) name814 (
		_w1987_,
		_w1992_,
		_w1994_,
		_w1995_
	);
	LUT4 #(
		.INIT('hfeaa)
	) name815 (
		_w1845_,
		_w1922_,
		_w1986_,
		_w1995_,
		_w1996_
	);
	LUT4 #(
		.INIT('heee4)
	) name816 (
		\g1092_reg/NET0131 ,
		\g2391_reg/NET0131 ,
		_w1381_,
		_w1388_,
		_w1997_
	);
	LUT4 #(
		.INIT('heee4)
	) name817 (
		\g1088_reg/NET0131 ,
		\g2392_reg/NET0131 ,
		_w1381_,
		_w1388_,
		_w1998_
	);
	LUT2 #(
		.INIT('h2)
	) name818 (
		\g1004_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w1999_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		\g1004_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		_w2000_
	);
	LUT3 #(
		.INIT('h0b)
	) name820 (
		_w1992_,
		_w1994_,
		_w2000_,
		_w2001_
	);
	LUT4 #(
		.INIT('hfef0)
	) name821 (
		_w1922_,
		_w1986_,
		_w1999_,
		_w2001_,
		_w2002_
	);
	LUT2 #(
		.INIT('h2)
	) name822 (
		\g1002_reg/NET0131 ,
		\g7961_pad ,
		_w2003_
	);
	LUT2 #(
		.INIT('h1)
	) name823 (
		\g1002_reg/NET0131 ,
		\g7961_pad ,
		_w2004_
	);
	LUT3 #(
		.INIT('h0b)
	) name824 (
		_w1992_,
		_w1994_,
		_w2004_,
		_w2005_
	);
	LUT4 #(
		.INIT('hfef0)
	) name825 (
		_w1922_,
		_w1986_,
		_w2003_,
		_w2005_,
		_w2006_
	);
	LUT2 #(
		.INIT('h2)
	) name826 (
		\g1088_reg/NET0131 ,
		\g1550_reg/NET0131 ,
		_w2007_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name827 (
		\g1092_reg/NET0131 ,
		\g1551_reg/NET0131 ,
		\g1552_reg/NET0131 ,
		\g7961_pad ,
		_w2008_
	);
	LUT2 #(
		.INIT('h4)
	) name828 (
		_w2007_,
		_w2008_,
		_w2009_
	);
	LUT3 #(
		.INIT('h8a)
	) name829 (
		\g1563_reg/NET0131 ,
		_w2007_,
		_w2008_,
		_w2010_
	);
	LUT2 #(
		.INIT('h2)
	) name830 (
		\g1088_reg/NET0131 ,
		\g1556_reg/NET0131 ,
		_w2011_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name831 (
		\g1092_reg/NET0131 ,
		\g1557_reg/NET0131 ,
		\g1558_reg/NET0131 ,
		\g7961_pad ,
		_w2012_
	);
	LUT2 #(
		.INIT('h4)
	) name832 (
		_w2011_,
		_w2012_,
		_w2013_
	);
	LUT2 #(
		.INIT('h8)
	) name833 (
		\g1603_reg/NET0131 ,
		\g7961_pad ,
		_w2014_
	);
	LUT4 #(
		.INIT('h153f)
	) name834 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1606_reg/NET0131 ,
		\g1609_reg/NET0131 ,
		_w2015_
	);
	LUT2 #(
		.INIT('h4)
	) name835 (
		_w2014_,
		_w2015_,
		_w2016_
	);
	LUT4 #(
		.INIT('h4b44)
	) name836 (
		_w2011_,
		_w2012_,
		_w2014_,
		_w2015_,
		_w2017_
	);
	LUT2 #(
		.INIT('h8)
	) name837 (
		\g1594_reg/NET0131 ,
		\g7961_pad ,
		_w2018_
	);
	LUT4 #(
		.INIT('h153f)
	) name838 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1597_reg/NET0131 ,
		\g1600_reg/NET0131 ,
		_w2019_
	);
	LUT2 #(
		.INIT('h4)
	) name839 (
		_w2018_,
		_w2019_,
		_w2020_
	);
	LUT3 #(
		.INIT('h9a)
	) name840 (
		\g1501_reg/NET0131 ,
		_w2018_,
		_w2019_,
		_w2021_
	);
	LUT2 #(
		.INIT('h8)
	) name841 (
		\g1088_reg/NET0131 ,
		\g1591_reg/NET0131 ,
		_w2022_
	);
	LUT4 #(
		.INIT('h135f)
	) name842 (
		\g1092_reg/NET0131 ,
		\g1585_reg/NET0131 ,
		\g1588_reg/NET0131 ,
		\g7961_pad ,
		_w2023_
	);
	LUT2 #(
		.INIT('h4)
	) name843 (
		_w2022_,
		_w2023_,
		_w2024_
	);
	LUT3 #(
		.INIT('h9a)
	) name844 (
		\g1491_reg/NET0131 ,
		_w2022_,
		_w2023_,
		_w2025_
	);
	LUT4 #(
		.INIT('h135f)
	) name845 (
		\g1088_reg/NET0131 ,
		\g1567_reg/NET0131 ,
		\g1573_reg/NET0131 ,
		\g7961_pad ,
		_w2026_
	);
	LUT2 #(
		.INIT('h8)
	) name846 (
		\g1092_reg/NET0131 ,
		\g1570_reg/NET0131 ,
		_w2027_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w2026_,
		_w2027_,
		_w2028_
	);
	LUT3 #(
		.INIT('ha6)
	) name848 (
		\g1471_reg/NET0131 ,
		_w2026_,
		_w2027_,
		_w2029_
	);
	LUT2 #(
		.INIT('h8)
	) name849 (
		\g1576_reg/NET0131 ,
		\g7961_pad ,
		_w2030_
	);
	LUT4 #(
		.INIT('h153f)
	) name850 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		\g1582_reg/NET0131 ,
		_w2031_
	);
	LUT2 #(
		.INIT('h4)
	) name851 (
		_w2030_,
		_w2031_,
		_w2032_
	);
	LUT3 #(
		.INIT('h9a)
	) name852 (
		\g1481_reg/NET0131 ,
		_w2030_,
		_w2031_,
		_w2033_
	);
	LUT4 #(
		.INIT('h0777)
	) name853 (
		_w2021_,
		_w2025_,
		_w2029_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h8)
	) name854 (
		_w2017_,
		_w2034_,
		_w2035_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w2017_,
		_w2033_,
		_w2036_
	);
	LUT3 #(
		.INIT('h13)
	) name856 (
		_w2021_,
		_w2025_,
		_w2029_,
		_w2037_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w2017_,
		_w2021_,
		_w2038_
	);
	LUT3 #(
		.INIT('h13)
	) name858 (
		_w2025_,
		_w2029_,
		_w2033_,
		_w2039_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name859 (
		_w2036_,
		_w2037_,
		_w2038_,
		_w2039_,
		_w2040_
	);
	LUT3 #(
		.INIT('h8a)
	) name860 (
		_w2010_,
		_w2035_,
		_w2040_,
		_w2041_
	);
	LUT4 #(
		.INIT('hf531)
	) name861 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1529_reg/NET0131 ,
		\g1531_reg/NET0131 ,
		_w2042_
	);
	LUT2 #(
		.INIT('h4)
	) name862 (
		\g1530_reg/NET0131 ,
		\g7961_pad ,
		_w2043_
	);
	LUT3 #(
		.INIT('ha6)
	) name863 (
		\g1491_reg/NET0131 ,
		_w2042_,
		_w2043_,
		_w2044_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name864 (
		\g1088_reg/NET0131 ,
		\g1514_reg/NET0131 ,
		\g1515_reg/NET0131 ,
		\g7961_pad ,
		_w2045_
	);
	LUT2 #(
		.INIT('h2)
	) name865 (
		\g1092_reg/NET0131 ,
		\g1516_reg/NET0131 ,
		_w2046_
	);
	LUT3 #(
		.INIT('ha6)
	) name866 (
		\g1476_reg/NET0131 ,
		_w2045_,
		_w2046_,
		_w2047_
	);
	LUT4 #(
		.INIT('hf531)
	) name867 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1535_reg/NET0131 ,
		\g1537_reg/NET0131 ,
		_w2048_
	);
	LUT2 #(
		.INIT('h4)
	) name868 (
		\g1536_reg/NET0131 ,
		\g7961_pad ,
		_w2049_
	);
	LUT3 #(
		.INIT('ha6)
	) name869 (
		\g1501_reg/NET0131 ,
		_w2048_,
		_w2049_,
		_w2050_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name870 (
		\g1088_reg/NET0131 ,
		\g1538_reg/NET0131 ,
		\g1539_reg/NET0131 ,
		\g7961_pad ,
		_w2051_
	);
	LUT2 #(
		.INIT('h2)
	) name871 (
		\g1092_reg/NET0131 ,
		\g1540_reg/NET0131 ,
		_w2052_
	);
	LUT3 #(
		.INIT('ha6)
	) name872 (
		\g1506_reg/NET0131 ,
		_w2051_,
		_w2052_,
		_w2053_
	);
	LUT4 #(
		.INIT('h8000)
	) name873 (
		_w2044_,
		_w2047_,
		_w2050_,
		_w2053_,
		_w2054_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name874 (
		\g1088_reg/NET0131 ,
		\g1526_reg/NET0131 ,
		\g1527_reg/NET0131 ,
		\g7961_pad ,
		_w2055_
	);
	LUT2 #(
		.INIT('h2)
	) name875 (
		\g1092_reg/NET0131 ,
		\g1528_reg/NET0131 ,
		_w2056_
	);
	LUT3 #(
		.INIT('ha6)
	) name876 (
		\g1486_reg/NET0131 ,
		_w2055_,
		_w2056_,
		_w2057_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name877 (
		\g1088_reg/NET0131 ,
		\g1511_reg/NET0131 ,
		\g1512_reg/NET0131 ,
		\g7961_pad ,
		_w2058_
	);
	LUT2 #(
		.INIT('h2)
	) name878 (
		\g1092_reg/NET0131 ,
		\g1513_reg/NET0131 ,
		_w2059_
	);
	LUT3 #(
		.INIT('ha6)
	) name879 (
		\g1471_reg/NET0131 ,
		_w2058_,
		_w2059_,
		_w2060_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name880 (
		\g1092_reg/NET0131 ,
		\g1524_reg/NET0131 ,
		\g1525_reg/NET0131 ,
		\g7961_pad ,
		_w2061_
	);
	LUT2 #(
		.INIT('h2)
	) name881 (
		\g1088_reg/NET0131 ,
		\g1523_reg/NET0131 ,
		_w2062_
	);
	LUT3 #(
		.INIT('ha6)
	) name882 (
		\g1481_reg/NET0131 ,
		_w2061_,
		_w2062_,
		_w2063_
	);
	LUT4 #(
		.INIT('h8000)
	) name883 (
		_w2010_,
		_w2057_,
		_w2060_,
		_w2063_,
		_w2064_
	);
	LUT4 #(
		.INIT('hf531)
	) name884 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1532_reg/NET0131 ,
		\g1534_reg/NET0131 ,
		_w2065_
	);
	LUT2 #(
		.INIT('h4)
	) name885 (
		\g1533_reg/NET0131 ,
		\g7961_pad ,
		_w2066_
	);
	LUT3 #(
		.INIT('ha6)
	) name886 (
		\g1496_reg/NET0131 ,
		_w2065_,
		_w2066_,
		_w2067_
	);
	LUT2 #(
		.INIT('h2)
	) name887 (
		\g1088_reg/NET0131 ,
		\g1553_reg/NET0131 ,
		_w2068_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name888 (
		\g1092_reg/NET0131 ,
		\g1554_reg/NET0131 ,
		\g1555_reg/NET0131 ,
		\g7961_pad ,
		_w2069_
	);
	LUT2 #(
		.INIT('h4)
	) name889 (
		_w2068_,
		_w2069_,
		_w2070_
	);
	LUT2 #(
		.INIT('h4)
	) name890 (
		\g1545_reg/NET0131 ,
		\g7961_pad ,
		_w2071_
	);
	LUT4 #(
		.INIT('hf531)
	) name891 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1544_reg/NET0131 ,
		\g1546_reg/NET0131 ,
		_w2072_
	);
	LUT4 #(
		.INIT('h4b44)
	) name892 (
		_w2068_,
		_w2069_,
		_w2071_,
		_w2072_,
		_w2073_
	);
	LUT2 #(
		.INIT('h4)
	) name893 (
		\g1542_reg/NET0131 ,
		\g7961_pad ,
		_w2074_
	);
	LUT4 #(
		.INIT('hf531)
	) name894 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1541_reg/NET0131 ,
		\g1543_reg/NET0131 ,
		_w2075_
	);
	LUT4 #(
		.INIT('h4b44)
	) name895 (
		_w2011_,
		_w2012_,
		_w2074_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h2)
	) name896 (
		\g1088_reg/NET0131 ,
		\g1702_reg/NET0131 ,
		_w2077_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name897 (
		\g1092_reg/NET0131 ,
		\g1703_reg/NET0131 ,
		\g1704_reg/NET0131 ,
		\g7961_pad ,
		_w2078_
	);
	LUT2 #(
		.INIT('h4)
	) name898 (
		_w2077_,
		_w2078_,
		_w2079_
	);
	LUT4 #(
		.INIT('h0002)
	) name899 (
		_w2067_,
		_w2073_,
		_w2076_,
		_w2079_,
		_w2080_
	);
	LUT4 #(
		.INIT('h8000)
	) name900 (
		\g1563_reg/NET0131 ,
		_w2054_,
		_w2064_,
		_w2080_,
		_w2081_
	);
	LUT4 #(
		.INIT('h7500)
	) name901 (
		_w2010_,
		_w2035_,
		_w2040_,
		_w2081_,
		_w2082_
	);
	LUT4 #(
		.INIT('h135f)
	) name902 (
		\g1088_reg/NET0131 ,
		\g1630_reg/NET0131 ,
		\g1636_reg/NET0131 ,
		\g7961_pad ,
		_w2083_
	);
	LUT2 #(
		.INIT('h8)
	) name903 (
		\g1092_reg/NET0131 ,
		\g1633_reg/NET0131 ,
		_w2084_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		_w2083_,
		_w2084_,
		_w2085_
	);
	LUT3 #(
		.INIT('ha6)
	) name905 (
		\g1496_reg/NET0131 ,
		_w2083_,
		_w2084_,
		_w2086_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		\g1612_reg/NET0131 ,
		\g7961_pad ,
		_w2087_
	);
	LUT4 #(
		.INIT('h153f)
	) name907 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1615_reg/NET0131 ,
		\g1618_reg/NET0131 ,
		_w2088_
	);
	LUT2 #(
		.INIT('h4)
	) name908 (
		_w2087_,
		_w2088_,
		_w2089_
	);
	LUT3 #(
		.INIT('h9a)
	) name909 (
		\g1476_reg/NET0131 ,
		_w2087_,
		_w2088_,
		_w2090_
	);
	LUT2 #(
		.INIT('h8)
	) name910 (
		\g1639_reg/NET0131 ,
		\g7961_pad ,
		_w2091_
	);
	LUT4 #(
		.INIT('h153f)
	) name911 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1642_reg/NET0131 ,
		\g1645_reg/NET0131 ,
		_w2092_
	);
	LUT2 #(
		.INIT('h4)
	) name912 (
		_w2091_,
		_w2092_,
		_w2093_
	);
	LUT3 #(
		.INIT('h9a)
	) name913 (
		\g1506_reg/NET0131 ,
		_w2091_,
		_w2092_,
		_w2094_
	);
	LUT4 #(
		.INIT('h153f)
	) name914 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1624_reg/NET0131 ,
		\g1627_reg/NET0131 ,
		_w2095_
	);
	LUT2 #(
		.INIT('h8)
	) name915 (
		\g1621_reg/NET0131 ,
		\g7961_pad ,
		_w2096_
	);
	LUT2 #(
		.INIT('h2)
	) name916 (
		_w2095_,
		_w2096_,
		_w2097_
	);
	LUT3 #(
		.INIT('ha6)
	) name917 (
		\g1486_reg/NET0131 ,
		_w2095_,
		_w2096_,
		_w2098_
	);
	LUT4 #(
		.INIT('hc800)
	) name918 (
		_w2086_,
		_w2090_,
		_w2094_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h8)
	) name919 (
		\g1648_reg/NET0131 ,
		\g7961_pad ,
		_w2100_
	);
	LUT4 #(
		.INIT('h153f)
	) name920 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1651_reg/NET0131 ,
		\g1654_reg/NET0131 ,
		_w2101_
	);
	LUT2 #(
		.INIT('h4)
	) name921 (
		_w2100_,
		_w2101_,
		_w2102_
	);
	LUT4 #(
		.INIT('h4b44)
	) name922 (
		_w2068_,
		_w2069_,
		_w2100_,
		_w2101_,
		_w2103_
	);
	LUT3 #(
		.INIT('h70)
	) name923 (
		_w2086_,
		_w2094_,
		_w2103_,
		_w2104_
	);
	LUT2 #(
		.INIT('h4)
	) name924 (
		_w2099_,
		_w2104_,
		_w2105_
	);
	LUT4 #(
		.INIT('h0015)
	) name925 (
		_w2086_,
		_w2090_,
		_w2094_,
		_w2098_,
		_w2106_
	);
	LUT2 #(
		.INIT('h2)
	) name926 (
		_w2094_,
		_w2103_,
		_w2107_
	);
	LUT3 #(
		.INIT('h13)
	) name927 (
		_w2086_,
		_w2090_,
		_w2098_,
		_w2108_
	);
	LUT3 #(
		.INIT('h45)
	) name928 (
		_w2106_,
		_w2107_,
		_w2108_,
		_w2109_
	);
	LUT3 #(
		.INIT('h8a)
	) name929 (
		_w2010_,
		_w2105_,
		_w2109_,
		_w2110_
	);
	LUT2 #(
		.INIT('h2)
	) name930 (
		\g1092_reg/NET0131 ,
		\g1700_reg/NET0131 ,
		_w2111_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name931 (
		\g1088_reg/NET0131 ,
		\g1699_reg/NET0131 ,
		\g1701_reg/NET0131 ,
		\g7961_pad ,
		_w2112_
	);
	LUT2 #(
		.INIT('h4)
	) name932 (
		_w2111_,
		_w2112_,
		_w2113_
	);
	LUT3 #(
		.INIT('h20)
	) name933 (
		\g1563_reg/NET0131 ,
		_w2007_,
		_w2008_,
		_w2114_
	);
	LUT4 #(
		.INIT('h4000)
	) name934 (
		_w2017_,
		_w2033_,
		_w2086_,
		_w2098_,
		_w2115_
	);
	LUT4 #(
		.INIT('h8000)
	) name935 (
		_w2021_,
		_w2025_,
		_w2029_,
		_w2090_,
		_w2116_
	);
	LUT4 #(
		.INIT('h8000)
	) name936 (
		\g1563_reg/NET0131 ,
		_w2107_,
		_w2115_,
		_w2116_,
		_w2117_
	);
	LUT3 #(
		.INIT('h02)
	) name937 (
		_w2113_,
		_w2114_,
		_w2117_,
		_w2118_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		\g1088_reg/NET0131 ,
		\g1695_reg/NET0131 ,
		_w2119_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name939 (
		\g1092_reg/NET0131 ,
		\g1693_reg/NET0131 ,
		\g1694_reg/NET0131 ,
		\g7961_pad ,
		_w2120_
	);
	LUT2 #(
		.INIT('h4)
	) name940 (
		_w2119_,
		_w2120_,
		_w2121_
	);
	LUT3 #(
		.INIT('hd0)
	) name941 (
		\g1088_reg/NET0131 ,
		\g1550_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w2122_
	);
	LUT2 #(
		.INIT('h8)
	) name942 (
		_w2008_,
		_w2122_,
		_w2123_
	);
	LUT4 #(
		.INIT('h45cf)
	) name943 (
		_w2008_,
		_w2111_,
		_w2112_,
		_w2122_,
		_w2124_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w2121_,
		_w2124_,
		_w2125_
	);
	LUT4 #(
		.INIT('h0080)
	) name945 (
		_w2054_,
		_w2064_,
		_w2080_,
		_w2121_,
		_w2126_
	);
	LUT2 #(
		.INIT('h4)
	) name946 (
		\g1696_reg/NET0131 ,
		\g7961_pad ,
		_w2127_
	);
	LUT4 #(
		.INIT('hf351)
	) name947 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1697_reg/NET0131 ,
		\g1698_reg/NET0131 ,
		_w2128_
	);
	LUT2 #(
		.INIT('h4)
	) name948 (
		_w2127_,
		_w2128_,
		_w2129_
	);
	LUT3 #(
		.INIT('h80)
	) name949 (
		\g1696_reg/NET0131 ,
		\g7961_pad ,
		_w2128_,
		_w2130_
	);
	LUT3 #(
		.INIT('he0)
	) name950 (
		_w2125_,
		_w2126_,
		_w2130_,
		_w2131_
	);
	LUT4 #(
		.INIT('hef00)
	) name951 (
		_w2082_,
		_w2110_,
		_w2118_,
		_w2131_,
		_w2132_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name952 (
		_w2099_,
		_w2104_,
		_w2107_,
		_w2108_,
		_w2133_
	);
	LUT3 #(
		.INIT('h80)
	) name953 (
		_w2107_,
		_w2115_,
		_w2116_,
		_w2134_
	);
	LUT3 #(
		.INIT('h20)
	) name954 (
		_w2010_,
		_w2106_,
		_w2113_,
		_w2135_
	);
	LUT3 #(
		.INIT('h20)
	) name955 (
		_w2133_,
		_w2134_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h2)
	) name956 (
		\g1088_reg/NET0131 ,
		\g1783_reg/NET0131 ,
		_w2137_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name957 (
		\g1092_reg/NET0131 ,
		\g1784_reg/NET0131 ,
		\g1785_reg/NET0131 ,
		\g7961_pad ,
		_w2138_
	);
	LUT2 #(
		.INIT('h4)
	) name958 (
		_w2137_,
		_w2138_,
		_w2139_
	);
	LUT4 #(
		.INIT('h0002)
	) name959 (
		_w2067_,
		_w2073_,
		_w2076_,
		_w2139_,
		_w2140_
	);
	LUT3 #(
		.INIT('h80)
	) name960 (
		_w2054_,
		_w2064_,
		_w2140_,
		_w2141_
	);
	LUT4 #(
		.INIT('h070f)
	) name961 (
		_w2054_,
		_w2064_,
		_w2121_,
		_w2140_,
		_w2142_
	);
	LUT4 #(
		.INIT('h0400)
	) name962 (
		_w2111_,
		_w2112_,
		_w2119_,
		_w2120_,
		_w2143_
	);
	LUT2 #(
		.INIT('h2)
	) name963 (
		_w2129_,
		_w2143_,
		_w2144_
	);
	LUT4 #(
		.INIT('h7f00)
	) name964 (
		_w2054_,
		_w2064_,
		_w2140_,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h2)
	) name965 (
		\g7961_pad ,
		_w2145_,
		_w2146_
	);
	LUT4 #(
		.INIT('h1f00)
	) name966 (
		_w2041_,
		_w2136_,
		_w2142_,
		_w2146_,
		_w2147_
	);
	LUT2 #(
		.INIT('h1)
	) name967 (
		\g1696_reg/NET0131 ,
		\g7961_pad ,
		_w2148_
	);
	LUT3 #(
		.INIT('h01)
	) name968 (
		_w2132_,
		_w2147_,
		_w2148_,
		_w2149_
	);
	LUT3 #(
		.INIT('h20)
	) name969 (
		\g1092_reg/NET0131 ,
		_w2127_,
		_w2128_,
		_w2150_
	);
	LUT3 #(
		.INIT('he0)
	) name970 (
		_w2125_,
		_w2126_,
		_w2150_,
		_w2151_
	);
	LUT4 #(
		.INIT('hef00)
	) name971 (
		_w2082_,
		_w2110_,
		_w2118_,
		_w2151_,
		_w2152_
	);
	LUT2 #(
		.INIT('h2)
	) name972 (
		\g1092_reg/NET0131 ,
		_w2145_,
		_w2153_
	);
	LUT4 #(
		.INIT('h1f00)
	) name973 (
		_w2041_,
		_w2136_,
		_w2142_,
		_w2153_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name974 (
		\g1092_reg/NET0131 ,
		\g1697_reg/NET0131 ,
		_w2155_
	);
	LUT3 #(
		.INIT('h01)
	) name975 (
		_w2152_,
		_w2154_,
		_w2155_,
		_w2156_
	);
	LUT3 #(
		.INIT('h20)
	) name976 (
		\g1088_reg/NET0131 ,
		_w2127_,
		_w2128_,
		_w2157_
	);
	LUT3 #(
		.INIT('he0)
	) name977 (
		_w2125_,
		_w2126_,
		_w2157_,
		_w2158_
	);
	LUT4 #(
		.INIT('hef00)
	) name978 (
		_w2082_,
		_w2110_,
		_w2118_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h2)
	) name979 (
		\g1088_reg/NET0131 ,
		_w2145_,
		_w2160_
	);
	LUT4 #(
		.INIT('h1f00)
	) name980 (
		_w2041_,
		_w2136_,
		_w2142_,
		_w2160_,
		_w2161_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		\g1088_reg/NET0131 ,
		\g1698_reg/NET0131 ,
		_w2162_
	);
	LUT3 #(
		.INIT('h01)
	) name982 (
		_w2159_,
		_w2161_,
		_w2162_,
		_w2163_
	);
	LUT3 #(
		.INIT('h51)
	) name983 (
		\g1186_reg/NET0131 ,
		\g1234_reg/NET0131 ,
		\g5657_pad ,
		_w2164_
	);
	LUT3 #(
		.INIT('h80)
	) name984 (
		\g499_reg/NET0131 ,
		\g544_reg/NET0131 ,
		\g5657_pad ,
		_w2165_
	);
	LUT3 #(
		.INIT('h51)
	) name985 (
		_w1508_,
		_w2164_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w2167_
	);
	LUT3 #(
		.INIT('h02)
	) name987 (
		\g1186_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w2168_
	);
	LUT4 #(
		.INIT('hae00)
	) name988 (
		_w1508_,
		_w2164_,
		_w2165_,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h2)
	) name989 (
		\g1018_reg/NET0131 ,
		\g1425_reg/NET0131 ,
		_w2170_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name990 (
		\g1024_reg/NET0131 ,
		\g1423_reg/NET0131 ,
		\g1424_reg/NET0131 ,
		\g5657_pad ,
		_w2171_
	);
	LUT2 #(
		.INIT('h2)
	) name991 (
		\g1024_reg/NET0131 ,
		\g1417_reg/NET0131 ,
		_w2172_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name992 (
		\g1018_reg/NET0131 ,
		\g1418_reg/NET0131 ,
		\g1419_reg/NET0131 ,
		\g5657_pad ,
		_w2173_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name993 (
		_w2170_,
		_w2171_,
		_w2172_,
		_w2173_,
		_w2174_
	);
	LUT2 #(
		.INIT('h4)
	) name994 (
		\g1391_reg/NET0131 ,
		\g5657_pad ,
		_w2175_
	);
	LUT4 #(
		.INIT('hf351)
	) name995 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1390_reg/NET0131 ,
		\g1392_reg/NET0131 ,
		_w2176_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		_w2175_,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h4)
	) name997 (
		\g1400_reg/NET0131 ,
		\g5657_pad ,
		_w2178_
	);
	LUT4 #(
		.INIT('hf351)
	) name998 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1399_reg/NET0131 ,
		\g1401_reg/NET0131 ,
		_w2179_
	);
	LUT4 #(
		.INIT('h0b00)
	) name999 (
		_w2175_,
		_w2176_,
		_w2178_,
		_w2179_,
		_w2180_
	);
	LUT2 #(
		.INIT('h8)
	) name1000 (
		_w2174_,
		_w2180_,
		_w2181_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		\g1409_reg/NET0131 ,
		\g5657_pad ,
		_w2182_
	);
	LUT4 #(
		.INIT('hf351)
	) name1002 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1408_reg/NET0131 ,
		\g1410_reg/NET0131 ,
		_w2183_
	);
	LUT2 #(
		.INIT('h4)
	) name1003 (
		_w2182_,
		_w2183_,
		_w2184_
	);
	LUT2 #(
		.INIT('h4)
	) name1004 (
		\g1397_reg/NET0131 ,
		\g5657_pad ,
		_w2185_
	);
	LUT4 #(
		.INIT('hf351)
	) name1005 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1396_reg/NET0131 ,
		\g1398_reg/NET0131 ,
		_w2186_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1006 (
		_w2182_,
		_w2183_,
		_w2185_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h4)
	) name1007 (
		\g1385_reg/NET0131 ,
		\g5657_pad ,
		_w2188_
	);
	LUT4 #(
		.INIT('hf351)
	) name1008 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1384_reg/NET0131 ,
		\g1386_reg/NET0131 ,
		_w2189_
	);
	LUT2 #(
		.INIT('h4)
	) name1009 (
		\g1388_reg/NET0131 ,
		\g5657_pad ,
		_w2190_
	);
	LUT4 #(
		.INIT('hf351)
	) name1010 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1387_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w2191_
	);
	LUT4 #(
		.INIT('h4044)
	) name1011 (
		_w2188_,
		_w2189_,
		_w2190_,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h4)
	) name1012 (
		\g1403_reg/NET0131 ,
		\g5657_pad ,
		_w2193_
	);
	LUT4 #(
		.INIT('hf351)
	) name1013 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1402_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		_w2194_
	);
	LUT2 #(
		.INIT('h4)
	) name1014 (
		\g1394_reg/NET0131 ,
		\g5657_pad ,
		_w2195_
	);
	LUT4 #(
		.INIT('hf351)
	) name1015 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1393_reg/NET0131 ,
		\g1395_reg/NET0131 ,
		_w2196_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		_w2195_,
		_w2196_,
		_w2197_
	);
	LUT4 #(
		.INIT('h4044)
	) name1017 (
		_w2193_,
		_w2194_,
		_w2195_,
		_w2196_,
		_w2198_
	);
	LUT2 #(
		.INIT('h4)
	) name1018 (
		\g1412_reg/NET0131 ,
		\g5657_pad ,
		_w2199_
	);
	LUT4 #(
		.INIT('hf351)
	) name1019 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1411_reg/NET0131 ,
		\g1413_reg/NET0131 ,
		_w2200_
	);
	LUT2 #(
		.INIT('h4)
	) name1020 (
		_w2199_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h4)
	) name1021 (
		\g1406_reg/NET0131 ,
		\g5657_pad ,
		_w2202_
	);
	LUT4 #(
		.INIT('hf351)
	) name1022 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1405_reg/NET0131 ,
		\g1407_reg/NET0131 ,
		_w2203_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1023 (
		_w2199_,
		_w2200_,
		_w2202_,
		_w2203_,
		_w2204_
	);
	LUT4 #(
		.INIT('h8000)
	) name1024 (
		_w2187_,
		_w2192_,
		_w2198_,
		_w2204_,
		_w2205_
	);
	LUT2 #(
		.INIT('h8)
	) name1025 (
		\g1300_reg/NET0131 ,
		\g5657_pad ,
		_w2206_
	);
	LUT4 #(
		.INIT('h135f)
	) name1026 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1303_reg/NET0131 ,
		\g1306_reg/NET0131 ,
		_w2207_
	);
	LUT2 #(
		.INIT('h4)
	) name1027 (
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT4 #(
		.INIT('hea15)
	) name1028 (
		_w2177_,
		_w2181_,
		_w2205_,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h8)
	) name1029 (
		\g1018_reg/NET0131 ,
		\g1294_reg/NET0131 ,
		_w2210_
	);
	LUT4 #(
		.INIT('h135f)
	) name1030 (
		\g1024_reg/NET0131 ,
		\g1291_reg/NET0131 ,
		\g1297_reg/NET0131 ,
		\g5657_pad ,
		_w2211_
	);
	LUT2 #(
		.INIT('h4)
	) name1031 (
		_w2210_,
		_w2211_,
		_w2212_
	);
	LUT3 #(
		.INIT('h08)
	) name1032 (
		_w2174_,
		_w2180_,
		_w2212_,
		_w2213_
	);
	LUT4 #(
		.INIT('hec13)
	) name1033 (
		_w2181_,
		_w2197_,
		_w2205_,
		_w2212_,
		_w2214_
	);
	LUT3 #(
		.INIT('h28)
	) name1034 (
		_w2169_,
		_w2209_,
		_w2214_,
		_w2215_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1035 (
		_w2188_,
		_w2189_,
		_w2206_,
		_w2207_,
		_w2216_
	);
	LUT2 #(
		.INIT('h2)
	) name1036 (
		_w2169_,
		_w2216_,
		_w2217_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1037 (
		_w2190_,
		_w2191_,
		_w2210_,
		_w2211_,
		_w2218_
	);
	LUT3 #(
		.INIT('h70)
	) name1038 (
		_w2181_,
		_w2205_,
		_w2218_,
		_w2219_
	);
	LUT4 #(
		.INIT('h4044)
	) name1039 (
		_w2190_,
		_w2191_,
		_w2210_,
		_w2211_,
		_w2220_
	);
	LUT4 #(
		.INIT('h002a)
	) name1040 (
		_w2169_,
		_w2205_,
		_w2213_,
		_w2220_,
		_w2221_
	);
	LUT2 #(
		.INIT('h4)
	) name1041 (
		_w2219_,
		_w2221_,
		_w2222_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1042 (
		_w2193_,
		_w2194_,
		_w2206_,
		_w2207_,
		_w2223_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1043 (
		_w2202_,
		_w2203_,
		_w2210_,
		_w2211_,
		_w2224_
	);
	LUT3 #(
		.INIT('hd7)
	) name1044 (
		_w2169_,
		_w2223_,
		_w2224_,
		_w2225_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1045 (
		_w2178_,
		_w2179_,
		_w2210_,
		_w2211_,
		_w2226_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1046 (
		_w2185_,
		_w2186_,
		_w2206_,
		_w2207_,
		_w2227_
	);
	LUT4 #(
		.INIT('h3993)
	) name1047 (
		_w2169_,
		_w2225_,
		_w2226_,
		_w2227_,
		_w2228_
	);
	LUT4 #(
		.INIT('h6996)
	) name1048 (
		_w2215_,
		_w2217_,
		_w2222_,
		_w2228_,
		_w2229_
	);
	LUT4 #(
		.INIT('hec13)
	) name1049 (
		_w2181_,
		_w2201_,
		_w2205_,
		_w2212_,
		_w2230_
	);
	LUT4 #(
		.INIT('hec13)
	) name1050 (
		_w2181_,
		_w2184_,
		_w2205_,
		_w2208_,
		_w2231_
	);
	LUT2 #(
		.INIT('h8)
	) name1051 (
		\g1243_reg/NET0131 ,
		_w2169_,
		_w2232_
	);
	LUT3 #(
		.INIT('h04)
	) name1052 (
		\g1196_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w2233_
	);
	LUT2 #(
		.INIT('h4)
	) name1053 (
		\g1224_reg/NET0131 ,
		\g3229_pad ,
		_w2234_
	);
	LUT4 #(
		.INIT('h0302)
	) name1054 (
		\g1227_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		\g3229_pad ,
		_w2235_
	);
	LUT3 #(
		.INIT('h20)
	) name1055 (
		_w2233_,
		_w2234_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h4)
	) name1056 (
		_w2166_,
		_w2236_,
		_w2237_
	);
	LUT4 #(
		.INIT('h009f)
	) name1057 (
		_w2230_,
		_w2231_,
		_w2232_,
		_w2237_,
		_w2238_
	);
	LUT3 #(
		.INIT('h8f)
	) name1058 (
		\g1196_reg/NET0131 ,
		_w2229_,
		_w2238_,
		_w2239_
	);
	LUT2 #(
		.INIT('h2)
	) name1059 (
		_w1534_,
		_w1605_,
		_w2240_
	);
	LUT2 #(
		.INIT('h4)
	) name1060 (
		_w1583_,
		_w2240_,
		_w2241_
	);
	LUT3 #(
		.INIT('h32)
	) name1061 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		_w2242_
	);
	LUT4 #(
		.INIT('h0054)
	) name1062 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1910_reg/NET0131 ,
		_w2243_
	);
	LUT2 #(
		.INIT('h8)
	) name1063 (
		_w1607_,
		_w2243_,
		_w2244_
	);
	LUT3 #(
		.INIT('h8c)
	) name1064 (
		_w1604_,
		_w2242_,
		_w2244_,
		_w2245_
	);
	LUT3 #(
		.INIT('h45)
	) name1065 (
		_w1613_,
		_w2241_,
		_w2245_,
		_w2246_
	);
	LUT2 #(
		.INIT('h4)
	) name1066 (
		\g2115_reg/NET0131 ,
		\g5657_pad ,
		_w2247_
	);
	LUT4 #(
		.INIT('hf351)
	) name1067 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2114_reg/NET0131 ,
		\g2116_reg/NET0131 ,
		_w2248_
	);
	LUT3 #(
		.INIT('h8a)
	) name1068 (
		\g1880_reg/NET0131 ,
		_w2247_,
		_w2248_,
		_w2249_
	);
	LUT3 #(
		.INIT('h80)
	) name1069 (
		\g1880_reg/NET0131 ,
		_w1539_,
		_w1544_,
		_w2250_
	);
	LUT3 #(
		.INIT('h13)
	) name1070 (
		_w1571_,
		_w2249_,
		_w2250_,
		_w2251_
	);
	LUT4 #(
		.INIT('hef00)
	) name1071 (
		_w1509_,
		_w1510_,
		_w1511_,
		_w1607_,
		_w2252_
	);
	LUT3 #(
		.INIT('hb0)
	) name1072 (
		_w2241_,
		_w2245_,
		_w2252_,
		_w2253_
	);
	LUT3 #(
		.INIT('h15)
	) name1073 (
		_w2246_,
		_w2251_,
		_w2253_,
		_w2254_
	);
	LUT2 #(
		.INIT('h4)
	) name1074 (
		_w1588_,
		_w2240_,
		_w2255_
	);
	LUT4 #(
		.INIT('h0054)
	) name1075 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1909_reg/NET0131 ,
		_w2256_
	);
	LUT2 #(
		.INIT('h8)
	) name1076 (
		_w1607_,
		_w2256_,
		_w2257_
	);
	LUT3 #(
		.INIT('h8c)
	) name1077 (
		_w1604_,
		_w2242_,
		_w2257_,
		_w2258_
	);
	LUT3 #(
		.INIT('h45)
	) name1078 (
		_w1613_,
		_w2255_,
		_w2258_,
		_w2259_
	);
	LUT3 #(
		.INIT('h8a)
	) name1079 (
		_w2252_,
		_w2255_,
		_w2258_,
		_w2260_
	);
	LUT3 #(
		.INIT('h23)
	) name1080 (
		_w2251_,
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h4)
	) name1081 (
		_w1587_,
		_w2240_,
		_w2262_
	);
	LUT4 #(
		.INIT('h0054)
	) name1082 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1911_reg/NET0131 ,
		_w2263_
	);
	LUT2 #(
		.INIT('h8)
	) name1083 (
		_w1607_,
		_w2263_,
		_w2264_
	);
	LUT3 #(
		.INIT('h8c)
	) name1084 (
		_w1604_,
		_w2242_,
		_w2264_,
		_w2265_
	);
	LUT3 #(
		.INIT('h45)
	) name1085 (
		_w1613_,
		_w2262_,
		_w2265_,
		_w2266_
	);
	LUT3 #(
		.INIT('h8a)
	) name1086 (
		_w2252_,
		_w2262_,
		_w2265_,
		_w2267_
	);
	LUT3 #(
		.INIT('h13)
	) name1087 (
		_w2251_,
		_w2266_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('h4)
	) name1088 (
		_w1586_,
		_w2240_,
		_w2269_
	);
	LUT4 #(
		.INIT('h0054)
	) name1089 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1912_reg/NET0131 ,
		_w2270_
	);
	LUT2 #(
		.INIT('h8)
	) name1090 (
		_w1607_,
		_w2270_,
		_w2271_
	);
	LUT3 #(
		.INIT('h8c)
	) name1091 (
		_w1604_,
		_w2242_,
		_w2271_,
		_w2272_
	);
	LUT3 #(
		.INIT('h45)
	) name1092 (
		_w1613_,
		_w2269_,
		_w2272_,
		_w2273_
	);
	LUT3 #(
		.INIT('h8a)
	) name1093 (
		_w2252_,
		_w2269_,
		_w2272_,
		_w2274_
	);
	LUT3 #(
		.INIT('h23)
	) name1094 (
		_w2251_,
		_w2273_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h4)
	) name1095 (
		_w1607_,
		_w1613_,
		_w2276_
	);
	LUT4 #(
		.INIT('h1000)
	) name1096 (
		_w1509_,
		_w1510_,
		_w1511_,
		_w1613_,
		_w2277_
	);
	LUT2 #(
		.INIT('h1)
	) name1097 (
		_w2276_,
		_w2277_,
		_w2278_
	);
	LUT3 #(
		.INIT('h54)
	) name1098 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		_w2279_
	);
	LUT2 #(
		.INIT('h2)
	) name1099 (
		_w1534_,
		_w2279_,
		_w2280_
	);
	LUT4 #(
		.INIT('h0054)
	) name1100 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1913_reg/NET0131 ,
		_w2281_
	);
	LUT2 #(
		.INIT('h8)
	) name1101 (
		_w1607_,
		_w2281_,
		_w2282_
	);
	LUT3 #(
		.INIT('h8c)
	) name1102 (
		_w1604_,
		_w2242_,
		_w2282_,
		_w2283_
	);
	LUT4 #(
		.INIT('h7f33)
	) name1103 (
		_w1575_,
		_w2278_,
		_w2280_,
		_w2283_,
		_w2284_
	);
	LUT4 #(
		.INIT('h0054)
	) name1104 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1914_reg/NET0131 ,
		_w2285_
	);
	LUT2 #(
		.INIT('h8)
	) name1105 (
		_w1607_,
		_w2285_,
		_w2286_
	);
	LUT3 #(
		.INIT('h8c)
	) name1106 (
		_w1604_,
		_w2242_,
		_w2286_,
		_w2287_
	);
	LUT4 #(
		.INIT('h7f33)
	) name1107 (
		_w1579_,
		_w2278_,
		_w2280_,
		_w2287_,
		_w2288_
	);
	LUT3 #(
		.INIT('hc4)
	) name1108 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g168_reg/NET0131 ,
		_w2289_
	);
	LUT4 #(
		.INIT('hb000)
	) name1109 (
		_w1698_,
		_w1699_,
		_w1735_,
		_w2289_,
		_w2290_
	);
	LUT4 #(
		.INIT('h4044)
	) name1110 (
		_w1695_,
		_w1696_,
		_w1745_,
		_w1746_,
		_w2291_
	);
	LUT2 #(
		.INIT('h4)
	) name1111 (
		_w1750_,
		_w2291_,
		_w2292_
	);
	LUT4 #(
		.INIT('h8000)
	) name1112 (
		_w1724_,
		_w1727_,
		_w1744_,
		_w2292_,
		_w2293_
	);
	LUT4 #(
		.INIT('h4000)
	) name1113 (
		_w1700_,
		_w1704_,
		_w1707_,
		_w1710_,
		_w2294_
	);
	LUT3 #(
		.INIT('h15)
	) name1114 (
		_w2290_,
		_w2293_,
		_w2294_,
		_w2295_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name1115 (
		_w1695_,
		_w1696_,
		_w1789_,
		_w1790_,
		_w2296_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1116 (
		_w1755_,
		_w1756_,
		_w1763_,
		_w1764_,
		_w2297_
	);
	LUT4 #(
		.INIT('hdd0d)
	) name1117 (
		_w1767_,
		_w1768_,
		_w1776_,
		_w1777_,
		_w2298_
	);
	LUT4 #(
		.INIT('h8000)
	) name1118 (
		_w1821_,
		_w2296_,
		_w2297_,
		_w2298_,
		_w2299_
	);
	LUT4 #(
		.INIT('h0200)
	) name1119 (
		_w1772_,
		_w1773_,
		_w1785_,
		_w1786_,
		_w2300_
	);
	LUT4 #(
		.INIT('h0020)
	) name1120 (
		_w1759_,
		_w1760_,
		_w1781_,
		_w1782_,
		_w2301_
	);
	LUT3 #(
		.INIT('h80)
	) name1121 (
		_w1795_,
		_w2300_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h8)
	) name1122 (
		_w2299_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h1)
	) name1123 (
		_w1830_,
		_w2303_,
		_w2304_
	);
	LUT3 #(
		.INIT('h15)
	) name1124 (
		\g105_reg/NET0131 ,
		_w2295_,
		_w2304_,
		_w2305_
	);
	LUT4 #(
		.INIT('h0040)
	) name1125 (
		_w1801_,
		_w1804_,
		_w1809_,
		_w1814_,
		_w2306_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1126 (
		_w1698_,
		_w1699_,
		_w1745_,
		_w1746_,
		_w2307_
	);
	LUT4 #(
		.INIT('h4044)
	) name1127 (
		_w1695_,
		_w1696_,
		_w1748_,
		_w1749_,
		_w2308_
	);
	LUT2 #(
		.INIT('h8)
	) name1128 (
		_w2307_,
		_w2308_,
		_w2309_
	);
	LUT4 #(
		.INIT('h8000)
	) name1129 (
		_w1724_,
		_w1727_,
		_w1744_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h8)
	) name1130 (
		_w1711_,
		_w2310_,
		_w2311_
	);
	LUT3 #(
		.INIT('h40)
	) name1131 (
		\g105_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w2312_
	);
	LUT3 #(
		.INIT('hd0)
	) name1132 (
		_w1737_,
		_w2306_,
		_w2312_,
		_w2313_
	);
	LUT3 #(
		.INIT('hd0)
	) name1133 (
		_w1737_,
		_w2306_,
		_w2311_,
		_w2314_
	);
	LUT4 #(
		.INIT('h0111)
	) name1134 (
		_w1830_,
		_w2290_,
		_w2293_,
		_w2294_,
		_w2315_
	);
	LUT4 #(
		.INIT('h0020)
	) name1135 (
		_w1776_,
		_w1777_,
		_w1789_,
		_w1790_,
		_w2316_
	);
	LUT4 #(
		.INIT('h0400)
	) name1136 (
		_w1755_,
		_w1756_,
		_w1763_,
		_w1764_,
		_w2317_
	);
	LUT4 #(
		.INIT('h0040)
	) name1137 (
		_w1695_,
		_w1696_,
		_w1767_,
		_w1768_,
		_w2318_
	);
	LUT3 #(
		.INIT('h80)
	) name1138 (
		_w2316_,
		_w2317_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h4)
	) name1139 (
		_w1697_,
		_w1821_,
		_w2320_
	);
	LUT4 #(
		.INIT('hc800)
	) name1140 (
		_w2299_,
		_w2302_,
		_w2319_,
		_w2320_,
		_w2321_
	);
	LUT4 #(
		.INIT('h4404)
	) name1141 (
		_w1695_,
		_w1696_,
		_w1781_,
		_w1782_,
		_w2322_
	);
	LUT4 #(
		.INIT('h00b0)
	) name1142 (
		_w1695_,
		_w1696_,
		_w1781_,
		_w1782_,
		_w2323_
	);
	LUT3 #(
		.INIT('h02)
	) name1143 (
		_w1821_,
		_w2322_,
		_w2323_,
		_w2324_
	);
	LUT4 #(
		.INIT('h44b4)
	) name1144 (
		_w1695_,
		_w1696_,
		_w1767_,
		_w1768_,
		_w2325_
	);
	LUT2 #(
		.INIT('h2)
	) name1145 (
		_w1791_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h8)
	) name1146 (
		_w2324_,
		_w2326_,
		_w2327_
	);
	LUT4 #(
		.INIT('ha080)
	) name1147 (
		_w1821_,
		_w2299_,
		_w2302_,
		_w2319_,
		_w2328_
	);
	LUT4 #(
		.INIT('h0090)
	) name1148 (
		_w1697_,
		_w1783_,
		_w1821_,
		_w2325_,
		_w2329_
	);
	LUT2 #(
		.INIT('h1)
	) name1149 (
		_w1791_,
		_w2329_,
		_w2330_
	);
	LUT4 #(
		.INIT('haaab)
	) name1150 (
		_w2321_,
		_w2327_,
		_w2328_,
		_w2330_,
		_w2331_
	);
	LUT2 #(
		.INIT('h8)
	) name1151 (
		_w2315_,
		_w2331_,
		_w2332_
	);
	LUT4 #(
		.INIT('h1011)
	) name1152 (
		_w2305_,
		_w2313_,
		_w2314_,
		_w2332_,
		_w2333_
	);
	LUT3 #(
		.INIT('he2)
	) name1153 (
		\g195_reg/NET0131 ,
		\g7961_pad ,
		_w2333_,
		_w2334_
	);
	LUT3 #(
		.INIT('he4)
	) name1154 (
		\g1092_reg/NET0131 ,
		\g198_reg/NET0131 ,
		_w2333_,
		_w2335_
	);
	LUT3 #(
		.INIT('he4)
	) name1155 (
		\g1088_reg/NET0131 ,
		\g201_reg/NET0131 ,
		_w2333_,
		_w2336_
	);
	LUT4 #(
		.INIT('h4044)
	) name1156 (
		_w1846_,
		_w1847_,
		_w1849_,
		_w1850_,
		_w2337_
	);
	LUT3 #(
		.INIT('h32)
	) name1157 (
		_w1855_,
		_w1859_,
		_w2337_,
		_w2338_
	);
	LUT3 #(
		.INIT('h22)
	) name1158 (
		_w1855_,
		_w1859_,
		_w2337_,
		_w2339_
	);
	LUT2 #(
		.INIT('h8)
	) name1159 (
		_w1911_,
		_w2338_,
		_w2340_
	);
	LUT3 #(
		.INIT('h13)
	) name1160 (
		_w1894_,
		_w2339_,
		_w2340_,
		_w2341_
	);
	LUT4 #(
		.INIT('h0103)
	) name1161 (
		_w1894_,
		_w1918_,
		_w2339_,
		_w2340_,
		_w2342_
	);
	LUT2 #(
		.INIT('h1)
	) name1162 (
		\g793_reg/NET0131 ,
		_w2342_,
		_w2343_
	);
	LUT4 #(
		.INIT('h4044)
	) name1163 (
		_w1846_,
		_w1847_,
		_w1857_,
		_w1858_,
		_w2344_
	);
	LUT3 #(
		.INIT('h40)
	) name1164 (
		_w1907_,
		_w1910_,
		_w2344_,
		_w2345_
	);
	LUT2 #(
		.INIT('h8)
	) name1165 (
		_w1904_,
		_w2345_,
		_w2346_
	);
	LUT4 #(
		.INIT('h0200)
	) name1166 (
		_w1894_,
		_w1975_,
		_w1978_,
		_w2346_,
		_w2347_
	);
	LUT3 #(
		.INIT('h10)
	) name1167 (
		\g793_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w2348_
	);
	LUT3 #(
		.INIT('h40)
	) name1168 (
		_w1950_,
		_w2347_,
		_w2348_,
		_w2349_
	);
	LUT3 #(
		.INIT('h20)
	) name1169 (
		_w1851_,
		_w1950_,
		_w2347_,
		_w2350_
	);
	LUT2 #(
		.INIT('h4)
	) name1170 (
		_w1848_,
		_w1919_,
		_w2351_
	);
	LUT4 #(
		.INIT('h0400)
	) name1171 (
		_w1935_,
		_w1936_,
		_w1970_,
		_w1971_,
		_w2352_
	);
	LUT4 #(
		.INIT('h0400)
	) name1172 (
		_w1923_,
		_w1924_,
		_w1965_,
		_w1966_,
		_w2353_
	);
	LUT3 #(
		.INIT('h80)
	) name1173 (
		_w1942_,
		_w2352_,
		_w2353_,
		_w2354_
	);
	LUT4 #(
		.INIT('h0400)
	) name1174 (
		_w1953_,
		_w1954_,
		_w1957_,
		_w1958_,
		_w2355_
	);
	LUT4 #(
		.INIT('h0400)
	) name1175 (
		_w1927_,
		_w1928_,
		_w1931_,
		_w1932_,
		_w2356_
	);
	LUT4 #(
		.INIT('h0400)
	) name1176 (
		_w1846_,
		_w1847_,
		_w1961_,
		_w1962_,
		_w2357_
	);
	LUT3 #(
		.INIT('h80)
	) name1177 (
		_w2355_,
		_w2356_,
		_w2357_,
		_w2358_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1178 (
		_w1846_,
		_w1847_,
		_w1931_,
		_w1932_,
		_w2359_
	);
	LUT2 #(
		.INIT('h8)
	) name1179 (
		_w1919_,
		_w2359_,
		_w2360_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1180 (
		_w1953_,
		_w1954_,
		_w1957_,
		_w1958_,
		_w2361_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1181 (
		_w1927_,
		_w1928_,
		_w1961_,
		_w1962_,
		_w2362_
	);
	LUT4 #(
		.INIT('h8000)
	) name1182 (
		_w1919_,
		_w2359_,
		_w2361_,
		_w2362_,
		_w2363_
	);
	LUT4 #(
		.INIT('h8880)
	) name1183 (
		_w2351_,
		_w2354_,
		_w2358_,
		_w2363_,
		_w2364_
	);
	LUT4 #(
		.INIT('h8880)
	) name1184 (
		_w1919_,
		_w2354_,
		_w2358_,
		_w2363_,
		_w2365_
	);
	LUT4 #(
		.INIT('h8004)
	) name1185 (
		_w1848_,
		_w1919_,
		_w1942_,
		_w1963_,
		_w2366_
	);
	LUT2 #(
		.INIT('h6)
	) name1186 (
		_w1933_,
		_w2366_,
		_w2367_
	);
	LUT3 #(
		.INIT('h45)
	) name1187 (
		_w2364_,
		_w2365_,
		_w2367_,
		_w2368_
	);
	LUT2 #(
		.INIT('h2)
	) name1188 (
		_w2342_,
		_w2368_,
		_w2369_
	);
	LUT4 #(
		.INIT('h1011)
	) name1189 (
		_w2343_,
		_w2349_,
		_w2350_,
		_w2369_,
		_w2370_
	);
	LUT3 #(
		.INIT('he4)
	) name1190 (
		\g7961_pad ,
		\g882_reg/NET0131 ,
		_w2370_,
		_w2371_
	);
	LUT3 #(
		.INIT('he4)
	) name1191 (
		\g1092_reg/NET0131 ,
		\g885_reg/NET0131 ,
		_w2370_,
		_w2372_
	);
	LUT3 #(
		.INIT('he4)
	) name1192 (
		\g1088_reg/NET0131 ,
		\g888_reg/NET0131 ,
		_w2370_,
		_w2373_
	);
	LUT2 #(
		.INIT('h1)
	) name1193 (
		\g789_reg/NET0131 ,
		_w2342_,
		_w2374_
	);
	LUT3 #(
		.INIT('h10)
	) name1194 (
		\g789_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w2375_
	);
	LUT3 #(
		.INIT('h40)
	) name1195 (
		_w1950_,
		_w2347_,
		_w2375_,
		_w2376_
	);
	LUT4 #(
		.INIT('hbb4b)
	) name1196 (
		_w1846_,
		_w1847_,
		_w1940_,
		_w1941_,
		_w2377_
	);
	LUT3 #(
		.INIT('h6c)
	) name1197 (
		_w1919_,
		_w1963_,
		_w2377_,
		_w2378_
	);
	LUT3 #(
		.INIT('h45)
	) name1198 (
		_w2364_,
		_w2365_,
		_w2378_,
		_w2379_
	);
	LUT2 #(
		.INIT('h2)
	) name1199 (
		_w2342_,
		_w2379_,
		_w2380_
	);
	LUT4 #(
		.INIT('h0203)
	) name1200 (
		_w2350_,
		_w2374_,
		_w2376_,
		_w2380_,
		_w2381_
	);
	LUT3 #(
		.INIT('he4)
	) name1201 (
		\g7961_pad ,
		\g918_reg/NET0131 ,
		_w2381_,
		_w2382_
	);
	LUT3 #(
		.INIT('he4)
	) name1202 (
		\g1092_reg/NET0131 ,
		\g921_reg/NET0131 ,
		_w2381_,
		_w2383_
	);
	LUT3 #(
		.INIT('he4)
	) name1203 (
		\g1088_reg/NET0131 ,
		\g924_reg/NET0131 ,
		_w2381_,
		_w2384_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		\g797_reg/NET0131 ,
		_w2342_,
		_w2385_
	);
	LUT3 #(
		.INIT('h10)
	) name1205 (
		\g797_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w2386_
	);
	LUT3 #(
		.INIT('h40)
	) name1206 (
		_w1950_,
		_w2347_,
		_w2386_,
		_w2387_
	);
	LUT3 #(
		.INIT('hb0)
	) name1207 (
		_w1848_,
		_w1919_,
		_w1933_,
		_w2388_
	);
	LUT3 #(
		.INIT('h4b)
	) name1208 (
		_w1848_,
		_w1919_,
		_w1933_,
		_w2389_
	);
	LUT4 #(
		.INIT('h5a6a)
	) name1209 (
		_w1955_,
		_w2360_,
		_w2366_,
		_w2388_,
		_w2390_
	);
	LUT3 #(
		.INIT('h45)
	) name1210 (
		_w2364_,
		_w2365_,
		_w2390_,
		_w2391_
	);
	LUT2 #(
		.INIT('h2)
	) name1211 (
		_w2342_,
		_w2391_,
		_w2392_
	);
	LUT4 #(
		.INIT('h0203)
	) name1212 (
		_w2350_,
		_w2385_,
		_w2387_,
		_w2392_,
		_w2393_
	);
	LUT3 #(
		.INIT('he4)
	) name1213 (
		\g7961_pad ,
		\g927_reg/NET0131 ,
		_w2393_,
		_w2394_
	);
	LUT3 #(
		.INIT('he4)
	) name1214 (
		\g1088_reg/NET0131 ,
		\g933_reg/NET0131 ,
		_w2393_,
		_w2395_
	);
	LUT3 #(
		.INIT('he4)
	) name1215 (
		\g1092_reg/NET0131 ,
		\g930_reg/NET0131 ,
		_w2393_,
		_w2396_
	);
	LUT2 #(
		.INIT('h4)
	) name1216 (
		\g7961_pad ,
		\g954_reg/NET0131 ,
		_w2397_
	);
	LUT2 #(
		.INIT('h8)
	) name1217 (
		_w2342_,
		_w2364_,
		_w2398_
	);
	LUT2 #(
		.INIT('h2)
	) name1218 (
		_w1876_,
		_w2342_,
		_w2399_
	);
	LUT4 #(
		.INIT('h0400)
	) name1219 (
		_w1849_,
		_w1850_,
		_w1874_,
		_w1875_,
		_w2400_
	);
	LUT3 #(
		.INIT('h40)
	) name1220 (
		_w1950_,
		_w2347_,
		_w2400_,
		_w2401_
	);
	LUT4 #(
		.INIT('h000b)
	) name1221 (
		_w2350_,
		_w2398_,
		_w2399_,
		_w2401_,
		_w2402_
	);
	LUT2 #(
		.INIT('h1)
	) name1222 (
		\g7961_pad ,
		\g954_reg/NET0131 ,
		_w2403_
	);
	LUT3 #(
		.INIT('hb4)
	) name1223 (
		_w1848_,
		_w1919_,
		_w1955_,
		_w2404_
	);
	LUT4 #(
		.INIT('hb004)
	) name1224 (
		_w1848_,
		_w1919_,
		_w1925_,
		_w1955_,
		_w2405_
	);
	LUT3 #(
		.INIT('h20)
	) name1225 (
		_w2366_,
		_w2389_,
		_w2405_,
		_w2406_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1226 (
		_w1846_,
		_w1847_,
		_w1935_,
		_w1936_,
		_w2407_
	);
	LUT3 #(
		.INIT('h13)
	) name1227 (
		_w1919_,
		_w2352_,
		_w2407_,
		_w2408_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1228 (
		_w1923_,
		_w1924_,
		_w1970_,
		_w1971_,
		_w2409_
	);
	LUT4 #(
		.INIT('h00ec)
	) name1229 (
		_w1919_,
		_w2352_,
		_w2407_,
		_w2409_,
		_w2410_
	);
	LUT3 #(
		.INIT('hb4)
	) name1230 (
		_w1848_,
		_w1919_,
		_w1967_,
		_w2411_
	);
	LUT2 #(
		.INIT('h8)
	) name1231 (
		_w2410_,
		_w2411_,
		_w2412_
	);
	LUT3 #(
		.INIT('hb4)
	) name1232 (
		_w1848_,
		_w1919_,
		_w1929_,
		_w2413_
	);
	LUT3 #(
		.INIT('h80)
	) name1233 (
		_w2410_,
		_w2411_,
		_w2413_,
		_w2414_
	);
	LUT3 #(
		.INIT('h15)
	) name1234 (
		_w1959_,
		_w2406_,
		_w2414_,
		_w2415_
	);
	LUT3 #(
		.INIT('h80)
	) name1235 (
		_w1959_,
		_w2406_,
		_w2414_,
		_w2416_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w1918_,
		_w2365_,
		_w2417_
	);
	LUT2 #(
		.INIT('h8)
	) name1237 (
		_w2341_,
		_w2417_,
		_w2418_
	);
	LUT4 #(
		.INIT('h0200)
	) name1238 (
		_w2341_,
		_w2415_,
		_w2416_,
		_w2417_,
		_w2419_
	);
	LUT3 #(
		.INIT('h23)
	) name1239 (
		_w2350_,
		_w2403_,
		_w2419_,
		_w2420_
	);
	LUT3 #(
		.INIT('hea)
	) name1240 (
		_w2397_,
		_w2402_,
		_w2420_,
		_w2421_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		\g1092_reg/NET0131 ,
		\g957_reg/NET0131 ,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		\g1092_reg/NET0131 ,
		\g957_reg/NET0131 ,
		_w2423_
	);
	LUT3 #(
		.INIT('h0b)
	) name1243 (
		_w2350_,
		_w2419_,
		_w2423_,
		_w2424_
	);
	LUT3 #(
		.INIT('hec)
	) name1244 (
		_w2402_,
		_w2422_,
		_w2424_,
		_w2425_
	);
	LUT2 #(
		.INIT('h4)
	) name1245 (
		\g1088_reg/NET0131 ,
		\g960_reg/NET0131 ,
		_w2426_
	);
	LUT2 #(
		.INIT('h1)
	) name1246 (
		\g1088_reg/NET0131 ,
		\g960_reg/NET0131 ,
		_w2427_
	);
	LUT3 #(
		.INIT('h0b)
	) name1247 (
		_w2350_,
		_w2419_,
		_w2427_,
		_w2428_
	);
	LUT3 #(
		.INIT('hec)
	) name1248 (
		_w2402_,
		_w2426_,
		_w2428_,
		_w2429_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1249 (
		_w2077_,
		_w2078_,
		_w2127_,
		_w2128_,
		_w2430_
	);
	LUT4 #(
		.INIT('h0002)
	) name1250 (
		_w2067_,
		_w2073_,
		_w2076_,
		_w2121_,
		_w2431_
	);
	LUT4 #(
		.INIT('h8000)
	) name1251 (
		_w2054_,
		_w2064_,
		_w2113_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h8)
	) name1252 (
		_w2430_,
		_w2432_,
		_w2433_
	);
	LUT3 #(
		.INIT('h10)
	) name1253 (
		_w2041_,
		_w2110_,
		_w2433_,
		_w2434_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1254 (
		_w2111_,
		_w2112_,
		_w2127_,
		_w2128_,
		_w2435_
	);
	LUT3 #(
		.INIT('h54)
	) name1255 (
		_w2121_,
		_w2123_,
		_w2435_,
		_w2436_
	);
	LUT3 #(
		.INIT('h44)
	) name1256 (
		_w2121_,
		_w2123_,
		_w2435_,
		_w2437_
	);
	LUT4 #(
		.INIT('h8000)
	) name1257 (
		_w2054_,
		_w2064_,
		_w2080_,
		_w2436_,
		_w2438_
	);
	LUT3 #(
		.INIT('h01)
	) name1258 (
		_w2141_,
		_w2437_,
		_w2438_,
		_w2439_
	);
	LUT2 #(
		.INIT('h4)
	) name1259 (
		_w2129_,
		_w2143_,
		_w2440_
	);
	LUT4 #(
		.INIT('h0040)
	) name1260 (
		_w2018_,
		_w2019_,
		_w2083_,
		_w2084_,
		_w2441_
	);
	LUT4 #(
		.INIT('h0040)
	) name1261 (
		_w2022_,
		_w2023_,
		_w2026_,
		_w2027_,
		_w2442_
	);
	LUT3 #(
		.INIT('h80)
	) name1262 (
		_w2093_,
		_w2441_,
		_w2442_,
		_w2443_
	);
	LUT4 #(
		.INIT('h0400)
	) name1263 (
		_w2087_,
		_w2088_,
		_w2127_,
		_w2128_,
		_w2444_
	);
	LUT4 #(
		.INIT('h0040)
	) name1264 (
		_w2030_,
		_w2031_,
		_w2095_,
		_w2096_,
		_w2445_
	);
	LUT4 #(
		.INIT('h0400)
	) name1265 (
		_w2014_,
		_w2015_,
		_w2100_,
		_w2101_,
		_w2446_
	);
	LUT3 #(
		.INIT('h80)
	) name1266 (
		_w2444_,
		_w2445_,
		_w2446_,
		_w2447_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1267 (
		_w2014_,
		_w2015_,
		_w2127_,
		_w2128_,
		_w2448_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name1268 (
		_w2030_,
		_w2031_,
		_w2095_,
		_w2096_,
		_w2449_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1269 (
		_w2087_,
		_w2088_,
		_w2100_,
		_w2101_,
		_w2450_
	);
	LUT4 #(
		.INIT('h8000)
	) name1270 (
		_w2143_,
		_w2448_,
		_w2449_,
		_w2450_,
		_w2451_
	);
	LUT4 #(
		.INIT('h8880)
	) name1271 (
		_w2440_,
		_w2443_,
		_w2447_,
		_w2451_,
		_w2452_
	);
	LUT4 #(
		.INIT('h8880)
	) name1272 (
		_w2143_,
		_w2443_,
		_w2447_,
		_w2451_,
		_w2453_
	);
	LUT4 #(
		.INIT('h8100)
	) name1273 (
		_w2028_,
		_w2089_,
		_w2129_,
		_w2143_,
		_w2454_
	);
	LUT2 #(
		.INIT('h9)
	) name1274 (
		_w2032_,
		_w2454_,
		_w2455_
	);
	LUT3 #(
		.INIT('h54)
	) name1275 (
		_w2452_,
		_w2453_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h2)
	) name1276 (
		_w2439_,
		_w2456_,
		_w2457_
	);
	LUT3 #(
		.INIT('h20)
	) name1277 (
		\g7961_pad ,
		_w2434_,
		_w2457_,
		_w2458_
	);
	LUT4 #(
		.INIT('hef00)
	) name1278 (
		_w2041_,
		_w2110_,
		_w2433_,
		_w2439_,
		_w2459_
	);
	LUT2 #(
		.INIT('h4)
	) name1279 (
		\g1481_reg/NET0131 ,
		\g7961_pad ,
		_w2460_
	);
	LUT2 #(
		.INIT('h4)
	) name1280 (
		_w2459_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		\g1576_reg/NET0131 ,
		\g7961_pad ,
		_w2462_
	);
	LUT3 #(
		.INIT('h01)
	) name1282 (
		_w2458_,
		_w2461_,
		_w2462_,
		_w2463_
	);
	LUT2 #(
		.INIT('h1)
	) name1283 (
		\g2270_reg/NET0131 ,
		\g7961_pad ,
		_w2464_
	);
	LUT2 #(
		.INIT('h2)
	) name1284 (
		\g2270_reg/NET0131 ,
		\g7961_pad ,
		_w2465_
	);
	LUT4 #(
		.INIT('h0040)
	) name1285 (
		_w1279_,
		_w1282_,
		_w1343_,
		_w1345_,
		_w2466_
	);
	LUT3 #(
		.INIT('h80)
	) name1286 (
		_w1348_,
		_w1351_,
		_w1355_,
		_w2467_
	);
	LUT4 #(
		.INIT('h4044)
	) name1287 (
		_w1251_,
		_w1252_,
		_w1362_,
		_w1363_,
		_w2468_
	);
	LUT4 #(
		.INIT('h8000)
	) name1288 (
		_w1348_,
		_w1351_,
		_w1355_,
		_w2468_,
		_w2469_
	);
	LUT3 #(
		.INIT('h80)
	) name1289 (
		_w1326_,
		_w1337_,
		_w2469_,
		_w2470_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1290 (
		_w1356_,
		_w1357_,
		_w1366_,
		_w1367_,
		_w2471_
	);
	LUT4 #(
		.INIT('h8000)
	) name1291 (
		_w1326_,
		_w1337_,
		_w2469_,
		_w2471_,
		_w2472_
	);
	LUT3 #(
		.INIT('hd0)
	) name1292 (
		_w1333_,
		_w2466_,
		_w2472_,
		_w2473_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1293 (
		_w1251_,
		_w1252_,
		_w1366_,
		_w1367_,
		_w2474_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1294 (
		_w1356_,
		_w1357_,
		_w1362_,
		_w1363_,
		_w2475_
	);
	LUT2 #(
		.INIT('h8)
	) name1295 (
		_w2474_,
		_w2475_,
		_w2476_
	);
	LUT4 #(
		.INIT('h8000)
	) name1296 (
		_w1326_,
		_w1337_,
		_w2467_,
		_w2476_,
		_w2477_
	);
	LUT3 #(
		.INIT('hc4)
	) name1297 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g2246_reg/NET0131 ,
		_w2478_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1298 (
		_w1312_,
		_w1362_,
		_w1363_,
		_w2478_,
		_w2479_
	);
	LUT4 #(
		.INIT('h007f)
	) name1299 (
		_w1326_,
		_w1337_,
		_w1374_,
		_w2479_,
		_w2480_
	);
	LUT2 #(
		.INIT('h4)
	) name1300 (
		_w1368_,
		_w1369_,
		_w2481_
	);
	LUT4 #(
		.INIT('h0400)
	) name1301 (
		_w1254_,
		_w1255_,
		_w1288_,
		_w1289_,
		_w2482_
	);
	LUT4 #(
		.INIT('h0200)
	) name1302 (
		_w1263_,
		_w1264_,
		_w1283_,
		_w1284_,
		_w2483_
	);
	LUT3 #(
		.INIT('h80)
	) name1303 (
		_w1302_,
		_w2482_,
		_w2483_,
		_w2484_
	);
	LUT4 #(
		.INIT('h0040)
	) name1304 (
		_w1270_,
		_w1271_,
		_w1274_,
		_w1275_,
		_w2485_
	);
	LUT4 #(
		.INIT('h0400)
	) name1305 (
		_w1258_,
		_w1259_,
		_w1366_,
		_w1367_,
		_w2486_
	);
	LUT4 #(
		.INIT('h8000)
	) name1306 (
		_w1297_,
		_w1306_,
		_w2485_,
		_w2486_,
		_w2487_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1307 (
		_w1295_,
		_w1296_,
		_w1366_,
		_w1367_,
		_w2488_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name1308 (
		_w1270_,
		_w1271_,
		_w1274_,
		_w1275_,
		_w2489_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1309 (
		_w1258_,
		_w1259_,
		_w1304_,
		_w1305_,
		_w2490_
	);
	LUT4 #(
		.INIT('h8000)
	) name1310 (
		_w1369_,
		_w2488_,
		_w2489_,
		_w2490_,
		_w2491_
	);
	LUT4 #(
		.INIT('h8880)
	) name1311 (
		_w2481_,
		_w2484_,
		_w2487_,
		_w2491_,
		_w2492_
	);
	LUT3 #(
		.INIT('h40)
	) name1312 (
		_w2477_,
		_w2480_,
		_w2492_,
		_w2493_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1313 (
		_w1333_,
		_w2466_,
		_w2472_,
		_w2493_,
		_w2494_
	);
	LUT4 #(
		.INIT('h8100)
	) name1314 (
		_w1260_,
		_w1302_,
		_w1368_,
		_w1369_,
		_w2495_
	);
	LUT2 #(
		.INIT('h9)
	) name1315 (
		_w1306_,
		_w2495_,
		_w2496_
	);
	LUT4 #(
		.INIT('h8880)
	) name1316 (
		_w1369_,
		_w2484_,
		_w2487_,
		_w2491_,
		_w2497_
	);
	LUT3 #(
		.INIT('h04)
	) name1317 (
		_w2477_,
		_w2480_,
		_w2497_,
		_w2498_
	);
	LUT4 #(
		.INIT('h0004)
	) name1318 (
		_w2477_,
		_w2480_,
		_w2496_,
		_w2497_,
		_w2499_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1319 (
		_w1333_,
		_w2466_,
		_w2472_,
		_w2499_,
		_w2500_
	);
	LUT3 #(
		.INIT('h45)
	) name1320 (
		\g2175_reg/NET0131 ,
		_w2477_,
		_w2480_,
		_w2501_
	);
	LUT2 #(
		.INIT('h4)
	) name1321 (
		\g2175_reg/NET0131 ,
		_w2472_,
		_w2502_
	);
	LUT4 #(
		.INIT('h020f)
	) name1322 (
		_w1333_,
		_w2466_,
		_w2501_,
		_w2502_,
		_w2503_
	);
	LUT4 #(
		.INIT('h0100)
	) name1323 (
		_w2464_,
		_w2494_,
		_w2500_,
		_w2503_,
		_w2504_
	);
	LUT2 #(
		.INIT('he)
	) name1324 (
		_w2465_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h1)
	) name1325 (
		\g1088_reg/NET0131 ,
		\g2276_reg/NET0131 ,
		_w2506_
	);
	LUT2 #(
		.INIT('h4)
	) name1326 (
		\g1088_reg/NET0131 ,
		\g2276_reg/NET0131 ,
		_w2507_
	);
	LUT4 #(
		.INIT('h0010)
	) name1327 (
		_w2494_,
		_w2500_,
		_w2503_,
		_w2506_,
		_w2508_
	);
	LUT2 #(
		.INIT('he)
	) name1328 (
		_w2507_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h1)
	) name1329 (
		\g1092_reg/NET0131 ,
		\g2273_reg/NET0131 ,
		_w2510_
	);
	LUT2 #(
		.INIT('h4)
	) name1330 (
		\g1092_reg/NET0131 ,
		\g2273_reg/NET0131 ,
		_w2511_
	);
	LUT4 #(
		.INIT('h0010)
	) name1331 (
		_w2494_,
		_w2500_,
		_w2503_,
		_w2510_,
		_w2512_
	);
	LUT2 #(
		.INIT('he)
	) name1332 (
		_w2511_,
		_w2512_,
		_w2513_
	);
	LUT3 #(
		.INIT('h20)
	) name1333 (
		\g1092_reg/NET0131 ,
		_w2434_,
		_w2457_,
		_w2514_
	);
	LUT2 #(
		.INIT('h2)
	) name1334 (
		\g1092_reg/NET0131 ,
		\g1481_reg/NET0131 ,
		_w2515_
	);
	LUT2 #(
		.INIT('h4)
	) name1335 (
		_w2459_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h1)
	) name1336 (
		\g1092_reg/NET0131 ,
		\g1579_reg/NET0131 ,
		_w2517_
	);
	LUT3 #(
		.INIT('h01)
	) name1337 (
		_w2514_,
		_w2516_,
		_w2517_,
		_w2518_
	);
	LUT2 #(
		.INIT('h1)
	) name1338 (
		\g2306_reg/NET0131 ,
		\g7961_pad ,
		_w2519_
	);
	LUT2 #(
		.INIT('h2)
	) name1339 (
		\g2306_reg/NET0131 ,
		\g7961_pad ,
		_w2520_
	);
	LUT3 #(
		.INIT('h45)
	) name1340 (
		\g2170_reg/NET0131 ,
		_w2477_,
		_w2480_,
		_w2521_
	);
	LUT2 #(
		.INIT('h4)
	) name1341 (
		\g2170_reg/NET0131 ,
		_w2472_,
		_w2522_
	);
	LUT4 #(
		.INIT('h020f)
	) name1342 (
		_w1333_,
		_w2466_,
		_w2521_,
		_w2522_,
		_w2523_
	);
	LUT4 #(
		.INIT('h9655)
	) name1343 (
		_w1260_,
		_w1302_,
		_w1368_,
		_w1369_,
		_w2524_
	);
	LUT4 #(
		.INIT('h0004)
	) name1344 (
		_w2477_,
		_w2480_,
		_w2497_,
		_w2524_,
		_w2525_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1345 (
		_w1333_,
		_w2466_,
		_w2472_,
		_w2525_,
		_w2526_
	);
	LUT4 #(
		.INIT('h0010)
	) name1346 (
		_w2494_,
		_w2519_,
		_w2523_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('he)
	) name1347 (
		_w2520_,
		_w2527_,
		_w2528_
	);
	LUT3 #(
		.INIT('h20)
	) name1348 (
		\g1088_reg/NET0131 ,
		_w2434_,
		_w2457_,
		_w2529_
	);
	LUT2 #(
		.INIT('h2)
	) name1349 (
		\g1088_reg/NET0131 ,
		\g1481_reg/NET0131 ,
		_w2530_
	);
	LUT2 #(
		.INIT('h4)
	) name1350 (
		_w2459_,
		_w2530_,
		_w2531_
	);
	LUT2 #(
		.INIT('h1)
	) name1351 (
		\g1088_reg/NET0131 ,
		\g1582_reg/NET0131 ,
		_w2532_
	);
	LUT3 #(
		.INIT('h01)
	) name1352 (
		_w2529_,
		_w2531_,
		_w2532_,
		_w2533_
	);
	LUT2 #(
		.INIT('h1)
	) name1353 (
		\g1092_reg/NET0131 ,
		\g2309_reg/NET0131 ,
		_w2534_
	);
	LUT2 #(
		.INIT('h4)
	) name1354 (
		\g1092_reg/NET0131 ,
		\g2309_reg/NET0131 ,
		_w2535_
	);
	LUT4 #(
		.INIT('h0004)
	) name1355 (
		_w2494_,
		_w2523_,
		_w2526_,
		_w2534_,
		_w2536_
	);
	LUT2 #(
		.INIT('he)
	) name1356 (
		_w2535_,
		_w2536_,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name1357 (
		\g1088_reg/NET0131 ,
		\g2312_reg/NET0131 ,
		_w2538_
	);
	LUT2 #(
		.INIT('h4)
	) name1358 (
		\g1088_reg/NET0131 ,
		\g2312_reg/NET0131 ,
		_w2539_
	);
	LUT4 #(
		.INIT('h0004)
	) name1359 (
		_w2494_,
		_w2523_,
		_w2526_,
		_w2538_,
		_w2540_
	);
	LUT2 #(
		.INIT('he)
	) name1360 (
		_w2539_,
		_w2540_,
		_w2541_
	);
	LUT2 #(
		.INIT('h1)
	) name1361 (
		\g2315_reg/NET0131 ,
		\g7961_pad ,
		_w2542_
	);
	LUT2 #(
		.INIT('h2)
	) name1362 (
		\g2315_reg/NET0131 ,
		\g7961_pad ,
		_w2543_
	);
	LUT3 #(
		.INIT('h45)
	) name1363 (
		\g2180_reg/NET0131 ,
		_w2477_,
		_w2480_,
		_w2544_
	);
	LUT2 #(
		.INIT('h4)
	) name1364 (
		\g2180_reg/NET0131 ,
		_w2472_,
		_w2545_
	);
	LUT4 #(
		.INIT('h020f)
	) name1365 (
		_w1333_,
		_w2466_,
		_w2544_,
		_w2545_,
		_w2546_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1366 (
		_w1274_,
		_w1275_,
		_w1304_,
		_w1305_,
		_w2547_
	);
	LUT4 #(
		.INIT('hebee)
	) name1367 (
		_w1276_,
		_w1306_,
		_w1368_,
		_w1369_,
		_w2548_
	);
	LUT3 #(
		.INIT('he0)
	) name1368 (
		_w1276_,
		_w2495_,
		_w2548_,
		_w2549_
	);
	LUT3 #(
		.INIT('h45)
	) name1369 (
		_w1306_,
		_w1368_,
		_w1369_,
		_w2550_
	);
	LUT4 #(
		.INIT('h4044)
	) name1370 (
		_w1304_,
		_w1305_,
		_w1366_,
		_w1367_,
		_w2551_
	);
	LUT2 #(
		.INIT('h8)
	) name1371 (
		_w1369_,
		_w2551_,
		_w2552_
	);
	LUT3 #(
		.INIT('h2a)
	) name1372 (
		_w1276_,
		_w1369_,
		_w2551_,
		_w2553_
	);
	LUT3 #(
		.INIT('h20)
	) name1373 (
		_w2495_,
		_w2550_,
		_w2553_,
		_w2554_
	);
	LUT2 #(
		.INIT('h2)
	) name1374 (
		_w2549_,
		_w2554_,
		_w2555_
	);
	LUT2 #(
		.INIT('h8)
	) name1375 (
		_w2498_,
		_w2555_,
		_w2556_
	);
	LUT3 #(
		.INIT('h8c)
	) name1376 (
		_w2473_,
		_w2546_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h1)
	) name1377 (
		_w2494_,
		_w2542_,
		_w2558_
	);
	LUT3 #(
		.INIT('hea)
	) name1378 (
		_w2543_,
		_w2557_,
		_w2558_,
		_w2559_
	);
	LUT2 #(
		.INIT('h1)
	) name1379 (
		\g1092_reg/NET0131 ,
		\g2318_reg/NET0131 ,
		_w2560_
	);
	LUT2 #(
		.INIT('h4)
	) name1380 (
		\g1092_reg/NET0131 ,
		\g2318_reg/NET0131 ,
		_w2561_
	);
	LUT2 #(
		.INIT('h1)
	) name1381 (
		_w2494_,
		_w2560_,
		_w2562_
	);
	LUT3 #(
		.INIT('hec)
	) name1382 (
		_w2557_,
		_w2561_,
		_w2562_,
		_w2563_
	);
	LUT3 #(
		.INIT('h15)
	) name1383 (
		\g101_reg/NET0131 ,
		_w2295_,
		_w2304_,
		_w2564_
	);
	LUT3 #(
		.INIT('h40)
	) name1384 (
		\g101_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w2565_
	);
	LUT3 #(
		.INIT('hd0)
	) name1385 (
		_w1737_,
		_w2306_,
		_w2565_,
		_w2566_
	);
	LUT4 #(
		.INIT('h8400)
	) name1386 (
		_w1697_,
		_w1769_,
		_w1783_,
		_w1821_,
		_w2567_
	);
	LUT4 #(
		.INIT('h1233)
	) name1387 (
		_w1697_,
		_w1769_,
		_w1783_,
		_w1821_,
		_w2568_
	);
	LUT4 #(
		.INIT('haaab)
	) name1388 (
		_w2321_,
		_w2328_,
		_w2567_,
		_w2568_,
		_w2569_
	);
	LUT2 #(
		.INIT('h8)
	) name1389 (
		_w2315_,
		_w2569_,
		_w2570_
	);
	LUT4 #(
		.INIT('h0203)
	) name1390 (
		_w2314_,
		_w2564_,
		_w2566_,
		_w2570_,
		_w2571_
	);
	LUT3 #(
		.INIT('he2)
	) name1391 (
		\g231_reg/NET0131 ,
		\g7961_pad ,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('h1)
	) name1392 (
		\g1088_reg/NET0131 ,
		\g2321_reg/NET0131 ,
		_w2573_
	);
	LUT2 #(
		.INIT('h4)
	) name1393 (
		\g1088_reg/NET0131 ,
		\g2321_reg/NET0131 ,
		_w2574_
	);
	LUT2 #(
		.INIT('h1)
	) name1394 (
		_w2494_,
		_w2573_,
		_w2575_
	);
	LUT3 #(
		.INIT('hec)
	) name1395 (
		_w2557_,
		_w2574_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h2)
	) name1396 (
		\g2342_reg/NET0131 ,
		\g7961_pad ,
		_w2577_
	);
	LUT3 #(
		.INIT('h8a)
	) name1397 (
		_w1269_,
		_w2477_,
		_w2480_,
		_w2578_
	);
	LUT2 #(
		.INIT('h8)
	) name1398 (
		_w1269_,
		_w2472_,
		_w2579_
	);
	LUT4 #(
		.INIT('h020f)
	) name1399 (
		_w1333_,
		_w2466_,
		_w2578_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h4)
	) name1400 (
		_w2494_,
		_w2580_,
		_w2581_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		\g2342_reg/NET0131 ,
		\g7961_pad ,
		_w2582_
	);
	LUT4 #(
		.INIT('h0a9a)
	) name1402 (
		_w1265_,
		_w1368_,
		_w1369_,
		_w2551_,
		_w2583_
	);
	LUT3 #(
		.INIT('h20)
	) name1403 (
		_w2495_,
		_w2550_,
		_w2583_,
		_w2584_
	);
	LUT4 #(
		.INIT('h8188)
	) name1404 (
		_w1276_,
		_w1285_,
		_w1368_,
		_w1369_,
		_w2585_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1405 (
		_w1254_,
		_w1255_,
		_w1288_,
		_w1289_,
		_w2586_
	);
	LUT4 #(
		.INIT('h8188)
	) name1406 (
		_w1256_,
		_w1290_,
		_w1368_,
		_w1369_,
		_w2587_
	);
	LUT2 #(
		.INIT('h8)
	) name1407 (
		_w2585_,
		_w2587_,
		_w2588_
	);
	LUT3 #(
		.INIT('h65)
	) name1408 (
		_w1297_,
		_w1368_,
		_w1369_,
		_w2589_
	);
	LUT4 #(
		.INIT('h5595)
	) name1409 (
		_w1272_,
		_w2584_,
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h2)
	) name1410 (
		_w2498_,
		_w2590_,
		_w2591_
	);
	LUT3 #(
		.INIT('h23)
	) name1411 (
		_w2473_,
		_w2582_,
		_w2591_,
		_w2592_
	);
	LUT3 #(
		.INIT('hea)
	) name1412 (
		_w2577_,
		_w2581_,
		_w2592_,
		_w2593_
	);
	LUT2 #(
		.INIT('h4)
	) name1413 (
		\g1092_reg/NET0131 ,
		\g2345_reg/NET0131 ,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		\g1092_reg/NET0131 ,
		\g2345_reg/NET0131 ,
		_w2595_
	);
	LUT3 #(
		.INIT('h0b)
	) name1415 (
		_w2473_,
		_w2591_,
		_w2595_,
		_w2596_
	);
	LUT3 #(
		.INIT('hec)
	) name1416 (
		_w2581_,
		_w2594_,
		_w2596_,
		_w2597_
	);
	LUT2 #(
		.INIT('h4)
	) name1417 (
		\g1088_reg/NET0131 ,
		\g2348_reg/NET0131 ,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name1418 (
		\g1088_reg/NET0131 ,
		\g2348_reg/NET0131 ,
		_w2599_
	);
	LUT3 #(
		.INIT('h0b)
	) name1419 (
		_w2473_,
		_w2591_,
		_w2599_,
		_w2600_
	);
	LUT3 #(
		.INIT('hec)
	) name1420 (
		_w2581_,
		_w2598_,
		_w2600_,
		_w2601_
	);
	LUT3 #(
		.INIT('he4)
	) name1421 (
		\g1092_reg/NET0131 ,
		\g234_reg/NET0131 ,
		_w2571_,
		_w2602_
	);
	LUT3 #(
		.INIT('he4)
	) name1422 (
		\g1088_reg/NET0131 ,
		\g237_reg/NET0131 ,
		_w2571_,
		_w2603_
	);
	LUT4 #(
		.INIT('h69cc)
	) name1423 (
		_w2028_,
		_w2089_,
		_w2129_,
		_w2143_,
		_w2604_
	);
	LUT3 #(
		.INIT('h45)
	) name1424 (
		_w2452_,
		_w2453_,
		_w2604_,
		_w2605_
	);
	LUT2 #(
		.INIT('h2)
	) name1425 (
		_w2439_,
		_w2605_,
		_w2606_
	);
	LUT3 #(
		.INIT('h20)
	) name1426 (
		\g7961_pad ,
		_w2434_,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h4)
	) name1427 (
		\g1476_reg/NET0131 ,
		\g7961_pad ,
		_w2608_
	);
	LUT2 #(
		.INIT('h4)
	) name1428 (
		_w2459_,
		_w2608_,
		_w2609_
	);
	LUT2 #(
		.INIT('h1)
	) name1429 (
		\g1612_reg/NET0131 ,
		\g7961_pad ,
		_w2610_
	);
	LUT3 #(
		.INIT('h01)
	) name1430 (
		_w2607_,
		_w2609_,
		_w2610_,
		_w2611_
	);
	LUT3 #(
		.INIT('h20)
	) name1431 (
		\g1092_reg/NET0131 ,
		_w2434_,
		_w2606_,
		_w2612_
	);
	LUT2 #(
		.INIT('h2)
	) name1432 (
		\g1092_reg/NET0131 ,
		\g1476_reg/NET0131 ,
		_w2613_
	);
	LUT2 #(
		.INIT('h4)
	) name1433 (
		_w2459_,
		_w2613_,
		_w2614_
	);
	LUT2 #(
		.INIT('h1)
	) name1434 (
		\g1092_reg/NET0131 ,
		\g1615_reg/NET0131 ,
		_w2615_
	);
	LUT3 #(
		.INIT('h01)
	) name1435 (
		_w2612_,
		_w2614_,
		_w2615_,
		_w2616_
	);
	LUT3 #(
		.INIT('h20)
	) name1436 (
		\g1088_reg/NET0131 ,
		_w2434_,
		_w2606_,
		_w2617_
	);
	LUT2 #(
		.INIT('h2)
	) name1437 (
		\g1088_reg/NET0131 ,
		\g1476_reg/NET0131 ,
		_w2618_
	);
	LUT2 #(
		.INIT('h4)
	) name1438 (
		_w2459_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h1)
	) name1439 (
		\g1088_reg/NET0131 ,
		\g1618_reg/NET0131 ,
		_w2620_
	);
	LUT3 #(
		.INIT('h01)
	) name1440 (
		_w2617_,
		_w2619_,
		_w2620_,
		_w2621_
	);
	LUT4 #(
		.INIT('hedee)
	) name1441 (
		_w2032_,
		_w2097_,
		_w2129_,
		_w2143_,
		_w2622_
	);
	LUT3 #(
		.INIT('he0)
	) name1442 (
		_w2097_,
		_w2454_,
		_w2622_,
		_w2623_
	);
	LUT4 #(
		.INIT('h4044)
	) name1443 (
		_w2030_,
		_w2031_,
		_w2127_,
		_w2128_,
		_w2624_
	);
	LUT2 #(
		.INIT('h8)
	) name1444 (
		_w2143_,
		_w2624_,
		_w2625_
	);
	LUT4 #(
		.INIT('h2022)
	) name1445 (
		_w2095_,
		_w2096_,
		_w2127_,
		_w2128_,
		_w2626_
	);
	LUT3 #(
		.INIT('h13)
	) name1446 (
		_w2143_,
		_w2445_,
		_w2626_,
		_w2627_
	);
	LUT3 #(
		.INIT('h02)
	) name1447 (
		_w2454_,
		_w2625_,
		_w2627_,
		_w2628_
	);
	LUT4 #(
		.INIT('h5545)
	) name1448 (
		_w2452_,
		_w2453_,
		_w2623_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h2)
	) name1449 (
		_w2439_,
		_w2629_,
		_w2630_
	);
	LUT3 #(
		.INIT('h20)
	) name1450 (
		\g7961_pad ,
		_w2434_,
		_w2630_,
		_w2631_
	);
	LUT2 #(
		.INIT('h4)
	) name1451 (
		\g1486_reg/NET0131 ,
		\g7961_pad ,
		_w2632_
	);
	LUT2 #(
		.INIT('h4)
	) name1452 (
		_w2459_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h1)
	) name1453 (
		\g1621_reg/NET0131 ,
		\g7961_pad ,
		_w2634_
	);
	LUT3 #(
		.INIT('h01)
	) name1454 (
		_w2631_,
		_w2633_,
		_w2634_,
		_w2635_
	);
	LUT3 #(
		.INIT('h20)
	) name1455 (
		\g1092_reg/NET0131 ,
		_w2434_,
		_w2630_,
		_w2636_
	);
	LUT2 #(
		.INIT('h2)
	) name1456 (
		\g1092_reg/NET0131 ,
		\g1486_reg/NET0131 ,
		_w2637_
	);
	LUT2 #(
		.INIT('h4)
	) name1457 (
		_w2459_,
		_w2637_,
		_w2638_
	);
	LUT2 #(
		.INIT('h1)
	) name1458 (
		\g1092_reg/NET0131 ,
		\g1624_reg/NET0131 ,
		_w2639_
	);
	LUT3 #(
		.INIT('h01)
	) name1459 (
		_w2636_,
		_w2638_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h1)
	) name1460 (
		_w1830_,
		_w2328_,
		_w2641_
	);
	LUT3 #(
		.INIT('h15)
	) name1461 (
		\g109_reg/NET0131 ,
		_w2295_,
		_w2641_,
		_w2642_
	);
	LUT3 #(
		.INIT('h40)
	) name1462 (
		\g109_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w2643_
	);
	LUT3 #(
		.INIT('hd0)
	) name1463 (
		_w1737_,
		_w2306_,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name1464 (
		_w1697_,
		_w1830_,
		_w2645_
	);
	LUT2 #(
		.INIT('h8)
	) name1465 (
		_w2295_,
		_w2645_,
		_w2646_
	);
	LUT3 #(
		.INIT('h2a)
	) name1466 (
		\g7961_pad ,
		_w2295_,
		_w2645_,
		_w2647_
	);
	LUT3 #(
		.INIT('h80)
	) name1467 (
		\g7961_pad ,
		_w1711_,
		_w2310_,
		_w2648_
	);
	LUT3 #(
		.INIT('hd0)
	) name1468 (
		_w1737_,
		_w2306_,
		_w2648_,
		_w2649_
	);
	LUT4 #(
		.INIT('heee0)
	) name1469 (
		_w2642_,
		_w2644_,
		_w2647_,
		_w2649_,
		_w2650_
	);
	LUT3 #(
		.INIT('h63)
	) name1470 (
		_w1697_,
		_w1791_,
		_w1821_,
		_w2651_
	);
	LUT2 #(
		.INIT('h2)
	) name1471 (
		_w1778_,
		_w2325_,
		_w2652_
	);
	LUT3 #(
		.INIT('h20)
	) name1472 (
		_w2324_,
		_w2651_,
		_w2652_,
		_w2653_
	);
	LUT3 #(
		.INIT('h51)
	) name1473 (
		_w1778_,
		_w2329_,
		_w2651_,
		_w2654_
	);
	LUT4 #(
		.INIT('haaab)
	) name1474 (
		_w2321_,
		_w2328_,
		_w2653_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h8)
	) name1475 (
		_w2315_,
		_w2655_,
		_w2656_
	);
	LUT4 #(
		.INIT('he2ee)
	) name1476 (
		\g240_reg/NET0131 ,
		\g7961_pad ,
		_w2314_,
		_w2656_,
		_w2657_
	);
	LUT2 #(
		.INIT('h4)
	) name1477 (
		_w2650_,
		_w2657_,
		_w2658_
	);
	LUT3 #(
		.INIT('h20)
	) name1478 (
		\g1088_reg/NET0131 ,
		_w2434_,
		_w2630_,
		_w2659_
	);
	LUT2 #(
		.INIT('h2)
	) name1479 (
		\g1088_reg/NET0131 ,
		\g1486_reg/NET0131 ,
		_w2660_
	);
	LUT2 #(
		.INIT('h4)
	) name1480 (
		_w2459_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		\g1088_reg/NET0131 ,
		\g1627_reg/NET0131 ,
		_w2662_
	);
	LUT3 #(
		.INIT('h01)
	) name1482 (
		_w2659_,
		_w2661_,
		_w2662_,
		_w2663_
	);
	LUT3 #(
		.INIT('h2a)
	) name1483 (
		\g1092_reg/NET0131 ,
		_w2295_,
		_w2645_,
		_w2664_
	);
	LUT3 #(
		.INIT('h80)
	) name1484 (
		\g1092_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w2665_
	);
	LUT3 #(
		.INIT('hd0)
	) name1485 (
		_w1737_,
		_w2306_,
		_w2665_,
		_w2666_
	);
	LUT4 #(
		.INIT('heee0)
	) name1486 (
		_w2642_,
		_w2644_,
		_w2664_,
		_w2666_,
		_w2667_
	);
	LUT4 #(
		.INIT('he4ee)
	) name1487 (
		\g1092_reg/NET0131 ,
		\g243_reg/NET0131 ,
		_w2314_,
		_w2656_,
		_w2668_
	);
	LUT2 #(
		.INIT('h4)
	) name1488 (
		_w2667_,
		_w2668_,
		_w2669_
	);
	LUT2 #(
		.INIT('h4)
	) name1489 (
		\g1092_reg/NET0131 ,
		\g1651_reg/NET0131 ,
		_w2670_
	);
	LUT4 #(
		.INIT('h0100)
	) name1490 (
		_w2141_,
		_w2437_,
		_w2438_,
		_w2452_,
		_w2671_
	);
	LUT4 #(
		.INIT('hef00)
	) name1491 (
		_w2041_,
		_w2110_,
		_w2433_,
		_w2671_,
		_w2672_
	);
	LUT3 #(
		.INIT('h0d)
	) name1492 (
		_w2070_,
		_w2459_,
		_w2672_,
		_w2673_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		\g1092_reg/NET0131 ,
		\g1651_reg/NET0131 ,
		_w2674_
	);
	LUT4 #(
		.INIT('h0001)
	) name1494 (
		_w2141_,
		_w2437_,
		_w2438_,
		_w2453_,
		_w2675_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1495 (
		_w2095_,
		_w2096_,
		_w2127_,
		_w2128_,
		_w2676_
	);
	LUT3 #(
		.INIT('h13)
	) name1496 (
		_w2143_,
		_w2445_,
		_w2676_,
		_w2677_
	);
	LUT3 #(
		.INIT('h02)
	) name1497 (
		_w2454_,
		_w2625_,
		_w2677_,
		_w2678_
	);
	LUT3 #(
		.INIT('h45)
	) name1498 (
		_w2024_,
		_w2129_,
		_w2143_,
		_w2679_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1499 (
		_w2018_,
		_w2019_,
		_w2127_,
		_w2128_,
		_w2680_
	);
	LUT3 #(
		.INIT('h13)
	) name1500 (
		_w2143_,
		_w2441_,
		_w2680_,
		_w2681_
	);
	LUT4 #(
		.INIT('h4044)
	) name1501 (
		_w2022_,
		_w2023_,
		_w2127_,
		_w2128_,
		_w2682_
	);
	LUT4 #(
		.INIT('h2022)
	) name1502 (
		_w2083_,
		_w2084_,
		_w2127_,
		_w2128_,
		_w2683_
	);
	LUT3 #(
		.INIT('h57)
	) name1503 (
		_w2143_,
		_w2682_,
		_w2683_,
		_w2684_
	);
	LUT3 #(
		.INIT('h10)
	) name1504 (
		_w2679_,
		_w2681_,
		_w2684_,
		_w2685_
	);
	LUT3 #(
		.INIT('h9a)
	) name1505 (
		_w2093_,
		_w2129_,
		_w2143_,
		_w2686_
	);
	LUT4 #(
		.INIT('h8188)
	) name1506 (
		_w2016_,
		_w2093_,
		_w2129_,
		_w2143_,
		_w2687_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1507 (
		_w2102_,
		_w2678_,
		_w2685_,
		_w2687_,
		_w2688_
	);
	LUT2 #(
		.INIT('h8)
	) name1508 (
		_w2675_,
		_w2688_,
		_w2689_
	);
	LUT3 #(
		.INIT('h23)
	) name1509 (
		_w2434_,
		_w2674_,
		_w2689_,
		_w2690_
	);
	LUT3 #(
		.INIT('hea)
	) name1510 (
		_w2670_,
		_w2673_,
		_w2690_,
		_w2691_
	);
	LUT2 #(
		.INIT('h2)
	) name1511 (
		\g1648_reg/NET0131 ,
		\g7961_pad ,
		_w2692_
	);
	LUT2 #(
		.INIT('h1)
	) name1512 (
		\g1648_reg/NET0131 ,
		\g7961_pad ,
		_w2693_
	);
	LUT3 #(
		.INIT('h0b)
	) name1513 (
		_w2434_,
		_w2689_,
		_w2693_,
		_w2694_
	);
	LUT3 #(
		.INIT('hec)
	) name1514 (
		_w2673_,
		_w2692_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h4)
	) name1515 (
		\g1088_reg/NET0131 ,
		\g1654_reg/NET0131 ,
		_w2696_
	);
	LUT2 #(
		.INIT('h1)
	) name1516 (
		\g1088_reg/NET0131 ,
		\g1654_reg/NET0131 ,
		_w2697_
	);
	LUT3 #(
		.INIT('h0b)
	) name1517 (
		_w2434_,
		_w2689_,
		_w2697_,
		_w2698_
	);
	LUT3 #(
		.INIT('hec)
	) name1518 (
		_w2673_,
		_w2696_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h2)
	) name1519 (
		\g267_reg/NET0131 ,
		\g7961_pad ,
		_w2700_
	);
	LUT2 #(
		.INIT('h4)
	) name1520 (
		_w1830_,
		_w2321_,
		_w2701_
	);
	LUT2 #(
		.INIT('h8)
	) name1521 (
		_w2295_,
		_w2701_,
		_w2702_
	);
	LUT3 #(
		.INIT('h2a)
	) name1522 (
		_w1730_,
		_w2295_,
		_w2304_,
		_w2703_
	);
	LUT3 #(
		.INIT('h80)
	) name1523 (
		_w1711_,
		_w1730_,
		_w2310_,
		_w2704_
	);
	LUT3 #(
		.INIT('hd0)
	) name1524 (
		_w1737_,
		_w2306_,
		_w2704_,
		_w2705_
	);
	LUT4 #(
		.INIT('h000b)
	) name1525 (
		_w2314_,
		_w2702_,
		_w2703_,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('h1)
	) name1526 (
		\g267_reg/NET0131 ,
		\g7961_pad ,
		_w2707_
	);
	LUT3 #(
		.INIT('h9c)
	) name1527 (
		_w1697_,
		_w1778_,
		_w1821_,
		_w2708_
	);
	LUT4 #(
		.INIT('h81c0)
	) name1528 (
		_w1697_,
		_w1778_,
		_w1795_,
		_w1821_,
		_w2709_
	);
	LUT3 #(
		.INIT('h20)
	) name1529 (
		_w2329_,
		_w2651_,
		_w2709_,
		_w2710_
	);
	LUT4 #(
		.INIT('h2d22)
	) name1530 (
		_w1772_,
		_w1773_,
		_w1785_,
		_w1786_,
		_w2711_
	);
	LUT4 #(
		.INIT('h81c0)
	) name1531 (
		_w1697_,
		_w1774_,
		_w1787_,
		_w1821_,
		_w2712_
	);
	LUT4 #(
		.INIT('h8c00)
	) name1532 (
		_w1697_,
		_w1761_,
		_w1821_,
		_w2317_,
		_w2713_
	);
	LUT4 #(
		.INIT('h4044)
	) name1533 (
		_w1755_,
		_w1756_,
		_w1763_,
		_w1764_,
		_w2714_
	);
	LUT4 #(
		.INIT('h1000)
	) name1534 (
		_w1697_,
		_w1761_,
		_w1821_,
		_w2714_,
		_w2715_
	);
	LUT3 #(
		.INIT('ha8)
	) name1535 (
		_w2712_,
		_w2713_,
		_w2715_,
		_w2716_
	);
	LUT4 #(
		.INIT('h7e3f)
	) name1536 (
		_w1697_,
		_w1761_,
		_w1765_,
		_w1821_,
		_w2717_
	);
	LUT2 #(
		.INIT('h2)
	) name1537 (
		_w2712_,
		_w2717_,
		_w2718_
	);
	LUT4 #(
		.INIT('h2e2a)
	) name1538 (
		_w1757_,
		_w2710_,
		_w2716_,
		_w2718_,
		_w2719_
	);
	LUT3 #(
		.INIT('h80)
	) name1539 (
		_w2295_,
		_w2641_,
		_w2719_,
		_w2720_
	);
	LUT3 #(
		.INIT('h23)
	) name1540 (
		_w2314_,
		_w2707_,
		_w2720_,
		_w2721_
	);
	LUT3 #(
		.INIT('hea)
	) name1541 (
		_w2700_,
		_w2706_,
		_w2721_,
		_w2722_
	);
	LUT2 #(
		.INIT('h4)
	) name1542 (
		\g1092_reg/NET0131 ,
		\g270_reg/NET0131 ,
		_w2723_
	);
	LUT2 #(
		.INIT('h1)
	) name1543 (
		\g1092_reg/NET0131 ,
		\g270_reg/NET0131 ,
		_w2724_
	);
	LUT3 #(
		.INIT('h0b)
	) name1544 (
		_w2314_,
		_w2720_,
		_w2724_,
		_w2725_
	);
	LUT3 #(
		.INIT('hec)
	) name1545 (
		_w2706_,
		_w2723_,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h4)
	) name1546 (
		\g1088_reg/NET0131 ,
		\g273_reg/NET0131 ,
		_w2727_
	);
	LUT2 #(
		.INIT('h1)
	) name1547 (
		\g1088_reg/NET0131 ,
		\g273_reg/NET0131 ,
		_w2728_
	);
	LUT3 #(
		.INIT('h0b)
	) name1548 (
		_w2314_,
		_w2720_,
		_w2728_,
		_w2729_
	);
	LUT3 #(
		.INIT('hec)
	) name1549 (
		_w2706_,
		_w2727_,
		_w2729_,
		_w2730_
	);
	LUT3 #(
		.INIT('h70)
	) name1550 (
		_w1534_,
		_w1601_,
		_w1613_,
		_w2731_
	);
	LUT4 #(
		.INIT('h0054)
	) name1551 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1916_reg/NET0131 ,
		_w2732_
	);
	LUT3 #(
		.INIT('h4c)
	) name1552 (
		_w1607_,
		_w2242_,
		_w2732_,
		_w2733_
	);
	LUT4 #(
		.INIT('h1000)
	) name1553 (
		_w1509_,
		_w1510_,
		_w1511_,
		_w2242_,
		_w2734_
	);
	LUT2 #(
		.INIT('h1)
	) name1554 (
		_w2733_,
		_w2734_,
		_w2735_
	);
	LUT3 #(
		.INIT('h07)
	) name1555 (
		_w1582_,
		_w2240_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('he)
	) name1556 (
		_w2731_,
		_w2736_,
		_w2737_
	);
	LUT4 #(
		.INIT('h0054)
	) name1557 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1917_reg/NET0131 ,
		_w2738_
	);
	LUT3 #(
		.INIT('h4c)
	) name1558 (
		_w1607_,
		_w2242_,
		_w2738_,
		_w2739_
	);
	LUT4 #(
		.INIT('hbbb0)
	) name1559 (
		_w1580_,
		_w2240_,
		_w2734_,
		_w2739_,
		_w2740_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w1613_,
		_w2740_,
		_w2741_
	);
	LUT2 #(
		.INIT('h2)
	) name1561 (
		_w1534_,
		_w2740_,
		_w2742_
	);
	LUT3 #(
		.INIT('h13)
	) name1562 (
		_w1602_,
		_w2741_,
		_w2742_,
		_w2743_
	);
	LUT2 #(
		.INIT('h4)
	) name1563 (
		\g1088_reg/NET0131 ,
		\g915_reg/NET0131 ,
		_w2744_
	);
	LUT2 #(
		.INIT('h2)
	) name1564 (
		_w1900_,
		_w2342_,
		_w2745_
	);
	LUT4 #(
		.INIT('h0400)
	) name1565 (
		_w1849_,
		_w1850_,
		_w1898_,
		_w1899_,
		_w2746_
	);
	LUT3 #(
		.INIT('h40)
	) name1566 (
		_w1950_,
		_w2347_,
		_w2746_,
		_w2747_
	);
	LUT4 #(
		.INIT('h000b)
	) name1567 (
		_w2350_,
		_w2398_,
		_w2745_,
		_w2747_,
		_w2748_
	);
	LUT2 #(
		.INIT('h1)
	) name1568 (
		\g1088_reg/NET0131 ,
		\g915_reg/NET0131 ,
		_w2749_
	);
	LUT3 #(
		.INIT('h15)
	) name1569 (
		_w1929_,
		_w2406_,
		_w2412_,
		_w2750_
	);
	LUT3 #(
		.INIT('h80)
	) name1570 (
		_w1929_,
		_w2410_,
		_w2411_,
		_w2751_
	);
	LUT3 #(
		.INIT('h15)
	) name1571 (
		_w2365_,
		_w2406_,
		_w2751_,
		_w2752_
	);
	LUT3 #(
		.INIT('h20)
	) name1572 (
		_w2342_,
		_w2750_,
		_w2752_,
		_w2753_
	);
	LUT3 #(
		.INIT('h23)
	) name1573 (
		_w2350_,
		_w2749_,
		_w2753_,
		_w2754_
	);
	LUT3 #(
		.INIT('hea)
	) name1574 (
		_w2744_,
		_w2748_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h4)
	) name1575 (
		\g7961_pad ,
		\g909_reg/NET0131 ,
		_w2756_
	);
	LUT2 #(
		.INIT('h1)
	) name1576 (
		\g7961_pad ,
		\g909_reg/NET0131 ,
		_w2757_
	);
	LUT3 #(
		.INIT('h0b)
	) name1577 (
		_w2350_,
		_w2753_,
		_w2757_,
		_w2758_
	);
	LUT3 #(
		.INIT('hec)
	) name1578 (
		_w2748_,
		_w2756_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h4)
	) name1579 (
		\g1092_reg/NET0131 ,
		\g912_reg/NET0131 ,
		_w2760_
	);
	LUT2 #(
		.INIT('h1)
	) name1580 (
		\g1092_reg/NET0131 ,
		\g912_reg/NET0131 ,
		_w2761_
	);
	LUT3 #(
		.INIT('h0b)
	) name1581 (
		_w2350_,
		_w2753_,
		_w2761_,
		_w2762_
	);
	LUT3 #(
		.INIT('hec)
	) name1582 (
		_w2748_,
		_w2760_,
		_w2762_,
		_w2763_
	);
	LUT2 #(
		.INIT('h2)
	) name1583 (
		\g222_reg/NET0131 ,
		\g7961_pad ,
		_w2764_
	);
	LUT3 #(
		.INIT('h2a)
	) name1584 (
		_w1740_,
		_w2295_,
		_w2304_,
		_w2765_
	);
	LUT3 #(
		.INIT('h80)
	) name1585 (
		_w1711_,
		_w1740_,
		_w2310_,
		_w2766_
	);
	LUT3 #(
		.INIT('hd0)
	) name1586 (
		_w1737_,
		_w2306_,
		_w2766_,
		_w2767_
	);
	LUT4 #(
		.INIT('h000b)
	) name1587 (
		_w2314_,
		_w2702_,
		_w2765_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h1)
	) name1588 (
		\g222_reg/NET0131 ,
		\g7961_pad ,
		_w2769_
	);
	LUT3 #(
		.INIT('h9c)
	) name1589 (
		_w1697_,
		_w1761_,
		_w1821_,
		_w2770_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name1590 (
		_w1765_,
		_w2710_,
		_w2712_,
		_w2770_,
		_w2771_
	);
	LUT3 #(
		.INIT('h80)
	) name1591 (
		_w2295_,
		_w2641_,
		_w2771_,
		_w2772_
	);
	LUT3 #(
		.INIT('h23)
	) name1592 (
		_w2314_,
		_w2769_,
		_w2772_,
		_w2773_
	);
	LUT3 #(
		.INIT('hea)
	) name1593 (
		_w2764_,
		_w2768_,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h4)
	) name1594 (
		\g1092_reg/NET0131 ,
		\g225_reg/NET0131 ,
		_w2775_
	);
	LUT2 #(
		.INIT('h1)
	) name1595 (
		\g1092_reg/NET0131 ,
		\g225_reg/NET0131 ,
		_w2776_
	);
	LUT3 #(
		.INIT('h0b)
	) name1596 (
		_w2314_,
		_w2772_,
		_w2776_,
		_w2777_
	);
	LUT3 #(
		.INIT('hec)
	) name1597 (
		_w2768_,
		_w2775_,
		_w2777_,
		_w2778_
	);
	LUT2 #(
		.INIT('h4)
	) name1598 (
		\g1088_reg/NET0131 ,
		\g228_reg/NET0131 ,
		_w2779_
	);
	LUT2 #(
		.INIT('h1)
	) name1599 (
		\g1088_reg/NET0131 ,
		\g228_reg/NET0131 ,
		_w2780_
	);
	LUT3 #(
		.INIT('h0b)
	) name1600 (
		_w2314_,
		_w2772_,
		_w2780_,
		_w2781_
	);
	LUT3 #(
		.INIT('hec)
	) name1601 (
		_w2768_,
		_w2779_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h1)
	) name1602 (
		\g2297_reg/NET0131 ,
		\g7961_pad ,
		_w2783_
	);
	LUT2 #(
		.INIT('h2)
	) name1603 (
		\g2297_reg/NET0131 ,
		\g7961_pad ,
		_w2784_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1604 (
		_w1297_,
		_w1368_,
		_w1369_,
		_w2482_,
		_w2785_
	);
	LUT4 #(
		.INIT('h2000)
	) name1605 (
		_w1297_,
		_w1368_,
		_w1369_,
		_w2586_,
		_w2786_
	);
	LUT3 #(
		.INIT('ha8)
	) name1606 (
		_w2585_,
		_w2785_,
		_w2786_,
		_w2787_
	);
	LUT4 #(
		.INIT('h22ea)
	) name1607 (
		_w1297_,
		_w2584_,
		_w2588_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h8)
	) name1608 (
		_w2498_,
		_w2788_,
		_w2789_
	);
	LUT3 #(
		.INIT('h23)
	) name1609 (
		_w2473_,
		_w2494_,
		_w2789_,
		_w2790_
	);
	LUT3 #(
		.INIT('h8a)
	) name1610 (
		_w1294_,
		_w2477_,
		_w2480_,
		_w2791_
	);
	LUT2 #(
		.INIT('h8)
	) name1611 (
		_w1294_,
		_w2472_,
		_w2792_
	);
	LUT4 #(
		.INIT('h020f)
	) name1612 (
		_w1333_,
		_w2466_,
		_w2791_,
		_w2792_,
		_w2793_
	);
	LUT2 #(
		.INIT('h4)
	) name1613 (
		_w2783_,
		_w2793_,
		_w2794_
	);
	LUT3 #(
		.INIT('hea)
	) name1614 (
		_w2784_,
		_w2790_,
		_w2794_,
		_w2795_
	);
	LUT2 #(
		.INIT('h1)
	) name1615 (
		\g1092_reg/NET0131 ,
		\g2300_reg/NET0131 ,
		_w2796_
	);
	LUT2 #(
		.INIT('h4)
	) name1616 (
		\g1092_reg/NET0131 ,
		\g2300_reg/NET0131 ,
		_w2797_
	);
	LUT2 #(
		.INIT('h2)
	) name1617 (
		_w2793_,
		_w2796_,
		_w2798_
	);
	LUT3 #(
		.INIT('hec)
	) name1618 (
		_w2790_,
		_w2797_,
		_w2798_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name1619 (
		\g1088_reg/NET0131 ,
		\g2303_reg/NET0131 ,
		_w2800_
	);
	LUT2 #(
		.INIT('h4)
	) name1620 (
		\g1088_reg/NET0131 ,
		\g2303_reg/NET0131 ,
		_w2801_
	);
	LUT2 #(
		.INIT('h2)
	) name1621 (
		_w2793_,
		_w2800_,
		_w2802_
	);
	LUT3 #(
		.INIT('hec)
	) name1622 (
		_w2790_,
		_w2801_,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h2)
	) name1623 (
		\g1603_reg/NET0131 ,
		\g7961_pad ,
		_w2804_
	);
	LUT3 #(
		.INIT('h0d)
	) name1624 (
		_w2013_,
		_w2459_,
		_w2672_,
		_w2805_
	);
	LUT2 #(
		.INIT('h1)
	) name1625 (
		\g1603_reg/NET0131 ,
		\g7961_pad ,
		_w2806_
	);
	LUT4 #(
		.INIT('h1555)
	) name1626 (
		_w2016_,
		_w2678_,
		_w2685_,
		_w2686_,
		_w2807_
	);
	LUT4 #(
		.INIT('h8288)
	) name1627 (
		_w2016_,
		_w2093_,
		_w2129_,
		_w2143_,
		_w2808_
	);
	LUT4 #(
		.INIT('h1555)
	) name1628 (
		_w2453_,
		_w2678_,
		_w2685_,
		_w2808_,
		_w2809_
	);
	LUT3 #(
		.INIT('h20)
	) name1629 (
		_w2439_,
		_w2807_,
		_w2809_,
		_w2810_
	);
	LUT3 #(
		.INIT('h23)
	) name1630 (
		_w2434_,
		_w2806_,
		_w2810_,
		_w2811_
	);
	LUT3 #(
		.INIT('hea)
	) name1631 (
		_w2804_,
		_w2805_,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h4)
	) name1632 (
		\g1092_reg/NET0131 ,
		\g1606_reg/NET0131 ,
		_w2813_
	);
	LUT2 #(
		.INIT('h1)
	) name1633 (
		\g1092_reg/NET0131 ,
		\g1606_reg/NET0131 ,
		_w2814_
	);
	LUT3 #(
		.INIT('h0b)
	) name1634 (
		_w2434_,
		_w2810_,
		_w2814_,
		_w2815_
	);
	LUT3 #(
		.INIT('hec)
	) name1635 (
		_w2805_,
		_w2813_,
		_w2815_,
		_w2816_
	);
	LUT2 #(
		.INIT('h4)
	) name1636 (
		\g1088_reg/NET0131 ,
		\g1609_reg/NET0131 ,
		_w2817_
	);
	LUT2 #(
		.INIT('h1)
	) name1637 (
		\g1088_reg/NET0131 ,
		\g1609_reg/NET0131 ,
		_w2818_
	);
	LUT3 #(
		.INIT('h0b)
	) name1638 (
		_w2434_,
		_w2810_,
		_w2818_,
		_w2819_
	);
	LUT3 #(
		.INIT('hec)
	) name1639 (
		_w2805_,
		_w2817_,
		_w2819_,
		_w2820_
	);
	LUT4 #(
		.INIT('h0002)
	) name1640 (
		\g499_reg/NET0131 ,
		\g544_reg/NET0131 ,
		\g559_reg/NET0131 ,
		\g563_pad ,
		_w2821_
	);
	LUT2 #(
		.INIT('h2)
	) name1641 (
		\g5657_pad ,
		\g705_reg/NET0131 ,
		_w2822_
	);
	LUT4 #(
		.INIT('hf351)
	) name1642 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g704_reg/NET0131 ,
		\g706_reg/NET0131 ,
		_w2823_
	);
	LUT2 #(
		.INIT('h4)
	) name1643 (
		_w2822_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h2)
	) name1644 (
		\g5657_pad ,
		\g714_reg/NET0131 ,
		_w2825_
	);
	LUT4 #(
		.INIT('hf351)
	) name1645 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g713_reg/NET0131 ,
		\g715_reg/NET0131 ,
		_w2826_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1646 (
		_w2822_,
		_w2823_,
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h2)
	) name1647 (
		\g5657_pad ,
		\g720_reg/NET0131 ,
		_w2828_
	);
	LUT4 #(
		.INIT('hf351)
	) name1648 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g719_reg/NET0131 ,
		\g721_reg/NET0131 ,
		_w2829_
	);
	LUT2 #(
		.INIT('h2)
	) name1649 (
		\g5657_pad ,
		\g738_reg/NET0131 ,
		_w2830_
	);
	LUT4 #(
		.INIT('hf351)
	) name1650 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g737_reg/NET0131 ,
		\g739_reg/NET0131 ,
		_w2831_
	);
	LUT4 #(
		.INIT('h4044)
	) name1651 (
		_w2828_,
		_w2829_,
		_w2830_,
		_w2831_,
		_w2832_
	);
	LUT2 #(
		.INIT('h8)
	) name1652 (
		_w2827_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h2)
	) name1653 (
		\g5657_pad ,
		\g723_reg/NET0131 ,
		_w2834_
	);
	LUT4 #(
		.INIT('hf351)
	) name1654 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g722_reg/NET0131 ,
		\g724_reg/NET0131 ,
		_w2835_
	);
	LUT2 #(
		.INIT('h4)
	) name1655 (
		_w2834_,
		_w2835_,
		_w2836_
	);
	LUT2 #(
		.INIT('h2)
	) name1656 (
		\g5657_pad ,
		\g702_reg/NET0131 ,
		_w2837_
	);
	LUT4 #(
		.INIT('hf351)
	) name1657 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g701_reg/NET0131 ,
		\g703_reg/NET0131 ,
		_w2838_
	);
	LUT2 #(
		.INIT('h4)
	) name1658 (
		_w2837_,
		_w2838_,
		_w2839_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1659 (
		_w2834_,
		_w2835_,
		_w2837_,
		_w2838_,
		_w2840_
	);
	LUT2 #(
		.INIT('h2)
	) name1660 (
		\g5657_pad ,
		\g708_reg/NET0131 ,
		_w2841_
	);
	LUT4 #(
		.INIT('hf351)
	) name1661 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g707_reg/NET0131 ,
		\g709_reg/NET0131 ,
		_w2842_
	);
	LUT2 #(
		.INIT('h4)
	) name1662 (
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h2)
	) name1663 (
		\g5657_pad ,
		\g699_reg/NET0131 ,
		_w2844_
	);
	LUT4 #(
		.INIT('hf351)
	) name1664 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g698_reg/NET0131 ,
		\g700_reg/NET0131 ,
		_w2845_
	);
	LUT4 #(
		.INIT('h0b00)
	) name1665 (
		_w2841_,
		_w2842_,
		_w2844_,
		_w2845_,
		_w2846_
	);
	LUT2 #(
		.INIT('h2)
	) name1666 (
		\g5657_pad ,
		\g726_reg/NET0131 ,
		_w2847_
	);
	LUT4 #(
		.INIT('hf351)
	) name1667 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g725_reg/NET0131 ,
		\g727_reg/NET0131 ,
		_w2848_
	);
	LUT2 #(
		.INIT('h4)
	) name1668 (
		_w2847_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name1669 (
		\g1024_reg/NET0131 ,
		\g731_reg/NET0131 ,
		_w2850_
	);
	LUT4 #(
		.INIT('hf351)
	) name1670 (
		\g1018_reg/NET0131 ,
		\g5657_pad ,
		\g732_reg/NET0131 ,
		\g733_reg/NET0131 ,
		_w2851_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name1671 (
		_w2847_,
		_w2848_,
		_w2850_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h2)
	) name1672 (
		\g5657_pad ,
		\g711_reg/NET0131 ,
		_w2853_
	);
	LUT4 #(
		.INIT('hf351)
	) name1673 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g710_reg/NET0131 ,
		\g712_reg/NET0131 ,
		_w2854_
	);
	LUT2 #(
		.INIT('h2)
	) name1674 (
		\g5657_pad ,
		\g717_reg/NET0131 ,
		_w2855_
	);
	LUT4 #(
		.INIT('hf351)
	) name1675 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g716_reg/NET0131 ,
		\g718_reg/NET0131 ,
		_w2856_
	);
	LUT4 #(
		.INIT('h0400)
	) name1676 (
		_w2853_,
		_w2854_,
		_w2855_,
		_w2856_,
		_w2857_
	);
	LUT4 #(
		.INIT('h8000)
	) name1677 (
		_w2840_,
		_w2846_,
		_w2852_,
		_w2857_,
		_w2858_
	);
	LUT2 #(
		.INIT('h8)
	) name1678 (
		\g1024_reg/NET0131 ,
		\g611_reg/NET0131 ,
		_w2859_
	);
	LUT4 #(
		.INIT('h153f)
	) name1679 (
		\g1018_reg/NET0131 ,
		\g5657_pad ,
		\g605_reg/NET0131 ,
		\g608_reg/NET0131 ,
		_w2860_
	);
	LUT2 #(
		.INIT('h4)
	) name1680 (
		_w2859_,
		_w2860_,
		_w2861_
	);
	LUT4 #(
		.INIT('hec13)
	) name1681 (
		_w2833_,
		_w2843_,
		_w2858_,
		_w2861_,
		_w2862_
	);
	LUT2 #(
		.INIT('h8)
	) name1682 (
		\g1018_reg/NET0131 ,
		\g617_reg/NET0131 ,
		_w2863_
	);
	LUT4 #(
		.INIT('h153f)
	) name1683 (
		\g1024_reg/NET0131 ,
		\g5657_pad ,
		\g614_reg/NET0131 ,
		\g620_reg/NET0131 ,
		_w2864_
	);
	LUT2 #(
		.INIT('h4)
	) name1684 (
		_w2863_,
		_w2864_,
		_w2865_
	);
	LUT4 #(
		.INIT('hea15)
	) name1685 (
		_w2824_,
		_w2833_,
		_w2858_,
		_w2865_,
		_w2866_
	);
	LUT3 #(
		.INIT('hd7)
	) name1686 (
		_w2821_,
		_w2862_,
		_w2866_,
		_w2867_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1687 (
		_w2844_,
		_w2845_,
		_w2863_,
		_w2864_,
		_w2868_
	);
	LUT2 #(
		.INIT('h2)
	) name1688 (
		_w2821_,
		_w2868_,
		_w2869_
	);
	LUT4 #(
		.INIT('hec13)
	) name1689 (
		_w2833_,
		_w2839_,
		_w2858_,
		_w2861_,
		_w2870_
	);
	LUT2 #(
		.INIT('h8)
	) name1690 (
		_w2821_,
		_w2868_,
		_w2871_
	);
	LUT3 #(
		.INIT('h7d)
	) name1691 (
		_w2821_,
		_w2868_,
		_w2870_,
		_w2872_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1692 (
		_w2853_,
		_w2854_,
		_w2863_,
		_w2864_,
		_w2873_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1693 (
		_w2825_,
		_w2826_,
		_w2859_,
		_w2860_,
		_w2874_
	);
	LUT3 #(
		.INIT('hd7)
	) name1694 (
		_w2821_,
		_w2873_,
		_w2874_,
		_w2875_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1695 (
		_w2828_,
		_w2829_,
		_w2859_,
		_w2860_,
		_w2876_
	);
	LUT4 #(
		.INIT('h4b44)
	) name1696 (
		_w2855_,
		_w2856_,
		_w2863_,
		_w2864_,
		_w2877_
	);
	LUT3 #(
		.INIT('hd7)
	) name1697 (
		_w2821_,
		_w2876_,
		_w2877_,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name1698 (
		_w2875_,
		_w2878_,
		_w2879_
	);
	LUT4 #(
		.INIT('he200)
	) name1699 (
		_w2869_,
		_w2870_,
		_w2871_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h4)
	) name1700 (
		_w2875_,
		_w2878_,
		_w2881_
	);
	LUT4 #(
		.INIT('he200)
	) name1701 (
		_w2869_,
		_w2870_,
		_w2871_,
		_w2881_,
		_w2882_
	);
	LUT3 #(
		.INIT('h1b)
	) name1702 (
		_w2867_,
		_w2880_,
		_w2882_,
		_w2883_
	);
	LUT4 #(
		.INIT('hd7ff)
	) name1703 (
		_w2821_,
		_w2862_,
		_w2866_,
		_w2881_,
		_w2884_
	);
	LUT4 #(
		.INIT('h7f33)
	) name1704 (
		_w2867_,
		_w2872_,
		_w2879_,
		_w2884_,
		_w2885_
	);
	LUT2 #(
		.INIT('h8)
	) name1705 (
		_w2883_,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h8)
	) name1706 (
		_w2875_,
		_w2878_,
		_w2887_
	);
	LUT4 #(
		.INIT('he200)
	) name1707 (
		_w2869_,
		_w2870_,
		_w2871_,
		_w2887_,
		_w2888_
	);
	LUT2 #(
		.INIT('h2)
	) name1708 (
		_w2875_,
		_w2878_,
		_w2889_
	);
	LUT4 #(
		.INIT('he200)
	) name1709 (
		_w2869_,
		_w2870_,
		_w2871_,
		_w2889_,
		_w2890_
	);
	LUT3 #(
		.INIT('h1b)
	) name1710 (
		_w2867_,
		_w2888_,
		_w2890_,
		_w2891_
	);
	LUT4 #(
		.INIT('hd7ff)
	) name1711 (
		_w2821_,
		_w2862_,
		_w2866_,
		_w2889_,
		_w2892_
	);
	LUT4 #(
		.INIT('h7f33)
	) name1712 (
		_w2867_,
		_w2872_,
		_w2887_,
		_w2892_,
		_w2893_
	);
	LUT3 #(
		.INIT('h80)
	) name1713 (
		\g1196_reg/NET0131 ,
		_w2891_,
		_w2893_,
		_w2894_
	);
	LUT4 #(
		.INIT('hec13)
	) name1714 (
		_w2833_,
		_w2836_,
		_w2858_,
		_w2865_,
		_w2895_
	);
	LUT4 #(
		.INIT('hec13)
	) name1715 (
		_w2833_,
		_w2849_,
		_w2858_,
		_w2861_,
		_w2896_
	);
	LUT2 #(
		.INIT('h8)
	) name1716 (
		\g1243_reg/NET0131 ,
		_w2821_,
		_w2897_
	);
	LUT3 #(
		.INIT('h04)
	) name1717 (
		\g499_reg/NET0131 ,
		\g548_reg/NET0131 ,
		\g5657_pad ,
		_w2898_
	);
	LUT4 #(
		.INIT('h0007)
	) name1718 (
		\g499_reg/NET0131 ,
		\g544_reg/NET0131 ,
		\g559_reg/NET0131 ,
		\g563_pad ,
		_w2899_
	);
	LUT2 #(
		.INIT('h4)
	) name1719 (
		_w2898_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('h4)
	) name1720 (
		\g499_reg/NET0131 ,
		\g5657_pad ,
		_w2901_
	);
	LUT3 #(
		.INIT('h04)
	) name1721 (
		_w2898_,
		_w2899_,
		_w2901_,
		_w2902_
	);
	LUT3 #(
		.INIT('h10)
	) name1722 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g525_reg/NET0131 ,
		_w2903_
	);
	LUT3 #(
		.INIT('hd8)
	) name1723 (
		\g3229_pad ,
		\g538_reg/NET0131 ,
		\g541_reg/NET0131 ,
		_w2904_
	);
	LUT2 #(
		.INIT('h8)
	) name1724 (
		_w2903_,
		_w2904_,
		_w2905_
	);
	LUT2 #(
		.INIT('h8)
	) name1725 (
		_w2902_,
		_w2905_,
		_w2906_
	);
	LUT4 #(
		.INIT('h009f)
	) name1726 (
		_w2895_,
		_w2896_,
		_w2897_,
		_w2906_,
		_w2907_
	);
	LUT3 #(
		.INIT('h8f)
	) name1727 (
		_w2886_,
		_w2894_,
		_w2907_,
		_w2908_
	);
	LUT4 #(
		.INIT('h0c5c)
	) name1728 (
		\g1092_reg/NET0131 ,
		\g1679_reg/NET0131 ,
		\g1680_reg/NET0131 ,
		\g1686_reg/NET0131 ,
		_w2909_
	);
	LUT4 #(
		.INIT('h4500)
	) name1729 (
		_w1684_,
		_w1687_,
		_w1688_,
		_w1690_,
		_w2910_
	);
	LUT2 #(
		.INIT('h1)
	) name1730 (
		_w2909_,
		_w2910_,
		_w2911_
	);
	LUT3 #(
		.INIT('h10)
	) name1731 (
		\g1563_reg/NET0131 ,
		_w1745_,
		_w1746_,
		_w2912_
	);
	LUT3 #(
		.INIT('h8a)
	) name1732 (
		\g1563_reg/NET0131 ,
		\g315_reg/NET0131 ,
		\g7961_pad ,
		_w2913_
	);
	LUT4 #(
		.INIT('h8a00)
	) name1733 (
		_w1696_,
		_w1734_,
		_w1735_,
		_w2913_,
		_w2914_
	);
	LUT2 #(
		.INIT('h8)
	) name1734 (
		_w1747_,
		_w2914_,
		_w2915_
	);
	LUT3 #(
		.INIT('h23)
	) name1735 (
		_w2306_,
		_w2912_,
		_w2915_,
		_w2916_
	);
	LUT4 #(
		.INIT('h2aaa)
	) name1736 (
		_w1737_,
		_w1771_,
		_w1780_,
		_w1797_,
		_w2917_
	);
	LUT2 #(
		.INIT('h4)
	) name1737 (
		_w1697_,
		_w2917_,
		_w2918_
	);
	LUT3 #(
		.INIT('h04)
	) name1738 (
		_w1697_,
		_w1737_,
		_w1747_,
		_w2919_
	);
	LUT3 #(
		.INIT('h23)
	) name1739 (
		_w2306_,
		_w2918_,
		_w2919_,
		_w2920_
	);
	LUT2 #(
		.INIT('h1)
	) name1740 (
		_w1700_,
		_w1830_,
		_w2921_
	);
	LUT3 #(
		.INIT('h70)
	) name1741 (
		_w2916_,
		_w2920_,
		_w2921_,
		_w2922_
	);
	LUT2 #(
		.INIT('h8)
	) name1742 (
		_w1333_,
		_w1368_,
		_w2923_
	);
	LUT3 #(
		.INIT('ha8)
	) name1743 (
		\g1563_reg/NET0131 ,
		_w1313_,
		_w1368_,
		_w2924_
	);
	LUT4 #(
		.INIT('h8000)
	) name1744 (
		\g1563_reg/NET0131 ,
		_w1287_,
		_w1299_,
		_w1308_,
		_w2925_
	);
	LUT2 #(
		.INIT('h1)
	) name1745 (
		_w2924_,
		_w2925_,
		_w2926_
	);
	LUT3 #(
		.INIT('h51)
	) name1746 (
		_w1253_,
		_w1333_,
		_w1368_,
		_w2927_
	);
	LUT4 #(
		.INIT('h4000)
	) name1747 (
		_w1253_,
		_w1287_,
		_w1299_,
		_w1308_,
		_w2928_
	);
	LUT4 #(
		.INIT('h070f)
	) name1748 (
		_w1326_,
		_w1337_,
		_w1364_,
		_w1374_,
		_w2929_
	);
	LUT3 #(
		.INIT('h10)
	) name1749 (
		_w2927_,
		_w2928_,
		_w2929_,
		_w2930_
	);
	LUT4 #(
		.INIT('hf400)
	) name1750 (
		_w2466_,
		_w2923_,
		_w2926_,
		_w2930_,
		_w2931_
	);
	LUT3 #(
		.INIT('h10)
	) name1751 (
		\g1563_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w2932_
	);
	LUT2 #(
		.INIT('h1)
	) name1752 (
		_w1975_,
		_w1978_,
		_w2933_
	);
	LUT4 #(
		.INIT('h0400)
	) name1753 (
		_w1846_,
		_w1847_,
		_w1849_,
		_w1850_,
		_w2934_
	);
	LUT4 #(
		.INIT('h1033)
	) name1754 (
		_w1950_,
		_w2932_,
		_w2933_,
		_w2934_,
		_w2935_
	);
	LUT2 #(
		.INIT('h4)
	) name1755 (
		_w1848_,
		_w1891_,
		_w2936_
	);
	LUT4 #(
		.INIT('h7f00)
	) name1756 (
		_w1947_,
		_w1982_,
		_w1983_,
		_w2936_,
		_w2937_
	);
	LUT2 #(
		.INIT('h1)
	) name1757 (
		_w1859_,
		_w1918_,
		_w2938_
	);
	LUT3 #(
		.INIT('hd0)
	) name1758 (
		_w2935_,
		_w2937_,
		_w2938_,
		_w2939_
	);
	LUT3 #(
		.INIT('h8a)
	) name1759 (
		\g1563_reg/NET0131 ,
		\g1696_reg/NET0131 ,
		\g7961_pad ,
		_w2940_
	);
	LUT4 #(
		.INIT('hb000)
	) name1760 (
		_w2007_,
		_w2008_,
		_w2128_,
		_w2940_,
		_w2941_
	);
	LUT3 #(
		.INIT('hb0)
	) name1761 (
		_w2105_,
		_w2109_,
		_w2941_,
		_w2942_
	);
	LUT3 #(
		.INIT('hb0)
	) name1762 (
		_w2035_,
		_w2040_,
		_w2941_,
		_w2943_
	);
	LUT3 #(
		.INIT('ha8)
	) name1763 (
		\g1563_reg/NET0131 ,
		_w2009_,
		_w2129_,
		_w2944_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		_w2117_,
		_w2944_,
		_w2945_
	);
	LUT3 #(
		.INIT('h31)
	) name1765 (
		_w2010_,
		_w2113_,
		_w2129_,
		_w2946_
	);
	LUT4 #(
		.INIT('h2000)
	) name1766 (
		_w2107_,
		_w2113_,
		_w2115_,
		_w2116_,
		_w2947_
	);
	LUT3 #(
		.INIT('h02)
	) name1767 (
		_w2142_,
		_w2946_,
		_w2947_,
		_w2948_
	);
	LUT4 #(
		.INIT('hfe00)
	) name1768 (
		_w2942_,
		_w2943_,
		_w2945_,
		_w2948_,
		_w2949_
	);
	LUT2 #(
		.INIT('h8)
	) name1769 (
		\g2580_reg/NET0131 ,
		\g2581_reg/NET0131 ,
		_w2950_
	);
	LUT2 #(
		.INIT('h2)
	) name1770 (
		\g1192_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		_w2951_
	);
	LUT3 #(
		.INIT('h08)
	) name1771 (
		\g1018_reg/NET0131 ,
		\g1192_reg/NET0131 ,
		\g1193_reg/NET0131 ,
		_w2952_
	);
	LUT4 #(
		.INIT('h0020)
	) name1772 (
		\g1018_reg/NET0131 ,
		\g1192_reg/NET0131 ,
		\g506_reg/NET0131 ,
		\g507_reg/NET0131 ,
		_w2953_
	);
	LUT3 #(
		.INIT('h0e)
	) name1773 (
		\g1018_reg/NET0131 ,
		\g16399_pad ,
		\g1886_reg/NET0131 ,
		_w2954_
	);
	LUT2 #(
		.INIT('h8)
	) name1774 (
		\g1886_reg/NET0131 ,
		\g1887_reg/NET0131 ,
		_w2955_
	);
	LUT3 #(
		.INIT('h2a)
	) name1775 (
		\g1018_reg/NET0131 ,
		\g1886_reg/NET0131 ,
		\g1887_reg/NET0131 ,
		_w2956_
	);
	LUT4 #(
		.INIT('hef00)
	) name1776 (
		_w2952_,
		_w2953_,
		_w2954_,
		_w2956_,
		_w2957_
	);
	LUT3 #(
		.INIT('h0e)
	) name1777 (
		\g1018_reg/NET0131 ,
		\g16437_pad ,
		\g2580_reg/NET0131 ,
		_w2958_
	);
	LUT3 #(
		.INIT('hba)
	) name1778 (
		_w2950_,
		_w2957_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h2)
	) name1779 (
		\g805_reg/NET0131 ,
		_w2342_,
		_w2960_
	);
	LUT3 #(
		.INIT('h20)
	) name1780 (
		\g805_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w2961_
	);
	LUT3 #(
		.INIT('h40)
	) name1781 (
		_w1950_,
		_w2347_,
		_w2961_,
		_w2962_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name1782 (
		_w1972_,
		_w2366_,
		_w2389_,
		_w2405_,
		_w2963_
	);
	LUT2 #(
		.INIT('h1)
	) name1783 (
		_w2365_,
		_w2963_,
		_w2964_
	);
	LUT2 #(
		.INIT('h8)
	) name1784 (
		_w2342_,
		_w2964_,
		_w2965_
	);
	LUT4 #(
		.INIT('hfdfc)
	) name1785 (
		_w2350_,
		_w2960_,
		_w2962_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h1)
	) name1786 (
		\g117_reg/NET0131 ,
		_w2315_,
		_w2967_
	);
	LUT3 #(
		.INIT('h40)
	) name1787 (
		\g117_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w2968_
	);
	LUT3 #(
		.INIT('hd0)
	) name1788 (
		_w1737_,
		_w2306_,
		_w2968_,
		_w2969_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name1789 (
		_w1774_,
		_w2329_,
		_w2651_,
		_w2709_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name1790 (
		_w2328_,
		_w2970_,
		_w2971_
	);
	LUT2 #(
		.INIT('h2)
	) name1791 (
		_w2315_,
		_w2971_,
		_w2972_
	);
	LUT4 #(
		.INIT('h0203)
	) name1792 (
		_w2314_,
		_w2967_,
		_w2969_,
		_w2972_,
		_w2973_
	);
	LUT3 #(
		.INIT('h80)
	) name1793 (
		_w2169_,
		_w2174_,
		_w2180_,
		_w2974_
	);
	LUT2 #(
		.INIT('h2)
	) name1794 (
		\g1018_reg/NET0131 ,
		\g1422_reg/NET0131 ,
		_w2975_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name1795 (
		\g1024_reg/NET0131 ,
		\g1420_reg/NET0131 ,
		\g1421_reg/NET0131 ,
		\g5657_pad ,
		_w2976_
	);
	LUT3 #(
		.INIT('h8a)
	) name1796 (
		_w2168_,
		_w2975_,
		_w2976_,
		_w2977_
	);
	LUT3 #(
		.INIT('h8a)
	) name1797 (
		_w1613_,
		_w2166_,
		_w2977_,
		_w2978_
	);
	LUT3 #(
		.INIT('h70)
	) name1798 (
		_w2205_,
		_w2974_,
		_w2978_,
		_w2979_
	);
	LUT3 #(
		.INIT('h54)
	) name1799 (
		\g1196_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w2980_
	);
	LUT2 #(
		.INIT('h2)
	) name1800 (
		_w2168_,
		_w2980_,
		_w2981_
	);
	LUT3 #(
		.INIT('h10)
	) name1801 (
		_w2166_,
		_w2224_,
		_w2981_,
		_w2982_
	);
	LUT2 #(
		.INIT('h1)
	) name1802 (
		\g1196_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		_w2983_
	);
	LUT3 #(
		.INIT('h01)
	) name1803 (
		\g1215_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w2984_
	);
	LUT3 #(
		.INIT('h13)
	) name1804 (
		_w2980_,
		_w2983_,
		_w2984_,
		_w2985_
	);
	LUT4 #(
		.INIT('hfc54)
	) name1805 (
		\g1186_reg/NET0131 ,
		\g1196_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		_w2986_
	);
	LUT3 #(
		.INIT('hd0)
	) name1806 (
		_w2164_,
		_w2165_,
		_w2986_,
		_w2987_
	);
	LUT3 #(
		.INIT('h54)
	) name1807 (
		\g1243_reg/NET0131 ,
		_w2985_,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h4)
	) name1808 (
		_w2982_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('he)
	) name1809 (
		_w2979_,
		_w2989_,
		_w2990_
	);
	LUT3 #(
		.INIT('h80)
	) name1810 (
		\g1186_reg/NET0131 ,
		_w2174_,
		_w2180_,
		_w2991_
	);
	LUT4 #(
		.INIT('hae00)
	) name1811 (
		_w1508_,
		_w2164_,
		_w2165_,
		_w2167_,
		_w2992_
	);
	LUT3 #(
		.INIT('h8a)
	) name1812 (
		\g1186_reg/NET0131 ,
		_w2975_,
		_w2976_,
		_w2993_
	);
	LUT2 #(
		.INIT('h2)
	) name1813 (
		_w2992_,
		_w2993_,
		_w2994_
	);
	LUT4 #(
		.INIT('h80aa)
	) name1814 (
		_w1613_,
		_w2205_,
		_w2991_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h2)
	) name1815 (
		_w2168_,
		_w2233_,
		_w2996_
	);
	LUT3 #(
		.INIT('h10)
	) name1816 (
		_w2166_,
		_w2226_,
		_w2996_,
		_w2997_
	);
	LUT3 #(
		.INIT('h01)
	) name1817 (
		\g1217_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w2998_
	);
	LUT3 #(
		.INIT('h13)
	) name1818 (
		_w2980_,
		_w2983_,
		_w2998_,
		_w2999_
	);
	LUT3 #(
		.INIT('h54)
	) name1819 (
		\g1243_reg/NET0131 ,
		_w2987_,
		_w2999_,
		_w3000_
	);
	LUT2 #(
		.INIT('h4)
	) name1820 (
		_w2997_,
		_w3000_,
		_w3001_
	);
	LUT2 #(
		.INIT('he)
	) name1821 (
		_w2995_,
		_w3001_,
		_w3002_
	);
	LUT3 #(
		.INIT('h10)
	) name1822 (
		_w2166_,
		_w2227_,
		_w2996_,
		_w3003_
	);
	LUT3 #(
		.INIT('h01)
	) name1823 (
		\g1218_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w3004_
	);
	LUT3 #(
		.INIT('h13)
	) name1824 (
		_w2980_,
		_w2983_,
		_w3004_,
		_w3005_
	);
	LUT3 #(
		.INIT('h54)
	) name1825 (
		\g1243_reg/NET0131 ,
		_w2987_,
		_w3005_,
		_w3006_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		_w3003_,
		_w3006_,
		_w3007_
	);
	LUT2 #(
		.INIT('he)
	) name1827 (
		_w2979_,
		_w3007_,
		_w3008_
	);
	LUT4 #(
		.INIT('h4440)
	) name1828 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w3009_
	);
	LUT4 #(
		.INIT('h3100)
	) name1829 (
		\g1186_reg/NET0131 ,
		\g1196_reg/NET0131 ,
		\g1230_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w3010_
	);
	LUT4 #(
		.INIT('h020f)
	) name1830 (
		_w2164_,
		_w2165_,
		_w3009_,
		_w3010_,
		_w3011_
	);
	LUT3 #(
		.INIT('h0e)
	) name1831 (
		\g1196_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w3012_
	);
	LUT3 #(
		.INIT('h01)
	) name1832 (
		\g1219_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w3013_
	);
	LUT3 #(
		.INIT('h4c)
	) name1833 (
		_w2980_,
		_w3012_,
		_w3013_,
		_w3014_
	);
	LUT4 #(
		.INIT('h5100)
	) name1834 (
		_w1508_,
		_w2164_,
		_w2165_,
		_w3012_,
		_w3015_
	);
	LUT3 #(
		.INIT('h02)
	) name1835 (
		_w3011_,
		_w3014_,
		_w3015_,
		_w3016_
	);
	LUT3 #(
		.INIT('h40)
	) name1836 (
		_w2166_,
		_w2981_,
		_w3011_,
		_w3017_
	);
	LUT3 #(
		.INIT('h13)
	) name1837 (
		_w2214_,
		_w3016_,
		_w3017_,
		_w3018_
	);
	LUT3 #(
		.INIT('h01)
	) name1838 (
		\g1220_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w3019_
	);
	LUT3 #(
		.INIT('h4c)
	) name1839 (
		_w2980_,
		_w3012_,
		_w3019_,
		_w3020_
	);
	LUT3 #(
		.INIT('h02)
	) name1840 (
		_w3011_,
		_w3015_,
		_w3020_,
		_w3021_
	);
	LUT3 #(
		.INIT('h07)
	) name1841 (
		_w2209_,
		_w3017_,
		_w3021_,
		_w3022_
	);
	LUT3 #(
		.INIT('h10)
	) name1842 (
		_w2166_,
		_w2223_,
		_w2981_,
		_w3023_
	);
	LUT3 #(
		.INIT('h01)
	) name1843 (
		\g1216_reg/NET0131 ,
		\g1245_reg/NET0131 ,
		\g1249_pad ,
		_w3024_
	);
	LUT3 #(
		.INIT('h4c)
	) name1844 (
		_w2980_,
		_w3012_,
		_w3024_,
		_w3025_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		_w3015_,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h1)
	) name1846 (
		_w3023_,
		_w3026_,
		_w3027_
	);
	LUT2 #(
		.INIT('he)
	) name1847 (
		_w2995_,
		_w3027_,
		_w3028_
	);
	LUT3 #(
		.INIT('h9a)
	) name1848 (
		_w2024_,
		_w2129_,
		_w2143_,
		_w3029_
	);
	LUT4 #(
		.INIT('h0200)
	) name1849 (
		_w2454_,
		_w2625_,
		_w2677_,
		_w3029_,
		_w3030_
	);
	LUT4 #(
		.INIT('h8488)
	) name1850 (
		_w2024_,
		_w2085_,
		_w2129_,
		_w2143_,
		_w3031_
	);
	LUT4 #(
		.INIT('h0200)
	) name1851 (
		_w2454_,
		_w2625_,
		_w2677_,
		_w3031_,
		_w3032_
	);
	LUT4 #(
		.INIT('h3301)
	) name1852 (
		_w2085_,
		_w2453_,
		_w3030_,
		_w3032_,
		_w3033_
	);
	LUT4 #(
		.INIT('hba8a)
	) name1853 (
		\g1496_reg/NET0131 ,
		_w2434_,
		_w2439_,
		_w3033_,
		_w3034_
	);
	LUT2 #(
		.INIT('h8)
	) name1854 (
		_w2315_,
		_w2328_,
		_w3035_
	);
	LUT2 #(
		.INIT('h4)
	) name1855 (
		_w2314_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h1)
	) name1856 (
		\g97_reg/NET0131 ,
		_w2315_,
		_w3037_
	);
	LUT3 #(
		.INIT('h40)
	) name1857 (
		\g97_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w3038_
	);
	LUT3 #(
		.INIT('hd0)
	) name1858 (
		_w1737_,
		_w2306_,
		_w3038_,
		_w3039_
	);
	LUT2 #(
		.INIT('h6)
	) name1859 (
		_w1783_,
		_w1821_,
		_w3040_
	);
	LUT3 #(
		.INIT('h10)
	) name1860 (
		_w1830_,
		_w2328_,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h8)
	) name1861 (
		_w2295_,
		_w3041_,
		_w3042_
	);
	LUT4 #(
		.INIT('h0203)
	) name1862 (
		_w2314_,
		_w3037_,
		_w3039_,
		_w3042_,
		_w3043_
	);
	LUT2 #(
		.INIT('h4)
	) name1863 (
		_w3036_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		\g113_reg/NET0131 ,
		_w2315_,
		_w3045_
	);
	LUT3 #(
		.INIT('h40)
	) name1865 (
		\g113_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w3046_
	);
	LUT3 #(
		.INIT('hd0)
	) name1866 (
		_w1737_,
		_w2306_,
		_w3046_,
		_w3047_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name1867 (
		_w1795_,
		_w2329_,
		_w2651_,
		_w2708_,
		_w3048_
	);
	LUT3 #(
		.INIT('h80)
	) name1868 (
		_w2295_,
		_w2641_,
		_w3048_,
		_w3049_
	);
	LUT4 #(
		.INIT('h0203)
	) name1869 (
		_w2314_,
		_w3045_,
		_w3047_,
		_w3049_,
		_w3050_
	);
	LUT2 #(
		.INIT('h4)
	) name1870 (
		_w3036_,
		_w3050_,
		_w3051_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		\g785_reg/NET0131 ,
		_w2342_,
		_w3052_
	);
	LUT3 #(
		.INIT('h20)
	) name1872 (
		\g785_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w3053_
	);
	LUT3 #(
		.INIT('h40)
	) name1873 (
		_w1950_,
		_w2347_,
		_w3053_,
		_w3054_
	);
	LUT2 #(
		.INIT('h6)
	) name1874 (
		_w1919_,
		_w1942_,
		_w3055_
	);
	LUT2 #(
		.INIT('h1)
	) name1875 (
		_w2365_,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h8)
	) name1876 (
		_w2342_,
		_w3056_,
		_w3057_
	);
	LUT4 #(
		.INIT('hfdfc)
	) name1877 (
		_w2350_,
		_w3052_,
		_w3054_,
		_w3057_,
		_w3058_
	);
	LUT2 #(
		.INIT('h6)
	) name1878 (
		_w2028_,
		_w2143_,
		_w3059_
	);
	LUT2 #(
		.INIT('h1)
	) name1879 (
		_w2453_,
		_w3059_,
		_w3060_
	);
	LUT4 #(
		.INIT('hba8a)
	) name1880 (
		\g1471_reg/NET0131 ,
		_w2434_,
		_w2439_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		\g801_reg/NET0131 ,
		_w2342_,
		_w3062_
	);
	LUT3 #(
		.INIT('h20)
	) name1882 (
		\g801_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w3063_
	);
	LUT3 #(
		.INIT('h40)
	) name1883 (
		_w1950_,
		_w2347_,
		_w3063_,
		_w3064_
	);
	LUT4 #(
		.INIT('ha6aa)
	) name1884 (
		_w1925_,
		_w2366_,
		_w2389_,
		_w2404_,
		_w3065_
	);
	LUT2 #(
		.INIT('h1)
	) name1885 (
		_w2365_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h8)
	) name1886 (
		_w2342_,
		_w3066_,
		_w3067_
	);
	LUT4 #(
		.INIT('hfdfc)
	) name1887 (
		_w2350_,
		_w3062_,
		_w3064_,
		_w3067_,
		_w3068_
	);
	LUT3 #(
		.INIT('h8a)
	) name1888 (
		\g2165_reg/NET0131 ,
		_w2477_,
		_w2480_,
		_w3069_
	);
	LUT2 #(
		.INIT('h8)
	) name1889 (
		\g2165_reg/NET0131 ,
		_w2472_,
		_w3070_
	);
	LUT4 #(
		.INIT('h020f)
	) name1890 (
		_w1333_,
		_w2466_,
		_w3069_,
		_w3070_,
		_w3071_
	);
	LUT2 #(
		.INIT('h9)
	) name1891 (
		_w1302_,
		_w1369_,
		_w3072_
	);
	LUT2 #(
		.INIT('h4)
	) name1892 (
		_w2472_,
		_w3072_,
		_w3073_
	);
	LUT3 #(
		.INIT('h84)
	) name1893 (
		_w1302_,
		_w1333_,
		_w1369_,
		_w3074_
	);
	LUT4 #(
		.INIT('hc4c0)
	) name1894 (
		_w2466_,
		_w2498_,
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('hd)
	) name1895 (
		_w3071_,
		_w3075_,
		_w3076_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1896 (
		_w1333_,
		_w2466_,
		_w2472_,
		_w2498_,
		_w3077_
	);
	LUT3 #(
		.INIT('h8a)
	) name1897 (
		\g2185_reg/NET0131 ,
		_w2477_,
		_w2480_,
		_w3078_
	);
	LUT2 #(
		.INIT('h8)
	) name1898 (
		\g2185_reg/NET0131 ,
		_w2472_,
		_w3079_
	);
	LUT4 #(
		.INIT('h020f)
	) name1899 (
		_w1333_,
		_w2466_,
		_w3078_,
		_w3079_,
		_w3080_
	);
	LUT4 #(
		.INIT('h0200)
	) name1900 (
		_w1274_,
		_w1275_,
		_w1304_,
		_w1305_,
		_w3081_
	);
	LUT3 #(
		.INIT('hb0)
	) name1901 (
		_w1368_,
		_w1369_,
		_w3081_,
		_w3082_
	);
	LUT3 #(
		.INIT('h40)
	) name1902 (
		_w1368_,
		_w1369_,
		_w2547_,
		_w3083_
	);
	LUT4 #(
		.INIT('h9995)
	) name1903 (
		_w1285_,
		_w2495_,
		_w3082_,
		_w3083_,
		_w3084_
	);
	LUT4 #(
		.INIT('h0004)
	) name1904 (
		_w2477_,
		_w2480_,
		_w2497_,
		_w3084_,
		_w3085_
	);
	LUT4 #(
		.INIT('h2f00)
	) name1905 (
		_w1333_,
		_w2466_,
		_w2472_,
		_w3085_,
		_w3086_
	);
	LUT3 #(
		.INIT('h0b)
	) name1906 (
		_w3077_,
		_w3080_,
		_w3086_,
		_w3087_
	);
	LUT3 #(
		.INIT('h8a)
	) name1907 (
		\g2195_reg/NET0131 ,
		_w2477_,
		_w2480_,
		_w3088_
	);
	LUT2 #(
		.INIT('h8)
	) name1908 (
		\g2195_reg/NET0131 ,
		_w2472_,
		_w3089_
	);
	LUT4 #(
		.INIT('h020f)
	) name1909 (
		_w1333_,
		_w2466_,
		_w3088_,
		_w3089_,
		_w3090_
	);
	LUT3 #(
		.INIT('h95)
	) name1910 (
		_w1290_,
		_w2584_,
		_w2585_,
		_w3091_
	);
	LUT2 #(
		.INIT('h8)
	) name1911 (
		_w2498_,
		_w3091_,
		_w3092_
	);
	LUT3 #(
		.INIT('h73)
	) name1912 (
		_w2473_,
		_w3090_,
		_w3092_,
		_w3093_
	);
	LUT4 #(
		.INIT('h5559)
	) name1913 (
		_w2024_,
		_w2454_,
		_w2625_,
		_w2677_,
		_w3094_
	);
	LUT2 #(
		.INIT('h4)
	) name1914 (
		_w2453_,
		_w3094_,
		_w3095_
	);
	LUT4 #(
		.INIT('hba8a)
	) name1915 (
		\g1491_reg/NET0131 ,
		_w2434_,
		_w2439_,
		_w3095_,
		_w3096_
	);
	LUT4 #(
		.INIT('h7e77)
	) name1916 (
		_w2024_,
		_w2085_,
		_w2129_,
		_w2143_,
		_w3097_
	);
	LUT4 #(
		.INIT('h1121)
	) name1917 (
		_w2020_,
		_w2453_,
		_w2678_,
		_w3097_,
		_w3098_
	);
	LUT4 #(
		.INIT('hba8a)
	) name1918 (
		\g1501_reg/NET0131 ,
		_w2434_,
		_w2439_,
		_w3098_,
		_w3099_
	);
	LUT2 #(
		.INIT('h2)
	) name1919 (
		\g809_reg/NET0131 ,
		_w2342_,
		_w3100_
	);
	LUT3 #(
		.INIT('h20)
	) name1920 (
		\g809_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w3101_
	);
	LUT3 #(
		.INIT('h40)
	) name1921 (
		_w1950_,
		_w2347_,
		_w3101_,
		_w3102_
	);
	LUT4 #(
		.INIT('h000b)
	) name1922 (
		_w2350_,
		_w2418_,
		_w3100_,
		_w3102_,
		_w3103_
	);
	LUT3 #(
		.INIT('h0b)
	) name1923 (
		_w1848_,
		_w1919_,
		_w1972_,
		_w3104_
	);
	LUT4 #(
		.INIT('h00f4)
	) name1924 (
		_w1848_,
		_w1919_,
		_w1972_,
		_w2409_,
		_w3105_
	);
	LUT4 #(
		.INIT('h2000)
	) name1925 (
		_w2366_,
		_w2389_,
		_w2405_,
		_w3105_,
		_w3106_
	);
	LUT2 #(
		.INIT('h1)
	) name1926 (
		_w1937_,
		_w3106_,
		_w3107_
	);
	LUT2 #(
		.INIT('h2)
	) name1927 (
		_w1937_,
		_w2409_,
		_w3108_
	);
	LUT2 #(
		.INIT('h4)
	) name1928 (
		_w3104_,
		_w3108_,
		_w3109_
	);
	LUT2 #(
		.INIT('h8)
	) name1929 (
		_w2406_,
		_w3109_,
		_w3110_
	);
	LUT4 #(
		.INIT('h0008)
	) name1930 (
		_w2341_,
		_w2417_,
		_w3107_,
		_w3110_,
		_w3111_
	);
	LUT2 #(
		.INIT('h4)
	) name1931 (
		_w2350_,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h1)
	) name1932 (
		_w3103_,
		_w3112_,
		_w3113_
	);
	LUT3 #(
		.INIT('h8a)
	) name1933 (
		\g2200_reg/NET0131 ,
		_w2477_,
		_w2480_,
		_w3114_
	);
	LUT2 #(
		.INIT('h8)
	) name1934 (
		\g2200_reg/NET0131 ,
		_w2472_,
		_w3115_
	);
	LUT4 #(
		.INIT('h020f)
	) name1935 (
		_w1333_,
		_w2466_,
		_w3114_,
		_w3115_,
		_w3116_
	);
	LUT3 #(
		.INIT('h9a)
	) name1936 (
		_w1290_,
		_w1368_,
		_w1369_,
		_w3117_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		_w2585_,
		_w3117_,
		_w3118_
	);
	LUT3 #(
		.INIT('h95)
	) name1938 (
		_w1256_,
		_w2584_,
		_w3118_,
		_w3119_
	);
	LUT2 #(
		.INIT('h8)
	) name1939 (
		_w2498_,
		_w3119_,
		_w3120_
	);
	LUT3 #(
		.INIT('h73)
	) name1940 (
		_w2473_,
		_w3116_,
		_w3120_,
		_w3121_
	);
	LUT3 #(
		.INIT('h2a)
	) name1941 (
		_w2093_,
		_w2678_,
		_w2685_,
		_w3122_
	);
	LUT4 #(
		.INIT('h2322)
	) name1942 (
		_w2024_,
		_w2093_,
		_w2129_,
		_w2143_,
		_w3123_
	);
	LUT3 #(
		.INIT('h40)
	) name1943 (
		_w2681_,
		_w2684_,
		_w3123_,
		_w3124_
	);
	LUT3 #(
		.INIT('h15)
	) name1944 (
		_w2453_,
		_w2678_,
		_w3124_,
		_w3125_
	);
	LUT2 #(
		.INIT('h4)
	) name1945 (
		_w3122_,
		_w3125_,
		_w3126_
	);
	LUT4 #(
		.INIT('hba8a)
	) name1946 (
		\g1506_reg/NET0131 ,
		_w2434_,
		_w2439_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('h2)
	) name1947 (
		\g813_reg/NET0131 ,
		_w2342_,
		_w3128_
	);
	LUT3 #(
		.INIT('h20)
	) name1948 (
		\g813_reg/NET0131 ,
		_w1849_,
		_w1850_,
		_w3129_
	);
	LUT3 #(
		.INIT('h40)
	) name1949 (
		_w1950_,
		_w2347_,
		_w3129_,
		_w3130_
	);
	LUT4 #(
		.INIT('h2000)
	) name1950 (
		_w2366_,
		_w2389_,
		_w2405_,
		_w2410_,
		_w3131_
	);
	LUT2 #(
		.INIT('h2)
	) name1951 (
		_w1967_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h1)
	) name1952 (
		_w1967_,
		_w2409_,
		_w3133_
	);
	LUT2 #(
		.INIT('h4)
	) name1953 (
		_w2408_,
		_w3133_,
		_w3134_
	);
	LUT2 #(
		.INIT('h8)
	) name1954 (
		_w2406_,
		_w3134_,
		_w3135_
	);
	LUT4 #(
		.INIT('h0008)
	) name1955 (
		_w2341_,
		_w2417_,
		_w3132_,
		_w3135_,
		_w3136_
	);
	LUT4 #(
		.INIT('hfdfc)
	) name1956 (
		_w2350_,
		_w3128_,
		_w3130_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h2)
	) name1957 (
		\g125_reg/NET0131 ,
		_w2315_,
		_w3138_
	);
	LUT3 #(
		.INIT('h80)
	) name1958 (
		\g125_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w3139_
	);
	LUT3 #(
		.INIT('hd0)
	) name1959 (
		_w1737_,
		_w2306_,
		_w3139_,
		_w3140_
	);
	LUT4 #(
		.INIT('h2130)
	) name1960 (
		_w1697_,
		_w1761_,
		_w1774_,
		_w1821_,
		_w3141_
	);
	LUT2 #(
		.INIT('h4)
	) name1961 (
		_w2711_,
		_w3141_,
		_w3142_
	);
	LUT4 #(
		.INIT('h11d5)
	) name1962 (
		_w1761_,
		_w2710_,
		_w2712_,
		_w3142_,
		_w3143_
	);
	LUT3 #(
		.INIT('h80)
	) name1963 (
		_w2295_,
		_w2641_,
		_w3143_,
		_w3144_
	);
	LUT4 #(
		.INIT('hfdfc)
	) name1964 (
		_w2314_,
		_w3138_,
		_w3140_,
		_w3144_,
		_w3145_
	);
	LUT3 #(
		.INIT('hfe)
	) name1965 (
		_w1507_,
		_w1512_,
		_w1516_,
		_w3146_
	);
	LUT3 #(
		.INIT('h2a)
	) name1966 (
		_w1613_,
		_w2169_,
		_w2230_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name1967 (
		_w2218_,
		_w2233_,
		_w3148_
	);
	LUT3 #(
		.INIT('h08)
	) name1968 (
		_w2174_,
		_w2180_,
		_w2233_,
		_w3149_
	);
	LUT3 #(
		.INIT('h13)
	) name1969 (
		_w2205_,
		_w3148_,
		_w3149_,
		_w3150_
	);
	LUT4 #(
		.INIT('h0504)
	) name1970 (
		\g1196_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1222_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w3151_
	);
	LUT2 #(
		.INIT('h8)
	) name1971 (
		_w2167_,
		_w3151_,
		_w3152_
	);
	LUT3 #(
		.INIT('h8c)
	) name1972 (
		_w2166_,
		_w3012_,
		_w3152_,
		_w3153_
	);
	LUT3 #(
		.INIT('hd0)
	) name1973 (
		_w2221_,
		_w3150_,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('he)
	) name1974 (
		_w3147_,
		_w3154_,
		_w3155_
	);
	LUT3 #(
		.INIT('h10)
	) name1975 (
		_w2166_,
		_w2216_,
		_w2996_,
		_w3156_
	);
	LUT4 #(
		.INIT('h0504)
	) name1976 (
		\g1196_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1223_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w3157_
	);
	LUT2 #(
		.INIT('h8)
	) name1977 (
		_w2167_,
		_w3157_,
		_w3158_
	);
	LUT3 #(
		.INIT('h8c)
	) name1978 (
		_w2166_,
		_w3012_,
		_w3158_,
		_w3159_
	);
	LUT3 #(
		.INIT('h45)
	) name1979 (
		_w1613_,
		_w3156_,
		_w3159_,
		_w3160_
	);
	LUT3 #(
		.INIT('h8a)
	) name1980 (
		_w2169_,
		_w3156_,
		_w3159_,
		_w3161_
	);
	LUT3 #(
		.INIT('h13)
	) name1981 (
		_w2231_,
		_w3160_,
		_w3161_,
		_w3162_
	);
	LUT3 #(
		.INIT('hf4)
	) name1982 (
		_w1687_,
		_w1688_,
		_w1689_,
		_w3163_
	);
	LUT2 #(
		.INIT('h4)
	) name1983 (
		_w1830_,
		_w2320_,
		_w3164_
	);
	LUT3 #(
		.INIT('h04)
	) name1984 (
		_w1700_,
		_w1737_,
		_w2291_,
		_w3165_
	);
	LUT2 #(
		.INIT('h4)
	) name1985 (
		_w1830_,
		_w3165_,
		_w3166_
	);
	LUT3 #(
		.INIT('hdc)
	) name1986 (
		_w2306_,
		_w3164_,
		_w3166_,
		_w3167_
	);
	LUT2 #(
		.INIT('h4)
	) name1987 (
		_w1918_,
		_w2351_,
		_w3168_
	);
	LUT2 #(
		.INIT('h1)
	) name1988 (
		_w1859_,
		_w2337_,
		_w3169_
	);
	LUT2 #(
		.INIT('h4)
	) name1989 (
		_w1918_,
		_w3169_,
		_w3170_
	);
	LUT4 #(
		.INIT('hfbf0)
	) name1990 (
		_w1950_,
		_w2933_,
		_w3168_,
		_w3170_,
		_w3171_
	);
	LUT3 #(
		.INIT('h02)
	) name1991 (
		_w1333_,
		_w1364_,
		_w2474_,
		_w3172_
	);
	LUT4 #(
		.INIT('h5150)
	) name1992 (
		_w1375_,
		_w2466_,
		_w2481_,
		_w3172_,
		_w3173_
	);
	LUT3 #(
		.INIT('h02)
	) name1993 (
		_w2010_,
		_w2121_,
		_w2435_,
		_w3174_
	);
	LUT3 #(
		.INIT('hb0)
	) name1994 (
		_w2105_,
		_w2109_,
		_w3174_,
		_w3175_
	);
	LUT3 #(
		.INIT('hb0)
	) name1995 (
		_w2035_,
		_w2040_,
		_w3174_,
		_w3176_
	);
	LUT4 #(
		.INIT('h5554)
	) name1996 (
		_w2141_,
		_w2440_,
		_w3175_,
		_w3176_,
		_w3177_
	);
	LUT3 #(
		.INIT('h54)
	) name1997 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g525_reg/NET0131 ,
		_w3178_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		_w2821_,
		_w3178_,
		_w3179_
	);
	LUT3 #(
		.INIT('h32)
	) name1999 (
		\g1196_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		\g525_reg/NET0131 ,
		_w3180_
	);
	LUT3 #(
		.INIT('h23)
	) name2000 (
		\g499_reg/NET0131 ,
		\g530_reg/NET0131 ,
		\g5657_pad ,
		_w3181_
	);
	LUT4 #(
		.INIT('h4000)
	) name2001 (
		_w2898_,
		_w2899_,
		_w3178_,
		_w3181_,
		_w3182_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2002 (
		_w2877_,
		_w3179_,
		_w3180_,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h1)
	) name2003 (
		_w1613_,
		_w3183_,
		_w3184_
	);
	LUT2 #(
		.INIT('h2)
	) name2004 (
		\g5657_pad ,
		\g735_reg/NET0131 ,
		_w3185_
	);
	LUT4 #(
		.INIT('hf351)
	) name2005 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g734_reg/NET0131 ,
		\g736_reg/NET0131 ,
		_w3186_
	);
	LUT3 #(
		.INIT('h8a)
	) name2006 (
		\g499_reg/NET0131 ,
		_w3185_,
		_w3186_,
		_w3187_
	);
	LUT3 #(
		.INIT('h80)
	) name2007 (
		\g499_reg/NET0131 ,
		_w2827_,
		_w2832_,
		_w3188_
	);
	LUT3 #(
		.INIT('h13)
	) name2008 (
		_w2858_,
		_w3187_,
		_w3188_,
		_w3189_
	);
	LUT2 #(
		.INIT('h2)
	) name2009 (
		_w2902_,
		_w3183_,
		_w3190_
	);
	LUT3 #(
		.INIT('h15)
	) name2010 (
		_w3184_,
		_w3189_,
		_w3190_,
		_w3191_
	);
	LUT3 #(
		.INIT('h23)
	) name2011 (
		\g499_reg/NET0131 ,
		\g531_reg/NET0131 ,
		\g5657_pad ,
		_w3192_
	);
	LUT4 #(
		.INIT('h4000)
	) name2012 (
		_w2898_,
		_w2899_,
		_w3178_,
		_w3192_,
		_w3193_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2013 (
		_w2874_,
		_w3179_,
		_w3180_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h1)
	) name2014 (
		_w1613_,
		_w3194_,
		_w3195_
	);
	LUT2 #(
		.INIT('h2)
	) name2015 (
		_w2902_,
		_w3194_,
		_w3196_
	);
	LUT3 #(
		.INIT('h13)
	) name2016 (
		_w3189_,
		_w3195_,
		_w3196_,
		_w3197_
	);
	LUT3 #(
		.INIT('h23)
	) name2017 (
		\g499_reg/NET0131 ,
		\g529_reg/NET0131 ,
		\g5657_pad ,
		_w3198_
	);
	LUT4 #(
		.INIT('h4000)
	) name2018 (
		_w2898_,
		_w2899_,
		_w3178_,
		_w3198_,
		_w3199_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2019 (
		_w2876_,
		_w3179_,
		_w3180_,
		_w3199_,
		_w3200_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w1613_,
		_w3200_,
		_w3201_
	);
	LUT2 #(
		.INIT('h2)
	) name2021 (
		_w2900_,
		_w3200_,
		_w3202_
	);
	LUT3 #(
		.INIT('h23)
	) name2022 (
		_w3189_,
		_w3201_,
		_w3202_,
		_w3203_
	);
	LUT3 #(
		.INIT('h23)
	) name2023 (
		\g499_reg/NET0131 ,
		\g532_reg/NET0131 ,
		\g5657_pad ,
		_w3204_
	);
	LUT4 #(
		.INIT('h4000)
	) name2024 (
		_w2898_,
		_w2899_,
		_w3178_,
		_w3204_,
		_w3205_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2025 (
		_w2873_,
		_w3179_,
		_w3180_,
		_w3205_,
		_w3206_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		_w1613_,
		_w3206_,
		_w3207_
	);
	LUT2 #(
		.INIT('h2)
	) name2027 (
		_w2900_,
		_w3206_,
		_w3208_
	);
	LUT3 #(
		.INIT('h23)
	) name2028 (
		_w3189_,
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT4 #(
		.INIT('haa8a)
	) name2029 (
		_w1613_,
		_w2898_,
		_w2899_,
		_w2901_,
		_w3210_
	);
	LUT3 #(
		.INIT('h23)
	) name2030 (
		\g499_reg/NET0131 ,
		\g533_reg/NET0131 ,
		\g5657_pad ,
		_w3211_
	);
	LUT4 #(
		.INIT('h4000)
	) name2031 (
		_w2898_,
		_w2899_,
		_w3178_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h2)
	) name2032 (
		_w3180_,
		_w3212_,
		_w3213_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name2033 (
		_w2862_,
		_w3179_,
		_w3210_,
		_w3213_,
		_w3214_
	);
	LUT3 #(
		.INIT('h23)
	) name2034 (
		\g499_reg/NET0131 ,
		\g534_reg/NET0131 ,
		\g5657_pad ,
		_w3215_
	);
	LUT4 #(
		.INIT('h4000)
	) name2035 (
		_w2898_,
		_w2899_,
		_w3178_,
		_w3215_,
		_w3216_
	);
	LUT2 #(
		.INIT('h2)
	) name2036 (
		_w3180_,
		_w3216_,
		_w3217_
	);
	LUT4 #(
		.INIT('hf7f0)
	) name2037 (
		_w2866_,
		_w3179_,
		_w3210_,
		_w3217_,
		_w3218_
	);
	LUT4 #(
		.INIT('hff10)
	) name2038 (
		_w2952_,
		_w2953_,
		_w2954_,
		_w2955_,
		_w3219_
	);
	LUT2 #(
		.INIT('h8)
	) name2039 (
		\g1018_reg/NET0131 ,
		\g1038_reg/NET0131 ,
		_w3220_
	);
	LUT4 #(
		.INIT('h135f)
	) name2040 (
		\g1024_reg/NET0131 ,
		\g1036_reg/NET0131 ,
		\g1040_reg/NET0131 ,
		\g5657_pad ,
		_w3221_
	);
	LUT2 #(
		.INIT('h4)
	) name2041 (
		_w3220_,
		_w3221_,
		_w3222_
	);
	LUT2 #(
		.INIT('h8)
	) name2042 (
		\g1024_reg/NET0131 ,
		\g1055_reg/NET0131 ,
		_w3223_
	);
	LUT4 #(
		.INIT('h135f)
	) name2043 (
		\g1018_reg/NET0131 ,
		\g1051_reg/NET0131 ,
		\g1053_reg/NET0131 ,
		\g5657_pad ,
		_w3224_
	);
	LUT4 #(
		.INIT('h0400)
	) name2044 (
		_w3220_,
		_w3221_,
		_w3223_,
		_w3224_,
		_w3225_
	);
	LUT2 #(
		.INIT('h4)
	) name2045 (
		\g1262_reg/NET0131 ,
		\g5657_pad ,
		_w3226_
	);
	LUT4 #(
		.INIT('hf351)
	) name2046 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1261_reg/NET0131 ,
		\g1263_reg/NET0131 ,
		_w3227_
	);
	LUT2 #(
		.INIT('h4)
	) name2047 (
		_w3226_,
		_w3227_,
		_w3228_
	);
	LUT2 #(
		.INIT('h2)
	) name2048 (
		\g1024_reg/NET0131 ,
		\g1264_reg/NET0131 ,
		_w3229_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2049 (
		\g1018_reg/NET0131 ,
		\g1265_reg/NET0131 ,
		\g1266_reg/NET0131 ,
		\g5657_pad ,
		_w3230_
	);
	LUT2 #(
		.INIT('h4)
	) name2050 (
		_w3229_,
		_w3230_,
		_w3231_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2051 (
		_w3226_,
		_w3227_,
		_w3229_,
		_w3230_,
		_w3232_
	);
	LUT2 #(
		.INIT('h8)
	) name2052 (
		_w3225_,
		_w3232_,
		_w3233_
	);
	LUT2 #(
		.INIT('h8)
	) name2053 (
		\g1024_reg/NET0131 ,
		\g1070_reg/NET0131 ,
		_w3234_
	);
	LUT4 #(
		.INIT('h135f)
	) name2054 (
		\g1018_reg/NET0131 ,
		\g1066_reg/NET0131 ,
		\g1068_reg/NET0131 ,
		\g5657_pad ,
		_w3235_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2055 (
		_w3223_,
		_w3224_,
		_w3234_,
		_w3235_,
		_w3236_
	);
	LUT2 #(
		.INIT('h2)
	) name2056 (
		\g1018_reg/NET0131 ,
		\g1269_reg/NET0131 ,
		_w3237_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2057 (
		\g1024_reg/NET0131 ,
		\g1267_reg/NET0131 ,
		\g1268_reg/NET0131 ,
		\g5657_pad ,
		_w3238_
	);
	LUT2 #(
		.INIT('h4)
	) name2058 (
		_w3237_,
		_w3238_,
		_w3239_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2059 (
		_w3220_,
		_w3221_,
		_w3237_,
		_w3238_,
		_w3240_
	);
	LUT3 #(
		.INIT('h80)
	) name2060 (
		_w3228_,
		_w3236_,
		_w3240_,
		_w3241_
	);
	LUT4 #(
		.INIT('h0400)
	) name2061 (
		_w3220_,
		_w3221_,
		_w3234_,
		_w3235_,
		_w3242_
	);
	LUT4 #(
		.INIT('h4044)
	) name2062 (
		_w3223_,
		_w3224_,
		_w3237_,
		_w3238_,
		_w3243_
	);
	LUT3 #(
		.INIT('h10)
	) name2063 (
		_w3228_,
		_w3242_,
		_w3243_,
		_w3244_
	);
	LUT3 #(
		.INIT('h01)
	) name2064 (
		_w3233_,
		_w3241_,
		_w3244_,
		_w3245_
	);
	LUT4 #(
		.INIT('h0400)
	) name2065 (
		_w3220_,
		_w3221_,
		_w3229_,
		_w3230_,
		_w3246_
	);
	LUT3 #(
		.INIT('h80)
	) name2066 (
		_w3228_,
		_w3236_,
		_w3246_,
		_w3247_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\g1024_reg/NET0131 ,
		\g1270_reg/NET0131 ,
		_w3248_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2068 (
		\g1018_reg/NET0131 ,
		\g1271_reg/NET0131 ,
		\g1272_reg/NET0131 ,
		\g5657_pad ,
		_w3249_
	);
	LUT2 #(
		.INIT('h4)
	) name2069 (
		_w3248_,
		_w3249_,
		_w3250_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2070 (
		_w3220_,
		_w3221_,
		_w3248_,
		_w3249_,
		_w3251_
	);
	LUT2 #(
		.INIT('h8)
	) name2071 (
		\g1011_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		_w3252_
	);
	LUT4 #(
		.INIT('h135f)
	) name2072 (
		\g1018_reg/NET0131 ,
		\g1081_reg/NET0131 ,
		\g1083_reg/NET0131 ,
		\g5657_pad ,
		_w3253_
	);
	LUT2 #(
		.INIT('h4)
	) name2073 (
		_w3252_,
		_w3253_,
		_w3254_
	);
	LUT4 #(
		.INIT('h0400)
	) name2074 (
		_w3226_,
		_w3227_,
		_w3252_,
		_w3253_,
		_w3255_
	);
	LUT3 #(
		.INIT('hd0)
	) name2075 (
		_w3239_,
		_w3251_,
		_w3255_,
		_w3256_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2076 (
		_w3220_,
		_w3221_,
		_w3234_,
		_w3235_,
		_w3257_
	);
	LUT3 #(
		.INIT('h10)
	) name2077 (
		_w3231_,
		_w3243_,
		_w3257_,
		_w3258_
	);
	LUT3 #(
		.INIT('h01)
	) name2078 (
		_w3247_,
		_w3256_,
		_w3258_,
		_w3259_
	);
	LUT2 #(
		.INIT('h8)
	) name2079 (
		\g1018_reg/NET0131 ,
		\g1253_reg/NET0131 ,
		_w3260_
	);
	LUT4 #(
		.INIT('h0777)
	) name2080 (
		\g1024_reg/NET0131 ,
		\g1176_reg/NET0131 ,
		\g1251_reg/NET0131 ,
		\g5657_pad ,
		_w3261_
	);
	LUT2 #(
		.INIT('h4)
	) name2081 (
		_w3260_,
		_w3261_,
		_w3262_
	);
	LUT2 #(
		.INIT('h8)
	) name2082 (
		\g1228_reg/NET0131 ,
		\g185_reg/NET0131 ,
		_w3263_
	);
	LUT3 #(
		.INIT('hb0)
	) name2083 (
		_w3260_,
		_w3261_,
		_w3263_,
		_w3264_
	);
	LUT2 #(
		.INIT('h8)
	) name2084 (
		\g1018_reg/NET0131 ,
		\g1285_reg/NET0131 ,
		_w3265_
	);
	LUT4 #(
		.INIT('h135f)
	) name2085 (
		\g1024_reg/NET0131 ,
		\g1282_reg/NET0131 ,
		\g1288_reg/NET0131 ,
		\g5657_pad ,
		_w3266_
	);
	LUT2 #(
		.INIT('h4)
	) name2086 (
		_w3265_,
		_w3266_,
		_w3267_
	);
	LUT2 #(
		.INIT('h4)
	) name2087 (
		_w3264_,
		_w3267_,
		_w3268_
	);
	LUT4 #(
		.INIT('h4044)
	) name2088 (
		_w3234_,
		_w3235_,
		_w3248_,
		_w3249_,
		_w3269_
	);
	LUT4 #(
		.INIT('h0400)
	) name2089 (
		_w3229_,
		_w3230_,
		_w3237_,
		_w3238_,
		_w3270_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2090 (
		_w3223_,
		_w3224_,
		_w3234_,
		_w3235_,
		_w3271_
	);
	LUT3 #(
		.INIT('h15)
	) name2091 (
		_w3269_,
		_w3270_,
		_w3271_,
		_w3272_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2092 (
		_w3226_,
		_w3227_,
		_w3252_,
		_w3253_,
		_w3273_
	);
	LUT3 #(
		.INIT('h8a)
	) name2093 (
		_w3222_,
		_w3250_,
		_w3273_,
		_w3274_
	);
	LUT4 #(
		.INIT('h4044)
	) name2094 (
		_w3223_,
		_w3224_,
		_w3234_,
		_w3235_,
		_w3275_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2095 (
		_w3226_,
		_w3227_,
		_w3248_,
		_w3249_,
		_w3276_
	);
	LUT2 #(
		.INIT('h8)
	) name2096 (
		_w3275_,
		_w3276_,
		_w3277_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2097 (
		_w3223_,
		_w3224_,
		_w3252_,
		_w3253_,
		_w3278_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2098 (
		_w3229_,
		_w3230_,
		_w3237_,
		_w3238_,
		_w3279_
	);
	LUT3 #(
		.INIT('h15)
	) name2099 (
		_w3222_,
		_w3278_,
		_w3279_,
		_w3280_
	);
	LUT4 #(
		.INIT('h7077)
	) name2100 (
		_w3272_,
		_w3274_,
		_w3277_,
		_w3280_,
		_w3281_
	);
	LUT4 #(
		.INIT('h0080)
	) name2101 (
		_w3245_,
		_w3259_,
		_w3268_,
		_w3281_,
		_w3282_
	);
	LUT4 #(
		.INIT('h27af)
	) name2102 (
		_w3231_,
		_w3239_,
		_w3242_,
		_w3254_,
		_w3283_
	);
	LUT4 #(
		.INIT('h4044)
	) name2103 (
		_w3226_,
		_w3227_,
		_w3229_,
		_w3230_,
		_w3284_
	);
	LUT2 #(
		.INIT('h8)
	) name2104 (
		_w3275_,
		_w3284_,
		_w3285_
	);
	LUT3 #(
		.INIT('h0e)
	) name2105 (
		_w3228_,
		_w3283_,
		_w3285_,
		_w3286_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2106 (
		_w3220_,
		_w3221_,
		_w3226_,
		_w3227_,
		_w3287_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2107 (
		_w3226_,
		_w3227_,
		_w3237_,
		_w3238_,
		_w3288_
	);
	LUT4 #(
		.INIT('h4022)
	) name2108 (
		_w3222_,
		_w3228_,
		_w3231_,
		_w3239_,
		_w3289_
	);
	LUT4 #(
		.INIT('h135f)
	) name2109 (
		_w3225_,
		_w3243_,
		_w3279_,
		_w3287_,
		_w3290_
	);
	LUT3 #(
		.INIT('h70)
	) name2110 (
		_w3278_,
		_w3289_,
		_w3290_,
		_w3291_
	);
	LUT3 #(
		.INIT('h80)
	) name2111 (
		_w3236_,
		_w3246_,
		_w3276_,
		_w3292_
	);
	LUT4 #(
		.INIT('h0400)
	) name2112 (
		_w3226_,
		_w3227_,
		_w3229_,
		_w3230_,
		_w3293_
	);
	LUT3 #(
		.INIT('h80)
	) name2113 (
		_w3250_,
		_w3257_,
		_w3293_,
		_w3294_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2114 (
		_w3220_,
		_w3221_,
		_w3248_,
		_w3249_,
		_w3295_
	);
	LUT2 #(
		.INIT('h8)
	) name2115 (
		_w3236_,
		_w3295_,
		_w3296_
	);
	LUT2 #(
		.INIT('h8)
	) name2116 (
		\g1255_reg/NET0131 ,
		\g5657_pad ,
		_w3297_
	);
	LUT4 #(
		.INIT('h135f)
	) name2117 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1257_reg/NET0131 ,
		\g1259_reg/NET0131 ,
		_w3298_
	);
	LUT2 #(
		.INIT('h4)
	) name2118 (
		_w3297_,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('h8)
	) name2119 (
		\g1210_reg/NET0131 ,
		\g185_reg/NET0131 ,
		_w3300_
	);
	LUT3 #(
		.INIT('hb0)
	) name2120 (
		_w3297_,
		_w3298_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h8)
	) name2121 (
		\g1024_reg/NET0131 ,
		\g1279_reg/NET0131 ,
		_w3302_
	);
	LUT4 #(
		.INIT('h135f)
	) name2122 (
		\g1018_reg/NET0131 ,
		\g1273_reg/NET0131 ,
		\g1276_reg/NET0131 ,
		\g5657_pad ,
		_w3303_
	);
	LUT2 #(
		.INIT('h4)
	) name2123 (
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2124 (
		_w3264_,
		_w3267_,
		_w3301_,
		_w3304_,
		_w3305_
	);
	LUT4 #(
		.INIT('h0001)
	) name2125 (
		_w3292_,
		_w3294_,
		_w3296_,
		_w3305_,
		_w3306_
	);
	LUT3 #(
		.INIT('h80)
	) name2126 (
		_w3286_,
		_w3291_,
		_w3306_,
		_w3307_
	);
	LUT3 #(
		.INIT('h40)
	) name2127 (
		\g3010_reg/NET0131 ,
		\g3013_reg/NET0131 ,
		\g3024_reg/NET0131 ,
		_w3308_
	);
	LUT4 #(
		.INIT('h0040)
	) name2128 (
		\g2993_reg/NET0131 ,
		\g2998_reg/NET0131 ,
		\g3002_reg/NET0131 ,
		\g3006_reg/NET0131 ,
		_w3309_
	);
	LUT2 #(
		.INIT('h1)
	) name2129 (
		\g3032_reg/NET0131 ,
		\g3036_reg/NET0131 ,
		_w3310_
	);
	LUT2 #(
		.INIT('h8)
	) name2130 (
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		_w3311_
	);
	LUT3 #(
		.INIT('h80)
	) name2131 (
		\g1024_reg/NET0131 ,
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		_w3312_
	);
	LUT4 #(
		.INIT('h8000)
	) name2132 (
		_w3308_,
		_w3309_,
		_w3310_,
		_w3312_,
		_w3313_
	);
	LUT4 #(
		.INIT('h0008)
	) name2133 (
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		\g3032_reg/NET0131 ,
		\g3036_reg/NET0131 ,
		_w3314_
	);
	LUT3 #(
		.INIT('h80)
	) name2134 (
		_w3308_,
		_w3309_,
		_w3314_,
		_w3315_
	);
	LUT3 #(
		.INIT('h7f)
	) name2135 (
		_w3308_,
		_w3309_,
		_w3314_,
		_w3316_
	);
	LUT3 #(
		.INIT('h20)
	) name2136 (
		\g1024_reg/NET0131 ,
		_w2206_,
		_w2207_,
		_w3317_
	);
	LUT2 #(
		.INIT('h1)
	) name2137 (
		\g1024_reg/NET0131 ,
		\g1306_reg/NET0131 ,
		_w3318_
	);
	LUT3 #(
		.INIT('h0b)
	) name2138 (
		_w3315_,
		_w3317_,
		_w3318_,
		_w3319_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2139 (
		_w3282_,
		_w3307_,
		_w3313_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h8)
	) name2140 (
		\g1018_reg/NET0131 ,
		\g2426_reg/NET0131 ,
		_w3321_
	);
	LUT4 #(
		.INIT('h135f)
	) name2141 (
		\g1024_reg/NET0131 ,
		\g2424_reg/NET0131 ,
		\g2428_reg/NET0131 ,
		\g5657_pad ,
		_w3322_
	);
	LUT2 #(
		.INIT('h4)
	) name2142 (
		_w3321_,
		_w3322_,
		_w3323_
	);
	LUT2 #(
		.INIT('h8)
	) name2143 (
		\g1018_reg/NET0131 ,
		\g2441_reg/NET0131 ,
		_w3324_
	);
	LUT4 #(
		.INIT('h135f)
	) name2144 (
		\g1024_reg/NET0131 ,
		\g2439_reg/NET0131 ,
		\g2443_reg/NET0131 ,
		\g5657_pad ,
		_w3325_
	);
	LUT2 #(
		.INIT('h4)
	) name2145 (
		_w3324_,
		_w3325_,
		_w3326_
	);
	LUT4 #(
		.INIT('h0400)
	) name2146 (
		_w3321_,
		_w3322_,
		_w3324_,
		_w3325_,
		_w3327_
	);
	LUT2 #(
		.INIT('h4)
	) name2147 (
		\g2653_reg/NET0131 ,
		\g5657_pad ,
		_w3328_
	);
	LUT4 #(
		.INIT('hf351)
	) name2148 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2652_reg/NET0131 ,
		\g2654_reg/NET0131 ,
		_w3329_
	);
	LUT2 #(
		.INIT('h4)
	) name2149 (
		_w3328_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h4)
	) name2150 (
		\g2650_reg/NET0131 ,
		\g5657_pad ,
		_w3331_
	);
	LUT4 #(
		.INIT('hf351)
	) name2151 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2649_reg/NET0131 ,
		\g2651_reg/NET0131 ,
		_w3332_
	);
	LUT2 #(
		.INIT('h4)
	) name2152 (
		_w3331_,
		_w3332_,
		_w3333_
	);
	LUT4 #(
		.INIT('h4044)
	) name2153 (
		_w3328_,
		_w3329_,
		_w3331_,
		_w3332_,
		_w3334_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2154 (
		_w3321_,
		_w3322_,
		_w3324_,
		_w3325_,
		_w3335_
	);
	LUT2 #(
		.INIT('h2)
	) name2155 (
		\g1018_reg/NET0131 ,
		\g2657_reg/NET0131 ,
		_w3336_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name2156 (
		\g1024_reg/NET0131 ,
		\g2655_reg/NET0131 ,
		\g2656_reg/NET0131 ,
		\g5657_pad ,
		_w3337_
	);
	LUT2 #(
		.INIT('h4)
	) name2157 (
		_w3336_,
		_w3337_,
		_w3338_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2158 (
		_w3331_,
		_w3332_,
		_w3336_,
		_w3337_,
		_w3339_
	);
	LUT4 #(
		.INIT('h3b7f)
	) name2159 (
		_w3323_,
		_w3326_,
		_w3334_,
		_w3339_,
		_w3340_
	);
	LUT2 #(
		.INIT('h8)
	) name2160 (
		\g1018_reg/NET0131 ,
		\g2456_reg/NET0131 ,
		_w3341_
	);
	LUT4 #(
		.INIT('h135f)
	) name2161 (
		\g1024_reg/NET0131 ,
		\g2454_reg/NET0131 ,
		\g2458_reg/NET0131 ,
		\g5657_pad ,
		_w3342_
	);
	LUT2 #(
		.INIT('h4)
	) name2162 (
		_w3341_,
		_w3342_,
		_w3343_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2163 (
		_w3321_,
		_w3322_,
		_w3341_,
		_w3342_,
		_w3344_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2164 (
		_w3324_,
		_w3325_,
		_w3328_,
		_w3329_,
		_w3345_
	);
	LUT2 #(
		.INIT('h8)
	) name2165 (
		_w3344_,
		_w3345_,
		_w3346_
	);
	LUT4 #(
		.INIT('h0400)
	) name2166 (
		_w3321_,
		_w3322_,
		_w3341_,
		_w3342_,
		_w3347_
	);
	LUT2 #(
		.INIT('h4)
	) name2167 (
		\g2659_reg/NET0131 ,
		\g5657_pad ,
		_w3348_
	);
	LUT4 #(
		.INIT('hf351)
	) name2168 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2658_reg/NET0131 ,
		\g2660_reg/NET0131 ,
		_w3349_
	);
	LUT2 #(
		.INIT('h4)
	) name2169 (
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT4 #(
		.INIT('h4044)
	) name2170 (
		_w3321_,
		_w3322_,
		_w3331_,
		_w3332_,
		_w3351_
	);
	LUT2 #(
		.INIT('h8)
	) name2171 (
		\g1018_reg/NET0131 ,
		\g2471_reg/NET0131 ,
		_w3352_
	);
	LUT4 #(
		.INIT('h0777)
	) name2172 (
		\g1024_reg/NET0131 ,
		\g2399_reg/NET0131 ,
		\g2469_reg/NET0131 ,
		\g5657_pad ,
		_w3353_
	);
	LUT2 #(
		.INIT('h4)
	) name2173 (
		_w3352_,
		_w3353_,
		_w3354_
	);
	LUT4 #(
		.INIT('hddcd)
	) name2174 (
		_w3347_,
		_w3350_,
		_w3351_,
		_w3354_,
		_w3355_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2175 (
		_w3321_,
		_w3322_,
		_w3331_,
		_w3332_,
		_w3356_
	);
	LUT4 #(
		.INIT('h0400)
	) name2176 (
		_w3348_,
		_w3349_,
		_w3352_,
		_w3353_,
		_w3357_
	);
	LUT2 #(
		.INIT('h8)
	) name2177 (
		_w3356_,
		_w3357_,
		_w3358_
	);
	LUT4 #(
		.INIT('h0020)
	) name2178 (
		_w3340_,
		_w3346_,
		_w3355_,
		_w3358_,
		_w3359_
	);
	LUT4 #(
		.INIT('h4044)
	) name2179 (
		_w3324_,
		_w3325_,
		_w3341_,
		_w3342_,
		_w3360_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2180 (
		_w3331_,
		_w3332_,
		_w3348_,
		_w3349_,
		_w3361_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name2181 (
		_w3323_,
		_w3339_,
		_w3360_,
		_w3361_,
		_w3362_
	);
	LUT4 #(
		.INIT('h4044)
	) name2182 (
		_w3331_,
		_w3332_,
		_w3336_,
		_w3337_,
		_w3363_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2183 (
		_w3324_,
		_w3325_,
		_w3341_,
		_w3342_,
		_w3364_
	);
	LUT4 #(
		.INIT('hd0c0)
	) name2184 (
		_w3323_,
		_w3354_,
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h1)
	) name2185 (
		_w3362_,
		_w3365_,
		_w3366_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2186 (
		_w3324_,
		_w3325_,
		_w3352_,
		_w3353_,
		_w3367_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2187 (
		_w3328_,
		_w3329_,
		_w3336_,
		_w3337_,
		_w3368_
	);
	LUT4 #(
		.INIT('h5400)
	) name2188 (
		_w3323_,
		_w3343_,
		_w3367_,
		_w3368_,
		_w3369_
	);
	LUT4 #(
		.INIT('h0400)
	) name2189 (
		_w3328_,
		_w3329_,
		_w3336_,
		_w3337_,
		_w3370_
	);
	LUT3 #(
		.INIT('h40)
	) name2190 (
		_w3326_,
		_w3347_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h8)
	) name2191 (
		\g1024_reg/NET0131 ,
		\g2564_reg/NET0131 ,
		_w3372_
	);
	LUT4 #(
		.INIT('h135f)
	) name2192 (
		\g1018_reg/NET0131 ,
		\g2639_reg/NET0131 ,
		\g2641_reg/NET0131 ,
		\g5657_pad ,
		_w3373_
	);
	LUT2 #(
		.INIT('h4)
	) name2193 (
		_w3372_,
		_w3373_,
		_w3374_
	);
	LUT2 #(
		.INIT('h8)
	) name2194 (
		\g185_reg/NET0131 ,
		\g2616_reg/NET0131 ,
		_w3375_
	);
	LUT3 #(
		.INIT('hb0)
	) name2195 (
		_w3372_,
		_w3373_,
		_w3375_,
		_w3376_
	);
	LUT2 #(
		.INIT('h8)
	) name2196 (
		\g1024_reg/NET0131 ,
		\g2676_reg/NET0131 ,
		_w3377_
	);
	LUT4 #(
		.INIT('h135f)
	) name2197 (
		\g1018_reg/NET0131 ,
		\g2670_reg/NET0131 ,
		\g2673_reg/NET0131 ,
		\g5657_pad ,
		_w3378_
	);
	LUT2 #(
		.INIT('h4)
	) name2198 (
		_w3377_,
		_w3378_,
		_w3379_
	);
	LUT2 #(
		.INIT('h4)
	) name2199 (
		_w3376_,
		_w3379_,
		_w3380_
	);
	LUT4 #(
		.INIT('h0400)
	) name2200 (
		_w3328_,
		_w3329_,
		_w3331_,
		_w3332_,
		_w3381_
	);
	LUT3 #(
		.INIT('h80)
	) name2201 (
		_w3323_,
		_w3364_,
		_w3381_,
		_w3382_
	);
	LUT4 #(
		.INIT('h0010)
	) name2202 (
		_w3369_,
		_w3371_,
		_w3380_,
		_w3382_,
		_w3383_
	);
	LUT3 #(
		.INIT('h80)
	) name2203 (
		_w3359_,
		_w3366_,
		_w3383_,
		_w3384_
	);
	LUT4 #(
		.INIT('hd1dd)
	) name2204 (
		_w3327_,
		_w3330_,
		_w3333_,
		_w3354_,
		_w3385_
	);
	LUT2 #(
		.INIT('h2)
	) name2205 (
		_w3338_,
		_w3385_,
		_w3386_
	);
	LUT4 #(
		.INIT('hb9fd)
	) name2206 (
		_w3323_,
		_w3333_,
		_w3338_,
		_w3370_,
		_w3387_
	);
	LUT4 #(
		.INIT('habef)
	) name2207 (
		_w3330_,
		_w3333_,
		_w3347_,
		_w3360_,
		_w3388_
	);
	LUT2 #(
		.INIT('h8)
	) name2208 (
		_w3335_,
		_w3363_,
		_w3389_
	);
	LUT4 #(
		.INIT('h00d0)
	) name2209 (
		_w3367_,
		_w3387_,
		_w3388_,
		_w3389_,
		_w3390_
	);
	LUT4 #(
		.INIT('h7aff)
	) name2210 (
		_w3323_,
		_w3334_,
		_w3350_,
		_w3364_,
		_w3391_
	);
	LUT3 #(
		.INIT('h80)
	) name2211 (
		_w3344_,
		_w3350_,
		_w3381_,
		_w3392_
	);
	LUT2 #(
		.INIT('h8)
	) name2212 (
		\g2643_reg/NET0131 ,
		\g5657_pad ,
		_w3393_
	);
	LUT4 #(
		.INIT('h135f)
	) name2213 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2645_reg/NET0131 ,
		\g2647_reg/NET0131 ,
		_w3394_
	);
	LUT2 #(
		.INIT('h4)
	) name2214 (
		_w3393_,
		_w3394_,
		_w3395_
	);
	LUT2 #(
		.INIT('h8)
	) name2215 (
		\g185_reg/NET0131 ,
		\g2598_reg/NET0131 ,
		_w3396_
	);
	LUT3 #(
		.INIT('hb0)
	) name2216 (
		_w3393_,
		_w3394_,
		_w3396_,
		_w3397_
	);
	LUT2 #(
		.INIT('h8)
	) name2217 (
		\g1024_reg/NET0131 ,
		\g2667_reg/NET0131 ,
		_w3398_
	);
	LUT4 #(
		.INIT('h135f)
	) name2218 (
		\g1018_reg/NET0131 ,
		\g2661_reg/NET0131 ,
		\g2664_reg/NET0131 ,
		\g5657_pad ,
		_w3399_
	);
	LUT2 #(
		.INIT('h4)
	) name2219 (
		_w3398_,
		_w3399_,
		_w3400_
	);
	LUT2 #(
		.INIT('h4)
	) name2220 (
		_w3397_,
		_w3400_,
		_w3401_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2221 (
		_w3376_,
		_w3379_,
		_w3397_,
		_w3400_,
		_w3402_
	);
	LUT3 #(
		.INIT('h02)
	) name2222 (
		_w3391_,
		_w3392_,
		_w3402_,
		_w3403_
	);
	LUT3 #(
		.INIT('h40)
	) name2223 (
		_w3386_,
		_w3390_,
		_w3403_,
		_w3404_
	);
	LUT3 #(
		.INIT('h80)
	) name2224 (
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		\g5657_pad ,
		_w3405_
	);
	LUT4 #(
		.INIT('h8000)
	) name2225 (
		_w3308_,
		_w3309_,
		_w3310_,
		_w3405_,
		_w3406_
	);
	LUT3 #(
		.INIT('h40)
	) name2226 (
		\g2688_reg/NET0131 ,
		\g5657_pad ,
		_w1418_,
		_w3407_
	);
	LUT2 #(
		.INIT('h1)
	) name2227 (
		\g2688_reg/NET0131 ,
		\g5657_pad ,
		_w3408_
	);
	LUT3 #(
		.INIT('h0b)
	) name2228 (
		_w3315_,
		_w3407_,
		_w3408_,
		_w3409_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2229 (
		_w3384_,
		_w3404_,
		_w3406_,
		_w3409_,
		_w3410_
	);
	LUT3 #(
		.INIT('h80)
	) name2230 (
		\g1018_reg/NET0131 ,
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		_w3411_
	);
	LUT4 #(
		.INIT('h8000)
	) name2231 (
		_w3308_,
		_w3309_,
		_w3310_,
		_w3411_,
		_w3412_
	);
	LUT3 #(
		.INIT('h20)
	) name2232 (
		\g1018_reg/NET0131 ,
		_w1417_,
		_w1418_,
		_w3413_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		\g1018_reg/NET0131 ,
		\g2691_reg/NET0131 ,
		_w3414_
	);
	LUT3 #(
		.INIT('h0b)
	) name2234 (
		_w3315_,
		_w3413_,
		_w3414_,
		_w3415_
	);
	LUT4 #(
		.INIT('h4f00)
	) name2235 (
		_w3384_,
		_w3404_,
		_w3412_,
		_w3415_,
		_w3416_
	);
	LUT3 #(
		.INIT('h20)
	) name2236 (
		\g1024_reg/NET0131 ,
		_w1417_,
		_w1418_,
		_w3417_
	);
	LUT2 #(
		.INIT('h1)
	) name2237 (
		\g1024_reg/NET0131 ,
		\g2694_reg/NET0131 ,
		_w3418_
	);
	LUT3 #(
		.INIT('h0b)
	) name2238 (
		_w3315_,
		_w3417_,
		_w3418_,
		_w3419_
	);
	LUT4 #(
		.INIT('h7500)
	) name2239 (
		_w3313_,
		_w3384_,
		_w3404_,
		_w3419_,
		_w3420_
	);
	LUT3 #(
		.INIT('h2a)
	) name2240 (
		_w1613_,
		_w2821_,
		_w2896_,
		_w3421_
	);
	LUT3 #(
		.INIT('h23)
	) name2241 (
		\g499_reg/NET0131 ,
		\g536_reg/NET0131 ,
		\g5657_pad ,
		_w3422_
	);
	LUT4 #(
		.INIT('h4000)
	) name2242 (
		_w2898_,
		_w2899_,
		_w3178_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h2)
	) name2243 (
		_w3180_,
		_w3423_,
		_w3424_
	);
	LUT3 #(
		.INIT('h70)
	) name2244 (
		_w2870_,
		_w3179_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('he)
	) name2245 (
		_w3421_,
		_w3425_,
		_w3426_
	);
	LUT3 #(
		.INIT('h23)
	) name2246 (
		\g499_reg/NET0131 ,
		\g537_reg/NET0131 ,
		\g5657_pad ,
		_w3427_
	);
	LUT4 #(
		.INIT('h4000)
	) name2247 (
		_w2898_,
		_w2899_,
		_w3178_,
		_w3427_,
		_w3428_
	);
	LUT4 #(
		.INIT('h00b0)
	) name2248 (
		_w2868_,
		_w3179_,
		_w3180_,
		_w3428_,
		_w3429_
	);
	LUT2 #(
		.INIT('h1)
	) name2249 (
		_w1613_,
		_w3429_,
		_w3430_
	);
	LUT2 #(
		.INIT('h2)
	) name2250 (
		_w2821_,
		_w3429_,
		_w3431_
	);
	LUT3 #(
		.INIT('h13)
	) name2251 (
		_w2895_,
		_w3430_,
		_w3431_,
		_w3432_
	);
	LUT4 #(
		.INIT('habaa)
	) name2252 (
		_w1504_,
		_w1509_,
		_w1510_,
		_w1511_,
		_w3433_
	);
	LUT2 #(
		.INIT('h1)
	) name2253 (
		\g2679_reg/NET0131 ,
		\g5657_pad ,
		_w3434_
	);
	LUT2 #(
		.INIT('h2)
	) name2254 (
		_w3391_,
		_w3392_,
		_w3435_
	);
	LUT3 #(
		.INIT('hd0)
	) name2255 (
		_w3338_,
		_w3385_,
		_w3401_,
		_w3436_
	);
	LUT3 #(
		.INIT('h80)
	) name2256 (
		_w3390_,
		_w3435_,
		_w3436_,
		_w3437_
	);
	LUT3 #(
		.INIT('h01)
	) name2257 (
		_w3369_,
		_w3371_,
		_w3382_,
		_w3438_
	);
	LUT2 #(
		.INIT('h2)
	) name2258 (
		_w3315_,
		_w3402_,
		_w3439_
	);
	LUT4 #(
		.INIT('h8000)
	) name2259 (
		_w3359_,
		_w3366_,
		_w3438_,
		_w3439_,
		_w3440_
	);
	LUT2 #(
		.INIT('h2)
	) name2260 (
		\g2679_reg/NET0131 ,
		\g5657_pad ,
		_w3441_
	);
	LUT3 #(
		.INIT('h0e)
	) name2261 (
		_w1459_,
		_w3315_,
		_w3441_,
		_w3442_
	);
	LUT4 #(
		.INIT('h1055)
	) name2262 (
		_w3434_,
		_w3437_,
		_w3440_,
		_w3442_,
		_w3443_
	);
	LUT2 #(
		.INIT('h1)
	) name2263 (
		\g1018_reg/NET0131 ,
		\g2682_reg/NET0131 ,
		_w3444_
	);
	LUT2 #(
		.INIT('h4)
	) name2264 (
		\g1018_reg/NET0131 ,
		\g2682_reg/NET0131 ,
		_w3445_
	);
	LUT3 #(
		.INIT('h0e)
	) name2265 (
		_w1459_,
		_w3315_,
		_w3445_,
		_w3446_
	);
	LUT4 #(
		.INIT('h040f)
	) name2266 (
		_w3437_,
		_w3440_,
		_w3444_,
		_w3446_,
		_w3447_
	);
	LUT2 #(
		.INIT('h1)
	) name2267 (
		\g1024_reg/NET0131 ,
		\g2685_reg/NET0131 ,
		_w3448_
	);
	LUT2 #(
		.INIT('h4)
	) name2268 (
		\g1024_reg/NET0131 ,
		\g2685_reg/NET0131 ,
		_w3449_
	);
	LUT3 #(
		.INIT('h0e)
	) name2269 (
		_w1459_,
		_w3315_,
		_w3449_,
		_w3450_
	);
	LUT4 #(
		.INIT('h040f)
	) name2270 (
		_w3437_,
		_w3440_,
		_w3448_,
		_w3450_,
		_w3451_
	);
	LUT2 #(
		.INIT('h4)
	) name2271 (
		_w1700_,
		_w2291_,
		_w3452_
	);
	LUT3 #(
		.INIT('h8c)
	) name2272 (
		_w1700_,
		_w1737_,
		_w2291_,
		_w3453_
	);
	LUT4 #(
		.INIT('h8000)
	) name2273 (
		_w1711_,
		_w1724_,
		_w1727_,
		_w1744_,
		_w3454_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2274 (
		_w1695_,
		_w1696_,
		_w1745_,
		_w1746_,
		_w3455_
	);
	LUT2 #(
		.INIT('h1)
	) name2275 (
		_w1700_,
		_w3455_,
		_w3456_
	);
	LUT2 #(
		.INIT('h8)
	) name2276 (
		_w3454_,
		_w3456_,
		_w3457_
	);
	LUT3 #(
		.INIT('h4f)
	) name2277 (
		_w2306_,
		_w3453_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h4)
	) name2278 (
		_w1364_,
		_w2474_,
		_w3459_
	);
	LUT3 #(
		.INIT('h20)
	) name2279 (
		_w1355_,
		_w1364_,
		_w2474_,
		_w3460_
	);
	LUT4 #(
		.INIT('h8000)
	) name2280 (
		_w1326_,
		_w1337_,
		_w1352_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h1)
	) name2281 (
		_w2470_,
		_w3461_,
		_w3462_
	);
	LUT2 #(
		.INIT('h2)
	) name2282 (
		_w1333_,
		_w3461_,
		_w3463_
	);
	LUT3 #(
		.INIT('hdc)
	) name2283 (
		_w2466_,
		_w3462_,
		_w3463_,
		_w3464_
	);
	LUT4 #(
		.INIT('h0400)
	) name2284 (
		_w1859_,
		_w1897_,
		_w1903_,
		_w1910_,
		_w3465_
	);
	LUT2 #(
		.INIT('h8)
	) name2285 (
		_w2337_,
		_w3465_,
		_w3466_
	);
	LUT2 #(
		.INIT('h8)
	) name2286 (
		_w1894_,
		_w3466_,
		_w3467_
	);
	LUT4 #(
		.INIT('h8000)
	) name2287 (
		_w1873_,
		_w1887_,
		_w1893_,
		_w3465_,
		_w3468_
	);
	LUT3 #(
		.INIT('h10)
	) name2288 (
		_w1975_,
		_w1978_,
		_w3468_,
		_w3469_
	);
	LUT4 #(
		.INIT('h0d0f)
	) name2289 (
		_w1851_,
		_w1950_,
		_w3467_,
		_w3469_,
		_w3470_
	);
	LUT3 #(
		.INIT('h02)
	) name2290 (
		_w2067_,
		_w2073_,
		_w2076_,
		_w3471_
	);
	LUT2 #(
		.INIT('h4)
	) name2291 (
		_w2121_,
		_w2435_,
		_w3472_
	);
	LUT4 #(
		.INIT('h8000)
	) name2292 (
		_w2054_,
		_w2064_,
		_w3471_,
		_w3472_,
		_w3473_
	);
	LUT4 #(
		.INIT('h00ef)
	) name2293 (
		_w2041_,
		_w2110_,
		_w2432_,
		_w3473_,
		_w3474_
	);
	LUT4 #(
		.INIT('h4000)
	) name2294 (
		\g1345_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2612_reg/NET0131 ,
		\g5657_pad ,
		_w3475_
	);
	LUT2 #(
		.INIT('h2)
	) name2295 (
		\g2809_reg/NET0131 ,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h2)
	) name2296 (
		\g1024_reg/NET0131 ,
		\g2802_reg/NET0131 ,
		_w3477_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2297 (
		\g1018_reg/NET0131 ,
		\g2803_reg/NET0131 ,
		\g2804_reg/NET0131 ,
		\g5657_pad ,
		_w3478_
	);
	LUT4 #(
		.INIT('h0400)
	) name2298 (
		_w1446_,
		_w1447_,
		_w3477_,
		_w3478_,
		_w3479_
	);
	LUT3 #(
		.INIT('h1d)
	) name2299 (
		\g2809_reg/NET0131 ,
		_w3475_,
		_w3479_,
		_w3480_
	);
	LUT3 #(
		.INIT('h45)
	) name2300 (
		\g1319_reg/NET0131 ,
		_w1449_,
		_w1450_,
		_w3481_
	);
	LUT3 #(
		.INIT('h8a)
	) name2301 (
		\g1339_reg/NET0131 ,
		\g2779_reg/NET0131 ,
		\g5657_pad ,
		_w3482_
	);
	LUT2 #(
		.INIT('h8)
	) name2302 (
		_w1424_,
		_w3482_,
		_w3483_
	);
	LUT3 #(
		.INIT('h45)
	) name2303 (
		\g1378_reg/NET0131 ,
		_w1451_,
		_w1452_,
		_w3484_
	);
	LUT3 #(
		.INIT('h45)
	) name2304 (
		\g1332_reg/NET0131 ,
		_w1437_,
		_w1438_,
		_w3485_
	);
	LUT4 #(
		.INIT('h0001)
	) name2305 (
		_w3481_,
		_w3483_,
		_w3484_,
		_w3485_,
		_w3486_
	);
	LUT3 #(
		.INIT('h45)
	) name2306 (
		\g1346_reg/NET0131 ,
		_w1431_,
		_w1432_,
		_w3487_
	);
	LUT3 #(
		.INIT('h45)
	) name2307 (
		\g1352_reg/NET0131 ,
		_w1426_,
		_w1427_,
		_w3488_
	);
	LUT3 #(
		.INIT('h8a)
	) name2308 (
		\g1352_reg/NET0131 ,
		\g2791_reg/NET0131 ,
		\g5657_pad ,
		_w3489_
	);
	LUT2 #(
		.INIT('h8)
	) name2309 (
		_w1427_,
		_w3489_,
		_w3490_
	);
	LUT3 #(
		.INIT('h45)
	) name2310 (
		\g1372_reg/NET0131 ,
		_w1420_,
		_w1421_,
		_w3491_
	);
	LUT4 #(
		.INIT('h0001)
	) name2311 (
		_w3487_,
		_w3488_,
		_w3490_,
		_w3491_,
		_w3492_
	);
	LUT3 #(
		.INIT('h45)
	) name2312 (
		\g1339_reg/NET0131 ,
		_w1423_,
		_w1424_,
		_w3493_
	);
	LUT3 #(
		.INIT('h8a)
	) name2313 (
		\g1365_reg/NET0131 ,
		\g2794_reg/NET0131 ,
		\g5657_pad ,
		_w3494_
	);
	LUT2 #(
		.INIT('h8)
	) name2314 (
		_w1435_,
		_w3494_,
		_w3495_
	);
	LUT3 #(
		.INIT('h8a)
	) name2315 (
		\g1372_reg/NET0131 ,
		\g2797_reg/NET0131 ,
		\g5657_pad ,
		_w3496_
	);
	LUT3 #(
		.INIT('h8a)
	) name2316 (
		\g1378_reg/NET0131 ,
		\g2800_reg/NET0131 ,
		\g5657_pad ,
		_w3497_
	);
	LUT4 #(
		.INIT('h135f)
	) name2317 (
		_w1421_,
		_w1452_,
		_w3496_,
		_w3497_,
		_w3498_
	);
	LUT3 #(
		.INIT('h45)
	) name2318 (
		\g1326_reg/NET0131 ,
		_w1440_,
		_w1441_,
		_w3499_
	);
	LUT4 #(
		.INIT('h0010)
	) name2319 (
		_w3493_,
		_w3495_,
		_w3498_,
		_w3499_,
		_w3500_
	);
	LUT3 #(
		.INIT('h45)
	) name2320 (
		\g1365_reg/NET0131 ,
		_w1434_,
		_w1435_,
		_w3501_
	);
	LUT3 #(
		.INIT('h45)
	) name2321 (
		\g1358_reg/NET0131 ,
		_w1429_,
		_w1430_,
		_w3502_
	);
	LUT3 #(
		.INIT('h8a)
	) name2322 (
		\g1319_reg/NET0131 ,
		\g2776_reg/NET0131 ,
		\g5657_pad ,
		_w3503_
	);
	LUT3 #(
		.INIT('h8a)
	) name2323 (
		\g1332_reg/NET0131 ,
		\g2782_reg/NET0131 ,
		\g5657_pad ,
		_w3504_
	);
	LUT4 #(
		.INIT('h153f)
	) name2324 (
		_w1438_,
		_w1450_,
		_w3503_,
		_w3504_,
		_w3505_
	);
	LUT3 #(
		.INIT('h8a)
	) name2325 (
		\g1346_reg/NET0131 ,
		\g2785_reg/NET0131 ,
		\g5657_pad ,
		_w3506_
	);
	LUT2 #(
		.INIT('h8)
	) name2326 (
		_w1432_,
		_w3506_,
		_w3507_
	);
	LUT4 #(
		.INIT('h0010)
	) name2327 (
		_w3501_,
		_w3502_,
		_w3505_,
		_w3507_,
		_w3508_
	);
	LUT4 #(
		.INIT('h8000)
	) name2328 (
		_w3486_,
		_w3492_,
		_w3500_,
		_w3508_,
		_w3509_
	);
	LUT3 #(
		.INIT('h8a)
	) name2329 (
		\g1358_reg/NET0131 ,
		\g2788_reg/NET0131 ,
		\g5657_pad ,
		_w3510_
	);
	LUT3 #(
		.INIT('h8a)
	) name2330 (
		\g1326_reg/NET0131 ,
		\g2773_reg/NET0131 ,
		\g5657_pad ,
		_w3511_
	);
	LUT4 #(
		.INIT('h135f)
	) name2331 (
		_w1430_,
		_w1441_,
		_w3510_,
		_w3511_,
		_w3512_
	);
	LUT2 #(
		.INIT('h4)
	) name2332 (
		_w3476_,
		_w3512_,
		_w3513_
	);
	LUT3 #(
		.INIT('h15)
	) name2333 (
		_w3480_,
		_w3509_,
		_w3513_,
		_w3514_
	);
	LUT4 #(
		.INIT('h2000)
	) name2334 (
		\g1018_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2612_reg/NET0131 ,
		_w3515_
	);
	LUT2 #(
		.INIT('h2)
	) name2335 (
		\g2810_reg/NET0131 ,
		_w3515_,
		_w3516_
	);
	LUT3 #(
		.INIT('h35)
	) name2336 (
		\g2810_reg/NET0131 ,
		_w3479_,
		_w3515_,
		_w3517_
	);
	LUT2 #(
		.INIT('h2)
	) name2337 (
		_w3512_,
		_w3516_,
		_w3518_
	);
	LUT3 #(
		.INIT('h13)
	) name2338 (
		_w3509_,
		_w3517_,
		_w3518_,
		_w3519_
	);
	LUT2 #(
		.INIT('h8)
	) name2339 (
		\g1211_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		_w3520_
	);
	LUT2 #(
		.INIT('h2)
	) name2340 (
		\g1024_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w3521_
	);
	LUT4 #(
		.INIT('h0080)
	) name2341 (
		\g1024_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w3522_
	);
	LUT2 #(
		.INIT('h2)
	) name2342 (
		\g1420_reg/NET0131 ,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h2)
	) name2343 (
		\g1024_reg/NET0131 ,
		\g1414_reg/NET0131 ,
		_w3524_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2344 (
		\g1018_reg/NET0131 ,
		\g1415_reg/NET0131 ,
		\g1416_reg/NET0131 ,
		\g5657_pad ,
		_w3525_
	);
	LUT4 #(
		.INIT('h0400)
	) name2345 (
		_w2172_,
		_w2173_,
		_w3524_,
		_w3525_,
		_w3526_
	);
	LUT3 #(
		.INIT('h1d)
	) name2346 (
		\g1420_reg/NET0131 ,
		_w3522_,
		_w3526_,
		_w3527_
	);
	LUT3 #(
		.INIT('h45)
	) name2347 (
		\g1346_reg/NET0131 ,
		_w2185_,
		_w2186_,
		_w3528_
	);
	LUT3 #(
		.INIT('h8a)
	) name2348 (
		\g1319_reg/NET0131 ,
		\g1388_reg/NET0131 ,
		\g5657_pad ,
		_w3529_
	);
	LUT2 #(
		.INIT('h8)
	) name2349 (
		_w2191_,
		_w3529_,
		_w3530_
	);
	LUT3 #(
		.INIT('h45)
	) name2350 (
		\g1332_reg/NET0131 ,
		_w2195_,
		_w2196_,
		_w3531_
	);
	LUT3 #(
		.INIT('h45)
	) name2351 (
		\g1358_reg/NET0131 ,
		_w2178_,
		_w2179_,
		_w3532_
	);
	LUT4 #(
		.INIT('h0001)
	) name2352 (
		_w3528_,
		_w3530_,
		_w3531_,
		_w3532_,
		_w3533_
	);
	LUT3 #(
		.INIT('h45)
	) name2353 (
		\g1339_reg/NET0131 ,
		_w2175_,
		_w2176_,
		_w3534_
	);
	LUT3 #(
		.INIT('h45)
	) name2354 (
		\g1372_reg/NET0131 ,
		_w2182_,
		_w2183_,
		_w3535_
	);
	LUT3 #(
		.INIT('h8a)
	) name2355 (
		\g1372_reg/NET0131 ,
		\g1409_reg/NET0131 ,
		\g5657_pad ,
		_w3536_
	);
	LUT2 #(
		.INIT('h8)
	) name2356 (
		_w2183_,
		_w3536_,
		_w3537_
	);
	LUT3 #(
		.INIT('h45)
	) name2357 (
		\g1365_reg/NET0131 ,
		_w2202_,
		_w2203_,
		_w3538_
	);
	LUT4 #(
		.INIT('h0001)
	) name2358 (
		_w3534_,
		_w3535_,
		_w3537_,
		_w3538_,
		_w3539_
	);
	LUT3 #(
		.INIT('h45)
	) name2359 (
		\g1319_reg/NET0131 ,
		_w2190_,
		_w2191_,
		_w3540_
	);
	LUT3 #(
		.INIT('h8a)
	) name2360 (
		\g1378_reg/NET0131 ,
		\g1412_reg/NET0131 ,
		\g5657_pad ,
		_w3541_
	);
	LUT2 #(
		.INIT('h8)
	) name2361 (
		_w2200_,
		_w3541_,
		_w3542_
	);
	LUT3 #(
		.INIT('h8a)
	) name2362 (
		\g1365_reg/NET0131 ,
		\g1406_reg/NET0131 ,
		\g5657_pad ,
		_w3543_
	);
	LUT3 #(
		.INIT('h8a)
	) name2363 (
		\g1332_reg/NET0131 ,
		\g1394_reg/NET0131 ,
		\g5657_pad ,
		_w3544_
	);
	LUT4 #(
		.INIT('h153f)
	) name2364 (
		_w2196_,
		_w2203_,
		_w3543_,
		_w3544_,
		_w3545_
	);
	LUT3 #(
		.INIT('h45)
	) name2365 (
		\g1326_reg/NET0131 ,
		_w2188_,
		_w2189_,
		_w3546_
	);
	LUT4 #(
		.INIT('h0010)
	) name2366 (
		_w3540_,
		_w3542_,
		_w3545_,
		_w3546_,
		_w3547_
	);
	LUT3 #(
		.INIT('h45)
	) name2367 (
		\g1378_reg/NET0131 ,
		_w2199_,
		_w2200_,
		_w3548_
	);
	LUT3 #(
		.INIT('h45)
	) name2368 (
		\g1352_reg/NET0131 ,
		_w2193_,
		_w2194_,
		_w3549_
	);
	LUT3 #(
		.INIT('h8a)
	) name2369 (
		\g1346_reg/NET0131 ,
		\g1397_reg/NET0131 ,
		\g5657_pad ,
		_w3550_
	);
	LUT3 #(
		.INIT('h8a)
	) name2370 (
		\g1358_reg/NET0131 ,
		\g1400_reg/NET0131 ,
		\g5657_pad ,
		_w3551_
	);
	LUT4 #(
		.INIT('h153f)
	) name2371 (
		_w2179_,
		_w2186_,
		_w3550_,
		_w3551_,
		_w3552_
	);
	LUT3 #(
		.INIT('h8a)
	) name2372 (
		\g1339_reg/NET0131 ,
		\g1391_reg/NET0131 ,
		\g5657_pad ,
		_w3553_
	);
	LUT2 #(
		.INIT('h8)
	) name2373 (
		_w2176_,
		_w3553_,
		_w3554_
	);
	LUT4 #(
		.INIT('h0010)
	) name2374 (
		_w3548_,
		_w3549_,
		_w3552_,
		_w3554_,
		_w3555_
	);
	LUT4 #(
		.INIT('h8000)
	) name2375 (
		_w3533_,
		_w3539_,
		_w3547_,
		_w3555_,
		_w3556_
	);
	LUT3 #(
		.INIT('h8a)
	) name2376 (
		\g1352_reg/NET0131 ,
		\g1403_reg/NET0131 ,
		\g5657_pad ,
		_w3557_
	);
	LUT3 #(
		.INIT('h8a)
	) name2377 (
		\g1326_reg/NET0131 ,
		\g1385_reg/NET0131 ,
		\g5657_pad ,
		_w3558_
	);
	LUT4 #(
		.INIT('h153f)
	) name2378 (
		_w2189_,
		_w2194_,
		_w3557_,
		_w3558_,
		_w3559_
	);
	LUT2 #(
		.INIT('h4)
	) name2379 (
		_w3523_,
		_w3559_,
		_w3560_
	);
	LUT3 #(
		.INIT('h15)
	) name2380 (
		_w3527_,
		_w3556_,
		_w3560_,
		_w3561_
	);
	LUT4 #(
		.INIT('h0080)
	) name2381 (
		\g1018_reg/NET0131 ,
		\g1211_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w3562_
	);
	LUT2 #(
		.INIT('h2)
	) name2382 (
		\g1422_reg/NET0131 ,
		_w3562_,
		_w3563_
	);
	LUT3 #(
		.INIT('h35)
	) name2383 (
		\g1422_reg/NET0131 ,
		_w3526_,
		_w3562_,
		_w3564_
	);
	LUT2 #(
		.INIT('h2)
	) name2384 (
		_w3559_,
		_w3563_,
		_w3565_
	);
	LUT3 #(
		.INIT('h13)
	) name2385 (
		_w3556_,
		_w3564_,
		_w3565_,
		_w3566_
	);
	LUT4 #(
		.INIT('h0800)
	) name2386 (
		\g1211_reg/NET0131 ,
		\g1224_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g5657_pad ,
		_w3567_
	);
	LUT2 #(
		.INIT('h2)
	) name2387 (
		\g1421_reg/NET0131 ,
		_w3567_,
		_w3568_
	);
	LUT3 #(
		.INIT('h35)
	) name2388 (
		\g1421_reg/NET0131 ,
		_w3526_,
		_w3567_,
		_w3569_
	);
	LUT2 #(
		.INIT('h2)
	) name2389 (
		_w3559_,
		_w3568_,
		_w3570_
	);
	LUT3 #(
		.INIT('h13)
	) name2390 (
		_w3556_,
		_w3569_,
		_w3570_,
		_w3571_
	);
	LUT4 #(
		.INIT('h2000)
	) name2391 (
		\g1024_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1918_reg/NET0131 ,
		_w3572_
	);
	LUT2 #(
		.INIT('h2)
	) name2392 (
		\g2114_reg/NET0131 ,
		_w3572_,
		_w3573_
	);
	LUT2 #(
		.INIT('h2)
	) name2393 (
		\g1024_reg/NET0131 ,
		\g2108_reg/NET0131 ,
		_w3574_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2394 (
		\g1018_reg/NET0131 ,
		\g2109_reg/NET0131 ,
		\g2110_reg/NET0131 ,
		\g5657_pad ,
		_w3575_
	);
	LUT4 #(
		.INIT('h0400)
	) name2395 (
		_w1537_,
		_w1538_,
		_w3574_,
		_w3575_,
		_w3576_
	);
	LUT3 #(
		.INIT('h1d)
	) name2396 (
		\g2114_reg/NET0131 ,
		_w3572_,
		_w3576_,
		_w3577_
	);
	LUT3 #(
		.INIT('h45)
	) name2397 (
		\g1346_reg/NET0131 ,
		_w1554_,
		_w1555_,
		_w3578_
	);
	LUT3 #(
		.INIT('h8a)
	) name2398 (
		\g1319_reg/NET0131 ,
		\g2082_reg/NET0131 ,
		\g5657_pad ,
		_w3579_
	);
	LUT2 #(
		.INIT('h8)
	) name2399 (
		_w1561_,
		_w3579_,
		_w3580_
	);
	LUT3 #(
		.INIT('h45)
	) name2400 (
		\g1358_reg/NET0131 ,
		_w1549_,
		_w1550_,
		_w3581_
	);
	LUT3 #(
		.INIT('h45)
	) name2401 (
		\g1332_reg/NET0131 ,
		_w1557_,
		_w1558_,
		_w3582_
	);
	LUT4 #(
		.INIT('h0001)
	) name2402 (
		_w3578_,
		_w3580_,
		_w3581_,
		_w3582_,
		_w3583_
	);
	LUT3 #(
		.INIT('h45)
	) name2403 (
		\g1339_reg/NET0131 ,
		_w1564_,
		_w1565_,
		_w3584_
	);
	LUT3 #(
		.INIT('h45)
	) name2404 (
		\g1378_reg/NET0131 ,
		_w1567_,
		_w1568_,
		_w3585_
	);
	LUT3 #(
		.INIT('h8a)
	) name2405 (
		\g1378_reg/NET0131 ,
		\g2106_reg/NET0131 ,
		\g5657_pad ,
		_w3586_
	);
	LUT2 #(
		.INIT('h8)
	) name2406 (
		_w1568_,
		_w3586_,
		_w3587_
	);
	LUT3 #(
		.INIT('h45)
	) name2407 (
		\g1372_reg/NET0131 ,
		_w1546_,
		_w1547_,
		_w3588_
	);
	LUT4 #(
		.INIT('h0001)
	) name2408 (
		_w3584_,
		_w3585_,
		_w3587_,
		_w3588_,
		_w3589_
	);
	LUT3 #(
		.INIT('h45)
	) name2409 (
		\g1319_reg/NET0131 ,
		_w1560_,
		_w1561_,
		_w3590_
	);
	LUT3 #(
		.INIT('h8a)
	) name2410 (
		\g1352_reg/NET0131 ,
		\g2097_reg/NET0131 ,
		\g5657_pad ,
		_w3591_
	);
	LUT2 #(
		.INIT('h8)
	) name2411 (
		_w1541_,
		_w3591_,
		_w3592_
	);
	LUT3 #(
		.INIT('h8a)
	) name2412 (
		\g1372_reg/NET0131 ,
		\g2103_reg/NET0131 ,
		\g5657_pad ,
		_w3593_
	);
	LUT3 #(
		.INIT('h8a)
	) name2413 (
		\g1358_reg/NET0131 ,
		\g2094_reg/NET0131 ,
		\g5657_pad ,
		_w3594_
	);
	LUT4 #(
		.INIT('h135f)
	) name2414 (
		_w1547_,
		_w1550_,
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT3 #(
		.INIT('h45)
	) name2415 (
		\g1326_reg/NET0131 ,
		_w1552_,
		_w1553_,
		_w3596_
	);
	LUT4 #(
		.INIT('h0010)
	) name2416 (
		_w3590_,
		_w3592_,
		_w3595_,
		_w3596_,
		_w3597_
	);
	LUT3 #(
		.INIT('h45)
	) name2417 (
		\g1352_reg/NET0131 ,
		_w1540_,
		_w1541_,
		_w3598_
	);
	LUT3 #(
		.INIT('h45)
	) name2418 (
		\g1365_reg/NET0131 ,
		_w1535_,
		_w1536_,
		_w3599_
	);
	LUT3 #(
		.INIT('h8a)
	) name2419 (
		\g1346_reg/NET0131 ,
		\g2091_reg/NET0131 ,
		\g5657_pad ,
		_w3600_
	);
	LUT3 #(
		.INIT('h8a)
	) name2420 (
		\g1332_reg/NET0131 ,
		\g2088_reg/NET0131 ,
		\g5657_pad ,
		_w3601_
	);
	LUT4 #(
		.INIT('h135f)
	) name2421 (
		_w1555_,
		_w1558_,
		_w3600_,
		_w3601_,
		_w3602_
	);
	LUT3 #(
		.INIT('h8a)
	) name2422 (
		\g1339_reg/NET0131 ,
		\g2085_reg/NET0131 ,
		\g5657_pad ,
		_w3603_
	);
	LUT2 #(
		.INIT('h8)
	) name2423 (
		_w1565_,
		_w3603_,
		_w3604_
	);
	LUT4 #(
		.INIT('h0010)
	) name2424 (
		_w3598_,
		_w3599_,
		_w3602_,
		_w3604_,
		_w3605_
	);
	LUT4 #(
		.INIT('h8000)
	) name2425 (
		_w3583_,
		_w3589_,
		_w3597_,
		_w3605_,
		_w3606_
	);
	LUT3 #(
		.INIT('h8a)
	) name2426 (
		\g1365_reg/NET0131 ,
		\g2100_reg/NET0131 ,
		\g5657_pad ,
		_w3607_
	);
	LUT3 #(
		.INIT('h8a)
	) name2427 (
		\g1326_reg/NET0131 ,
		\g2079_reg/NET0131 ,
		\g5657_pad ,
		_w3608_
	);
	LUT4 #(
		.INIT('h135f)
	) name2428 (
		_w1536_,
		_w1553_,
		_w3607_,
		_w3608_,
		_w3609_
	);
	LUT2 #(
		.INIT('h4)
	) name2429 (
		_w3573_,
		_w3609_,
		_w3610_
	);
	LUT3 #(
		.INIT('h15)
	) name2430 (
		_w3577_,
		_w3606_,
		_w3610_,
		_w3611_
	);
	LUT4 #(
		.INIT('h2000)
	) name2431 (
		\g1024_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g525_reg/NET0131 ,
		\g538_reg/NET0131 ,
		_w3612_
	);
	LUT2 #(
		.INIT('h2)
	) name2432 (
		\g734_reg/NET0131 ,
		_w3612_,
		_w3613_
	);
	LUT2 #(
		.INIT('h2)
	) name2433 (
		\g1024_reg/NET0131 ,
		\g728_reg/NET0131 ,
		_w3614_
	);
	LUT4 #(
		.INIT('hf351)
	) name2434 (
		\g1018_reg/NET0131 ,
		\g5657_pad ,
		\g729_reg/NET0131 ,
		\g730_reg/NET0131 ,
		_w3615_
	);
	LUT4 #(
		.INIT('h0400)
	) name2435 (
		_w2850_,
		_w2851_,
		_w3614_,
		_w3615_,
		_w3616_
	);
	LUT3 #(
		.INIT('h1d)
	) name2436 (
		\g734_reg/NET0131 ,
		_w3612_,
		_w3616_,
		_w3617_
	);
	LUT3 #(
		.INIT('h45)
	) name2437 (
		\g1326_reg/NET0131 ,
		_w2844_,
		_w2845_,
		_w3618_
	);
	LUT3 #(
		.INIT('ha2)
	) name2438 (
		\g1319_reg/NET0131 ,
		\g5657_pad ,
		\g702_reg/NET0131 ,
		_w3619_
	);
	LUT2 #(
		.INIT('h8)
	) name2439 (
		_w2838_,
		_w3619_,
		_w3620_
	);
	LUT3 #(
		.INIT('h45)
	) name2440 (
		\g1358_reg/NET0131 ,
		_w2825_,
		_w2826_,
		_w3621_
	);
	LUT3 #(
		.INIT('h45)
	) name2441 (
		\g1352_reg/NET0131 ,
		_w2855_,
		_w2856_,
		_w3622_
	);
	LUT4 #(
		.INIT('h0001)
	) name2442 (
		_w3618_,
		_w3620_,
		_w3621_,
		_w3622_,
		_w3623_
	);
	LUT3 #(
		.INIT('h45)
	) name2443 (
		\g1339_reg/NET0131 ,
		_w2822_,
		_w2823_,
		_w3624_
	);
	LUT3 #(
		.INIT('h45)
	) name2444 (
		\g1378_reg/NET0131 ,
		_w2847_,
		_w2848_,
		_w3625_
	);
	LUT3 #(
		.INIT('ha2)
	) name2445 (
		\g1378_reg/NET0131 ,
		\g5657_pad ,
		\g726_reg/NET0131 ,
		_w3626_
	);
	LUT2 #(
		.INIT('h8)
	) name2446 (
		_w2848_,
		_w3626_,
		_w3627_
	);
	LUT3 #(
		.INIT('h45)
	) name2447 (
		\g1372_reg/NET0131 ,
		_w2834_,
		_w2835_,
		_w3628_
	);
	LUT4 #(
		.INIT('h0001)
	) name2448 (
		_w3624_,
		_w3625_,
		_w3627_,
		_w3628_,
		_w3629_
	);
	LUT3 #(
		.INIT('h45)
	) name2449 (
		\g1319_reg/NET0131 ,
		_w2837_,
		_w2838_,
		_w3630_
	);
	LUT3 #(
		.INIT('ha2)
	) name2450 (
		\g1332_reg/NET0131 ,
		\g5657_pad ,
		\g708_reg/NET0131 ,
		_w3631_
	);
	LUT2 #(
		.INIT('h8)
	) name2451 (
		_w2842_,
		_w3631_,
		_w3632_
	);
	LUT3 #(
		.INIT('ha2)
	) name2452 (
		\g1372_reg/NET0131 ,
		\g5657_pad ,
		\g723_reg/NET0131 ,
		_w3633_
	);
	LUT3 #(
		.INIT('ha2)
	) name2453 (
		\g1358_reg/NET0131 ,
		\g5657_pad ,
		\g714_reg/NET0131 ,
		_w3634_
	);
	LUT4 #(
		.INIT('h153f)
	) name2454 (
		_w2826_,
		_w2835_,
		_w3633_,
		_w3634_,
		_w3635_
	);
	LUT3 #(
		.INIT('h45)
	) name2455 (
		\g1346_reg/NET0131 ,
		_w2853_,
		_w2854_,
		_w3636_
	);
	LUT4 #(
		.INIT('h0010)
	) name2456 (
		_w3630_,
		_w3632_,
		_w3635_,
		_w3636_,
		_w3637_
	);
	LUT3 #(
		.INIT('h45)
	) name2457 (
		\g1332_reg/NET0131 ,
		_w2841_,
		_w2842_,
		_w3638_
	);
	LUT3 #(
		.INIT('h45)
	) name2458 (
		\g1365_reg/NET0131 ,
		_w2828_,
		_w2829_,
		_w3639_
	);
	LUT3 #(
		.INIT('ha2)
	) name2459 (
		\g1326_reg/NET0131 ,
		\g5657_pad ,
		\g699_reg/NET0131 ,
		_w3640_
	);
	LUT3 #(
		.INIT('ha2)
	) name2460 (
		\g1352_reg/NET0131 ,
		\g5657_pad ,
		\g717_reg/NET0131 ,
		_w3641_
	);
	LUT4 #(
		.INIT('h135f)
	) name2461 (
		_w2845_,
		_w2856_,
		_w3640_,
		_w3641_,
		_w3642_
	);
	LUT3 #(
		.INIT('ha2)
	) name2462 (
		\g1339_reg/NET0131 ,
		\g5657_pad ,
		\g705_reg/NET0131 ,
		_w3643_
	);
	LUT2 #(
		.INIT('h8)
	) name2463 (
		_w2823_,
		_w3643_,
		_w3644_
	);
	LUT4 #(
		.INIT('h0010)
	) name2464 (
		_w3638_,
		_w3639_,
		_w3642_,
		_w3644_,
		_w3645_
	);
	LUT4 #(
		.INIT('h8000)
	) name2465 (
		_w3623_,
		_w3629_,
		_w3637_,
		_w3645_,
		_w3646_
	);
	LUT3 #(
		.INIT('ha2)
	) name2466 (
		\g1365_reg/NET0131 ,
		\g5657_pad ,
		\g720_reg/NET0131 ,
		_w3647_
	);
	LUT3 #(
		.INIT('ha2)
	) name2467 (
		\g1346_reg/NET0131 ,
		\g5657_pad ,
		\g711_reg/NET0131 ,
		_w3648_
	);
	LUT4 #(
		.INIT('h135f)
	) name2468 (
		_w2829_,
		_w2854_,
		_w3647_,
		_w3648_,
		_w3649_
	);
	LUT2 #(
		.INIT('h4)
	) name2469 (
		_w3613_,
		_w3649_,
		_w3650_
	);
	LUT3 #(
		.INIT('h15)
	) name2470 (
		_w3617_,
		_w3646_,
		_w3650_,
		_w3651_
	);
	LUT4 #(
		.INIT('h4000)
	) name2471 (
		\g1345_reg/NET0131 ,
		\g525_reg/NET0131 ,
		\g538_reg/NET0131 ,
		\g5657_pad ,
		_w3652_
	);
	LUT2 #(
		.INIT('h2)
	) name2472 (
		\g735_reg/NET0131 ,
		_w3652_,
		_w3653_
	);
	LUT3 #(
		.INIT('h35)
	) name2473 (
		\g735_reg/NET0131 ,
		_w3616_,
		_w3652_,
		_w3654_
	);
	LUT2 #(
		.INIT('h2)
	) name2474 (
		_w3649_,
		_w3653_,
		_w3655_
	);
	LUT3 #(
		.INIT('h13)
	) name2475 (
		_w3646_,
		_w3654_,
		_w3655_,
		_w3656_
	);
	LUT4 #(
		.INIT('h2000)
	) name2476 (
		\g1018_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g525_reg/NET0131 ,
		\g538_reg/NET0131 ,
		_w3657_
	);
	LUT2 #(
		.INIT('h2)
	) name2477 (
		\g736_reg/NET0131 ,
		_w3657_,
		_w3658_
	);
	LUT3 #(
		.INIT('h35)
	) name2478 (
		\g736_reg/NET0131 ,
		_w3616_,
		_w3657_,
		_w3659_
	);
	LUT2 #(
		.INIT('h2)
	) name2479 (
		_w3649_,
		_w3658_,
		_w3660_
	);
	LUT3 #(
		.INIT('h13)
	) name2480 (
		_w3646_,
		_w3659_,
		_w3660_,
		_w3661_
	);
	LUT4 #(
		.INIT('h2000)
	) name2481 (
		\g1018_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1918_reg/NET0131 ,
		_w3662_
	);
	LUT2 #(
		.INIT('h2)
	) name2482 (
		\g2116_reg/NET0131 ,
		_w3662_,
		_w3663_
	);
	LUT3 #(
		.INIT('h35)
	) name2483 (
		\g2116_reg/NET0131 ,
		_w3576_,
		_w3662_,
		_w3664_
	);
	LUT2 #(
		.INIT('h2)
	) name2484 (
		_w3609_,
		_w3663_,
		_w3665_
	);
	LUT3 #(
		.INIT('h13)
	) name2485 (
		_w3606_,
		_w3664_,
		_w3665_,
		_w3666_
	);
	LUT4 #(
		.INIT('h4000)
	) name2486 (
		\g1345_reg/NET0131 ,
		\g1905_reg/NET0131 ,
		\g1918_reg/NET0131 ,
		\g5657_pad ,
		_w3667_
	);
	LUT2 #(
		.INIT('h2)
	) name2487 (
		\g2115_reg/NET0131 ,
		_w3667_,
		_w3668_
	);
	LUT3 #(
		.INIT('h35)
	) name2488 (
		\g2115_reg/NET0131 ,
		_w3576_,
		_w3667_,
		_w3669_
	);
	LUT2 #(
		.INIT('h2)
	) name2489 (
		_w3609_,
		_w3668_,
		_w3670_
	);
	LUT3 #(
		.INIT('h13)
	) name2490 (
		_w3606_,
		_w3669_,
		_w3670_,
		_w3671_
	);
	LUT4 #(
		.INIT('h2000)
	) name2491 (
		\g1024_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g2599_reg/NET0131 ,
		\g2612_reg/NET0131 ,
		_w3672_
	);
	LUT2 #(
		.INIT('h2)
	) name2492 (
		\g2808_reg/NET0131 ,
		_w3672_,
		_w3673_
	);
	LUT3 #(
		.INIT('h35)
	) name2493 (
		\g2808_reg/NET0131 ,
		_w3479_,
		_w3672_,
		_w3674_
	);
	LUT2 #(
		.INIT('h2)
	) name2494 (
		_w3512_,
		_w3673_,
		_w3675_
	);
	LUT3 #(
		.INIT('h13)
	) name2495 (
		_w3509_,
		_w3674_,
		_w3675_,
		_w3676_
	);
	LUT2 #(
		.INIT('h1)
	) name2496 (
		_w1578_,
		_w3315_,
		_w3677_
	);
	LUT2 #(
		.INIT('h8)
	) name2497 (
		\g1018_reg/NET0131 ,
		\g1747_reg/NET0131 ,
		_w3678_
	);
	LUT4 #(
		.INIT('h135f)
	) name2498 (
		\g1024_reg/NET0131 ,
		\g1745_reg/NET0131 ,
		\g1749_reg/NET0131 ,
		\g5657_pad ,
		_w3679_
	);
	LUT2 #(
		.INIT('h4)
	) name2499 (
		_w3678_,
		_w3679_,
		_w3680_
	);
	LUT2 #(
		.INIT('h8)
	) name2500 (
		\g1018_reg/NET0131 ,
		\g1762_reg/NET0131 ,
		_w3681_
	);
	LUT4 #(
		.INIT('h135f)
	) name2501 (
		\g1024_reg/NET0131 ,
		\g1760_reg/NET0131 ,
		\g1764_reg/NET0131 ,
		\g5657_pad ,
		_w3682_
	);
	LUT2 #(
		.INIT('h4)
	) name2502 (
		_w3681_,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h8)
	) name2503 (
		\g1018_reg/NET0131 ,
		\g1732_reg/NET0131 ,
		_w3684_
	);
	LUT4 #(
		.INIT('h135f)
	) name2504 (
		\g1024_reg/NET0131 ,
		\g1730_reg/NET0131 ,
		\g1734_reg/NET0131 ,
		\g5657_pad ,
		_w3685_
	);
	LUT2 #(
		.INIT('h4)
	) name2505 (
		_w3684_,
		_w3685_,
		_w3686_
	);
	LUT4 #(
		.INIT('h0400)
	) name2506 (
		_w3681_,
		_w3682_,
		_w3684_,
		_w3685_,
		_w3687_
	);
	LUT2 #(
		.INIT('h4)
	) name2507 (
		\g1959_reg/NET0131 ,
		\g5657_pad ,
		_w3688_
	);
	LUT4 #(
		.INIT('hf351)
	) name2508 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1958_reg/NET0131 ,
		\g1960_reg/NET0131 ,
		_w3689_
	);
	LUT2 #(
		.INIT('h4)
	) name2509 (
		_w3688_,
		_w3689_,
		_w3690_
	);
	LUT2 #(
		.INIT('h2)
	) name2510 (
		\g1024_reg/NET0131 ,
		\g1961_reg/NET0131 ,
		_w3691_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2511 (
		\g1018_reg/NET0131 ,
		\g1962_reg/NET0131 ,
		\g1963_reg/NET0131 ,
		\g5657_pad ,
		_w3692_
	);
	LUT2 #(
		.INIT('h4)
	) name2512 (
		_w3691_,
		_w3692_,
		_w3693_
	);
	LUT4 #(
		.INIT('h0400)
	) name2513 (
		_w3688_,
		_w3689_,
		_w3691_,
		_w3692_,
		_w3694_
	);
	LUT2 #(
		.INIT('h8)
	) name2514 (
		_w3687_,
		_w3694_,
		_w3695_
	);
	LUT4 #(
		.INIT('h4044)
	) name2515 (
		_w3681_,
		_w3682_,
		_w3684_,
		_w3685_,
		_w3696_
	);
	LUT2 #(
		.INIT('h4)
	) name2516 (
		\g1956_reg/NET0131 ,
		\g5657_pad ,
		_w3697_
	);
	LUT4 #(
		.INIT('hf351)
	) name2517 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1955_reg/NET0131 ,
		\g1957_reg/NET0131 ,
		_w3698_
	);
	LUT2 #(
		.INIT('h4)
	) name2518 (
		_w3697_,
		_w3698_,
		_w3699_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2519 (
		_w3691_,
		_w3692_,
		_w3697_,
		_w3698_,
		_w3700_
	);
	LUT4 #(
		.INIT('hecfd)
	) name2520 (
		_w3683_,
		_w3686_,
		_w3690_,
		_w3700_,
		_w3701_
	);
	LUT3 #(
		.INIT('h45)
	) name2521 (
		_w3680_,
		_w3695_,
		_w3701_,
		_w3702_
	);
	LUT4 #(
		.INIT('h0400)
	) name2522 (
		_w3688_,
		_w3689_,
		_w3697_,
		_w3698_,
		_w3703_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2523 (
		_w3678_,
		_w3679_,
		_w3681_,
		_w3682_,
		_w3704_
	);
	LUT3 #(
		.INIT('h80)
	) name2524 (
		_w3686_,
		_w3703_,
		_w3704_,
		_w3705_
	);
	LUT2 #(
		.INIT('h8)
	) name2525 (
		\g1018_reg/NET0131 ,
		\g1777_reg/NET0131 ,
		_w3706_
	);
	LUT4 #(
		.INIT('h0777)
	) name2526 (
		\g1024_reg/NET0131 ,
		\g1705_reg/NET0131 ,
		\g1775_reg/NET0131 ,
		\g5657_pad ,
		_w3707_
	);
	LUT2 #(
		.INIT('h4)
	) name2527 (
		_w3706_,
		_w3707_,
		_w3708_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2528 (
		_w3678_,
		_w3679_,
		_w3706_,
		_w3707_,
		_w3709_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2529 (
		_w3688_,
		_w3689_,
		_w3691_,
		_w3692_,
		_w3710_
	);
	LUT4 #(
		.INIT('h3200)
	) name2530 (
		_w3683_,
		_w3686_,
		_w3709_,
		_w3710_,
		_w3711_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2531 (
		_w3684_,
		_w3685_,
		_w3697_,
		_w3698_,
		_w3712_
	);
	LUT2 #(
		.INIT('h2)
	) name2532 (
		\g1024_reg/NET0131 ,
		\g1964_reg/NET0131 ,
		_w3713_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2533 (
		\g1018_reg/NET0131 ,
		\g1965_reg/NET0131 ,
		\g1966_reg/NET0131 ,
		\g5657_pad ,
		_w3714_
	);
	LUT2 #(
		.INIT('h4)
	) name2534 (
		_w3713_,
		_w3714_,
		_w3715_
	);
	LUT4 #(
		.INIT('h3777)
	) name2535 (
		_w3700_,
		_w3708_,
		_w3712_,
		_w3715_,
		_w3716_
	);
	LUT4 #(
		.INIT('h0400)
	) name2536 (
		_w3678_,
		_w3679_,
		_w3684_,
		_w3685_,
		_w3717_
	);
	LUT4 #(
		.INIT('h4044)
	) name2537 (
		_w3688_,
		_w3689_,
		_w3697_,
		_w3698_,
		_w3718_
	);
	LUT4 #(
		.INIT('h0ddd)
	) name2538 (
		_w3687_,
		_w3715_,
		_w3717_,
		_w3718_,
		_w3719_
	);
	LUT4 #(
		.INIT('h1000)
	) name2539 (
		_w3705_,
		_w3711_,
		_w3716_,
		_w3719_,
		_w3720_
	);
	LUT4 #(
		.INIT('he8f8)
	) name2540 (
		_w3683_,
		_w3686_,
		_w3693_,
		_w3715_,
		_w3721_
	);
	LUT4 #(
		.INIT('h4044)
	) name2541 (
		_w3678_,
		_w3679_,
		_w3697_,
		_w3698_,
		_w3722_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2542 (
		_w3706_,
		_w3707_,
		_w3713_,
		_w3714_,
		_w3723_
	);
	LUT4 #(
		.INIT('h4044)
	) name2543 (
		_w3684_,
		_w3685_,
		_w3697_,
		_w3698_,
		_w3724_
	);
	LUT2 #(
		.INIT('h8)
	) name2544 (
		_w3723_,
		_w3724_,
		_w3725_
	);
	LUT2 #(
		.INIT('h8)
	) name2545 (
		\g1018_reg/NET0131 ,
		\g1947_reg/NET0131 ,
		_w3726_
	);
	LUT4 #(
		.INIT('h0777)
	) name2546 (
		\g1024_reg/NET0131 ,
		\g1870_reg/NET0131 ,
		\g1945_reg/NET0131 ,
		\g5657_pad ,
		_w3727_
	);
	LUT2 #(
		.INIT('h4)
	) name2547 (
		_w3726_,
		_w3727_,
		_w3728_
	);
	LUT2 #(
		.INIT('h8)
	) name2548 (
		\g185_reg/NET0131 ,
		\g1922_reg/NET0131 ,
		_w3729_
	);
	LUT3 #(
		.INIT('hb0)
	) name2549 (
		_w3726_,
		_w3727_,
		_w3729_,
		_w3730_
	);
	LUT2 #(
		.INIT('h8)
	) name2550 (
		\g1018_reg/NET0131 ,
		\g1979_reg/NET0131 ,
		_w3731_
	);
	LUT4 #(
		.INIT('h135f)
	) name2551 (
		\g1024_reg/NET0131 ,
		\g1976_reg/NET0131 ,
		\g1982_reg/NET0131 ,
		\g5657_pad ,
		_w3732_
	);
	LUT2 #(
		.INIT('h4)
	) name2552 (
		_w3731_,
		_w3732_,
		_w3733_
	);
	LUT4 #(
		.INIT('h0700)
	) name2553 (
		_w3723_,
		_w3724_,
		_w3730_,
		_w3733_,
		_w3734_
	);
	LUT3 #(
		.INIT('hb0)
	) name2554 (
		_w3721_,
		_w3722_,
		_w3734_,
		_w3735_
	);
	LUT3 #(
		.INIT('h40)
	) name2555 (
		_w3702_,
		_w3720_,
		_w3735_,
		_w3736_
	);
	LUT4 #(
		.INIT('h8000)
	) name2556 (
		_w3686_,
		_w3704_,
		_w3715_,
		_w3718_,
		_w3737_
	);
	LUT3 #(
		.INIT('h80)
	) name2557 (
		_w3696_,
		_w3703_,
		_w3715_,
		_w3738_
	);
	LUT4 #(
		.INIT('h0400)
	) name2558 (
		_w3691_,
		_w3692_,
		_w3706_,
		_w3707_,
		_w3739_
	);
	LUT4 #(
		.INIT('hf1fd)
	) name2559 (
		_w3687_,
		_w3690_,
		_w3699_,
		_w3739_,
		_w3740_
	);
	LUT3 #(
		.INIT('h10)
	) name2560 (
		_w3737_,
		_w3738_,
		_w3740_,
		_w3741_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2561 (
		_w3691_,
		_w3692_,
		_w3697_,
		_w3698_,
		_w3742_
	);
	LUT4 #(
		.INIT('h400a)
	) name2562 (
		_w3686_,
		_w3690_,
		_w3693_,
		_w3699_,
		_w3743_
	);
	LUT4 #(
		.INIT('h57df)
	) name2563 (
		_w3680_,
		_w3686_,
		_w3700_,
		_w3710_,
		_w3744_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2564 (
		_w3688_,
		_w3689_,
		_w3697_,
		_w3698_,
		_w3745_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2565 (
		_w3684_,
		_w3685_,
		_w3713_,
		_w3714_,
		_w3746_
	);
	LUT4 #(
		.INIT('hcedf)
	) name2566 (
		_w3680_,
		_w3683_,
		_w3745_,
		_w3746_,
		_w3747_
	);
	LUT4 #(
		.INIT('h7000)
	) name2567 (
		_w3709_,
		_w3743_,
		_w3744_,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h8)
	) name2568 (
		\g1949_reg/NET0131 ,
		\g5657_pad ,
		_w3749_
	);
	LUT4 #(
		.INIT('h135f)
	) name2569 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1951_reg/NET0131 ,
		\g1953_reg/NET0131 ,
		_w3750_
	);
	LUT2 #(
		.INIT('h4)
	) name2570 (
		_w3749_,
		_w3750_,
		_w3751_
	);
	LUT2 #(
		.INIT('h8)
	) name2571 (
		\g185_reg/NET0131 ,
		\g1904_reg/NET0131 ,
		_w3752_
	);
	LUT3 #(
		.INIT('hb0)
	) name2572 (
		_w3749_,
		_w3750_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h8)
	) name2573 (
		\g1024_reg/NET0131 ,
		\g1973_reg/NET0131 ,
		_w3754_
	);
	LUT4 #(
		.INIT('h135f)
	) name2574 (
		\g1018_reg/NET0131 ,
		\g1967_reg/NET0131 ,
		\g1970_reg/NET0131 ,
		\g5657_pad ,
		_w3755_
	);
	LUT2 #(
		.INIT('h4)
	) name2575 (
		_w3754_,
		_w3755_,
		_w3756_
	);
	LUT2 #(
		.INIT('h4)
	) name2576 (
		_w3753_,
		_w3756_,
		_w3757_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2577 (
		_w3730_,
		_w3733_,
		_w3753_,
		_w3756_,
		_w3758_
	);
	LUT2 #(
		.INIT('h2)
	) name2578 (
		_w3315_,
		_w3758_,
		_w3759_
	);
	LUT3 #(
		.INIT('h80)
	) name2579 (
		_w3741_,
		_w3748_,
		_w3759_,
		_w3760_
	);
	LUT3 #(
		.INIT('hba)
	) name2580 (
		_w3677_,
		_w3736_,
		_w3760_,
		_w3761_
	);
	LUT2 #(
		.INIT('h1)
	) name2581 (
		_w2865_,
		_w3315_,
		_w3762_
	);
	LUT2 #(
		.INIT('h2)
	) name2582 (
		\g5657_pad ,
		\g576_reg/NET0131 ,
		_w3763_
	);
	LUT4 #(
		.INIT('hf351)
	) name2583 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g575_reg/NET0131 ,
		\g577_reg/NET0131 ,
		_w3764_
	);
	LUT2 #(
		.INIT('h4)
	) name2584 (
		_w3763_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h2)
	) name2585 (
		\g1024_reg/NET0131 ,
		\g578_reg/NET0131 ,
		_w3766_
	);
	LUT4 #(
		.INIT('hf351)
	) name2586 (
		\g1018_reg/NET0131 ,
		\g5657_pad ,
		\g579_reg/NET0131 ,
		\g580_reg/NET0131 ,
		_w3767_
	);
	LUT2 #(
		.INIT('h4)
	) name2587 (
		_w3766_,
		_w3767_,
		_w3768_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2588 (
		_w3763_,
		_w3764_,
		_w3766_,
		_w3767_,
		_w3769_
	);
	LUT2 #(
		.INIT('h8)
	) name2589 (
		\g1018_reg/NET0131 ,
		\g366_reg/NET0131 ,
		_w3770_
	);
	LUT4 #(
		.INIT('h135f)
	) name2590 (
		\g1024_reg/NET0131 ,
		\g364_reg/NET0131 ,
		\g368_reg/NET0131 ,
		\g5657_pad ,
		_w3771_
	);
	LUT2 #(
		.INIT('h4)
	) name2591 (
		_w3770_,
		_w3771_,
		_w3772_
	);
	LUT2 #(
		.INIT('h8)
	) name2592 (
		\g1018_reg/NET0131 ,
		\g351_reg/NET0131 ,
		_w3773_
	);
	LUT4 #(
		.INIT('h135f)
	) name2593 (
		\g1024_reg/NET0131 ,
		\g349_reg/NET0131 ,
		\g353_reg/NET0131 ,
		\g5657_pad ,
		_w3774_
	);
	LUT2 #(
		.INIT('h4)
	) name2594 (
		_w3773_,
		_w3774_,
		_w3775_
	);
	LUT4 #(
		.INIT('h0400)
	) name2595 (
		_w3770_,
		_w3771_,
		_w3773_,
		_w3774_,
		_w3776_
	);
	LUT2 #(
		.INIT('h2)
	) name2596 (
		\g1024_reg/NET0131 ,
		\g581_reg/NET0131 ,
		_w3777_
	);
	LUT4 #(
		.INIT('hf351)
	) name2597 (
		\g1018_reg/NET0131 ,
		\g5657_pad ,
		\g582_reg/NET0131 ,
		\g583_reg/NET0131 ,
		_w3778_
	);
	LUT2 #(
		.INIT('h4)
	) name2598 (
		_w3777_,
		_w3778_,
		_w3779_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2599 (
		_w3763_,
		_w3764_,
		_w3777_,
		_w3778_,
		_w3780_
	);
	LUT4 #(
		.INIT('h4044)
	) name2600 (
		_w3770_,
		_w3771_,
		_w3773_,
		_w3774_,
		_w3781_
	);
	LUT4 #(
		.INIT('h737f)
	) name2601 (
		_w3769_,
		_w3772_,
		_w3775_,
		_w3780_,
		_w3782_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2602 (
		_w3770_,
		_w3771_,
		_w3773_,
		_w3774_,
		_w3783_
	);
	LUT2 #(
		.INIT('h8)
	) name2603 (
		\g1018_reg/NET0131 ,
		\g381_reg/NET0131 ,
		_w3784_
	);
	LUT4 #(
		.INIT('h135f)
	) name2604 (
		\g1024_reg/NET0131 ,
		\g379_reg/NET0131 ,
		\g383_reg/NET0131 ,
		\g5657_pad ,
		_w3785_
	);
	LUT2 #(
		.INIT('h4)
	) name2605 (
		_w3784_,
		_w3785_,
		_w3786_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2606 (
		_w3766_,
		_w3767_,
		_w3784_,
		_w3785_,
		_w3787_
	);
	LUT2 #(
		.INIT('h2)
	) name2607 (
		\g5657_pad ,
		\g585_reg/NET0131 ,
		_w3788_
	);
	LUT4 #(
		.INIT('hf351)
	) name2608 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g584_reg/NET0131 ,
		\g586_reg/NET0131 ,
		_w3789_
	);
	LUT2 #(
		.INIT('h4)
	) name2609 (
		_w3788_,
		_w3789_,
		_w3790_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2610 (
		_w3773_,
		_w3774_,
		_w3788_,
		_w3789_,
		_w3791_
	);
	LUT2 #(
		.INIT('h8)
	) name2611 (
		\g1018_reg/NET0131 ,
		\g396_reg/NET0131 ,
		_w3792_
	);
	LUT4 #(
		.INIT('h0777)
	) name2612 (
		\g1024_reg/NET0131 ,
		\g324_reg/NET0131 ,
		\g394_reg/NET0131 ,
		\g5657_pad ,
		_w3793_
	);
	LUT2 #(
		.INIT('h4)
	) name2613 (
		_w3792_,
		_w3793_,
		_w3794_
	);
	LUT4 #(
		.INIT('h0400)
	) name2614 (
		_w3763_,
		_w3764_,
		_w3792_,
		_w3793_,
		_w3795_
	);
	LUT4 #(
		.INIT('h0777)
	) name2615 (
		_w3783_,
		_w3787_,
		_w3791_,
		_w3795_,
		_w3796_
	);
	LUT4 #(
		.INIT('h4044)
	) name2616 (
		_w3770_,
		_w3771_,
		_w3784_,
		_w3785_,
		_w3797_
	);
	LUT4 #(
		.INIT('h5100)
	) name2617 (
		_w3765_,
		_w3779_,
		_w3791_,
		_w3797_,
		_w3798_
	);
	LUT4 #(
		.INIT('h0400)
	) name2618 (
		_w3763_,
		_w3764_,
		_w3766_,
		_w3767_,
		_w3799_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2619 (
		_w3770_,
		_w3771_,
		_w3773_,
		_w3774_,
		_w3800_
	);
	LUT3 #(
		.INIT('h40)
	) name2620 (
		_w3786_,
		_w3799_,
		_w3800_,
		_w3801_
	);
	LUT4 #(
		.INIT('h0008)
	) name2621 (
		_w3782_,
		_w3796_,
		_w3798_,
		_w3801_,
		_w3802_
	);
	LUT4 #(
		.INIT('h4044)
	) name2622 (
		_w3763_,
		_w3764_,
		_w3777_,
		_w3778_,
		_w3803_
	);
	LUT4 #(
		.INIT('hf200)
	) name2623 (
		_w3783_,
		_w3786_,
		_w3794_,
		_w3803_,
		_w3804_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2624 (
		_w3766_,
		_w3767_,
		_w3777_,
		_w3778_,
		_w3805_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2625 (
		_w3773_,
		_w3774_,
		_w3784_,
		_w3785_,
		_w3806_
	);
	LUT4 #(
		.INIT('hf020)
	) name2626 (
		_w3783_,
		_w3794_,
		_w3805_,
		_w3806_,
		_w3807_
	);
	LUT2 #(
		.INIT('h1)
	) name2627 (
		_w3804_,
		_w3807_,
		_w3808_
	);
	LUT2 #(
		.INIT('h8)
	) name2628 (
		\g1018_reg/NET0131 ,
		\g567_reg/NET0131 ,
		_w3809_
	);
	LUT4 #(
		.INIT('h0777)
	) name2629 (
		\g1024_reg/NET0131 ,
		\g489_reg/NET0131 ,
		\g5657_pad ,
		\g565_reg/NET0131 ,
		_w3810_
	);
	LUT2 #(
		.INIT('h4)
	) name2630 (
		_w3809_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h8)
	) name2631 (
		\g185_reg/NET0131 ,
		\g542_reg/NET0131 ,
		_w3812_
	);
	LUT3 #(
		.INIT('hb0)
	) name2632 (
		_w3809_,
		_w3810_,
		_w3812_,
		_w3813_
	);
	LUT2 #(
		.INIT('h8)
	) name2633 (
		\g1024_reg/NET0131 ,
		\g602_reg/NET0131 ,
		_w3814_
	);
	LUT4 #(
		.INIT('h153f)
	) name2634 (
		\g1018_reg/NET0131 ,
		\g5657_pad ,
		\g596_reg/NET0131 ,
		\g599_reg/NET0131 ,
		_w3815_
	);
	LUT2 #(
		.INIT('h4)
	) name2635 (
		_w3814_,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h4)
	) name2636 (
		_w3813_,
		_w3816_,
		_w3817_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2637 (
		_w3770_,
		_w3771_,
		_w3784_,
		_w3785_,
		_w3818_
	);
	LUT4 #(
		.INIT('h0400)
	) name2638 (
		_w3766_,
		_w3767_,
		_w3777_,
		_w3778_,
		_w3819_
	);
	LUT3 #(
		.INIT('h80)
	) name2639 (
		_w3775_,
		_w3818_,
		_w3819_,
		_w3820_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2640 (
		_w3763_,
		_w3764_,
		_w3792_,
		_w3793_,
		_w3821_
	);
	LUT4 #(
		.INIT('h4044)
	) name2641 (
		_w3773_,
		_w3774_,
		_w3788_,
		_w3789_,
		_w3822_
	);
	LUT3 #(
		.INIT('he0)
	) name2642 (
		_w3786_,
		_w3821_,
		_w3822_,
		_w3823_
	);
	LUT3 #(
		.INIT('h02)
	) name2643 (
		_w3817_,
		_w3820_,
		_w3823_,
		_w3824_
	);
	LUT3 #(
		.INIT('h80)
	) name2644 (
		_w3802_,
		_w3808_,
		_w3824_,
		_w3825_
	);
	LUT4 #(
		.INIT('h4044)
	) name2645 (
		_w3763_,
		_w3764_,
		_w3766_,
		_w3767_,
		_w3826_
	);
	LUT4 #(
		.INIT('h135f)
	) name2646 (
		_w3781_,
		_w3797_,
		_w3803_,
		_w3826_,
		_w3827_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2647 (
		_w3784_,
		_w3785_,
		_w3788_,
		_w3789_,
		_w3828_
	);
	LUT3 #(
		.INIT('h80)
	) name2648 (
		_w3769_,
		_w3800_,
		_w3828_,
		_w3829_
	);
	LUT3 #(
		.INIT('h20)
	) name2649 (
		_w3780_,
		_w3794_,
		_w3800_,
		_w3830_
	);
	LUT3 #(
		.INIT('h80)
	) name2650 (
		_w3790_,
		_w3799_,
		_w3806_,
		_w3831_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2651 (
		_w3763_,
		_w3764_,
		_w3773_,
		_w3774_,
		_w3832_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2652 (
		_w3784_,
		_w3785_,
		_w3788_,
		_w3789_,
		_w3833_
	);
	LUT4 #(
		.INIT('h153f)
	) name2653 (
		_w3783_,
		_w3787_,
		_w3832_,
		_w3833_,
		_w3834_
	);
	LUT4 #(
		.INIT('h0100)
	) name2654 (
		_w3829_,
		_w3830_,
		_w3831_,
		_w3834_,
		_w3835_
	);
	LUT3 #(
		.INIT('h20)
	) name2655 (
		_w3783_,
		_w3794_,
		_w3799_,
		_w3836_
	);
	LUT4 #(
		.INIT('h8bcf)
	) name2656 (
		_w3765_,
		_w3768_,
		_w3776_,
		_w3794_,
		_w3837_
	);
	LUT3 #(
		.INIT('h8a)
	) name2657 (
		_w3779_,
		_w3836_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h8)
	) name2658 (
		\g5657_pad ,
		\g569_reg/NET0131 ,
		_w3839_
	);
	LUT4 #(
		.INIT('h135f)
	) name2659 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g571_reg/NET0131 ,
		\g573_reg/NET0131 ,
		_w3840_
	);
	LUT2 #(
		.INIT('h4)
	) name2660 (
		_w3839_,
		_w3840_,
		_w3841_
	);
	LUT2 #(
		.INIT('h8)
	) name2661 (
		\g185_reg/NET0131 ,
		\g524_reg/NET0131 ,
		_w3842_
	);
	LUT3 #(
		.INIT('hb0)
	) name2662 (
		_w3839_,
		_w3840_,
		_w3842_,
		_w3843_
	);
	LUT2 #(
		.INIT('h8)
	) name2663 (
		\g1018_reg/NET0131 ,
		\g590_reg/NET0131 ,
		_w3844_
	);
	LUT4 #(
		.INIT('h153f)
	) name2664 (
		\g1024_reg/NET0131 ,
		\g5657_pad ,
		\g587_reg/NET0131 ,
		\g593_reg/NET0131 ,
		_w3845_
	);
	LUT2 #(
		.INIT('h4)
	) name2665 (
		_w3844_,
		_w3845_,
		_w3846_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		_w3843_,
		_w3846_,
		_w3847_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2667 (
		_w3813_,
		_w3816_,
		_w3843_,
		_w3846_,
		_w3848_
	);
	LUT2 #(
		.INIT('h2)
	) name2668 (
		_w3315_,
		_w3848_,
		_w3849_
	);
	LUT4 #(
		.INIT('h0800)
	) name2669 (
		_w3827_,
		_w3835_,
		_w3838_,
		_w3849_,
		_w3850_
	);
	LUT3 #(
		.INIT('hba)
	) name2670 (
		_w3762_,
		_w3825_,
		_w3850_,
		_w3851_
	);
	LUT2 #(
		.INIT('h2)
	) name2671 (
		_w2208_,
		_w3315_,
		_w3852_
	);
	LUT4 #(
		.INIT('h004f)
	) name2672 (
		_w3282_,
		_w3307_,
		_w3315_,
		_w3852_,
		_w3853_
	);
	LUT4 #(
		.INIT('h5303)
	) name2673 (
		\g1092_reg/NET0131 ,
		\g298_reg/NET0131 ,
		\g299_reg/NET0131 ,
		\g305_reg/NET0131 ,
		_w3854_
	);
	LUT2 #(
		.INIT('h1)
	) name2674 (
		_w1574_,
		_w3315_,
		_w3855_
	);
	LUT4 #(
		.INIT('h1000)
	) name2675 (
		_w3737_,
		_w3738_,
		_w3740_,
		_w3757_,
		_w3856_
	);
	LUT3 #(
		.INIT('h4c)
	) name2676 (
		_w3748_,
		_w3759_,
		_w3856_,
		_w3857_
	);
	LUT3 #(
		.INIT('h0b)
	) name2677 (
		_w3721_,
		_w3722_,
		_w3725_,
		_w3858_
	);
	LUT3 #(
		.INIT('h40)
	) name2678 (
		_w3702_,
		_w3720_,
		_w3858_,
		_w3859_
	);
	LUT3 #(
		.INIT('hea)
	) name2679 (
		_w3855_,
		_w3857_,
		_w3859_,
		_w3860_
	);
	LUT2 #(
		.INIT('h1)
	) name2680 (
		_w2212_,
		_w3315_,
		_w3861_
	);
	LUT3 #(
		.INIT('h01)
	) name2681 (
		_w3292_,
		_w3294_,
		_w3296_,
		_w3862_
	);
	LUT4 #(
		.INIT('h0700)
	) name2682 (
		_w3275_,
		_w3284_,
		_w3301_,
		_w3304_,
		_w3863_
	);
	LUT3 #(
		.INIT('he0)
	) name2683 (
		_w3228_,
		_w3283_,
		_w3863_,
		_w3864_
	);
	LUT3 #(
		.INIT('h80)
	) name2684 (
		_w3291_,
		_w3862_,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h4)
	) name2685 (
		_w3305_,
		_w3315_,
		_w3866_
	);
	LUT4 #(
		.INIT('h0800)
	) name2686 (
		_w3245_,
		_w3259_,
		_w3281_,
		_w3866_,
		_w3867_
	);
	LUT3 #(
		.INIT('hba)
	) name2687 (
		_w3861_,
		_w3865_,
		_w3867_,
		_w3868_
	);
	LUT2 #(
		.INIT('h1)
	) name2688 (
		_w2861_,
		_w3315_,
		_w3869_
	);
	LUT4 #(
		.INIT('h7500)
	) name2689 (
		_w3779_,
		_w3836_,
		_w3837_,
		_w3847_,
		_w3870_
	);
	LUT3 #(
		.INIT('h80)
	) name2690 (
		_w3827_,
		_w3835_,
		_w3870_,
		_w3871_
	);
	LUT4 #(
		.INIT('h0002)
	) name2691 (
		_w3315_,
		_w3820_,
		_w3823_,
		_w3848_,
		_w3872_
	);
	LUT3 #(
		.INIT('h80)
	) name2692 (
		_w3802_,
		_w3808_,
		_w3872_,
		_w3873_
	);
	LUT3 #(
		.INIT('hba)
	) name2693 (
		_w3869_,
		_w3871_,
		_w3873_,
		_w3874_
	);
	LUT2 #(
		.INIT('h8)
	) name2694 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w3875_
	);
	LUT3 #(
		.INIT('h8c)
	) name2695 (
		_w1700_,
		_w1736_,
		_w2291_,
		_w3876_
	);
	LUT4 #(
		.INIT('h0080)
	) name2696 (
		_w1771_,
		_w1780_,
		_w1797_,
		_w3452_,
		_w3877_
	);
	LUT3 #(
		.INIT('h02)
	) name2697 (
		_w3875_,
		_w3876_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h8)
	) name2698 (
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w3879_
	);
	LUT3 #(
		.INIT('h10)
	) name2699 (
		_w3876_,
		_w3877_,
		_w3879_,
		_w3880_
	);
	LUT2 #(
		.INIT('h8)
	) name2700 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w3881_
	);
	LUT3 #(
		.INIT('h10)
	) name2701 (
		_w3876_,
		_w3877_,
		_w3881_,
		_w3882_
	);
	LUT4 #(
		.INIT('h0080)
	) name2702 (
		_w1287_,
		_w1299_,
		_w1308_,
		_w3459_,
		_w3883_
	);
	LUT4 #(
		.INIT('h7500)
	) name2703 (
		_w1313_,
		_w1364_,
		_w2474_,
		_w3875_,
		_w3884_
	);
	LUT2 #(
		.INIT('h4)
	) name2704 (
		_w3883_,
		_w3884_,
		_w3885_
	);
	LUT4 #(
		.INIT('h7500)
	) name2705 (
		_w1313_,
		_w1364_,
		_w2474_,
		_w3879_,
		_w3886_
	);
	LUT2 #(
		.INIT('h4)
	) name2706 (
		_w3883_,
		_w3886_,
		_w3887_
	);
	LUT4 #(
		.INIT('h7500)
	) name2707 (
		_w1313_,
		_w1364_,
		_w2474_,
		_w3881_,
		_w3888_
	);
	LUT2 #(
		.INIT('h4)
	) name2708 (
		_w3883_,
		_w3888_,
		_w3889_
	);
	LUT2 #(
		.INIT('h4)
	) name2709 (
		_w1859_,
		_w2337_,
		_w3890_
	);
	LUT4 #(
		.INIT('h80c0)
	) name2710 (
		_w1859_,
		_w1926_,
		_w1938_,
		_w2337_,
		_w3891_
	);
	LUT4 #(
		.INIT('h7300)
	) name2711 (
		_w1859_,
		_w1890_,
		_w2337_,
		_w3875_,
		_w3892_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2712 (
		_w1982_,
		_w1983_,
		_w3891_,
		_w3892_,
		_w3893_
	);
	LUT4 #(
		.INIT('h7300)
	) name2713 (
		_w1859_,
		_w1890_,
		_w2337_,
		_w3879_,
		_w3894_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2714 (
		_w1982_,
		_w1983_,
		_w3891_,
		_w3894_,
		_w3895_
	);
	LUT4 #(
		.INIT('h7300)
	) name2715 (
		_w1859_,
		_w1890_,
		_w2337_,
		_w3881_,
		_w3896_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2716 (
		_w1982_,
		_w1983_,
		_w3891_,
		_w3896_,
		_w3897_
	);
	LUT4 #(
		.INIT('h2022)
	) name2717 (
		_w2094_,
		_w2103_,
		_w2121_,
		_w2435_,
		_w3898_
	);
	LUT4 #(
		.INIT('h7500)
	) name2718 (
		_w2009_,
		_w2121_,
		_w2435_,
		_w3875_,
		_w3899_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2719 (
		_w2115_,
		_w2116_,
		_w3898_,
		_w3899_,
		_w3900_
	);
	LUT4 #(
		.INIT('h7500)
	) name2720 (
		_w2009_,
		_w2121_,
		_w2435_,
		_w3879_,
		_w3901_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2721 (
		_w2115_,
		_w2116_,
		_w3898_,
		_w3901_,
		_w3902_
	);
	LUT4 #(
		.INIT('h7500)
	) name2722 (
		_w2009_,
		_w2121_,
		_w2435_,
		_w3881_,
		_w3903_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2723 (
		_w2115_,
		_w2116_,
		_w3898_,
		_w3903_,
		_w3904_
	);
	LUT3 #(
		.INIT('h23)
	) name2724 (
		\g1018_reg/NET0131 ,
		\g1192_reg/NET0131 ,
		\g16355_pad ,
		_w3905_
	);
	LUT3 #(
		.INIT('ha2)
	) name2725 (
		\g1018_reg/NET0131 ,
		\g506_reg/NET0131 ,
		\g507_reg/NET0131 ,
		_w3906_
	);
	LUT3 #(
		.INIT('h51)
	) name2726 (
		_w2951_,
		_w3905_,
		_w3906_,
		_w3907_
	);
	LUT3 #(
		.INIT('h08)
	) name2727 (
		\g1024_reg/NET0131 ,
		\g1326_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w3908_
	);
	LUT4 #(
		.INIT('h8000)
	) name2728 (
		\g1319_reg/NET0131 ,
		\g1332_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		\g1346_reg/NET0131 ,
		_w3909_
	);
	LUT2 #(
		.INIT('h8)
	) name2729 (
		_w3908_,
		_w3909_,
		_w3910_
	);
	LUT3 #(
		.INIT('h80)
	) name2730 (
		\g1352_reg/NET0131 ,
		\g1358_reg/NET0131 ,
		\g1365_reg/NET0131 ,
		_w3911_
	);
	LUT2 #(
		.INIT('h8)
	) name2731 (
		\g1372_reg/NET0131 ,
		\g1378_reg/NET0131 ,
		_w3912_
	);
	LUT4 #(
		.INIT('h8000)
	) name2732 (
		_w3908_,
		_w3909_,
		_w3911_,
		_w3912_,
		_w3913_
	);
	LUT2 #(
		.INIT('h8)
	) name2733 (
		\g1018_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		_w3914_
	);
	LUT3 #(
		.INIT('h70)
	) name2734 (
		\g1018_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		\g1378_reg/NET0131 ,
		_w3915_
	);
	LUT3 #(
		.INIT('h70)
	) name2735 (
		\g1018_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		\g1372_reg/NET0131 ,
		_w3916_
	);
	LUT4 #(
		.INIT('h8000)
	) name2736 (
		_w3908_,
		_w3909_,
		_w3911_,
		_w3916_,
		_w3917_
	);
	LUT3 #(
		.INIT('h54)
	) name2737 (
		_w3913_,
		_w3915_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h8)
	) name2738 (
		\g1092_reg/NET0131 ,
		\g1098_reg/NET0131 ,
		_w3919_
	);
	LUT4 #(
		.INIT('h135f)
	) name2739 (
		\g1088_reg/NET0131 ,
		\g1095_reg/NET0131 ,
		\g1101_reg/NET0131 ,
		\g7961_pad ,
		_w3920_
	);
	LUT2 #(
		.INIT('h2)
	) name2740 (
		\g1088_reg/NET0131 ,
		\g1113_reg/NET0131 ,
		_w3921_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2741 (
		\g1092_reg/NET0131 ,
		\g1114_reg/NET0131 ,
		\g1115_reg/NET0131 ,
		\g7961_pad ,
		_w3922_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2742 (
		_w3919_,
		_w3920_,
		_w3921_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h8)
	) name2743 (
		\g1092_reg/NET0131 ,
		\g1107_reg/NET0131 ,
		_w3924_
	);
	LUT4 #(
		.INIT('h135f)
	) name2744 (
		\g1088_reg/NET0131 ,
		\g1104_reg/NET0131 ,
		\g1110_reg/NET0131 ,
		\g7961_pad ,
		_w3925_
	);
	LUT2 #(
		.INIT('h4)
	) name2745 (
		_w3924_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('hb)
	) name2746 (
		_w3924_,
		_w3925_,
		_w3927_
	);
	LUT3 #(
		.INIT('h07)
	) name2747 (
		\g1563_reg/NET0131 ,
		_w3923_,
		_w3926_,
		_w3928_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2748 (
		_w1874_,
		_w1875_,
		_w1898_,
		_w1899_,
		_w3929_
	);
	LUT4 #(
		.INIT('h8000)
	) name2749 (
		\g793_reg/NET0131 ,
		\g797_reg/NET0131 ,
		\g805_reg/NET0131 ,
		\g809_reg/NET0131 ,
		_w3930_
	);
	LUT4 #(
		.INIT('h8000)
	) name2750 (
		\g785_reg/NET0131 ,
		\g789_reg/NET0131 ,
		\g801_reg/NET0131 ,
		\g813_reg/NET0131 ,
		_w3931_
	);
	LUT2 #(
		.INIT('h8)
	) name2751 (
		_w3930_,
		_w3931_,
		_w3932_
	);
	LUT2 #(
		.INIT('h7)
	) name2752 (
		_w3930_,
		_w3931_,
		_w3933_
	);
	LUT3 #(
		.INIT('h80)
	) name2753 (
		\g1563_reg/NET0131 ,
		_w3930_,
		_w3931_,
		_w3934_
	);
	LUT4 #(
		.INIT('he000)
	) name2754 (
		_w1890_,
		_w3923_,
		_w3929_,
		_w3934_,
		_w3935_
	);
	LUT2 #(
		.INIT('he)
	) name2755 (
		_w3928_,
		_w3935_,
		_w3936_
	);
	LUT2 #(
		.INIT('h8)
	) name2756 (
		\g1092_reg/NET0131 ,
		\g411_reg/NET0131 ,
		_w3937_
	);
	LUT4 #(
		.INIT('h135f)
	) name2757 (
		\g1088_reg/NET0131 ,
		\g408_reg/NET0131 ,
		\g414_reg/NET0131 ,
		\g7961_pad ,
		_w3938_
	);
	LUT2 #(
		.INIT('h2)
	) name2758 (
		\g1088_reg/NET0131 ,
		\g426_reg/NET0131 ,
		_w3939_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2759 (
		\g1092_reg/NET0131 ,
		\g427_reg/NET0131 ,
		\g428_reg/NET0131 ,
		\g7961_pad ,
		_w3940_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2760 (
		_w3937_,
		_w3938_,
		_w3939_,
		_w3940_,
		_w3941_
	);
	LUT2 #(
		.INIT('h8)
	) name2761 (
		\g1092_reg/NET0131 ,
		\g420_reg/NET0131 ,
		_w3942_
	);
	LUT4 #(
		.INIT('h135f)
	) name2762 (
		\g1088_reg/NET0131 ,
		\g417_reg/NET0131 ,
		\g423_reg/NET0131 ,
		\g7961_pad ,
		_w3943_
	);
	LUT2 #(
		.INIT('h4)
	) name2763 (
		_w3942_,
		_w3943_,
		_w3944_
	);
	LUT2 #(
		.INIT('hb)
	) name2764 (
		_w3942_,
		_w3943_,
		_w3945_
	);
	LUT3 #(
		.INIT('h07)
	) name2765 (
		\g1563_reg/NET0131 ,
		_w3941_,
		_w3944_,
		_w3946_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2766 (
		_w1728_,
		_w1729_,
		_w1738_,
		_w1739_,
		_w3947_
	);
	LUT4 #(
		.INIT('h8000)
	) name2767 (
		\g109_reg/NET0131 ,
		\g117_reg/NET0131 ,
		\g121_reg/NET0131 ,
		\g97_reg/NET0131 ,
		_w3948_
	);
	LUT4 #(
		.INIT('h8000)
	) name2768 (
		\g101_reg/NET0131 ,
		\g105_reg/NET0131 ,
		\g113_reg/NET0131 ,
		\g125_reg/NET0131 ,
		_w3949_
	);
	LUT2 #(
		.INIT('h8)
	) name2769 (
		_w3948_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h7)
	) name2770 (
		_w3948_,
		_w3949_,
		_w3951_
	);
	LUT3 #(
		.INIT('h80)
	) name2771 (
		\g1563_reg/NET0131 ,
		_w3948_,
		_w3949_,
		_w3952_
	);
	LUT4 #(
		.INIT('he000)
	) name2772 (
		_w1736_,
		_w3941_,
		_w3947_,
		_w3952_,
		_w3953_
	);
	LUT2 #(
		.INIT('he)
	) name2773 (
		_w3946_,
		_w3953_,
		_w3954_
	);
	LUT2 #(
		.INIT('h8)
	) name2774 (
		\g1092_reg/NET0131 ,
		\g2486_reg/NET0131 ,
		_w3955_
	);
	LUT4 #(
		.INIT('h135f)
	) name2775 (
		\g1088_reg/NET0131 ,
		\g2483_reg/NET0131 ,
		\g2489_reg/NET0131 ,
		\g7961_pad ,
		_w3956_
	);
	LUT2 #(
		.INIT('h2)
	) name2776 (
		\g1088_reg/NET0131 ,
		\g2501_reg/NET0131 ,
		_w3957_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2777 (
		\g1092_reg/NET0131 ,
		\g2502_reg/NET0131 ,
		\g2503_reg/NET0131 ,
		\g7961_pad ,
		_w3958_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2778 (
		_w3955_,
		_w3956_,
		_w3957_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h8)
	) name2779 (
		\g1092_reg/NET0131 ,
		\g2495_reg/NET0131 ,
		_w3960_
	);
	LUT4 #(
		.INIT('h135f)
	) name2780 (
		\g1088_reg/NET0131 ,
		\g2492_reg/NET0131 ,
		\g2498_reg/NET0131 ,
		\g7961_pad ,
		_w3961_
	);
	LUT2 #(
		.INIT('h4)
	) name2781 (
		_w3960_,
		_w3961_,
		_w3962_
	);
	LUT2 #(
		.INIT('hb)
	) name2782 (
		_w3960_,
		_w3961_,
		_w3963_
	);
	LUT3 #(
		.INIT('h07)
	) name2783 (
		\g1563_reg/NET0131 ,
		_w3959_,
		_w3962_,
		_w3964_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2784 (
		_w1267_,
		_w1268_,
		_w1292_,
		_w1293_,
		_w3965_
	);
	LUT4 #(
		.INIT('h8000)
	) name2785 (
		\g2175_reg/NET0131 ,
		\g2180_reg/NET0131 ,
		\g2190_reg/NET0131 ,
		\g2195_reg/NET0131 ,
		_w3966_
	);
	LUT4 #(
		.INIT('h8000)
	) name2786 (
		\g2165_reg/NET0131 ,
		\g2170_reg/NET0131 ,
		\g2185_reg/NET0131 ,
		\g2200_reg/NET0131 ,
		_w3967_
	);
	LUT2 #(
		.INIT('h8)
	) name2787 (
		_w3966_,
		_w3967_,
		_w3968_
	);
	LUT3 #(
		.INIT('h80)
	) name2788 (
		\g1563_reg/NET0131 ,
		_w3966_,
		_w3967_,
		_w3969_
	);
	LUT4 #(
		.INIT('he000)
	) name2789 (
		_w1313_,
		_w3959_,
		_w3965_,
		_w3969_,
		_w3970_
	);
	LUT2 #(
		.INIT('he)
	) name2790 (
		_w3964_,
		_w3970_,
		_w3971_
	);
	LUT2 #(
		.INIT('h2)
	) name2791 (
		\g1088_reg/NET0131 ,
		\g1807_reg/NET0131 ,
		_w3972_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name2792 (
		\g1092_reg/NET0131 ,
		\g1808_reg/NET0131 ,
		\g1809_reg/NET0131 ,
		\g7961_pad ,
		_w3973_
	);
	LUT2 #(
		.INIT('h8)
	) name2793 (
		\g1092_reg/NET0131 ,
		\g1792_reg/NET0131 ,
		_w3974_
	);
	LUT4 #(
		.INIT('h135f)
	) name2794 (
		\g1088_reg/NET0131 ,
		\g1789_reg/NET0131 ,
		\g1795_reg/NET0131 ,
		\g7961_pad ,
		_w3975_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2795 (
		_w3972_,
		_w3973_,
		_w3974_,
		_w3975_,
		_w3976_
	);
	LUT2 #(
		.INIT('h8)
	) name2796 (
		\g1092_reg/NET0131 ,
		\g1801_reg/NET0131 ,
		_w3977_
	);
	LUT4 #(
		.INIT('h135f)
	) name2797 (
		\g1088_reg/NET0131 ,
		\g1798_reg/NET0131 ,
		\g1804_reg/NET0131 ,
		\g7961_pad ,
		_w3978_
	);
	LUT2 #(
		.INIT('h4)
	) name2798 (
		_w3977_,
		_w3978_,
		_w3979_
	);
	LUT2 #(
		.INIT('hb)
	) name2799 (
		_w3977_,
		_w3978_,
		_w3980_
	);
	LUT3 #(
		.INIT('h07)
	) name2800 (
		\g1563_reg/NET0131 ,
		_w3976_,
		_w3979_,
		_w3981_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2801 (
		_w2011_,
		_w2012_,
		_w2068_,
		_w2069_,
		_w3982_
	);
	LUT4 #(
		.INIT('h8000)
	) name2802 (
		\g1481_reg/NET0131 ,
		\g1486_reg/NET0131 ,
		\g1496_reg/NET0131 ,
		\g1501_reg/NET0131 ,
		_w3983_
	);
	LUT4 #(
		.INIT('h8000)
	) name2803 (
		\g1471_reg/NET0131 ,
		\g1476_reg/NET0131 ,
		\g1491_reg/NET0131 ,
		\g1506_reg/NET0131 ,
		_w3984_
	);
	LUT2 #(
		.INIT('h8)
	) name2804 (
		_w3983_,
		_w3984_,
		_w3985_
	);
	LUT2 #(
		.INIT('h7)
	) name2805 (
		_w3983_,
		_w3984_,
		_w3986_
	);
	LUT3 #(
		.INIT('h80)
	) name2806 (
		\g1563_reg/NET0131 ,
		_w3983_,
		_w3984_,
		_w3987_
	);
	LUT4 #(
		.INIT('he000)
	) name2807 (
		_w2009_,
		_w3976_,
		_w3982_,
		_w3987_,
		_w3988_
	);
	LUT2 #(
		.INIT('he)
	) name2808 (
		_w3981_,
		_w3988_,
		_w3989_
	);
	LUT4 #(
		.INIT('h2000)
	) name2809 (
		_w1897_,
		_w1903_,
		_w1910_,
		_w1916_,
		_w3990_
	);
	LUT4 #(
		.INIT('h7fff)
	) name2810 (
		_w1873_,
		_w1887_,
		_w1893_,
		_w3990_,
		_w3991_
	);
	LUT2 #(
		.INIT('h7)
	) name2811 (
		_w1828_,
		_w3454_,
		_w3992_
	);
	LUT4 #(
		.INIT('h8000)
	) name2812 (
		_w1348_,
		_w1351_,
		_w1355_,
		_w1373_,
		_w3993_
	);
	LUT3 #(
		.INIT('h7f)
	) name2813 (
		_w1326_,
		_w1337_,
		_w3993_,
		_w3994_
	);
	LUT4 #(
		.INIT('h0200)
	) name2814 (
		_w2067_,
		_w2073_,
		_w2076_,
		_w2139_,
		_w3995_
	);
	LUT3 #(
		.INIT('h7f)
	) name2815 (
		_w2054_,
		_w2064_,
		_w3995_,
		_w3996_
	);
	LUT3 #(
		.INIT('h45)
	) name2816 (
		\g1563_reg/NET0131 ,
		_w3919_,
		_w3920_,
		_w3997_
	);
	LUT4 #(
		.INIT('h0d00)
	) name2817 (
		_w1852_,
		_w1853_,
		_w3924_,
		_w3925_,
		_w3998_
	);
	LUT3 #(
		.INIT('h08)
	) name2818 (
		_w3929_,
		_w3932_,
		_w3998_,
		_w3999_
	);
	LUT3 #(
		.INIT('h8a)
	) name2819 (
		\g1563_reg/NET0131 ,
		_w3924_,
		_w3925_,
		_w4000_
	);
	LUT3 #(
		.INIT('h07)
	) name2820 (
		_w3929_,
		_w3934_,
		_w4000_,
		_w4001_
	);
	LUT4 #(
		.INIT('hcccd)
	) name2821 (
		_w3923_,
		_w3997_,
		_w3999_,
		_w4001_,
		_w4002_
	);
	LUT3 #(
		.INIT('h45)
	) name2822 (
		\g1563_reg/NET0131 ,
		_w3937_,
		_w3938_,
		_w4003_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2823 (
		_w1734_,
		_w1735_,
		_w3942_,
		_w3943_,
		_w4004_
	);
	LUT3 #(
		.INIT('h08)
	) name2824 (
		_w3947_,
		_w3950_,
		_w4004_,
		_w4005_
	);
	LUT3 #(
		.INIT('h8a)
	) name2825 (
		\g1563_reg/NET0131 ,
		_w3942_,
		_w3943_,
		_w4006_
	);
	LUT3 #(
		.INIT('h07)
	) name2826 (
		_w3947_,
		_w3952_,
		_w4006_,
		_w4007_
	);
	LUT4 #(
		.INIT('hcccd)
	) name2827 (
		_w3941_,
		_w4003_,
		_w4005_,
		_w4007_,
		_w4008_
	);
	LUT3 #(
		.INIT('h45)
	) name2828 (
		\g1563_reg/NET0131 ,
		_w3955_,
		_w3956_,
		_w4009_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2829 (
		_w1311_,
		_w1312_,
		_w3960_,
		_w3961_,
		_w4010_
	);
	LUT3 #(
		.INIT('h08)
	) name2830 (
		_w3965_,
		_w3968_,
		_w4010_,
		_w4011_
	);
	LUT3 #(
		.INIT('h8a)
	) name2831 (
		\g1563_reg/NET0131 ,
		_w3960_,
		_w3961_,
		_w4012_
	);
	LUT3 #(
		.INIT('h07)
	) name2832 (
		_w3965_,
		_w3969_,
		_w4012_,
		_w4013_
	);
	LUT4 #(
		.INIT('hcccd)
	) name2833 (
		_w3959_,
		_w4009_,
		_w4011_,
		_w4013_,
		_w4014_
	);
	LUT3 #(
		.INIT('h45)
	) name2834 (
		\g1563_reg/NET0131 ,
		_w3974_,
		_w3975_,
		_w4015_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2835 (
		_w2007_,
		_w2008_,
		_w3977_,
		_w3978_,
		_w4016_
	);
	LUT3 #(
		.INIT('h08)
	) name2836 (
		_w3982_,
		_w3985_,
		_w4016_,
		_w4017_
	);
	LUT3 #(
		.INIT('h8a)
	) name2837 (
		\g1563_reg/NET0131 ,
		_w3977_,
		_w3978_,
		_w4018_
	);
	LUT3 #(
		.INIT('h07)
	) name2838 (
		_w3982_,
		_w3987_,
		_w4018_,
		_w4019_
	);
	LUT4 #(
		.INIT('hcccd)
	) name2839 (
		_w3976_,
		_w4015_,
		_w4017_,
		_w4019_,
		_w4020_
	);
	LUT3 #(
		.INIT('h45)
	) name2840 (
		_w3315_,
		_w3753_,
		_w3756_,
		_w4021_
	);
	LUT3 #(
		.INIT('h45)
	) name2841 (
		_w3315_,
		_w3730_,
		_w3733_,
		_w4022_
	);
	LUT3 #(
		.INIT('h45)
	) name2842 (
		_w3315_,
		_w3843_,
		_w3846_,
		_w4023_
	);
	LUT3 #(
		.INIT('h45)
	) name2843 (
		_w3315_,
		_w3813_,
		_w3816_,
		_w4024_
	);
	LUT3 #(
		.INIT('h0b)
	) name2844 (
		_w3301_,
		_w3304_,
		_w3315_,
		_w4025_
	);
	LUT3 #(
		.INIT('h0b)
	) name2845 (
		_w3264_,
		_w3267_,
		_w3315_,
		_w4026_
	);
	LUT3 #(
		.INIT('h45)
	) name2846 (
		_w3315_,
		_w3397_,
		_w3400_,
		_w4027_
	);
	LUT3 #(
		.INIT('h45)
	) name2847 (
		_w3315_,
		_w3376_,
		_w3379_,
		_w4028_
	);
	LUT4 #(
		.INIT('h7f00)
	) name2848 (
		_w3908_,
		_w3909_,
		_w3911_,
		_w3916_,
		_w4029_
	);
	LUT3 #(
		.INIT('h07)
	) name2849 (
		\g1018_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		\g1372_reg/NET0131 ,
		_w4030_
	);
	LUT4 #(
		.INIT('h8000)
	) name2850 (
		_w3908_,
		_w3909_,
		_w3911_,
		_w4030_,
		_w4031_
	);
	LUT2 #(
		.INIT('he)
	) name2851 (
		_w4029_,
		_w4031_,
		_w4032_
	);
	LUT3 #(
		.INIT('h73)
	) name2852 (
		_w1391_,
		_w1396_,
		_w1398_,
		_w4033_
	);
	LUT2 #(
		.INIT('h2)
	) name2853 (
		\g1088_reg/NET0131 ,
		_w3923_,
		_w4034_
	);
	LUT3 #(
		.INIT('h10)
	) name2854 (
		_w3999_,
		_w4001_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h2)
	) name2855 (
		\g7961_pad ,
		_w3923_,
		_w4036_
	);
	LUT3 #(
		.INIT('h10)
	) name2856 (
		_w3999_,
		_w4001_,
		_w4036_,
		_w4037_
	);
	LUT2 #(
		.INIT('h2)
	) name2857 (
		\g1092_reg/NET0131 ,
		_w3923_,
		_w4038_
	);
	LUT3 #(
		.INIT('h10)
	) name2858 (
		_w3999_,
		_w4001_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h2)
	) name2859 (
		\g1088_reg/NET0131 ,
		_w3941_,
		_w4040_
	);
	LUT3 #(
		.INIT('h10)
	) name2860 (
		_w4005_,
		_w4007_,
		_w4040_,
		_w4041_
	);
	LUT2 #(
		.INIT('h2)
	) name2861 (
		\g7961_pad ,
		_w3941_,
		_w4042_
	);
	LUT3 #(
		.INIT('h10)
	) name2862 (
		_w4005_,
		_w4007_,
		_w4042_,
		_w4043_
	);
	LUT2 #(
		.INIT('h2)
	) name2863 (
		\g1092_reg/NET0131 ,
		_w3941_,
		_w4044_
	);
	LUT3 #(
		.INIT('h10)
	) name2864 (
		_w4005_,
		_w4007_,
		_w4044_,
		_w4045_
	);
	LUT2 #(
		.INIT('h2)
	) name2865 (
		\g1088_reg/NET0131 ,
		_w3959_,
		_w4046_
	);
	LUT3 #(
		.INIT('h10)
	) name2866 (
		_w4011_,
		_w4013_,
		_w4046_,
		_w4047_
	);
	LUT2 #(
		.INIT('h2)
	) name2867 (
		\g7961_pad ,
		_w3959_,
		_w4048_
	);
	LUT3 #(
		.INIT('h10)
	) name2868 (
		_w4011_,
		_w4013_,
		_w4048_,
		_w4049_
	);
	LUT2 #(
		.INIT('h2)
	) name2869 (
		\g1092_reg/NET0131 ,
		_w3959_,
		_w4050_
	);
	LUT3 #(
		.INIT('h10)
	) name2870 (
		_w4011_,
		_w4013_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h2)
	) name2871 (
		\g1088_reg/NET0131 ,
		_w3976_,
		_w4052_
	);
	LUT3 #(
		.INIT('h10)
	) name2872 (
		_w4017_,
		_w4019_,
		_w4052_,
		_w4053_
	);
	LUT2 #(
		.INIT('h2)
	) name2873 (
		\g7961_pad ,
		_w3976_,
		_w4054_
	);
	LUT3 #(
		.INIT('h10)
	) name2874 (
		_w4017_,
		_w4019_,
		_w4054_,
		_w4055_
	);
	LUT2 #(
		.INIT('h2)
	) name2875 (
		\g1092_reg/NET0131 ,
		_w3976_,
		_w4056_
	);
	LUT3 #(
		.INIT('h10)
	) name2876 (
		_w4017_,
		_w4019_,
		_w4056_,
		_w4057_
	);
	LUT3 #(
		.INIT('h2a)
	) name2877 (
		\g1426_reg/NET0131 ,
		\g267_reg/NET0131 ,
		\g7961_pad ,
		_w4058_
	);
	LUT2 #(
		.INIT('h8)
	) name2878 (
		_w1756_,
		_w4058_,
		_w4059_
	);
	LUT3 #(
		.INIT('h51)
	) name2879 (
		\g1457_reg/NET0131 ,
		_w1789_,
		_w1790_,
		_w4060_
	);
	LUT3 #(
		.INIT('h2a)
	) name2880 (
		\g1457_reg/NET0131 ,
		\g195_reg/NET0131 ,
		\g7961_pad ,
		_w4061_
	);
	LUT3 #(
		.INIT('h4c)
	) name2881 (
		\g1088_reg/NET0131 ,
		\g1448_reg/NET0131 ,
		\g210_reg/NET0131 ,
		_w4062_
	);
	LUT4 #(
		.INIT('h135f)
	) name2882 (
		_w1789_,
		_w1794_,
		_w4061_,
		_w4062_,
		_w4063_
	);
	LUT3 #(
		.INIT('h10)
	) name2883 (
		_w4059_,
		_w4060_,
		_w4063_,
		_w4064_
	);
	LUT3 #(
		.INIT('h2a)
	) name2884 (
		\g1435_reg/NET0131 ,
		\g258_reg/NET0131 ,
		\g7961_pad ,
		_w4065_
	);
	LUT3 #(
		.INIT('h4c)
	) name2885 (
		\g1088_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		\g192_reg/NET0131 ,
		_w4066_
	);
	LUT4 #(
		.INIT('h135f)
	) name2886 (
		_w1759_,
		_w1781_,
		_w4065_,
		_w4066_,
		_w4067_
	);
	LUT3 #(
		.INIT('h51)
	) name2887 (
		\g1435_reg/NET0131 ,
		_w1759_,
		_w1760_,
		_w4068_
	);
	LUT3 #(
		.INIT('h45)
	) name2888 (
		\g1426_reg/NET0131 ,
		_w1755_,
		_w1756_,
		_w4069_
	);
	LUT3 #(
		.INIT('h02)
	) name2889 (
		_w4067_,
		_w4068_,
		_w4069_,
		_w4070_
	);
	LUT2 #(
		.INIT('h1)
	) name2890 (
		\g2896_reg/NET0131 ,
		\g2900_reg/NET0131 ,
		_w4071_
	);
	LUT3 #(
		.INIT('h01)
	) name2891 (
		\g2892_reg/NET0131 ,
		\g2903_reg/NET0131 ,
		\g2908_reg/NET0131 ,
		_w4072_
	);
	LUT2 #(
		.INIT('h8)
	) name2892 (
		_w4071_,
		_w4072_,
		_w4073_
	);
	LUT4 #(
		.INIT('h0b00)
	) name2893 (
		_w1695_,
		_w1696_,
		_w1698_,
		_w1699_,
		_w4074_
	);
	LUT2 #(
		.INIT('h4)
	) name2894 (
		_w1747_,
		_w4074_,
		_w4075_
	);
	LUT3 #(
		.INIT('h23)
	) name2895 (
		_w1747_,
		_w4073_,
		_w4074_,
		_w4076_
	);
	LUT3 #(
		.INIT('h2a)
	) name2896 (
		\g1453_reg/NET0131 ,
		\g240_reg/NET0131 ,
		\g7961_pad ,
		_w4077_
	);
	LUT3 #(
		.INIT('h2a)
	) name2897 (
		\g1439_reg/NET0131 ,
		\g213_reg/NET0131 ,
		\g7961_pad ,
		_w4078_
	);
	LUT4 #(
		.INIT('h135f)
	) name2898 (
		_w1776_,
		_w1786_,
		_w4077_,
		_w4078_,
		_w4079_
	);
	LUT3 #(
		.INIT('h45)
	) name2899 (
		\g1439_reg/NET0131 ,
		_w1785_,
		_w1786_,
		_w4080_
	);
	LUT3 #(
		.INIT('h51)
	) name2900 (
		\g1453_reg/NET0131 ,
		_w1776_,
		_w1777_,
		_w4081_
	);
	LUT3 #(
		.INIT('h02)
	) name2901 (
		_w4079_,
		_w4080_,
		_w4081_,
		_w4082_
	);
	LUT4 #(
		.INIT('h8000)
	) name2902 (
		_w4064_,
		_w4070_,
		_w4076_,
		_w4082_,
		_w4083_
	);
	LUT3 #(
		.INIT('h59)
	) name2903 (
		\g1462_reg/NET0131 ,
		_w1767_,
		_w1768_,
		_w4084_
	);
	LUT3 #(
		.INIT('h65)
	) name2904 (
		\g1430_reg/NET0131 ,
		_w1763_,
		_w1764_,
		_w4085_
	);
	LUT2 #(
		.INIT('h1)
	) name2905 (
		_w4084_,
		_w4085_,
		_w4086_
	);
	LUT3 #(
		.INIT('h45)
	) name2906 (
		\g1448_reg/NET0131 ,
		_w1793_,
		_w1794_,
		_w4087_
	);
	LUT3 #(
		.INIT('h51)
	) name2907 (
		\g1466_reg/NET0131 ,
		_w1781_,
		_w1782_,
		_w4088_
	);
	LUT3 #(
		.INIT('h59)
	) name2908 (
		\g1444_reg/NET0131 ,
		_w1772_,
		_w1773_,
		_w4089_
	);
	LUT3 #(
		.INIT('h01)
	) name2909 (
		_w4087_,
		_w4088_,
		_w4089_,
		_w4090_
	);
	LUT2 #(
		.INIT('h8)
	) name2910 (
		_w4086_,
		_w4090_,
		_w4091_
	);
	LUT4 #(
		.INIT('h8000)
	) name2911 (
		_w1795_,
		_w1821_,
		_w2300_,
		_w2301_,
		_w4092_
	);
	LUT2 #(
		.INIT('h8)
	) name2912 (
		_w2319_,
		_w4092_,
		_w4093_
	);
	LUT3 #(
		.INIT('h07)
	) name2913 (
		_w4083_,
		_w4091_,
		_w4093_,
		_w4094_
	);
	LUT3 #(
		.INIT('h2a)
	) name2914 (
		\g1426_reg/NET0131 ,
		\g7961_pad ,
		\g954_reg/NET0131 ,
		_w4095_
	);
	LUT3 #(
		.INIT('h2a)
	) name2915 (
		\g1453_reg/NET0131 ,
		\g7961_pad ,
		\g927_reg/NET0131 ,
		_w4096_
	);
	LUT4 #(
		.INIT('h153f)
	) name2916 (
		_w1954_,
		_w1958_,
		_w4095_,
		_w4096_,
		_w4097_
	);
	LUT3 #(
		.INIT('h45)
	) name2917 (
		\g1439_reg/NET0131 ,
		_w1935_,
		_w1936_,
		_w4098_
	);
	LUT3 #(
		.INIT('h45)
	) name2918 (
		\g1448_reg/NET0131 ,
		_w1923_,
		_w1924_,
		_w4099_
	);
	LUT3 #(
		.INIT('h02)
	) name2919 (
		_w4097_,
		_w4098_,
		_w4099_,
		_w4100_
	);
	LUT3 #(
		.INIT('h2a)
	) name2920 (
		\g1439_reg/NET0131 ,
		\g7961_pad ,
		\g900_reg/NET0131 ,
		_w4101_
	);
	LUT3 #(
		.INIT('h2a)
	) name2921 (
		\g1457_reg/NET0131 ,
		\g7961_pad ,
		\g882_reg/NET0131 ,
		_w4102_
	);
	LUT4 #(
		.INIT('h153f)
	) name2922 (
		_w1932_,
		_w1936_,
		_w4101_,
		_w4102_,
		_w4103_
	);
	LUT3 #(
		.INIT('h2a)
	) name2923 (
		\g1462_reg/NET0131 ,
		\g7961_pad ,
		\g918_reg/NET0131 ,
		_w4104_
	);
	LUT2 #(
		.INIT('h8)
	) name2924 (
		_w1962_,
		_w4104_,
		_w4105_
	);
	LUT2 #(
		.INIT('h2)
	) name2925 (
		_w4103_,
		_w4105_,
		_w4106_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2926 (
		_w1846_,
		_w1847_,
		_w1849_,
		_w1850_,
		_w4107_
	);
	LUT2 #(
		.INIT('h8)
	) name2927 (
		_w1859_,
		_w4107_,
		_w4108_
	);
	LUT3 #(
		.INIT('h4c)
	) name2928 (
		\g1088_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		\g879_reg/NET0131 ,
		_w4109_
	);
	LUT4 #(
		.INIT('h153f)
	) name2929 (
		_w1940_,
		_w4071_,
		_w4072_,
		_w4109_,
		_w4110_
	);
	LUT3 #(
		.INIT('h70)
	) name2930 (
		_w1859_,
		_w4107_,
		_w4110_,
		_w4111_
	);
	LUT3 #(
		.INIT('h80)
	) name2931 (
		_w4100_,
		_w4106_,
		_w4111_,
		_w4112_
	);
	LUT3 #(
		.INIT('h4c)
	) name2932 (
		\g1088_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		\g942_reg/NET0131 ,
		_w4113_
	);
	LUT2 #(
		.INIT('h8)
	) name2933 (
		_w1971_,
		_w4113_,
		_w4114_
	);
	LUT3 #(
		.INIT('h45)
	) name2934 (
		\g1426_reg/NET0131 ,
		_w1957_,
		_w1958_,
		_w4115_
	);
	LUT3 #(
		.INIT('h45)
	) name2935 (
		\g1430_reg/NET0131 ,
		_w1927_,
		_w1928_,
		_w4116_
	);
	LUT3 #(
		.INIT('h45)
	) name2936 (
		\g1457_reg/NET0131 ,
		_w1931_,
		_w1932_,
		_w4117_
	);
	LUT4 #(
		.INIT('h0001)
	) name2937 (
		_w4114_,
		_w4115_,
		_w4116_,
		_w4117_,
		_w4118_
	);
	LUT3 #(
		.INIT('h4c)
	) name2938 (
		\g1088_reg/NET0131 ,
		\g1448_reg/NET0131 ,
		\g897_reg/NET0131 ,
		_w4119_
	);
	LUT2 #(
		.INIT('h8)
	) name2939 (
		_w1924_,
		_w4119_,
		_w4120_
	);
	LUT3 #(
		.INIT('h45)
	) name2940 (
		\g1435_reg/NET0131 ,
		_w1965_,
		_w1966_,
		_w4121_
	);
	LUT3 #(
		.INIT('h4c)
	) name2941 (
		\g1092_reg/NET0131 ,
		\g1435_reg/NET0131 ,
		\g948_reg/NET0131 ,
		_w4122_
	);
	LUT3 #(
		.INIT('h2a)
	) name2942 (
		\g1430_reg/NET0131 ,
		\g7961_pad ,
		\g909_reg/NET0131 ,
		_w4123_
	);
	LUT4 #(
		.INIT('h153f)
	) name2943 (
		_w1928_,
		_w1966_,
		_w4122_,
		_w4123_,
		_w4124_
	);
	LUT3 #(
		.INIT('h10)
	) name2944 (
		_w4120_,
		_w4121_,
		_w4124_,
		_w4125_
	);
	LUT3 #(
		.INIT('h45)
	) name2945 (
		\g1453_reg/NET0131 ,
		_w1953_,
		_w1954_,
		_w4126_
	);
	LUT3 #(
		.INIT('h45)
	) name2946 (
		\g1444_reg/NET0131 ,
		_w1970_,
		_w1971_,
		_w4127_
	);
	LUT3 #(
		.INIT('h45)
	) name2947 (
		\g1462_reg/NET0131 ,
		_w1961_,
		_w1962_,
		_w4128_
	);
	LUT3 #(
		.INIT('h51)
	) name2948 (
		\g1466_reg/NET0131 ,
		_w1940_,
		_w1941_,
		_w4129_
	);
	LUT4 #(
		.INIT('h0001)
	) name2949 (
		_w4126_,
		_w4127_,
		_w4128_,
		_w4129_,
		_w4130_
	);
	LUT3 #(
		.INIT('h80)
	) name2950 (
		_w4118_,
		_w4125_,
		_w4130_,
		_w4131_
	);
	LUT4 #(
		.INIT('h8000)
	) name2951 (
		_w1919_,
		_w1942_,
		_w2352_,
		_w2353_,
		_w4132_
	);
	LUT2 #(
		.INIT('h8)
	) name2952 (
		_w2358_,
		_w4132_,
		_w4133_
	);
	LUT3 #(
		.INIT('h07)
	) name2953 (
		_w4112_,
		_w4131_,
		_w4133_,
		_w4134_
	);
	LUT3 #(
		.INIT('h4c)
	) name2954 (
		\g1092_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		\g2291_reg/NET0131 ,
		_w4135_
	);
	LUT2 #(
		.INIT('h8)
	) name2955 (
		_w1289_,
		_w4135_,
		_w4136_
	);
	LUT3 #(
		.INIT('h45)
	) name2956 (
		\g1426_reg/NET0131 ,
		_w1270_,
		_w1271_,
		_w4137_
	);
	LUT3 #(
		.INIT('h45)
	) name2957 (
		\g1439_reg/NET0131 ,
		_w1288_,
		_w1289_,
		_w4138_
	);
	LUT3 #(
		.INIT('h2a)
	) name2958 (
		\g1430_reg/NET0131 ,
		\g2297_reg/NET0131 ,
		\g7961_pad ,
		_w4139_
	);
	LUT2 #(
		.INIT('h8)
	) name2959 (
		_w1296_,
		_w4139_,
		_w4140_
	);
	LUT4 #(
		.INIT('h0001)
	) name2960 (
		_w4136_,
		_w4137_,
		_w4138_,
		_w4140_,
		_w4141_
	);
	LUT3 #(
		.INIT('h2a)
	) name2961 (
		\g1457_reg/NET0131 ,
		\g2270_reg/NET0131 ,
		\g7961_pad ,
		_w4142_
	);
	LUT3 #(
		.INIT('h2a)
	) name2962 (
		\g1426_reg/NET0131 ,
		\g2342_reg/NET0131 ,
		\g7961_pad ,
		_w4143_
	);
	LUT4 #(
		.INIT('h153f)
	) name2963 (
		_w1271_,
		_w1305_,
		_w4142_,
		_w4143_,
		_w4144_
	);
	LUT3 #(
		.INIT('h45)
	) name2964 (
		\g1457_reg/NET0131 ,
		_w1304_,
		_w1305_,
		_w4145_
	);
	LUT3 #(
		.INIT('h51)
	) name2965 (
		\g1444_reg/NET0131 ,
		_w1263_,
		_w1264_,
		_w4146_
	);
	LUT3 #(
		.INIT('h02)
	) name2966 (
		_w4144_,
		_w4145_,
		_w4146_,
		_w4147_
	);
	LUT2 #(
		.INIT('h8)
	) name2967 (
		_w4141_,
		_w4147_,
		_w4148_
	);
	LUT3 #(
		.INIT('h4c)
	) name2968 (
		\g1092_reg/NET0131 ,
		\g1435_reg/NET0131 ,
		\g2336_reg/NET0131 ,
		_w4149_
	);
	LUT3 #(
		.INIT('h2a)
	) name2969 (
		\g1453_reg/NET0131 ,
		\g2315_reg/NET0131 ,
		\g7961_pad ,
		_w4150_
	);
	LUT4 #(
		.INIT('h135f)
	) name2970 (
		_w1255_,
		_w1274_,
		_w4149_,
		_w4150_,
		_w4151_
	);
	LUT3 #(
		.INIT('h51)
	) name2971 (
		\g1466_reg/NET0131 ,
		_w1300_,
		_w1301_,
		_w4152_
	);
	LUT3 #(
		.INIT('h45)
	) name2972 (
		\g1430_reg/NET0131 ,
		_w1295_,
		_w1296_,
		_w4153_
	);
	LUT3 #(
		.INIT('h02)
	) name2973 (
		_w4151_,
		_w4152_,
		_w4153_,
		_w4154_
	);
	LUT3 #(
		.INIT('h45)
	) name2974 (
		\g1462_reg/NET0131 ,
		_w1258_,
		_w1259_,
		_w4155_
	);
	LUT3 #(
		.INIT('h45)
	) name2975 (
		\g1435_reg/NET0131 ,
		_w1254_,
		_w1255_,
		_w4156_
	);
	LUT3 #(
		.INIT('h4c)
	) name2976 (
		\g1092_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		\g2327_reg/NET0131 ,
		_w4157_
	);
	LUT2 #(
		.INIT('h8)
	) name2977 (
		_w1263_,
		_w4157_,
		_w4158_
	);
	LUT3 #(
		.INIT('h51)
	) name2978 (
		\g1453_reg/NET0131 ,
		_w1274_,
		_w1275_,
		_w4159_
	);
	LUT4 #(
		.INIT('h0001)
	) name2979 (
		_w4155_,
		_w4156_,
		_w4158_,
		_w4159_,
		_w4160_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name2980 (
		_w1251_,
		_w1252_,
		_w1366_,
		_w1367_,
		_w4161_
	);
	LUT2 #(
		.INIT('h8)
	) name2981 (
		_w1364_,
		_w4161_,
		_w4162_
	);
	LUT3 #(
		.INIT('h13)
	) name2982 (
		_w1364_,
		_w4073_,
		_w4161_,
		_w4163_
	);
	LUT3 #(
		.INIT('h2a)
	) name2983 (
		\g1462_reg/NET0131 ,
		\g2306_reg/NET0131 ,
		\g7961_pad ,
		_w4164_
	);
	LUT3 #(
		.INIT('h4c)
	) name2984 (
		\g1092_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		\g2264_reg/NET0131 ,
		_w4165_
	);
	LUT4 #(
		.INIT('h135f)
	) name2985 (
		_w1259_,
		_w1300_,
		_w4164_,
		_w4165_,
		_w4166_
	);
	LUT3 #(
		.INIT('h9a)
	) name2986 (
		\g1448_reg/NET0131 ,
		_w1283_,
		_w1284_,
		_w4167_
	);
	LUT2 #(
		.INIT('h8)
	) name2987 (
		_w4166_,
		_w4167_,
		_w4168_
	);
	LUT4 #(
		.INIT('h8000)
	) name2988 (
		_w4154_,
		_w4160_,
		_w4163_,
		_w4168_,
		_w4169_
	);
	LUT4 #(
		.INIT('h8000)
	) name2989 (
		_w1302_,
		_w1369_,
		_w2482_,
		_w2483_,
		_w4170_
	);
	LUT2 #(
		.INIT('h8)
	) name2990 (
		_w2487_,
		_w4170_,
		_w4171_
	);
	LUT3 #(
		.INIT('h07)
	) name2991 (
		_w4148_,
		_w4169_,
		_w4171_,
		_w4172_
	);
	LUT3 #(
		.INIT('h4c)
	) name2992 (
		\g1092_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		\g1570_reg/NET0131 ,
		_w4173_
	);
	LUT2 #(
		.INIT('h8)
	) name2993 (
		_w2026_,
		_w4173_,
		_w4174_
	);
	LUT3 #(
		.INIT('h45)
	) name2994 (
		\g1448_reg/NET0131 ,
		_w2022_,
		_w2023_,
		_w4175_
	);
	LUT3 #(
		.INIT('h51)
	) name2995 (
		\g1453_reg/NET0131 ,
		_w2095_,
		_w2096_,
		_w4176_
	);
	LUT3 #(
		.INIT('h45)
	) name2996 (
		\g1462_reg/NET0131 ,
		_w2087_,
		_w2088_,
		_w4177_
	);
	LUT4 #(
		.INIT('h0001)
	) name2997 (
		_w4174_,
		_w4175_,
		_w4176_,
		_w4177_,
		_w4178_
	);
	LUT3 #(
		.INIT('h4c)
	) name2998 (
		\g1088_reg/NET0131 ,
		\g1448_reg/NET0131 ,
		\g1591_reg/NET0131 ,
		_w4179_
	);
	LUT3 #(
		.INIT('h2a)
	) name2999 (
		\g1430_reg/NET0131 ,
		\g1603_reg/NET0131 ,
		\g7961_pad ,
		_w4180_
	);
	LUT4 #(
		.INIT('h153f)
	) name3000 (
		_w2015_,
		_w2023_,
		_w4179_,
		_w4180_,
		_w4181_
	);
	LUT3 #(
		.INIT('h45)
	) name3001 (
		\g1439_reg/NET0131 ,
		_w2018_,
		_w2019_,
		_w4182_
	);
	LUT3 #(
		.INIT('h45)
	) name3002 (
		\g1426_reg/NET0131 ,
		_w2100_,
		_w2101_,
		_w4183_
	);
	LUT3 #(
		.INIT('h02)
	) name3003 (
		_w4181_,
		_w4182_,
		_w4183_,
		_w4184_
	);
	LUT2 #(
		.INIT('h8)
	) name3004 (
		_w4178_,
		_w4184_,
		_w4185_
	);
	LUT3 #(
		.INIT('h2a)
	) name3005 (
		\g1426_reg/NET0131 ,
		\g1648_reg/NET0131 ,
		\g7961_pad ,
		_w4186_
	);
	LUT2 #(
		.INIT('h8)
	) name3006 (
		_w2101_,
		_w4186_,
		_w4187_
	);
	LUT3 #(
		.INIT('h45)
	) name3007 (
		\g1435_reg/NET0131 ,
		_w2091_,
		_w2092_,
		_w4188_
	);
	LUT3 #(
		.INIT('h2a)
	) name3008 (
		\g1435_reg/NET0131 ,
		\g1639_reg/NET0131 ,
		\g7961_pad ,
		_w4189_
	);
	LUT3 #(
		.INIT('h2a)
	) name3009 (
		\g1453_reg/NET0131 ,
		\g1621_reg/NET0131 ,
		\g7961_pad ,
		_w4190_
	);
	LUT4 #(
		.INIT('h135f)
	) name3010 (
		_w2092_,
		_w2095_,
		_w4189_,
		_w4190_,
		_w4191_
	);
	LUT3 #(
		.INIT('h10)
	) name3011 (
		_w4187_,
		_w4188_,
		_w4191_,
		_w4192_
	);
	LUT3 #(
		.INIT('h45)
	) name3012 (
		\g1430_reg/NET0131 ,
		_w2014_,
		_w2015_,
		_w4193_
	);
	LUT3 #(
		.INIT('h51)
	) name3013 (
		\g1466_reg/NET0131 ,
		_w2026_,
		_w2027_,
		_w4194_
	);
	LUT3 #(
		.INIT('h45)
	) name3014 (
		\g1457_reg/NET0131 ,
		_w2030_,
		_w2031_,
		_w4195_
	);
	LUT3 #(
		.INIT('h51)
	) name3015 (
		\g1444_reg/NET0131 ,
		_w2083_,
		_w2084_,
		_w4196_
	);
	LUT4 #(
		.INIT('h0001)
	) name3016 (
		_w4193_,
		_w4194_,
		_w4195_,
		_w4196_,
		_w4197_
	);
	LUT4 #(
		.INIT('hb0bb)
	) name3017 (
		_w2111_,
		_w2112_,
		_w2127_,
		_w2128_,
		_w4198_
	);
	LUT2 #(
		.INIT('h8)
	) name3018 (
		_w2121_,
		_w4198_,
		_w4199_
	);
	LUT3 #(
		.INIT('h13)
	) name3019 (
		_w2121_,
		_w4073_,
		_w4198_,
		_w4200_
	);
	LUT3 #(
		.INIT('h2a)
	) name3020 (
		\g1439_reg/NET0131 ,
		\g1594_reg/NET0131 ,
		\g7961_pad ,
		_w4201_
	);
	LUT3 #(
		.INIT('h2a)
	) name3021 (
		\g1462_reg/NET0131 ,
		\g1612_reg/NET0131 ,
		\g7961_pad ,
		_w4202_
	);
	LUT4 #(
		.INIT('h135f)
	) name3022 (
		_w2019_,
		_w2088_,
		_w4201_,
		_w4202_,
		_w4203_
	);
	LUT3 #(
		.INIT('h2a)
	) name3023 (
		\g1457_reg/NET0131 ,
		\g1576_reg/NET0131 ,
		\g7961_pad ,
		_w4204_
	);
	LUT3 #(
		.INIT('h4c)
	) name3024 (
		\g1092_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		\g1633_reg/NET0131 ,
		_w4205_
	);
	LUT4 #(
		.INIT('h135f)
	) name3025 (
		_w2031_,
		_w2083_,
		_w4204_,
		_w4205_,
		_w4206_
	);
	LUT2 #(
		.INIT('h8)
	) name3026 (
		_w4203_,
		_w4206_,
		_w4207_
	);
	LUT4 #(
		.INIT('h8000)
	) name3027 (
		_w4192_,
		_w4197_,
		_w4200_,
		_w4207_,
		_w4208_
	);
	LUT4 #(
		.INIT('h8000)
	) name3028 (
		_w2093_,
		_w2143_,
		_w2441_,
		_w2442_,
		_w4209_
	);
	LUT2 #(
		.INIT('h8)
	) name3029 (
		_w2447_,
		_w4209_,
		_w4210_
	);
	LUT3 #(
		.INIT('h07)
	) name3030 (
		_w4185_,
		_w4208_,
		_w4210_,
		_w4211_
	);
	LUT2 #(
		.INIT('h2)
	) name3031 (
		\g1092_reg/NET0131 ,
		\g1561_reg/NET0131 ,
		_w4212_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3032 (
		\g1088_reg/NET0131 ,
		\g1559_reg/NET0131 ,
		\g1560_reg/NET0131 ,
		\g7961_pad ,
		_w4213_
	);
	LUT4 #(
		.INIT('h8088)
	) name3033 (
		_w3983_,
		_w3984_,
		_w4212_,
		_w4213_,
		_w4214_
	);
	LUT2 #(
		.INIT('h8)
	) name3034 (
		\g1810_reg/NET0131 ,
		\g7961_pad ,
		_w4215_
	);
	LUT3 #(
		.INIT('h15)
	) name3035 (
		\g1563_reg/NET0131 ,
		\g1810_reg/NET0131 ,
		\g7961_pad ,
		_w4216_
	);
	LUT4 #(
		.INIT('h040c)
	) name3036 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1813_reg/NET0131 ,
		\g1816_reg/NET0131 ,
		_w4217_
	);
	LUT2 #(
		.INIT('h1)
	) name3037 (
		\g1092_reg/NET0131 ,
		\g1813_reg/NET0131 ,
		_w4218_
	);
	LUT3 #(
		.INIT('h07)
	) name3038 (
		_w4216_,
		_w4217_,
		_w4218_,
		_w4219_
	);
	LUT3 #(
		.INIT('hd0)
	) name3039 (
		_w3881_,
		_w4214_,
		_w4219_,
		_w4220_
	);
	LUT2 #(
		.INIT('h2)
	) name3040 (
		\g1092_reg/NET0131 ,
		\g867_reg/NET0131 ,
		_w4221_
	);
	LUT4 #(
		.INIT('hf531)
	) name3041 (
		\g1088_reg/NET0131 ,
		\g7961_pad ,
		\g865_reg/NET0131 ,
		\g866_reg/NET0131 ,
		_w4222_
	);
	LUT4 #(
		.INIT('h8088)
	) name3042 (
		_w3930_,
		_w3931_,
		_w4221_,
		_w4222_,
		_w4223_
	);
	LUT4 #(
		.INIT('h153f)
	) name3043 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1119_reg/NET0131 ,
		\g1122_reg/NET0131 ,
		_w4224_
	);
	LUT3 #(
		.INIT('h10)
	) name3044 (
		\g1116_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w4225_
	);
	LUT2 #(
		.INIT('h1)
	) name3045 (
		\g1116_reg/NET0131 ,
		\g7961_pad ,
		_w4226_
	);
	LUT3 #(
		.INIT('h07)
	) name3046 (
		_w4224_,
		_w4225_,
		_w4226_,
		_w4227_
	);
	LUT3 #(
		.INIT('hd0)
	) name3047 (
		_w3879_,
		_w4223_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h8)
	) name3048 (
		\g1116_reg/NET0131 ,
		\g7961_pad ,
		_w4229_
	);
	LUT3 #(
		.INIT('h13)
	) name3049 (
		\g1116_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w4230_
	);
	LUT4 #(
		.INIT('h040c)
	) name3050 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1119_reg/NET0131 ,
		\g1122_reg/NET0131 ,
		_w4231_
	);
	LUT2 #(
		.INIT('h1)
	) name3051 (
		\g1092_reg/NET0131 ,
		\g1119_reg/NET0131 ,
		_w4232_
	);
	LUT3 #(
		.INIT('h07)
	) name3052 (
		_w4230_,
		_w4231_,
		_w4232_,
		_w4233_
	);
	LUT3 #(
		.INIT('hd0)
	) name3053 (
		_w3881_,
		_w4223_,
		_w4233_,
		_w4234_
	);
	LUT4 #(
		.INIT('h002a)
	) name3054 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1119_reg/NET0131 ,
		\g1122_reg/NET0131 ,
		_w4235_
	);
	LUT2 #(
		.INIT('h1)
	) name3055 (
		\g1088_reg/NET0131 ,
		\g1122_reg/NET0131 ,
		_w4236_
	);
	LUT3 #(
		.INIT('h07)
	) name3056 (
		_w4230_,
		_w4235_,
		_w4236_,
		_w4237_
	);
	LUT3 #(
		.INIT('hd0)
	) name3057 (
		_w3875_,
		_w4223_,
		_w4237_,
		_w4238_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		\g1088_reg/NET0131 ,
		\g1828_reg/NET0131 ,
		_w4239_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3059 (
		\g1092_reg/NET0131 ,
		\g1829_reg/NET0131 ,
		\g1830_reg/NET0131 ,
		\g7961_pad ,
		_w4240_
	);
	LUT2 #(
		.INIT('h4)
	) name3060 (
		_w4239_,
		_w4240_,
		_w4241_
	);
	LUT2 #(
		.INIT('h8)
	) name3061 (
		\g1092_reg/NET0131 ,
		\g1822_reg/NET0131 ,
		_w4242_
	);
	LUT4 #(
		.INIT('h135f)
	) name3062 (
		\g1088_reg/NET0131 ,
		\g1819_reg/NET0131 ,
		\g1825_reg/NET0131 ,
		\g7961_pad ,
		_w4243_
	);
	LUT2 #(
		.INIT('h4)
	) name3063 (
		_w4242_,
		_w4243_,
		_w4244_
	);
	LUT2 #(
		.INIT('hb)
	) name3064 (
		_w4242_,
		_w4243_,
		_w4245_
	);
	LUT4 #(
		.INIT('h153f)
	) name3065 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1813_reg/NET0131 ,
		\g1816_reg/NET0131 ,
		_w4246_
	);
	LUT2 #(
		.INIT('h4)
	) name3066 (
		_w4215_,
		_w4246_,
		_w4247_
	);
	LUT4 #(
		.INIT('h1000)
	) name3067 (
		_w4215_,
		_w4242_,
		_w4243_,
		_w4246_,
		_w4248_
	);
	LUT2 #(
		.INIT('h2)
	) name3068 (
		_w4241_,
		_w4248_,
		_w4249_
	);
	LUT3 #(
		.INIT('h20)
	) name3069 (
		\g1563_reg/NET0131 ,
		_w4215_,
		_w4246_,
		_w4250_
	);
	LUT3 #(
		.INIT('h20)
	) name3070 (
		\g1563_reg/NET0131 ,
		_w4242_,
		_w4243_,
		_w4251_
	);
	LUT3 #(
		.INIT('h1b)
	) name3071 (
		_w4214_,
		_w4250_,
		_w4251_,
		_w4252_
	);
	LUT2 #(
		.INIT('hd)
	) name3072 (
		_w4249_,
		_w4252_,
		_w4253_
	);
	LUT4 #(
		.INIT('h8002)
	) name3073 (
		\g1563_reg/NET0131 ,
		_w4214_,
		_w4244_,
		_w4247_,
		_w4254_
	);
	LUT4 #(
		.INIT('haa08)
	) name3074 (
		\g1088_reg/NET0131 ,
		_w4249_,
		_w4252_,
		_w4254_,
		_w4255_
	);
	LUT4 #(
		.INIT('haa08)
	) name3075 (
		\g7961_pad ,
		_w4249_,
		_w4252_,
		_w4254_,
		_w4256_
	);
	LUT4 #(
		.INIT('haa08)
	) name3076 (
		\g1092_reg/NET0131 ,
		_w4249_,
		_w4252_,
		_w4254_,
		_w4257_
	);
	LUT2 #(
		.INIT('h8)
	) name3077 (
		\g1092_reg/NET0131 ,
		\g432_reg/NET0131 ,
		_w4258_
	);
	LUT4 #(
		.INIT('h135f)
	) name3078 (
		\g1088_reg/NET0131 ,
		\g429_reg/NET0131 ,
		\g435_reg/NET0131 ,
		\g7961_pad ,
		_w4259_
	);
	LUT2 #(
		.INIT('h4)
	) name3079 (
		_w4258_,
		_w4259_,
		_w4260_
	);
	LUT2 #(
		.INIT('h8)
	) name3080 (
		\g1092_reg/NET0131 ,
		\g441_reg/NET0131 ,
		_w4261_
	);
	LUT4 #(
		.INIT('h135f)
	) name3081 (
		\g1088_reg/NET0131 ,
		\g438_reg/NET0131 ,
		\g444_reg/NET0131 ,
		\g7961_pad ,
		_w4262_
	);
	LUT2 #(
		.INIT('h4)
	) name3082 (
		_w4261_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('hb)
	) name3083 (
		_w4261_,
		_w4262_,
		_w4264_
	);
	LUT2 #(
		.INIT('h2)
	) name3084 (
		\g1092_reg/NET0131 ,
		\g179_reg/NET0131 ,
		_w4265_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3085 (
		\g1088_reg/NET0131 ,
		\g177_reg/NET0131 ,
		\g178_reg/NET0131 ,
		\g7961_pad ,
		_w4266_
	);
	LUT4 #(
		.INIT('h8088)
	) name3086 (
		_w3948_,
		_w3949_,
		_w4265_,
		_w4266_,
		_w4267_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3087 (
		\g1092_reg/NET0131 ,
		\g448_reg/NET0131 ,
		\g449_reg/NET0131 ,
		\g7961_pad ,
		_w4268_
	);
	LUT2 #(
		.INIT('h2)
	) name3088 (
		\g1088_reg/NET0131 ,
		\g447_reg/NET0131 ,
		_w4269_
	);
	LUT3 #(
		.INIT('hc4)
	) name3089 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g447_reg/NET0131 ,
		_w4270_
	);
	LUT2 #(
		.INIT('h8)
	) name3090 (
		_w4268_,
		_w4270_,
		_w4271_
	);
	LUT4 #(
		.INIT('h4200)
	) name3091 (
		_w4260_,
		_w4263_,
		_w4267_,
		_w4271_,
		_w4272_
	);
	LUT4 #(
		.INIT('hbdff)
	) name3092 (
		_w4260_,
		_w4263_,
		_w4267_,
		_w4271_,
		_w4273_
	);
	LUT4 #(
		.INIT('h8002)
	) name3093 (
		\g1563_reg/NET0131 ,
		_w4260_,
		_w4263_,
		_w4267_,
		_w4274_
	);
	LUT3 #(
		.INIT('ha8)
	) name3094 (
		\g7961_pad ,
		_w4272_,
		_w4274_,
		_w4275_
	);
	LUT3 #(
		.INIT('h80)
	) name3095 (
		\g1088_reg/NET0131 ,
		\g1462_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		_w4276_
	);
	LUT3 #(
		.INIT('h80)
	) name3096 (
		\g1448_reg/NET0131 ,
		\g1453_reg/NET0131 ,
		\g1457_reg/NET0131 ,
		_w4277_
	);
	LUT4 #(
		.INIT('h7000)
	) name3097 (
		_w4071_,
		_w4072_,
		_w4276_,
		_w4277_,
		_w4278_
	);
	LUT3 #(
		.INIT('h80)
	) name3098 (
		\g1435_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		_w4279_
	);
	LUT2 #(
		.INIT('h8)
	) name3099 (
		\g1426_reg/NET0131 ,
		\g1430_reg/NET0131 ,
		_w4280_
	);
	LUT2 #(
		.INIT('h8)
	) name3100 (
		_w4279_,
		_w4280_,
		_w4281_
	);
	LUT4 #(
		.INIT('h0008)
	) name3101 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g2896_reg/NET0131 ,
		\g2900_reg/NET0131 ,
		_w4282_
	);
	LUT2 #(
		.INIT('h8)
	) name3102 (
		_w4072_,
		_w4282_,
		_w4283_
	);
	LUT3 #(
		.INIT('h2a)
	) name3103 (
		\g1426_reg/NET0131 ,
		_w4072_,
		_w4282_,
		_w4284_
	);
	LUT4 #(
		.INIT('h8000)
	) name3104 (
		\g1430_reg/NET0131 ,
		\g1435_reg/NET0131 ,
		\g1439_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		_w4285_
	);
	LUT3 #(
		.INIT('h70)
	) name3105 (
		_w4072_,
		_w4282_,
		_w4285_,
		_w4286_
	);
	LUT4 #(
		.INIT('h7270)
	) name3106 (
		_w4278_,
		_w4281_,
		_w4284_,
		_w4286_,
		_w4287_
	);
	LUT3 #(
		.INIT('ha8)
	) name3107 (
		\g1088_reg/NET0131 ,
		_w4272_,
		_w4274_,
		_w4288_
	);
	LUT3 #(
		.INIT('ha8)
	) name3108 (
		\g1092_reg/NET0131 ,
		_w4272_,
		_w4274_,
		_w4289_
	);
	LUT2 #(
		.INIT('h2)
	) name3109 (
		\g1088_reg/NET0131 ,
		\g1134_reg/NET0131 ,
		_w4290_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3110 (
		\g1092_reg/NET0131 ,
		\g1135_reg/NET0131 ,
		\g1136_reg/NET0131 ,
		\g7961_pad ,
		_w4291_
	);
	LUT2 #(
		.INIT('h4)
	) name3111 (
		_w4290_,
		_w4291_,
		_w4292_
	);
	LUT2 #(
		.INIT('h8)
	) name3112 (
		\g1092_reg/NET0131 ,
		\g1128_reg/NET0131 ,
		_w4293_
	);
	LUT4 #(
		.INIT('h135f)
	) name3113 (
		\g1088_reg/NET0131 ,
		\g1125_reg/NET0131 ,
		\g1131_reg/NET0131 ,
		\g7961_pad ,
		_w4294_
	);
	LUT2 #(
		.INIT('h4)
	) name3114 (
		_w4293_,
		_w4294_,
		_w4295_
	);
	LUT2 #(
		.INIT('hb)
	) name3115 (
		_w4293_,
		_w4294_,
		_w4296_
	);
	LUT2 #(
		.INIT('h2)
	) name3116 (
		_w4224_,
		_w4229_,
		_w4297_
	);
	LUT4 #(
		.INIT('h0200)
	) name3117 (
		_w4224_,
		_w4229_,
		_w4293_,
		_w4294_,
		_w4298_
	);
	LUT2 #(
		.INIT('h2)
	) name3118 (
		_w4292_,
		_w4298_,
		_w4299_
	);
	LUT3 #(
		.INIT('h08)
	) name3119 (
		\g1563_reg/NET0131 ,
		_w4224_,
		_w4229_,
		_w4300_
	);
	LUT3 #(
		.INIT('h20)
	) name3120 (
		\g1563_reg/NET0131 ,
		_w4293_,
		_w4294_,
		_w4301_
	);
	LUT3 #(
		.INIT('h1b)
	) name3121 (
		_w4223_,
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('hd)
	) name3122 (
		_w4299_,
		_w4302_,
		_w4303_
	);
	LUT4 #(
		.INIT('h8002)
	) name3123 (
		\g1563_reg/NET0131 ,
		_w4223_,
		_w4295_,
		_w4297_,
		_w4304_
	);
	LUT4 #(
		.INIT('haa08)
	) name3124 (
		\g1088_reg/NET0131 ,
		_w4299_,
		_w4302_,
		_w4304_,
		_w4305_
	);
	LUT4 #(
		.INIT('haa08)
	) name3125 (
		\g7961_pad ,
		_w4299_,
		_w4302_,
		_w4304_,
		_w4306_
	);
	LUT4 #(
		.INIT('haa08)
	) name3126 (
		\g1092_reg/NET0131 ,
		_w4299_,
		_w4302_,
		_w4304_,
		_w4307_
	);
	LUT2 #(
		.INIT('h8)
	) name3127 (
		\g1092_reg/NET0131 ,
		\g2507_reg/NET0131 ,
		_w4308_
	);
	LUT4 #(
		.INIT('h135f)
	) name3128 (
		\g1088_reg/NET0131 ,
		\g2504_reg/NET0131 ,
		\g2510_reg/NET0131 ,
		\g7961_pad ,
		_w4309_
	);
	LUT2 #(
		.INIT('h4)
	) name3129 (
		_w4308_,
		_w4309_,
		_w4310_
	);
	LUT2 #(
		.INIT('h8)
	) name3130 (
		\g1092_reg/NET0131 ,
		\g2516_reg/NET0131 ,
		_w4311_
	);
	LUT4 #(
		.INIT('h135f)
	) name3131 (
		\g1088_reg/NET0131 ,
		\g2513_reg/NET0131 ,
		\g2519_reg/NET0131 ,
		\g7961_pad ,
		_w4312_
	);
	LUT2 #(
		.INIT('h4)
	) name3132 (
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('hb)
	) name3133 (
		_w4311_,
		_w4312_,
		_w4314_
	);
	LUT2 #(
		.INIT('h4)
	) name3134 (
		\g2254_reg/NET0131 ,
		\g7961_pad ,
		_w4315_
	);
	LUT4 #(
		.INIT('hf531)
	) name3135 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2253_reg/NET0131 ,
		\g2255_reg/NET0131 ,
		_w4316_
	);
	LUT4 #(
		.INIT('h8088)
	) name3136 (
		_w3966_,
		_w3967_,
		_w4315_,
		_w4316_,
		_w4317_
	);
	LUT4 #(
		.INIT('hc4f5)
	) name3137 (
		\g1092_reg/NET0131 ,
		\g2523_reg/NET0131 ,
		\g2524_reg/NET0131 ,
		\g7961_pad ,
		_w4318_
	);
	LUT2 #(
		.INIT('h2)
	) name3138 (
		\g1088_reg/NET0131 ,
		\g2522_reg/NET0131 ,
		_w4319_
	);
	LUT3 #(
		.INIT('hc4)
	) name3139 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g2522_reg/NET0131 ,
		_w4320_
	);
	LUT2 #(
		.INIT('h8)
	) name3140 (
		_w4318_,
		_w4320_,
		_w4321_
	);
	LUT4 #(
		.INIT('h4200)
	) name3141 (
		_w4310_,
		_w4313_,
		_w4317_,
		_w4321_,
		_w4322_
	);
	LUT4 #(
		.INIT('hbdff)
	) name3142 (
		_w4310_,
		_w4313_,
		_w4317_,
		_w4321_,
		_w4323_
	);
	LUT4 #(
		.INIT('h8002)
	) name3143 (
		\g1563_reg/NET0131 ,
		_w4310_,
		_w4313_,
		_w4317_,
		_w4324_
	);
	LUT3 #(
		.INIT('ha8)
	) name3144 (
		\g1088_reg/NET0131 ,
		_w4322_,
		_w4324_,
		_w4325_
	);
	LUT3 #(
		.INIT('ha8)
	) name3145 (
		\g7961_pad ,
		_w4322_,
		_w4324_,
		_w4326_
	);
	LUT3 #(
		.INIT('ha8)
	) name3146 (
		\g1092_reg/NET0131 ,
		_w4322_,
		_w4324_,
		_w4327_
	);
	LUT3 #(
		.INIT('h80)
	) name3147 (
		\g1092_reg/NET0131 ,
		_w1848_,
		_w1919_,
		_w4328_
	);
	LUT3 #(
		.INIT('h2a)
	) name3148 (
		\g1092_reg/NET0131 ,
		_w4071_,
		_w4072_,
		_w4329_
	);
	LUT3 #(
		.INIT('h70)
	) name3149 (
		_w1859_,
		_w4107_,
		_w4329_,
		_w4330_
	);
	LUT2 #(
		.INIT('he)
	) name3150 (
		_w4328_,
		_w4330_,
		_w4331_
	);
	LUT2 #(
		.INIT('h4)
	) name3151 (
		\g1056_reg/NET0131 ,
		\g7961_pad ,
		_w4332_
	);
	LUT4 #(
		.INIT('h8acf)
	) name3152 (
		\g1045_reg/NET0131 ,
		\g1048_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w4333_
	);
	LUT2 #(
		.INIT('h4)
	) name3153 (
		_w4332_,
		_w4333_,
		_w4334_
	);
	LUT2 #(
		.INIT('h4)
	) name3154 (
		\g1085_reg/NET0131 ,
		\g7961_pad ,
		_w4335_
	);
	LUT4 #(
		.INIT('h8acf)
	) name3155 (
		\g1075_reg/NET0131 ,
		\g1078_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w4336_
	);
	LUT2 #(
		.INIT('h4)
	) name3156 (
		_w4335_,
		_w4336_,
		_w4337_
	);
	LUT4 #(
		.INIT('h0400)
	) name3157 (
		_w4332_,
		_w4333_,
		_w4335_,
		_w4336_,
		_w4338_
	);
	LUT2 #(
		.INIT('h4)
	) name3158 (
		\g1041_reg/NET0131 ,
		\g7961_pad ,
		_w4339_
	);
	LUT4 #(
		.INIT('h8acf)
	) name3159 (
		\g1030_reg/NET0131 ,
		\g1033_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w4340_
	);
	LUT2 #(
		.INIT('h4)
	) name3160 (
		_w4339_,
		_w4340_,
		_w4341_
	);
	LUT3 #(
		.INIT('h8a)
	) name3161 (
		\g3229_pad ,
		_w4339_,
		_w4340_,
		_w4342_
	);
	LUT3 #(
		.INIT('h23)
	) name3162 (
		\g1041_reg/NET0131 ,
		\g3229_pad ,
		\g7961_pad ,
		_w4343_
	);
	LUT2 #(
		.INIT('h8)
	) name3163 (
		_w4340_,
		_w4343_,
		_w4344_
	);
	LUT3 #(
		.INIT('h65)
	) name3164 (
		\g3229_pad ,
		_w4339_,
		_w4340_,
		_w4345_
	);
	LUT4 #(
		.INIT('h0444)
	) name3165 (
		_w4332_,
		_w4333_,
		_w4340_,
		_w4343_,
		_w4346_
	);
	LUT4 #(
		.INIT('hccc5)
	) name3166 (
		_w4334_,
		_w4338_,
		_w4342_,
		_w4344_,
		_w4347_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3167 (
		\g1060_reg/NET0131 ,
		_w4328_,
		_w4330_,
		_w4347_,
		_w4348_
	);
	LUT3 #(
		.INIT('h80)
	) name3168 (
		\g1088_reg/NET0131 ,
		_w1848_,
		_w1919_,
		_w4349_
	);
	LUT3 #(
		.INIT('h2a)
	) name3169 (
		\g1088_reg/NET0131 ,
		_w4071_,
		_w4072_,
		_w4350_
	);
	LUT3 #(
		.INIT('h70)
	) name3170 (
		_w1859_,
		_w4107_,
		_w4350_,
		_w4351_
	);
	LUT2 #(
		.INIT('he)
	) name3171 (
		_w4349_,
		_w4351_,
		_w4352_
	);
	LUT4 #(
		.INIT('h333a)
	) name3172 (
		\g1063_reg/NET0131 ,
		_w4347_,
		_w4349_,
		_w4351_,
		_w4353_
	);
	LUT3 #(
		.INIT('h80)
	) name3173 (
		\g7961_pad ,
		_w1848_,
		_w1919_,
		_w4354_
	);
	LUT3 #(
		.INIT('h2a)
	) name3174 (
		\g7961_pad ,
		_w4071_,
		_w4072_,
		_w4355_
	);
	LUT3 #(
		.INIT('h70)
	) name3175 (
		_w1859_,
		_w4107_,
		_w4355_,
		_w4356_
	);
	LUT2 #(
		.INIT('he)
	) name3176 (
		_w4354_,
		_w4356_,
		_w4357_
	);
	LUT4 #(
		.INIT('h333a)
	) name3177 (
		\g1071_reg/NET0131 ,
		_w4347_,
		_w4354_,
		_w4356_,
		_w4358_
	);
	LUT4 #(
		.INIT('h135f)
	) name3178 (
		\g1024_reg/NET0131 ,
		\g1871_reg/NET0131 ,
		\g1877_reg/NET0131 ,
		\g5657_pad ,
		_w4359_
	);
	LUT2 #(
		.INIT('h8)
	) name3179 (
		\g1018_reg/NET0131 ,
		\g1874_reg/NET0131 ,
		_w4360_
	);
	LUT3 #(
		.INIT('h4c)
	) name3180 (
		\g1018_reg/NET0131 ,
		\g1196_reg/NET0131 ,
		\g1874_reg/NET0131 ,
		_w4361_
	);
	LUT4 #(
		.INIT('hb000)
	) name3181 (
		_w1576_,
		_w1577_,
		_w4359_,
		_w4361_,
		_w4362_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name3182 (
		_w1572_,
		_w1573_,
		_w4359_,
		_w4360_,
		_w4363_
	);
	LUT2 #(
		.INIT('h1)
	) name3183 (
		\g3002_reg/NET0131 ,
		\g3006_reg/NET0131 ,
		_w4364_
	);
	LUT3 #(
		.INIT('h01)
	) name3184 (
		\g3010_reg/NET0131 ,
		\g3013_reg/NET0131 ,
		\g3024_reg/NET0131 ,
		_w4365_
	);
	LUT2 #(
		.INIT('h8)
	) name3185 (
		_w4364_,
		_w4365_,
		_w4366_
	);
	LUT4 #(
		.INIT('h7775)
	) name3186 (
		\g1024_reg/NET0131 ,
		_w4362_,
		_w4363_,
		_w4366_,
		_w4367_
	);
	LUT4 #(
		.INIT('h888a)
	) name3187 (
		\g1024_reg/NET0131 ,
		_w4362_,
		_w4363_,
		_w4366_,
		_w4368_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3188 (
		_w3697_,
		_w3698_,
		_w3713_,
		_w3714_,
		_w4369_
	);
	LUT3 #(
		.INIT('h01)
	) name3189 (
		\g3229_pad ,
		_w3710_,
		_w4369_,
		_w4370_
	);
	LUT4 #(
		.INIT('h0008)
	) name3190 (
		\g3229_pad ,
		_w3715_,
		_w3718_,
		_w3742_,
		_w4371_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3191 (
		\g1955_reg/NET0131 ,
		_w4367_,
		_w4370_,
		_w4371_,
		_w4372_
	);
	LUT4 #(
		.INIT('h7775)
	) name3192 (
		\g5657_pad ,
		_w4362_,
		_w4363_,
		_w4366_,
		_w4373_
	);
	LUT4 #(
		.INIT('h888a)
	) name3193 (
		\g5657_pad ,
		_w4362_,
		_w4363_,
		_w4366_,
		_w4374_
	);
	LUT4 #(
		.INIT('haafc)
	) name3194 (
		\g1956_reg/NET0131 ,
		_w4370_,
		_w4371_,
		_w4373_,
		_w4375_
	);
	LUT4 #(
		.INIT('h7775)
	) name3195 (
		\g1018_reg/NET0131 ,
		_w4362_,
		_w4363_,
		_w4366_,
		_w4376_
	);
	LUT4 #(
		.INIT('h888a)
	) name3196 (
		\g1018_reg/NET0131 ,
		_w4362_,
		_w4363_,
		_w4366_,
		_w4377_
	);
	LUT4 #(
		.INIT('haafc)
	) name3197 (
		\g1957_reg/NET0131 ,
		_w4370_,
		_w4371_,
		_w4376_,
		_w4378_
	);
	LUT3 #(
		.INIT('h80)
	) name3198 (
		\g1092_reg/NET0131 ,
		_w1697_,
		_w1821_,
		_w4379_
	);
	LUT3 #(
		.INIT('hb0)
	) name3199 (
		_w1747_,
		_w4074_,
		_w4329_,
		_w4380_
	);
	LUT2 #(
		.INIT('he)
	) name3200 (
		_w4379_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h4)
	) name3201 (
		\g398_reg/NET0131 ,
		\g7961_pad ,
		_w4382_
	);
	LUT4 #(
		.INIT('hf351)
	) name3202 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g388_reg/NET0131 ,
		\g391_reg/NET0131 ,
		_w4383_
	);
	LUT2 #(
		.INIT('h4)
	) name3203 (
		_w4382_,
		_w4383_,
		_w4384_
	);
	LUT2 #(
		.INIT('h4)
	) name3204 (
		\g354_reg/NET0131 ,
		\g7961_pad ,
		_w4385_
	);
	LUT4 #(
		.INIT('hf351)
	) name3205 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g343_reg/NET0131 ,
		\g346_reg/NET0131 ,
		_w4386_
	);
	LUT2 #(
		.INIT('h4)
	) name3206 (
		_w4385_,
		_w4386_,
		_w4387_
	);
	LUT2 #(
		.INIT('h4)
	) name3207 (
		\g369_reg/NET0131 ,
		\g7961_pad ,
		_w4388_
	);
	LUT4 #(
		.INIT('hf351)
	) name3208 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g358_reg/NET0131 ,
		\g361_reg/NET0131 ,
		_w4389_
	);
	LUT2 #(
		.INIT('h4)
	) name3209 (
		_w4388_,
		_w4389_,
		_w4390_
	);
	LUT2 #(
		.INIT('h2)
	) name3210 (
		\g1092_reg/NET0131 ,
		\g373_reg/NET0131 ,
		_w4391_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3211 (
		\g1088_reg/NET0131 ,
		\g376_reg/NET0131 ,
		\g384_reg/NET0131 ,
		\g7961_pad ,
		_w4392_
	);
	LUT2 #(
		.INIT('h4)
	) name3212 (
		_w4391_,
		_w4392_,
		_w4393_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3213 (
		_w4388_,
		_w4389_,
		_w4391_,
		_w4392_,
		_w4394_
	);
	LUT3 #(
		.INIT('h8a)
	) name3214 (
		\g3229_pad ,
		_w4385_,
		_w4386_,
		_w4395_
	);
	LUT4 #(
		.INIT('h88d1)
	) name3215 (
		\g3229_pad ,
		_w4384_,
		_w4387_,
		_w4394_,
		_w4396_
	);
	LUT4 #(
		.INIT('hfe02)
	) name3216 (
		\g343_reg/NET0131 ,
		_w4379_,
		_w4380_,
		_w4396_,
		_w4397_
	);
	LUT3 #(
		.INIT('h80)
	) name3217 (
		\g1088_reg/NET0131 ,
		_w1697_,
		_w1821_,
		_w4398_
	);
	LUT3 #(
		.INIT('hb0)
	) name3218 (
		_w1747_,
		_w4074_,
		_w4350_,
		_w4399_
	);
	LUT2 #(
		.INIT('he)
	) name3219 (
		_w4398_,
		_w4399_,
		_w4400_
	);
	LUT4 #(
		.INIT('hccca)
	) name3220 (
		\g346_reg/NET0131 ,
		_w4396_,
		_w4398_,
		_w4399_,
		_w4401_
	);
	LUT3 #(
		.INIT('h80)
	) name3221 (
		\g7961_pad ,
		_w1697_,
		_w1821_,
		_w4402_
	);
	LUT3 #(
		.INIT('hb0)
	) name3222 (
		_w1747_,
		_w4074_,
		_w4355_,
		_w4403_
	);
	LUT2 #(
		.INIT('he)
	) name3223 (
		_w4402_,
		_w4403_,
		_w4404_
	);
	LUT4 #(
		.INIT('hccca)
	) name3224 (
		\g354_reg/NET0131 ,
		_w4396_,
		_w4402_,
		_w4403_,
		_w4405_
	);
	LUT3 #(
		.INIT('h45)
	) name3225 (
		\g3229_pad ,
		\g354_reg/NET0131 ,
		\g7961_pad ,
		_w4406_
	);
	LUT2 #(
		.INIT('h8)
	) name3226 (
		_w4386_,
		_w4406_,
		_w4407_
	);
	LUT4 #(
		.INIT('h1030)
	) name3227 (
		_w4386_,
		_w4388_,
		_w4389_,
		_w4406_,
		_w4408_
	);
	LUT3 #(
		.INIT('h65)
	) name3228 (
		\g3229_pad ,
		_w4385_,
		_w4386_,
		_w4409_
	);
	LUT4 #(
		.INIT('h0400)
	) name3229 (
		_w4382_,
		_w4383_,
		_w4388_,
		_w4389_,
		_w4410_
	);
	LUT4 #(
		.INIT('hfd01)
	) name3230 (
		_w4390_,
		_w4395_,
		_w4407_,
		_w4410_,
		_w4411_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3231 (
		\g373_reg/NET0131 ,
		_w4379_,
		_w4380_,
		_w4411_,
		_w4412_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3232 (
		\g376_reg/NET0131 ,
		_w4398_,
		_w4399_,
		_w4411_,
		_w4413_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3233 (
		\g384_reg/NET0131 ,
		_w4402_,
		_w4403_,
		_w4411_,
		_w4414_
	);
	LUT4 #(
		.INIT('h135f)
	) name3234 (
		\g1024_reg/NET0131 ,
		\g490_reg/NET0131 ,
		\g496_reg/NET0131 ,
		\g5657_pad ,
		_w4415_
	);
	LUT2 #(
		.INIT('h8)
	) name3235 (
		\g1018_reg/NET0131 ,
		\g493_reg/NET0131 ,
		_w4416_
	);
	LUT3 #(
		.INIT('h4c)
	) name3236 (
		\g1018_reg/NET0131 ,
		\g1196_reg/NET0131 ,
		\g493_reg/NET0131 ,
		_w4417_
	);
	LUT4 #(
		.INIT('hb000)
	) name3237 (
		_w2863_,
		_w2864_,
		_w4415_,
		_w4417_,
		_w4418_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name3238 (
		_w2859_,
		_w2860_,
		_w4415_,
		_w4416_,
		_w4419_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3239 (
		\g1024_reg/NET0131 ,
		_w4366_,
		_w4418_,
		_w4419_,
		_w4420_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3240 (
		\g1024_reg/NET0131 ,
		_w4366_,
		_w4418_,
		_w4419_,
		_w4421_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3241 (
		_w3763_,
		_w3764_,
		_w3788_,
		_w3789_,
		_w4422_
	);
	LUT3 #(
		.INIT('h01)
	) name3242 (
		\g3229_pad ,
		_w3805_,
		_w4422_,
		_w4423_
	);
	LUT4 #(
		.INIT('h0200)
	) name3243 (
		\g3229_pad ,
		_w3769_,
		_w3780_,
		_w3790_,
		_w4424_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3244 (
		\g575_reg/NET0131 ,
		_w4420_,
		_w4423_,
		_w4424_,
		_w4425_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3245 (
		\g5657_pad ,
		_w4366_,
		_w4418_,
		_w4419_,
		_w4426_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3246 (
		\g5657_pad ,
		_w4366_,
		_w4418_,
		_w4419_,
		_w4427_
	);
	LUT4 #(
		.INIT('haafc)
	) name3247 (
		\g576_reg/NET0131 ,
		_w4423_,
		_w4424_,
		_w4426_,
		_w4428_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3248 (
		\g1018_reg/NET0131 ,
		_w4366_,
		_w4418_,
		_w4419_,
		_w4429_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3249 (
		\g1018_reg/NET0131 ,
		_w4366_,
		_w4418_,
		_w4419_,
		_w4430_
	);
	LUT4 #(
		.INIT('haafc)
	) name3250 (
		\g577_reg/NET0131 ,
		_w4423_,
		_w4424_,
		_w4429_,
		_w4431_
	);
	LUT4 #(
		.INIT('hfe0e)
	) name3251 (
		\g1018_reg/NET0131 ,
		\g16297_pad ,
		\g506_reg/NET0131 ,
		\g507_reg/NET0131 ,
		_w4432_
	);
	LUT4 #(
		.INIT('h135f)
	) name3252 (
		\g1024_reg/NET0131 ,
		\g1177_reg/NET0131 ,
		\g1183_reg/NET0131 ,
		\g5657_pad ,
		_w4433_
	);
	LUT2 #(
		.INIT('h8)
	) name3253 (
		\g1018_reg/NET0131 ,
		\g1180_reg/NET0131 ,
		_w4434_
	);
	LUT3 #(
		.INIT('h70)
	) name3254 (
		\g1018_reg/NET0131 ,
		\g1180_reg/NET0131 ,
		\g1196_reg/NET0131 ,
		_w4435_
	);
	LUT4 #(
		.INIT('hb000)
	) name3255 (
		_w2206_,
		_w2207_,
		_w4433_,
		_w4435_,
		_w4436_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name3256 (
		_w2210_,
		_w2211_,
		_w4433_,
		_w4434_,
		_w4437_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3257 (
		\g1024_reg/NET0131 ,
		_w4366_,
		_w4436_,
		_w4437_,
		_w4438_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3258 (
		\g1024_reg/NET0131 ,
		_w4366_,
		_w4436_,
		_w4437_,
		_w4439_
	);
	LUT3 #(
		.INIT('h01)
	) name3259 (
		\g3229_pad ,
		_w3276_,
		_w3279_,
		_w4440_
	);
	LUT4 #(
		.INIT('h0020)
	) name3260 (
		\g3229_pad ,
		_w3232_,
		_w3250_,
		_w3288_,
		_w4441_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3261 (
		\g1261_reg/NET0131 ,
		_w4438_,
		_w4440_,
		_w4441_,
		_w4442_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3262 (
		\g5657_pad ,
		_w4366_,
		_w4436_,
		_w4437_,
		_w4443_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3263 (
		\g5657_pad ,
		_w4366_,
		_w4436_,
		_w4437_,
		_w4444_
	);
	LUT4 #(
		.INIT('haafc)
	) name3264 (
		\g1262_reg/NET0131 ,
		_w4440_,
		_w4441_,
		_w4443_,
		_w4445_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3265 (
		\g1018_reg/NET0131 ,
		_w4366_,
		_w4436_,
		_w4437_,
		_w4446_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3266 (
		\g1018_reg/NET0131 ,
		_w4366_,
		_w4436_,
		_w4437_,
		_w4447_
	);
	LUT4 #(
		.INIT('haafc)
	) name3267 (
		\g1263_reg/NET0131 ,
		_w4440_,
		_w4441_,
		_w4446_,
		_w4448_
	);
	LUT4 #(
		.INIT('hb4bb)
	) name3268 (
		_w3226_,
		_w3227_,
		_w3229_,
		_w3230_,
		_w4449_
	);
	LUT4 #(
		.INIT('h4044)
	) name3269 (
		_w3229_,
		_w3230_,
		_w3248_,
		_w3249_,
		_w4450_
	);
	LUT3 #(
		.INIT('hf9)
	) name3270 (
		\g3229_pad ,
		_w4449_,
		_w4450_,
		_w4451_
	);
	LUT3 #(
		.INIT('hb8)
	) name3271 (
		\g1267_reg/NET0131 ,
		_w4438_,
		_w4451_,
		_w4452_
	);
	LUT3 #(
		.INIT('h80)
	) name3272 (
		\g1092_reg/NET0131 ,
		_w1368_,
		_w1369_,
		_w4453_
	);
	LUT3 #(
		.INIT('h70)
	) name3273 (
		_w1364_,
		_w4161_,
		_w4329_,
		_w4454_
	);
	LUT2 #(
		.INIT('he)
	) name3274 (
		_w4453_,
		_w4454_,
		_w4455_
	);
	LUT2 #(
		.INIT('h4)
	) name3275 (
		\g2473_reg/NET0131 ,
		\g7961_pad ,
		_w4456_
	);
	LUT4 #(
		.INIT('hf351)
	) name3276 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2463_reg/NET0131 ,
		\g2466_reg/NET0131 ,
		_w4457_
	);
	LUT2 #(
		.INIT('h4)
	) name3277 (
		_w4456_,
		_w4457_,
		_w4458_
	);
	LUT2 #(
		.INIT('h4)
	) name3278 (
		\g2429_reg/NET0131 ,
		\g7961_pad ,
		_w4459_
	);
	LUT4 #(
		.INIT('hf351)
	) name3279 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2418_reg/NET0131 ,
		\g2421_reg/NET0131 ,
		_w4460_
	);
	LUT2 #(
		.INIT('h4)
	) name3280 (
		_w4459_,
		_w4460_,
		_w4461_
	);
	LUT2 #(
		.INIT('h4)
	) name3281 (
		\g2444_reg/NET0131 ,
		\g7961_pad ,
		_w4462_
	);
	LUT4 #(
		.INIT('hf351)
	) name3282 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2433_reg/NET0131 ,
		\g2436_reg/NET0131 ,
		_w4463_
	);
	LUT2 #(
		.INIT('h4)
	) name3283 (
		_w4462_,
		_w4463_,
		_w4464_
	);
	LUT2 #(
		.INIT('h2)
	) name3284 (
		\g1092_reg/NET0131 ,
		\g2448_reg/NET0131 ,
		_w4465_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3285 (
		\g1088_reg/NET0131 ,
		\g2451_reg/NET0131 ,
		\g2459_reg/NET0131 ,
		\g7961_pad ,
		_w4466_
	);
	LUT2 #(
		.INIT('h4)
	) name3286 (
		_w4465_,
		_w4466_,
		_w4467_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3287 (
		_w4462_,
		_w4463_,
		_w4465_,
		_w4466_,
		_w4468_
	);
	LUT3 #(
		.INIT('h8a)
	) name3288 (
		\g3229_pad ,
		_w4459_,
		_w4460_,
		_w4469_
	);
	LUT4 #(
		.INIT('h88d1)
	) name3289 (
		\g3229_pad ,
		_w4458_,
		_w4461_,
		_w4468_,
		_w4470_
	);
	LUT4 #(
		.INIT('hfe02)
	) name3290 (
		\g2418_reg/NET0131 ,
		_w4453_,
		_w4454_,
		_w4470_,
		_w4471_
	);
	LUT3 #(
		.INIT('hb8)
	) name3291 (
		\g1268_reg/NET0131 ,
		_w4443_,
		_w4451_,
		_w4472_
	);
	LUT3 #(
		.INIT('hb8)
	) name3292 (
		\g1269_reg/NET0131 ,
		_w4446_,
		_w4451_,
		_w4473_
	);
	LUT3 #(
		.INIT('h80)
	) name3293 (
		\g1088_reg/NET0131 ,
		_w1368_,
		_w1369_,
		_w4474_
	);
	LUT3 #(
		.INIT('h70)
	) name3294 (
		_w1364_,
		_w4161_,
		_w4350_,
		_w4475_
	);
	LUT2 #(
		.INIT('he)
	) name3295 (
		_w4474_,
		_w4475_,
		_w4476_
	);
	LUT4 #(
		.INIT('hccca)
	) name3296 (
		\g2421_reg/NET0131 ,
		_w4470_,
		_w4474_,
		_w4475_,
		_w4477_
	);
	LUT3 #(
		.INIT('h80)
	) name3297 (
		\g7961_pad ,
		_w1368_,
		_w1369_,
		_w4478_
	);
	LUT3 #(
		.INIT('h70)
	) name3298 (
		_w1364_,
		_w4161_,
		_w4355_,
		_w4479_
	);
	LUT2 #(
		.INIT('he)
	) name3299 (
		_w4478_,
		_w4479_,
		_w4480_
	);
	LUT4 #(
		.INIT('hccca)
	) name3300 (
		\g2429_reg/NET0131 ,
		_w4470_,
		_w4478_,
		_w4479_,
		_w4481_
	);
	LUT3 #(
		.INIT('h23)
	) name3301 (
		\g2429_reg/NET0131 ,
		\g3229_pad ,
		\g7961_pad ,
		_w4482_
	);
	LUT2 #(
		.INIT('h8)
	) name3302 (
		_w4460_,
		_w4482_,
		_w4483_
	);
	LUT4 #(
		.INIT('h1030)
	) name3303 (
		_w4460_,
		_w4462_,
		_w4463_,
		_w4482_,
		_w4484_
	);
	LUT3 #(
		.INIT('h65)
	) name3304 (
		\g3229_pad ,
		_w4459_,
		_w4460_,
		_w4485_
	);
	LUT4 #(
		.INIT('h0400)
	) name3305 (
		_w4456_,
		_w4457_,
		_w4462_,
		_w4463_,
		_w4486_
	);
	LUT4 #(
		.INIT('hfd01)
	) name3306 (
		_w4464_,
		_w4469_,
		_w4483_,
		_w4486_,
		_w4487_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3307 (
		\g2448_reg/NET0131 ,
		_w4453_,
		_w4454_,
		_w4487_,
		_w4488_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3308 (
		\g2451_reg/NET0131 ,
		_w4474_,
		_w4475_,
		_w4487_,
		_w4489_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3309 (
		\g2459_reg/NET0131 ,
		_w4478_,
		_w4479_,
		_w4487_,
		_w4490_
	);
	LUT2 #(
		.INIT('h4)
	) name3310 (
		\g1060_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		_w4491_
	);
	LUT4 #(
		.INIT('h8caf)
	) name3311 (
		\g1063_reg/NET0131 ,
		\g1071_reg/NET0131 ,
		\g1088_reg/NET0131 ,
		\g7961_pad ,
		_w4492_
	);
	LUT2 #(
		.INIT('h4)
	) name3312 (
		_w4491_,
		_w4492_,
		_w4493_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3313 (
		_w4332_,
		_w4333_,
		_w4491_,
		_w4492_,
		_w4494_
	);
	LUT4 #(
		.INIT('h88d1)
	) name3314 (
		\g3229_pad ,
		_w4337_,
		_w4341_,
		_w4494_,
		_w4495_
	);
	LUT4 #(
		.INIT('hfe02)
	) name3315 (
		\g1030_reg/NET0131 ,
		_w4328_,
		_w4330_,
		_w4495_,
		_w4496_
	);
	LUT4 #(
		.INIT('h135f)
	) name3316 (
		\g1024_reg/NET0131 ,
		\g2565_reg/NET0131 ,
		\g2571_reg/NET0131 ,
		\g5657_pad ,
		_w4497_
	);
	LUT2 #(
		.INIT('h8)
	) name3317 (
		\g1018_reg/NET0131 ,
		\g2568_reg/NET0131 ,
		_w4498_
	);
	LUT3 #(
		.INIT('h4c)
	) name3318 (
		\g1018_reg/NET0131 ,
		\g1196_reg/NET0131 ,
		\g2568_reg/NET0131 ,
		_w4499_
	);
	LUT4 #(
		.INIT('hb000)
	) name3319 (
		_w1417_,
		_w1418_,
		_w4497_,
		_w4499_,
		_w4500_
	);
	LUT4 #(
		.INIT('hbb0b)
	) name3320 (
		_w1457_,
		_w1458_,
		_w4497_,
		_w4498_,
		_w4501_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3321 (
		\g1024_reg/NET0131 ,
		_w4366_,
		_w4500_,
		_w4501_,
		_w4502_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3322 (
		\g1024_reg/NET0131 ,
		_w4366_,
		_w4500_,
		_w4501_,
		_w4503_
	);
	LUT3 #(
		.INIT('h01)
	) name3323 (
		\g3229_pad ,
		_w3361_,
		_w3368_,
		_w4504_
	);
	LUT4 #(
		.INIT('h0200)
	) name3324 (
		\g3229_pad ,
		_w3334_,
		_w3339_,
		_w3350_,
		_w4505_
	);
	LUT4 #(
		.INIT('hbbb8)
	) name3325 (
		\g2649_reg/NET0131 ,
		_w4502_,
		_w4504_,
		_w4505_,
		_w4506_
	);
	LUT3 #(
		.INIT('h80)
	) name3326 (
		\g1092_reg/NET0131 ,
		_w2129_,
		_w2143_,
		_w4507_
	);
	LUT3 #(
		.INIT('h70)
	) name3327 (
		_w2121_,
		_w4198_,
		_w4329_,
		_w4508_
	);
	LUT2 #(
		.INIT('he)
	) name3328 (
		_w4507_,
		_w4508_,
		_w4509_
	);
	LUT2 #(
		.INIT('h4)
	) name3329 (
		\g1779_reg/NET0131 ,
		\g7961_pad ,
		_w4510_
	);
	LUT4 #(
		.INIT('hf351)
	) name3330 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1769_reg/NET0131 ,
		\g1772_reg/NET0131 ,
		_w4511_
	);
	LUT2 #(
		.INIT('h4)
	) name3331 (
		_w4510_,
		_w4511_,
		_w4512_
	);
	LUT2 #(
		.INIT('h4)
	) name3332 (
		\g1735_reg/NET0131 ,
		\g7961_pad ,
		_w4513_
	);
	LUT4 #(
		.INIT('hf351)
	) name3333 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1724_reg/NET0131 ,
		\g1727_reg/NET0131 ,
		_w4514_
	);
	LUT2 #(
		.INIT('h4)
	) name3334 (
		_w4513_,
		_w4514_,
		_w4515_
	);
	LUT2 #(
		.INIT('h4)
	) name3335 (
		\g1750_reg/NET0131 ,
		\g7961_pad ,
		_w4516_
	);
	LUT4 #(
		.INIT('hf351)
	) name3336 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1739_reg/NET0131 ,
		\g1742_reg/NET0131 ,
		_w4517_
	);
	LUT2 #(
		.INIT('h4)
	) name3337 (
		_w4516_,
		_w4517_,
		_w4518_
	);
	LUT2 #(
		.INIT('h2)
	) name3338 (
		\g1092_reg/NET0131 ,
		\g1754_reg/NET0131 ,
		_w4519_
	);
	LUT4 #(
		.INIT('hd0dd)
	) name3339 (
		\g1088_reg/NET0131 ,
		\g1757_reg/NET0131 ,
		\g1765_reg/NET0131 ,
		\g7961_pad ,
		_w4520_
	);
	LUT2 #(
		.INIT('h4)
	) name3340 (
		_w4519_,
		_w4520_,
		_w4521_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3341 (
		_w4516_,
		_w4517_,
		_w4519_,
		_w4520_,
		_w4522_
	);
	LUT3 #(
		.INIT('h8a)
	) name3342 (
		\g3229_pad ,
		_w4513_,
		_w4514_,
		_w4523_
	);
	LUT4 #(
		.INIT('h88d1)
	) name3343 (
		\g3229_pad ,
		_w4512_,
		_w4515_,
		_w4522_,
		_w4524_
	);
	LUT4 #(
		.INIT('hfe02)
	) name3344 (
		\g1724_reg/NET0131 ,
		_w4507_,
		_w4508_,
		_w4524_,
		_w4525_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3345 (
		\g5657_pad ,
		_w4366_,
		_w4500_,
		_w4501_,
		_w4526_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3346 (
		\g5657_pad ,
		_w4366_,
		_w4500_,
		_w4501_,
		_w4527_
	);
	LUT4 #(
		.INIT('haafc)
	) name3347 (
		\g2650_reg/NET0131 ,
		_w4504_,
		_w4505_,
		_w4526_,
		_w4528_
	);
	LUT4 #(
		.INIT('h5f5d)
	) name3348 (
		\g1018_reg/NET0131 ,
		_w4366_,
		_w4500_,
		_w4501_,
		_w4529_
	);
	LUT4 #(
		.INIT('ha0a2)
	) name3349 (
		\g1018_reg/NET0131 ,
		_w4366_,
		_w4500_,
		_w4501_,
		_w4530_
	);
	LUT4 #(
		.INIT('haafc)
	) name3350 (
		\g2651_reg/NET0131 ,
		_w4504_,
		_w4505_,
		_w4529_,
		_w4531_
	);
	LUT3 #(
		.INIT('h23)
	) name3351 (
		\g2659_reg/NET0131 ,
		\g3229_pad ,
		\g5657_pad ,
		_w4532_
	);
	LUT2 #(
		.INIT('h8)
	) name3352 (
		_w3349_,
		_w4532_,
		_w4533_
	);
	LUT4 #(
		.INIT('h3efe)
	) name3353 (
		\g3229_pad ,
		_w3330_,
		_w3333_,
		_w4533_,
		_w4534_
	);
	LUT3 #(
		.INIT('h8c)
	) name3354 (
		\g2650_reg/NET0131 ,
		\g3229_pad ,
		\g5657_pad ,
		_w4535_
	);
	LUT4 #(
		.INIT('hb000)
	) name3355 (
		_w3328_,
		_w3329_,
		_w3332_,
		_w4535_,
		_w4536_
	);
	LUT3 #(
		.INIT('h8c)
	) name3356 (
		\g2659_reg/NET0131 ,
		\g3229_pad ,
		\g5657_pad ,
		_w4537_
	);
	LUT2 #(
		.INIT('h8)
	) name3357 (
		_w3349_,
		_w4537_,
		_w4538_
	);
	LUT3 #(
		.INIT('h13)
	) name3358 (
		_w3334_,
		_w4536_,
		_w4538_,
		_w4539_
	);
	LUT4 #(
		.INIT('hb888)
	) name3359 (
		\g2655_reg/NET0131 ,
		_w4502_,
		_w4534_,
		_w4539_,
		_w4540_
	);
	LUT4 #(
		.INIT('hb888)
	) name3360 (
		\g2656_reg/NET0131 ,
		_w4526_,
		_w4534_,
		_w4539_,
		_w4541_
	);
	LUT4 #(
		.INIT('hb888)
	) name3361 (
		\g2657_reg/NET0131 ,
		_w4529_,
		_w4534_,
		_w4539_,
		_w4542_
	);
	LUT3 #(
		.INIT('h80)
	) name3362 (
		\g1088_reg/NET0131 ,
		_w2129_,
		_w2143_,
		_w4543_
	);
	LUT3 #(
		.INIT('h70)
	) name3363 (
		_w2121_,
		_w4198_,
		_w4350_,
		_w4544_
	);
	LUT2 #(
		.INIT('he)
	) name3364 (
		_w4543_,
		_w4544_,
		_w4545_
	);
	LUT4 #(
		.INIT('hccca)
	) name3365 (
		\g1727_reg/NET0131 ,
		_w4524_,
		_w4543_,
		_w4544_,
		_w4546_
	);
	LUT3 #(
		.INIT('h80)
	) name3366 (
		\g7961_pad ,
		_w2129_,
		_w2143_,
		_w4547_
	);
	LUT3 #(
		.INIT('h70)
	) name3367 (
		_w2121_,
		_w4198_,
		_w4355_,
		_w4548_
	);
	LUT2 #(
		.INIT('he)
	) name3368 (
		_w4547_,
		_w4548_,
		_w4549_
	);
	LUT4 #(
		.INIT('hccca)
	) name3369 (
		\g1735_reg/NET0131 ,
		_w4524_,
		_w4547_,
		_w4548_,
		_w4550_
	);
	LUT3 #(
		.INIT('h23)
	) name3370 (
		\g1735_reg/NET0131 ,
		\g3229_pad ,
		\g7961_pad ,
		_w4551_
	);
	LUT2 #(
		.INIT('h8)
	) name3371 (
		_w4514_,
		_w4551_,
		_w4552_
	);
	LUT4 #(
		.INIT('h1030)
	) name3372 (
		_w4514_,
		_w4516_,
		_w4517_,
		_w4551_,
		_w4553_
	);
	LUT3 #(
		.INIT('h65)
	) name3373 (
		\g3229_pad ,
		_w4513_,
		_w4514_,
		_w4554_
	);
	LUT4 #(
		.INIT('h0400)
	) name3374 (
		_w4510_,
		_w4511_,
		_w4516_,
		_w4517_,
		_w4555_
	);
	LUT4 #(
		.INIT('hfd01)
	) name3375 (
		_w4518_,
		_w4523_,
		_w4552_,
		_w4555_,
		_w4556_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3376 (
		\g1754_reg/NET0131 ,
		_w4507_,
		_w4508_,
		_w4556_,
		_w4557_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3377 (
		\g1757_reg/NET0131 ,
		_w4543_,
		_w4544_,
		_w4556_,
		_w4558_
	);
	LUT4 #(
		.INIT('h02fe)
	) name3378 (
		\g1765_reg/NET0131 ,
		_w4547_,
		_w4548_,
		_w4556_,
		_w4559_
	);
	LUT4 #(
		.INIT('hfe02)
	) name3379 (
		\g1033_reg/NET0131 ,
		_w4349_,
		_w4351_,
		_w4495_,
		_w4560_
	);
	LUT4 #(
		.INIT('hfe02)
	) name3380 (
		\g1041_reg/NET0131 ,
		_w4354_,
		_w4356_,
		_w4495_,
		_w4561_
	);
	LUT4 #(
		.INIT('h0322)
	) name3381 (
		_w4214_,
		_w4241_,
		_w4244_,
		_w4247_,
		_w4562_
	);
	LUT2 #(
		.INIT('h2)
	) name3382 (
		_w4214_,
		_w4244_,
		_w4563_
	);
	LUT4 #(
		.INIT('hb393)
	) name3383 (
		\g1563_reg/NET0131 ,
		_w4244_,
		_w4562_,
		_w4563_,
		_w4564_
	);
	LUT4 #(
		.INIT('h0322)
	) name3384 (
		_w4223_,
		_w4292_,
		_w4295_,
		_w4297_,
		_w4565_
	);
	LUT2 #(
		.INIT('h2)
	) name3385 (
		_w4223_,
		_w4295_,
		_w4566_
	);
	LUT4 #(
		.INIT('hb393)
	) name3386 (
		\g1563_reg/NET0131 ,
		_w4295_,
		_w4565_,
		_w4566_,
		_w4567_
	);
	LUT3 #(
		.INIT('ha2)
	) name3387 (
		\g1563_reg/NET0131 ,
		_w4268_,
		_w4269_,
		_w4568_
	);
	LUT4 #(
		.INIT('h7133)
	) name3388 (
		_w4260_,
		_w4263_,
		_w4267_,
		_w4568_,
		_w4569_
	);
	LUT3 #(
		.INIT('ha2)
	) name3389 (
		\g1563_reg/NET0131 ,
		_w4318_,
		_w4319_,
		_w4570_
	);
	LUT4 #(
		.INIT('h7133)
	) name3390 (
		_w4310_,
		_w4313_,
		_w4317_,
		_w4570_,
		_w4571_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3391 (
		_w3919_,
		_w3920_,
		_w3921_,
		_w3922_,
		_w4572_
	);
	LUT3 #(
		.INIT('hef)
	) name3392 (
		_w3999_,
		_w4001_,
		_w4572_,
		_w4573_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3393 (
		_w3937_,
		_w3938_,
		_w3939_,
		_w3940_,
		_w4574_
	);
	LUT3 #(
		.INIT('hef)
	) name3394 (
		_w4005_,
		_w4007_,
		_w4574_,
		_w4575_
	);
	LUT4 #(
		.INIT('h0b00)
	) name3395 (
		_w3955_,
		_w3956_,
		_w3957_,
		_w3958_,
		_w4576_
	);
	LUT3 #(
		.INIT('hef)
	) name3396 (
		_w4011_,
		_w4013_,
		_w4576_,
		_w4577_
	);
	LUT4 #(
		.INIT('h4044)
	) name3397 (
		_w3972_,
		_w3973_,
		_w3974_,
		_w3975_,
		_w4578_
	);
	LUT3 #(
		.INIT('hef)
	) name3398 (
		_w4017_,
		_w4019_,
		_w4578_,
		_w4579_
	);
	LUT4 #(
		.INIT('h4000)
	) name3399 (
		\g3010_reg/NET0131 ,
		\g3013_reg/NET0131 ,
		\g3024_reg/NET0131 ,
		\g3080_reg/NET0131 ,
		_w4580_
	);
	LUT3 #(
		.INIT('h04)
	) name3400 (
		\g3028_reg/NET0131 ,
		\g3032_reg/NET0131 ,
		\g3036_reg/NET0131 ,
		_w4581_
	);
	LUT3 #(
		.INIT('h02)
	) name3401 (
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		\g3234_pad ,
		_w4582_
	);
	LUT4 #(
		.INIT('h0800)
	) name3402 (
		_w3309_,
		_w4580_,
		_w4581_,
		_w4582_,
		_w4583_
	);
	LUT2 #(
		.INIT('h2)
	) name3403 (
		\g3028_reg/NET0131 ,
		\g3234_pad ,
		_w4584_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3404 (
		\g3018_reg/NET0131 ,
		_w3309_,
		_w4580_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('he)
	) name3405 (
		_w4583_,
		_w4585_,
		_w4586_
	);
	LUT3 #(
		.INIT('h0e)
	) name3406 (
		\g1425_reg/NET0131 ,
		_w3562_,
		_w3914_,
		_w4587_
	);
	LUT3 #(
		.INIT('h0e)
	) name3407 (
		\g739_reg/NET0131 ,
		_w3657_,
		_w3914_,
		_w4588_
	);
	LUT3 #(
		.INIT('h13)
	) name3408 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g432_reg/NET0131 ,
		_w4589_
	);
	LUT2 #(
		.INIT('h8)
	) name3409 (
		_w4259_,
		_w4589_,
		_w4590_
	);
	LUT3 #(
		.INIT('h0d)
	) name3410 (
		\g1563_reg/NET0131 ,
		_w4267_,
		_w4590_,
		_w4591_
	);
	LUT3 #(
		.INIT('h13)
	) name3411 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g2507_reg/NET0131 ,
		_w4592_
	);
	LUT2 #(
		.INIT('h8)
	) name3412 (
		_w4309_,
		_w4592_,
		_w4593_
	);
	LUT3 #(
		.INIT('h0d)
	) name3413 (
		\g1563_reg/NET0131 ,
		_w4317_,
		_w4593_,
		_w4594_
	);
	LUT2 #(
		.INIT('h8)
	) name3414 (
		_w4216_,
		_w4246_,
		_w4595_
	);
	LUT3 #(
		.INIT('h0d)
	) name3415 (
		\g1563_reg/NET0131 ,
		_w4214_,
		_w4595_,
		_w4596_
	);
	LUT3 #(
		.INIT('h80)
	) name3416 (
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		\g3036_reg/NET0131 ,
		_w4597_
	);
	LUT3 #(
		.INIT('h80)
	) name3417 (
		_w3309_,
		_w4580_,
		_w4597_,
		_w4598_
	);
	LUT4 #(
		.INIT('h0020)
	) name3418 (
		\g3018_reg/NET0131 ,
		\g3028_reg/NET0131 ,
		\g3032_reg/NET0131 ,
		\g3036_reg/NET0131 ,
		_w4599_
	);
	LUT4 #(
		.INIT('h1555)
	) name3419 (
		\g3234_pad ,
		_w3309_,
		_w4580_,
		_w4599_,
		_w4600_
	);
	LUT4 #(
		.INIT('h1555)
	) name3420 (
		\g3036_reg/NET0131 ,
		_w3309_,
		_w3311_,
		_w4580_,
		_w4601_
	);
	LUT3 #(
		.INIT('h04)
	) name3421 (
		_w4598_,
		_w4600_,
		_w4601_,
		_w4602_
	);
	LUT4 #(
		.INIT('h6aaa)
	) name3422 (
		\g3032_reg/NET0131 ,
		_w3309_,
		_w4580_,
		_w4597_,
		_w4603_
	);
	LUT2 #(
		.INIT('h8)
	) name3423 (
		_w4600_,
		_w4603_,
		_w4604_
	);
	LUT2 #(
		.INIT('h8)
	) name3424 (
		\g1352_reg/NET0131 ,
		\g1358_reg/NET0131 ,
		_w4605_
	);
	LUT3 #(
		.INIT('h80)
	) name3425 (
		_w3908_,
		_w3909_,
		_w4605_,
		_w4606_
	);
	LUT4 #(
		.INIT('h1555)
	) name3426 (
		\g1365_reg/NET0131 ,
		_w3908_,
		_w3909_,
		_w4605_,
		_w4607_
	);
	LUT4 #(
		.INIT('h007f)
	) name3427 (
		_w3908_,
		_w3909_,
		_w3911_,
		_w3914_,
		_w4608_
	);
	LUT2 #(
		.INIT('h4)
	) name3428 (
		_w4607_,
		_w4608_,
		_w4609_
	);
	LUT2 #(
		.INIT('h2)
	) name3429 (
		\g3018_reg/NET0131 ,
		\g3234_pad ,
		_w4610_
	);
	LUT4 #(
		.INIT('h0800)
	) name3430 (
		_w3309_,
		_w4580_,
		_w4581_,
		_w4610_,
		_w4611_
	);
	LUT2 #(
		.INIT('h1)
	) name3431 (
		\g3018_reg/NET0131 ,
		\g3234_pad ,
		_w4612_
	);
	LUT3 #(
		.INIT('h70)
	) name3432 (
		_w3309_,
		_w4580_,
		_w4612_,
		_w4613_
	);
	LUT2 #(
		.INIT('h1)
	) name3433 (
		_w4611_,
		_w4613_,
		_w4614_
	);
	LUT3 #(
		.INIT('h15)
	) name3434 (
		\g3234_pad ,
		_w3309_,
		_w4580_,
		_w4615_
	);
	LUT4 #(
		.INIT('h8000)
	) name3435 (
		\g2993_reg/NET0131 ,
		\g2998_reg/NET0131 ,
		\g3006_reg/NET0131 ,
		\g3080_reg/NET0131 ,
		_w4616_
	);
	LUT2 #(
		.INIT('h8)
	) name3436 (
		\g3002_reg/NET0131 ,
		\g3013_reg/NET0131 ,
		_w4617_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3437 (
		\g3010_reg/NET0131 ,
		\g3024_reg/NET0131 ,
		_w4616_,
		_w4617_,
		_w4618_
	);
	LUT2 #(
		.INIT('h8)
	) name3438 (
		_w4615_,
		_w4618_,
		_w4619_
	);
	LUT3 #(
		.INIT('h0d)
	) name3439 (
		\g1024_reg/NET0131 ,
		\g1964_reg/NET0131 ,
		\g3229_pad ,
		_w4620_
	);
	LUT2 #(
		.INIT('h8)
	) name3440 (
		_w3714_,
		_w4620_,
		_w4621_
	);
	LUT4 #(
		.INIT('h3efe)
	) name3441 (
		\g3229_pad ,
		_w3690_,
		_w3699_,
		_w4621_,
		_w4622_
	);
	LUT3 #(
		.INIT('h8c)
	) name3442 (
		\g1956_reg/NET0131 ,
		\g3229_pad ,
		\g5657_pad ,
		_w4623_
	);
	LUT4 #(
		.INIT('hb000)
	) name3443 (
		_w3688_,
		_w3689_,
		_w3698_,
		_w4623_,
		_w4624_
	);
	LUT3 #(
		.INIT('hd0)
	) name3444 (
		\g1024_reg/NET0131 ,
		\g1964_reg/NET0131 ,
		\g3229_pad ,
		_w4625_
	);
	LUT2 #(
		.INIT('h8)
	) name3445 (
		_w3714_,
		_w4625_,
		_w4626_
	);
	LUT3 #(
		.INIT('h13)
	) name3446 (
		_w3718_,
		_w4624_,
		_w4626_,
		_w4627_
	);
	LUT2 #(
		.INIT('h8)
	) name3447 (
		_w4622_,
		_w4627_,
		_w4628_
	);
	LUT4 #(
		.INIT('h006a)
	) name3448 (
		\g1430_reg/NET0131 ,
		_w4278_,
		_w4279_,
		_w4283_,
		_w4629_
	);
	LUT2 #(
		.INIT('h8)
	) name3449 (
		\g1439_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		_w4630_
	);
	LUT3 #(
		.INIT('h15)
	) name3450 (
		\g1435_reg/NET0131 ,
		_w4278_,
		_w4630_,
		_w4631_
	);
	LUT3 #(
		.INIT('h07)
	) name3451 (
		_w4278_,
		_w4279_,
		_w4283_,
		_w4632_
	);
	LUT2 #(
		.INIT('h4)
	) name3452 (
		_w4631_,
		_w4632_,
		_w4633_
	);
	LUT3 #(
		.INIT('h06)
	) name3453 (
		\g1444_reg/NET0131 ,
		_w4278_,
		_w4283_,
		_w4634_
	);
	LUT4 #(
		.INIT('h8000)
	) name3454 (
		\g1088_reg/NET0131 ,
		\g1457_reg/NET0131 ,
		\g1462_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		_w4635_
	);
	LUT4 #(
		.INIT('h4055)
	) name3455 (
		\g1453_reg/NET0131 ,
		_w4071_,
		_w4072_,
		_w4635_,
		_w4636_
	);
	LUT2 #(
		.INIT('h8)
	) name3456 (
		\g1453_reg/NET0131 ,
		\g1457_reg/NET0131 ,
		_w4637_
	);
	LUT4 #(
		.INIT('h7000)
	) name3457 (
		_w4071_,
		_w4072_,
		_w4276_,
		_w4637_,
		_w4638_
	);
	LUT3 #(
		.INIT('h01)
	) name3458 (
		_w4283_,
		_w4636_,
		_w4638_,
		_w4639_
	);
	LUT3 #(
		.INIT('h70)
	) name3459 (
		_w4071_,
		_w4072_,
		_w4276_,
		_w4640_
	);
	LUT4 #(
		.INIT('h407f)
	) name3460 (
		_w3875_,
		_w4071_,
		_w4072_,
		_w4276_,
		_w4641_
	);
	LUT3 #(
		.INIT('h13)
	) name3461 (
		\g1088_reg/NET0131 ,
		\g1462_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		_w4642_
	);
	LUT3 #(
		.INIT('h01)
	) name3462 (
		\g1462_reg/NET0131 ,
		\g2896_reg/NET0131 ,
		\g2900_reg/NET0131 ,
		_w4643_
	);
	LUT3 #(
		.INIT('h13)
	) name3463 (
		_w4072_,
		_w4642_,
		_w4643_,
		_w4644_
	);
	LUT2 #(
		.INIT('h8)
	) name3464 (
		_w4641_,
		_w4644_,
		_w4645_
	);
	LUT3 #(
		.INIT('h51)
	) name3465 (
		\g3229_pad ,
		\g5657_pad ,
		\g585_reg/NET0131 ,
		_w4646_
	);
	LUT2 #(
		.INIT('h8)
	) name3466 (
		_w3789_,
		_w4646_,
		_w4647_
	);
	LUT4 #(
		.INIT('h3efe)
	) name3467 (
		\g3229_pad ,
		_w3765_,
		_w3768_,
		_w4647_,
		_w4648_
	);
	LUT3 #(
		.INIT('ha2)
	) name3468 (
		\g3229_pad ,
		\g5657_pad ,
		\g576_reg/NET0131 ,
		_w4649_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3469 (
		_w3764_,
		_w3766_,
		_w3767_,
		_w4649_,
		_w4650_
	);
	LUT3 #(
		.INIT('ha2)
	) name3470 (
		\g3229_pad ,
		\g5657_pad ,
		\g585_reg/NET0131 ,
		_w4651_
	);
	LUT2 #(
		.INIT('h8)
	) name3471 (
		_w3789_,
		_w4651_,
		_w4652_
	);
	LUT3 #(
		.INIT('h13)
	) name3472 (
		_w3769_,
		_w4650_,
		_w4652_,
		_w4653_
	);
	LUT2 #(
		.INIT('h8)
	) name3473 (
		_w4648_,
		_w4653_,
		_w4654_
	);
	LUT4 #(
		.INIT('h0800)
	) name3474 (
		\g1024_reg/NET0131 ,
		\g1326_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g1358_reg/NET0131 ,
		_w4655_
	);
	LUT4 #(
		.INIT('h0e0a)
	) name3475 (
		\g1352_reg/NET0131 ,
		_w3909_,
		_w3914_,
		_w4655_,
		_w4656_
	);
	LUT2 #(
		.INIT('h4)
	) name3476 (
		_w4606_,
		_w4656_,
		_w4657_
	);
	LUT2 #(
		.INIT('h8)
	) name3477 (
		\g2892_reg/NET0131 ,
		\g2903_reg/NET0131 ,
		_w4658_
	);
	LUT4 #(
		.INIT('h8000)
	) name3478 (
		\g2892_reg/NET0131 ,
		\g2903_reg/NET0131 ,
		\g2908_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		_w4659_
	);
	LUT2 #(
		.INIT('h4)
	) name3479 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		_w4660_
	);
	LUT4 #(
		.INIT('h0004)
	) name3480 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		\g2896_reg/NET0131 ,
		\g2900_reg/NET0131 ,
		_w4661_
	);
	LUT3 #(
		.INIT('h04)
	) name3481 (
		\g2917_reg/NET0131 ,
		\g2920_reg/NET0131 ,
		\g2924_reg/NET0131 ,
		_w4662_
	);
	LUT4 #(
		.INIT('h0020)
	) name3482 (
		\g2912_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		\g2920_reg/NET0131 ,
		\g2924_reg/NET0131 ,
		_w4663_
	);
	LUT4 #(
		.INIT('h1555)
	) name3483 (
		\g2814_reg/NET0131 ,
		_w4659_,
		_w4661_,
		_w4663_,
		_w4664_
	);
	LUT3 #(
		.INIT('h80)
	) name3484 (
		\g2912_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		\g2924_reg/NET0131 ,
		_w4665_
	);
	LUT4 #(
		.INIT('h8000)
	) name3485 (
		_w4071_,
		_w4659_,
		_w4660_,
		_w4665_,
		_w4666_
	);
	LUT4 #(
		.INIT('h8000)
	) name3486 (
		\g2912_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		\g2920_reg/NET0131 ,
		\g2924_reg/NET0131 ,
		_w4667_
	);
	LUT3 #(
		.INIT('h80)
	) name3487 (
		_w4659_,
		_w4661_,
		_w4667_,
		_w4668_
	);
	LUT4 #(
		.INIT('h00c8)
	) name3488 (
		\g2920_reg/NET0131 ,
		_w4664_,
		_w4666_,
		_w4668_,
		_w4669_
	);
	LUT3 #(
		.INIT('h0e)
	) name3489 (
		\g2813_reg/NET0131 ,
		_w3515_,
		_w3914_,
		_w4670_
	);
	LUT2 #(
		.INIT('h8)
	) name3490 (
		\g1024_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		_w4671_
	);
	LUT3 #(
		.INIT('h0e)
	) name3491 (
		\g1423_reg/NET0131 ,
		_w3522_,
		_w4671_,
		_w4672_
	);
	LUT2 #(
		.INIT('h8)
	) name3492 (
		\g1316_reg/NET0131 ,
		\g5657_pad ,
		_w4673_
	);
	LUT3 #(
		.INIT('h0e)
	) name3493 (
		\g1424_reg/NET0131 ,
		_w3567_,
		_w4673_,
		_w4674_
	);
	LUT3 #(
		.INIT('h0e)
	) name3494 (
		\g737_reg/NET0131 ,
		_w3612_,
		_w4671_,
		_w4675_
	);
	LUT3 #(
		.INIT('h0e)
	) name3495 (
		\g2119_reg/NET0131 ,
		_w3662_,
		_w3914_,
		_w4676_
	);
	LUT3 #(
		.INIT('h0e)
	) name3496 (
		\g738_reg/NET0131 ,
		_w3652_,
		_w4673_,
		_w4677_
	);
	LUT4 #(
		.INIT('h006a)
	) name3497 (
		\g1439_reg/NET0131 ,
		\g1444_reg/NET0131 ,
		_w4278_,
		_w4283_,
		_w4678_
	);
	LUT4 #(
		.INIT('h0302)
	) name3498 (
		\g1448_reg/NET0131 ,
		_w4278_,
		_w4283_,
		_w4638_,
		_w4679_
	);
	LUT4 #(
		.INIT('hc666)
	) name3499 (
		\g1088_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		_w4071_,
		_w4072_,
		_w4680_
	);
	LUT2 #(
		.INIT('h4)
	) name3500 (
		_w4283_,
		_w4680_,
		_w4681_
	);
	LUT3 #(
		.INIT('h2a)
	) name3501 (
		\g1457_reg/NET0131 ,
		_w4072_,
		_w4282_,
		_w4682_
	);
	LUT4 #(
		.INIT('h2000)
	) name3502 (
		\g1088_reg/NET0131 ,
		\g1457_reg/NET0131 ,
		\g1462_reg/NET0131 ,
		\g1466_reg/NET0131 ,
		_w4683_
	);
	LUT3 #(
		.INIT('h70)
	) name3503 (
		_w4071_,
		_w4072_,
		_w4683_,
		_w4684_
	);
	LUT3 #(
		.INIT('hf4)
	) name3504 (
		_w4640_,
		_w4682_,
		_w4684_,
		_w4685_
	);
	LUT3 #(
		.INIT('h70)
	) name3505 (
		\g1018_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		\g1346_reg/NET0131 ,
		_w4686_
	);
	LUT4 #(
		.INIT('h0080)
	) name3506 (
		\g1024_reg/NET0131 ,
		\g1319_reg/NET0131 ,
		\g1326_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w4687_
	);
	LUT4 #(
		.INIT('h7000)
	) name3507 (
		\g1018_reg/NET0131 ,
		\g1316_reg/NET0131 ,
		\g1332_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w4688_
	);
	LUT3 #(
		.INIT('h15)
	) name3508 (
		_w4686_,
		_w4687_,
		_w4688_,
		_w4689_
	);
	LUT2 #(
		.INIT('h1)
	) name3509 (
		_w3910_,
		_w4689_,
		_w4690_
	);
	LUT3 #(
		.INIT('h15)
	) name3510 (
		\g1358_reg/NET0131 ,
		_w3908_,
		_w3909_,
		_w4691_
	);
	LUT3 #(
		.INIT('h13)
	) name3511 (
		_w3909_,
		_w3914_,
		_w4655_,
		_w4692_
	);
	LUT2 #(
		.INIT('h4)
	) name3512 (
		_w4691_,
		_w4692_,
		_w4693_
	);
	LUT3 #(
		.INIT('h23)
	) name3513 (
		\g2650_reg/NET0131 ,
		\g3229_pad ,
		\g5657_pad ,
		_w4694_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3514 (
		_w3332_,
		_w3336_,
		_w3337_,
		_w4694_,
		_w4695_
	);
	LUT4 #(
		.INIT('h0007)
	) name3515 (
		\g3229_pad ,
		_w3339_,
		_w3368_,
		_w4695_,
		_w4696_
	);
	LUT3 #(
		.INIT('hab)
	) name3516 (
		_w4362_,
		_w4363_,
		_w4366_,
		_w4697_
	);
	LUT3 #(
		.INIT('hcd)
	) name3517 (
		_w4366_,
		_w4418_,
		_w4419_,
		_w4698_
	);
	LUT3 #(
		.INIT('hcd)
	) name3518 (
		_w4366_,
		_w4436_,
		_w4437_,
		_w4699_
	);
	LUT3 #(
		.INIT('hcd)
	) name3519 (
		_w4366_,
		_w4500_,
		_w4501_,
		_w4700_
	);
	LUT3 #(
		.INIT('hbf)
	) name3520 (
		_w4342_,
		_w4346_,
		_w4493_,
		_w4701_
	);
	LUT3 #(
		.INIT('h0d)
	) name3521 (
		\g1024_reg/NET0131 ,
		\g1961_reg/NET0131 ,
		\g3229_pad ,
		_w4702_
	);
	LUT2 #(
		.INIT('h8)
	) name3522 (
		_w3692_,
		_w4702_,
		_w4703_
	);
	LUT3 #(
		.INIT('hd0)
	) name3523 (
		\g1024_reg/NET0131 ,
		\g1961_reg/NET0131 ,
		\g3229_pad ,
		_w4704_
	);
	LUT2 #(
		.INIT('h8)
	) name3524 (
		_w3692_,
		_w4704_,
		_w4705_
	);
	LUT4 #(
		.INIT('h57df)
	) name3525 (
		_w3690_,
		_w3699_,
		_w4703_,
		_w4705_,
		_w4706_
	);
	LUT3 #(
		.INIT('hdf)
	) name3526 (
		_w4393_,
		_w4395_,
		_w4408_,
		_w4707_
	);
	LUT3 #(
		.INIT('h31)
	) name3527 (
		\g1024_reg/NET0131 ,
		\g3229_pad ,
		\g581_reg/NET0131 ,
		_w4708_
	);
	LUT2 #(
		.INIT('h8)
	) name3528 (
		_w3778_,
		_w4708_,
		_w4709_
	);
	LUT3 #(
		.INIT('hc4)
	) name3529 (
		\g1024_reg/NET0131 ,
		\g3229_pad ,
		\g581_reg/NET0131 ,
		_w4710_
	);
	LUT2 #(
		.INIT('h8)
	) name3530 (
		_w3778_,
		_w4710_,
		_w4711_
	);
	LUT4 #(
		.INIT('h37bf)
	) name3531 (
		_w3765_,
		_w3768_,
		_w4709_,
		_w4711_,
		_w4712_
	);
	LUT3 #(
		.INIT('h0d)
	) name3532 (
		\g1024_reg/NET0131 ,
		\g1264_reg/NET0131 ,
		\g3229_pad ,
		_w4713_
	);
	LUT4 #(
		.INIT('hb000)
	) name3533 (
		_w3226_,
		_w3227_,
		_w3230_,
		_w4713_,
		_w4714_
	);
	LUT3 #(
		.INIT('hd0)
	) name3534 (
		\g1018_reg/NET0131 ,
		\g1269_reg/NET0131 ,
		\g3229_pad ,
		_w4715_
	);
	LUT2 #(
		.INIT('h8)
	) name3535 (
		_w3238_,
		_w4715_,
		_w4716_
	);
	LUT4 #(
		.INIT('h135f)
	) name3536 (
		_w3239_,
		_w3293_,
		_w4714_,
		_w4716_,
		_w4717_
	);
	LUT3 #(
		.INIT('hdf)
	) name3537 (
		_w4467_,
		_w4469_,
		_w4484_,
		_w4718_
	);
	LUT3 #(
		.INIT('hd0)
	) name3538 (
		\g1018_reg/NET0131 ,
		\g2657_reg/NET0131 ,
		\g3229_pad ,
		_w4719_
	);
	LUT2 #(
		.INIT('h8)
	) name3539 (
		_w3337_,
		_w4719_,
		_w4720_
	);
	LUT3 #(
		.INIT('h0d)
	) name3540 (
		\g1018_reg/NET0131 ,
		\g2657_reg/NET0131 ,
		\g3229_pad ,
		_w4721_
	);
	LUT2 #(
		.INIT('h8)
	) name3541 (
		_w3337_,
		_w4721_,
		_w4722_
	);
	LUT4 #(
		.INIT('h5d7f)
	) name3542 (
		_w3330_,
		_w3333_,
		_w4720_,
		_w4722_,
		_w4723_
	);
	LUT3 #(
		.INIT('hdf)
	) name3543 (
		_w4521_,
		_w4523_,
		_w4553_,
		_w4724_
	);
	LUT4 #(
		.INIT('h5ccc)
	) name3544 (
		\g1326_reg/NET0131 ,
		\g1384_reg/NET0131 ,
		_w3520_,
		_w3521_,
		_w4725_
	);
	LUT3 #(
		.INIT('h5c)
	) name3545 (
		\g1326_reg/NET0131 ,
		\g1385_reg/NET0131 ,
		_w3567_,
		_w4726_
	);
	LUT3 #(
		.INIT('h0e)
	) name3546 (
		\g2811_reg/NET0131 ,
		_w3672_,
		_w4671_,
		_w4727_
	);
	LUT3 #(
		.INIT('h5c)
	) name3547 (
		\g1326_reg/NET0131 ,
		\g1386_reg/NET0131 ,
		_w3562_,
		_w4728_
	);
	LUT3 #(
		.INIT('h0e)
	) name3548 (
		\g2812_reg/NET0131 ,
		_w3475_,
		_w4673_,
		_w4729_
	);
	LUT3 #(
		.INIT('h5c)
	) name3549 (
		\g1319_reg/NET0131 ,
		\g1387_reg/NET0131 ,
		_w3522_,
		_w4730_
	);
	LUT3 #(
		.INIT('h5c)
	) name3550 (
		\g1319_reg/NET0131 ,
		\g1388_reg/NET0131 ,
		_w3567_,
		_w4731_
	);
	LUT3 #(
		.INIT('h5c)
	) name3551 (
		\g1319_reg/NET0131 ,
		\g1389_reg/NET0131 ,
		_w3562_,
		_w4732_
	);
	LUT3 #(
		.INIT('h5c)
	) name3552 (
		\g1339_reg/NET0131 ,
		\g1390_reg/NET0131 ,
		_w3522_,
		_w4733_
	);
	LUT3 #(
		.INIT('h5c)
	) name3553 (
		\g1339_reg/NET0131 ,
		\g1391_reg/NET0131 ,
		_w3567_,
		_w4734_
	);
	LUT3 #(
		.INIT('h5c)
	) name3554 (
		\g1339_reg/NET0131 ,
		\g1392_reg/NET0131 ,
		_w3562_,
		_w4735_
	);
	LUT3 #(
		.INIT('h5c)
	) name3555 (
		\g1332_reg/NET0131 ,
		\g1393_reg/NET0131 ,
		_w3522_,
		_w4736_
	);
	LUT3 #(
		.INIT('h5c)
	) name3556 (
		\g1332_reg/NET0131 ,
		\g1394_reg/NET0131 ,
		_w3567_,
		_w4737_
	);
	LUT3 #(
		.INIT('h5c)
	) name3557 (
		\g1332_reg/NET0131 ,
		\g1395_reg/NET0131 ,
		_w3562_,
		_w4738_
	);
	LUT3 #(
		.INIT('h5c)
	) name3558 (
		\g1346_reg/NET0131 ,
		\g1396_reg/NET0131 ,
		_w3522_,
		_w4739_
	);
	LUT3 #(
		.INIT('h5c)
	) name3559 (
		\g1346_reg/NET0131 ,
		\g1397_reg/NET0131 ,
		_w3567_,
		_w4740_
	);
	LUT3 #(
		.INIT('h5c)
	) name3560 (
		\g1346_reg/NET0131 ,
		\g1398_reg/NET0131 ,
		_w3562_,
		_w4741_
	);
	LUT3 #(
		.INIT('h5c)
	) name3561 (
		\g1358_reg/NET0131 ,
		\g1399_reg/NET0131 ,
		_w3522_,
		_w4742_
	);
	LUT3 #(
		.INIT('h5c)
	) name3562 (
		\g1358_reg/NET0131 ,
		\g1400_reg/NET0131 ,
		_w3567_,
		_w4743_
	);
	LUT3 #(
		.INIT('h5c)
	) name3563 (
		\g1358_reg/NET0131 ,
		\g1401_reg/NET0131 ,
		_w3562_,
		_w4744_
	);
	LUT3 #(
		.INIT('h5c)
	) name3564 (
		\g1352_reg/NET0131 ,
		\g1402_reg/NET0131 ,
		_w3522_,
		_w4745_
	);
	LUT3 #(
		.INIT('h5c)
	) name3565 (
		\g1352_reg/NET0131 ,
		\g1403_reg/NET0131 ,
		_w3567_,
		_w4746_
	);
	LUT3 #(
		.INIT('h5c)
	) name3566 (
		\g1352_reg/NET0131 ,
		\g1404_reg/NET0131 ,
		_w3562_,
		_w4747_
	);
	LUT3 #(
		.INIT('h5c)
	) name3567 (
		\g1365_reg/NET0131 ,
		\g1405_reg/NET0131 ,
		_w3522_,
		_w4748_
	);
	LUT3 #(
		.INIT('h5c)
	) name3568 (
		\g1365_reg/NET0131 ,
		\g1406_reg/NET0131 ,
		_w3567_,
		_w4749_
	);
	LUT3 #(
		.INIT('h5c)
	) name3569 (
		\g1365_reg/NET0131 ,
		\g1407_reg/NET0131 ,
		_w3562_,
		_w4750_
	);
	LUT3 #(
		.INIT('h5c)
	) name3570 (
		\g1372_reg/NET0131 ,
		\g1408_reg/NET0131 ,
		_w3522_,
		_w4751_
	);
	LUT3 #(
		.INIT('h5c)
	) name3571 (
		\g1372_reg/NET0131 ,
		\g1409_reg/NET0131 ,
		_w3567_,
		_w4752_
	);
	LUT3 #(
		.INIT('h5c)
	) name3572 (
		\g1372_reg/NET0131 ,
		\g1410_reg/NET0131 ,
		_w3562_,
		_w4753_
	);
	LUT3 #(
		.INIT('h5c)
	) name3573 (
		\g1378_reg/NET0131 ,
		\g1411_reg/NET0131 ,
		_w3522_,
		_w4754_
	);
	LUT3 #(
		.INIT('h5c)
	) name3574 (
		\g1378_reg/NET0131 ,
		\g1412_reg/NET0131 ,
		_w3567_,
		_w4755_
	);
	LUT3 #(
		.INIT('h5c)
	) name3575 (
		\g1378_reg/NET0131 ,
		\g1413_reg/NET0131 ,
		_w3562_,
		_w4756_
	);
	LUT4 #(
		.INIT('h7f08)
	) name3576 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g2200_reg/NET0131 ,
		\g2232_reg/NET0131 ,
		_w4757_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3577 (
		\g1088_reg/NET0131 ,
		\g1471_reg/NET0131 ,
		\g1511_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4758_
	);
	LUT4 #(
		.INIT('h5ccc)
	) name3578 (
		\g1471_reg/NET0131 ,
		\g1512_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w4759_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3579 (
		\g1092_reg/NET0131 ,
		\g1471_reg/NET0131 ,
		\g1513_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4760_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3580 (
		\g1088_reg/NET0131 ,
		\g1491_reg/NET0131 ,
		\g1529_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4761_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3581 (
		\g1092_reg/NET0131 ,
		\g1491_reg/NET0131 ,
		\g1531_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4762_
	);
	LUT4 #(
		.INIT('h5ccc)
	) name3582 (
		\g1491_reg/NET0131 ,
		\g1530_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w4763_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3583 (
		\g1088_reg/NET0131 ,
		\g1496_reg/NET0131 ,
		\g1532_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4764_
	);
	LUT4 #(
		.INIT('h5ccc)
	) name3584 (
		\g1496_reg/NET0131 ,
		\g1533_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w4765_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3585 (
		\g1092_reg/NET0131 ,
		\g1496_reg/NET0131 ,
		\g1534_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4766_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3586 (
		\g1088_reg/NET0131 ,
		\g1501_reg/NET0131 ,
		\g1535_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4767_
	);
	LUT4 #(
		.INIT('h5ccc)
	) name3587 (
		\g1501_reg/NET0131 ,
		\g1536_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w4768_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3588 (
		\g1092_reg/NET0131 ,
		\g1501_reg/NET0131 ,
		\g1537_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4769_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3589 (
		\g1088_reg/NET0131 ,
		\g1506_reg/NET0131 ,
		\g1538_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4770_
	);
	LUT4 #(
		.INIT('h5ccc)
	) name3590 (
		\g1506_reg/NET0131 ,
		\g1539_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w4771_
	);
	LUT3 #(
		.INIT('h5c)
	) name3591 (
		\g1326_reg/NET0131 ,
		\g698_reg/NET0131 ,
		_w3612_,
		_w4772_
	);
	LUT3 #(
		.INIT('h5c)
	) name3592 (
		\g1326_reg/NET0131 ,
		\g699_reg/NET0131 ,
		_w3652_,
		_w4773_
	);
	LUT3 #(
		.INIT('h5c)
	) name3593 (
		\g1326_reg/NET0131 ,
		\g700_reg/NET0131 ,
		_w3657_,
		_w4774_
	);
	LUT3 #(
		.INIT('h5c)
	) name3594 (
		\g1319_reg/NET0131 ,
		\g701_reg/NET0131 ,
		_w3612_,
		_w4775_
	);
	LUT3 #(
		.INIT('h5c)
	) name3595 (
		\g1319_reg/NET0131 ,
		\g702_reg/NET0131 ,
		_w3652_,
		_w4776_
	);
	LUT3 #(
		.INIT('h5c)
	) name3596 (
		\g1319_reg/NET0131 ,
		\g703_reg/NET0131 ,
		_w3657_,
		_w4777_
	);
	LUT3 #(
		.INIT('h5c)
	) name3597 (
		\g1339_reg/NET0131 ,
		\g704_reg/NET0131 ,
		_w3612_,
		_w4778_
	);
	LUT3 #(
		.INIT('h5c)
	) name3598 (
		\g1339_reg/NET0131 ,
		\g705_reg/NET0131 ,
		_w3652_,
		_w4779_
	);
	LUT3 #(
		.INIT('h5c)
	) name3599 (
		\g1339_reg/NET0131 ,
		\g706_reg/NET0131 ,
		_w3657_,
		_w4780_
	);
	LUT3 #(
		.INIT('h5c)
	) name3600 (
		\g1332_reg/NET0131 ,
		\g707_reg/NET0131 ,
		_w3612_,
		_w4781_
	);
	LUT3 #(
		.INIT('h5c)
	) name3601 (
		\g1332_reg/NET0131 ,
		\g708_reg/NET0131 ,
		_w3652_,
		_w4782_
	);
	LUT3 #(
		.INIT('h5c)
	) name3602 (
		\g1332_reg/NET0131 ,
		\g709_reg/NET0131 ,
		_w3657_,
		_w4783_
	);
	LUT3 #(
		.INIT('h5c)
	) name3603 (
		\g1346_reg/NET0131 ,
		\g710_reg/NET0131 ,
		_w3612_,
		_w4784_
	);
	LUT3 #(
		.INIT('h5c)
	) name3604 (
		\g1346_reg/NET0131 ,
		\g711_reg/NET0131 ,
		_w3652_,
		_w4785_
	);
	LUT3 #(
		.INIT('h5c)
	) name3605 (
		\g1346_reg/NET0131 ,
		\g712_reg/NET0131 ,
		_w3657_,
		_w4786_
	);
	LUT3 #(
		.INIT('h5c)
	) name3606 (
		\g1358_reg/NET0131 ,
		\g713_reg/NET0131 ,
		_w3612_,
		_w4787_
	);
	LUT3 #(
		.INIT('h5c)
	) name3607 (
		\g1358_reg/NET0131 ,
		\g714_reg/NET0131 ,
		_w3652_,
		_w4788_
	);
	LUT3 #(
		.INIT('h5c)
	) name3608 (
		\g1358_reg/NET0131 ,
		\g715_reg/NET0131 ,
		_w3657_,
		_w4789_
	);
	LUT3 #(
		.INIT('h5c)
	) name3609 (
		\g1352_reg/NET0131 ,
		\g716_reg/NET0131 ,
		_w3612_,
		_w4790_
	);
	LUT3 #(
		.INIT('h5c)
	) name3610 (
		\g1352_reg/NET0131 ,
		\g717_reg/NET0131 ,
		_w3652_,
		_w4791_
	);
	LUT3 #(
		.INIT('h5c)
	) name3611 (
		\g1352_reg/NET0131 ,
		\g718_reg/NET0131 ,
		_w3657_,
		_w4792_
	);
	LUT3 #(
		.INIT('h5c)
	) name3612 (
		\g1365_reg/NET0131 ,
		\g719_reg/NET0131 ,
		_w3612_,
		_w4793_
	);
	LUT3 #(
		.INIT('h5c)
	) name3613 (
		\g1365_reg/NET0131 ,
		\g720_reg/NET0131 ,
		_w3652_,
		_w4794_
	);
	LUT3 #(
		.INIT('h5c)
	) name3614 (
		\g1365_reg/NET0131 ,
		\g721_reg/NET0131 ,
		_w3657_,
		_w4795_
	);
	LUT3 #(
		.INIT('h5c)
	) name3615 (
		\g1372_reg/NET0131 ,
		\g722_reg/NET0131 ,
		_w3612_,
		_w4796_
	);
	LUT3 #(
		.INIT('h5c)
	) name3616 (
		\g1372_reg/NET0131 ,
		\g723_reg/NET0131 ,
		_w3652_,
		_w4797_
	);
	LUT3 #(
		.INIT('h5c)
	) name3617 (
		\g1372_reg/NET0131 ,
		\g724_reg/NET0131 ,
		_w3657_,
		_w4798_
	);
	LUT3 #(
		.INIT('h5c)
	) name3618 (
		\g1378_reg/NET0131 ,
		\g725_reg/NET0131 ,
		_w3612_,
		_w4799_
	);
	LUT3 #(
		.INIT('h5c)
	) name3619 (
		\g1378_reg/NET0131 ,
		\g726_reg/NET0131 ,
		_w3652_,
		_w4800_
	);
	LUT3 #(
		.INIT('h5c)
	) name3620 (
		\g1378_reg/NET0131 ,
		\g727_reg/NET0131 ,
		_w3657_,
		_w4801_
	);
	LUT3 #(
		.INIT('h0e)
	) name3621 (
		\g2118_reg/NET0131 ,
		_w3667_,
		_w4673_,
		_w4802_
	);
	LUT4 #(
		.INIT('h7f08)
	) name3622 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g2195_reg/NET0131 ,
		\g2229_reg/NET0131 ,
		_w4803_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3623 (
		\g1092_reg/NET0131 ,
		\g1506_reg/NET0131 ,
		\g1540_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4804_
	);
	LUT3 #(
		.INIT('h0e)
	) name3624 (
		\g2117_reg/NET0131 ,
		_w3572_,
		_w4671_,
		_w4805_
	);
	LUT2 #(
		.INIT('h2)
	) name3625 (
		\g1846_reg/NET0131 ,
		\g7961_pad ,
		_w4806_
	);
	LUT2 #(
		.INIT('h1)
	) name3626 (
		\g1846_reg/NET0131 ,
		\g7961_pad ,
		_w4807_
	);
	LUT3 #(
		.INIT('h04)
	) name3627 (
		_w2127_,
		_w2128_,
		_w4807_,
		_w4808_
	);
	LUT3 #(
		.INIT('hec)
	) name3628 (
		_w2143_,
		_w4806_,
		_w4808_,
		_w4809_
	);
	LUT2 #(
		.INIT('h4)
	) name3629 (
		\g1092_reg/NET0131 ,
		\g1849_reg/NET0131 ,
		_w4810_
	);
	LUT2 #(
		.INIT('h1)
	) name3630 (
		\g1092_reg/NET0131 ,
		\g1849_reg/NET0131 ,
		_w4811_
	);
	LUT3 #(
		.INIT('h04)
	) name3631 (
		_w2127_,
		_w2128_,
		_w4811_,
		_w4812_
	);
	LUT3 #(
		.INIT('hec)
	) name3632 (
		_w2143_,
		_w4810_,
		_w4812_,
		_w4813_
	);
	LUT2 #(
		.INIT('h4)
	) name3633 (
		\g1088_reg/NET0131 ,
		\g1852_reg/NET0131 ,
		_w4814_
	);
	LUT2 #(
		.INIT('h1)
	) name3634 (
		\g1088_reg/NET0131 ,
		\g1852_reg/NET0131 ,
		_w4815_
	);
	LUT3 #(
		.INIT('h04)
	) name3635 (
		_w2127_,
		_w2128_,
		_w4815_,
		_w4816_
	);
	LUT3 #(
		.INIT('hec)
	) name3636 (
		_w2143_,
		_w4814_,
		_w4816_,
		_w4817_
	);
	LUT2 #(
		.INIT('h2)
	) name3637 (
		\g465_reg/NET0131 ,
		\g7961_pad ,
		_w4818_
	);
	LUT2 #(
		.INIT('h1)
	) name3638 (
		\g465_reg/NET0131 ,
		\g7961_pad ,
		_w4819_
	);
	LUT3 #(
		.INIT('h04)
	) name3639 (
		_w1695_,
		_w1696_,
		_w4819_,
		_w4820_
	);
	LUT3 #(
		.INIT('hec)
	) name3640 (
		_w1821_,
		_w4818_,
		_w4820_,
		_w4821_
	);
	LUT2 #(
		.INIT('h4)
	) name3641 (
		\g1092_reg/NET0131 ,
		\g468_reg/NET0131 ,
		_w4822_
	);
	LUT2 #(
		.INIT('h1)
	) name3642 (
		\g1092_reg/NET0131 ,
		\g468_reg/NET0131 ,
		_w4823_
	);
	LUT3 #(
		.INIT('h04)
	) name3643 (
		_w1695_,
		_w1696_,
		_w4823_,
		_w4824_
	);
	LUT3 #(
		.INIT('hec)
	) name3644 (
		_w1821_,
		_w4822_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h4)
	) name3645 (
		\g1088_reg/NET0131 ,
		\g471_reg/NET0131 ,
		_w4826_
	);
	LUT2 #(
		.INIT('h1)
	) name3646 (
		\g1088_reg/NET0131 ,
		\g471_reg/NET0131 ,
		_w4827_
	);
	LUT3 #(
		.INIT('h04)
	) name3647 (
		_w1695_,
		_w1696_,
		_w4827_,
		_w4828_
	);
	LUT3 #(
		.INIT('hec)
	) name3648 (
		_w1821_,
		_w4826_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h2)
	) name3649 (
		\g2540_reg/NET0131 ,
		\g7961_pad ,
		_w4830_
	);
	LUT4 #(
		.INIT('hddd0)
	) name3650 (
		\g1092_reg/NET0131 ,
		\g2394_reg/NET0131 ,
		\g2540_reg/NET0131 ,
		\g7961_pad ,
		_w4831_
	);
	LUT4 #(
		.INIT('h2000)
	) name3651 (
		_w1252_,
		_w1362_,
		_w1363_,
		_w4831_,
		_w4832_
	);
	LUT3 #(
		.INIT('hec)
	) name3652 (
		_w1368_,
		_w4830_,
		_w4832_,
		_w4833_
	);
	LUT2 #(
		.INIT('h4)
	) name3653 (
		\g1092_reg/NET0131 ,
		\g2543_reg/NET0131 ,
		_w4834_
	);
	LUT3 #(
		.INIT('hd8)
	) name3654 (
		\g1092_reg/NET0131 ,
		\g2394_reg/NET0131 ,
		\g2543_reg/NET0131 ,
		_w4835_
	);
	LUT4 #(
		.INIT('h2000)
	) name3655 (
		_w1252_,
		_w1362_,
		_w1363_,
		_w4835_,
		_w4836_
	);
	LUT3 #(
		.INIT('hec)
	) name3656 (
		_w1368_,
		_w4834_,
		_w4836_,
		_w4837_
	);
	LUT2 #(
		.INIT('h4)
	) name3657 (
		\g1088_reg/NET0131 ,
		\g2546_reg/NET0131 ,
		_w4838_
	);
	LUT4 #(
		.INIT('hf3a2)
	) name3658 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g2394_reg/NET0131 ,
		\g2546_reg/NET0131 ,
		_w4839_
	);
	LUT4 #(
		.INIT('h2000)
	) name3659 (
		_w1252_,
		_w1362_,
		_w1363_,
		_w4839_,
		_w4840_
	);
	LUT3 #(
		.INIT('hec)
	) name3660 (
		_w1368_,
		_w4838_,
		_w4840_,
		_w4841_
	);
	LUT3 #(
		.INIT('h70)
	) name3661 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g847_reg/NET0131 ,
		_w4842_
	);
	LUT3 #(
		.INIT('h80)
	) name3662 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g862_reg/NET0131 ,
		_w4843_
	);
	LUT3 #(
		.INIT('hec)
	) name3663 (
		_w1899_,
		_w4842_,
		_w4843_,
		_w4844_
	);
	LUT3 #(
		.INIT('h70)
	) name3664 (
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		\g848_reg/NET0131 ,
		_w4845_
	);
	LUT4 #(
		.INIT('hc040)
	) name3665 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		\g862_reg/NET0131 ,
		_w4846_
	);
	LUT3 #(
		.INIT('hec)
	) name3666 (
		_w1899_,
		_w4845_,
		_w4846_,
		_w4847_
	);
	LUT3 #(
		.INIT('h70)
	) name3667 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g849_reg/NET0131 ,
		_w4848_
	);
	LUT4 #(
		.INIT('hc040)
	) name3668 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g862_reg/NET0131 ,
		_w4849_
	);
	LUT3 #(
		.INIT('hec)
	) name3669 (
		_w1899_,
		_w4848_,
		_w4849_,
		_w4850_
	);
	LUT3 #(
		.INIT('h70)
	) name3670 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g850_reg/NET0131 ,
		_w4851_
	);
	LUT3 #(
		.INIT('h80)
	) name3671 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g859_reg/NET0131 ,
		_w4852_
	);
	LUT3 #(
		.INIT('hec)
	) name3672 (
		_w1875_,
		_w4851_,
		_w4852_,
		_w4853_
	);
	LUT3 #(
		.INIT('h70)
	) name3673 (
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		\g851_reg/NET0131 ,
		_w4854_
	);
	LUT4 #(
		.INIT('hc040)
	) name3674 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		\g859_reg/NET0131 ,
		_w4855_
	);
	LUT3 #(
		.INIT('hec)
	) name3675 (
		_w1875_,
		_w4854_,
		_w4855_,
		_w4856_
	);
	LUT3 #(
		.INIT('h70)
	) name3676 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g852_reg/NET0131 ,
		_w4857_
	);
	LUT4 #(
		.INIT('hc040)
	) name3677 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g859_reg/NET0131 ,
		_w4858_
	);
	LUT3 #(
		.INIT('hec)
	) name3678 (
		_w1875_,
		_w4857_,
		_w4858_,
		_w4859_
	);
	LUT3 #(
		.INIT('h70)
	) name3679 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g159_reg/NET0131 ,
		_w4860_
	);
	LUT3 #(
		.INIT('h80)
	) name3680 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g174_reg/NET0131 ,
		_w4861_
	);
	LUT3 #(
		.INIT('hec)
	) name3681 (
		_w1739_,
		_w4860_,
		_w4861_,
		_w4862_
	);
	LUT3 #(
		.INIT('h4c)
	) name3682 (
		\g1563_reg/NET0131 ,
		\g160_reg/NET0131 ,
		\g7961_pad ,
		_w4863_
	);
	LUT4 #(
		.INIT('hc400)
	) name3683 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g174_reg/NET0131 ,
		\g7961_pad ,
		_w4864_
	);
	LUT3 #(
		.INIT('hec)
	) name3684 (
		_w1739_,
		_w4863_,
		_w4864_,
		_w4865_
	);
	LUT3 #(
		.INIT('h70)
	) name3685 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g161_reg/NET0131 ,
		_w4866_
	);
	LUT4 #(
		.INIT('hc040)
	) name3686 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g174_reg/NET0131 ,
		_w4867_
	);
	LUT3 #(
		.INIT('hec)
	) name3687 (
		_w1739_,
		_w4866_,
		_w4867_,
		_w4868_
	);
	LUT3 #(
		.INIT('h70)
	) name3688 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g162_reg/NET0131 ,
		_w4869_
	);
	LUT3 #(
		.INIT('h80)
	) name3689 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g171_reg/NET0131 ,
		_w4870_
	);
	LUT3 #(
		.INIT('hec)
	) name3690 (
		_w1729_,
		_w4869_,
		_w4870_,
		_w4871_
	);
	LUT3 #(
		.INIT('h4c)
	) name3691 (
		\g1563_reg/NET0131 ,
		\g163_reg/NET0131 ,
		\g7961_pad ,
		_w4872_
	);
	LUT4 #(
		.INIT('hc400)
	) name3692 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g171_reg/NET0131 ,
		\g7961_pad ,
		_w4873_
	);
	LUT3 #(
		.INIT('hec)
	) name3693 (
		_w1729_,
		_w4872_,
		_w4873_,
		_w4874_
	);
	LUT3 #(
		.INIT('h70)
	) name3694 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g164_reg/NET0131 ,
		_w4875_
	);
	LUT4 #(
		.INIT('hc040)
	) name3695 (
		\g1088_reg/NET0131 ,
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g171_reg/NET0131 ,
		_w4876_
	);
	LUT3 #(
		.INIT('hec)
	) name3696 (
		_w1729_,
		_w4875_,
		_w4876_,
		_w4877_
	);
	LUT4 #(
		.INIT('h7f08)
	) name3697 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g805_reg/NET0131 ,
		\g838_reg/NET0131 ,
		_w4878_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3698 (
		\g1088_reg/NET0131 ,
		\g117_reg/NET0131 ,
		\g150_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4879_
	);
	LUT4 #(
		.INIT('h5ccc)
	) name3699 (
		\g117_reg/NET0131 ,
		\g151_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		_w4880_
	);
	LUT4 #(
		.INIT('h72f0)
	) name3700 (
		\g1092_reg/NET0131 ,
		\g117_reg/NET0131 ,
		\g152_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		_w4881_
	);
	LUT4 #(
		.INIT('h7f08)
	) name3701 (
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		\g805_reg/NET0131 ,
		\g839_reg/NET0131 ,
		_w4882_
	);
	LUT4 #(
		.INIT('h7f08)
	) name3702 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g805_reg/NET0131 ,
		\g840_reg/NET0131 ,
		_w4883_
	);
	LUT4 #(
		.INIT('h7f08)
	) name3703 (
		\g1088_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g813_reg/NET0131 ,
		\g844_reg/NET0131 ,
		_w4884_
	);
	LUT4 #(
		.INIT('h7f08)
	) name3704 (
		\g1563_reg/NET0131 ,
		\g7961_pad ,
		\g813_reg/NET0131 ,
		\g845_reg/NET0131 ,
		_w4885_
	);
	LUT4 #(
		.INIT('h7f08)
	) name3705 (
		\g1092_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g813_reg/NET0131 ,
		\g846_reg/NET0131 ,
		_w4886_
	);
	LUT4 #(
		.INIT('h7f20)
	) name3706 (
		\g1088_reg/NET0131 ,
		\g125_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g156_reg/NET0131 ,
		_w4887_
	);
	LUT4 #(
		.INIT('h74f0)
	) name3707 (
		\g125_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g157_reg/NET0131 ,
		\g7961_pad ,
		_w4888_
	);
	LUT4 #(
		.INIT('h7f20)
	) name3708 (
		\g1092_reg/NET0131 ,
		\g125_reg/NET0131 ,
		\g1563_reg/NET0131 ,
		\g158_reg/NET0131 ,
		_w4889_
	);
	LUT3 #(
		.INIT('h4c)
	) name3709 (
		\g1024_reg/NET0131 ,
		\g1196_reg/NET0131 ,
		\g2000_reg/NET0131 ,
		_w4890_
	);
	LUT4 #(
		.INIT('h0800)
	) name3710 (
		_w1577_,
		_w4359_,
		_w4360_,
		_w4890_,
		_w4891_
	);
	LUT3 #(
		.INIT('h4c)
	) name3711 (
		\g1018_reg/NET0131 ,
		\g1196_reg/NET0131 ,
		\g617_reg/NET0131 ,
		_w4892_
	);
	LUT4 #(
		.INIT('h0800)
	) name3712 (
		_w2864_,
		_w4415_,
		_w4416_,
		_w4892_,
		_w4893_
	);
	LUT3 #(
		.INIT('h2a)
	) name3713 (
		\g1196_reg/NET0131 ,
		\g1300_reg/NET0131 ,
		\g5657_pad ,
		_w4894_
	);
	LUT4 #(
		.INIT('h0800)
	) name3714 (
		_w2207_,
		_w4433_,
		_w4434_,
		_w4894_,
		_w4895_
	);
	LUT3 #(
		.INIT('h2a)
	) name3715 (
		\g1196_reg/NET0131 ,
		\g2688_reg/NET0131 ,
		\g5657_pad ,
		_w4896_
	);
	LUT4 #(
		.INIT('h0800)
	) name3716 (
		_w1418_,
		_w4497_,
		_w4498_,
		_w4896_,
		_w4897_
	);
	LUT4 #(
		.INIT('h060a)
	) name3717 (
		\g1332_reg/NET0131 ,
		\g1339_reg/NET0131 ,
		_w3914_,
		_w4687_,
		_w4898_
	);
	LUT3 #(
		.INIT('h6a)
	) name3718 (
		\g3010_reg/NET0131 ,
		_w4616_,
		_w4617_,
		_w4899_
	);
	LUT2 #(
		.INIT('h8)
	) name3719 (
		_w4615_,
		_w4899_,
		_w4900_
	);
	LUT3 #(
		.INIT('h32)
	) name3720 (
		_w4393_,
		_w4394_,
		_w4409_,
		_w4901_
	);
	LUT3 #(
		.INIT('h23)
	) name3721 (
		\g1956_reg/NET0131 ,
		\g3229_pad ,
		\g5657_pad ,
		_w4902_
	);
	LUT2 #(
		.INIT('h8)
	) name3722 (
		_w3698_,
		_w4902_,
		_w4903_
	);
	LUT3 #(
		.INIT('h8a)
	) name3723 (
		\g3229_pad ,
		_w3697_,
		_w3698_,
		_w4904_
	);
	LUT4 #(
		.INIT('h888b)
	) name3724 (
		_w3690_,
		_w3693_,
		_w4903_,
		_w4904_,
		_w4905_
	);
	LUT3 #(
		.INIT('h23)
	) name3725 (
		\g1262_reg/NET0131 ,
		\g3229_pad ,
		\g5657_pad ,
		_w4906_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3726 (
		_w3227_,
		_w3237_,
		_w3238_,
		_w4906_,
		_w4907_
	);
	LUT4 #(
		.INIT('h0013)
	) name3727 (
		\g3229_pad ,
		_w3279_,
		_w3288_,
		_w4907_,
		_w4908_
	);
	LUT3 #(
		.INIT('h32)
	) name3728 (
		_w4467_,
		_w4468_,
		_w4485_,
		_w4909_
	);
	LUT3 #(
		.INIT('h51)
	) name3729 (
		\g3229_pad ,
		\g5657_pad ,
		\g576_reg/NET0131 ,
		_w4910_
	);
	LUT4 #(
		.INIT('h8a00)
	) name3730 (
		_w3764_,
		_w3777_,
		_w3778_,
		_w4910_,
		_w4911_
	);
	LUT4 #(
		.INIT('h0007)
	) name3731 (
		\g3229_pad ,
		_w3780_,
		_w3805_,
		_w4911_,
		_w4912_
	);
	LUT3 #(
		.INIT('h32)
	) name3732 (
		_w4521_,
		_w4522_,
		_w4554_,
		_w4913_
	);
	LUT3 #(
		.INIT('h12)
	) name3733 (
		\g1339_reg/NET0131 ,
		_w3914_,
		_w4687_,
		_w4914_
	);
	LUT3 #(
		.INIT('h0e)
	) name3734 (
		_w4345_,
		_w4493_,
		_w4494_,
		_w4915_
	);
	LUT3 #(
		.INIT('h15)
	) name3735 (
		\g2814_reg/NET0131 ,
		_w4659_,
		_w4661_,
		_w4916_
	);
	LUT4 #(
		.INIT('h8000)
	) name3736 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		\g2896_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		_w4917_
	);
	LUT4 #(
		.INIT('h6ccc)
	) name3737 (
		\g2900_reg/NET0131 ,
		\g2908_reg/NET0131 ,
		_w4658_,
		_w4917_,
		_w4918_
	);
	LUT2 #(
		.INIT('h8)
	) name3738 (
		_w4916_,
		_w4918_,
		_w4919_
	);
	LUT3 #(
		.INIT('h5c)
	) name3739 (
		\g1326_reg/NET0131 ,
		\g2080_reg/NET0131 ,
		_w3662_,
		_w4920_
	);
	LUT3 #(
		.INIT('h5c)
	) name3740 (
		\g1372_reg/NET0131 ,
		\g2103_reg/NET0131 ,
		_w3667_,
		_w4921_
	);
	LUT3 #(
		.INIT('h5c)
	) name3741 (
		\g1346_reg/NET0131 ,
		\g2092_reg/NET0131 ,
		_w3662_,
		_w4922_
	);
	LUT3 #(
		.INIT('h5c)
	) name3742 (
		\g1326_reg/NET0131 ,
		\g2078_reg/NET0131 ,
		_w3572_,
		_w4923_
	);
	LUT3 #(
		.INIT('h5c)
	) name3743 (
		\g1326_reg/NET0131 ,
		\g2079_reg/NET0131 ,
		_w3667_,
		_w4924_
	);
	LUT3 #(
		.INIT('h5c)
	) name3744 (
		\g1319_reg/NET0131 ,
		\g2081_reg/NET0131 ,
		_w3572_,
		_w4925_
	);
	LUT3 #(
		.INIT('h5c)
	) name3745 (
		\g1319_reg/NET0131 ,
		\g2082_reg/NET0131 ,
		_w3667_,
		_w4926_
	);
	LUT3 #(
		.INIT('h5c)
	) name3746 (
		\g1319_reg/NET0131 ,
		\g2083_reg/NET0131 ,
		_w3662_,
		_w4927_
	);
	LUT3 #(
		.INIT('h5c)
	) name3747 (
		\g1339_reg/NET0131 ,
		\g2084_reg/NET0131 ,
		_w3572_,
		_w4928_
	);
	LUT3 #(
		.INIT('h5c)
	) name3748 (
		\g1339_reg/NET0131 ,
		\g2085_reg/NET0131 ,
		_w3667_,
		_w4929_
	);
	LUT3 #(
		.INIT('h5c)
	) name3749 (
		\g1332_reg/NET0131 ,
		\g2087_reg/NET0131 ,
		_w3572_,
		_w4930_
	);
	LUT3 #(
		.INIT('h5c)
	) name3750 (
		\g1332_reg/NET0131 ,
		\g2089_reg/NET0131 ,
		_w3662_,
		_w4931_
	);
	LUT3 #(
		.INIT('h5c)
	) name3751 (
		\g1358_reg/NET0131 ,
		\g2093_reg/NET0131 ,
		_w3572_,
		_w4932_
	);
	LUT3 #(
		.INIT('h5c)
	) name3752 (
		\g1358_reg/NET0131 ,
		\g2095_reg/NET0131 ,
		_w3662_,
		_w4933_
	);
	LUT3 #(
		.INIT('h5c)
	) name3753 (
		\g1352_reg/NET0131 ,
		\g2097_reg/NET0131 ,
		_w3667_,
		_w4934_
	);
	LUT3 #(
		.INIT('h5c)
	) name3754 (
		\g1365_reg/NET0131 ,
		\g2099_reg/NET0131 ,
		_w3572_,
		_w4935_
	);
	LUT3 #(
		.INIT('h5c)
	) name3755 (
		\g1365_reg/NET0131 ,
		\g2100_reg/NET0131 ,
		_w3667_,
		_w4936_
	);
	LUT3 #(
		.INIT('h5c)
	) name3756 (
		\g1365_reg/NET0131 ,
		\g2101_reg/NET0131 ,
		_w3662_,
		_w4937_
	);
	LUT3 #(
		.INIT('h5c)
	) name3757 (
		\g1372_reg/NET0131 ,
		\g2102_reg/NET0131 ,
		_w3572_,
		_w4938_
	);
	LUT3 #(
		.INIT('h5c)
	) name3758 (
		\g1372_reg/NET0131 ,
		\g2104_reg/NET0131 ,
		_w3662_,
		_w4939_
	);
	LUT3 #(
		.INIT('h5c)
	) name3759 (
		\g1378_reg/NET0131 ,
		\g2106_reg/NET0131 ,
		_w3667_,
		_w4940_
	);
	LUT3 #(
		.INIT('h5c)
	) name3760 (
		\g1378_reg/NET0131 ,
		\g2107_reg/NET0131 ,
		_w3662_,
		_w4941_
	);
	LUT3 #(
		.INIT('h5c)
	) name3761 (
		\g1346_reg/NET0131 ,
		\g2091_reg/NET0131 ,
		_w3667_,
		_w4942_
	);
	LUT3 #(
		.INIT('h5c)
	) name3762 (
		\g1346_reg/NET0131 ,
		\g2090_reg/NET0131 ,
		_w3572_,
		_w4943_
	);
	LUT3 #(
		.INIT('h5c)
	) name3763 (
		\g1339_reg/NET0131 ,
		\g2086_reg/NET0131 ,
		_w3662_,
		_w4944_
	);
	LUT3 #(
		.INIT('h5c)
	) name3764 (
		\g1358_reg/NET0131 ,
		\g2788_reg/NET0131 ,
		_w3475_,
		_w4945_
	);
	LUT3 #(
		.INIT('h5c)
	) name3765 (
		\g1378_reg/NET0131 ,
		\g2105_reg/NET0131 ,
		_w3572_,
		_w4946_
	);
	LUT3 #(
		.INIT('h5c)
	) name3766 (
		\g1332_reg/NET0131 ,
		\g2088_reg/NET0131 ,
		_w3667_,
		_w4947_
	);
	LUT3 #(
		.INIT('h5c)
	) name3767 (
		\g1352_reg/NET0131 ,
		\g2098_reg/NET0131 ,
		_w3662_,
		_w4948_
	);
	LUT3 #(
		.INIT('h5c)
	) name3768 (
		\g1358_reg/NET0131 ,
		\g2094_reg/NET0131 ,
		_w3667_,
		_w4949_
	);
	LUT3 #(
		.INIT('h5c)
	) name3769 (
		\g1326_reg/NET0131 ,
		\g2772_reg/NET0131 ,
		_w3672_,
		_w4950_
	);
	LUT3 #(
		.INIT('h5c)
	) name3770 (
		\g1326_reg/NET0131 ,
		\g2773_reg/NET0131 ,
		_w3475_,
		_w4951_
	);
	LUT3 #(
		.INIT('h5c)
	) name3771 (
		\g1326_reg/NET0131 ,
		\g2774_reg/NET0131 ,
		_w3515_,
		_w4952_
	);
	LUT3 #(
		.INIT('h5c)
	) name3772 (
		\g1319_reg/NET0131 ,
		\g2775_reg/NET0131 ,
		_w3672_,
		_w4953_
	);
	LUT3 #(
		.INIT('h5c)
	) name3773 (
		\g1319_reg/NET0131 ,
		\g2776_reg/NET0131 ,
		_w3475_,
		_w4954_
	);
	LUT3 #(
		.INIT('h5c)
	) name3774 (
		\g1319_reg/NET0131 ,
		\g2777_reg/NET0131 ,
		_w3515_,
		_w4955_
	);
	LUT3 #(
		.INIT('h5c)
	) name3775 (
		\g1339_reg/NET0131 ,
		\g2778_reg/NET0131 ,
		_w3672_,
		_w4956_
	);
	LUT3 #(
		.INIT('h5c)
	) name3776 (
		\g1339_reg/NET0131 ,
		\g2779_reg/NET0131 ,
		_w3475_,
		_w4957_
	);
	LUT3 #(
		.INIT('h5c)
	) name3777 (
		\g1339_reg/NET0131 ,
		\g2780_reg/NET0131 ,
		_w3515_,
		_w4958_
	);
	LUT3 #(
		.INIT('h5c)
	) name3778 (
		\g1332_reg/NET0131 ,
		\g2781_reg/NET0131 ,
		_w3672_,
		_w4959_
	);
	LUT3 #(
		.INIT('h5c)
	) name3779 (
		\g1332_reg/NET0131 ,
		\g2782_reg/NET0131 ,
		_w3475_,
		_w4960_
	);
	LUT3 #(
		.INIT('h5c)
	) name3780 (
		\g1332_reg/NET0131 ,
		\g2783_reg/NET0131 ,
		_w3515_,
		_w4961_
	);
	LUT3 #(
		.INIT('h5c)
	) name3781 (
		\g1346_reg/NET0131 ,
		\g2784_reg/NET0131 ,
		_w3672_,
		_w4962_
	);
	LUT3 #(
		.INIT('h5c)
	) name3782 (
		\g1346_reg/NET0131 ,
		\g2785_reg/NET0131 ,
		_w3475_,
		_w4963_
	);
	LUT3 #(
		.INIT('h5c)
	) name3783 (
		\g1346_reg/NET0131 ,
		\g2786_reg/NET0131 ,
		_w3515_,
		_w4964_
	);
	LUT3 #(
		.INIT('h5c)
	) name3784 (
		\g1358_reg/NET0131 ,
		\g2787_reg/NET0131 ,
		_w3672_,
		_w4965_
	);
	LUT3 #(
		.INIT('h5c)
	) name3785 (
		\g1358_reg/NET0131 ,
		\g2789_reg/NET0131 ,
		_w3515_,
		_w4966_
	);
	LUT3 #(
		.INIT('h5c)
	) name3786 (
		\g1352_reg/NET0131 ,
		\g2790_reg/NET0131 ,
		_w3672_,
		_w4967_
	);
	LUT3 #(
		.INIT('h5c)
	) name3787 (
		\g1352_reg/NET0131 ,
		\g2791_reg/NET0131 ,
		_w3475_,
		_w4968_
	);
	LUT3 #(
		.INIT('h5c)
	) name3788 (
		\g1352_reg/NET0131 ,
		\g2792_reg/NET0131 ,
		_w3515_,
		_w4969_
	);
	LUT3 #(
		.INIT('h5c)
	) name3789 (
		\g1365_reg/NET0131 ,
		\g2793_reg/NET0131 ,
		_w3672_,
		_w4970_
	);
	LUT3 #(
		.INIT('h5c)
	) name3790 (
		\g1352_reg/NET0131 ,
		\g2096_reg/NET0131 ,
		_w3572_,
		_w4971_
	);
	LUT3 #(
		.INIT('h5c)
	) name3791 (
		\g1365_reg/NET0131 ,
		\g2794_reg/NET0131 ,
		_w3475_,
		_w4972_
	);
	LUT3 #(
		.INIT('h5c)
	) name3792 (
		\g1365_reg/NET0131 ,
		\g2795_reg/NET0131 ,
		_w3515_,
		_w4973_
	);
	LUT3 #(
		.INIT('h5c)
	) name3793 (
		\g1372_reg/NET0131 ,
		\g2796_reg/NET0131 ,
		_w3672_,
		_w4974_
	);
	LUT3 #(
		.INIT('h5c)
	) name3794 (
		\g1372_reg/NET0131 ,
		\g2797_reg/NET0131 ,
		_w3475_,
		_w4975_
	);
	LUT3 #(
		.INIT('h5c)
	) name3795 (
		\g1372_reg/NET0131 ,
		\g2798_reg/NET0131 ,
		_w3515_,
		_w4976_
	);
	LUT3 #(
		.INIT('h5c)
	) name3796 (
		\g1378_reg/NET0131 ,
		\g2799_reg/NET0131 ,
		_w3672_,
		_w4977_
	);
	LUT3 #(
		.INIT('h5c)
	) name3797 (
		\g1378_reg/NET0131 ,
		\g2800_reg/NET0131 ,
		_w3475_,
		_w4978_
	);
	LUT3 #(
		.INIT('h5c)
	) name3798 (
		\g1378_reg/NET0131 ,
		\g2801_reg/NET0131 ,
		_w3515_,
		_w4979_
	);
	LUT2 #(
		.INIT('h1)
	) name3799 (
		\g1164_reg/NET0131 ,
		\g7961_pad ,
		_w4980_
	);
	LUT3 #(
		.INIT('h0b)
	) name3800 (
		_w1857_,
		_w1858_,
		_w4980_,
		_w4981_
	);
	LUT2 #(
		.INIT('h2)
	) name3801 (
		\g1164_reg/NET0131 ,
		\g7961_pad ,
		_w4982_
	);
	LUT3 #(
		.INIT('hf8)
	) name3802 (
		_w2337_,
		_w4981_,
		_w4982_,
		_w4983_
	);
	LUT3 #(
		.INIT('h6a)
	) name3803 (
		\g2900_reg/NET0131 ,
		_w4658_,
		_w4917_,
		_w4984_
	);
	LUT2 #(
		.INIT('h8)
	) name3804 (
		_w4916_,
		_w4984_,
		_w4985_
	);
	LUT2 #(
		.INIT('h8)
	) name3805 (
		\g2912_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		_w4986_
	);
	LUT4 #(
		.INIT('h1555)
	) name3806 (
		\g2924_reg/NET0131 ,
		_w4659_,
		_w4661_,
		_w4986_,
		_w4987_
	);
	LUT3 #(
		.INIT('h02)
	) name3807 (
		_w4664_,
		_w4666_,
		_w4987_,
		_w4988_
	);
	LUT4 #(
		.INIT('h3313)
	) name3808 (
		\g1024_reg/NET0131 ,
		\g1319_reg/NET0131 ,
		\g1326_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w4989_
	);
	LUT3 #(
		.INIT('h01)
	) name3809 (
		_w3914_,
		_w4687_,
		_w4989_,
		_w4990_
	);
	LUT3 #(
		.INIT('h04)
	) name3810 (
		\g2814_reg/NET0131 ,
		\g2912_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		_w4991_
	);
	LUT4 #(
		.INIT('h0800)
	) name3811 (
		_w4659_,
		_w4661_,
		_w4662_,
		_w4991_,
		_w4992_
	);
	LUT2 #(
		.INIT('h4)
	) name3812 (
		\g2814_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		_w4993_
	);
	LUT4 #(
		.INIT('h7f00)
	) name3813 (
		\g2912_reg/NET0131 ,
		_w4659_,
		_w4661_,
		_w4993_,
		_w4994_
	);
	LUT2 #(
		.INIT('he)
	) name3814 (
		_w4992_,
		_w4994_,
		_w4995_
	);
	LUT4 #(
		.INIT('h9669)
	) name3815 (
		\g2963_reg/NET0131 ,
		\g2966_reg/NET0131 ,
		\g2975_reg/NET0131 ,
		\g2978_reg/NET0131 ,
		_w4996_
	);
	LUT2 #(
		.INIT('h9)
	) name3816 (
		\g2969_reg/NET0131 ,
		\g2972_reg/NET0131 ,
		_w4997_
	);
	LUT2 #(
		.INIT('h2)
	) name3817 (
		\g3139_reg/NET0131 ,
		\g3231_pad ,
		_w4998_
	);
	LUT2 #(
		.INIT('h9)
	) name3818 (
		\g2874_reg/NET0131 ,
		\g2981_reg/NET0131 ,
		_w4999_
	);
	LUT4 #(
		.INIT('h6996)
	) name3819 (
		_w4996_,
		_w4997_,
		_w4998_,
		_w4999_,
		_w5000_
	);
	LUT3 #(
		.INIT('h96)
	) name3820 (
		\g2935_reg/NET0131 ,
		\g2938_reg/NET0131 ,
		\g2959_reg/NET0131 ,
		_w5001_
	);
	LUT3 #(
		.INIT('h69)
	) name3821 (
		\g2941_reg/NET0131 ,
		\g2944_reg/NET0131 ,
		\g2956_reg/NET0131 ,
		_w5002_
	);
	LUT2 #(
		.INIT('h9)
	) name3822 (
		\g2947_reg/NET0131 ,
		\g2953_reg/NET0131 ,
		_w5003_
	);
	LUT4 #(
		.INIT('h9969)
	) name3823 (
		\g2947_reg/NET0131 ,
		\g2953_reg/NET0131 ,
		\g3139_reg/NET0131 ,
		\g3231_pad ,
		_w5004_
	);
	LUT3 #(
		.INIT('h69)
	) name3824 (
		_w5001_,
		_w5002_,
		_w5004_,
		_w5005_
	);
	LUT4 #(
		.INIT('h6996)
	) name3825 (
		\g2934_reg/NET0131 ,
		_w5001_,
		_w5002_,
		_w5003_,
		_w5006_
	);
	LUT4 #(
		.INIT('h9669)
	) name3826 (
		\g2962_reg/NET0131 ,
		_w4996_,
		_w4997_,
		_w4999_,
		_w5007_
	);
	LUT2 #(
		.INIT('h4)
	) name3827 (
		\g2814_reg/NET0131 ,
		\g2912_reg/NET0131 ,
		_w5008_
	);
	LUT4 #(
		.INIT('h0800)
	) name3828 (
		_w4659_,
		_w4661_,
		_w4662_,
		_w5008_,
		_w5009_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		\g2814_reg/NET0131 ,
		\g2912_reg/NET0131 ,
		_w5010_
	);
	LUT3 #(
		.INIT('h70)
	) name3830 (
		_w4659_,
		_w4661_,
		_w5010_,
		_w5011_
	);
	LUT2 #(
		.INIT('h1)
	) name3831 (
		_w5009_,
		_w5011_,
		_w5012_
	);
	LUT2 #(
		.INIT('h6)
	) name3832 (
		\g3002_reg/NET0131 ,
		_w4616_,
		_w5013_
	);
	LUT2 #(
		.INIT('h8)
	) name3833 (
		_w4615_,
		_w5013_,
		_w5014_
	);
	LUT3 #(
		.INIT('h6c)
	) name3834 (
		\g2993_reg/NET0131 ,
		\g2998_reg/NET0131 ,
		\g3080_reg/NET0131 ,
		_w5015_
	);
	LUT4 #(
		.INIT('hbfaa)
	) name3835 (
		\g3234_pad ,
		_w3309_,
		_w4580_,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name3836 (
		\g1869_reg/NET0131 ,
		\g5657_pad ,
		_w5017_
	);
	LUT4 #(
		.INIT('hf531)
	) name3837 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1867_reg/NET0131 ,
		\g1868_reg/NET0131 ,
		_w5018_
	);
	LUT2 #(
		.INIT('h4)
	) name3838 (
		_w5017_,
		_w5018_,
		_w5019_
	);
	LUT2 #(
		.INIT('h4)
	) name3839 (
		\g488_reg/NET0131 ,
		\g5657_pad ,
		_w5020_
	);
	LUT4 #(
		.INIT('hf531)
	) name3840 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g486_reg/NET0131 ,
		\g487_reg/NET0131 ,
		_w5021_
	);
	LUT2 #(
		.INIT('h4)
	) name3841 (
		_w5020_,
		_w5021_,
		_w5022_
	);
	LUT2 #(
		.INIT('h4)
	) name3842 (
		\g1860_reg/NET0131 ,
		\g5657_pad ,
		_w5023_
	);
	LUT4 #(
		.INIT('hf531)
	) name3843 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1858_reg/NET0131 ,
		\g1859_reg/NET0131 ,
		_w5024_
	);
	LUT2 #(
		.INIT('h4)
	) name3844 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT3 #(
		.INIT('h10)
	) name3845 (
		\g2912_reg/NET0131 ,
		\g2920_reg/NET0131 ,
		\g2924_reg/NET0131 ,
		_w5026_
	);
	LUT4 #(
		.INIT('h0008)
	) name3846 (
		\g1088_reg/NET0131 ,
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		_w5027_
	);
	LUT4 #(
		.INIT('h8000)
	) name3847 (
		_w4071_,
		_w4072_,
		_w5026_,
		_w5027_,
		_w5028_
	);
	LUT4 #(
		.INIT('h0200)
	) name3848 (
		\g801_reg/NET0131 ,
		\g805_reg/NET0131 ,
		\g809_reg/NET0131 ,
		\g813_reg/NET0131 ,
		_w5029_
	);
	LUT3 #(
		.INIT('he2)
	) name3849 (
		\g856_reg/NET0131 ,
		_w5028_,
		_w5029_,
		_w5030_
	);
	LUT4 #(
		.INIT('h0200)
	) name3850 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		\g7961_pad ,
		_w5031_
	);
	LUT4 #(
		.INIT('h8000)
	) name3851 (
		_w4071_,
		_w4072_,
		_w5026_,
		_w5031_,
		_w5032_
	);
	LUT3 #(
		.INIT('hca)
	) name3852 (
		\g857_reg/NET0131 ,
		_w5029_,
		_w5032_,
		_w5033_
	);
	LUT4 #(
		.INIT('h0008)
	) name3853 (
		\g1092_reg/NET0131 ,
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		_w5034_
	);
	LUT4 #(
		.INIT('h8000)
	) name3854 (
		_w4071_,
		_w4072_,
		_w5026_,
		_w5034_,
		_w5035_
	);
	LUT3 #(
		.INIT('hca)
	) name3855 (
		\g858_reg/NET0131 ,
		_w5029_,
		_w5035_,
		_w5036_
	);
	LUT2 #(
		.INIT('h4)
	) name3856 (
		\g479_reg/NET0131 ,
		\g5657_pad ,
		_w5037_
	);
	LUT4 #(
		.INIT('hf531)
	) name3857 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g477_reg/NET0131 ,
		\g478_reg/NET0131 ,
		_w5038_
	);
	LUT2 #(
		.INIT('h4)
	) name3858 (
		_w5037_,
		_w5038_,
		_w5039_
	);
	LUT4 #(
		.INIT('h0200)
	) name3859 (
		\g2185_reg/NET0131 ,
		\g2190_reg/NET0131 ,
		\g2195_reg/NET0131 ,
		\g2200_reg/NET0131 ,
		_w5040_
	);
	LUT3 #(
		.INIT('he2)
	) name3860 (
		\g2244_reg/NET0131 ,
		_w5028_,
		_w5040_,
		_w5041_
	);
	LUT3 #(
		.INIT('he2)
	) name3861 (
		\g2245_reg/NET0131 ,
		_w5032_,
		_w5040_,
		_w5042_
	);
	LUT3 #(
		.INIT('he2)
	) name3862 (
		\g2246_reg/NET0131 ,
		_w5035_,
		_w5040_,
		_w5043_
	);
	LUT2 #(
		.INIT('h4)
	) name3863 (
		\g1166_reg/NET0131 ,
		\g5657_pad ,
		_w5044_
	);
	LUT4 #(
		.INIT('hf531)
	) name3864 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1164_reg/NET0131 ,
		\g1165_reg/NET0131 ,
		_w5045_
	);
	LUT2 #(
		.INIT('h4)
	) name3865 (
		_w5044_,
		_w5045_,
		_w5046_
	);
	LUT2 #(
		.INIT('h4)
	) name3866 (
		\g464_reg/NET0131 ,
		\g5657_pad ,
		_w5047_
	);
	LUT4 #(
		.INIT('hf531)
	) name3867 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g480_reg/NET0131 ,
		\g484_reg/NET0131 ,
		_w5048_
	);
	LUT2 #(
		.INIT('h4)
	) name3868 (
		_w5047_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h4)
	) name3869 (
		\g1151_reg/NET0131 ,
		\g5657_pad ,
		_w5050_
	);
	LUT4 #(
		.INIT('hf531)
	) name3870 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1167_reg/NET0131 ,
		\g1171_reg/NET0131 ,
		_w5051_
	);
	LUT2 #(
		.INIT('h4)
	) name3871 (
		_w5050_,
		_w5051_,
		_w5052_
	);
	LUT2 #(
		.INIT('h4)
	) name3872 (
		\g1175_reg/NET0131 ,
		\g5657_pad ,
		_w5053_
	);
	LUT4 #(
		.INIT('hf531)
	) name3873 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1173_reg/NET0131 ,
		\g1174_reg/NET0131 ,
		_w5054_
	);
	LUT2 #(
		.INIT('h4)
	) name3874 (
		_w5053_,
		_w5054_,
		_w5055_
	);
	LUT3 #(
		.INIT('h06)
	) name3875 (
		\g2993_reg/NET0131 ,
		\g3080_reg/NET0131 ,
		\g3234_pad ,
		_w5056_
	);
	LUT2 #(
		.INIT('h4)
	) name3876 (
		\g2554_reg/NET0131 ,
		\g5657_pad ,
		_w5057_
	);
	LUT4 #(
		.INIT('hf531)
	) name3877 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2552_reg/NET0131 ,
		\g2553_reg/NET0131 ,
		_w5058_
	);
	LUT2 #(
		.INIT('h4)
	) name3878 (
		_w5057_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h4)
	) name3879 (
		\g2539_reg/NET0131 ,
		\g5657_pad ,
		_w5060_
	);
	LUT4 #(
		.INIT('hf531)
	) name3880 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2555_reg/NET0131 ,
		\g2559_reg/NET0131 ,
		_w5061_
	);
	LUT2 #(
		.INIT('h4)
	) name3881 (
		_w5060_,
		_w5061_,
		_w5062_
	);
	LUT2 #(
		.INIT('h4)
	) name3882 (
		\g2563_reg/NET0131 ,
		\g5657_pad ,
		_w5063_
	);
	LUT4 #(
		.INIT('hf531)
	) name3883 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g2561_reg/NET0131 ,
		\g2562_reg/NET0131 ,
		_w5064_
	);
	LUT2 #(
		.INIT('h4)
	) name3884 (
		_w5063_,
		_w5064_,
		_w5065_
	);
	LUT2 #(
		.INIT('h4)
	) name3885 (
		\g1845_reg/NET0131 ,
		\g5657_pad ,
		_w5066_
	);
	LUT4 #(
		.INIT('hf531)
	) name3886 (
		\g1018_reg/NET0131 ,
		\g1024_reg/NET0131 ,
		\g1861_reg/NET0131 ,
		\g1865_reg/NET0131 ,
		_w5067_
	);
	LUT2 #(
		.INIT('h4)
	) name3887 (
		_w5066_,
		_w5067_,
		_w5068_
	);
	LUT3 #(
		.INIT('h3a)
	) name3888 (
		\g2253_reg/NET0131 ,
		_w3968_,
		_w5028_,
		_w5069_
	);
	LUT3 #(
		.INIT('h3a)
	) name3889 (
		\g2254_reg/NET0131 ,
		_w3968_,
		_w5032_,
		_w5070_
	);
	LUT3 #(
		.INIT('h3a)
	) name3890 (
		\g2255_reg/NET0131 ,
		_w3968_,
		_w5035_,
		_w5071_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3891 (
		\g2993_reg/NET0131 ,
		\g2998_reg/NET0131 ,
		\g3006_reg/NET0131 ,
		\g3080_reg/NET0131 ,
		_w5072_
	);
	LUT4 #(
		.INIT('h1500)
	) name3892 (
		\g3234_pad ,
		_w3309_,
		_w4580_,
		_w5072_,
		_w5073_
	);
	LUT3 #(
		.INIT('h41)
	) name3893 (
		\g2814_reg/NET0131 ,
		\g2883_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		_w5074_
	);
	LUT3 #(
		.INIT('h8f)
	) name3894 (
		_w4659_,
		_w4661_,
		_w5074_,
		_w5075_
	);
	LUT2 #(
		.INIT('h6)
	) name3895 (
		\g2892_reg/NET0131 ,
		_w4917_,
		_w5076_
	);
	LUT2 #(
		.INIT('h8)
	) name3896 (
		_w4916_,
		_w5076_,
		_w5077_
	);
	LUT3 #(
		.INIT('h6c)
	) name3897 (
		\g2892_reg/NET0131 ,
		\g2903_reg/NET0131 ,
		_w4917_,
		_w5078_
	);
	LUT2 #(
		.INIT('h8)
	) name3898 (
		_w4916_,
		_w5078_,
		_w5079_
	);
	LUT3 #(
		.INIT('h6c)
	) name3899 (
		\g3002_reg/NET0131 ,
		\g3013_reg/NET0131 ,
		_w4616_,
		_w5080_
	);
	LUT2 #(
		.INIT('h8)
	) name3900 (
		_w4615_,
		_w5080_,
		_w5081_
	);
	LUT3 #(
		.INIT('h06)
	) name3901 (
		\g1326_reg/NET0131 ,
		_w3521_,
		_w3914_,
		_w5082_
	);
	LUT3 #(
		.INIT('h6c)
	) name3902 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		_w5083_
	);
	LUT4 #(
		.INIT('h1500)
	) name3903 (
		\g2814_reg/NET0131 ,
		_w4659_,
		_w4661_,
		_w5083_,
		_w5084_
	);
	LUT4 #(
		.INIT('h78f0)
	) name3904 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		\g2896_reg/NET0131 ,
		\g2950_reg/NET0131 ,
		_w5085_
	);
	LUT4 #(
		.INIT('h1500)
	) name3905 (
		\g2814_reg/NET0131 ,
		_w4659_,
		_w4661_,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('he)
	) name3906 (
		\g2933_reg/NET0131 ,
		\g51_pad ,
		_w5087_
	);
	LUT3 #(
		.INIT('h02)
	) name3907 (
		\g2883_reg/NET0131 ,
		\g2888_reg/NET0131 ,
		\g2917_reg/NET0131 ,
		_w5088_
	);
	LUT4 #(
		.INIT('h8000)
	) name3908 (
		_w4071_,
		_w4072_,
		_w5026_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('he)
	) name3909 (
		\g3079_reg/NET0131 ,
		\g3234_pad ,
		_w5090_
	);
	LUT2 #(
		.INIT('h4)
	) name3910 (
		\g1024_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		_w5091_
	);
	LUT4 #(
		.INIT('h000e)
	) name3911 (
		\g1024_reg/NET0131 ,
		\g1345_reg/NET0131 ,
		\g3002_reg/NET0131 ,
		\g3006_reg/NET0131 ,
		_w5092_
	);
	LUT3 #(
		.INIT('hec)
	) name3912 (
		_w4365_,
		_w5091_,
		_w5092_,
		_w5093_
	);
	LUT3 #(
		.INIT('h72)
	) name3913 (
		\g1024_reg/NET0131 ,
		\g1240_reg/NET0131 ,
		\g1243_reg/NET0131 ,
		_w5094_
	);
	LUT3 #(
		.INIT('h5c)
	) name3914 (
		\g291_reg/NET0131 ,
		\g305_reg/NET0131 ,
		\g3229_pad ,
		_w5095_
	);
	LUT3 #(
		.INIT('h72)
	) name3915 (
		\g3229_pad ,
		\g978_reg/NET0131 ,
		\g992_reg/NET0131 ,
		_w5096_
	);
	LUT3 #(
		.INIT('h3b)
	) name3916 (
		\g2814_reg/NET0131 ,
		\g2879_reg/NET0131 ,
		\g2929_reg/NET0131 ,
		_w5097_
	);
	LUT3 #(
		.INIT('h5c)
	) name3917 (
		\g1672_reg/NET0131 ,
		\g1686_reg/NET0131 ,
		\g3229_pad ,
		_w5098_
	);
	LUT3 #(
		.INIT('h5c)
	) name3918 (
		\g2366_reg/NET0131 ,
		\g2380_reg/NET0131 ,
		\g3229_pad ,
		_w5099_
	);
	LUT2 #(
		.INIT('h2)
	) name3919 (
		\g2817_reg/NET0131 ,
		\g51_pad ,
		_w5100_
	);
	LUT2 #(
		.INIT('h2)
	) name3920 (
		\g3054_reg/NET0131 ,
		\g3234_pad ,
		_w5101_
	);
	LUT4 #(
		.INIT('h0200)
	) name3921 (
		\g113_reg/NET0131 ,
		\g117_reg/NET0131 ,
		\g121_reg/NET0131 ,
		\g125_reg/NET0131 ,
		_w5102_
	);
	LUT4 #(
		.INIT('h0200)
	) name3922 (
		\g1491_reg/NET0131 ,
		\g1496_reg/NET0131 ,
		\g1501_reg/NET0131 ,
		\g1506_reg/NET0131 ,
		_w5103_
	);
	LUT2 #(
		.INIT('h2)
	) name3923 (
		\g2950_reg/NET0131 ,
		\g51_pad ,
		_w5104_
	);
	LUT2 #(
		.INIT('h2)
	) name3924 (
		\g3080_reg/NET0131 ,
		\g3234_pad ,
		_w5105_
	);
	LUT2 #(
		.INIT('h2)
	) name3925 (
		\g121_reg/NET0131 ,
		_w2315_,
		_w5106_
	);
	LUT3 #(
		.INIT('h80)
	) name3926 (
		\g121_reg/NET0131 ,
		_w1711_,
		_w2310_,
		_w5107_
	);
	LUT3 #(
		.INIT('hd0)
	) name3927 (
		_w1737_,
		_w2306_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h1)
	) name3928 (
		_w5106_,
		_w5108_,
		_w5109_
	);
	LUT3 #(
		.INIT('h9c)
	) name3929 (
		_w1697_,
		_w1774_,
		_w1821_,
		_w5110_
	);
	LUT3 #(
		.INIT('h6a)
	) name3930 (
		_w1787_,
		_w2710_,
		_w5110_,
		_w5111_
	);
	LUT2 #(
		.INIT('h2)
	) name3931 (
		_w2315_,
		_w2328_,
		_w5112_
	);
	LUT3 #(
		.INIT('h10)
	) name3932 (
		_w2314_,
		_w5111_,
		_w5112_,
		_w5113_
	);
	LUT2 #(
		.INIT('hd)
	) name3933 (
		_w5109_,
		_w5113_,
		_w5114_
	);
	LUT4 #(
		.INIT('h88d8)
	) name3934 (
		\g499_reg/NET0131 ,
		\g544_reg/NET0131 ,
		\g548_reg/NET0131 ,
		\g5657_pad ,
		_w5115_
	);
	LUT3 #(
		.INIT('h8a)
	) name3935 (
		\g2190_reg/NET0131 ,
		_w2477_,
		_w2480_,
		_w5116_
	);
	LUT2 #(
		.INIT('h8)
	) name3936 (
		\g2190_reg/NET0131 ,
		_w2472_,
		_w5117_
	);
	LUT4 #(
		.INIT('h020f)
	) name3937 (
		_w1333_,
		_w2466_,
		_w5116_,
		_w5117_,
		_w5118_
	);
	LUT3 #(
		.INIT('h02)
	) name3938 (
		_w2495_,
		_w2550_,
		_w2552_,
		_w5119_
	);
	LUT3 #(
		.INIT('h95)
	) name3939 (
		_w1265_,
		_w2585_,
		_w5119_,
		_w5120_
	);
	LUT2 #(
		.INIT('h8)
	) name3940 (
		_w2498_,
		_w5120_,
		_w5121_
	);
	LUT3 #(
		.INIT('h73)
	) name3941 (
		_w2473_,
		_w5118_,
		_w5121_,
		_w5122_
	);
	LUT2 #(
		.INIT('h1)
	) name3942 (
		\g1088_reg/NET0131 ,
		\g246_reg/NET0131 ,
		_w5123_
	);
	LUT2 #(
		.INIT('h4)
	) name3943 (
		\g1088_reg/NET0131 ,
		\g246_reg/NET0131 ,
		_w5124_
	);
	LUT4 #(
		.INIT('ha8fc)
	) name3944 (
		_w2314_,
		_w2642_,
		_w2644_,
		_w2646_,
		_w5125_
	);
	LUT3 #(
		.INIT('h0b)
	) name3945 (
		_w2314_,
		_w2656_,
		_w5123_,
		_w5126_
	);
	LUT3 #(
		.INIT('hba)
	) name3946 (
		_w5124_,
		_w5125_,
		_w5126_,
		_w5127_
	);
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g101_reg/P0001  = _w16_ ;
	assign \g105_reg/P0001  = _w31_ ;
	assign \g109_reg/P0001  = _w51_ ;
	assign \g1138_reg/P0001  = _w69_ ;
	assign \g113_reg/P0001  = _w71_ ;
	assign \g1140_reg/P0001  = _w73_ ;
	assign \g117_reg/P0001  = _w86_ ;
	assign \g121_reg/P0001  = _w101_ ;
	assign \g125_reg/P0001  = _w120_ ;
	assign \g1471_reg/P0001  = _w222_ ;
	assign \g1476_reg/P0001  = _w224_ ;
	assign \g1481_reg/P0001  = _w227_ ;
	assign \g1486_reg/P0001  = _w229_ ;
	assign \g1491_reg/P0001  = _w232_ ;
	assign \g1496_reg/P0001  = _w234_ ;
	assign \g1501_reg/P0001  = _w237_ ;
	assign \g1506_reg/P0001  = _w239_ ;
	assign \g16496_pad  = _w1250_ ;
	assign \g1660_reg/P0001  = _w333_ ;
	assign \g1662_reg/P0001  = _w335_ ;
	assign \g1664_reg/P0001  = _w337_ ;
	assign \g1666_reg/P0001  = _w339_ ;
	assign \g1668_reg/P0001  = _w341_ ;
	assign \g1670_reg/P0001  = _w343_ ;
	assign \g1672_reg/P0001  = _w345_ ;
	assign \g18/_0_  = _w1389_ ;
	assign \g1832_reg/P0001  = _w419_ ;
	assign \g1834_reg/P0001  = _w421_ ;
	assign \g2165_reg/P0001  = _w541_ ;
	assign \g2170_reg/P0001  = _w544_ ;
	assign \g2175_reg/P0001  = _w546_ ;
	assign \g2180_reg/P0001  = _w548_ ;
	assign \g2185_reg/P0001  = _w550_ ;
	assign \g2190_reg/P0001  = _w552_ ;
	assign \g2195_reg/P0001  = _w554_ ;
	assign \g2200_reg/P0001  = _w557_ ;
	assign \g2354_reg/P0001  = _w636_ ;
	assign \g2356_reg/P0001  = _w638_ ;
	assign \g2358_reg/P0001  = _w640_ ;
	assign \g2360_reg/P0001  = _w642_ ;
	assign \g2362_reg/P0001  = _w644_ ;
	assign \g2364_reg/P0001  = _w646_ ;
	assign \g2366_reg/P0001  = _w648_ ;
	assign \g2526_reg/P0001  = _w715_ ;
	assign \g2528_reg/P0001  = _w717_ ;
	assign \g25489_pad  = _w1395_ ;
	assign \g279_reg/P0001  = _w820_ ;
	assign \g281_reg/P0001  = _w838_ ;
	assign \g283_reg/P0001  = _w840_ ;
	assign \g285_reg/P0001  = _w842_ ;
	assign \g2879_reg/NET0131_syn_2  = _w845_ ;
	assign \g287_reg/P0001  = _w847_ ;
	assign \g289_reg/P0001  = _w853_ ;
	assign \g291_reg/P0001  = _w860_ ;
	assign \g451_reg/P0001  = _w1012_ ;
	assign \g453_reg/P0001  = _w1014_ ;
	assign \g59421/_3_  = _w1399_ ;
	assign \g59425/_1_  = _w1403_ ;
	assign \g59435/_0_  = _w1407_ ;
	assign \g59436/_0_  = _w1409_ ;
	assign \g59441/_3_  = _w1410_ ;
	assign \g59442/_0_  = _w1414_ ;
	assign \g59445/_0_  = _w1415_ ;
	assign \g59453/_0_  = _w1524_ ;
	assign \g59462/_3_  = _w1525_ ;
	assign \g59466/_3_  = _w1526_ ;
	assign \g59467/_3_  = _w1527_ ;
	assign \g59468/_3_  = _w1528_ ;
	assign \g59469/_3_  = _w1529_ ;
	assign \g59470/_3_  = _w1530_ ;
	assign \g59471/_3_  = _w1531_ ;
	assign \g59472/_3_  = _w1532_ ;
	assign \g59473/_3_  = _w1533_ ;
	assign \g59489/_0_  = _w1612_ ;
	assign \g59498/_0_  = _w1628_ ;
	assign \g59499/_0_  = _w1634_ ;
	assign \g59500/_0_  = _w1640_ ;
	assign \g59502/_2_  = _w1648_ ;
	assign \g59503/_0_  = _w1652_ ;
	assign \g59505/_2_  = _w1658_ ;
	assign \g59507/_0_  = _w1667_ ;
	assign \g59508/_0_  = _w1674_ ;
	assign \g59533/_3_  = _w1675_ ;
	assign \g59534/_3_  = _w1676_ ;
	assign \g59535/_3_  = _w1677_ ;
	assign \g59536/_3_  = _w1678_ ;
	assign \g59537/_3_  = _w1679_ ;
	assign \g59538/_3_  = _w1680_ ;
	assign \g59539/_3_  = _w1681_ ;
	assign \g59540/_3_  = _w1682_ ;
	assign \g59548/_0_  = _w1693_ ;
	assign \g59550/_0_  = _w1834_ ;
	assign \g59551/_0_  = _w1839_ ;
	assign \g59552/_0_  = _w1844_ ;
	assign \g59554/_0_  = _w1996_ ;
	assign \g59555/_0_  = _w1997_ ;
	assign \g59556/_0_  = _w1998_ ;
	assign \g59557/_0_  = _w2002_ ;
	assign \g59558/_0_  = _w2006_ ;
	assign \g59559/_0_  = _w2149_ ;
	assign \g59560/_0_  = _w2156_ ;
	assign \g59561/_0_  = _w2163_ ;
	assign \g59639/_0_  = _w2239_ ;
	assign \g59694/_2_  = _w2254_ ;
	assign \g59695/_0_  = _w2261_ ;
	assign \g59697/_2_  = _w2268_ ;
	assign \g59698/_0_  = _w2275_ ;
	assign \g59699/_0_  = _w2284_ ;
	assign \g59700/_0_  = _w2288_ ;
	assign \g59705/_0_  = _w2334_ ;
	assign \g59706/_0_  = _w2335_ ;
	assign \g59707/_0_  = _w2336_ ;
	assign \g59708/_0_  = _w2371_ ;
	assign \g59709/_0_  = _w2372_ ;
	assign \g59710/_0_  = _w2373_ ;
	assign \g59711/_0_  = _w2382_ ;
	assign \g59712/_0_  = _w2383_ ;
	assign \g59713/_0_  = _w2384_ ;
	assign \g59714/_0_  = _w2394_ ;
	assign \g59715/_0_  = _w2395_ ;
	assign \g59716/_0_  = _w2396_ ;
	assign \g59717/_0_  = _w2421_ ;
	assign \g59718/_0_  = _w2425_ ;
	assign \g59719/_0_  = _w2429_ ;
	assign \g59720/_0_  = _w2463_ ;
	assign \g59721/_0_  = _w2505_ ;
	assign \g59722/_0_  = _w2509_ ;
	assign \g59723/_0_  = _w2513_ ;
	assign \g59724/_0_  = _w2518_ ;
	assign \g59725/_0_  = _w2528_ ;
	assign \g59726/_0_  = _w2533_ ;
	assign \g59727/_0_  = _w2537_ ;
	assign \g59728/_0_  = _w2541_ ;
	assign \g59729/_0_  = _w2559_ ;
	assign \g59730/_0_  = _w2563_ ;
	assign \g59731/_0_  = _w2572_ ;
	assign \g59732/_0_  = _w2576_ ;
	assign \g59733/_0_  = _w2593_ ;
	assign \g59734/_0_  = _w2597_ ;
	assign \g59735/_0_  = _w2601_ ;
	assign \g59736/_0_  = _w2602_ ;
	assign \g59737/_0_  = _w2603_ ;
	assign \g59738/_0_  = _w2611_ ;
	assign \g59739/_0_  = _w2616_ ;
	assign \g59740/_0_  = _w2621_ ;
	assign \g59741/_0_  = _w2635_ ;
	assign \g59742/_0_  = _w2640_ ;
	assign \g59743/_0_  = _w2658_ ;
	assign \g59744/_0_  = _w2663_ ;
	assign \g59745/_0_  = _w2669_ ;
	assign \g59747/_0_  = _w2691_ ;
	assign \g59748/_0_  = _w2695_ ;
	assign \g59749/_0_  = _w2699_ ;
	assign \g59750/_0_  = _w2722_ ;
	assign \g59751/_0_  = _w2726_ ;
	assign \g59752/_0_  = _w2730_ ;
	assign \g59753/_0_  = _w2737_ ;
	assign \g59754/_0_  = _w2743_ ;
	assign \g59755/_0_  = _w2755_ ;
	assign \g59756/_0_  = _w2759_ ;
	assign \g59757/_0_  = _w2763_ ;
	assign \g59758/_0_  = _w2774_ ;
	assign \g59759/_0_  = _w2778_ ;
	assign \g59760/_0_  = _w2782_ ;
	assign \g59761/_0_  = _w2795_ ;
	assign \g59762/_0_  = _w2799_ ;
	assign \g59763/_0_  = _w2803_ ;
	assign \g59764/_0_  = _w2812_ ;
	assign \g59765/_0_  = _w2816_ ;
	assign \g59766/_0_  = _w2820_ ;
	assign \g59915/_0_  = _w2908_ ;
	assign \g59952/_2_  = _w2911_ ;
	assign \g60046/_0_  = _w2922_ ;
	assign \g60048/_0_  = _w2931_ ;
	assign \g60049/_0_  = _w2939_ ;
	assign \g60051/_0_  = _w2949_ ;
	assign \g60063/_0_  = _w2959_ ;
	assign \g60103/_0_  = _w2966_ ;
	assign \g60104/_0_  = _w2973_ ;
	assign \g60105/_0_  = _w2990_ ;
	assign \g60107/_2_  = _w3002_ ;
	assign \g60108/_0_  = _w3008_ ;
	assign \g60109/_0_  = _w3018_ ;
	assign \g60110/_0_  = _w3022_ ;
	assign \g60112/_2_  = _w3028_ ;
	assign \g60119/_0_  = _w3034_ ;
	assign \g60120/_0_  = _w3044_ ;
	assign \g60121/_0_  = _w3051_ ;
	assign \g60122/_0_  = _w3058_ ;
	assign \g60123/_0_  = _w3061_ ;
	assign \g60124/_0_  = _w3068_ ;
	assign \g60126/_0_  = _w3076_ ;
	assign \g60127/_0_  = _w3087_ ;
	assign \g60128/_0_  = _w3093_ ;
	assign \g60129/_0_  = _w3096_ ;
	assign \g60130/_0_  = _w3099_ ;
	assign \g60135/_0_  = _w3113_ ;
	assign \g60136/_0_  = _w3121_ ;
	assign \g60137/_0_  = _w3127_ ;
	assign \g60138/_0_  = _w3137_ ;
	assign \g60139/_0_  = _w3145_ ;
	assign \g60143/_3_  = _w3146_ ;
	assign \g60144/_0_  = _w3155_ ;
	assign \g60145/_0_  = _w3162_ ;
	assign \g60339/_0_  = _w3163_ ;
	assign \g60404/_0_  = _w3167_ ;
	assign \g60427/_0_  = _w3171_ ;
	assign \g60428/_0_  = _w3173_ ;
	assign \g60429/_0_  = _w3177_ ;
	assign \g60434/_0_  = _w3191_ ;
	assign \g60435/_0_  = _w3197_ ;
	assign \g60437/_0_  = _w3203_ ;
	assign \g60438/_0_  = _w3209_ ;
	assign \g60439/_0_  = _w3214_ ;
	assign \g60440/_0_  = _w3218_ ;
	assign \g60441/_0_  = _w3219_ ;
	assign \g60448/_0_  = _w3320_ ;
	assign \g60451/_0_  = _w3410_ ;
	assign \g60452/_0_  = _w3416_ ;
	assign \g60453/_0_  = _w3420_ ;
	assign \g60459/_0_  = _w3426_ ;
	assign \g60460/_0_  = _w3432_ ;
	assign \g60523/_0_  = _w3433_ ;
	assign \g60534/_0_  = _w3443_ ;
	assign \g60535/_0_  = _w3447_ ;
	assign \g60536/_0_  = _w3451_ ;
	assign \g60585/_0_  = _w3458_ ;
	assign \g60586/_0_  = _w3464_ ;
	assign \g60587/_0_  = _w3470_ ;
	assign \g60588/_0_  = _w3474_ ;
	assign \g60591/_0_  = _w3514_ ;
	assign \g60592/_0_  = _w3519_ ;
	assign \g60599/_0_  = _w3561_ ;
	assign \g60601/_0_  = _w3566_ ;
	assign \g60602/_0_  = _w3571_ ;
	assign \g60603/_0_  = _w3611_ ;
	assign \g60604/_0_  = _w3651_ ;
	assign \g60605/_0_  = _w3656_ ;
	assign \g60606/_0_  = _w3661_ ;
	assign \g60607/_0_  = _w3666_ ;
	assign \g60608/_0_  = _w3671_ ;
	assign \g60609/_0_  = _w3676_ ;
	assign \g60613/_0_  = _w3761_ ;
	assign \g60614/_0_  = _w3851_ ;
	assign \g60615/_0_  = _w3853_ ;
	assign \g60694/_0_  = _w3854_ ;
	assign \g60708/_0_  = _w3860_ ;
	assign \g60709/_0_  = _w3868_ ;
	assign \g60710/_0_  = _w3874_ ;
	assign \g60785/_0_  = _w3878_ ;
	assign \g60787/_0_  = _w3880_ ;
	assign \g60788/_0_  = _w3882_ ;
	assign \g60799/_0_  = _w3885_ ;
	assign \g60801/_0_  = _w3887_ ;
	assign \g60802/_0_  = _w3889_ ;
	assign \g60803/_1__syn_2  = _w3893_ ;
	assign \g60805/_1__syn_2  = _w3895_ ;
	assign \g60806/_1__syn_2  = _w3897_ ;
	assign \g60808/_0_  = _w3900_ ;
	assign \g60810/_0_  = _w3902_ ;
	assign \g60811/_0_  = _w3904_ ;
	assign \g60825/_3_  = _w3907_ ;
	assign \g60896/_0_  = _w3918_ ;
	assign \g60980/_0_  = _w3936_ ;
	assign \g60981/_0_  = _w3954_ ;
	assign \g60985/_0_  = _w3971_ ;
	assign \g60986/_0_  = _w3989_ ;
	assign \g61012/_0_  = _w3991_ ;
	assign \g61013/_0_  = _w3992_ ;
	assign \g61015/_0_  = _w3994_ ;
	assign \g61017/_0_  = _w3996_ ;
	assign \g61122/_0_  = _w4002_ ;
	assign \g61123/_0_  = _w4008_ ;
	assign \g61124/_0_  = _w4014_ ;
	assign \g61125/_0_  = _w4020_ ;
	assign \g61222/_0_  = _w4021_ ;
	assign \g61223/_0_  = _w4022_ ;
	assign \g61224/_0_  = _w4023_ ;
	assign \g61225/_0_  = _w4024_ ;
	assign \g61228/_0_  = _w4025_ ;
	assign \g61229/_0_  = _w4026_ ;
	assign \g61230/_0_  = _w4027_ ;
	assign \g61231/_0_  = _w4028_ ;
	assign \g61281/_0_  = _w4032_ ;
	assign \g61293/_1_  = _w4033_ ;
	assign \g61307/_0__syn_2  = _w4035_ ;
	assign \g61309/_0__syn_2  = _w4037_ ;
	assign \g61310/_0__syn_2  = _w4039_ ;
	assign \g61311/_1_  = _w4041_ ;
	assign \g61312/_1_  = _w4043_ ;
	assign \g61313/_1_  = _w4045_ ;
	assign \g61324/_1_  = _w4047_ ;
	assign \g61325/_1_  = _w4049_ ;
	assign \g61326/_1_  = _w4051_ ;
	assign \g61328/_1_  = _w4053_ ;
	assign \g61329/_1_  = _w4055_ ;
	assign \g61330/_1_  = _w4057_ ;
	assign \g61332/_1_  = _w4094_ ;
	assign \g61333/_1_  = _w4134_ ;
	assign \g61334/_1_  = _w4172_ ;
	assign \g61335/_1_  = _w4211_ ;
	assign \g61336/_0_  = _w4220_ ;
	assign \g61338/_0_  = _w4228_ ;
	assign \g61339/_0_  = _w4234_ ;
	assign \g61340/_0_  = _w4238_ ;
	assign \g61377/_1_  = _w4255_ ;
	assign \g61378/_1_  = _w4256_ ;
	assign \g61379/_1_  = _w4257_ ;
	assign \g61388/_1_  = _w4275_ ;
	assign \g61391/_0_  = _w4287_ ;
	assign \g61394/_1_  = _w4288_ ;
	assign \g61395/_1_  = _w4289_ ;
	assign \g61396/_1_  = _w4305_ ;
	assign \g61398/_1_  = _w4306_ ;
	assign \g61399/_1_  = _w4307_ ;
	assign \g61421/_1_  = _w4325_ ;
	assign \g61422/_1_  = _w4326_ ;
	assign \g61423/_1_  = _w4327_ ;
	assign \g61524/_0_  = _w4348_ ;
	assign \g61525/_0_  = _w4353_ ;
	assign \g61526/_0_  = _w4358_ ;
	assign \g61527/_0_  = _w4372_ ;
	assign \g61528/_0_  = _w4375_ ;
	assign \g61529/_0_  = _w4378_ ;
	assign \g61530/_0_  = _w4397_ ;
	assign \g61531/_0_  = _w4401_ ;
	assign \g61532/_0_  = _w4405_ ;
	assign \g61533/_0_  = _w4412_ ;
	assign \g61534/_0_  = _w4413_ ;
	assign \g61535/_0_  = _w4414_ ;
	assign \g61536/_0_  = _w4425_ ;
	assign \g61537/_0_  = _w4428_ ;
	assign \g61538/_0_  = _w4431_ ;
	assign \g61539/_0_  = _w4432_ ;
	assign \g61540/_0_  = _w4442_ ;
	assign \g61541/_0_  = _w4445_ ;
	assign \g61542/_0_  = _w4448_ ;
	assign \g61543/_0_  = _w4452_ ;
	assign \g61544/_0_  = _w4471_ ;
	assign \g61545/_0_  = _w4472_ ;
	assign \g61546/_0_  = _w4473_ ;
	assign \g61547/_0_  = _w4477_ ;
	assign \g61548/_0_  = _w4481_ ;
	assign \g61549/_0_  = _w4488_ ;
	assign \g61550/_0_  = _w4489_ ;
	assign \g61551/_0_  = _w4490_ ;
	assign \g61552/_0_  = _w4496_ ;
	assign \g61553/_0_  = _w4506_ ;
	assign \g61554/_0_  = _w4525_ ;
	assign \g61555/_0_  = _w4528_ ;
	assign \g61556/_0_  = _w4531_ ;
	assign \g61557/_0_  = _w4540_ ;
	assign \g61558/_0_  = _w4541_ ;
	assign \g61559/_0_  = _w4542_ ;
	assign \g61560/_0_  = _w4546_ ;
	assign \g61561/_0_  = _w4550_ ;
	assign \g61562/_0_  = _w4557_ ;
	assign \g61563/_0_  = _w4558_ ;
	assign \g61564/_0_  = _w4559_ ;
	assign \g61565/_0_  = _w4560_ ;
	assign \g61566/_0_  = _w4561_ ;
	assign \g61620/_0_  = _w4564_ ;
	assign \g61621/_0_  = _w4567_ ;
	assign \g61622/_0_  = _w4569_ ;
	assign \g61623/_0_  = _w4571_ ;
	assign \g61753/_0_  = _w4573_ ;
	assign \g61764/_0_  = _w4575_ ;
	assign \g61786/_0_  = _w4577_ ;
	assign \g61795/_0_  = _w4579_ ;
	assign \g61801/_0_  = _w4586_ ;
	assign \g61803/_0_  = _w4587_ ;
	assign \g61808/_0_  = _w4588_ ;
	assign \g61848/_0_  = _w4591_ ;
	assign \g61850/_0_  = _w4594_ ;
	assign \g61851/_0_  = _w4596_ ;
	assign \g62097/_0_  = _w4602_ ;
	assign \g62102/_0_  = _w4604_ ;
	assign \g62115/_0_  = _w4609_ ;
	assign \g62119/_0_  = _w4253_ ;
	assign \g62130/_1_  = _w4404_ ;
	assign \g62131/_0_  = _w4614_ ;
	assign \g62132/_0_  = _w4619_ ;
	assign \g62139/_1_  = _w4427_ ;
	assign \g62140/_1_  = _w4368_ ;
	assign \g62141/_1_  = _w4374_ ;
	assign \g62144/_0_  = _w4628_ ;
	assign \g62145/_0_  = _w4629_ ;
	assign \g62146/_0_  = _w4633_ ;
	assign \g62147/_0_  = _w4634_ ;
	assign \g62150/_0_  = _w4639_ ;
	assign \g62151/_1_  = _w4381_ ;
	assign \g62152/_0_  = _w4645_ ;
	assign \g62153/_1_  = _w4400_ ;
	assign \g62156/_1_  = _w4377_ ;
	assign \g62157/_0_  = _w4273_ ;
	assign \g62159/_0_  = _w4303_ ;
	assign \g62161/_0_  = _w4654_ ;
	assign \g62187/_1_  = _w4439_ ;
	assign \g62190/_1_  = _w4444_ ;
	assign \g62191/_1_  = _w4421_ ;
	assign \g62192/_1_  = _w4447_ ;
	assign \g62194/_1_  = _w4455_ ;
	assign \g62195/_1_  = _w4476_ ;
	assign \g62196/_1_  = _w4480_ ;
	assign \g62203/_0_  = _w4323_ ;
	assign \g62204/_1_  = _w4430_ ;
	assign \g62207/_0__syn_2  = _w4503_ ;
	assign \g62208/_1_  = _w4509_ ;
	assign \g62209/_1_  = _w4527_ ;
	assign \g62210/_1_  = _w4530_ ;
	assign \g62211/_1_  = _w4545_ ;
	assign \g62212/_1_  = _w4549_ ;
	assign \g62217/_0_  = _w4657_ ;
	assign \g62286/_0_  = _w4669_ ;
	assign \g62287/_0_  = _w4670_ ;
	assign \g62288/_0_  = _w4672_ ;
	assign \g62289/_0_  = _w4674_ ;
	assign \g62290/_0_  = _w4675_ ;
	assign \g62291/_0_  = _w4676_ ;
	assign \g62292/_0_  = _w4677_ ;
	assign \g62435/_0_  = _w4678_ ;
	assign \g62436/_0_  = _w4679_ ;
	assign \g62439/_0_  = _w4681_ ;
	assign \g62456/_0_  = _w4685_ ;
	assign \g62486/_1_  = _w4331_ ;
	assign \g62492/_1_  = _w4352_ ;
	assign \g62494/_0_  = _w4690_ ;
	assign \g62495/_1_  = _w4357_ ;
	assign \g62497/_0_  = _w4693_ ;
	assign \g62537/_0_  = _w4696_ ;
	assign \g62544/_0_  = _w4697_ ;
	assign \g62546/_0_  = _w4698_ ;
	assign \g62547/_0_  = _w4699_ ;
	assign \g62549/_3_  = _w4700_ ;
	assign \g62552/_0_  = _w4701_ ;
	assign \g62554/_0_  = _w4706_ ;
	assign \g62555/_0_  = _w4707_ ;
	assign \g62556/_0_  = _w4712_ ;
	assign \g62558/_0_  = _w4717_ ;
	assign \g62559/_0_  = _w4718_ ;
	assign \g62561/_0_  = _w4723_ ;
	assign \g62562/_0_  = _w4724_ ;
	assign \g62566/_0_  = _w4725_ ;
	assign \g62567/_0_  = _w4726_ ;
	assign \g62568/_0_  = _w4727_ ;
	assign \g62569/_0_  = _w4728_ ;
	assign \g62570/_0_  = _w4729_ ;
	assign \g62571/_0_  = _w4730_ ;
	assign \g62572/_0_  = _w4731_ ;
	assign \g62573/_0_  = _w4732_ ;
	assign \g62574/_0_  = _w4733_ ;
	assign \g62575/_0_  = _w4734_ ;
	assign \g62576/_0_  = _w4735_ ;
	assign \g62577/_0_  = _w4736_ ;
	assign \g62578/_0_  = _w4737_ ;
	assign \g62579/_0_  = _w4738_ ;
	assign \g62580/_0_  = _w4739_ ;
	assign \g62581/_0_  = _w4740_ ;
	assign \g62582/_0_  = _w4741_ ;
	assign \g62583/_0_  = _w4742_ ;
	assign \g62584/_0_  = _w4743_ ;
	assign \g62585/_0_  = _w4744_ ;
	assign \g62586/_0_  = _w4745_ ;
	assign \g62587/_0_  = _w4746_ ;
	assign \g62588/_0_  = _w4747_ ;
	assign \g62589/_0_  = _w4748_ ;
	assign \g62590/_0_  = _w4749_ ;
	assign \g62591/_0_  = _w4750_ ;
	assign \g62592/_0_  = _w4751_ ;
	assign \g62593/_0_  = _w4752_ ;
	assign \g62594/_0_  = _w4753_ ;
	assign \g62595/_0_  = _w4754_ ;
	assign \g62596/_0_  = _w4755_ ;
	assign \g62597/_0_  = _w4756_ ;
	assign \g62602/_0_  = _w4757_ ;
	assign \g62607/_0_  = _w4758_ ;
	assign \g62608/_0_  = _w4759_ ;
	assign \g62609/_0_  = _w4760_ ;
	assign \g62619/_0_  = _w4761_ ;
	assign \g62620/_0_  = _w4762_ ;
	assign \g62621/_0_  = _w4763_ ;
	assign \g62622/_0_  = _w4764_ ;
	assign \g62623/_0_  = _w4765_ ;
	assign \g62624/_0_  = _w4766_ ;
	assign \g62626/_0_  = _w4767_ ;
	assign \g62627/_0_  = _w4768_ ;
	assign \g62628/_0_  = _w4769_ ;
	assign \g62629/_0_  = _w4770_ ;
	assign \g62630/_0_  = _w4771_ ;
	assign \g62631/_0_  = _w4772_ ;
	assign \g62632/_0_  = _w4773_ ;
	assign \g62633/_0_  = _w4774_ ;
	assign \g62634/_0_  = _w4775_ ;
	assign \g62635/_0_  = _w4776_ ;
	assign \g62636/_0_  = _w4777_ ;
	assign \g62637/_0_  = _w4778_ ;
	assign \g62638/_0_  = _w4779_ ;
	assign \g62639/_0_  = _w4780_ ;
	assign \g62640/_0_  = _w4781_ ;
	assign \g62641/_0_  = _w4782_ ;
	assign \g62642/_0_  = _w4783_ ;
	assign \g62643/_0_  = _w4784_ ;
	assign \g62644/_0_  = _w4785_ ;
	assign \g62645/_0_  = _w4786_ ;
	assign \g62646/_0_  = _w4787_ ;
	assign \g62647/_0_  = _w4788_ ;
	assign \g62648/_0_  = _w4789_ ;
	assign \g62649/_0_  = _w4790_ ;
	assign \g62650/_0_  = _w4791_ ;
	assign \g62651/_0_  = _w4792_ ;
	assign \g62652/_0_  = _w4793_ ;
	assign \g62653/_0_  = _w4794_ ;
	assign \g62654/_0_  = _w4795_ ;
	assign \g62655/_0_  = _w4796_ ;
	assign \g62656/_0_  = _w4797_ ;
	assign \g62657/_0_  = _w4798_ ;
	assign \g62658/_0_  = _w4799_ ;
	assign \g62659/_0_  = _w4800_ ;
	assign \g62660/_0_  = _w4801_ ;
	assign \g62661/_0_  = _w4802_ ;
	assign \g62674/_0_  = _w4803_ ;
	assign \g62682/_0_  = _w4804_ ;
	assign \g62683/_0_  = _w4805_ ;
	assign \g62689/_0_  = _w4809_ ;
	assign \g62690/_0_  = _w4813_ ;
	assign \g62691/_0_  = _w4817_ ;
	assign \g62694/_0_  = _w4821_ ;
	assign \g62695/_0_  = _w4825_ ;
	assign \g62696/_0_  = _w4829_ ;
	assign \g62698/_0_  = _w4833_ ;
	assign \g62699/_0_  = _w4837_ ;
	assign \g62700/_0_  = _w4841_ ;
	assign \g62723/_0_  = _w4844_ ;
	assign \g62724/_0_  = _w4847_ ;
	assign \g62725/_0_  = _w4850_ ;
	assign \g62726/_0_  = _w4853_ ;
	assign \g62727/_0_  = _w4856_ ;
	assign \g62728/_0_  = _w4859_ ;
	assign \g62735/_0_  = _w4862_ ;
	assign \g62736/_0_  = _w4865_ ;
	assign \g62737/_0_  = _w4868_ ;
	assign \g62738/_0_  = _w4871_ ;
	assign \g62739/_0_  = _w4874_ ;
	assign \g62740/_0_  = _w4877_ ;
	assign \g62754/_0_  = _w4878_ ;
	assign \g62762/_0_  = _w4879_ ;
	assign \g62763/_0_  = _w4880_ ;
	assign \g62764/_0_  = _w4881_ ;
	assign \g62780/_0_  = _w4882_ ;
	assign \g62781/_0_  = _w4883_ ;
	assign \g62785/_0_  = _w4884_ ;
	assign \g62786/_0_  = _w4885_ ;
	assign \g62787/_0_  = _w4886_ ;
	assign \g62791/_0_  = _w4887_ ;
	assign \g62792/_0_  = _w4888_ ;
	assign \g62794/_0_  = _w4889_ ;
	assign \g62804/_0_  = _w4891_ ;
	assign \g62806/_0_  = _w4893_ ;
	assign \g62807/_0_  = _w4895_ ;
	assign \g62811/_0_  = _w4897_ ;
	assign \g62968/_0_  = _w4898_ ;
	assign \g63005/_0_  = _w4900_ ;
	assign \g63041/_0_  = _w4901_ ;
	assign \g63116/_0_  = _w4905_ ;
	assign \g63157/_0_  = _w4908_ ;
	assign \g63164/_0_  = _w4909_ ;
	assign \g63170/_0_  = _w4912_ ;
	assign \g63189/_0_  = _w4913_ ;
	assign \g63202/_0_  = _w4914_ ;
	assign \g63206/_0_  = _w4915_ ;
	assign \g63207/_0_  = _w4919_ ;
	assign \g63265/_0_  = _w4920_ ;
	assign \g63266/_0_  = _w4921_ ;
	assign \g63269/_0_  = _w4922_ ;
	assign \g63271/_0_  = _w4923_ ;
	assign \g63272/_0_  = _w4924_ ;
	assign \g63273/_0_  = _w4925_ ;
	assign \g63274/_0_  = _w4926_ ;
	assign \g63275/_0_  = _w4927_ ;
	assign \g63276/_0_  = _w4928_ ;
	assign \g63277/_0_  = _w4929_ ;
	assign \g63278/_0_  = _w4930_ ;
	assign \g63280/_0_  = _w4931_ ;
	assign \g63281/_0_  = _w4932_ ;
	assign \g63282/_0_  = _w4933_ ;
	assign \g63283/_0_  = _w4934_ ;
	assign \g63284/_0_  = _w4935_ ;
	assign \g63285/_0_  = _w4936_ ;
	assign \g63286/_0_  = _w4937_ ;
	assign \g63287/_0_  = _w4938_ ;
	assign \g63288/_0_  = _w4939_ ;
	assign \g63289/_0_  = _w4940_ ;
	assign \g63290/_0_  = _w4941_ ;
	assign \g63292/_0_  = _w4942_ ;
	assign \g63293/_0_  = _w4943_ ;
	assign \g63294/_0_  = _w4944_ ;
	assign \g63295/_0_  = _w4945_ ;
	assign \g63296/_0_  = _w4946_ ;
	assign \g63297/_0_  = _w4947_ ;
	assign \g63298/_0_  = _w4948_ ;
	assign \g63299/_0_  = _w4949_ ;
	assign \g63302/_0_  = _w4950_ ;
	assign \g63303/_0_  = _w4951_ ;
	assign \g63304/_0_  = _w4952_ ;
	assign \g63305/_0_  = _w4953_ ;
	assign \g63306/_0_  = _w4954_ ;
	assign \g63307/_0_  = _w4955_ ;
	assign \g63308/_0_  = _w4956_ ;
	assign \g63309/_0_  = _w4957_ ;
	assign \g63310/_0_  = _w4958_ ;
	assign \g63311/_0_  = _w4959_ ;
	assign \g63312/_0_  = _w4960_ ;
	assign \g63313/_0_  = _w4961_ ;
	assign \g63314/_0_  = _w4962_ ;
	assign \g63315/_0_  = _w4963_ ;
	assign \g63316/_0_  = _w4964_ ;
	assign \g63317/_0_  = _w4965_ ;
	assign \g63318/_0_  = _w4966_ ;
	assign \g63319/_0_  = _w4967_ ;
	assign \g63320/_0_  = _w4968_ ;
	assign \g63321/_0_  = _w4969_ ;
	assign \g63322/_0_  = _w4970_ ;
	assign \g63323/_0_  = _w4971_ ;
	assign \g63324/_0_  = _w4972_ ;
	assign \g63325/_0_  = _w4973_ ;
	assign \g63326/_0_  = _w4974_ ;
	assign \g63327/_0_  = _w4975_ ;
	assign \g63328/_0_  = _w4976_ ;
	assign \g63329/_0_  = _w4977_ ;
	assign \g63330/_0_  = _w4978_ ;
	assign \g63331/_0_  = _w4979_ ;
	assign \g63339/_0_  = _w4983_ ;
	assign \g63505/_0_  = _w4985_ ;
	assign \g63525/_0_  = _w4075_ ;
	assign \g63543/_1_  = _w3452_ ;
	assign \g63602/_0_  = _w4988_ ;
	assign \g63653/_0_  = _w3459_ ;
	assign \g63663/_1_  = _w3472_ ;
	assign \g63677/_0_  = _w4162_ ;
	assign \g63694/_0_  = _w4199_ ;
	assign \g63729/_0_  = _w4990_ ;
	assign \g63766/_0_  = _w4995_ ;
	assign \g63771/_1_  = _w3875_ ;
	assign \g63773/_1_  = _w3881_ ;
	assign \g63784/_1_  = _w3879_ ;
	assign \g63964/_0_  = _w5000_ ;
	assign \g63965/_0_  = _w5005_ ;
	assign \g63966/_0_  = _w5006_ ;
	assign \g63967/_0_  = _w5007_ ;
	assign \g64257/_1_  = _w1920_ ;
	assign \g64266/_0_  = _w5012_ ;
	assign \g64275/_0_  = _w5014_ ;
	assign \g64400/_0_  = _w3890_ ;
	assign \g64416/_0_  = _w4108_ ;
	assign \g64470/_3_  = _w5016_ ;
	assign \g64473/_0_  = _w5019_ ;
	assign \g64474/_0_  = _w5022_ ;
	assign \g64475/_0_  = _w5025_ ;
	assign \g64479/_0_  = _w5030_ ;
	assign \g64480/_0_  = _w5033_ ;
	assign \g64481/_0_  = _w5036_ ;
	assign \g64483/_0_  = _w5039_ ;
	assign \g64484/_0_  = _w5041_ ;
	assign \g64485/_0_  = _w5042_ ;
	assign \g64486/_0_  = _w5043_ ;
	assign \g64493/_0_  = _w5046_ ;
	assign \g64494/_0_  = _w5049_ ;
	assign \g64495/_0_  = _w5052_ ;
	assign \g64496/_0_  = _w5055_ ;
	assign \g64505/_3_  = _w5056_ ;
	assign \g64507/_0_  = _w5059_ ;
	assign \g64508/_0_  = _w5062_ ;
	assign \g64510/_0_  = _w5065_ ;
	assign \g64511/_0_  = _w5068_ ;
	assign \g64544/_0_  = _w5069_ ;
	assign \g64545/_0_  = _w5070_ ;
	assign \g64546/_0_  = _w5071_ ;
	assign \g64639/_0_  = _w5073_ ;
	assign \g64641/_0_  = _w5075_ ;
	assign \g64642/_0_  = _w5077_ ;
	assign \g64645/_0_  = _w5079_ ;
	assign \g64650/_0_  = _w5081_ ;
	assign \g64737/_0_  = _w5082_ ;
	assign \g64738/_0_  = _w5084_ ;
	assign \g65066/_0_  = _w3841_ ;
	assign \g65070/_0_  = _w2865_ ;
	assign \g65090/_0_  = _w1574_ ;
	assign \g65102/_0_  = _w3926_ ;
	assign \g65102/_3_  = _w3927_ ;
	assign \g65126/_3_  = _w4245_ ;
	assign \g65147/_3_  = _w4264_ ;
	assign \g65163/_0_  = _w3751_ ;
	assign \g65176/_3_  = _w4296_ ;
	assign \g65178/_0_  = _w3374_ ;
	assign \g65182/_0_  = _w3728_ ;
	assign \g65190/_1_  = _w1578_ ;
	assign \g65191/_0_  = _w3299_ ;
	assign \g65196/_0_  = _w3262_ ;
	assign \g65268/_0_  = _w1459_ ;
	assign \g65275/_0_  = _w2208_ ;
	assign \g65290/_0_  = _w3962_ ;
	assign \g65290/_3_  = _w3963_ ;
	assign \g65291/_0_  = _w2212_ ;
	assign \g65292/_0_  = _w2861_ ;
	assign \g65298/_0_  = _w3944_ ;
	assign \g65298/_3_  = _w3945_ ;
	assign \g65314/_0_  = _w3979_ ;
	assign \g65314/_3_  = _w3980_ ;
	assign \g65319/_3_  = _w4314_ ;
	assign \g65335/_0_  = _w3811_ ;
	assign \g65342/_0_  = _w1419_ ;
	assign \g65348/_0_  = _w3395_ ;
	assign \g65422/_0_  = _w5086_ ;
	assign \g65465/_1_  = _w5032_ ;
	assign \g65469/_1_  = _w5035_ ;
	assign \g65478/_1_  = _w5028_ ;
	assign \g65507/_0_  = _w3316_ ;
	assign \g65548/_0_  = _w3933_ ;
	assign \g65699/_1_  = _w1294_ ;
	assign \g65713/_1_  = _w2013_ ;
	assign \g65835/_0_  = _w5087_ ;
	assign \g65860/_0_  = _w5089_ ;
	assign \g65863/_0_  = _w5090_ ;
	assign \g66094/_1_  = _w3951_ ;
	assign \g66102/_0_  = _w5093_ ;
	assign \g66107/_0_  = _w5094_ ;
	assign \g66130/_3_  = _w5095_ ;
	assign \g66131/_3_  = _w5096_ ;
	assign \g66228/_1_  = _w4671_ ;
	assign \g66348/_1_  = _w1400_ ;
	assign \g66543/_0_  = _w5097_ ;
	assign \g66549/_1_  = _w3986_ ;
	assign \g66640/_3_  = _w5098_ ;
	assign \g66641/_3_  = _w5099_ ;
	assign \g66950/_1_  = _w3914_ ;
	assign \g67111/_0_  = _w5100_ ;
	assign \g67219/_0_  = _w5101_ ;
	assign \g67263/_0_  = _w5102_ ;
	assign \g67909/_1_  = _w4673_ ;
	assign \g68049/_0_  = _w5103_ ;
	assign \g68220/_0_  = _w1137_ ;
	assign \g68413/_0_  = _w1135_ ;
	assign \g68511/_0_  = _w1245_ ;
	assign \g68536/_0_  = _w1130_ ;
	assign \g68543/_1_  = _w1397_ ;
	assign \g68554/_0_  = _w5104_ ;
	assign \g68559/_0_  = _w5105_ ;
	assign \g70915/_0_  = _w5114_ ;
	assign \g71108/_1_  = _w2166_ ;
	assign \g71115/_2_  = _w5115_ ;
	assign \g71244_dup/_0_  = _w2070_ ;
	assign \g71368/_0_  = _w5122_ ;
	assign \g71581/_0_  = _w5127_ ;
	assign \g71720/_0_  = _w1269_ ;
	assign \g785_reg/P0001  = _w1126_ ;
	assign \g789_reg/P0001  = _w1128_ ;
	assign \g797_reg/P0001  = _w1133_ ;
	assign \g809_reg/P0001  = _w1139_ ;
	assign \g813_reg/P0001  = _w1141_ ;
	assign \g966_reg/P0001  = _w1231_ ;
	assign \g968_reg/P0001  = _w1233_ ;
	assign \g970_reg/P0001  = _w1235_ ;
	assign \g972_reg/P0001  = _w1237_ ;
	assign \g974_reg/P0001  = _w1239_ ;
	assign \g976_reg/P0001  = _w1241_ ;
	assign \g978_reg/P0001  = _w1243_ ;
endmodule;