module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , s_pad , t_pad , u_pad , v_pad , w_pad , x_pad , y_pad , z_pad , \a0_pad  , \b0_pad  , \c0_pad  , \d0_pad  , \e0_pad  , \f0_pad  , \g0_pad  , \h0_pad  );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input s_pad ;
  input t_pad ;
  input u_pad ;
  input v_pad ;
  input w_pad ;
  input x_pad ;
  input y_pad ;
  input z_pad ;
  output \a0_pad  ;
  output \b0_pad  ;
  output \c0_pad  ;
  output \d0_pad  ;
  output \e0_pad  ;
  output \f0_pad  ;
  output \g0_pad  ;
  output \h0_pad  ;
  wire n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 ;
  assign n18 = ~a_pad & i_pad ;
  assign n19 = ~i_pad & ~s_pad ;
  assign n20 = ~n18 & ~n19 ;
  assign n21 = ~b_pad & i_pad ;
  assign n22 = ~i_pad & ~t_pad ;
  assign n23 = ~n21 & ~n22 ;
  assign n24 = ~c_pad & i_pad ;
  assign n25 = ~i_pad & ~u_pad ;
  assign n26 = ~n24 & ~n25 ;
  assign n27 = ~d_pad & i_pad ;
  assign n28 = ~i_pad & ~v_pad ;
  assign n29 = ~n27 & ~n28 ;
  assign n30 = ~e_pad & i_pad ;
  assign n31 = ~i_pad & ~w_pad ;
  assign n32 = ~n30 & ~n31 ;
  assign n33 = ~f_pad & i_pad ;
  assign n34 = ~i_pad & ~x_pad ;
  assign n35 = ~n33 & ~n34 ;
  assign n36 = ~g_pad & i_pad ;
  assign n37 = ~i_pad & ~y_pad ;
  assign n38 = ~n36 & ~n37 ;
  assign n39 = ~h_pad & i_pad ;
  assign n40 = ~i_pad & ~z_pad ;
  assign n41 = ~n39 & ~n40 ;
  assign \a0_pad  = n20 ;
  assign \b0_pad  = n23 ;
  assign \c0_pad  = n26 ;
  assign \d0_pad  = n29 ;
  assign \e0_pad  = n32 ;
  assign \f0_pad  = n35 ;
  assign \g0_pad  = n38 ;
  assign \h0_pad  = n41 ;
endmodule
