module top (\a[0] , \a[1] , \a[2] , \a[3] , \a[4] , \a[5] , \a[6] , \a[7] , \a[8] , \a[9] , \a[10] , \a[11] , \a[12] , \a[13] , \a[14] , \a[15] , \a[16] , \a[17] , \a[18] , \a[19] , \a[20] , \a[21] , \a[22] , \a[23] , \a[24] , \a[25] , \a[26] , \a[27] , \a[28] , \a[29] , \a[30] , \a[31] , \a[32] , \a[33] , \a[34] , \a[35] , \a[36] , \a[37] , \a[38] , \a[39] , \a[40] , \a[41] , \a[42] , \a[43] , \a[44] , \a[45] , \a[46] , \a[47] , \a[48] , \a[49] , \a[50] , \a[51] , \a[52] , \a[53] , \a[54] , \a[55] , \a[56] , \a[57] , \a[58] , \a[59] , \a[60] , \a[61] , \a[62] , \a[63] , \a[64] , \a[65] , \a[66] , \a[67] , \a[68] , \a[69] , \a[70] , \a[71] , \a[72] , \a[73] , \a[74] , \a[75] , \a[76] , \a[77] , \a[78] , \a[79] , \a[80] , \a[81] , \a[82] , \a[83] , \a[84] , \a[85] , \a[86] , \a[87] , \a[88] , \a[89] , \a[90] , \a[91] , \a[92] , \a[93] , \a[94] , \a[95] , \a[96] , \a[97] , \a[98] , \a[99] , \a[100] , \a[101] , \a[102] , \a[103] , \a[104] , \a[105] , \a[106] , \a[107] , \a[108] , \a[109] , \a[110] , \a[111] , \a[112] , \a[113] , \a[114] , \a[115] , \a[116] , \a[117] , \a[118] , \a[119] , \a[120] , \a[121] , \a[122] , \a[123] , \a[124] , \a[125] , \a[126] , \a[127] , \b[0] , \b[1] , \b[2] , \b[3] , \b[4] , \b[5] , \b[6] , \b[7] , \b[8] , \b[9] , \b[10] , \b[11] , \b[12] , \b[13] , \b[14] , \b[15] , \b[16] , \b[17] , \b[18] , \b[19] , \b[20] , \b[21] , \b[22] , \b[23] , \b[24] , \b[25] , \b[26] , \b[27] , \b[28] , \b[29] , \b[30] , \b[31] , \b[32] , \b[33] , \b[34] , \b[35] , \b[36] , \b[37] , \b[38] , \b[39] , \b[40] , \b[41] , \b[42] , \b[43] , \b[44] , \b[45] , \b[46] , \b[47] , \b[48] , \b[49] , \b[50] , \b[51] , \b[52] , \b[53] , \b[54] , \b[55] , \b[56] , \b[57] , \b[58] , \b[59] , \b[60] , \b[61] , \b[62] , \b[63] , \b[64] , \b[65] , \b[66] , \b[67] , \b[68] , \b[69] , \b[70] , \b[71] , \b[72] , \b[73] , \b[74] , \b[75] , \b[76] , \b[77] , \b[78] , \b[79] , \b[80] , \b[81] , \b[82] , \b[83] , \b[84] , \b[85] , \b[86] , \b[87] , \b[88] , \b[89] , \b[90] , \b[91] , \b[92] , \b[93] , \b[94] , \b[95] , \b[96] , \b[97] , \b[98] , \b[99] , \b[100] , \b[101] , \b[102] , \b[103] , \b[104] , \b[105] , \b[106] , \b[107] , \b[108] , \b[109] , \b[110] , \b[111] , \b[112] , \b[113] , \b[114] , \b[115] , \b[116] , \b[117] , \b[118] , \b[119] , \b[120] , \b[121] , \b[122] , \b[123] , \b[124] , \b[125] , \b[126] , \b[127] , \f[0] , \f[1] , \f[2] , \f[3] , \f[4] , \f[5] , \f[6] , \f[7] , \f[8] , \f[9] , \f[10] , \f[11] , \f[12] , \f[13] , \f[14] , \f[15] , \f[16] , \f[17] , \f[18] , \f[19] , \f[20] , \f[21] , \f[22] , \f[23] , \f[24] , \f[25] , \f[26] , \f[27] , \f[28] , \f[29] , \f[30] , \f[31] , \f[32] , \f[33] , \f[34] , \f[35] , \f[36] , \f[37] , \f[38] , \f[39] , \f[40] , \f[41] , \f[42] , \f[43] , \f[44] , \f[45] , \f[46] , \f[47] , \f[48] , \f[49] , \f[50] , \f[51] , \f[52] , \f[53] , \f[54] , \f[55] , \f[56] , \f[57] , \f[58] , \f[59] , \f[60] , \f[61] , \f[62] , \f[63] , \f[64] , \f[65] , \f[66] , \f[67] , \f[68] , \f[69] , \f[70] , \f[71] , \f[72] , \f[73] , \f[74] , \f[75] , \f[76] , \f[77] , \f[78] , \f[79] , \f[80] , \f[81] , \f[82] , \f[83] , \f[84] , \f[85] , \f[86] , \f[87] , \f[88] , \f[89] , \f[90] , \f[91] , \f[92] , \f[93] , \f[94] , \f[95] , \f[96] , \f[97] , \f[98] , \f[99] , \f[100] , \f[101] , \f[102] , \f[103] , \f[104] , \f[105] , \f[106] , \f[107] , \f[108] , \f[109] , \f[110] , \f[111] , \f[112] , \f[113] , \f[114] , \f[115] , \f[116] , \f[117] , \f[118] , \f[119] , \f[120] , \f[121] , \f[122] , \f[123] , \f[124] , \f[125] , \f[126] , \f[127] , cOut);
	input \a[0]  ;
	input \a[1]  ;
	input \a[2]  ;
	input \a[3]  ;
	input \a[4]  ;
	input \a[5]  ;
	input \a[6]  ;
	input \a[7]  ;
	input \a[8]  ;
	input \a[9]  ;
	input \a[10]  ;
	input \a[11]  ;
	input \a[12]  ;
	input \a[13]  ;
	input \a[14]  ;
	input \a[15]  ;
	input \a[16]  ;
	input \a[17]  ;
	input \a[18]  ;
	input \a[19]  ;
	input \a[20]  ;
	input \a[21]  ;
	input \a[22]  ;
	input \a[23]  ;
	input \a[24]  ;
	input \a[25]  ;
	input \a[26]  ;
	input \a[27]  ;
	input \a[28]  ;
	input \a[29]  ;
	input \a[30]  ;
	input \a[31]  ;
	input \a[32]  ;
	input \a[33]  ;
	input \a[34]  ;
	input \a[35]  ;
	input \a[36]  ;
	input \a[37]  ;
	input \a[38]  ;
	input \a[39]  ;
	input \a[40]  ;
	input \a[41]  ;
	input \a[42]  ;
	input \a[43]  ;
	input \a[44]  ;
	input \a[45]  ;
	input \a[46]  ;
	input \a[47]  ;
	input \a[48]  ;
	input \a[49]  ;
	input \a[50]  ;
	input \a[51]  ;
	input \a[52]  ;
	input \a[53]  ;
	input \a[54]  ;
	input \a[55]  ;
	input \a[56]  ;
	input \a[57]  ;
	input \a[58]  ;
	input \a[59]  ;
	input \a[60]  ;
	input \a[61]  ;
	input \a[62]  ;
	input \a[63]  ;
	input \a[64]  ;
	input \a[65]  ;
	input \a[66]  ;
	input \a[67]  ;
	input \a[68]  ;
	input \a[69]  ;
	input \a[70]  ;
	input \a[71]  ;
	input \a[72]  ;
	input \a[73]  ;
	input \a[74]  ;
	input \a[75]  ;
	input \a[76]  ;
	input \a[77]  ;
	input \a[78]  ;
	input \a[79]  ;
	input \a[80]  ;
	input \a[81]  ;
	input \a[82]  ;
	input \a[83]  ;
	input \a[84]  ;
	input \a[85]  ;
	input \a[86]  ;
	input \a[87]  ;
	input \a[88]  ;
	input \a[89]  ;
	input \a[90]  ;
	input \a[91]  ;
	input \a[92]  ;
	input \a[93]  ;
	input \a[94]  ;
	input \a[95]  ;
	input \a[96]  ;
	input \a[97]  ;
	input \a[98]  ;
	input \a[99]  ;
	input \a[100]  ;
	input \a[101]  ;
	input \a[102]  ;
	input \a[103]  ;
	input \a[104]  ;
	input \a[105]  ;
	input \a[106]  ;
	input \a[107]  ;
	input \a[108]  ;
	input \a[109]  ;
	input \a[110]  ;
	input \a[111]  ;
	input \a[112]  ;
	input \a[113]  ;
	input \a[114]  ;
	input \a[115]  ;
	input \a[116]  ;
	input \a[117]  ;
	input \a[118]  ;
	input \a[119]  ;
	input \a[120]  ;
	input \a[121]  ;
	input \a[122]  ;
	input \a[123]  ;
	input \a[124]  ;
	input \a[125]  ;
	input \a[126]  ;
	input \a[127]  ;
	input \b[0]  ;
	input \b[1]  ;
	input \b[2]  ;
	input \b[3]  ;
	input \b[4]  ;
	input \b[5]  ;
	input \b[6]  ;
	input \b[7]  ;
	input \b[8]  ;
	input \b[9]  ;
	input \b[10]  ;
	input \b[11]  ;
	input \b[12]  ;
	input \b[13]  ;
	input \b[14]  ;
	input \b[15]  ;
	input \b[16]  ;
	input \b[17]  ;
	input \b[18]  ;
	input \b[19]  ;
	input \b[20]  ;
	input \b[21]  ;
	input \b[22]  ;
	input \b[23]  ;
	input \b[24]  ;
	input \b[25]  ;
	input \b[26]  ;
	input \b[27]  ;
	input \b[28]  ;
	input \b[29]  ;
	input \b[30]  ;
	input \b[31]  ;
	input \b[32]  ;
	input \b[33]  ;
	input \b[34]  ;
	input \b[35]  ;
	input \b[36]  ;
	input \b[37]  ;
	input \b[38]  ;
	input \b[39]  ;
	input \b[40]  ;
	input \b[41]  ;
	input \b[42]  ;
	input \b[43]  ;
	input \b[44]  ;
	input \b[45]  ;
	input \b[46]  ;
	input \b[47]  ;
	input \b[48]  ;
	input \b[49]  ;
	input \b[50]  ;
	input \b[51]  ;
	input \b[52]  ;
	input \b[53]  ;
	input \b[54]  ;
	input \b[55]  ;
	input \b[56]  ;
	input \b[57]  ;
	input \b[58]  ;
	input \b[59]  ;
	input \b[60]  ;
	input \b[61]  ;
	input \b[62]  ;
	input \b[63]  ;
	input \b[64]  ;
	input \b[65]  ;
	input \b[66]  ;
	input \b[67]  ;
	input \b[68]  ;
	input \b[69]  ;
	input \b[70]  ;
	input \b[71]  ;
	input \b[72]  ;
	input \b[73]  ;
	input \b[74]  ;
	input \b[75]  ;
	input \b[76]  ;
	input \b[77]  ;
	input \b[78]  ;
	input \b[79]  ;
	input \b[80]  ;
	input \b[81]  ;
	input \b[82]  ;
	input \b[83]  ;
	input \b[84]  ;
	input \b[85]  ;
	input \b[86]  ;
	input \b[87]  ;
	input \b[88]  ;
	input \b[89]  ;
	input \b[90]  ;
	input \b[91]  ;
	input \b[92]  ;
	input \b[93]  ;
	input \b[94]  ;
	input \b[95]  ;
	input \b[96]  ;
	input \b[97]  ;
	input \b[98]  ;
	input \b[99]  ;
	input \b[100]  ;
	input \b[101]  ;
	input \b[102]  ;
	input \b[103]  ;
	input \b[104]  ;
	input \b[105]  ;
	input \b[106]  ;
	input \b[107]  ;
	input \b[108]  ;
	input \b[109]  ;
	input \b[110]  ;
	input \b[111]  ;
	input \b[112]  ;
	input \b[113]  ;
	input \b[114]  ;
	input \b[115]  ;
	input \b[116]  ;
	input \b[117]  ;
	input \b[118]  ;
	input \b[119]  ;
	input \b[120]  ;
	input \b[121]  ;
	input \b[122]  ;
	input \b[123]  ;
	input \b[124]  ;
	input \b[125]  ;
	input \b[126]  ;
	input \b[127]  ;
	output \f[0]  ;
	output \f[1]  ;
	output \f[2]  ;
	output \f[3]  ;
	output \f[4]  ;
	output \f[5]  ;
	output \f[6]  ;
	output \f[7]  ;
	output \f[8]  ;
	output \f[9]  ;
	output \f[10]  ;
	output \f[11]  ;
	output \f[12]  ;
	output \f[13]  ;
	output \f[14]  ;
	output \f[15]  ;
	output \f[16]  ;
	output \f[17]  ;
	output \f[18]  ;
	output \f[19]  ;
	output \f[20]  ;
	output \f[21]  ;
	output \f[22]  ;
	output \f[23]  ;
	output \f[24]  ;
	output \f[25]  ;
	output \f[26]  ;
	output \f[27]  ;
	output \f[28]  ;
	output \f[29]  ;
	output \f[30]  ;
	output \f[31]  ;
	output \f[32]  ;
	output \f[33]  ;
	output \f[34]  ;
	output \f[35]  ;
	output \f[36]  ;
	output \f[37]  ;
	output \f[38]  ;
	output \f[39]  ;
	output \f[40]  ;
	output \f[41]  ;
	output \f[42]  ;
	output \f[43]  ;
	output \f[44]  ;
	output \f[45]  ;
	output \f[46]  ;
	output \f[47]  ;
	output \f[48]  ;
	output \f[49]  ;
	output \f[50]  ;
	output \f[51]  ;
	output \f[52]  ;
	output \f[53]  ;
	output \f[54]  ;
	output \f[55]  ;
	output \f[56]  ;
	output \f[57]  ;
	output \f[58]  ;
	output \f[59]  ;
	output \f[60]  ;
	output \f[61]  ;
	output \f[62]  ;
	output \f[63]  ;
	output \f[64]  ;
	output \f[65]  ;
	output \f[66]  ;
	output \f[67]  ;
	output \f[68]  ;
	output \f[69]  ;
	output \f[70]  ;
	output \f[71]  ;
	output \f[72]  ;
	output \f[73]  ;
	output \f[74]  ;
	output \f[75]  ;
	output \f[76]  ;
	output \f[77]  ;
	output \f[78]  ;
	output \f[79]  ;
	output \f[80]  ;
	output \f[81]  ;
	output \f[82]  ;
	output \f[83]  ;
	output \f[84]  ;
	output \f[85]  ;
	output \f[86]  ;
	output \f[87]  ;
	output \f[88]  ;
	output \f[89]  ;
	output \f[90]  ;
	output \f[91]  ;
	output \f[92]  ;
	output \f[93]  ;
	output \f[94]  ;
	output \f[95]  ;
	output \f[96]  ;
	output \f[97]  ;
	output \f[98]  ;
	output \f[99]  ;
	output \f[100]  ;
	output \f[101]  ;
	output \f[102]  ;
	output \f[103]  ;
	output \f[104]  ;
	output \f[105]  ;
	output \f[106]  ;
	output \f[107]  ;
	output \f[108]  ;
	output \f[109]  ;
	output \f[110]  ;
	output \f[111]  ;
	output \f[112]  ;
	output \f[113]  ;
	output \f[114]  ;
	output \f[115]  ;
	output \f[116]  ;
	output \f[117]  ;
	output \f[118]  ;
	output \f[119]  ;
	output \f[120]  ;
	output \f[121]  ;
	output \f[122]  ;
	output \f[123]  ;
	output \f[124]  ;
	output \f[125]  ;
	output \f[126]  ;
	output \f[127]  ;
	output cOut ;
	wire _w1275_ ;
	wire _w1274_ ;
	wire _w1273_ ;
	wire _w1272_ ;
	wire _w1271_ ;
	wire _w1270_ ;
	wire _w1269_ ;
	wire _w1268_ ;
	wire _w1267_ ;
	wire _w1266_ ;
	wire _w1265_ ;
	wire _w1264_ ;
	wire _w1263_ ;
	wire _w1262_ ;
	wire _w1261_ ;
	wire _w1260_ ;
	wire _w1259_ ;
	wire _w1258_ ;
	wire _w1257_ ;
	wire _w1256_ ;
	wire _w1255_ ;
	wire _w1254_ ;
	wire _w1253_ ;
	wire _w1252_ ;
	wire _w1251_ ;
	wire _w1250_ ;
	wire _w1249_ ;
	wire _w1248_ ;
	wire _w1247_ ;
	wire _w1246_ ;
	wire _w1245_ ;
	wire _w1244_ ;
	wire _w1243_ ;
	wire _w1242_ ;
	wire _w1241_ ;
	wire _w1240_ ;
	wire _w1239_ ;
	wire _w1238_ ;
	wire _w1237_ ;
	wire _w1236_ ;
	wire _w1235_ ;
	wire _w1234_ ;
	wire _w1233_ ;
	wire _w1232_ ;
	wire _w1231_ ;
	wire _w1230_ ;
	wire _w1229_ ;
	wire _w1228_ ;
	wire _w1227_ ;
	wire _w1226_ ;
	wire _w1225_ ;
	wire _w1224_ ;
	wire _w1223_ ;
	wire _w1222_ ;
	wire _w1221_ ;
	wire _w1220_ ;
	wire _w1219_ ;
	wire _w1218_ ;
	wire _w1217_ ;
	wire _w1216_ ;
	wire _w1215_ ;
	wire _w1214_ ;
	wire _w1213_ ;
	wire _w1212_ ;
	wire _w1211_ ;
	wire _w1210_ ;
	wire _w1209_ ;
	wire _w1208_ ;
	wire _w1207_ ;
	wire _w1206_ ;
	wire _w1205_ ;
	wire _w1204_ ;
	wire _w1203_ ;
	wire _w1202_ ;
	wire _w1201_ ;
	wire _w1200_ ;
	wire _w1199_ ;
	wire _w1198_ ;
	wire _w1197_ ;
	wire _w1196_ ;
	wire _w1195_ ;
	wire _w1194_ ;
	wire _w1193_ ;
	wire _w1192_ ;
	wire _w1191_ ;
	wire _w1190_ ;
	wire _w1189_ ;
	wire _w1188_ ;
	wire _w1187_ ;
	wire _w1186_ ;
	wire _w1185_ ;
	wire _w1184_ ;
	wire _w1183_ ;
	wire _w1182_ ;
	wire _w1181_ ;
	wire _w1180_ ;
	wire _w1179_ ;
	wire _w1178_ ;
	wire _w1177_ ;
	wire _w1176_ ;
	wire _w1175_ ;
	wire _w1174_ ;
	wire _w1173_ ;
	wire _w1172_ ;
	wire _w1171_ ;
	wire _w1170_ ;
	wire _w1169_ ;
	wire _w1168_ ;
	wire _w1167_ ;
	wire _w1166_ ;
	wire _w1165_ ;
	wire _w1164_ ;
	wire _w1163_ ;
	wire _w1162_ ;
	wire _w1161_ ;
	wire _w1160_ ;
	wire _w1159_ ;
	wire _w1158_ ;
	wire _w1157_ ;
	wire _w1156_ ;
	wire _w1155_ ;
	wire _w1154_ ;
	wire _w1153_ ;
	wire _w1152_ ;
	wire _w1151_ ;
	wire _w1150_ ;
	wire _w1149_ ;
	wire _w1148_ ;
	wire _w1147_ ;
	wire _w1146_ ;
	wire _w1145_ ;
	wire _w1144_ ;
	wire _w1143_ ;
	wire _w1142_ ;
	wire _w1141_ ;
	wire _w1140_ ;
	wire _w1139_ ;
	wire _w1138_ ;
	wire _w1137_ ;
	wire _w1136_ ;
	wire _w1135_ ;
	wire _w1134_ ;
	wire _w1133_ ;
	wire _w1132_ ;
	wire _w1131_ ;
	wire _w1130_ ;
	wire _w1129_ ;
	wire _w1128_ ;
	wire _w1127_ ;
	wire _w1126_ ;
	wire _w1125_ ;
	wire _w1124_ ;
	wire _w1123_ ;
	wire _w1122_ ;
	wire _w1121_ ;
	wire _w1120_ ;
	wire _w1119_ ;
	wire _w1118_ ;
	wire _w1117_ ;
	wire _w1116_ ;
	wire _w1115_ ;
	wire _w1114_ ;
	wire _w1113_ ;
	wire _w1112_ ;
	wire _w1111_ ;
	wire _w1110_ ;
	wire _w1109_ ;
	wire _w1108_ ;
	wire _w1107_ ;
	wire _w1106_ ;
	wire _w1105_ ;
	wire _w1104_ ;
	wire _w1103_ ;
	wire _w1102_ ;
	wire _w1101_ ;
	wire _w1100_ ;
	wire _w1099_ ;
	wire _w1098_ ;
	wire _w1097_ ;
	wire _w1096_ ;
	wire _w1095_ ;
	wire _w1094_ ;
	wire _w1093_ ;
	wire _w1092_ ;
	wire _w1091_ ;
	wire _w1090_ ;
	wire _w1089_ ;
	wire _w1088_ ;
	wire _w1087_ ;
	wire _w1086_ ;
	wire _w1085_ ;
	wire _w1084_ ;
	wire _w1083_ ;
	wire _w1082_ ;
	wire _w1081_ ;
	wire _w1080_ ;
	wire _w1079_ ;
	wire _w1078_ ;
	wire _w1077_ ;
	wire _w1076_ ;
	wire _w1075_ ;
	wire _w1074_ ;
	wire _w1073_ ;
	wire _w1072_ ;
	wire _w1071_ ;
	wire _w1070_ ;
	wire _w1069_ ;
	wire _w1068_ ;
	wire _w1067_ ;
	wire _w1066_ ;
	wire _w1065_ ;
	wire _w1064_ ;
	wire _w1063_ ;
	wire _w1062_ ;
	wire _w1061_ ;
	wire _w1060_ ;
	wire _w1059_ ;
	wire _w1058_ ;
	wire _w1057_ ;
	wire _w1056_ ;
	wire _w1055_ ;
	wire _w1054_ ;
	wire _w1053_ ;
	wire _w1052_ ;
	wire _w1051_ ;
	wire _w1050_ ;
	wire _w1049_ ;
	wire _w1048_ ;
	wire _w1047_ ;
	wire _w1046_ ;
	wire _w1045_ ;
	wire _w1044_ ;
	wire _w1043_ ;
	wire _w1042_ ;
	wire _w1041_ ;
	wire _w1040_ ;
	wire _w1039_ ;
	wire _w1038_ ;
	wire _w1037_ ;
	wire _w1036_ ;
	wire _w1035_ ;
	wire _w1034_ ;
	wire _w1033_ ;
	wire _w1032_ ;
	wire _w1031_ ;
	wire _w1030_ ;
	wire _w1029_ ;
	wire _w1028_ ;
	wire _w1027_ ;
	wire _w1026_ ;
	wire _w1025_ ;
	wire _w1024_ ;
	wire _w1023_ ;
	wire _w1022_ ;
	wire _w1021_ ;
	wire _w1020_ ;
	wire _w1019_ ;
	wire _w1018_ ;
	wire _w1017_ ;
	wire _w1016_ ;
	wire _w1015_ ;
	wire _w1014_ ;
	wire _w1013_ ;
	wire _w1012_ ;
	wire _w1011_ ;
	wire _w1010_ ;
	wire _w1009_ ;
	wire _w1008_ ;
	wire _w1007_ ;
	wire _w1006_ ;
	wire _w1005_ ;
	wire _w1004_ ;
	wire _w1003_ ;
	wire _w1002_ ;
	wire _w1001_ ;
	wire _w1000_ ;
	wire _w999_ ;
	wire _w998_ ;
	wire _w997_ ;
	wire _w996_ ;
	wire _w995_ ;
	wire _w994_ ;
	wire _w993_ ;
	wire _w992_ ;
	wire _w991_ ;
	wire _w990_ ;
	wire _w989_ ;
	wire _w988_ ;
	wire _w987_ ;
	wire _w986_ ;
	wire _w985_ ;
	wire _w984_ ;
	wire _w983_ ;
	wire _w982_ ;
	wire _w981_ ;
	wire _w980_ ;
	wire _w979_ ;
	wire _w978_ ;
	wire _w977_ ;
	wire _w976_ ;
	wire _w975_ ;
	wire _w974_ ;
	wire _w973_ ;
	wire _w972_ ;
	wire _w971_ ;
	wire _w970_ ;
	wire _w969_ ;
	wire _w968_ ;
	wire _w967_ ;
	wire _w966_ ;
	wire _w965_ ;
	wire _w964_ ;
	wire _w963_ ;
	wire _w962_ ;
	wire _w961_ ;
	wire _w960_ ;
	wire _w959_ ;
	wire _w958_ ;
	wire _w957_ ;
	wire _w956_ ;
	wire _w955_ ;
	wire _w954_ ;
	wire _w953_ ;
	wire _w952_ ;
	wire _w951_ ;
	wire _w950_ ;
	wire _w949_ ;
	wire _w948_ ;
	wire _w947_ ;
	wire _w946_ ;
	wire _w945_ ;
	wire _w944_ ;
	wire _w943_ ;
	wire _w942_ ;
	wire _w941_ ;
	wire _w940_ ;
	wire _w939_ ;
	wire _w938_ ;
	wire _w937_ ;
	wire _w936_ ;
	wire _w935_ ;
	wire _w934_ ;
	wire _w933_ ;
	wire _w932_ ;
	wire _w931_ ;
	wire _w930_ ;
	wire _w929_ ;
	wire _w928_ ;
	wire _w927_ ;
	wire _w926_ ;
	wire _w925_ ;
	wire _w924_ ;
	wire _w923_ ;
	wire _w922_ ;
	wire _w921_ ;
	wire _w920_ ;
	wire _w919_ ;
	wire _w918_ ;
	wire _w917_ ;
	wire _w916_ ;
	wire _w915_ ;
	wire _w914_ ;
	wire _w913_ ;
	wire _w912_ ;
	wire _w911_ ;
	wire _w910_ ;
	wire _w909_ ;
	wire _w908_ ;
	wire _w907_ ;
	wire _w906_ ;
	wire _w905_ ;
	wire _w904_ ;
	wire _w903_ ;
	wire _w902_ ;
	wire _w901_ ;
	wire _w900_ ;
	wire _w899_ ;
	wire _w898_ ;
	wire _w897_ ;
	wire _w896_ ;
	wire _w895_ ;
	wire _w894_ ;
	wire _w893_ ;
	wire _w892_ ;
	wire _w891_ ;
	wire _w890_ ;
	wire _w889_ ;
	wire _w888_ ;
	wire _w887_ ;
	wire _w886_ ;
	wire _w885_ ;
	wire _w884_ ;
	wire _w883_ ;
	wire _w882_ ;
	wire _w881_ ;
	wire _w880_ ;
	wire _w879_ ;
	wire _w878_ ;
	wire _w877_ ;
	wire _w876_ ;
	wire _w875_ ;
	wire _w874_ ;
	wire _w873_ ;
	wire _w872_ ;
	wire _w871_ ;
	wire _w870_ ;
	wire _w869_ ;
	wire _w868_ ;
	wire _w867_ ;
	wire _w866_ ;
	wire _w865_ ;
	wire _w864_ ;
	wire _w863_ ;
	wire _w862_ ;
	wire _w861_ ;
	wire _w860_ ;
	wire _w859_ ;
	wire _w858_ ;
	wire _w857_ ;
	wire _w856_ ;
	wire _w855_ ;
	wire _w854_ ;
	wire _w853_ ;
	wire _w852_ ;
	wire _w851_ ;
	wire _w850_ ;
	wire _w849_ ;
	wire _w848_ ;
	wire _w847_ ;
	wire _w846_ ;
	wire _w845_ ;
	wire _w844_ ;
	wire _w843_ ;
	wire _w842_ ;
	wire _w841_ ;
	wire _w840_ ;
	wire _w839_ ;
	wire _w838_ ;
	wire _w837_ ;
	wire _w836_ ;
	wire _w835_ ;
	wire _w834_ ;
	wire _w833_ ;
	wire _w832_ ;
	wire _w831_ ;
	wire _w830_ ;
	wire _w829_ ;
	wire _w828_ ;
	wire _w827_ ;
	wire _w826_ ;
	wire _w825_ ;
	wire _w824_ ;
	wire _w823_ ;
	wire _w822_ ;
	wire _w821_ ;
	wire _w820_ ;
	wire _w819_ ;
	wire _w818_ ;
	wire _w817_ ;
	wire _w816_ ;
	wire _w815_ ;
	wire _w814_ ;
	wire _w813_ ;
	wire _w812_ ;
	wire _w811_ ;
	wire _w810_ ;
	wire _w809_ ;
	wire _w808_ ;
	wire _w807_ ;
	wire _w806_ ;
	wire _w805_ ;
	wire _w804_ ;
	wire _w803_ ;
	wire _w802_ ;
	wire _w801_ ;
	wire _w800_ ;
	wire _w799_ ;
	wire _w798_ ;
	wire _w513_ ;
	wire _w512_ ;
	wire _w511_ ;
	wire _w510_ ;
	wire _w509_ ;
	wire _w508_ ;
	wire _w507_ ;
	wire _w506_ ;
	wire _w505_ ;
	wire _w504_ ;
	wire _w503_ ;
	wire _w502_ ;
	wire _w501_ ;
	wire _w500_ ;
	wire _w499_ ;
	wire _w498_ ;
	wire _w497_ ;
	wire _w496_ ;
	wire _w495_ ;
	wire _w494_ ;
	wire _w493_ ;
	wire _w492_ ;
	wire _w491_ ;
	wire _w490_ ;
	wire _w489_ ;
	wire _w488_ ;
	wire _w487_ ;
	wire _w486_ ;
	wire _w485_ ;
	wire _w484_ ;
	wire _w483_ ;
	wire _w482_ ;
	wire _w481_ ;
	wire _w480_ ;
	wire _w479_ ;
	wire _w478_ ;
	wire _w477_ ;
	wire _w476_ ;
	wire _w475_ ;
	wire _w474_ ;
	wire _w473_ ;
	wire _w472_ ;
	wire _w471_ ;
	wire _w470_ ;
	wire _w469_ ;
	wire _w468_ ;
	wire _w467_ ;
	wire _w466_ ;
	wire _w465_ ;
	wire _w464_ ;
	wire _w463_ ;
	wire _w462_ ;
	wire _w461_ ;
	wire _w460_ ;
	wire _w459_ ;
	wire _w458_ ;
	wire _w457_ ;
	wire _w456_ ;
	wire _w455_ ;
	wire _w454_ ;
	wire _w453_ ;
	wire _w452_ ;
	wire _w451_ ;
	wire _w450_ ;
	wire _w449_ ;
	wire _w448_ ;
	wire _w447_ ;
	wire _w446_ ;
	wire _w445_ ;
	wire _w444_ ;
	wire _w443_ ;
	wire _w442_ ;
	wire _w441_ ;
	wire _w440_ ;
	wire _w439_ ;
	wire _w438_ ;
	wire _w437_ ;
	wire _w436_ ;
	wire _w435_ ;
	wire _w434_ ;
	wire _w433_ ;
	wire _w432_ ;
	wire _w431_ ;
	wire _w430_ ;
	wire _w429_ ;
	wire _w428_ ;
	wire _w427_ ;
	wire _w426_ ;
	wire _w425_ ;
	wire _w424_ ;
	wire _w423_ ;
	wire _w422_ ;
	wire _w421_ ;
	wire _w420_ ;
	wire _w419_ ;
	wire _w418_ ;
	wire _w417_ ;
	wire _w416_ ;
	wire _w415_ ;
	wire _w414_ ;
	wire _w413_ ;
	wire _w412_ ;
	wire _w411_ ;
	wire _w410_ ;
	wire _w409_ ;
	wire _w408_ ;
	wire _w407_ ;
	wire _w406_ ;
	wire _w405_ ;
	wire _w404_ ;
	wire _w403_ ;
	wire _w402_ ;
	wire _w401_ ;
	wire _w400_ ;
	wire _w399_ ;
	wire _w398_ ;
	wire _w397_ ;
	wire _w396_ ;
	wire _w395_ ;
	wire _w394_ ;
	wire _w393_ ;
	wire _w392_ ;
	wire _w391_ ;
	wire _w390_ ;
	wire _w389_ ;
	wire _w388_ ;
	wire _w387_ ;
	wire _w386_ ;
	wire _w385_ ;
	wire _w384_ ;
	wire _w315_ ;
	wire _w314_ ;
	wire _w313_ ;
	wire _w312_ ;
	wire _w311_ ;
	wire _w310_ ;
	wire _w309_ ;
	wire _w308_ ;
	wire _w307_ ;
	wire _w306_ ;
	wire _w305_ ;
	wire _w304_ ;
	wire _w303_ ;
	wire _w302_ ;
	wire _w301_ ;
	wire _w300_ ;
	wire _w299_ ;
	wire _w298_ ;
	wire _w297_ ;
	wire _w296_ ;
	wire _w295_ ;
	wire _w294_ ;
	wire _w293_ ;
	wire _w292_ ;
	wire _w291_ ;
	wire _w290_ ;
	wire _w289_ ;
	wire _w288_ ;
	wire _w287_ ;
	wire _w286_ ;
	wire _w269_ ;
	wire _w268_ ;
	wire _w267_ ;
	wire _w266_ ;
	wire _w265_ ;
	wire _w264_ ;
	wire _w263_ ;
	wire _w262_ ;
	wire _w261_ ;
	wire _w260_ ;
	wire _w259_ ;
	wire _w258_ ;
	wire _w257_ ;
	wire _w270_ ;
	wire _w271_ ;
	wire _w272_ ;
	wire _w273_ ;
	wire _w274_ ;
	wire _w275_ ;
	wire _w276_ ;
	wire _w277_ ;
	wire _w278_ ;
	wire _w279_ ;
	wire _w280_ ;
	wire _w281_ ;
	wire _w282_ ;
	wire _w283_ ;
	wire _w284_ ;
	wire _w285_ ;
	wire _w316_ ;
	wire _w317_ ;
	wire _w318_ ;
	wire _w319_ ;
	wire _w320_ ;
	wire _w321_ ;
	wire _w322_ ;
	wire _w323_ ;
	wire _w324_ ;
	wire _w325_ ;
	wire _w326_ ;
	wire _w327_ ;
	wire _w328_ ;
	wire _w329_ ;
	wire _w330_ ;
	wire _w331_ ;
	wire _w332_ ;
	wire _w333_ ;
	wire _w334_ ;
	wire _w335_ ;
	wire _w336_ ;
	wire _w337_ ;
	wire _w338_ ;
	wire _w339_ ;
	wire _w340_ ;
	wire _w341_ ;
	wire _w342_ ;
	wire _w343_ ;
	wire _w344_ ;
	wire _w345_ ;
	wire _w346_ ;
	wire _w347_ ;
	wire _w348_ ;
	wire _w349_ ;
	wire _w350_ ;
	wire _w351_ ;
	wire _w352_ ;
	wire _w353_ ;
	wire _w354_ ;
	wire _w355_ ;
	wire _w356_ ;
	wire _w357_ ;
	wire _w358_ ;
	wire _w359_ ;
	wire _w360_ ;
	wire _w361_ ;
	wire _w362_ ;
	wire _w363_ ;
	wire _w364_ ;
	wire _w365_ ;
	wire _w366_ ;
	wire _w367_ ;
	wire _w368_ ;
	wire _w369_ ;
	wire _w370_ ;
	wire _w371_ ;
	wire _w372_ ;
	wire _w373_ ;
	wire _w374_ ;
	wire _w375_ ;
	wire _w376_ ;
	wire _w377_ ;
	wire _w378_ ;
	wire _w379_ ;
	wire _w380_ ;
	wire _w381_ ;
	wire _w382_ ;
	wire _w383_ ;
	wire _w514_ ;
	wire _w515_ ;
	wire _w516_ ;
	wire _w517_ ;
	wire _w518_ ;
	wire _w519_ ;
	wire _w520_ ;
	wire _w521_ ;
	wire _w522_ ;
	wire _w523_ ;
	wire _w524_ ;
	wire _w525_ ;
	wire _w526_ ;
	wire _w527_ ;
	wire _w528_ ;
	wire _w529_ ;
	wire _w530_ ;
	wire _w531_ ;
	wire _w532_ ;
	wire _w533_ ;
	wire _w534_ ;
	wire _w535_ ;
	wire _w536_ ;
	wire _w537_ ;
	wire _w538_ ;
	wire _w539_ ;
	wire _w540_ ;
	wire _w541_ ;
	wire _w542_ ;
	wire _w543_ ;
	wire _w544_ ;
	wire _w545_ ;
	wire _w546_ ;
	wire _w547_ ;
	wire _w548_ ;
	wire _w549_ ;
	wire _w550_ ;
	wire _w551_ ;
	wire _w552_ ;
	wire _w553_ ;
	wire _w554_ ;
	wire _w555_ ;
	wire _w556_ ;
	wire _w557_ ;
	wire _w558_ ;
	wire _w559_ ;
	wire _w560_ ;
	wire _w561_ ;
	wire _w562_ ;
	wire _w563_ ;
	wire _w564_ ;
	wire _w565_ ;
	wire _w566_ ;
	wire _w567_ ;
	wire _w568_ ;
	wire _w569_ ;
	wire _w570_ ;
	wire _w571_ ;
	wire _w572_ ;
	wire _w573_ ;
	wire _w574_ ;
	wire _w575_ ;
	wire _w576_ ;
	wire _w577_ ;
	wire _w578_ ;
	wire _w579_ ;
	wire _w580_ ;
	wire _w581_ ;
	wire _w582_ ;
	wire _w583_ ;
	wire _w584_ ;
	wire _w585_ ;
	wire _w586_ ;
	wire _w587_ ;
	wire _w588_ ;
	wire _w589_ ;
	wire _w590_ ;
	wire _w591_ ;
	wire _w592_ ;
	wire _w593_ ;
	wire _w594_ ;
	wire _w595_ ;
	wire _w596_ ;
	wire _w597_ ;
	wire _w598_ ;
	wire _w599_ ;
	wire _w600_ ;
	wire _w601_ ;
	wire _w602_ ;
	wire _w603_ ;
	wire _w604_ ;
	wire _w605_ ;
	wire _w606_ ;
	wire _w607_ ;
	wire _w608_ ;
	wire _w609_ ;
	wire _w610_ ;
	wire _w611_ ;
	wire _w612_ ;
	wire _w613_ ;
	wire _w614_ ;
	wire _w615_ ;
	wire _w616_ ;
	wire _w617_ ;
	wire _w618_ ;
	wire _w619_ ;
	wire _w620_ ;
	wire _w621_ ;
	wire _w622_ ;
	wire _w623_ ;
	wire _w624_ ;
	wire _w625_ ;
	wire _w626_ ;
	wire _w627_ ;
	wire _w628_ ;
	wire _w629_ ;
	wire _w630_ ;
	wire _w631_ ;
	wire _w632_ ;
	wire _w633_ ;
	wire _w634_ ;
	wire _w635_ ;
	wire _w636_ ;
	wire _w637_ ;
	wire _w638_ ;
	wire _w639_ ;
	wire _w640_ ;
	wire _w641_ ;
	wire _w642_ ;
	wire _w643_ ;
	wire _w644_ ;
	wire _w645_ ;
	wire _w646_ ;
	wire _w647_ ;
	wire _w648_ ;
	wire _w649_ ;
	wire _w650_ ;
	wire _w651_ ;
	wire _w652_ ;
	wire _w653_ ;
	wire _w654_ ;
	wire _w655_ ;
	wire _w656_ ;
	wire _w657_ ;
	wire _w658_ ;
	wire _w659_ ;
	wire _w660_ ;
	wire _w661_ ;
	wire _w662_ ;
	wire _w663_ ;
	wire _w664_ ;
	wire _w665_ ;
	wire _w666_ ;
	wire _w667_ ;
	wire _w668_ ;
	wire _w669_ ;
	wire _w670_ ;
	wire _w671_ ;
	wire _w672_ ;
	wire _w673_ ;
	wire _w674_ ;
	wire _w675_ ;
	wire _w676_ ;
	wire _w677_ ;
	wire _w678_ ;
	wire _w679_ ;
	wire _w680_ ;
	wire _w681_ ;
	wire _w682_ ;
	wire _w683_ ;
	wire _w684_ ;
	wire _w685_ ;
	wire _w686_ ;
	wire _w687_ ;
	wire _w688_ ;
	wire _w689_ ;
	wire _w690_ ;
	wire _w691_ ;
	wire _w692_ ;
	wire _w693_ ;
	wire _w694_ ;
	wire _w695_ ;
	wire _w696_ ;
	wire _w697_ ;
	wire _w698_ ;
	wire _w699_ ;
	wire _w700_ ;
	wire _w701_ ;
	wire _w702_ ;
	wire _w703_ ;
	wire _w704_ ;
	wire _w705_ ;
	wire _w706_ ;
	wire _w707_ ;
	wire _w708_ ;
	wire _w709_ ;
	wire _w710_ ;
	wire _w711_ ;
	wire _w712_ ;
	wire _w713_ ;
	wire _w714_ ;
	wire _w715_ ;
	wire _w716_ ;
	wire _w717_ ;
	wire _w718_ ;
	wire _w719_ ;
	wire _w720_ ;
	wire _w721_ ;
	wire _w722_ ;
	wire _w723_ ;
	wire _w724_ ;
	wire _w725_ ;
	wire _w726_ ;
	wire _w727_ ;
	wire _w728_ ;
	wire _w729_ ;
	wire _w730_ ;
	wire _w731_ ;
	wire _w732_ ;
	wire _w733_ ;
	wire _w734_ ;
	wire _w735_ ;
	wire _w736_ ;
	wire _w737_ ;
	wire _w738_ ;
	wire _w739_ ;
	wire _w740_ ;
	wire _w741_ ;
	wire _w742_ ;
	wire _w743_ ;
	wire _w744_ ;
	wire _w745_ ;
	wire _w746_ ;
	wire _w747_ ;
	wire _w748_ ;
	wire _w749_ ;
	wire _w750_ ;
	wire _w751_ ;
	wire _w752_ ;
	wire _w753_ ;
	wire _w754_ ;
	wire _w755_ ;
	wire _w756_ ;
	wire _w757_ ;
	wire _w758_ ;
	wire _w759_ ;
	wire _w760_ ;
	wire _w761_ ;
	wire _w762_ ;
	wire _w763_ ;
	wire _w764_ ;
	wire _w765_ ;
	wire _w766_ ;
	wire _w767_ ;
	wire _w768_ ;
	wire _w769_ ;
	wire _w770_ ;
	wire _w771_ ;
	wire _w772_ ;
	wire _w773_ ;
	wire _w774_ ;
	wire _w775_ ;
	wire _w776_ ;
	wire _w777_ ;
	wire _w778_ ;
	wire _w779_ ;
	wire _w780_ ;
	wire _w781_ ;
	wire _w782_ ;
	wire _w783_ ;
	wire _w784_ ;
	wire _w785_ ;
	wire _w786_ ;
	wire _w787_ ;
	wire _w788_ ;
	wire _w789_ ;
	wire _w790_ ;
	wire _w791_ ;
	wire _w792_ ;
	wire _w793_ ;
	wire _w794_ ;
	wire _w795_ ;
	wire _w796_ ;
	wire _w797_ ;
	LUT2 #(
		.INIT('h8)
	) name0 (
		\a[0] ,
		\b[0] ,
		_w257_
	);
	LUT2 #(
		.INIT('h1)
	) name1 (
		\a[0] ,
		\b[0] ,
		_w258_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		_w257_,
		_w258_,
		_w259_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		\a[1] ,
		\b[1] ,
		_w260_
	);
	LUT2 #(
		.INIT('h8)
	) name4 (
		\a[1] ,
		\b[1] ,
		_w261_
	);
	LUT2 #(
		.INIT('h1)
	) name5 (
		_w260_,
		_w261_,
		_w262_
	);
	LUT2 #(
		.INIT('h2)
	) name6 (
		_w257_,
		_w262_,
		_w263_
	);
	LUT2 #(
		.INIT('h4)
	) name7 (
		_w257_,
		_w262_,
		_w264_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w263_,
		_w264_,
		_w265_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		\a[2] ,
		\b[2] ,
		_w266_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		\a[2] ,
		\b[2] ,
		_w267_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w266_,
		_w267_,
		_w268_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w257_,
		_w261_,
		_w269_
	);
	LUT2 #(
		.INIT('h1)
	) name13 (
		_w260_,
		_w269_,
		_w270_
	);
	LUT2 #(
		.INIT('h4)
	) name14 (
		_w268_,
		_w270_,
		_w271_
	);
	LUT2 #(
		.INIT('h2)
	) name15 (
		_w268_,
		_w270_,
		_w272_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w271_,
		_w272_,
		_w273_
	);
	LUT2 #(
		.INIT('h1)
	) name17 (
		\a[3] ,
		\b[3] ,
		_w274_
	);
	LUT2 #(
		.INIT('h8)
	) name18 (
		\a[3] ,
		\b[3] ,
		_w275_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w274_,
		_w275_,
		_w276_
	);
	LUT2 #(
		.INIT('h1)
	) name20 (
		_w267_,
		_w270_,
		_w277_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w266_,
		_w277_,
		_w278_
	);
	LUT2 #(
		.INIT('h4)
	) name22 (
		_w276_,
		_w278_,
		_w279_
	);
	LUT2 #(
		.INIT('h2)
	) name23 (
		_w276_,
		_w278_,
		_w280_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w279_,
		_w280_,
		_w281_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		\a[4] ,
		\b[4] ,
		_w282_
	);
	LUT2 #(
		.INIT('h8)
	) name26 (
		\a[4] ,
		\b[4] ,
		_w283_
	);
	LUT2 #(
		.INIT('h1)
	) name27 (
		_w282_,
		_w283_,
		_w284_
	);
	LUT2 #(
		.INIT('h1)
	) name28 (
		_w275_,
		_w278_,
		_w285_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w274_,
		_w285_,
		_w286_
	);
	LUT2 #(
		.INIT('h4)
	) name30 (
		_w284_,
		_w286_,
		_w287_
	);
	LUT2 #(
		.INIT('h2)
	) name31 (
		_w284_,
		_w286_,
		_w288_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w287_,
		_w288_,
		_w289_
	);
	LUT2 #(
		.INIT('h1)
	) name33 (
		\a[5] ,
		\b[5] ,
		_w290_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		\a[5] ,
		\b[5] ,
		_w291_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w290_,
		_w291_,
		_w292_
	);
	LUT2 #(
		.INIT('h1)
	) name36 (
		_w283_,
		_w286_,
		_w293_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w282_,
		_w293_,
		_w294_
	);
	LUT2 #(
		.INIT('h4)
	) name38 (
		_w292_,
		_w294_,
		_w295_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		_w292_,
		_w294_,
		_w296_
	);
	LUT2 #(
		.INIT('h1)
	) name40 (
		_w295_,
		_w296_,
		_w297_
	);
	LUT2 #(
		.INIT('h1)
	) name41 (
		\a[6] ,
		\b[6] ,
		_w298_
	);
	LUT2 #(
		.INIT('h8)
	) name42 (
		\a[6] ,
		\b[6] ,
		_w299_
	);
	LUT2 #(
		.INIT('h1)
	) name43 (
		_w298_,
		_w299_,
		_w300_
	);
	LUT2 #(
		.INIT('h1)
	) name44 (
		_w291_,
		_w294_,
		_w301_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w290_,
		_w301_,
		_w302_
	);
	LUT2 #(
		.INIT('h4)
	) name46 (
		_w300_,
		_w302_,
		_w303_
	);
	LUT2 #(
		.INIT('h2)
	) name47 (
		_w300_,
		_w302_,
		_w304_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w303_,
		_w304_,
		_w305_
	);
	LUT2 #(
		.INIT('h1)
	) name49 (
		\a[7] ,
		\b[7] ,
		_w306_
	);
	LUT2 #(
		.INIT('h8)
	) name50 (
		\a[7] ,
		\b[7] ,
		_w307_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w306_,
		_w307_,
		_w308_
	);
	LUT2 #(
		.INIT('h1)
	) name52 (
		_w299_,
		_w302_,
		_w309_
	);
	LUT2 #(
		.INIT('h1)
	) name53 (
		_w298_,
		_w309_,
		_w310_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		_w308_,
		_w310_,
		_w311_
	);
	LUT2 #(
		.INIT('h2)
	) name55 (
		_w308_,
		_w310_,
		_w312_
	);
	LUT2 #(
		.INIT('h1)
	) name56 (
		_w311_,
		_w312_,
		_w313_
	);
	LUT2 #(
		.INIT('h1)
	) name57 (
		\a[8] ,
		\b[8] ,
		_w314_
	);
	LUT2 #(
		.INIT('h8)
	) name58 (
		\a[8] ,
		\b[8] ,
		_w315_
	);
	LUT2 #(
		.INIT('h1)
	) name59 (
		_w314_,
		_w315_,
		_w316_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w307_,
		_w310_,
		_w317_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w306_,
		_w317_,
		_w318_
	);
	LUT2 #(
		.INIT('h4)
	) name62 (
		_w316_,
		_w318_,
		_w319_
	);
	LUT2 #(
		.INIT('h2)
	) name63 (
		_w316_,
		_w318_,
		_w320_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w319_,
		_w320_,
		_w321_
	);
	LUT2 #(
		.INIT('h1)
	) name65 (
		\a[9] ,
		\b[9] ,
		_w322_
	);
	LUT2 #(
		.INIT('h8)
	) name66 (
		\a[9] ,
		\b[9] ,
		_w323_
	);
	LUT2 #(
		.INIT('h1)
	) name67 (
		_w322_,
		_w323_,
		_w324_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w315_,
		_w318_,
		_w325_
	);
	LUT2 #(
		.INIT('h1)
	) name69 (
		_w314_,
		_w325_,
		_w326_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		_w324_,
		_w326_,
		_w327_
	);
	LUT2 #(
		.INIT('h2)
	) name71 (
		_w324_,
		_w326_,
		_w328_
	);
	LUT2 #(
		.INIT('h1)
	) name72 (
		_w327_,
		_w328_,
		_w329_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		\a[10] ,
		\b[10] ,
		_w330_
	);
	LUT2 #(
		.INIT('h8)
	) name74 (
		\a[10] ,
		\b[10] ,
		_w331_
	);
	LUT2 #(
		.INIT('h1)
	) name75 (
		_w330_,
		_w331_,
		_w332_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w323_,
		_w326_,
		_w333_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w322_,
		_w333_,
		_w334_
	);
	LUT2 #(
		.INIT('h4)
	) name78 (
		_w332_,
		_w334_,
		_w335_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		_w332_,
		_w334_,
		_w336_
	);
	LUT2 #(
		.INIT('h1)
	) name80 (
		_w335_,
		_w336_,
		_w337_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		\a[11] ,
		\b[11] ,
		_w338_
	);
	LUT2 #(
		.INIT('h8)
	) name82 (
		\a[11] ,
		\b[11] ,
		_w339_
	);
	LUT2 #(
		.INIT('h1)
	) name83 (
		_w338_,
		_w339_,
		_w340_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w331_,
		_w334_,
		_w341_
	);
	LUT2 #(
		.INIT('h1)
	) name85 (
		_w330_,
		_w341_,
		_w342_
	);
	LUT2 #(
		.INIT('h4)
	) name86 (
		_w340_,
		_w342_,
		_w343_
	);
	LUT2 #(
		.INIT('h2)
	) name87 (
		_w340_,
		_w342_,
		_w344_
	);
	LUT2 #(
		.INIT('h1)
	) name88 (
		_w343_,
		_w344_,
		_w345_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		\a[12] ,
		\b[12] ,
		_w346_
	);
	LUT2 #(
		.INIT('h8)
	) name90 (
		\a[12] ,
		\b[12] ,
		_w347_
	);
	LUT2 #(
		.INIT('h1)
	) name91 (
		_w346_,
		_w347_,
		_w348_
	);
	LUT2 #(
		.INIT('h1)
	) name92 (
		_w339_,
		_w342_,
		_w349_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w338_,
		_w349_,
		_w350_
	);
	LUT2 #(
		.INIT('h4)
	) name94 (
		_w348_,
		_w350_,
		_w351_
	);
	LUT2 #(
		.INIT('h2)
	) name95 (
		_w348_,
		_w350_,
		_w352_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w351_,
		_w352_,
		_w353_
	);
	LUT2 #(
		.INIT('h1)
	) name97 (
		\a[13] ,
		\b[13] ,
		_w354_
	);
	LUT2 #(
		.INIT('h8)
	) name98 (
		\a[13] ,
		\b[13] ,
		_w355_
	);
	LUT2 #(
		.INIT('h1)
	) name99 (
		_w354_,
		_w355_,
		_w356_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w347_,
		_w350_,
		_w357_
	);
	LUT2 #(
		.INIT('h1)
	) name101 (
		_w346_,
		_w357_,
		_w358_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w356_,
		_w358_,
		_w359_
	);
	LUT2 #(
		.INIT('h2)
	) name103 (
		_w356_,
		_w358_,
		_w360_
	);
	LUT2 #(
		.INIT('h1)
	) name104 (
		_w359_,
		_w360_,
		_w361_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		\a[14] ,
		\b[14] ,
		_w362_
	);
	LUT2 #(
		.INIT('h8)
	) name106 (
		\a[14] ,
		\b[14] ,
		_w363_
	);
	LUT2 #(
		.INIT('h1)
	) name107 (
		_w362_,
		_w363_,
		_w364_
	);
	LUT2 #(
		.INIT('h1)
	) name108 (
		_w355_,
		_w358_,
		_w365_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w354_,
		_w365_,
		_w366_
	);
	LUT2 #(
		.INIT('h4)
	) name110 (
		_w364_,
		_w366_,
		_w367_
	);
	LUT2 #(
		.INIT('h2)
	) name111 (
		_w364_,
		_w366_,
		_w368_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w367_,
		_w368_,
		_w369_
	);
	LUT2 #(
		.INIT('h1)
	) name113 (
		\a[15] ,
		\b[15] ,
		_w370_
	);
	LUT2 #(
		.INIT('h8)
	) name114 (
		\a[15] ,
		\b[15] ,
		_w371_
	);
	LUT2 #(
		.INIT('h1)
	) name115 (
		_w370_,
		_w371_,
		_w372_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w363_,
		_w366_,
		_w373_
	);
	LUT2 #(
		.INIT('h1)
	) name117 (
		_w362_,
		_w373_,
		_w374_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w372_,
		_w374_,
		_w375_
	);
	LUT2 #(
		.INIT('h2)
	) name119 (
		_w372_,
		_w374_,
		_w376_
	);
	LUT2 #(
		.INIT('h1)
	) name120 (
		_w375_,
		_w376_,
		_w377_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		\a[16] ,
		\b[16] ,
		_w378_
	);
	LUT2 #(
		.INIT('h8)
	) name122 (
		\a[16] ,
		\b[16] ,
		_w379_
	);
	LUT2 #(
		.INIT('h1)
	) name123 (
		_w378_,
		_w379_,
		_w380_
	);
	LUT2 #(
		.INIT('h1)
	) name124 (
		_w371_,
		_w374_,
		_w381_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w370_,
		_w381_,
		_w382_
	);
	LUT2 #(
		.INIT('h4)
	) name126 (
		_w380_,
		_w382_,
		_w383_
	);
	LUT2 #(
		.INIT('h2)
	) name127 (
		_w380_,
		_w382_,
		_w384_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w383_,
		_w384_,
		_w385_
	);
	LUT2 #(
		.INIT('h1)
	) name129 (
		\a[17] ,
		\b[17] ,
		_w386_
	);
	LUT2 #(
		.INIT('h8)
	) name130 (
		\a[17] ,
		\b[17] ,
		_w387_
	);
	LUT2 #(
		.INIT('h1)
	) name131 (
		_w386_,
		_w387_,
		_w388_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w379_,
		_w382_,
		_w389_
	);
	LUT2 #(
		.INIT('h1)
	) name133 (
		_w378_,
		_w389_,
		_w390_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w388_,
		_w390_,
		_w391_
	);
	LUT2 #(
		.INIT('h2)
	) name135 (
		_w388_,
		_w390_,
		_w392_
	);
	LUT2 #(
		.INIT('h1)
	) name136 (
		_w391_,
		_w392_,
		_w393_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		\a[18] ,
		\b[18] ,
		_w394_
	);
	LUT2 #(
		.INIT('h8)
	) name138 (
		\a[18] ,
		\b[18] ,
		_w395_
	);
	LUT2 #(
		.INIT('h1)
	) name139 (
		_w394_,
		_w395_,
		_w396_
	);
	LUT2 #(
		.INIT('h1)
	) name140 (
		_w387_,
		_w390_,
		_w397_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w386_,
		_w397_,
		_w398_
	);
	LUT2 #(
		.INIT('h4)
	) name142 (
		_w396_,
		_w398_,
		_w399_
	);
	LUT2 #(
		.INIT('h2)
	) name143 (
		_w396_,
		_w398_,
		_w400_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w399_,
		_w400_,
		_w401_
	);
	LUT2 #(
		.INIT('h1)
	) name145 (
		\a[19] ,
		\b[19] ,
		_w402_
	);
	LUT2 #(
		.INIT('h8)
	) name146 (
		\a[19] ,
		\b[19] ,
		_w403_
	);
	LUT2 #(
		.INIT('h1)
	) name147 (
		_w402_,
		_w403_,
		_w404_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w395_,
		_w398_,
		_w405_
	);
	LUT2 #(
		.INIT('h1)
	) name149 (
		_w394_,
		_w405_,
		_w406_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w404_,
		_w406_,
		_w407_
	);
	LUT2 #(
		.INIT('h2)
	) name151 (
		_w404_,
		_w406_,
		_w408_
	);
	LUT2 #(
		.INIT('h1)
	) name152 (
		_w407_,
		_w408_,
		_w409_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		\a[20] ,
		\b[20] ,
		_w410_
	);
	LUT2 #(
		.INIT('h8)
	) name154 (
		\a[20] ,
		\b[20] ,
		_w411_
	);
	LUT2 #(
		.INIT('h1)
	) name155 (
		_w410_,
		_w411_,
		_w412_
	);
	LUT2 #(
		.INIT('h1)
	) name156 (
		_w403_,
		_w406_,
		_w413_
	);
	LUT2 #(
		.INIT('h1)
	) name157 (
		_w402_,
		_w413_,
		_w414_
	);
	LUT2 #(
		.INIT('h4)
	) name158 (
		_w412_,
		_w414_,
		_w415_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		_w412_,
		_w414_,
		_w416_
	);
	LUT2 #(
		.INIT('h1)
	) name160 (
		_w415_,
		_w416_,
		_w417_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		\a[21] ,
		\b[21] ,
		_w418_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		\a[21] ,
		\b[21] ,
		_w419_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w418_,
		_w419_,
		_w420_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w411_,
		_w414_,
		_w421_
	);
	LUT2 #(
		.INIT('h1)
	) name165 (
		_w410_,
		_w421_,
		_w422_
	);
	LUT2 #(
		.INIT('h4)
	) name166 (
		_w420_,
		_w422_,
		_w423_
	);
	LUT2 #(
		.INIT('h2)
	) name167 (
		_w420_,
		_w422_,
		_w424_
	);
	LUT2 #(
		.INIT('h1)
	) name168 (
		_w423_,
		_w424_,
		_w425_
	);
	LUT2 #(
		.INIT('h1)
	) name169 (
		\a[22] ,
		\b[22] ,
		_w426_
	);
	LUT2 #(
		.INIT('h8)
	) name170 (
		\a[22] ,
		\b[22] ,
		_w427_
	);
	LUT2 #(
		.INIT('h1)
	) name171 (
		_w426_,
		_w427_,
		_w428_
	);
	LUT2 #(
		.INIT('h1)
	) name172 (
		_w419_,
		_w422_,
		_w429_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w418_,
		_w429_,
		_w430_
	);
	LUT2 #(
		.INIT('h4)
	) name174 (
		_w428_,
		_w430_,
		_w431_
	);
	LUT2 #(
		.INIT('h2)
	) name175 (
		_w428_,
		_w430_,
		_w432_
	);
	LUT2 #(
		.INIT('h1)
	) name176 (
		_w431_,
		_w432_,
		_w433_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		\a[23] ,
		\b[23] ,
		_w434_
	);
	LUT2 #(
		.INIT('h8)
	) name178 (
		\a[23] ,
		\b[23] ,
		_w435_
	);
	LUT2 #(
		.INIT('h1)
	) name179 (
		_w434_,
		_w435_,
		_w436_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w427_,
		_w430_,
		_w437_
	);
	LUT2 #(
		.INIT('h1)
	) name181 (
		_w426_,
		_w437_,
		_w438_
	);
	LUT2 #(
		.INIT('h4)
	) name182 (
		_w436_,
		_w438_,
		_w439_
	);
	LUT2 #(
		.INIT('h2)
	) name183 (
		_w436_,
		_w438_,
		_w440_
	);
	LUT2 #(
		.INIT('h1)
	) name184 (
		_w439_,
		_w440_,
		_w441_
	);
	LUT2 #(
		.INIT('h1)
	) name185 (
		\a[24] ,
		\b[24] ,
		_w442_
	);
	LUT2 #(
		.INIT('h8)
	) name186 (
		\a[24] ,
		\b[24] ,
		_w443_
	);
	LUT2 #(
		.INIT('h1)
	) name187 (
		_w442_,
		_w443_,
		_w444_
	);
	LUT2 #(
		.INIT('h1)
	) name188 (
		_w435_,
		_w438_,
		_w445_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w434_,
		_w445_,
		_w446_
	);
	LUT2 #(
		.INIT('h4)
	) name190 (
		_w444_,
		_w446_,
		_w447_
	);
	LUT2 #(
		.INIT('h2)
	) name191 (
		_w444_,
		_w446_,
		_w448_
	);
	LUT2 #(
		.INIT('h1)
	) name192 (
		_w447_,
		_w448_,
		_w449_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		\a[25] ,
		\b[25] ,
		_w450_
	);
	LUT2 #(
		.INIT('h8)
	) name194 (
		\a[25] ,
		\b[25] ,
		_w451_
	);
	LUT2 #(
		.INIT('h1)
	) name195 (
		_w450_,
		_w451_,
		_w452_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w443_,
		_w446_,
		_w453_
	);
	LUT2 #(
		.INIT('h1)
	) name197 (
		_w442_,
		_w453_,
		_w454_
	);
	LUT2 #(
		.INIT('h4)
	) name198 (
		_w452_,
		_w454_,
		_w455_
	);
	LUT2 #(
		.INIT('h2)
	) name199 (
		_w452_,
		_w454_,
		_w456_
	);
	LUT2 #(
		.INIT('h1)
	) name200 (
		_w455_,
		_w456_,
		_w457_
	);
	LUT2 #(
		.INIT('h1)
	) name201 (
		\a[26] ,
		\b[26] ,
		_w458_
	);
	LUT2 #(
		.INIT('h8)
	) name202 (
		\a[26] ,
		\b[26] ,
		_w459_
	);
	LUT2 #(
		.INIT('h1)
	) name203 (
		_w458_,
		_w459_,
		_w460_
	);
	LUT2 #(
		.INIT('h1)
	) name204 (
		_w451_,
		_w454_,
		_w461_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w450_,
		_w461_,
		_w462_
	);
	LUT2 #(
		.INIT('h4)
	) name206 (
		_w460_,
		_w462_,
		_w463_
	);
	LUT2 #(
		.INIT('h2)
	) name207 (
		_w460_,
		_w462_,
		_w464_
	);
	LUT2 #(
		.INIT('h1)
	) name208 (
		_w463_,
		_w464_,
		_w465_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		\a[27] ,
		\b[27] ,
		_w466_
	);
	LUT2 #(
		.INIT('h8)
	) name210 (
		\a[27] ,
		\b[27] ,
		_w467_
	);
	LUT2 #(
		.INIT('h1)
	) name211 (
		_w466_,
		_w467_,
		_w468_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w459_,
		_w462_,
		_w469_
	);
	LUT2 #(
		.INIT('h1)
	) name213 (
		_w458_,
		_w469_,
		_w470_
	);
	LUT2 #(
		.INIT('h4)
	) name214 (
		_w468_,
		_w470_,
		_w471_
	);
	LUT2 #(
		.INIT('h2)
	) name215 (
		_w468_,
		_w470_,
		_w472_
	);
	LUT2 #(
		.INIT('h1)
	) name216 (
		_w471_,
		_w472_,
		_w473_
	);
	LUT2 #(
		.INIT('h1)
	) name217 (
		\a[28] ,
		\b[28] ,
		_w474_
	);
	LUT2 #(
		.INIT('h8)
	) name218 (
		\a[28] ,
		\b[28] ,
		_w475_
	);
	LUT2 #(
		.INIT('h1)
	) name219 (
		_w474_,
		_w475_,
		_w476_
	);
	LUT2 #(
		.INIT('h1)
	) name220 (
		_w467_,
		_w470_,
		_w477_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w466_,
		_w477_,
		_w478_
	);
	LUT2 #(
		.INIT('h4)
	) name222 (
		_w476_,
		_w478_,
		_w479_
	);
	LUT2 #(
		.INIT('h2)
	) name223 (
		_w476_,
		_w478_,
		_w480_
	);
	LUT2 #(
		.INIT('h1)
	) name224 (
		_w479_,
		_w480_,
		_w481_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		\a[29] ,
		\b[29] ,
		_w482_
	);
	LUT2 #(
		.INIT('h8)
	) name226 (
		\a[29] ,
		\b[29] ,
		_w483_
	);
	LUT2 #(
		.INIT('h1)
	) name227 (
		_w482_,
		_w483_,
		_w484_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w475_,
		_w478_,
		_w485_
	);
	LUT2 #(
		.INIT('h1)
	) name229 (
		_w474_,
		_w485_,
		_w486_
	);
	LUT2 #(
		.INIT('h4)
	) name230 (
		_w484_,
		_w486_,
		_w487_
	);
	LUT2 #(
		.INIT('h2)
	) name231 (
		_w484_,
		_w486_,
		_w488_
	);
	LUT2 #(
		.INIT('h1)
	) name232 (
		_w487_,
		_w488_,
		_w489_
	);
	LUT2 #(
		.INIT('h1)
	) name233 (
		\a[30] ,
		\b[30] ,
		_w490_
	);
	LUT2 #(
		.INIT('h8)
	) name234 (
		\a[30] ,
		\b[30] ,
		_w491_
	);
	LUT2 #(
		.INIT('h1)
	) name235 (
		_w490_,
		_w491_,
		_w492_
	);
	LUT2 #(
		.INIT('h1)
	) name236 (
		_w483_,
		_w486_,
		_w493_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w482_,
		_w493_,
		_w494_
	);
	LUT2 #(
		.INIT('h4)
	) name238 (
		_w492_,
		_w494_,
		_w495_
	);
	LUT2 #(
		.INIT('h2)
	) name239 (
		_w492_,
		_w494_,
		_w496_
	);
	LUT2 #(
		.INIT('h1)
	) name240 (
		_w495_,
		_w496_,
		_w497_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		\a[31] ,
		\b[31] ,
		_w498_
	);
	LUT2 #(
		.INIT('h8)
	) name242 (
		\a[31] ,
		\b[31] ,
		_w499_
	);
	LUT2 #(
		.INIT('h1)
	) name243 (
		_w498_,
		_w499_,
		_w500_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w491_,
		_w494_,
		_w501_
	);
	LUT2 #(
		.INIT('h1)
	) name245 (
		_w490_,
		_w501_,
		_w502_
	);
	LUT2 #(
		.INIT('h4)
	) name246 (
		_w500_,
		_w502_,
		_w503_
	);
	LUT2 #(
		.INIT('h2)
	) name247 (
		_w500_,
		_w502_,
		_w504_
	);
	LUT2 #(
		.INIT('h1)
	) name248 (
		_w503_,
		_w504_,
		_w505_
	);
	LUT2 #(
		.INIT('h1)
	) name249 (
		\a[32] ,
		\b[32] ,
		_w506_
	);
	LUT2 #(
		.INIT('h8)
	) name250 (
		\a[32] ,
		\b[32] ,
		_w507_
	);
	LUT2 #(
		.INIT('h1)
	) name251 (
		_w506_,
		_w507_,
		_w508_
	);
	LUT2 #(
		.INIT('h1)
	) name252 (
		_w499_,
		_w502_,
		_w509_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w498_,
		_w509_,
		_w510_
	);
	LUT2 #(
		.INIT('h4)
	) name254 (
		_w508_,
		_w510_,
		_w511_
	);
	LUT2 #(
		.INIT('h2)
	) name255 (
		_w508_,
		_w510_,
		_w512_
	);
	LUT2 #(
		.INIT('h1)
	) name256 (
		_w511_,
		_w512_,
		_w513_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		\a[33] ,
		\b[33] ,
		_w514_
	);
	LUT2 #(
		.INIT('h8)
	) name258 (
		\a[33] ,
		\b[33] ,
		_w515_
	);
	LUT2 #(
		.INIT('h1)
	) name259 (
		_w514_,
		_w515_,
		_w516_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w507_,
		_w510_,
		_w517_
	);
	LUT2 #(
		.INIT('h1)
	) name261 (
		_w506_,
		_w517_,
		_w518_
	);
	LUT2 #(
		.INIT('h4)
	) name262 (
		_w516_,
		_w518_,
		_w519_
	);
	LUT2 #(
		.INIT('h2)
	) name263 (
		_w516_,
		_w518_,
		_w520_
	);
	LUT2 #(
		.INIT('h1)
	) name264 (
		_w519_,
		_w520_,
		_w521_
	);
	LUT2 #(
		.INIT('h1)
	) name265 (
		\a[34] ,
		\b[34] ,
		_w522_
	);
	LUT2 #(
		.INIT('h8)
	) name266 (
		\a[34] ,
		\b[34] ,
		_w523_
	);
	LUT2 #(
		.INIT('h1)
	) name267 (
		_w522_,
		_w523_,
		_w524_
	);
	LUT2 #(
		.INIT('h1)
	) name268 (
		_w515_,
		_w518_,
		_w525_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w514_,
		_w525_,
		_w526_
	);
	LUT2 #(
		.INIT('h4)
	) name270 (
		_w524_,
		_w526_,
		_w527_
	);
	LUT2 #(
		.INIT('h2)
	) name271 (
		_w524_,
		_w526_,
		_w528_
	);
	LUT2 #(
		.INIT('h1)
	) name272 (
		_w527_,
		_w528_,
		_w529_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		\a[35] ,
		\b[35] ,
		_w530_
	);
	LUT2 #(
		.INIT('h8)
	) name274 (
		\a[35] ,
		\b[35] ,
		_w531_
	);
	LUT2 #(
		.INIT('h1)
	) name275 (
		_w530_,
		_w531_,
		_w532_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w523_,
		_w526_,
		_w533_
	);
	LUT2 #(
		.INIT('h1)
	) name277 (
		_w522_,
		_w533_,
		_w534_
	);
	LUT2 #(
		.INIT('h4)
	) name278 (
		_w532_,
		_w534_,
		_w535_
	);
	LUT2 #(
		.INIT('h2)
	) name279 (
		_w532_,
		_w534_,
		_w536_
	);
	LUT2 #(
		.INIT('h1)
	) name280 (
		_w535_,
		_w536_,
		_w537_
	);
	LUT2 #(
		.INIT('h1)
	) name281 (
		\a[36] ,
		\b[36] ,
		_w538_
	);
	LUT2 #(
		.INIT('h8)
	) name282 (
		\a[36] ,
		\b[36] ,
		_w539_
	);
	LUT2 #(
		.INIT('h1)
	) name283 (
		_w538_,
		_w539_,
		_w540_
	);
	LUT2 #(
		.INIT('h1)
	) name284 (
		_w531_,
		_w534_,
		_w541_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w530_,
		_w541_,
		_w542_
	);
	LUT2 #(
		.INIT('h4)
	) name286 (
		_w540_,
		_w542_,
		_w543_
	);
	LUT2 #(
		.INIT('h2)
	) name287 (
		_w540_,
		_w542_,
		_w544_
	);
	LUT2 #(
		.INIT('h1)
	) name288 (
		_w543_,
		_w544_,
		_w545_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		\a[37] ,
		\b[37] ,
		_w546_
	);
	LUT2 #(
		.INIT('h8)
	) name290 (
		\a[37] ,
		\b[37] ,
		_w547_
	);
	LUT2 #(
		.INIT('h1)
	) name291 (
		_w546_,
		_w547_,
		_w548_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w539_,
		_w542_,
		_w549_
	);
	LUT2 #(
		.INIT('h1)
	) name293 (
		_w538_,
		_w549_,
		_w550_
	);
	LUT2 #(
		.INIT('h4)
	) name294 (
		_w548_,
		_w550_,
		_w551_
	);
	LUT2 #(
		.INIT('h2)
	) name295 (
		_w548_,
		_w550_,
		_w552_
	);
	LUT2 #(
		.INIT('h1)
	) name296 (
		_w551_,
		_w552_,
		_w553_
	);
	LUT2 #(
		.INIT('h1)
	) name297 (
		\a[38] ,
		\b[38] ,
		_w554_
	);
	LUT2 #(
		.INIT('h8)
	) name298 (
		\a[38] ,
		\b[38] ,
		_w555_
	);
	LUT2 #(
		.INIT('h1)
	) name299 (
		_w554_,
		_w555_,
		_w556_
	);
	LUT2 #(
		.INIT('h1)
	) name300 (
		_w547_,
		_w550_,
		_w557_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w546_,
		_w557_,
		_w558_
	);
	LUT2 #(
		.INIT('h4)
	) name302 (
		_w556_,
		_w558_,
		_w559_
	);
	LUT2 #(
		.INIT('h2)
	) name303 (
		_w556_,
		_w558_,
		_w560_
	);
	LUT2 #(
		.INIT('h1)
	) name304 (
		_w559_,
		_w560_,
		_w561_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		\a[39] ,
		\b[39] ,
		_w562_
	);
	LUT2 #(
		.INIT('h8)
	) name306 (
		\a[39] ,
		\b[39] ,
		_w563_
	);
	LUT2 #(
		.INIT('h1)
	) name307 (
		_w562_,
		_w563_,
		_w564_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w555_,
		_w558_,
		_w565_
	);
	LUT2 #(
		.INIT('h1)
	) name309 (
		_w554_,
		_w565_,
		_w566_
	);
	LUT2 #(
		.INIT('h4)
	) name310 (
		_w564_,
		_w566_,
		_w567_
	);
	LUT2 #(
		.INIT('h2)
	) name311 (
		_w564_,
		_w566_,
		_w568_
	);
	LUT2 #(
		.INIT('h1)
	) name312 (
		_w567_,
		_w568_,
		_w569_
	);
	LUT2 #(
		.INIT('h1)
	) name313 (
		\a[40] ,
		\b[40] ,
		_w570_
	);
	LUT2 #(
		.INIT('h8)
	) name314 (
		\a[40] ,
		\b[40] ,
		_w571_
	);
	LUT2 #(
		.INIT('h1)
	) name315 (
		_w570_,
		_w571_,
		_w572_
	);
	LUT2 #(
		.INIT('h1)
	) name316 (
		_w563_,
		_w566_,
		_w573_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w562_,
		_w573_,
		_w574_
	);
	LUT2 #(
		.INIT('h4)
	) name318 (
		_w572_,
		_w574_,
		_w575_
	);
	LUT2 #(
		.INIT('h2)
	) name319 (
		_w572_,
		_w574_,
		_w576_
	);
	LUT2 #(
		.INIT('h1)
	) name320 (
		_w575_,
		_w576_,
		_w577_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		\a[41] ,
		\b[41] ,
		_w578_
	);
	LUT2 #(
		.INIT('h8)
	) name322 (
		\a[41] ,
		\b[41] ,
		_w579_
	);
	LUT2 #(
		.INIT('h1)
	) name323 (
		_w578_,
		_w579_,
		_w580_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w571_,
		_w574_,
		_w581_
	);
	LUT2 #(
		.INIT('h1)
	) name325 (
		_w570_,
		_w581_,
		_w582_
	);
	LUT2 #(
		.INIT('h4)
	) name326 (
		_w580_,
		_w582_,
		_w583_
	);
	LUT2 #(
		.INIT('h2)
	) name327 (
		_w580_,
		_w582_,
		_w584_
	);
	LUT2 #(
		.INIT('h1)
	) name328 (
		_w583_,
		_w584_,
		_w585_
	);
	LUT2 #(
		.INIT('h1)
	) name329 (
		\a[42] ,
		\b[42] ,
		_w586_
	);
	LUT2 #(
		.INIT('h8)
	) name330 (
		\a[42] ,
		\b[42] ,
		_w587_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w586_,
		_w587_,
		_w588_
	);
	LUT2 #(
		.INIT('h1)
	) name332 (
		_w579_,
		_w582_,
		_w589_
	);
	LUT2 #(
		.INIT('h1)
	) name333 (
		_w578_,
		_w589_,
		_w590_
	);
	LUT2 #(
		.INIT('h4)
	) name334 (
		_w588_,
		_w590_,
		_w591_
	);
	LUT2 #(
		.INIT('h2)
	) name335 (
		_w588_,
		_w590_,
		_w592_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w591_,
		_w592_,
		_w593_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		\a[43] ,
		\b[43] ,
		_w594_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		\a[43] ,
		\b[43] ,
		_w595_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w594_,
		_w595_,
		_w596_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w587_,
		_w590_,
		_w597_
	);
	LUT2 #(
		.INIT('h1)
	) name341 (
		_w586_,
		_w597_,
		_w598_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		_w596_,
		_w598_,
		_w599_
	);
	LUT2 #(
		.INIT('h2)
	) name343 (
		_w596_,
		_w598_,
		_w600_
	);
	LUT2 #(
		.INIT('h1)
	) name344 (
		_w599_,
		_w600_,
		_w601_
	);
	LUT2 #(
		.INIT('h1)
	) name345 (
		\a[44] ,
		\b[44] ,
		_w602_
	);
	LUT2 #(
		.INIT('h8)
	) name346 (
		\a[44] ,
		\b[44] ,
		_w603_
	);
	LUT2 #(
		.INIT('h1)
	) name347 (
		_w602_,
		_w603_,
		_w604_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		_w595_,
		_w598_,
		_w605_
	);
	LUT2 #(
		.INIT('h1)
	) name349 (
		_w594_,
		_w605_,
		_w606_
	);
	LUT2 #(
		.INIT('h4)
	) name350 (
		_w604_,
		_w606_,
		_w607_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w604_,
		_w606_,
		_w608_
	);
	LUT2 #(
		.INIT('h1)
	) name352 (
		_w607_,
		_w608_,
		_w609_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		\a[45] ,
		\b[45] ,
		_w610_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		\a[45] ,
		\b[45] ,
		_w611_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		_w610_,
		_w611_,
		_w612_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w603_,
		_w606_,
		_w613_
	);
	LUT2 #(
		.INIT('h1)
	) name357 (
		_w602_,
		_w613_,
		_w614_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		_w612_,
		_w614_,
		_w615_
	);
	LUT2 #(
		.INIT('h2)
	) name359 (
		_w612_,
		_w614_,
		_w616_
	);
	LUT2 #(
		.INIT('h1)
	) name360 (
		_w615_,
		_w616_,
		_w617_
	);
	LUT2 #(
		.INIT('h1)
	) name361 (
		\a[46] ,
		\b[46] ,
		_w618_
	);
	LUT2 #(
		.INIT('h8)
	) name362 (
		\a[46] ,
		\b[46] ,
		_w619_
	);
	LUT2 #(
		.INIT('h1)
	) name363 (
		_w618_,
		_w619_,
		_w620_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		_w611_,
		_w614_,
		_w621_
	);
	LUT2 #(
		.INIT('h1)
	) name365 (
		_w610_,
		_w621_,
		_w622_
	);
	LUT2 #(
		.INIT('h4)
	) name366 (
		_w620_,
		_w622_,
		_w623_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		_w620_,
		_w622_,
		_w624_
	);
	LUT2 #(
		.INIT('h1)
	) name368 (
		_w623_,
		_w624_,
		_w625_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		\a[47] ,
		\b[47] ,
		_w626_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		\a[47] ,
		\b[47] ,
		_w627_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w626_,
		_w627_,
		_w628_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w619_,
		_w622_,
		_w629_
	);
	LUT2 #(
		.INIT('h1)
	) name373 (
		_w618_,
		_w629_,
		_w630_
	);
	LUT2 #(
		.INIT('h4)
	) name374 (
		_w628_,
		_w630_,
		_w631_
	);
	LUT2 #(
		.INIT('h2)
	) name375 (
		_w628_,
		_w630_,
		_w632_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w631_,
		_w632_,
		_w633_
	);
	LUT2 #(
		.INIT('h1)
	) name377 (
		\a[48] ,
		\b[48] ,
		_w634_
	);
	LUT2 #(
		.INIT('h8)
	) name378 (
		\a[48] ,
		\b[48] ,
		_w635_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w634_,
		_w635_,
		_w636_
	);
	LUT2 #(
		.INIT('h1)
	) name380 (
		_w627_,
		_w630_,
		_w637_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w626_,
		_w637_,
		_w638_
	);
	LUT2 #(
		.INIT('h4)
	) name382 (
		_w636_,
		_w638_,
		_w639_
	);
	LUT2 #(
		.INIT('h2)
	) name383 (
		_w636_,
		_w638_,
		_w640_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w639_,
		_w640_,
		_w641_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		\a[49] ,
		\b[49] ,
		_w642_
	);
	LUT2 #(
		.INIT('h8)
	) name386 (
		\a[49] ,
		\b[49] ,
		_w643_
	);
	LUT2 #(
		.INIT('h1)
	) name387 (
		_w642_,
		_w643_,
		_w644_
	);
	LUT2 #(
		.INIT('h1)
	) name388 (
		_w635_,
		_w638_,
		_w645_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w634_,
		_w645_,
		_w646_
	);
	LUT2 #(
		.INIT('h4)
	) name390 (
		_w644_,
		_w646_,
		_w647_
	);
	LUT2 #(
		.INIT('h2)
	) name391 (
		_w644_,
		_w646_,
		_w648_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w647_,
		_w648_,
		_w649_
	);
	LUT2 #(
		.INIT('h1)
	) name393 (
		\a[50] ,
		\b[50] ,
		_w650_
	);
	LUT2 #(
		.INIT('h8)
	) name394 (
		\a[50] ,
		\b[50] ,
		_w651_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w650_,
		_w651_,
		_w652_
	);
	LUT2 #(
		.INIT('h1)
	) name396 (
		_w643_,
		_w646_,
		_w653_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w642_,
		_w653_,
		_w654_
	);
	LUT2 #(
		.INIT('h4)
	) name398 (
		_w652_,
		_w654_,
		_w655_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		_w652_,
		_w654_,
		_w656_
	);
	LUT2 #(
		.INIT('h1)
	) name400 (
		_w655_,
		_w656_,
		_w657_
	);
	LUT2 #(
		.INIT('h1)
	) name401 (
		\a[51] ,
		\b[51] ,
		_w658_
	);
	LUT2 #(
		.INIT('h8)
	) name402 (
		\a[51] ,
		\b[51] ,
		_w659_
	);
	LUT2 #(
		.INIT('h1)
	) name403 (
		_w658_,
		_w659_,
		_w660_
	);
	LUT2 #(
		.INIT('h1)
	) name404 (
		_w651_,
		_w654_,
		_w661_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w650_,
		_w661_,
		_w662_
	);
	LUT2 #(
		.INIT('h4)
	) name406 (
		_w660_,
		_w662_,
		_w663_
	);
	LUT2 #(
		.INIT('h2)
	) name407 (
		_w660_,
		_w662_,
		_w664_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w663_,
		_w664_,
		_w665_
	);
	LUT2 #(
		.INIT('h1)
	) name409 (
		\a[52] ,
		\b[52] ,
		_w666_
	);
	LUT2 #(
		.INIT('h8)
	) name410 (
		\a[52] ,
		\b[52] ,
		_w667_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w666_,
		_w667_,
		_w668_
	);
	LUT2 #(
		.INIT('h1)
	) name412 (
		_w659_,
		_w662_,
		_w669_
	);
	LUT2 #(
		.INIT('h1)
	) name413 (
		_w658_,
		_w669_,
		_w670_
	);
	LUT2 #(
		.INIT('h4)
	) name414 (
		_w668_,
		_w670_,
		_w671_
	);
	LUT2 #(
		.INIT('h2)
	) name415 (
		_w668_,
		_w670_,
		_w672_
	);
	LUT2 #(
		.INIT('h1)
	) name416 (
		_w671_,
		_w672_,
		_w673_
	);
	LUT2 #(
		.INIT('h1)
	) name417 (
		\a[53] ,
		\b[53] ,
		_w674_
	);
	LUT2 #(
		.INIT('h8)
	) name418 (
		\a[53] ,
		\b[53] ,
		_w675_
	);
	LUT2 #(
		.INIT('h1)
	) name419 (
		_w674_,
		_w675_,
		_w676_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w667_,
		_w670_,
		_w677_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		_w666_,
		_w677_,
		_w678_
	);
	LUT2 #(
		.INIT('h4)
	) name422 (
		_w676_,
		_w678_,
		_w679_
	);
	LUT2 #(
		.INIT('h2)
	) name423 (
		_w676_,
		_w678_,
		_w680_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w679_,
		_w680_,
		_w681_
	);
	LUT2 #(
		.INIT('h1)
	) name425 (
		\a[54] ,
		\b[54] ,
		_w682_
	);
	LUT2 #(
		.INIT('h8)
	) name426 (
		\a[54] ,
		\b[54] ,
		_w683_
	);
	LUT2 #(
		.INIT('h1)
	) name427 (
		_w682_,
		_w683_,
		_w684_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w675_,
		_w678_,
		_w685_
	);
	LUT2 #(
		.INIT('h1)
	) name429 (
		_w674_,
		_w685_,
		_w686_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		_w684_,
		_w686_,
		_w687_
	);
	LUT2 #(
		.INIT('h2)
	) name431 (
		_w684_,
		_w686_,
		_w688_
	);
	LUT2 #(
		.INIT('h1)
	) name432 (
		_w687_,
		_w688_,
		_w689_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		\a[55] ,
		\b[55] ,
		_w690_
	);
	LUT2 #(
		.INIT('h8)
	) name434 (
		\a[55] ,
		\b[55] ,
		_w691_
	);
	LUT2 #(
		.INIT('h1)
	) name435 (
		_w690_,
		_w691_,
		_w692_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w683_,
		_w686_,
		_w693_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w682_,
		_w693_,
		_w694_
	);
	LUT2 #(
		.INIT('h4)
	) name438 (
		_w692_,
		_w694_,
		_w695_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		_w692_,
		_w694_,
		_w696_
	);
	LUT2 #(
		.INIT('h1)
	) name440 (
		_w695_,
		_w696_,
		_w697_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		\a[56] ,
		\b[56] ,
		_w698_
	);
	LUT2 #(
		.INIT('h8)
	) name442 (
		\a[56] ,
		\b[56] ,
		_w699_
	);
	LUT2 #(
		.INIT('h1)
	) name443 (
		_w698_,
		_w699_,
		_w700_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w691_,
		_w694_,
		_w701_
	);
	LUT2 #(
		.INIT('h1)
	) name445 (
		_w690_,
		_w701_,
		_w702_
	);
	LUT2 #(
		.INIT('h4)
	) name446 (
		_w700_,
		_w702_,
		_w703_
	);
	LUT2 #(
		.INIT('h2)
	) name447 (
		_w700_,
		_w702_,
		_w704_
	);
	LUT2 #(
		.INIT('h1)
	) name448 (
		_w703_,
		_w704_,
		_w705_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		\a[57] ,
		\b[57] ,
		_w706_
	);
	LUT2 #(
		.INIT('h8)
	) name450 (
		\a[57] ,
		\b[57] ,
		_w707_
	);
	LUT2 #(
		.INIT('h1)
	) name451 (
		_w706_,
		_w707_,
		_w708_
	);
	LUT2 #(
		.INIT('h1)
	) name452 (
		_w699_,
		_w702_,
		_w709_
	);
	LUT2 #(
		.INIT('h1)
	) name453 (
		_w698_,
		_w709_,
		_w710_
	);
	LUT2 #(
		.INIT('h4)
	) name454 (
		_w708_,
		_w710_,
		_w711_
	);
	LUT2 #(
		.INIT('h2)
	) name455 (
		_w708_,
		_w710_,
		_w712_
	);
	LUT2 #(
		.INIT('h1)
	) name456 (
		_w711_,
		_w712_,
		_w713_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		\a[58] ,
		\b[58] ,
		_w714_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		\a[58] ,
		\b[58] ,
		_w715_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w714_,
		_w715_,
		_w716_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w707_,
		_w710_,
		_w717_
	);
	LUT2 #(
		.INIT('h1)
	) name461 (
		_w706_,
		_w717_,
		_w718_
	);
	LUT2 #(
		.INIT('h4)
	) name462 (
		_w716_,
		_w718_,
		_w719_
	);
	LUT2 #(
		.INIT('h2)
	) name463 (
		_w716_,
		_w718_,
		_w720_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		_w719_,
		_w720_,
		_w721_
	);
	LUT2 #(
		.INIT('h1)
	) name465 (
		\a[59] ,
		\b[59] ,
		_w722_
	);
	LUT2 #(
		.INIT('h8)
	) name466 (
		\a[59] ,
		\b[59] ,
		_w723_
	);
	LUT2 #(
		.INIT('h1)
	) name467 (
		_w722_,
		_w723_,
		_w724_
	);
	LUT2 #(
		.INIT('h1)
	) name468 (
		_w715_,
		_w718_,
		_w725_
	);
	LUT2 #(
		.INIT('h1)
	) name469 (
		_w714_,
		_w725_,
		_w726_
	);
	LUT2 #(
		.INIT('h4)
	) name470 (
		_w724_,
		_w726_,
		_w727_
	);
	LUT2 #(
		.INIT('h2)
	) name471 (
		_w724_,
		_w726_,
		_w728_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w727_,
		_w728_,
		_w729_
	);
	LUT2 #(
		.INIT('h1)
	) name473 (
		\a[60] ,
		\b[60] ,
		_w730_
	);
	LUT2 #(
		.INIT('h8)
	) name474 (
		\a[60] ,
		\b[60] ,
		_w731_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w730_,
		_w731_,
		_w732_
	);
	LUT2 #(
		.INIT('h1)
	) name476 (
		_w723_,
		_w726_,
		_w733_
	);
	LUT2 #(
		.INIT('h1)
	) name477 (
		_w722_,
		_w733_,
		_w734_
	);
	LUT2 #(
		.INIT('h4)
	) name478 (
		_w732_,
		_w734_,
		_w735_
	);
	LUT2 #(
		.INIT('h2)
	) name479 (
		_w732_,
		_w734_,
		_w736_
	);
	LUT2 #(
		.INIT('h1)
	) name480 (
		_w735_,
		_w736_,
		_w737_
	);
	LUT2 #(
		.INIT('h1)
	) name481 (
		\a[61] ,
		\b[61] ,
		_w738_
	);
	LUT2 #(
		.INIT('h8)
	) name482 (
		\a[61] ,
		\b[61] ,
		_w739_
	);
	LUT2 #(
		.INIT('h1)
	) name483 (
		_w738_,
		_w739_,
		_w740_
	);
	LUT2 #(
		.INIT('h1)
	) name484 (
		_w731_,
		_w734_,
		_w741_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w730_,
		_w741_,
		_w742_
	);
	LUT2 #(
		.INIT('h4)
	) name486 (
		_w740_,
		_w742_,
		_w743_
	);
	LUT2 #(
		.INIT('h2)
	) name487 (
		_w740_,
		_w742_,
		_w744_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w743_,
		_w744_,
		_w745_
	);
	LUT2 #(
		.INIT('h1)
	) name489 (
		\a[62] ,
		\b[62] ,
		_w746_
	);
	LUT2 #(
		.INIT('h8)
	) name490 (
		\a[62] ,
		\b[62] ,
		_w747_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w746_,
		_w747_,
		_w748_
	);
	LUT2 #(
		.INIT('h1)
	) name492 (
		_w739_,
		_w742_,
		_w749_
	);
	LUT2 #(
		.INIT('h1)
	) name493 (
		_w738_,
		_w749_,
		_w750_
	);
	LUT2 #(
		.INIT('h4)
	) name494 (
		_w748_,
		_w750_,
		_w751_
	);
	LUT2 #(
		.INIT('h2)
	) name495 (
		_w748_,
		_w750_,
		_w752_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w751_,
		_w752_,
		_w753_
	);
	LUT2 #(
		.INIT('h1)
	) name497 (
		\a[63] ,
		\b[63] ,
		_w754_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\a[63] ,
		\b[63] ,
		_w755_
	);
	LUT2 #(
		.INIT('h1)
	) name499 (
		_w754_,
		_w755_,
		_w756_
	);
	LUT2 #(
		.INIT('h1)
	) name500 (
		_w747_,
		_w750_,
		_w757_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w746_,
		_w757_,
		_w758_
	);
	LUT2 #(
		.INIT('h4)
	) name502 (
		_w756_,
		_w758_,
		_w759_
	);
	LUT2 #(
		.INIT('h2)
	) name503 (
		_w756_,
		_w758_,
		_w760_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w759_,
		_w760_,
		_w761_
	);
	LUT2 #(
		.INIT('h1)
	) name505 (
		\a[64] ,
		\b[64] ,
		_w762_
	);
	LUT2 #(
		.INIT('h8)
	) name506 (
		\a[64] ,
		\b[64] ,
		_w763_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w762_,
		_w763_,
		_w764_
	);
	LUT2 #(
		.INIT('h1)
	) name508 (
		_w755_,
		_w758_,
		_w765_
	);
	LUT2 #(
		.INIT('h1)
	) name509 (
		_w754_,
		_w765_,
		_w766_
	);
	LUT2 #(
		.INIT('h4)
	) name510 (
		_w764_,
		_w766_,
		_w767_
	);
	LUT2 #(
		.INIT('h2)
	) name511 (
		_w764_,
		_w766_,
		_w768_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w767_,
		_w768_,
		_w769_
	);
	LUT2 #(
		.INIT('h1)
	) name513 (
		\a[65] ,
		\b[65] ,
		_w770_
	);
	LUT2 #(
		.INIT('h8)
	) name514 (
		\a[65] ,
		\b[65] ,
		_w771_
	);
	LUT2 #(
		.INIT('h1)
	) name515 (
		_w770_,
		_w771_,
		_w772_
	);
	LUT2 #(
		.INIT('h1)
	) name516 (
		_w763_,
		_w766_,
		_w773_
	);
	LUT2 #(
		.INIT('h1)
	) name517 (
		_w762_,
		_w773_,
		_w774_
	);
	LUT2 #(
		.INIT('h4)
	) name518 (
		_w772_,
		_w774_,
		_w775_
	);
	LUT2 #(
		.INIT('h2)
	) name519 (
		_w772_,
		_w774_,
		_w776_
	);
	LUT2 #(
		.INIT('h1)
	) name520 (
		_w775_,
		_w776_,
		_w777_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		\a[66] ,
		\b[66] ,
		_w778_
	);
	LUT2 #(
		.INIT('h8)
	) name522 (
		\a[66] ,
		\b[66] ,
		_w779_
	);
	LUT2 #(
		.INIT('h1)
	) name523 (
		_w778_,
		_w779_,
		_w780_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		_w771_,
		_w774_,
		_w781_
	);
	LUT2 #(
		.INIT('h1)
	) name525 (
		_w770_,
		_w781_,
		_w782_
	);
	LUT2 #(
		.INIT('h4)
	) name526 (
		_w780_,
		_w782_,
		_w783_
	);
	LUT2 #(
		.INIT('h2)
	) name527 (
		_w780_,
		_w782_,
		_w784_
	);
	LUT2 #(
		.INIT('h1)
	) name528 (
		_w783_,
		_w784_,
		_w785_
	);
	LUT2 #(
		.INIT('h1)
	) name529 (
		\a[67] ,
		\b[67] ,
		_w786_
	);
	LUT2 #(
		.INIT('h8)
	) name530 (
		\a[67] ,
		\b[67] ,
		_w787_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w786_,
		_w787_,
		_w788_
	);
	LUT2 #(
		.INIT('h1)
	) name532 (
		_w779_,
		_w782_,
		_w789_
	);
	LUT2 #(
		.INIT('h1)
	) name533 (
		_w778_,
		_w789_,
		_w790_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		_w788_,
		_w790_,
		_w791_
	);
	LUT2 #(
		.INIT('h2)
	) name535 (
		_w788_,
		_w790_,
		_w792_
	);
	LUT2 #(
		.INIT('h1)
	) name536 (
		_w791_,
		_w792_,
		_w793_
	);
	LUT2 #(
		.INIT('h1)
	) name537 (
		\a[68] ,
		\b[68] ,
		_w794_
	);
	LUT2 #(
		.INIT('h8)
	) name538 (
		\a[68] ,
		\b[68] ,
		_w795_
	);
	LUT2 #(
		.INIT('h1)
	) name539 (
		_w794_,
		_w795_,
		_w796_
	);
	LUT2 #(
		.INIT('h1)
	) name540 (
		_w787_,
		_w790_,
		_w797_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		_w786_,
		_w797_,
		_w798_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w796_,
		_w798_,
		_w799_
	);
	LUT2 #(
		.INIT('h2)
	) name543 (
		_w796_,
		_w798_,
		_w800_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		_w799_,
		_w800_,
		_w801_
	);
	LUT2 #(
		.INIT('h1)
	) name545 (
		\a[69] ,
		\b[69] ,
		_w802_
	);
	LUT2 #(
		.INIT('h8)
	) name546 (
		\a[69] ,
		\b[69] ,
		_w803_
	);
	LUT2 #(
		.INIT('h1)
	) name547 (
		_w802_,
		_w803_,
		_w804_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w795_,
		_w798_,
		_w805_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		_w794_,
		_w805_,
		_w806_
	);
	LUT2 #(
		.INIT('h4)
	) name550 (
		_w804_,
		_w806_,
		_w807_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		_w804_,
		_w806_,
		_w808_
	);
	LUT2 #(
		.INIT('h1)
	) name552 (
		_w807_,
		_w808_,
		_w809_
	);
	LUT2 #(
		.INIT('h1)
	) name553 (
		\a[70] ,
		\b[70] ,
		_w810_
	);
	LUT2 #(
		.INIT('h8)
	) name554 (
		\a[70] ,
		\b[70] ,
		_w811_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w810_,
		_w811_,
		_w812_
	);
	LUT2 #(
		.INIT('h1)
	) name556 (
		_w803_,
		_w806_,
		_w813_
	);
	LUT2 #(
		.INIT('h1)
	) name557 (
		_w802_,
		_w813_,
		_w814_
	);
	LUT2 #(
		.INIT('h4)
	) name558 (
		_w812_,
		_w814_,
		_w815_
	);
	LUT2 #(
		.INIT('h2)
	) name559 (
		_w812_,
		_w814_,
		_w816_
	);
	LUT2 #(
		.INIT('h1)
	) name560 (
		_w815_,
		_w816_,
		_w817_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		\a[71] ,
		\b[71] ,
		_w818_
	);
	LUT2 #(
		.INIT('h8)
	) name562 (
		\a[71] ,
		\b[71] ,
		_w819_
	);
	LUT2 #(
		.INIT('h1)
	) name563 (
		_w818_,
		_w819_,
		_w820_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		_w811_,
		_w814_,
		_w821_
	);
	LUT2 #(
		.INIT('h1)
	) name565 (
		_w810_,
		_w821_,
		_w822_
	);
	LUT2 #(
		.INIT('h4)
	) name566 (
		_w820_,
		_w822_,
		_w823_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		_w820_,
		_w822_,
		_w824_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w823_,
		_w824_,
		_w825_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		\a[72] ,
		\b[72] ,
		_w826_
	);
	LUT2 #(
		.INIT('h8)
	) name570 (
		\a[72] ,
		\b[72] ,
		_w827_
	);
	LUT2 #(
		.INIT('h1)
	) name571 (
		_w826_,
		_w827_,
		_w828_
	);
	LUT2 #(
		.INIT('h1)
	) name572 (
		_w819_,
		_w822_,
		_w829_
	);
	LUT2 #(
		.INIT('h1)
	) name573 (
		_w818_,
		_w829_,
		_w830_
	);
	LUT2 #(
		.INIT('h4)
	) name574 (
		_w828_,
		_w830_,
		_w831_
	);
	LUT2 #(
		.INIT('h2)
	) name575 (
		_w828_,
		_w830_,
		_w832_
	);
	LUT2 #(
		.INIT('h1)
	) name576 (
		_w831_,
		_w832_,
		_w833_
	);
	LUT2 #(
		.INIT('h1)
	) name577 (
		\a[73] ,
		\b[73] ,
		_w834_
	);
	LUT2 #(
		.INIT('h8)
	) name578 (
		\a[73] ,
		\b[73] ,
		_w835_
	);
	LUT2 #(
		.INIT('h1)
	) name579 (
		_w834_,
		_w835_,
		_w836_
	);
	LUT2 #(
		.INIT('h1)
	) name580 (
		_w827_,
		_w830_,
		_w837_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w826_,
		_w837_,
		_w838_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		_w836_,
		_w838_,
		_w839_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		_w836_,
		_w838_,
		_w840_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		_w839_,
		_w840_,
		_w841_
	);
	LUT2 #(
		.INIT('h1)
	) name585 (
		\a[74] ,
		\b[74] ,
		_w842_
	);
	LUT2 #(
		.INIT('h8)
	) name586 (
		\a[74] ,
		\b[74] ,
		_w843_
	);
	LUT2 #(
		.INIT('h1)
	) name587 (
		_w842_,
		_w843_,
		_w844_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w835_,
		_w838_,
		_w845_
	);
	LUT2 #(
		.INIT('h1)
	) name589 (
		_w834_,
		_w845_,
		_w846_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		_w844_,
		_w846_,
		_w847_
	);
	LUT2 #(
		.INIT('h2)
	) name591 (
		_w844_,
		_w846_,
		_w848_
	);
	LUT2 #(
		.INIT('h1)
	) name592 (
		_w847_,
		_w848_,
		_w849_
	);
	LUT2 #(
		.INIT('h1)
	) name593 (
		\a[75] ,
		\b[75] ,
		_w850_
	);
	LUT2 #(
		.INIT('h8)
	) name594 (
		\a[75] ,
		\b[75] ,
		_w851_
	);
	LUT2 #(
		.INIT('h1)
	) name595 (
		_w850_,
		_w851_,
		_w852_
	);
	LUT2 #(
		.INIT('h1)
	) name596 (
		_w843_,
		_w846_,
		_w853_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		_w842_,
		_w853_,
		_w854_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		_w852_,
		_w854_,
		_w855_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		_w852_,
		_w854_,
		_w856_
	);
	LUT2 #(
		.INIT('h1)
	) name600 (
		_w855_,
		_w856_,
		_w857_
	);
	LUT2 #(
		.INIT('h1)
	) name601 (
		\a[76] ,
		\b[76] ,
		_w858_
	);
	LUT2 #(
		.INIT('h8)
	) name602 (
		\a[76] ,
		\b[76] ,
		_w859_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w858_,
		_w859_,
		_w860_
	);
	LUT2 #(
		.INIT('h1)
	) name604 (
		_w851_,
		_w854_,
		_w861_
	);
	LUT2 #(
		.INIT('h1)
	) name605 (
		_w850_,
		_w861_,
		_w862_
	);
	LUT2 #(
		.INIT('h4)
	) name606 (
		_w860_,
		_w862_,
		_w863_
	);
	LUT2 #(
		.INIT('h2)
	) name607 (
		_w860_,
		_w862_,
		_w864_
	);
	LUT2 #(
		.INIT('h1)
	) name608 (
		_w863_,
		_w864_,
		_w865_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		\a[77] ,
		\b[77] ,
		_w866_
	);
	LUT2 #(
		.INIT('h8)
	) name610 (
		\a[77] ,
		\b[77] ,
		_w867_
	);
	LUT2 #(
		.INIT('h1)
	) name611 (
		_w866_,
		_w867_,
		_w868_
	);
	LUT2 #(
		.INIT('h1)
	) name612 (
		_w859_,
		_w862_,
		_w869_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		_w858_,
		_w869_,
		_w870_
	);
	LUT2 #(
		.INIT('h4)
	) name614 (
		_w868_,
		_w870_,
		_w871_
	);
	LUT2 #(
		.INIT('h2)
	) name615 (
		_w868_,
		_w870_,
		_w872_
	);
	LUT2 #(
		.INIT('h1)
	) name616 (
		_w871_,
		_w872_,
		_w873_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		\a[78] ,
		\b[78] ,
		_w874_
	);
	LUT2 #(
		.INIT('h8)
	) name618 (
		\a[78] ,
		\b[78] ,
		_w875_
	);
	LUT2 #(
		.INIT('h1)
	) name619 (
		_w874_,
		_w875_,
		_w876_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		_w867_,
		_w870_,
		_w877_
	);
	LUT2 #(
		.INIT('h1)
	) name621 (
		_w866_,
		_w877_,
		_w878_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		_w876_,
		_w878_,
		_w879_
	);
	LUT2 #(
		.INIT('h2)
	) name623 (
		_w876_,
		_w878_,
		_w880_
	);
	LUT2 #(
		.INIT('h1)
	) name624 (
		_w879_,
		_w880_,
		_w881_
	);
	LUT2 #(
		.INIT('h1)
	) name625 (
		\a[79] ,
		\b[79] ,
		_w882_
	);
	LUT2 #(
		.INIT('h8)
	) name626 (
		\a[79] ,
		\b[79] ,
		_w883_
	);
	LUT2 #(
		.INIT('h1)
	) name627 (
		_w882_,
		_w883_,
		_w884_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		_w875_,
		_w878_,
		_w885_
	);
	LUT2 #(
		.INIT('h1)
	) name629 (
		_w874_,
		_w885_,
		_w886_
	);
	LUT2 #(
		.INIT('h4)
	) name630 (
		_w884_,
		_w886_,
		_w887_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		_w884_,
		_w886_,
		_w888_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w887_,
		_w888_,
		_w889_
	);
	LUT2 #(
		.INIT('h1)
	) name633 (
		\a[80] ,
		\b[80] ,
		_w890_
	);
	LUT2 #(
		.INIT('h8)
	) name634 (
		\a[80] ,
		\b[80] ,
		_w891_
	);
	LUT2 #(
		.INIT('h1)
	) name635 (
		_w890_,
		_w891_,
		_w892_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w883_,
		_w886_,
		_w893_
	);
	LUT2 #(
		.INIT('h1)
	) name637 (
		_w882_,
		_w893_,
		_w894_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		_w892_,
		_w894_,
		_w895_
	);
	LUT2 #(
		.INIT('h2)
	) name639 (
		_w892_,
		_w894_,
		_w896_
	);
	LUT2 #(
		.INIT('h1)
	) name640 (
		_w895_,
		_w896_,
		_w897_
	);
	LUT2 #(
		.INIT('h1)
	) name641 (
		\a[81] ,
		\b[81] ,
		_w898_
	);
	LUT2 #(
		.INIT('h8)
	) name642 (
		\a[81] ,
		\b[81] ,
		_w899_
	);
	LUT2 #(
		.INIT('h1)
	) name643 (
		_w898_,
		_w899_,
		_w900_
	);
	LUT2 #(
		.INIT('h1)
	) name644 (
		_w891_,
		_w894_,
		_w901_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		_w890_,
		_w901_,
		_w902_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		_w900_,
		_w902_,
		_w903_
	);
	LUT2 #(
		.INIT('h2)
	) name647 (
		_w900_,
		_w902_,
		_w904_
	);
	LUT2 #(
		.INIT('h1)
	) name648 (
		_w903_,
		_w904_,
		_w905_
	);
	LUT2 #(
		.INIT('h1)
	) name649 (
		\a[82] ,
		\b[82] ,
		_w906_
	);
	LUT2 #(
		.INIT('h8)
	) name650 (
		\a[82] ,
		\b[82] ,
		_w907_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w906_,
		_w907_,
		_w908_
	);
	LUT2 #(
		.INIT('h1)
	) name652 (
		_w899_,
		_w902_,
		_w909_
	);
	LUT2 #(
		.INIT('h1)
	) name653 (
		_w898_,
		_w909_,
		_w910_
	);
	LUT2 #(
		.INIT('h4)
	) name654 (
		_w908_,
		_w910_,
		_w911_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		_w908_,
		_w910_,
		_w912_
	);
	LUT2 #(
		.INIT('h1)
	) name656 (
		_w911_,
		_w912_,
		_w913_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		\a[83] ,
		\b[83] ,
		_w914_
	);
	LUT2 #(
		.INIT('h8)
	) name658 (
		\a[83] ,
		\b[83] ,
		_w915_
	);
	LUT2 #(
		.INIT('h1)
	) name659 (
		_w914_,
		_w915_,
		_w916_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		_w907_,
		_w910_,
		_w917_
	);
	LUT2 #(
		.INIT('h1)
	) name661 (
		_w906_,
		_w917_,
		_w918_
	);
	LUT2 #(
		.INIT('h4)
	) name662 (
		_w916_,
		_w918_,
		_w919_
	);
	LUT2 #(
		.INIT('h2)
	) name663 (
		_w916_,
		_w918_,
		_w920_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w919_,
		_w920_,
		_w921_
	);
	LUT2 #(
		.INIT('h1)
	) name665 (
		\a[84] ,
		\b[84] ,
		_w922_
	);
	LUT2 #(
		.INIT('h8)
	) name666 (
		\a[84] ,
		\b[84] ,
		_w923_
	);
	LUT2 #(
		.INIT('h1)
	) name667 (
		_w922_,
		_w923_,
		_w924_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w915_,
		_w918_,
		_w925_
	);
	LUT2 #(
		.INIT('h1)
	) name669 (
		_w914_,
		_w925_,
		_w926_
	);
	LUT2 #(
		.INIT('h4)
	) name670 (
		_w924_,
		_w926_,
		_w927_
	);
	LUT2 #(
		.INIT('h2)
	) name671 (
		_w924_,
		_w926_,
		_w928_
	);
	LUT2 #(
		.INIT('h1)
	) name672 (
		_w927_,
		_w928_,
		_w929_
	);
	LUT2 #(
		.INIT('h1)
	) name673 (
		\a[85] ,
		\b[85] ,
		_w930_
	);
	LUT2 #(
		.INIT('h8)
	) name674 (
		\a[85] ,
		\b[85] ,
		_w931_
	);
	LUT2 #(
		.INIT('h1)
	) name675 (
		_w930_,
		_w931_,
		_w932_
	);
	LUT2 #(
		.INIT('h1)
	) name676 (
		_w923_,
		_w926_,
		_w933_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		_w922_,
		_w933_,
		_w934_
	);
	LUT2 #(
		.INIT('h4)
	) name678 (
		_w932_,
		_w934_,
		_w935_
	);
	LUT2 #(
		.INIT('h2)
	) name679 (
		_w932_,
		_w934_,
		_w936_
	);
	LUT2 #(
		.INIT('h1)
	) name680 (
		_w935_,
		_w936_,
		_w937_
	);
	LUT2 #(
		.INIT('h1)
	) name681 (
		\a[86] ,
		\b[86] ,
		_w938_
	);
	LUT2 #(
		.INIT('h8)
	) name682 (
		\a[86] ,
		\b[86] ,
		_w939_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w938_,
		_w939_,
		_w940_
	);
	LUT2 #(
		.INIT('h1)
	) name684 (
		_w931_,
		_w934_,
		_w941_
	);
	LUT2 #(
		.INIT('h1)
	) name685 (
		_w930_,
		_w941_,
		_w942_
	);
	LUT2 #(
		.INIT('h4)
	) name686 (
		_w940_,
		_w942_,
		_w943_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		_w940_,
		_w942_,
		_w944_
	);
	LUT2 #(
		.INIT('h1)
	) name688 (
		_w943_,
		_w944_,
		_w945_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		\a[87] ,
		\b[87] ,
		_w946_
	);
	LUT2 #(
		.INIT('h8)
	) name690 (
		\a[87] ,
		\b[87] ,
		_w947_
	);
	LUT2 #(
		.INIT('h1)
	) name691 (
		_w946_,
		_w947_,
		_w948_
	);
	LUT2 #(
		.INIT('h1)
	) name692 (
		_w939_,
		_w942_,
		_w949_
	);
	LUT2 #(
		.INIT('h1)
	) name693 (
		_w938_,
		_w949_,
		_w950_
	);
	LUT2 #(
		.INIT('h4)
	) name694 (
		_w948_,
		_w950_,
		_w951_
	);
	LUT2 #(
		.INIT('h2)
	) name695 (
		_w948_,
		_w950_,
		_w952_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w951_,
		_w952_,
		_w953_
	);
	LUT2 #(
		.INIT('h1)
	) name697 (
		\a[88] ,
		\b[88] ,
		_w954_
	);
	LUT2 #(
		.INIT('h8)
	) name698 (
		\a[88] ,
		\b[88] ,
		_w955_
	);
	LUT2 #(
		.INIT('h1)
	) name699 (
		_w954_,
		_w955_,
		_w956_
	);
	LUT2 #(
		.INIT('h1)
	) name700 (
		_w947_,
		_w950_,
		_w957_
	);
	LUT2 #(
		.INIT('h1)
	) name701 (
		_w946_,
		_w957_,
		_w958_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		_w956_,
		_w958_,
		_w959_
	);
	LUT2 #(
		.INIT('h2)
	) name703 (
		_w956_,
		_w958_,
		_w960_
	);
	LUT2 #(
		.INIT('h1)
	) name704 (
		_w959_,
		_w960_,
		_w961_
	);
	LUT2 #(
		.INIT('h1)
	) name705 (
		\a[89] ,
		\b[89] ,
		_w962_
	);
	LUT2 #(
		.INIT('h8)
	) name706 (
		\a[89] ,
		\b[89] ,
		_w963_
	);
	LUT2 #(
		.INIT('h1)
	) name707 (
		_w962_,
		_w963_,
		_w964_
	);
	LUT2 #(
		.INIT('h1)
	) name708 (
		_w955_,
		_w958_,
		_w965_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		_w954_,
		_w965_,
		_w966_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		_w964_,
		_w966_,
		_w967_
	);
	LUT2 #(
		.INIT('h2)
	) name711 (
		_w964_,
		_w966_,
		_w968_
	);
	LUT2 #(
		.INIT('h1)
	) name712 (
		_w967_,
		_w968_,
		_w969_
	);
	LUT2 #(
		.INIT('h1)
	) name713 (
		\a[90] ,
		\b[90] ,
		_w970_
	);
	LUT2 #(
		.INIT('h8)
	) name714 (
		\a[90] ,
		\b[90] ,
		_w971_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w970_,
		_w971_,
		_w972_
	);
	LUT2 #(
		.INIT('h1)
	) name716 (
		_w963_,
		_w966_,
		_w973_
	);
	LUT2 #(
		.INIT('h1)
	) name717 (
		_w962_,
		_w973_,
		_w974_
	);
	LUT2 #(
		.INIT('h4)
	) name718 (
		_w972_,
		_w974_,
		_w975_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		_w972_,
		_w974_,
		_w976_
	);
	LUT2 #(
		.INIT('h1)
	) name720 (
		_w975_,
		_w976_,
		_w977_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		\a[91] ,
		\b[91] ,
		_w978_
	);
	LUT2 #(
		.INIT('h8)
	) name722 (
		\a[91] ,
		\b[91] ,
		_w979_
	);
	LUT2 #(
		.INIT('h1)
	) name723 (
		_w978_,
		_w979_,
		_w980_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		_w971_,
		_w974_,
		_w981_
	);
	LUT2 #(
		.INIT('h1)
	) name725 (
		_w970_,
		_w981_,
		_w982_
	);
	LUT2 #(
		.INIT('h4)
	) name726 (
		_w980_,
		_w982_,
		_w983_
	);
	LUT2 #(
		.INIT('h2)
	) name727 (
		_w980_,
		_w982_,
		_w984_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		_w983_,
		_w984_,
		_w985_
	);
	LUT2 #(
		.INIT('h1)
	) name729 (
		\a[92] ,
		\b[92] ,
		_w986_
	);
	LUT2 #(
		.INIT('h8)
	) name730 (
		\a[92] ,
		\b[92] ,
		_w987_
	);
	LUT2 #(
		.INIT('h1)
	) name731 (
		_w986_,
		_w987_,
		_w988_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w979_,
		_w982_,
		_w989_
	);
	LUT2 #(
		.INIT('h1)
	) name733 (
		_w978_,
		_w989_,
		_w990_
	);
	LUT2 #(
		.INIT('h4)
	) name734 (
		_w988_,
		_w990_,
		_w991_
	);
	LUT2 #(
		.INIT('h2)
	) name735 (
		_w988_,
		_w990_,
		_w992_
	);
	LUT2 #(
		.INIT('h1)
	) name736 (
		_w991_,
		_w992_,
		_w993_
	);
	LUT2 #(
		.INIT('h1)
	) name737 (
		\a[93] ,
		\b[93] ,
		_w994_
	);
	LUT2 #(
		.INIT('h8)
	) name738 (
		\a[93] ,
		\b[93] ,
		_w995_
	);
	LUT2 #(
		.INIT('h1)
	) name739 (
		_w994_,
		_w995_,
		_w996_
	);
	LUT2 #(
		.INIT('h1)
	) name740 (
		_w987_,
		_w990_,
		_w997_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		_w986_,
		_w997_,
		_w998_
	);
	LUT2 #(
		.INIT('h4)
	) name742 (
		_w996_,
		_w998_,
		_w999_
	);
	LUT2 #(
		.INIT('h2)
	) name743 (
		_w996_,
		_w998_,
		_w1000_
	);
	LUT2 #(
		.INIT('h1)
	) name744 (
		_w999_,
		_w1000_,
		_w1001_
	);
	LUT2 #(
		.INIT('h1)
	) name745 (
		\a[94] ,
		\b[94] ,
		_w1002_
	);
	LUT2 #(
		.INIT('h8)
	) name746 (
		\a[94] ,
		\b[94] ,
		_w1003_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w1002_,
		_w1003_,
		_w1004_
	);
	LUT2 #(
		.INIT('h1)
	) name748 (
		_w995_,
		_w998_,
		_w1005_
	);
	LUT2 #(
		.INIT('h1)
	) name749 (
		_w994_,
		_w1005_,
		_w1006_
	);
	LUT2 #(
		.INIT('h4)
	) name750 (
		_w1004_,
		_w1006_,
		_w1007_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		_w1004_,
		_w1006_,
		_w1008_
	);
	LUT2 #(
		.INIT('h1)
	) name752 (
		_w1007_,
		_w1008_,
		_w1009_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		\a[95] ,
		\b[95] ,
		_w1010_
	);
	LUT2 #(
		.INIT('h8)
	) name754 (
		\a[95] ,
		\b[95] ,
		_w1011_
	);
	LUT2 #(
		.INIT('h1)
	) name755 (
		_w1010_,
		_w1011_,
		_w1012_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		_w1003_,
		_w1006_,
		_w1013_
	);
	LUT2 #(
		.INIT('h1)
	) name757 (
		_w1002_,
		_w1013_,
		_w1014_
	);
	LUT2 #(
		.INIT('h4)
	) name758 (
		_w1012_,
		_w1014_,
		_w1015_
	);
	LUT2 #(
		.INIT('h2)
	) name759 (
		_w1012_,
		_w1014_,
		_w1016_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w1015_,
		_w1016_,
		_w1017_
	);
	LUT2 #(
		.INIT('h1)
	) name761 (
		\a[96] ,
		\b[96] ,
		_w1018_
	);
	LUT2 #(
		.INIT('h8)
	) name762 (
		\a[96] ,
		\b[96] ,
		_w1019_
	);
	LUT2 #(
		.INIT('h1)
	) name763 (
		_w1018_,
		_w1019_,
		_w1020_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w1011_,
		_w1014_,
		_w1021_
	);
	LUT2 #(
		.INIT('h1)
	) name765 (
		_w1010_,
		_w1021_,
		_w1022_
	);
	LUT2 #(
		.INIT('h4)
	) name766 (
		_w1020_,
		_w1022_,
		_w1023_
	);
	LUT2 #(
		.INIT('h2)
	) name767 (
		_w1020_,
		_w1022_,
		_w1024_
	);
	LUT2 #(
		.INIT('h1)
	) name768 (
		_w1023_,
		_w1024_,
		_w1025_
	);
	LUT2 #(
		.INIT('h1)
	) name769 (
		\a[97] ,
		\b[97] ,
		_w1026_
	);
	LUT2 #(
		.INIT('h8)
	) name770 (
		\a[97] ,
		\b[97] ,
		_w1027_
	);
	LUT2 #(
		.INIT('h1)
	) name771 (
		_w1026_,
		_w1027_,
		_w1028_
	);
	LUT2 #(
		.INIT('h1)
	) name772 (
		_w1019_,
		_w1022_,
		_w1029_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		_w1018_,
		_w1029_,
		_w1030_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		_w1028_,
		_w1030_,
		_w1031_
	);
	LUT2 #(
		.INIT('h2)
	) name775 (
		_w1028_,
		_w1030_,
		_w1032_
	);
	LUT2 #(
		.INIT('h1)
	) name776 (
		_w1031_,
		_w1032_,
		_w1033_
	);
	LUT2 #(
		.INIT('h1)
	) name777 (
		\a[98] ,
		\b[98] ,
		_w1034_
	);
	LUT2 #(
		.INIT('h8)
	) name778 (
		\a[98] ,
		\b[98] ,
		_w1035_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		_w1034_,
		_w1035_,
		_w1036_
	);
	LUT2 #(
		.INIT('h1)
	) name780 (
		_w1027_,
		_w1030_,
		_w1037_
	);
	LUT2 #(
		.INIT('h1)
	) name781 (
		_w1026_,
		_w1037_,
		_w1038_
	);
	LUT2 #(
		.INIT('h4)
	) name782 (
		_w1036_,
		_w1038_,
		_w1039_
	);
	LUT2 #(
		.INIT('h2)
	) name783 (
		_w1036_,
		_w1038_,
		_w1040_
	);
	LUT2 #(
		.INIT('h1)
	) name784 (
		_w1039_,
		_w1040_,
		_w1041_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		\a[99] ,
		\b[99] ,
		_w1042_
	);
	LUT2 #(
		.INIT('h8)
	) name786 (
		\a[99] ,
		\b[99] ,
		_w1043_
	);
	LUT2 #(
		.INIT('h1)
	) name787 (
		_w1042_,
		_w1043_,
		_w1044_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		_w1035_,
		_w1038_,
		_w1045_
	);
	LUT2 #(
		.INIT('h1)
	) name789 (
		_w1034_,
		_w1045_,
		_w1046_
	);
	LUT2 #(
		.INIT('h4)
	) name790 (
		_w1044_,
		_w1046_,
		_w1047_
	);
	LUT2 #(
		.INIT('h2)
	) name791 (
		_w1044_,
		_w1046_,
		_w1048_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w1047_,
		_w1048_,
		_w1049_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		\a[100] ,
		\b[100] ,
		_w1050_
	);
	LUT2 #(
		.INIT('h8)
	) name794 (
		\a[100] ,
		\b[100] ,
		_w1051_
	);
	LUT2 #(
		.INIT('h1)
	) name795 (
		_w1050_,
		_w1051_,
		_w1052_
	);
	LUT2 #(
		.INIT('h1)
	) name796 (
		_w1043_,
		_w1046_,
		_w1053_
	);
	LUT2 #(
		.INIT('h1)
	) name797 (
		_w1042_,
		_w1053_,
		_w1054_
	);
	LUT2 #(
		.INIT('h4)
	) name798 (
		_w1052_,
		_w1054_,
		_w1055_
	);
	LUT2 #(
		.INIT('h2)
	) name799 (
		_w1052_,
		_w1054_,
		_w1056_
	);
	LUT2 #(
		.INIT('h1)
	) name800 (
		_w1055_,
		_w1056_,
		_w1057_
	);
	LUT2 #(
		.INIT('h1)
	) name801 (
		\a[101] ,
		\b[101] ,
		_w1058_
	);
	LUT2 #(
		.INIT('h8)
	) name802 (
		\a[101] ,
		\b[101] ,
		_w1059_
	);
	LUT2 #(
		.INIT('h1)
	) name803 (
		_w1058_,
		_w1059_,
		_w1060_
	);
	LUT2 #(
		.INIT('h1)
	) name804 (
		_w1051_,
		_w1054_,
		_w1061_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		_w1050_,
		_w1061_,
		_w1062_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		_w1060_,
		_w1062_,
		_w1063_
	);
	LUT2 #(
		.INIT('h2)
	) name807 (
		_w1060_,
		_w1062_,
		_w1064_
	);
	LUT2 #(
		.INIT('h1)
	) name808 (
		_w1063_,
		_w1064_,
		_w1065_
	);
	LUT2 #(
		.INIT('h1)
	) name809 (
		\a[102] ,
		\b[102] ,
		_w1066_
	);
	LUT2 #(
		.INIT('h8)
	) name810 (
		\a[102] ,
		\b[102] ,
		_w1067_
	);
	LUT2 #(
		.INIT('h1)
	) name811 (
		_w1066_,
		_w1067_,
		_w1068_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w1059_,
		_w1062_,
		_w1069_
	);
	LUT2 #(
		.INIT('h1)
	) name813 (
		_w1058_,
		_w1069_,
		_w1070_
	);
	LUT2 #(
		.INIT('h4)
	) name814 (
		_w1068_,
		_w1070_,
		_w1071_
	);
	LUT2 #(
		.INIT('h2)
	) name815 (
		_w1068_,
		_w1070_,
		_w1072_
	);
	LUT2 #(
		.INIT('h1)
	) name816 (
		_w1071_,
		_w1072_,
		_w1073_
	);
	LUT2 #(
		.INIT('h1)
	) name817 (
		\a[103] ,
		\b[103] ,
		_w1074_
	);
	LUT2 #(
		.INIT('h8)
	) name818 (
		\a[103] ,
		\b[103] ,
		_w1075_
	);
	LUT2 #(
		.INIT('h1)
	) name819 (
		_w1074_,
		_w1075_,
		_w1076_
	);
	LUT2 #(
		.INIT('h1)
	) name820 (
		_w1067_,
		_w1070_,
		_w1077_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w1066_,
		_w1077_,
		_w1078_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		_w1076_,
		_w1078_,
		_w1079_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		_w1076_,
		_w1078_,
		_w1080_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		_w1079_,
		_w1080_,
		_w1081_
	);
	LUT2 #(
		.INIT('h1)
	) name825 (
		\a[104] ,
		\b[104] ,
		_w1082_
	);
	LUT2 #(
		.INIT('h8)
	) name826 (
		\a[104] ,
		\b[104] ,
		_w1083_
	);
	LUT2 #(
		.INIT('h1)
	) name827 (
		_w1082_,
		_w1083_,
		_w1084_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		_w1075_,
		_w1078_,
		_w1085_
	);
	LUT2 #(
		.INIT('h1)
	) name829 (
		_w1074_,
		_w1085_,
		_w1086_
	);
	LUT2 #(
		.INIT('h4)
	) name830 (
		_w1084_,
		_w1086_,
		_w1087_
	);
	LUT2 #(
		.INIT('h2)
	) name831 (
		_w1084_,
		_w1086_,
		_w1088_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		_w1087_,
		_w1088_,
		_w1089_
	);
	LUT2 #(
		.INIT('h1)
	) name833 (
		\a[105] ,
		\b[105] ,
		_w1090_
	);
	LUT2 #(
		.INIT('h8)
	) name834 (
		\a[105] ,
		\b[105] ,
		_w1091_
	);
	LUT2 #(
		.INIT('h1)
	) name835 (
		_w1090_,
		_w1091_,
		_w1092_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w1083_,
		_w1086_,
		_w1093_
	);
	LUT2 #(
		.INIT('h1)
	) name837 (
		_w1082_,
		_w1093_,
		_w1094_
	);
	LUT2 #(
		.INIT('h4)
	) name838 (
		_w1092_,
		_w1094_,
		_w1095_
	);
	LUT2 #(
		.INIT('h2)
	) name839 (
		_w1092_,
		_w1094_,
		_w1096_
	);
	LUT2 #(
		.INIT('h1)
	) name840 (
		_w1095_,
		_w1096_,
		_w1097_
	);
	LUT2 #(
		.INIT('h1)
	) name841 (
		\a[106] ,
		\b[106] ,
		_w1098_
	);
	LUT2 #(
		.INIT('h8)
	) name842 (
		\a[106] ,
		\b[106] ,
		_w1099_
	);
	LUT2 #(
		.INIT('h1)
	) name843 (
		_w1098_,
		_w1099_,
		_w1100_
	);
	LUT2 #(
		.INIT('h1)
	) name844 (
		_w1091_,
		_w1094_,
		_w1101_
	);
	LUT2 #(
		.INIT('h1)
	) name845 (
		_w1090_,
		_w1101_,
		_w1102_
	);
	LUT2 #(
		.INIT('h4)
	) name846 (
		_w1100_,
		_w1102_,
		_w1103_
	);
	LUT2 #(
		.INIT('h2)
	) name847 (
		_w1100_,
		_w1102_,
		_w1104_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w1103_,
		_w1104_,
		_w1105_
	);
	LUT2 #(
		.INIT('h1)
	) name849 (
		\a[107] ,
		\b[107] ,
		_w1106_
	);
	LUT2 #(
		.INIT('h8)
	) name850 (
		\a[107] ,
		\b[107] ,
		_w1107_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w1106_,
		_w1107_,
		_w1108_
	);
	LUT2 #(
		.INIT('h1)
	) name852 (
		_w1099_,
		_w1102_,
		_w1109_
	);
	LUT2 #(
		.INIT('h1)
	) name853 (
		_w1098_,
		_w1109_,
		_w1110_
	);
	LUT2 #(
		.INIT('h4)
	) name854 (
		_w1108_,
		_w1110_,
		_w1111_
	);
	LUT2 #(
		.INIT('h2)
	) name855 (
		_w1108_,
		_w1110_,
		_w1112_
	);
	LUT2 #(
		.INIT('h1)
	) name856 (
		_w1111_,
		_w1112_,
		_w1113_
	);
	LUT2 #(
		.INIT('h1)
	) name857 (
		\a[108] ,
		\b[108] ,
		_w1114_
	);
	LUT2 #(
		.INIT('h8)
	) name858 (
		\a[108] ,
		\b[108] ,
		_w1115_
	);
	LUT2 #(
		.INIT('h1)
	) name859 (
		_w1114_,
		_w1115_,
		_w1116_
	);
	LUT2 #(
		.INIT('h1)
	) name860 (
		_w1107_,
		_w1110_,
		_w1117_
	);
	LUT2 #(
		.INIT('h1)
	) name861 (
		_w1106_,
		_w1117_,
		_w1118_
	);
	LUT2 #(
		.INIT('h4)
	) name862 (
		_w1116_,
		_w1118_,
		_w1119_
	);
	LUT2 #(
		.INIT('h2)
	) name863 (
		_w1116_,
		_w1118_,
		_w1120_
	);
	LUT2 #(
		.INIT('h1)
	) name864 (
		_w1119_,
		_w1120_,
		_w1121_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		\a[109] ,
		\b[109] ,
		_w1122_
	);
	LUT2 #(
		.INIT('h8)
	) name866 (
		\a[109] ,
		\b[109] ,
		_w1123_
	);
	LUT2 #(
		.INIT('h1)
	) name867 (
		_w1122_,
		_w1123_,
		_w1124_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w1115_,
		_w1118_,
		_w1125_
	);
	LUT2 #(
		.INIT('h1)
	) name869 (
		_w1114_,
		_w1125_,
		_w1126_
	);
	LUT2 #(
		.INIT('h4)
	) name870 (
		_w1124_,
		_w1126_,
		_w1127_
	);
	LUT2 #(
		.INIT('h2)
	) name871 (
		_w1124_,
		_w1126_,
		_w1128_
	);
	LUT2 #(
		.INIT('h1)
	) name872 (
		_w1127_,
		_w1128_,
		_w1129_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		\a[110] ,
		\b[110] ,
		_w1130_
	);
	LUT2 #(
		.INIT('h8)
	) name874 (
		\a[110] ,
		\b[110] ,
		_w1131_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		_w1130_,
		_w1131_,
		_w1132_
	);
	LUT2 #(
		.INIT('h1)
	) name876 (
		_w1123_,
		_w1126_,
		_w1133_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w1122_,
		_w1133_,
		_w1134_
	);
	LUT2 #(
		.INIT('h4)
	) name878 (
		_w1132_,
		_w1134_,
		_w1135_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		_w1132_,
		_w1134_,
		_w1136_
	);
	LUT2 #(
		.INIT('h1)
	) name880 (
		_w1135_,
		_w1136_,
		_w1137_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		\a[111] ,
		\b[111] ,
		_w1138_
	);
	LUT2 #(
		.INIT('h8)
	) name882 (
		\a[111] ,
		\b[111] ,
		_w1139_
	);
	LUT2 #(
		.INIT('h1)
	) name883 (
		_w1138_,
		_w1139_,
		_w1140_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w1131_,
		_w1134_,
		_w1141_
	);
	LUT2 #(
		.INIT('h1)
	) name885 (
		_w1130_,
		_w1141_,
		_w1142_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		_w1140_,
		_w1142_,
		_w1143_
	);
	LUT2 #(
		.INIT('h2)
	) name887 (
		_w1140_,
		_w1142_,
		_w1144_
	);
	LUT2 #(
		.INIT('h1)
	) name888 (
		_w1143_,
		_w1144_,
		_w1145_
	);
	LUT2 #(
		.INIT('h1)
	) name889 (
		\a[112] ,
		\b[112] ,
		_w1146_
	);
	LUT2 #(
		.INIT('h8)
	) name890 (
		\a[112] ,
		\b[112] ,
		_w1147_
	);
	LUT2 #(
		.INIT('h1)
	) name891 (
		_w1146_,
		_w1147_,
		_w1148_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w1139_,
		_w1142_,
		_w1149_
	);
	LUT2 #(
		.INIT('h1)
	) name893 (
		_w1138_,
		_w1149_,
		_w1150_
	);
	LUT2 #(
		.INIT('h4)
	) name894 (
		_w1148_,
		_w1150_,
		_w1151_
	);
	LUT2 #(
		.INIT('h2)
	) name895 (
		_w1148_,
		_w1150_,
		_w1152_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w1151_,
		_w1152_,
		_w1153_
	);
	LUT2 #(
		.INIT('h1)
	) name897 (
		\a[113] ,
		\b[113] ,
		_w1154_
	);
	LUT2 #(
		.INIT('h8)
	) name898 (
		\a[113] ,
		\b[113] ,
		_w1155_
	);
	LUT2 #(
		.INIT('h1)
	) name899 (
		_w1154_,
		_w1155_,
		_w1156_
	);
	LUT2 #(
		.INIT('h1)
	) name900 (
		_w1147_,
		_w1150_,
		_w1157_
	);
	LUT2 #(
		.INIT('h1)
	) name901 (
		_w1146_,
		_w1157_,
		_w1158_
	);
	LUT2 #(
		.INIT('h4)
	) name902 (
		_w1156_,
		_w1158_,
		_w1159_
	);
	LUT2 #(
		.INIT('h2)
	) name903 (
		_w1156_,
		_w1158_,
		_w1160_
	);
	LUT2 #(
		.INIT('h1)
	) name904 (
		_w1159_,
		_w1160_,
		_w1161_
	);
	LUT2 #(
		.INIT('h1)
	) name905 (
		\a[114] ,
		\b[114] ,
		_w1162_
	);
	LUT2 #(
		.INIT('h8)
	) name906 (
		\a[114] ,
		\b[114] ,
		_w1163_
	);
	LUT2 #(
		.INIT('h1)
	) name907 (
		_w1162_,
		_w1163_,
		_w1164_
	);
	LUT2 #(
		.INIT('h1)
	) name908 (
		_w1155_,
		_w1158_,
		_w1165_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		_w1154_,
		_w1165_,
		_w1166_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		_w1164_,
		_w1166_,
		_w1167_
	);
	LUT2 #(
		.INIT('h2)
	) name911 (
		_w1164_,
		_w1166_,
		_w1168_
	);
	LUT2 #(
		.INIT('h1)
	) name912 (
		_w1167_,
		_w1168_,
		_w1169_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		\a[115] ,
		\b[115] ,
		_w1170_
	);
	LUT2 #(
		.INIT('h8)
	) name914 (
		\a[115] ,
		\b[115] ,
		_w1171_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w1170_,
		_w1171_,
		_w1172_
	);
	LUT2 #(
		.INIT('h1)
	) name916 (
		_w1163_,
		_w1166_,
		_w1173_
	);
	LUT2 #(
		.INIT('h1)
	) name917 (
		_w1162_,
		_w1173_,
		_w1174_
	);
	LUT2 #(
		.INIT('h4)
	) name918 (
		_w1172_,
		_w1174_,
		_w1175_
	);
	LUT2 #(
		.INIT('h2)
	) name919 (
		_w1172_,
		_w1174_,
		_w1176_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w1175_,
		_w1176_,
		_w1177_
	);
	LUT2 #(
		.INIT('h1)
	) name921 (
		\a[116] ,
		\b[116] ,
		_w1178_
	);
	LUT2 #(
		.INIT('h8)
	) name922 (
		\a[116] ,
		\b[116] ,
		_w1179_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		_w1178_,
		_w1179_,
		_w1180_
	);
	LUT2 #(
		.INIT('h1)
	) name924 (
		_w1171_,
		_w1174_,
		_w1181_
	);
	LUT2 #(
		.INIT('h1)
	) name925 (
		_w1170_,
		_w1181_,
		_w1182_
	);
	LUT2 #(
		.INIT('h4)
	) name926 (
		_w1180_,
		_w1182_,
		_w1183_
	);
	LUT2 #(
		.INIT('h2)
	) name927 (
		_w1180_,
		_w1182_,
		_w1184_
	);
	LUT2 #(
		.INIT('h1)
	) name928 (
		_w1183_,
		_w1184_,
		_w1185_
	);
	LUT2 #(
		.INIT('h1)
	) name929 (
		\a[117] ,
		\b[117] ,
		_w1186_
	);
	LUT2 #(
		.INIT('h8)
	) name930 (
		\a[117] ,
		\b[117] ,
		_w1187_
	);
	LUT2 #(
		.INIT('h1)
	) name931 (
		_w1186_,
		_w1187_,
		_w1188_
	);
	LUT2 #(
		.INIT('h1)
	) name932 (
		_w1179_,
		_w1182_,
		_w1189_
	);
	LUT2 #(
		.INIT('h1)
	) name933 (
		_w1178_,
		_w1189_,
		_w1190_
	);
	LUT2 #(
		.INIT('h4)
	) name934 (
		_w1188_,
		_w1190_,
		_w1191_
	);
	LUT2 #(
		.INIT('h2)
	) name935 (
		_w1188_,
		_w1190_,
		_w1192_
	);
	LUT2 #(
		.INIT('h1)
	) name936 (
		_w1191_,
		_w1192_,
		_w1193_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		\a[118] ,
		\b[118] ,
		_w1194_
	);
	LUT2 #(
		.INIT('h8)
	) name938 (
		\a[118] ,
		\b[118] ,
		_w1195_
	);
	LUT2 #(
		.INIT('h1)
	) name939 (
		_w1194_,
		_w1195_,
		_w1196_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w1187_,
		_w1190_,
		_w1197_
	);
	LUT2 #(
		.INIT('h1)
	) name941 (
		_w1186_,
		_w1197_,
		_w1198_
	);
	LUT2 #(
		.INIT('h4)
	) name942 (
		_w1196_,
		_w1198_,
		_w1199_
	);
	LUT2 #(
		.INIT('h2)
	) name943 (
		_w1196_,
		_w1198_,
		_w1200_
	);
	LUT2 #(
		.INIT('h1)
	) name944 (
		_w1199_,
		_w1200_,
		_w1201_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		\a[119] ,
		\b[119] ,
		_w1202_
	);
	LUT2 #(
		.INIT('h8)
	) name946 (
		\a[119] ,
		\b[119] ,
		_w1203_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w1202_,
		_w1203_,
		_w1204_
	);
	LUT2 #(
		.INIT('h1)
	) name948 (
		_w1195_,
		_w1198_,
		_w1205_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w1194_,
		_w1205_,
		_w1206_
	);
	LUT2 #(
		.INIT('h4)
	) name950 (
		_w1204_,
		_w1206_,
		_w1207_
	);
	LUT2 #(
		.INIT('h2)
	) name951 (
		_w1204_,
		_w1206_,
		_w1208_
	);
	LUT2 #(
		.INIT('h1)
	) name952 (
		_w1207_,
		_w1208_,
		_w1209_
	);
	LUT2 #(
		.INIT('h1)
	) name953 (
		\a[120] ,
		\b[120] ,
		_w1210_
	);
	LUT2 #(
		.INIT('h8)
	) name954 (
		\a[120] ,
		\b[120] ,
		_w1211_
	);
	LUT2 #(
		.INIT('h1)
	) name955 (
		_w1210_,
		_w1211_,
		_w1212_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		_w1203_,
		_w1206_,
		_w1213_
	);
	LUT2 #(
		.INIT('h1)
	) name957 (
		_w1202_,
		_w1213_,
		_w1214_
	);
	LUT2 #(
		.INIT('h4)
	) name958 (
		_w1212_,
		_w1214_,
		_w1215_
	);
	LUT2 #(
		.INIT('h2)
	) name959 (
		_w1212_,
		_w1214_,
		_w1216_
	);
	LUT2 #(
		.INIT('h1)
	) name960 (
		_w1215_,
		_w1216_,
		_w1217_
	);
	LUT2 #(
		.INIT('h1)
	) name961 (
		\a[121] ,
		\b[121] ,
		_w1218_
	);
	LUT2 #(
		.INIT('h8)
	) name962 (
		\a[121] ,
		\b[121] ,
		_w1219_
	);
	LUT2 #(
		.INIT('h1)
	) name963 (
		_w1218_,
		_w1219_,
		_w1220_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		_w1211_,
		_w1214_,
		_w1221_
	);
	LUT2 #(
		.INIT('h1)
	) name965 (
		_w1210_,
		_w1221_,
		_w1222_
	);
	LUT2 #(
		.INIT('h4)
	) name966 (
		_w1220_,
		_w1222_,
		_w1223_
	);
	LUT2 #(
		.INIT('h2)
	) name967 (
		_w1220_,
		_w1222_,
		_w1224_
	);
	LUT2 #(
		.INIT('h1)
	) name968 (
		_w1223_,
		_w1224_,
		_w1225_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		\a[122] ,
		\b[122] ,
		_w1226_
	);
	LUT2 #(
		.INIT('h8)
	) name970 (
		\a[122] ,
		\b[122] ,
		_w1227_
	);
	LUT2 #(
		.INIT('h1)
	) name971 (
		_w1226_,
		_w1227_,
		_w1228_
	);
	LUT2 #(
		.INIT('h1)
	) name972 (
		_w1219_,
		_w1222_,
		_w1229_
	);
	LUT2 #(
		.INIT('h1)
	) name973 (
		_w1218_,
		_w1229_,
		_w1230_
	);
	LUT2 #(
		.INIT('h4)
	) name974 (
		_w1228_,
		_w1230_,
		_w1231_
	);
	LUT2 #(
		.INIT('h2)
	) name975 (
		_w1228_,
		_w1230_,
		_w1232_
	);
	LUT2 #(
		.INIT('h1)
	) name976 (
		_w1231_,
		_w1232_,
		_w1233_
	);
	LUT2 #(
		.INIT('h1)
	) name977 (
		\a[123] ,
		\b[123] ,
		_w1234_
	);
	LUT2 #(
		.INIT('h8)
	) name978 (
		\a[123] ,
		\b[123] ,
		_w1235_
	);
	LUT2 #(
		.INIT('h1)
	) name979 (
		_w1234_,
		_w1235_,
		_w1236_
	);
	LUT2 #(
		.INIT('h1)
	) name980 (
		_w1227_,
		_w1230_,
		_w1237_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w1226_,
		_w1237_,
		_w1238_
	);
	LUT2 #(
		.INIT('h4)
	) name982 (
		_w1236_,
		_w1238_,
		_w1239_
	);
	LUT2 #(
		.INIT('h2)
	) name983 (
		_w1236_,
		_w1238_,
		_w1240_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		_w1239_,
		_w1240_,
		_w1241_
	);
	LUT2 #(
		.INIT('h1)
	) name985 (
		\a[124] ,
		\b[124] ,
		_w1242_
	);
	LUT2 #(
		.INIT('h8)
	) name986 (
		\a[124] ,
		\b[124] ,
		_w1243_
	);
	LUT2 #(
		.INIT('h1)
	) name987 (
		_w1242_,
		_w1243_,
		_w1244_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w1235_,
		_w1238_,
		_w1245_
	);
	LUT2 #(
		.INIT('h1)
	) name989 (
		_w1234_,
		_w1245_,
		_w1246_
	);
	LUT2 #(
		.INIT('h4)
	) name990 (
		_w1244_,
		_w1246_,
		_w1247_
	);
	LUT2 #(
		.INIT('h2)
	) name991 (
		_w1244_,
		_w1246_,
		_w1248_
	);
	LUT2 #(
		.INIT('h1)
	) name992 (
		_w1247_,
		_w1248_,
		_w1249_
	);
	LUT2 #(
		.INIT('h1)
	) name993 (
		\a[125] ,
		\b[125] ,
		_w1250_
	);
	LUT2 #(
		.INIT('h8)
	) name994 (
		\a[125] ,
		\b[125] ,
		_w1251_
	);
	LUT2 #(
		.INIT('h1)
	) name995 (
		_w1250_,
		_w1251_,
		_w1252_
	);
	LUT2 #(
		.INIT('h1)
	) name996 (
		_w1243_,
		_w1246_,
		_w1253_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w1242_,
		_w1253_,
		_w1254_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w1252_,
		_w1254_,
		_w1255_
	);
	LUT2 #(
		.INIT('h2)
	) name999 (
		_w1252_,
		_w1254_,
		_w1256_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		_w1255_,
		_w1256_,
		_w1257_
	);
	LUT2 #(
		.INIT('h1)
	) name1001 (
		\a[126] ,
		\b[126] ,
		_w1258_
	);
	LUT2 #(
		.INIT('h8)
	) name1002 (
		\a[126] ,
		\b[126] ,
		_w1259_
	);
	LUT2 #(
		.INIT('h1)
	) name1003 (
		_w1258_,
		_w1259_,
		_w1260_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		_w1251_,
		_w1254_,
		_w1261_
	);
	LUT2 #(
		.INIT('h1)
	) name1005 (
		_w1250_,
		_w1261_,
		_w1262_
	);
	LUT2 #(
		.INIT('h4)
	) name1006 (
		_w1260_,
		_w1262_,
		_w1263_
	);
	LUT2 #(
		.INIT('h2)
	) name1007 (
		_w1260_,
		_w1262_,
		_w1264_
	);
	LUT2 #(
		.INIT('h1)
	) name1008 (
		_w1263_,
		_w1264_,
		_w1265_
	);
	LUT2 #(
		.INIT('h1)
	) name1009 (
		\a[127] ,
		\b[127] ,
		_w1266_
	);
	LUT2 #(
		.INIT('h8)
	) name1010 (
		\a[127] ,
		\b[127] ,
		_w1267_
	);
	LUT2 #(
		.INIT('h1)
	) name1011 (
		_w1266_,
		_w1267_,
		_w1268_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w1259_,
		_w1262_,
		_w1269_
	);
	LUT2 #(
		.INIT('h1)
	) name1013 (
		_w1258_,
		_w1269_,
		_w1270_
	);
	LUT2 #(
		.INIT('h2)
	) name1014 (
		_w1268_,
		_w1270_,
		_w1271_
	);
	LUT2 #(
		.INIT('h4)
	) name1015 (
		_w1268_,
		_w1270_,
		_w1272_
	);
	LUT2 #(
		.INIT('h1)
	) name1016 (
		_w1271_,
		_w1272_,
		_w1273_
	);
	LUT2 #(
		.INIT('h1)
	) name1017 (
		_w1267_,
		_w1270_,
		_w1274_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		_w1266_,
		_w1274_,
		_w1275_
	);
	assign \f[0]  = _w259_ ;
	assign \f[1]  = _w265_ ;
	assign \f[2]  = _w273_ ;
	assign \f[3]  = _w281_ ;
	assign \f[4]  = _w289_ ;
	assign \f[5]  = _w297_ ;
	assign \f[6]  = _w305_ ;
	assign \f[7]  = _w313_ ;
	assign \f[8]  = _w321_ ;
	assign \f[9]  = _w329_ ;
	assign \f[10]  = _w337_ ;
	assign \f[11]  = _w345_ ;
	assign \f[12]  = _w353_ ;
	assign \f[13]  = _w361_ ;
	assign \f[14]  = _w369_ ;
	assign \f[15]  = _w377_ ;
	assign \f[16]  = _w385_ ;
	assign \f[17]  = _w393_ ;
	assign \f[18]  = _w401_ ;
	assign \f[19]  = _w409_ ;
	assign \f[20]  = _w417_ ;
	assign \f[21]  = _w425_ ;
	assign \f[22]  = _w433_ ;
	assign \f[23]  = _w441_ ;
	assign \f[24]  = _w449_ ;
	assign \f[25]  = _w457_ ;
	assign \f[26]  = _w465_ ;
	assign \f[27]  = _w473_ ;
	assign \f[28]  = _w481_ ;
	assign \f[29]  = _w489_ ;
	assign \f[30]  = _w497_ ;
	assign \f[31]  = _w505_ ;
	assign \f[32]  = _w513_ ;
	assign \f[33]  = _w521_ ;
	assign \f[34]  = _w529_ ;
	assign \f[35]  = _w537_ ;
	assign \f[36]  = _w545_ ;
	assign \f[37]  = _w553_ ;
	assign \f[38]  = _w561_ ;
	assign \f[39]  = _w569_ ;
	assign \f[40]  = _w577_ ;
	assign \f[41]  = _w585_ ;
	assign \f[42]  = _w593_ ;
	assign \f[43]  = _w601_ ;
	assign \f[44]  = _w609_ ;
	assign \f[45]  = _w617_ ;
	assign \f[46]  = _w625_ ;
	assign \f[47]  = _w633_ ;
	assign \f[48]  = _w641_ ;
	assign \f[49]  = _w649_ ;
	assign \f[50]  = _w657_ ;
	assign \f[51]  = _w665_ ;
	assign \f[52]  = _w673_ ;
	assign \f[53]  = _w681_ ;
	assign \f[54]  = _w689_ ;
	assign \f[55]  = _w697_ ;
	assign \f[56]  = _w705_ ;
	assign \f[57]  = _w713_ ;
	assign \f[58]  = _w721_ ;
	assign \f[59]  = _w729_ ;
	assign \f[60]  = _w737_ ;
	assign \f[61]  = _w745_ ;
	assign \f[62]  = _w753_ ;
	assign \f[63]  = _w761_ ;
	assign \f[64]  = _w769_ ;
	assign \f[65]  = _w777_ ;
	assign \f[66]  = _w785_ ;
	assign \f[67]  = _w793_ ;
	assign \f[68]  = _w801_ ;
	assign \f[69]  = _w809_ ;
	assign \f[70]  = _w817_ ;
	assign \f[71]  = _w825_ ;
	assign \f[72]  = _w833_ ;
	assign \f[73]  = _w841_ ;
	assign \f[74]  = _w849_ ;
	assign \f[75]  = _w857_ ;
	assign \f[76]  = _w865_ ;
	assign \f[77]  = _w873_ ;
	assign \f[78]  = _w881_ ;
	assign \f[79]  = _w889_ ;
	assign \f[80]  = _w897_ ;
	assign \f[81]  = _w905_ ;
	assign \f[82]  = _w913_ ;
	assign \f[83]  = _w921_ ;
	assign \f[84]  = _w929_ ;
	assign \f[85]  = _w937_ ;
	assign \f[86]  = _w945_ ;
	assign \f[87]  = _w953_ ;
	assign \f[88]  = _w961_ ;
	assign \f[89]  = _w969_ ;
	assign \f[90]  = _w977_ ;
	assign \f[91]  = _w985_ ;
	assign \f[92]  = _w993_ ;
	assign \f[93]  = _w1001_ ;
	assign \f[94]  = _w1009_ ;
	assign \f[95]  = _w1017_ ;
	assign \f[96]  = _w1025_ ;
	assign \f[97]  = _w1033_ ;
	assign \f[98]  = _w1041_ ;
	assign \f[99]  = _w1049_ ;
	assign \f[100]  = _w1057_ ;
	assign \f[101]  = _w1065_ ;
	assign \f[102]  = _w1073_ ;
	assign \f[103]  = _w1081_ ;
	assign \f[104]  = _w1089_ ;
	assign \f[105]  = _w1097_ ;
	assign \f[106]  = _w1105_ ;
	assign \f[107]  = _w1113_ ;
	assign \f[108]  = _w1121_ ;
	assign \f[109]  = _w1129_ ;
	assign \f[110]  = _w1137_ ;
	assign \f[111]  = _w1145_ ;
	assign \f[112]  = _w1153_ ;
	assign \f[113]  = _w1161_ ;
	assign \f[114]  = _w1169_ ;
	assign \f[115]  = _w1177_ ;
	assign \f[116]  = _w1185_ ;
	assign \f[117]  = _w1193_ ;
	assign \f[118]  = _w1201_ ;
	assign \f[119]  = _w1209_ ;
	assign \f[120]  = _w1217_ ;
	assign \f[121]  = _w1225_ ;
	assign \f[122]  = _w1233_ ;
	assign \f[123]  = _w1241_ ;
	assign \f[124]  = _w1249_ ;
	assign \f[125]  = _w1257_ ;
	assign \f[126]  = _w1265_ ;
	assign \f[127]  = _w1273_ ;
	assign cOut = _w1275_ ;
endmodule;