module top (\DATA_0_0_pad , \DATA_0_10_pad , \DATA_0_11_pad , \DATA_0_12_pad , \DATA_0_13_pad , \DATA_0_14_pad , \DATA_0_15_pad , \DATA_0_16_pad , \DATA_0_17_pad , \DATA_0_18_pad , \DATA_0_19_pad , \DATA_0_1_pad , \DATA_0_20_pad , \DATA_0_21_pad , \DATA_0_22_pad , \DATA_0_23_pad , \DATA_0_24_pad , \DATA_0_25_pad , \DATA_0_26_pad , \DATA_0_27_pad , \DATA_0_28_pad , \DATA_0_29_pad , \DATA_0_2_pad , \DATA_0_30_pad , \DATA_0_31_pad , \DATA_0_3_pad , \DATA_0_4_pad , \DATA_0_5_pad , \DATA_0_6_pad , \DATA_0_7_pad , \DATA_0_8_pad , \DATA_0_9_pad , RESET_pad, \TM0_pad , \TM1_pad , \WX10829_reg/NET0131 , \WX10831_reg/NET0131 , \WX10833_reg/NET0131 , \WX10835_reg/NET0131 , \WX10837_reg/NET0131 , \WX10839_reg/NET0131 , \WX10841_reg/NET0131 , \WX10843_reg/NET0131 , \WX10845_reg/NET0131 , \WX10847_reg/NET0131 , \WX10849_reg/NET0131 , \WX10851_reg/NET0131 , \WX10853_reg/NET0131 , \WX10855_reg/NET0131 , \WX10857_reg/NET0131 , \WX10859_reg/NET0131 , \WX10861_reg/NET0131 , \WX10863_reg/NET0131 , \WX10865_reg/NET0131 , \WX10867_reg/NET0131 , \WX10869_reg/NET0131 , \WX10871_reg/NET0131 , \WX10873_reg/NET0131 , \WX10875_reg/NET0131 , \WX10877_reg/NET0131 , \WX10879_reg/NET0131 , \WX10881_reg/NET0131 , \WX10883_reg/NET0131 , \WX10885_reg/NET0131 , \WX10887_reg/NET0131 , \WX10889_reg/NET0131 , \WX10891_reg/NET0131 , \WX10989_reg/NET0131 , \WX10991_reg/NET0131 , \WX10993_reg/NET0131 , \WX10995_reg/NET0131 , \WX10997_reg/NET0131 , \WX10999_reg/NET0131 , \WX11001_reg/NET0131 , \WX11003_reg/NET0131 , \WX11005_reg/NET0131 , \WX11007_reg/NET0131 , \WX11009_reg/NET0131 , \WX11011_reg/NET0131 , \WX11013_reg/NET0131 , \WX11015_reg/NET0131 , \WX11017_reg/NET0131 , \WX11019_reg/NET0131 , \WX11021_reg/NET0131 , \WX11023_reg/NET0131 , \WX11025_reg/NET0131 , \WX11027_reg/NET0131 , \WX11029_reg/NET0131 , \WX11031_reg/NET0131 , \WX11033_reg/NET0131 , \WX11035_reg/NET0131 , \WX11037_reg/NET0131 , \WX11039_reg/NET0131 , \WX11041_reg/NET0131 , \WX11043_reg/NET0131 , \WX11045_reg/NET0131 , \WX11047_reg/NET0131 , \WX11049_reg/NET0131 , \WX11051_reg/NET0131 , \WX11053_reg/NET0131 , \WX11055_reg/NET0131 , \WX11057_reg/NET0131 , \WX11059_reg/NET0131 , \WX11061_reg/NET0131 , \WX11063_reg/NET0131 , \WX11065_reg/NET0131 , \WX11067_reg/NET0131 , \WX11069_reg/NET0131 , \WX11071_reg/NET0131 , \WX11073_reg/NET0131 , \WX11075_reg/NET0131 , \WX11077_reg/NET0131 , \WX11079_reg/NET0131 , \WX11081_reg/NET0131 , \WX11083_reg/NET0131 , \WX11085_reg/NET0131 , \WX11087_reg/NET0131 , \WX11089_reg/NET0131 , \WX11091_reg/NET0131 , \WX11093_reg/NET0131 , \WX11095_reg/NET0131 , \WX11097_reg/NET0131 , \WX11099_reg/NET0131 , \WX11101_reg/NET0131 , \WX11103_reg/NET0131 , \WX11105_reg/NET0131 , \WX11107_reg/NET0131 , \WX11109_reg/NET0131 , \WX11111_reg/NET0131 , \WX11113_reg/NET0131 , \WX11115_reg/NET0131 , \WX11117_reg/NET0131 , \WX11119_reg/NET0131 , \WX11121_reg/NET0131 , \WX11123_reg/NET0131 , \WX11125_reg/NET0131 , \WX11127_reg/NET0131 , \WX11129_reg/NET0131 , \WX11131_reg/NET0131 , \WX11133_reg/NET0131 , \WX11135_reg/NET0131 , \WX11137_reg/NET0131 , \WX11139_reg/NET0131 , \WX11141_reg/NET0131 , \WX11143_reg/NET0131 , \WX11145_reg/NET0131 , \WX11147_reg/NET0131 , \WX11149_reg/NET0131 , \WX11151_reg/NET0131 , \WX11153_reg/NET0131 , \WX11155_reg/NET0131 , \WX11157_reg/NET0131 , \WX11159_reg/NET0131 , \WX11161_reg/NET0131 , \WX11163_reg/NET0131 , \WX11165_reg/NET0131 , \WX11167_reg/NET0131 , \WX11169_reg/NET0131 , \WX11171_reg/NET0131 , \WX11173_reg/NET0131 , \WX11175_reg/NET0131 , \WX11177_reg/NET0131 , \WX11179_reg/NET0131 , \WX11181_reg/NET0131 , \WX11183_reg/NET0131 , \WX11185_reg/NET0131 , \WX11187_reg/NET0131 , \WX11189_reg/NET0131 , \WX11191_reg/NET0131 , \WX11193_reg/NET0131 , \WX11195_reg/NET0131 , \WX11197_reg/NET0131 , \WX11199_reg/NET0131 , \WX11201_reg/NET0131 , \WX11203_reg/NET0131 , \WX11205_reg/NET0131 , \WX11207_reg/NET0131 , \WX11209_reg/NET0131 , \WX11211_reg/NET0131 , \WX11213_reg/NET0131 , \WX11215_reg/NET0131 , \WX11217_reg/NET0131 , \WX11219_reg/NET0131 , \WX11221_reg/NET0131 , \WX11223_reg/NET0131 , \WX11225_reg/NET0131 , \WX11227_reg/NET0131 , \WX11229_reg/NET0131 , \WX11231_reg/NET0131 , \WX11233_reg/NET0131 , \WX11235_reg/NET0131 , \WX11237_reg/NET0131 , \WX11239_reg/NET0131 , \WX11241_reg/NET0131 , \WX11243_reg/NET0131 , \WX1938_reg/NET0131 , \WX1940_reg/NET0131 , \WX1942_reg/NET0131 , \WX1944_reg/NET0131 , \WX1946_reg/NET0131 , \WX1948_reg/NET0131 , \WX1950_reg/NET0131 , \WX1952_reg/NET0131 , \WX1954_reg/NET0131 , \WX1956_reg/NET0131 , \WX1958_reg/NET0131 , \WX1960_reg/NET0131 , \WX1962_reg/NET0131 , \WX1964_reg/NET0131 , \WX1966_reg/NET0131 , \WX1968_reg/NET0131 , \WX1970_reg/NET0131 , \WX1972_reg/NET0131 , \WX1974_reg/NET0131 , \WX1976_reg/NET0131 , \WX1978_reg/NET0131 , \WX1980_reg/NET0131 , \WX1982_reg/NET0131 , \WX1984_reg/NET0131 , \WX1986_reg/NET0131 , \WX1988_reg/NET0131 , \WX1990_reg/NET0131 , \WX1992_reg/NET0131 , \WX1994_reg/NET0131 , \WX1996_reg/NET0131 , \WX1998_reg/NET0131 , \WX2000_reg/NET0131 , \WX2002_reg/NET0131 , \WX2004_reg/NET0131 , \WX2006_reg/NET0131 , \WX2008_reg/NET0131 , \WX2010_reg/NET0131 , \WX2012_reg/NET0131 , \WX2014_reg/NET0131 , \WX2016_reg/NET0131 , \WX2018_reg/NET0131 , \WX2020_reg/NET0131 , \WX2022_reg/NET0131 , \WX2024_reg/NET0131 , \WX2026_reg/NET0131 , \WX2028_reg/NET0131 , \WX2030_reg/NET0131 , \WX2032_reg/NET0131 , \WX2034_reg/NET0131 , \WX2036_reg/NET0131 , \WX2038_reg/NET0131 , \WX2040_reg/NET0131 , \WX2042_reg/NET0131 , \WX2044_reg/NET0131 , \WX2046_reg/NET0131 , \WX2048_reg/NET0131 , \WX2050_reg/NET0131 , \WX2052_reg/NET0131 , \WX2054_reg/NET0131 , \WX2056_reg/NET0131 , \WX2058_reg/NET0131 , \WX2060_reg/NET0131 , \WX2062_reg/NET0131 , \WX2064_reg/NET0131 , \WX2066_reg/NET0131 , \WX2068_reg/NET0131 , \WX2070_reg/NET0131 , \WX2072_reg/NET0131 , \WX2074_reg/NET0131 , \WX2076_reg/NET0131 , \WX2078_reg/NET0131 , \WX2080_reg/NET0131 , \WX2082_reg/NET0131 , \WX2084_reg/NET0131 , \WX2086_reg/NET0131 , \WX2088_reg/NET0131 , \WX2090_reg/NET0131 , \WX2092_reg/NET0131 , \WX2094_reg/NET0131 , \WX2096_reg/NET0131 , \WX2098_reg/NET0131 , \WX2100_reg/NET0131 , \WX2102_reg/NET0131 , \WX2104_reg/NET0131 , \WX2106_reg/NET0131 , \WX2108_reg/NET0131 , \WX2110_reg/NET0131 , \WX2112_reg/NET0131 , \WX2114_reg/NET0131 , \WX2116_reg/NET0131 , \WX2118_reg/NET0131 , \WX2120_reg/NET0131 , \WX2122_reg/NET0131 , \WX2124_reg/NET0131 , \WX2126_reg/NET0131 , \WX2128_reg/NET0131 , \WX2130_reg/NET0131 , \WX2132_reg/NET0131 , \WX2134_reg/NET0131 , \WX2136_reg/NET0131 , \WX2138_reg/NET0131 , \WX2140_reg/NET0131 , \WX2142_reg/NET0131 , \WX2144_reg/NET0131 , \WX2146_reg/NET0131 , \WX2148_reg/NET0131 , \WX2150_reg/NET0131 , \WX2152_reg/NET0131 , \WX2154_reg/NET0131 , \WX2156_reg/NET0131 , \WX2158_reg/NET0131 , \WX2160_reg/NET0131 , \WX2162_reg/NET0131 , \WX2164_reg/NET0131 , \WX2166_reg/NET0131 , \WX2168_reg/NET0131 , \WX2170_reg/NET0131 , \WX2172_reg/NET0131 , \WX2174_reg/NET0131 , \WX2176_reg/NET0131 , \WX2178_reg/NET0131 , \WX2180_reg/NET0131 , \WX2182_reg/NET0131 , \WX2184_reg/NET0131 , \WX2186_reg/NET0131 , \WX2188_reg/NET0131 , \WX2190_reg/NET0131 , \WX2192_reg/NET0131 , \WX3231_reg/NET0131 , \WX3233_reg/NET0131 , \WX3235_reg/NET0131 , \WX3237_reg/NET0131 , \WX3239_reg/NET0131 , \WX3241_reg/NET0131 , \WX3243_reg/NET0131 , \WX3245_reg/NET0131 , \WX3247_reg/NET0131 , \WX3249_reg/NET0131 , \WX3251_reg/NET0131 , \WX3253_reg/NET0131 , \WX3255_reg/NET0131 , \WX3257_reg/NET0131 , \WX3259_reg/NET0131 , \WX3261_reg/NET0131 , \WX3263_reg/NET0131 , \WX3265_reg/NET0131 , \WX3267_reg/NET0131 , \WX3269_reg/NET0131 , \WX3271_reg/NET0131 , \WX3273_reg/NET0131 , \WX3275_reg/NET0131 , \WX3277_reg/NET0131 , \WX3279_reg/NET0131 , \WX3281_reg/NET0131 , \WX3283_reg/NET0131 , \WX3285_reg/NET0131 , \WX3287_reg/NET0131 , \WX3289_reg/NET0131 , \WX3291_reg/NET0131 , \WX3293_reg/NET0131 , \WX3295_reg/NET0131 , \WX3297_reg/NET0131 , \WX3299_reg/NET0131 , \WX3301_reg/NET0131 , \WX3303_reg/NET0131 , \WX3305_reg/NET0131 , \WX3307_reg/NET0131 , \WX3309_reg/NET0131 , \WX3311_reg/NET0131 , \WX3313_reg/NET0131 , \WX3315_reg/NET0131 , \WX3317_reg/NET0131 , \WX3319_reg/NET0131 , \WX3321_reg/NET0131 , \WX3323_reg/NET0131 , \WX3325_reg/NET0131 , \WX3327_reg/NET0131 , \WX3329_reg/NET0131 , \WX3331_reg/NET0131 , \WX3333_reg/NET0131 , \WX3335_reg/NET0131 , \WX3337_reg/NET0131 , \WX3339_reg/NET0131 , \WX3341_reg/NET0131 , \WX3343_reg/NET0131 , \WX3345_reg/NET0131 , \WX3347_reg/NET0131 , \WX3349_reg/NET0131 , \WX3351_reg/NET0131 , \WX3353_reg/NET0131 , \WX3355_reg/NET0131 , \WX3357_reg/NET0131 , \WX3359_reg/NET0131 , \WX3361_reg/NET0131 , \WX3363_reg/NET0131 , \WX3365_reg/NET0131 , \WX3367_reg/NET0131 , \WX3369_reg/NET0131 , \WX3371_reg/NET0131 , \WX3373_reg/NET0131 , \WX3375_reg/NET0131 , \WX3377_reg/NET0131 , \WX3379_reg/NET0131 , \WX3381_reg/NET0131 , \WX3383_reg/NET0131 , \WX3385_reg/NET0131 , \WX3387_reg/NET0131 , \WX3389_reg/NET0131 , \WX3391_reg/NET0131 , \WX3393_reg/NET0131 , \WX3395_reg/NET0131 , \WX3397_reg/NET0131 , \WX3399_reg/NET0131 , \WX3401_reg/NET0131 , \WX3403_reg/NET0131 , \WX3405_reg/NET0131 , \WX3407_reg/NET0131 , \WX3409_reg/NET0131 , \WX3411_reg/NET0131 , \WX3413_reg/NET0131 , \WX3415_reg/NET0131 , \WX3417_reg/NET0131 , \WX3419_reg/NET0131 , \WX3421_reg/NET0131 , \WX3423_reg/NET0131 , \WX3425_reg/NET0131 , \WX3427_reg/NET0131 , \WX3429_reg/NET0131 , \WX3431_reg/NET0131 , \WX3433_reg/NET0131 , \WX3435_reg/NET0131 , \WX3437_reg/NET0131 , \WX3439_reg/NET0131 , \WX3441_reg/NET0131 , \WX3443_reg/NET0131 , \WX3445_reg/NET0131 , \WX3447_reg/NET0131 , \WX3449_reg/NET0131 , \WX3451_reg/NET0131 , \WX3453_reg/NET0131 , \WX3455_reg/NET0131 , \WX3457_reg/NET0131 , \WX3459_reg/NET0131 , \WX3461_reg/NET0131 , \WX3463_reg/NET0131 , \WX3465_reg/NET0131 , \WX3467_reg/NET0131 , \WX3469_reg/NET0131 , \WX3471_reg/NET0131 , \WX3473_reg/NET0131 , \WX3475_reg/NET0131 , \WX3477_reg/NET0131 , \WX3479_reg/NET0131 , \WX3481_reg/NET0131 , \WX3483_reg/NET0131 , \WX3485_reg/NET0131 , \WX4524_reg/NET0131 , \WX4526_reg/NET0131 , \WX4528_reg/NET0131 , \WX4530_reg/NET0131 , \WX4532_reg/NET0131 , \WX4534_reg/NET0131 , \WX4536_reg/NET0131 , \WX4538_reg/NET0131 , \WX4540_reg/NET0131 , \WX4542_reg/NET0131 , \WX4544_reg/NET0131 , \WX4546_reg/NET0131 , \WX4548_reg/NET0131 , \WX4550_reg/NET0131 , \WX4552_reg/NET0131 , \WX4554_reg/NET0131 , \WX4556_reg/NET0131 , \WX4558_reg/NET0131 , \WX4560_reg/NET0131 , \WX4562_reg/NET0131 , \WX4564_reg/NET0131 , \WX4566_reg/NET0131 , \WX4568_reg/NET0131 , \WX4570_reg/NET0131 , \WX4572_reg/NET0131 , \WX4574_reg/NET0131 , \WX4576_reg/NET0131 , \WX4578_reg/NET0131 , \WX4580_reg/NET0131 , \WX4582_reg/NET0131 , \WX4584_reg/NET0131 , \WX4586_reg/NET0131 , \WX4588_reg/NET0131 , \WX4590_reg/NET0131 , \WX4592_reg/NET0131 , \WX4594_reg/NET0131 , \WX4596_reg/NET0131 , \WX4598_reg/NET0131 , \WX4600_reg/NET0131 , \WX4602_reg/NET0131 , \WX4604_reg/NET0131 , \WX4606_reg/NET0131 , \WX4608_reg/NET0131 , \WX4610_reg/NET0131 , \WX4612_reg/NET0131 , \WX4614_reg/NET0131 , \WX4616_reg/NET0131 , \WX4618_reg/NET0131 , \WX4620_reg/NET0131 , \WX4622_reg/NET0131 , \WX4624_reg/NET0131 , \WX4626_reg/NET0131 , \WX4628_reg/NET0131 , \WX4630_reg/NET0131 , \WX4632_reg/NET0131 , \WX4634_reg/NET0131 , \WX4636_reg/NET0131 , \WX4638_reg/NET0131 , \WX4640_reg/NET0131 , \WX4642_reg/NET0131 , \WX4644_reg/NET0131 , \WX4646_reg/NET0131 , \WX4648_reg/NET0131 , \WX4650_reg/NET0131 , \WX4652_reg/NET0131 , \WX4654_reg/NET0131 , \WX4656_reg/NET0131 , \WX4658_reg/NET0131 , \WX4660_reg/NET0131 , \WX4662_reg/NET0131 , \WX4664_reg/NET0131 , \WX4666_reg/NET0131 , \WX4668_reg/NET0131 , \WX4670_reg/NET0131 , \WX4672_reg/NET0131 , \WX4674_reg/NET0131 , \WX4676_reg/NET0131 , \WX4678_reg/NET0131 , \WX4680_reg/NET0131 , \WX4682_reg/NET0131 , \WX4684_reg/NET0131 , \WX4686_reg/NET0131 , \WX4688_reg/NET0131 , \WX4690_reg/NET0131 , \WX4692_reg/NET0131 , \WX4694_reg/NET0131 , \WX4696_reg/NET0131 , \WX4698_reg/NET0131 , \WX4700_reg/NET0131 , \WX4702_reg/NET0131 , \WX4704_reg/NET0131 , \WX4706_reg/NET0131 , \WX4708_reg/NET0131 , \WX4710_reg/NET0131 , \WX4712_reg/NET0131 , \WX4714_reg/NET0131 , \WX4716_reg/NET0131 , \WX4718_reg/NET0131 , \WX4720_reg/NET0131 , \WX4722_reg/NET0131 , \WX4724_reg/NET0131 , \WX4726_reg/NET0131 , \WX4728_reg/NET0131 , \WX4730_reg/NET0131 , \WX4732_reg/NET0131 , \WX4734_reg/NET0131 , \WX4736_reg/NET0131 , \WX4738_reg/NET0131 , \WX4740_reg/NET0131 , \WX4742_reg/NET0131 , \WX4744_reg/NET0131 , \WX4746_reg/NET0131 , \WX4748_reg/NET0131 , \WX4750_reg/NET0131 , \WX4752_reg/NET0131 , \WX4754_reg/NET0131 , \WX4756_reg/NET0131 , \WX4758_reg/NET0131 , \WX4760_reg/NET0131 , \WX4762_reg/NET0131 , \WX4764_reg/NET0131 , \WX4766_reg/NET0131 , \WX4768_reg/NET0131 , \WX4770_reg/NET0131 , \WX4772_reg/NET0131 , \WX4774_reg/NET0131 , \WX4776_reg/NET0131 , \WX4778_reg/NET0131 , \WX5817_reg/NET0131 , \WX5819_reg/NET0131 , \WX5821_reg/NET0131 , \WX5823_reg/NET0131 , \WX5825_reg/NET0131 , \WX5827_reg/NET0131 , \WX5829_reg/NET0131 , \WX5831_reg/NET0131 , \WX5833_reg/NET0131 , \WX5835_reg/NET0131 , \WX5837_reg/NET0131 , \WX5839_reg/NET0131 , \WX5841_reg/NET0131 , \WX5843_reg/NET0131 , \WX5845_reg/NET0131 , \WX5847_reg/NET0131 , \WX5849_reg/NET0131 , \WX5851_reg/NET0131 , \WX5853_reg/NET0131 , \WX5855_reg/NET0131 , \WX5857_reg/NET0131 , \WX5859_reg/NET0131 , \WX5861_reg/NET0131 , \WX5863_reg/NET0131 , \WX5865_reg/NET0131 , \WX5867_reg/NET0131 , \WX5869_reg/NET0131 , \WX5871_reg/NET0131 , \WX5873_reg/NET0131 , \WX5875_reg/NET0131 , \WX5877_reg/NET0131 , \WX5879_reg/NET0131 , \WX5881_reg/NET0131 , \WX5883_reg/NET0131 , \WX5885_reg/NET0131 , \WX5887_reg/NET0131 , \WX5889_reg/NET0131 , \WX5891_reg/NET0131 , \WX5893_reg/NET0131 , \WX5895_reg/NET0131 , \WX5897_reg/NET0131 , \WX5899_reg/NET0131 , \WX5901_reg/NET0131 , \WX5903_reg/NET0131 , \WX5905_reg/NET0131 , \WX5907_reg/NET0131 , \WX5909_reg/NET0131 , \WX5911_reg/NET0131 , \WX5913_reg/NET0131 , \WX5915_reg/NET0131 , \WX5917_reg/NET0131 , \WX5919_reg/NET0131 , \WX5921_reg/NET0131 , \WX5923_reg/NET0131 , \WX5925_reg/NET0131 , \WX5927_reg/NET0131 , \WX5929_reg/NET0131 , \WX5931_reg/NET0131 , \WX5933_reg/NET0131 , \WX5935_reg/NET0131 , \WX5937_reg/NET0131 , \WX5939_reg/NET0131 , \WX5941_reg/NET0131 , \WX5943_reg/NET0131 , \WX5945_reg/NET0131 , \WX5947_reg/NET0131 , \WX5949_reg/NET0131 , \WX5951_reg/NET0131 , \WX5953_reg/NET0131 , \WX5955_reg/NET0131 , \WX5957_reg/NET0131 , \WX5959_reg/NET0131 , \WX5961_reg/NET0131 , \WX5963_reg/NET0131 , \WX5965_reg/NET0131 , \WX5967_reg/NET0131 , \WX5969_reg/NET0131 , \WX5971_reg/NET0131 , \WX5973_reg/NET0131 , \WX5975_reg/NET0131 , \WX5977_reg/NET0131 , \WX5979_reg/NET0131 , \WX5981_reg/NET0131 , \WX5983_reg/NET0131 , \WX5985_reg/NET0131 , \WX5987_reg/NET0131 , \WX5989_reg/NET0131 , \WX5991_reg/NET0131 , \WX5993_reg/NET0131 , \WX5995_reg/NET0131 , \WX5997_reg/NET0131 , \WX5999_reg/NET0131 , \WX6001_reg/NET0131 , \WX6003_reg/NET0131 , \WX6005_reg/NET0131 , \WX6007_reg/NET0131 , \WX6009_reg/NET0131 , \WX6011_reg/NET0131 , \WX6013_reg/NET0131 , \WX6015_reg/NET0131 , \WX6017_reg/NET0131 , \WX6019_reg/NET0131 , \WX6021_reg/NET0131 , \WX6023_reg/NET0131 , \WX6025_reg/NET0131 , \WX6027_reg/NET0131 , \WX6029_reg/NET0131 , \WX6031_reg/NET0131 , \WX6033_reg/NET0131 , \WX6035_reg/NET0131 , \WX6037_reg/NET0131 , \WX6039_reg/NET0131 , \WX6041_reg/NET0131 , \WX6043_reg/NET0131 , \WX6045_reg/NET0131 , \WX6047_reg/NET0131 , \WX6049_reg/NET0131 , \WX6051_reg/NET0131 , \WX6053_reg/NET0131 , \WX6055_reg/NET0131 , \WX6057_reg/NET0131 , \WX6059_reg/NET0131 , \WX6061_reg/NET0131 , \WX6063_reg/NET0131 , \WX6065_reg/NET0131 , \WX6067_reg/NET0131 , \WX6069_reg/NET0131 , \WX6071_reg/NET0131 , \WX645_reg/NET0131 , \WX647_reg/NET0131 , \WX649_reg/NET0131 , \WX651_reg/NET0131 , \WX653_reg/NET0131 , \WX655_reg/NET0131 , \WX657_reg/NET0131 , \WX659_reg/NET0131 , \WX661_reg/NET0131 , \WX663_reg/NET0131 , \WX665_reg/NET0131 , \WX667_reg/NET0131 , \WX669_reg/NET0131 , \WX671_reg/NET0131 , \WX673_reg/NET0131 , \WX675_reg/NET0131 , \WX677_reg/NET0131 , \WX679_reg/NET0131 , \WX681_reg/NET0131 , \WX683_reg/NET0131 , \WX685_reg/NET0131 , \WX687_reg/NET0131 , \WX689_reg/NET0131 , \WX691_reg/NET0131 , \WX693_reg/NET0131 , \WX695_reg/NET0131 , \WX697_reg/NET0131 , \WX699_reg/NET0131 , \WX701_reg/NET0131 , \WX703_reg/NET0131 , \WX705_reg/NET0131 , \WX707_reg/NET0131 , \WX709_reg/NET0131 , \WX7110_reg/NET0131 , \WX7112_reg/NET0131 , \WX7114_reg/NET0131 , \WX7116_reg/NET0131 , \WX7118_reg/NET0131 , \WX711_reg/NET0131 , \WX7120_reg/NET0131 , \WX7122_reg/NET0131 , \WX7124_reg/NET0131 , \WX7126_reg/NET0131 , \WX7128_reg/NET0131 , \WX7130_reg/NET0131 , \WX7132_reg/NET0131 , \WX7134_reg/NET0131 , \WX7136_reg/NET0131 , \WX7138_reg/NET0131 , \WX713_reg/NET0131 , \WX7140_reg/NET0131 , \WX7142_reg/NET0131 , \WX7144_reg/NET0131 , \WX7146_reg/NET0131 , \WX7148_reg/NET0131 , \WX7150_reg/NET0131 , \WX7152_reg/NET0131 , \WX7154_reg/NET0131 , \WX7156_reg/NET0131 , \WX7158_reg/NET0131 , \WX715_reg/NET0131 , \WX7160_reg/NET0131 , \WX7162_reg/NET0131 , \WX7164_reg/NET0131 , \WX7166_reg/NET0131 , \WX7168_reg/NET0131 , \WX7170_reg/NET0131 , \WX7172_reg/NET0131 , \WX7174_reg/NET0131 , \WX7176_reg/NET0131 , \WX7178_reg/NET0131 , \WX717_reg/NET0131 , \WX7180_reg/NET0131 , \WX7182_reg/NET0131 , \WX7184_reg/NET0131 , \WX7186_reg/NET0131 , \WX7188_reg/NET0131 , \WX7190_reg/NET0131 , \WX7192_reg/NET0131 , \WX7194_reg/NET0131 , \WX7196_reg/NET0131 , \WX7198_reg/NET0131 , \WX719_reg/NET0131 , \WX7200_reg/NET0131 , \WX7202_reg/NET0131 , \WX7204_reg/NET0131 , \WX7206_reg/NET0131 , \WX7208_reg/NET0131 , \WX7210_reg/NET0131 , \WX7212_reg/NET0131 , \WX7214_reg/NET0131 , \WX7216_reg/NET0131 , \WX7218_reg/NET0131 , \WX721_reg/NET0131 , \WX7220_reg/NET0131 , \WX7222_reg/NET0131 , \WX7224_reg/NET0131 , \WX7226_reg/NET0131 , \WX7228_reg/NET0131 , \WX7230_reg/NET0131 , \WX7232_reg/NET0131 , \WX7234_reg/NET0131 , \WX7236_reg/NET0131 , \WX7238_reg/NET0131 , \WX723_reg/NET0131 , \WX7240_reg/NET0131 , \WX7242_reg/NET0131 , \WX7244_reg/NET0131 , \WX7246_reg/NET0131 , \WX7248_reg/NET0131 , \WX7250_reg/NET0131 , \WX7252_reg/NET0131 , \WX7254_reg/NET0131 , \WX7256_reg/NET0131 , \WX7258_reg/NET0131 , \WX725_reg/NET0131 , \WX7260_reg/NET0131 , \WX7262_reg/NET0131 , \WX7264_reg/NET0131 , \WX7266_reg/NET0131 , \WX7268_reg/NET0131 , \WX7270_reg/NET0131 , \WX7272_reg/NET0131 , \WX7274_reg/NET0131 , \WX7276_reg/NET0131 , \WX7278_reg/NET0131 , \WX727_reg/NET0131 , \WX7280_reg/NET0131 , \WX7282_reg/NET0131 , \WX7284_reg/NET0131 , \WX7286_reg/NET0131 , \WX7288_reg/NET0131 , \WX7290_reg/NET0131 , \WX7292_reg/NET0131 , \WX7294_reg/NET0131 , \WX7296_reg/NET0131 , \WX7298_reg/NET0131 , \WX729_reg/NET0131 , \WX7300_reg/NET0131 , \WX7302_reg/NET0131 , \WX7304_reg/NET0131 , \WX7306_reg/NET0131 , \WX7308_reg/NET0131 , \WX7310_reg/NET0131 , \WX7312_reg/NET0131 , \WX7314_reg/NET0131 , \WX7316_reg/NET0131 , \WX7318_reg/NET0131 , \WX731_reg/NET0131 , \WX7320_reg/NET0131 , \WX7322_reg/NET0131 , \WX7324_reg/NET0131 , \WX7326_reg/NET0131 , \WX7328_reg/NET0131 , \WX7330_reg/NET0131 , \WX7332_reg/NET0131 , \WX7334_reg/NET0131 , \WX7336_reg/NET0131 , \WX7338_reg/NET0131 , \WX733_reg/NET0131 , \WX7340_reg/NET0131 , \WX7342_reg/NET0131 , \WX7344_reg/NET0131 , \WX7346_reg/NET0131 , \WX7348_reg/NET0131 , \WX7350_reg/NET0131 , \WX7352_reg/NET0131 , \WX7354_reg/NET0131 , \WX7356_reg/NET0131 , \WX7358_reg/NET0131 , \WX735_reg/NET0131 , \WX7360_reg/NET0131 , \WX7362_reg/NET0131 , \WX7364_reg/NET0131 , \WX737_reg/NET0131 , \WX739_reg/NET0131 , \WX741_reg/NET0131 , \WX743_reg/NET0131 , \WX745_reg/NET0131 , \WX747_reg/NET0131 , \WX749_reg/NET0131 , \WX751_reg/NET0131 , \WX753_reg/NET0131 , \WX755_reg/NET0131 , \WX757_reg/NET0131 , \WX759_reg/NET0131 , \WX761_reg/NET0131 , \WX763_reg/NET0131 , \WX765_reg/NET0131 , \WX767_reg/NET0131 , \WX769_reg/NET0131 , \WX771_reg/NET0131 , \WX773_reg/NET0131 , \WX775_reg/NET0131 , \WX777_reg/NET0131 , \WX779_reg/NET0131 , \WX781_reg/NET0131 , \WX783_reg/NET0131 , \WX785_reg/NET0131 , \WX787_reg/NET0131 , \WX789_reg/NET0131 , \WX791_reg/NET0131 , \WX793_reg/NET0131 , \WX795_reg/NET0131 , \WX797_reg/NET0131 , \WX799_reg/NET0131 , \WX801_reg/NET0131 , \WX803_reg/NET0131 , \WX805_reg/NET0131 , \WX807_reg/NET0131 , \WX809_reg/NET0131 , \WX811_reg/NET0131 , \WX813_reg/NET0131 , \WX815_reg/NET0131 , \WX817_reg/NET0131 , \WX819_reg/NET0131 , \WX821_reg/NET0131 , \WX823_reg/NET0131 , \WX825_reg/NET0131 , \WX827_reg/NET0131 , \WX829_reg/NET0131 , \WX831_reg/NET0131 , \WX833_reg/NET0131 , \WX835_reg/NET0131 , \WX837_reg/NET0131 , \WX839_reg/NET0131 , \WX8403_reg/NET0131 , \WX8405_reg/NET0131 , \WX8407_reg/NET0131 , \WX8409_reg/NET0131 , \WX8411_reg/NET0131 , \WX8413_reg/NET0131 , \WX8415_reg/NET0131 , \WX8417_reg/NET0131 , \WX8419_reg/NET0131 , \WX841_reg/NET0131 , \WX8421_reg/NET0131 , \WX8423_reg/NET0131 , \WX8425_reg/NET0131 , \WX8427_reg/NET0131 , \WX8429_reg/NET0131 , \WX8431_reg/NET0131 , \WX8433_reg/NET0131 , \WX8435_reg/NET0131 , \WX8437_reg/NET0131 , \WX8439_reg/NET0131 , \WX843_reg/NET0131 , \WX8441_reg/NET0131 , \WX8443_reg/NET0131 , \WX8445_reg/NET0131 , \WX8447_reg/NET0131 , \WX8449_reg/NET0131 , \WX8451_reg/NET0131 , \WX8453_reg/NET0131 , \WX8455_reg/NET0131 , \WX8457_reg/NET0131 , \WX8459_reg/NET0131 , \WX845_reg/NET0131 , \WX8461_reg/NET0131 , \WX8463_reg/NET0131 , \WX8465_reg/NET0131 , \WX8467_reg/NET0131 , \WX8469_reg/NET0131 , \WX8471_reg/NET0131 , \WX8473_reg/NET0131 , \WX8475_reg/NET0131 , \WX8477_reg/NET0131 , \WX8479_reg/NET0131 , \WX847_reg/NET0131 , \WX8481_reg/NET0131 , \WX8483_reg/NET0131 , \WX8485_reg/NET0131 , \WX8487_reg/NET0131 , \WX8489_reg/NET0131 , \WX8491_reg/NET0131 , \WX8493_reg/NET0131 , \WX8495_reg/NET0131 , \WX8497_reg/NET0131 , \WX8499_reg/NET0131 , \WX849_reg/NET0131 , \WX8501_reg/NET0131 , \WX8503_reg/NET0131 , \WX8505_reg/NET0131 , \WX8507_reg/NET0131 , \WX8509_reg/NET0131 , \WX8511_reg/NET0131 , \WX8513_reg/NET0131 , \WX8515_reg/NET0131 , \WX8517_reg/NET0131 , \WX8519_reg/NET0131 , \WX851_reg/NET0131 , \WX8521_reg/NET0131 , \WX8523_reg/NET0131 , \WX8525_reg/NET0131 , \WX8527_reg/NET0131 , \WX8529_reg/NET0131 , \WX8531_reg/NET0131 , \WX8533_reg/NET0131 , \WX8535_reg/NET0131 , \WX8537_reg/NET0131 , \WX8539_reg/NET0131 , \WX853_reg/NET0131 , \WX8541_reg/NET0131 , \WX8543_reg/NET0131 , \WX8545_reg/NET0131 , \WX8547_reg/NET0131 , \WX8549_reg/NET0131 , \WX8551_reg/NET0131 , \WX8553_reg/NET0131 , \WX8555_reg/NET0131 , \WX8557_reg/NET0131 , \WX8559_reg/NET0131 , \WX855_reg/NET0131 , \WX8561_reg/NET0131 , \WX8563_reg/NET0131 , \WX8565_reg/NET0131 , \WX8567_reg/NET0131 , \WX8569_reg/NET0131 , \WX8571_reg/NET0131 , \WX8573_reg/NET0131 , \WX8575_reg/NET0131 , \WX8577_reg/NET0131 , \WX8579_reg/NET0131 , \WX857_reg/NET0131 , \WX8581_reg/NET0131 , \WX8583_reg/NET0131 , \WX8585_reg/NET0131 , \WX8587_reg/NET0131 , \WX8589_reg/NET0131 , \WX8591_reg/NET0131 , \WX8593_reg/NET0131 , \WX8595_reg/NET0131 , \WX8597_reg/NET0131 , \WX8599_reg/NET0131 , \WX859_reg/NET0131 , \WX8601_reg/NET0131 , \WX8603_reg/NET0131 , \WX8605_reg/NET0131 , \WX8607_reg/NET0131 , \WX8609_reg/NET0131 , \WX8611_reg/NET0131 , \WX8613_reg/NET0131 , \WX8615_reg/NET0131 , \WX8617_reg/NET0131 , \WX8619_reg/NET0131 , \WX861_reg/NET0131 , \WX8621_reg/NET0131 , \WX8623_reg/NET0131 , \WX8625_reg/NET0131 , \WX8627_reg/NET0131 , \WX8629_reg/NET0131 , \WX8631_reg/NET0131 , \WX8633_reg/NET0131 , \WX8635_reg/NET0131 , \WX8637_reg/NET0131 , \WX8639_reg/NET0131 , \WX863_reg/NET0131 , \WX8641_reg/NET0131 , \WX8643_reg/NET0131 , \WX8645_reg/NET0131 , \WX8647_reg/NET0131 , \WX8649_reg/NET0131 , \WX8651_reg/NET0131 , \WX8653_reg/NET0131 , \WX8655_reg/NET0131 , \WX8657_reg/NET0131 , \WX865_reg/NET0131 , \WX867_reg/NET0131 , \WX869_reg/NET0131 , \WX871_reg/NET0131 , \WX873_reg/NET0131 , \WX875_reg/NET0131 , \WX877_reg/NET0131 , \WX879_reg/NET0131 , \WX881_reg/NET0131 , \WX883_reg/NET0131 , \WX885_reg/NET0131 , \WX887_reg/NET0131 , \WX889_reg/NET0131 , \WX891_reg/NET0131 , \WX893_reg/NET0131 , \WX895_reg/NET0131 , \WX897_reg/NET0131 , \WX899_reg/NET0131 , \WX9696_reg/NET0131 , \WX9698_reg/NET0131 , \WX9700_reg/NET0131 , \WX9702_reg/NET0131 , \WX9704_reg/NET0131 , \WX9706_reg/NET0131 , \WX9708_reg/NET0131 , \WX9710_reg/NET0131 , \WX9712_reg/NET0131 , \WX9714_reg/NET0131 , \WX9716_reg/NET0131 , \WX9718_reg/NET0131 , \WX9720_reg/NET0131 , \WX9722_reg/NET0131 , \WX9724_reg/NET0131 , \WX9726_reg/NET0131 , \WX9728_reg/NET0131 , \WX9730_reg/NET0131 , \WX9732_reg/NET0131 , \WX9734_reg/NET0131 , \WX9736_reg/NET0131 , \WX9738_reg/NET0131 , \WX9740_reg/NET0131 , \WX9742_reg/NET0131 , \WX9744_reg/NET0131 , \WX9746_reg/NET0131 , \WX9748_reg/NET0131 , \WX9750_reg/NET0131 , \WX9752_reg/NET0131 , \WX9754_reg/NET0131 , \WX9756_reg/NET0131 , \WX9758_reg/NET0131 , \WX9760_reg/NET0131 , \WX9762_reg/NET0131 , \WX9764_reg/NET0131 , \WX9766_reg/NET0131 , \WX9768_reg/NET0131 , \WX9770_reg/NET0131 , \WX9772_reg/NET0131 , \WX9774_reg/NET0131 , \WX9776_reg/NET0131 , \WX9778_reg/NET0131 , \WX9780_reg/NET0131 , \WX9782_reg/NET0131 , \WX9784_reg/NET0131 , \WX9786_reg/NET0131 , \WX9788_reg/NET0131 , \WX9790_reg/NET0131 , \WX9792_reg/NET0131 , \WX9794_reg/NET0131 , \WX9796_reg/NET0131 , \WX9798_reg/NET0131 , \WX9800_reg/NET0131 , \WX9802_reg/NET0131 , \WX9804_reg/NET0131 , \WX9806_reg/NET0131 , \WX9808_reg/NET0131 , \WX9810_reg/NET0131 , \WX9812_reg/NET0131 , \WX9814_reg/NET0131 , \WX9816_reg/NET0131 , \WX9818_reg/NET0131 , \WX9820_reg/NET0131 , \WX9822_reg/NET0131 , \WX9824_reg/NET0131 , \WX9826_reg/NET0131 , \WX9828_reg/NET0131 , \WX9830_reg/NET0131 , \WX9832_reg/NET0131 , \WX9834_reg/NET0131 , \WX9836_reg/NET0131 , \WX9838_reg/NET0131 , \WX9840_reg/NET0131 , \WX9842_reg/NET0131 , \WX9844_reg/NET0131 , \WX9846_reg/NET0131 , \WX9848_reg/NET0131 , \WX9850_reg/NET0131 , \WX9852_reg/NET0131 , \WX9854_reg/NET0131 , \WX9856_reg/NET0131 , \WX9858_reg/NET0131 , \WX9860_reg/NET0131 , \WX9862_reg/NET0131 , \WX9864_reg/NET0131 , \WX9866_reg/NET0131 , \WX9868_reg/NET0131 , \WX9870_reg/NET0131 , \WX9872_reg/NET0131 , \WX9874_reg/NET0131 , \WX9876_reg/NET0131 , \WX9878_reg/NET0131 , \WX9880_reg/NET0131 , \WX9882_reg/NET0131 , \WX9884_reg/NET0131 , \WX9886_reg/NET0131 , \WX9888_reg/NET0131 , \WX9890_reg/NET0131 , \WX9892_reg/NET0131 , \WX9894_reg/NET0131 , \WX9896_reg/NET0131 , \WX9898_reg/NET0131 , \WX9900_reg/NET0131 , \WX9902_reg/NET0131 , \WX9904_reg/NET0131 , \WX9906_reg/NET0131 , \WX9908_reg/NET0131 , \WX9910_reg/NET0131 , \WX9912_reg/NET0131 , \WX9914_reg/NET0131 , \WX9916_reg/NET0131 , \WX9918_reg/NET0131 , \WX9920_reg/NET0131 , \WX9922_reg/NET0131 , \WX9924_reg/NET0131 , \WX9926_reg/NET0131 , \WX9928_reg/NET0131 , \WX9930_reg/NET0131 , \WX9932_reg/NET0131 , \WX9934_reg/NET0131 , \WX9936_reg/NET0131 , \WX9938_reg/NET0131 , \WX9940_reg/NET0131 , \WX9942_reg/NET0131 , \WX9944_reg/NET0131 , \WX9946_reg/NET0131 , \WX9948_reg/NET0131 , \WX9950_reg/NET0131 , \_2077__reg/NET0131 , \_2078__reg/NET0131 , \_2079__reg/NET0131 , \_2080__reg/NET0131 , \_2081__reg/NET0131 , \_2082__reg/NET0131 , \_2083__reg/NET0131 , \_2084__reg/NET0131 , \_2085__reg/NET0131 , \_2086__reg/NET0131 , \_2087__reg/NET0131 , \_2088__reg/NET0131 , \_2089__reg/NET0131 , \_2090__reg/NET0131 , \_2091__reg/NET0131 , \_2092__reg/NET0131 , \_2093__reg/NET0131 , \_2094__reg/NET0131 , \_2095__reg/NET0131 , \_2096__reg/NET0131 , \_2097__reg/NET0131 , \_2098__reg/NET0131 , \_2099__reg/NET0131 , \_2100__reg/NET0131 , \_2101__reg/NET0131 , \_2102__reg/NET0131 , \_2103__reg/NET0131 , \_2104__reg/NET0131 , \_2105__reg/NET0131 , \_2106__reg/NET0131 , \_2107__reg/NET0131 , \_2108__reg/NET0131 , \_2109__reg/NET0131 , \_2110__reg/NET0131 , \_2111__reg/NET0131 , \_2112__reg/NET0131 , \_2113__reg/NET0131 , \_2114__reg/NET0131 , \_2115__reg/NET0131 , \_2116__reg/NET0131 , \_2117__reg/NET0131 , \_2118__reg/NET0131 , \_2119__reg/NET0131 , \_2120__reg/NET0131 , \_2121__reg/NET0131 , \_2122__reg/NET0131 , \_2123__reg/NET0131 , \_2124__reg/NET0131 , \_2125__reg/NET0131 , \_2126__reg/NET0131 , \_2127__reg/NET0131 , \_2128__reg/NET0131 , \_2129__reg/NET0131 , \_2130__reg/NET0131 , \_2131__reg/NET0131 , \_2132__reg/NET0131 , \_2133__reg/NET0131 , \_2134__reg/NET0131 , \_2135__reg/NET0131 , \_2136__reg/NET0131 , \_2137__reg/NET0131 , \_2138__reg/NET0131 , \_2139__reg/NET0131 , \_2140__reg/NET0131 , \_2141__reg/NET0131 , \_2142__reg/NET0131 , \_2143__reg/NET0131 , \_2144__reg/NET0131 , \_2145__reg/NET0131 , \_2146__reg/NET0131 , \_2147__reg/NET0131 , \_2148__reg/NET0131 , \_2149__reg/NET0131 , \_2150__reg/NET0131 , \_2151__reg/NET0131 , \_2152__reg/NET0131 , \_2153__reg/NET0131 , \_2154__reg/NET0131 , \_2155__reg/NET0131 , \_2156__reg/NET0131 , \_2157__reg/NET0131 , \_2158__reg/NET0131 , \_2159__reg/NET0131 , \_2160__reg/NET0131 , \_2161__reg/NET0131 , \_2162__reg/NET0131 , \_2163__reg/NET0131 , \_2164__reg/NET0131 , \_2165__reg/NET0131 , \_2166__reg/NET0131 , \_2167__reg/NET0131 , \_2168__reg/NET0131 , \_2169__reg/NET0131 , \_2170__reg/NET0131 , \_2171__reg/NET0131 , \_2172__reg/NET0131 , \_2173__reg/NET0131 , \_2174__reg/NET0131 , \_2175__reg/NET0131 , \_2176__reg/NET0131 , \_2177__reg/NET0131 , \_2178__reg/NET0131 , \_2179__reg/NET0131 , \_2180__reg/NET0131 , \_2181__reg/NET0131 , \_2182__reg/NET0131 , \_2183__reg/NET0131 , \_2184__reg/NET0131 , \_2185__reg/NET0131 , \_2186__reg/NET0131 , \_2187__reg/NET0131 , \_2188__reg/NET0131 , \_2189__reg/NET0131 , \_2190__reg/NET0131 , \_2191__reg/NET0131 , \_2192__reg/NET0131 , \_2193__reg/NET0131 , \_2194__reg/NET0131 , \_2195__reg/NET0131 , \_2196__reg/NET0131 , \_2197__reg/NET0131 , \_2198__reg/NET0131 , \_2199__reg/NET0131 , \_2200__reg/NET0131 , \_2201__reg/NET0131 , \_2202__reg/NET0131 , \_2203__reg/NET0131 , \_2204__reg/NET0131 , \_2205__reg/NET0131 , \_2206__reg/NET0131 , \_2207__reg/NET0131 , \_2208__reg/NET0131 , \_2209__reg/NET0131 , \_2210__reg/NET0131 , \_2211__reg/NET0131 , \_2212__reg/NET0131 , \_2213__reg/NET0131 , \_2214__reg/NET0131 , \_2215__reg/NET0131 , \_2216__reg/NET0131 , \_2217__reg/NET0131 , \_2218__reg/NET0131 , \_2219__reg/NET0131 , \_2220__reg/NET0131 , \_2221__reg/NET0131 , \_2222__reg/NET0131 , \_2223__reg/NET0131 , \_2224__reg/NET0131 , \_2225__reg/NET0131 , \_2226__reg/NET0131 , \_2227__reg/NET0131 , \_2228__reg/NET0131 , \_2229__reg/NET0131 , \_2230__reg/NET0131 , \_2231__reg/NET0131 , \_2232__reg/NET0131 , \_2233__reg/NET0131 , \_2234__reg/NET0131 , \_2235__reg/NET0131 , \_2236__reg/NET0131 , \_2237__reg/NET0131 , \_2238__reg/NET0131 , \_2239__reg/NET0131 , \_2240__reg/NET0131 , \_2241__reg/NET0131 , \_2242__reg/NET0131 , \_2243__reg/NET0131 , \_2244__reg/NET0131 , \_2245__reg/NET0131 , \_2246__reg/NET0131 , \_2247__reg/NET0131 , \_2248__reg/NET0131 , \_2249__reg/NET0131 , \_2250__reg/NET0131 , \_2251__reg/NET0131 , \_2252__reg/NET0131 , \_2253__reg/NET0131 , \_2254__reg/NET0131 , \_2255__reg/NET0131 , \_2256__reg/NET0131 , \_2257__reg/NET0131 , \_2258__reg/NET0131 , \_2259__reg/NET0131 , \_2260__reg/NET0131 , \_2261__reg/NET0131 , \_2262__reg/NET0131 , \_2263__reg/NET0131 , \_2264__reg/NET0131 , \_2265__reg/NET0131 , \_2266__reg/NET0131 , \_2267__reg/NET0131 , \_2268__reg/NET0131 , \_2269__reg/NET0131 , \_2270__reg/NET0131 , \_2271__reg/NET0131 , \_2272__reg/NET0131 , \_2273__reg/NET0131 , \_2274__reg/NET0131 , \_2275__reg/NET0131 , \_2276__reg/NET0131 , \_2277__reg/NET0131 , \_2278__reg/NET0131 , \_2279__reg/NET0131 , \_2280__reg/NET0131 , \_2281__reg/NET0131 , \_2282__reg/NET0131 , \_2283__reg/NET0131 , \_2284__reg/NET0131 , \_2285__reg/NET0131 , \_2286__reg/NET0131 , \_2287__reg/NET0131 , \_2288__reg/NET0131 , \_2289__reg/NET0131 , \_2290__reg/NET0131 , \_2291__reg/NET0131 , \_2292__reg/NET0131 , \_2293__reg/NET0131 , \_2294__reg/NET0131 , \_2295__reg/NET0131 , \_2296__reg/NET0131 , \_2297__reg/NET0131 , \_2298__reg/NET0131 , \_2299__reg/NET0131 , \_2300__reg/NET0131 , \_2301__reg/NET0131 , \_2302__reg/NET0131 , \_2303__reg/NET0131 , \_2304__reg/NET0131 , \_2305__reg/NET0131 , \_2306__reg/NET0131 , \_2307__reg/NET0131 , \_2308__reg/NET0131 , \_2309__reg/NET0131 , \_2310__reg/NET0131 , \_2311__reg/NET0131 , \_2312__reg/NET0131 , \_2313__reg/NET0131 , \_2314__reg/NET0131 , \_2315__reg/NET0131 , \_2316__reg/NET0131 , \_2317__reg/NET0131 , \_2318__reg/NET0131 , \_2319__reg/NET0131 , \_2320__reg/NET0131 , \_2321__reg/NET0131 , \_2322__reg/NET0131 , \_2323__reg/NET0131 , \_2324__reg/NET0131 , \_2325__reg/NET0131 , \_2326__reg/NET0131 , \_2327__reg/NET0131 , \_2328__reg/NET0131 , \_2329__reg/NET0131 , \_2330__reg/NET0131 , \_2331__reg/NET0131 , \_2332__reg/NET0131 , \_2333__reg/NET0131 , \_2334__reg/NET0131 , \_2335__reg/NET0131 , \_2336__reg/NET0131 , \_2337__reg/NET0131 , \_2338__reg/NET0131 , \_2339__reg/NET0131 , \_2340__reg/NET0131 , \_2341__reg/NET0131 , \_2342__reg/NET0131 , \_2343__reg/NET0131 , \_2344__reg/NET0131 , \_2345__reg/NET0131 , \_2346__reg/NET0131 , \_2347__reg/NET0131 , \_2348__reg/NET0131 , \_2349__reg/NET0131 , \_2350__reg/NET0131 , \_2351__reg/NET0131 , \_2352__reg/NET0131 , \_2353__reg/NET0131 , \_2354__reg/NET0131 , \_2355__reg/NET0131 , \_2356__reg/NET0131 , \_2357__reg/NET0131 , \_2358__reg/NET0131 , \_2359__reg/NET0131 , \_2360__reg/NET0131 , \_2361__reg/NET0131 , \_2362__reg/NET0131 , \_2363__reg/NET0131 , \_2364__reg/NET0131 , \DATA_9_0_pad , \DATA_9_10_pad , \DATA_9_11_pad , \DATA_9_12_pad , \DATA_9_13_pad , \DATA_9_14_pad , \DATA_9_15_pad , \DATA_9_16_pad , \DATA_9_17_pad , \DATA_9_18_pad , \DATA_9_19_pad , \DATA_9_1_pad , \DATA_9_20_pad , \DATA_9_21_pad , \DATA_9_22_pad , \DATA_9_23_pad , \DATA_9_24_pad , \DATA_9_25_pad , \DATA_9_26_pad , \DATA_9_27_pad , \DATA_9_28_pad , \DATA_9_29_pad , \DATA_9_2_pad , \DATA_9_30_pad , \DATA_9_31_pad , \DATA_9_3_pad , \DATA_9_4_pad , \DATA_9_5_pad , \DATA_9_6_pad , \DATA_9_7_pad , \DATA_9_8_pad , \DATA_9_9_pad , \_al_n0 , \_al_n1 , \g19/_0_ , \g35/_0_ , \g36/_0_ , \g40/_0_ , \g55780/_0_ , \g55783/_0_ , \g55795/_0_ , \g55796/_0_ , \g55797/_0_ , \g55798/_0_ , \g55799/_0_ , \g55800/_0_ , \g55801/_0_ , \g55802/_0_ , \g55803/_0_ , \g55834/_0_ , \g55835/_0_ , \g55836/_0_ , \g55837/_0_ , \g55838/_0_ , \g55839/_0_ , \g55840/_0_ , \g55841/_0_ , \g55842/_0_ , \g55856/_0_ , \g55894/_0_ , \g55895/_0_ , \g55896/_0_ , \g55897/_0_ , \g55898/_0_ , \g55899/_0_ , \g55900/_0_ , \g55901/_0_ , \g55902/_0_ , \g55916/_0_ , \g55953/_0_ , \g55954/_0_ , \g55955/_0_ , \g55956/_0_ , \g55957/_0_ , \g55958/_0_ , \g55959/_0_ , \g55960/_0_ , \g55961/_0_ , \g55975/_0_ , \g56012/_0_ , \g56013/_0_ , \g56014/_0_ , \g56015/_0_ , \g56016/_0_ , \g56017/_0_ , \g56018/_0_ , \g56019/_0_ , \g56020/_0_ , \g56034/_0_ , \g56071/_0_ , \g56072/_0_ , \g56073/_0_ , \g56074/_0_ , \g56075/_0_ , \g56076/_0_ , \g56077/_0_ , \g56078/_0_ , \g56079/_0_ , \g56093/_0_ , \g56130/_0_ , \g56131/_0_ , \g56132/_0_ , \g56133/_0_ , \g56134/_0_ , \g56135/_0_ , \g56136/_0_ , \g56137/_0_ , \g56138/_0_ , \g56152/_0_ , \g56189/_0_ , \g56190/_0_ , \g56191/_0_ , \g56192/_0_ , \g56193/_0_ , \g56194/_0_ , \g56195/_0_ , \g56196/_0_ , \g56197/_0_ , \g56211/_0_ , \g56248/_0_ , \g56249/_0_ , \g56250/_0_ , \g56251/_0_ , \g56252/_0_ , \g56253/_0_ , \g56254/_0_ , \g56255/_0_ , \g56256/_0_ , \g56270/_0_ , \g56307/_0_ , \g56308/_0_ , \g56309/_0_ , \g56310/_0_ , \g56311/_0_ , \g56312/_0_ , \g56313/_0_ , \g56314/_0_ , \g56315/_0_ , \g56329/_0_ , \g56366/_0_ , \g56367/_0_ , \g56368/_0_ , \g56369/_0_ , \g56370/_0_ , \g56371/_0_ , \g56372/_0_ , \g56373/_0_ , \g56374/_0_ , \g56388/_0_ , \g56425/_0_ , \g56426/_0_ , \g56427/_0_ , \g56428/_0_ , \g56429/_0_ , \g56430/_0_ , \g56431/_0_ , \g56432/_0_ , \g56433/_0_ , \g56447/_0_ , \g56484/_0_ , \g56485/_0_ , \g56486/_0_ , \g56487/_0_ , \g56488/_0_ , \g56489/_0_ , \g56490/_0_ , \g56491/_0_ , \g56492/_0_ , \g56507/_0_ , \g56543/_0_ , \g56544/_0_ , \g56545/_0_ , \g56546/_0_ , \g56547/_0_ , \g56548/_0_ , \g56549/_0_ , \g56551/_0_ , \g56567/_0_ , \g56602/_0_ , \g56603/_0_ , \g56604/_0_ , \g56605/_0_ , \g56606/_0_ , \g56607/_0_ , \g56608/_0_ , \g56610/_0_ , \g56627/_0_ , \g56661/_0_ , \g56662/_0_ , \g56663/_0_ , \g56664/_0_ , \g56665/_0_ , \g56666/_0_ , \g56667/_0_ , \g56668/_0_ , \g56686/_0_ , \g56720/_0_ , \g56721/_0_ , \g56722/_0_ , \g56723/_0_ , \g56724/_0_ , \g56725/_0_ , \g56726/_0_ , \g56727/_0_ , \g56728/_0_ , \g56745/_0_ , \g56779/_0_ , \g56780/_0_ , \g56781/_0_ , \g56782/_0_ , \g56783/_0_ , \g56784/_0_ , \g56785/_0_ , \g56804/_0_ , \g56838/_0_ , \g56839/_0_ , \g56840/_0_ , \g56841/_0_ , \g56842/_0_ , \g56843/_0_ , \g56844/_0_ , \g56845/_0_ , \g56846/_0_ , \g56863/_0_ , \g56897/_0_ , \g56898/_0_ , \g56899/_0_ , \g56900/_0_ , \g56901/_0_ , \g56902/_0_ , \g56903/_0_ , \g56905/_0_ , \g56921/_0_ , \g56956/_0_ , \g56957/_0_ , \g56958/_0_ , \g56959/_0_ , \g56960/_0_ , \g56961/_0_ , \g56962/_0_ , \g56964/_0_ , \g56980/_0_ , \g57015/_0_ , \g57016/_0_ , \g57017/_0_ , \g57018/_0_ , \g57019/_0_ , \g57020/_0_ , \g57021/_0_ , \g57023/_0_ , \g57040/_0_ , \g57074/_0_ , \g57075/_0_ , \g57076/_0_ , \g57077/_0_ , \g57078/_0_ , \g57079/_0_ , \g57080/_0_ , \g57081/_0_ , \g57099/_0_ , \g57133/_0_ , \g57134/_0_ , \g57135/_0_ , \g57136/_0_ , \g57137/_0_ , \g57138/_0_ , \g57139/_0_ , \g57140/_0_ , \g57141/_0_ , \g57159/_0_ , \g57193/_0_ , \g57195/_0_ , \g57196/_0_ , \g57197/_0_ , \g57198/_0_ , \g57199/_0_ , \g57200/_0_ , \g57202/_0_ , \g57219/_0_ , \g57254/_0_ , \g57255/_0_ , \g57256/_0_ , \g57257/_0_ , \g57258/_0_ , \g57259/_0_ , \g57260/_0_ , \g57262/_0_ , \g57263/_0_ , \g57285/_0_ , \g57318/_0_ , \g57319/_0_ , \g57320/_0_ , \g57321/_0_ , \g57322/_0_ , \g57323/_0_ , \g57324/_0_ , \g57325/_0_ , \g57326/_0_ , \g57328/_0_ , \g57329/_0_ , \g57330/_0_ , \g57350/_0_ , \g57387/_0_ , \g57388/_0_ , \g57390/_0_ , \g57391/_0_ , \g57392/_0_ , \g57393/_0_ , \g57395/_0_ , \g57396/_0_ , \g57439/_0_ , \g57476/_0_ , \g57477/_0_ , \g57478/_0_ , \g57479/_0_ , \g57480/_0_ , \g57481/_0_ , \g57482/_0_ , \g57483/_0_ , \g57484/_0_ , \g57485/_0_ , \g57486/_0_ , \g57487/_0_ , \g57488/_0_ , \g57489/_0_ , \g57490/_0_ , \g57491/_0_ , \g57492/_0_ , \g57493/_0_ , \g57494/_0_ , \g57495/_0_ , \g57496/_0_ , \g57497/_0_ , \g57498/_0_ , \g57499/_0_ , \g57500/_0_ , \g57501/_0_ , \g57502/_0_ , \g57503/_0_ , \g57504/_0_ , \g57505/_0_ , \g57524/_0_ , \g57537/_0_ , \g57541/_0_ , \g57543/_0_ , \g58163/_0_ , \g58572/_0_ , \g58573/_0_ , \g58574/_0_ , \g58575/_0_ , \g58576/_0_ , \g58577/_0_ , \g58578/_0_ , \g58579/_0_ , \g58580/_0_ , \g58581/_0_ , \g58582/_0_ , \g58583/_0_ , \g58584/_0_ , \g58585/_0_ , \g58586/_0_ , \g58587/_0_ , \g58588/_0_ , \g58589/_0_ , \g58590/_0_ , \g58591/_0_ , \g58592/_0_ , \g58593/_0_ , \g58594/_0_ , \g58595/_0_ , \g58596/_0_ , \g58597/_0_ , \g58598/_0_ , \g58600/_0_ , \g58602/_0_ , \g58604/_0_ , \g58615/_0_ , \g59240/_0_ , \g59241/_0_ , \g59242/_0_ , \g59243/_0_ , \g59244/_0_ , \g59245/_0_ , \g59246/_0_ , \g59247/_0_ , \g59248/_0_ , \g59249/_0_ , \g59250/_0_ , \g59251/_0_ , \g59252/_0_ , \g59253/_0_ , \g59254/_0_ , \g59255/_0_ , \g59256/_0_ , \g59257/_0_ , \g59258/_0_ , \g59259/_0_ , \g59260/_0_ , \g59261/_0_ , \g59262/_0_ , \g59263/_0_ , \g59264/_0_ , \g59265/_0_ , \g59266/_0_ , \g59267/_0_ , \g59268/_0_ , \g59269/_0_ , \g59270/_0_ , \g59271/_0_ , \g59272/_0_ , \g59273/_0_ , \g59274/_0_ , \g59275/_0_ , \g59276/_0_ , \g59277/_0_ , \g59278/_0_ , \g59279/_0_ , \g59280/_0_ , \g59281/_0_ , \g59282/_0_ , \g59283/_0_ , \g59284/_0_ , \g59285/_0_ , \g59286/_0_ , \g59287/_0_ , \g59288/_0_ , \g59289/_0_ , \g59290/_0_ , \g59291/_0_ , \g59292/_0_ , \g59293/_0_ , \g59294/_0_ , \g59295/_0_ , \g59296/_0_ , \g59297/_0_ , \g59298/_0_ , \g59299/_0_ , \g59300/_0_ , \g59301/_0_ , \g59302/_0_ , \g59303/_0_ , \g59304/_0_ , \g59305/_0_ , \g59306/_0_ , \g59307/_0_ , \g59308/_0_ , \g59309/_0_ , \g59310/_0_ , \g59311/_0_ , \g59312/_0_ , \g59313/_0_ , \g59314/_0_ , \g59315/_0_ , \g59316/_0_ , \g59317/_0_ , \g59318/_0_ , \g59319/_0_ , \g59320/_0_ , \g59321/_0_ , \g59322/_0_ , \g59323/_0_ , \g59324/_0_ , \g59325/_0_ , \g59326/_0_ , \g59327/_0_ , \g59328/_0_ , \g59329/_0_ , \g59330/_0_ , \g59331/_0_ , \g59332/_0_ , \g59333/_0_ , \g59334/_0_ , \g59335/_0_ , \g59336/_0_ , \g59337/_0_ , \g59338/_0_ , \g59339/_0_ , \g59340/_0_ , \g59341/_0_ , \g59342/_0_ , \g59343/_0_ , \g59344/_0_ , \g59345/_0_ , \g59346/_0_ , \g59347/_0_ , \g59348/_0_ , \g59349/_0_ , \g59350/_0_ , \g59351/_0_ , \g59352/_0_ , \g59353/_0_ , \g59354/_0_ , \g59355/_0_ , \g59356/_0_ , \g59357/_0_ , \g59358/_0_ , \g59359/_0_ , \g59360/_0_ , \g59361/_0_ , \g59362/_0_ , \g59363/_0_ , \g59364/_0_ , \g59365/_0_ , \g59366/_0_ , \g59367/_0_ , \g59368/_0_ , \g59369/_0_ , \g59370/_0_ , \g59371/_0_ , \g59372/_0_ , \g59373/_0_ , \g59374/_0_ , \g59375/_0_ , \g59376/_0_ , \g59377/_0_ , \g59378/_0_ , \g59379/_0_ , \g59380/_0_ , \g59381/_0_ , \g59382/_0_ , \g59383/_0_ , \g59384/_0_ , \g59385/_0_ , \g59386/_0_ , \g59387/_0_ , \g59388/_0_ , \g59389/_0_ , \g59390/_0_ , \g59391/_0_ , \g59392/_0_ , \g59393/_0_ , \g59394/_0_ , \g59395/_0_ , \g59396/_0_ , \g59397/_0_ , \g59398/_0_ , \g59399/_0_ , \g59400/_0_ , \g59401/_0_ , \g59402/_0_ , \g59403/_0_ , \g59404/_0_ , \g59405/_0_ , \g59406/_0_ , \g59407/_0_ , \g59408/_0_ , \g59409/_0_ , \g59410/_0_ , \g59411/_0_ , \g59412/_0_ , \g59413/_0_ , \g59414/_0_ , \g59415/_0_ , \g59416/_0_ , \g59417/_0_ , \g59418/_0_ , \g59419/_0_ , \g59420/_0_ , \g59421/_0_ , \g59422/_0_ , \g59423/_0_ , \g59424/_0_ , \g59425/_0_ , \g59426/_0_ , \g59427/_0_ , \g59428/_0_ , \g59429/_0_ , \g59430/_0_ , \g59431/_0_ , \g59432/_0_ , \g59433/_0_ , \g59434/_0_ , \g59435/_0_ , \g59436/_0_ , \g59437/_0_ , \g59438/_0_ , \g59439/_0_ , \g59440/_0_ , \g59441/_0_ , \g59442/_0_ , \g59443/_0_ , \g59444/_0_ , \g59445/_0_ , \g59446/_0_ , \g59447/_0_ , \g59448/_0_ , \g59449/_0_ , \g59450/_0_ , \g59451/_0_ , \g59452/_0_ , \g59453/_0_ , \g59454/_0_ , \g59455/_0_ , \g59456/_0_ , \g59457/_0_ , \g59458/_0_ , \g59459/_0_ , \g59460/_0_ , \g59461/_0_ , \g59462/_0_ , \g59463/_0_ , \g59464/_0_ , \g59465/_0_ , \g59466/_0_ , \g59467/_0_ , \g59468/_0_ , \g59469/_0_ , \g59470/_0_ , \g59471/_0_ , \g59472/_0_ , \g59473/_0_ , \g59474/_0_ , \g59475/_0_ , \g59476/_0_ , \g59477/_0_ , \g59478/_0_ , \g59479/_0_ , \g59480/_0_ , \g59481/_0_ , \g59482/_0_ , \g59483/_0_ , \g59484/_0_ , \g59485/_0_ , \g59486/_0_ , \g59487/_0_ , \g59488/_0_ , \g59489/_0_ , \g59490/_0_ , \g59491/_0_ , \g59492/_0_ , \g59493/_0_ , \g59494/_0_ , \g59495/_0_ , \g59496/_0_ , \g59497/_0_ , \g59498/_0_ , \g59500/_0_ , \g59503/_0_ , \g59512/_0_ , \g61336/_0_ , \g61521/_0_ , \g61523/_0_ , \g61524/_0_ , \g61526/_0_ , \g61527/_0_ , \g61528/_0_ , \g61529/_0_ , \g61530/_0_ , \g61531/_0_ , \g61532/_0_ , \g61533/_0_ , \g61535/_0_ , \g61537/_0_ , \g61539/_0_ , \g61540/_0_ , \g61541/_0_ , \g61542/_0_ , \g61546/_0_ , \g61550/_0_ , \g61551/_0_ , \g61552/_0_ , \g61554/_0_ , \g61555/_0_ , \g61556/_0_ , \g61558/_0_ , \g61559/_0_ , \g61561/_0_ , \g61562/_0_ , \g61563/_0_ , \g61564/_0_ , \g61565/_0_ , \g61566/_0_ , \g61568/_0_ , \g61570/_0_ , \g61571/_0_ , \g61572/_0_ , \g61573/_0_ , \g61577/_0_ , \g61578/_0_ , \g61579/_0_ , \g61580/_0_ , \g61581/_0_ , \g61582/_0_ , \g61583/_0_ , \g61584/_0_ , \g61585/_0_ , \g61586/_0_ , \g61587/_0_ , \g61588/_0_ , \g61589/_0_ , \g61591/_0_ , \g61592/_0_ , \g61594/_0_ , \g61595/_0_ , \g61596/_0_ , \g61597/_0_ , \g61598/_0_ , \g61599/_0_ , \g61600/_0_ , \g61601/_0_ , \g61605/_0_ , \g61606/_0_ , \g61607/_0_ , \g61608/_0_ , \g61609/_0_ , \g61610/_0_ , \g61611/_0_ , \g61612/_0_ , \g61613/_0_ , \g61615/_0_ , \g61616/_0_ , \g61617/_0_ , \g61618/_0_ , \g61619/_0_ , \g61620/_0_ , \g61621/_0_ , \g61623/_0_ , \g61624/_0_ , \g61625/_0_ , \g61626/_0_ , \g61627/_0_ , \g61629/_0_ , \g61630/_0_ , \g61631/_0_ , \g61632/_0_ , \g61633/_0_ , \g61634/_0_ , \g61636/_0_ , \g61638/_0_ , \g61639/_0_ , \g61640/_0_ , \g61641/_0_ , \g61642/_0_ , \g61644/_0_ , \g61647/_0_ , \g61648/_0_ , \g61649/_0_ , \g61650/_0_ , \g61653/_0_ , \g61654/_0_ , \g61655/_0_ , \g61656/_0_ , \g61658/_0_ , \g61661/_0_ , \g61662/_0_ , \g61663/_0_ , \g61664/_0_ , \g61666/_0_ , \g61667/_0_ , \g61668/_0_ , \g61670/_0_ , \g61671/_0_ , \g61672/_0_ , \g61673/_0_ , \g61675/_0_ , \g61676/_0_ , \g61680/_0_ , \g61681/_0_ , \g61682/_0_ , \g61683/_0_ , \g61684/_0_ , \g61686/_0_ , \g61687/_0_ , \g61688/_0_ , \g61689/_0_ , \g61690/_0_ , \g61691/_0_ , \g61693/_0_ , \g61694/_0_ , \g61696/_0_ , \g61697/_0_ , \g61698/_0_ , \g61699/_0_ , \g61700/_0_ , \g61701/_0_ , \g61702/_0_ , \g61703/_0_ , \g61704/_0_ , \g61705/_0_ , \g61706/_0_ , \g61707/_0_ , \g61708/_0_ , \g61711/_0_ , \g61712/_0_ , \g61714/_0_ , \g61716/_0_ , \g61717/_0_ , \g61719/_0_ , \g61720/_0_ , \g61721/_0_ , \g61724/_0_ , \g61725/_0_ , \g61728/_0_ , \g61729/_0_ , \g61731/_0_ , \g61732/_0_ , \g61733/_0_ , \g61736/_0_ , \g61737/_0_ , \g61739/_0_ , \g61740/_0_ , \g61741/_0_ , \g61743/_0_ , \g61744/_0_ , \g61745/_0_ , \g61746/_0_ , \g61747/_0_ , \g61748/_0_ , \g61749/_0_ , \g61750/_0_ , \g61751/_0_ , \g61752/_0_ , \g61753/_0_ , \g61754/_0_ , \g61755/_0_ , \g61757/_0_ , \g61758/_0_ , \g61759/_0_ , \g61760/_0_ , \g61761/_0_ , \g61762/_0_ , \g61763/_0_ , \g61764/_0_ , \g61765/_0_ , \g61766/_0_ , \g61767/_0_ , \g61768/_0_ , \g61769/_0_ , \g61770/_0_ , \g61771/_0_ , \g61772/_0_ , \g61773/_0_ , \g61774/_0_ , \g61775/_0_ , \g61776/_0_ , \g61777/_0_ , \g61778/_0_ , \g61780/_0_ , \g61781/_0_ , \g61783/_0_ , \g61784/_0_ , \g61786/_0_ , \g61787/_0_ , \g61790/_0_ , \g61791/_0_ , \g61794/_0_ , \g61795/_0_ , \g61796/_0_ , \g61797/_0_ , \g61798/_0_ , \g61799/_0_ , \g61800/_0_ , \g61801/_0_ , \g61802/_0_ , \g61803/_0_ , \g61805/_0_ , \g61806/_0_ , \g61807/_0_ , \g61808/_0_ , \g61809/_0_ , \g61810/_0_ , \g61811/_0_ , \g61812/_0_ , \g61813/_0_ , \g61816/_0_ , \g61817/_0_ , \g61818/_0_ , \g61820/_0_ , \g61822/_0_ , \g61823/_0_ , \g61825/_0_ , \g61826/_0_ , \g61827/_0_ , \g61828/_0_ , \g61829/_0_ , \g61832/_0_ , \g61834/_0_ , \g61835/_0_ , \g61837/_0_ , \g61838/_0_ , \g61839/_0_ , \g61840/_0_ , \g61844/_0_ , \g61847/_0_ , \g61848/_0_ , \g61849/_0_ , \g61850/_0_ , \g61851/_0_ , \g61853/_0_ , \g61854/_0_ , \g61855/_0_ , \g61856/_0_ , \g61858/_0_ , \g61859/_0_ , \g61861/_0_ , \g61862/_0_ , \g61863/_0_ , \g61864/_0_ , \g61865/_0_ , \g61866/_0_ , \g61867/_0_ , \g61868/_0_ , \g61869/_0_ , \g61870/_0_ , \g61871/_0_ , \g61873/_0_ , \g61874/_0_ , \g61875/_0_ , \g61877/_0_ , \g61878/_0_ , \g61879/_0_ , \g61880/_0_ , \g61881/_0_ , \g61883/_0_ , \g61884/_0_ , \g61886/_0_ , \g61887/_0_ , \g61890/_0_ , \g61891/_0_ , \g61892/_0_ , \g61893/_0_ , \g61894/_0_ , \g61895/_0_ , \g61900/_0_ , \g61901/_0_ , \g61902/_0_ , \g61904/_0_ , \g61905/_0_ , \g61906/_0_ , \g61907/_0_ , \g61914/_0_ , \g61915/_0_ , \g61917/_0_ , \g61919/_0_ , \g61921/_0_ , \g61924/_0_ , \g61925/_0_ , \g61926/_0_ , \g61927/_0_ , \g61928/_0_ , \g61929/_0_ , \g61930/_0_ , \g61931/_0_ , \g61932/_0_ , \g61933/_0_ , \g61934/_0_ , \g61935/_0_ , \g61936/_0_ , \g61937/_0_ , \g61938/_0_ , \g61939/_0_ , \g61943/_0_ , \g61944/_0_ , \g61945/_0_ , \g61947/_0_ , \g61948/_0_ , \g61949/_0_ , \g61950/_0_ , \g61951/_0_ , \g61952/_0_ , \g61953/_0_ , \g61955/_0_ , \g61956/_0_ , \g61957/_0_ , \g61958/_0_ , \g61959/_0_ , \g61960/_0_ , \g61961/_0_ , \g61962/_0_ , \g61963/_0_ , \g61964/_0_ , \g61965/_0_ , \g61966/_0_ , \g61967/_0_ , \g61968/_0_ , \g61969/_0_ , \g61970/_0_ , \g61971/_0_ , \g61972/_0_ , \g61973/_0_ , \g61974/_0_ , \g61976/_0_ , \g61978/_0_ , \g61980/_0_ , \g61981/_0_ , \g61982/_0_ , \g61983/_0_ , \g61984/_0_ , \g61985/_0_ , \g61986/_0_ , \g61987/_0_ , \g61988/_0_ , \g61989/_0_ , \g61990/_0_ , \g61992/_0_ , \g61994/_0_ , \g61995/_0_ , \g61996/_0_ , \g61997/_0_ , \g61998/_0_ , \g62000/_0_ , \g62001/_0_ , \g62002/_0_ , \g62003/_0_ , \g62004/_0_ , \g62005/_0_ , \g62007/_0_ , \g62008/_0_ , \g62009/_0_ , \g62010/_0_ , \g62011/_0_ , \g62012/_0_ , \g62013/_0_ , \g62014/_0_ , \g62015/_0_ , \g62016/_0_ , \g62017/_0_ , \g62018/_0_ , \g62019/_0_ , \g62020/_0_ , \g62021/_0_ , \g62022/_0_ , \g62023/_0_ , \g62024/_0_ , \g62025/_0_ , \g62026/_0_ , \g62027/_0_ , \g62030/_0_ , \g62033/_0_ , \g62034/_0_ , \g62036/_0_ , \g62038/_0_ , \g62041/_0_ , \g62042/_0_ , \g62043/_0_ , \g62044/_0_ , \g62045/_0_ , \g62046/_0_ , \g62047/_0_ , \g62048/_0_ , \g62050/_0_ , \g62051/_0_ , \g62052/_0_ , \g62055/_0_ , \g62057/_0_ , \g62058/_0_ , \g62059/_0_ , \g62060/_0_ , \g62061/_0_ , \g62062/_0_ , \g62064/_0_ , \g62065/_0_ , \g62066/_0_ , \g62067/_0_ , \g62068/_0_ , \g62072/_0_ , \g62073/_0_ , \g62074/_0_ , \g62075/_0_ , \g62076/_0_ , \g62077/_0_ , \g62078/_0_ , \g62080/_0_ , \g62081/_0_ , \g62082/_0_ , \g62084/_0_ , \g62085/_0_ , \g62086/_0_ , \g62087/_0_ , \g62088/_0_ , \g62089/_0_ , \g62090/_0_ , \g62091/_0_ , \g62092/_0_ , \g62094/_0_ , \g62096/_0_ , \g62097/_0_ , \g62098/_0_ , \g62099/_0_ , \g62100/_0_ , \g62101/_0_ , \g62102/_0_ , \g62104/_0_ , \g62106/_0_ , \g62107/_0_ , \g62108/_0_ , \g62110/_0_ , \g62112/_0_ , \g62113/_0_ , \g62114/_0_ , \g62116/_0_ , \g62117/_0_ , \g62118/_0_ , \g62119/_0_ , \g62120/_0_ , \g62121/_0_ , \g62122/_0_ , \g62124/_0_ , \g62126/_0_ , \g62127/_0_ , \g62128/_0_ , \g62129/_0_ , \g62130/_0_ , \g62131/_0_ , \g62132/_0_ , \g62133/_0_ , \g62135/_0_ , \g62136/_0_ , \g62137/_0_ , \g62138/_0_ , \g62140/_0_ , \g62143/_0_ , \g62144/_0_ , \g62149/_0_ , \g62150/_0_ , \g62151/_0_ , \g62153/_0_ , \g62155/_0_ , \g62156/_0_ , \g62158/_0_ , \g62160/_0_ , \g62161/_0_ , \g62162/_0_ , \g62164/_0_ , \g62165/_0_ , \g62166/_0_ , \g62167/_0_ , \g62168/_0_ , \g62169/_0_ , \g62172/_0_ , \g62173/_0_ , \g62175/_0_ , \g62176/_0_ , \g62177/_0_ , \g62178/_0_ , \g62179/_0_ , \g62180/_0_ , \g62181/_0_ , \g62182/_0_ , \g62183/_0_ , \g62184/_0_ , \g62185/_0_ , \g62186/_0_ , \g62188/_0_ , \g62189/_0_ , \g62190/_0_ , \g62191/_0_ , \g62193/_0_ , \g62194/_0_ , \g62195/_0_ , \g62196/_0_ , \g62197/_0_ , \g62200/_0_ , \g62201/_0_ , \g62202/_0_ , \g62203/_0_ , \g62205/_0_ , \g62206/_0_ , \g62207/_0_ , \g62208/_0_ , \g62209/_0_ , \g62210/_0_ , \g62211/_0_ , \g62215/_0_ , \g62218/_0_ , \g62219/_0_ , \g62221/_0_ , \g62222/_0_ , \g62223/_0_ , \g62224/_0_ , \g62225/_0_ , \g62226/_0_ , \g62229/_0_ , \g62230/_0_ , \g62231/_0_ , \g62233/_0_ , \g62236/_0_ , \g62237/_0_ , \g62238/_0_ , \g62240/_0_ , \g62241/_0_ , \g62243/_0_ , \g62244/_0_ , \g62245/_0_ , \g62247/_0_ , \g62248/_0_ , \g62250/_0_ , \g62252/_0_ , \g62253/_0_ , \g62255/_0_ , \g62256/_0_ , \g62257/_0_ , \g62258/_0_ , \g62259/_0_ , \g62260/_0_ , \g62261/_0_ , \g62262/_0_ , \g62263/_0_ , \g62264/_0_ , \g62265/_0_ , \g62267/_0_ , \g62269/_0_ , \g62270/_0_ , \g62272/_0_ , \g62274/_0_ , \g62277/_0_ , \g62279/_0_ , \g62280/_0_ , \g62281/_0_ , \g62283/_0_ , \g62284/_0_ , \g62285/_0_ , \g62286/_0_ , \g62288/_0_ , \g62289/_0_ , \g62290/_0_ , \g62294/_0_ , \g62295/_0_ , \g62296/_0_ , \g62297/_0_ , \g62298/_0_ , \g62299/_0_ , \g62303/_0_ , \g62305/_0_ , \g62306/_0_ , \g62307/_0_ , \g62309/_0_ , \g62311/_0_ , \g62312/_0_ , \g62313/_0_ , \g62314/_0_ , \g62315/_0_ , \g62316/_0_ , \g62317/_0_ , \g62318/_0_ , \g62319/_0_ , \g62320/_0_ , \g62322/_0_ , \g62324/_0_ , \g62325/_0_ , \g62326/_0_ , \g62327/_0_ , \g62329/_0_ , \g62330/_0_ , \g62331/_0_ , \g62332/_0_ , \g62333/_0_ , \g62335/_0_ , \g62336/_0_ , \g62338/_0_ , \g62341/_0_ , \g62342/_0_ , \g62344/_0_ , \g62345/_0_ , \g62348/_0_ , \g62349/_0_ , \g62350/_0_ , \g62353/_0_ , \g62354/_0_ , \g62355/_0_ , \g62356/_0_ , \g62359/_0_ , \g62362/_0_ , \g62363/_0_ , \g62364/_0_ , \g62365/_0_ , \g62366/_0_ , \g62367/_0_ , \g62368/_0_ , \g62369/_0_ , \g62370/_0_ , \g62371/_0_ , \g62372/_0_ , \g62373/_0_ , \g62374/_0_ , \g62376/_0_ , \g62467/_0_ , \g62468/_0_ , \g62469/_0_ , \g62470/_0_ , \g62471/_0_ , \g62472/_0_ , \g62473/_0_ , \g62474/_0_ , \g62475/_0_ , \g62478/_0_ , \g62480/_0_ , \g62481/_0_ , \g62482/_0_ , \g62483/_0_ , \g62484/_0_ , \g62485/_0_ , \g62486/_0_ , \g62487/_0_ , \g62488/_0_ , \g62489/_0_ , \g62490/_0_ , \g62491/_0_ , \g62492/_0_ , \g62493/_0_ , \g62494/_0_ , \g62495/_0_ , \g62496/_0_ , \g62497/_0_ , \g62498/_0_ , \g62499/_0_ , \g62500/_0_ , \g62501/_0_ , \g62502/_0_ , \g62503/_0_ , \g62504/_0_ , \g62509/_0_ , \g62510/_0_ , \g62511/_0_ , \g62512/_0_ , \g62513/_0_ , \g62514/_0_ , \g62515/_0_ , \g62516/_0_ , \g62517/_0_ , \g62518/_0_ , \g62519/_0_ , \g62520/_0_ , \g62521/_0_ , \g62523/_0_ , \g62526/_0_ , \g62528/_0_ , \g62529/_0_ , \g62531/_0_ , \g62532/_0_ , \g62533/_0_ , \g62534/_0_ , \g62535/_0_ , \g62536/_0_ , \g62537/_0_ , \g62539/_0_ , \g62540/_0_ , \g62541/_0_ , \g62542/_0_ , \g62543/_0_ , \g62544/_0_ , \g62545/_0_ , \g62547/_0_ , \g62548/_0_ , \g62549/_0_ , \g62550/_0_ , \g62551/_0_ , \g62552/_0_ , \g62553/_0_ , \g62554/_0_ , \g62555/_0_ , \g62556/_0_ , \g62557/_0_ , \g62560/_0_ , \g62562/_0_ , \g62563/_0_ , \g62564/_0_ , \g62565/_0_ , \g62566/_0_ , \g62567/_0_ , \g62569/_0_ , \g62570/_0_ , \g62571/_0_ , \g62572/_0_ , \g62573/_0_ , \g62574/_0_ , \g62576/_0_ , \g62577/_0_ , \g62581/_0_ , \g62582/_0_ , \g62584/_0_ , \g62585/_0_ , \g62586/_0_ , \g62588/_0_ , \g62589/_0_ , \g62593/_0_ , \g62594/_0_ , \g62595/_0_ , \g62596/_0_ , \g62597/_0_ , \g62598/_0_ , \g62599/_0_ , \g62600/_0_ , \g62601/_0_ , \g62602/_0_ , \g62603/_0_ , \g62604/_0_ , \g62605/_0_ , \g62606/_0_ , \g62607/_0_ , \g62608/_0_ , \g62609/_0_ , \g62610/_0_ , \g62612/_0_ , \g62613/_0_ , \g62614/_0_ , \g62615/_0_ , \g62617/_0_ , \g62618/_0_ , \g62620/_0_ , \g62621/_0_ , \g62622/_0_ , \g62624/_0_ , \g62625/_0_ , \g62626/_0_ , \g62627/_0_ , \g62629/_0_ , \g62630/_0_ , \g62632/_0_ , \g62633/_0_ , \g62635/_0_ , \g62636/_0_ , \g62637/_0_ , \g62638/_0_ , \g62640/_0_ , \g62641/_0_ , \g62642/_0_ , \g62643/_0_ , \g62644/_0_ , \g62646/_0_ , \g62647/_0_ , \g62649/_0_ , \g62650/_0_ , \g62651/_0_ , \g62653/_0_ , \g62655/_0_ , \g62656/_0_ , \g62657/_0_ , \g62658/_0_ , \g62660/_0_ , \g62661/_0_ , \g62662/_0_ , \g62663/_0_ , \g62664/_0_ , \g62665/_0_ , \g62667/_0_ , \g62669/_0_ , \g62670/_0_ , \g62671/_0_ , \g62672/_0_ , \g62674/_0_ , \g62675/_0_ , \g62676/_0_ , \g62677/_0_ , \g62678/_0_ , \g62679/_0_ , \g62680/_0_ , \g62681/_0_ , \g62682/_0_ , \g62684/_0_ , \g62685/_0_ , \g62686/_0_ , \g62687/_0_ , \g62690/_0_ , \g62693/_0_ , \g62698/_0_ , \g62699/_0_ , \g62700/_0_ , \g62701/_0_ , \g62702/_0_ , \g62703/_0_ , \g62704/_0_ , \g62709/_0_ , \g62710/_0_ , \g62711/_0_ , \g62714/_0_ , \g62715/_0_ , \g62717/_0_ , \g62718/_0_ , \g62719/_0_ , \g62720/_0_ , \g62721/_0_ , \g62723/_0_ , \g62725/_0_ , \g62726/_0_ , \g62729/_0_ , \g62731/_0_ , \g62733/_0_ , \g62738/_0_ , \g62741/_0_ , \g62742/_0_ , \g62744/_0_ , \g62745/_0_ , \g62746/_0_ , \g62747/_0_ , \g62748/_0_ , \g62749/_0_ , \g62753/_0_ , \g62755/_0_ , \g62756/_0_ , \g62758/_0_ , \g62759/_0_ , \g62760/_0_ , \g62761/_0_ , \g62763/_0_ , \g62766/_0_ , \g62767/_0_ , \g62768/_0_ , \g65554/_0_ , \g65561/_0_ , \g65569/_0_ , \g65580/_0_ , \g65599/_0_ , \g65606/_0_ , \g65636/_0_ , \g65864/_0_ );
	input \DATA_0_0_pad  ;
	input \DATA_0_10_pad  ;
	input \DATA_0_11_pad  ;
	input \DATA_0_12_pad  ;
	input \DATA_0_13_pad  ;
	input \DATA_0_14_pad  ;
	input \DATA_0_15_pad  ;
	input \DATA_0_16_pad  ;
	input \DATA_0_17_pad  ;
	input \DATA_0_18_pad  ;
	input \DATA_0_19_pad  ;
	input \DATA_0_1_pad  ;
	input \DATA_0_20_pad  ;
	input \DATA_0_21_pad  ;
	input \DATA_0_22_pad  ;
	input \DATA_0_23_pad  ;
	input \DATA_0_24_pad  ;
	input \DATA_0_25_pad  ;
	input \DATA_0_26_pad  ;
	input \DATA_0_27_pad  ;
	input \DATA_0_28_pad  ;
	input \DATA_0_29_pad  ;
	input \DATA_0_2_pad  ;
	input \DATA_0_30_pad  ;
	input \DATA_0_31_pad  ;
	input \DATA_0_3_pad  ;
	input \DATA_0_4_pad  ;
	input \DATA_0_5_pad  ;
	input \DATA_0_6_pad  ;
	input \DATA_0_7_pad  ;
	input \DATA_0_8_pad  ;
	input \DATA_0_9_pad  ;
	input RESET_pad ;
	input \TM0_pad  ;
	input \TM1_pad  ;
	input \WX10829_reg/NET0131  ;
	input \WX10831_reg/NET0131  ;
	input \WX10833_reg/NET0131  ;
	input \WX10835_reg/NET0131  ;
	input \WX10837_reg/NET0131  ;
	input \WX10839_reg/NET0131  ;
	input \WX10841_reg/NET0131  ;
	input \WX10843_reg/NET0131  ;
	input \WX10845_reg/NET0131  ;
	input \WX10847_reg/NET0131  ;
	input \WX10849_reg/NET0131  ;
	input \WX10851_reg/NET0131  ;
	input \WX10853_reg/NET0131  ;
	input \WX10855_reg/NET0131  ;
	input \WX10857_reg/NET0131  ;
	input \WX10859_reg/NET0131  ;
	input \WX10861_reg/NET0131  ;
	input \WX10863_reg/NET0131  ;
	input \WX10865_reg/NET0131  ;
	input \WX10867_reg/NET0131  ;
	input \WX10869_reg/NET0131  ;
	input \WX10871_reg/NET0131  ;
	input \WX10873_reg/NET0131  ;
	input \WX10875_reg/NET0131  ;
	input \WX10877_reg/NET0131  ;
	input \WX10879_reg/NET0131  ;
	input \WX10881_reg/NET0131  ;
	input \WX10883_reg/NET0131  ;
	input \WX10885_reg/NET0131  ;
	input \WX10887_reg/NET0131  ;
	input \WX10889_reg/NET0131  ;
	input \WX10891_reg/NET0131  ;
	input \WX10989_reg/NET0131  ;
	input \WX10991_reg/NET0131  ;
	input \WX10993_reg/NET0131  ;
	input \WX10995_reg/NET0131  ;
	input \WX10997_reg/NET0131  ;
	input \WX10999_reg/NET0131  ;
	input \WX11001_reg/NET0131  ;
	input \WX11003_reg/NET0131  ;
	input \WX11005_reg/NET0131  ;
	input \WX11007_reg/NET0131  ;
	input \WX11009_reg/NET0131  ;
	input \WX11011_reg/NET0131  ;
	input \WX11013_reg/NET0131  ;
	input \WX11015_reg/NET0131  ;
	input \WX11017_reg/NET0131  ;
	input \WX11019_reg/NET0131  ;
	input \WX11021_reg/NET0131  ;
	input \WX11023_reg/NET0131  ;
	input \WX11025_reg/NET0131  ;
	input \WX11027_reg/NET0131  ;
	input \WX11029_reg/NET0131  ;
	input \WX11031_reg/NET0131  ;
	input \WX11033_reg/NET0131  ;
	input \WX11035_reg/NET0131  ;
	input \WX11037_reg/NET0131  ;
	input \WX11039_reg/NET0131  ;
	input \WX11041_reg/NET0131  ;
	input \WX11043_reg/NET0131  ;
	input \WX11045_reg/NET0131  ;
	input \WX11047_reg/NET0131  ;
	input \WX11049_reg/NET0131  ;
	input \WX11051_reg/NET0131  ;
	input \WX11053_reg/NET0131  ;
	input \WX11055_reg/NET0131  ;
	input \WX11057_reg/NET0131  ;
	input \WX11059_reg/NET0131  ;
	input \WX11061_reg/NET0131  ;
	input \WX11063_reg/NET0131  ;
	input \WX11065_reg/NET0131  ;
	input \WX11067_reg/NET0131  ;
	input \WX11069_reg/NET0131  ;
	input \WX11071_reg/NET0131  ;
	input \WX11073_reg/NET0131  ;
	input \WX11075_reg/NET0131  ;
	input \WX11077_reg/NET0131  ;
	input \WX11079_reg/NET0131  ;
	input \WX11081_reg/NET0131  ;
	input \WX11083_reg/NET0131  ;
	input \WX11085_reg/NET0131  ;
	input \WX11087_reg/NET0131  ;
	input \WX11089_reg/NET0131  ;
	input \WX11091_reg/NET0131  ;
	input \WX11093_reg/NET0131  ;
	input \WX11095_reg/NET0131  ;
	input \WX11097_reg/NET0131  ;
	input \WX11099_reg/NET0131  ;
	input \WX11101_reg/NET0131  ;
	input \WX11103_reg/NET0131  ;
	input \WX11105_reg/NET0131  ;
	input \WX11107_reg/NET0131  ;
	input \WX11109_reg/NET0131  ;
	input \WX11111_reg/NET0131  ;
	input \WX11113_reg/NET0131  ;
	input \WX11115_reg/NET0131  ;
	input \WX11117_reg/NET0131  ;
	input \WX11119_reg/NET0131  ;
	input \WX11121_reg/NET0131  ;
	input \WX11123_reg/NET0131  ;
	input \WX11125_reg/NET0131  ;
	input \WX11127_reg/NET0131  ;
	input \WX11129_reg/NET0131  ;
	input \WX11131_reg/NET0131  ;
	input \WX11133_reg/NET0131  ;
	input \WX11135_reg/NET0131  ;
	input \WX11137_reg/NET0131  ;
	input \WX11139_reg/NET0131  ;
	input \WX11141_reg/NET0131  ;
	input \WX11143_reg/NET0131  ;
	input \WX11145_reg/NET0131  ;
	input \WX11147_reg/NET0131  ;
	input \WX11149_reg/NET0131  ;
	input \WX11151_reg/NET0131  ;
	input \WX11153_reg/NET0131  ;
	input \WX11155_reg/NET0131  ;
	input \WX11157_reg/NET0131  ;
	input \WX11159_reg/NET0131  ;
	input \WX11161_reg/NET0131  ;
	input \WX11163_reg/NET0131  ;
	input \WX11165_reg/NET0131  ;
	input \WX11167_reg/NET0131  ;
	input \WX11169_reg/NET0131  ;
	input \WX11171_reg/NET0131  ;
	input \WX11173_reg/NET0131  ;
	input \WX11175_reg/NET0131  ;
	input \WX11177_reg/NET0131  ;
	input \WX11179_reg/NET0131  ;
	input \WX11181_reg/NET0131  ;
	input \WX11183_reg/NET0131  ;
	input \WX11185_reg/NET0131  ;
	input \WX11187_reg/NET0131  ;
	input \WX11189_reg/NET0131  ;
	input \WX11191_reg/NET0131  ;
	input \WX11193_reg/NET0131  ;
	input \WX11195_reg/NET0131  ;
	input \WX11197_reg/NET0131  ;
	input \WX11199_reg/NET0131  ;
	input \WX11201_reg/NET0131  ;
	input \WX11203_reg/NET0131  ;
	input \WX11205_reg/NET0131  ;
	input \WX11207_reg/NET0131  ;
	input \WX11209_reg/NET0131  ;
	input \WX11211_reg/NET0131  ;
	input \WX11213_reg/NET0131  ;
	input \WX11215_reg/NET0131  ;
	input \WX11217_reg/NET0131  ;
	input \WX11219_reg/NET0131  ;
	input \WX11221_reg/NET0131  ;
	input \WX11223_reg/NET0131  ;
	input \WX11225_reg/NET0131  ;
	input \WX11227_reg/NET0131  ;
	input \WX11229_reg/NET0131  ;
	input \WX11231_reg/NET0131  ;
	input \WX11233_reg/NET0131  ;
	input \WX11235_reg/NET0131  ;
	input \WX11237_reg/NET0131  ;
	input \WX11239_reg/NET0131  ;
	input \WX11241_reg/NET0131  ;
	input \WX11243_reg/NET0131  ;
	input \WX1938_reg/NET0131  ;
	input \WX1940_reg/NET0131  ;
	input \WX1942_reg/NET0131  ;
	input \WX1944_reg/NET0131  ;
	input \WX1946_reg/NET0131  ;
	input \WX1948_reg/NET0131  ;
	input \WX1950_reg/NET0131  ;
	input \WX1952_reg/NET0131  ;
	input \WX1954_reg/NET0131  ;
	input \WX1956_reg/NET0131  ;
	input \WX1958_reg/NET0131  ;
	input \WX1960_reg/NET0131  ;
	input \WX1962_reg/NET0131  ;
	input \WX1964_reg/NET0131  ;
	input \WX1966_reg/NET0131  ;
	input \WX1968_reg/NET0131  ;
	input \WX1970_reg/NET0131  ;
	input \WX1972_reg/NET0131  ;
	input \WX1974_reg/NET0131  ;
	input \WX1976_reg/NET0131  ;
	input \WX1978_reg/NET0131  ;
	input \WX1980_reg/NET0131  ;
	input \WX1982_reg/NET0131  ;
	input \WX1984_reg/NET0131  ;
	input \WX1986_reg/NET0131  ;
	input \WX1988_reg/NET0131  ;
	input \WX1990_reg/NET0131  ;
	input \WX1992_reg/NET0131  ;
	input \WX1994_reg/NET0131  ;
	input \WX1996_reg/NET0131  ;
	input \WX1998_reg/NET0131  ;
	input \WX2000_reg/NET0131  ;
	input \WX2002_reg/NET0131  ;
	input \WX2004_reg/NET0131  ;
	input \WX2006_reg/NET0131  ;
	input \WX2008_reg/NET0131  ;
	input \WX2010_reg/NET0131  ;
	input \WX2012_reg/NET0131  ;
	input \WX2014_reg/NET0131  ;
	input \WX2016_reg/NET0131  ;
	input \WX2018_reg/NET0131  ;
	input \WX2020_reg/NET0131  ;
	input \WX2022_reg/NET0131  ;
	input \WX2024_reg/NET0131  ;
	input \WX2026_reg/NET0131  ;
	input \WX2028_reg/NET0131  ;
	input \WX2030_reg/NET0131  ;
	input \WX2032_reg/NET0131  ;
	input \WX2034_reg/NET0131  ;
	input \WX2036_reg/NET0131  ;
	input \WX2038_reg/NET0131  ;
	input \WX2040_reg/NET0131  ;
	input \WX2042_reg/NET0131  ;
	input \WX2044_reg/NET0131  ;
	input \WX2046_reg/NET0131  ;
	input \WX2048_reg/NET0131  ;
	input \WX2050_reg/NET0131  ;
	input \WX2052_reg/NET0131  ;
	input \WX2054_reg/NET0131  ;
	input \WX2056_reg/NET0131  ;
	input \WX2058_reg/NET0131  ;
	input \WX2060_reg/NET0131  ;
	input \WX2062_reg/NET0131  ;
	input \WX2064_reg/NET0131  ;
	input \WX2066_reg/NET0131  ;
	input \WX2068_reg/NET0131  ;
	input \WX2070_reg/NET0131  ;
	input \WX2072_reg/NET0131  ;
	input \WX2074_reg/NET0131  ;
	input \WX2076_reg/NET0131  ;
	input \WX2078_reg/NET0131  ;
	input \WX2080_reg/NET0131  ;
	input \WX2082_reg/NET0131  ;
	input \WX2084_reg/NET0131  ;
	input \WX2086_reg/NET0131  ;
	input \WX2088_reg/NET0131  ;
	input \WX2090_reg/NET0131  ;
	input \WX2092_reg/NET0131  ;
	input \WX2094_reg/NET0131  ;
	input \WX2096_reg/NET0131  ;
	input \WX2098_reg/NET0131  ;
	input \WX2100_reg/NET0131  ;
	input \WX2102_reg/NET0131  ;
	input \WX2104_reg/NET0131  ;
	input \WX2106_reg/NET0131  ;
	input \WX2108_reg/NET0131  ;
	input \WX2110_reg/NET0131  ;
	input \WX2112_reg/NET0131  ;
	input \WX2114_reg/NET0131  ;
	input \WX2116_reg/NET0131  ;
	input \WX2118_reg/NET0131  ;
	input \WX2120_reg/NET0131  ;
	input \WX2122_reg/NET0131  ;
	input \WX2124_reg/NET0131  ;
	input \WX2126_reg/NET0131  ;
	input \WX2128_reg/NET0131  ;
	input \WX2130_reg/NET0131  ;
	input \WX2132_reg/NET0131  ;
	input \WX2134_reg/NET0131  ;
	input \WX2136_reg/NET0131  ;
	input \WX2138_reg/NET0131  ;
	input \WX2140_reg/NET0131  ;
	input \WX2142_reg/NET0131  ;
	input \WX2144_reg/NET0131  ;
	input \WX2146_reg/NET0131  ;
	input \WX2148_reg/NET0131  ;
	input \WX2150_reg/NET0131  ;
	input \WX2152_reg/NET0131  ;
	input \WX2154_reg/NET0131  ;
	input \WX2156_reg/NET0131  ;
	input \WX2158_reg/NET0131  ;
	input \WX2160_reg/NET0131  ;
	input \WX2162_reg/NET0131  ;
	input \WX2164_reg/NET0131  ;
	input \WX2166_reg/NET0131  ;
	input \WX2168_reg/NET0131  ;
	input \WX2170_reg/NET0131  ;
	input \WX2172_reg/NET0131  ;
	input \WX2174_reg/NET0131  ;
	input \WX2176_reg/NET0131  ;
	input \WX2178_reg/NET0131  ;
	input \WX2180_reg/NET0131  ;
	input \WX2182_reg/NET0131  ;
	input \WX2184_reg/NET0131  ;
	input \WX2186_reg/NET0131  ;
	input \WX2188_reg/NET0131  ;
	input \WX2190_reg/NET0131  ;
	input \WX2192_reg/NET0131  ;
	input \WX3231_reg/NET0131  ;
	input \WX3233_reg/NET0131  ;
	input \WX3235_reg/NET0131  ;
	input \WX3237_reg/NET0131  ;
	input \WX3239_reg/NET0131  ;
	input \WX3241_reg/NET0131  ;
	input \WX3243_reg/NET0131  ;
	input \WX3245_reg/NET0131  ;
	input \WX3247_reg/NET0131  ;
	input \WX3249_reg/NET0131  ;
	input \WX3251_reg/NET0131  ;
	input \WX3253_reg/NET0131  ;
	input \WX3255_reg/NET0131  ;
	input \WX3257_reg/NET0131  ;
	input \WX3259_reg/NET0131  ;
	input \WX3261_reg/NET0131  ;
	input \WX3263_reg/NET0131  ;
	input \WX3265_reg/NET0131  ;
	input \WX3267_reg/NET0131  ;
	input \WX3269_reg/NET0131  ;
	input \WX3271_reg/NET0131  ;
	input \WX3273_reg/NET0131  ;
	input \WX3275_reg/NET0131  ;
	input \WX3277_reg/NET0131  ;
	input \WX3279_reg/NET0131  ;
	input \WX3281_reg/NET0131  ;
	input \WX3283_reg/NET0131  ;
	input \WX3285_reg/NET0131  ;
	input \WX3287_reg/NET0131  ;
	input \WX3289_reg/NET0131  ;
	input \WX3291_reg/NET0131  ;
	input \WX3293_reg/NET0131  ;
	input \WX3295_reg/NET0131  ;
	input \WX3297_reg/NET0131  ;
	input \WX3299_reg/NET0131  ;
	input \WX3301_reg/NET0131  ;
	input \WX3303_reg/NET0131  ;
	input \WX3305_reg/NET0131  ;
	input \WX3307_reg/NET0131  ;
	input \WX3309_reg/NET0131  ;
	input \WX3311_reg/NET0131  ;
	input \WX3313_reg/NET0131  ;
	input \WX3315_reg/NET0131  ;
	input \WX3317_reg/NET0131  ;
	input \WX3319_reg/NET0131  ;
	input \WX3321_reg/NET0131  ;
	input \WX3323_reg/NET0131  ;
	input \WX3325_reg/NET0131  ;
	input \WX3327_reg/NET0131  ;
	input \WX3329_reg/NET0131  ;
	input \WX3331_reg/NET0131  ;
	input \WX3333_reg/NET0131  ;
	input \WX3335_reg/NET0131  ;
	input \WX3337_reg/NET0131  ;
	input \WX3339_reg/NET0131  ;
	input \WX3341_reg/NET0131  ;
	input \WX3343_reg/NET0131  ;
	input \WX3345_reg/NET0131  ;
	input \WX3347_reg/NET0131  ;
	input \WX3349_reg/NET0131  ;
	input \WX3351_reg/NET0131  ;
	input \WX3353_reg/NET0131  ;
	input \WX3355_reg/NET0131  ;
	input \WX3357_reg/NET0131  ;
	input \WX3359_reg/NET0131  ;
	input \WX3361_reg/NET0131  ;
	input \WX3363_reg/NET0131  ;
	input \WX3365_reg/NET0131  ;
	input \WX3367_reg/NET0131  ;
	input \WX3369_reg/NET0131  ;
	input \WX3371_reg/NET0131  ;
	input \WX3373_reg/NET0131  ;
	input \WX3375_reg/NET0131  ;
	input \WX3377_reg/NET0131  ;
	input \WX3379_reg/NET0131  ;
	input \WX3381_reg/NET0131  ;
	input \WX3383_reg/NET0131  ;
	input \WX3385_reg/NET0131  ;
	input \WX3387_reg/NET0131  ;
	input \WX3389_reg/NET0131  ;
	input \WX3391_reg/NET0131  ;
	input \WX3393_reg/NET0131  ;
	input \WX3395_reg/NET0131  ;
	input \WX3397_reg/NET0131  ;
	input \WX3399_reg/NET0131  ;
	input \WX3401_reg/NET0131  ;
	input \WX3403_reg/NET0131  ;
	input \WX3405_reg/NET0131  ;
	input \WX3407_reg/NET0131  ;
	input \WX3409_reg/NET0131  ;
	input \WX3411_reg/NET0131  ;
	input \WX3413_reg/NET0131  ;
	input \WX3415_reg/NET0131  ;
	input \WX3417_reg/NET0131  ;
	input \WX3419_reg/NET0131  ;
	input \WX3421_reg/NET0131  ;
	input \WX3423_reg/NET0131  ;
	input \WX3425_reg/NET0131  ;
	input \WX3427_reg/NET0131  ;
	input \WX3429_reg/NET0131  ;
	input \WX3431_reg/NET0131  ;
	input \WX3433_reg/NET0131  ;
	input \WX3435_reg/NET0131  ;
	input \WX3437_reg/NET0131  ;
	input \WX3439_reg/NET0131  ;
	input \WX3441_reg/NET0131  ;
	input \WX3443_reg/NET0131  ;
	input \WX3445_reg/NET0131  ;
	input \WX3447_reg/NET0131  ;
	input \WX3449_reg/NET0131  ;
	input \WX3451_reg/NET0131  ;
	input \WX3453_reg/NET0131  ;
	input \WX3455_reg/NET0131  ;
	input \WX3457_reg/NET0131  ;
	input \WX3459_reg/NET0131  ;
	input \WX3461_reg/NET0131  ;
	input \WX3463_reg/NET0131  ;
	input \WX3465_reg/NET0131  ;
	input \WX3467_reg/NET0131  ;
	input \WX3469_reg/NET0131  ;
	input \WX3471_reg/NET0131  ;
	input \WX3473_reg/NET0131  ;
	input \WX3475_reg/NET0131  ;
	input \WX3477_reg/NET0131  ;
	input \WX3479_reg/NET0131  ;
	input \WX3481_reg/NET0131  ;
	input \WX3483_reg/NET0131  ;
	input \WX3485_reg/NET0131  ;
	input \WX4524_reg/NET0131  ;
	input \WX4526_reg/NET0131  ;
	input \WX4528_reg/NET0131  ;
	input \WX4530_reg/NET0131  ;
	input \WX4532_reg/NET0131  ;
	input \WX4534_reg/NET0131  ;
	input \WX4536_reg/NET0131  ;
	input \WX4538_reg/NET0131  ;
	input \WX4540_reg/NET0131  ;
	input \WX4542_reg/NET0131  ;
	input \WX4544_reg/NET0131  ;
	input \WX4546_reg/NET0131  ;
	input \WX4548_reg/NET0131  ;
	input \WX4550_reg/NET0131  ;
	input \WX4552_reg/NET0131  ;
	input \WX4554_reg/NET0131  ;
	input \WX4556_reg/NET0131  ;
	input \WX4558_reg/NET0131  ;
	input \WX4560_reg/NET0131  ;
	input \WX4562_reg/NET0131  ;
	input \WX4564_reg/NET0131  ;
	input \WX4566_reg/NET0131  ;
	input \WX4568_reg/NET0131  ;
	input \WX4570_reg/NET0131  ;
	input \WX4572_reg/NET0131  ;
	input \WX4574_reg/NET0131  ;
	input \WX4576_reg/NET0131  ;
	input \WX4578_reg/NET0131  ;
	input \WX4580_reg/NET0131  ;
	input \WX4582_reg/NET0131  ;
	input \WX4584_reg/NET0131  ;
	input \WX4586_reg/NET0131  ;
	input \WX4588_reg/NET0131  ;
	input \WX4590_reg/NET0131  ;
	input \WX4592_reg/NET0131  ;
	input \WX4594_reg/NET0131  ;
	input \WX4596_reg/NET0131  ;
	input \WX4598_reg/NET0131  ;
	input \WX4600_reg/NET0131  ;
	input \WX4602_reg/NET0131  ;
	input \WX4604_reg/NET0131  ;
	input \WX4606_reg/NET0131  ;
	input \WX4608_reg/NET0131  ;
	input \WX4610_reg/NET0131  ;
	input \WX4612_reg/NET0131  ;
	input \WX4614_reg/NET0131  ;
	input \WX4616_reg/NET0131  ;
	input \WX4618_reg/NET0131  ;
	input \WX4620_reg/NET0131  ;
	input \WX4622_reg/NET0131  ;
	input \WX4624_reg/NET0131  ;
	input \WX4626_reg/NET0131  ;
	input \WX4628_reg/NET0131  ;
	input \WX4630_reg/NET0131  ;
	input \WX4632_reg/NET0131  ;
	input \WX4634_reg/NET0131  ;
	input \WX4636_reg/NET0131  ;
	input \WX4638_reg/NET0131  ;
	input \WX4640_reg/NET0131  ;
	input \WX4642_reg/NET0131  ;
	input \WX4644_reg/NET0131  ;
	input \WX4646_reg/NET0131  ;
	input \WX4648_reg/NET0131  ;
	input \WX4650_reg/NET0131  ;
	input \WX4652_reg/NET0131  ;
	input \WX4654_reg/NET0131  ;
	input \WX4656_reg/NET0131  ;
	input \WX4658_reg/NET0131  ;
	input \WX4660_reg/NET0131  ;
	input \WX4662_reg/NET0131  ;
	input \WX4664_reg/NET0131  ;
	input \WX4666_reg/NET0131  ;
	input \WX4668_reg/NET0131  ;
	input \WX4670_reg/NET0131  ;
	input \WX4672_reg/NET0131  ;
	input \WX4674_reg/NET0131  ;
	input \WX4676_reg/NET0131  ;
	input \WX4678_reg/NET0131  ;
	input \WX4680_reg/NET0131  ;
	input \WX4682_reg/NET0131  ;
	input \WX4684_reg/NET0131  ;
	input \WX4686_reg/NET0131  ;
	input \WX4688_reg/NET0131  ;
	input \WX4690_reg/NET0131  ;
	input \WX4692_reg/NET0131  ;
	input \WX4694_reg/NET0131  ;
	input \WX4696_reg/NET0131  ;
	input \WX4698_reg/NET0131  ;
	input \WX4700_reg/NET0131  ;
	input \WX4702_reg/NET0131  ;
	input \WX4704_reg/NET0131  ;
	input \WX4706_reg/NET0131  ;
	input \WX4708_reg/NET0131  ;
	input \WX4710_reg/NET0131  ;
	input \WX4712_reg/NET0131  ;
	input \WX4714_reg/NET0131  ;
	input \WX4716_reg/NET0131  ;
	input \WX4718_reg/NET0131  ;
	input \WX4720_reg/NET0131  ;
	input \WX4722_reg/NET0131  ;
	input \WX4724_reg/NET0131  ;
	input \WX4726_reg/NET0131  ;
	input \WX4728_reg/NET0131  ;
	input \WX4730_reg/NET0131  ;
	input \WX4732_reg/NET0131  ;
	input \WX4734_reg/NET0131  ;
	input \WX4736_reg/NET0131  ;
	input \WX4738_reg/NET0131  ;
	input \WX4740_reg/NET0131  ;
	input \WX4742_reg/NET0131  ;
	input \WX4744_reg/NET0131  ;
	input \WX4746_reg/NET0131  ;
	input \WX4748_reg/NET0131  ;
	input \WX4750_reg/NET0131  ;
	input \WX4752_reg/NET0131  ;
	input \WX4754_reg/NET0131  ;
	input \WX4756_reg/NET0131  ;
	input \WX4758_reg/NET0131  ;
	input \WX4760_reg/NET0131  ;
	input \WX4762_reg/NET0131  ;
	input \WX4764_reg/NET0131  ;
	input \WX4766_reg/NET0131  ;
	input \WX4768_reg/NET0131  ;
	input \WX4770_reg/NET0131  ;
	input \WX4772_reg/NET0131  ;
	input \WX4774_reg/NET0131  ;
	input \WX4776_reg/NET0131  ;
	input \WX4778_reg/NET0131  ;
	input \WX5817_reg/NET0131  ;
	input \WX5819_reg/NET0131  ;
	input \WX5821_reg/NET0131  ;
	input \WX5823_reg/NET0131  ;
	input \WX5825_reg/NET0131  ;
	input \WX5827_reg/NET0131  ;
	input \WX5829_reg/NET0131  ;
	input \WX5831_reg/NET0131  ;
	input \WX5833_reg/NET0131  ;
	input \WX5835_reg/NET0131  ;
	input \WX5837_reg/NET0131  ;
	input \WX5839_reg/NET0131  ;
	input \WX5841_reg/NET0131  ;
	input \WX5843_reg/NET0131  ;
	input \WX5845_reg/NET0131  ;
	input \WX5847_reg/NET0131  ;
	input \WX5849_reg/NET0131  ;
	input \WX5851_reg/NET0131  ;
	input \WX5853_reg/NET0131  ;
	input \WX5855_reg/NET0131  ;
	input \WX5857_reg/NET0131  ;
	input \WX5859_reg/NET0131  ;
	input \WX5861_reg/NET0131  ;
	input \WX5863_reg/NET0131  ;
	input \WX5865_reg/NET0131  ;
	input \WX5867_reg/NET0131  ;
	input \WX5869_reg/NET0131  ;
	input \WX5871_reg/NET0131  ;
	input \WX5873_reg/NET0131  ;
	input \WX5875_reg/NET0131  ;
	input \WX5877_reg/NET0131  ;
	input \WX5879_reg/NET0131  ;
	input \WX5881_reg/NET0131  ;
	input \WX5883_reg/NET0131  ;
	input \WX5885_reg/NET0131  ;
	input \WX5887_reg/NET0131  ;
	input \WX5889_reg/NET0131  ;
	input \WX5891_reg/NET0131  ;
	input \WX5893_reg/NET0131  ;
	input \WX5895_reg/NET0131  ;
	input \WX5897_reg/NET0131  ;
	input \WX5899_reg/NET0131  ;
	input \WX5901_reg/NET0131  ;
	input \WX5903_reg/NET0131  ;
	input \WX5905_reg/NET0131  ;
	input \WX5907_reg/NET0131  ;
	input \WX5909_reg/NET0131  ;
	input \WX5911_reg/NET0131  ;
	input \WX5913_reg/NET0131  ;
	input \WX5915_reg/NET0131  ;
	input \WX5917_reg/NET0131  ;
	input \WX5919_reg/NET0131  ;
	input \WX5921_reg/NET0131  ;
	input \WX5923_reg/NET0131  ;
	input \WX5925_reg/NET0131  ;
	input \WX5927_reg/NET0131  ;
	input \WX5929_reg/NET0131  ;
	input \WX5931_reg/NET0131  ;
	input \WX5933_reg/NET0131  ;
	input \WX5935_reg/NET0131  ;
	input \WX5937_reg/NET0131  ;
	input \WX5939_reg/NET0131  ;
	input \WX5941_reg/NET0131  ;
	input \WX5943_reg/NET0131  ;
	input \WX5945_reg/NET0131  ;
	input \WX5947_reg/NET0131  ;
	input \WX5949_reg/NET0131  ;
	input \WX5951_reg/NET0131  ;
	input \WX5953_reg/NET0131  ;
	input \WX5955_reg/NET0131  ;
	input \WX5957_reg/NET0131  ;
	input \WX5959_reg/NET0131  ;
	input \WX5961_reg/NET0131  ;
	input \WX5963_reg/NET0131  ;
	input \WX5965_reg/NET0131  ;
	input \WX5967_reg/NET0131  ;
	input \WX5969_reg/NET0131  ;
	input \WX5971_reg/NET0131  ;
	input \WX5973_reg/NET0131  ;
	input \WX5975_reg/NET0131  ;
	input \WX5977_reg/NET0131  ;
	input \WX5979_reg/NET0131  ;
	input \WX5981_reg/NET0131  ;
	input \WX5983_reg/NET0131  ;
	input \WX5985_reg/NET0131  ;
	input \WX5987_reg/NET0131  ;
	input \WX5989_reg/NET0131  ;
	input \WX5991_reg/NET0131  ;
	input \WX5993_reg/NET0131  ;
	input \WX5995_reg/NET0131  ;
	input \WX5997_reg/NET0131  ;
	input \WX5999_reg/NET0131  ;
	input \WX6001_reg/NET0131  ;
	input \WX6003_reg/NET0131  ;
	input \WX6005_reg/NET0131  ;
	input \WX6007_reg/NET0131  ;
	input \WX6009_reg/NET0131  ;
	input \WX6011_reg/NET0131  ;
	input \WX6013_reg/NET0131  ;
	input \WX6015_reg/NET0131  ;
	input \WX6017_reg/NET0131  ;
	input \WX6019_reg/NET0131  ;
	input \WX6021_reg/NET0131  ;
	input \WX6023_reg/NET0131  ;
	input \WX6025_reg/NET0131  ;
	input \WX6027_reg/NET0131  ;
	input \WX6029_reg/NET0131  ;
	input \WX6031_reg/NET0131  ;
	input \WX6033_reg/NET0131  ;
	input \WX6035_reg/NET0131  ;
	input \WX6037_reg/NET0131  ;
	input \WX6039_reg/NET0131  ;
	input \WX6041_reg/NET0131  ;
	input \WX6043_reg/NET0131  ;
	input \WX6045_reg/NET0131  ;
	input \WX6047_reg/NET0131  ;
	input \WX6049_reg/NET0131  ;
	input \WX6051_reg/NET0131  ;
	input \WX6053_reg/NET0131  ;
	input \WX6055_reg/NET0131  ;
	input \WX6057_reg/NET0131  ;
	input \WX6059_reg/NET0131  ;
	input \WX6061_reg/NET0131  ;
	input \WX6063_reg/NET0131  ;
	input \WX6065_reg/NET0131  ;
	input \WX6067_reg/NET0131  ;
	input \WX6069_reg/NET0131  ;
	input \WX6071_reg/NET0131  ;
	input \WX645_reg/NET0131  ;
	input \WX647_reg/NET0131  ;
	input \WX649_reg/NET0131  ;
	input \WX651_reg/NET0131  ;
	input \WX653_reg/NET0131  ;
	input \WX655_reg/NET0131  ;
	input \WX657_reg/NET0131  ;
	input \WX659_reg/NET0131  ;
	input \WX661_reg/NET0131  ;
	input \WX663_reg/NET0131  ;
	input \WX665_reg/NET0131  ;
	input \WX667_reg/NET0131  ;
	input \WX669_reg/NET0131  ;
	input \WX671_reg/NET0131  ;
	input \WX673_reg/NET0131  ;
	input \WX675_reg/NET0131  ;
	input \WX677_reg/NET0131  ;
	input \WX679_reg/NET0131  ;
	input \WX681_reg/NET0131  ;
	input \WX683_reg/NET0131  ;
	input \WX685_reg/NET0131  ;
	input \WX687_reg/NET0131  ;
	input \WX689_reg/NET0131  ;
	input \WX691_reg/NET0131  ;
	input \WX693_reg/NET0131  ;
	input \WX695_reg/NET0131  ;
	input \WX697_reg/NET0131  ;
	input \WX699_reg/NET0131  ;
	input \WX701_reg/NET0131  ;
	input \WX703_reg/NET0131  ;
	input \WX705_reg/NET0131  ;
	input \WX707_reg/NET0131  ;
	input \WX709_reg/NET0131  ;
	input \WX7110_reg/NET0131  ;
	input \WX7112_reg/NET0131  ;
	input \WX7114_reg/NET0131  ;
	input \WX7116_reg/NET0131  ;
	input \WX7118_reg/NET0131  ;
	input \WX711_reg/NET0131  ;
	input \WX7120_reg/NET0131  ;
	input \WX7122_reg/NET0131  ;
	input \WX7124_reg/NET0131  ;
	input \WX7126_reg/NET0131  ;
	input \WX7128_reg/NET0131  ;
	input \WX7130_reg/NET0131  ;
	input \WX7132_reg/NET0131  ;
	input \WX7134_reg/NET0131  ;
	input \WX7136_reg/NET0131  ;
	input \WX7138_reg/NET0131  ;
	input \WX713_reg/NET0131  ;
	input \WX7140_reg/NET0131  ;
	input \WX7142_reg/NET0131  ;
	input \WX7144_reg/NET0131  ;
	input \WX7146_reg/NET0131  ;
	input \WX7148_reg/NET0131  ;
	input \WX7150_reg/NET0131  ;
	input \WX7152_reg/NET0131  ;
	input \WX7154_reg/NET0131  ;
	input \WX7156_reg/NET0131  ;
	input \WX7158_reg/NET0131  ;
	input \WX715_reg/NET0131  ;
	input \WX7160_reg/NET0131  ;
	input \WX7162_reg/NET0131  ;
	input \WX7164_reg/NET0131  ;
	input \WX7166_reg/NET0131  ;
	input \WX7168_reg/NET0131  ;
	input \WX7170_reg/NET0131  ;
	input \WX7172_reg/NET0131  ;
	input \WX7174_reg/NET0131  ;
	input \WX7176_reg/NET0131  ;
	input \WX7178_reg/NET0131  ;
	input \WX717_reg/NET0131  ;
	input \WX7180_reg/NET0131  ;
	input \WX7182_reg/NET0131  ;
	input \WX7184_reg/NET0131  ;
	input \WX7186_reg/NET0131  ;
	input \WX7188_reg/NET0131  ;
	input \WX7190_reg/NET0131  ;
	input \WX7192_reg/NET0131  ;
	input \WX7194_reg/NET0131  ;
	input \WX7196_reg/NET0131  ;
	input \WX7198_reg/NET0131  ;
	input \WX719_reg/NET0131  ;
	input \WX7200_reg/NET0131  ;
	input \WX7202_reg/NET0131  ;
	input \WX7204_reg/NET0131  ;
	input \WX7206_reg/NET0131  ;
	input \WX7208_reg/NET0131  ;
	input \WX7210_reg/NET0131  ;
	input \WX7212_reg/NET0131  ;
	input \WX7214_reg/NET0131  ;
	input \WX7216_reg/NET0131  ;
	input \WX7218_reg/NET0131  ;
	input \WX721_reg/NET0131  ;
	input \WX7220_reg/NET0131  ;
	input \WX7222_reg/NET0131  ;
	input \WX7224_reg/NET0131  ;
	input \WX7226_reg/NET0131  ;
	input \WX7228_reg/NET0131  ;
	input \WX7230_reg/NET0131  ;
	input \WX7232_reg/NET0131  ;
	input \WX7234_reg/NET0131  ;
	input \WX7236_reg/NET0131  ;
	input \WX7238_reg/NET0131  ;
	input \WX723_reg/NET0131  ;
	input \WX7240_reg/NET0131  ;
	input \WX7242_reg/NET0131  ;
	input \WX7244_reg/NET0131  ;
	input \WX7246_reg/NET0131  ;
	input \WX7248_reg/NET0131  ;
	input \WX7250_reg/NET0131  ;
	input \WX7252_reg/NET0131  ;
	input \WX7254_reg/NET0131  ;
	input \WX7256_reg/NET0131  ;
	input \WX7258_reg/NET0131  ;
	input \WX725_reg/NET0131  ;
	input \WX7260_reg/NET0131  ;
	input \WX7262_reg/NET0131  ;
	input \WX7264_reg/NET0131  ;
	input \WX7266_reg/NET0131  ;
	input \WX7268_reg/NET0131  ;
	input \WX7270_reg/NET0131  ;
	input \WX7272_reg/NET0131  ;
	input \WX7274_reg/NET0131  ;
	input \WX7276_reg/NET0131  ;
	input \WX7278_reg/NET0131  ;
	input \WX727_reg/NET0131  ;
	input \WX7280_reg/NET0131  ;
	input \WX7282_reg/NET0131  ;
	input \WX7284_reg/NET0131  ;
	input \WX7286_reg/NET0131  ;
	input \WX7288_reg/NET0131  ;
	input \WX7290_reg/NET0131  ;
	input \WX7292_reg/NET0131  ;
	input \WX7294_reg/NET0131  ;
	input \WX7296_reg/NET0131  ;
	input \WX7298_reg/NET0131  ;
	input \WX729_reg/NET0131  ;
	input \WX7300_reg/NET0131  ;
	input \WX7302_reg/NET0131  ;
	input \WX7304_reg/NET0131  ;
	input \WX7306_reg/NET0131  ;
	input \WX7308_reg/NET0131  ;
	input \WX7310_reg/NET0131  ;
	input \WX7312_reg/NET0131  ;
	input \WX7314_reg/NET0131  ;
	input \WX7316_reg/NET0131  ;
	input \WX7318_reg/NET0131  ;
	input \WX731_reg/NET0131  ;
	input \WX7320_reg/NET0131  ;
	input \WX7322_reg/NET0131  ;
	input \WX7324_reg/NET0131  ;
	input \WX7326_reg/NET0131  ;
	input \WX7328_reg/NET0131  ;
	input \WX7330_reg/NET0131  ;
	input \WX7332_reg/NET0131  ;
	input \WX7334_reg/NET0131  ;
	input \WX7336_reg/NET0131  ;
	input \WX7338_reg/NET0131  ;
	input \WX733_reg/NET0131  ;
	input \WX7340_reg/NET0131  ;
	input \WX7342_reg/NET0131  ;
	input \WX7344_reg/NET0131  ;
	input \WX7346_reg/NET0131  ;
	input \WX7348_reg/NET0131  ;
	input \WX7350_reg/NET0131  ;
	input \WX7352_reg/NET0131  ;
	input \WX7354_reg/NET0131  ;
	input \WX7356_reg/NET0131  ;
	input \WX7358_reg/NET0131  ;
	input \WX735_reg/NET0131  ;
	input \WX7360_reg/NET0131  ;
	input \WX7362_reg/NET0131  ;
	input \WX7364_reg/NET0131  ;
	input \WX737_reg/NET0131  ;
	input \WX739_reg/NET0131  ;
	input \WX741_reg/NET0131  ;
	input \WX743_reg/NET0131  ;
	input \WX745_reg/NET0131  ;
	input \WX747_reg/NET0131  ;
	input \WX749_reg/NET0131  ;
	input \WX751_reg/NET0131  ;
	input \WX753_reg/NET0131  ;
	input \WX755_reg/NET0131  ;
	input \WX757_reg/NET0131  ;
	input \WX759_reg/NET0131  ;
	input \WX761_reg/NET0131  ;
	input \WX763_reg/NET0131  ;
	input \WX765_reg/NET0131  ;
	input \WX767_reg/NET0131  ;
	input \WX769_reg/NET0131  ;
	input \WX771_reg/NET0131  ;
	input \WX773_reg/NET0131  ;
	input \WX775_reg/NET0131  ;
	input \WX777_reg/NET0131  ;
	input \WX779_reg/NET0131  ;
	input \WX781_reg/NET0131  ;
	input \WX783_reg/NET0131  ;
	input \WX785_reg/NET0131  ;
	input \WX787_reg/NET0131  ;
	input \WX789_reg/NET0131  ;
	input \WX791_reg/NET0131  ;
	input \WX793_reg/NET0131  ;
	input \WX795_reg/NET0131  ;
	input \WX797_reg/NET0131  ;
	input \WX799_reg/NET0131  ;
	input \WX801_reg/NET0131  ;
	input \WX803_reg/NET0131  ;
	input \WX805_reg/NET0131  ;
	input \WX807_reg/NET0131  ;
	input \WX809_reg/NET0131  ;
	input \WX811_reg/NET0131  ;
	input \WX813_reg/NET0131  ;
	input \WX815_reg/NET0131  ;
	input \WX817_reg/NET0131  ;
	input \WX819_reg/NET0131  ;
	input \WX821_reg/NET0131  ;
	input \WX823_reg/NET0131  ;
	input \WX825_reg/NET0131  ;
	input \WX827_reg/NET0131  ;
	input \WX829_reg/NET0131  ;
	input \WX831_reg/NET0131  ;
	input \WX833_reg/NET0131  ;
	input \WX835_reg/NET0131  ;
	input \WX837_reg/NET0131  ;
	input \WX839_reg/NET0131  ;
	input \WX8403_reg/NET0131  ;
	input \WX8405_reg/NET0131  ;
	input \WX8407_reg/NET0131  ;
	input \WX8409_reg/NET0131  ;
	input \WX8411_reg/NET0131  ;
	input \WX8413_reg/NET0131  ;
	input \WX8415_reg/NET0131  ;
	input \WX8417_reg/NET0131  ;
	input \WX8419_reg/NET0131  ;
	input \WX841_reg/NET0131  ;
	input \WX8421_reg/NET0131  ;
	input \WX8423_reg/NET0131  ;
	input \WX8425_reg/NET0131  ;
	input \WX8427_reg/NET0131  ;
	input \WX8429_reg/NET0131  ;
	input \WX8431_reg/NET0131  ;
	input \WX8433_reg/NET0131  ;
	input \WX8435_reg/NET0131  ;
	input \WX8437_reg/NET0131  ;
	input \WX8439_reg/NET0131  ;
	input \WX843_reg/NET0131  ;
	input \WX8441_reg/NET0131  ;
	input \WX8443_reg/NET0131  ;
	input \WX8445_reg/NET0131  ;
	input \WX8447_reg/NET0131  ;
	input \WX8449_reg/NET0131  ;
	input \WX8451_reg/NET0131  ;
	input \WX8453_reg/NET0131  ;
	input \WX8455_reg/NET0131  ;
	input \WX8457_reg/NET0131  ;
	input \WX8459_reg/NET0131  ;
	input \WX845_reg/NET0131  ;
	input \WX8461_reg/NET0131  ;
	input \WX8463_reg/NET0131  ;
	input \WX8465_reg/NET0131  ;
	input \WX8467_reg/NET0131  ;
	input \WX8469_reg/NET0131  ;
	input \WX8471_reg/NET0131  ;
	input \WX8473_reg/NET0131  ;
	input \WX8475_reg/NET0131  ;
	input \WX8477_reg/NET0131  ;
	input \WX8479_reg/NET0131  ;
	input \WX847_reg/NET0131  ;
	input \WX8481_reg/NET0131  ;
	input \WX8483_reg/NET0131  ;
	input \WX8485_reg/NET0131  ;
	input \WX8487_reg/NET0131  ;
	input \WX8489_reg/NET0131  ;
	input \WX8491_reg/NET0131  ;
	input \WX8493_reg/NET0131  ;
	input \WX8495_reg/NET0131  ;
	input \WX8497_reg/NET0131  ;
	input \WX8499_reg/NET0131  ;
	input \WX849_reg/NET0131  ;
	input \WX8501_reg/NET0131  ;
	input \WX8503_reg/NET0131  ;
	input \WX8505_reg/NET0131  ;
	input \WX8507_reg/NET0131  ;
	input \WX8509_reg/NET0131  ;
	input \WX8511_reg/NET0131  ;
	input \WX8513_reg/NET0131  ;
	input \WX8515_reg/NET0131  ;
	input \WX8517_reg/NET0131  ;
	input \WX8519_reg/NET0131  ;
	input \WX851_reg/NET0131  ;
	input \WX8521_reg/NET0131  ;
	input \WX8523_reg/NET0131  ;
	input \WX8525_reg/NET0131  ;
	input \WX8527_reg/NET0131  ;
	input \WX8529_reg/NET0131  ;
	input \WX8531_reg/NET0131  ;
	input \WX8533_reg/NET0131  ;
	input \WX8535_reg/NET0131  ;
	input \WX8537_reg/NET0131  ;
	input \WX8539_reg/NET0131  ;
	input \WX853_reg/NET0131  ;
	input \WX8541_reg/NET0131  ;
	input \WX8543_reg/NET0131  ;
	input \WX8545_reg/NET0131  ;
	input \WX8547_reg/NET0131  ;
	input \WX8549_reg/NET0131  ;
	input \WX8551_reg/NET0131  ;
	input \WX8553_reg/NET0131  ;
	input \WX8555_reg/NET0131  ;
	input \WX8557_reg/NET0131  ;
	input \WX8559_reg/NET0131  ;
	input \WX855_reg/NET0131  ;
	input \WX8561_reg/NET0131  ;
	input \WX8563_reg/NET0131  ;
	input \WX8565_reg/NET0131  ;
	input \WX8567_reg/NET0131  ;
	input \WX8569_reg/NET0131  ;
	input \WX8571_reg/NET0131  ;
	input \WX8573_reg/NET0131  ;
	input \WX8575_reg/NET0131  ;
	input \WX8577_reg/NET0131  ;
	input \WX8579_reg/NET0131  ;
	input \WX857_reg/NET0131  ;
	input \WX8581_reg/NET0131  ;
	input \WX8583_reg/NET0131  ;
	input \WX8585_reg/NET0131  ;
	input \WX8587_reg/NET0131  ;
	input \WX8589_reg/NET0131  ;
	input \WX8591_reg/NET0131  ;
	input \WX8593_reg/NET0131  ;
	input \WX8595_reg/NET0131  ;
	input \WX8597_reg/NET0131  ;
	input \WX8599_reg/NET0131  ;
	input \WX859_reg/NET0131  ;
	input \WX8601_reg/NET0131  ;
	input \WX8603_reg/NET0131  ;
	input \WX8605_reg/NET0131  ;
	input \WX8607_reg/NET0131  ;
	input \WX8609_reg/NET0131  ;
	input \WX8611_reg/NET0131  ;
	input \WX8613_reg/NET0131  ;
	input \WX8615_reg/NET0131  ;
	input \WX8617_reg/NET0131  ;
	input \WX8619_reg/NET0131  ;
	input \WX861_reg/NET0131  ;
	input \WX8621_reg/NET0131  ;
	input \WX8623_reg/NET0131  ;
	input \WX8625_reg/NET0131  ;
	input \WX8627_reg/NET0131  ;
	input \WX8629_reg/NET0131  ;
	input \WX8631_reg/NET0131  ;
	input \WX8633_reg/NET0131  ;
	input \WX8635_reg/NET0131  ;
	input \WX8637_reg/NET0131  ;
	input \WX8639_reg/NET0131  ;
	input \WX863_reg/NET0131  ;
	input \WX8641_reg/NET0131  ;
	input \WX8643_reg/NET0131  ;
	input \WX8645_reg/NET0131  ;
	input \WX8647_reg/NET0131  ;
	input \WX8649_reg/NET0131  ;
	input \WX8651_reg/NET0131  ;
	input \WX8653_reg/NET0131  ;
	input \WX8655_reg/NET0131  ;
	input \WX8657_reg/NET0131  ;
	input \WX865_reg/NET0131  ;
	input \WX867_reg/NET0131  ;
	input \WX869_reg/NET0131  ;
	input \WX871_reg/NET0131  ;
	input \WX873_reg/NET0131  ;
	input \WX875_reg/NET0131  ;
	input \WX877_reg/NET0131  ;
	input \WX879_reg/NET0131  ;
	input \WX881_reg/NET0131  ;
	input \WX883_reg/NET0131  ;
	input \WX885_reg/NET0131  ;
	input \WX887_reg/NET0131  ;
	input \WX889_reg/NET0131  ;
	input \WX891_reg/NET0131  ;
	input \WX893_reg/NET0131  ;
	input \WX895_reg/NET0131  ;
	input \WX897_reg/NET0131  ;
	input \WX899_reg/NET0131  ;
	input \WX9696_reg/NET0131  ;
	input \WX9698_reg/NET0131  ;
	input \WX9700_reg/NET0131  ;
	input \WX9702_reg/NET0131  ;
	input \WX9704_reg/NET0131  ;
	input \WX9706_reg/NET0131  ;
	input \WX9708_reg/NET0131  ;
	input \WX9710_reg/NET0131  ;
	input \WX9712_reg/NET0131  ;
	input \WX9714_reg/NET0131  ;
	input \WX9716_reg/NET0131  ;
	input \WX9718_reg/NET0131  ;
	input \WX9720_reg/NET0131  ;
	input \WX9722_reg/NET0131  ;
	input \WX9724_reg/NET0131  ;
	input \WX9726_reg/NET0131  ;
	input \WX9728_reg/NET0131  ;
	input \WX9730_reg/NET0131  ;
	input \WX9732_reg/NET0131  ;
	input \WX9734_reg/NET0131  ;
	input \WX9736_reg/NET0131  ;
	input \WX9738_reg/NET0131  ;
	input \WX9740_reg/NET0131  ;
	input \WX9742_reg/NET0131  ;
	input \WX9744_reg/NET0131  ;
	input \WX9746_reg/NET0131  ;
	input \WX9748_reg/NET0131  ;
	input \WX9750_reg/NET0131  ;
	input \WX9752_reg/NET0131  ;
	input \WX9754_reg/NET0131  ;
	input \WX9756_reg/NET0131  ;
	input \WX9758_reg/NET0131  ;
	input \WX9760_reg/NET0131  ;
	input \WX9762_reg/NET0131  ;
	input \WX9764_reg/NET0131  ;
	input \WX9766_reg/NET0131  ;
	input \WX9768_reg/NET0131  ;
	input \WX9770_reg/NET0131  ;
	input \WX9772_reg/NET0131  ;
	input \WX9774_reg/NET0131  ;
	input \WX9776_reg/NET0131  ;
	input \WX9778_reg/NET0131  ;
	input \WX9780_reg/NET0131  ;
	input \WX9782_reg/NET0131  ;
	input \WX9784_reg/NET0131  ;
	input \WX9786_reg/NET0131  ;
	input \WX9788_reg/NET0131  ;
	input \WX9790_reg/NET0131  ;
	input \WX9792_reg/NET0131  ;
	input \WX9794_reg/NET0131  ;
	input \WX9796_reg/NET0131  ;
	input \WX9798_reg/NET0131  ;
	input \WX9800_reg/NET0131  ;
	input \WX9802_reg/NET0131  ;
	input \WX9804_reg/NET0131  ;
	input \WX9806_reg/NET0131  ;
	input \WX9808_reg/NET0131  ;
	input \WX9810_reg/NET0131  ;
	input \WX9812_reg/NET0131  ;
	input \WX9814_reg/NET0131  ;
	input \WX9816_reg/NET0131  ;
	input \WX9818_reg/NET0131  ;
	input \WX9820_reg/NET0131  ;
	input \WX9822_reg/NET0131  ;
	input \WX9824_reg/NET0131  ;
	input \WX9826_reg/NET0131  ;
	input \WX9828_reg/NET0131  ;
	input \WX9830_reg/NET0131  ;
	input \WX9832_reg/NET0131  ;
	input \WX9834_reg/NET0131  ;
	input \WX9836_reg/NET0131  ;
	input \WX9838_reg/NET0131  ;
	input \WX9840_reg/NET0131  ;
	input \WX9842_reg/NET0131  ;
	input \WX9844_reg/NET0131  ;
	input \WX9846_reg/NET0131  ;
	input \WX9848_reg/NET0131  ;
	input \WX9850_reg/NET0131  ;
	input \WX9852_reg/NET0131  ;
	input \WX9854_reg/NET0131  ;
	input \WX9856_reg/NET0131  ;
	input \WX9858_reg/NET0131  ;
	input \WX9860_reg/NET0131  ;
	input \WX9862_reg/NET0131  ;
	input \WX9864_reg/NET0131  ;
	input \WX9866_reg/NET0131  ;
	input \WX9868_reg/NET0131  ;
	input \WX9870_reg/NET0131  ;
	input \WX9872_reg/NET0131  ;
	input \WX9874_reg/NET0131  ;
	input \WX9876_reg/NET0131  ;
	input \WX9878_reg/NET0131  ;
	input \WX9880_reg/NET0131  ;
	input \WX9882_reg/NET0131  ;
	input \WX9884_reg/NET0131  ;
	input \WX9886_reg/NET0131  ;
	input \WX9888_reg/NET0131  ;
	input \WX9890_reg/NET0131  ;
	input \WX9892_reg/NET0131  ;
	input \WX9894_reg/NET0131  ;
	input \WX9896_reg/NET0131  ;
	input \WX9898_reg/NET0131  ;
	input \WX9900_reg/NET0131  ;
	input \WX9902_reg/NET0131  ;
	input \WX9904_reg/NET0131  ;
	input \WX9906_reg/NET0131  ;
	input \WX9908_reg/NET0131  ;
	input \WX9910_reg/NET0131  ;
	input \WX9912_reg/NET0131  ;
	input \WX9914_reg/NET0131  ;
	input \WX9916_reg/NET0131  ;
	input \WX9918_reg/NET0131  ;
	input \WX9920_reg/NET0131  ;
	input \WX9922_reg/NET0131  ;
	input \WX9924_reg/NET0131  ;
	input \WX9926_reg/NET0131  ;
	input \WX9928_reg/NET0131  ;
	input \WX9930_reg/NET0131  ;
	input \WX9932_reg/NET0131  ;
	input \WX9934_reg/NET0131  ;
	input \WX9936_reg/NET0131  ;
	input \WX9938_reg/NET0131  ;
	input \WX9940_reg/NET0131  ;
	input \WX9942_reg/NET0131  ;
	input \WX9944_reg/NET0131  ;
	input \WX9946_reg/NET0131  ;
	input \WX9948_reg/NET0131  ;
	input \WX9950_reg/NET0131  ;
	input \_2077__reg/NET0131  ;
	input \_2078__reg/NET0131  ;
	input \_2079__reg/NET0131  ;
	input \_2080__reg/NET0131  ;
	input \_2081__reg/NET0131  ;
	input \_2082__reg/NET0131  ;
	input \_2083__reg/NET0131  ;
	input \_2084__reg/NET0131  ;
	input \_2085__reg/NET0131  ;
	input \_2086__reg/NET0131  ;
	input \_2087__reg/NET0131  ;
	input \_2088__reg/NET0131  ;
	input \_2089__reg/NET0131  ;
	input \_2090__reg/NET0131  ;
	input \_2091__reg/NET0131  ;
	input \_2092__reg/NET0131  ;
	input \_2093__reg/NET0131  ;
	input \_2094__reg/NET0131  ;
	input \_2095__reg/NET0131  ;
	input \_2096__reg/NET0131  ;
	input \_2097__reg/NET0131  ;
	input \_2098__reg/NET0131  ;
	input \_2099__reg/NET0131  ;
	input \_2100__reg/NET0131  ;
	input \_2101__reg/NET0131  ;
	input \_2102__reg/NET0131  ;
	input \_2103__reg/NET0131  ;
	input \_2104__reg/NET0131  ;
	input \_2105__reg/NET0131  ;
	input \_2106__reg/NET0131  ;
	input \_2107__reg/NET0131  ;
	input \_2108__reg/NET0131  ;
	input \_2109__reg/NET0131  ;
	input \_2110__reg/NET0131  ;
	input \_2111__reg/NET0131  ;
	input \_2112__reg/NET0131  ;
	input \_2113__reg/NET0131  ;
	input \_2114__reg/NET0131  ;
	input \_2115__reg/NET0131  ;
	input \_2116__reg/NET0131  ;
	input \_2117__reg/NET0131  ;
	input \_2118__reg/NET0131  ;
	input \_2119__reg/NET0131  ;
	input \_2120__reg/NET0131  ;
	input \_2121__reg/NET0131  ;
	input \_2122__reg/NET0131  ;
	input \_2123__reg/NET0131  ;
	input \_2124__reg/NET0131  ;
	input \_2125__reg/NET0131  ;
	input \_2126__reg/NET0131  ;
	input \_2127__reg/NET0131  ;
	input \_2128__reg/NET0131  ;
	input \_2129__reg/NET0131  ;
	input \_2130__reg/NET0131  ;
	input \_2131__reg/NET0131  ;
	input \_2132__reg/NET0131  ;
	input \_2133__reg/NET0131  ;
	input \_2134__reg/NET0131  ;
	input \_2135__reg/NET0131  ;
	input \_2136__reg/NET0131  ;
	input \_2137__reg/NET0131  ;
	input \_2138__reg/NET0131  ;
	input \_2139__reg/NET0131  ;
	input \_2140__reg/NET0131  ;
	input \_2141__reg/NET0131  ;
	input \_2142__reg/NET0131  ;
	input \_2143__reg/NET0131  ;
	input \_2144__reg/NET0131  ;
	input \_2145__reg/NET0131  ;
	input \_2146__reg/NET0131  ;
	input \_2147__reg/NET0131  ;
	input \_2148__reg/NET0131  ;
	input \_2149__reg/NET0131  ;
	input \_2150__reg/NET0131  ;
	input \_2151__reg/NET0131  ;
	input \_2152__reg/NET0131  ;
	input \_2153__reg/NET0131  ;
	input \_2154__reg/NET0131  ;
	input \_2155__reg/NET0131  ;
	input \_2156__reg/NET0131  ;
	input \_2157__reg/NET0131  ;
	input \_2158__reg/NET0131  ;
	input \_2159__reg/NET0131  ;
	input \_2160__reg/NET0131  ;
	input \_2161__reg/NET0131  ;
	input \_2162__reg/NET0131  ;
	input \_2163__reg/NET0131  ;
	input \_2164__reg/NET0131  ;
	input \_2165__reg/NET0131  ;
	input \_2166__reg/NET0131  ;
	input \_2167__reg/NET0131  ;
	input \_2168__reg/NET0131  ;
	input \_2169__reg/NET0131  ;
	input \_2170__reg/NET0131  ;
	input \_2171__reg/NET0131  ;
	input \_2172__reg/NET0131  ;
	input \_2173__reg/NET0131  ;
	input \_2174__reg/NET0131  ;
	input \_2175__reg/NET0131  ;
	input \_2176__reg/NET0131  ;
	input \_2177__reg/NET0131  ;
	input \_2178__reg/NET0131  ;
	input \_2179__reg/NET0131  ;
	input \_2180__reg/NET0131  ;
	input \_2181__reg/NET0131  ;
	input \_2182__reg/NET0131  ;
	input \_2183__reg/NET0131  ;
	input \_2184__reg/NET0131  ;
	input \_2185__reg/NET0131  ;
	input \_2186__reg/NET0131  ;
	input \_2187__reg/NET0131  ;
	input \_2188__reg/NET0131  ;
	input \_2189__reg/NET0131  ;
	input \_2190__reg/NET0131  ;
	input \_2191__reg/NET0131  ;
	input \_2192__reg/NET0131  ;
	input \_2193__reg/NET0131  ;
	input \_2194__reg/NET0131  ;
	input \_2195__reg/NET0131  ;
	input \_2196__reg/NET0131  ;
	input \_2197__reg/NET0131  ;
	input \_2198__reg/NET0131  ;
	input \_2199__reg/NET0131  ;
	input \_2200__reg/NET0131  ;
	input \_2201__reg/NET0131  ;
	input \_2202__reg/NET0131  ;
	input \_2203__reg/NET0131  ;
	input \_2204__reg/NET0131  ;
	input \_2205__reg/NET0131  ;
	input \_2206__reg/NET0131  ;
	input \_2207__reg/NET0131  ;
	input \_2208__reg/NET0131  ;
	input \_2209__reg/NET0131  ;
	input \_2210__reg/NET0131  ;
	input \_2211__reg/NET0131  ;
	input \_2212__reg/NET0131  ;
	input \_2213__reg/NET0131  ;
	input \_2214__reg/NET0131  ;
	input \_2215__reg/NET0131  ;
	input \_2216__reg/NET0131  ;
	input \_2217__reg/NET0131  ;
	input \_2218__reg/NET0131  ;
	input \_2219__reg/NET0131  ;
	input \_2220__reg/NET0131  ;
	input \_2221__reg/NET0131  ;
	input \_2222__reg/NET0131  ;
	input \_2223__reg/NET0131  ;
	input \_2224__reg/NET0131  ;
	input \_2225__reg/NET0131  ;
	input \_2226__reg/NET0131  ;
	input \_2227__reg/NET0131  ;
	input \_2228__reg/NET0131  ;
	input \_2229__reg/NET0131  ;
	input \_2230__reg/NET0131  ;
	input \_2231__reg/NET0131  ;
	input \_2232__reg/NET0131  ;
	input \_2233__reg/NET0131  ;
	input \_2234__reg/NET0131  ;
	input \_2235__reg/NET0131  ;
	input \_2236__reg/NET0131  ;
	input \_2237__reg/NET0131  ;
	input \_2238__reg/NET0131  ;
	input \_2239__reg/NET0131  ;
	input \_2240__reg/NET0131  ;
	input \_2241__reg/NET0131  ;
	input \_2242__reg/NET0131  ;
	input \_2243__reg/NET0131  ;
	input \_2244__reg/NET0131  ;
	input \_2245__reg/NET0131  ;
	input \_2246__reg/NET0131  ;
	input \_2247__reg/NET0131  ;
	input \_2248__reg/NET0131  ;
	input \_2249__reg/NET0131  ;
	input \_2250__reg/NET0131  ;
	input \_2251__reg/NET0131  ;
	input \_2252__reg/NET0131  ;
	input \_2253__reg/NET0131  ;
	input \_2254__reg/NET0131  ;
	input \_2255__reg/NET0131  ;
	input \_2256__reg/NET0131  ;
	input \_2257__reg/NET0131  ;
	input \_2258__reg/NET0131  ;
	input \_2259__reg/NET0131  ;
	input \_2260__reg/NET0131  ;
	input \_2261__reg/NET0131  ;
	input \_2262__reg/NET0131  ;
	input \_2263__reg/NET0131  ;
	input \_2264__reg/NET0131  ;
	input \_2265__reg/NET0131  ;
	input \_2266__reg/NET0131  ;
	input \_2267__reg/NET0131  ;
	input \_2268__reg/NET0131  ;
	input \_2269__reg/NET0131  ;
	input \_2270__reg/NET0131  ;
	input \_2271__reg/NET0131  ;
	input \_2272__reg/NET0131  ;
	input \_2273__reg/NET0131  ;
	input \_2274__reg/NET0131  ;
	input \_2275__reg/NET0131  ;
	input \_2276__reg/NET0131  ;
	input \_2277__reg/NET0131  ;
	input \_2278__reg/NET0131  ;
	input \_2279__reg/NET0131  ;
	input \_2280__reg/NET0131  ;
	input \_2281__reg/NET0131  ;
	input \_2282__reg/NET0131  ;
	input \_2283__reg/NET0131  ;
	input \_2284__reg/NET0131  ;
	input \_2285__reg/NET0131  ;
	input \_2286__reg/NET0131  ;
	input \_2287__reg/NET0131  ;
	input \_2288__reg/NET0131  ;
	input \_2289__reg/NET0131  ;
	input \_2290__reg/NET0131  ;
	input \_2291__reg/NET0131  ;
	input \_2292__reg/NET0131  ;
	input \_2293__reg/NET0131  ;
	input \_2294__reg/NET0131  ;
	input \_2295__reg/NET0131  ;
	input \_2296__reg/NET0131  ;
	input \_2297__reg/NET0131  ;
	input \_2298__reg/NET0131  ;
	input \_2299__reg/NET0131  ;
	input \_2300__reg/NET0131  ;
	input \_2301__reg/NET0131  ;
	input \_2302__reg/NET0131  ;
	input \_2303__reg/NET0131  ;
	input \_2304__reg/NET0131  ;
	input \_2305__reg/NET0131  ;
	input \_2306__reg/NET0131  ;
	input \_2307__reg/NET0131  ;
	input \_2308__reg/NET0131  ;
	input \_2309__reg/NET0131  ;
	input \_2310__reg/NET0131  ;
	input \_2311__reg/NET0131  ;
	input \_2312__reg/NET0131  ;
	input \_2313__reg/NET0131  ;
	input \_2314__reg/NET0131  ;
	input \_2315__reg/NET0131  ;
	input \_2316__reg/NET0131  ;
	input \_2317__reg/NET0131  ;
	input \_2318__reg/NET0131  ;
	input \_2319__reg/NET0131  ;
	input \_2320__reg/NET0131  ;
	input \_2321__reg/NET0131  ;
	input \_2322__reg/NET0131  ;
	input \_2323__reg/NET0131  ;
	input \_2324__reg/NET0131  ;
	input \_2325__reg/NET0131  ;
	input \_2326__reg/NET0131  ;
	input \_2327__reg/NET0131  ;
	input \_2328__reg/NET0131  ;
	input \_2329__reg/NET0131  ;
	input \_2330__reg/NET0131  ;
	input \_2331__reg/NET0131  ;
	input \_2332__reg/NET0131  ;
	input \_2333__reg/NET0131  ;
	input \_2334__reg/NET0131  ;
	input \_2335__reg/NET0131  ;
	input \_2336__reg/NET0131  ;
	input \_2337__reg/NET0131  ;
	input \_2338__reg/NET0131  ;
	input \_2339__reg/NET0131  ;
	input \_2340__reg/NET0131  ;
	input \_2341__reg/NET0131  ;
	input \_2342__reg/NET0131  ;
	input \_2343__reg/NET0131  ;
	input \_2344__reg/NET0131  ;
	input \_2345__reg/NET0131  ;
	input \_2346__reg/NET0131  ;
	input \_2347__reg/NET0131  ;
	input \_2348__reg/NET0131  ;
	input \_2349__reg/NET0131  ;
	input \_2350__reg/NET0131  ;
	input \_2351__reg/NET0131  ;
	input \_2352__reg/NET0131  ;
	input \_2353__reg/NET0131  ;
	input \_2354__reg/NET0131  ;
	input \_2355__reg/NET0131  ;
	input \_2356__reg/NET0131  ;
	input \_2357__reg/NET0131  ;
	input \_2358__reg/NET0131  ;
	input \_2359__reg/NET0131  ;
	input \_2360__reg/NET0131  ;
	input \_2361__reg/NET0131  ;
	input \_2362__reg/NET0131  ;
	input \_2363__reg/NET0131  ;
	input \_2364__reg/NET0131  ;
	output \DATA_9_0_pad  ;
	output \DATA_9_10_pad  ;
	output \DATA_9_11_pad  ;
	output \DATA_9_12_pad  ;
	output \DATA_9_13_pad  ;
	output \DATA_9_14_pad  ;
	output \DATA_9_15_pad  ;
	output \DATA_9_16_pad  ;
	output \DATA_9_17_pad  ;
	output \DATA_9_18_pad  ;
	output \DATA_9_19_pad  ;
	output \DATA_9_1_pad  ;
	output \DATA_9_20_pad  ;
	output \DATA_9_21_pad  ;
	output \DATA_9_22_pad  ;
	output \DATA_9_23_pad  ;
	output \DATA_9_24_pad  ;
	output \DATA_9_25_pad  ;
	output \DATA_9_26_pad  ;
	output \DATA_9_27_pad  ;
	output \DATA_9_28_pad  ;
	output \DATA_9_29_pad  ;
	output \DATA_9_2_pad  ;
	output \DATA_9_30_pad  ;
	output \DATA_9_31_pad  ;
	output \DATA_9_3_pad  ;
	output \DATA_9_4_pad  ;
	output \DATA_9_5_pad  ;
	output \DATA_9_6_pad  ;
	output \DATA_9_7_pad  ;
	output \DATA_9_8_pad  ;
	output \DATA_9_9_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g19/_0_  ;
	output \g35/_0_  ;
	output \g36/_0_  ;
	output \g40/_0_  ;
	output \g55780/_0_  ;
	output \g55783/_0_  ;
	output \g55795/_0_  ;
	output \g55796/_0_  ;
	output \g55797/_0_  ;
	output \g55798/_0_  ;
	output \g55799/_0_  ;
	output \g55800/_0_  ;
	output \g55801/_0_  ;
	output \g55802/_0_  ;
	output \g55803/_0_  ;
	output \g55834/_0_  ;
	output \g55835/_0_  ;
	output \g55836/_0_  ;
	output \g55837/_0_  ;
	output \g55838/_0_  ;
	output \g55839/_0_  ;
	output \g55840/_0_  ;
	output \g55841/_0_  ;
	output \g55842/_0_  ;
	output \g55856/_0_  ;
	output \g55894/_0_  ;
	output \g55895/_0_  ;
	output \g55896/_0_  ;
	output \g55897/_0_  ;
	output \g55898/_0_  ;
	output \g55899/_0_  ;
	output \g55900/_0_  ;
	output \g55901/_0_  ;
	output \g55902/_0_  ;
	output \g55916/_0_  ;
	output \g55953/_0_  ;
	output \g55954/_0_  ;
	output \g55955/_0_  ;
	output \g55956/_0_  ;
	output \g55957/_0_  ;
	output \g55958/_0_  ;
	output \g55959/_0_  ;
	output \g55960/_0_  ;
	output \g55961/_0_  ;
	output \g55975/_0_  ;
	output \g56012/_0_  ;
	output \g56013/_0_  ;
	output \g56014/_0_  ;
	output \g56015/_0_  ;
	output \g56016/_0_  ;
	output \g56017/_0_  ;
	output \g56018/_0_  ;
	output \g56019/_0_  ;
	output \g56020/_0_  ;
	output \g56034/_0_  ;
	output \g56071/_0_  ;
	output \g56072/_0_  ;
	output \g56073/_0_  ;
	output \g56074/_0_  ;
	output \g56075/_0_  ;
	output \g56076/_0_  ;
	output \g56077/_0_  ;
	output \g56078/_0_  ;
	output \g56079/_0_  ;
	output \g56093/_0_  ;
	output \g56130/_0_  ;
	output \g56131/_0_  ;
	output \g56132/_0_  ;
	output \g56133/_0_  ;
	output \g56134/_0_  ;
	output \g56135/_0_  ;
	output \g56136/_0_  ;
	output \g56137/_0_  ;
	output \g56138/_0_  ;
	output \g56152/_0_  ;
	output \g56189/_0_  ;
	output \g56190/_0_  ;
	output \g56191/_0_  ;
	output \g56192/_0_  ;
	output \g56193/_0_  ;
	output \g56194/_0_  ;
	output \g56195/_0_  ;
	output \g56196/_0_  ;
	output \g56197/_0_  ;
	output \g56211/_0_  ;
	output \g56248/_0_  ;
	output \g56249/_0_  ;
	output \g56250/_0_  ;
	output \g56251/_0_  ;
	output \g56252/_0_  ;
	output \g56253/_0_  ;
	output \g56254/_0_  ;
	output \g56255/_0_  ;
	output \g56256/_0_  ;
	output \g56270/_0_  ;
	output \g56307/_0_  ;
	output \g56308/_0_  ;
	output \g56309/_0_  ;
	output \g56310/_0_  ;
	output \g56311/_0_  ;
	output \g56312/_0_  ;
	output \g56313/_0_  ;
	output \g56314/_0_  ;
	output \g56315/_0_  ;
	output \g56329/_0_  ;
	output \g56366/_0_  ;
	output \g56367/_0_  ;
	output \g56368/_0_  ;
	output \g56369/_0_  ;
	output \g56370/_0_  ;
	output \g56371/_0_  ;
	output \g56372/_0_  ;
	output \g56373/_0_  ;
	output \g56374/_0_  ;
	output \g56388/_0_  ;
	output \g56425/_0_  ;
	output \g56426/_0_  ;
	output \g56427/_0_  ;
	output \g56428/_0_  ;
	output \g56429/_0_  ;
	output \g56430/_0_  ;
	output \g56431/_0_  ;
	output \g56432/_0_  ;
	output \g56433/_0_  ;
	output \g56447/_0_  ;
	output \g56484/_0_  ;
	output \g56485/_0_  ;
	output \g56486/_0_  ;
	output \g56487/_0_  ;
	output \g56488/_0_  ;
	output \g56489/_0_  ;
	output \g56490/_0_  ;
	output \g56491/_0_  ;
	output \g56492/_0_  ;
	output \g56507/_0_  ;
	output \g56543/_0_  ;
	output \g56544/_0_  ;
	output \g56545/_0_  ;
	output \g56546/_0_  ;
	output \g56547/_0_  ;
	output \g56548/_0_  ;
	output \g56549/_0_  ;
	output \g56551/_0_  ;
	output \g56567/_0_  ;
	output \g56602/_0_  ;
	output \g56603/_0_  ;
	output \g56604/_0_  ;
	output \g56605/_0_  ;
	output \g56606/_0_  ;
	output \g56607/_0_  ;
	output \g56608/_0_  ;
	output \g56610/_0_  ;
	output \g56627/_0_  ;
	output \g56661/_0_  ;
	output \g56662/_0_  ;
	output \g56663/_0_  ;
	output \g56664/_0_  ;
	output \g56665/_0_  ;
	output \g56666/_0_  ;
	output \g56667/_0_  ;
	output \g56668/_0_  ;
	output \g56686/_0_  ;
	output \g56720/_0_  ;
	output \g56721/_0_  ;
	output \g56722/_0_  ;
	output \g56723/_0_  ;
	output \g56724/_0_  ;
	output \g56725/_0_  ;
	output \g56726/_0_  ;
	output \g56727/_0_  ;
	output \g56728/_0_  ;
	output \g56745/_0_  ;
	output \g56779/_0_  ;
	output \g56780/_0_  ;
	output \g56781/_0_  ;
	output \g56782/_0_  ;
	output \g56783/_0_  ;
	output \g56784/_0_  ;
	output \g56785/_0_  ;
	output \g56804/_0_  ;
	output \g56838/_0_  ;
	output \g56839/_0_  ;
	output \g56840/_0_  ;
	output \g56841/_0_  ;
	output \g56842/_0_  ;
	output \g56843/_0_  ;
	output \g56844/_0_  ;
	output \g56845/_0_  ;
	output \g56846/_0_  ;
	output \g56863/_0_  ;
	output \g56897/_0_  ;
	output \g56898/_0_  ;
	output \g56899/_0_  ;
	output \g56900/_0_  ;
	output \g56901/_0_  ;
	output \g56902/_0_  ;
	output \g56903/_0_  ;
	output \g56905/_0_  ;
	output \g56921/_0_  ;
	output \g56956/_0_  ;
	output \g56957/_0_  ;
	output \g56958/_0_  ;
	output \g56959/_0_  ;
	output \g56960/_0_  ;
	output \g56961/_0_  ;
	output \g56962/_0_  ;
	output \g56964/_0_  ;
	output \g56980/_0_  ;
	output \g57015/_0_  ;
	output \g57016/_0_  ;
	output \g57017/_0_  ;
	output \g57018/_0_  ;
	output \g57019/_0_  ;
	output \g57020/_0_  ;
	output \g57021/_0_  ;
	output \g57023/_0_  ;
	output \g57040/_0_  ;
	output \g57074/_0_  ;
	output \g57075/_0_  ;
	output \g57076/_0_  ;
	output \g57077/_0_  ;
	output \g57078/_0_  ;
	output \g57079/_0_  ;
	output \g57080/_0_  ;
	output \g57081/_0_  ;
	output \g57099/_0_  ;
	output \g57133/_0_  ;
	output \g57134/_0_  ;
	output \g57135/_0_  ;
	output \g57136/_0_  ;
	output \g57137/_0_  ;
	output \g57138/_0_  ;
	output \g57139/_0_  ;
	output \g57140/_0_  ;
	output \g57141/_0_  ;
	output \g57159/_0_  ;
	output \g57193/_0_  ;
	output \g57195/_0_  ;
	output \g57196/_0_  ;
	output \g57197/_0_  ;
	output \g57198/_0_  ;
	output \g57199/_0_  ;
	output \g57200/_0_  ;
	output \g57202/_0_  ;
	output \g57219/_0_  ;
	output \g57254/_0_  ;
	output \g57255/_0_  ;
	output \g57256/_0_  ;
	output \g57257/_0_  ;
	output \g57258/_0_  ;
	output \g57259/_0_  ;
	output \g57260/_0_  ;
	output \g57262/_0_  ;
	output \g57263/_0_  ;
	output \g57285/_0_  ;
	output \g57318/_0_  ;
	output \g57319/_0_  ;
	output \g57320/_0_  ;
	output \g57321/_0_  ;
	output \g57322/_0_  ;
	output \g57323/_0_  ;
	output \g57324/_0_  ;
	output \g57325/_0_  ;
	output \g57326/_0_  ;
	output \g57328/_0_  ;
	output \g57329/_0_  ;
	output \g57330/_0_  ;
	output \g57350/_0_  ;
	output \g57387/_0_  ;
	output \g57388/_0_  ;
	output \g57390/_0_  ;
	output \g57391/_0_  ;
	output \g57392/_0_  ;
	output \g57393/_0_  ;
	output \g57395/_0_  ;
	output \g57396/_0_  ;
	output \g57439/_0_  ;
	output \g57476/_0_  ;
	output \g57477/_0_  ;
	output \g57478/_0_  ;
	output \g57479/_0_  ;
	output \g57480/_0_  ;
	output \g57481/_0_  ;
	output \g57482/_0_  ;
	output \g57483/_0_  ;
	output \g57484/_0_  ;
	output \g57485/_0_  ;
	output \g57486/_0_  ;
	output \g57487/_0_  ;
	output \g57488/_0_  ;
	output \g57489/_0_  ;
	output \g57490/_0_  ;
	output \g57491/_0_  ;
	output \g57492/_0_  ;
	output \g57493/_0_  ;
	output \g57494/_0_  ;
	output \g57495/_0_  ;
	output \g57496/_0_  ;
	output \g57497/_0_  ;
	output \g57498/_0_  ;
	output \g57499/_0_  ;
	output \g57500/_0_  ;
	output \g57501/_0_  ;
	output \g57502/_0_  ;
	output \g57503/_0_  ;
	output \g57504/_0_  ;
	output \g57505/_0_  ;
	output \g57524/_0_  ;
	output \g57537/_0_  ;
	output \g57541/_0_  ;
	output \g57543/_0_  ;
	output \g58163/_0_  ;
	output \g58572/_0_  ;
	output \g58573/_0_  ;
	output \g58574/_0_  ;
	output \g58575/_0_  ;
	output \g58576/_0_  ;
	output \g58577/_0_  ;
	output \g58578/_0_  ;
	output \g58579/_0_  ;
	output \g58580/_0_  ;
	output \g58581/_0_  ;
	output \g58582/_0_  ;
	output \g58583/_0_  ;
	output \g58584/_0_  ;
	output \g58585/_0_  ;
	output \g58586/_0_  ;
	output \g58587/_0_  ;
	output \g58588/_0_  ;
	output \g58589/_0_  ;
	output \g58590/_0_  ;
	output \g58591/_0_  ;
	output \g58592/_0_  ;
	output \g58593/_0_  ;
	output \g58594/_0_  ;
	output \g58595/_0_  ;
	output \g58596/_0_  ;
	output \g58597/_0_  ;
	output \g58598/_0_  ;
	output \g58600/_0_  ;
	output \g58602/_0_  ;
	output \g58604/_0_  ;
	output \g58615/_0_  ;
	output \g59240/_0_  ;
	output \g59241/_0_  ;
	output \g59242/_0_  ;
	output \g59243/_0_  ;
	output \g59244/_0_  ;
	output \g59245/_0_  ;
	output \g59246/_0_  ;
	output \g59247/_0_  ;
	output \g59248/_0_  ;
	output \g59249/_0_  ;
	output \g59250/_0_  ;
	output \g59251/_0_  ;
	output \g59252/_0_  ;
	output \g59253/_0_  ;
	output \g59254/_0_  ;
	output \g59255/_0_  ;
	output \g59256/_0_  ;
	output \g59257/_0_  ;
	output \g59258/_0_  ;
	output \g59259/_0_  ;
	output \g59260/_0_  ;
	output \g59261/_0_  ;
	output \g59262/_0_  ;
	output \g59263/_0_  ;
	output \g59264/_0_  ;
	output \g59265/_0_  ;
	output \g59266/_0_  ;
	output \g59267/_0_  ;
	output \g59268/_0_  ;
	output \g59269/_0_  ;
	output \g59270/_0_  ;
	output \g59271/_0_  ;
	output \g59272/_0_  ;
	output \g59273/_0_  ;
	output \g59274/_0_  ;
	output \g59275/_0_  ;
	output \g59276/_0_  ;
	output \g59277/_0_  ;
	output \g59278/_0_  ;
	output \g59279/_0_  ;
	output \g59280/_0_  ;
	output \g59281/_0_  ;
	output \g59282/_0_  ;
	output \g59283/_0_  ;
	output \g59284/_0_  ;
	output \g59285/_0_  ;
	output \g59286/_0_  ;
	output \g59287/_0_  ;
	output \g59288/_0_  ;
	output \g59289/_0_  ;
	output \g59290/_0_  ;
	output \g59291/_0_  ;
	output \g59292/_0_  ;
	output \g59293/_0_  ;
	output \g59294/_0_  ;
	output \g59295/_0_  ;
	output \g59296/_0_  ;
	output \g59297/_0_  ;
	output \g59298/_0_  ;
	output \g59299/_0_  ;
	output \g59300/_0_  ;
	output \g59301/_0_  ;
	output \g59302/_0_  ;
	output \g59303/_0_  ;
	output \g59304/_0_  ;
	output \g59305/_0_  ;
	output \g59306/_0_  ;
	output \g59307/_0_  ;
	output \g59308/_0_  ;
	output \g59309/_0_  ;
	output \g59310/_0_  ;
	output \g59311/_0_  ;
	output \g59312/_0_  ;
	output \g59313/_0_  ;
	output \g59314/_0_  ;
	output \g59315/_0_  ;
	output \g59316/_0_  ;
	output \g59317/_0_  ;
	output \g59318/_0_  ;
	output \g59319/_0_  ;
	output \g59320/_0_  ;
	output \g59321/_0_  ;
	output \g59322/_0_  ;
	output \g59323/_0_  ;
	output \g59324/_0_  ;
	output \g59325/_0_  ;
	output \g59326/_0_  ;
	output \g59327/_0_  ;
	output \g59328/_0_  ;
	output \g59329/_0_  ;
	output \g59330/_0_  ;
	output \g59331/_0_  ;
	output \g59332/_0_  ;
	output \g59333/_0_  ;
	output \g59334/_0_  ;
	output \g59335/_0_  ;
	output \g59336/_0_  ;
	output \g59337/_0_  ;
	output \g59338/_0_  ;
	output \g59339/_0_  ;
	output \g59340/_0_  ;
	output \g59341/_0_  ;
	output \g59342/_0_  ;
	output \g59343/_0_  ;
	output \g59344/_0_  ;
	output \g59345/_0_  ;
	output \g59346/_0_  ;
	output \g59347/_0_  ;
	output \g59348/_0_  ;
	output \g59349/_0_  ;
	output \g59350/_0_  ;
	output \g59351/_0_  ;
	output \g59352/_0_  ;
	output \g59353/_0_  ;
	output \g59354/_0_  ;
	output \g59355/_0_  ;
	output \g59356/_0_  ;
	output \g59357/_0_  ;
	output \g59358/_0_  ;
	output \g59359/_0_  ;
	output \g59360/_0_  ;
	output \g59361/_0_  ;
	output \g59362/_0_  ;
	output \g59363/_0_  ;
	output \g59364/_0_  ;
	output \g59365/_0_  ;
	output \g59366/_0_  ;
	output \g59367/_0_  ;
	output \g59368/_0_  ;
	output \g59369/_0_  ;
	output \g59370/_0_  ;
	output \g59371/_0_  ;
	output \g59372/_0_  ;
	output \g59373/_0_  ;
	output \g59374/_0_  ;
	output \g59375/_0_  ;
	output \g59376/_0_  ;
	output \g59377/_0_  ;
	output \g59378/_0_  ;
	output \g59379/_0_  ;
	output \g59380/_0_  ;
	output \g59381/_0_  ;
	output \g59382/_0_  ;
	output \g59383/_0_  ;
	output \g59384/_0_  ;
	output \g59385/_0_  ;
	output \g59386/_0_  ;
	output \g59387/_0_  ;
	output \g59388/_0_  ;
	output \g59389/_0_  ;
	output \g59390/_0_  ;
	output \g59391/_0_  ;
	output \g59392/_0_  ;
	output \g59393/_0_  ;
	output \g59394/_0_  ;
	output \g59395/_0_  ;
	output \g59396/_0_  ;
	output \g59397/_0_  ;
	output \g59398/_0_  ;
	output \g59399/_0_  ;
	output \g59400/_0_  ;
	output \g59401/_0_  ;
	output \g59402/_0_  ;
	output \g59403/_0_  ;
	output \g59404/_0_  ;
	output \g59405/_0_  ;
	output \g59406/_0_  ;
	output \g59407/_0_  ;
	output \g59408/_0_  ;
	output \g59409/_0_  ;
	output \g59410/_0_  ;
	output \g59411/_0_  ;
	output \g59412/_0_  ;
	output \g59413/_0_  ;
	output \g59414/_0_  ;
	output \g59415/_0_  ;
	output \g59416/_0_  ;
	output \g59417/_0_  ;
	output \g59418/_0_  ;
	output \g59419/_0_  ;
	output \g59420/_0_  ;
	output \g59421/_0_  ;
	output \g59422/_0_  ;
	output \g59423/_0_  ;
	output \g59424/_0_  ;
	output \g59425/_0_  ;
	output \g59426/_0_  ;
	output \g59427/_0_  ;
	output \g59428/_0_  ;
	output \g59429/_0_  ;
	output \g59430/_0_  ;
	output \g59431/_0_  ;
	output \g59432/_0_  ;
	output \g59433/_0_  ;
	output \g59434/_0_  ;
	output \g59435/_0_  ;
	output \g59436/_0_  ;
	output \g59437/_0_  ;
	output \g59438/_0_  ;
	output \g59439/_0_  ;
	output \g59440/_0_  ;
	output \g59441/_0_  ;
	output \g59442/_0_  ;
	output \g59443/_0_  ;
	output \g59444/_0_  ;
	output \g59445/_0_  ;
	output \g59446/_0_  ;
	output \g59447/_0_  ;
	output \g59448/_0_  ;
	output \g59449/_0_  ;
	output \g59450/_0_  ;
	output \g59451/_0_  ;
	output \g59452/_0_  ;
	output \g59453/_0_  ;
	output \g59454/_0_  ;
	output \g59455/_0_  ;
	output \g59456/_0_  ;
	output \g59457/_0_  ;
	output \g59458/_0_  ;
	output \g59459/_0_  ;
	output \g59460/_0_  ;
	output \g59461/_0_  ;
	output \g59462/_0_  ;
	output \g59463/_0_  ;
	output \g59464/_0_  ;
	output \g59465/_0_  ;
	output \g59466/_0_  ;
	output \g59467/_0_  ;
	output \g59468/_0_  ;
	output \g59469/_0_  ;
	output \g59470/_0_  ;
	output \g59471/_0_  ;
	output \g59472/_0_  ;
	output \g59473/_0_  ;
	output \g59474/_0_  ;
	output \g59475/_0_  ;
	output \g59476/_0_  ;
	output \g59477/_0_  ;
	output \g59478/_0_  ;
	output \g59479/_0_  ;
	output \g59480/_0_  ;
	output \g59481/_0_  ;
	output \g59482/_0_  ;
	output \g59483/_0_  ;
	output \g59484/_0_  ;
	output \g59485/_0_  ;
	output \g59486/_0_  ;
	output \g59487/_0_  ;
	output \g59488/_0_  ;
	output \g59489/_0_  ;
	output \g59490/_0_  ;
	output \g59491/_0_  ;
	output \g59492/_0_  ;
	output \g59493/_0_  ;
	output \g59494/_0_  ;
	output \g59495/_0_  ;
	output \g59496/_0_  ;
	output \g59497/_0_  ;
	output \g59498/_0_  ;
	output \g59500/_0_  ;
	output \g59503/_0_  ;
	output \g59512/_0_  ;
	output \g61336/_0_  ;
	output \g61521/_0_  ;
	output \g61523/_0_  ;
	output \g61524/_0_  ;
	output \g61526/_0_  ;
	output \g61527/_0_  ;
	output \g61528/_0_  ;
	output \g61529/_0_  ;
	output \g61530/_0_  ;
	output \g61531/_0_  ;
	output \g61532/_0_  ;
	output \g61533/_0_  ;
	output \g61535/_0_  ;
	output \g61537/_0_  ;
	output \g61539/_0_  ;
	output \g61540/_0_  ;
	output \g61541/_0_  ;
	output \g61542/_0_  ;
	output \g61546/_0_  ;
	output \g61550/_0_  ;
	output \g61551/_0_  ;
	output \g61552/_0_  ;
	output \g61554/_0_  ;
	output \g61555/_0_  ;
	output \g61556/_0_  ;
	output \g61558/_0_  ;
	output \g61559/_0_  ;
	output \g61561/_0_  ;
	output \g61562/_0_  ;
	output \g61563/_0_  ;
	output \g61564/_0_  ;
	output \g61565/_0_  ;
	output \g61566/_0_  ;
	output \g61568/_0_  ;
	output \g61570/_0_  ;
	output \g61571/_0_  ;
	output \g61572/_0_  ;
	output \g61573/_0_  ;
	output \g61577/_0_  ;
	output \g61578/_0_  ;
	output \g61579/_0_  ;
	output \g61580/_0_  ;
	output \g61581/_0_  ;
	output \g61582/_0_  ;
	output \g61583/_0_  ;
	output \g61584/_0_  ;
	output \g61585/_0_  ;
	output \g61586/_0_  ;
	output \g61587/_0_  ;
	output \g61588/_0_  ;
	output \g61589/_0_  ;
	output \g61591/_0_  ;
	output \g61592/_0_  ;
	output \g61594/_0_  ;
	output \g61595/_0_  ;
	output \g61596/_0_  ;
	output \g61597/_0_  ;
	output \g61598/_0_  ;
	output \g61599/_0_  ;
	output \g61600/_0_  ;
	output \g61601/_0_  ;
	output \g61605/_0_  ;
	output \g61606/_0_  ;
	output \g61607/_0_  ;
	output \g61608/_0_  ;
	output \g61609/_0_  ;
	output \g61610/_0_  ;
	output \g61611/_0_  ;
	output \g61612/_0_  ;
	output \g61613/_0_  ;
	output \g61615/_0_  ;
	output \g61616/_0_  ;
	output \g61617/_0_  ;
	output \g61618/_0_  ;
	output \g61619/_0_  ;
	output \g61620/_0_  ;
	output \g61621/_0_  ;
	output \g61623/_0_  ;
	output \g61624/_0_  ;
	output \g61625/_0_  ;
	output \g61626/_0_  ;
	output \g61627/_0_  ;
	output \g61629/_0_  ;
	output \g61630/_0_  ;
	output \g61631/_0_  ;
	output \g61632/_0_  ;
	output \g61633/_0_  ;
	output \g61634/_0_  ;
	output \g61636/_0_  ;
	output \g61638/_0_  ;
	output \g61639/_0_  ;
	output \g61640/_0_  ;
	output \g61641/_0_  ;
	output \g61642/_0_  ;
	output \g61644/_0_  ;
	output \g61647/_0_  ;
	output \g61648/_0_  ;
	output \g61649/_0_  ;
	output \g61650/_0_  ;
	output \g61653/_0_  ;
	output \g61654/_0_  ;
	output \g61655/_0_  ;
	output \g61656/_0_  ;
	output \g61658/_0_  ;
	output \g61661/_0_  ;
	output \g61662/_0_  ;
	output \g61663/_0_  ;
	output \g61664/_0_  ;
	output \g61666/_0_  ;
	output \g61667/_0_  ;
	output \g61668/_0_  ;
	output \g61670/_0_  ;
	output \g61671/_0_  ;
	output \g61672/_0_  ;
	output \g61673/_0_  ;
	output \g61675/_0_  ;
	output \g61676/_0_  ;
	output \g61680/_0_  ;
	output \g61681/_0_  ;
	output \g61682/_0_  ;
	output \g61683/_0_  ;
	output \g61684/_0_  ;
	output \g61686/_0_  ;
	output \g61687/_0_  ;
	output \g61688/_0_  ;
	output \g61689/_0_  ;
	output \g61690/_0_  ;
	output \g61691/_0_  ;
	output \g61693/_0_  ;
	output \g61694/_0_  ;
	output \g61696/_0_  ;
	output \g61697/_0_  ;
	output \g61698/_0_  ;
	output \g61699/_0_  ;
	output \g61700/_0_  ;
	output \g61701/_0_  ;
	output \g61702/_0_  ;
	output \g61703/_0_  ;
	output \g61704/_0_  ;
	output \g61705/_0_  ;
	output \g61706/_0_  ;
	output \g61707/_0_  ;
	output \g61708/_0_  ;
	output \g61711/_0_  ;
	output \g61712/_0_  ;
	output \g61714/_0_  ;
	output \g61716/_0_  ;
	output \g61717/_0_  ;
	output \g61719/_0_  ;
	output \g61720/_0_  ;
	output \g61721/_0_  ;
	output \g61724/_0_  ;
	output \g61725/_0_  ;
	output \g61728/_0_  ;
	output \g61729/_0_  ;
	output \g61731/_0_  ;
	output \g61732/_0_  ;
	output \g61733/_0_  ;
	output \g61736/_0_  ;
	output \g61737/_0_  ;
	output \g61739/_0_  ;
	output \g61740/_0_  ;
	output \g61741/_0_  ;
	output \g61743/_0_  ;
	output \g61744/_0_  ;
	output \g61745/_0_  ;
	output \g61746/_0_  ;
	output \g61747/_0_  ;
	output \g61748/_0_  ;
	output \g61749/_0_  ;
	output \g61750/_0_  ;
	output \g61751/_0_  ;
	output \g61752/_0_  ;
	output \g61753/_0_  ;
	output \g61754/_0_  ;
	output \g61755/_0_  ;
	output \g61757/_0_  ;
	output \g61758/_0_  ;
	output \g61759/_0_  ;
	output \g61760/_0_  ;
	output \g61761/_0_  ;
	output \g61762/_0_  ;
	output \g61763/_0_  ;
	output \g61764/_0_  ;
	output \g61765/_0_  ;
	output \g61766/_0_  ;
	output \g61767/_0_  ;
	output \g61768/_0_  ;
	output \g61769/_0_  ;
	output \g61770/_0_  ;
	output \g61771/_0_  ;
	output \g61772/_0_  ;
	output \g61773/_0_  ;
	output \g61774/_0_  ;
	output \g61775/_0_  ;
	output \g61776/_0_  ;
	output \g61777/_0_  ;
	output \g61778/_0_  ;
	output \g61780/_0_  ;
	output \g61781/_0_  ;
	output \g61783/_0_  ;
	output \g61784/_0_  ;
	output \g61786/_0_  ;
	output \g61787/_0_  ;
	output \g61790/_0_  ;
	output \g61791/_0_  ;
	output \g61794/_0_  ;
	output \g61795/_0_  ;
	output \g61796/_0_  ;
	output \g61797/_0_  ;
	output \g61798/_0_  ;
	output \g61799/_0_  ;
	output \g61800/_0_  ;
	output \g61801/_0_  ;
	output \g61802/_0_  ;
	output \g61803/_0_  ;
	output \g61805/_0_  ;
	output \g61806/_0_  ;
	output \g61807/_0_  ;
	output \g61808/_0_  ;
	output \g61809/_0_  ;
	output \g61810/_0_  ;
	output \g61811/_0_  ;
	output \g61812/_0_  ;
	output \g61813/_0_  ;
	output \g61816/_0_  ;
	output \g61817/_0_  ;
	output \g61818/_0_  ;
	output \g61820/_0_  ;
	output \g61822/_0_  ;
	output \g61823/_0_  ;
	output \g61825/_0_  ;
	output \g61826/_0_  ;
	output \g61827/_0_  ;
	output \g61828/_0_  ;
	output \g61829/_0_  ;
	output \g61832/_0_  ;
	output \g61834/_0_  ;
	output \g61835/_0_  ;
	output \g61837/_0_  ;
	output \g61838/_0_  ;
	output \g61839/_0_  ;
	output \g61840/_0_  ;
	output \g61844/_0_  ;
	output \g61847/_0_  ;
	output \g61848/_0_  ;
	output \g61849/_0_  ;
	output \g61850/_0_  ;
	output \g61851/_0_  ;
	output \g61853/_0_  ;
	output \g61854/_0_  ;
	output \g61855/_0_  ;
	output \g61856/_0_  ;
	output \g61858/_0_  ;
	output \g61859/_0_  ;
	output \g61861/_0_  ;
	output \g61862/_0_  ;
	output \g61863/_0_  ;
	output \g61864/_0_  ;
	output \g61865/_0_  ;
	output \g61866/_0_  ;
	output \g61867/_0_  ;
	output \g61868/_0_  ;
	output \g61869/_0_  ;
	output \g61870/_0_  ;
	output \g61871/_0_  ;
	output \g61873/_0_  ;
	output \g61874/_0_  ;
	output \g61875/_0_  ;
	output \g61877/_0_  ;
	output \g61878/_0_  ;
	output \g61879/_0_  ;
	output \g61880/_0_  ;
	output \g61881/_0_  ;
	output \g61883/_0_  ;
	output \g61884/_0_  ;
	output \g61886/_0_  ;
	output \g61887/_0_  ;
	output \g61890/_0_  ;
	output \g61891/_0_  ;
	output \g61892/_0_  ;
	output \g61893/_0_  ;
	output \g61894/_0_  ;
	output \g61895/_0_  ;
	output \g61900/_0_  ;
	output \g61901/_0_  ;
	output \g61902/_0_  ;
	output \g61904/_0_  ;
	output \g61905/_0_  ;
	output \g61906/_0_  ;
	output \g61907/_0_  ;
	output \g61914/_0_  ;
	output \g61915/_0_  ;
	output \g61917/_0_  ;
	output \g61919/_0_  ;
	output \g61921/_0_  ;
	output \g61924/_0_  ;
	output \g61925/_0_  ;
	output \g61926/_0_  ;
	output \g61927/_0_  ;
	output \g61928/_0_  ;
	output \g61929/_0_  ;
	output \g61930/_0_  ;
	output \g61931/_0_  ;
	output \g61932/_0_  ;
	output \g61933/_0_  ;
	output \g61934/_0_  ;
	output \g61935/_0_  ;
	output \g61936/_0_  ;
	output \g61937/_0_  ;
	output \g61938/_0_  ;
	output \g61939/_0_  ;
	output \g61943/_0_  ;
	output \g61944/_0_  ;
	output \g61945/_0_  ;
	output \g61947/_0_  ;
	output \g61948/_0_  ;
	output \g61949/_0_  ;
	output \g61950/_0_  ;
	output \g61951/_0_  ;
	output \g61952/_0_  ;
	output \g61953/_0_  ;
	output \g61955/_0_  ;
	output \g61956/_0_  ;
	output \g61957/_0_  ;
	output \g61958/_0_  ;
	output \g61959/_0_  ;
	output \g61960/_0_  ;
	output \g61961/_0_  ;
	output \g61962/_0_  ;
	output \g61963/_0_  ;
	output \g61964/_0_  ;
	output \g61965/_0_  ;
	output \g61966/_0_  ;
	output \g61967/_0_  ;
	output \g61968/_0_  ;
	output \g61969/_0_  ;
	output \g61970/_0_  ;
	output \g61971/_0_  ;
	output \g61972/_0_  ;
	output \g61973/_0_  ;
	output \g61974/_0_  ;
	output \g61976/_0_  ;
	output \g61978/_0_  ;
	output \g61980/_0_  ;
	output \g61981/_0_  ;
	output \g61982/_0_  ;
	output \g61983/_0_  ;
	output \g61984/_0_  ;
	output \g61985/_0_  ;
	output \g61986/_0_  ;
	output \g61987/_0_  ;
	output \g61988/_0_  ;
	output \g61989/_0_  ;
	output \g61990/_0_  ;
	output \g61992/_0_  ;
	output \g61994/_0_  ;
	output \g61995/_0_  ;
	output \g61996/_0_  ;
	output \g61997/_0_  ;
	output \g61998/_0_  ;
	output \g62000/_0_  ;
	output \g62001/_0_  ;
	output \g62002/_0_  ;
	output \g62003/_0_  ;
	output \g62004/_0_  ;
	output \g62005/_0_  ;
	output \g62007/_0_  ;
	output \g62008/_0_  ;
	output \g62009/_0_  ;
	output \g62010/_0_  ;
	output \g62011/_0_  ;
	output \g62012/_0_  ;
	output \g62013/_0_  ;
	output \g62014/_0_  ;
	output \g62015/_0_  ;
	output \g62016/_0_  ;
	output \g62017/_0_  ;
	output \g62018/_0_  ;
	output \g62019/_0_  ;
	output \g62020/_0_  ;
	output \g62021/_0_  ;
	output \g62022/_0_  ;
	output \g62023/_0_  ;
	output \g62024/_0_  ;
	output \g62025/_0_  ;
	output \g62026/_0_  ;
	output \g62027/_0_  ;
	output \g62030/_0_  ;
	output \g62033/_0_  ;
	output \g62034/_0_  ;
	output \g62036/_0_  ;
	output \g62038/_0_  ;
	output \g62041/_0_  ;
	output \g62042/_0_  ;
	output \g62043/_0_  ;
	output \g62044/_0_  ;
	output \g62045/_0_  ;
	output \g62046/_0_  ;
	output \g62047/_0_  ;
	output \g62048/_0_  ;
	output \g62050/_0_  ;
	output \g62051/_0_  ;
	output \g62052/_0_  ;
	output \g62055/_0_  ;
	output \g62057/_0_  ;
	output \g62058/_0_  ;
	output \g62059/_0_  ;
	output \g62060/_0_  ;
	output \g62061/_0_  ;
	output \g62062/_0_  ;
	output \g62064/_0_  ;
	output \g62065/_0_  ;
	output \g62066/_0_  ;
	output \g62067/_0_  ;
	output \g62068/_0_  ;
	output \g62072/_0_  ;
	output \g62073/_0_  ;
	output \g62074/_0_  ;
	output \g62075/_0_  ;
	output \g62076/_0_  ;
	output \g62077/_0_  ;
	output \g62078/_0_  ;
	output \g62080/_0_  ;
	output \g62081/_0_  ;
	output \g62082/_0_  ;
	output \g62084/_0_  ;
	output \g62085/_0_  ;
	output \g62086/_0_  ;
	output \g62087/_0_  ;
	output \g62088/_0_  ;
	output \g62089/_0_  ;
	output \g62090/_0_  ;
	output \g62091/_0_  ;
	output \g62092/_0_  ;
	output \g62094/_0_  ;
	output \g62096/_0_  ;
	output \g62097/_0_  ;
	output \g62098/_0_  ;
	output \g62099/_0_  ;
	output \g62100/_0_  ;
	output \g62101/_0_  ;
	output \g62102/_0_  ;
	output \g62104/_0_  ;
	output \g62106/_0_  ;
	output \g62107/_0_  ;
	output \g62108/_0_  ;
	output \g62110/_0_  ;
	output \g62112/_0_  ;
	output \g62113/_0_  ;
	output \g62114/_0_  ;
	output \g62116/_0_  ;
	output \g62117/_0_  ;
	output \g62118/_0_  ;
	output \g62119/_0_  ;
	output \g62120/_0_  ;
	output \g62121/_0_  ;
	output \g62122/_0_  ;
	output \g62124/_0_  ;
	output \g62126/_0_  ;
	output \g62127/_0_  ;
	output \g62128/_0_  ;
	output \g62129/_0_  ;
	output \g62130/_0_  ;
	output \g62131/_0_  ;
	output \g62132/_0_  ;
	output \g62133/_0_  ;
	output \g62135/_0_  ;
	output \g62136/_0_  ;
	output \g62137/_0_  ;
	output \g62138/_0_  ;
	output \g62140/_0_  ;
	output \g62143/_0_  ;
	output \g62144/_0_  ;
	output \g62149/_0_  ;
	output \g62150/_0_  ;
	output \g62151/_0_  ;
	output \g62153/_0_  ;
	output \g62155/_0_  ;
	output \g62156/_0_  ;
	output \g62158/_0_  ;
	output \g62160/_0_  ;
	output \g62161/_0_  ;
	output \g62162/_0_  ;
	output \g62164/_0_  ;
	output \g62165/_0_  ;
	output \g62166/_0_  ;
	output \g62167/_0_  ;
	output \g62168/_0_  ;
	output \g62169/_0_  ;
	output \g62172/_0_  ;
	output \g62173/_0_  ;
	output \g62175/_0_  ;
	output \g62176/_0_  ;
	output \g62177/_0_  ;
	output \g62178/_0_  ;
	output \g62179/_0_  ;
	output \g62180/_0_  ;
	output \g62181/_0_  ;
	output \g62182/_0_  ;
	output \g62183/_0_  ;
	output \g62184/_0_  ;
	output \g62185/_0_  ;
	output \g62186/_0_  ;
	output \g62188/_0_  ;
	output \g62189/_0_  ;
	output \g62190/_0_  ;
	output \g62191/_0_  ;
	output \g62193/_0_  ;
	output \g62194/_0_  ;
	output \g62195/_0_  ;
	output \g62196/_0_  ;
	output \g62197/_0_  ;
	output \g62200/_0_  ;
	output \g62201/_0_  ;
	output \g62202/_0_  ;
	output \g62203/_0_  ;
	output \g62205/_0_  ;
	output \g62206/_0_  ;
	output \g62207/_0_  ;
	output \g62208/_0_  ;
	output \g62209/_0_  ;
	output \g62210/_0_  ;
	output \g62211/_0_  ;
	output \g62215/_0_  ;
	output \g62218/_0_  ;
	output \g62219/_0_  ;
	output \g62221/_0_  ;
	output \g62222/_0_  ;
	output \g62223/_0_  ;
	output \g62224/_0_  ;
	output \g62225/_0_  ;
	output \g62226/_0_  ;
	output \g62229/_0_  ;
	output \g62230/_0_  ;
	output \g62231/_0_  ;
	output \g62233/_0_  ;
	output \g62236/_0_  ;
	output \g62237/_0_  ;
	output \g62238/_0_  ;
	output \g62240/_0_  ;
	output \g62241/_0_  ;
	output \g62243/_0_  ;
	output \g62244/_0_  ;
	output \g62245/_0_  ;
	output \g62247/_0_  ;
	output \g62248/_0_  ;
	output \g62250/_0_  ;
	output \g62252/_0_  ;
	output \g62253/_0_  ;
	output \g62255/_0_  ;
	output \g62256/_0_  ;
	output \g62257/_0_  ;
	output \g62258/_0_  ;
	output \g62259/_0_  ;
	output \g62260/_0_  ;
	output \g62261/_0_  ;
	output \g62262/_0_  ;
	output \g62263/_0_  ;
	output \g62264/_0_  ;
	output \g62265/_0_  ;
	output \g62267/_0_  ;
	output \g62269/_0_  ;
	output \g62270/_0_  ;
	output \g62272/_0_  ;
	output \g62274/_0_  ;
	output \g62277/_0_  ;
	output \g62279/_0_  ;
	output \g62280/_0_  ;
	output \g62281/_0_  ;
	output \g62283/_0_  ;
	output \g62284/_0_  ;
	output \g62285/_0_  ;
	output \g62286/_0_  ;
	output \g62288/_0_  ;
	output \g62289/_0_  ;
	output \g62290/_0_  ;
	output \g62294/_0_  ;
	output \g62295/_0_  ;
	output \g62296/_0_  ;
	output \g62297/_0_  ;
	output \g62298/_0_  ;
	output \g62299/_0_  ;
	output \g62303/_0_  ;
	output \g62305/_0_  ;
	output \g62306/_0_  ;
	output \g62307/_0_  ;
	output \g62309/_0_  ;
	output \g62311/_0_  ;
	output \g62312/_0_  ;
	output \g62313/_0_  ;
	output \g62314/_0_  ;
	output \g62315/_0_  ;
	output \g62316/_0_  ;
	output \g62317/_0_  ;
	output \g62318/_0_  ;
	output \g62319/_0_  ;
	output \g62320/_0_  ;
	output \g62322/_0_  ;
	output \g62324/_0_  ;
	output \g62325/_0_  ;
	output \g62326/_0_  ;
	output \g62327/_0_  ;
	output \g62329/_0_  ;
	output \g62330/_0_  ;
	output \g62331/_0_  ;
	output \g62332/_0_  ;
	output \g62333/_0_  ;
	output \g62335/_0_  ;
	output \g62336/_0_  ;
	output \g62338/_0_  ;
	output \g62341/_0_  ;
	output \g62342/_0_  ;
	output \g62344/_0_  ;
	output \g62345/_0_  ;
	output \g62348/_0_  ;
	output \g62349/_0_  ;
	output \g62350/_0_  ;
	output \g62353/_0_  ;
	output \g62354/_0_  ;
	output \g62355/_0_  ;
	output \g62356/_0_  ;
	output \g62359/_0_  ;
	output \g62362/_0_  ;
	output \g62363/_0_  ;
	output \g62364/_0_  ;
	output \g62365/_0_  ;
	output \g62366/_0_  ;
	output \g62367/_0_  ;
	output \g62368/_0_  ;
	output \g62369/_0_  ;
	output \g62370/_0_  ;
	output \g62371/_0_  ;
	output \g62372/_0_  ;
	output \g62373/_0_  ;
	output \g62374/_0_  ;
	output \g62376/_0_  ;
	output \g62467/_0_  ;
	output \g62468/_0_  ;
	output \g62469/_0_  ;
	output \g62470/_0_  ;
	output \g62471/_0_  ;
	output \g62472/_0_  ;
	output \g62473/_0_  ;
	output \g62474/_0_  ;
	output \g62475/_0_  ;
	output \g62478/_0_  ;
	output \g62480/_0_  ;
	output \g62481/_0_  ;
	output \g62482/_0_  ;
	output \g62483/_0_  ;
	output \g62484/_0_  ;
	output \g62485/_0_  ;
	output \g62486/_0_  ;
	output \g62487/_0_  ;
	output \g62488/_0_  ;
	output \g62489/_0_  ;
	output \g62490/_0_  ;
	output \g62491/_0_  ;
	output \g62492/_0_  ;
	output \g62493/_0_  ;
	output \g62494/_0_  ;
	output \g62495/_0_  ;
	output \g62496/_0_  ;
	output \g62497/_0_  ;
	output \g62498/_0_  ;
	output \g62499/_0_  ;
	output \g62500/_0_  ;
	output \g62501/_0_  ;
	output \g62502/_0_  ;
	output \g62503/_0_  ;
	output \g62504/_0_  ;
	output \g62509/_0_  ;
	output \g62510/_0_  ;
	output \g62511/_0_  ;
	output \g62512/_0_  ;
	output \g62513/_0_  ;
	output \g62514/_0_  ;
	output \g62515/_0_  ;
	output \g62516/_0_  ;
	output \g62517/_0_  ;
	output \g62518/_0_  ;
	output \g62519/_0_  ;
	output \g62520/_0_  ;
	output \g62521/_0_  ;
	output \g62523/_0_  ;
	output \g62526/_0_  ;
	output \g62528/_0_  ;
	output \g62529/_0_  ;
	output \g62531/_0_  ;
	output \g62532/_0_  ;
	output \g62533/_0_  ;
	output \g62534/_0_  ;
	output \g62535/_0_  ;
	output \g62536/_0_  ;
	output \g62537/_0_  ;
	output \g62539/_0_  ;
	output \g62540/_0_  ;
	output \g62541/_0_  ;
	output \g62542/_0_  ;
	output \g62543/_0_  ;
	output \g62544/_0_  ;
	output \g62545/_0_  ;
	output \g62547/_0_  ;
	output \g62548/_0_  ;
	output \g62549/_0_  ;
	output \g62550/_0_  ;
	output \g62551/_0_  ;
	output \g62552/_0_  ;
	output \g62553/_0_  ;
	output \g62554/_0_  ;
	output \g62555/_0_  ;
	output \g62556/_0_  ;
	output \g62557/_0_  ;
	output \g62560/_0_  ;
	output \g62562/_0_  ;
	output \g62563/_0_  ;
	output \g62564/_0_  ;
	output \g62565/_0_  ;
	output \g62566/_0_  ;
	output \g62567/_0_  ;
	output \g62569/_0_  ;
	output \g62570/_0_  ;
	output \g62571/_0_  ;
	output \g62572/_0_  ;
	output \g62573/_0_  ;
	output \g62574/_0_  ;
	output \g62576/_0_  ;
	output \g62577/_0_  ;
	output \g62581/_0_  ;
	output \g62582/_0_  ;
	output \g62584/_0_  ;
	output \g62585/_0_  ;
	output \g62586/_0_  ;
	output \g62588/_0_  ;
	output \g62589/_0_  ;
	output \g62593/_0_  ;
	output \g62594/_0_  ;
	output \g62595/_0_  ;
	output \g62596/_0_  ;
	output \g62597/_0_  ;
	output \g62598/_0_  ;
	output \g62599/_0_  ;
	output \g62600/_0_  ;
	output \g62601/_0_  ;
	output \g62602/_0_  ;
	output \g62603/_0_  ;
	output \g62604/_0_  ;
	output \g62605/_0_  ;
	output \g62606/_0_  ;
	output \g62607/_0_  ;
	output \g62608/_0_  ;
	output \g62609/_0_  ;
	output \g62610/_0_  ;
	output \g62612/_0_  ;
	output \g62613/_0_  ;
	output \g62614/_0_  ;
	output \g62615/_0_  ;
	output \g62617/_0_  ;
	output \g62618/_0_  ;
	output \g62620/_0_  ;
	output \g62621/_0_  ;
	output \g62622/_0_  ;
	output \g62624/_0_  ;
	output \g62625/_0_  ;
	output \g62626/_0_  ;
	output \g62627/_0_  ;
	output \g62629/_0_  ;
	output \g62630/_0_  ;
	output \g62632/_0_  ;
	output \g62633/_0_  ;
	output \g62635/_0_  ;
	output \g62636/_0_  ;
	output \g62637/_0_  ;
	output \g62638/_0_  ;
	output \g62640/_0_  ;
	output \g62641/_0_  ;
	output \g62642/_0_  ;
	output \g62643/_0_  ;
	output \g62644/_0_  ;
	output \g62646/_0_  ;
	output \g62647/_0_  ;
	output \g62649/_0_  ;
	output \g62650/_0_  ;
	output \g62651/_0_  ;
	output \g62653/_0_  ;
	output \g62655/_0_  ;
	output \g62656/_0_  ;
	output \g62657/_0_  ;
	output \g62658/_0_  ;
	output \g62660/_0_  ;
	output \g62661/_0_  ;
	output \g62662/_0_  ;
	output \g62663/_0_  ;
	output \g62664/_0_  ;
	output \g62665/_0_  ;
	output \g62667/_0_  ;
	output \g62669/_0_  ;
	output \g62670/_0_  ;
	output \g62671/_0_  ;
	output \g62672/_0_  ;
	output \g62674/_0_  ;
	output \g62675/_0_  ;
	output \g62676/_0_  ;
	output \g62677/_0_  ;
	output \g62678/_0_  ;
	output \g62679/_0_  ;
	output \g62680/_0_  ;
	output \g62681/_0_  ;
	output \g62682/_0_  ;
	output \g62684/_0_  ;
	output \g62685/_0_  ;
	output \g62686/_0_  ;
	output \g62687/_0_  ;
	output \g62690/_0_  ;
	output \g62693/_0_  ;
	output \g62698/_0_  ;
	output \g62699/_0_  ;
	output \g62700/_0_  ;
	output \g62701/_0_  ;
	output \g62702/_0_  ;
	output \g62703/_0_  ;
	output \g62704/_0_  ;
	output \g62709/_0_  ;
	output \g62710/_0_  ;
	output \g62711/_0_  ;
	output \g62714/_0_  ;
	output \g62715/_0_  ;
	output \g62717/_0_  ;
	output \g62718/_0_  ;
	output \g62719/_0_  ;
	output \g62720/_0_  ;
	output \g62721/_0_  ;
	output \g62723/_0_  ;
	output \g62725/_0_  ;
	output \g62726/_0_  ;
	output \g62729/_0_  ;
	output \g62731/_0_  ;
	output \g62733/_0_  ;
	output \g62738/_0_  ;
	output \g62741/_0_  ;
	output \g62742/_0_  ;
	output \g62744/_0_  ;
	output \g62745/_0_  ;
	output \g62746/_0_  ;
	output \g62747/_0_  ;
	output \g62748/_0_  ;
	output \g62749/_0_  ;
	output \g62753/_0_  ;
	output \g62755/_0_  ;
	output \g62756/_0_  ;
	output \g62758/_0_  ;
	output \g62759/_0_  ;
	output \g62760/_0_  ;
	output \g62761/_0_  ;
	output \g62763/_0_  ;
	output \g62766/_0_  ;
	output \g62767/_0_  ;
	output \g62768/_0_  ;
	output \g65554/_0_  ;
	output \g65561/_0_  ;
	output \g65569/_0_  ;
	output \g65580/_0_  ;
	output \g65599/_0_  ;
	output \g65606/_0_  ;
	output \g65636/_0_  ;
	output \g65864/_0_  ;
	wire _w8710_ ;
	wire _w8709_ ;
	wire _w8708_ ;
	wire _w8707_ ;
	wire _w8706_ ;
	wire _w8705_ ;
	wire _w8704_ ;
	wire _w8703_ ;
	wire _w8702_ ;
	wire _w8701_ ;
	wire _w8700_ ;
	wire _w8699_ ;
	wire _w8698_ ;
	wire _w8697_ ;
	wire _w8696_ ;
	wire _w8695_ ;
	wire _w8694_ ;
	wire _w8693_ ;
	wire _w8692_ ;
	wire _w8691_ ;
	wire _w8690_ ;
	wire _w8689_ ;
	wire _w8688_ ;
	wire _w8687_ ;
	wire _w8686_ ;
	wire _w8685_ ;
	wire _w8684_ ;
	wire _w8683_ ;
	wire _w8682_ ;
	wire _w8681_ ;
	wire _w8680_ ;
	wire _w8679_ ;
	wire _w8678_ ;
	wire _w8677_ ;
	wire _w8676_ ;
	wire _w8675_ ;
	wire _w8674_ ;
	wire _w8673_ ;
	wire _w8672_ ;
	wire _w8671_ ;
	wire _w8670_ ;
	wire _w8669_ ;
	wire _w8668_ ;
	wire _w8667_ ;
	wire _w8666_ ;
	wire _w8665_ ;
	wire _w8664_ ;
	wire _w8663_ ;
	wire _w8662_ ;
	wire _w8661_ ;
	wire _w8660_ ;
	wire _w8659_ ;
	wire _w8658_ ;
	wire _w8657_ ;
	wire _w8656_ ;
	wire _w8655_ ;
	wire _w8654_ ;
	wire _w8653_ ;
	wire _w8652_ ;
	wire _w8651_ ;
	wire _w8650_ ;
	wire _w8649_ ;
	wire _w8648_ ;
	wire _w8647_ ;
	wire _w8646_ ;
	wire _w8645_ ;
	wire _w8644_ ;
	wire _w8643_ ;
	wire _w8642_ ;
	wire _w8641_ ;
	wire _w8640_ ;
	wire _w8639_ ;
	wire _w8638_ ;
	wire _w8637_ ;
	wire _w8636_ ;
	wire _w8635_ ;
	wire _w8634_ ;
	wire _w8633_ ;
	wire _w8632_ ;
	wire _w8631_ ;
	wire _w8630_ ;
	wire _w8629_ ;
	wire _w8628_ ;
	wire _w8627_ ;
	wire _w8626_ ;
	wire _w8625_ ;
	wire _w8624_ ;
	wire _w8623_ ;
	wire _w8622_ ;
	wire _w8621_ ;
	wire _w8620_ ;
	wire _w8619_ ;
	wire _w8618_ ;
	wire _w8617_ ;
	wire _w8616_ ;
	wire _w8615_ ;
	wire _w8614_ ;
	wire _w8613_ ;
	wire _w8612_ ;
	wire _w8611_ ;
	wire _w8610_ ;
	wire _w8609_ ;
	wire _w8608_ ;
	wire _w8607_ ;
	wire _w8606_ ;
	wire _w8605_ ;
	wire _w8604_ ;
	wire _w8603_ ;
	wire _w8602_ ;
	wire _w8601_ ;
	wire _w8600_ ;
	wire _w8599_ ;
	wire _w8598_ ;
	wire _w8597_ ;
	wire _w8596_ ;
	wire _w8595_ ;
	wire _w8594_ ;
	wire _w8593_ ;
	wire _w8592_ ;
	wire _w8591_ ;
	wire _w8590_ ;
	wire _w8589_ ;
	wire _w8588_ ;
	wire _w8587_ ;
	wire _w8586_ ;
	wire _w8585_ ;
	wire _w8584_ ;
	wire _w8583_ ;
	wire _w8582_ ;
	wire _w8581_ ;
	wire _w8580_ ;
	wire _w8579_ ;
	wire _w8578_ ;
	wire _w8577_ ;
	wire _w8576_ ;
	wire _w8575_ ;
	wire _w8574_ ;
	wire _w8573_ ;
	wire _w8572_ ;
	wire _w8571_ ;
	wire _w8570_ ;
	wire _w8569_ ;
	wire _w8568_ ;
	wire _w8567_ ;
	wire _w8566_ ;
	wire _w8565_ ;
	wire _w8564_ ;
	wire _w8563_ ;
	wire _w8562_ ;
	wire _w8561_ ;
	wire _w8560_ ;
	wire _w8559_ ;
	wire _w8558_ ;
	wire _w8557_ ;
	wire _w8556_ ;
	wire _w8555_ ;
	wire _w8554_ ;
	wire _w8553_ ;
	wire _w8552_ ;
	wire _w8551_ ;
	wire _w8550_ ;
	wire _w8549_ ;
	wire _w8548_ ;
	wire _w8547_ ;
	wire _w8546_ ;
	wire _w8545_ ;
	wire _w8544_ ;
	wire _w8543_ ;
	wire _w8542_ ;
	wire _w8541_ ;
	wire _w8540_ ;
	wire _w8539_ ;
	wire _w8538_ ;
	wire _w8537_ ;
	wire _w8536_ ;
	wire _w8535_ ;
	wire _w8534_ ;
	wire _w8533_ ;
	wire _w8532_ ;
	wire _w8531_ ;
	wire _w8530_ ;
	wire _w8529_ ;
	wire _w8528_ ;
	wire _w8527_ ;
	wire _w8526_ ;
	wire _w8525_ ;
	wire _w8524_ ;
	wire _w8523_ ;
	wire _w8522_ ;
	wire _w8521_ ;
	wire _w8520_ ;
	wire _w8519_ ;
	wire _w8518_ ;
	wire _w8517_ ;
	wire _w8516_ ;
	wire _w8515_ ;
	wire _w8514_ ;
	wire _w8513_ ;
	wire _w8512_ ;
	wire _w8511_ ;
	wire _w8510_ ;
	wire _w8509_ ;
	wire _w8508_ ;
	wire _w8507_ ;
	wire _w8506_ ;
	wire _w8505_ ;
	wire _w8504_ ;
	wire _w8503_ ;
	wire _w8502_ ;
	wire _w8501_ ;
	wire _w8500_ ;
	wire _w8499_ ;
	wire _w8498_ ;
	wire _w8497_ ;
	wire _w8496_ ;
	wire _w8495_ ;
	wire _w8494_ ;
	wire _w8493_ ;
	wire _w8492_ ;
	wire _w8491_ ;
	wire _w8490_ ;
	wire _w8489_ ;
	wire _w8488_ ;
	wire _w8487_ ;
	wire _w8486_ ;
	wire _w8485_ ;
	wire _w8484_ ;
	wire _w8483_ ;
	wire _w8482_ ;
	wire _w8481_ ;
	wire _w8480_ ;
	wire _w8479_ ;
	wire _w8478_ ;
	wire _w8477_ ;
	wire _w8476_ ;
	wire _w8475_ ;
	wire _w8474_ ;
	wire _w8473_ ;
	wire _w8472_ ;
	wire _w8471_ ;
	wire _w8470_ ;
	wire _w8469_ ;
	wire _w8468_ ;
	wire _w8467_ ;
	wire _w8466_ ;
	wire _w8465_ ;
	wire _w8464_ ;
	wire _w8463_ ;
	wire _w8462_ ;
	wire _w8461_ ;
	wire _w8460_ ;
	wire _w8459_ ;
	wire _w8458_ ;
	wire _w8457_ ;
	wire _w8456_ ;
	wire _w8455_ ;
	wire _w8454_ ;
	wire _w8453_ ;
	wire _w8452_ ;
	wire _w8451_ ;
	wire _w8450_ ;
	wire _w8449_ ;
	wire _w8448_ ;
	wire _w8447_ ;
	wire _w8446_ ;
	wire _w8445_ ;
	wire _w8444_ ;
	wire _w8443_ ;
	wire _w8442_ ;
	wire _w8441_ ;
	wire _w8440_ ;
	wire _w8439_ ;
	wire _w8438_ ;
	wire _w8437_ ;
	wire _w8436_ ;
	wire _w8435_ ;
	wire _w8434_ ;
	wire _w8433_ ;
	wire _w8432_ ;
	wire _w8431_ ;
	wire _w8430_ ;
	wire _w8429_ ;
	wire _w8428_ ;
	wire _w8427_ ;
	wire _w8426_ ;
	wire _w8425_ ;
	wire _w8424_ ;
	wire _w8423_ ;
	wire _w8422_ ;
	wire _w8421_ ;
	wire _w8420_ ;
	wire _w8419_ ;
	wire _w8418_ ;
	wire _w8417_ ;
	wire _w8416_ ;
	wire _w8415_ ;
	wire _w8414_ ;
	wire _w8413_ ;
	wire _w8412_ ;
	wire _w8411_ ;
	wire _w8410_ ;
	wire _w8409_ ;
	wire _w8408_ ;
	wire _w8407_ ;
	wire _w8406_ ;
	wire _w8405_ ;
	wire _w8404_ ;
	wire _w8403_ ;
	wire _w8402_ ;
	wire _w8401_ ;
	wire _w8400_ ;
	wire _w8399_ ;
	wire _w8398_ ;
	wire _w8397_ ;
	wire _w8396_ ;
	wire _w8395_ ;
	wire _w8394_ ;
	wire _w8393_ ;
	wire _w8392_ ;
	wire _w8391_ ;
	wire _w8390_ ;
	wire _w8389_ ;
	wire _w8388_ ;
	wire _w8387_ ;
	wire _w8386_ ;
	wire _w8385_ ;
	wire _w8384_ ;
	wire _w8383_ ;
	wire _w8382_ ;
	wire _w8381_ ;
	wire _w8380_ ;
	wire _w8379_ ;
	wire _w8378_ ;
	wire _w8377_ ;
	wire _w8376_ ;
	wire _w8375_ ;
	wire _w8374_ ;
	wire _w8373_ ;
	wire _w8372_ ;
	wire _w8371_ ;
	wire _w8370_ ;
	wire _w8369_ ;
	wire _w8368_ ;
	wire _w8367_ ;
	wire _w8366_ ;
	wire _w8365_ ;
	wire _w8364_ ;
	wire _w8363_ ;
	wire _w8362_ ;
	wire _w8361_ ;
	wire _w8360_ ;
	wire _w8359_ ;
	wire _w8358_ ;
	wire _w8357_ ;
	wire _w8356_ ;
	wire _w8355_ ;
	wire _w8354_ ;
	wire _w8353_ ;
	wire _w8352_ ;
	wire _w8351_ ;
	wire _w8350_ ;
	wire _w8349_ ;
	wire _w8348_ ;
	wire _w8347_ ;
	wire _w8346_ ;
	wire _w8345_ ;
	wire _w8344_ ;
	wire _w8343_ ;
	wire _w8342_ ;
	wire _w8341_ ;
	wire _w8340_ ;
	wire _w8339_ ;
	wire _w8338_ ;
	wire _w8337_ ;
	wire _w8336_ ;
	wire _w8335_ ;
	wire _w8334_ ;
	wire _w8333_ ;
	wire _w8332_ ;
	wire _w8331_ ;
	wire _w8330_ ;
	wire _w8329_ ;
	wire _w8328_ ;
	wire _w8327_ ;
	wire _w8326_ ;
	wire _w8325_ ;
	wire _w8324_ ;
	wire _w8323_ ;
	wire _w8322_ ;
	wire _w8321_ ;
	wire _w8320_ ;
	wire _w8319_ ;
	wire _w8318_ ;
	wire _w8317_ ;
	wire _w8316_ ;
	wire _w8315_ ;
	wire _w8314_ ;
	wire _w8313_ ;
	wire _w8312_ ;
	wire _w8311_ ;
	wire _w8310_ ;
	wire _w8309_ ;
	wire _w8308_ ;
	wire _w8307_ ;
	wire _w8306_ ;
	wire _w8305_ ;
	wire _w8304_ ;
	wire _w8303_ ;
	wire _w8302_ ;
	wire _w8301_ ;
	wire _w8300_ ;
	wire _w8299_ ;
	wire _w8298_ ;
	wire _w8297_ ;
	wire _w8296_ ;
	wire _w8295_ ;
	wire _w8294_ ;
	wire _w8293_ ;
	wire _w8292_ ;
	wire _w8291_ ;
	wire _w8290_ ;
	wire _w8289_ ;
	wire _w8288_ ;
	wire _w8287_ ;
	wire _w8286_ ;
	wire _w8285_ ;
	wire _w8284_ ;
	wire _w8283_ ;
	wire _w8282_ ;
	wire _w8281_ ;
	wire _w8280_ ;
	wire _w8279_ ;
	wire _w8278_ ;
	wire _w8277_ ;
	wire _w8276_ ;
	wire _w8275_ ;
	wire _w8274_ ;
	wire _w8273_ ;
	wire _w8272_ ;
	wire _w8271_ ;
	wire _w8270_ ;
	wire _w8269_ ;
	wire _w8268_ ;
	wire _w8267_ ;
	wire _w8266_ ;
	wire _w8265_ ;
	wire _w8264_ ;
	wire _w8263_ ;
	wire _w8262_ ;
	wire _w8261_ ;
	wire _w8260_ ;
	wire _w8259_ ;
	wire _w8258_ ;
	wire _w8257_ ;
	wire _w8256_ ;
	wire _w8255_ ;
	wire _w8254_ ;
	wire _w8253_ ;
	wire _w8252_ ;
	wire _w8251_ ;
	wire _w8250_ ;
	wire _w8249_ ;
	wire _w8248_ ;
	wire _w8247_ ;
	wire _w8246_ ;
	wire _w8245_ ;
	wire _w8244_ ;
	wire _w8243_ ;
	wire _w8242_ ;
	wire _w8241_ ;
	wire _w8240_ ;
	wire _w8239_ ;
	wire _w8238_ ;
	wire _w8237_ ;
	wire _w8236_ ;
	wire _w8235_ ;
	wire _w8234_ ;
	wire _w8233_ ;
	wire _w8232_ ;
	wire _w8231_ ;
	wire _w8230_ ;
	wire _w8229_ ;
	wire _w8228_ ;
	wire _w8227_ ;
	wire _w8226_ ;
	wire _w8225_ ;
	wire _w8224_ ;
	wire _w8223_ ;
	wire _w8222_ ;
	wire _w8221_ ;
	wire _w8220_ ;
	wire _w8219_ ;
	wire _w8218_ ;
	wire _w8217_ ;
	wire _w8216_ ;
	wire _w8215_ ;
	wire _w8214_ ;
	wire _w8213_ ;
	wire _w8212_ ;
	wire _w8211_ ;
	wire _w8210_ ;
	wire _w8209_ ;
	wire _w8208_ ;
	wire _w8207_ ;
	wire _w8206_ ;
	wire _w8205_ ;
	wire _w8204_ ;
	wire _w8203_ ;
	wire _w8202_ ;
	wire _w8201_ ;
	wire _w8200_ ;
	wire _w8199_ ;
	wire _w8198_ ;
	wire _w8197_ ;
	wire _w8196_ ;
	wire _w8195_ ;
	wire _w8194_ ;
	wire _w8193_ ;
	wire _w8192_ ;
	wire _w8191_ ;
	wire _w8190_ ;
	wire _w8189_ ;
	wire _w8188_ ;
	wire _w8187_ ;
	wire _w8186_ ;
	wire _w8185_ ;
	wire _w8184_ ;
	wire _w8183_ ;
	wire _w8182_ ;
	wire _w8181_ ;
	wire _w8180_ ;
	wire _w8179_ ;
	wire _w8178_ ;
	wire _w8177_ ;
	wire _w8176_ ;
	wire _w8175_ ;
	wire _w8174_ ;
	wire _w8173_ ;
	wire _w8172_ ;
	wire _w8171_ ;
	wire _w8170_ ;
	wire _w8169_ ;
	wire _w8168_ ;
	wire _w8167_ ;
	wire _w8166_ ;
	wire _w8165_ ;
	wire _w8164_ ;
	wire _w8163_ ;
	wire _w8162_ ;
	wire _w8161_ ;
	wire _w8160_ ;
	wire _w8159_ ;
	wire _w8158_ ;
	wire _w8157_ ;
	wire _w8156_ ;
	wire _w8155_ ;
	wire _w8154_ ;
	wire _w8153_ ;
	wire _w8152_ ;
	wire _w8151_ ;
	wire _w8150_ ;
	wire _w8149_ ;
	wire _w8148_ ;
	wire _w8147_ ;
	wire _w8146_ ;
	wire _w8145_ ;
	wire _w8144_ ;
	wire _w8143_ ;
	wire _w8142_ ;
	wire _w8141_ ;
	wire _w8140_ ;
	wire _w8139_ ;
	wire _w8138_ ;
	wire _w8137_ ;
	wire _w8136_ ;
	wire _w8135_ ;
	wire _w8134_ ;
	wire _w8133_ ;
	wire _w8132_ ;
	wire _w8131_ ;
	wire _w8130_ ;
	wire _w8129_ ;
	wire _w8128_ ;
	wire _w8127_ ;
	wire _w8126_ ;
	wire _w8125_ ;
	wire _w8124_ ;
	wire _w8123_ ;
	wire _w8122_ ;
	wire _w8121_ ;
	wire _w8120_ ;
	wire _w8119_ ;
	wire _w8118_ ;
	wire _w8117_ ;
	wire _w8116_ ;
	wire _w8115_ ;
	wire _w8114_ ;
	wire _w8113_ ;
	wire _w8112_ ;
	wire _w8111_ ;
	wire _w8110_ ;
	wire _w8109_ ;
	wire _w8108_ ;
	wire _w8107_ ;
	wire _w8106_ ;
	wire _w8105_ ;
	wire _w8104_ ;
	wire _w8103_ ;
	wire _w8102_ ;
	wire _w8101_ ;
	wire _w8100_ ;
	wire _w8099_ ;
	wire _w8098_ ;
	wire _w8097_ ;
	wire _w8096_ ;
	wire _w8095_ ;
	wire _w8094_ ;
	wire _w8093_ ;
	wire _w8092_ ;
	wire _w8091_ ;
	wire _w8090_ ;
	wire _w8089_ ;
	wire _w8088_ ;
	wire _w8087_ ;
	wire _w8086_ ;
	wire _w8085_ ;
	wire _w8084_ ;
	wire _w8083_ ;
	wire _w8082_ ;
	wire _w8081_ ;
	wire _w8080_ ;
	wire _w8079_ ;
	wire _w8078_ ;
	wire _w8077_ ;
	wire _w8076_ ;
	wire _w8075_ ;
	wire _w8074_ ;
	wire _w8073_ ;
	wire _w8072_ ;
	wire _w8071_ ;
	wire _w8070_ ;
	wire _w8069_ ;
	wire _w8068_ ;
	wire _w8067_ ;
	wire _w8066_ ;
	wire _w8065_ ;
	wire _w8064_ ;
	wire _w8063_ ;
	wire _w8062_ ;
	wire _w8061_ ;
	wire _w8060_ ;
	wire _w8059_ ;
	wire _w8058_ ;
	wire _w8057_ ;
	wire _w8056_ ;
	wire _w8055_ ;
	wire _w8054_ ;
	wire _w8053_ ;
	wire _w8052_ ;
	wire _w8051_ ;
	wire _w8050_ ;
	wire _w8049_ ;
	wire _w8048_ ;
	wire _w8047_ ;
	wire _w8046_ ;
	wire _w8045_ ;
	wire _w8044_ ;
	wire _w8043_ ;
	wire _w8042_ ;
	wire _w8041_ ;
	wire _w8040_ ;
	wire _w8039_ ;
	wire _w8038_ ;
	wire _w8037_ ;
	wire _w8036_ ;
	wire _w8035_ ;
	wire _w8034_ ;
	wire _w8033_ ;
	wire _w8032_ ;
	wire _w8031_ ;
	wire _w8030_ ;
	wire _w8029_ ;
	wire _w8028_ ;
	wire _w8027_ ;
	wire _w8026_ ;
	wire _w8025_ ;
	wire _w8024_ ;
	wire _w8023_ ;
	wire _w8022_ ;
	wire _w8021_ ;
	wire _w8020_ ;
	wire _w8019_ ;
	wire _w8018_ ;
	wire _w8017_ ;
	wire _w8016_ ;
	wire _w8015_ ;
	wire _w8014_ ;
	wire _w8013_ ;
	wire _w8012_ ;
	wire _w8011_ ;
	wire _w8010_ ;
	wire _w8009_ ;
	wire _w8008_ ;
	wire _w8007_ ;
	wire _w8006_ ;
	wire _w8005_ ;
	wire _w8004_ ;
	wire _w8003_ ;
	wire _w8002_ ;
	wire _w8001_ ;
	wire _w8000_ ;
	wire _w7999_ ;
	wire _w7998_ ;
	wire _w7997_ ;
	wire _w7996_ ;
	wire _w7995_ ;
	wire _w7994_ ;
	wire _w7993_ ;
	wire _w7992_ ;
	wire _w7991_ ;
	wire _w7990_ ;
	wire _w7989_ ;
	wire _w7988_ ;
	wire _w7987_ ;
	wire _w7986_ ;
	wire _w7985_ ;
	wire _w7984_ ;
	wire _w7983_ ;
	wire _w7982_ ;
	wire _w7981_ ;
	wire _w7980_ ;
	wire _w7979_ ;
	wire _w7978_ ;
	wire _w7977_ ;
	wire _w7976_ ;
	wire _w7975_ ;
	wire _w7974_ ;
	wire _w7973_ ;
	wire _w7972_ ;
	wire _w7971_ ;
	wire _w7970_ ;
	wire _w7969_ ;
	wire _w7968_ ;
	wire _w7967_ ;
	wire _w7966_ ;
	wire _w7965_ ;
	wire _w7964_ ;
	wire _w7963_ ;
	wire _w7962_ ;
	wire _w7961_ ;
	wire _w7960_ ;
	wire _w7959_ ;
	wire _w7958_ ;
	wire _w7957_ ;
	wire _w7956_ ;
	wire _w7955_ ;
	wire _w7954_ ;
	wire _w7953_ ;
	wire _w7952_ ;
	wire _w7951_ ;
	wire _w7950_ ;
	wire _w7949_ ;
	wire _w7948_ ;
	wire _w7947_ ;
	wire _w7946_ ;
	wire _w7945_ ;
	wire _w7944_ ;
	wire _w7943_ ;
	wire _w7942_ ;
	wire _w7941_ ;
	wire _w7940_ ;
	wire _w7939_ ;
	wire _w7938_ ;
	wire _w7937_ ;
	wire _w7936_ ;
	wire _w7935_ ;
	wire _w7934_ ;
	wire _w7933_ ;
	wire _w7932_ ;
	wire _w7931_ ;
	wire _w7930_ ;
	wire _w7929_ ;
	wire _w7928_ ;
	wire _w7927_ ;
	wire _w7926_ ;
	wire _w7925_ ;
	wire _w7924_ ;
	wire _w7923_ ;
	wire _w7922_ ;
	wire _w7921_ ;
	wire _w7920_ ;
	wire _w7919_ ;
	wire _w7918_ ;
	wire _w7917_ ;
	wire _w7916_ ;
	wire _w7915_ ;
	wire _w7914_ ;
	wire _w7913_ ;
	wire _w7912_ ;
	wire _w7911_ ;
	wire _w7910_ ;
	wire _w7909_ ;
	wire _w7908_ ;
	wire _w7907_ ;
	wire _w7906_ ;
	wire _w7905_ ;
	wire _w7904_ ;
	wire _w7903_ ;
	wire _w7902_ ;
	wire _w7901_ ;
	wire _w7900_ ;
	wire _w7899_ ;
	wire _w7898_ ;
	wire _w7897_ ;
	wire _w7896_ ;
	wire _w7895_ ;
	wire _w7894_ ;
	wire _w7893_ ;
	wire _w7892_ ;
	wire _w7891_ ;
	wire _w7890_ ;
	wire _w7889_ ;
	wire _w7888_ ;
	wire _w7887_ ;
	wire _w7886_ ;
	wire _w7885_ ;
	wire _w7884_ ;
	wire _w7883_ ;
	wire _w7882_ ;
	wire _w7881_ ;
	wire _w7880_ ;
	wire _w7879_ ;
	wire _w7878_ ;
	wire _w7877_ ;
	wire _w7876_ ;
	wire _w7875_ ;
	wire _w7874_ ;
	wire _w7873_ ;
	wire _w7872_ ;
	wire _w7871_ ;
	wire _w7870_ ;
	wire _w7869_ ;
	wire _w7868_ ;
	wire _w7867_ ;
	wire _w7866_ ;
	wire _w7865_ ;
	wire _w7864_ ;
	wire _w7863_ ;
	wire _w7862_ ;
	wire _w7861_ ;
	wire _w7860_ ;
	wire _w7859_ ;
	wire _w7858_ ;
	wire _w7857_ ;
	wire _w7856_ ;
	wire _w7855_ ;
	wire _w7854_ ;
	wire _w7853_ ;
	wire _w7852_ ;
	wire _w7851_ ;
	wire _w7850_ ;
	wire _w7849_ ;
	wire _w7848_ ;
	wire _w7847_ ;
	wire _w7846_ ;
	wire _w7845_ ;
	wire _w7844_ ;
	wire _w7843_ ;
	wire _w7842_ ;
	wire _w7841_ ;
	wire _w7840_ ;
	wire _w7839_ ;
	wire _w7838_ ;
	wire _w7837_ ;
	wire _w7836_ ;
	wire _w7835_ ;
	wire _w7834_ ;
	wire _w7833_ ;
	wire _w7832_ ;
	wire _w7831_ ;
	wire _w7830_ ;
	wire _w7829_ ;
	wire _w7828_ ;
	wire _w7827_ ;
	wire _w7826_ ;
	wire _w7825_ ;
	wire _w7824_ ;
	wire _w7823_ ;
	wire _w7822_ ;
	wire _w7821_ ;
	wire _w7820_ ;
	wire _w7819_ ;
	wire _w7818_ ;
	wire _w7817_ ;
	wire _w7816_ ;
	wire _w7815_ ;
	wire _w7814_ ;
	wire _w7813_ ;
	wire _w7812_ ;
	wire _w7811_ ;
	wire _w7810_ ;
	wire _w7809_ ;
	wire _w7808_ ;
	wire _w7807_ ;
	wire _w7806_ ;
	wire _w7805_ ;
	wire _w7804_ ;
	wire _w7803_ ;
	wire _w7802_ ;
	wire _w7801_ ;
	wire _w7800_ ;
	wire _w7799_ ;
	wire _w7798_ ;
	wire _w7797_ ;
	wire _w7796_ ;
	wire _w7795_ ;
	wire _w7794_ ;
	wire _w7793_ ;
	wire _w7792_ ;
	wire _w7791_ ;
	wire _w7790_ ;
	wire _w7789_ ;
	wire _w7788_ ;
	wire _w7787_ ;
	wire _w7786_ ;
	wire _w7785_ ;
	wire _w7784_ ;
	wire _w7783_ ;
	wire _w7782_ ;
	wire _w7781_ ;
	wire _w7780_ ;
	wire _w7779_ ;
	wire _w7778_ ;
	wire _w7777_ ;
	wire _w7776_ ;
	wire _w7775_ ;
	wire _w7774_ ;
	wire _w7773_ ;
	wire _w7772_ ;
	wire _w7771_ ;
	wire _w7770_ ;
	wire _w7769_ ;
	wire _w7768_ ;
	wire _w7767_ ;
	wire _w7766_ ;
	wire _w7765_ ;
	wire _w7764_ ;
	wire _w7763_ ;
	wire _w7762_ ;
	wire _w7761_ ;
	wire _w7760_ ;
	wire _w7759_ ;
	wire _w7758_ ;
	wire _w7757_ ;
	wire _w7756_ ;
	wire _w7755_ ;
	wire _w7754_ ;
	wire _w7753_ ;
	wire _w7752_ ;
	wire _w7751_ ;
	wire _w7750_ ;
	wire _w7749_ ;
	wire _w7748_ ;
	wire _w7747_ ;
	wire _w7746_ ;
	wire _w7745_ ;
	wire _w7744_ ;
	wire _w7743_ ;
	wire _w7742_ ;
	wire _w7741_ ;
	wire _w7740_ ;
	wire _w7739_ ;
	wire _w7738_ ;
	wire _w7737_ ;
	wire _w7736_ ;
	wire _w7735_ ;
	wire _w7734_ ;
	wire _w7733_ ;
	wire _w7732_ ;
	wire _w7731_ ;
	wire _w7730_ ;
	wire _w7729_ ;
	wire _w7728_ ;
	wire _w7727_ ;
	wire _w7726_ ;
	wire _w7725_ ;
	wire _w7724_ ;
	wire _w7723_ ;
	wire _w7722_ ;
	wire _w7721_ ;
	wire _w7720_ ;
	wire _w7719_ ;
	wire _w7718_ ;
	wire _w7717_ ;
	wire _w7716_ ;
	wire _w7715_ ;
	wire _w7714_ ;
	wire _w7713_ ;
	wire _w7712_ ;
	wire _w7711_ ;
	wire _w7710_ ;
	wire _w7709_ ;
	wire _w7708_ ;
	wire _w7707_ ;
	wire _w7706_ ;
	wire _w7705_ ;
	wire _w7704_ ;
	wire _w7703_ ;
	wire _w7702_ ;
	wire _w7701_ ;
	wire _w7700_ ;
	wire _w7699_ ;
	wire _w7698_ ;
	wire _w7697_ ;
	wire _w7696_ ;
	wire _w7695_ ;
	wire _w7694_ ;
	wire _w7693_ ;
	wire _w7692_ ;
	wire _w7691_ ;
	wire _w7690_ ;
	wire _w7689_ ;
	wire _w7688_ ;
	wire _w7687_ ;
	wire _w7686_ ;
	wire _w7685_ ;
	wire _w7684_ ;
	wire _w7683_ ;
	wire _w7682_ ;
	wire _w7681_ ;
	wire _w7680_ ;
	wire _w7679_ ;
	wire _w7678_ ;
	wire _w7677_ ;
	wire _w7676_ ;
	wire _w7675_ ;
	wire _w7674_ ;
	wire _w7673_ ;
	wire _w7672_ ;
	wire _w7671_ ;
	wire _w7670_ ;
	wire _w7669_ ;
	wire _w7668_ ;
	wire _w7667_ ;
	wire _w7666_ ;
	wire _w7665_ ;
	wire _w7664_ ;
	wire _w7663_ ;
	wire _w7662_ ;
	wire _w7661_ ;
	wire _w7660_ ;
	wire _w7659_ ;
	wire _w7658_ ;
	wire _w7657_ ;
	wire _w7656_ ;
	wire _w7655_ ;
	wire _w7654_ ;
	wire _w7653_ ;
	wire _w7652_ ;
	wire _w7651_ ;
	wire _w7650_ ;
	wire _w7649_ ;
	wire _w7648_ ;
	wire _w7647_ ;
	wire _w7646_ ;
	wire _w7645_ ;
	wire _w7644_ ;
	wire _w7643_ ;
	wire _w7642_ ;
	wire _w7641_ ;
	wire _w7640_ ;
	wire _w7639_ ;
	wire _w7638_ ;
	wire _w7637_ ;
	wire _w7636_ ;
	wire _w7635_ ;
	wire _w7634_ ;
	wire _w7633_ ;
	wire _w7632_ ;
	wire _w7631_ ;
	wire _w7630_ ;
	wire _w7629_ ;
	wire _w7628_ ;
	wire _w7627_ ;
	wire _w7626_ ;
	wire _w7625_ ;
	wire _w7624_ ;
	wire _w7623_ ;
	wire _w7622_ ;
	wire _w7621_ ;
	wire _w7620_ ;
	wire _w7619_ ;
	wire _w7618_ ;
	wire _w7617_ ;
	wire _w7616_ ;
	wire _w7615_ ;
	wire _w7614_ ;
	wire _w7613_ ;
	wire _w7612_ ;
	wire _w7611_ ;
	wire _w7610_ ;
	wire _w7609_ ;
	wire _w7608_ ;
	wire _w7607_ ;
	wire _w7606_ ;
	wire _w7605_ ;
	wire _w7604_ ;
	wire _w7603_ ;
	wire _w7602_ ;
	wire _w7601_ ;
	wire _w7600_ ;
	wire _w7599_ ;
	wire _w7598_ ;
	wire _w7597_ ;
	wire _w7596_ ;
	wire _w7595_ ;
	wire _w7594_ ;
	wire _w7593_ ;
	wire _w7592_ ;
	wire _w7591_ ;
	wire _w7590_ ;
	wire _w7589_ ;
	wire _w7588_ ;
	wire _w7587_ ;
	wire _w7586_ ;
	wire _w7585_ ;
	wire _w7584_ ;
	wire _w7583_ ;
	wire _w7582_ ;
	wire _w7581_ ;
	wire _w7580_ ;
	wire _w7579_ ;
	wire _w7578_ ;
	wire _w7577_ ;
	wire _w7576_ ;
	wire _w7575_ ;
	wire _w7574_ ;
	wire _w7573_ ;
	wire _w7572_ ;
	wire _w7571_ ;
	wire _w7570_ ;
	wire _w7569_ ;
	wire _w7568_ ;
	wire _w7567_ ;
	wire _w7566_ ;
	wire _w7565_ ;
	wire _w7564_ ;
	wire _w7563_ ;
	wire _w7562_ ;
	wire _w7561_ ;
	wire _w7560_ ;
	wire _w7559_ ;
	wire _w7558_ ;
	wire _w7557_ ;
	wire _w7556_ ;
	wire _w7555_ ;
	wire _w7554_ ;
	wire _w7553_ ;
	wire _w7552_ ;
	wire _w7551_ ;
	wire _w7550_ ;
	wire _w7549_ ;
	wire _w7548_ ;
	wire _w7547_ ;
	wire _w7546_ ;
	wire _w7545_ ;
	wire _w7544_ ;
	wire _w7543_ ;
	wire _w7542_ ;
	wire _w7541_ ;
	wire _w7540_ ;
	wire _w7539_ ;
	wire _w7538_ ;
	wire _w7537_ ;
	wire _w7536_ ;
	wire _w7535_ ;
	wire _w7534_ ;
	wire _w7533_ ;
	wire _w7532_ ;
	wire _w7531_ ;
	wire _w7530_ ;
	wire _w7529_ ;
	wire _w7528_ ;
	wire _w7527_ ;
	wire _w7526_ ;
	wire _w7525_ ;
	wire _w7524_ ;
	wire _w7523_ ;
	wire _w7522_ ;
	wire _w7521_ ;
	wire _w7520_ ;
	wire _w7519_ ;
	wire _w7518_ ;
	wire _w7517_ ;
	wire _w7516_ ;
	wire _w7515_ ;
	wire _w7514_ ;
	wire _w7513_ ;
	wire _w7512_ ;
	wire _w7511_ ;
	wire _w7510_ ;
	wire _w7509_ ;
	wire _w7508_ ;
	wire _w7507_ ;
	wire _w7506_ ;
	wire _w7505_ ;
	wire _w7504_ ;
	wire _w7503_ ;
	wire _w7502_ ;
	wire _w7501_ ;
	wire _w7500_ ;
	wire _w7499_ ;
	wire _w7498_ ;
	wire _w7497_ ;
	wire _w7496_ ;
	wire _w7495_ ;
	wire _w7494_ ;
	wire _w7493_ ;
	wire _w7492_ ;
	wire _w7491_ ;
	wire _w7490_ ;
	wire _w7489_ ;
	wire _w7488_ ;
	wire _w7487_ ;
	wire _w7486_ ;
	wire _w7485_ ;
	wire _w7484_ ;
	wire _w7483_ ;
	wire _w7482_ ;
	wire _w7481_ ;
	wire _w7480_ ;
	wire _w7479_ ;
	wire _w7478_ ;
	wire _w7477_ ;
	wire _w7476_ ;
	wire _w7475_ ;
	wire _w7474_ ;
	wire _w7473_ ;
	wire _w7472_ ;
	wire _w7471_ ;
	wire _w7470_ ;
	wire _w7469_ ;
	wire _w7468_ ;
	wire _w7467_ ;
	wire _w7466_ ;
	wire _w7465_ ;
	wire _w7464_ ;
	wire _w7463_ ;
	wire _w7462_ ;
	wire _w7461_ ;
	wire _w7460_ ;
	wire _w7459_ ;
	wire _w7458_ ;
	wire _w7457_ ;
	wire _w7456_ ;
	wire _w7455_ ;
	wire _w7454_ ;
	wire _w7453_ ;
	wire _w7452_ ;
	wire _w7451_ ;
	wire _w7450_ ;
	wire _w7449_ ;
	wire _w7448_ ;
	wire _w7447_ ;
	wire _w7446_ ;
	wire _w7445_ ;
	wire _w7444_ ;
	wire _w7443_ ;
	wire _w7442_ ;
	wire _w7441_ ;
	wire _w7440_ ;
	wire _w7439_ ;
	wire _w7438_ ;
	wire _w7437_ ;
	wire _w7436_ ;
	wire _w7435_ ;
	wire _w7434_ ;
	wire _w7433_ ;
	wire _w7432_ ;
	wire _w7431_ ;
	wire _w7430_ ;
	wire _w7429_ ;
	wire _w7428_ ;
	wire _w7427_ ;
	wire _w7426_ ;
	wire _w7425_ ;
	wire _w7424_ ;
	wire _w7423_ ;
	wire _w7422_ ;
	wire _w7421_ ;
	wire _w7420_ ;
	wire _w7419_ ;
	wire _w7418_ ;
	wire _w7417_ ;
	wire _w7416_ ;
	wire _w7415_ ;
	wire _w7414_ ;
	wire _w7413_ ;
	wire _w7412_ ;
	wire _w7411_ ;
	wire _w7410_ ;
	wire _w7409_ ;
	wire _w7408_ ;
	wire _w7407_ ;
	wire _w7406_ ;
	wire _w7405_ ;
	wire _w7404_ ;
	wire _w7403_ ;
	wire _w7402_ ;
	wire _w7401_ ;
	wire _w7400_ ;
	wire _w7399_ ;
	wire _w7398_ ;
	wire _w7397_ ;
	wire _w7396_ ;
	wire _w7395_ ;
	wire _w7394_ ;
	wire _w7393_ ;
	wire _w7392_ ;
	wire _w7391_ ;
	wire _w7390_ ;
	wire _w7389_ ;
	wire _w7388_ ;
	wire _w7387_ ;
	wire _w7386_ ;
	wire _w7385_ ;
	wire _w7384_ ;
	wire _w7383_ ;
	wire _w7382_ ;
	wire _w7381_ ;
	wire _w7380_ ;
	wire _w7379_ ;
	wire _w7378_ ;
	wire _w7377_ ;
	wire _w7376_ ;
	wire _w7375_ ;
	wire _w7374_ ;
	wire _w7373_ ;
	wire _w7372_ ;
	wire _w7371_ ;
	wire _w7370_ ;
	wire _w7369_ ;
	wire _w7368_ ;
	wire _w7367_ ;
	wire _w7366_ ;
	wire _w7365_ ;
	wire _w7364_ ;
	wire _w7363_ ;
	wire _w7362_ ;
	wire _w7361_ ;
	wire _w7360_ ;
	wire _w7359_ ;
	wire _w7358_ ;
	wire _w7357_ ;
	wire _w7356_ ;
	wire _w7355_ ;
	wire _w7354_ ;
	wire _w7353_ ;
	wire _w7352_ ;
	wire _w7351_ ;
	wire _w7350_ ;
	wire _w7349_ ;
	wire _w7348_ ;
	wire _w7347_ ;
	wire _w7346_ ;
	wire _w7345_ ;
	wire _w7344_ ;
	wire _w7343_ ;
	wire _w7342_ ;
	wire _w7341_ ;
	wire _w7340_ ;
	wire _w7339_ ;
	wire _w7338_ ;
	wire _w7337_ ;
	wire _w7336_ ;
	wire _w7335_ ;
	wire _w7334_ ;
	wire _w7333_ ;
	wire _w7332_ ;
	wire _w7331_ ;
	wire _w7330_ ;
	wire _w7329_ ;
	wire _w7328_ ;
	wire _w7327_ ;
	wire _w7326_ ;
	wire _w7325_ ;
	wire _w7324_ ;
	wire _w7323_ ;
	wire _w7322_ ;
	wire _w7321_ ;
	wire _w7320_ ;
	wire _w7319_ ;
	wire _w7318_ ;
	wire _w7317_ ;
	wire _w7316_ ;
	wire _w7315_ ;
	wire _w7314_ ;
	wire _w7313_ ;
	wire _w7312_ ;
	wire _w7311_ ;
	wire _w7310_ ;
	wire _w7309_ ;
	wire _w7308_ ;
	wire _w7307_ ;
	wire _w7306_ ;
	wire _w7305_ ;
	wire _w7304_ ;
	wire _w7303_ ;
	wire _w7302_ ;
	wire _w7301_ ;
	wire _w7300_ ;
	wire _w7299_ ;
	wire _w7298_ ;
	wire _w7297_ ;
	wire _w7296_ ;
	wire _w7295_ ;
	wire _w7294_ ;
	wire _w7293_ ;
	wire _w7292_ ;
	wire _w7291_ ;
	wire _w7290_ ;
	wire _w7289_ ;
	wire _w7288_ ;
	wire _w7287_ ;
	wire _w7286_ ;
	wire _w7285_ ;
	wire _w7284_ ;
	wire _w7283_ ;
	wire _w7282_ ;
	wire _w7281_ ;
	wire _w7280_ ;
	wire _w7279_ ;
	wire _w7278_ ;
	wire _w7277_ ;
	wire _w7276_ ;
	wire _w7275_ ;
	wire _w7274_ ;
	wire _w7273_ ;
	wire _w7272_ ;
	wire _w7271_ ;
	wire _w7270_ ;
	wire _w7269_ ;
	wire _w7268_ ;
	wire _w7267_ ;
	wire _w7266_ ;
	wire _w7265_ ;
	wire _w7264_ ;
	wire _w7263_ ;
	wire _w7262_ ;
	wire _w7261_ ;
	wire _w7260_ ;
	wire _w7259_ ;
	wire _w7258_ ;
	wire _w7257_ ;
	wire _w7256_ ;
	wire _w7255_ ;
	wire _w7254_ ;
	wire _w7253_ ;
	wire _w7252_ ;
	wire _w7251_ ;
	wire _w7250_ ;
	wire _w7249_ ;
	wire _w7248_ ;
	wire _w7247_ ;
	wire _w7246_ ;
	wire _w7245_ ;
	wire _w7244_ ;
	wire _w7243_ ;
	wire _w7242_ ;
	wire _w7241_ ;
	wire _w7240_ ;
	wire _w7239_ ;
	wire _w7238_ ;
	wire _w7237_ ;
	wire _w7236_ ;
	wire _w7235_ ;
	wire _w7234_ ;
	wire _w7233_ ;
	wire _w7232_ ;
	wire _w7231_ ;
	wire _w7230_ ;
	wire _w7229_ ;
	wire _w7228_ ;
	wire _w7227_ ;
	wire _w7226_ ;
	wire _w7225_ ;
	wire _w7224_ ;
	wire _w7223_ ;
	wire _w7222_ ;
	wire _w7221_ ;
	wire _w7220_ ;
	wire _w7219_ ;
	wire _w7218_ ;
	wire _w7217_ ;
	wire _w7216_ ;
	wire _w7215_ ;
	wire _w7214_ ;
	wire _w7213_ ;
	wire _w7212_ ;
	wire _w7211_ ;
	wire _w7210_ ;
	wire _w7209_ ;
	wire _w7208_ ;
	wire _w7207_ ;
	wire _w7206_ ;
	wire _w7205_ ;
	wire _w7204_ ;
	wire _w7203_ ;
	wire _w7202_ ;
	wire _w7201_ ;
	wire _w7200_ ;
	wire _w7199_ ;
	wire _w7198_ ;
	wire _w7197_ ;
	wire _w7196_ ;
	wire _w7195_ ;
	wire _w7194_ ;
	wire _w7193_ ;
	wire _w7192_ ;
	wire _w7191_ ;
	wire _w7190_ ;
	wire _w7189_ ;
	wire _w7188_ ;
	wire _w7187_ ;
	wire _w7186_ ;
	wire _w7185_ ;
	wire _w7184_ ;
	wire _w7183_ ;
	wire _w7182_ ;
	wire _w7181_ ;
	wire _w7180_ ;
	wire _w7179_ ;
	wire _w7178_ ;
	wire _w7177_ ;
	wire _w7176_ ;
	wire _w7175_ ;
	wire _w7174_ ;
	wire _w7173_ ;
	wire _w7172_ ;
	wire _w7171_ ;
	wire _w7170_ ;
	wire _w7169_ ;
	wire _w7168_ ;
	wire _w7167_ ;
	wire _w7166_ ;
	wire _w7165_ ;
	wire _w7164_ ;
	wire _w7163_ ;
	wire _w7162_ ;
	wire _w7161_ ;
	wire _w7160_ ;
	wire _w7159_ ;
	wire _w7158_ ;
	wire _w7157_ ;
	wire _w7156_ ;
	wire _w7155_ ;
	wire _w7154_ ;
	wire _w7153_ ;
	wire _w7152_ ;
	wire _w7151_ ;
	wire _w7150_ ;
	wire _w7149_ ;
	wire _w7148_ ;
	wire _w7147_ ;
	wire _w7146_ ;
	wire _w7145_ ;
	wire _w7144_ ;
	wire _w7143_ ;
	wire _w7142_ ;
	wire _w7141_ ;
	wire _w7140_ ;
	wire _w7139_ ;
	wire _w7138_ ;
	wire _w7137_ ;
	wire _w7136_ ;
	wire _w7135_ ;
	wire _w7134_ ;
	wire _w7133_ ;
	wire _w7132_ ;
	wire _w7131_ ;
	wire _w7130_ ;
	wire _w7129_ ;
	wire _w7128_ ;
	wire _w7127_ ;
	wire _w7126_ ;
	wire _w7125_ ;
	wire _w7124_ ;
	wire _w7123_ ;
	wire _w7122_ ;
	wire _w7121_ ;
	wire _w7120_ ;
	wire _w7119_ ;
	wire _w7118_ ;
	wire _w7117_ ;
	wire _w7116_ ;
	wire _w7115_ ;
	wire _w7114_ ;
	wire _w7113_ ;
	wire _w7112_ ;
	wire _w7111_ ;
	wire _w7110_ ;
	wire _w7109_ ;
	wire _w7108_ ;
	wire _w7107_ ;
	wire _w7106_ ;
	wire _w7105_ ;
	wire _w7104_ ;
	wire _w7103_ ;
	wire _w7102_ ;
	wire _w7101_ ;
	wire _w7100_ ;
	wire _w7099_ ;
	wire _w7098_ ;
	wire _w7097_ ;
	wire _w7096_ ;
	wire _w7095_ ;
	wire _w7094_ ;
	wire _w7093_ ;
	wire _w7092_ ;
	wire _w7091_ ;
	wire _w7090_ ;
	wire _w7089_ ;
	wire _w7088_ ;
	wire _w7087_ ;
	wire _w7086_ ;
	wire _w7085_ ;
	wire _w7084_ ;
	wire _w7083_ ;
	wire _w7082_ ;
	wire _w7081_ ;
	wire _w7080_ ;
	wire _w7079_ ;
	wire _w7078_ ;
	wire _w7077_ ;
	wire _w7076_ ;
	wire _w7075_ ;
	wire _w7074_ ;
	wire _w7073_ ;
	wire _w7072_ ;
	wire _w7071_ ;
	wire _w7070_ ;
	wire _w7069_ ;
	wire _w7068_ ;
	wire _w7067_ ;
	wire _w7066_ ;
	wire _w7065_ ;
	wire _w7064_ ;
	wire _w7063_ ;
	wire _w7062_ ;
	wire _w7061_ ;
	wire _w7060_ ;
	wire _w7059_ ;
	wire _w7058_ ;
	wire _w7057_ ;
	wire _w7056_ ;
	wire _w7055_ ;
	wire _w7054_ ;
	wire _w7053_ ;
	wire _w7052_ ;
	wire _w7051_ ;
	wire _w7050_ ;
	wire _w7049_ ;
	wire _w7048_ ;
	wire _w7047_ ;
	wire _w7046_ ;
	wire _w7045_ ;
	wire _w7044_ ;
	wire _w7043_ ;
	wire _w7042_ ;
	wire _w7041_ ;
	wire _w7040_ ;
	wire _w7039_ ;
	wire _w7038_ ;
	wire _w7037_ ;
	wire _w7036_ ;
	wire _w7035_ ;
	wire _w7034_ ;
	wire _w7033_ ;
	wire _w7032_ ;
	wire _w7031_ ;
	wire _w7030_ ;
	wire _w7029_ ;
	wire _w7028_ ;
	wire _w7027_ ;
	wire _w7026_ ;
	wire _w7025_ ;
	wire _w7024_ ;
	wire _w7023_ ;
	wire _w7022_ ;
	wire _w7021_ ;
	wire _w7020_ ;
	wire _w7019_ ;
	wire _w7018_ ;
	wire _w7017_ ;
	wire _w7016_ ;
	wire _w7015_ ;
	wire _w7014_ ;
	wire _w7013_ ;
	wire _w7012_ ;
	wire _w7011_ ;
	wire _w7010_ ;
	wire _w7009_ ;
	wire _w7008_ ;
	wire _w7007_ ;
	wire _w7006_ ;
	wire _w7005_ ;
	wire _w7004_ ;
	wire _w7003_ ;
	wire _w7002_ ;
	wire _w7001_ ;
	wire _w7000_ ;
	wire _w6999_ ;
	wire _w6998_ ;
	wire _w6997_ ;
	wire _w6996_ ;
	wire _w6995_ ;
	wire _w6994_ ;
	wire _w6993_ ;
	wire _w6992_ ;
	wire _w6991_ ;
	wire _w6990_ ;
	wire _w6989_ ;
	wire _w6988_ ;
	wire _w6987_ ;
	wire _w6986_ ;
	wire _w6985_ ;
	wire _w6984_ ;
	wire _w6983_ ;
	wire _w6982_ ;
	wire _w6981_ ;
	wire _w6980_ ;
	wire _w6979_ ;
	wire _w6978_ ;
	wire _w6977_ ;
	wire _w6976_ ;
	wire _w6975_ ;
	wire _w6974_ ;
	wire _w6973_ ;
	wire _w6972_ ;
	wire _w6971_ ;
	wire _w6970_ ;
	wire _w6969_ ;
	wire _w6968_ ;
	wire _w6967_ ;
	wire _w6966_ ;
	wire _w6965_ ;
	wire _w6964_ ;
	wire _w6963_ ;
	wire _w6962_ ;
	wire _w6961_ ;
	wire _w6960_ ;
	wire _w6959_ ;
	wire _w6958_ ;
	wire _w6957_ ;
	wire _w6956_ ;
	wire _w6955_ ;
	wire _w6954_ ;
	wire _w6953_ ;
	wire _w6952_ ;
	wire _w6951_ ;
	wire _w6950_ ;
	wire _w6949_ ;
	wire _w6948_ ;
	wire _w6947_ ;
	wire _w6946_ ;
	wire _w6945_ ;
	wire _w6944_ ;
	wire _w6943_ ;
	wire _w6942_ ;
	wire _w6941_ ;
	wire _w6940_ ;
	wire _w6939_ ;
	wire _w6938_ ;
	wire _w6937_ ;
	wire _w6936_ ;
	wire _w6935_ ;
	wire _w6934_ ;
	wire _w6933_ ;
	wire _w6932_ ;
	wire _w6931_ ;
	wire _w6930_ ;
	wire _w6929_ ;
	wire _w6928_ ;
	wire _w6927_ ;
	wire _w6926_ ;
	wire _w6925_ ;
	wire _w6924_ ;
	wire _w6923_ ;
	wire _w6922_ ;
	wire _w6921_ ;
	wire _w6920_ ;
	wire _w6919_ ;
	wire _w6918_ ;
	wire _w6917_ ;
	wire _w6916_ ;
	wire _w6915_ ;
	wire _w6914_ ;
	wire _w6913_ ;
	wire _w6912_ ;
	wire _w6911_ ;
	wire _w6910_ ;
	wire _w6909_ ;
	wire _w6908_ ;
	wire _w6907_ ;
	wire _w6906_ ;
	wire _w6905_ ;
	wire _w6904_ ;
	wire _w6903_ ;
	wire _w6902_ ;
	wire _w6901_ ;
	wire _w6900_ ;
	wire _w6899_ ;
	wire _w6898_ ;
	wire _w6897_ ;
	wire _w6896_ ;
	wire _w6895_ ;
	wire _w6894_ ;
	wire _w6893_ ;
	wire _w6892_ ;
	wire _w6891_ ;
	wire _w6890_ ;
	wire _w6889_ ;
	wire _w6888_ ;
	wire _w6887_ ;
	wire _w6886_ ;
	wire _w6885_ ;
	wire _w6884_ ;
	wire _w6883_ ;
	wire _w6882_ ;
	wire _w6881_ ;
	wire _w6880_ ;
	wire _w6879_ ;
	wire _w6878_ ;
	wire _w6877_ ;
	wire _w6876_ ;
	wire _w6875_ ;
	wire _w6874_ ;
	wire _w6873_ ;
	wire _w6872_ ;
	wire _w6871_ ;
	wire _w6870_ ;
	wire _w6869_ ;
	wire _w6868_ ;
	wire _w6867_ ;
	wire _w6866_ ;
	wire _w6865_ ;
	wire _w6864_ ;
	wire _w6863_ ;
	wire _w6862_ ;
	wire _w6861_ ;
	wire _w6860_ ;
	wire _w6859_ ;
	wire _w6858_ ;
	wire _w6857_ ;
	wire _w6856_ ;
	wire _w6855_ ;
	wire _w6854_ ;
	wire _w6853_ ;
	wire _w6852_ ;
	wire _w6851_ ;
	wire _w6850_ ;
	wire _w6849_ ;
	wire _w6848_ ;
	wire _w6847_ ;
	wire _w6846_ ;
	wire _w6845_ ;
	wire _w6844_ ;
	wire _w6843_ ;
	wire _w6842_ ;
	wire _w6841_ ;
	wire _w6840_ ;
	wire _w6839_ ;
	wire _w6838_ ;
	wire _w6837_ ;
	wire _w6836_ ;
	wire _w6835_ ;
	wire _w6834_ ;
	wire _w6833_ ;
	wire _w6832_ ;
	wire _w6831_ ;
	wire _w6830_ ;
	wire _w6829_ ;
	wire _w6828_ ;
	wire _w6827_ ;
	wire _w6826_ ;
	wire _w6825_ ;
	wire _w6824_ ;
	wire _w6823_ ;
	wire _w6822_ ;
	wire _w6821_ ;
	wire _w6820_ ;
	wire _w6819_ ;
	wire _w6818_ ;
	wire _w6817_ ;
	wire _w6816_ ;
	wire _w6815_ ;
	wire _w6814_ ;
	wire _w6813_ ;
	wire _w6812_ ;
	wire _w6811_ ;
	wire _w6810_ ;
	wire _w6809_ ;
	wire _w6808_ ;
	wire _w6807_ ;
	wire _w6806_ ;
	wire _w6805_ ;
	wire _w6804_ ;
	wire _w6803_ ;
	wire _w6802_ ;
	wire _w6801_ ;
	wire _w6800_ ;
	wire _w6799_ ;
	wire _w6798_ ;
	wire _w6797_ ;
	wire _w6796_ ;
	wire _w6795_ ;
	wire _w6794_ ;
	wire _w6793_ ;
	wire _w6792_ ;
	wire _w6791_ ;
	wire _w6790_ ;
	wire _w6789_ ;
	wire _w6788_ ;
	wire _w6787_ ;
	wire _w6786_ ;
	wire _w6785_ ;
	wire _w6784_ ;
	wire _w6783_ ;
	wire _w6782_ ;
	wire _w6781_ ;
	wire _w6780_ ;
	wire _w6779_ ;
	wire _w6778_ ;
	wire _w6777_ ;
	wire _w6776_ ;
	wire _w6775_ ;
	wire _w6774_ ;
	wire _w6773_ ;
	wire _w6772_ ;
	wire _w6771_ ;
	wire _w6770_ ;
	wire _w6769_ ;
	wire _w6768_ ;
	wire _w6767_ ;
	wire _w6766_ ;
	wire _w6765_ ;
	wire _w6764_ ;
	wire _w6763_ ;
	wire _w6762_ ;
	wire _w6761_ ;
	wire _w6760_ ;
	wire _w6759_ ;
	wire _w6758_ ;
	wire _w6757_ ;
	wire _w6756_ ;
	wire _w6755_ ;
	wire _w6754_ ;
	wire _w6753_ ;
	wire _w6752_ ;
	wire _w6751_ ;
	wire _w6750_ ;
	wire _w6749_ ;
	wire _w6748_ ;
	wire _w6747_ ;
	wire _w6746_ ;
	wire _w6745_ ;
	wire _w6744_ ;
	wire _w6743_ ;
	wire _w6742_ ;
	wire _w6741_ ;
	wire _w6740_ ;
	wire _w6739_ ;
	wire _w6738_ ;
	wire _w6737_ ;
	wire _w6736_ ;
	wire _w6735_ ;
	wire _w6734_ ;
	wire _w6733_ ;
	wire _w6732_ ;
	wire _w6731_ ;
	wire _w6730_ ;
	wire _w6729_ ;
	wire _w6728_ ;
	wire _w6727_ ;
	wire _w6726_ ;
	wire _w6725_ ;
	wire _w6724_ ;
	wire _w6723_ ;
	wire _w6722_ ;
	wire _w6721_ ;
	wire _w6720_ ;
	wire _w6719_ ;
	wire _w6718_ ;
	wire _w6717_ ;
	wire _w6716_ ;
	wire _w6715_ ;
	wire _w6714_ ;
	wire _w6713_ ;
	wire _w6712_ ;
	wire _w6711_ ;
	wire _w6710_ ;
	wire _w6709_ ;
	wire _w6708_ ;
	wire _w6707_ ;
	wire _w6706_ ;
	wire _w6705_ ;
	wire _w6704_ ;
	wire _w6703_ ;
	wire _w6702_ ;
	wire _w6701_ ;
	wire _w6700_ ;
	wire _w6699_ ;
	wire _w6698_ ;
	wire _w6697_ ;
	wire _w6696_ ;
	wire _w6695_ ;
	wire _w6694_ ;
	wire _w6693_ ;
	wire _w6692_ ;
	wire _w6691_ ;
	wire _w6690_ ;
	wire _w6689_ ;
	wire _w6688_ ;
	wire _w6687_ ;
	wire _w6686_ ;
	wire _w6685_ ;
	wire _w6684_ ;
	wire _w6683_ ;
	wire _w6682_ ;
	wire _w6681_ ;
	wire _w6680_ ;
	wire _w6679_ ;
	wire _w6678_ ;
	wire _w6677_ ;
	wire _w6676_ ;
	wire _w6675_ ;
	wire _w6674_ ;
	wire _w6673_ ;
	wire _w6672_ ;
	wire _w6671_ ;
	wire _w6670_ ;
	wire _w6669_ ;
	wire _w6668_ ;
	wire _w6667_ ;
	wire _w6666_ ;
	wire _w6665_ ;
	wire _w6664_ ;
	wire _w6663_ ;
	wire _w6662_ ;
	wire _w6661_ ;
	wire _w6660_ ;
	wire _w6659_ ;
	wire _w6658_ ;
	wire _w6657_ ;
	wire _w6656_ ;
	wire _w6655_ ;
	wire _w6654_ ;
	wire _w6653_ ;
	wire _w6652_ ;
	wire _w6651_ ;
	wire _w6650_ ;
	wire _w6649_ ;
	wire _w6648_ ;
	wire _w6647_ ;
	wire _w6646_ ;
	wire _w6645_ ;
	wire _w6644_ ;
	wire _w6643_ ;
	wire _w6642_ ;
	wire _w6641_ ;
	wire _w6640_ ;
	wire _w6639_ ;
	wire _w6638_ ;
	wire _w6637_ ;
	wire _w6636_ ;
	wire _w6635_ ;
	wire _w6634_ ;
	wire _w6633_ ;
	wire _w6632_ ;
	wire _w6631_ ;
	wire _w6630_ ;
	wire _w6629_ ;
	wire _w6628_ ;
	wire _w6627_ ;
	wire _w6626_ ;
	wire _w6625_ ;
	wire _w6624_ ;
	wire _w6623_ ;
	wire _w6622_ ;
	wire _w6621_ ;
	wire _w6620_ ;
	wire _w6619_ ;
	wire _w6618_ ;
	wire _w6617_ ;
	wire _w6616_ ;
	wire _w6615_ ;
	wire _w6614_ ;
	wire _w6613_ ;
	wire _w6612_ ;
	wire _w6611_ ;
	wire _w6610_ ;
	wire _w6609_ ;
	wire _w6608_ ;
	wire _w6607_ ;
	wire _w6606_ ;
	wire _w6605_ ;
	wire _w6604_ ;
	wire _w6603_ ;
	wire _w6602_ ;
	wire _w6601_ ;
	wire _w6600_ ;
	wire _w6599_ ;
	wire _w6598_ ;
	wire _w6597_ ;
	wire _w6596_ ;
	wire _w6595_ ;
	wire _w3864_ ;
	wire _w3863_ ;
	wire _w3862_ ;
	wire _w3861_ ;
	wire _w3860_ ;
	wire _w3859_ ;
	wire _w3858_ ;
	wire _w3857_ ;
	wire _w3856_ ;
	wire _w3855_ ;
	wire _w3854_ ;
	wire _w3853_ ;
	wire _w3852_ ;
	wire _w3851_ ;
	wire _w3850_ ;
	wire _w3849_ ;
	wire _w3848_ ;
	wire _w3847_ ;
	wire _w3846_ ;
	wire _w3845_ ;
	wire _w3844_ ;
	wire _w3843_ ;
	wire _w3842_ ;
	wire _w3841_ ;
	wire _w3840_ ;
	wire _w3839_ ;
	wire _w3838_ ;
	wire _w3837_ ;
	wire _w3836_ ;
	wire _w3835_ ;
	wire _w3834_ ;
	wire _w3833_ ;
	wire _w3832_ ;
	wire _w3831_ ;
	wire _w3830_ ;
	wire _w3829_ ;
	wire _w3828_ ;
	wire _w3827_ ;
	wire _w3826_ ;
	wire _w3825_ ;
	wire _w3824_ ;
	wire _w3823_ ;
	wire _w3822_ ;
	wire _w3821_ ;
	wire _w3820_ ;
	wire _w3819_ ;
	wire _w3818_ ;
	wire _w3817_ ;
	wire _w3816_ ;
	wire _w3815_ ;
	wire _w3814_ ;
	wire _w3813_ ;
	wire _w3812_ ;
	wire _w3811_ ;
	wire _w3810_ ;
	wire _w3809_ ;
	wire _w3808_ ;
	wire _w3807_ ;
	wire _w3806_ ;
	wire _w3805_ ;
	wire _w3804_ ;
	wire _w3803_ ;
	wire _w3802_ ;
	wire _w3801_ ;
	wire _w3800_ ;
	wire _w3799_ ;
	wire _w3798_ ;
	wire _w3797_ ;
	wire _w3796_ ;
	wire _w3795_ ;
	wire _w3794_ ;
	wire _w3793_ ;
	wire _w3792_ ;
	wire _w3791_ ;
	wire _w3790_ ;
	wire _w3789_ ;
	wire _w3788_ ;
	wire _w3787_ ;
	wire _w3786_ ;
	wire _w3785_ ;
	wire _w3784_ ;
	wire _w3783_ ;
	wire _w3782_ ;
	wire _w3781_ ;
	wire _w3780_ ;
	wire _w3779_ ;
	wire _w3778_ ;
	wire _w3777_ ;
	wire _w3776_ ;
	wire _w3775_ ;
	wire _w3774_ ;
	wire _w3773_ ;
	wire _w3772_ ;
	wire _w3771_ ;
	wire _w3770_ ;
	wire _w3769_ ;
	wire _w3768_ ;
	wire _w3767_ ;
	wire _w3766_ ;
	wire _w3765_ ;
	wire _w3764_ ;
	wire _w3763_ ;
	wire _w3762_ ;
	wire _w3761_ ;
	wire _w3760_ ;
	wire _w3759_ ;
	wire _w3758_ ;
	wire _w3757_ ;
	wire _w3756_ ;
	wire _w3755_ ;
	wire _w3754_ ;
	wire _w3753_ ;
	wire _w3752_ ;
	wire _w3751_ ;
	wire _w3750_ ;
	wire _w3749_ ;
	wire _w3748_ ;
	wire _w3747_ ;
	wire _w3746_ ;
	wire _w3745_ ;
	wire _w3744_ ;
	wire _w3743_ ;
	wire _w3742_ ;
	wire _w3741_ ;
	wire _w3740_ ;
	wire _w3739_ ;
	wire _w3738_ ;
	wire _w3737_ ;
	wire _w3736_ ;
	wire _w3735_ ;
	wire _w3734_ ;
	wire _w3733_ ;
	wire _w3732_ ;
	wire _w3731_ ;
	wire _w3730_ ;
	wire _w3729_ ;
	wire _w3728_ ;
	wire _w3727_ ;
	wire _w3726_ ;
	wire _w3725_ ;
	wire _w3724_ ;
	wire _w3723_ ;
	wire _w3722_ ;
	wire _w3721_ ;
	wire _w3720_ ;
	wire _w3719_ ;
	wire _w3718_ ;
	wire _w3717_ ;
	wire _w3716_ ;
	wire _w3715_ ;
	wire _w3714_ ;
	wire _w3713_ ;
	wire _w3712_ ;
	wire _w3711_ ;
	wire _w3710_ ;
	wire _w3709_ ;
	wire _w3708_ ;
	wire _w3707_ ;
	wire _w3706_ ;
	wire _w3705_ ;
	wire _w3704_ ;
	wire _w3703_ ;
	wire _w3702_ ;
	wire _w3701_ ;
	wire _w3700_ ;
	wire _w3699_ ;
	wire _w3698_ ;
	wire _w3697_ ;
	wire _w3696_ ;
	wire _w3695_ ;
	wire _w3694_ ;
	wire _w3693_ ;
	wire _w3692_ ;
	wire _w3691_ ;
	wire _w3690_ ;
	wire _w3689_ ;
	wire _w3688_ ;
	wire _w3687_ ;
	wire _w3686_ ;
	wire _w3685_ ;
	wire _w3684_ ;
	wire _w3683_ ;
	wire _w3682_ ;
	wire _w3681_ ;
	wire _w3680_ ;
	wire _w3679_ ;
	wire _w3678_ ;
	wire _w3677_ ;
	wire _w3676_ ;
	wire _w3675_ ;
	wire _w3674_ ;
	wire _w3673_ ;
	wire _w3672_ ;
	wire _w3671_ ;
	wire _w3670_ ;
	wire _w3669_ ;
	wire _w3668_ ;
	wire _w3667_ ;
	wire _w3666_ ;
	wire _w3665_ ;
	wire _w3664_ ;
	wire _w3663_ ;
	wire _w3662_ ;
	wire _w3661_ ;
	wire _w3660_ ;
	wire _w3659_ ;
	wire _w3658_ ;
	wire _w3657_ ;
	wire _w3656_ ;
	wire _w3655_ ;
	wire _w3654_ ;
	wire _w3653_ ;
	wire _w3652_ ;
	wire _w3651_ ;
	wire _w3650_ ;
	wire _w3649_ ;
	wire _w3648_ ;
	wire _w3647_ ;
	wire _w3646_ ;
	wire _w3645_ ;
	wire _w3644_ ;
	wire _w3643_ ;
	wire _w3642_ ;
	wire _w3641_ ;
	wire _w3640_ ;
	wire _w3639_ ;
	wire _w3638_ ;
	wire _w3637_ ;
	wire _w3636_ ;
	wire _w3635_ ;
	wire _w3634_ ;
	wire _w3633_ ;
	wire _w3632_ ;
	wire _w3631_ ;
	wire _w3630_ ;
	wire _w3629_ ;
	wire _w3628_ ;
	wire _w3627_ ;
	wire _w3626_ ;
	wire _w3625_ ;
	wire _w3624_ ;
	wire _w3623_ ;
	wire _w3622_ ;
	wire _w3621_ ;
	wire _w3620_ ;
	wire _w3619_ ;
	wire _w3618_ ;
	wire _w3617_ ;
	wire _w3616_ ;
	wire _w3615_ ;
	wire _w3614_ ;
	wire _w3613_ ;
	wire _w3612_ ;
	wire _w3611_ ;
	wire _w3610_ ;
	wire _w3609_ ;
	wire _w3608_ ;
	wire _w3607_ ;
	wire _w3606_ ;
	wire _w3605_ ;
	wire _w3604_ ;
	wire _w3603_ ;
	wire _w3602_ ;
	wire _w3601_ ;
	wire _w3600_ ;
	wire _w3599_ ;
	wire _w3598_ ;
	wire _w3597_ ;
	wire _w3596_ ;
	wire _w3595_ ;
	wire _w3594_ ;
	wire _w3593_ ;
	wire _w3592_ ;
	wire _w3591_ ;
	wire _w3590_ ;
	wire _w3589_ ;
	wire _w3588_ ;
	wire _w3587_ ;
	wire _w3586_ ;
	wire _w3585_ ;
	wire _w3584_ ;
	wire _w3583_ ;
	wire _w3582_ ;
	wire _w3581_ ;
	wire _w3580_ ;
	wire _w3579_ ;
	wire _w3578_ ;
	wire _w3577_ ;
	wire _w3576_ ;
	wire _w3575_ ;
	wire _w3574_ ;
	wire _w3573_ ;
	wire _w3572_ ;
	wire _w3571_ ;
	wire _w3570_ ;
	wire _w3569_ ;
	wire _w3568_ ;
	wire _w3567_ ;
	wire _w3566_ ;
	wire _w3565_ ;
	wire _w3564_ ;
	wire _w3563_ ;
	wire _w3562_ ;
	wire _w3561_ ;
	wire _w3560_ ;
	wire _w3559_ ;
	wire _w3558_ ;
	wire _w3557_ ;
	wire _w3556_ ;
	wire _w3555_ ;
	wire _w3554_ ;
	wire _w3553_ ;
	wire _w3552_ ;
	wire _w3551_ ;
	wire _w3550_ ;
	wire _w3549_ ;
	wire _w3548_ ;
	wire _w3547_ ;
	wire _w3546_ ;
	wire _w3545_ ;
	wire _w3544_ ;
	wire _w3543_ ;
	wire _w3542_ ;
	wire _w3541_ ;
	wire _w3540_ ;
	wire _w3539_ ;
	wire _w3538_ ;
	wire _w3537_ ;
	wire _w3536_ ;
	wire _w3535_ ;
	wire _w3534_ ;
	wire _w3533_ ;
	wire _w3532_ ;
	wire _w3531_ ;
	wire _w3530_ ;
	wire _w3529_ ;
	wire _w3528_ ;
	wire _w3527_ ;
	wire _w3526_ ;
	wire _w3525_ ;
	wire _w3524_ ;
	wire _w3523_ ;
	wire _w3522_ ;
	wire _w3521_ ;
	wire _w3520_ ;
	wire _w3519_ ;
	wire _w3518_ ;
	wire _w3517_ ;
	wire _w3516_ ;
	wire _w3515_ ;
	wire _w3514_ ;
	wire _w3513_ ;
	wire _w3512_ ;
	wire _w3511_ ;
	wire _w3510_ ;
	wire _w3509_ ;
	wire _w3508_ ;
	wire _w3507_ ;
	wire _w3506_ ;
	wire _w3505_ ;
	wire _w3504_ ;
	wire _w3503_ ;
	wire _w3502_ ;
	wire _w3501_ ;
	wire _w3500_ ;
	wire _w3499_ ;
	wire _w3498_ ;
	wire _w3497_ ;
	wire _w3496_ ;
	wire _w3495_ ;
	wire _w3494_ ;
	wire _w3493_ ;
	wire _w3492_ ;
	wire _w3491_ ;
	wire _w3490_ ;
	wire _w3489_ ;
	wire _w3488_ ;
	wire _w3487_ ;
	wire _w3486_ ;
	wire _w3485_ ;
	wire _w3484_ ;
	wire _w3483_ ;
	wire _w3482_ ;
	wire _w3481_ ;
	wire _w3480_ ;
	wire _w3479_ ;
	wire _w3478_ ;
	wire _w3477_ ;
	wire _w3476_ ;
	wire _w3475_ ;
	wire _w3474_ ;
	wire _w3473_ ;
	wire _w3472_ ;
	wire _w3471_ ;
	wire _w3470_ ;
	wire _w3469_ ;
	wire _w3468_ ;
	wire _w3467_ ;
	wire _w3466_ ;
	wire _w3465_ ;
	wire _w3464_ ;
	wire _w3463_ ;
	wire _w3462_ ;
	wire _w3461_ ;
	wire _w3460_ ;
	wire _w3459_ ;
	wire _w3458_ ;
	wire _w3457_ ;
	wire _w3456_ ;
	wire _w3455_ ;
	wire _w3454_ ;
	wire _w3453_ ;
	wire _w3452_ ;
	wire _w3451_ ;
	wire _w3450_ ;
	wire _w3449_ ;
	wire _w3448_ ;
	wire _w3447_ ;
	wire _w3446_ ;
	wire _w3445_ ;
	wire _w3444_ ;
	wire _w3443_ ;
	wire _w3442_ ;
	wire _w3441_ ;
	wire _w3440_ ;
	wire _w3439_ ;
	wire _w3438_ ;
	wire _w3437_ ;
	wire _w3436_ ;
	wire _w3435_ ;
	wire _w3434_ ;
	wire _w3433_ ;
	wire _w3432_ ;
	wire _w3431_ ;
	wire _w3430_ ;
	wire _w3429_ ;
	wire _w3428_ ;
	wire _w3427_ ;
	wire _w3426_ ;
	wire _w3425_ ;
	wire _w3424_ ;
	wire _w3423_ ;
	wire _w3422_ ;
	wire _w3421_ ;
	wire _w3420_ ;
	wire _w3419_ ;
	wire _w3418_ ;
	wire _w3417_ ;
	wire _w3416_ ;
	wire _w3415_ ;
	wire _w3414_ ;
	wire _w3413_ ;
	wire _w3412_ ;
	wire _w3411_ ;
	wire _w3410_ ;
	wire _w3409_ ;
	wire _w3408_ ;
	wire _w3407_ ;
	wire _w3406_ ;
	wire _w3405_ ;
	wire _w3404_ ;
	wire _w3403_ ;
	wire _w3402_ ;
	wire _w3401_ ;
	wire _w3400_ ;
	wire _w3399_ ;
	wire _w3398_ ;
	wire _w3397_ ;
	wire _w3396_ ;
	wire _w3395_ ;
	wire _w3394_ ;
	wire _w3393_ ;
	wire _w3392_ ;
	wire _w3391_ ;
	wire _w3390_ ;
	wire _w3389_ ;
	wire _w3388_ ;
	wire _w3387_ ;
	wire _w3386_ ;
	wire _w3385_ ;
	wire _w3384_ ;
	wire _w3383_ ;
	wire _w3382_ ;
	wire _w3381_ ;
	wire _w3380_ ;
	wire _w3379_ ;
	wire _w3378_ ;
	wire _w3377_ ;
	wire _w3376_ ;
	wire _w3375_ ;
	wire _w3374_ ;
	wire _w3373_ ;
	wire _w3372_ ;
	wire _w3371_ ;
	wire _w3370_ ;
	wire _w3369_ ;
	wire _w3368_ ;
	wire _w3367_ ;
	wire _w3366_ ;
	wire _w3365_ ;
	wire _w3364_ ;
	wire _w3363_ ;
	wire _w3362_ ;
	wire _w3361_ ;
	wire _w3360_ ;
	wire _w3359_ ;
	wire _w3358_ ;
	wire _w3357_ ;
	wire _w3356_ ;
	wire _w3355_ ;
	wire _w3354_ ;
	wire _w3353_ ;
	wire _w3352_ ;
	wire _w3351_ ;
	wire _w3350_ ;
	wire _w3349_ ;
	wire _w3348_ ;
	wire _w3347_ ;
	wire _w3346_ ;
	wire _w3345_ ;
	wire _w3344_ ;
	wire _w3343_ ;
	wire _w3342_ ;
	wire _w3341_ ;
	wire _w3340_ ;
	wire _w3339_ ;
	wire _w3338_ ;
	wire _w3337_ ;
	wire _w3336_ ;
	wire _w3335_ ;
	wire _w3334_ ;
	wire _w3333_ ;
	wire _w3332_ ;
	wire _w3331_ ;
	wire _w3330_ ;
	wire _w3329_ ;
	wire _w3328_ ;
	wire _w3327_ ;
	wire _w3326_ ;
	wire _w3325_ ;
	wire _w3324_ ;
	wire _w3323_ ;
	wire _w3322_ ;
	wire _w3321_ ;
	wire _w3320_ ;
	wire _w3319_ ;
	wire _w3318_ ;
	wire _w3317_ ;
	wire _w3316_ ;
	wire _w3315_ ;
	wire _w3314_ ;
	wire _w3313_ ;
	wire _w3312_ ;
	wire _w3311_ ;
	wire _w3310_ ;
	wire _w3309_ ;
	wire _w3308_ ;
	wire _w3307_ ;
	wire _w3306_ ;
	wire _w3305_ ;
	wire _w3304_ ;
	wire _w3303_ ;
	wire _w3302_ ;
	wire _w3301_ ;
	wire _w3300_ ;
	wire _w3299_ ;
	wire _w3298_ ;
	wire _w3297_ ;
	wire _w3296_ ;
	wire _w3295_ ;
	wire _w3294_ ;
	wire _w3293_ ;
	wire _w3292_ ;
	wire _w3291_ ;
	wire _w3290_ ;
	wire _w3289_ ;
	wire _w3288_ ;
	wire _w3287_ ;
	wire _w3286_ ;
	wire _w3285_ ;
	wire _w3284_ ;
	wire _w3283_ ;
	wire _w3282_ ;
	wire _w3281_ ;
	wire _w3280_ ;
	wire _w3279_ ;
	wire _w3278_ ;
	wire _w3277_ ;
	wire _w3276_ ;
	wire _w3275_ ;
	wire _w3274_ ;
	wire _w3273_ ;
	wire _w3272_ ;
	wire _w3271_ ;
	wire _w3270_ ;
	wire _w3269_ ;
	wire _w3268_ ;
	wire _w3267_ ;
	wire _w3266_ ;
	wire _w3265_ ;
	wire _w3264_ ;
	wire _w3263_ ;
	wire _w3262_ ;
	wire _w3261_ ;
	wire _w3260_ ;
	wire _w3259_ ;
	wire _w3258_ ;
	wire _w3257_ ;
	wire _w3256_ ;
	wire _w3255_ ;
	wire _w3254_ ;
	wire _w3253_ ;
	wire _w3252_ ;
	wire _w3251_ ;
	wire _w3250_ ;
	wire _w3249_ ;
	wire _w3248_ ;
	wire _w3247_ ;
	wire _w3246_ ;
	wire _w3245_ ;
	wire _w3244_ ;
	wire _w3243_ ;
	wire _w3242_ ;
	wire _w3241_ ;
	wire _w3240_ ;
	wire _w3239_ ;
	wire _w3238_ ;
	wire _w3237_ ;
	wire _w3236_ ;
	wire _w3235_ ;
	wire _w3234_ ;
	wire _w3233_ ;
	wire _w3232_ ;
	wire _w3231_ ;
	wire _w3230_ ;
	wire _w3229_ ;
	wire _w3228_ ;
	wire _w3227_ ;
	wire _w3226_ ;
	wire _w3225_ ;
	wire _w3224_ ;
	wire _w3223_ ;
	wire _w3222_ ;
	wire _w3221_ ;
	wire _w3220_ ;
	wire _w3219_ ;
	wire _w3218_ ;
	wire _w3217_ ;
	wire _w3216_ ;
	wire _w3215_ ;
	wire _w3214_ ;
	wire _w3213_ ;
	wire _w3212_ ;
	wire _w3211_ ;
	wire _w3210_ ;
	wire _w3209_ ;
	wire _w3208_ ;
	wire _w3207_ ;
	wire _w3206_ ;
	wire _w3205_ ;
	wire _w3204_ ;
	wire _w3203_ ;
	wire _w3202_ ;
	wire _w3201_ ;
	wire _w3200_ ;
	wire _w3199_ ;
	wire _w3198_ ;
	wire _w3197_ ;
	wire _w3196_ ;
	wire _w3195_ ;
	wire _w3194_ ;
	wire _w3193_ ;
	wire _w3192_ ;
	wire _w3191_ ;
	wire _w3190_ ;
	wire _w3189_ ;
	wire _w3188_ ;
	wire _w3187_ ;
	wire _w3186_ ;
	wire _w3185_ ;
	wire _w3184_ ;
	wire _w3183_ ;
	wire _w3182_ ;
	wire _w3181_ ;
	wire _w3180_ ;
	wire _w3179_ ;
	wire _w3178_ ;
	wire _w3177_ ;
	wire _w3176_ ;
	wire _w3175_ ;
	wire _w3174_ ;
	wire _w3173_ ;
	wire _w3172_ ;
	wire _w3171_ ;
	wire _w3170_ ;
	wire _w3169_ ;
	wire _w3168_ ;
	wire _w3167_ ;
	wire _w3166_ ;
	wire _w3165_ ;
	wire _w3164_ ;
	wire _w3163_ ;
	wire _w3162_ ;
	wire _w3161_ ;
	wire _w3160_ ;
	wire _w3159_ ;
	wire _w3158_ ;
	wire _w3157_ ;
	wire _w3156_ ;
	wire _w3155_ ;
	wire _w3154_ ;
	wire _w3153_ ;
	wire _w3152_ ;
	wire _w3151_ ;
	wire _w3150_ ;
	wire _w3149_ ;
	wire _w3148_ ;
	wire _w3147_ ;
	wire _w3146_ ;
	wire _w3145_ ;
	wire _w3144_ ;
	wire _w3143_ ;
	wire _w3142_ ;
	wire _w3141_ ;
	wire _w3140_ ;
	wire _w3139_ ;
	wire _w3138_ ;
	wire _w3137_ ;
	wire _w3136_ ;
	wire _w3135_ ;
	wire _w3134_ ;
	wire _w3133_ ;
	wire _w3132_ ;
	wire _w3131_ ;
	wire _w3130_ ;
	wire _w3129_ ;
	wire _w3128_ ;
	wire _w3127_ ;
	wire _w3126_ ;
	wire _w3125_ ;
	wire _w3124_ ;
	wire _w3123_ ;
	wire _w3122_ ;
	wire _w3121_ ;
	wire _w3120_ ;
	wire _w3119_ ;
	wire _w3118_ ;
	wire _w3117_ ;
	wire _w3116_ ;
	wire _w3115_ ;
	wire _w3114_ ;
	wire _w3113_ ;
	wire _w3112_ ;
	wire _w3111_ ;
	wire _w3110_ ;
	wire _w3109_ ;
	wire _w3108_ ;
	wire _w3107_ ;
	wire _w3106_ ;
	wire _w3105_ ;
	wire _w3104_ ;
	wire _w3103_ ;
	wire _w3102_ ;
	wire _w3101_ ;
	wire _w3100_ ;
	wire _w3099_ ;
	wire _w3098_ ;
	wire _w3097_ ;
	wire _w3096_ ;
	wire _w3095_ ;
	wire _w3094_ ;
	wire _w3093_ ;
	wire _w3092_ ;
	wire _w3091_ ;
	wire _w3090_ ;
	wire _w3089_ ;
	wire _w3088_ ;
	wire _w3087_ ;
	wire _w3086_ ;
	wire _w3085_ ;
	wire _w3084_ ;
	wire _w3083_ ;
	wire _w3082_ ;
	wire _w3081_ ;
	wire _w3080_ ;
	wire _w3079_ ;
	wire _w3078_ ;
	wire _w3077_ ;
	wire _w3076_ ;
	wire _w3075_ ;
	wire _w3074_ ;
	wire _w3073_ ;
	wire _w3072_ ;
	wire _w3071_ ;
	wire _w3070_ ;
	wire _w3069_ ;
	wire _w3068_ ;
	wire _w3067_ ;
	wire _w3066_ ;
	wire _w3065_ ;
	wire _w3064_ ;
	wire _w3063_ ;
	wire _w3062_ ;
	wire _w3061_ ;
	wire _w3060_ ;
	wire _w3059_ ;
	wire _w3058_ ;
	wire _w3057_ ;
	wire _w3056_ ;
	wire _w3055_ ;
	wire _w3054_ ;
	wire _w3053_ ;
	wire _w3052_ ;
	wire _w3051_ ;
	wire _w3050_ ;
	wire _w3049_ ;
	wire _w3048_ ;
	wire _w3047_ ;
	wire _w3046_ ;
	wire _w3045_ ;
	wire _w3044_ ;
	wire _w3043_ ;
	wire _w3042_ ;
	wire _w3041_ ;
	wire _w3040_ ;
	wire _w3039_ ;
	wire _w3038_ ;
	wire _w3037_ ;
	wire _w3036_ ;
	wire _w3035_ ;
	wire _w3034_ ;
	wire _w3033_ ;
	wire _w3032_ ;
	wire _w3031_ ;
	wire _w3030_ ;
	wire _w3029_ ;
	wire _w3028_ ;
	wire _w3027_ ;
	wire _w3026_ ;
	wire _w3025_ ;
	wire _w3024_ ;
	wire _w3023_ ;
	wire _w3022_ ;
	wire _w3021_ ;
	wire _w3020_ ;
	wire _w3019_ ;
	wire _w3018_ ;
	wire _w3017_ ;
	wire _w3016_ ;
	wire _w3015_ ;
	wire _w3014_ ;
	wire _w3013_ ;
	wire _w3012_ ;
	wire _w3011_ ;
	wire _w3010_ ;
	wire _w3009_ ;
	wire _w3008_ ;
	wire _w3007_ ;
	wire _w3006_ ;
	wire _w3005_ ;
	wire _w3004_ ;
	wire _w3003_ ;
	wire _w3002_ ;
	wire _w3001_ ;
	wire _w3000_ ;
	wire _w2999_ ;
	wire _w2998_ ;
	wire _w2997_ ;
	wire _w2996_ ;
	wire _w2995_ ;
	wire _w2994_ ;
	wire _w2993_ ;
	wire _w2992_ ;
	wire _w2991_ ;
	wire _w2990_ ;
	wire _w2989_ ;
	wire _w2988_ ;
	wire _w2987_ ;
	wire _w2986_ ;
	wire _w2985_ ;
	wire _w2984_ ;
	wire _w2983_ ;
	wire _w2982_ ;
	wire _w2981_ ;
	wire _w2980_ ;
	wire _w2979_ ;
	wire _w2978_ ;
	wire _w2977_ ;
	wire _w2976_ ;
	wire _w2975_ ;
	wire _w2974_ ;
	wire _w2973_ ;
	wire _w2972_ ;
	wire _w2971_ ;
	wire _w2970_ ;
	wire _w2969_ ;
	wire _w2968_ ;
	wire _w2967_ ;
	wire _w2966_ ;
	wire _w2965_ ;
	wire _w2964_ ;
	wire _w2963_ ;
	wire _w2962_ ;
	wire _w2961_ ;
	wire _w2960_ ;
	wire _w2959_ ;
	wire _w2958_ ;
	wire _w2957_ ;
	wire _w2956_ ;
	wire _w2955_ ;
	wire _w2954_ ;
	wire _w2953_ ;
	wire _w2952_ ;
	wire _w2951_ ;
	wire _w2950_ ;
	wire _w2949_ ;
	wire _w2948_ ;
	wire _w2947_ ;
	wire _w2946_ ;
	wire _w2945_ ;
	wire _w2944_ ;
	wire _w2943_ ;
	wire _w2942_ ;
	wire _w2941_ ;
	wire _w2940_ ;
	wire _w2939_ ;
	wire _w2938_ ;
	wire _w2937_ ;
	wire _w2936_ ;
	wire _w2935_ ;
	wire _w2934_ ;
	wire _w2933_ ;
	wire _w2932_ ;
	wire _w2931_ ;
	wire _w2930_ ;
	wire _w2929_ ;
	wire _w2928_ ;
	wire _w2927_ ;
	wire _w2926_ ;
	wire _w2925_ ;
	wire _w2924_ ;
	wire _w2923_ ;
	wire _w2922_ ;
	wire _w2921_ ;
	wire _w2920_ ;
	wire _w2919_ ;
	wire _w2918_ ;
	wire _w2917_ ;
	wire _w2916_ ;
	wire _w2915_ ;
	wire _w2914_ ;
	wire _w2913_ ;
	wire _w2912_ ;
	wire _w2911_ ;
	wire _w2910_ ;
	wire _w2909_ ;
	wire _w2908_ ;
	wire _w2907_ ;
	wire _w2906_ ;
	wire _w2905_ ;
	wire _w2904_ ;
	wire _w2903_ ;
	wire _w2902_ ;
	wire _w2901_ ;
	wire _w2900_ ;
	wire _w2899_ ;
	wire _w2898_ ;
	wire _w2897_ ;
	wire _w2896_ ;
	wire _w2895_ ;
	wire _w2894_ ;
	wire _w2893_ ;
	wire _w2892_ ;
	wire _w2891_ ;
	wire _w2890_ ;
	wire _w2889_ ;
	wire _w2888_ ;
	wire _w2887_ ;
	wire _w2886_ ;
	wire _w2885_ ;
	wire _w2884_ ;
	wire _w2883_ ;
	wire _w2882_ ;
	wire _w2881_ ;
	wire _w2880_ ;
	wire _w2879_ ;
	wire _w2878_ ;
	wire _w2877_ ;
	wire _w2876_ ;
	wire _w2875_ ;
	wire _w2874_ ;
	wire _w2873_ ;
	wire _w2872_ ;
	wire _w2871_ ;
	wire _w2870_ ;
	wire _w2869_ ;
	wire _w2868_ ;
	wire _w2867_ ;
	wire _w2866_ ;
	wire _w2865_ ;
	wire _w2864_ ;
	wire _w2863_ ;
	wire _w2862_ ;
	wire _w2861_ ;
	wire _w2860_ ;
	wire _w2859_ ;
	wire _w2858_ ;
	wire _w2857_ ;
	wire _w2856_ ;
	wire _w2855_ ;
	wire _w2854_ ;
	wire _w2853_ ;
	wire _w2852_ ;
	wire _w2851_ ;
	wire _w2850_ ;
	wire _w2849_ ;
	wire _w2848_ ;
	wire _w2847_ ;
	wire _w2846_ ;
	wire _w2845_ ;
	wire _w2844_ ;
	wire _w2843_ ;
	wire _w2842_ ;
	wire _w2841_ ;
	wire _w2840_ ;
	wire _w2839_ ;
	wire _w2838_ ;
	wire _w2837_ ;
	wire _w2836_ ;
	wire _w2835_ ;
	wire _w2834_ ;
	wire _w2833_ ;
	wire _w2832_ ;
	wire _w2831_ ;
	wire _w2830_ ;
	wire _w2829_ ;
	wire _w2828_ ;
	wire _w2827_ ;
	wire _w2826_ ;
	wire _w2825_ ;
	wire _w2824_ ;
	wire _w2823_ ;
	wire _w2822_ ;
	wire _w2821_ ;
	wire _w2820_ ;
	wire _w2819_ ;
	wire _w2818_ ;
	wire _w2817_ ;
	wire _w2816_ ;
	wire _w2815_ ;
	wire _w2814_ ;
	wire _w2813_ ;
	wire _w2812_ ;
	wire _w2811_ ;
	wire _w2810_ ;
	wire _w2809_ ;
	wire _w2808_ ;
	wire _w2807_ ;
	wire _w2806_ ;
	wire _w2805_ ;
	wire _w2804_ ;
	wire _w2803_ ;
	wire _w2802_ ;
	wire _w2801_ ;
	wire _w2800_ ;
	wire _w2799_ ;
	wire _w2798_ ;
	wire _w2797_ ;
	wire _w2796_ ;
	wire _w2795_ ;
	wire _w2794_ ;
	wire _w2793_ ;
	wire _w2792_ ;
	wire _w2791_ ;
	wire _w2790_ ;
	wire _w2789_ ;
	wire _w2788_ ;
	wire _w2787_ ;
	wire _w2786_ ;
	wire _w2785_ ;
	wire _w2784_ ;
	wire _w2783_ ;
	wire _w2782_ ;
	wire _w2781_ ;
	wire _w2780_ ;
	wire _w2779_ ;
	wire _w2778_ ;
	wire _w2777_ ;
	wire _w2776_ ;
	wire _w2775_ ;
	wire _w2774_ ;
	wire _w2773_ ;
	wire _w2772_ ;
	wire _w2771_ ;
	wire _w2770_ ;
	wire _w2769_ ;
	wire _w2768_ ;
	wire _w2767_ ;
	wire _w2766_ ;
	wire _w2765_ ;
	wire _w2764_ ;
	wire _w2763_ ;
	wire _w2762_ ;
	wire _w2761_ ;
	wire _w2760_ ;
	wire _w2759_ ;
	wire _w2758_ ;
	wire _w2757_ ;
	wire _w2756_ ;
	wire _w2755_ ;
	wire _w2754_ ;
	wire _w2753_ ;
	wire _w2752_ ;
	wire _w2751_ ;
	wire _w2750_ ;
	wire _w2749_ ;
	wire _w2748_ ;
	wire _w2747_ ;
	wire _w2746_ ;
	wire _w2745_ ;
	wire _w2744_ ;
	wire _w2743_ ;
	wire _w2742_ ;
	wire _w2741_ ;
	wire _w2740_ ;
	wire _w2739_ ;
	wire _w2738_ ;
	wire _w2737_ ;
	wire _w2736_ ;
	wire _w2735_ ;
	wire _w2734_ ;
	wire _w2733_ ;
	wire _w2732_ ;
	wire _w2731_ ;
	wire _w2730_ ;
	wire _w2729_ ;
	wire _w2728_ ;
	wire _w2727_ ;
	wire _w2726_ ;
	wire _w2725_ ;
	wire _w2724_ ;
	wire _w2723_ ;
	wire _w2722_ ;
	wire _w2721_ ;
	wire _w2720_ ;
	wire _w2719_ ;
	wire _w2718_ ;
	wire _w2717_ ;
	wire _w2716_ ;
	wire _w2715_ ;
	wire _w2714_ ;
	wire _w2713_ ;
	wire _w2712_ ;
	wire _w2711_ ;
	wire _w2710_ ;
	wire _w2709_ ;
	wire _w2708_ ;
	wire _w2707_ ;
	wire _w2706_ ;
	wire _w2705_ ;
	wire _w2704_ ;
	wire _w2703_ ;
	wire _w2702_ ;
	wire _w2701_ ;
	wire _w2700_ ;
	wire _w2699_ ;
	wire _w2698_ ;
	wire _w2697_ ;
	wire _w2696_ ;
	wire _w2695_ ;
	wire _w2694_ ;
	wire _w2693_ ;
	wire _w2692_ ;
	wire _w2691_ ;
	wire _w2690_ ;
	wire _w2689_ ;
	wire _w2688_ ;
	wire _w2687_ ;
	wire _w2686_ ;
	wire _w2685_ ;
	wire _w2684_ ;
	wire _w2683_ ;
	wire _w2682_ ;
	wire _w2681_ ;
	wire _w2680_ ;
	wire _w2679_ ;
	wire _w2678_ ;
	wire _w2677_ ;
	wire _w2676_ ;
	wire _w2675_ ;
	wire _w2674_ ;
	wire _w2673_ ;
	wire _w2672_ ;
	wire _w2671_ ;
	wire _w2670_ ;
	wire _w2669_ ;
	wire _w2668_ ;
	wire _w2667_ ;
	wire _w2666_ ;
	wire _w2665_ ;
	wire _w2664_ ;
	wire _w2663_ ;
	wire _w2662_ ;
	wire _w2661_ ;
	wire _w2660_ ;
	wire _w2659_ ;
	wire _w2658_ ;
	wire _w2657_ ;
	wire _w2656_ ;
	wire _w2655_ ;
	wire _w2654_ ;
	wire _w2653_ ;
	wire _w2652_ ;
	wire _w2651_ ;
	wire _w2650_ ;
	wire _w2649_ ;
	wire _w2648_ ;
	wire _w2647_ ;
	wire _w2646_ ;
	wire _w2645_ ;
	wire _w2644_ ;
	wire _w2643_ ;
	wire _w2642_ ;
	wire _w2641_ ;
	wire _w2640_ ;
	wire _w2639_ ;
	wire _w2638_ ;
	wire _w2637_ ;
	wire _w2636_ ;
	wire _w2635_ ;
	wire _w2634_ ;
	wire _w2633_ ;
	wire _w2632_ ;
	wire _w2631_ ;
	wire _w2630_ ;
	wire _w2629_ ;
	wire _w2628_ ;
	wire _w2627_ ;
	wire _w2626_ ;
	wire _w2625_ ;
	wire _w2624_ ;
	wire _w2623_ ;
	wire _w2622_ ;
	wire _w2621_ ;
	wire _w2620_ ;
	wire _w2619_ ;
	wire _w2618_ ;
	wire _w2617_ ;
	wire _w2048_ ;
	wire _w2047_ ;
	wire _w2046_ ;
	wire _w2045_ ;
	wire _w2044_ ;
	wire _w2043_ ;
	wire _w2042_ ;
	wire _w2041_ ;
	wire _w2040_ ;
	wire _w2039_ ;
	wire _w2038_ ;
	wire _w2037_ ;
	wire _w2036_ ;
	wire _w2035_ ;
	wire _w2034_ ;
	wire _w2033_ ;
	wire _w2032_ ;
	wire _w2031_ ;
	wire _w2030_ ;
	wire _w2029_ ;
	wire _w2028_ ;
	wire _w2027_ ;
	wire _w2026_ ;
	wire _w2025_ ;
	wire _w2024_ ;
	wire _w2023_ ;
	wire _w2022_ ;
	wire _w2021_ ;
	wire _w2020_ ;
	wire _w2019_ ;
	wire _w2018_ ;
	wire _w2017_ ;
	wire _w2016_ ;
	wire _w2015_ ;
	wire _w2014_ ;
	wire _w2013_ ;
	wire _w2012_ ;
	wire _w2011_ ;
	wire _w2010_ ;
	wire _w2009_ ;
	wire _w2008_ ;
	wire _w2007_ ;
	wire _w2006_ ;
	wire _w2005_ ;
	wire _w2004_ ;
	wire _w2003_ ;
	wire _w2002_ ;
	wire _w2001_ ;
	wire _w2000_ ;
	wire _w1999_ ;
	wire _w1998_ ;
	wire _w1997_ ;
	wire _w1996_ ;
	wire _w1995_ ;
	wire _w1994_ ;
	wire _w1993_ ;
	wire _w1992_ ;
	wire _w1991_ ;
	wire _w1990_ ;
	wire _w1989_ ;
	wire _w1988_ ;
	wire _w1987_ ;
	wire _w1986_ ;
	wire _w1985_ ;
	wire _w1984_ ;
	wire _w1983_ ;
	wire _w1982_ ;
	wire _w1981_ ;
	wire _w1980_ ;
	wire _w1979_ ;
	wire _w1978_ ;
	wire _w1977_ ;
	wire _w1976_ ;
	wire _w1975_ ;
	wire _w1974_ ;
	wire _w1973_ ;
	wire _w1972_ ;
	wire _w1971_ ;
	wire _w1970_ ;
	wire _w1969_ ;
	wire _w1968_ ;
	wire _w1967_ ;
	wire _w1966_ ;
	wire _w1965_ ;
	wire _w1964_ ;
	wire _w1963_ ;
	wire _w1962_ ;
	wire _w1961_ ;
	wire _w1960_ ;
	wire _w1959_ ;
	wire _w1958_ ;
	wire _w1957_ ;
	wire _w1956_ ;
	wire _w1955_ ;
	wire _w1954_ ;
	wire _w1953_ ;
	wire _w1952_ ;
	wire _w1951_ ;
	wire _w1950_ ;
	wire _w1949_ ;
	wire _w1948_ ;
	wire _w1947_ ;
	wire _w1946_ ;
	wire _w1945_ ;
	wire _w1944_ ;
	wire _w1943_ ;
	wire _w1942_ ;
	wire _w1941_ ;
	wire _w1940_ ;
	wire _w1939_ ;
	wire _w1938_ ;
	wire _w1937_ ;
	wire _w1936_ ;
	wire _w1935_ ;
	wire _w1934_ ;
	wire _w1933_ ;
	wire _w1932_ ;
	wire _w1931_ ;
	wire _w1930_ ;
	wire _w1929_ ;
	wire _w1928_ ;
	wire _w1927_ ;
	wire _w1926_ ;
	wire _w1925_ ;
	wire _w1924_ ;
	wire _w1923_ ;
	wire _w1922_ ;
	wire _w1921_ ;
	wire _w1920_ ;
	wire _w1919_ ;
	wire _w1918_ ;
	wire _w1917_ ;
	wire _w1916_ ;
	wire _w1915_ ;
	wire _w1914_ ;
	wire _w1913_ ;
	wire _w1912_ ;
	wire _w1911_ ;
	wire _w1910_ ;
	wire _w1909_ ;
	wire _w1908_ ;
	wire _w1907_ ;
	wire _w1906_ ;
	wire _w1905_ ;
	wire _w1904_ ;
	wire _w1903_ ;
	wire _w1902_ ;
	wire _w1901_ ;
	wire _w1900_ ;
	wire _w1899_ ;
	wire _w1898_ ;
	wire _w1897_ ;
	wire _w1896_ ;
	wire _w1895_ ;
	wire _w1894_ ;
	wire _w1893_ ;
	wire _w1892_ ;
	wire _w1891_ ;
	wire _w1890_ ;
	wire _w1889_ ;
	wire _w1888_ ;
	wire _w1887_ ;
	wire _w1886_ ;
	wire _w1885_ ;
	wire _w1884_ ;
	wire _w1883_ ;
	wire _w1882_ ;
	wire _w1881_ ;
	wire _w1880_ ;
	wire _w1879_ ;
	wire _w1878_ ;
	wire _w1877_ ;
	wire _w1876_ ;
	wire _w1875_ ;
	wire _w1874_ ;
	wire _w1873_ ;
	wire _w1872_ ;
	wire _w1871_ ;
	wire _w1870_ ;
	wire _w1869_ ;
	wire _w1868_ ;
	wire _w1867_ ;
	wire _w1866_ ;
	wire _w1865_ ;
	wire _w1864_ ;
	wire _w1863_ ;
	wire _w1862_ ;
	wire _w1861_ ;
	wire _w1860_ ;
	wire _w1859_ ;
	wire _w1858_ ;
	wire _w1857_ ;
	wire _w1856_ ;
	wire _w1855_ ;
	wire _w1854_ ;
	wire _w1853_ ;
	wire _w1852_ ;
	wire _w1851_ ;
	wire _w1850_ ;
	wire _w1849_ ;
	wire _w1848_ ;
	wire _w1847_ ;
	wire _w1846_ ;
	wire _w1845_ ;
	wire _w1844_ ;
	wire _w1843_ ;
	wire _w1842_ ;
	wire _w1841_ ;
	wire _w1840_ ;
	wire _w1839_ ;
	wire _w1838_ ;
	wire _w1837_ ;
	wire _w1836_ ;
	wire _w1835_ ;
	wire _w1834_ ;
	wire _w1833_ ;
	wire _w1832_ ;
	wire _w1831_ ;
	wire _w1830_ ;
	wire _w1829_ ;
	wire _w1828_ ;
	wire _w1827_ ;
	wire _w1826_ ;
	wire _w1825_ ;
	wire _w1824_ ;
	wire _w1823_ ;
	wire _w1822_ ;
	wire _w1821_ ;
	wire _w1820_ ;
	wire _w1819_ ;
	wire _w1818_ ;
	wire _w1817_ ;
	wire _w1816_ ;
	wire _w1815_ ;
	wire _w1814_ ;
	wire _w1813_ ;
	wire _w1812_ ;
	wire _w1811_ ;
	wire _w1810_ ;
	wire _w1809_ ;
	wire _w1808_ ;
	wire _w1807_ ;
	wire _w1806_ ;
	wire _w1805_ ;
	wire _w1804_ ;
	wire _w1803_ ;
	wire _w1802_ ;
	wire _w1801_ ;
	wire _w1800_ ;
	wire _w1799_ ;
	wire _w1798_ ;
	wire _w1797_ ;
	wire _w1796_ ;
	wire _w1795_ ;
	wire _w1794_ ;
	wire _w1793_ ;
	wire _w1792_ ;
	wire _w1791_ ;
	wire _w1790_ ;
	wire _w1789_ ;
	wire _w1788_ ;
	wire _w1787_ ;
	wire _w1786_ ;
	wire _w1785_ ;
	wire _w1784_ ;
	wire _w1783_ ;
	wire _w1782_ ;
	wire _w1781_ ;
	wire _w1780_ ;
	wire _w1779_ ;
	wire _w1778_ ;
	wire _w1777_ ;
	wire _w1776_ ;
	wire _w1775_ ;
	wire _w1774_ ;
	wire _w1773_ ;
	wire _w1772_ ;
	wire _w1771_ ;
	wire _w1770_ ;
	wire _w1769_ ;
	wire _w1768_ ;
	wire _w1767_ ;
	wire _w1766_ ;
	wire _w1765_ ;
	wire _w1634_ ;
	wire _w1633_ ;
	wire _w1632_ ;
	wire _w1631_ ;
	wire _w1630_ ;
	wire _w1629_ ;
	wire _w1628_ ;
	wire _w1627_ ;
	wire _w1626_ ;
	wire _w1625_ ;
	wire _w1624_ ;
	wire _w1623_ ;
	wire _w1622_ ;
	wire _w1621_ ;
	wire _w1620_ ;
	wire _w1619_ ;
	wire _w1618_ ;
	wire _w1617_ ;
	wire _w1616_ ;
	wire _w1615_ ;
	wire _w1614_ ;
	wire _w1613_ ;
	wire _w1612_ ;
	wire _w1611_ ;
	wire _w1610_ ;
	wire _w1609_ ;
	wire _w1608_ ;
	wire _w1607_ ;
	wire _w1606_ ;
	wire _w1605_ ;
	wire _w1604_ ;
	wire _w1603_ ;
	wire _w1602_ ;
	wire _w1601_ ;
	wire _w1600_ ;
	wire _w1599_ ;
	wire _w1598_ ;
	wire _w1597_ ;
	wire _w1596_ ;
	wire _w1595_ ;
	wire _w1594_ ;
	wire _w1593_ ;
	wire _w1592_ ;
	wire _w1591_ ;
	wire _w1590_ ;
	wire _w1589_ ;
	wire _w1588_ ;
	wire _w1587_ ;
	wire _w1586_ ;
	wire _w1585_ ;
	wire _w1584_ ;
	wire _w1583_ ;
	wire _w1582_ ;
	wire _w1581_ ;
	wire _w1580_ ;
	wire _w1579_ ;
	wire _w1578_ ;
	wire _w1577_ ;
	wire _w1576_ ;
	wire _w1575_ ;
	wire _w1574_ ;
	wire _w1573_ ;
	wire _w1572_ ;
	wire _w1571_ ;
	wire _w1570_ ;
	wire _w1569_ ;
	wire _w1568_ ;
	wire _w1567_ ;
	wire _w1536_ ;
	wire _w1535_ ;
	wire _w1534_ ;
	wire _w1533_ ;
	wire _w1532_ ;
	wire _w1531_ ;
	wire _w1530_ ;
	wire _w1529_ ;
	wire _w1528_ ;
	wire _w1527_ ;
	wire _w1526_ ;
	wire _w1525_ ;
	wire _w1524_ ;
	wire _w1523_ ;
	wire _w1522_ ;
	wire _w1521_ ;
	wire _w1508_ ;
	wire _w1509_ ;
	wire _w1510_ ;
	wire _w1511_ ;
	wire _w1512_ ;
	wire _w1513_ ;
	wire _w1514_ ;
	wire _w1515_ ;
	wire _w1516_ ;
	wire _w1517_ ;
	wire _w1518_ ;
	wire _w1519_ ;
	wire _w1520_ ;
	wire _w1537_ ;
	wire _w1538_ ;
	wire _w1539_ ;
	wire _w1540_ ;
	wire _w1541_ ;
	wire _w1542_ ;
	wire _w1543_ ;
	wire _w1544_ ;
	wire _w1545_ ;
	wire _w1546_ ;
	wire _w1547_ ;
	wire _w1548_ ;
	wire _w1549_ ;
	wire _w1550_ ;
	wire _w1551_ ;
	wire _w1552_ ;
	wire _w1553_ ;
	wire _w1554_ ;
	wire _w1555_ ;
	wire _w1556_ ;
	wire _w1557_ ;
	wire _w1558_ ;
	wire _w1559_ ;
	wire _w1560_ ;
	wire _w1561_ ;
	wire _w1562_ ;
	wire _w1563_ ;
	wire _w1564_ ;
	wire _w1565_ ;
	wire _w1566_ ;
	wire _w1635_ ;
	wire _w1636_ ;
	wire _w1637_ ;
	wire _w1638_ ;
	wire _w1639_ ;
	wire _w1640_ ;
	wire _w1641_ ;
	wire _w1642_ ;
	wire _w1643_ ;
	wire _w1644_ ;
	wire _w1645_ ;
	wire _w1646_ ;
	wire _w1647_ ;
	wire _w1648_ ;
	wire _w1649_ ;
	wire _w1650_ ;
	wire _w1651_ ;
	wire _w1652_ ;
	wire _w1653_ ;
	wire _w1654_ ;
	wire _w1655_ ;
	wire _w1656_ ;
	wire _w1657_ ;
	wire _w1658_ ;
	wire _w1659_ ;
	wire _w1660_ ;
	wire _w1661_ ;
	wire _w1662_ ;
	wire _w1663_ ;
	wire _w1664_ ;
	wire _w1665_ ;
	wire _w1666_ ;
	wire _w1667_ ;
	wire _w1668_ ;
	wire _w1669_ ;
	wire _w1670_ ;
	wire _w1671_ ;
	wire _w1672_ ;
	wire _w1673_ ;
	wire _w1674_ ;
	wire _w1675_ ;
	wire _w1676_ ;
	wire _w1677_ ;
	wire _w1678_ ;
	wire _w1679_ ;
	wire _w1680_ ;
	wire _w1681_ ;
	wire _w1682_ ;
	wire _w1683_ ;
	wire _w1684_ ;
	wire _w1685_ ;
	wire _w1686_ ;
	wire _w1687_ ;
	wire _w1688_ ;
	wire _w1689_ ;
	wire _w1690_ ;
	wire _w1691_ ;
	wire _w1692_ ;
	wire _w1693_ ;
	wire _w1694_ ;
	wire _w1695_ ;
	wire _w1696_ ;
	wire _w1697_ ;
	wire _w1698_ ;
	wire _w1699_ ;
	wire _w1700_ ;
	wire _w1701_ ;
	wire _w1702_ ;
	wire _w1703_ ;
	wire _w1704_ ;
	wire _w1705_ ;
	wire _w1706_ ;
	wire _w1707_ ;
	wire _w1708_ ;
	wire _w1709_ ;
	wire _w1710_ ;
	wire _w1711_ ;
	wire _w1712_ ;
	wire _w1713_ ;
	wire _w1714_ ;
	wire _w1715_ ;
	wire _w1716_ ;
	wire _w1717_ ;
	wire _w1718_ ;
	wire _w1719_ ;
	wire _w1720_ ;
	wire _w1721_ ;
	wire _w1722_ ;
	wire _w1723_ ;
	wire _w1724_ ;
	wire _w1725_ ;
	wire _w1726_ ;
	wire _w1727_ ;
	wire _w1728_ ;
	wire _w1729_ ;
	wire _w1730_ ;
	wire _w1731_ ;
	wire _w1732_ ;
	wire _w1733_ ;
	wire _w1734_ ;
	wire _w1735_ ;
	wire _w1736_ ;
	wire _w1737_ ;
	wire _w1738_ ;
	wire _w1739_ ;
	wire _w1740_ ;
	wire _w1741_ ;
	wire _w1742_ ;
	wire _w1743_ ;
	wire _w1744_ ;
	wire _w1745_ ;
	wire _w1746_ ;
	wire _w1747_ ;
	wire _w1748_ ;
	wire _w1749_ ;
	wire _w1750_ ;
	wire _w1751_ ;
	wire _w1752_ ;
	wire _w1753_ ;
	wire _w1754_ ;
	wire _w1755_ ;
	wire _w1756_ ;
	wire _w1757_ ;
	wire _w1758_ ;
	wire _w1759_ ;
	wire _w1760_ ;
	wire _w1761_ ;
	wire _w1762_ ;
	wire _w1763_ ;
	wire _w1764_ ;
	wire _w2049_ ;
	wire _w2050_ ;
	wire _w2051_ ;
	wire _w2052_ ;
	wire _w2053_ ;
	wire _w2054_ ;
	wire _w2055_ ;
	wire _w2056_ ;
	wire _w2057_ ;
	wire _w2058_ ;
	wire _w2059_ ;
	wire _w2060_ ;
	wire _w2061_ ;
	wire _w2062_ ;
	wire _w2063_ ;
	wire _w2064_ ;
	wire _w2065_ ;
	wire _w2066_ ;
	wire _w2067_ ;
	wire _w2068_ ;
	wire _w2069_ ;
	wire _w2070_ ;
	wire _w2071_ ;
	wire _w2072_ ;
	wire _w2073_ ;
	wire _w2074_ ;
	wire _w2075_ ;
	wire _w2076_ ;
	wire _w2077_ ;
	wire _w2078_ ;
	wire _w2079_ ;
	wire _w2080_ ;
	wire _w2081_ ;
	wire _w2082_ ;
	wire _w2083_ ;
	wire _w2084_ ;
	wire _w2085_ ;
	wire _w2086_ ;
	wire _w2087_ ;
	wire _w2088_ ;
	wire _w2089_ ;
	wire _w2090_ ;
	wire _w2091_ ;
	wire _w2092_ ;
	wire _w2093_ ;
	wire _w2094_ ;
	wire _w2095_ ;
	wire _w2096_ ;
	wire _w2097_ ;
	wire _w2098_ ;
	wire _w2099_ ;
	wire _w2100_ ;
	wire _w2101_ ;
	wire _w2102_ ;
	wire _w2103_ ;
	wire _w2104_ ;
	wire _w2105_ ;
	wire _w2106_ ;
	wire _w2107_ ;
	wire _w2108_ ;
	wire _w2109_ ;
	wire _w2110_ ;
	wire _w2111_ ;
	wire _w2112_ ;
	wire _w2113_ ;
	wire _w2114_ ;
	wire _w2115_ ;
	wire _w2116_ ;
	wire _w2117_ ;
	wire _w2118_ ;
	wire _w2119_ ;
	wire _w2120_ ;
	wire _w2121_ ;
	wire _w2122_ ;
	wire _w2123_ ;
	wire _w2124_ ;
	wire _w2125_ ;
	wire _w2126_ ;
	wire _w2127_ ;
	wire _w2128_ ;
	wire _w2129_ ;
	wire _w2130_ ;
	wire _w2131_ ;
	wire _w2132_ ;
	wire _w2133_ ;
	wire _w2134_ ;
	wire _w2135_ ;
	wire _w2136_ ;
	wire _w2137_ ;
	wire _w2138_ ;
	wire _w2139_ ;
	wire _w2140_ ;
	wire _w2141_ ;
	wire _w2142_ ;
	wire _w2143_ ;
	wire _w2144_ ;
	wire _w2145_ ;
	wire _w2146_ ;
	wire _w2147_ ;
	wire _w2148_ ;
	wire _w2149_ ;
	wire _w2150_ ;
	wire _w2151_ ;
	wire _w2152_ ;
	wire _w2153_ ;
	wire _w2154_ ;
	wire _w2155_ ;
	wire _w2156_ ;
	wire _w2157_ ;
	wire _w2158_ ;
	wire _w2159_ ;
	wire _w2160_ ;
	wire _w2161_ ;
	wire _w2162_ ;
	wire _w2163_ ;
	wire _w2164_ ;
	wire _w2165_ ;
	wire _w2166_ ;
	wire _w2167_ ;
	wire _w2168_ ;
	wire _w2169_ ;
	wire _w2170_ ;
	wire _w2171_ ;
	wire _w2172_ ;
	wire _w2173_ ;
	wire _w2174_ ;
	wire _w2175_ ;
	wire _w2176_ ;
	wire _w2177_ ;
	wire _w2178_ ;
	wire _w2179_ ;
	wire _w2180_ ;
	wire _w2181_ ;
	wire _w2182_ ;
	wire _w2183_ ;
	wire _w2184_ ;
	wire _w2185_ ;
	wire _w2186_ ;
	wire _w2187_ ;
	wire _w2188_ ;
	wire _w2189_ ;
	wire _w2190_ ;
	wire _w2191_ ;
	wire _w2192_ ;
	wire _w2193_ ;
	wire _w2194_ ;
	wire _w2195_ ;
	wire _w2196_ ;
	wire _w2197_ ;
	wire _w2198_ ;
	wire _w2199_ ;
	wire _w2200_ ;
	wire _w2201_ ;
	wire _w2202_ ;
	wire _w2203_ ;
	wire _w2204_ ;
	wire _w2205_ ;
	wire _w2206_ ;
	wire _w2207_ ;
	wire _w2208_ ;
	wire _w2209_ ;
	wire _w2210_ ;
	wire _w2211_ ;
	wire _w2212_ ;
	wire _w2213_ ;
	wire _w2214_ ;
	wire _w2215_ ;
	wire _w2216_ ;
	wire _w2217_ ;
	wire _w2218_ ;
	wire _w2219_ ;
	wire _w2220_ ;
	wire _w2221_ ;
	wire _w2222_ ;
	wire _w2223_ ;
	wire _w2224_ ;
	wire _w2225_ ;
	wire _w2226_ ;
	wire _w2227_ ;
	wire _w2228_ ;
	wire _w2229_ ;
	wire _w2230_ ;
	wire _w2231_ ;
	wire _w2232_ ;
	wire _w2233_ ;
	wire _w2234_ ;
	wire _w2235_ ;
	wire _w2236_ ;
	wire _w2237_ ;
	wire _w2238_ ;
	wire _w2239_ ;
	wire _w2240_ ;
	wire _w2241_ ;
	wire _w2242_ ;
	wire _w2243_ ;
	wire _w2244_ ;
	wire _w2245_ ;
	wire _w2246_ ;
	wire _w2247_ ;
	wire _w2248_ ;
	wire _w2249_ ;
	wire _w2250_ ;
	wire _w2251_ ;
	wire _w2252_ ;
	wire _w2253_ ;
	wire _w2254_ ;
	wire _w2255_ ;
	wire _w2256_ ;
	wire _w2257_ ;
	wire _w2258_ ;
	wire _w2259_ ;
	wire _w2260_ ;
	wire _w2261_ ;
	wire _w2262_ ;
	wire _w2263_ ;
	wire _w2264_ ;
	wire _w2265_ ;
	wire _w2266_ ;
	wire _w2267_ ;
	wire _w2268_ ;
	wire _w2269_ ;
	wire _w2270_ ;
	wire _w2271_ ;
	wire _w2272_ ;
	wire _w2273_ ;
	wire _w2274_ ;
	wire _w2275_ ;
	wire _w2276_ ;
	wire _w2277_ ;
	wire _w2278_ ;
	wire _w2279_ ;
	wire _w2280_ ;
	wire _w2281_ ;
	wire _w2282_ ;
	wire _w2283_ ;
	wire _w2284_ ;
	wire _w2285_ ;
	wire _w2286_ ;
	wire _w2287_ ;
	wire _w2288_ ;
	wire _w2289_ ;
	wire _w2290_ ;
	wire _w2291_ ;
	wire _w2292_ ;
	wire _w2293_ ;
	wire _w2294_ ;
	wire _w2295_ ;
	wire _w2296_ ;
	wire _w2297_ ;
	wire _w2298_ ;
	wire _w2299_ ;
	wire _w2300_ ;
	wire _w2301_ ;
	wire _w2302_ ;
	wire _w2303_ ;
	wire _w2304_ ;
	wire _w2305_ ;
	wire _w2306_ ;
	wire _w2307_ ;
	wire _w2308_ ;
	wire _w2309_ ;
	wire _w2310_ ;
	wire _w2311_ ;
	wire _w2312_ ;
	wire _w2313_ ;
	wire _w2314_ ;
	wire _w2315_ ;
	wire _w2316_ ;
	wire _w2317_ ;
	wire _w2318_ ;
	wire _w2319_ ;
	wire _w2320_ ;
	wire _w2321_ ;
	wire _w2322_ ;
	wire _w2323_ ;
	wire _w2324_ ;
	wire _w2325_ ;
	wire _w2326_ ;
	wire _w2327_ ;
	wire _w2328_ ;
	wire _w2329_ ;
	wire _w2330_ ;
	wire _w2331_ ;
	wire _w2332_ ;
	wire _w2333_ ;
	wire _w2334_ ;
	wire _w2335_ ;
	wire _w2336_ ;
	wire _w2337_ ;
	wire _w2338_ ;
	wire _w2339_ ;
	wire _w2340_ ;
	wire _w2341_ ;
	wire _w2342_ ;
	wire _w2343_ ;
	wire _w2344_ ;
	wire _w2345_ ;
	wire _w2346_ ;
	wire _w2347_ ;
	wire _w2348_ ;
	wire _w2349_ ;
	wire _w2350_ ;
	wire _w2351_ ;
	wire _w2352_ ;
	wire _w2353_ ;
	wire _w2354_ ;
	wire _w2355_ ;
	wire _w2356_ ;
	wire _w2357_ ;
	wire _w2358_ ;
	wire _w2359_ ;
	wire _w2360_ ;
	wire _w2361_ ;
	wire _w2362_ ;
	wire _w2363_ ;
	wire _w2364_ ;
	wire _w2365_ ;
	wire _w2366_ ;
	wire _w2367_ ;
	wire _w2368_ ;
	wire _w2369_ ;
	wire _w2370_ ;
	wire _w2371_ ;
	wire _w2372_ ;
	wire _w2373_ ;
	wire _w2374_ ;
	wire _w2375_ ;
	wire _w2376_ ;
	wire _w2377_ ;
	wire _w2378_ ;
	wire _w2379_ ;
	wire _w2380_ ;
	wire _w2381_ ;
	wire _w2382_ ;
	wire _w2383_ ;
	wire _w2384_ ;
	wire _w2385_ ;
	wire _w2386_ ;
	wire _w2387_ ;
	wire _w2388_ ;
	wire _w2389_ ;
	wire _w2390_ ;
	wire _w2391_ ;
	wire _w2392_ ;
	wire _w2393_ ;
	wire _w2394_ ;
	wire _w2395_ ;
	wire _w2396_ ;
	wire _w2397_ ;
	wire _w2398_ ;
	wire _w2399_ ;
	wire _w2400_ ;
	wire _w2401_ ;
	wire _w2402_ ;
	wire _w2403_ ;
	wire _w2404_ ;
	wire _w2405_ ;
	wire _w2406_ ;
	wire _w2407_ ;
	wire _w2408_ ;
	wire _w2409_ ;
	wire _w2410_ ;
	wire _w2411_ ;
	wire _w2412_ ;
	wire _w2413_ ;
	wire _w2414_ ;
	wire _w2415_ ;
	wire _w2416_ ;
	wire _w2417_ ;
	wire _w2418_ ;
	wire _w2419_ ;
	wire _w2420_ ;
	wire _w2421_ ;
	wire _w2422_ ;
	wire _w2423_ ;
	wire _w2424_ ;
	wire _w2425_ ;
	wire _w2426_ ;
	wire _w2427_ ;
	wire _w2428_ ;
	wire _w2429_ ;
	wire _w2430_ ;
	wire _w2431_ ;
	wire _w2432_ ;
	wire _w2433_ ;
	wire _w2434_ ;
	wire _w2435_ ;
	wire _w2436_ ;
	wire _w2437_ ;
	wire _w2438_ ;
	wire _w2439_ ;
	wire _w2440_ ;
	wire _w2441_ ;
	wire _w2442_ ;
	wire _w2443_ ;
	wire _w2444_ ;
	wire _w2445_ ;
	wire _w2446_ ;
	wire _w2447_ ;
	wire _w2448_ ;
	wire _w2449_ ;
	wire _w2450_ ;
	wire _w2451_ ;
	wire _w2452_ ;
	wire _w2453_ ;
	wire _w2454_ ;
	wire _w2455_ ;
	wire _w2456_ ;
	wire _w2457_ ;
	wire _w2458_ ;
	wire _w2459_ ;
	wire _w2460_ ;
	wire _w2461_ ;
	wire _w2462_ ;
	wire _w2463_ ;
	wire _w2464_ ;
	wire _w2465_ ;
	wire _w2466_ ;
	wire _w2467_ ;
	wire _w2468_ ;
	wire _w2469_ ;
	wire _w2470_ ;
	wire _w2471_ ;
	wire _w2472_ ;
	wire _w2473_ ;
	wire _w2474_ ;
	wire _w2475_ ;
	wire _w2476_ ;
	wire _w2477_ ;
	wire _w2478_ ;
	wire _w2479_ ;
	wire _w2480_ ;
	wire _w2481_ ;
	wire _w2482_ ;
	wire _w2483_ ;
	wire _w2484_ ;
	wire _w2485_ ;
	wire _w2486_ ;
	wire _w2487_ ;
	wire _w2488_ ;
	wire _w2489_ ;
	wire _w2490_ ;
	wire _w2491_ ;
	wire _w2492_ ;
	wire _w2493_ ;
	wire _w2494_ ;
	wire _w2495_ ;
	wire _w2496_ ;
	wire _w2497_ ;
	wire _w2498_ ;
	wire _w2499_ ;
	wire _w2500_ ;
	wire _w2501_ ;
	wire _w2502_ ;
	wire _w2503_ ;
	wire _w2504_ ;
	wire _w2505_ ;
	wire _w2506_ ;
	wire _w2507_ ;
	wire _w2508_ ;
	wire _w2509_ ;
	wire _w2510_ ;
	wire _w2511_ ;
	wire _w2512_ ;
	wire _w2513_ ;
	wire _w2514_ ;
	wire _w2515_ ;
	wire _w2516_ ;
	wire _w2517_ ;
	wire _w2518_ ;
	wire _w2519_ ;
	wire _w2520_ ;
	wire _w2521_ ;
	wire _w2522_ ;
	wire _w2523_ ;
	wire _w2524_ ;
	wire _w2525_ ;
	wire _w2526_ ;
	wire _w2527_ ;
	wire _w2528_ ;
	wire _w2529_ ;
	wire _w2530_ ;
	wire _w2531_ ;
	wire _w2532_ ;
	wire _w2533_ ;
	wire _w2534_ ;
	wire _w2535_ ;
	wire _w2536_ ;
	wire _w2537_ ;
	wire _w2538_ ;
	wire _w2539_ ;
	wire _w2540_ ;
	wire _w2541_ ;
	wire _w2542_ ;
	wire _w2543_ ;
	wire _w2544_ ;
	wire _w2545_ ;
	wire _w2546_ ;
	wire _w2547_ ;
	wire _w2548_ ;
	wire _w2549_ ;
	wire _w2550_ ;
	wire _w2551_ ;
	wire _w2552_ ;
	wire _w2553_ ;
	wire _w2554_ ;
	wire _w2555_ ;
	wire _w2556_ ;
	wire _w2557_ ;
	wire _w2558_ ;
	wire _w2559_ ;
	wire _w2560_ ;
	wire _w2561_ ;
	wire _w2562_ ;
	wire _w2563_ ;
	wire _w2564_ ;
	wire _w2565_ ;
	wire _w2566_ ;
	wire _w2567_ ;
	wire _w2568_ ;
	wire _w2569_ ;
	wire _w2570_ ;
	wire _w2571_ ;
	wire _w2572_ ;
	wire _w2573_ ;
	wire _w2574_ ;
	wire _w2575_ ;
	wire _w2576_ ;
	wire _w2577_ ;
	wire _w2578_ ;
	wire _w2579_ ;
	wire _w2580_ ;
	wire _w2581_ ;
	wire _w2582_ ;
	wire _w2583_ ;
	wire _w2584_ ;
	wire _w2585_ ;
	wire _w2586_ ;
	wire _w2587_ ;
	wire _w2588_ ;
	wire _w2589_ ;
	wire _w2590_ ;
	wire _w2591_ ;
	wire _w2592_ ;
	wire _w2593_ ;
	wire _w2594_ ;
	wire _w2595_ ;
	wire _w2596_ ;
	wire _w2597_ ;
	wire _w2598_ ;
	wire _w2599_ ;
	wire _w2600_ ;
	wire _w2601_ ;
	wire _w2602_ ;
	wire _w2603_ ;
	wire _w2604_ ;
	wire _w2605_ ;
	wire _w2606_ ;
	wire _w2607_ ;
	wire _w2608_ ;
	wire _w2609_ ;
	wire _w2610_ ;
	wire _w2611_ ;
	wire _w2612_ ;
	wire _w2613_ ;
	wire _w2614_ ;
	wire _w2615_ ;
	wire _w2616_ ;
	wire _w3865_ ;
	wire _w3866_ ;
	wire _w3867_ ;
	wire _w3868_ ;
	wire _w3869_ ;
	wire _w3870_ ;
	wire _w3871_ ;
	wire _w3872_ ;
	wire _w3873_ ;
	wire _w3874_ ;
	wire _w3875_ ;
	wire _w3876_ ;
	wire _w3877_ ;
	wire _w3878_ ;
	wire _w3879_ ;
	wire _w3880_ ;
	wire _w3881_ ;
	wire _w3882_ ;
	wire _w3883_ ;
	wire _w3884_ ;
	wire _w3885_ ;
	wire _w3886_ ;
	wire _w3887_ ;
	wire _w3888_ ;
	wire _w3889_ ;
	wire _w3890_ ;
	wire _w3891_ ;
	wire _w3892_ ;
	wire _w3893_ ;
	wire _w3894_ ;
	wire _w3895_ ;
	wire _w3896_ ;
	wire _w3897_ ;
	wire _w3898_ ;
	wire _w3899_ ;
	wire _w3900_ ;
	wire _w3901_ ;
	wire _w3902_ ;
	wire _w3903_ ;
	wire _w3904_ ;
	wire _w3905_ ;
	wire _w3906_ ;
	wire _w3907_ ;
	wire _w3908_ ;
	wire _w3909_ ;
	wire _w3910_ ;
	wire _w3911_ ;
	wire _w3912_ ;
	wire _w3913_ ;
	wire _w3914_ ;
	wire _w3915_ ;
	wire _w3916_ ;
	wire _w3917_ ;
	wire _w3918_ ;
	wire _w3919_ ;
	wire _w3920_ ;
	wire _w3921_ ;
	wire _w3922_ ;
	wire _w3923_ ;
	wire _w3924_ ;
	wire _w3925_ ;
	wire _w3926_ ;
	wire _w3927_ ;
	wire _w3928_ ;
	wire _w3929_ ;
	wire _w3930_ ;
	wire _w3931_ ;
	wire _w3932_ ;
	wire _w3933_ ;
	wire _w3934_ ;
	wire _w3935_ ;
	wire _w3936_ ;
	wire _w3937_ ;
	wire _w3938_ ;
	wire _w3939_ ;
	wire _w3940_ ;
	wire _w3941_ ;
	wire _w3942_ ;
	wire _w3943_ ;
	wire _w3944_ ;
	wire _w3945_ ;
	wire _w3946_ ;
	wire _w3947_ ;
	wire _w3948_ ;
	wire _w3949_ ;
	wire _w3950_ ;
	wire _w3951_ ;
	wire _w3952_ ;
	wire _w3953_ ;
	wire _w3954_ ;
	wire _w3955_ ;
	wire _w3956_ ;
	wire _w3957_ ;
	wire _w3958_ ;
	wire _w3959_ ;
	wire _w3960_ ;
	wire _w3961_ ;
	wire _w3962_ ;
	wire _w3963_ ;
	wire _w3964_ ;
	wire _w3965_ ;
	wire _w3966_ ;
	wire _w3967_ ;
	wire _w3968_ ;
	wire _w3969_ ;
	wire _w3970_ ;
	wire _w3971_ ;
	wire _w3972_ ;
	wire _w3973_ ;
	wire _w3974_ ;
	wire _w3975_ ;
	wire _w3976_ ;
	wire _w3977_ ;
	wire _w3978_ ;
	wire _w3979_ ;
	wire _w3980_ ;
	wire _w3981_ ;
	wire _w3982_ ;
	wire _w3983_ ;
	wire _w3984_ ;
	wire _w3985_ ;
	wire _w3986_ ;
	wire _w3987_ ;
	wire _w3988_ ;
	wire _w3989_ ;
	wire _w3990_ ;
	wire _w3991_ ;
	wire _w3992_ ;
	wire _w3993_ ;
	wire _w3994_ ;
	wire _w3995_ ;
	wire _w3996_ ;
	wire _w3997_ ;
	wire _w3998_ ;
	wire _w3999_ ;
	wire _w4000_ ;
	wire _w4001_ ;
	wire _w4002_ ;
	wire _w4003_ ;
	wire _w4004_ ;
	wire _w4005_ ;
	wire _w4006_ ;
	wire _w4007_ ;
	wire _w4008_ ;
	wire _w4009_ ;
	wire _w4010_ ;
	wire _w4011_ ;
	wire _w4012_ ;
	wire _w4013_ ;
	wire _w4014_ ;
	wire _w4015_ ;
	wire _w4016_ ;
	wire _w4017_ ;
	wire _w4018_ ;
	wire _w4019_ ;
	wire _w4020_ ;
	wire _w4021_ ;
	wire _w4022_ ;
	wire _w4023_ ;
	wire _w4024_ ;
	wire _w4025_ ;
	wire _w4026_ ;
	wire _w4027_ ;
	wire _w4028_ ;
	wire _w4029_ ;
	wire _w4030_ ;
	wire _w4031_ ;
	wire _w4032_ ;
	wire _w4033_ ;
	wire _w4034_ ;
	wire _w4035_ ;
	wire _w4036_ ;
	wire _w4037_ ;
	wire _w4038_ ;
	wire _w4039_ ;
	wire _w4040_ ;
	wire _w4041_ ;
	wire _w4042_ ;
	wire _w4043_ ;
	wire _w4044_ ;
	wire _w4045_ ;
	wire _w4046_ ;
	wire _w4047_ ;
	wire _w4048_ ;
	wire _w4049_ ;
	wire _w4050_ ;
	wire _w4051_ ;
	wire _w4052_ ;
	wire _w4053_ ;
	wire _w4054_ ;
	wire _w4055_ ;
	wire _w4056_ ;
	wire _w4057_ ;
	wire _w4058_ ;
	wire _w4059_ ;
	wire _w4060_ ;
	wire _w4061_ ;
	wire _w4062_ ;
	wire _w4063_ ;
	wire _w4064_ ;
	wire _w4065_ ;
	wire _w4066_ ;
	wire _w4067_ ;
	wire _w4068_ ;
	wire _w4069_ ;
	wire _w4070_ ;
	wire _w4071_ ;
	wire _w4072_ ;
	wire _w4073_ ;
	wire _w4074_ ;
	wire _w4075_ ;
	wire _w4076_ ;
	wire _w4077_ ;
	wire _w4078_ ;
	wire _w4079_ ;
	wire _w4080_ ;
	wire _w4081_ ;
	wire _w4082_ ;
	wire _w4083_ ;
	wire _w4084_ ;
	wire _w4085_ ;
	wire _w4086_ ;
	wire _w4087_ ;
	wire _w4088_ ;
	wire _w4089_ ;
	wire _w4090_ ;
	wire _w4091_ ;
	wire _w4092_ ;
	wire _w4093_ ;
	wire _w4094_ ;
	wire _w4095_ ;
	wire _w4096_ ;
	wire _w4097_ ;
	wire _w4098_ ;
	wire _w4099_ ;
	wire _w4100_ ;
	wire _w4101_ ;
	wire _w4102_ ;
	wire _w4103_ ;
	wire _w4104_ ;
	wire _w4105_ ;
	wire _w4106_ ;
	wire _w4107_ ;
	wire _w4108_ ;
	wire _w4109_ ;
	wire _w4110_ ;
	wire _w4111_ ;
	wire _w4112_ ;
	wire _w4113_ ;
	wire _w4114_ ;
	wire _w4115_ ;
	wire _w4116_ ;
	wire _w4117_ ;
	wire _w4118_ ;
	wire _w4119_ ;
	wire _w4120_ ;
	wire _w4121_ ;
	wire _w4122_ ;
	wire _w4123_ ;
	wire _w4124_ ;
	wire _w4125_ ;
	wire _w4126_ ;
	wire _w4127_ ;
	wire _w4128_ ;
	wire _w4129_ ;
	wire _w4130_ ;
	wire _w4131_ ;
	wire _w4132_ ;
	wire _w4133_ ;
	wire _w4134_ ;
	wire _w4135_ ;
	wire _w4136_ ;
	wire _w4137_ ;
	wire _w4138_ ;
	wire _w4139_ ;
	wire _w4140_ ;
	wire _w4141_ ;
	wire _w4142_ ;
	wire _w4143_ ;
	wire _w4144_ ;
	wire _w4145_ ;
	wire _w4146_ ;
	wire _w4147_ ;
	wire _w4148_ ;
	wire _w4149_ ;
	wire _w4150_ ;
	wire _w4151_ ;
	wire _w4152_ ;
	wire _w4153_ ;
	wire _w4154_ ;
	wire _w4155_ ;
	wire _w4156_ ;
	wire _w4157_ ;
	wire _w4158_ ;
	wire _w4159_ ;
	wire _w4160_ ;
	wire _w4161_ ;
	wire _w4162_ ;
	wire _w4163_ ;
	wire _w4164_ ;
	wire _w4165_ ;
	wire _w4166_ ;
	wire _w4167_ ;
	wire _w4168_ ;
	wire _w4169_ ;
	wire _w4170_ ;
	wire _w4171_ ;
	wire _w4172_ ;
	wire _w4173_ ;
	wire _w4174_ ;
	wire _w4175_ ;
	wire _w4176_ ;
	wire _w4177_ ;
	wire _w4178_ ;
	wire _w4179_ ;
	wire _w4180_ ;
	wire _w4181_ ;
	wire _w4182_ ;
	wire _w4183_ ;
	wire _w4184_ ;
	wire _w4185_ ;
	wire _w4186_ ;
	wire _w4187_ ;
	wire _w4188_ ;
	wire _w4189_ ;
	wire _w4190_ ;
	wire _w4191_ ;
	wire _w4192_ ;
	wire _w4193_ ;
	wire _w4194_ ;
	wire _w4195_ ;
	wire _w4196_ ;
	wire _w4197_ ;
	wire _w4198_ ;
	wire _w4199_ ;
	wire _w4200_ ;
	wire _w4201_ ;
	wire _w4202_ ;
	wire _w4203_ ;
	wire _w4204_ ;
	wire _w4205_ ;
	wire _w4206_ ;
	wire _w4207_ ;
	wire _w4208_ ;
	wire _w4209_ ;
	wire _w4210_ ;
	wire _w4211_ ;
	wire _w4212_ ;
	wire _w4213_ ;
	wire _w4214_ ;
	wire _w4215_ ;
	wire _w4216_ ;
	wire _w4217_ ;
	wire _w4218_ ;
	wire _w4219_ ;
	wire _w4220_ ;
	wire _w4221_ ;
	wire _w4222_ ;
	wire _w4223_ ;
	wire _w4224_ ;
	wire _w4225_ ;
	wire _w4226_ ;
	wire _w4227_ ;
	wire _w4228_ ;
	wire _w4229_ ;
	wire _w4230_ ;
	wire _w4231_ ;
	wire _w4232_ ;
	wire _w4233_ ;
	wire _w4234_ ;
	wire _w4235_ ;
	wire _w4236_ ;
	wire _w4237_ ;
	wire _w4238_ ;
	wire _w4239_ ;
	wire _w4240_ ;
	wire _w4241_ ;
	wire _w4242_ ;
	wire _w4243_ ;
	wire _w4244_ ;
	wire _w4245_ ;
	wire _w4246_ ;
	wire _w4247_ ;
	wire _w4248_ ;
	wire _w4249_ ;
	wire _w4250_ ;
	wire _w4251_ ;
	wire _w4252_ ;
	wire _w4253_ ;
	wire _w4254_ ;
	wire _w4255_ ;
	wire _w4256_ ;
	wire _w4257_ ;
	wire _w4258_ ;
	wire _w4259_ ;
	wire _w4260_ ;
	wire _w4261_ ;
	wire _w4262_ ;
	wire _w4263_ ;
	wire _w4264_ ;
	wire _w4265_ ;
	wire _w4266_ ;
	wire _w4267_ ;
	wire _w4268_ ;
	wire _w4269_ ;
	wire _w4270_ ;
	wire _w4271_ ;
	wire _w4272_ ;
	wire _w4273_ ;
	wire _w4274_ ;
	wire _w4275_ ;
	wire _w4276_ ;
	wire _w4277_ ;
	wire _w4278_ ;
	wire _w4279_ ;
	wire _w4280_ ;
	wire _w4281_ ;
	wire _w4282_ ;
	wire _w4283_ ;
	wire _w4284_ ;
	wire _w4285_ ;
	wire _w4286_ ;
	wire _w4287_ ;
	wire _w4288_ ;
	wire _w4289_ ;
	wire _w4290_ ;
	wire _w4291_ ;
	wire _w4292_ ;
	wire _w4293_ ;
	wire _w4294_ ;
	wire _w4295_ ;
	wire _w4296_ ;
	wire _w4297_ ;
	wire _w4298_ ;
	wire _w4299_ ;
	wire _w4300_ ;
	wire _w4301_ ;
	wire _w4302_ ;
	wire _w4303_ ;
	wire _w4304_ ;
	wire _w4305_ ;
	wire _w4306_ ;
	wire _w4307_ ;
	wire _w4308_ ;
	wire _w4309_ ;
	wire _w4310_ ;
	wire _w4311_ ;
	wire _w4312_ ;
	wire _w4313_ ;
	wire _w4314_ ;
	wire _w4315_ ;
	wire _w4316_ ;
	wire _w4317_ ;
	wire _w4318_ ;
	wire _w4319_ ;
	wire _w4320_ ;
	wire _w4321_ ;
	wire _w4322_ ;
	wire _w4323_ ;
	wire _w4324_ ;
	wire _w4325_ ;
	wire _w4326_ ;
	wire _w4327_ ;
	wire _w4328_ ;
	wire _w4329_ ;
	wire _w4330_ ;
	wire _w4331_ ;
	wire _w4332_ ;
	wire _w4333_ ;
	wire _w4334_ ;
	wire _w4335_ ;
	wire _w4336_ ;
	wire _w4337_ ;
	wire _w4338_ ;
	wire _w4339_ ;
	wire _w4340_ ;
	wire _w4341_ ;
	wire _w4342_ ;
	wire _w4343_ ;
	wire _w4344_ ;
	wire _w4345_ ;
	wire _w4346_ ;
	wire _w4347_ ;
	wire _w4348_ ;
	wire _w4349_ ;
	wire _w4350_ ;
	wire _w4351_ ;
	wire _w4352_ ;
	wire _w4353_ ;
	wire _w4354_ ;
	wire _w4355_ ;
	wire _w4356_ ;
	wire _w4357_ ;
	wire _w4358_ ;
	wire _w4359_ ;
	wire _w4360_ ;
	wire _w4361_ ;
	wire _w4362_ ;
	wire _w4363_ ;
	wire _w4364_ ;
	wire _w4365_ ;
	wire _w4366_ ;
	wire _w4367_ ;
	wire _w4368_ ;
	wire _w4369_ ;
	wire _w4370_ ;
	wire _w4371_ ;
	wire _w4372_ ;
	wire _w4373_ ;
	wire _w4374_ ;
	wire _w4375_ ;
	wire _w4376_ ;
	wire _w4377_ ;
	wire _w4378_ ;
	wire _w4379_ ;
	wire _w4380_ ;
	wire _w4381_ ;
	wire _w4382_ ;
	wire _w4383_ ;
	wire _w4384_ ;
	wire _w4385_ ;
	wire _w4386_ ;
	wire _w4387_ ;
	wire _w4388_ ;
	wire _w4389_ ;
	wire _w4390_ ;
	wire _w4391_ ;
	wire _w4392_ ;
	wire _w4393_ ;
	wire _w4394_ ;
	wire _w4395_ ;
	wire _w4396_ ;
	wire _w4397_ ;
	wire _w4398_ ;
	wire _w4399_ ;
	wire _w4400_ ;
	wire _w4401_ ;
	wire _w4402_ ;
	wire _w4403_ ;
	wire _w4404_ ;
	wire _w4405_ ;
	wire _w4406_ ;
	wire _w4407_ ;
	wire _w4408_ ;
	wire _w4409_ ;
	wire _w4410_ ;
	wire _w4411_ ;
	wire _w4412_ ;
	wire _w4413_ ;
	wire _w4414_ ;
	wire _w4415_ ;
	wire _w4416_ ;
	wire _w4417_ ;
	wire _w4418_ ;
	wire _w4419_ ;
	wire _w4420_ ;
	wire _w4421_ ;
	wire _w4422_ ;
	wire _w4423_ ;
	wire _w4424_ ;
	wire _w4425_ ;
	wire _w4426_ ;
	wire _w4427_ ;
	wire _w4428_ ;
	wire _w4429_ ;
	wire _w4430_ ;
	wire _w4431_ ;
	wire _w4432_ ;
	wire _w4433_ ;
	wire _w4434_ ;
	wire _w4435_ ;
	wire _w4436_ ;
	wire _w4437_ ;
	wire _w4438_ ;
	wire _w4439_ ;
	wire _w4440_ ;
	wire _w4441_ ;
	wire _w4442_ ;
	wire _w4443_ ;
	wire _w4444_ ;
	wire _w4445_ ;
	wire _w4446_ ;
	wire _w4447_ ;
	wire _w4448_ ;
	wire _w4449_ ;
	wire _w4450_ ;
	wire _w4451_ ;
	wire _w4452_ ;
	wire _w4453_ ;
	wire _w4454_ ;
	wire _w4455_ ;
	wire _w4456_ ;
	wire _w4457_ ;
	wire _w4458_ ;
	wire _w4459_ ;
	wire _w4460_ ;
	wire _w4461_ ;
	wire _w4462_ ;
	wire _w4463_ ;
	wire _w4464_ ;
	wire _w4465_ ;
	wire _w4466_ ;
	wire _w4467_ ;
	wire _w4468_ ;
	wire _w4469_ ;
	wire _w4470_ ;
	wire _w4471_ ;
	wire _w4472_ ;
	wire _w4473_ ;
	wire _w4474_ ;
	wire _w4475_ ;
	wire _w4476_ ;
	wire _w4477_ ;
	wire _w4478_ ;
	wire _w4479_ ;
	wire _w4480_ ;
	wire _w4481_ ;
	wire _w4482_ ;
	wire _w4483_ ;
	wire _w4484_ ;
	wire _w4485_ ;
	wire _w4486_ ;
	wire _w4487_ ;
	wire _w4488_ ;
	wire _w4489_ ;
	wire _w4490_ ;
	wire _w4491_ ;
	wire _w4492_ ;
	wire _w4493_ ;
	wire _w4494_ ;
	wire _w4495_ ;
	wire _w4496_ ;
	wire _w4497_ ;
	wire _w4498_ ;
	wire _w4499_ ;
	wire _w4500_ ;
	wire _w4501_ ;
	wire _w4502_ ;
	wire _w4503_ ;
	wire _w4504_ ;
	wire _w4505_ ;
	wire _w4506_ ;
	wire _w4507_ ;
	wire _w4508_ ;
	wire _w4509_ ;
	wire _w4510_ ;
	wire _w4511_ ;
	wire _w4512_ ;
	wire _w4513_ ;
	wire _w4514_ ;
	wire _w4515_ ;
	wire _w4516_ ;
	wire _w4517_ ;
	wire _w4518_ ;
	wire _w4519_ ;
	wire _w4520_ ;
	wire _w4521_ ;
	wire _w4522_ ;
	wire _w4523_ ;
	wire _w4524_ ;
	wire _w4525_ ;
	wire _w4526_ ;
	wire _w4527_ ;
	wire _w4528_ ;
	wire _w4529_ ;
	wire _w4530_ ;
	wire _w4531_ ;
	wire _w4532_ ;
	wire _w4533_ ;
	wire _w4534_ ;
	wire _w4535_ ;
	wire _w4536_ ;
	wire _w4537_ ;
	wire _w4538_ ;
	wire _w4539_ ;
	wire _w4540_ ;
	wire _w4541_ ;
	wire _w4542_ ;
	wire _w4543_ ;
	wire _w4544_ ;
	wire _w4545_ ;
	wire _w4546_ ;
	wire _w4547_ ;
	wire _w4548_ ;
	wire _w4549_ ;
	wire _w4550_ ;
	wire _w4551_ ;
	wire _w4552_ ;
	wire _w4553_ ;
	wire _w4554_ ;
	wire _w4555_ ;
	wire _w4556_ ;
	wire _w4557_ ;
	wire _w4558_ ;
	wire _w4559_ ;
	wire _w4560_ ;
	wire _w4561_ ;
	wire _w4562_ ;
	wire _w4563_ ;
	wire _w4564_ ;
	wire _w4565_ ;
	wire _w4566_ ;
	wire _w4567_ ;
	wire _w4568_ ;
	wire _w4569_ ;
	wire _w4570_ ;
	wire _w4571_ ;
	wire _w4572_ ;
	wire _w4573_ ;
	wire _w4574_ ;
	wire _w4575_ ;
	wire _w4576_ ;
	wire _w4577_ ;
	wire _w4578_ ;
	wire _w4579_ ;
	wire _w4580_ ;
	wire _w4581_ ;
	wire _w4582_ ;
	wire _w4583_ ;
	wire _w4584_ ;
	wire _w4585_ ;
	wire _w4586_ ;
	wire _w4587_ ;
	wire _w4588_ ;
	wire _w4589_ ;
	wire _w4590_ ;
	wire _w4591_ ;
	wire _w4592_ ;
	wire _w4593_ ;
	wire _w4594_ ;
	wire _w4595_ ;
	wire _w4596_ ;
	wire _w4597_ ;
	wire _w4598_ ;
	wire _w4599_ ;
	wire _w4600_ ;
	wire _w4601_ ;
	wire _w4602_ ;
	wire _w4603_ ;
	wire _w4604_ ;
	wire _w4605_ ;
	wire _w4606_ ;
	wire _w4607_ ;
	wire _w4608_ ;
	wire _w4609_ ;
	wire _w4610_ ;
	wire _w4611_ ;
	wire _w4612_ ;
	wire _w4613_ ;
	wire _w4614_ ;
	wire _w4615_ ;
	wire _w4616_ ;
	wire _w4617_ ;
	wire _w4618_ ;
	wire _w4619_ ;
	wire _w4620_ ;
	wire _w4621_ ;
	wire _w4622_ ;
	wire _w4623_ ;
	wire _w4624_ ;
	wire _w4625_ ;
	wire _w4626_ ;
	wire _w4627_ ;
	wire _w4628_ ;
	wire _w4629_ ;
	wire _w4630_ ;
	wire _w4631_ ;
	wire _w4632_ ;
	wire _w4633_ ;
	wire _w4634_ ;
	wire _w4635_ ;
	wire _w4636_ ;
	wire _w4637_ ;
	wire _w4638_ ;
	wire _w4639_ ;
	wire _w4640_ ;
	wire _w4641_ ;
	wire _w4642_ ;
	wire _w4643_ ;
	wire _w4644_ ;
	wire _w4645_ ;
	wire _w4646_ ;
	wire _w4647_ ;
	wire _w4648_ ;
	wire _w4649_ ;
	wire _w4650_ ;
	wire _w4651_ ;
	wire _w4652_ ;
	wire _w4653_ ;
	wire _w4654_ ;
	wire _w4655_ ;
	wire _w4656_ ;
	wire _w4657_ ;
	wire _w4658_ ;
	wire _w4659_ ;
	wire _w4660_ ;
	wire _w4661_ ;
	wire _w4662_ ;
	wire _w4663_ ;
	wire _w4664_ ;
	wire _w4665_ ;
	wire _w4666_ ;
	wire _w4667_ ;
	wire _w4668_ ;
	wire _w4669_ ;
	wire _w4670_ ;
	wire _w4671_ ;
	wire _w4672_ ;
	wire _w4673_ ;
	wire _w4674_ ;
	wire _w4675_ ;
	wire _w4676_ ;
	wire _w4677_ ;
	wire _w4678_ ;
	wire _w4679_ ;
	wire _w4680_ ;
	wire _w4681_ ;
	wire _w4682_ ;
	wire _w4683_ ;
	wire _w4684_ ;
	wire _w4685_ ;
	wire _w4686_ ;
	wire _w4687_ ;
	wire _w4688_ ;
	wire _w4689_ ;
	wire _w4690_ ;
	wire _w4691_ ;
	wire _w4692_ ;
	wire _w4693_ ;
	wire _w4694_ ;
	wire _w4695_ ;
	wire _w4696_ ;
	wire _w4697_ ;
	wire _w4698_ ;
	wire _w4699_ ;
	wire _w4700_ ;
	wire _w4701_ ;
	wire _w4702_ ;
	wire _w4703_ ;
	wire _w4704_ ;
	wire _w4705_ ;
	wire _w4706_ ;
	wire _w4707_ ;
	wire _w4708_ ;
	wire _w4709_ ;
	wire _w4710_ ;
	wire _w4711_ ;
	wire _w4712_ ;
	wire _w4713_ ;
	wire _w4714_ ;
	wire _w4715_ ;
	wire _w4716_ ;
	wire _w4717_ ;
	wire _w4718_ ;
	wire _w4719_ ;
	wire _w4720_ ;
	wire _w4721_ ;
	wire _w4722_ ;
	wire _w4723_ ;
	wire _w4724_ ;
	wire _w4725_ ;
	wire _w4726_ ;
	wire _w4727_ ;
	wire _w4728_ ;
	wire _w4729_ ;
	wire _w4730_ ;
	wire _w4731_ ;
	wire _w4732_ ;
	wire _w4733_ ;
	wire _w4734_ ;
	wire _w4735_ ;
	wire _w4736_ ;
	wire _w4737_ ;
	wire _w4738_ ;
	wire _w4739_ ;
	wire _w4740_ ;
	wire _w4741_ ;
	wire _w4742_ ;
	wire _w4743_ ;
	wire _w4744_ ;
	wire _w4745_ ;
	wire _w4746_ ;
	wire _w4747_ ;
	wire _w4748_ ;
	wire _w4749_ ;
	wire _w4750_ ;
	wire _w4751_ ;
	wire _w4752_ ;
	wire _w4753_ ;
	wire _w4754_ ;
	wire _w4755_ ;
	wire _w4756_ ;
	wire _w4757_ ;
	wire _w4758_ ;
	wire _w4759_ ;
	wire _w4760_ ;
	wire _w4761_ ;
	wire _w4762_ ;
	wire _w4763_ ;
	wire _w4764_ ;
	wire _w4765_ ;
	wire _w4766_ ;
	wire _w4767_ ;
	wire _w4768_ ;
	wire _w4769_ ;
	wire _w4770_ ;
	wire _w4771_ ;
	wire _w4772_ ;
	wire _w4773_ ;
	wire _w4774_ ;
	wire _w4775_ ;
	wire _w4776_ ;
	wire _w4777_ ;
	wire _w4778_ ;
	wire _w4779_ ;
	wire _w4780_ ;
	wire _w4781_ ;
	wire _w4782_ ;
	wire _w4783_ ;
	wire _w4784_ ;
	wire _w4785_ ;
	wire _w4786_ ;
	wire _w4787_ ;
	wire _w4788_ ;
	wire _w4789_ ;
	wire _w4790_ ;
	wire _w4791_ ;
	wire _w4792_ ;
	wire _w4793_ ;
	wire _w4794_ ;
	wire _w4795_ ;
	wire _w4796_ ;
	wire _w4797_ ;
	wire _w4798_ ;
	wire _w4799_ ;
	wire _w4800_ ;
	wire _w4801_ ;
	wire _w4802_ ;
	wire _w4803_ ;
	wire _w4804_ ;
	wire _w4805_ ;
	wire _w4806_ ;
	wire _w4807_ ;
	wire _w4808_ ;
	wire _w4809_ ;
	wire _w4810_ ;
	wire _w4811_ ;
	wire _w4812_ ;
	wire _w4813_ ;
	wire _w4814_ ;
	wire _w4815_ ;
	wire _w4816_ ;
	wire _w4817_ ;
	wire _w4818_ ;
	wire _w4819_ ;
	wire _w4820_ ;
	wire _w4821_ ;
	wire _w4822_ ;
	wire _w4823_ ;
	wire _w4824_ ;
	wire _w4825_ ;
	wire _w4826_ ;
	wire _w4827_ ;
	wire _w4828_ ;
	wire _w4829_ ;
	wire _w4830_ ;
	wire _w4831_ ;
	wire _w4832_ ;
	wire _w4833_ ;
	wire _w4834_ ;
	wire _w4835_ ;
	wire _w4836_ ;
	wire _w4837_ ;
	wire _w4838_ ;
	wire _w4839_ ;
	wire _w4840_ ;
	wire _w4841_ ;
	wire _w4842_ ;
	wire _w4843_ ;
	wire _w4844_ ;
	wire _w4845_ ;
	wire _w4846_ ;
	wire _w4847_ ;
	wire _w4848_ ;
	wire _w4849_ ;
	wire _w4850_ ;
	wire _w4851_ ;
	wire _w4852_ ;
	wire _w4853_ ;
	wire _w4854_ ;
	wire _w4855_ ;
	wire _w4856_ ;
	wire _w4857_ ;
	wire _w4858_ ;
	wire _w4859_ ;
	wire _w4860_ ;
	wire _w4861_ ;
	wire _w4862_ ;
	wire _w4863_ ;
	wire _w4864_ ;
	wire _w4865_ ;
	wire _w4866_ ;
	wire _w4867_ ;
	wire _w4868_ ;
	wire _w4869_ ;
	wire _w4870_ ;
	wire _w4871_ ;
	wire _w4872_ ;
	wire _w4873_ ;
	wire _w4874_ ;
	wire _w4875_ ;
	wire _w4876_ ;
	wire _w4877_ ;
	wire _w4878_ ;
	wire _w4879_ ;
	wire _w4880_ ;
	wire _w4881_ ;
	wire _w4882_ ;
	wire _w4883_ ;
	wire _w4884_ ;
	wire _w4885_ ;
	wire _w4886_ ;
	wire _w4887_ ;
	wire _w4888_ ;
	wire _w4889_ ;
	wire _w4890_ ;
	wire _w4891_ ;
	wire _w4892_ ;
	wire _w4893_ ;
	wire _w4894_ ;
	wire _w4895_ ;
	wire _w4896_ ;
	wire _w4897_ ;
	wire _w4898_ ;
	wire _w4899_ ;
	wire _w4900_ ;
	wire _w4901_ ;
	wire _w4902_ ;
	wire _w4903_ ;
	wire _w4904_ ;
	wire _w4905_ ;
	wire _w4906_ ;
	wire _w4907_ ;
	wire _w4908_ ;
	wire _w4909_ ;
	wire _w4910_ ;
	wire _w4911_ ;
	wire _w4912_ ;
	wire _w4913_ ;
	wire _w4914_ ;
	wire _w4915_ ;
	wire _w4916_ ;
	wire _w4917_ ;
	wire _w4918_ ;
	wire _w4919_ ;
	wire _w4920_ ;
	wire _w4921_ ;
	wire _w4922_ ;
	wire _w4923_ ;
	wire _w4924_ ;
	wire _w4925_ ;
	wire _w4926_ ;
	wire _w4927_ ;
	wire _w4928_ ;
	wire _w4929_ ;
	wire _w4930_ ;
	wire _w4931_ ;
	wire _w4932_ ;
	wire _w4933_ ;
	wire _w4934_ ;
	wire _w4935_ ;
	wire _w4936_ ;
	wire _w4937_ ;
	wire _w4938_ ;
	wire _w4939_ ;
	wire _w4940_ ;
	wire _w4941_ ;
	wire _w4942_ ;
	wire _w4943_ ;
	wire _w4944_ ;
	wire _w4945_ ;
	wire _w4946_ ;
	wire _w4947_ ;
	wire _w4948_ ;
	wire _w4949_ ;
	wire _w4950_ ;
	wire _w4951_ ;
	wire _w4952_ ;
	wire _w4953_ ;
	wire _w4954_ ;
	wire _w4955_ ;
	wire _w4956_ ;
	wire _w4957_ ;
	wire _w4958_ ;
	wire _w4959_ ;
	wire _w4960_ ;
	wire _w4961_ ;
	wire _w4962_ ;
	wire _w4963_ ;
	wire _w4964_ ;
	wire _w4965_ ;
	wire _w4966_ ;
	wire _w4967_ ;
	wire _w4968_ ;
	wire _w4969_ ;
	wire _w4970_ ;
	wire _w4971_ ;
	wire _w4972_ ;
	wire _w4973_ ;
	wire _w4974_ ;
	wire _w4975_ ;
	wire _w4976_ ;
	wire _w4977_ ;
	wire _w4978_ ;
	wire _w4979_ ;
	wire _w4980_ ;
	wire _w4981_ ;
	wire _w4982_ ;
	wire _w4983_ ;
	wire _w4984_ ;
	wire _w4985_ ;
	wire _w4986_ ;
	wire _w4987_ ;
	wire _w4988_ ;
	wire _w4989_ ;
	wire _w4990_ ;
	wire _w4991_ ;
	wire _w4992_ ;
	wire _w4993_ ;
	wire _w4994_ ;
	wire _w4995_ ;
	wire _w4996_ ;
	wire _w4997_ ;
	wire _w4998_ ;
	wire _w4999_ ;
	wire _w5000_ ;
	wire _w5001_ ;
	wire _w5002_ ;
	wire _w5003_ ;
	wire _w5004_ ;
	wire _w5005_ ;
	wire _w5006_ ;
	wire _w5007_ ;
	wire _w5008_ ;
	wire _w5009_ ;
	wire _w5010_ ;
	wire _w5011_ ;
	wire _w5012_ ;
	wire _w5013_ ;
	wire _w5014_ ;
	wire _w5015_ ;
	wire _w5016_ ;
	wire _w5017_ ;
	wire _w5018_ ;
	wire _w5019_ ;
	wire _w5020_ ;
	wire _w5021_ ;
	wire _w5022_ ;
	wire _w5023_ ;
	wire _w5024_ ;
	wire _w5025_ ;
	wire _w5026_ ;
	wire _w5027_ ;
	wire _w5028_ ;
	wire _w5029_ ;
	wire _w5030_ ;
	wire _w5031_ ;
	wire _w5032_ ;
	wire _w5033_ ;
	wire _w5034_ ;
	wire _w5035_ ;
	wire _w5036_ ;
	wire _w5037_ ;
	wire _w5038_ ;
	wire _w5039_ ;
	wire _w5040_ ;
	wire _w5041_ ;
	wire _w5042_ ;
	wire _w5043_ ;
	wire _w5044_ ;
	wire _w5045_ ;
	wire _w5046_ ;
	wire _w5047_ ;
	wire _w5048_ ;
	wire _w5049_ ;
	wire _w5050_ ;
	wire _w5051_ ;
	wire _w5052_ ;
	wire _w5053_ ;
	wire _w5054_ ;
	wire _w5055_ ;
	wire _w5056_ ;
	wire _w5057_ ;
	wire _w5058_ ;
	wire _w5059_ ;
	wire _w5060_ ;
	wire _w5061_ ;
	wire _w5062_ ;
	wire _w5063_ ;
	wire _w5064_ ;
	wire _w5065_ ;
	wire _w5066_ ;
	wire _w5067_ ;
	wire _w5068_ ;
	wire _w5069_ ;
	wire _w5070_ ;
	wire _w5071_ ;
	wire _w5072_ ;
	wire _w5073_ ;
	wire _w5074_ ;
	wire _w5075_ ;
	wire _w5076_ ;
	wire _w5077_ ;
	wire _w5078_ ;
	wire _w5079_ ;
	wire _w5080_ ;
	wire _w5081_ ;
	wire _w5082_ ;
	wire _w5083_ ;
	wire _w5084_ ;
	wire _w5085_ ;
	wire _w5086_ ;
	wire _w5087_ ;
	wire _w5088_ ;
	wire _w5089_ ;
	wire _w5090_ ;
	wire _w5091_ ;
	wire _w5092_ ;
	wire _w5093_ ;
	wire _w5094_ ;
	wire _w5095_ ;
	wire _w5096_ ;
	wire _w5097_ ;
	wire _w5098_ ;
	wire _w5099_ ;
	wire _w5100_ ;
	wire _w5101_ ;
	wire _w5102_ ;
	wire _w5103_ ;
	wire _w5104_ ;
	wire _w5105_ ;
	wire _w5106_ ;
	wire _w5107_ ;
	wire _w5108_ ;
	wire _w5109_ ;
	wire _w5110_ ;
	wire _w5111_ ;
	wire _w5112_ ;
	wire _w5113_ ;
	wire _w5114_ ;
	wire _w5115_ ;
	wire _w5116_ ;
	wire _w5117_ ;
	wire _w5118_ ;
	wire _w5119_ ;
	wire _w5120_ ;
	wire _w5121_ ;
	wire _w5122_ ;
	wire _w5123_ ;
	wire _w5124_ ;
	wire _w5125_ ;
	wire _w5126_ ;
	wire _w5127_ ;
	wire _w5128_ ;
	wire _w5129_ ;
	wire _w5130_ ;
	wire _w5131_ ;
	wire _w5132_ ;
	wire _w5133_ ;
	wire _w5134_ ;
	wire _w5135_ ;
	wire _w5136_ ;
	wire _w5137_ ;
	wire _w5138_ ;
	wire _w5139_ ;
	wire _w5140_ ;
	wire _w5141_ ;
	wire _w5142_ ;
	wire _w5143_ ;
	wire _w5144_ ;
	wire _w5145_ ;
	wire _w5146_ ;
	wire _w5147_ ;
	wire _w5148_ ;
	wire _w5149_ ;
	wire _w5150_ ;
	wire _w5151_ ;
	wire _w5152_ ;
	wire _w5153_ ;
	wire _w5154_ ;
	wire _w5155_ ;
	wire _w5156_ ;
	wire _w5157_ ;
	wire _w5158_ ;
	wire _w5159_ ;
	wire _w5160_ ;
	wire _w5161_ ;
	wire _w5162_ ;
	wire _w5163_ ;
	wire _w5164_ ;
	wire _w5165_ ;
	wire _w5166_ ;
	wire _w5167_ ;
	wire _w5168_ ;
	wire _w5169_ ;
	wire _w5170_ ;
	wire _w5171_ ;
	wire _w5172_ ;
	wire _w5173_ ;
	wire _w5174_ ;
	wire _w5175_ ;
	wire _w5176_ ;
	wire _w5177_ ;
	wire _w5178_ ;
	wire _w5179_ ;
	wire _w5180_ ;
	wire _w5181_ ;
	wire _w5182_ ;
	wire _w5183_ ;
	wire _w5184_ ;
	wire _w5185_ ;
	wire _w5186_ ;
	wire _w5187_ ;
	wire _w5188_ ;
	wire _w5189_ ;
	wire _w5190_ ;
	wire _w5191_ ;
	wire _w5192_ ;
	wire _w5193_ ;
	wire _w5194_ ;
	wire _w5195_ ;
	wire _w5196_ ;
	wire _w5197_ ;
	wire _w5198_ ;
	wire _w5199_ ;
	wire _w5200_ ;
	wire _w5201_ ;
	wire _w5202_ ;
	wire _w5203_ ;
	wire _w5204_ ;
	wire _w5205_ ;
	wire _w5206_ ;
	wire _w5207_ ;
	wire _w5208_ ;
	wire _w5209_ ;
	wire _w5210_ ;
	wire _w5211_ ;
	wire _w5212_ ;
	wire _w5213_ ;
	wire _w5214_ ;
	wire _w5215_ ;
	wire _w5216_ ;
	wire _w5217_ ;
	wire _w5218_ ;
	wire _w5219_ ;
	wire _w5220_ ;
	wire _w5221_ ;
	wire _w5222_ ;
	wire _w5223_ ;
	wire _w5224_ ;
	wire _w5225_ ;
	wire _w5226_ ;
	wire _w5227_ ;
	wire _w5228_ ;
	wire _w5229_ ;
	wire _w5230_ ;
	wire _w5231_ ;
	wire _w5232_ ;
	wire _w5233_ ;
	wire _w5234_ ;
	wire _w5235_ ;
	wire _w5236_ ;
	wire _w5237_ ;
	wire _w5238_ ;
	wire _w5239_ ;
	wire _w5240_ ;
	wire _w5241_ ;
	wire _w5242_ ;
	wire _w5243_ ;
	wire _w5244_ ;
	wire _w5245_ ;
	wire _w5246_ ;
	wire _w5247_ ;
	wire _w5248_ ;
	wire _w5249_ ;
	wire _w5250_ ;
	wire _w5251_ ;
	wire _w5252_ ;
	wire _w5253_ ;
	wire _w5254_ ;
	wire _w5255_ ;
	wire _w5256_ ;
	wire _w5257_ ;
	wire _w5258_ ;
	wire _w5259_ ;
	wire _w5260_ ;
	wire _w5261_ ;
	wire _w5262_ ;
	wire _w5263_ ;
	wire _w5264_ ;
	wire _w5265_ ;
	wire _w5266_ ;
	wire _w5267_ ;
	wire _w5268_ ;
	wire _w5269_ ;
	wire _w5270_ ;
	wire _w5271_ ;
	wire _w5272_ ;
	wire _w5273_ ;
	wire _w5274_ ;
	wire _w5275_ ;
	wire _w5276_ ;
	wire _w5277_ ;
	wire _w5278_ ;
	wire _w5279_ ;
	wire _w5280_ ;
	wire _w5281_ ;
	wire _w5282_ ;
	wire _w5283_ ;
	wire _w5284_ ;
	wire _w5285_ ;
	wire _w5286_ ;
	wire _w5287_ ;
	wire _w5288_ ;
	wire _w5289_ ;
	wire _w5290_ ;
	wire _w5291_ ;
	wire _w5292_ ;
	wire _w5293_ ;
	wire _w5294_ ;
	wire _w5295_ ;
	wire _w5296_ ;
	wire _w5297_ ;
	wire _w5298_ ;
	wire _w5299_ ;
	wire _w5300_ ;
	wire _w5301_ ;
	wire _w5302_ ;
	wire _w5303_ ;
	wire _w5304_ ;
	wire _w5305_ ;
	wire _w5306_ ;
	wire _w5307_ ;
	wire _w5308_ ;
	wire _w5309_ ;
	wire _w5310_ ;
	wire _w5311_ ;
	wire _w5312_ ;
	wire _w5313_ ;
	wire _w5314_ ;
	wire _w5315_ ;
	wire _w5316_ ;
	wire _w5317_ ;
	wire _w5318_ ;
	wire _w5319_ ;
	wire _w5320_ ;
	wire _w5321_ ;
	wire _w5322_ ;
	wire _w5323_ ;
	wire _w5324_ ;
	wire _w5325_ ;
	wire _w5326_ ;
	wire _w5327_ ;
	wire _w5328_ ;
	wire _w5329_ ;
	wire _w5330_ ;
	wire _w5331_ ;
	wire _w5332_ ;
	wire _w5333_ ;
	wire _w5334_ ;
	wire _w5335_ ;
	wire _w5336_ ;
	wire _w5337_ ;
	wire _w5338_ ;
	wire _w5339_ ;
	wire _w5340_ ;
	wire _w5341_ ;
	wire _w5342_ ;
	wire _w5343_ ;
	wire _w5344_ ;
	wire _w5345_ ;
	wire _w5346_ ;
	wire _w5347_ ;
	wire _w5348_ ;
	wire _w5349_ ;
	wire _w5350_ ;
	wire _w5351_ ;
	wire _w5352_ ;
	wire _w5353_ ;
	wire _w5354_ ;
	wire _w5355_ ;
	wire _w5356_ ;
	wire _w5357_ ;
	wire _w5358_ ;
	wire _w5359_ ;
	wire _w5360_ ;
	wire _w5361_ ;
	wire _w5362_ ;
	wire _w5363_ ;
	wire _w5364_ ;
	wire _w5365_ ;
	wire _w5366_ ;
	wire _w5367_ ;
	wire _w5368_ ;
	wire _w5369_ ;
	wire _w5370_ ;
	wire _w5371_ ;
	wire _w5372_ ;
	wire _w5373_ ;
	wire _w5374_ ;
	wire _w5375_ ;
	wire _w5376_ ;
	wire _w5377_ ;
	wire _w5378_ ;
	wire _w5379_ ;
	wire _w5380_ ;
	wire _w5381_ ;
	wire _w5382_ ;
	wire _w5383_ ;
	wire _w5384_ ;
	wire _w5385_ ;
	wire _w5386_ ;
	wire _w5387_ ;
	wire _w5388_ ;
	wire _w5389_ ;
	wire _w5390_ ;
	wire _w5391_ ;
	wire _w5392_ ;
	wire _w5393_ ;
	wire _w5394_ ;
	wire _w5395_ ;
	wire _w5396_ ;
	wire _w5397_ ;
	wire _w5398_ ;
	wire _w5399_ ;
	wire _w5400_ ;
	wire _w5401_ ;
	wire _w5402_ ;
	wire _w5403_ ;
	wire _w5404_ ;
	wire _w5405_ ;
	wire _w5406_ ;
	wire _w5407_ ;
	wire _w5408_ ;
	wire _w5409_ ;
	wire _w5410_ ;
	wire _w5411_ ;
	wire _w5412_ ;
	wire _w5413_ ;
	wire _w5414_ ;
	wire _w5415_ ;
	wire _w5416_ ;
	wire _w5417_ ;
	wire _w5418_ ;
	wire _w5419_ ;
	wire _w5420_ ;
	wire _w5421_ ;
	wire _w5422_ ;
	wire _w5423_ ;
	wire _w5424_ ;
	wire _w5425_ ;
	wire _w5426_ ;
	wire _w5427_ ;
	wire _w5428_ ;
	wire _w5429_ ;
	wire _w5430_ ;
	wire _w5431_ ;
	wire _w5432_ ;
	wire _w5433_ ;
	wire _w5434_ ;
	wire _w5435_ ;
	wire _w5436_ ;
	wire _w5437_ ;
	wire _w5438_ ;
	wire _w5439_ ;
	wire _w5440_ ;
	wire _w5441_ ;
	wire _w5442_ ;
	wire _w5443_ ;
	wire _w5444_ ;
	wire _w5445_ ;
	wire _w5446_ ;
	wire _w5447_ ;
	wire _w5448_ ;
	wire _w5449_ ;
	wire _w5450_ ;
	wire _w5451_ ;
	wire _w5452_ ;
	wire _w5453_ ;
	wire _w5454_ ;
	wire _w5455_ ;
	wire _w5456_ ;
	wire _w5457_ ;
	wire _w5458_ ;
	wire _w5459_ ;
	wire _w5460_ ;
	wire _w5461_ ;
	wire _w5462_ ;
	wire _w5463_ ;
	wire _w5464_ ;
	wire _w5465_ ;
	wire _w5466_ ;
	wire _w5467_ ;
	wire _w5468_ ;
	wire _w5469_ ;
	wire _w5470_ ;
	wire _w5471_ ;
	wire _w5472_ ;
	wire _w5473_ ;
	wire _w5474_ ;
	wire _w5475_ ;
	wire _w5476_ ;
	wire _w5477_ ;
	wire _w5478_ ;
	wire _w5479_ ;
	wire _w5480_ ;
	wire _w5481_ ;
	wire _w5482_ ;
	wire _w5483_ ;
	wire _w5484_ ;
	wire _w5485_ ;
	wire _w5486_ ;
	wire _w5487_ ;
	wire _w5488_ ;
	wire _w5489_ ;
	wire _w5490_ ;
	wire _w5491_ ;
	wire _w5492_ ;
	wire _w5493_ ;
	wire _w5494_ ;
	wire _w5495_ ;
	wire _w5496_ ;
	wire _w5497_ ;
	wire _w5498_ ;
	wire _w5499_ ;
	wire _w5500_ ;
	wire _w5501_ ;
	wire _w5502_ ;
	wire _w5503_ ;
	wire _w5504_ ;
	wire _w5505_ ;
	wire _w5506_ ;
	wire _w5507_ ;
	wire _w5508_ ;
	wire _w5509_ ;
	wire _w5510_ ;
	wire _w5511_ ;
	wire _w5512_ ;
	wire _w5513_ ;
	wire _w5514_ ;
	wire _w5515_ ;
	wire _w5516_ ;
	wire _w5517_ ;
	wire _w5518_ ;
	wire _w5519_ ;
	wire _w5520_ ;
	wire _w5521_ ;
	wire _w5522_ ;
	wire _w5523_ ;
	wire _w5524_ ;
	wire _w5525_ ;
	wire _w5526_ ;
	wire _w5527_ ;
	wire _w5528_ ;
	wire _w5529_ ;
	wire _w5530_ ;
	wire _w5531_ ;
	wire _w5532_ ;
	wire _w5533_ ;
	wire _w5534_ ;
	wire _w5535_ ;
	wire _w5536_ ;
	wire _w5537_ ;
	wire _w5538_ ;
	wire _w5539_ ;
	wire _w5540_ ;
	wire _w5541_ ;
	wire _w5542_ ;
	wire _w5543_ ;
	wire _w5544_ ;
	wire _w5545_ ;
	wire _w5546_ ;
	wire _w5547_ ;
	wire _w5548_ ;
	wire _w5549_ ;
	wire _w5550_ ;
	wire _w5551_ ;
	wire _w5552_ ;
	wire _w5553_ ;
	wire _w5554_ ;
	wire _w5555_ ;
	wire _w5556_ ;
	wire _w5557_ ;
	wire _w5558_ ;
	wire _w5559_ ;
	wire _w5560_ ;
	wire _w5561_ ;
	wire _w5562_ ;
	wire _w5563_ ;
	wire _w5564_ ;
	wire _w5565_ ;
	wire _w5566_ ;
	wire _w5567_ ;
	wire _w5568_ ;
	wire _w5569_ ;
	wire _w5570_ ;
	wire _w5571_ ;
	wire _w5572_ ;
	wire _w5573_ ;
	wire _w5574_ ;
	wire _w5575_ ;
	wire _w5576_ ;
	wire _w5577_ ;
	wire _w5578_ ;
	wire _w5579_ ;
	wire _w5580_ ;
	wire _w5581_ ;
	wire _w5582_ ;
	wire _w5583_ ;
	wire _w5584_ ;
	wire _w5585_ ;
	wire _w5586_ ;
	wire _w5587_ ;
	wire _w5588_ ;
	wire _w5589_ ;
	wire _w5590_ ;
	wire _w5591_ ;
	wire _w5592_ ;
	wire _w5593_ ;
	wire _w5594_ ;
	wire _w5595_ ;
	wire _w5596_ ;
	wire _w5597_ ;
	wire _w5598_ ;
	wire _w5599_ ;
	wire _w5600_ ;
	wire _w5601_ ;
	wire _w5602_ ;
	wire _w5603_ ;
	wire _w5604_ ;
	wire _w5605_ ;
	wire _w5606_ ;
	wire _w5607_ ;
	wire _w5608_ ;
	wire _w5609_ ;
	wire _w5610_ ;
	wire _w5611_ ;
	wire _w5612_ ;
	wire _w5613_ ;
	wire _w5614_ ;
	wire _w5615_ ;
	wire _w5616_ ;
	wire _w5617_ ;
	wire _w5618_ ;
	wire _w5619_ ;
	wire _w5620_ ;
	wire _w5621_ ;
	wire _w5622_ ;
	wire _w5623_ ;
	wire _w5624_ ;
	wire _w5625_ ;
	wire _w5626_ ;
	wire _w5627_ ;
	wire _w5628_ ;
	wire _w5629_ ;
	wire _w5630_ ;
	wire _w5631_ ;
	wire _w5632_ ;
	wire _w5633_ ;
	wire _w5634_ ;
	wire _w5635_ ;
	wire _w5636_ ;
	wire _w5637_ ;
	wire _w5638_ ;
	wire _w5639_ ;
	wire _w5640_ ;
	wire _w5641_ ;
	wire _w5642_ ;
	wire _w5643_ ;
	wire _w5644_ ;
	wire _w5645_ ;
	wire _w5646_ ;
	wire _w5647_ ;
	wire _w5648_ ;
	wire _w5649_ ;
	wire _w5650_ ;
	wire _w5651_ ;
	wire _w5652_ ;
	wire _w5653_ ;
	wire _w5654_ ;
	wire _w5655_ ;
	wire _w5656_ ;
	wire _w5657_ ;
	wire _w5658_ ;
	wire _w5659_ ;
	wire _w5660_ ;
	wire _w5661_ ;
	wire _w5662_ ;
	wire _w5663_ ;
	wire _w5664_ ;
	wire _w5665_ ;
	wire _w5666_ ;
	wire _w5667_ ;
	wire _w5668_ ;
	wire _w5669_ ;
	wire _w5670_ ;
	wire _w5671_ ;
	wire _w5672_ ;
	wire _w5673_ ;
	wire _w5674_ ;
	wire _w5675_ ;
	wire _w5676_ ;
	wire _w5677_ ;
	wire _w5678_ ;
	wire _w5679_ ;
	wire _w5680_ ;
	wire _w5681_ ;
	wire _w5682_ ;
	wire _w5683_ ;
	wire _w5684_ ;
	wire _w5685_ ;
	wire _w5686_ ;
	wire _w5687_ ;
	wire _w5688_ ;
	wire _w5689_ ;
	wire _w5690_ ;
	wire _w5691_ ;
	wire _w5692_ ;
	wire _w5693_ ;
	wire _w5694_ ;
	wire _w5695_ ;
	wire _w5696_ ;
	wire _w5697_ ;
	wire _w5698_ ;
	wire _w5699_ ;
	wire _w5700_ ;
	wire _w5701_ ;
	wire _w5702_ ;
	wire _w5703_ ;
	wire _w5704_ ;
	wire _w5705_ ;
	wire _w5706_ ;
	wire _w5707_ ;
	wire _w5708_ ;
	wire _w5709_ ;
	wire _w5710_ ;
	wire _w5711_ ;
	wire _w5712_ ;
	wire _w5713_ ;
	wire _w5714_ ;
	wire _w5715_ ;
	wire _w5716_ ;
	wire _w5717_ ;
	wire _w5718_ ;
	wire _w5719_ ;
	wire _w5720_ ;
	wire _w5721_ ;
	wire _w5722_ ;
	wire _w5723_ ;
	wire _w5724_ ;
	wire _w5725_ ;
	wire _w5726_ ;
	wire _w5727_ ;
	wire _w5728_ ;
	wire _w5729_ ;
	wire _w5730_ ;
	wire _w5731_ ;
	wire _w5732_ ;
	wire _w5733_ ;
	wire _w5734_ ;
	wire _w5735_ ;
	wire _w5736_ ;
	wire _w5737_ ;
	wire _w5738_ ;
	wire _w5739_ ;
	wire _w5740_ ;
	wire _w5741_ ;
	wire _w5742_ ;
	wire _w5743_ ;
	wire _w5744_ ;
	wire _w5745_ ;
	wire _w5746_ ;
	wire _w5747_ ;
	wire _w5748_ ;
	wire _w5749_ ;
	wire _w5750_ ;
	wire _w5751_ ;
	wire _w5752_ ;
	wire _w5753_ ;
	wire _w5754_ ;
	wire _w5755_ ;
	wire _w5756_ ;
	wire _w5757_ ;
	wire _w5758_ ;
	wire _w5759_ ;
	wire _w5760_ ;
	wire _w5761_ ;
	wire _w5762_ ;
	wire _w5763_ ;
	wire _w5764_ ;
	wire _w5765_ ;
	wire _w5766_ ;
	wire _w5767_ ;
	wire _w5768_ ;
	wire _w5769_ ;
	wire _w5770_ ;
	wire _w5771_ ;
	wire _w5772_ ;
	wire _w5773_ ;
	wire _w5774_ ;
	wire _w5775_ ;
	wire _w5776_ ;
	wire _w5777_ ;
	wire _w5778_ ;
	wire _w5779_ ;
	wire _w5780_ ;
	wire _w5781_ ;
	wire _w5782_ ;
	wire _w5783_ ;
	wire _w5784_ ;
	wire _w5785_ ;
	wire _w5786_ ;
	wire _w5787_ ;
	wire _w5788_ ;
	wire _w5789_ ;
	wire _w5790_ ;
	wire _w5791_ ;
	wire _w5792_ ;
	wire _w5793_ ;
	wire _w5794_ ;
	wire _w5795_ ;
	wire _w5796_ ;
	wire _w5797_ ;
	wire _w5798_ ;
	wire _w5799_ ;
	wire _w5800_ ;
	wire _w5801_ ;
	wire _w5802_ ;
	wire _w5803_ ;
	wire _w5804_ ;
	wire _w5805_ ;
	wire _w5806_ ;
	wire _w5807_ ;
	wire _w5808_ ;
	wire _w5809_ ;
	wire _w5810_ ;
	wire _w5811_ ;
	wire _w5812_ ;
	wire _w5813_ ;
	wire _w5814_ ;
	wire _w5815_ ;
	wire _w5816_ ;
	wire _w5817_ ;
	wire _w5818_ ;
	wire _w5819_ ;
	wire _w5820_ ;
	wire _w5821_ ;
	wire _w5822_ ;
	wire _w5823_ ;
	wire _w5824_ ;
	wire _w5825_ ;
	wire _w5826_ ;
	wire _w5827_ ;
	wire _w5828_ ;
	wire _w5829_ ;
	wire _w5830_ ;
	wire _w5831_ ;
	wire _w5832_ ;
	wire _w5833_ ;
	wire _w5834_ ;
	wire _w5835_ ;
	wire _w5836_ ;
	wire _w5837_ ;
	wire _w5838_ ;
	wire _w5839_ ;
	wire _w5840_ ;
	wire _w5841_ ;
	wire _w5842_ ;
	wire _w5843_ ;
	wire _w5844_ ;
	wire _w5845_ ;
	wire _w5846_ ;
	wire _w5847_ ;
	wire _w5848_ ;
	wire _w5849_ ;
	wire _w5850_ ;
	wire _w5851_ ;
	wire _w5852_ ;
	wire _w5853_ ;
	wire _w5854_ ;
	wire _w5855_ ;
	wire _w5856_ ;
	wire _w5857_ ;
	wire _w5858_ ;
	wire _w5859_ ;
	wire _w5860_ ;
	wire _w5861_ ;
	wire _w5862_ ;
	wire _w5863_ ;
	wire _w5864_ ;
	wire _w5865_ ;
	wire _w5866_ ;
	wire _w5867_ ;
	wire _w5868_ ;
	wire _w5869_ ;
	wire _w5870_ ;
	wire _w5871_ ;
	wire _w5872_ ;
	wire _w5873_ ;
	wire _w5874_ ;
	wire _w5875_ ;
	wire _w5876_ ;
	wire _w5877_ ;
	wire _w5878_ ;
	wire _w5879_ ;
	wire _w5880_ ;
	wire _w5881_ ;
	wire _w5882_ ;
	wire _w5883_ ;
	wire _w5884_ ;
	wire _w5885_ ;
	wire _w5886_ ;
	wire _w5887_ ;
	wire _w5888_ ;
	wire _w5889_ ;
	wire _w5890_ ;
	wire _w5891_ ;
	wire _w5892_ ;
	wire _w5893_ ;
	wire _w5894_ ;
	wire _w5895_ ;
	wire _w5896_ ;
	wire _w5897_ ;
	wire _w5898_ ;
	wire _w5899_ ;
	wire _w5900_ ;
	wire _w5901_ ;
	wire _w5902_ ;
	wire _w5903_ ;
	wire _w5904_ ;
	wire _w5905_ ;
	wire _w5906_ ;
	wire _w5907_ ;
	wire _w5908_ ;
	wire _w5909_ ;
	wire _w5910_ ;
	wire _w5911_ ;
	wire _w5912_ ;
	wire _w5913_ ;
	wire _w5914_ ;
	wire _w5915_ ;
	wire _w5916_ ;
	wire _w5917_ ;
	wire _w5918_ ;
	wire _w5919_ ;
	wire _w5920_ ;
	wire _w5921_ ;
	wire _w5922_ ;
	wire _w5923_ ;
	wire _w5924_ ;
	wire _w5925_ ;
	wire _w5926_ ;
	wire _w5927_ ;
	wire _w5928_ ;
	wire _w5929_ ;
	wire _w5930_ ;
	wire _w5931_ ;
	wire _w5932_ ;
	wire _w5933_ ;
	wire _w5934_ ;
	wire _w5935_ ;
	wire _w5936_ ;
	wire _w5937_ ;
	wire _w5938_ ;
	wire _w5939_ ;
	wire _w5940_ ;
	wire _w5941_ ;
	wire _w5942_ ;
	wire _w5943_ ;
	wire _w5944_ ;
	wire _w5945_ ;
	wire _w5946_ ;
	wire _w5947_ ;
	wire _w5948_ ;
	wire _w5949_ ;
	wire _w5950_ ;
	wire _w5951_ ;
	wire _w5952_ ;
	wire _w5953_ ;
	wire _w5954_ ;
	wire _w5955_ ;
	wire _w5956_ ;
	wire _w5957_ ;
	wire _w5958_ ;
	wire _w5959_ ;
	wire _w5960_ ;
	wire _w5961_ ;
	wire _w5962_ ;
	wire _w5963_ ;
	wire _w5964_ ;
	wire _w5965_ ;
	wire _w5966_ ;
	wire _w5967_ ;
	wire _w5968_ ;
	wire _w5969_ ;
	wire _w5970_ ;
	wire _w5971_ ;
	wire _w5972_ ;
	wire _w5973_ ;
	wire _w5974_ ;
	wire _w5975_ ;
	wire _w5976_ ;
	wire _w5977_ ;
	wire _w5978_ ;
	wire _w5979_ ;
	wire _w5980_ ;
	wire _w5981_ ;
	wire _w5982_ ;
	wire _w5983_ ;
	wire _w5984_ ;
	wire _w5985_ ;
	wire _w5986_ ;
	wire _w5987_ ;
	wire _w5988_ ;
	wire _w5989_ ;
	wire _w5990_ ;
	wire _w5991_ ;
	wire _w5992_ ;
	wire _w5993_ ;
	wire _w5994_ ;
	wire _w5995_ ;
	wire _w5996_ ;
	wire _w5997_ ;
	wire _w5998_ ;
	wire _w5999_ ;
	wire _w6000_ ;
	wire _w6001_ ;
	wire _w6002_ ;
	wire _w6003_ ;
	wire _w6004_ ;
	wire _w6005_ ;
	wire _w6006_ ;
	wire _w6007_ ;
	wire _w6008_ ;
	wire _w6009_ ;
	wire _w6010_ ;
	wire _w6011_ ;
	wire _w6012_ ;
	wire _w6013_ ;
	wire _w6014_ ;
	wire _w6015_ ;
	wire _w6016_ ;
	wire _w6017_ ;
	wire _w6018_ ;
	wire _w6019_ ;
	wire _w6020_ ;
	wire _w6021_ ;
	wire _w6022_ ;
	wire _w6023_ ;
	wire _w6024_ ;
	wire _w6025_ ;
	wire _w6026_ ;
	wire _w6027_ ;
	wire _w6028_ ;
	wire _w6029_ ;
	wire _w6030_ ;
	wire _w6031_ ;
	wire _w6032_ ;
	wire _w6033_ ;
	wire _w6034_ ;
	wire _w6035_ ;
	wire _w6036_ ;
	wire _w6037_ ;
	wire _w6038_ ;
	wire _w6039_ ;
	wire _w6040_ ;
	wire _w6041_ ;
	wire _w6042_ ;
	wire _w6043_ ;
	wire _w6044_ ;
	wire _w6045_ ;
	wire _w6046_ ;
	wire _w6047_ ;
	wire _w6048_ ;
	wire _w6049_ ;
	wire _w6050_ ;
	wire _w6051_ ;
	wire _w6052_ ;
	wire _w6053_ ;
	wire _w6054_ ;
	wire _w6055_ ;
	wire _w6056_ ;
	wire _w6057_ ;
	wire _w6058_ ;
	wire _w6059_ ;
	wire _w6060_ ;
	wire _w6061_ ;
	wire _w6062_ ;
	wire _w6063_ ;
	wire _w6064_ ;
	wire _w6065_ ;
	wire _w6066_ ;
	wire _w6067_ ;
	wire _w6068_ ;
	wire _w6069_ ;
	wire _w6070_ ;
	wire _w6071_ ;
	wire _w6072_ ;
	wire _w6073_ ;
	wire _w6074_ ;
	wire _w6075_ ;
	wire _w6076_ ;
	wire _w6077_ ;
	wire _w6078_ ;
	wire _w6079_ ;
	wire _w6080_ ;
	wire _w6081_ ;
	wire _w6082_ ;
	wire _w6083_ ;
	wire _w6084_ ;
	wire _w6085_ ;
	wire _w6086_ ;
	wire _w6087_ ;
	wire _w6088_ ;
	wire _w6089_ ;
	wire _w6090_ ;
	wire _w6091_ ;
	wire _w6092_ ;
	wire _w6093_ ;
	wire _w6094_ ;
	wire _w6095_ ;
	wire _w6096_ ;
	wire _w6097_ ;
	wire _w6098_ ;
	wire _w6099_ ;
	wire _w6100_ ;
	wire _w6101_ ;
	wire _w6102_ ;
	wire _w6103_ ;
	wire _w6104_ ;
	wire _w6105_ ;
	wire _w6106_ ;
	wire _w6107_ ;
	wire _w6108_ ;
	wire _w6109_ ;
	wire _w6110_ ;
	wire _w6111_ ;
	wire _w6112_ ;
	wire _w6113_ ;
	wire _w6114_ ;
	wire _w6115_ ;
	wire _w6116_ ;
	wire _w6117_ ;
	wire _w6118_ ;
	wire _w6119_ ;
	wire _w6120_ ;
	wire _w6121_ ;
	wire _w6122_ ;
	wire _w6123_ ;
	wire _w6124_ ;
	wire _w6125_ ;
	wire _w6126_ ;
	wire _w6127_ ;
	wire _w6128_ ;
	wire _w6129_ ;
	wire _w6130_ ;
	wire _w6131_ ;
	wire _w6132_ ;
	wire _w6133_ ;
	wire _w6134_ ;
	wire _w6135_ ;
	wire _w6136_ ;
	wire _w6137_ ;
	wire _w6138_ ;
	wire _w6139_ ;
	wire _w6140_ ;
	wire _w6141_ ;
	wire _w6142_ ;
	wire _w6143_ ;
	wire _w6144_ ;
	wire _w6145_ ;
	wire _w6146_ ;
	wire _w6147_ ;
	wire _w6148_ ;
	wire _w6149_ ;
	wire _w6150_ ;
	wire _w6151_ ;
	wire _w6152_ ;
	wire _w6153_ ;
	wire _w6154_ ;
	wire _w6155_ ;
	wire _w6156_ ;
	wire _w6157_ ;
	wire _w6158_ ;
	wire _w6159_ ;
	wire _w6160_ ;
	wire _w6161_ ;
	wire _w6162_ ;
	wire _w6163_ ;
	wire _w6164_ ;
	wire _w6165_ ;
	wire _w6166_ ;
	wire _w6167_ ;
	wire _w6168_ ;
	wire _w6169_ ;
	wire _w6170_ ;
	wire _w6171_ ;
	wire _w6172_ ;
	wire _w6173_ ;
	wire _w6174_ ;
	wire _w6175_ ;
	wire _w6176_ ;
	wire _w6177_ ;
	wire _w6178_ ;
	wire _w6179_ ;
	wire _w6180_ ;
	wire _w6181_ ;
	wire _w6182_ ;
	wire _w6183_ ;
	wire _w6184_ ;
	wire _w6185_ ;
	wire _w6186_ ;
	wire _w6187_ ;
	wire _w6188_ ;
	wire _w6189_ ;
	wire _w6190_ ;
	wire _w6191_ ;
	wire _w6192_ ;
	wire _w6193_ ;
	wire _w6194_ ;
	wire _w6195_ ;
	wire _w6196_ ;
	wire _w6197_ ;
	wire _w6198_ ;
	wire _w6199_ ;
	wire _w6200_ ;
	wire _w6201_ ;
	wire _w6202_ ;
	wire _w6203_ ;
	wire _w6204_ ;
	wire _w6205_ ;
	wire _w6206_ ;
	wire _w6207_ ;
	wire _w6208_ ;
	wire _w6209_ ;
	wire _w6210_ ;
	wire _w6211_ ;
	wire _w6212_ ;
	wire _w6213_ ;
	wire _w6214_ ;
	wire _w6215_ ;
	wire _w6216_ ;
	wire _w6217_ ;
	wire _w6218_ ;
	wire _w6219_ ;
	wire _w6220_ ;
	wire _w6221_ ;
	wire _w6222_ ;
	wire _w6223_ ;
	wire _w6224_ ;
	wire _w6225_ ;
	wire _w6226_ ;
	wire _w6227_ ;
	wire _w6228_ ;
	wire _w6229_ ;
	wire _w6230_ ;
	wire _w6231_ ;
	wire _w6232_ ;
	wire _w6233_ ;
	wire _w6234_ ;
	wire _w6235_ ;
	wire _w6236_ ;
	wire _w6237_ ;
	wire _w6238_ ;
	wire _w6239_ ;
	wire _w6240_ ;
	wire _w6241_ ;
	wire _w6242_ ;
	wire _w6243_ ;
	wire _w6244_ ;
	wire _w6245_ ;
	wire _w6246_ ;
	wire _w6247_ ;
	wire _w6248_ ;
	wire _w6249_ ;
	wire _w6250_ ;
	wire _w6251_ ;
	wire _w6252_ ;
	wire _w6253_ ;
	wire _w6254_ ;
	wire _w6255_ ;
	wire _w6256_ ;
	wire _w6257_ ;
	wire _w6258_ ;
	wire _w6259_ ;
	wire _w6260_ ;
	wire _w6261_ ;
	wire _w6262_ ;
	wire _w6263_ ;
	wire _w6264_ ;
	wire _w6265_ ;
	wire _w6266_ ;
	wire _w6267_ ;
	wire _w6268_ ;
	wire _w6269_ ;
	wire _w6270_ ;
	wire _w6271_ ;
	wire _w6272_ ;
	wire _w6273_ ;
	wire _w6274_ ;
	wire _w6275_ ;
	wire _w6276_ ;
	wire _w6277_ ;
	wire _w6278_ ;
	wire _w6279_ ;
	wire _w6280_ ;
	wire _w6281_ ;
	wire _w6282_ ;
	wire _w6283_ ;
	wire _w6284_ ;
	wire _w6285_ ;
	wire _w6286_ ;
	wire _w6287_ ;
	wire _w6288_ ;
	wire _w6289_ ;
	wire _w6290_ ;
	wire _w6291_ ;
	wire _w6292_ ;
	wire _w6293_ ;
	wire _w6294_ ;
	wire _w6295_ ;
	wire _w6296_ ;
	wire _w6297_ ;
	wire _w6298_ ;
	wire _w6299_ ;
	wire _w6300_ ;
	wire _w6301_ ;
	wire _w6302_ ;
	wire _w6303_ ;
	wire _w6304_ ;
	wire _w6305_ ;
	wire _w6306_ ;
	wire _w6307_ ;
	wire _w6308_ ;
	wire _w6309_ ;
	wire _w6310_ ;
	wire _w6311_ ;
	wire _w6312_ ;
	wire _w6313_ ;
	wire _w6314_ ;
	wire _w6315_ ;
	wire _w6316_ ;
	wire _w6317_ ;
	wire _w6318_ ;
	wire _w6319_ ;
	wire _w6320_ ;
	wire _w6321_ ;
	wire _w6322_ ;
	wire _w6323_ ;
	wire _w6324_ ;
	wire _w6325_ ;
	wire _w6326_ ;
	wire _w6327_ ;
	wire _w6328_ ;
	wire _w6329_ ;
	wire _w6330_ ;
	wire _w6331_ ;
	wire _w6332_ ;
	wire _w6333_ ;
	wire _w6334_ ;
	wire _w6335_ ;
	wire _w6336_ ;
	wire _w6337_ ;
	wire _w6338_ ;
	wire _w6339_ ;
	wire _w6340_ ;
	wire _w6341_ ;
	wire _w6342_ ;
	wire _w6343_ ;
	wire _w6344_ ;
	wire _w6345_ ;
	wire _w6346_ ;
	wire _w6347_ ;
	wire _w6348_ ;
	wire _w6349_ ;
	wire _w6350_ ;
	wire _w6351_ ;
	wire _w6352_ ;
	wire _w6353_ ;
	wire _w6354_ ;
	wire _w6355_ ;
	wire _w6356_ ;
	wire _w6357_ ;
	wire _w6358_ ;
	wire _w6359_ ;
	wire _w6360_ ;
	wire _w6361_ ;
	wire _w6362_ ;
	wire _w6363_ ;
	wire _w6364_ ;
	wire _w6365_ ;
	wire _w6366_ ;
	wire _w6367_ ;
	wire _w6368_ ;
	wire _w6369_ ;
	wire _w6370_ ;
	wire _w6371_ ;
	wire _w6372_ ;
	wire _w6373_ ;
	wire _w6374_ ;
	wire _w6375_ ;
	wire _w6376_ ;
	wire _w6377_ ;
	wire _w6378_ ;
	wire _w6379_ ;
	wire _w6380_ ;
	wire _w6381_ ;
	wire _w6382_ ;
	wire _w6383_ ;
	wire _w6384_ ;
	wire _w6385_ ;
	wire _w6386_ ;
	wire _w6387_ ;
	wire _w6388_ ;
	wire _w6389_ ;
	wire _w6390_ ;
	wire _w6391_ ;
	wire _w6392_ ;
	wire _w6393_ ;
	wire _w6394_ ;
	wire _w6395_ ;
	wire _w6396_ ;
	wire _w6397_ ;
	wire _w6398_ ;
	wire _w6399_ ;
	wire _w6400_ ;
	wire _w6401_ ;
	wire _w6402_ ;
	wire _w6403_ ;
	wire _w6404_ ;
	wire _w6405_ ;
	wire _w6406_ ;
	wire _w6407_ ;
	wire _w6408_ ;
	wire _w6409_ ;
	wire _w6410_ ;
	wire _w6411_ ;
	wire _w6412_ ;
	wire _w6413_ ;
	wire _w6414_ ;
	wire _w6415_ ;
	wire _w6416_ ;
	wire _w6417_ ;
	wire _w6418_ ;
	wire _w6419_ ;
	wire _w6420_ ;
	wire _w6421_ ;
	wire _w6422_ ;
	wire _w6423_ ;
	wire _w6424_ ;
	wire _w6425_ ;
	wire _w6426_ ;
	wire _w6427_ ;
	wire _w6428_ ;
	wire _w6429_ ;
	wire _w6430_ ;
	wire _w6431_ ;
	wire _w6432_ ;
	wire _w6433_ ;
	wire _w6434_ ;
	wire _w6435_ ;
	wire _w6436_ ;
	wire _w6437_ ;
	wire _w6438_ ;
	wire _w6439_ ;
	wire _w6440_ ;
	wire _w6441_ ;
	wire _w6442_ ;
	wire _w6443_ ;
	wire _w6444_ ;
	wire _w6445_ ;
	wire _w6446_ ;
	wire _w6447_ ;
	wire _w6448_ ;
	wire _w6449_ ;
	wire _w6450_ ;
	wire _w6451_ ;
	wire _w6452_ ;
	wire _w6453_ ;
	wire _w6454_ ;
	wire _w6455_ ;
	wire _w6456_ ;
	wire _w6457_ ;
	wire _w6458_ ;
	wire _w6459_ ;
	wire _w6460_ ;
	wire _w6461_ ;
	wire _w6462_ ;
	wire _w6463_ ;
	wire _w6464_ ;
	wire _w6465_ ;
	wire _w6466_ ;
	wire _w6467_ ;
	wire _w6468_ ;
	wire _w6469_ ;
	wire _w6470_ ;
	wire _w6471_ ;
	wire _w6472_ ;
	wire _w6473_ ;
	wire _w6474_ ;
	wire _w6475_ ;
	wire _w6476_ ;
	wire _w6477_ ;
	wire _w6478_ ;
	wire _w6479_ ;
	wire _w6480_ ;
	wire _w6481_ ;
	wire _w6482_ ;
	wire _w6483_ ;
	wire _w6484_ ;
	wire _w6485_ ;
	wire _w6486_ ;
	wire _w6487_ ;
	wire _w6488_ ;
	wire _w6489_ ;
	wire _w6490_ ;
	wire _w6491_ ;
	wire _w6492_ ;
	wire _w6493_ ;
	wire _w6494_ ;
	wire _w6495_ ;
	wire _w6496_ ;
	wire _w6497_ ;
	wire _w6498_ ;
	wire _w6499_ ;
	wire _w6500_ ;
	wire _w6501_ ;
	wire _w6502_ ;
	wire _w6503_ ;
	wire _w6504_ ;
	wire _w6505_ ;
	wire _w6506_ ;
	wire _w6507_ ;
	wire _w6508_ ;
	wire _w6509_ ;
	wire _w6510_ ;
	wire _w6511_ ;
	wire _w6512_ ;
	wire _w6513_ ;
	wire _w6514_ ;
	wire _w6515_ ;
	wire _w6516_ ;
	wire _w6517_ ;
	wire _w6518_ ;
	wire _w6519_ ;
	wire _w6520_ ;
	wire _w6521_ ;
	wire _w6522_ ;
	wire _w6523_ ;
	wire _w6524_ ;
	wire _w6525_ ;
	wire _w6526_ ;
	wire _w6527_ ;
	wire _w6528_ ;
	wire _w6529_ ;
	wire _w6530_ ;
	wire _w6531_ ;
	wire _w6532_ ;
	wire _w6533_ ;
	wire _w6534_ ;
	wire _w6535_ ;
	wire _w6536_ ;
	wire _w6537_ ;
	wire _w6538_ ;
	wire _w6539_ ;
	wire _w6540_ ;
	wire _w6541_ ;
	wire _w6542_ ;
	wire _w6543_ ;
	wire _w6544_ ;
	wire _w6545_ ;
	wire _w6546_ ;
	wire _w6547_ ;
	wire _w6548_ ;
	wire _w6549_ ;
	wire _w6550_ ;
	wire _w6551_ ;
	wire _w6552_ ;
	wire _w6553_ ;
	wire _w6554_ ;
	wire _w6555_ ;
	wire _w6556_ ;
	wire _w6557_ ;
	wire _w6558_ ;
	wire _w6559_ ;
	wire _w6560_ ;
	wire _w6561_ ;
	wire _w6562_ ;
	wire _w6563_ ;
	wire _w6564_ ;
	wire _w6565_ ;
	wire _w6566_ ;
	wire _w6567_ ;
	wire _w6568_ ;
	wire _w6569_ ;
	wire _w6570_ ;
	wire _w6571_ ;
	wire _w6572_ ;
	wire _w6573_ ;
	wire _w6574_ ;
	wire _w6575_ ;
	wire _w6576_ ;
	wire _w6577_ ;
	wire _w6578_ ;
	wire _w6579_ ;
	wire _w6580_ ;
	wire _w6581_ ;
	wire _w6582_ ;
	wire _w6583_ ;
	wire _w6584_ ;
	wire _w6585_ ;
	wire _w6586_ ;
	wire _w6587_ ;
	wire _w6588_ ;
	wire _w6589_ ;
	wire _w6590_ ;
	wire _w6591_ ;
	wire _w6592_ ;
	wire _w6593_ ;
	wire _w6594_ ;
	LUT2 #(
		.INIT('h2)
	) name0 (
		\TM0_pad ,
		\WX10891_reg/NET0131 ,
		_w1508_
	);
	LUT2 #(
		.INIT('h2)
	) name1 (
		\WX835_reg/NET0131 ,
		\WX899_reg/NET0131 ,
		_w1509_
	);
	LUT2 #(
		.INIT('h4)
	) name2 (
		\WX835_reg/NET0131 ,
		\WX899_reg/NET0131 ,
		_w1510_
	);
	LUT2 #(
		.INIT('h1)
	) name3 (
		_w1509_,
		_w1510_,
		_w1511_
	);
	LUT2 #(
		.INIT('h2)
	) name4 (
		\WX707_reg/NET0131 ,
		\WX771_reg/NET0131 ,
		_w1512_
	);
	LUT2 #(
		.INIT('h4)
	) name5 (
		\WX707_reg/NET0131 ,
		\WX771_reg/NET0131 ,
		_w1513_
	);
	LUT2 #(
		.INIT('h1)
	) name6 (
		_w1512_,
		_w1513_,
		_w1514_
	);
	LUT2 #(
		.INIT('h8)
	) name7 (
		_w1511_,
		_w1514_,
		_w1515_
	);
	LUT2 #(
		.INIT('h1)
	) name8 (
		_w1511_,
		_w1514_,
		_w1516_
	);
	LUT2 #(
		.INIT('h1)
	) name9 (
		_w1515_,
		_w1516_,
		_w1517_
	);
	LUT2 #(
		.INIT('h8)
	) name10 (
		_w1508_,
		_w1517_,
		_w1518_
	);
	LUT2 #(
		.INIT('h1)
	) name11 (
		_w1508_,
		_w1517_,
		_w1519_
	);
	LUT2 #(
		.INIT('h1)
	) name12 (
		_w1518_,
		_w1519_,
		_w1520_
	);
	LUT2 #(
		.INIT('h2)
	) name13 (
		\TM0_pad ,
		\WX10871_reg/NET0131 ,
		_w1521_
	);
	LUT2 #(
		.INIT('h2)
	) name14 (
		\WX815_reg/NET0131 ,
		\WX879_reg/NET0131 ,
		_w1522_
	);
	LUT2 #(
		.INIT('h4)
	) name15 (
		\WX815_reg/NET0131 ,
		\WX879_reg/NET0131 ,
		_w1523_
	);
	LUT2 #(
		.INIT('h1)
	) name16 (
		_w1522_,
		_w1523_,
		_w1524_
	);
	LUT2 #(
		.INIT('h2)
	) name17 (
		\WX687_reg/NET0131 ,
		\WX751_reg/NET0131 ,
		_w1525_
	);
	LUT2 #(
		.INIT('h4)
	) name18 (
		\WX687_reg/NET0131 ,
		\WX751_reg/NET0131 ,
		_w1526_
	);
	LUT2 #(
		.INIT('h1)
	) name19 (
		_w1525_,
		_w1526_,
		_w1527_
	);
	LUT2 #(
		.INIT('h8)
	) name20 (
		_w1524_,
		_w1527_,
		_w1528_
	);
	LUT2 #(
		.INIT('h1)
	) name21 (
		_w1524_,
		_w1527_,
		_w1529_
	);
	LUT2 #(
		.INIT('h1)
	) name22 (
		_w1528_,
		_w1529_,
		_w1530_
	);
	LUT2 #(
		.INIT('h8)
	) name23 (
		_w1521_,
		_w1530_,
		_w1531_
	);
	LUT2 #(
		.INIT('h1)
	) name24 (
		_w1521_,
		_w1530_,
		_w1532_
	);
	LUT2 #(
		.INIT('h1)
	) name25 (
		_w1531_,
		_w1532_,
		_w1533_
	);
	LUT2 #(
		.INIT('h2)
	) name26 (
		\TM0_pad ,
		\WX10869_reg/NET0131 ,
		_w1534_
	);
	LUT2 #(
		.INIT('h2)
	) name27 (
		\WX813_reg/NET0131 ,
		\WX877_reg/NET0131 ,
		_w1535_
	);
	LUT2 #(
		.INIT('h4)
	) name28 (
		\WX813_reg/NET0131 ,
		\WX877_reg/NET0131 ,
		_w1536_
	);
	LUT2 #(
		.INIT('h1)
	) name29 (
		_w1535_,
		_w1536_,
		_w1537_
	);
	LUT2 #(
		.INIT('h2)
	) name30 (
		\WX685_reg/NET0131 ,
		\WX749_reg/NET0131 ,
		_w1538_
	);
	LUT2 #(
		.INIT('h4)
	) name31 (
		\WX685_reg/NET0131 ,
		\WX749_reg/NET0131 ,
		_w1539_
	);
	LUT2 #(
		.INIT('h1)
	) name32 (
		_w1538_,
		_w1539_,
		_w1540_
	);
	LUT2 #(
		.INIT('h8)
	) name33 (
		_w1537_,
		_w1540_,
		_w1541_
	);
	LUT2 #(
		.INIT('h1)
	) name34 (
		_w1537_,
		_w1540_,
		_w1542_
	);
	LUT2 #(
		.INIT('h1)
	) name35 (
		_w1541_,
		_w1542_,
		_w1543_
	);
	LUT2 #(
		.INIT('h8)
	) name36 (
		_w1534_,
		_w1543_,
		_w1544_
	);
	LUT2 #(
		.INIT('h1)
	) name37 (
		_w1534_,
		_w1543_,
		_w1545_
	);
	LUT2 #(
		.INIT('h1)
	) name38 (
		_w1544_,
		_w1545_,
		_w1546_
	);
	LUT2 #(
		.INIT('h2)
	) name39 (
		\TM0_pad ,
		\WX10867_reg/NET0131 ,
		_w1547_
	);
	LUT2 #(
		.INIT('h2)
	) name40 (
		\WX811_reg/NET0131 ,
		\WX875_reg/NET0131 ,
		_w1548_
	);
	LUT2 #(
		.INIT('h4)
	) name41 (
		\WX811_reg/NET0131 ,
		\WX875_reg/NET0131 ,
		_w1549_
	);
	LUT2 #(
		.INIT('h1)
	) name42 (
		_w1548_,
		_w1549_,
		_w1550_
	);
	LUT2 #(
		.INIT('h2)
	) name43 (
		\WX683_reg/NET0131 ,
		\WX747_reg/NET0131 ,
		_w1551_
	);
	LUT2 #(
		.INIT('h4)
	) name44 (
		\WX683_reg/NET0131 ,
		\WX747_reg/NET0131 ,
		_w1552_
	);
	LUT2 #(
		.INIT('h1)
	) name45 (
		_w1551_,
		_w1552_,
		_w1553_
	);
	LUT2 #(
		.INIT('h8)
	) name46 (
		_w1550_,
		_w1553_,
		_w1554_
	);
	LUT2 #(
		.INIT('h1)
	) name47 (
		_w1550_,
		_w1553_,
		_w1555_
	);
	LUT2 #(
		.INIT('h1)
	) name48 (
		_w1554_,
		_w1555_,
		_w1556_
	);
	LUT2 #(
		.INIT('h8)
	) name49 (
		_w1547_,
		_w1556_,
		_w1557_
	);
	LUT2 #(
		.INIT('h1)
	) name50 (
		_w1547_,
		_w1556_,
		_w1558_
	);
	LUT2 #(
		.INIT('h1)
	) name51 (
		_w1557_,
		_w1558_,
		_w1559_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		\TM0_pad ,
		\WX10865_reg/NET0131 ,
		_w1560_
	);
	LUT2 #(
		.INIT('h2)
	) name53 (
		\WX809_reg/NET0131 ,
		\WX873_reg/NET0131 ,
		_w1561_
	);
	LUT2 #(
		.INIT('h4)
	) name54 (
		\WX809_reg/NET0131 ,
		\WX873_reg/NET0131 ,
		_w1562_
	);
	LUT2 #(
		.INIT('h1)
	) name55 (
		_w1561_,
		_w1562_,
		_w1563_
	);
	LUT2 #(
		.INIT('h2)
	) name56 (
		\WX681_reg/NET0131 ,
		\WX745_reg/NET0131 ,
		_w1564_
	);
	LUT2 #(
		.INIT('h4)
	) name57 (
		\WX681_reg/NET0131 ,
		\WX745_reg/NET0131 ,
		_w1565_
	);
	LUT2 #(
		.INIT('h1)
	) name58 (
		_w1564_,
		_w1565_,
		_w1566_
	);
	LUT2 #(
		.INIT('h8)
	) name59 (
		_w1563_,
		_w1566_,
		_w1567_
	);
	LUT2 #(
		.INIT('h1)
	) name60 (
		_w1563_,
		_w1566_,
		_w1568_
	);
	LUT2 #(
		.INIT('h1)
	) name61 (
		_w1567_,
		_w1568_,
		_w1569_
	);
	LUT2 #(
		.INIT('h8)
	) name62 (
		_w1560_,
		_w1569_,
		_w1570_
	);
	LUT2 #(
		.INIT('h1)
	) name63 (
		_w1560_,
		_w1569_,
		_w1571_
	);
	LUT2 #(
		.INIT('h1)
	) name64 (
		_w1570_,
		_w1571_,
		_w1572_
	);
	LUT2 #(
		.INIT('h2)
	) name65 (
		\TM0_pad ,
		\WX10863_reg/NET0131 ,
		_w1573_
	);
	LUT2 #(
		.INIT('h2)
	) name66 (
		\WX807_reg/NET0131 ,
		\WX871_reg/NET0131 ,
		_w1574_
	);
	LUT2 #(
		.INIT('h4)
	) name67 (
		\WX807_reg/NET0131 ,
		\WX871_reg/NET0131 ,
		_w1575_
	);
	LUT2 #(
		.INIT('h1)
	) name68 (
		_w1574_,
		_w1575_,
		_w1576_
	);
	LUT2 #(
		.INIT('h2)
	) name69 (
		\WX679_reg/NET0131 ,
		\WX743_reg/NET0131 ,
		_w1577_
	);
	LUT2 #(
		.INIT('h4)
	) name70 (
		\WX679_reg/NET0131 ,
		\WX743_reg/NET0131 ,
		_w1578_
	);
	LUT2 #(
		.INIT('h1)
	) name71 (
		_w1577_,
		_w1578_,
		_w1579_
	);
	LUT2 #(
		.INIT('h8)
	) name72 (
		_w1576_,
		_w1579_,
		_w1580_
	);
	LUT2 #(
		.INIT('h1)
	) name73 (
		_w1576_,
		_w1579_,
		_w1581_
	);
	LUT2 #(
		.INIT('h1)
	) name74 (
		_w1580_,
		_w1581_,
		_w1582_
	);
	LUT2 #(
		.INIT('h8)
	) name75 (
		_w1573_,
		_w1582_,
		_w1583_
	);
	LUT2 #(
		.INIT('h1)
	) name76 (
		_w1573_,
		_w1582_,
		_w1584_
	);
	LUT2 #(
		.INIT('h1)
	) name77 (
		_w1583_,
		_w1584_,
		_w1585_
	);
	LUT2 #(
		.INIT('h2)
	) name78 (
		\TM0_pad ,
		\WX10861_reg/NET0131 ,
		_w1586_
	);
	LUT2 #(
		.INIT('h2)
	) name79 (
		\WX805_reg/NET0131 ,
		\WX869_reg/NET0131 ,
		_w1587_
	);
	LUT2 #(
		.INIT('h4)
	) name80 (
		\WX805_reg/NET0131 ,
		\WX869_reg/NET0131 ,
		_w1588_
	);
	LUT2 #(
		.INIT('h1)
	) name81 (
		_w1587_,
		_w1588_,
		_w1589_
	);
	LUT2 #(
		.INIT('h2)
	) name82 (
		\WX677_reg/NET0131 ,
		\WX741_reg/NET0131 ,
		_w1590_
	);
	LUT2 #(
		.INIT('h4)
	) name83 (
		\WX677_reg/NET0131 ,
		\WX741_reg/NET0131 ,
		_w1591_
	);
	LUT2 #(
		.INIT('h1)
	) name84 (
		_w1590_,
		_w1591_,
		_w1592_
	);
	LUT2 #(
		.INIT('h8)
	) name85 (
		_w1589_,
		_w1592_,
		_w1593_
	);
	LUT2 #(
		.INIT('h1)
	) name86 (
		_w1589_,
		_w1592_,
		_w1594_
	);
	LUT2 #(
		.INIT('h1)
	) name87 (
		_w1593_,
		_w1594_,
		_w1595_
	);
	LUT2 #(
		.INIT('h8)
	) name88 (
		_w1586_,
		_w1595_,
		_w1596_
	);
	LUT2 #(
		.INIT('h1)
	) name89 (
		_w1586_,
		_w1595_,
		_w1597_
	);
	LUT2 #(
		.INIT('h1)
	) name90 (
		_w1596_,
		_w1597_,
		_w1598_
	);
	LUT2 #(
		.INIT('h2)
	) name91 (
		\WX803_reg/NET0131 ,
		\WX867_reg/NET0131 ,
		_w1599_
	);
	LUT2 #(
		.INIT('h4)
	) name92 (
		\WX803_reg/NET0131 ,
		\WX867_reg/NET0131 ,
		_w1600_
	);
	LUT2 #(
		.INIT('h1)
	) name93 (
		_w1599_,
		_w1600_,
		_w1601_
	);
	LUT2 #(
		.INIT('h2)
	) name94 (
		\WX739_reg/NET0131 ,
		_w1601_,
		_w1602_
	);
	LUT2 #(
		.INIT('h4)
	) name95 (
		\WX739_reg/NET0131 ,
		_w1601_,
		_w1603_
	);
	LUT2 #(
		.INIT('h1)
	) name96 (
		_w1602_,
		_w1603_,
		_w1604_
	);
	LUT2 #(
		.INIT('h8)
	) name97 (
		\TM0_pad ,
		\WX10859_reg/NET0131 ,
		_w1605_
	);
	LUT2 #(
		.INIT('h1)
	) name98 (
		\TM1_pad ,
		\WX675_reg/NET0131 ,
		_w1606_
	);
	LUT2 #(
		.INIT('h8)
	) name99 (
		\TM1_pad ,
		\WX675_reg/NET0131 ,
		_w1607_
	);
	LUT2 #(
		.INIT('h1)
	) name100 (
		_w1606_,
		_w1607_,
		_w1608_
	);
	LUT2 #(
		.INIT('h2)
	) name101 (
		_w1605_,
		_w1608_,
		_w1609_
	);
	LUT2 #(
		.INIT('h4)
	) name102 (
		_w1605_,
		_w1608_,
		_w1610_
	);
	LUT2 #(
		.INIT('h1)
	) name103 (
		_w1609_,
		_w1610_,
		_w1611_
	);
	LUT2 #(
		.INIT('h8)
	) name104 (
		_w1604_,
		_w1611_,
		_w1612_
	);
	LUT2 #(
		.INIT('h1)
	) name105 (
		_w1604_,
		_w1611_,
		_w1613_
	);
	LUT2 #(
		.INIT('h1)
	) name106 (
		_w1612_,
		_w1613_,
		_w1614_
	);
	LUT2 #(
		.INIT('h2)
	) name107 (
		\WX801_reg/NET0131 ,
		\WX865_reg/NET0131 ,
		_w1615_
	);
	LUT2 #(
		.INIT('h4)
	) name108 (
		\WX801_reg/NET0131 ,
		\WX865_reg/NET0131 ,
		_w1616_
	);
	LUT2 #(
		.INIT('h1)
	) name109 (
		_w1615_,
		_w1616_,
		_w1617_
	);
	LUT2 #(
		.INIT('h2)
	) name110 (
		\WX737_reg/NET0131 ,
		_w1617_,
		_w1618_
	);
	LUT2 #(
		.INIT('h4)
	) name111 (
		\WX737_reg/NET0131 ,
		_w1617_,
		_w1619_
	);
	LUT2 #(
		.INIT('h1)
	) name112 (
		_w1618_,
		_w1619_,
		_w1620_
	);
	LUT2 #(
		.INIT('h8)
	) name113 (
		\TM0_pad ,
		\WX10857_reg/NET0131 ,
		_w1621_
	);
	LUT2 #(
		.INIT('h1)
	) name114 (
		\TM1_pad ,
		\WX673_reg/NET0131 ,
		_w1622_
	);
	LUT2 #(
		.INIT('h8)
	) name115 (
		\TM1_pad ,
		\WX673_reg/NET0131 ,
		_w1623_
	);
	LUT2 #(
		.INIT('h1)
	) name116 (
		_w1622_,
		_w1623_,
		_w1624_
	);
	LUT2 #(
		.INIT('h2)
	) name117 (
		_w1621_,
		_w1624_,
		_w1625_
	);
	LUT2 #(
		.INIT('h4)
	) name118 (
		_w1621_,
		_w1624_,
		_w1626_
	);
	LUT2 #(
		.INIT('h1)
	) name119 (
		_w1625_,
		_w1626_,
		_w1627_
	);
	LUT2 #(
		.INIT('h8)
	) name120 (
		_w1620_,
		_w1627_,
		_w1628_
	);
	LUT2 #(
		.INIT('h1)
	) name121 (
		_w1620_,
		_w1627_,
		_w1629_
	);
	LUT2 #(
		.INIT('h1)
	) name122 (
		_w1628_,
		_w1629_,
		_w1630_
	);
	LUT2 #(
		.INIT('h2)
	) name123 (
		\WX799_reg/NET0131 ,
		\WX863_reg/NET0131 ,
		_w1631_
	);
	LUT2 #(
		.INIT('h4)
	) name124 (
		\WX799_reg/NET0131 ,
		\WX863_reg/NET0131 ,
		_w1632_
	);
	LUT2 #(
		.INIT('h1)
	) name125 (
		_w1631_,
		_w1632_,
		_w1633_
	);
	LUT2 #(
		.INIT('h2)
	) name126 (
		\WX735_reg/NET0131 ,
		_w1633_,
		_w1634_
	);
	LUT2 #(
		.INIT('h4)
	) name127 (
		\WX735_reg/NET0131 ,
		_w1633_,
		_w1635_
	);
	LUT2 #(
		.INIT('h1)
	) name128 (
		_w1634_,
		_w1635_,
		_w1636_
	);
	LUT2 #(
		.INIT('h8)
	) name129 (
		\TM0_pad ,
		\WX10855_reg/NET0131 ,
		_w1637_
	);
	LUT2 #(
		.INIT('h1)
	) name130 (
		\TM1_pad ,
		\WX671_reg/NET0131 ,
		_w1638_
	);
	LUT2 #(
		.INIT('h8)
	) name131 (
		\TM1_pad ,
		\WX671_reg/NET0131 ,
		_w1639_
	);
	LUT2 #(
		.INIT('h1)
	) name132 (
		_w1638_,
		_w1639_,
		_w1640_
	);
	LUT2 #(
		.INIT('h2)
	) name133 (
		_w1637_,
		_w1640_,
		_w1641_
	);
	LUT2 #(
		.INIT('h4)
	) name134 (
		_w1637_,
		_w1640_,
		_w1642_
	);
	LUT2 #(
		.INIT('h1)
	) name135 (
		_w1641_,
		_w1642_,
		_w1643_
	);
	LUT2 #(
		.INIT('h8)
	) name136 (
		_w1636_,
		_w1643_,
		_w1644_
	);
	LUT2 #(
		.INIT('h1)
	) name137 (
		_w1636_,
		_w1643_,
		_w1645_
	);
	LUT2 #(
		.INIT('h1)
	) name138 (
		_w1644_,
		_w1645_,
		_w1646_
	);
	LUT2 #(
		.INIT('h2)
	) name139 (
		\WX797_reg/NET0131 ,
		\WX861_reg/NET0131 ,
		_w1647_
	);
	LUT2 #(
		.INIT('h4)
	) name140 (
		\WX797_reg/NET0131 ,
		\WX861_reg/NET0131 ,
		_w1648_
	);
	LUT2 #(
		.INIT('h1)
	) name141 (
		_w1647_,
		_w1648_,
		_w1649_
	);
	LUT2 #(
		.INIT('h2)
	) name142 (
		\WX733_reg/NET0131 ,
		_w1649_,
		_w1650_
	);
	LUT2 #(
		.INIT('h4)
	) name143 (
		\WX733_reg/NET0131 ,
		_w1649_,
		_w1651_
	);
	LUT2 #(
		.INIT('h1)
	) name144 (
		_w1650_,
		_w1651_,
		_w1652_
	);
	LUT2 #(
		.INIT('h8)
	) name145 (
		\TM0_pad ,
		\WX10853_reg/NET0131 ,
		_w1653_
	);
	LUT2 #(
		.INIT('h1)
	) name146 (
		\TM1_pad ,
		\WX669_reg/NET0131 ,
		_w1654_
	);
	LUT2 #(
		.INIT('h8)
	) name147 (
		\TM1_pad ,
		\WX669_reg/NET0131 ,
		_w1655_
	);
	LUT2 #(
		.INIT('h1)
	) name148 (
		_w1654_,
		_w1655_,
		_w1656_
	);
	LUT2 #(
		.INIT('h2)
	) name149 (
		_w1653_,
		_w1656_,
		_w1657_
	);
	LUT2 #(
		.INIT('h4)
	) name150 (
		_w1653_,
		_w1656_,
		_w1658_
	);
	LUT2 #(
		.INIT('h1)
	) name151 (
		_w1657_,
		_w1658_,
		_w1659_
	);
	LUT2 #(
		.INIT('h8)
	) name152 (
		_w1652_,
		_w1659_,
		_w1660_
	);
	LUT2 #(
		.INIT('h1)
	) name153 (
		_w1652_,
		_w1659_,
		_w1661_
	);
	LUT2 #(
		.INIT('h1)
	) name154 (
		_w1660_,
		_w1661_,
		_w1662_
	);
	LUT2 #(
		.INIT('h2)
	) name155 (
		\TM0_pad ,
		\WX10889_reg/NET0131 ,
		_w1663_
	);
	LUT2 #(
		.INIT('h2)
	) name156 (
		\WX833_reg/NET0131 ,
		\WX897_reg/NET0131 ,
		_w1664_
	);
	LUT2 #(
		.INIT('h4)
	) name157 (
		\WX833_reg/NET0131 ,
		\WX897_reg/NET0131 ,
		_w1665_
	);
	LUT2 #(
		.INIT('h1)
	) name158 (
		_w1664_,
		_w1665_,
		_w1666_
	);
	LUT2 #(
		.INIT('h2)
	) name159 (
		\WX705_reg/NET0131 ,
		\WX769_reg/NET0131 ,
		_w1667_
	);
	LUT2 #(
		.INIT('h4)
	) name160 (
		\WX705_reg/NET0131 ,
		\WX769_reg/NET0131 ,
		_w1668_
	);
	LUT2 #(
		.INIT('h1)
	) name161 (
		_w1667_,
		_w1668_,
		_w1669_
	);
	LUT2 #(
		.INIT('h8)
	) name162 (
		_w1666_,
		_w1669_,
		_w1670_
	);
	LUT2 #(
		.INIT('h1)
	) name163 (
		_w1666_,
		_w1669_,
		_w1671_
	);
	LUT2 #(
		.INIT('h1)
	) name164 (
		_w1670_,
		_w1671_,
		_w1672_
	);
	LUT2 #(
		.INIT('h8)
	) name165 (
		_w1663_,
		_w1672_,
		_w1673_
	);
	LUT2 #(
		.INIT('h1)
	) name166 (
		_w1663_,
		_w1672_,
		_w1674_
	);
	LUT2 #(
		.INIT('h1)
	) name167 (
		_w1673_,
		_w1674_,
		_w1675_
	);
	LUT2 #(
		.INIT('h2)
	) name168 (
		\WX795_reg/NET0131 ,
		\WX859_reg/NET0131 ,
		_w1676_
	);
	LUT2 #(
		.INIT('h4)
	) name169 (
		\WX795_reg/NET0131 ,
		\WX859_reg/NET0131 ,
		_w1677_
	);
	LUT2 #(
		.INIT('h1)
	) name170 (
		_w1676_,
		_w1677_,
		_w1678_
	);
	LUT2 #(
		.INIT('h2)
	) name171 (
		\WX731_reg/NET0131 ,
		_w1678_,
		_w1679_
	);
	LUT2 #(
		.INIT('h4)
	) name172 (
		\WX731_reg/NET0131 ,
		_w1678_,
		_w1680_
	);
	LUT2 #(
		.INIT('h1)
	) name173 (
		_w1679_,
		_w1680_,
		_w1681_
	);
	LUT2 #(
		.INIT('h8)
	) name174 (
		\TM0_pad ,
		\WX10851_reg/NET0131 ,
		_w1682_
	);
	LUT2 #(
		.INIT('h1)
	) name175 (
		\TM1_pad ,
		\WX667_reg/NET0131 ,
		_w1683_
	);
	LUT2 #(
		.INIT('h8)
	) name176 (
		\TM1_pad ,
		\WX667_reg/NET0131 ,
		_w1684_
	);
	LUT2 #(
		.INIT('h1)
	) name177 (
		_w1683_,
		_w1684_,
		_w1685_
	);
	LUT2 #(
		.INIT('h2)
	) name178 (
		_w1682_,
		_w1685_,
		_w1686_
	);
	LUT2 #(
		.INIT('h4)
	) name179 (
		_w1682_,
		_w1685_,
		_w1687_
	);
	LUT2 #(
		.INIT('h1)
	) name180 (
		_w1686_,
		_w1687_,
		_w1688_
	);
	LUT2 #(
		.INIT('h8)
	) name181 (
		_w1681_,
		_w1688_,
		_w1689_
	);
	LUT2 #(
		.INIT('h1)
	) name182 (
		_w1681_,
		_w1688_,
		_w1690_
	);
	LUT2 #(
		.INIT('h1)
	) name183 (
		_w1689_,
		_w1690_,
		_w1691_
	);
	LUT2 #(
		.INIT('h2)
	) name184 (
		\WX793_reg/NET0131 ,
		\WX857_reg/NET0131 ,
		_w1692_
	);
	LUT2 #(
		.INIT('h4)
	) name185 (
		\WX793_reg/NET0131 ,
		\WX857_reg/NET0131 ,
		_w1693_
	);
	LUT2 #(
		.INIT('h1)
	) name186 (
		_w1692_,
		_w1693_,
		_w1694_
	);
	LUT2 #(
		.INIT('h2)
	) name187 (
		\WX729_reg/NET0131 ,
		_w1694_,
		_w1695_
	);
	LUT2 #(
		.INIT('h4)
	) name188 (
		\WX729_reg/NET0131 ,
		_w1694_,
		_w1696_
	);
	LUT2 #(
		.INIT('h1)
	) name189 (
		_w1695_,
		_w1696_,
		_w1697_
	);
	LUT2 #(
		.INIT('h8)
	) name190 (
		\TM0_pad ,
		\WX10849_reg/NET0131 ,
		_w1698_
	);
	LUT2 #(
		.INIT('h1)
	) name191 (
		\TM1_pad ,
		\WX665_reg/NET0131 ,
		_w1699_
	);
	LUT2 #(
		.INIT('h8)
	) name192 (
		\TM1_pad ,
		\WX665_reg/NET0131 ,
		_w1700_
	);
	LUT2 #(
		.INIT('h1)
	) name193 (
		_w1699_,
		_w1700_,
		_w1701_
	);
	LUT2 #(
		.INIT('h2)
	) name194 (
		_w1698_,
		_w1701_,
		_w1702_
	);
	LUT2 #(
		.INIT('h4)
	) name195 (
		_w1698_,
		_w1701_,
		_w1703_
	);
	LUT2 #(
		.INIT('h1)
	) name196 (
		_w1702_,
		_w1703_,
		_w1704_
	);
	LUT2 #(
		.INIT('h8)
	) name197 (
		_w1697_,
		_w1704_,
		_w1705_
	);
	LUT2 #(
		.INIT('h1)
	) name198 (
		_w1697_,
		_w1704_,
		_w1706_
	);
	LUT2 #(
		.INIT('h1)
	) name199 (
		_w1705_,
		_w1706_,
		_w1707_
	);
	LUT2 #(
		.INIT('h2)
	) name200 (
		\WX791_reg/NET0131 ,
		\WX855_reg/NET0131 ,
		_w1708_
	);
	LUT2 #(
		.INIT('h4)
	) name201 (
		\WX791_reg/NET0131 ,
		\WX855_reg/NET0131 ,
		_w1709_
	);
	LUT2 #(
		.INIT('h1)
	) name202 (
		_w1708_,
		_w1709_,
		_w1710_
	);
	LUT2 #(
		.INIT('h2)
	) name203 (
		\WX727_reg/NET0131 ,
		_w1710_,
		_w1711_
	);
	LUT2 #(
		.INIT('h4)
	) name204 (
		\WX727_reg/NET0131 ,
		_w1710_,
		_w1712_
	);
	LUT2 #(
		.INIT('h1)
	) name205 (
		_w1711_,
		_w1712_,
		_w1713_
	);
	LUT2 #(
		.INIT('h8)
	) name206 (
		\TM0_pad ,
		\WX10847_reg/NET0131 ,
		_w1714_
	);
	LUT2 #(
		.INIT('h1)
	) name207 (
		\TM1_pad ,
		\WX663_reg/NET0131 ,
		_w1715_
	);
	LUT2 #(
		.INIT('h8)
	) name208 (
		\TM1_pad ,
		\WX663_reg/NET0131 ,
		_w1716_
	);
	LUT2 #(
		.INIT('h1)
	) name209 (
		_w1715_,
		_w1716_,
		_w1717_
	);
	LUT2 #(
		.INIT('h2)
	) name210 (
		_w1714_,
		_w1717_,
		_w1718_
	);
	LUT2 #(
		.INIT('h4)
	) name211 (
		_w1714_,
		_w1717_,
		_w1719_
	);
	LUT2 #(
		.INIT('h1)
	) name212 (
		_w1718_,
		_w1719_,
		_w1720_
	);
	LUT2 #(
		.INIT('h8)
	) name213 (
		_w1713_,
		_w1720_,
		_w1721_
	);
	LUT2 #(
		.INIT('h1)
	) name214 (
		_w1713_,
		_w1720_,
		_w1722_
	);
	LUT2 #(
		.INIT('h1)
	) name215 (
		_w1721_,
		_w1722_,
		_w1723_
	);
	LUT2 #(
		.INIT('h2)
	) name216 (
		\WX789_reg/NET0131 ,
		\WX853_reg/NET0131 ,
		_w1724_
	);
	LUT2 #(
		.INIT('h4)
	) name217 (
		\WX789_reg/NET0131 ,
		\WX853_reg/NET0131 ,
		_w1725_
	);
	LUT2 #(
		.INIT('h1)
	) name218 (
		_w1724_,
		_w1725_,
		_w1726_
	);
	LUT2 #(
		.INIT('h2)
	) name219 (
		\WX725_reg/NET0131 ,
		_w1726_,
		_w1727_
	);
	LUT2 #(
		.INIT('h4)
	) name220 (
		\WX725_reg/NET0131 ,
		_w1726_,
		_w1728_
	);
	LUT2 #(
		.INIT('h1)
	) name221 (
		_w1727_,
		_w1728_,
		_w1729_
	);
	LUT2 #(
		.INIT('h8)
	) name222 (
		\TM0_pad ,
		\WX10845_reg/NET0131 ,
		_w1730_
	);
	LUT2 #(
		.INIT('h1)
	) name223 (
		\TM1_pad ,
		\WX661_reg/NET0131 ,
		_w1731_
	);
	LUT2 #(
		.INIT('h8)
	) name224 (
		\TM1_pad ,
		\WX661_reg/NET0131 ,
		_w1732_
	);
	LUT2 #(
		.INIT('h1)
	) name225 (
		_w1731_,
		_w1732_,
		_w1733_
	);
	LUT2 #(
		.INIT('h2)
	) name226 (
		_w1730_,
		_w1733_,
		_w1734_
	);
	LUT2 #(
		.INIT('h4)
	) name227 (
		_w1730_,
		_w1733_,
		_w1735_
	);
	LUT2 #(
		.INIT('h1)
	) name228 (
		_w1734_,
		_w1735_,
		_w1736_
	);
	LUT2 #(
		.INIT('h8)
	) name229 (
		_w1729_,
		_w1736_,
		_w1737_
	);
	LUT2 #(
		.INIT('h1)
	) name230 (
		_w1729_,
		_w1736_,
		_w1738_
	);
	LUT2 #(
		.INIT('h1)
	) name231 (
		_w1737_,
		_w1738_,
		_w1739_
	);
	LUT2 #(
		.INIT('h2)
	) name232 (
		\WX787_reg/NET0131 ,
		\WX851_reg/NET0131 ,
		_w1740_
	);
	LUT2 #(
		.INIT('h4)
	) name233 (
		\WX787_reg/NET0131 ,
		\WX851_reg/NET0131 ,
		_w1741_
	);
	LUT2 #(
		.INIT('h1)
	) name234 (
		_w1740_,
		_w1741_,
		_w1742_
	);
	LUT2 #(
		.INIT('h2)
	) name235 (
		\WX723_reg/NET0131 ,
		_w1742_,
		_w1743_
	);
	LUT2 #(
		.INIT('h4)
	) name236 (
		\WX723_reg/NET0131 ,
		_w1742_,
		_w1744_
	);
	LUT2 #(
		.INIT('h1)
	) name237 (
		_w1743_,
		_w1744_,
		_w1745_
	);
	LUT2 #(
		.INIT('h8)
	) name238 (
		\TM0_pad ,
		\WX10843_reg/NET0131 ,
		_w1746_
	);
	LUT2 #(
		.INIT('h1)
	) name239 (
		\TM1_pad ,
		\WX659_reg/NET0131 ,
		_w1747_
	);
	LUT2 #(
		.INIT('h8)
	) name240 (
		\TM1_pad ,
		\WX659_reg/NET0131 ,
		_w1748_
	);
	LUT2 #(
		.INIT('h1)
	) name241 (
		_w1747_,
		_w1748_,
		_w1749_
	);
	LUT2 #(
		.INIT('h2)
	) name242 (
		_w1746_,
		_w1749_,
		_w1750_
	);
	LUT2 #(
		.INIT('h4)
	) name243 (
		_w1746_,
		_w1749_,
		_w1751_
	);
	LUT2 #(
		.INIT('h1)
	) name244 (
		_w1750_,
		_w1751_,
		_w1752_
	);
	LUT2 #(
		.INIT('h8)
	) name245 (
		_w1745_,
		_w1752_,
		_w1753_
	);
	LUT2 #(
		.INIT('h1)
	) name246 (
		_w1745_,
		_w1752_,
		_w1754_
	);
	LUT2 #(
		.INIT('h1)
	) name247 (
		_w1753_,
		_w1754_,
		_w1755_
	);
	LUT2 #(
		.INIT('h2)
	) name248 (
		\WX785_reg/NET0131 ,
		\WX849_reg/NET0131 ,
		_w1756_
	);
	LUT2 #(
		.INIT('h4)
	) name249 (
		\WX785_reg/NET0131 ,
		\WX849_reg/NET0131 ,
		_w1757_
	);
	LUT2 #(
		.INIT('h1)
	) name250 (
		_w1756_,
		_w1757_,
		_w1758_
	);
	LUT2 #(
		.INIT('h2)
	) name251 (
		\WX721_reg/NET0131 ,
		_w1758_,
		_w1759_
	);
	LUT2 #(
		.INIT('h4)
	) name252 (
		\WX721_reg/NET0131 ,
		_w1758_,
		_w1760_
	);
	LUT2 #(
		.INIT('h1)
	) name253 (
		_w1759_,
		_w1760_,
		_w1761_
	);
	LUT2 #(
		.INIT('h8)
	) name254 (
		\TM0_pad ,
		\WX10841_reg/NET0131 ,
		_w1762_
	);
	LUT2 #(
		.INIT('h1)
	) name255 (
		\TM1_pad ,
		\WX657_reg/NET0131 ,
		_w1763_
	);
	LUT2 #(
		.INIT('h8)
	) name256 (
		\TM1_pad ,
		\WX657_reg/NET0131 ,
		_w1764_
	);
	LUT2 #(
		.INIT('h1)
	) name257 (
		_w1763_,
		_w1764_,
		_w1765_
	);
	LUT2 #(
		.INIT('h2)
	) name258 (
		_w1762_,
		_w1765_,
		_w1766_
	);
	LUT2 #(
		.INIT('h4)
	) name259 (
		_w1762_,
		_w1765_,
		_w1767_
	);
	LUT2 #(
		.INIT('h1)
	) name260 (
		_w1766_,
		_w1767_,
		_w1768_
	);
	LUT2 #(
		.INIT('h8)
	) name261 (
		_w1761_,
		_w1768_,
		_w1769_
	);
	LUT2 #(
		.INIT('h1)
	) name262 (
		_w1761_,
		_w1768_,
		_w1770_
	);
	LUT2 #(
		.INIT('h1)
	) name263 (
		_w1769_,
		_w1770_,
		_w1771_
	);
	LUT2 #(
		.INIT('h2)
	) name264 (
		\WX783_reg/NET0131 ,
		\WX847_reg/NET0131 ,
		_w1772_
	);
	LUT2 #(
		.INIT('h4)
	) name265 (
		\WX783_reg/NET0131 ,
		\WX847_reg/NET0131 ,
		_w1773_
	);
	LUT2 #(
		.INIT('h1)
	) name266 (
		_w1772_,
		_w1773_,
		_w1774_
	);
	LUT2 #(
		.INIT('h2)
	) name267 (
		\WX719_reg/NET0131 ,
		_w1774_,
		_w1775_
	);
	LUT2 #(
		.INIT('h4)
	) name268 (
		\WX719_reg/NET0131 ,
		_w1774_,
		_w1776_
	);
	LUT2 #(
		.INIT('h1)
	) name269 (
		_w1775_,
		_w1776_,
		_w1777_
	);
	LUT2 #(
		.INIT('h8)
	) name270 (
		\TM0_pad ,
		\WX10839_reg/NET0131 ,
		_w1778_
	);
	LUT2 #(
		.INIT('h1)
	) name271 (
		\TM1_pad ,
		\WX655_reg/NET0131 ,
		_w1779_
	);
	LUT2 #(
		.INIT('h8)
	) name272 (
		\TM1_pad ,
		\WX655_reg/NET0131 ,
		_w1780_
	);
	LUT2 #(
		.INIT('h1)
	) name273 (
		_w1779_,
		_w1780_,
		_w1781_
	);
	LUT2 #(
		.INIT('h2)
	) name274 (
		_w1778_,
		_w1781_,
		_w1782_
	);
	LUT2 #(
		.INIT('h4)
	) name275 (
		_w1778_,
		_w1781_,
		_w1783_
	);
	LUT2 #(
		.INIT('h1)
	) name276 (
		_w1782_,
		_w1783_,
		_w1784_
	);
	LUT2 #(
		.INIT('h8)
	) name277 (
		_w1777_,
		_w1784_,
		_w1785_
	);
	LUT2 #(
		.INIT('h1)
	) name278 (
		_w1777_,
		_w1784_,
		_w1786_
	);
	LUT2 #(
		.INIT('h1)
	) name279 (
		_w1785_,
		_w1786_,
		_w1787_
	);
	LUT2 #(
		.INIT('h2)
	) name280 (
		\WX781_reg/NET0131 ,
		\WX845_reg/NET0131 ,
		_w1788_
	);
	LUT2 #(
		.INIT('h4)
	) name281 (
		\WX781_reg/NET0131 ,
		\WX845_reg/NET0131 ,
		_w1789_
	);
	LUT2 #(
		.INIT('h1)
	) name282 (
		_w1788_,
		_w1789_,
		_w1790_
	);
	LUT2 #(
		.INIT('h2)
	) name283 (
		\WX717_reg/NET0131 ,
		_w1790_,
		_w1791_
	);
	LUT2 #(
		.INIT('h4)
	) name284 (
		\WX717_reg/NET0131 ,
		_w1790_,
		_w1792_
	);
	LUT2 #(
		.INIT('h1)
	) name285 (
		_w1791_,
		_w1792_,
		_w1793_
	);
	LUT2 #(
		.INIT('h8)
	) name286 (
		\TM0_pad ,
		\WX10837_reg/NET0131 ,
		_w1794_
	);
	LUT2 #(
		.INIT('h1)
	) name287 (
		\TM1_pad ,
		\WX653_reg/NET0131 ,
		_w1795_
	);
	LUT2 #(
		.INIT('h8)
	) name288 (
		\TM1_pad ,
		\WX653_reg/NET0131 ,
		_w1796_
	);
	LUT2 #(
		.INIT('h1)
	) name289 (
		_w1795_,
		_w1796_,
		_w1797_
	);
	LUT2 #(
		.INIT('h2)
	) name290 (
		_w1794_,
		_w1797_,
		_w1798_
	);
	LUT2 #(
		.INIT('h4)
	) name291 (
		_w1794_,
		_w1797_,
		_w1799_
	);
	LUT2 #(
		.INIT('h1)
	) name292 (
		_w1798_,
		_w1799_,
		_w1800_
	);
	LUT2 #(
		.INIT('h8)
	) name293 (
		_w1793_,
		_w1800_,
		_w1801_
	);
	LUT2 #(
		.INIT('h1)
	) name294 (
		_w1793_,
		_w1800_,
		_w1802_
	);
	LUT2 #(
		.INIT('h1)
	) name295 (
		_w1801_,
		_w1802_,
		_w1803_
	);
	LUT2 #(
		.INIT('h2)
	) name296 (
		\WX779_reg/NET0131 ,
		\WX843_reg/NET0131 ,
		_w1804_
	);
	LUT2 #(
		.INIT('h4)
	) name297 (
		\WX779_reg/NET0131 ,
		\WX843_reg/NET0131 ,
		_w1805_
	);
	LUT2 #(
		.INIT('h1)
	) name298 (
		_w1804_,
		_w1805_,
		_w1806_
	);
	LUT2 #(
		.INIT('h2)
	) name299 (
		\WX715_reg/NET0131 ,
		_w1806_,
		_w1807_
	);
	LUT2 #(
		.INIT('h4)
	) name300 (
		\WX715_reg/NET0131 ,
		_w1806_,
		_w1808_
	);
	LUT2 #(
		.INIT('h1)
	) name301 (
		_w1807_,
		_w1808_,
		_w1809_
	);
	LUT2 #(
		.INIT('h8)
	) name302 (
		\TM0_pad ,
		\WX10835_reg/NET0131 ,
		_w1810_
	);
	LUT2 #(
		.INIT('h1)
	) name303 (
		\TM1_pad ,
		\WX651_reg/NET0131 ,
		_w1811_
	);
	LUT2 #(
		.INIT('h8)
	) name304 (
		\TM1_pad ,
		\WX651_reg/NET0131 ,
		_w1812_
	);
	LUT2 #(
		.INIT('h1)
	) name305 (
		_w1811_,
		_w1812_,
		_w1813_
	);
	LUT2 #(
		.INIT('h2)
	) name306 (
		_w1810_,
		_w1813_,
		_w1814_
	);
	LUT2 #(
		.INIT('h4)
	) name307 (
		_w1810_,
		_w1813_,
		_w1815_
	);
	LUT2 #(
		.INIT('h1)
	) name308 (
		_w1814_,
		_w1815_,
		_w1816_
	);
	LUT2 #(
		.INIT('h8)
	) name309 (
		_w1809_,
		_w1816_,
		_w1817_
	);
	LUT2 #(
		.INIT('h1)
	) name310 (
		_w1809_,
		_w1816_,
		_w1818_
	);
	LUT2 #(
		.INIT('h1)
	) name311 (
		_w1817_,
		_w1818_,
		_w1819_
	);
	LUT2 #(
		.INIT('h2)
	) name312 (
		\WX777_reg/NET0131 ,
		\WX841_reg/NET0131 ,
		_w1820_
	);
	LUT2 #(
		.INIT('h4)
	) name313 (
		\WX777_reg/NET0131 ,
		\WX841_reg/NET0131 ,
		_w1821_
	);
	LUT2 #(
		.INIT('h1)
	) name314 (
		_w1820_,
		_w1821_,
		_w1822_
	);
	LUT2 #(
		.INIT('h2)
	) name315 (
		\WX713_reg/NET0131 ,
		_w1822_,
		_w1823_
	);
	LUT2 #(
		.INIT('h4)
	) name316 (
		\WX713_reg/NET0131 ,
		_w1822_,
		_w1824_
	);
	LUT2 #(
		.INIT('h1)
	) name317 (
		_w1823_,
		_w1824_,
		_w1825_
	);
	LUT2 #(
		.INIT('h8)
	) name318 (
		\TM0_pad ,
		\WX10833_reg/NET0131 ,
		_w1826_
	);
	LUT2 #(
		.INIT('h1)
	) name319 (
		\TM1_pad ,
		\WX649_reg/NET0131 ,
		_w1827_
	);
	LUT2 #(
		.INIT('h8)
	) name320 (
		\TM1_pad ,
		\WX649_reg/NET0131 ,
		_w1828_
	);
	LUT2 #(
		.INIT('h1)
	) name321 (
		_w1827_,
		_w1828_,
		_w1829_
	);
	LUT2 #(
		.INIT('h2)
	) name322 (
		_w1826_,
		_w1829_,
		_w1830_
	);
	LUT2 #(
		.INIT('h4)
	) name323 (
		_w1826_,
		_w1829_,
		_w1831_
	);
	LUT2 #(
		.INIT('h1)
	) name324 (
		_w1830_,
		_w1831_,
		_w1832_
	);
	LUT2 #(
		.INIT('h8)
	) name325 (
		_w1825_,
		_w1832_,
		_w1833_
	);
	LUT2 #(
		.INIT('h1)
	) name326 (
		_w1825_,
		_w1832_,
		_w1834_
	);
	LUT2 #(
		.INIT('h1)
	) name327 (
		_w1833_,
		_w1834_,
		_w1835_
	);
	LUT2 #(
		.INIT('h2)
	) name328 (
		\TM0_pad ,
		\WX10887_reg/NET0131 ,
		_w1836_
	);
	LUT2 #(
		.INIT('h2)
	) name329 (
		\WX831_reg/NET0131 ,
		\WX895_reg/NET0131 ,
		_w1837_
	);
	LUT2 #(
		.INIT('h4)
	) name330 (
		\WX831_reg/NET0131 ,
		\WX895_reg/NET0131 ,
		_w1838_
	);
	LUT2 #(
		.INIT('h1)
	) name331 (
		_w1837_,
		_w1838_,
		_w1839_
	);
	LUT2 #(
		.INIT('h2)
	) name332 (
		\WX703_reg/NET0131 ,
		\WX767_reg/NET0131 ,
		_w1840_
	);
	LUT2 #(
		.INIT('h4)
	) name333 (
		\WX703_reg/NET0131 ,
		\WX767_reg/NET0131 ,
		_w1841_
	);
	LUT2 #(
		.INIT('h1)
	) name334 (
		_w1840_,
		_w1841_,
		_w1842_
	);
	LUT2 #(
		.INIT('h8)
	) name335 (
		_w1839_,
		_w1842_,
		_w1843_
	);
	LUT2 #(
		.INIT('h1)
	) name336 (
		_w1839_,
		_w1842_,
		_w1844_
	);
	LUT2 #(
		.INIT('h1)
	) name337 (
		_w1843_,
		_w1844_,
		_w1845_
	);
	LUT2 #(
		.INIT('h8)
	) name338 (
		_w1836_,
		_w1845_,
		_w1846_
	);
	LUT2 #(
		.INIT('h1)
	) name339 (
		_w1836_,
		_w1845_,
		_w1847_
	);
	LUT2 #(
		.INIT('h1)
	) name340 (
		_w1846_,
		_w1847_,
		_w1848_
	);
	LUT2 #(
		.INIT('h2)
	) name341 (
		\WX775_reg/NET0131 ,
		\WX839_reg/NET0131 ,
		_w1849_
	);
	LUT2 #(
		.INIT('h4)
	) name342 (
		\WX775_reg/NET0131 ,
		\WX839_reg/NET0131 ,
		_w1850_
	);
	LUT2 #(
		.INIT('h1)
	) name343 (
		_w1849_,
		_w1850_,
		_w1851_
	);
	LUT2 #(
		.INIT('h2)
	) name344 (
		\WX711_reg/NET0131 ,
		_w1851_,
		_w1852_
	);
	LUT2 #(
		.INIT('h4)
	) name345 (
		\WX711_reg/NET0131 ,
		_w1851_,
		_w1853_
	);
	LUT2 #(
		.INIT('h1)
	) name346 (
		_w1852_,
		_w1853_,
		_w1854_
	);
	LUT2 #(
		.INIT('h8)
	) name347 (
		\TM0_pad ,
		\WX10831_reg/NET0131 ,
		_w1855_
	);
	LUT2 #(
		.INIT('h1)
	) name348 (
		\TM1_pad ,
		\WX647_reg/NET0131 ,
		_w1856_
	);
	LUT2 #(
		.INIT('h8)
	) name349 (
		\TM1_pad ,
		\WX647_reg/NET0131 ,
		_w1857_
	);
	LUT2 #(
		.INIT('h1)
	) name350 (
		_w1856_,
		_w1857_,
		_w1858_
	);
	LUT2 #(
		.INIT('h2)
	) name351 (
		_w1855_,
		_w1858_,
		_w1859_
	);
	LUT2 #(
		.INIT('h4)
	) name352 (
		_w1855_,
		_w1858_,
		_w1860_
	);
	LUT2 #(
		.INIT('h1)
	) name353 (
		_w1859_,
		_w1860_,
		_w1861_
	);
	LUT2 #(
		.INIT('h8)
	) name354 (
		_w1854_,
		_w1861_,
		_w1862_
	);
	LUT2 #(
		.INIT('h1)
	) name355 (
		_w1854_,
		_w1861_,
		_w1863_
	);
	LUT2 #(
		.INIT('h1)
	) name356 (
		_w1862_,
		_w1863_,
		_w1864_
	);
	LUT2 #(
		.INIT('h2)
	) name357 (
		\WX773_reg/NET0131 ,
		\WX837_reg/NET0131 ,
		_w1865_
	);
	LUT2 #(
		.INIT('h4)
	) name358 (
		\WX773_reg/NET0131 ,
		\WX837_reg/NET0131 ,
		_w1866_
	);
	LUT2 #(
		.INIT('h1)
	) name359 (
		_w1865_,
		_w1866_,
		_w1867_
	);
	LUT2 #(
		.INIT('h2)
	) name360 (
		\WX709_reg/NET0131 ,
		_w1867_,
		_w1868_
	);
	LUT2 #(
		.INIT('h4)
	) name361 (
		\WX709_reg/NET0131 ,
		_w1867_,
		_w1869_
	);
	LUT2 #(
		.INIT('h1)
	) name362 (
		_w1868_,
		_w1869_,
		_w1870_
	);
	LUT2 #(
		.INIT('h8)
	) name363 (
		\TM0_pad ,
		\WX10829_reg/NET0131 ,
		_w1871_
	);
	LUT2 #(
		.INIT('h1)
	) name364 (
		\TM1_pad ,
		\WX645_reg/NET0131 ,
		_w1872_
	);
	LUT2 #(
		.INIT('h8)
	) name365 (
		\TM1_pad ,
		\WX645_reg/NET0131 ,
		_w1873_
	);
	LUT2 #(
		.INIT('h1)
	) name366 (
		_w1872_,
		_w1873_,
		_w1874_
	);
	LUT2 #(
		.INIT('h2)
	) name367 (
		_w1871_,
		_w1874_,
		_w1875_
	);
	LUT2 #(
		.INIT('h4)
	) name368 (
		_w1871_,
		_w1874_,
		_w1876_
	);
	LUT2 #(
		.INIT('h1)
	) name369 (
		_w1875_,
		_w1876_,
		_w1877_
	);
	LUT2 #(
		.INIT('h8)
	) name370 (
		_w1870_,
		_w1877_,
		_w1878_
	);
	LUT2 #(
		.INIT('h1)
	) name371 (
		_w1870_,
		_w1877_,
		_w1879_
	);
	LUT2 #(
		.INIT('h1)
	) name372 (
		_w1878_,
		_w1879_,
		_w1880_
	);
	LUT2 #(
		.INIT('h2)
	) name373 (
		\TM0_pad ,
		\WX10885_reg/NET0131 ,
		_w1881_
	);
	LUT2 #(
		.INIT('h2)
	) name374 (
		\WX829_reg/NET0131 ,
		\WX893_reg/NET0131 ,
		_w1882_
	);
	LUT2 #(
		.INIT('h4)
	) name375 (
		\WX829_reg/NET0131 ,
		\WX893_reg/NET0131 ,
		_w1883_
	);
	LUT2 #(
		.INIT('h1)
	) name376 (
		_w1882_,
		_w1883_,
		_w1884_
	);
	LUT2 #(
		.INIT('h2)
	) name377 (
		\WX701_reg/NET0131 ,
		\WX765_reg/NET0131 ,
		_w1885_
	);
	LUT2 #(
		.INIT('h4)
	) name378 (
		\WX701_reg/NET0131 ,
		\WX765_reg/NET0131 ,
		_w1886_
	);
	LUT2 #(
		.INIT('h1)
	) name379 (
		_w1885_,
		_w1886_,
		_w1887_
	);
	LUT2 #(
		.INIT('h8)
	) name380 (
		_w1884_,
		_w1887_,
		_w1888_
	);
	LUT2 #(
		.INIT('h1)
	) name381 (
		_w1884_,
		_w1887_,
		_w1889_
	);
	LUT2 #(
		.INIT('h1)
	) name382 (
		_w1888_,
		_w1889_,
		_w1890_
	);
	LUT2 #(
		.INIT('h8)
	) name383 (
		_w1881_,
		_w1890_,
		_w1891_
	);
	LUT2 #(
		.INIT('h1)
	) name384 (
		_w1881_,
		_w1890_,
		_w1892_
	);
	LUT2 #(
		.INIT('h1)
	) name385 (
		_w1891_,
		_w1892_,
		_w1893_
	);
	LUT2 #(
		.INIT('h2)
	) name386 (
		\TM0_pad ,
		\WX10883_reg/NET0131 ,
		_w1894_
	);
	LUT2 #(
		.INIT('h2)
	) name387 (
		\WX827_reg/NET0131 ,
		\WX891_reg/NET0131 ,
		_w1895_
	);
	LUT2 #(
		.INIT('h4)
	) name388 (
		\WX827_reg/NET0131 ,
		\WX891_reg/NET0131 ,
		_w1896_
	);
	LUT2 #(
		.INIT('h1)
	) name389 (
		_w1895_,
		_w1896_,
		_w1897_
	);
	LUT2 #(
		.INIT('h2)
	) name390 (
		\WX699_reg/NET0131 ,
		\WX763_reg/NET0131 ,
		_w1898_
	);
	LUT2 #(
		.INIT('h4)
	) name391 (
		\WX699_reg/NET0131 ,
		\WX763_reg/NET0131 ,
		_w1899_
	);
	LUT2 #(
		.INIT('h1)
	) name392 (
		_w1898_,
		_w1899_,
		_w1900_
	);
	LUT2 #(
		.INIT('h8)
	) name393 (
		_w1897_,
		_w1900_,
		_w1901_
	);
	LUT2 #(
		.INIT('h1)
	) name394 (
		_w1897_,
		_w1900_,
		_w1902_
	);
	LUT2 #(
		.INIT('h1)
	) name395 (
		_w1901_,
		_w1902_,
		_w1903_
	);
	LUT2 #(
		.INIT('h8)
	) name396 (
		_w1894_,
		_w1903_,
		_w1904_
	);
	LUT2 #(
		.INIT('h1)
	) name397 (
		_w1894_,
		_w1903_,
		_w1905_
	);
	LUT2 #(
		.INIT('h1)
	) name398 (
		_w1904_,
		_w1905_,
		_w1906_
	);
	LUT2 #(
		.INIT('h2)
	) name399 (
		\TM0_pad ,
		\WX10881_reg/NET0131 ,
		_w1907_
	);
	LUT2 #(
		.INIT('h2)
	) name400 (
		\WX825_reg/NET0131 ,
		\WX889_reg/NET0131 ,
		_w1908_
	);
	LUT2 #(
		.INIT('h4)
	) name401 (
		\WX825_reg/NET0131 ,
		\WX889_reg/NET0131 ,
		_w1909_
	);
	LUT2 #(
		.INIT('h1)
	) name402 (
		_w1908_,
		_w1909_,
		_w1910_
	);
	LUT2 #(
		.INIT('h2)
	) name403 (
		\WX697_reg/NET0131 ,
		\WX761_reg/NET0131 ,
		_w1911_
	);
	LUT2 #(
		.INIT('h4)
	) name404 (
		\WX697_reg/NET0131 ,
		\WX761_reg/NET0131 ,
		_w1912_
	);
	LUT2 #(
		.INIT('h1)
	) name405 (
		_w1911_,
		_w1912_,
		_w1913_
	);
	LUT2 #(
		.INIT('h8)
	) name406 (
		_w1910_,
		_w1913_,
		_w1914_
	);
	LUT2 #(
		.INIT('h1)
	) name407 (
		_w1910_,
		_w1913_,
		_w1915_
	);
	LUT2 #(
		.INIT('h1)
	) name408 (
		_w1914_,
		_w1915_,
		_w1916_
	);
	LUT2 #(
		.INIT('h8)
	) name409 (
		_w1907_,
		_w1916_,
		_w1917_
	);
	LUT2 #(
		.INIT('h1)
	) name410 (
		_w1907_,
		_w1916_,
		_w1918_
	);
	LUT2 #(
		.INIT('h1)
	) name411 (
		_w1917_,
		_w1918_,
		_w1919_
	);
	LUT2 #(
		.INIT('h2)
	) name412 (
		\TM0_pad ,
		\WX10879_reg/NET0131 ,
		_w1920_
	);
	LUT2 #(
		.INIT('h2)
	) name413 (
		\WX823_reg/NET0131 ,
		\WX887_reg/NET0131 ,
		_w1921_
	);
	LUT2 #(
		.INIT('h4)
	) name414 (
		\WX823_reg/NET0131 ,
		\WX887_reg/NET0131 ,
		_w1922_
	);
	LUT2 #(
		.INIT('h1)
	) name415 (
		_w1921_,
		_w1922_,
		_w1923_
	);
	LUT2 #(
		.INIT('h2)
	) name416 (
		\WX695_reg/NET0131 ,
		\WX759_reg/NET0131 ,
		_w1924_
	);
	LUT2 #(
		.INIT('h4)
	) name417 (
		\WX695_reg/NET0131 ,
		\WX759_reg/NET0131 ,
		_w1925_
	);
	LUT2 #(
		.INIT('h1)
	) name418 (
		_w1924_,
		_w1925_,
		_w1926_
	);
	LUT2 #(
		.INIT('h8)
	) name419 (
		_w1923_,
		_w1926_,
		_w1927_
	);
	LUT2 #(
		.INIT('h1)
	) name420 (
		_w1923_,
		_w1926_,
		_w1928_
	);
	LUT2 #(
		.INIT('h1)
	) name421 (
		_w1927_,
		_w1928_,
		_w1929_
	);
	LUT2 #(
		.INIT('h8)
	) name422 (
		_w1920_,
		_w1929_,
		_w1930_
	);
	LUT2 #(
		.INIT('h1)
	) name423 (
		_w1920_,
		_w1929_,
		_w1931_
	);
	LUT2 #(
		.INIT('h1)
	) name424 (
		_w1930_,
		_w1931_,
		_w1932_
	);
	LUT2 #(
		.INIT('h2)
	) name425 (
		\TM0_pad ,
		\WX10877_reg/NET0131 ,
		_w1933_
	);
	LUT2 #(
		.INIT('h2)
	) name426 (
		\WX821_reg/NET0131 ,
		\WX885_reg/NET0131 ,
		_w1934_
	);
	LUT2 #(
		.INIT('h4)
	) name427 (
		\WX821_reg/NET0131 ,
		\WX885_reg/NET0131 ,
		_w1935_
	);
	LUT2 #(
		.INIT('h1)
	) name428 (
		_w1934_,
		_w1935_,
		_w1936_
	);
	LUT2 #(
		.INIT('h2)
	) name429 (
		\WX693_reg/NET0131 ,
		\WX757_reg/NET0131 ,
		_w1937_
	);
	LUT2 #(
		.INIT('h4)
	) name430 (
		\WX693_reg/NET0131 ,
		\WX757_reg/NET0131 ,
		_w1938_
	);
	LUT2 #(
		.INIT('h1)
	) name431 (
		_w1937_,
		_w1938_,
		_w1939_
	);
	LUT2 #(
		.INIT('h8)
	) name432 (
		_w1936_,
		_w1939_,
		_w1940_
	);
	LUT2 #(
		.INIT('h1)
	) name433 (
		_w1936_,
		_w1939_,
		_w1941_
	);
	LUT2 #(
		.INIT('h1)
	) name434 (
		_w1940_,
		_w1941_,
		_w1942_
	);
	LUT2 #(
		.INIT('h8)
	) name435 (
		_w1933_,
		_w1942_,
		_w1943_
	);
	LUT2 #(
		.INIT('h1)
	) name436 (
		_w1933_,
		_w1942_,
		_w1944_
	);
	LUT2 #(
		.INIT('h1)
	) name437 (
		_w1943_,
		_w1944_,
		_w1945_
	);
	LUT2 #(
		.INIT('h2)
	) name438 (
		\TM0_pad ,
		\WX10875_reg/NET0131 ,
		_w1946_
	);
	LUT2 #(
		.INIT('h2)
	) name439 (
		\WX819_reg/NET0131 ,
		\WX883_reg/NET0131 ,
		_w1947_
	);
	LUT2 #(
		.INIT('h4)
	) name440 (
		\WX819_reg/NET0131 ,
		\WX883_reg/NET0131 ,
		_w1948_
	);
	LUT2 #(
		.INIT('h1)
	) name441 (
		_w1947_,
		_w1948_,
		_w1949_
	);
	LUT2 #(
		.INIT('h2)
	) name442 (
		\WX691_reg/NET0131 ,
		\WX755_reg/NET0131 ,
		_w1950_
	);
	LUT2 #(
		.INIT('h4)
	) name443 (
		\WX691_reg/NET0131 ,
		\WX755_reg/NET0131 ,
		_w1951_
	);
	LUT2 #(
		.INIT('h1)
	) name444 (
		_w1950_,
		_w1951_,
		_w1952_
	);
	LUT2 #(
		.INIT('h8)
	) name445 (
		_w1949_,
		_w1952_,
		_w1953_
	);
	LUT2 #(
		.INIT('h1)
	) name446 (
		_w1949_,
		_w1952_,
		_w1954_
	);
	LUT2 #(
		.INIT('h1)
	) name447 (
		_w1953_,
		_w1954_,
		_w1955_
	);
	LUT2 #(
		.INIT('h8)
	) name448 (
		_w1946_,
		_w1955_,
		_w1956_
	);
	LUT2 #(
		.INIT('h1)
	) name449 (
		_w1946_,
		_w1955_,
		_w1957_
	);
	LUT2 #(
		.INIT('h1)
	) name450 (
		_w1956_,
		_w1957_,
		_w1958_
	);
	LUT2 #(
		.INIT('h2)
	) name451 (
		\TM0_pad ,
		\WX10873_reg/NET0131 ,
		_w1959_
	);
	LUT2 #(
		.INIT('h2)
	) name452 (
		\WX817_reg/NET0131 ,
		\WX881_reg/NET0131 ,
		_w1960_
	);
	LUT2 #(
		.INIT('h4)
	) name453 (
		\WX817_reg/NET0131 ,
		\WX881_reg/NET0131 ,
		_w1961_
	);
	LUT2 #(
		.INIT('h1)
	) name454 (
		_w1960_,
		_w1961_,
		_w1962_
	);
	LUT2 #(
		.INIT('h2)
	) name455 (
		\WX689_reg/NET0131 ,
		\WX753_reg/NET0131 ,
		_w1963_
	);
	LUT2 #(
		.INIT('h4)
	) name456 (
		\WX689_reg/NET0131 ,
		\WX753_reg/NET0131 ,
		_w1964_
	);
	LUT2 #(
		.INIT('h1)
	) name457 (
		_w1963_,
		_w1964_,
		_w1965_
	);
	LUT2 #(
		.INIT('h8)
	) name458 (
		_w1962_,
		_w1965_,
		_w1966_
	);
	LUT2 #(
		.INIT('h1)
	) name459 (
		_w1962_,
		_w1965_,
		_w1967_
	);
	LUT2 #(
		.INIT('h1)
	) name460 (
		_w1966_,
		_w1967_,
		_w1968_
	);
	LUT2 #(
		.INIT('h8)
	) name461 (
		_w1959_,
		_w1968_,
		_w1969_
	);
	LUT2 #(
		.INIT('h1)
	) name462 (
		_w1959_,
		_w1968_,
		_w1970_
	);
	LUT2 #(
		.INIT('h1)
	) name463 (
		_w1969_,
		_w1970_,
		_w1971_
	);
	LUT2 #(
		.INIT('h1)
	) name464 (
		\TM0_pad ,
		_w1595_,
		_w1972_
	);
	LUT2 #(
		.INIT('h8)
	) name465 (
		RESET_pad,
		\TM1_pad ,
		_w1973_
	);
	LUT2 #(
		.INIT('h4)
	) name466 (
		_w1586_,
		_w1973_,
		_w1974_
	);
	LUT2 #(
		.INIT('h4)
	) name467 (
		_w1972_,
		_w1974_,
		_w1975_
	);
	LUT2 #(
		.INIT('h2)
	) name468 (
		RESET_pad,
		\TM1_pad ,
		_w1976_
	);
	LUT2 #(
		.INIT('h2)
	) name469 (
		\TM0_pad ,
		\_2092__reg/NET0131 ,
		_w1977_
	);
	LUT2 #(
		.INIT('h2)
	) name470 (
		\WX2098_reg/NET0131 ,
		\WX2162_reg/NET0131 ,
		_w1978_
	);
	LUT2 #(
		.INIT('h4)
	) name471 (
		\WX2098_reg/NET0131 ,
		\WX2162_reg/NET0131 ,
		_w1979_
	);
	LUT2 #(
		.INIT('h1)
	) name472 (
		_w1978_,
		_w1979_,
		_w1980_
	);
	LUT2 #(
		.INIT('h2)
	) name473 (
		\WX1970_reg/NET0131 ,
		\WX2034_reg/NET0131 ,
		_w1981_
	);
	LUT2 #(
		.INIT('h4)
	) name474 (
		\WX1970_reg/NET0131 ,
		\WX2034_reg/NET0131 ,
		_w1982_
	);
	LUT2 #(
		.INIT('h1)
	) name475 (
		_w1981_,
		_w1982_,
		_w1983_
	);
	LUT2 #(
		.INIT('h4)
	) name476 (
		_w1980_,
		_w1983_,
		_w1984_
	);
	LUT2 #(
		.INIT('h2)
	) name477 (
		_w1980_,
		_w1983_,
		_w1985_
	);
	LUT2 #(
		.INIT('h1)
	) name478 (
		\TM0_pad ,
		_w1984_,
		_w1986_
	);
	LUT2 #(
		.INIT('h4)
	) name479 (
		_w1985_,
		_w1986_,
		_w1987_
	);
	LUT2 #(
		.INIT('h2)
	) name480 (
		_w1976_,
		_w1977_,
		_w1988_
	);
	LUT2 #(
		.INIT('h4)
	) name481 (
		_w1987_,
		_w1988_,
		_w1989_
	);
	LUT2 #(
		.INIT('h1)
	) name482 (
		_w1975_,
		_w1989_,
		_w1990_
	);
	LUT2 #(
		.INIT('h2)
	) name483 (
		\WX9830_reg/NET0131 ,
		\WX9894_reg/NET0131 ,
		_w1991_
	);
	LUT2 #(
		.INIT('h4)
	) name484 (
		\WX9830_reg/NET0131 ,
		\WX9894_reg/NET0131 ,
		_w1992_
	);
	LUT2 #(
		.INIT('h1)
	) name485 (
		_w1991_,
		_w1992_,
		_w1993_
	);
	LUT2 #(
		.INIT('h2)
	) name486 (
		\WX9766_reg/NET0131 ,
		_w1993_,
		_w1994_
	);
	LUT2 #(
		.INIT('h4)
	) name487 (
		\WX9766_reg/NET0131 ,
		_w1993_,
		_w1995_
	);
	LUT2 #(
		.INIT('h1)
	) name488 (
		_w1994_,
		_w1995_,
		_w1996_
	);
	LUT2 #(
		.INIT('h2)
	) name489 (
		\TM1_pad ,
		\WX9702_reg/NET0131 ,
		_w1997_
	);
	LUT2 #(
		.INIT('h4)
	) name490 (
		\TM1_pad ,
		\WX9702_reg/NET0131 ,
		_w1998_
	);
	LUT2 #(
		.INIT('h1)
	) name491 (
		_w1997_,
		_w1998_,
		_w1999_
	);
	LUT2 #(
		.INIT('h4)
	) name492 (
		_w1996_,
		_w1999_,
		_w2000_
	);
	LUT2 #(
		.INIT('h2)
	) name493 (
		_w1996_,
		_w1999_,
		_w2001_
	);
	LUT2 #(
		.INIT('h1)
	) name494 (
		\TM0_pad ,
		_w2000_,
		_w2002_
	);
	LUT2 #(
		.INIT('h4)
	) name495 (
		_w2001_,
		_w2002_,
		_w2003_
	);
	LUT2 #(
		.INIT('h1)
	) name496 (
		_w1810_,
		_w2003_,
		_w2004_
	);
	LUT2 #(
		.INIT('h2)
	) name497 (
		_w1973_,
		_w2004_,
		_w2005_
	);
	LUT2 #(
		.INIT('h8)
	) name498 (
		\TM0_pad ,
		\_2329__reg/NET0131 ,
		_w2006_
	);
	LUT2 #(
		.INIT('h2)
	) name499 (
		\WX11123_reg/NET0131 ,
		\WX11187_reg/NET0131 ,
		_w2007_
	);
	LUT2 #(
		.INIT('h4)
	) name500 (
		\WX11123_reg/NET0131 ,
		\WX11187_reg/NET0131 ,
		_w2008_
	);
	LUT2 #(
		.INIT('h1)
	) name501 (
		_w2007_,
		_w2008_,
		_w2009_
	);
	LUT2 #(
		.INIT('h2)
	) name502 (
		\WX11059_reg/NET0131 ,
		_w2009_,
		_w2010_
	);
	LUT2 #(
		.INIT('h4)
	) name503 (
		\WX11059_reg/NET0131 ,
		_w2009_,
		_w2011_
	);
	LUT2 #(
		.INIT('h1)
	) name504 (
		_w2010_,
		_w2011_,
		_w2012_
	);
	LUT2 #(
		.INIT('h2)
	) name505 (
		\TM1_pad ,
		\WX10995_reg/NET0131 ,
		_w2013_
	);
	LUT2 #(
		.INIT('h4)
	) name506 (
		\TM1_pad ,
		\WX10995_reg/NET0131 ,
		_w2014_
	);
	LUT2 #(
		.INIT('h1)
	) name507 (
		_w2013_,
		_w2014_,
		_w2015_
	);
	LUT2 #(
		.INIT('h4)
	) name508 (
		_w2012_,
		_w2015_,
		_w2016_
	);
	LUT2 #(
		.INIT('h2)
	) name509 (
		_w2012_,
		_w2015_,
		_w2017_
	);
	LUT2 #(
		.INIT('h1)
	) name510 (
		\TM0_pad ,
		_w2016_,
		_w2018_
	);
	LUT2 #(
		.INIT('h4)
	) name511 (
		_w2017_,
		_w2018_,
		_w2019_
	);
	LUT2 #(
		.INIT('h1)
	) name512 (
		_w2006_,
		_w2019_,
		_w2020_
	);
	LUT2 #(
		.INIT('h2)
	) name513 (
		_w1976_,
		_w2020_,
		_w2021_
	);
	LUT2 #(
		.INIT('h1)
	) name514 (
		_w2005_,
		_w2021_,
		_w2022_
	);
	LUT2 #(
		.INIT('h4)
	) name515 (
		_w1946_,
		_w1973_,
		_w2023_
	);
	LUT2 #(
		.INIT('h2)
	) name516 (
		\WX11163_reg/NET0131 ,
		\WX11227_reg/NET0131 ,
		_w2024_
	);
	LUT2 #(
		.INIT('h4)
	) name517 (
		\WX11163_reg/NET0131 ,
		\WX11227_reg/NET0131 ,
		_w2025_
	);
	LUT2 #(
		.INIT('h1)
	) name518 (
		_w2024_,
		_w2025_,
		_w2026_
	);
	LUT2 #(
		.INIT('h2)
	) name519 (
		\WX11035_reg/NET0131 ,
		\WX11099_reg/NET0131 ,
		_w2027_
	);
	LUT2 #(
		.INIT('h4)
	) name520 (
		\WX11035_reg/NET0131 ,
		\WX11099_reg/NET0131 ,
		_w2028_
	);
	LUT2 #(
		.INIT('h1)
	) name521 (
		_w2027_,
		_w2028_,
		_w2029_
	);
	LUT2 #(
		.INIT('h4)
	) name522 (
		_w2026_,
		_w2029_,
		_w2030_
	);
	LUT2 #(
		.INIT('h2)
	) name523 (
		_w2026_,
		_w2029_,
		_w2031_
	);
	LUT2 #(
		.INIT('h1)
	) name524 (
		\TM0_pad ,
		_w2030_,
		_w2032_
	);
	LUT2 #(
		.INIT('h4)
	) name525 (
		_w2031_,
		_w2032_,
		_w2033_
	);
	LUT2 #(
		.INIT('h2)
	) name526 (
		_w2023_,
		_w2033_,
		_w2034_
	);
	LUT2 #(
		.INIT('h1)
	) name527 (
		\DATA_0_8_pad ,
		\TM0_pad ,
		_w2035_
	);
	LUT2 #(
		.INIT('h2)
	) name528 (
		\TM0_pad ,
		\_2341__reg/NET0131 ,
		_w2036_
	);
	LUT2 #(
		.INIT('h2)
	) name529 (
		_w1976_,
		_w2035_,
		_w2037_
	);
	LUT2 #(
		.INIT('h4)
	) name530 (
		_w2036_,
		_w2037_,
		_w2038_
	);
	LUT2 #(
		.INIT('h1)
	) name531 (
		_w2034_,
		_w2038_,
		_w2039_
	);
	LUT2 #(
		.INIT('h4)
	) name532 (
		_w1560_,
		_w1973_,
		_w2040_
	);
	LUT2 #(
		.INIT('h2)
	) name533 (
		\WX11153_reg/NET0131 ,
		\WX11217_reg/NET0131 ,
		_w2041_
	);
	LUT2 #(
		.INIT('h4)
	) name534 (
		\WX11153_reg/NET0131 ,
		\WX11217_reg/NET0131 ,
		_w2042_
	);
	LUT2 #(
		.INIT('h1)
	) name535 (
		_w2041_,
		_w2042_,
		_w2043_
	);
	LUT2 #(
		.INIT('h2)
	) name536 (
		\WX11025_reg/NET0131 ,
		\WX11089_reg/NET0131 ,
		_w2044_
	);
	LUT2 #(
		.INIT('h4)
	) name537 (
		\WX11025_reg/NET0131 ,
		\WX11089_reg/NET0131 ,
		_w2045_
	);
	LUT2 #(
		.INIT('h1)
	) name538 (
		_w2044_,
		_w2045_,
		_w2046_
	);
	LUT2 #(
		.INIT('h4)
	) name539 (
		_w2043_,
		_w2046_,
		_w2047_
	);
	LUT2 #(
		.INIT('h2)
	) name540 (
		_w2043_,
		_w2046_,
		_w2048_
	);
	LUT2 #(
		.INIT('h1)
	) name541 (
		\TM0_pad ,
		_w2047_,
		_w2049_
	);
	LUT2 #(
		.INIT('h4)
	) name542 (
		_w2048_,
		_w2049_,
		_w2050_
	);
	LUT2 #(
		.INIT('h2)
	) name543 (
		_w2040_,
		_w2050_,
		_w2051_
	);
	LUT2 #(
		.INIT('h1)
	) name544 (
		\DATA_0_13_pad ,
		\TM0_pad ,
		_w2052_
	);
	LUT2 #(
		.INIT('h2)
	) name545 (
		\TM0_pad ,
		\_2346__reg/NET0131 ,
		_w2053_
	);
	LUT2 #(
		.INIT('h2)
	) name546 (
		_w1976_,
		_w2052_,
		_w2054_
	);
	LUT2 #(
		.INIT('h4)
	) name547 (
		_w2053_,
		_w2054_,
		_w2055_
	);
	LUT2 #(
		.INIT('h1)
	) name548 (
		_w2051_,
		_w2055_,
		_w2056_
	);
	LUT2 #(
		.INIT('h1)
	) name549 (
		\TM0_pad ,
		_w1864_,
		_w2057_
	);
	LUT2 #(
		.INIT('h1)
	) name550 (
		_w1855_,
		_w2057_,
		_w2058_
	);
	LUT2 #(
		.INIT('h2)
	) name551 (
		_w1973_,
		_w2058_,
		_w2059_
	);
	LUT2 #(
		.INIT('h8)
	) name552 (
		\TM0_pad ,
		\_2107__reg/NET0131 ,
		_w2060_
	);
	LUT2 #(
		.INIT('h2)
	) name553 (
		\WX2068_reg/NET0131 ,
		\WX2132_reg/NET0131 ,
		_w2061_
	);
	LUT2 #(
		.INIT('h4)
	) name554 (
		\WX2068_reg/NET0131 ,
		\WX2132_reg/NET0131 ,
		_w2062_
	);
	LUT2 #(
		.INIT('h1)
	) name555 (
		_w2061_,
		_w2062_,
		_w2063_
	);
	LUT2 #(
		.INIT('h2)
	) name556 (
		\WX2004_reg/NET0131 ,
		_w2063_,
		_w2064_
	);
	LUT2 #(
		.INIT('h4)
	) name557 (
		\WX2004_reg/NET0131 ,
		_w2063_,
		_w2065_
	);
	LUT2 #(
		.INIT('h1)
	) name558 (
		_w2064_,
		_w2065_,
		_w2066_
	);
	LUT2 #(
		.INIT('h2)
	) name559 (
		\TM1_pad ,
		\WX1940_reg/NET0131 ,
		_w2067_
	);
	LUT2 #(
		.INIT('h4)
	) name560 (
		\TM1_pad ,
		\WX1940_reg/NET0131 ,
		_w2068_
	);
	LUT2 #(
		.INIT('h1)
	) name561 (
		_w2067_,
		_w2068_,
		_w2069_
	);
	LUT2 #(
		.INIT('h4)
	) name562 (
		_w2066_,
		_w2069_,
		_w2070_
	);
	LUT2 #(
		.INIT('h2)
	) name563 (
		_w2066_,
		_w2069_,
		_w2071_
	);
	LUT2 #(
		.INIT('h1)
	) name564 (
		\TM0_pad ,
		_w2070_,
		_w2072_
	);
	LUT2 #(
		.INIT('h4)
	) name565 (
		_w2071_,
		_w2072_,
		_w2073_
	);
	LUT2 #(
		.INIT('h1)
	) name566 (
		_w2060_,
		_w2073_,
		_w2074_
	);
	LUT2 #(
		.INIT('h2)
	) name567 (
		_w1976_,
		_w2074_,
		_w2075_
	);
	LUT2 #(
		.INIT('h1)
	) name568 (
		_w2059_,
		_w2075_,
		_w2076_
	);
	LUT2 #(
		.INIT('h1)
	) name569 (
		\TM0_pad ,
		_w1835_,
		_w2077_
	);
	LUT2 #(
		.INIT('h1)
	) name570 (
		_w1826_,
		_w2077_,
		_w2078_
	);
	LUT2 #(
		.INIT('h2)
	) name571 (
		_w1973_,
		_w2078_,
		_w2079_
	);
	LUT2 #(
		.INIT('h8)
	) name572 (
		\TM0_pad ,
		\_2106__reg/NET0131 ,
		_w2080_
	);
	LUT2 #(
		.INIT('h2)
	) name573 (
		\WX2070_reg/NET0131 ,
		\WX2134_reg/NET0131 ,
		_w2081_
	);
	LUT2 #(
		.INIT('h4)
	) name574 (
		\WX2070_reg/NET0131 ,
		\WX2134_reg/NET0131 ,
		_w2082_
	);
	LUT2 #(
		.INIT('h1)
	) name575 (
		_w2081_,
		_w2082_,
		_w2083_
	);
	LUT2 #(
		.INIT('h2)
	) name576 (
		\WX2006_reg/NET0131 ,
		_w2083_,
		_w2084_
	);
	LUT2 #(
		.INIT('h4)
	) name577 (
		\WX2006_reg/NET0131 ,
		_w2083_,
		_w2085_
	);
	LUT2 #(
		.INIT('h1)
	) name578 (
		_w2084_,
		_w2085_,
		_w2086_
	);
	LUT2 #(
		.INIT('h2)
	) name579 (
		\TM1_pad ,
		\WX1942_reg/NET0131 ,
		_w2087_
	);
	LUT2 #(
		.INIT('h4)
	) name580 (
		\TM1_pad ,
		\WX1942_reg/NET0131 ,
		_w2088_
	);
	LUT2 #(
		.INIT('h1)
	) name581 (
		_w2087_,
		_w2088_,
		_w2089_
	);
	LUT2 #(
		.INIT('h4)
	) name582 (
		_w2086_,
		_w2089_,
		_w2090_
	);
	LUT2 #(
		.INIT('h2)
	) name583 (
		_w2086_,
		_w2089_,
		_w2091_
	);
	LUT2 #(
		.INIT('h1)
	) name584 (
		\TM0_pad ,
		_w2090_,
		_w2092_
	);
	LUT2 #(
		.INIT('h4)
	) name585 (
		_w2091_,
		_w2092_,
		_w2093_
	);
	LUT2 #(
		.INIT('h1)
	) name586 (
		_w2080_,
		_w2093_,
		_w2094_
	);
	LUT2 #(
		.INIT('h2)
	) name587 (
		_w1976_,
		_w2094_,
		_w2095_
	);
	LUT2 #(
		.INIT('h1)
	) name588 (
		_w2079_,
		_w2095_,
		_w2096_
	);
	LUT2 #(
		.INIT('h2)
	) name589 (
		\WX3391_reg/NET0131 ,
		\WX3455_reg/NET0131 ,
		_w2097_
	);
	LUT2 #(
		.INIT('h4)
	) name590 (
		\WX3391_reg/NET0131 ,
		\WX3455_reg/NET0131 ,
		_w2098_
	);
	LUT2 #(
		.INIT('h1)
	) name591 (
		_w2097_,
		_w2098_,
		_w2099_
	);
	LUT2 #(
		.INIT('h2)
	) name592 (
		\WX3263_reg/NET0131 ,
		\WX3327_reg/NET0131 ,
		_w2100_
	);
	LUT2 #(
		.INIT('h4)
	) name593 (
		\WX3263_reg/NET0131 ,
		\WX3327_reg/NET0131 ,
		_w2101_
	);
	LUT2 #(
		.INIT('h1)
	) name594 (
		_w2100_,
		_w2101_,
		_w2102_
	);
	LUT2 #(
		.INIT('h4)
	) name595 (
		_w2099_,
		_w2102_,
		_w2103_
	);
	LUT2 #(
		.INIT('h2)
	) name596 (
		_w2099_,
		_w2102_,
		_w2104_
	);
	LUT2 #(
		.INIT('h1)
	) name597 (
		\TM0_pad ,
		_w2103_,
		_w2105_
	);
	LUT2 #(
		.INIT('h4)
	) name598 (
		_w2104_,
		_w2105_,
		_w2106_
	);
	LUT2 #(
		.INIT('h2)
	) name599 (
		_w1974_,
		_w2106_,
		_w2107_
	);
	LUT2 #(
		.INIT('h2)
	) name600 (
		\TM0_pad ,
		\_2156__reg/NET0131 ,
		_w2108_
	);
	LUT2 #(
		.INIT('h2)
	) name601 (
		\WX4684_reg/NET0131 ,
		\WX4748_reg/NET0131 ,
		_w2109_
	);
	LUT2 #(
		.INIT('h4)
	) name602 (
		\WX4684_reg/NET0131 ,
		\WX4748_reg/NET0131 ,
		_w2110_
	);
	LUT2 #(
		.INIT('h1)
	) name603 (
		_w2109_,
		_w2110_,
		_w2111_
	);
	LUT2 #(
		.INIT('h2)
	) name604 (
		\WX4556_reg/NET0131 ,
		\WX4620_reg/NET0131 ,
		_w2112_
	);
	LUT2 #(
		.INIT('h4)
	) name605 (
		\WX4556_reg/NET0131 ,
		\WX4620_reg/NET0131 ,
		_w2113_
	);
	LUT2 #(
		.INIT('h1)
	) name606 (
		_w2112_,
		_w2113_,
		_w2114_
	);
	LUT2 #(
		.INIT('h4)
	) name607 (
		_w2111_,
		_w2114_,
		_w2115_
	);
	LUT2 #(
		.INIT('h2)
	) name608 (
		_w2111_,
		_w2114_,
		_w2116_
	);
	LUT2 #(
		.INIT('h1)
	) name609 (
		\TM0_pad ,
		_w2115_,
		_w2117_
	);
	LUT2 #(
		.INIT('h4)
	) name610 (
		_w2116_,
		_w2117_,
		_w2118_
	);
	LUT2 #(
		.INIT('h2)
	) name611 (
		_w1976_,
		_w2108_,
		_w2119_
	);
	LUT2 #(
		.INIT('h4)
	) name612 (
		_w2118_,
		_w2119_,
		_w2120_
	);
	LUT2 #(
		.INIT('h1)
	) name613 (
		_w2107_,
		_w2120_,
		_w2121_
	);
	LUT2 #(
		.INIT('h8)
	) name614 (
		\TM0_pad ,
		\_2139__reg/NET0131 ,
		_w2122_
	);
	LUT2 #(
		.INIT('h2)
	) name615 (
		\WX3361_reg/NET0131 ,
		\WX3425_reg/NET0131 ,
		_w2123_
	);
	LUT2 #(
		.INIT('h4)
	) name616 (
		\WX3361_reg/NET0131 ,
		\WX3425_reg/NET0131 ,
		_w2124_
	);
	LUT2 #(
		.INIT('h1)
	) name617 (
		_w2123_,
		_w2124_,
		_w2125_
	);
	LUT2 #(
		.INIT('h2)
	) name618 (
		\WX3297_reg/NET0131 ,
		_w2125_,
		_w2126_
	);
	LUT2 #(
		.INIT('h4)
	) name619 (
		\WX3297_reg/NET0131 ,
		_w2125_,
		_w2127_
	);
	LUT2 #(
		.INIT('h1)
	) name620 (
		_w2126_,
		_w2127_,
		_w2128_
	);
	LUT2 #(
		.INIT('h2)
	) name621 (
		\TM1_pad ,
		\WX3233_reg/NET0131 ,
		_w2129_
	);
	LUT2 #(
		.INIT('h4)
	) name622 (
		\TM1_pad ,
		\WX3233_reg/NET0131 ,
		_w2130_
	);
	LUT2 #(
		.INIT('h1)
	) name623 (
		_w2129_,
		_w2130_,
		_w2131_
	);
	LUT2 #(
		.INIT('h4)
	) name624 (
		_w2128_,
		_w2131_,
		_w2132_
	);
	LUT2 #(
		.INIT('h2)
	) name625 (
		_w2128_,
		_w2131_,
		_w2133_
	);
	LUT2 #(
		.INIT('h1)
	) name626 (
		\TM0_pad ,
		_w2132_,
		_w2134_
	);
	LUT2 #(
		.INIT('h4)
	) name627 (
		_w2133_,
		_w2134_,
		_w2135_
	);
	LUT2 #(
		.INIT('h1)
	) name628 (
		_w2122_,
		_w2135_,
		_w2136_
	);
	LUT2 #(
		.INIT('h2)
	) name629 (
		_w1976_,
		_w2136_,
		_w2137_
	);
	LUT2 #(
		.INIT('h1)
	) name630 (
		_w1855_,
		_w2073_,
		_w2138_
	);
	LUT2 #(
		.INIT('h2)
	) name631 (
		_w1973_,
		_w2138_,
		_w2139_
	);
	LUT2 #(
		.INIT('h1)
	) name632 (
		_w2137_,
		_w2139_,
		_w2140_
	);
	LUT2 #(
		.INIT('h8)
	) name633 (
		\TM0_pad ,
		\_2288__reg/NET0131 ,
		_w2141_
	);
	LUT2 #(
		.INIT('h2)
	) name634 (
		\WX9848_reg/NET0131 ,
		\WX9912_reg/NET0131 ,
		_w2142_
	);
	LUT2 #(
		.INIT('h4)
	) name635 (
		\WX9848_reg/NET0131 ,
		\WX9912_reg/NET0131 ,
		_w2143_
	);
	LUT2 #(
		.INIT('h1)
	) name636 (
		_w2142_,
		_w2143_,
		_w2144_
	);
	LUT2 #(
		.INIT('h2)
	) name637 (
		\WX9784_reg/NET0131 ,
		_w2144_,
		_w2145_
	);
	LUT2 #(
		.INIT('h4)
	) name638 (
		\WX9784_reg/NET0131 ,
		_w2144_,
		_w2146_
	);
	LUT2 #(
		.INIT('h1)
	) name639 (
		_w2145_,
		_w2146_,
		_w2147_
	);
	LUT2 #(
		.INIT('h2)
	) name640 (
		\TM1_pad ,
		\WX9720_reg/NET0131 ,
		_w2148_
	);
	LUT2 #(
		.INIT('h4)
	) name641 (
		\TM1_pad ,
		\WX9720_reg/NET0131 ,
		_w2149_
	);
	LUT2 #(
		.INIT('h1)
	) name642 (
		_w2148_,
		_w2149_,
		_w2150_
	);
	LUT2 #(
		.INIT('h4)
	) name643 (
		_w2147_,
		_w2150_,
		_w2151_
	);
	LUT2 #(
		.INIT('h2)
	) name644 (
		_w2147_,
		_w2150_,
		_w2152_
	);
	LUT2 #(
		.INIT('h1)
	) name645 (
		\TM0_pad ,
		_w2151_,
		_w2153_
	);
	LUT2 #(
		.INIT('h4)
	) name646 (
		_w2152_,
		_w2153_,
		_w2154_
	);
	LUT2 #(
		.INIT('h1)
	) name647 (
		_w2141_,
		_w2154_,
		_w2155_
	);
	LUT2 #(
		.INIT('h2)
	) name648 (
		_w1976_,
		_w2155_,
		_w2156_
	);
	LUT2 #(
		.INIT('h2)
	) name649 (
		\WX8555_reg/NET0131 ,
		\WX8619_reg/NET0131 ,
		_w2157_
	);
	LUT2 #(
		.INIT('h4)
	) name650 (
		\WX8555_reg/NET0131 ,
		\WX8619_reg/NET0131 ,
		_w2158_
	);
	LUT2 #(
		.INIT('h1)
	) name651 (
		_w2157_,
		_w2158_,
		_w2159_
	);
	LUT2 #(
		.INIT('h2)
	) name652 (
		\WX8491_reg/NET0131 ,
		_w2159_,
		_w2160_
	);
	LUT2 #(
		.INIT('h4)
	) name653 (
		\WX8491_reg/NET0131 ,
		_w2159_,
		_w2161_
	);
	LUT2 #(
		.INIT('h1)
	) name654 (
		_w2160_,
		_w2161_,
		_w2162_
	);
	LUT2 #(
		.INIT('h2)
	) name655 (
		\TM1_pad ,
		\WX8427_reg/NET0131 ,
		_w2163_
	);
	LUT2 #(
		.INIT('h4)
	) name656 (
		\TM1_pad ,
		\WX8427_reg/NET0131 ,
		_w2164_
	);
	LUT2 #(
		.INIT('h1)
	) name657 (
		_w2163_,
		_w2164_,
		_w2165_
	);
	LUT2 #(
		.INIT('h4)
	) name658 (
		_w2162_,
		_w2165_,
		_w2166_
	);
	LUT2 #(
		.INIT('h2)
	) name659 (
		_w2162_,
		_w2165_,
		_w2167_
	);
	LUT2 #(
		.INIT('h1)
	) name660 (
		\TM0_pad ,
		_w2166_,
		_w2168_
	);
	LUT2 #(
		.INIT('h4)
	) name661 (
		_w2167_,
		_w2168_,
		_w2169_
	);
	LUT2 #(
		.INIT('h1)
	) name662 (
		_w1653_,
		_w2169_,
		_w2170_
	);
	LUT2 #(
		.INIT('h2)
	) name663 (
		_w1973_,
		_w2170_,
		_w2171_
	);
	LUT2 #(
		.INIT('h1)
	) name664 (
		_w2156_,
		_w2171_,
		_w2172_
	);
	LUT2 #(
		.INIT('h8)
	) name665 (
		\TM0_pad ,
		\_2321__reg/NET0131 ,
		_w2173_
	);
	LUT2 #(
		.INIT('h2)
	) name666 (
		\WX11139_reg/NET0131 ,
		\WX11203_reg/NET0131 ,
		_w2174_
	);
	LUT2 #(
		.INIT('h4)
	) name667 (
		\WX11139_reg/NET0131 ,
		\WX11203_reg/NET0131 ,
		_w2175_
	);
	LUT2 #(
		.INIT('h1)
	) name668 (
		_w2174_,
		_w2175_,
		_w2176_
	);
	LUT2 #(
		.INIT('h2)
	) name669 (
		\WX11075_reg/NET0131 ,
		_w2176_,
		_w2177_
	);
	LUT2 #(
		.INIT('h4)
	) name670 (
		\WX11075_reg/NET0131 ,
		_w2176_,
		_w2178_
	);
	LUT2 #(
		.INIT('h1)
	) name671 (
		_w2177_,
		_w2178_,
		_w2179_
	);
	LUT2 #(
		.INIT('h2)
	) name672 (
		\TM1_pad ,
		\WX11011_reg/NET0131 ,
		_w2180_
	);
	LUT2 #(
		.INIT('h4)
	) name673 (
		\TM1_pad ,
		\WX11011_reg/NET0131 ,
		_w2181_
	);
	LUT2 #(
		.INIT('h1)
	) name674 (
		_w2180_,
		_w2181_,
		_w2182_
	);
	LUT2 #(
		.INIT('h4)
	) name675 (
		_w2179_,
		_w2182_,
		_w2183_
	);
	LUT2 #(
		.INIT('h2)
	) name676 (
		_w2179_,
		_w2182_,
		_w2184_
	);
	LUT2 #(
		.INIT('h1)
	) name677 (
		\TM0_pad ,
		_w2183_,
		_w2185_
	);
	LUT2 #(
		.INIT('h4)
	) name678 (
		_w2184_,
		_w2185_,
		_w2186_
	);
	LUT2 #(
		.INIT('h1)
	) name679 (
		_w2173_,
		_w2186_,
		_w2187_
	);
	LUT2 #(
		.INIT('h2)
	) name680 (
		_w1976_,
		_w2187_,
		_w2188_
	);
	LUT2 #(
		.INIT('h2)
	) name681 (
		\WX9846_reg/NET0131 ,
		\WX9910_reg/NET0131 ,
		_w2189_
	);
	LUT2 #(
		.INIT('h4)
	) name682 (
		\WX9846_reg/NET0131 ,
		\WX9910_reg/NET0131 ,
		_w2190_
	);
	LUT2 #(
		.INIT('h1)
	) name683 (
		_w2189_,
		_w2190_,
		_w2191_
	);
	LUT2 #(
		.INIT('h2)
	) name684 (
		\WX9782_reg/NET0131 ,
		_w2191_,
		_w2192_
	);
	LUT2 #(
		.INIT('h4)
	) name685 (
		\WX9782_reg/NET0131 ,
		_w2191_,
		_w2193_
	);
	LUT2 #(
		.INIT('h1)
	) name686 (
		_w2192_,
		_w2193_,
		_w2194_
	);
	LUT2 #(
		.INIT('h2)
	) name687 (
		\TM1_pad ,
		\WX9718_reg/NET0131 ,
		_w2195_
	);
	LUT2 #(
		.INIT('h4)
	) name688 (
		\TM1_pad ,
		\WX9718_reg/NET0131 ,
		_w2196_
	);
	LUT2 #(
		.INIT('h1)
	) name689 (
		_w2195_,
		_w2196_,
		_w2197_
	);
	LUT2 #(
		.INIT('h4)
	) name690 (
		_w2194_,
		_w2197_,
		_w2198_
	);
	LUT2 #(
		.INIT('h2)
	) name691 (
		_w2194_,
		_w2197_,
		_w2199_
	);
	LUT2 #(
		.INIT('h1)
	) name692 (
		\TM0_pad ,
		_w2198_,
		_w2200_
	);
	LUT2 #(
		.INIT('h4)
	) name693 (
		_w2199_,
		_w2200_,
		_w2201_
	);
	LUT2 #(
		.INIT('h1)
	) name694 (
		_w1682_,
		_w2201_,
		_w2202_
	);
	LUT2 #(
		.INIT('h2)
	) name695 (
		_w1973_,
		_w2202_,
		_w2203_
	);
	LUT2 #(
		.INIT('h1)
	) name696 (
		_w2188_,
		_w2203_,
		_w2204_
	);
	LUT2 #(
		.INIT('h8)
	) name697 (
		\TM0_pad ,
		\_2189__reg/NET0131 ,
		_w2205_
	);
	LUT2 #(
		.INIT('h2)
	) name698 (
		\WX5975_reg/NET0131 ,
		\WX6039_reg/NET0131 ,
		_w2206_
	);
	LUT2 #(
		.INIT('h4)
	) name699 (
		\WX5975_reg/NET0131 ,
		\WX6039_reg/NET0131 ,
		_w2207_
	);
	LUT2 #(
		.INIT('h1)
	) name700 (
		_w2206_,
		_w2207_,
		_w2208_
	);
	LUT2 #(
		.INIT('h2)
	) name701 (
		\WX5911_reg/NET0131 ,
		_w2208_,
		_w2209_
	);
	LUT2 #(
		.INIT('h4)
	) name702 (
		\WX5911_reg/NET0131 ,
		_w2208_,
		_w2210_
	);
	LUT2 #(
		.INIT('h1)
	) name703 (
		_w2209_,
		_w2210_,
		_w2211_
	);
	LUT2 #(
		.INIT('h2)
	) name704 (
		\TM1_pad ,
		\WX5847_reg/NET0131 ,
		_w2212_
	);
	LUT2 #(
		.INIT('h4)
	) name705 (
		\TM1_pad ,
		\WX5847_reg/NET0131 ,
		_w2213_
	);
	LUT2 #(
		.INIT('h1)
	) name706 (
		_w2212_,
		_w2213_,
		_w2214_
	);
	LUT2 #(
		.INIT('h4)
	) name707 (
		_w2211_,
		_w2214_,
		_w2215_
	);
	LUT2 #(
		.INIT('h2)
	) name708 (
		_w2211_,
		_w2214_,
		_w2216_
	);
	LUT2 #(
		.INIT('h1)
	) name709 (
		\TM0_pad ,
		_w2215_,
		_w2217_
	);
	LUT2 #(
		.INIT('h4)
	) name710 (
		_w2216_,
		_w2217_,
		_w2218_
	);
	LUT2 #(
		.INIT('h1)
	) name711 (
		_w2205_,
		_w2218_,
		_w2219_
	);
	LUT2 #(
		.INIT('h2)
	) name712 (
		_w1976_,
		_w2219_,
		_w2220_
	);
	LUT2 #(
		.INIT('h2)
	) name713 (
		\WX4682_reg/NET0131 ,
		\WX4746_reg/NET0131 ,
		_w2221_
	);
	LUT2 #(
		.INIT('h4)
	) name714 (
		\WX4682_reg/NET0131 ,
		\WX4746_reg/NET0131 ,
		_w2222_
	);
	LUT2 #(
		.INIT('h1)
	) name715 (
		_w2221_,
		_w2222_,
		_w2223_
	);
	LUT2 #(
		.INIT('h2)
	) name716 (
		\WX4618_reg/NET0131 ,
		_w2223_,
		_w2224_
	);
	LUT2 #(
		.INIT('h4)
	) name717 (
		\WX4618_reg/NET0131 ,
		_w2223_,
		_w2225_
	);
	LUT2 #(
		.INIT('h1)
	) name718 (
		_w2224_,
		_w2225_,
		_w2226_
	);
	LUT2 #(
		.INIT('h2)
	) name719 (
		\TM1_pad ,
		\WX4554_reg/NET0131 ,
		_w2227_
	);
	LUT2 #(
		.INIT('h4)
	) name720 (
		\TM1_pad ,
		\WX4554_reg/NET0131 ,
		_w2228_
	);
	LUT2 #(
		.INIT('h1)
	) name721 (
		_w2227_,
		_w2228_,
		_w2229_
	);
	LUT2 #(
		.INIT('h4)
	) name722 (
		_w2226_,
		_w2229_,
		_w2230_
	);
	LUT2 #(
		.INIT('h2)
	) name723 (
		_w2226_,
		_w2229_,
		_w2231_
	);
	LUT2 #(
		.INIT('h1)
	) name724 (
		\TM0_pad ,
		_w2230_,
		_w2232_
	);
	LUT2 #(
		.INIT('h4)
	) name725 (
		_w2231_,
		_w2232_,
		_w2233_
	);
	LUT2 #(
		.INIT('h1)
	) name726 (
		_w1605_,
		_w2233_,
		_w2234_
	);
	LUT2 #(
		.INIT('h2)
	) name727 (
		_w1973_,
		_w2234_,
		_w2235_
	);
	LUT2 #(
		.INIT('h1)
	) name728 (
		_w2220_,
		_w2235_,
		_w2236_
	);
	LUT2 #(
		.INIT('h8)
	) name729 (
		\TM0_pad ,
		\_2222__reg/NET0131 ,
		_w2237_
	);
	LUT2 #(
		.INIT('h2)
	) name730 (
		\WX7266_reg/NET0131 ,
		\WX7330_reg/NET0131 ,
		_w2238_
	);
	LUT2 #(
		.INIT('h4)
	) name731 (
		\WX7266_reg/NET0131 ,
		\WX7330_reg/NET0131 ,
		_w2239_
	);
	LUT2 #(
		.INIT('h1)
	) name732 (
		_w2238_,
		_w2239_,
		_w2240_
	);
	LUT2 #(
		.INIT('h2)
	) name733 (
		\WX7202_reg/NET0131 ,
		_w2240_,
		_w2241_
	);
	LUT2 #(
		.INIT('h4)
	) name734 (
		\WX7202_reg/NET0131 ,
		_w2240_,
		_w2242_
	);
	LUT2 #(
		.INIT('h1)
	) name735 (
		_w2241_,
		_w2242_,
		_w2243_
	);
	LUT2 #(
		.INIT('h2)
	) name736 (
		\TM1_pad ,
		\WX7138_reg/NET0131 ,
		_w2244_
	);
	LUT2 #(
		.INIT('h4)
	) name737 (
		\TM1_pad ,
		\WX7138_reg/NET0131 ,
		_w2245_
	);
	LUT2 #(
		.INIT('h1)
	) name738 (
		_w2244_,
		_w2245_,
		_w2246_
	);
	LUT2 #(
		.INIT('h4)
	) name739 (
		_w2243_,
		_w2246_,
		_w2247_
	);
	LUT2 #(
		.INIT('h2)
	) name740 (
		_w2243_,
		_w2246_,
		_w2248_
	);
	LUT2 #(
		.INIT('h1)
	) name741 (
		\TM0_pad ,
		_w2247_,
		_w2249_
	);
	LUT2 #(
		.INIT('h4)
	) name742 (
		_w2248_,
		_w2249_,
		_w2250_
	);
	LUT2 #(
		.INIT('h1)
	) name743 (
		_w2237_,
		_w2250_,
		_w2251_
	);
	LUT2 #(
		.INIT('h2)
	) name744 (
		_w1976_,
		_w2251_,
		_w2252_
	);
	LUT2 #(
		.INIT('h2)
	) name745 (
		\WX5973_reg/NET0131 ,
		\WX6037_reg/NET0131 ,
		_w2253_
	);
	LUT2 #(
		.INIT('h4)
	) name746 (
		\WX5973_reg/NET0131 ,
		\WX6037_reg/NET0131 ,
		_w2254_
	);
	LUT2 #(
		.INIT('h1)
	) name747 (
		_w2253_,
		_w2254_,
		_w2255_
	);
	LUT2 #(
		.INIT('h2)
	) name748 (
		\WX5909_reg/NET0131 ,
		_w2255_,
		_w2256_
	);
	LUT2 #(
		.INIT('h4)
	) name749 (
		\WX5909_reg/NET0131 ,
		_w2255_,
		_w2257_
	);
	LUT2 #(
		.INIT('h1)
	) name750 (
		_w2256_,
		_w2257_,
		_w2258_
	);
	LUT2 #(
		.INIT('h2)
	) name751 (
		\TM1_pad ,
		\WX5845_reg/NET0131 ,
		_w2259_
	);
	LUT2 #(
		.INIT('h4)
	) name752 (
		\TM1_pad ,
		\WX5845_reg/NET0131 ,
		_w2260_
	);
	LUT2 #(
		.INIT('h1)
	) name753 (
		_w2259_,
		_w2260_,
		_w2261_
	);
	LUT2 #(
		.INIT('h4)
	) name754 (
		_w2258_,
		_w2261_,
		_w2262_
	);
	LUT2 #(
		.INIT('h2)
	) name755 (
		_w2258_,
		_w2261_,
		_w2263_
	);
	LUT2 #(
		.INIT('h1)
	) name756 (
		\TM0_pad ,
		_w2262_,
		_w2264_
	);
	LUT2 #(
		.INIT('h4)
	) name757 (
		_w2263_,
		_w2264_,
		_w2265_
	);
	LUT2 #(
		.INIT('h1)
	) name758 (
		_w1621_,
		_w2265_,
		_w2266_
	);
	LUT2 #(
		.INIT('h2)
	) name759 (
		_w1973_,
		_w2266_,
		_w2267_
	);
	LUT2 #(
		.INIT('h1)
	) name760 (
		_w2252_,
		_w2267_,
		_w2268_
	);
	LUT2 #(
		.INIT('h8)
	) name761 (
		\TM0_pad ,
		\_2255__reg/NET0131 ,
		_w2269_
	);
	LUT2 #(
		.INIT('h2)
	) name762 (
		\WX8557_reg/NET0131 ,
		\WX8621_reg/NET0131 ,
		_w2270_
	);
	LUT2 #(
		.INIT('h4)
	) name763 (
		\WX8557_reg/NET0131 ,
		\WX8621_reg/NET0131 ,
		_w2271_
	);
	LUT2 #(
		.INIT('h1)
	) name764 (
		_w2270_,
		_w2271_,
		_w2272_
	);
	LUT2 #(
		.INIT('h2)
	) name765 (
		\WX8493_reg/NET0131 ,
		_w2272_,
		_w2273_
	);
	LUT2 #(
		.INIT('h4)
	) name766 (
		\WX8493_reg/NET0131 ,
		_w2272_,
		_w2274_
	);
	LUT2 #(
		.INIT('h1)
	) name767 (
		_w2273_,
		_w2274_,
		_w2275_
	);
	LUT2 #(
		.INIT('h2)
	) name768 (
		\TM1_pad ,
		\WX8429_reg/NET0131 ,
		_w2276_
	);
	LUT2 #(
		.INIT('h4)
	) name769 (
		\TM1_pad ,
		\WX8429_reg/NET0131 ,
		_w2277_
	);
	LUT2 #(
		.INIT('h1)
	) name770 (
		_w2276_,
		_w2277_,
		_w2278_
	);
	LUT2 #(
		.INIT('h4)
	) name771 (
		_w2275_,
		_w2278_,
		_w2279_
	);
	LUT2 #(
		.INIT('h2)
	) name772 (
		_w2275_,
		_w2278_,
		_w2280_
	);
	LUT2 #(
		.INIT('h1)
	) name773 (
		\TM0_pad ,
		_w2279_,
		_w2281_
	);
	LUT2 #(
		.INIT('h4)
	) name774 (
		_w2280_,
		_w2281_,
		_w2282_
	);
	LUT2 #(
		.INIT('h1)
	) name775 (
		_w2269_,
		_w2282_,
		_w2283_
	);
	LUT2 #(
		.INIT('h2)
	) name776 (
		_w1976_,
		_w2283_,
		_w2284_
	);
	LUT2 #(
		.INIT('h2)
	) name777 (
		\WX7264_reg/NET0131 ,
		\WX7328_reg/NET0131 ,
		_w2285_
	);
	LUT2 #(
		.INIT('h4)
	) name778 (
		\WX7264_reg/NET0131 ,
		\WX7328_reg/NET0131 ,
		_w2286_
	);
	LUT2 #(
		.INIT('h1)
	) name779 (
		_w2285_,
		_w2286_,
		_w2287_
	);
	LUT2 #(
		.INIT('h2)
	) name780 (
		\WX7200_reg/NET0131 ,
		_w2287_,
		_w2288_
	);
	LUT2 #(
		.INIT('h4)
	) name781 (
		\WX7200_reg/NET0131 ,
		_w2287_,
		_w2289_
	);
	LUT2 #(
		.INIT('h1)
	) name782 (
		_w2288_,
		_w2289_,
		_w2290_
	);
	LUT2 #(
		.INIT('h2)
	) name783 (
		\TM1_pad ,
		\WX7136_reg/NET0131 ,
		_w2291_
	);
	LUT2 #(
		.INIT('h4)
	) name784 (
		\TM1_pad ,
		\WX7136_reg/NET0131 ,
		_w2292_
	);
	LUT2 #(
		.INIT('h1)
	) name785 (
		_w2291_,
		_w2292_,
		_w2293_
	);
	LUT2 #(
		.INIT('h4)
	) name786 (
		_w2290_,
		_w2293_,
		_w2294_
	);
	LUT2 #(
		.INIT('h2)
	) name787 (
		_w2290_,
		_w2293_,
		_w2295_
	);
	LUT2 #(
		.INIT('h1)
	) name788 (
		\TM0_pad ,
		_w2294_,
		_w2296_
	);
	LUT2 #(
		.INIT('h4)
	) name789 (
		_w2295_,
		_w2296_,
		_w2297_
	);
	LUT2 #(
		.INIT('h1)
	) name790 (
		_w1637_,
		_w2297_,
		_w2298_
	);
	LUT2 #(
		.INIT('h2)
	) name791 (
		_w1973_,
		_w2298_,
		_w2299_
	);
	LUT2 #(
		.INIT('h1)
	) name792 (
		_w2284_,
		_w2299_,
		_w2300_
	);
	LUT2 #(
		.INIT('h1)
	) name793 (
		\TM0_pad ,
		_w1819_,
		_w2301_
	);
	LUT2 #(
		.INIT('h1)
	) name794 (
		_w1810_,
		_w2301_,
		_w2302_
	);
	LUT2 #(
		.INIT('h2)
	) name795 (
		_w1973_,
		_w2302_,
		_w2303_
	);
	LUT2 #(
		.INIT('h8)
	) name796 (
		\TM0_pad ,
		\_2105__reg/NET0131 ,
		_w2304_
	);
	LUT2 #(
		.INIT('h2)
	) name797 (
		\WX2072_reg/NET0131 ,
		\WX2136_reg/NET0131 ,
		_w2305_
	);
	LUT2 #(
		.INIT('h4)
	) name798 (
		\WX2072_reg/NET0131 ,
		\WX2136_reg/NET0131 ,
		_w2306_
	);
	LUT2 #(
		.INIT('h1)
	) name799 (
		_w2305_,
		_w2306_,
		_w2307_
	);
	LUT2 #(
		.INIT('h2)
	) name800 (
		\WX2008_reg/NET0131 ,
		_w2307_,
		_w2308_
	);
	LUT2 #(
		.INIT('h4)
	) name801 (
		\WX2008_reg/NET0131 ,
		_w2307_,
		_w2309_
	);
	LUT2 #(
		.INIT('h1)
	) name802 (
		_w2308_,
		_w2309_,
		_w2310_
	);
	LUT2 #(
		.INIT('h2)
	) name803 (
		\TM1_pad ,
		\WX1944_reg/NET0131 ,
		_w2311_
	);
	LUT2 #(
		.INIT('h4)
	) name804 (
		\TM1_pad ,
		\WX1944_reg/NET0131 ,
		_w2312_
	);
	LUT2 #(
		.INIT('h1)
	) name805 (
		_w2311_,
		_w2312_,
		_w2313_
	);
	LUT2 #(
		.INIT('h4)
	) name806 (
		_w2310_,
		_w2313_,
		_w2314_
	);
	LUT2 #(
		.INIT('h2)
	) name807 (
		_w2310_,
		_w2313_,
		_w2315_
	);
	LUT2 #(
		.INIT('h1)
	) name808 (
		\TM0_pad ,
		_w2314_,
		_w2316_
	);
	LUT2 #(
		.INIT('h4)
	) name809 (
		_w2315_,
		_w2316_,
		_w2317_
	);
	LUT2 #(
		.INIT('h1)
	) name810 (
		_w2304_,
		_w2317_,
		_w2318_
	);
	LUT2 #(
		.INIT('h2)
	) name811 (
		_w1976_,
		_w2318_,
		_w2319_
	);
	LUT2 #(
		.INIT('h1)
	) name812 (
		_w2303_,
		_w2319_,
		_w2320_
	);
	LUT2 #(
		.INIT('h2)
	) name813 (
		\WX11119_reg/NET0131 ,
		\WX11183_reg/NET0131 ,
		_w2321_
	);
	LUT2 #(
		.INIT('h4)
	) name814 (
		\WX11119_reg/NET0131 ,
		\WX11183_reg/NET0131 ,
		_w2322_
	);
	LUT2 #(
		.INIT('h1)
	) name815 (
		_w2321_,
		_w2322_,
		_w2323_
	);
	LUT2 #(
		.INIT('h2)
	) name816 (
		\WX11055_reg/NET0131 ,
		_w2323_,
		_w2324_
	);
	LUT2 #(
		.INIT('h4)
	) name817 (
		\WX11055_reg/NET0131 ,
		_w2323_,
		_w2325_
	);
	LUT2 #(
		.INIT('h1)
	) name818 (
		_w2324_,
		_w2325_,
		_w2326_
	);
	LUT2 #(
		.INIT('h2)
	) name819 (
		\TM1_pad ,
		\WX10991_reg/NET0131 ,
		_w2327_
	);
	LUT2 #(
		.INIT('h4)
	) name820 (
		\TM1_pad ,
		\WX10991_reg/NET0131 ,
		_w2328_
	);
	LUT2 #(
		.INIT('h1)
	) name821 (
		_w2327_,
		_w2328_,
		_w2329_
	);
	LUT2 #(
		.INIT('h4)
	) name822 (
		_w2326_,
		_w2329_,
		_w2330_
	);
	LUT2 #(
		.INIT('h2)
	) name823 (
		_w2326_,
		_w2329_,
		_w2331_
	);
	LUT2 #(
		.INIT('h1)
	) name824 (
		\TM0_pad ,
		_w2330_,
		_w2332_
	);
	LUT2 #(
		.INIT('h4)
	) name825 (
		_w2331_,
		_w2332_,
		_w2333_
	);
	LUT2 #(
		.INIT('h1)
	) name826 (
		_w1855_,
		_w2333_,
		_w2334_
	);
	LUT2 #(
		.INIT('h2)
	) name827 (
		_w1973_,
		_w2334_,
		_w2335_
	);
	LUT2 #(
		.INIT('h1)
	) name828 (
		\DATA_0_30_pad ,
		\TM0_pad ,
		_w2336_
	);
	LUT2 #(
		.INIT('h2)
	) name829 (
		\TM0_pad ,
		\_2363__reg/NET0131 ,
		_w2337_
	);
	LUT2 #(
		.INIT('h2)
	) name830 (
		_w1976_,
		_w2336_,
		_w2338_
	);
	LUT2 #(
		.INIT('h4)
	) name831 (
		_w2337_,
		_w2338_,
		_w2339_
	);
	LUT2 #(
		.INIT('h1)
	) name832 (
		_w2335_,
		_w2339_,
		_w2340_
	);
	LUT2 #(
		.INIT('h4)
	) name833 (
		_w1573_,
		_w1973_,
		_w2341_
	);
	LUT2 #(
		.INIT('h2)
	) name834 (
		\WX3393_reg/NET0131 ,
		\WX3457_reg/NET0131 ,
		_w2342_
	);
	LUT2 #(
		.INIT('h4)
	) name835 (
		\WX3393_reg/NET0131 ,
		\WX3457_reg/NET0131 ,
		_w2343_
	);
	LUT2 #(
		.INIT('h1)
	) name836 (
		_w2342_,
		_w2343_,
		_w2344_
	);
	LUT2 #(
		.INIT('h2)
	) name837 (
		\WX3265_reg/NET0131 ,
		\WX3329_reg/NET0131 ,
		_w2345_
	);
	LUT2 #(
		.INIT('h4)
	) name838 (
		\WX3265_reg/NET0131 ,
		\WX3329_reg/NET0131 ,
		_w2346_
	);
	LUT2 #(
		.INIT('h1)
	) name839 (
		_w2345_,
		_w2346_,
		_w2347_
	);
	LUT2 #(
		.INIT('h4)
	) name840 (
		_w2344_,
		_w2347_,
		_w2348_
	);
	LUT2 #(
		.INIT('h2)
	) name841 (
		_w2344_,
		_w2347_,
		_w2349_
	);
	LUT2 #(
		.INIT('h1)
	) name842 (
		\TM0_pad ,
		_w2348_,
		_w2350_
	);
	LUT2 #(
		.INIT('h4)
	) name843 (
		_w2349_,
		_w2350_,
		_w2351_
	);
	LUT2 #(
		.INIT('h2)
	) name844 (
		_w2341_,
		_w2351_,
		_w2352_
	);
	LUT2 #(
		.INIT('h2)
	) name845 (
		\TM0_pad ,
		\_2155__reg/NET0131 ,
		_w2353_
	);
	LUT2 #(
		.INIT('h2)
	) name846 (
		\WX4686_reg/NET0131 ,
		\WX4750_reg/NET0131 ,
		_w2354_
	);
	LUT2 #(
		.INIT('h4)
	) name847 (
		\WX4686_reg/NET0131 ,
		\WX4750_reg/NET0131 ,
		_w2355_
	);
	LUT2 #(
		.INIT('h1)
	) name848 (
		_w2354_,
		_w2355_,
		_w2356_
	);
	LUT2 #(
		.INIT('h2)
	) name849 (
		\WX4558_reg/NET0131 ,
		\WX4622_reg/NET0131 ,
		_w2357_
	);
	LUT2 #(
		.INIT('h4)
	) name850 (
		\WX4558_reg/NET0131 ,
		\WX4622_reg/NET0131 ,
		_w2358_
	);
	LUT2 #(
		.INIT('h1)
	) name851 (
		_w2357_,
		_w2358_,
		_w2359_
	);
	LUT2 #(
		.INIT('h4)
	) name852 (
		_w2356_,
		_w2359_,
		_w2360_
	);
	LUT2 #(
		.INIT('h2)
	) name853 (
		_w2356_,
		_w2359_,
		_w2361_
	);
	LUT2 #(
		.INIT('h1)
	) name854 (
		\TM0_pad ,
		_w2360_,
		_w2362_
	);
	LUT2 #(
		.INIT('h4)
	) name855 (
		_w2361_,
		_w2362_,
		_w2363_
	);
	LUT2 #(
		.INIT('h2)
	) name856 (
		_w1976_,
		_w2353_,
		_w2364_
	);
	LUT2 #(
		.INIT('h4)
	) name857 (
		_w2363_,
		_w2364_,
		_w2365_
	);
	LUT2 #(
		.INIT('h1)
	) name858 (
		_w2352_,
		_w2365_,
		_w2366_
	);
	LUT2 #(
		.INIT('h8)
	) name859 (
		\TM0_pad ,
		\_2287__reg/NET0131 ,
		_w2367_
	);
	LUT2 #(
		.INIT('h2)
	) name860 (
		\WX9850_reg/NET0131 ,
		\WX9914_reg/NET0131 ,
		_w2368_
	);
	LUT2 #(
		.INIT('h4)
	) name861 (
		\WX9850_reg/NET0131 ,
		\WX9914_reg/NET0131 ,
		_w2369_
	);
	LUT2 #(
		.INIT('h1)
	) name862 (
		_w2368_,
		_w2369_,
		_w2370_
	);
	LUT2 #(
		.INIT('h2)
	) name863 (
		\WX9786_reg/NET0131 ,
		_w2370_,
		_w2371_
	);
	LUT2 #(
		.INIT('h4)
	) name864 (
		\WX9786_reg/NET0131 ,
		_w2370_,
		_w2372_
	);
	LUT2 #(
		.INIT('h1)
	) name865 (
		_w2371_,
		_w2372_,
		_w2373_
	);
	LUT2 #(
		.INIT('h2)
	) name866 (
		\TM1_pad ,
		\WX9722_reg/NET0131 ,
		_w2374_
	);
	LUT2 #(
		.INIT('h4)
	) name867 (
		\TM1_pad ,
		\WX9722_reg/NET0131 ,
		_w2375_
	);
	LUT2 #(
		.INIT('h1)
	) name868 (
		_w2374_,
		_w2375_,
		_w2376_
	);
	LUT2 #(
		.INIT('h4)
	) name869 (
		_w2373_,
		_w2376_,
		_w2377_
	);
	LUT2 #(
		.INIT('h2)
	) name870 (
		_w2373_,
		_w2376_,
		_w2378_
	);
	LUT2 #(
		.INIT('h1)
	) name871 (
		\TM0_pad ,
		_w2377_,
		_w2379_
	);
	LUT2 #(
		.INIT('h4)
	) name872 (
		_w2378_,
		_w2379_,
		_w2380_
	);
	LUT2 #(
		.INIT('h1)
	) name873 (
		_w2367_,
		_w2380_,
		_w2381_
	);
	LUT2 #(
		.INIT('h2)
	) name874 (
		_w1976_,
		_w2381_,
		_w2382_
	);
	LUT2 #(
		.INIT('h1)
	) name875 (
		_w1637_,
		_w2282_,
		_w2383_
	);
	LUT2 #(
		.INIT('h2)
	) name876 (
		_w1973_,
		_w2383_,
		_w2384_
	);
	LUT2 #(
		.INIT('h1)
	) name877 (
		_w2382_,
		_w2384_,
		_w2385_
	);
	LUT2 #(
		.INIT('h8)
	) name878 (
		\TM0_pad ,
		\_2138__reg/NET0131 ,
		_w2386_
	);
	LUT2 #(
		.INIT('h2)
	) name879 (
		\WX3363_reg/NET0131 ,
		\WX3427_reg/NET0131 ,
		_w2387_
	);
	LUT2 #(
		.INIT('h4)
	) name880 (
		\WX3363_reg/NET0131 ,
		\WX3427_reg/NET0131 ,
		_w2388_
	);
	LUT2 #(
		.INIT('h1)
	) name881 (
		_w2387_,
		_w2388_,
		_w2389_
	);
	LUT2 #(
		.INIT('h2)
	) name882 (
		\WX3299_reg/NET0131 ,
		_w2389_,
		_w2390_
	);
	LUT2 #(
		.INIT('h4)
	) name883 (
		\WX3299_reg/NET0131 ,
		_w2389_,
		_w2391_
	);
	LUT2 #(
		.INIT('h1)
	) name884 (
		_w2390_,
		_w2391_,
		_w2392_
	);
	LUT2 #(
		.INIT('h2)
	) name885 (
		\TM1_pad ,
		\WX3235_reg/NET0131 ,
		_w2393_
	);
	LUT2 #(
		.INIT('h4)
	) name886 (
		\TM1_pad ,
		\WX3235_reg/NET0131 ,
		_w2394_
	);
	LUT2 #(
		.INIT('h1)
	) name887 (
		_w2393_,
		_w2394_,
		_w2395_
	);
	LUT2 #(
		.INIT('h4)
	) name888 (
		_w2392_,
		_w2395_,
		_w2396_
	);
	LUT2 #(
		.INIT('h2)
	) name889 (
		_w2392_,
		_w2395_,
		_w2397_
	);
	LUT2 #(
		.INIT('h1)
	) name890 (
		\TM0_pad ,
		_w2396_,
		_w2398_
	);
	LUT2 #(
		.INIT('h4)
	) name891 (
		_w2397_,
		_w2398_,
		_w2399_
	);
	LUT2 #(
		.INIT('h1)
	) name892 (
		_w2386_,
		_w2399_,
		_w2400_
	);
	LUT2 #(
		.INIT('h2)
	) name893 (
		_w1976_,
		_w2400_,
		_w2401_
	);
	LUT2 #(
		.INIT('h1)
	) name894 (
		_w1826_,
		_w2093_,
		_w2402_
	);
	LUT2 #(
		.INIT('h2)
	) name895 (
		_w1973_,
		_w2402_,
		_w2403_
	);
	LUT2 #(
		.INIT('h1)
	) name896 (
		_w2401_,
		_w2403_,
		_w2404_
	);
	LUT2 #(
		.INIT('h8)
	) name897 (
		\TM0_pad ,
		\_2320__reg/NET0131 ,
		_w2405_
	);
	LUT2 #(
		.INIT('h2)
	) name898 (
		\WX11141_reg/NET0131 ,
		\WX11205_reg/NET0131 ,
		_w2406_
	);
	LUT2 #(
		.INIT('h4)
	) name899 (
		\WX11141_reg/NET0131 ,
		\WX11205_reg/NET0131 ,
		_w2407_
	);
	LUT2 #(
		.INIT('h1)
	) name900 (
		_w2406_,
		_w2407_,
		_w2408_
	);
	LUT2 #(
		.INIT('h2)
	) name901 (
		\WX11077_reg/NET0131 ,
		_w2408_,
		_w2409_
	);
	LUT2 #(
		.INIT('h4)
	) name902 (
		\WX11077_reg/NET0131 ,
		_w2408_,
		_w2410_
	);
	LUT2 #(
		.INIT('h1)
	) name903 (
		_w2409_,
		_w2410_,
		_w2411_
	);
	LUT2 #(
		.INIT('h2)
	) name904 (
		\TM1_pad ,
		\WX11013_reg/NET0131 ,
		_w2412_
	);
	LUT2 #(
		.INIT('h4)
	) name905 (
		\TM1_pad ,
		\WX11013_reg/NET0131 ,
		_w2413_
	);
	LUT2 #(
		.INIT('h1)
	) name906 (
		_w2412_,
		_w2413_,
		_w2414_
	);
	LUT2 #(
		.INIT('h4)
	) name907 (
		_w2411_,
		_w2414_,
		_w2415_
	);
	LUT2 #(
		.INIT('h2)
	) name908 (
		_w2411_,
		_w2414_,
		_w2416_
	);
	LUT2 #(
		.INIT('h1)
	) name909 (
		\TM0_pad ,
		_w2415_,
		_w2417_
	);
	LUT2 #(
		.INIT('h4)
	) name910 (
		_w2416_,
		_w2417_,
		_w2418_
	);
	LUT2 #(
		.INIT('h1)
	) name911 (
		_w2405_,
		_w2418_,
		_w2419_
	);
	LUT2 #(
		.INIT('h2)
	) name912 (
		_w1976_,
		_w2419_,
		_w2420_
	);
	LUT2 #(
		.INIT('h1)
	) name913 (
		_w1653_,
		_w2154_,
		_w2421_
	);
	LUT2 #(
		.INIT('h2)
	) name914 (
		_w1973_,
		_w2421_,
		_w2422_
	);
	LUT2 #(
		.INIT('h1)
	) name915 (
		_w2420_,
		_w2422_,
		_w2423_
	);
	LUT2 #(
		.INIT('h2)
	) name916 (
		_w1974_,
		_w2118_,
		_w2424_
	);
	LUT2 #(
		.INIT('h2)
	) name917 (
		\TM0_pad ,
		\_2188__reg/NET0131 ,
		_w2425_
	);
	LUT2 #(
		.INIT('h2)
	) name918 (
		\WX5977_reg/NET0131 ,
		\WX6041_reg/NET0131 ,
		_w2426_
	);
	LUT2 #(
		.INIT('h4)
	) name919 (
		\WX5977_reg/NET0131 ,
		\WX6041_reg/NET0131 ,
		_w2427_
	);
	LUT2 #(
		.INIT('h1)
	) name920 (
		_w2426_,
		_w2427_,
		_w2428_
	);
	LUT2 #(
		.INIT('h2)
	) name921 (
		\WX5849_reg/NET0131 ,
		\WX5913_reg/NET0131 ,
		_w2429_
	);
	LUT2 #(
		.INIT('h4)
	) name922 (
		\WX5849_reg/NET0131 ,
		\WX5913_reg/NET0131 ,
		_w2430_
	);
	LUT2 #(
		.INIT('h1)
	) name923 (
		_w2429_,
		_w2430_,
		_w2431_
	);
	LUT2 #(
		.INIT('h4)
	) name924 (
		_w2428_,
		_w2431_,
		_w2432_
	);
	LUT2 #(
		.INIT('h2)
	) name925 (
		_w2428_,
		_w2431_,
		_w2433_
	);
	LUT2 #(
		.INIT('h1)
	) name926 (
		\TM0_pad ,
		_w2432_,
		_w2434_
	);
	LUT2 #(
		.INIT('h4)
	) name927 (
		_w2433_,
		_w2434_,
		_w2435_
	);
	LUT2 #(
		.INIT('h2)
	) name928 (
		_w1976_,
		_w2425_,
		_w2436_
	);
	LUT2 #(
		.INIT('h4)
	) name929 (
		_w2435_,
		_w2436_,
		_w2437_
	);
	LUT2 #(
		.INIT('h1)
	) name930 (
		_w2424_,
		_w2437_,
		_w2438_
	);
	LUT2 #(
		.INIT('h8)
	) name931 (
		\TM0_pad ,
		\_2221__reg/NET0131 ,
		_w2439_
	);
	LUT2 #(
		.INIT('h2)
	) name932 (
		\WX7268_reg/NET0131 ,
		\WX7332_reg/NET0131 ,
		_w2440_
	);
	LUT2 #(
		.INIT('h4)
	) name933 (
		\WX7268_reg/NET0131 ,
		\WX7332_reg/NET0131 ,
		_w2441_
	);
	LUT2 #(
		.INIT('h1)
	) name934 (
		_w2440_,
		_w2441_,
		_w2442_
	);
	LUT2 #(
		.INIT('h2)
	) name935 (
		\WX7204_reg/NET0131 ,
		_w2442_,
		_w2443_
	);
	LUT2 #(
		.INIT('h4)
	) name936 (
		\WX7204_reg/NET0131 ,
		_w2442_,
		_w2444_
	);
	LUT2 #(
		.INIT('h1)
	) name937 (
		_w2443_,
		_w2444_,
		_w2445_
	);
	LUT2 #(
		.INIT('h2)
	) name938 (
		\TM1_pad ,
		\WX7140_reg/NET0131 ,
		_w2446_
	);
	LUT2 #(
		.INIT('h4)
	) name939 (
		\TM1_pad ,
		\WX7140_reg/NET0131 ,
		_w2447_
	);
	LUT2 #(
		.INIT('h1)
	) name940 (
		_w2446_,
		_w2447_,
		_w2448_
	);
	LUT2 #(
		.INIT('h4)
	) name941 (
		_w2445_,
		_w2448_,
		_w2449_
	);
	LUT2 #(
		.INIT('h2)
	) name942 (
		_w2445_,
		_w2448_,
		_w2450_
	);
	LUT2 #(
		.INIT('h1)
	) name943 (
		\TM0_pad ,
		_w2449_,
		_w2451_
	);
	LUT2 #(
		.INIT('h4)
	) name944 (
		_w2450_,
		_w2451_,
		_w2452_
	);
	LUT2 #(
		.INIT('h1)
	) name945 (
		_w2439_,
		_w2452_,
		_w2453_
	);
	LUT2 #(
		.INIT('h2)
	) name946 (
		_w1976_,
		_w2453_,
		_w2454_
	);
	LUT2 #(
		.INIT('h1)
	) name947 (
		_w1605_,
		_w2218_,
		_w2455_
	);
	LUT2 #(
		.INIT('h2)
	) name948 (
		_w1973_,
		_w2455_,
		_w2456_
	);
	LUT2 #(
		.INIT('h1)
	) name949 (
		_w2454_,
		_w2456_,
		_w2457_
	);
	LUT2 #(
		.INIT('h8)
	) name950 (
		\TM0_pad ,
		\_2254__reg/NET0131 ,
		_w2458_
	);
	LUT2 #(
		.INIT('h2)
	) name951 (
		\WX8559_reg/NET0131 ,
		\WX8623_reg/NET0131 ,
		_w2459_
	);
	LUT2 #(
		.INIT('h4)
	) name952 (
		\WX8559_reg/NET0131 ,
		\WX8623_reg/NET0131 ,
		_w2460_
	);
	LUT2 #(
		.INIT('h1)
	) name953 (
		_w2459_,
		_w2460_,
		_w2461_
	);
	LUT2 #(
		.INIT('h2)
	) name954 (
		\WX8495_reg/NET0131 ,
		_w2461_,
		_w2462_
	);
	LUT2 #(
		.INIT('h4)
	) name955 (
		\WX8495_reg/NET0131 ,
		_w2461_,
		_w2463_
	);
	LUT2 #(
		.INIT('h1)
	) name956 (
		_w2462_,
		_w2463_,
		_w2464_
	);
	LUT2 #(
		.INIT('h2)
	) name957 (
		\TM1_pad ,
		\WX8431_reg/NET0131 ,
		_w2465_
	);
	LUT2 #(
		.INIT('h4)
	) name958 (
		\TM1_pad ,
		\WX8431_reg/NET0131 ,
		_w2466_
	);
	LUT2 #(
		.INIT('h1)
	) name959 (
		_w2465_,
		_w2466_,
		_w2467_
	);
	LUT2 #(
		.INIT('h4)
	) name960 (
		_w2464_,
		_w2467_,
		_w2468_
	);
	LUT2 #(
		.INIT('h2)
	) name961 (
		_w2464_,
		_w2467_,
		_w2469_
	);
	LUT2 #(
		.INIT('h1)
	) name962 (
		\TM0_pad ,
		_w2468_,
		_w2470_
	);
	LUT2 #(
		.INIT('h4)
	) name963 (
		_w2469_,
		_w2470_,
		_w2471_
	);
	LUT2 #(
		.INIT('h1)
	) name964 (
		_w2458_,
		_w2471_,
		_w2472_
	);
	LUT2 #(
		.INIT('h2)
	) name965 (
		_w1976_,
		_w2472_,
		_w2473_
	);
	LUT2 #(
		.INIT('h1)
	) name966 (
		_w1621_,
		_w2250_,
		_w2474_
	);
	LUT2 #(
		.INIT('h2)
	) name967 (
		_w1973_,
		_w2474_,
		_w2475_
	);
	LUT2 #(
		.INIT('h1)
	) name968 (
		_w2473_,
		_w2475_,
		_w2476_
	);
	LUT2 #(
		.INIT('h1)
	) name969 (
		\TM0_pad ,
		_w1803_,
		_w2477_
	);
	LUT2 #(
		.INIT('h1)
	) name970 (
		_w1794_,
		_w2477_,
		_w2478_
	);
	LUT2 #(
		.INIT('h2)
	) name971 (
		_w1973_,
		_w2478_,
		_w2479_
	);
	LUT2 #(
		.INIT('h8)
	) name972 (
		\TM0_pad ,
		\_2104__reg/NET0131 ,
		_w2480_
	);
	LUT2 #(
		.INIT('h2)
	) name973 (
		\WX2074_reg/NET0131 ,
		\WX2138_reg/NET0131 ,
		_w2481_
	);
	LUT2 #(
		.INIT('h4)
	) name974 (
		\WX2074_reg/NET0131 ,
		\WX2138_reg/NET0131 ,
		_w2482_
	);
	LUT2 #(
		.INIT('h1)
	) name975 (
		_w2481_,
		_w2482_,
		_w2483_
	);
	LUT2 #(
		.INIT('h2)
	) name976 (
		\WX2010_reg/NET0131 ,
		_w2483_,
		_w2484_
	);
	LUT2 #(
		.INIT('h4)
	) name977 (
		\WX2010_reg/NET0131 ,
		_w2483_,
		_w2485_
	);
	LUT2 #(
		.INIT('h1)
	) name978 (
		_w2484_,
		_w2485_,
		_w2486_
	);
	LUT2 #(
		.INIT('h2)
	) name979 (
		\TM1_pad ,
		\WX1946_reg/NET0131 ,
		_w2487_
	);
	LUT2 #(
		.INIT('h4)
	) name980 (
		\TM1_pad ,
		\WX1946_reg/NET0131 ,
		_w2488_
	);
	LUT2 #(
		.INIT('h1)
	) name981 (
		_w2487_,
		_w2488_,
		_w2489_
	);
	LUT2 #(
		.INIT('h4)
	) name982 (
		_w2486_,
		_w2489_,
		_w2490_
	);
	LUT2 #(
		.INIT('h2)
	) name983 (
		_w2486_,
		_w2489_,
		_w2491_
	);
	LUT2 #(
		.INIT('h1)
	) name984 (
		\TM0_pad ,
		_w2490_,
		_w2492_
	);
	LUT2 #(
		.INIT('h4)
	) name985 (
		_w2491_,
		_w2492_,
		_w2493_
	);
	LUT2 #(
		.INIT('h1)
	) name986 (
		_w2480_,
		_w2493_,
		_w2494_
	);
	LUT2 #(
		.INIT('h2)
	) name987 (
		_w1976_,
		_w2494_,
		_w2495_
	);
	LUT2 #(
		.INIT('h1)
	) name988 (
		_w2479_,
		_w2495_,
		_w2496_
	);
	LUT2 #(
		.INIT('h2)
	) name989 (
		\WX11121_reg/NET0131 ,
		\WX11185_reg/NET0131 ,
		_w2497_
	);
	LUT2 #(
		.INIT('h4)
	) name990 (
		\WX11121_reg/NET0131 ,
		\WX11185_reg/NET0131 ,
		_w2498_
	);
	LUT2 #(
		.INIT('h1)
	) name991 (
		_w2497_,
		_w2498_,
		_w2499_
	);
	LUT2 #(
		.INIT('h2)
	) name992 (
		\WX11057_reg/NET0131 ,
		_w2499_,
		_w2500_
	);
	LUT2 #(
		.INIT('h4)
	) name993 (
		\WX11057_reg/NET0131 ,
		_w2499_,
		_w2501_
	);
	LUT2 #(
		.INIT('h1)
	) name994 (
		_w2500_,
		_w2501_,
		_w2502_
	);
	LUT2 #(
		.INIT('h2)
	) name995 (
		\TM1_pad ,
		\WX10993_reg/NET0131 ,
		_w2503_
	);
	LUT2 #(
		.INIT('h4)
	) name996 (
		\TM1_pad ,
		\WX10993_reg/NET0131 ,
		_w2504_
	);
	LUT2 #(
		.INIT('h1)
	) name997 (
		_w2503_,
		_w2504_,
		_w2505_
	);
	LUT2 #(
		.INIT('h4)
	) name998 (
		_w2502_,
		_w2505_,
		_w2506_
	);
	LUT2 #(
		.INIT('h2)
	) name999 (
		_w2502_,
		_w2505_,
		_w2507_
	);
	LUT2 #(
		.INIT('h1)
	) name1000 (
		\TM0_pad ,
		_w2506_,
		_w2508_
	);
	LUT2 #(
		.INIT('h4)
	) name1001 (
		_w2507_,
		_w2508_,
		_w2509_
	);
	LUT2 #(
		.INIT('h1)
	) name1002 (
		_w1826_,
		_w2509_,
		_w2510_
	);
	LUT2 #(
		.INIT('h2)
	) name1003 (
		_w1973_,
		_w2510_,
		_w2511_
	);
	LUT2 #(
		.INIT('h1)
	) name1004 (
		\DATA_0_29_pad ,
		\TM0_pad ,
		_w2512_
	);
	LUT2 #(
		.INIT('h2)
	) name1005 (
		\TM0_pad ,
		\_2362__reg/NET0131 ,
		_w2513_
	);
	LUT2 #(
		.INIT('h2)
	) name1006 (
		_w1976_,
		_w2512_,
		_w2514_
	);
	LUT2 #(
		.INIT('h4)
	) name1007 (
		_w2513_,
		_w2514_,
		_w2515_
	);
	LUT2 #(
		.INIT('h1)
	) name1008 (
		_w2511_,
		_w2515_,
		_w2516_
	);
	LUT2 #(
		.INIT('h8)
	) name1009 (
		RESET_pad,
		\WX10831_reg/NET0131 ,
		_w2517_
	);
	LUT2 #(
		.INIT('h2)
	) name1010 (
		\WX3395_reg/NET0131 ,
		\WX3459_reg/NET0131 ,
		_w2518_
	);
	LUT2 #(
		.INIT('h4)
	) name1011 (
		\WX3395_reg/NET0131 ,
		\WX3459_reg/NET0131 ,
		_w2519_
	);
	LUT2 #(
		.INIT('h1)
	) name1012 (
		_w2518_,
		_w2519_,
		_w2520_
	);
	LUT2 #(
		.INIT('h2)
	) name1013 (
		\WX3267_reg/NET0131 ,
		\WX3331_reg/NET0131 ,
		_w2521_
	);
	LUT2 #(
		.INIT('h4)
	) name1014 (
		\WX3267_reg/NET0131 ,
		\WX3331_reg/NET0131 ,
		_w2522_
	);
	LUT2 #(
		.INIT('h1)
	) name1015 (
		_w2521_,
		_w2522_,
		_w2523_
	);
	LUT2 #(
		.INIT('h4)
	) name1016 (
		_w2520_,
		_w2523_,
		_w2524_
	);
	LUT2 #(
		.INIT('h2)
	) name1017 (
		_w2520_,
		_w2523_,
		_w2525_
	);
	LUT2 #(
		.INIT('h1)
	) name1018 (
		\TM0_pad ,
		_w2524_,
		_w2526_
	);
	LUT2 #(
		.INIT('h4)
	) name1019 (
		_w2525_,
		_w2526_,
		_w2527_
	);
	LUT2 #(
		.INIT('h2)
	) name1020 (
		_w2040_,
		_w2527_,
		_w2528_
	);
	LUT2 #(
		.INIT('h2)
	) name1021 (
		\TM0_pad ,
		\_2154__reg/NET0131 ,
		_w2529_
	);
	LUT2 #(
		.INIT('h2)
	) name1022 (
		\WX4688_reg/NET0131 ,
		\WX4752_reg/NET0131 ,
		_w2530_
	);
	LUT2 #(
		.INIT('h4)
	) name1023 (
		\WX4688_reg/NET0131 ,
		\WX4752_reg/NET0131 ,
		_w2531_
	);
	LUT2 #(
		.INIT('h1)
	) name1024 (
		_w2530_,
		_w2531_,
		_w2532_
	);
	LUT2 #(
		.INIT('h2)
	) name1025 (
		\WX4560_reg/NET0131 ,
		\WX4624_reg/NET0131 ,
		_w2533_
	);
	LUT2 #(
		.INIT('h4)
	) name1026 (
		\WX4560_reg/NET0131 ,
		\WX4624_reg/NET0131 ,
		_w2534_
	);
	LUT2 #(
		.INIT('h1)
	) name1027 (
		_w2533_,
		_w2534_,
		_w2535_
	);
	LUT2 #(
		.INIT('h4)
	) name1028 (
		_w2532_,
		_w2535_,
		_w2536_
	);
	LUT2 #(
		.INIT('h2)
	) name1029 (
		_w2532_,
		_w2535_,
		_w2537_
	);
	LUT2 #(
		.INIT('h1)
	) name1030 (
		\TM0_pad ,
		_w2536_,
		_w2538_
	);
	LUT2 #(
		.INIT('h4)
	) name1031 (
		_w2537_,
		_w2538_,
		_w2539_
	);
	LUT2 #(
		.INIT('h2)
	) name1032 (
		_w1976_,
		_w2529_,
		_w2540_
	);
	LUT2 #(
		.INIT('h4)
	) name1033 (
		_w2539_,
		_w2540_,
		_w2541_
	);
	LUT2 #(
		.INIT('h1)
	) name1034 (
		_w2528_,
		_w2541_,
		_w2542_
	);
	LUT2 #(
		.INIT('h8)
	) name1035 (
		\TM0_pad ,
		\_2286__reg/NET0131 ,
		_w2543_
	);
	LUT2 #(
		.INIT('h2)
	) name1036 (
		\WX9852_reg/NET0131 ,
		\WX9916_reg/NET0131 ,
		_w2544_
	);
	LUT2 #(
		.INIT('h4)
	) name1037 (
		\WX9852_reg/NET0131 ,
		\WX9916_reg/NET0131 ,
		_w2545_
	);
	LUT2 #(
		.INIT('h1)
	) name1038 (
		_w2544_,
		_w2545_,
		_w2546_
	);
	LUT2 #(
		.INIT('h2)
	) name1039 (
		\WX9788_reg/NET0131 ,
		_w2546_,
		_w2547_
	);
	LUT2 #(
		.INIT('h4)
	) name1040 (
		\WX9788_reg/NET0131 ,
		_w2546_,
		_w2548_
	);
	LUT2 #(
		.INIT('h1)
	) name1041 (
		_w2547_,
		_w2548_,
		_w2549_
	);
	LUT2 #(
		.INIT('h2)
	) name1042 (
		\TM1_pad ,
		\WX9724_reg/NET0131 ,
		_w2550_
	);
	LUT2 #(
		.INIT('h4)
	) name1043 (
		\TM1_pad ,
		\WX9724_reg/NET0131 ,
		_w2551_
	);
	LUT2 #(
		.INIT('h1)
	) name1044 (
		_w2550_,
		_w2551_,
		_w2552_
	);
	LUT2 #(
		.INIT('h4)
	) name1045 (
		_w2549_,
		_w2552_,
		_w2553_
	);
	LUT2 #(
		.INIT('h2)
	) name1046 (
		_w2549_,
		_w2552_,
		_w2554_
	);
	LUT2 #(
		.INIT('h1)
	) name1047 (
		\TM0_pad ,
		_w2553_,
		_w2555_
	);
	LUT2 #(
		.INIT('h4)
	) name1048 (
		_w2554_,
		_w2555_,
		_w2556_
	);
	LUT2 #(
		.INIT('h1)
	) name1049 (
		_w2543_,
		_w2556_,
		_w2557_
	);
	LUT2 #(
		.INIT('h2)
	) name1050 (
		_w1976_,
		_w2557_,
		_w2558_
	);
	LUT2 #(
		.INIT('h1)
	) name1051 (
		_w1621_,
		_w2471_,
		_w2559_
	);
	LUT2 #(
		.INIT('h2)
	) name1052 (
		_w1973_,
		_w2559_,
		_w2560_
	);
	LUT2 #(
		.INIT('h1)
	) name1053 (
		_w2558_,
		_w2560_,
		_w2561_
	);
	LUT2 #(
		.INIT('h8)
	) name1054 (
		\TM0_pad ,
		\_2137__reg/NET0131 ,
		_w2562_
	);
	LUT2 #(
		.INIT('h2)
	) name1055 (
		\WX3365_reg/NET0131 ,
		\WX3429_reg/NET0131 ,
		_w2563_
	);
	LUT2 #(
		.INIT('h4)
	) name1056 (
		\WX3365_reg/NET0131 ,
		\WX3429_reg/NET0131 ,
		_w2564_
	);
	LUT2 #(
		.INIT('h1)
	) name1057 (
		_w2563_,
		_w2564_,
		_w2565_
	);
	LUT2 #(
		.INIT('h2)
	) name1058 (
		\WX3301_reg/NET0131 ,
		_w2565_,
		_w2566_
	);
	LUT2 #(
		.INIT('h4)
	) name1059 (
		\WX3301_reg/NET0131 ,
		_w2565_,
		_w2567_
	);
	LUT2 #(
		.INIT('h1)
	) name1060 (
		_w2566_,
		_w2567_,
		_w2568_
	);
	LUT2 #(
		.INIT('h2)
	) name1061 (
		\TM1_pad ,
		\WX3237_reg/NET0131 ,
		_w2569_
	);
	LUT2 #(
		.INIT('h4)
	) name1062 (
		\TM1_pad ,
		\WX3237_reg/NET0131 ,
		_w2570_
	);
	LUT2 #(
		.INIT('h1)
	) name1063 (
		_w2569_,
		_w2570_,
		_w2571_
	);
	LUT2 #(
		.INIT('h4)
	) name1064 (
		_w2568_,
		_w2571_,
		_w2572_
	);
	LUT2 #(
		.INIT('h2)
	) name1065 (
		_w2568_,
		_w2571_,
		_w2573_
	);
	LUT2 #(
		.INIT('h1)
	) name1066 (
		\TM0_pad ,
		_w2572_,
		_w2574_
	);
	LUT2 #(
		.INIT('h4)
	) name1067 (
		_w2573_,
		_w2574_,
		_w2575_
	);
	LUT2 #(
		.INIT('h1)
	) name1068 (
		_w2562_,
		_w2575_,
		_w2576_
	);
	LUT2 #(
		.INIT('h2)
	) name1069 (
		_w1976_,
		_w2576_,
		_w2577_
	);
	LUT2 #(
		.INIT('h1)
	) name1070 (
		_w1810_,
		_w2317_,
		_w2578_
	);
	LUT2 #(
		.INIT('h2)
	) name1071 (
		_w1973_,
		_w2578_,
		_w2579_
	);
	LUT2 #(
		.INIT('h1)
	) name1072 (
		_w2577_,
		_w2579_,
		_w2580_
	);
	LUT2 #(
		.INIT('h8)
	) name1073 (
		\TM0_pad ,
		\_2319__reg/NET0131 ,
		_w2581_
	);
	LUT2 #(
		.INIT('h2)
	) name1074 (
		\WX11143_reg/NET0131 ,
		\WX11207_reg/NET0131 ,
		_w2582_
	);
	LUT2 #(
		.INIT('h4)
	) name1075 (
		\WX11143_reg/NET0131 ,
		\WX11207_reg/NET0131 ,
		_w2583_
	);
	LUT2 #(
		.INIT('h1)
	) name1076 (
		_w2582_,
		_w2583_,
		_w2584_
	);
	LUT2 #(
		.INIT('h2)
	) name1077 (
		\WX11079_reg/NET0131 ,
		_w2584_,
		_w2585_
	);
	LUT2 #(
		.INIT('h4)
	) name1078 (
		\WX11079_reg/NET0131 ,
		_w2584_,
		_w2586_
	);
	LUT2 #(
		.INIT('h1)
	) name1079 (
		_w2585_,
		_w2586_,
		_w2587_
	);
	LUT2 #(
		.INIT('h2)
	) name1080 (
		\TM1_pad ,
		\WX11015_reg/NET0131 ,
		_w2588_
	);
	LUT2 #(
		.INIT('h4)
	) name1081 (
		\TM1_pad ,
		\WX11015_reg/NET0131 ,
		_w2589_
	);
	LUT2 #(
		.INIT('h1)
	) name1082 (
		_w2588_,
		_w2589_,
		_w2590_
	);
	LUT2 #(
		.INIT('h4)
	) name1083 (
		_w2587_,
		_w2590_,
		_w2591_
	);
	LUT2 #(
		.INIT('h2)
	) name1084 (
		_w2587_,
		_w2590_,
		_w2592_
	);
	LUT2 #(
		.INIT('h1)
	) name1085 (
		\TM0_pad ,
		_w2591_,
		_w2593_
	);
	LUT2 #(
		.INIT('h4)
	) name1086 (
		_w2592_,
		_w2593_,
		_w2594_
	);
	LUT2 #(
		.INIT('h1)
	) name1087 (
		_w2581_,
		_w2594_,
		_w2595_
	);
	LUT2 #(
		.INIT('h2)
	) name1088 (
		_w1976_,
		_w2595_,
		_w2596_
	);
	LUT2 #(
		.INIT('h1)
	) name1089 (
		_w1637_,
		_w2380_,
		_w2597_
	);
	LUT2 #(
		.INIT('h2)
	) name1090 (
		_w1973_,
		_w2597_,
		_w2598_
	);
	LUT2 #(
		.INIT('h1)
	) name1091 (
		_w2596_,
		_w2598_,
		_w2599_
	);
	LUT2 #(
		.INIT('h2)
	) name1092 (
		_w2341_,
		_w2363_,
		_w2600_
	);
	LUT2 #(
		.INIT('h2)
	) name1093 (
		\TM0_pad ,
		\_2187__reg/NET0131 ,
		_w2601_
	);
	LUT2 #(
		.INIT('h2)
	) name1094 (
		\WX5979_reg/NET0131 ,
		\WX6043_reg/NET0131 ,
		_w2602_
	);
	LUT2 #(
		.INIT('h4)
	) name1095 (
		\WX5979_reg/NET0131 ,
		\WX6043_reg/NET0131 ,
		_w2603_
	);
	LUT2 #(
		.INIT('h1)
	) name1096 (
		_w2602_,
		_w2603_,
		_w2604_
	);
	LUT2 #(
		.INIT('h2)
	) name1097 (
		\WX5851_reg/NET0131 ,
		\WX5915_reg/NET0131 ,
		_w2605_
	);
	LUT2 #(
		.INIT('h4)
	) name1098 (
		\WX5851_reg/NET0131 ,
		\WX5915_reg/NET0131 ,
		_w2606_
	);
	LUT2 #(
		.INIT('h1)
	) name1099 (
		_w2605_,
		_w2606_,
		_w2607_
	);
	LUT2 #(
		.INIT('h4)
	) name1100 (
		_w2604_,
		_w2607_,
		_w2608_
	);
	LUT2 #(
		.INIT('h2)
	) name1101 (
		_w2604_,
		_w2607_,
		_w2609_
	);
	LUT2 #(
		.INIT('h1)
	) name1102 (
		\TM0_pad ,
		_w2608_,
		_w2610_
	);
	LUT2 #(
		.INIT('h4)
	) name1103 (
		_w2609_,
		_w2610_,
		_w2611_
	);
	LUT2 #(
		.INIT('h2)
	) name1104 (
		_w1976_,
		_w2601_,
		_w2612_
	);
	LUT2 #(
		.INIT('h4)
	) name1105 (
		_w2611_,
		_w2612_,
		_w2613_
	);
	LUT2 #(
		.INIT('h1)
	) name1106 (
		_w2600_,
		_w2613_,
		_w2614_
	);
	LUT2 #(
		.INIT('h2)
	) name1107 (
		_w1974_,
		_w2435_,
		_w2615_
	);
	LUT2 #(
		.INIT('h2)
	) name1108 (
		\TM0_pad ,
		\_2220__reg/NET0131 ,
		_w2616_
	);
	LUT2 #(
		.INIT('h2)
	) name1109 (
		\WX7270_reg/NET0131 ,
		\WX7334_reg/NET0131 ,
		_w2617_
	);
	LUT2 #(
		.INIT('h4)
	) name1110 (
		\WX7270_reg/NET0131 ,
		\WX7334_reg/NET0131 ,
		_w2618_
	);
	LUT2 #(
		.INIT('h1)
	) name1111 (
		_w2617_,
		_w2618_,
		_w2619_
	);
	LUT2 #(
		.INIT('h2)
	) name1112 (
		\WX7142_reg/NET0131 ,
		\WX7206_reg/NET0131 ,
		_w2620_
	);
	LUT2 #(
		.INIT('h4)
	) name1113 (
		\WX7142_reg/NET0131 ,
		\WX7206_reg/NET0131 ,
		_w2621_
	);
	LUT2 #(
		.INIT('h1)
	) name1114 (
		_w2620_,
		_w2621_,
		_w2622_
	);
	LUT2 #(
		.INIT('h4)
	) name1115 (
		_w2619_,
		_w2622_,
		_w2623_
	);
	LUT2 #(
		.INIT('h2)
	) name1116 (
		_w2619_,
		_w2622_,
		_w2624_
	);
	LUT2 #(
		.INIT('h1)
	) name1117 (
		\TM0_pad ,
		_w2623_,
		_w2625_
	);
	LUT2 #(
		.INIT('h4)
	) name1118 (
		_w2624_,
		_w2625_,
		_w2626_
	);
	LUT2 #(
		.INIT('h2)
	) name1119 (
		_w1976_,
		_w2616_,
		_w2627_
	);
	LUT2 #(
		.INIT('h4)
	) name1120 (
		_w2626_,
		_w2627_,
		_w2628_
	);
	LUT2 #(
		.INIT('h1)
	) name1121 (
		_w2615_,
		_w2628_,
		_w2629_
	);
	LUT2 #(
		.INIT('h8)
	) name1122 (
		\TM0_pad ,
		\_2253__reg/NET0131 ,
		_w2630_
	);
	LUT2 #(
		.INIT('h2)
	) name1123 (
		\WX8561_reg/NET0131 ,
		\WX8625_reg/NET0131 ,
		_w2631_
	);
	LUT2 #(
		.INIT('h4)
	) name1124 (
		\WX8561_reg/NET0131 ,
		\WX8625_reg/NET0131 ,
		_w2632_
	);
	LUT2 #(
		.INIT('h1)
	) name1125 (
		_w2631_,
		_w2632_,
		_w2633_
	);
	LUT2 #(
		.INIT('h2)
	) name1126 (
		\WX8497_reg/NET0131 ,
		_w2633_,
		_w2634_
	);
	LUT2 #(
		.INIT('h4)
	) name1127 (
		\WX8497_reg/NET0131 ,
		_w2633_,
		_w2635_
	);
	LUT2 #(
		.INIT('h1)
	) name1128 (
		_w2634_,
		_w2635_,
		_w2636_
	);
	LUT2 #(
		.INIT('h2)
	) name1129 (
		\TM1_pad ,
		\WX8433_reg/NET0131 ,
		_w2637_
	);
	LUT2 #(
		.INIT('h4)
	) name1130 (
		\TM1_pad ,
		\WX8433_reg/NET0131 ,
		_w2638_
	);
	LUT2 #(
		.INIT('h1)
	) name1131 (
		_w2637_,
		_w2638_,
		_w2639_
	);
	LUT2 #(
		.INIT('h4)
	) name1132 (
		_w2636_,
		_w2639_,
		_w2640_
	);
	LUT2 #(
		.INIT('h2)
	) name1133 (
		_w2636_,
		_w2639_,
		_w2641_
	);
	LUT2 #(
		.INIT('h1)
	) name1134 (
		\TM0_pad ,
		_w2640_,
		_w2642_
	);
	LUT2 #(
		.INIT('h4)
	) name1135 (
		_w2641_,
		_w2642_,
		_w2643_
	);
	LUT2 #(
		.INIT('h1)
	) name1136 (
		_w2630_,
		_w2643_,
		_w2644_
	);
	LUT2 #(
		.INIT('h2)
	) name1137 (
		_w1976_,
		_w2644_,
		_w2645_
	);
	LUT2 #(
		.INIT('h1)
	) name1138 (
		_w1605_,
		_w2452_,
		_w2646_
	);
	LUT2 #(
		.INIT('h2)
	) name1139 (
		_w1973_,
		_w2646_,
		_w2647_
	);
	LUT2 #(
		.INIT('h1)
	) name1140 (
		_w2645_,
		_w2647_,
		_w2648_
	);
	LUT2 #(
		.INIT('h1)
	) name1141 (
		\TM0_pad ,
		_w1787_,
		_w2649_
	);
	LUT2 #(
		.INIT('h1)
	) name1142 (
		_w1778_,
		_w2649_,
		_w2650_
	);
	LUT2 #(
		.INIT('h2)
	) name1143 (
		_w1973_,
		_w2650_,
		_w2651_
	);
	LUT2 #(
		.INIT('h8)
	) name1144 (
		\TM0_pad ,
		\_2103__reg/NET0131 ,
		_w2652_
	);
	LUT2 #(
		.INIT('h2)
	) name1145 (
		\WX2076_reg/NET0131 ,
		\WX2140_reg/NET0131 ,
		_w2653_
	);
	LUT2 #(
		.INIT('h4)
	) name1146 (
		\WX2076_reg/NET0131 ,
		\WX2140_reg/NET0131 ,
		_w2654_
	);
	LUT2 #(
		.INIT('h1)
	) name1147 (
		_w2653_,
		_w2654_,
		_w2655_
	);
	LUT2 #(
		.INIT('h2)
	) name1148 (
		\WX2012_reg/NET0131 ,
		_w2655_,
		_w2656_
	);
	LUT2 #(
		.INIT('h4)
	) name1149 (
		\WX2012_reg/NET0131 ,
		_w2655_,
		_w2657_
	);
	LUT2 #(
		.INIT('h1)
	) name1150 (
		_w2656_,
		_w2657_,
		_w2658_
	);
	LUT2 #(
		.INIT('h2)
	) name1151 (
		\TM1_pad ,
		\WX1948_reg/NET0131 ,
		_w2659_
	);
	LUT2 #(
		.INIT('h4)
	) name1152 (
		\TM1_pad ,
		\WX1948_reg/NET0131 ,
		_w2660_
	);
	LUT2 #(
		.INIT('h1)
	) name1153 (
		_w2659_,
		_w2660_,
		_w2661_
	);
	LUT2 #(
		.INIT('h4)
	) name1154 (
		_w2658_,
		_w2661_,
		_w2662_
	);
	LUT2 #(
		.INIT('h2)
	) name1155 (
		_w2658_,
		_w2661_,
		_w2663_
	);
	LUT2 #(
		.INIT('h1)
	) name1156 (
		\TM0_pad ,
		_w2662_,
		_w2664_
	);
	LUT2 #(
		.INIT('h4)
	) name1157 (
		_w2663_,
		_w2664_,
		_w2665_
	);
	LUT2 #(
		.INIT('h1)
	) name1158 (
		_w2652_,
		_w2665_,
		_w2666_
	);
	LUT2 #(
		.INIT('h2)
	) name1159 (
		_w1976_,
		_w2666_,
		_w2667_
	);
	LUT2 #(
		.INIT('h1)
	) name1160 (
		_w2651_,
		_w2667_,
		_w2668_
	);
	LUT2 #(
		.INIT('h1)
	) name1161 (
		_w1810_,
		_w2019_,
		_w2669_
	);
	LUT2 #(
		.INIT('h2)
	) name1162 (
		_w1973_,
		_w2669_,
		_w2670_
	);
	LUT2 #(
		.INIT('h1)
	) name1163 (
		\DATA_0_28_pad ,
		\TM0_pad ,
		_w2671_
	);
	LUT2 #(
		.INIT('h2)
	) name1164 (
		\TM0_pad ,
		\_2361__reg/NET0131 ,
		_w2672_
	);
	LUT2 #(
		.INIT('h2)
	) name1165 (
		_w1976_,
		_w2671_,
		_w2673_
	);
	LUT2 #(
		.INIT('h4)
	) name1166 (
		_w2672_,
		_w2673_,
		_w2674_
	);
	LUT2 #(
		.INIT('h1)
	) name1167 (
		_w2670_,
		_w2674_,
		_w2675_
	);
	LUT2 #(
		.INIT('h8)
	) name1168 (
		RESET_pad,
		\WX10833_reg/NET0131 ,
		_w2676_
	);
	LUT2 #(
		.INIT('h4)
	) name1169 (
		_w1547_,
		_w1973_,
		_w2677_
	);
	LUT2 #(
		.INIT('h2)
	) name1170 (
		\WX3397_reg/NET0131 ,
		\WX3461_reg/NET0131 ,
		_w2678_
	);
	LUT2 #(
		.INIT('h4)
	) name1171 (
		\WX3397_reg/NET0131 ,
		\WX3461_reg/NET0131 ,
		_w2679_
	);
	LUT2 #(
		.INIT('h1)
	) name1172 (
		_w2678_,
		_w2679_,
		_w2680_
	);
	LUT2 #(
		.INIT('h2)
	) name1173 (
		\WX3269_reg/NET0131 ,
		\WX3333_reg/NET0131 ,
		_w2681_
	);
	LUT2 #(
		.INIT('h4)
	) name1174 (
		\WX3269_reg/NET0131 ,
		\WX3333_reg/NET0131 ,
		_w2682_
	);
	LUT2 #(
		.INIT('h1)
	) name1175 (
		_w2681_,
		_w2682_,
		_w2683_
	);
	LUT2 #(
		.INIT('h4)
	) name1176 (
		_w2680_,
		_w2683_,
		_w2684_
	);
	LUT2 #(
		.INIT('h2)
	) name1177 (
		_w2680_,
		_w2683_,
		_w2685_
	);
	LUT2 #(
		.INIT('h1)
	) name1178 (
		\TM0_pad ,
		_w2684_,
		_w2686_
	);
	LUT2 #(
		.INIT('h4)
	) name1179 (
		_w2685_,
		_w2686_,
		_w2687_
	);
	LUT2 #(
		.INIT('h2)
	) name1180 (
		_w2677_,
		_w2687_,
		_w2688_
	);
	LUT2 #(
		.INIT('h2)
	) name1181 (
		\TM0_pad ,
		\_2153__reg/NET0131 ,
		_w2689_
	);
	LUT2 #(
		.INIT('h2)
	) name1182 (
		\WX4690_reg/NET0131 ,
		\WX4754_reg/NET0131 ,
		_w2690_
	);
	LUT2 #(
		.INIT('h4)
	) name1183 (
		\WX4690_reg/NET0131 ,
		\WX4754_reg/NET0131 ,
		_w2691_
	);
	LUT2 #(
		.INIT('h1)
	) name1184 (
		_w2690_,
		_w2691_,
		_w2692_
	);
	LUT2 #(
		.INIT('h2)
	) name1185 (
		\WX4562_reg/NET0131 ,
		\WX4626_reg/NET0131 ,
		_w2693_
	);
	LUT2 #(
		.INIT('h4)
	) name1186 (
		\WX4562_reg/NET0131 ,
		\WX4626_reg/NET0131 ,
		_w2694_
	);
	LUT2 #(
		.INIT('h1)
	) name1187 (
		_w2693_,
		_w2694_,
		_w2695_
	);
	LUT2 #(
		.INIT('h4)
	) name1188 (
		_w2692_,
		_w2695_,
		_w2696_
	);
	LUT2 #(
		.INIT('h2)
	) name1189 (
		_w2692_,
		_w2695_,
		_w2697_
	);
	LUT2 #(
		.INIT('h1)
	) name1190 (
		\TM0_pad ,
		_w2696_,
		_w2698_
	);
	LUT2 #(
		.INIT('h4)
	) name1191 (
		_w2697_,
		_w2698_,
		_w2699_
	);
	LUT2 #(
		.INIT('h2)
	) name1192 (
		_w1976_,
		_w2689_,
		_w2700_
	);
	LUT2 #(
		.INIT('h4)
	) name1193 (
		_w2699_,
		_w2700_,
		_w2701_
	);
	LUT2 #(
		.INIT('h1)
	) name1194 (
		_w2688_,
		_w2701_,
		_w2702_
	);
	LUT2 #(
		.INIT('h8)
	) name1195 (
		\TM0_pad ,
		\_2285__reg/NET0131 ,
		_w2703_
	);
	LUT2 #(
		.INIT('h2)
	) name1196 (
		\WX9854_reg/NET0131 ,
		\WX9918_reg/NET0131 ,
		_w2704_
	);
	LUT2 #(
		.INIT('h4)
	) name1197 (
		\WX9854_reg/NET0131 ,
		\WX9918_reg/NET0131 ,
		_w2705_
	);
	LUT2 #(
		.INIT('h1)
	) name1198 (
		_w2704_,
		_w2705_,
		_w2706_
	);
	LUT2 #(
		.INIT('h2)
	) name1199 (
		\WX9790_reg/NET0131 ,
		_w2706_,
		_w2707_
	);
	LUT2 #(
		.INIT('h4)
	) name1200 (
		\WX9790_reg/NET0131 ,
		_w2706_,
		_w2708_
	);
	LUT2 #(
		.INIT('h1)
	) name1201 (
		_w2707_,
		_w2708_,
		_w2709_
	);
	LUT2 #(
		.INIT('h2)
	) name1202 (
		\TM1_pad ,
		\WX9726_reg/NET0131 ,
		_w2710_
	);
	LUT2 #(
		.INIT('h4)
	) name1203 (
		\TM1_pad ,
		\WX9726_reg/NET0131 ,
		_w2711_
	);
	LUT2 #(
		.INIT('h1)
	) name1204 (
		_w2710_,
		_w2711_,
		_w2712_
	);
	LUT2 #(
		.INIT('h4)
	) name1205 (
		_w2709_,
		_w2712_,
		_w2713_
	);
	LUT2 #(
		.INIT('h2)
	) name1206 (
		_w2709_,
		_w2712_,
		_w2714_
	);
	LUT2 #(
		.INIT('h1)
	) name1207 (
		\TM0_pad ,
		_w2713_,
		_w2715_
	);
	LUT2 #(
		.INIT('h4)
	) name1208 (
		_w2714_,
		_w2715_,
		_w2716_
	);
	LUT2 #(
		.INIT('h1)
	) name1209 (
		_w2703_,
		_w2716_,
		_w2717_
	);
	LUT2 #(
		.INIT('h2)
	) name1210 (
		_w1976_,
		_w2717_,
		_w2718_
	);
	LUT2 #(
		.INIT('h1)
	) name1211 (
		_w1605_,
		_w2643_,
		_w2719_
	);
	LUT2 #(
		.INIT('h2)
	) name1212 (
		_w1973_,
		_w2719_,
		_w2720_
	);
	LUT2 #(
		.INIT('h1)
	) name1213 (
		_w2718_,
		_w2720_,
		_w2721_
	);
	LUT2 #(
		.INIT('h8)
	) name1214 (
		\TM0_pad ,
		\_2136__reg/NET0131 ,
		_w2722_
	);
	LUT2 #(
		.INIT('h2)
	) name1215 (
		\WX3367_reg/NET0131 ,
		\WX3431_reg/NET0131 ,
		_w2723_
	);
	LUT2 #(
		.INIT('h4)
	) name1216 (
		\WX3367_reg/NET0131 ,
		\WX3431_reg/NET0131 ,
		_w2724_
	);
	LUT2 #(
		.INIT('h1)
	) name1217 (
		_w2723_,
		_w2724_,
		_w2725_
	);
	LUT2 #(
		.INIT('h2)
	) name1218 (
		\WX3303_reg/NET0131 ,
		_w2725_,
		_w2726_
	);
	LUT2 #(
		.INIT('h4)
	) name1219 (
		\WX3303_reg/NET0131 ,
		_w2725_,
		_w2727_
	);
	LUT2 #(
		.INIT('h1)
	) name1220 (
		_w2726_,
		_w2727_,
		_w2728_
	);
	LUT2 #(
		.INIT('h2)
	) name1221 (
		\TM1_pad ,
		\WX3239_reg/NET0131 ,
		_w2729_
	);
	LUT2 #(
		.INIT('h4)
	) name1222 (
		\TM1_pad ,
		\WX3239_reg/NET0131 ,
		_w2730_
	);
	LUT2 #(
		.INIT('h1)
	) name1223 (
		_w2729_,
		_w2730_,
		_w2731_
	);
	LUT2 #(
		.INIT('h4)
	) name1224 (
		_w2728_,
		_w2731_,
		_w2732_
	);
	LUT2 #(
		.INIT('h2)
	) name1225 (
		_w2728_,
		_w2731_,
		_w2733_
	);
	LUT2 #(
		.INIT('h1)
	) name1226 (
		\TM0_pad ,
		_w2732_,
		_w2734_
	);
	LUT2 #(
		.INIT('h4)
	) name1227 (
		_w2733_,
		_w2734_,
		_w2735_
	);
	LUT2 #(
		.INIT('h1)
	) name1228 (
		_w2722_,
		_w2735_,
		_w2736_
	);
	LUT2 #(
		.INIT('h2)
	) name1229 (
		_w1976_,
		_w2736_,
		_w2737_
	);
	LUT2 #(
		.INIT('h1)
	) name1230 (
		_w1794_,
		_w2493_,
		_w2738_
	);
	LUT2 #(
		.INIT('h2)
	) name1231 (
		_w1973_,
		_w2738_,
		_w2739_
	);
	LUT2 #(
		.INIT('h1)
	) name1232 (
		_w2737_,
		_w2739_,
		_w2740_
	);
	LUT2 #(
		.INIT('h8)
	) name1233 (
		\TM0_pad ,
		\_2318__reg/NET0131 ,
		_w2741_
	);
	LUT2 #(
		.INIT('h2)
	) name1234 (
		\WX11145_reg/NET0131 ,
		\WX11209_reg/NET0131 ,
		_w2742_
	);
	LUT2 #(
		.INIT('h4)
	) name1235 (
		\WX11145_reg/NET0131 ,
		\WX11209_reg/NET0131 ,
		_w2743_
	);
	LUT2 #(
		.INIT('h1)
	) name1236 (
		_w2742_,
		_w2743_,
		_w2744_
	);
	LUT2 #(
		.INIT('h2)
	) name1237 (
		\WX11081_reg/NET0131 ,
		_w2744_,
		_w2745_
	);
	LUT2 #(
		.INIT('h4)
	) name1238 (
		\WX11081_reg/NET0131 ,
		_w2744_,
		_w2746_
	);
	LUT2 #(
		.INIT('h1)
	) name1239 (
		_w2745_,
		_w2746_,
		_w2747_
	);
	LUT2 #(
		.INIT('h2)
	) name1240 (
		\TM1_pad ,
		\WX11017_reg/NET0131 ,
		_w2748_
	);
	LUT2 #(
		.INIT('h4)
	) name1241 (
		\TM1_pad ,
		\WX11017_reg/NET0131 ,
		_w2749_
	);
	LUT2 #(
		.INIT('h1)
	) name1242 (
		_w2748_,
		_w2749_,
		_w2750_
	);
	LUT2 #(
		.INIT('h4)
	) name1243 (
		_w2747_,
		_w2750_,
		_w2751_
	);
	LUT2 #(
		.INIT('h2)
	) name1244 (
		_w2747_,
		_w2750_,
		_w2752_
	);
	LUT2 #(
		.INIT('h1)
	) name1245 (
		\TM0_pad ,
		_w2751_,
		_w2753_
	);
	LUT2 #(
		.INIT('h4)
	) name1246 (
		_w2752_,
		_w2753_,
		_w2754_
	);
	LUT2 #(
		.INIT('h1)
	) name1247 (
		_w2741_,
		_w2754_,
		_w2755_
	);
	LUT2 #(
		.INIT('h2)
	) name1248 (
		_w1976_,
		_w2755_,
		_w2756_
	);
	LUT2 #(
		.INIT('h1)
	) name1249 (
		_w1621_,
		_w2556_,
		_w2757_
	);
	LUT2 #(
		.INIT('h2)
	) name1250 (
		_w1973_,
		_w2757_,
		_w2758_
	);
	LUT2 #(
		.INIT('h1)
	) name1251 (
		_w2756_,
		_w2758_,
		_w2759_
	);
	LUT2 #(
		.INIT('h2)
	) name1252 (
		_w2040_,
		_w2539_,
		_w2760_
	);
	LUT2 #(
		.INIT('h2)
	) name1253 (
		\TM0_pad ,
		\_2186__reg/NET0131 ,
		_w2761_
	);
	LUT2 #(
		.INIT('h2)
	) name1254 (
		\WX5981_reg/NET0131 ,
		\WX6045_reg/NET0131 ,
		_w2762_
	);
	LUT2 #(
		.INIT('h4)
	) name1255 (
		\WX5981_reg/NET0131 ,
		\WX6045_reg/NET0131 ,
		_w2763_
	);
	LUT2 #(
		.INIT('h1)
	) name1256 (
		_w2762_,
		_w2763_,
		_w2764_
	);
	LUT2 #(
		.INIT('h2)
	) name1257 (
		\WX5853_reg/NET0131 ,
		\WX5917_reg/NET0131 ,
		_w2765_
	);
	LUT2 #(
		.INIT('h4)
	) name1258 (
		\WX5853_reg/NET0131 ,
		\WX5917_reg/NET0131 ,
		_w2766_
	);
	LUT2 #(
		.INIT('h1)
	) name1259 (
		_w2765_,
		_w2766_,
		_w2767_
	);
	LUT2 #(
		.INIT('h4)
	) name1260 (
		_w2764_,
		_w2767_,
		_w2768_
	);
	LUT2 #(
		.INIT('h2)
	) name1261 (
		_w2764_,
		_w2767_,
		_w2769_
	);
	LUT2 #(
		.INIT('h1)
	) name1262 (
		\TM0_pad ,
		_w2768_,
		_w2770_
	);
	LUT2 #(
		.INIT('h4)
	) name1263 (
		_w2769_,
		_w2770_,
		_w2771_
	);
	LUT2 #(
		.INIT('h2)
	) name1264 (
		_w1976_,
		_w2761_,
		_w2772_
	);
	LUT2 #(
		.INIT('h4)
	) name1265 (
		_w2771_,
		_w2772_,
		_w2773_
	);
	LUT2 #(
		.INIT('h1)
	) name1266 (
		_w2760_,
		_w2773_,
		_w2774_
	);
	LUT2 #(
		.INIT('h2)
	) name1267 (
		_w2341_,
		_w2611_,
		_w2775_
	);
	LUT2 #(
		.INIT('h2)
	) name1268 (
		\TM0_pad ,
		\_2219__reg/NET0131 ,
		_w2776_
	);
	LUT2 #(
		.INIT('h2)
	) name1269 (
		\WX7272_reg/NET0131 ,
		\WX7336_reg/NET0131 ,
		_w2777_
	);
	LUT2 #(
		.INIT('h4)
	) name1270 (
		\WX7272_reg/NET0131 ,
		\WX7336_reg/NET0131 ,
		_w2778_
	);
	LUT2 #(
		.INIT('h1)
	) name1271 (
		_w2777_,
		_w2778_,
		_w2779_
	);
	LUT2 #(
		.INIT('h2)
	) name1272 (
		\WX7144_reg/NET0131 ,
		\WX7208_reg/NET0131 ,
		_w2780_
	);
	LUT2 #(
		.INIT('h4)
	) name1273 (
		\WX7144_reg/NET0131 ,
		\WX7208_reg/NET0131 ,
		_w2781_
	);
	LUT2 #(
		.INIT('h1)
	) name1274 (
		_w2780_,
		_w2781_,
		_w2782_
	);
	LUT2 #(
		.INIT('h4)
	) name1275 (
		_w2779_,
		_w2782_,
		_w2783_
	);
	LUT2 #(
		.INIT('h2)
	) name1276 (
		_w2779_,
		_w2782_,
		_w2784_
	);
	LUT2 #(
		.INIT('h1)
	) name1277 (
		\TM0_pad ,
		_w2783_,
		_w2785_
	);
	LUT2 #(
		.INIT('h4)
	) name1278 (
		_w2784_,
		_w2785_,
		_w2786_
	);
	LUT2 #(
		.INIT('h2)
	) name1279 (
		_w1976_,
		_w2776_,
		_w2787_
	);
	LUT2 #(
		.INIT('h4)
	) name1280 (
		_w2786_,
		_w2787_,
		_w2788_
	);
	LUT2 #(
		.INIT('h1)
	) name1281 (
		_w2775_,
		_w2788_,
		_w2789_
	);
	LUT2 #(
		.INIT('h2)
	) name1282 (
		_w1974_,
		_w2626_,
		_w2790_
	);
	LUT2 #(
		.INIT('h2)
	) name1283 (
		\TM0_pad ,
		\_2252__reg/NET0131 ,
		_w2791_
	);
	LUT2 #(
		.INIT('h2)
	) name1284 (
		\WX8563_reg/NET0131 ,
		\WX8627_reg/NET0131 ,
		_w2792_
	);
	LUT2 #(
		.INIT('h4)
	) name1285 (
		\WX8563_reg/NET0131 ,
		\WX8627_reg/NET0131 ,
		_w2793_
	);
	LUT2 #(
		.INIT('h1)
	) name1286 (
		_w2792_,
		_w2793_,
		_w2794_
	);
	LUT2 #(
		.INIT('h2)
	) name1287 (
		\WX8435_reg/NET0131 ,
		\WX8499_reg/NET0131 ,
		_w2795_
	);
	LUT2 #(
		.INIT('h4)
	) name1288 (
		\WX8435_reg/NET0131 ,
		\WX8499_reg/NET0131 ,
		_w2796_
	);
	LUT2 #(
		.INIT('h1)
	) name1289 (
		_w2795_,
		_w2796_,
		_w2797_
	);
	LUT2 #(
		.INIT('h4)
	) name1290 (
		_w2794_,
		_w2797_,
		_w2798_
	);
	LUT2 #(
		.INIT('h2)
	) name1291 (
		_w2794_,
		_w2797_,
		_w2799_
	);
	LUT2 #(
		.INIT('h1)
	) name1292 (
		\TM0_pad ,
		_w2798_,
		_w2800_
	);
	LUT2 #(
		.INIT('h4)
	) name1293 (
		_w2799_,
		_w2800_,
		_w2801_
	);
	LUT2 #(
		.INIT('h2)
	) name1294 (
		_w1976_,
		_w2791_,
		_w2802_
	);
	LUT2 #(
		.INIT('h4)
	) name1295 (
		_w2801_,
		_w2802_,
		_w2803_
	);
	LUT2 #(
		.INIT('h1)
	) name1296 (
		_w2790_,
		_w2803_,
		_w2804_
	);
	LUT2 #(
		.INIT('h1)
	) name1297 (
		\TM0_pad ,
		_w1771_,
		_w2805_
	);
	LUT2 #(
		.INIT('h1)
	) name1298 (
		_w1762_,
		_w2805_,
		_w2806_
	);
	LUT2 #(
		.INIT('h2)
	) name1299 (
		_w1973_,
		_w2806_,
		_w2807_
	);
	LUT2 #(
		.INIT('h8)
	) name1300 (
		\TM0_pad ,
		\_2102__reg/NET0131 ,
		_w2808_
	);
	LUT2 #(
		.INIT('h2)
	) name1301 (
		\WX2078_reg/NET0131 ,
		\WX2142_reg/NET0131 ,
		_w2809_
	);
	LUT2 #(
		.INIT('h4)
	) name1302 (
		\WX2078_reg/NET0131 ,
		\WX2142_reg/NET0131 ,
		_w2810_
	);
	LUT2 #(
		.INIT('h1)
	) name1303 (
		_w2809_,
		_w2810_,
		_w2811_
	);
	LUT2 #(
		.INIT('h2)
	) name1304 (
		\WX2014_reg/NET0131 ,
		_w2811_,
		_w2812_
	);
	LUT2 #(
		.INIT('h4)
	) name1305 (
		\WX2014_reg/NET0131 ,
		_w2811_,
		_w2813_
	);
	LUT2 #(
		.INIT('h1)
	) name1306 (
		_w2812_,
		_w2813_,
		_w2814_
	);
	LUT2 #(
		.INIT('h2)
	) name1307 (
		\TM1_pad ,
		\WX1950_reg/NET0131 ,
		_w2815_
	);
	LUT2 #(
		.INIT('h4)
	) name1308 (
		\TM1_pad ,
		\WX1950_reg/NET0131 ,
		_w2816_
	);
	LUT2 #(
		.INIT('h1)
	) name1309 (
		_w2815_,
		_w2816_,
		_w2817_
	);
	LUT2 #(
		.INIT('h4)
	) name1310 (
		_w2814_,
		_w2817_,
		_w2818_
	);
	LUT2 #(
		.INIT('h2)
	) name1311 (
		_w2814_,
		_w2817_,
		_w2819_
	);
	LUT2 #(
		.INIT('h1)
	) name1312 (
		\TM0_pad ,
		_w2818_,
		_w2820_
	);
	LUT2 #(
		.INIT('h4)
	) name1313 (
		_w2819_,
		_w2820_,
		_w2821_
	);
	LUT2 #(
		.INIT('h1)
	) name1314 (
		_w2808_,
		_w2821_,
		_w2822_
	);
	LUT2 #(
		.INIT('h2)
	) name1315 (
		_w1976_,
		_w2822_,
		_w2823_
	);
	LUT2 #(
		.INIT('h1)
	) name1316 (
		_w2807_,
		_w2823_,
		_w2824_
	);
	LUT2 #(
		.INIT('h2)
	) name1317 (
		\WX11125_reg/NET0131 ,
		\WX11189_reg/NET0131 ,
		_w2825_
	);
	LUT2 #(
		.INIT('h4)
	) name1318 (
		\WX11125_reg/NET0131 ,
		\WX11189_reg/NET0131 ,
		_w2826_
	);
	LUT2 #(
		.INIT('h1)
	) name1319 (
		_w2825_,
		_w2826_,
		_w2827_
	);
	LUT2 #(
		.INIT('h2)
	) name1320 (
		\WX11061_reg/NET0131 ,
		_w2827_,
		_w2828_
	);
	LUT2 #(
		.INIT('h4)
	) name1321 (
		\WX11061_reg/NET0131 ,
		_w2827_,
		_w2829_
	);
	LUT2 #(
		.INIT('h1)
	) name1322 (
		_w2828_,
		_w2829_,
		_w2830_
	);
	LUT2 #(
		.INIT('h2)
	) name1323 (
		\TM1_pad ,
		\WX10997_reg/NET0131 ,
		_w2831_
	);
	LUT2 #(
		.INIT('h4)
	) name1324 (
		\TM1_pad ,
		\WX10997_reg/NET0131 ,
		_w2832_
	);
	LUT2 #(
		.INIT('h1)
	) name1325 (
		_w2831_,
		_w2832_,
		_w2833_
	);
	LUT2 #(
		.INIT('h4)
	) name1326 (
		_w2830_,
		_w2833_,
		_w2834_
	);
	LUT2 #(
		.INIT('h2)
	) name1327 (
		_w2830_,
		_w2833_,
		_w2835_
	);
	LUT2 #(
		.INIT('h1)
	) name1328 (
		\TM0_pad ,
		_w2834_,
		_w2836_
	);
	LUT2 #(
		.INIT('h4)
	) name1329 (
		_w2835_,
		_w2836_,
		_w2837_
	);
	LUT2 #(
		.INIT('h1)
	) name1330 (
		_w1794_,
		_w2837_,
		_w2838_
	);
	LUT2 #(
		.INIT('h2)
	) name1331 (
		_w1973_,
		_w2838_,
		_w2839_
	);
	LUT2 #(
		.INIT('h1)
	) name1332 (
		\DATA_0_27_pad ,
		\TM0_pad ,
		_w2840_
	);
	LUT2 #(
		.INIT('h2)
	) name1333 (
		\TM0_pad ,
		\_2360__reg/NET0131 ,
		_w2841_
	);
	LUT2 #(
		.INIT('h2)
	) name1334 (
		_w1976_,
		_w2840_,
		_w2842_
	);
	LUT2 #(
		.INIT('h4)
	) name1335 (
		_w2841_,
		_w2842_,
		_w2843_
	);
	LUT2 #(
		.INIT('h1)
	) name1336 (
		_w2839_,
		_w2843_,
		_w2844_
	);
	LUT2 #(
		.INIT('h8)
	) name1337 (
		RESET_pad,
		\WX10835_reg/NET0131 ,
		_w2845_
	);
	LUT2 #(
		.INIT('h4)
	) name1338 (
		_w1534_,
		_w1973_,
		_w2846_
	);
	LUT2 #(
		.INIT('h2)
	) name1339 (
		\WX3399_reg/NET0131 ,
		\WX3463_reg/NET0131 ,
		_w2847_
	);
	LUT2 #(
		.INIT('h4)
	) name1340 (
		\WX3399_reg/NET0131 ,
		\WX3463_reg/NET0131 ,
		_w2848_
	);
	LUT2 #(
		.INIT('h1)
	) name1341 (
		_w2847_,
		_w2848_,
		_w2849_
	);
	LUT2 #(
		.INIT('h2)
	) name1342 (
		\WX3271_reg/NET0131 ,
		\WX3335_reg/NET0131 ,
		_w2850_
	);
	LUT2 #(
		.INIT('h4)
	) name1343 (
		\WX3271_reg/NET0131 ,
		\WX3335_reg/NET0131 ,
		_w2851_
	);
	LUT2 #(
		.INIT('h1)
	) name1344 (
		_w2850_,
		_w2851_,
		_w2852_
	);
	LUT2 #(
		.INIT('h4)
	) name1345 (
		_w2849_,
		_w2852_,
		_w2853_
	);
	LUT2 #(
		.INIT('h2)
	) name1346 (
		_w2849_,
		_w2852_,
		_w2854_
	);
	LUT2 #(
		.INIT('h1)
	) name1347 (
		\TM0_pad ,
		_w2853_,
		_w2855_
	);
	LUT2 #(
		.INIT('h4)
	) name1348 (
		_w2854_,
		_w2855_,
		_w2856_
	);
	LUT2 #(
		.INIT('h2)
	) name1349 (
		_w2846_,
		_w2856_,
		_w2857_
	);
	LUT2 #(
		.INIT('h2)
	) name1350 (
		\TM0_pad ,
		\_2152__reg/NET0131 ,
		_w2858_
	);
	LUT2 #(
		.INIT('h2)
	) name1351 (
		\WX4692_reg/NET0131 ,
		\WX4756_reg/NET0131 ,
		_w2859_
	);
	LUT2 #(
		.INIT('h4)
	) name1352 (
		\WX4692_reg/NET0131 ,
		\WX4756_reg/NET0131 ,
		_w2860_
	);
	LUT2 #(
		.INIT('h1)
	) name1353 (
		_w2859_,
		_w2860_,
		_w2861_
	);
	LUT2 #(
		.INIT('h2)
	) name1354 (
		\WX4564_reg/NET0131 ,
		\WX4628_reg/NET0131 ,
		_w2862_
	);
	LUT2 #(
		.INIT('h4)
	) name1355 (
		\WX4564_reg/NET0131 ,
		\WX4628_reg/NET0131 ,
		_w2863_
	);
	LUT2 #(
		.INIT('h1)
	) name1356 (
		_w2862_,
		_w2863_,
		_w2864_
	);
	LUT2 #(
		.INIT('h4)
	) name1357 (
		_w2861_,
		_w2864_,
		_w2865_
	);
	LUT2 #(
		.INIT('h2)
	) name1358 (
		_w2861_,
		_w2864_,
		_w2866_
	);
	LUT2 #(
		.INIT('h1)
	) name1359 (
		\TM0_pad ,
		_w2865_,
		_w2867_
	);
	LUT2 #(
		.INIT('h4)
	) name1360 (
		_w2866_,
		_w2867_,
		_w2868_
	);
	LUT2 #(
		.INIT('h2)
	) name1361 (
		_w1976_,
		_w2858_,
		_w2869_
	);
	LUT2 #(
		.INIT('h4)
	) name1362 (
		_w2868_,
		_w2869_,
		_w2870_
	);
	LUT2 #(
		.INIT('h1)
	) name1363 (
		_w2857_,
		_w2870_,
		_w2871_
	);
	LUT2 #(
		.INIT('h2)
	) name1364 (
		_w1974_,
		_w2801_,
		_w2872_
	);
	LUT2 #(
		.INIT('h2)
	) name1365 (
		\TM0_pad ,
		\_2284__reg/NET0131 ,
		_w2873_
	);
	LUT2 #(
		.INIT('h2)
	) name1366 (
		\WX9856_reg/NET0131 ,
		\WX9920_reg/NET0131 ,
		_w2874_
	);
	LUT2 #(
		.INIT('h4)
	) name1367 (
		\WX9856_reg/NET0131 ,
		\WX9920_reg/NET0131 ,
		_w2875_
	);
	LUT2 #(
		.INIT('h1)
	) name1368 (
		_w2874_,
		_w2875_,
		_w2876_
	);
	LUT2 #(
		.INIT('h2)
	) name1369 (
		\WX9728_reg/NET0131 ,
		\WX9792_reg/NET0131 ,
		_w2877_
	);
	LUT2 #(
		.INIT('h4)
	) name1370 (
		\WX9728_reg/NET0131 ,
		\WX9792_reg/NET0131 ,
		_w2878_
	);
	LUT2 #(
		.INIT('h1)
	) name1371 (
		_w2877_,
		_w2878_,
		_w2879_
	);
	LUT2 #(
		.INIT('h4)
	) name1372 (
		_w2876_,
		_w2879_,
		_w2880_
	);
	LUT2 #(
		.INIT('h2)
	) name1373 (
		_w2876_,
		_w2879_,
		_w2881_
	);
	LUT2 #(
		.INIT('h1)
	) name1374 (
		\TM0_pad ,
		_w2880_,
		_w2882_
	);
	LUT2 #(
		.INIT('h4)
	) name1375 (
		_w2881_,
		_w2882_,
		_w2883_
	);
	LUT2 #(
		.INIT('h2)
	) name1376 (
		_w1976_,
		_w2873_,
		_w2884_
	);
	LUT2 #(
		.INIT('h4)
	) name1377 (
		_w2883_,
		_w2884_,
		_w2885_
	);
	LUT2 #(
		.INIT('h1)
	) name1378 (
		_w2872_,
		_w2885_,
		_w2886_
	);
	LUT2 #(
		.INIT('h8)
	) name1379 (
		\TM0_pad ,
		\_2135__reg/NET0131 ,
		_w2887_
	);
	LUT2 #(
		.INIT('h2)
	) name1380 (
		\WX3369_reg/NET0131 ,
		\WX3433_reg/NET0131 ,
		_w2888_
	);
	LUT2 #(
		.INIT('h4)
	) name1381 (
		\WX3369_reg/NET0131 ,
		\WX3433_reg/NET0131 ,
		_w2889_
	);
	LUT2 #(
		.INIT('h1)
	) name1382 (
		_w2888_,
		_w2889_,
		_w2890_
	);
	LUT2 #(
		.INIT('h2)
	) name1383 (
		\WX3305_reg/NET0131 ,
		_w2890_,
		_w2891_
	);
	LUT2 #(
		.INIT('h4)
	) name1384 (
		\WX3305_reg/NET0131 ,
		_w2890_,
		_w2892_
	);
	LUT2 #(
		.INIT('h1)
	) name1385 (
		_w2891_,
		_w2892_,
		_w2893_
	);
	LUT2 #(
		.INIT('h2)
	) name1386 (
		\TM1_pad ,
		\WX3241_reg/NET0131 ,
		_w2894_
	);
	LUT2 #(
		.INIT('h4)
	) name1387 (
		\TM1_pad ,
		\WX3241_reg/NET0131 ,
		_w2895_
	);
	LUT2 #(
		.INIT('h1)
	) name1388 (
		_w2894_,
		_w2895_,
		_w2896_
	);
	LUT2 #(
		.INIT('h4)
	) name1389 (
		_w2893_,
		_w2896_,
		_w2897_
	);
	LUT2 #(
		.INIT('h2)
	) name1390 (
		_w2893_,
		_w2896_,
		_w2898_
	);
	LUT2 #(
		.INIT('h1)
	) name1391 (
		\TM0_pad ,
		_w2897_,
		_w2899_
	);
	LUT2 #(
		.INIT('h4)
	) name1392 (
		_w2898_,
		_w2899_,
		_w2900_
	);
	LUT2 #(
		.INIT('h1)
	) name1393 (
		_w2887_,
		_w2900_,
		_w2901_
	);
	LUT2 #(
		.INIT('h2)
	) name1394 (
		_w1976_,
		_w2901_,
		_w2902_
	);
	LUT2 #(
		.INIT('h1)
	) name1395 (
		_w1778_,
		_w2665_,
		_w2903_
	);
	LUT2 #(
		.INIT('h2)
	) name1396 (
		_w1973_,
		_w2903_,
		_w2904_
	);
	LUT2 #(
		.INIT('h1)
	) name1397 (
		_w2902_,
		_w2904_,
		_w2905_
	);
	LUT2 #(
		.INIT('h8)
	) name1398 (
		\TM0_pad ,
		\_2317__reg/NET0131 ,
		_w2906_
	);
	LUT2 #(
		.INIT('h2)
	) name1399 (
		\WX11147_reg/NET0131 ,
		\WX11211_reg/NET0131 ,
		_w2907_
	);
	LUT2 #(
		.INIT('h4)
	) name1400 (
		\WX11147_reg/NET0131 ,
		\WX11211_reg/NET0131 ,
		_w2908_
	);
	LUT2 #(
		.INIT('h1)
	) name1401 (
		_w2907_,
		_w2908_,
		_w2909_
	);
	LUT2 #(
		.INIT('h2)
	) name1402 (
		\WX11083_reg/NET0131 ,
		_w2909_,
		_w2910_
	);
	LUT2 #(
		.INIT('h4)
	) name1403 (
		\WX11083_reg/NET0131 ,
		_w2909_,
		_w2911_
	);
	LUT2 #(
		.INIT('h1)
	) name1404 (
		_w2910_,
		_w2911_,
		_w2912_
	);
	LUT2 #(
		.INIT('h2)
	) name1405 (
		\TM1_pad ,
		\WX11019_reg/NET0131 ,
		_w2913_
	);
	LUT2 #(
		.INIT('h4)
	) name1406 (
		\TM1_pad ,
		\WX11019_reg/NET0131 ,
		_w2914_
	);
	LUT2 #(
		.INIT('h1)
	) name1407 (
		_w2913_,
		_w2914_,
		_w2915_
	);
	LUT2 #(
		.INIT('h4)
	) name1408 (
		_w2912_,
		_w2915_,
		_w2916_
	);
	LUT2 #(
		.INIT('h2)
	) name1409 (
		_w2912_,
		_w2915_,
		_w2917_
	);
	LUT2 #(
		.INIT('h1)
	) name1410 (
		\TM0_pad ,
		_w2916_,
		_w2918_
	);
	LUT2 #(
		.INIT('h4)
	) name1411 (
		_w2917_,
		_w2918_,
		_w2919_
	);
	LUT2 #(
		.INIT('h1)
	) name1412 (
		_w2906_,
		_w2919_,
		_w2920_
	);
	LUT2 #(
		.INIT('h2)
	) name1413 (
		_w1976_,
		_w2920_,
		_w2921_
	);
	LUT2 #(
		.INIT('h1)
	) name1414 (
		_w1605_,
		_w2716_,
		_w2922_
	);
	LUT2 #(
		.INIT('h2)
	) name1415 (
		_w1973_,
		_w2922_,
		_w2923_
	);
	LUT2 #(
		.INIT('h1)
	) name1416 (
		_w2921_,
		_w2923_,
		_w2924_
	);
	LUT2 #(
		.INIT('h2)
	) name1417 (
		_w2677_,
		_w2699_,
		_w2925_
	);
	LUT2 #(
		.INIT('h2)
	) name1418 (
		\TM0_pad ,
		\_2185__reg/NET0131 ,
		_w2926_
	);
	LUT2 #(
		.INIT('h2)
	) name1419 (
		\WX5983_reg/NET0131 ,
		\WX6047_reg/NET0131 ,
		_w2927_
	);
	LUT2 #(
		.INIT('h4)
	) name1420 (
		\WX5983_reg/NET0131 ,
		\WX6047_reg/NET0131 ,
		_w2928_
	);
	LUT2 #(
		.INIT('h1)
	) name1421 (
		_w2927_,
		_w2928_,
		_w2929_
	);
	LUT2 #(
		.INIT('h2)
	) name1422 (
		\WX5855_reg/NET0131 ,
		\WX5919_reg/NET0131 ,
		_w2930_
	);
	LUT2 #(
		.INIT('h4)
	) name1423 (
		\WX5855_reg/NET0131 ,
		\WX5919_reg/NET0131 ,
		_w2931_
	);
	LUT2 #(
		.INIT('h1)
	) name1424 (
		_w2930_,
		_w2931_,
		_w2932_
	);
	LUT2 #(
		.INIT('h4)
	) name1425 (
		_w2929_,
		_w2932_,
		_w2933_
	);
	LUT2 #(
		.INIT('h2)
	) name1426 (
		_w2929_,
		_w2932_,
		_w2934_
	);
	LUT2 #(
		.INIT('h1)
	) name1427 (
		\TM0_pad ,
		_w2933_,
		_w2935_
	);
	LUT2 #(
		.INIT('h4)
	) name1428 (
		_w2934_,
		_w2935_,
		_w2936_
	);
	LUT2 #(
		.INIT('h2)
	) name1429 (
		_w1976_,
		_w2926_,
		_w2937_
	);
	LUT2 #(
		.INIT('h4)
	) name1430 (
		_w2936_,
		_w2937_,
		_w2938_
	);
	LUT2 #(
		.INIT('h1)
	) name1431 (
		_w2925_,
		_w2938_,
		_w2939_
	);
	LUT2 #(
		.INIT('h2)
	) name1432 (
		_w2040_,
		_w2771_,
		_w2940_
	);
	LUT2 #(
		.INIT('h2)
	) name1433 (
		\TM0_pad ,
		\_2218__reg/NET0131 ,
		_w2941_
	);
	LUT2 #(
		.INIT('h2)
	) name1434 (
		\WX7274_reg/NET0131 ,
		\WX7338_reg/NET0131 ,
		_w2942_
	);
	LUT2 #(
		.INIT('h4)
	) name1435 (
		\WX7274_reg/NET0131 ,
		\WX7338_reg/NET0131 ,
		_w2943_
	);
	LUT2 #(
		.INIT('h1)
	) name1436 (
		_w2942_,
		_w2943_,
		_w2944_
	);
	LUT2 #(
		.INIT('h2)
	) name1437 (
		\WX7146_reg/NET0131 ,
		\WX7210_reg/NET0131 ,
		_w2945_
	);
	LUT2 #(
		.INIT('h4)
	) name1438 (
		\WX7146_reg/NET0131 ,
		\WX7210_reg/NET0131 ,
		_w2946_
	);
	LUT2 #(
		.INIT('h1)
	) name1439 (
		_w2945_,
		_w2946_,
		_w2947_
	);
	LUT2 #(
		.INIT('h4)
	) name1440 (
		_w2944_,
		_w2947_,
		_w2948_
	);
	LUT2 #(
		.INIT('h2)
	) name1441 (
		_w2944_,
		_w2947_,
		_w2949_
	);
	LUT2 #(
		.INIT('h1)
	) name1442 (
		\TM0_pad ,
		_w2948_,
		_w2950_
	);
	LUT2 #(
		.INIT('h4)
	) name1443 (
		_w2949_,
		_w2950_,
		_w2951_
	);
	LUT2 #(
		.INIT('h2)
	) name1444 (
		_w1976_,
		_w2941_,
		_w2952_
	);
	LUT2 #(
		.INIT('h4)
	) name1445 (
		_w2951_,
		_w2952_,
		_w2953_
	);
	LUT2 #(
		.INIT('h1)
	) name1446 (
		_w2940_,
		_w2953_,
		_w2954_
	);
	LUT2 #(
		.INIT('h2)
	) name1447 (
		_w2341_,
		_w2786_,
		_w2955_
	);
	LUT2 #(
		.INIT('h2)
	) name1448 (
		\TM0_pad ,
		\_2251__reg/NET0131 ,
		_w2956_
	);
	LUT2 #(
		.INIT('h2)
	) name1449 (
		\WX8565_reg/NET0131 ,
		\WX8629_reg/NET0131 ,
		_w2957_
	);
	LUT2 #(
		.INIT('h4)
	) name1450 (
		\WX8565_reg/NET0131 ,
		\WX8629_reg/NET0131 ,
		_w2958_
	);
	LUT2 #(
		.INIT('h1)
	) name1451 (
		_w2957_,
		_w2958_,
		_w2959_
	);
	LUT2 #(
		.INIT('h2)
	) name1452 (
		\WX8437_reg/NET0131 ,
		\WX8501_reg/NET0131 ,
		_w2960_
	);
	LUT2 #(
		.INIT('h4)
	) name1453 (
		\WX8437_reg/NET0131 ,
		\WX8501_reg/NET0131 ,
		_w2961_
	);
	LUT2 #(
		.INIT('h1)
	) name1454 (
		_w2960_,
		_w2961_,
		_w2962_
	);
	LUT2 #(
		.INIT('h4)
	) name1455 (
		_w2959_,
		_w2962_,
		_w2963_
	);
	LUT2 #(
		.INIT('h2)
	) name1456 (
		_w2959_,
		_w2962_,
		_w2964_
	);
	LUT2 #(
		.INIT('h1)
	) name1457 (
		\TM0_pad ,
		_w2963_,
		_w2965_
	);
	LUT2 #(
		.INIT('h4)
	) name1458 (
		_w2964_,
		_w2965_,
		_w2966_
	);
	LUT2 #(
		.INIT('h2)
	) name1459 (
		_w1976_,
		_w2956_,
		_w2967_
	);
	LUT2 #(
		.INIT('h4)
	) name1460 (
		_w2966_,
		_w2967_,
		_w2968_
	);
	LUT2 #(
		.INIT('h1)
	) name1461 (
		_w2955_,
		_w2968_,
		_w2969_
	);
	LUT2 #(
		.INIT('h1)
	) name1462 (
		\TM0_pad ,
		_w1755_,
		_w2970_
	);
	LUT2 #(
		.INIT('h1)
	) name1463 (
		_w1746_,
		_w2970_,
		_w2971_
	);
	LUT2 #(
		.INIT('h2)
	) name1464 (
		_w1973_,
		_w2971_,
		_w2972_
	);
	LUT2 #(
		.INIT('h8)
	) name1465 (
		\TM0_pad ,
		\_2101__reg/NET0131 ,
		_w2973_
	);
	LUT2 #(
		.INIT('h2)
	) name1466 (
		\WX2080_reg/NET0131 ,
		\WX2144_reg/NET0131 ,
		_w2974_
	);
	LUT2 #(
		.INIT('h4)
	) name1467 (
		\WX2080_reg/NET0131 ,
		\WX2144_reg/NET0131 ,
		_w2975_
	);
	LUT2 #(
		.INIT('h1)
	) name1468 (
		_w2974_,
		_w2975_,
		_w2976_
	);
	LUT2 #(
		.INIT('h2)
	) name1469 (
		\WX2016_reg/NET0131 ,
		_w2976_,
		_w2977_
	);
	LUT2 #(
		.INIT('h4)
	) name1470 (
		\WX2016_reg/NET0131 ,
		_w2976_,
		_w2978_
	);
	LUT2 #(
		.INIT('h1)
	) name1471 (
		_w2977_,
		_w2978_,
		_w2979_
	);
	LUT2 #(
		.INIT('h2)
	) name1472 (
		\TM1_pad ,
		\WX1952_reg/NET0131 ,
		_w2980_
	);
	LUT2 #(
		.INIT('h4)
	) name1473 (
		\TM1_pad ,
		\WX1952_reg/NET0131 ,
		_w2981_
	);
	LUT2 #(
		.INIT('h1)
	) name1474 (
		_w2980_,
		_w2981_,
		_w2982_
	);
	LUT2 #(
		.INIT('h4)
	) name1475 (
		_w2979_,
		_w2982_,
		_w2983_
	);
	LUT2 #(
		.INIT('h2)
	) name1476 (
		_w2979_,
		_w2982_,
		_w2984_
	);
	LUT2 #(
		.INIT('h1)
	) name1477 (
		\TM0_pad ,
		_w2983_,
		_w2985_
	);
	LUT2 #(
		.INIT('h4)
	) name1478 (
		_w2984_,
		_w2985_,
		_w2986_
	);
	LUT2 #(
		.INIT('h1)
	) name1479 (
		_w2973_,
		_w2986_,
		_w2987_
	);
	LUT2 #(
		.INIT('h2)
	) name1480 (
		_w1976_,
		_w2987_,
		_w2988_
	);
	LUT2 #(
		.INIT('h1)
	) name1481 (
		_w2972_,
		_w2988_,
		_w2989_
	);
	LUT2 #(
		.INIT('h2)
	) name1482 (
		\WX11127_reg/NET0131 ,
		\WX11191_reg/NET0131 ,
		_w2990_
	);
	LUT2 #(
		.INIT('h4)
	) name1483 (
		\WX11127_reg/NET0131 ,
		\WX11191_reg/NET0131 ,
		_w2991_
	);
	LUT2 #(
		.INIT('h1)
	) name1484 (
		_w2990_,
		_w2991_,
		_w2992_
	);
	LUT2 #(
		.INIT('h2)
	) name1485 (
		\WX11063_reg/NET0131 ,
		_w2992_,
		_w2993_
	);
	LUT2 #(
		.INIT('h4)
	) name1486 (
		\WX11063_reg/NET0131 ,
		_w2992_,
		_w2994_
	);
	LUT2 #(
		.INIT('h1)
	) name1487 (
		_w2993_,
		_w2994_,
		_w2995_
	);
	LUT2 #(
		.INIT('h2)
	) name1488 (
		\TM1_pad ,
		\WX10999_reg/NET0131 ,
		_w2996_
	);
	LUT2 #(
		.INIT('h4)
	) name1489 (
		\TM1_pad ,
		\WX10999_reg/NET0131 ,
		_w2997_
	);
	LUT2 #(
		.INIT('h1)
	) name1490 (
		_w2996_,
		_w2997_,
		_w2998_
	);
	LUT2 #(
		.INIT('h4)
	) name1491 (
		_w2995_,
		_w2998_,
		_w2999_
	);
	LUT2 #(
		.INIT('h2)
	) name1492 (
		_w2995_,
		_w2998_,
		_w3000_
	);
	LUT2 #(
		.INIT('h1)
	) name1493 (
		\TM0_pad ,
		_w2999_,
		_w3001_
	);
	LUT2 #(
		.INIT('h4)
	) name1494 (
		_w3000_,
		_w3001_,
		_w3002_
	);
	LUT2 #(
		.INIT('h1)
	) name1495 (
		_w1778_,
		_w3002_,
		_w3003_
	);
	LUT2 #(
		.INIT('h2)
	) name1496 (
		_w1973_,
		_w3003_,
		_w3004_
	);
	LUT2 #(
		.INIT('h1)
	) name1497 (
		\DATA_0_26_pad ,
		\TM0_pad ,
		_w3005_
	);
	LUT2 #(
		.INIT('h2)
	) name1498 (
		\TM0_pad ,
		\_2359__reg/NET0131 ,
		_w3006_
	);
	LUT2 #(
		.INIT('h2)
	) name1499 (
		_w1976_,
		_w3005_,
		_w3007_
	);
	LUT2 #(
		.INIT('h4)
	) name1500 (
		_w3006_,
		_w3007_,
		_w3008_
	);
	LUT2 #(
		.INIT('h1)
	) name1501 (
		_w3004_,
		_w3008_,
		_w3009_
	);
	LUT2 #(
		.INIT('h8)
	) name1502 (
		RESET_pad,
		\WX10837_reg/NET0131 ,
		_w3010_
	);
	LUT2 #(
		.INIT('h4)
	) name1503 (
		_w1521_,
		_w1973_,
		_w3011_
	);
	LUT2 #(
		.INIT('h2)
	) name1504 (
		\WX3401_reg/NET0131 ,
		\WX3465_reg/NET0131 ,
		_w3012_
	);
	LUT2 #(
		.INIT('h4)
	) name1505 (
		\WX3401_reg/NET0131 ,
		\WX3465_reg/NET0131 ,
		_w3013_
	);
	LUT2 #(
		.INIT('h1)
	) name1506 (
		_w3012_,
		_w3013_,
		_w3014_
	);
	LUT2 #(
		.INIT('h2)
	) name1507 (
		\WX3273_reg/NET0131 ,
		\WX3337_reg/NET0131 ,
		_w3015_
	);
	LUT2 #(
		.INIT('h4)
	) name1508 (
		\WX3273_reg/NET0131 ,
		\WX3337_reg/NET0131 ,
		_w3016_
	);
	LUT2 #(
		.INIT('h1)
	) name1509 (
		_w3015_,
		_w3016_,
		_w3017_
	);
	LUT2 #(
		.INIT('h4)
	) name1510 (
		_w3014_,
		_w3017_,
		_w3018_
	);
	LUT2 #(
		.INIT('h2)
	) name1511 (
		_w3014_,
		_w3017_,
		_w3019_
	);
	LUT2 #(
		.INIT('h1)
	) name1512 (
		\TM0_pad ,
		_w3018_,
		_w3020_
	);
	LUT2 #(
		.INIT('h4)
	) name1513 (
		_w3019_,
		_w3020_,
		_w3021_
	);
	LUT2 #(
		.INIT('h2)
	) name1514 (
		_w3011_,
		_w3021_,
		_w3022_
	);
	LUT2 #(
		.INIT('h2)
	) name1515 (
		\TM0_pad ,
		\_2151__reg/NET0131 ,
		_w3023_
	);
	LUT2 #(
		.INIT('h2)
	) name1516 (
		\WX4694_reg/NET0131 ,
		\WX4758_reg/NET0131 ,
		_w3024_
	);
	LUT2 #(
		.INIT('h4)
	) name1517 (
		\WX4694_reg/NET0131 ,
		\WX4758_reg/NET0131 ,
		_w3025_
	);
	LUT2 #(
		.INIT('h1)
	) name1518 (
		_w3024_,
		_w3025_,
		_w3026_
	);
	LUT2 #(
		.INIT('h2)
	) name1519 (
		\WX4566_reg/NET0131 ,
		\WX4630_reg/NET0131 ,
		_w3027_
	);
	LUT2 #(
		.INIT('h4)
	) name1520 (
		\WX4566_reg/NET0131 ,
		\WX4630_reg/NET0131 ,
		_w3028_
	);
	LUT2 #(
		.INIT('h1)
	) name1521 (
		_w3027_,
		_w3028_,
		_w3029_
	);
	LUT2 #(
		.INIT('h4)
	) name1522 (
		_w3026_,
		_w3029_,
		_w3030_
	);
	LUT2 #(
		.INIT('h2)
	) name1523 (
		_w3026_,
		_w3029_,
		_w3031_
	);
	LUT2 #(
		.INIT('h1)
	) name1524 (
		\TM0_pad ,
		_w3030_,
		_w3032_
	);
	LUT2 #(
		.INIT('h4)
	) name1525 (
		_w3031_,
		_w3032_,
		_w3033_
	);
	LUT2 #(
		.INIT('h2)
	) name1526 (
		_w1976_,
		_w3023_,
		_w3034_
	);
	LUT2 #(
		.INIT('h4)
	) name1527 (
		_w3033_,
		_w3034_,
		_w3035_
	);
	LUT2 #(
		.INIT('h1)
	) name1528 (
		_w3022_,
		_w3035_,
		_w3036_
	);
	LUT2 #(
		.INIT('h2)
	) name1529 (
		_w2341_,
		_w2966_,
		_w3037_
	);
	LUT2 #(
		.INIT('h2)
	) name1530 (
		\TM0_pad ,
		\_2283__reg/NET0131 ,
		_w3038_
	);
	LUT2 #(
		.INIT('h2)
	) name1531 (
		\WX9858_reg/NET0131 ,
		\WX9922_reg/NET0131 ,
		_w3039_
	);
	LUT2 #(
		.INIT('h4)
	) name1532 (
		\WX9858_reg/NET0131 ,
		\WX9922_reg/NET0131 ,
		_w3040_
	);
	LUT2 #(
		.INIT('h1)
	) name1533 (
		_w3039_,
		_w3040_,
		_w3041_
	);
	LUT2 #(
		.INIT('h2)
	) name1534 (
		\WX9730_reg/NET0131 ,
		\WX9794_reg/NET0131 ,
		_w3042_
	);
	LUT2 #(
		.INIT('h4)
	) name1535 (
		\WX9730_reg/NET0131 ,
		\WX9794_reg/NET0131 ,
		_w3043_
	);
	LUT2 #(
		.INIT('h1)
	) name1536 (
		_w3042_,
		_w3043_,
		_w3044_
	);
	LUT2 #(
		.INIT('h4)
	) name1537 (
		_w3041_,
		_w3044_,
		_w3045_
	);
	LUT2 #(
		.INIT('h2)
	) name1538 (
		_w3041_,
		_w3044_,
		_w3046_
	);
	LUT2 #(
		.INIT('h1)
	) name1539 (
		\TM0_pad ,
		_w3045_,
		_w3047_
	);
	LUT2 #(
		.INIT('h4)
	) name1540 (
		_w3046_,
		_w3047_,
		_w3048_
	);
	LUT2 #(
		.INIT('h2)
	) name1541 (
		_w1976_,
		_w3038_,
		_w3049_
	);
	LUT2 #(
		.INIT('h4)
	) name1542 (
		_w3048_,
		_w3049_,
		_w3050_
	);
	LUT2 #(
		.INIT('h1)
	) name1543 (
		_w3037_,
		_w3050_,
		_w3051_
	);
	LUT2 #(
		.INIT('h8)
	) name1544 (
		\TM0_pad ,
		\_2134__reg/NET0131 ,
		_w3052_
	);
	LUT2 #(
		.INIT('h2)
	) name1545 (
		\WX3371_reg/NET0131 ,
		\WX3435_reg/NET0131 ,
		_w3053_
	);
	LUT2 #(
		.INIT('h4)
	) name1546 (
		\WX3371_reg/NET0131 ,
		\WX3435_reg/NET0131 ,
		_w3054_
	);
	LUT2 #(
		.INIT('h1)
	) name1547 (
		_w3053_,
		_w3054_,
		_w3055_
	);
	LUT2 #(
		.INIT('h2)
	) name1548 (
		\WX3307_reg/NET0131 ,
		_w3055_,
		_w3056_
	);
	LUT2 #(
		.INIT('h4)
	) name1549 (
		\WX3307_reg/NET0131 ,
		_w3055_,
		_w3057_
	);
	LUT2 #(
		.INIT('h1)
	) name1550 (
		_w3056_,
		_w3057_,
		_w3058_
	);
	LUT2 #(
		.INIT('h2)
	) name1551 (
		\TM1_pad ,
		\WX3243_reg/NET0131 ,
		_w3059_
	);
	LUT2 #(
		.INIT('h4)
	) name1552 (
		\TM1_pad ,
		\WX3243_reg/NET0131 ,
		_w3060_
	);
	LUT2 #(
		.INIT('h1)
	) name1553 (
		_w3059_,
		_w3060_,
		_w3061_
	);
	LUT2 #(
		.INIT('h4)
	) name1554 (
		_w3058_,
		_w3061_,
		_w3062_
	);
	LUT2 #(
		.INIT('h2)
	) name1555 (
		_w3058_,
		_w3061_,
		_w3063_
	);
	LUT2 #(
		.INIT('h1)
	) name1556 (
		\TM0_pad ,
		_w3062_,
		_w3064_
	);
	LUT2 #(
		.INIT('h4)
	) name1557 (
		_w3063_,
		_w3064_,
		_w3065_
	);
	LUT2 #(
		.INIT('h1)
	) name1558 (
		_w3052_,
		_w3065_,
		_w3066_
	);
	LUT2 #(
		.INIT('h2)
	) name1559 (
		_w1976_,
		_w3066_,
		_w3067_
	);
	LUT2 #(
		.INIT('h1)
	) name1560 (
		_w1762_,
		_w2821_,
		_w3068_
	);
	LUT2 #(
		.INIT('h2)
	) name1561 (
		_w1973_,
		_w3068_,
		_w3069_
	);
	LUT2 #(
		.INIT('h1)
	) name1562 (
		_w3067_,
		_w3069_,
		_w3070_
	);
	LUT2 #(
		.INIT('h2)
	) name1563 (
		_w1974_,
		_w2883_,
		_w3071_
	);
	LUT2 #(
		.INIT('h2)
	) name1564 (
		\TM0_pad ,
		\_2316__reg/NET0131 ,
		_w3072_
	);
	LUT2 #(
		.INIT('h2)
	) name1565 (
		\WX11149_reg/NET0131 ,
		\WX11213_reg/NET0131 ,
		_w3073_
	);
	LUT2 #(
		.INIT('h4)
	) name1566 (
		\WX11149_reg/NET0131 ,
		\WX11213_reg/NET0131 ,
		_w3074_
	);
	LUT2 #(
		.INIT('h1)
	) name1567 (
		_w3073_,
		_w3074_,
		_w3075_
	);
	LUT2 #(
		.INIT('h2)
	) name1568 (
		\WX11021_reg/NET0131 ,
		\WX11085_reg/NET0131 ,
		_w3076_
	);
	LUT2 #(
		.INIT('h4)
	) name1569 (
		\WX11021_reg/NET0131 ,
		\WX11085_reg/NET0131 ,
		_w3077_
	);
	LUT2 #(
		.INIT('h1)
	) name1570 (
		_w3076_,
		_w3077_,
		_w3078_
	);
	LUT2 #(
		.INIT('h4)
	) name1571 (
		_w3075_,
		_w3078_,
		_w3079_
	);
	LUT2 #(
		.INIT('h2)
	) name1572 (
		_w3075_,
		_w3078_,
		_w3080_
	);
	LUT2 #(
		.INIT('h1)
	) name1573 (
		\TM0_pad ,
		_w3079_,
		_w3081_
	);
	LUT2 #(
		.INIT('h4)
	) name1574 (
		_w3080_,
		_w3081_,
		_w3082_
	);
	LUT2 #(
		.INIT('h2)
	) name1575 (
		_w1976_,
		_w3072_,
		_w3083_
	);
	LUT2 #(
		.INIT('h4)
	) name1576 (
		_w3082_,
		_w3083_,
		_w3084_
	);
	LUT2 #(
		.INIT('h1)
	) name1577 (
		_w3071_,
		_w3084_,
		_w3085_
	);
	LUT2 #(
		.INIT('h2)
	) name1578 (
		_w2846_,
		_w2868_,
		_w3086_
	);
	LUT2 #(
		.INIT('h2)
	) name1579 (
		\TM0_pad ,
		\_2184__reg/NET0131 ,
		_w3087_
	);
	LUT2 #(
		.INIT('h2)
	) name1580 (
		\WX5985_reg/NET0131 ,
		\WX6049_reg/NET0131 ,
		_w3088_
	);
	LUT2 #(
		.INIT('h4)
	) name1581 (
		\WX5985_reg/NET0131 ,
		\WX6049_reg/NET0131 ,
		_w3089_
	);
	LUT2 #(
		.INIT('h1)
	) name1582 (
		_w3088_,
		_w3089_,
		_w3090_
	);
	LUT2 #(
		.INIT('h2)
	) name1583 (
		\WX5857_reg/NET0131 ,
		\WX5921_reg/NET0131 ,
		_w3091_
	);
	LUT2 #(
		.INIT('h4)
	) name1584 (
		\WX5857_reg/NET0131 ,
		\WX5921_reg/NET0131 ,
		_w3092_
	);
	LUT2 #(
		.INIT('h1)
	) name1585 (
		_w3091_,
		_w3092_,
		_w3093_
	);
	LUT2 #(
		.INIT('h4)
	) name1586 (
		_w3090_,
		_w3093_,
		_w3094_
	);
	LUT2 #(
		.INIT('h2)
	) name1587 (
		_w3090_,
		_w3093_,
		_w3095_
	);
	LUT2 #(
		.INIT('h1)
	) name1588 (
		\TM0_pad ,
		_w3094_,
		_w3096_
	);
	LUT2 #(
		.INIT('h4)
	) name1589 (
		_w3095_,
		_w3096_,
		_w3097_
	);
	LUT2 #(
		.INIT('h2)
	) name1590 (
		_w1976_,
		_w3087_,
		_w3098_
	);
	LUT2 #(
		.INIT('h4)
	) name1591 (
		_w3097_,
		_w3098_,
		_w3099_
	);
	LUT2 #(
		.INIT('h1)
	) name1592 (
		_w3086_,
		_w3099_,
		_w3100_
	);
	LUT2 #(
		.INIT('h2)
	) name1593 (
		_w2677_,
		_w2936_,
		_w3101_
	);
	LUT2 #(
		.INIT('h2)
	) name1594 (
		\TM0_pad ,
		\_2217__reg/NET0131 ,
		_w3102_
	);
	LUT2 #(
		.INIT('h2)
	) name1595 (
		\WX7276_reg/NET0131 ,
		\WX7340_reg/NET0131 ,
		_w3103_
	);
	LUT2 #(
		.INIT('h4)
	) name1596 (
		\WX7276_reg/NET0131 ,
		\WX7340_reg/NET0131 ,
		_w3104_
	);
	LUT2 #(
		.INIT('h1)
	) name1597 (
		_w3103_,
		_w3104_,
		_w3105_
	);
	LUT2 #(
		.INIT('h2)
	) name1598 (
		\WX7148_reg/NET0131 ,
		\WX7212_reg/NET0131 ,
		_w3106_
	);
	LUT2 #(
		.INIT('h4)
	) name1599 (
		\WX7148_reg/NET0131 ,
		\WX7212_reg/NET0131 ,
		_w3107_
	);
	LUT2 #(
		.INIT('h1)
	) name1600 (
		_w3106_,
		_w3107_,
		_w3108_
	);
	LUT2 #(
		.INIT('h4)
	) name1601 (
		_w3105_,
		_w3108_,
		_w3109_
	);
	LUT2 #(
		.INIT('h2)
	) name1602 (
		_w3105_,
		_w3108_,
		_w3110_
	);
	LUT2 #(
		.INIT('h1)
	) name1603 (
		\TM0_pad ,
		_w3109_,
		_w3111_
	);
	LUT2 #(
		.INIT('h4)
	) name1604 (
		_w3110_,
		_w3111_,
		_w3112_
	);
	LUT2 #(
		.INIT('h2)
	) name1605 (
		_w1976_,
		_w3102_,
		_w3113_
	);
	LUT2 #(
		.INIT('h4)
	) name1606 (
		_w3112_,
		_w3113_,
		_w3114_
	);
	LUT2 #(
		.INIT('h1)
	) name1607 (
		_w3101_,
		_w3114_,
		_w3115_
	);
	LUT2 #(
		.INIT('h2)
	) name1608 (
		_w2040_,
		_w2951_,
		_w3116_
	);
	LUT2 #(
		.INIT('h2)
	) name1609 (
		\TM0_pad ,
		\_2250__reg/NET0131 ,
		_w3117_
	);
	LUT2 #(
		.INIT('h2)
	) name1610 (
		\WX8567_reg/NET0131 ,
		\WX8631_reg/NET0131 ,
		_w3118_
	);
	LUT2 #(
		.INIT('h4)
	) name1611 (
		\WX8567_reg/NET0131 ,
		\WX8631_reg/NET0131 ,
		_w3119_
	);
	LUT2 #(
		.INIT('h1)
	) name1612 (
		_w3118_,
		_w3119_,
		_w3120_
	);
	LUT2 #(
		.INIT('h2)
	) name1613 (
		\WX8439_reg/NET0131 ,
		\WX8503_reg/NET0131 ,
		_w3121_
	);
	LUT2 #(
		.INIT('h4)
	) name1614 (
		\WX8439_reg/NET0131 ,
		\WX8503_reg/NET0131 ,
		_w3122_
	);
	LUT2 #(
		.INIT('h1)
	) name1615 (
		_w3121_,
		_w3122_,
		_w3123_
	);
	LUT2 #(
		.INIT('h4)
	) name1616 (
		_w3120_,
		_w3123_,
		_w3124_
	);
	LUT2 #(
		.INIT('h2)
	) name1617 (
		_w3120_,
		_w3123_,
		_w3125_
	);
	LUT2 #(
		.INIT('h1)
	) name1618 (
		\TM0_pad ,
		_w3124_,
		_w3126_
	);
	LUT2 #(
		.INIT('h4)
	) name1619 (
		_w3125_,
		_w3126_,
		_w3127_
	);
	LUT2 #(
		.INIT('h2)
	) name1620 (
		_w1976_,
		_w3117_,
		_w3128_
	);
	LUT2 #(
		.INIT('h4)
	) name1621 (
		_w3127_,
		_w3128_,
		_w3129_
	);
	LUT2 #(
		.INIT('h1)
	) name1622 (
		_w3116_,
		_w3129_,
		_w3130_
	);
	LUT2 #(
		.INIT('h1)
	) name1623 (
		\TM0_pad ,
		_w1739_,
		_w3131_
	);
	LUT2 #(
		.INIT('h1)
	) name1624 (
		_w1730_,
		_w3131_,
		_w3132_
	);
	LUT2 #(
		.INIT('h2)
	) name1625 (
		_w1973_,
		_w3132_,
		_w3133_
	);
	LUT2 #(
		.INIT('h8)
	) name1626 (
		\TM0_pad ,
		\_2100__reg/NET0131 ,
		_w3134_
	);
	LUT2 #(
		.INIT('h2)
	) name1627 (
		\WX2082_reg/NET0131 ,
		\WX2146_reg/NET0131 ,
		_w3135_
	);
	LUT2 #(
		.INIT('h4)
	) name1628 (
		\WX2082_reg/NET0131 ,
		\WX2146_reg/NET0131 ,
		_w3136_
	);
	LUT2 #(
		.INIT('h1)
	) name1629 (
		_w3135_,
		_w3136_,
		_w3137_
	);
	LUT2 #(
		.INIT('h2)
	) name1630 (
		\WX2018_reg/NET0131 ,
		_w3137_,
		_w3138_
	);
	LUT2 #(
		.INIT('h4)
	) name1631 (
		\WX2018_reg/NET0131 ,
		_w3137_,
		_w3139_
	);
	LUT2 #(
		.INIT('h1)
	) name1632 (
		_w3138_,
		_w3139_,
		_w3140_
	);
	LUT2 #(
		.INIT('h2)
	) name1633 (
		\TM1_pad ,
		\WX1954_reg/NET0131 ,
		_w3141_
	);
	LUT2 #(
		.INIT('h4)
	) name1634 (
		\TM1_pad ,
		\WX1954_reg/NET0131 ,
		_w3142_
	);
	LUT2 #(
		.INIT('h1)
	) name1635 (
		_w3141_,
		_w3142_,
		_w3143_
	);
	LUT2 #(
		.INIT('h4)
	) name1636 (
		_w3140_,
		_w3143_,
		_w3144_
	);
	LUT2 #(
		.INIT('h2)
	) name1637 (
		_w3140_,
		_w3143_,
		_w3145_
	);
	LUT2 #(
		.INIT('h1)
	) name1638 (
		\TM0_pad ,
		_w3144_,
		_w3146_
	);
	LUT2 #(
		.INIT('h4)
	) name1639 (
		_w3145_,
		_w3146_,
		_w3147_
	);
	LUT2 #(
		.INIT('h1)
	) name1640 (
		_w3134_,
		_w3147_,
		_w3148_
	);
	LUT2 #(
		.INIT('h2)
	) name1641 (
		_w1976_,
		_w3148_,
		_w3149_
	);
	LUT2 #(
		.INIT('h1)
	) name1642 (
		_w3133_,
		_w3149_,
		_w3150_
	);
	LUT2 #(
		.INIT('h2)
	) name1643 (
		\WX11129_reg/NET0131 ,
		\WX11193_reg/NET0131 ,
		_w3151_
	);
	LUT2 #(
		.INIT('h4)
	) name1644 (
		\WX11129_reg/NET0131 ,
		\WX11193_reg/NET0131 ,
		_w3152_
	);
	LUT2 #(
		.INIT('h1)
	) name1645 (
		_w3151_,
		_w3152_,
		_w3153_
	);
	LUT2 #(
		.INIT('h2)
	) name1646 (
		\WX11065_reg/NET0131 ,
		_w3153_,
		_w3154_
	);
	LUT2 #(
		.INIT('h4)
	) name1647 (
		\WX11065_reg/NET0131 ,
		_w3153_,
		_w3155_
	);
	LUT2 #(
		.INIT('h1)
	) name1648 (
		_w3154_,
		_w3155_,
		_w3156_
	);
	LUT2 #(
		.INIT('h2)
	) name1649 (
		\TM1_pad ,
		\WX11001_reg/NET0131 ,
		_w3157_
	);
	LUT2 #(
		.INIT('h4)
	) name1650 (
		\TM1_pad ,
		\WX11001_reg/NET0131 ,
		_w3158_
	);
	LUT2 #(
		.INIT('h1)
	) name1651 (
		_w3157_,
		_w3158_,
		_w3159_
	);
	LUT2 #(
		.INIT('h4)
	) name1652 (
		_w3156_,
		_w3159_,
		_w3160_
	);
	LUT2 #(
		.INIT('h2)
	) name1653 (
		_w3156_,
		_w3159_,
		_w3161_
	);
	LUT2 #(
		.INIT('h1)
	) name1654 (
		\TM0_pad ,
		_w3160_,
		_w3162_
	);
	LUT2 #(
		.INIT('h4)
	) name1655 (
		_w3161_,
		_w3162_,
		_w3163_
	);
	LUT2 #(
		.INIT('h1)
	) name1656 (
		_w1762_,
		_w3163_,
		_w3164_
	);
	LUT2 #(
		.INIT('h2)
	) name1657 (
		_w1973_,
		_w3164_,
		_w3165_
	);
	LUT2 #(
		.INIT('h1)
	) name1658 (
		\DATA_0_25_pad ,
		\TM0_pad ,
		_w3166_
	);
	LUT2 #(
		.INIT('h2)
	) name1659 (
		\TM0_pad ,
		\_2358__reg/NET0131 ,
		_w3167_
	);
	LUT2 #(
		.INIT('h2)
	) name1660 (
		_w1976_,
		_w3166_,
		_w3168_
	);
	LUT2 #(
		.INIT('h4)
	) name1661 (
		_w3167_,
		_w3168_,
		_w3169_
	);
	LUT2 #(
		.INIT('h1)
	) name1662 (
		_w3165_,
		_w3169_,
		_w3170_
	);
	LUT2 #(
		.INIT('h8)
	) name1663 (
		RESET_pad,
		\WX10839_reg/NET0131 ,
		_w3171_
	);
	LUT2 #(
		.INIT('h4)
	) name1664 (
		_w1959_,
		_w1973_,
		_w3172_
	);
	LUT2 #(
		.INIT('h2)
	) name1665 (
		\WX3403_reg/NET0131 ,
		\WX3467_reg/NET0131 ,
		_w3173_
	);
	LUT2 #(
		.INIT('h4)
	) name1666 (
		\WX3403_reg/NET0131 ,
		\WX3467_reg/NET0131 ,
		_w3174_
	);
	LUT2 #(
		.INIT('h1)
	) name1667 (
		_w3173_,
		_w3174_,
		_w3175_
	);
	LUT2 #(
		.INIT('h2)
	) name1668 (
		\WX3275_reg/NET0131 ,
		\WX3339_reg/NET0131 ,
		_w3176_
	);
	LUT2 #(
		.INIT('h4)
	) name1669 (
		\WX3275_reg/NET0131 ,
		\WX3339_reg/NET0131 ,
		_w3177_
	);
	LUT2 #(
		.INIT('h1)
	) name1670 (
		_w3176_,
		_w3177_,
		_w3178_
	);
	LUT2 #(
		.INIT('h4)
	) name1671 (
		_w3175_,
		_w3178_,
		_w3179_
	);
	LUT2 #(
		.INIT('h2)
	) name1672 (
		_w3175_,
		_w3178_,
		_w3180_
	);
	LUT2 #(
		.INIT('h1)
	) name1673 (
		\TM0_pad ,
		_w3179_,
		_w3181_
	);
	LUT2 #(
		.INIT('h4)
	) name1674 (
		_w3180_,
		_w3181_,
		_w3182_
	);
	LUT2 #(
		.INIT('h2)
	) name1675 (
		_w3172_,
		_w3182_,
		_w3183_
	);
	LUT2 #(
		.INIT('h2)
	) name1676 (
		\TM0_pad ,
		\_2150__reg/NET0131 ,
		_w3184_
	);
	LUT2 #(
		.INIT('h2)
	) name1677 (
		\WX4696_reg/NET0131 ,
		\WX4760_reg/NET0131 ,
		_w3185_
	);
	LUT2 #(
		.INIT('h4)
	) name1678 (
		\WX4696_reg/NET0131 ,
		\WX4760_reg/NET0131 ,
		_w3186_
	);
	LUT2 #(
		.INIT('h1)
	) name1679 (
		_w3185_,
		_w3186_,
		_w3187_
	);
	LUT2 #(
		.INIT('h2)
	) name1680 (
		\WX4568_reg/NET0131 ,
		\WX4632_reg/NET0131 ,
		_w3188_
	);
	LUT2 #(
		.INIT('h4)
	) name1681 (
		\WX4568_reg/NET0131 ,
		\WX4632_reg/NET0131 ,
		_w3189_
	);
	LUT2 #(
		.INIT('h1)
	) name1682 (
		_w3188_,
		_w3189_,
		_w3190_
	);
	LUT2 #(
		.INIT('h4)
	) name1683 (
		_w3187_,
		_w3190_,
		_w3191_
	);
	LUT2 #(
		.INIT('h2)
	) name1684 (
		_w3187_,
		_w3190_,
		_w3192_
	);
	LUT2 #(
		.INIT('h1)
	) name1685 (
		\TM0_pad ,
		_w3191_,
		_w3193_
	);
	LUT2 #(
		.INIT('h4)
	) name1686 (
		_w3192_,
		_w3193_,
		_w3194_
	);
	LUT2 #(
		.INIT('h2)
	) name1687 (
		_w1976_,
		_w3184_,
		_w3195_
	);
	LUT2 #(
		.INIT('h4)
	) name1688 (
		_w3194_,
		_w3195_,
		_w3196_
	);
	LUT2 #(
		.INIT('h1)
	) name1689 (
		_w3183_,
		_w3196_,
		_w3197_
	);
	LUT2 #(
		.INIT('h2)
	) name1690 (
		_w2040_,
		_w3127_,
		_w3198_
	);
	LUT2 #(
		.INIT('h2)
	) name1691 (
		\TM0_pad ,
		\_2282__reg/NET0131 ,
		_w3199_
	);
	LUT2 #(
		.INIT('h2)
	) name1692 (
		\WX9860_reg/NET0131 ,
		\WX9924_reg/NET0131 ,
		_w3200_
	);
	LUT2 #(
		.INIT('h4)
	) name1693 (
		\WX9860_reg/NET0131 ,
		\WX9924_reg/NET0131 ,
		_w3201_
	);
	LUT2 #(
		.INIT('h1)
	) name1694 (
		_w3200_,
		_w3201_,
		_w3202_
	);
	LUT2 #(
		.INIT('h2)
	) name1695 (
		\WX9732_reg/NET0131 ,
		\WX9796_reg/NET0131 ,
		_w3203_
	);
	LUT2 #(
		.INIT('h4)
	) name1696 (
		\WX9732_reg/NET0131 ,
		\WX9796_reg/NET0131 ,
		_w3204_
	);
	LUT2 #(
		.INIT('h1)
	) name1697 (
		_w3203_,
		_w3204_,
		_w3205_
	);
	LUT2 #(
		.INIT('h4)
	) name1698 (
		_w3202_,
		_w3205_,
		_w3206_
	);
	LUT2 #(
		.INIT('h2)
	) name1699 (
		_w3202_,
		_w3205_,
		_w3207_
	);
	LUT2 #(
		.INIT('h1)
	) name1700 (
		\TM0_pad ,
		_w3206_,
		_w3208_
	);
	LUT2 #(
		.INIT('h4)
	) name1701 (
		_w3207_,
		_w3208_,
		_w3209_
	);
	LUT2 #(
		.INIT('h2)
	) name1702 (
		_w1976_,
		_w3199_,
		_w3210_
	);
	LUT2 #(
		.INIT('h4)
	) name1703 (
		_w3209_,
		_w3210_,
		_w3211_
	);
	LUT2 #(
		.INIT('h1)
	) name1704 (
		_w3198_,
		_w3211_,
		_w3212_
	);
	LUT2 #(
		.INIT('h2)
	) name1705 (
		_w2341_,
		_w3048_,
		_w3213_
	);
	LUT2 #(
		.INIT('h2)
	) name1706 (
		\TM0_pad ,
		\_2315__reg/NET0131 ,
		_w3214_
	);
	LUT2 #(
		.INIT('h2)
	) name1707 (
		\WX11151_reg/NET0131 ,
		\WX11215_reg/NET0131 ,
		_w3215_
	);
	LUT2 #(
		.INIT('h4)
	) name1708 (
		\WX11151_reg/NET0131 ,
		\WX11215_reg/NET0131 ,
		_w3216_
	);
	LUT2 #(
		.INIT('h1)
	) name1709 (
		_w3215_,
		_w3216_,
		_w3217_
	);
	LUT2 #(
		.INIT('h2)
	) name1710 (
		\WX11023_reg/NET0131 ,
		\WX11087_reg/NET0131 ,
		_w3218_
	);
	LUT2 #(
		.INIT('h4)
	) name1711 (
		\WX11023_reg/NET0131 ,
		\WX11087_reg/NET0131 ,
		_w3219_
	);
	LUT2 #(
		.INIT('h1)
	) name1712 (
		_w3218_,
		_w3219_,
		_w3220_
	);
	LUT2 #(
		.INIT('h4)
	) name1713 (
		_w3217_,
		_w3220_,
		_w3221_
	);
	LUT2 #(
		.INIT('h2)
	) name1714 (
		_w3217_,
		_w3220_,
		_w3222_
	);
	LUT2 #(
		.INIT('h1)
	) name1715 (
		\TM0_pad ,
		_w3221_,
		_w3223_
	);
	LUT2 #(
		.INIT('h4)
	) name1716 (
		_w3222_,
		_w3223_,
		_w3224_
	);
	LUT2 #(
		.INIT('h2)
	) name1717 (
		_w1976_,
		_w3214_,
		_w3225_
	);
	LUT2 #(
		.INIT('h4)
	) name1718 (
		_w3224_,
		_w3225_,
		_w3226_
	);
	LUT2 #(
		.INIT('h1)
	) name1719 (
		_w3213_,
		_w3226_,
		_w3227_
	);
	LUT2 #(
		.INIT('h8)
	) name1720 (
		\TM0_pad ,
		\_2133__reg/NET0131 ,
		_w3228_
	);
	LUT2 #(
		.INIT('h2)
	) name1721 (
		\WX3373_reg/NET0131 ,
		\WX3437_reg/NET0131 ,
		_w3229_
	);
	LUT2 #(
		.INIT('h4)
	) name1722 (
		\WX3373_reg/NET0131 ,
		\WX3437_reg/NET0131 ,
		_w3230_
	);
	LUT2 #(
		.INIT('h1)
	) name1723 (
		_w3229_,
		_w3230_,
		_w3231_
	);
	LUT2 #(
		.INIT('h2)
	) name1724 (
		\WX3309_reg/NET0131 ,
		_w3231_,
		_w3232_
	);
	LUT2 #(
		.INIT('h4)
	) name1725 (
		\WX3309_reg/NET0131 ,
		_w3231_,
		_w3233_
	);
	LUT2 #(
		.INIT('h1)
	) name1726 (
		_w3232_,
		_w3233_,
		_w3234_
	);
	LUT2 #(
		.INIT('h2)
	) name1727 (
		\TM1_pad ,
		\WX3245_reg/NET0131 ,
		_w3235_
	);
	LUT2 #(
		.INIT('h4)
	) name1728 (
		\TM1_pad ,
		\WX3245_reg/NET0131 ,
		_w3236_
	);
	LUT2 #(
		.INIT('h1)
	) name1729 (
		_w3235_,
		_w3236_,
		_w3237_
	);
	LUT2 #(
		.INIT('h4)
	) name1730 (
		_w3234_,
		_w3237_,
		_w3238_
	);
	LUT2 #(
		.INIT('h2)
	) name1731 (
		_w3234_,
		_w3237_,
		_w3239_
	);
	LUT2 #(
		.INIT('h1)
	) name1732 (
		\TM0_pad ,
		_w3238_,
		_w3240_
	);
	LUT2 #(
		.INIT('h4)
	) name1733 (
		_w3239_,
		_w3240_,
		_w3241_
	);
	LUT2 #(
		.INIT('h1)
	) name1734 (
		_w3228_,
		_w3241_,
		_w3242_
	);
	LUT2 #(
		.INIT('h2)
	) name1735 (
		_w1976_,
		_w3242_,
		_w3243_
	);
	LUT2 #(
		.INIT('h1)
	) name1736 (
		_w1746_,
		_w2986_,
		_w3244_
	);
	LUT2 #(
		.INIT('h2)
	) name1737 (
		_w1973_,
		_w3244_,
		_w3245_
	);
	LUT2 #(
		.INIT('h1)
	) name1738 (
		_w3243_,
		_w3245_,
		_w3246_
	);
	LUT2 #(
		.INIT('h2)
	) name1739 (
		_w3011_,
		_w3033_,
		_w3247_
	);
	LUT2 #(
		.INIT('h2)
	) name1740 (
		\TM0_pad ,
		\_2183__reg/NET0131 ,
		_w3248_
	);
	LUT2 #(
		.INIT('h2)
	) name1741 (
		\WX5987_reg/NET0131 ,
		\WX6051_reg/NET0131 ,
		_w3249_
	);
	LUT2 #(
		.INIT('h4)
	) name1742 (
		\WX5987_reg/NET0131 ,
		\WX6051_reg/NET0131 ,
		_w3250_
	);
	LUT2 #(
		.INIT('h1)
	) name1743 (
		_w3249_,
		_w3250_,
		_w3251_
	);
	LUT2 #(
		.INIT('h2)
	) name1744 (
		\WX5859_reg/NET0131 ,
		\WX5923_reg/NET0131 ,
		_w3252_
	);
	LUT2 #(
		.INIT('h4)
	) name1745 (
		\WX5859_reg/NET0131 ,
		\WX5923_reg/NET0131 ,
		_w3253_
	);
	LUT2 #(
		.INIT('h1)
	) name1746 (
		_w3252_,
		_w3253_,
		_w3254_
	);
	LUT2 #(
		.INIT('h4)
	) name1747 (
		_w3251_,
		_w3254_,
		_w3255_
	);
	LUT2 #(
		.INIT('h2)
	) name1748 (
		_w3251_,
		_w3254_,
		_w3256_
	);
	LUT2 #(
		.INIT('h1)
	) name1749 (
		\TM0_pad ,
		_w3255_,
		_w3257_
	);
	LUT2 #(
		.INIT('h4)
	) name1750 (
		_w3256_,
		_w3257_,
		_w3258_
	);
	LUT2 #(
		.INIT('h2)
	) name1751 (
		_w1976_,
		_w3248_,
		_w3259_
	);
	LUT2 #(
		.INIT('h4)
	) name1752 (
		_w3258_,
		_w3259_,
		_w3260_
	);
	LUT2 #(
		.INIT('h1)
	) name1753 (
		_w3247_,
		_w3260_,
		_w3261_
	);
	LUT2 #(
		.INIT('h2)
	) name1754 (
		_w2846_,
		_w3097_,
		_w3262_
	);
	LUT2 #(
		.INIT('h2)
	) name1755 (
		\TM0_pad ,
		\_2216__reg/NET0131 ,
		_w3263_
	);
	LUT2 #(
		.INIT('h2)
	) name1756 (
		\WX7278_reg/NET0131 ,
		\WX7342_reg/NET0131 ,
		_w3264_
	);
	LUT2 #(
		.INIT('h4)
	) name1757 (
		\WX7278_reg/NET0131 ,
		\WX7342_reg/NET0131 ,
		_w3265_
	);
	LUT2 #(
		.INIT('h1)
	) name1758 (
		_w3264_,
		_w3265_,
		_w3266_
	);
	LUT2 #(
		.INIT('h2)
	) name1759 (
		\WX7150_reg/NET0131 ,
		\WX7214_reg/NET0131 ,
		_w3267_
	);
	LUT2 #(
		.INIT('h4)
	) name1760 (
		\WX7150_reg/NET0131 ,
		\WX7214_reg/NET0131 ,
		_w3268_
	);
	LUT2 #(
		.INIT('h1)
	) name1761 (
		_w3267_,
		_w3268_,
		_w3269_
	);
	LUT2 #(
		.INIT('h4)
	) name1762 (
		_w3266_,
		_w3269_,
		_w3270_
	);
	LUT2 #(
		.INIT('h2)
	) name1763 (
		_w3266_,
		_w3269_,
		_w3271_
	);
	LUT2 #(
		.INIT('h1)
	) name1764 (
		\TM0_pad ,
		_w3270_,
		_w3272_
	);
	LUT2 #(
		.INIT('h4)
	) name1765 (
		_w3271_,
		_w3272_,
		_w3273_
	);
	LUT2 #(
		.INIT('h2)
	) name1766 (
		_w1976_,
		_w3263_,
		_w3274_
	);
	LUT2 #(
		.INIT('h4)
	) name1767 (
		_w3273_,
		_w3274_,
		_w3275_
	);
	LUT2 #(
		.INIT('h1)
	) name1768 (
		_w3262_,
		_w3275_,
		_w3276_
	);
	LUT2 #(
		.INIT('h2)
	) name1769 (
		_w2677_,
		_w3112_,
		_w3277_
	);
	LUT2 #(
		.INIT('h2)
	) name1770 (
		\TM0_pad ,
		\_2249__reg/NET0131 ,
		_w3278_
	);
	LUT2 #(
		.INIT('h2)
	) name1771 (
		\WX8569_reg/NET0131 ,
		\WX8633_reg/NET0131 ,
		_w3279_
	);
	LUT2 #(
		.INIT('h4)
	) name1772 (
		\WX8569_reg/NET0131 ,
		\WX8633_reg/NET0131 ,
		_w3280_
	);
	LUT2 #(
		.INIT('h1)
	) name1773 (
		_w3279_,
		_w3280_,
		_w3281_
	);
	LUT2 #(
		.INIT('h2)
	) name1774 (
		\WX8441_reg/NET0131 ,
		\WX8505_reg/NET0131 ,
		_w3282_
	);
	LUT2 #(
		.INIT('h4)
	) name1775 (
		\WX8441_reg/NET0131 ,
		\WX8505_reg/NET0131 ,
		_w3283_
	);
	LUT2 #(
		.INIT('h1)
	) name1776 (
		_w3282_,
		_w3283_,
		_w3284_
	);
	LUT2 #(
		.INIT('h4)
	) name1777 (
		_w3281_,
		_w3284_,
		_w3285_
	);
	LUT2 #(
		.INIT('h2)
	) name1778 (
		_w3281_,
		_w3284_,
		_w3286_
	);
	LUT2 #(
		.INIT('h1)
	) name1779 (
		\TM0_pad ,
		_w3285_,
		_w3287_
	);
	LUT2 #(
		.INIT('h4)
	) name1780 (
		_w3286_,
		_w3287_,
		_w3288_
	);
	LUT2 #(
		.INIT('h2)
	) name1781 (
		_w1976_,
		_w3278_,
		_w3289_
	);
	LUT2 #(
		.INIT('h4)
	) name1782 (
		_w3288_,
		_w3289_,
		_w3290_
	);
	LUT2 #(
		.INIT('h1)
	) name1783 (
		_w3277_,
		_w3290_,
		_w3291_
	);
	LUT2 #(
		.INIT('h1)
	) name1784 (
		\TM0_pad ,
		_w1723_,
		_w3292_
	);
	LUT2 #(
		.INIT('h1)
	) name1785 (
		_w1714_,
		_w3292_,
		_w3293_
	);
	LUT2 #(
		.INIT('h2)
	) name1786 (
		_w1973_,
		_w3293_,
		_w3294_
	);
	LUT2 #(
		.INIT('h8)
	) name1787 (
		\TM0_pad ,
		\_2099__reg/NET0131 ,
		_w3295_
	);
	LUT2 #(
		.INIT('h2)
	) name1788 (
		\WX2084_reg/NET0131 ,
		\WX2148_reg/NET0131 ,
		_w3296_
	);
	LUT2 #(
		.INIT('h4)
	) name1789 (
		\WX2084_reg/NET0131 ,
		\WX2148_reg/NET0131 ,
		_w3297_
	);
	LUT2 #(
		.INIT('h1)
	) name1790 (
		_w3296_,
		_w3297_,
		_w3298_
	);
	LUT2 #(
		.INIT('h2)
	) name1791 (
		\WX2020_reg/NET0131 ,
		_w3298_,
		_w3299_
	);
	LUT2 #(
		.INIT('h4)
	) name1792 (
		\WX2020_reg/NET0131 ,
		_w3298_,
		_w3300_
	);
	LUT2 #(
		.INIT('h1)
	) name1793 (
		_w3299_,
		_w3300_,
		_w3301_
	);
	LUT2 #(
		.INIT('h2)
	) name1794 (
		\TM1_pad ,
		\WX1956_reg/NET0131 ,
		_w3302_
	);
	LUT2 #(
		.INIT('h4)
	) name1795 (
		\TM1_pad ,
		\WX1956_reg/NET0131 ,
		_w3303_
	);
	LUT2 #(
		.INIT('h1)
	) name1796 (
		_w3302_,
		_w3303_,
		_w3304_
	);
	LUT2 #(
		.INIT('h4)
	) name1797 (
		_w3301_,
		_w3304_,
		_w3305_
	);
	LUT2 #(
		.INIT('h2)
	) name1798 (
		_w3301_,
		_w3304_,
		_w3306_
	);
	LUT2 #(
		.INIT('h1)
	) name1799 (
		\TM0_pad ,
		_w3305_,
		_w3307_
	);
	LUT2 #(
		.INIT('h4)
	) name1800 (
		_w3306_,
		_w3307_,
		_w3308_
	);
	LUT2 #(
		.INIT('h1)
	) name1801 (
		_w3295_,
		_w3308_,
		_w3309_
	);
	LUT2 #(
		.INIT('h2)
	) name1802 (
		_w1976_,
		_w3309_,
		_w3310_
	);
	LUT2 #(
		.INIT('h1)
	) name1803 (
		_w3294_,
		_w3310_,
		_w3311_
	);
	LUT2 #(
		.INIT('h2)
	) name1804 (
		\WX11131_reg/NET0131 ,
		\WX11195_reg/NET0131 ,
		_w3312_
	);
	LUT2 #(
		.INIT('h4)
	) name1805 (
		\WX11131_reg/NET0131 ,
		\WX11195_reg/NET0131 ,
		_w3313_
	);
	LUT2 #(
		.INIT('h1)
	) name1806 (
		_w3312_,
		_w3313_,
		_w3314_
	);
	LUT2 #(
		.INIT('h2)
	) name1807 (
		\WX11067_reg/NET0131 ,
		_w3314_,
		_w3315_
	);
	LUT2 #(
		.INIT('h4)
	) name1808 (
		\WX11067_reg/NET0131 ,
		_w3314_,
		_w3316_
	);
	LUT2 #(
		.INIT('h1)
	) name1809 (
		_w3315_,
		_w3316_,
		_w3317_
	);
	LUT2 #(
		.INIT('h2)
	) name1810 (
		\TM1_pad ,
		\WX11003_reg/NET0131 ,
		_w3318_
	);
	LUT2 #(
		.INIT('h4)
	) name1811 (
		\TM1_pad ,
		\WX11003_reg/NET0131 ,
		_w3319_
	);
	LUT2 #(
		.INIT('h1)
	) name1812 (
		_w3318_,
		_w3319_,
		_w3320_
	);
	LUT2 #(
		.INIT('h4)
	) name1813 (
		_w3317_,
		_w3320_,
		_w3321_
	);
	LUT2 #(
		.INIT('h2)
	) name1814 (
		_w3317_,
		_w3320_,
		_w3322_
	);
	LUT2 #(
		.INIT('h1)
	) name1815 (
		\TM0_pad ,
		_w3321_,
		_w3323_
	);
	LUT2 #(
		.INIT('h4)
	) name1816 (
		_w3322_,
		_w3323_,
		_w3324_
	);
	LUT2 #(
		.INIT('h1)
	) name1817 (
		_w1746_,
		_w3324_,
		_w3325_
	);
	LUT2 #(
		.INIT('h2)
	) name1818 (
		_w1973_,
		_w3325_,
		_w3326_
	);
	LUT2 #(
		.INIT('h1)
	) name1819 (
		\DATA_0_24_pad ,
		\TM0_pad ,
		_w3327_
	);
	LUT2 #(
		.INIT('h2)
	) name1820 (
		\TM0_pad ,
		\_2357__reg/NET0131 ,
		_w3328_
	);
	LUT2 #(
		.INIT('h2)
	) name1821 (
		_w1976_,
		_w3327_,
		_w3329_
	);
	LUT2 #(
		.INIT('h4)
	) name1822 (
		_w3328_,
		_w3329_,
		_w3330_
	);
	LUT2 #(
		.INIT('h1)
	) name1823 (
		_w3326_,
		_w3330_,
		_w3331_
	);
	LUT2 #(
		.INIT('h8)
	) name1824 (
		RESET_pad,
		\WX10841_reg/NET0131 ,
		_w3332_
	);
	LUT2 #(
		.INIT('h2)
	) name1825 (
		\WX3405_reg/NET0131 ,
		\WX3469_reg/NET0131 ,
		_w3333_
	);
	LUT2 #(
		.INIT('h4)
	) name1826 (
		\WX3405_reg/NET0131 ,
		\WX3469_reg/NET0131 ,
		_w3334_
	);
	LUT2 #(
		.INIT('h1)
	) name1827 (
		_w3333_,
		_w3334_,
		_w3335_
	);
	LUT2 #(
		.INIT('h2)
	) name1828 (
		\WX3277_reg/NET0131 ,
		\WX3341_reg/NET0131 ,
		_w3336_
	);
	LUT2 #(
		.INIT('h4)
	) name1829 (
		\WX3277_reg/NET0131 ,
		\WX3341_reg/NET0131 ,
		_w3337_
	);
	LUT2 #(
		.INIT('h1)
	) name1830 (
		_w3336_,
		_w3337_,
		_w3338_
	);
	LUT2 #(
		.INIT('h4)
	) name1831 (
		_w3335_,
		_w3338_,
		_w3339_
	);
	LUT2 #(
		.INIT('h2)
	) name1832 (
		_w3335_,
		_w3338_,
		_w3340_
	);
	LUT2 #(
		.INIT('h1)
	) name1833 (
		\TM0_pad ,
		_w3339_,
		_w3341_
	);
	LUT2 #(
		.INIT('h4)
	) name1834 (
		_w3340_,
		_w3341_,
		_w3342_
	);
	LUT2 #(
		.INIT('h2)
	) name1835 (
		_w2023_,
		_w3342_,
		_w3343_
	);
	LUT2 #(
		.INIT('h2)
	) name1836 (
		\TM0_pad ,
		\_2149__reg/NET0131 ,
		_w3344_
	);
	LUT2 #(
		.INIT('h2)
	) name1837 (
		\WX4698_reg/NET0131 ,
		\WX4762_reg/NET0131 ,
		_w3345_
	);
	LUT2 #(
		.INIT('h4)
	) name1838 (
		\WX4698_reg/NET0131 ,
		\WX4762_reg/NET0131 ,
		_w3346_
	);
	LUT2 #(
		.INIT('h1)
	) name1839 (
		_w3345_,
		_w3346_,
		_w3347_
	);
	LUT2 #(
		.INIT('h2)
	) name1840 (
		\WX4570_reg/NET0131 ,
		\WX4634_reg/NET0131 ,
		_w3348_
	);
	LUT2 #(
		.INIT('h4)
	) name1841 (
		\WX4570_reg/NET0131 ,
		\WX4634_reg/NET0131 ,
		_w3349_
	);
	LUT2 #(
		.INIT('h1)
	) name1842 (
		_w3348_,
		_w3349_,
		_w3350_
	);
	LUT2 #(
		.INIT('h4)
	) name1843 (
		_w3347_,
		_w3350_,
		_w3351_
	);
	LUT2 #(
		.INIT('h2)
	) name1844 (
		_w3347_,
		_w3350_,
		_w3352_
	);
	LUT2 #(
		.INIT('h1)
	) name1845 (
		\TM0_pad ,
		_w3351_,
		_w3353_
	);
	LUT2 #(
		.INIT('h4)
	) name1846 (
		_w3352_,
		_w3353_,
		_w3354_
	);
	LUT2 #(
		.INIT('h2)
	) name1847 (
		_w1976_,
		_w3344_,
		_w3355_
	);
	LUT2 #(
		.INIT('h4)
	) name1848 (
		_w3354_,
		_w3355_,
		_w3356_
	);
	LUT2 #(
		.INIT('h1)
	) name1849 (
		_w3343_,
		_w3356_,
		_w3357_
	);
	LUT2 #(
		.INIT('h2)
	) name1850 (
		_w2677_,
		_w3288_,
		_w3358_
	);
	LUT2 #(
		.INIT('h2)
	) name1851 (
		\TM0_pad ,
		\_2281__reg/NET0131 ,
		_w3359_
	);
	LUT2 #(
		.INIT('h2)
	) name1852 (
		\WX9862_reg/NET0131 ,
		\WX9926_reg/NET0131 ,
		_w3360_
	);
	LUT2 #(
		.INIT('h4)
	) name1853 (
		\WX9862_reg/NET0131 ,
		\WX9926_reg/NET0131 ,
		_w3361_
	);
	LUT2 #(
		.INIT('h1)
	) name1854 (
		_w3360_,
		_w3361_,
		_w3362_
	);
	LUT2 #(
		.INIT('h2)
	) name1855 (
		\WX9734_reg/NET0131 ,
		\WX9798_reg/NET0131 ,
		_w3363_
	);
	LUT2 #(
		.INIT('h4)
	) name1856 (
		\WX9734_reg/NET0131 ,
		\WX9798_reg/NET0131 ,
		_w3364_
	);
	LUT2 #(
		.INIT('h1)
	) name1857 (
		_w3363_,
		_w3364_,
		_w3365_
	);
	LUT2 #(
		.INIT('h4)
	) name1858 (
		_w3362_,
		_w3365_,
		_w3366_
	);
	LUT2 #(
		.INIT('h2)
	) name1859 (
		_w3362_,
		_w3365_,
		_w3367_
	);
	LUT2 #(
		.INIT('h1)
	) name1860 (
		\TM0_pad ,
		_w3366_,
		_w3368_
	);
	LUT2 #(
		.INIT('h4)
	) name1861 (
		_w3367_,
		_w3368_,
		_w3369_
	);
	LUT2 #(
		.INIT('h2)
	) name1862 (
		_w1976_,
		_w3359_,
		_w3370_
	);
	LUT2 #(
		.INIT('h4)
	) name1863 (
		_w3369_,
		_w3370_,
		_w3371_
	);
	LUT2 #(
		.INIT('h1)
	) name1864 (
		_w3358_,
		_w3371_,
		_w3372_
	);
	LUT2 #(
		.INIT('h2)
	) name1865 (
		_w2040_,
		_w3209_,
		_w3373_
	);
	LUT2 #(
		.INIT('h2)
	) name1866 (
		\TM0_pad ,
		\_2314__reg/NET0131 ,
		_w3374_
	);
	LUT2 #(
		.INIT('h2)
	) name1867 (
		_w1976_,
		_w3374_,
		_w3375_
	);
	LUT2 #(
		.INIT('h4)
	) name1868 (
		_w2050_,
		_w3375_,
		_w3376_
	);
	LUT2 #(
		.INIT('h1)
	) name1869 (
		_w3373_,
		_w3376_,
		_w3377_
	);
	LUT2 #(
		.INIT('h8)
	) name1870 (
		\TM0_pad ,
		\_2132__reg/NET0131 ,
		_w3378_
	);
	LUT2 #(
		.INIT('h2)
	) name1871 (
		\WX3375_reg/NET0131 ,
		\WX3439_reg/NET0131 ,
		_w3379_
	);
	LUT2 #(
		.INIT('h4)
	) name1872 (
		\WX3375_reg/NET0131 ,
		\WX3439_reg/NET0131 ,
		_w3380_
	);
	LUT2 #(
		.INIT('h1)
	) name1873 (
		_w3379_,
		_w3380_,
		_w3381_
	);
	LUT2 #(
		.INIT('h2)
	) name1874 (
		\WX3311_reg/NET0131 ,
		_w3381_,
		_w3382_
	);
	LUT2 #(
		.INIT('h4)
	) name1875 (
		\WX3311_reg/NET0131 ,
		_w3381_,
		_w3383_
	);
	LUT2 #(
		.INIT('h1)
	) name1876 (
		_w3382_,
		_w3383_,
		_w3384_
	);
	LUT2 #(
		.INIT('h2)
	) name1877 (
		\TM1_pad ,
		\WX3247_reg/NET0131 ,
		_w3385_
	);
	LUT2 #(
		.INIT('h4)
	) name1878 (
		\TM1_pad ,
		\WX3247_reg/NET0131 ,
		_w3386_
	);
	LUT2 #(
		.INIT('h1)
	) name1879 (
		_w3385_,
		_w3386_,
		_w3387_
	);
	LUT2 #(
		.INIT('h4)
	) name1880 (
		_w3384_,
		_w3387_,
		_w3388_
	);
	LUT2 #(
		.INIT('h2)
	) name1881 (
		_w3384_,
		_w3387_,
		_w3389_
	);
	LUT2 #(
		.INIT('h1)
	) name1882 (
		\TM0_pad ,
		_w3388_,
		_w3390_
	);
	LUT2 #(
		.INIT('h4)
	) name1883 (
		_w3389_,
		_w3390_,
		_w3391_
	);
	LUT2 #(
		.INIT('h1)
	) name1884 (
		_w3378_,
		_w3391_,
		_w3392_
	);
	LUT2 #(
		.INIT('h2)
	) name1885 (
		_w1976_,
		_w3392_,
		_w3393_
	);
	LUT2 #(
		.INIT('h1)
	) name1886 (
		_w1730_,
		_w3147_,
		_w3394_
	);
	LUT2 #(
		.INIT('h2)
	) name1887 (
		_w1973_,
		_w3394_,
		_w3395_
	);
	LUT2 #(
		.INIT('h1)
	) name1888 (
		_w3393_,
		_w3395_,
		_w3396_
	);
	LUT2 #(
		.INIT('h2)
	) name1889 (
		_w3172_,
		_w3194_,
		_w3397_
	);
	LUT2 #(
		.INIT('h2)
	) name1890 (
		\TM0_pad ,
		\_2182__reg/NET0131 ,
		_w3398_
	);
	LUT2 #(
		.INIT('h2)
	) name1891 (
		\WX5989_reg/NET0131 ,
		\WX6053_reg/NET0131 ,
		_w3399_
	);
	LUT2 #(
		.INIT('h4)
	) name1892 (
		\WX5989_reg/NET0131 ,
		\WX6053_reg/NET0131 ,
		_w3400_
	);
	LUT2 #(
		.INIT('h1)
	) name1893 (
		_w3399_,
		_w3400_,
		_w3401_
	);
	LUT2 #(
		.INIT('h2)
	) name1894 (
		\WX5861_reg/NET0131 ,
		\WX5925_reg/NET0131 ,
		_w3402_
	);
	LUT2 #(
		.INIT('h4)
	) name1895 (
		\WX5861_reg/NET0131 ,
		\WX5925_reg/NET0131 ,
		_w3403_
	);
	LUT2 #(
		.INIT('h1)
	) name1896 (
		_w3402_,
		_w3403_,
		_w3404_
	);
	LUT2 #(
		.INIT('h4)
	) name1897 (
		_w3401_,
		_w3404_,
		_w3405_
	);
	LUT2 #(
		.INIT('h2)
	) name1898 (
		_w3401_,
		_w3404_,
		_w3406_
	);
	LUT2 #(
		.INIT('h1)
	) name1899 (
		\TM0_pad ,
		_w3405_,
		_w3407_
	);
	LUT2 #(
		.INIT('h4)
	) name1900 (
		_w3406_,
		_w3407_,
		_w3408_
	);
	LUT2 #(
		.INIT('h2)
	) name1901 (
		_w1976_,
		_w3398_,
		_w3409_
	);
	LUT2 #(
		.INIT('h4)
	) name1902 (
		_w3408_,
		_w3409_,
		_w3410_
	);
	LUT2 #(
		.INIT('h1)
	) name1903 (
		_w3397_,
		_w3410_,
		_w3411_
	);
	LUT2 #(
		.INIT('h2)
	) name1904 (
		_w3011_,
		_w3258_,
		_w3412_
	);
	LUT2 #(
		.INIT('h2)
	) name1905 (
		\TM0_pad ,
		\_2215__reg/NET0131 ,
		_w3413_
	);
	LUT2 #(
		.INIT('h2)
	) name1906 (
		\WX7280_reg/NET0131 ,
		\WX7344_reg/NET0131 ,
		_w3414_
	);
	LUT2 #(
		.INIT('h4)
	) name1907 (
		\WX7280_reg/NET0131 ,
		\WX7344_reg/NET0131 ,
		_w3415_
	);
	LUT2 #(
		.INIT('h1)
	) name1908 (
		_w3414_,
		_w3415_,
		_w3416_
	);
	LUT2 #(
		.INIT('h2)
	) name1909 (
		\WX7152_reg/NET0131 ,
		\WX7216_reg/NET0131 ,
		_w3417_
	);
	LUT2 #(
		.INIT('h4)
	) name1910 (
		\WX7152_reg/NET0131 ,
		\WX7216_reg/NET0131 ,
		_w3418_
	);
	LUT2 #(
		.INIT('h1)
	) name1911 (
		_w3417_,
		_w3418_,
		_w3419_
	);
	LUT2 #(
		.INIT('h4)
	) name1912 (
		_w3416_,
		_w3419_,
		_w3420_
	);
	LUT2 #(
		.INIT('h2)
	) name1913 (
		_w3416_,
		_w3419_,
		_w3421_
	);
	LUT2 #(
		.INIT('h1)
	) name1914 (
		\TM0_pad ,
		_w3420_,
		_w3422_
	);
	LUT2 #(
		.INIT('h4)
	) name1915 (
		_w3421_,
		_w3422_,
		_w3423_
	);
	LUT2 #(
		.INIT('h2)
	) name1916 (
		_w1976_,
		_w3413_,
		_w3424_
	);
	LUT2 #(
		.INIT('h4)
	) name1917 (
		_w3423_,
		_w3424_,
		_w3425_
	);
	LUT2 #(
		.INIT('h1)
	) name1918 (
		_w3412_,
		_w3425_,
		_w3426_
	);
	LUT2 #(
		.INIT('h2)
	) name1919 (
		_w2846_,
		_w3273_,
		_w3427_
	);
	LUT2 #(
		.INIT('h2)
	) name1920 (
		\TM0_pad ,
		\_2248__reg/NET0131 ,
		_w3428_
	);
	LUT2 #(
		.INIT('h2)
	) name1921 (
		\WX8571_reg/NET0131 ,
		\WX8635_reg/NET0131 ,
		_w3429_
	);
	LUT2 #(
		.INIT('h4)
	) name1922 (
		\WX8571_reg/NET0131 ,
		\WX8635_reg/NET0131 ,
		_w3430_
	);
	LUT2 #(
		.INIT('h1)
	) name1923 (
		_w3429_,
		_w3430_,
		_w3431_
	);
	LUT2 #(
		.INIT('h2)
	) name1924 (
		\WX8443_reg/NET0131 ,
		\WX8507_reg/NET0131 ,
		_w3432_
	);
	LUT2 #(
		.INIT('h4)
	) name1925 (
		\WX8443_reg/NET0131 ,
		\WX8507_reg/NET0131 ,
		_w3433_
	);
	LUT2 #(
		.INIT('h1)
	) name1926 (
		_w3432_,
		_w3433_,
		_w3434_
	);
	LUT2 #(
		.INIT('h4)
	) name1927 (
		_w3431_,
		_w3434_,
		_w3435_
	);
	LUT2 #(
		.INIT('h2)
	) name1928 (
		_w3431_,
		_w3434_,
		_w3436_
	);
	LUT2 #(
		.INIT('h1)
	) name1929 (
		\TM0_pad ,
		_w3435_,
		_w3437_
	);
	LUT2 #(
		.INIT('h4)
	) name1930 (
		_w3436_,
		_w3437_,
		_w3438_
	);
	LUT2 #(
		.INIT('h2)
	) name1931 (
		_w1976_,
		_w3428_,
		_w3439_
	);
	LUT2 #(
		.INIT('h4)
	) name1932 (
		_w3438_,
		_w3439_,
		_w3440_
	);
	LUT2 #(
		.INIT('h1)
	) name1933 (
		_w3427_,
		_w3440_,
		_w3441_
	);
	LUT2 #(
		.INIT('h1)
	) name1934 (
		\TM0_pad ,
		_w1707_,
		_w3442_
	);
	LUT2 #(
		.INIT('h1)
	) name1935 (
		_w1698_,
		_w3442_,
		_w3443_
	);
	LUT2 #(
		.INIT('h2)
	) name1936 (
		_w1973_,
		_w3443_,
		_w3444_
	);
	LUT2 #(
		.INIT('h8)
	) name1937 (
		\TM0_pad ,
		\_2098__reg/NET0131 ,
		_w3445_
	);
	LUT2 #(
		.INIT('h2)
	) name1938 (
		\WX2086_reg/NET0131 ,
		\WX2150_reg/NET0131 ,
		_w3446_
	);
	LUT2 #(
		.INIT('h4)
	) name1939 (
		\WX2086_reg/NET0131 ,
		\WX2150_reg/NET0131 ,
		_w3447_
	);
	LUT2 #(
		.INIT('h1)
	) name1940 (
		_w3446_,
		_w3447_,
		_w3448_
	);
	LUT2 #(
		.INIT('h2)
	) name1941 (
		\WX2022_reg/NET0131 ,
		_w3448_,
		_w3449_
	);
	LUT2 #(
		.INIT('h4)
	) name1942 (
		\WX2022_reg/NET0131 ,
		_w3448_,
		_w3450_
	);
	LUT2 #(
		.INIT('h1)
	) name1943 (
		_w3449_,
		_w3450_,
		_w3451_
	);
	LUT2 #(
		.INIT('h2)
	) name1944 (
		\TM1_pad ,
		\WX1958_reg/NET0131 ,
		_w3452_
	);
	LUT2 #(
		.INIT('h4)
	) name1945 (
		\TM1_pad ,
		\WX1958_reg/NET0131 ,
		_w3453_
	);
	LUT2 #(
		.INIT('h1)
	) name1946 (
		_w3452_,
		_w3453_,
		_w3454_
	);
	LUT2 #(
		.INIT('h4)
	) name1947 (
		_w3451_,
		_w3454_,
		_w3455_
	);
	LUT2 #(
		.INIT('h2)
	) name1948 (
		_w3451_,
		_w3454_,
		_w3456_
	);
	LUT2 #(
		.INIT('h1)
	) name1949 (
		\TM0_pad ,
		_w3455_,
		_w3457_
	);
	LUT2 #(
		.INIT('h4)
	) name1950 (
		_w3456_,
		_w3457_,
		_w3458_
	);
	LUT2 #(
		.INIT('h1)
	) name1951 (
		_w3445_,
		_w3458_,
		_w3459_
	);
	LUT2 #(
		.INIT('h2)
	) name1952 (
		_w1976_,
		_w3459_,
		_w3460_
	);
	LUT2 #(
		.INIT('h1)
	) name1953 (
		_w3444_,
		_w3460_,
		_w3461_
	);
	LUT2 #(
		.INIT('h2)
	) name1954 (
		\WX11133_reg/NET0131 ,
		\WX11197_reg/NET0131 ,
		_w3462_
	);
	LUT2 #(
		.INIT('h4)
	) name1955 (
		\WX11133_reg/NET0131 ,
		\WX11197_reg/NET0131 ,
		_w3463_
	);
	LUT2 #(
		.INIT('h1)
	) name1956 (
		_w3462_,
		_w3463_,
		_w3464_
	);
	LUT2 #(
		.INIT('h2)
	) name1957 (
		\WX11069_reg/NET0131 ,
		_w3464_,
		_w3465_
	);
	LUT2 #(
		.INIT('h4)
	) name1958 (
		\WX11069_reg/NET0131 ,
		_w3464_,
		_w3466_
	);
	LUT2 #(
		.INIT('h1)
	) name1959 (
		_w3465_,
		_w3466_,
		_w3467_
	);
	LUT2 #(
		.INIT('h2)
	) name1960 (
		\TM1_pad ,
		\WX11005_reg/NET0131 ,
		_w3468_
	);
	LUT2 #(
		.INIT('h4)
	) name1961 (
		\TM1_pad ,
		\WX11005_reg/NET0131 ,
		_w3469_
	);
	LUT2 #(
		.INIT('h1)
	) name1962 (
		_w3468_,
		_w3469_,
		_w3470_
	);
	LUT2 #(
		.INIT('h4)
	) name1963 (
		_w3467_,
		_w3470_,
		_w3471_
	);
	LUT2 #(
		.INIT('h2)
	) name1964 (
		_w3467_,
		_w3470_,
		_w3472_
	);
	LUT2 #(
		.INIT('h1)
	) name1965 (
		\TM0_pad ,
		_w3471_,
		_w3473_
	);
	LUT2 #(
		.INIT('h4)
	) name1966 (
		_w3472_,
		_w3473_,
		_w3474_
	);
	LUT2 #(
		.INIT('h1)
	) name1967 (
		_w1730_,
		_w3474_,
		_w3475_
	);
	LUT2 #(
		.INIT('h2)
	) name1968 (
		_w1973_,
		_w3475_,
		_w3476_
	);
	LUT2 #(
		.INIT('h1)
	) name1969 (
		\DATA_0_23_pad ,
		\TM0_pad ,
		_w3477_
	);
	LUT2 #(
		.INIT('h2)
	) name1970 (
		\TM0_pad ,
		\_2356__reg/NET0131 ,
		_w3478_
	);
	LUT2 #(
		.INIT('h2)
	) name1971 (
		_w1976_,
		_w3477_,
		_w3479_
	);
	LUT2 #(
		.INIT('h4)
	) name1972 (
		_w3478_,
		_w3479_,
		_w3480_
	);
	LUT2 #(
		.INIT('h1)
	) name1973 (
		_w3476_,
		_w3480_,
		_w3481_
	);
	LUT2 #(
		.INIT('h8)
	) name1974 (
		RESET_pad,
		\WX10843_reg/NET0131 ,
		_w3482_
	);
	LUT2 #(
		.INIT('h4)
	) name1975 (
		_w1933_,
		_w1973_,
		_w3483_
	);
	LUT2 #(
		.INIT('h2)
	) name1976 (
		\WX3407_reg/NET0131 ,
		\WX3471_reg/NET0131 ,
		_w3484_
	);
	LUT2 #(
		.INIT('h4)
	) name1977 (
		\WX3407_reg/NET0131 ,
		\WX3471_reg/NET0131 ,
		_w3485_
	);
	LUT2 #(
		.INIT('h1)
	) name1978 (
		_w3484_,
		_w3485_,
		_w3486_
	);
	LUT2 #(
		.INIT('h2)
	) name1979 (
		\WX3279_reg/NET0131 ,
		\WX3343_reg/NET0131 ,
		_w3487_
	);
	LUT2 #(
		.INIT('h4)
	) name1980 (
		\WX3279_reg/NET0131 ,
		\WX3343_reg/NET0131 ,
		_w3488_
	);
	LUT2 #(
		.INIT('h1)
	) name1981 (
		_w3487_,
		_w3488_,
		_w3489_
	);
	LUT2 #(
		.INIT('h4)
	) name1982 (
		_w3486_,
		_w3489_,
		_w3490_
	);
	LUT2 #(
		.INIT('h2)
	) name1983 (
		_w3486_,
		_w3489_,
		_w3491_
	);
	LUT2 #(
		.INIT('h1)
	) name1984 (
		\TM0_pad ,
		_w3490_,
		_w3492_
	);
	LUT2 #(
		.INIT('h4)
	) name1985 (
		_w3491_,
		_w3492_,
		_w3493_
	);
	LUT2 #(
		.INIT('h2)
	) name1986 (
		_w3483_,
		_w3493_,
		_w3494_
	);
	LUT2 #(
		.INIT('h2)
	) name1987 (
		\TM0_pad ,
		\_2148__reg/NET0131 ,
		_w3495_
	);
	LUT2 #(
		.INIT('h2)
	) name1988 (
		\WX4700_reg/NET0131 ,
		\WX4764_reg/NET0131 ,
		_w3496_
	);
	LUT2 #(
		.INIT('h4)
	) name1989 (
		\WX4700_reg/NET0131 ,
		\WX4764_reg/NET0131 ,
		_w3497_
	);
	LUT2 #(
		.INIT('h1)
	) name1990 (
		_w3496_,
		_w3497_,
		_w3498_
	);
	LUT2 #(
		.INIT('h2)
	) name1991 (
		\WX4572_reg/NET0131 ,
		\WX4636_reg/NET0131 ,
		_w3499_
	);
	LUT2 #(
		.INIT('h4)
	) name1992 (
		\WX4572_reg/NET0131 ,
		\WX4636_reg/NET0131 ,
		_w3500_
	);
	LUT2 #(
		.INIT('h1)
	) name1993 (
		_w3499_,
		_w3500_,
		_w3501_
	);
	LUT2 #(
		.INIT('h4)
	) name1994 (
		_w3498_,
		_w3501_,
		_w3502_
	);
	LUT2 #(
		.INIT('h2)
	) name1995 (
		_w3498_,
		_w3501_,
		_w3503_
	);
	LUT2 #(
		.INIT('h1)
	) name1996 (
		\TM0_pad ,
		_w3502_,
		_w3504_
	);
	LUT2 #(
		.INIT('h4)
	) name1997 (
		_w3503_,
		_w3504_,
		_w3505_
	);
	LUT2 #(
		.INIT('h2)
	) name1998 (
		_w1976_,
		_w3495_,
		_w3506_
	);
	LUT2 #(
		.INIT('h4)
	) name1999 (
		_w3505_,
		_w3506_,
		_w3507_
	);
	LUT2 #(
		.INIT('h1)
	) name2000 (
		_w3494_,
		_w3507_,
		_w3508_
	);
	LUT2 #(
		.INIT('h2)
	) name2001 (
		_w2846_,
		_w3438_,
		_w3509_
	);
	LUT2 #(
		.INIT('h2)
	) name2002 (
		\TM0_pad ,
		\_2280__reg/NET0131 ,
		_w3510_
	);
	LUT2 #(
		.INIT('h2)
	) name2003 (
		\WX9864_reg/NET0131 ,
		\WX9928_reg/NET0131 ,
		_w3511_
	);
	LUT2 #(
		.INIT('h4)
	) name2004 (
		\WX9864_reg/NET0131 ,
		\WX9928_reg/NET0131 ,
		_w3512_
	);
	LUT2 #(
		.INIT('h1)
	) name2005 (
		_w3511_,
		_w3512_,
		_w3513_
	);
	LUT2 #(
		.INIT('h2)
	) name2006 (
		\WX9736_reg/NET0131 ,
		\WX9800_reg/NET0131 ,
		_w3514_
	);
	LUT2 #(
		.INIT('h4)
	) name2007 (
		\WX9736_reg/NET0131 ,
		\WX9800_reg/NET0131 ,
		_w3515_
	);
	LUT2 #(
		.INIT('h1)
	) name2008 (
		_w3514_,
		_w3515_,
		_w3516_
	);
	LUT2 #(
		.INIT('h4)
	) name2009 (
		_w3513_,
		_w3516_,
		_w3517_
	);
	LUT2 #(
		.INIT('h2)
	) name2010 (
		_w3513_,
		_w3516_,
		_w3518_
	);
	LUT2 #(
		.INIT('h1)
	) name2011 (
		\TM0_pad ,
		_w3517_,
		_w3519_
	);
	LUT2 #(
		.INIT('h4)
	) name2012 (
		_w3518_,
		_w3519_,
		_w3520_
	);
	LUT2 #(
		.INIT('h2)
	) name2013 (
		_w1976_,
		_w3510_,
		_w3521_
	);
	LUT2 #(
		.INIT('h4)
	) name2014 (
		_w3520_,
		_w3521_,
		_w3522_
	);
	LUT2 #(
		.INIT('h1)
	) name2015 (
		_w3509_,
		_w3522_,
		_w3523_
	);
	LUT2 #(
		.INIT('h2)
	) name2016 (
		_w2677_,
		_w3369_,
		_w3524_
	);
	LUT2 #(
		.INIT('h2)
	) name2017 (
		\TM0_pad ,
		\_2313__reg/NET0131 ,
		_w3525_
	);
	LUT2 #(
		.INIT('h2)
	) name2018 (
		\WX11155_reg/NET0131 ,
		\WX11219_reg/NET0131 ,
		_w3526_
	);
	LUT2 #(
		.INIT('h4)
	) name2019 (
		\WX11155_reg/NET0131 ,
		\WX11219_reg/NET0131 ,
		_w3527_
	);
	LUT2 #(
		.INIT('h1)
	) name2020 (
		_w3526_,
		_w3527_,
		_w3528_
	);
	LUT2 #(
		.INIT('h2)
	) name2021 (
		\WX11027_reg/NET0131 ,
		\WX11091_reg/NET0131 ,
		_w3529_
	);
	LUT2 #(
		.INIT('h4)
	) name2022 (
		\WX11027_reg/NET0131 ,
		\WX11091_reg/NET0131 ,
		_w3530_
	);
	LUT2 #(
		.INIT('h1)
	) name2023 (
		_w3529_,
		_w3530_,
		_w3531_
	);
	LUT2 #(
		.INIT('h4)
	) name2024 (
		_w3528_,
		_w3531_,
		_w3532_
	);
	LUT2 #(
		.INIT('h2)
	) name2025 (
		_w3528_,
		_w3531_,
		_w3533_
	);
	LUT2 #(
		.INIT('h1)
	) name2026 (
		\TM0_pad ,
		_w3532_,
		_w3534_
	);
	LUT2 #(
		.INIT('h4)
	) name2027 (
		_w3533_,
		_w3534_,
		_w3535_
	);
	LUT2 #(
		.INIT('h2)
	) name2028 (
		_w1976_,
		_w3525_,
		_w3536_
	);
	LUT2 #(
		.INIT('h4)
	) name2029 (
		_w3535_,
		_w3536_,
		_w3537_
	);
	LUT2 #(
		.INIT('h1)
	) name2030 (
		_w3524_,
		_w3537_,
		_w3538_
	);
	LUT2 #(
		.INIT('h8)
	) name2031 (
		\TM0_pad ,
		\_2131__reg/NET0131 ,
		_w3539_
	);
	LUT2 #(
		.INIT('h2)
	) name2032 (
		\WX3377_reg/NET0131 ,
		\WX3441_reg/NET0131 ,
		_w3540_
	);
	LUT2 #(
		.INIT('h4)
	) name2033 (
		\WX3377_reg/NET0131 ,
		\WX3441_reg/NET0131 ,
		_w3541_
	);
	LUT2 #(
		.INIT('h1)
	) name2034 (
		_w3540_,
		_w3541_,
		_w3542_
	);
	LUT2 #(
		.INIT('h2)
	) name2035 (
		\WX3313_reg/NET0131 ,
		_w3542_,
		_w3543_
	);
	LUT2 #(
		.INIT('h4)
	) name2036 (
		\WX3313_reg/NET0131 ,
		_w3542_,
		_w3544_
	);
	LUT2 #(
		.INIT('h1)
	) name2037 (
		_w3543_,
		_w3544_,
		_w3545_
	);
	LUT2 #(
		.INIT('h2)
	) name2038 (
		\TM1_pad ,
		\WX3249_reg/NET0131 ,
		_w3546_
	);
	LUT2 #(
		.INIT('h4)
	) name2039 (
		\TM1_pad ,
		\WX3249_reg/NET0131 ,
		_w3547_
	);
	LUT2 #(
		.INIT('h1)
	) name2040 (
		_w3546_,
		_w3547_,
		_w3548_
	);
	LUT2 #(
		.INIT('h4)
	) name2041 (
		_w3545_,
		_w3548_,
		_w3549_
	);
	LUT2 #(
		.INIT('h2)
	) name2042 (
		_w3545_,
		_w3548_,
		_w3550_
	);
	LUT2 #(
		.INIT('h1)
	) name2043 (
		\TM0_pad ,
		_w3549_,
		_w3551_
	);
	LUT2 #(
		.INIT('h4)
	) name2044 (
		_w3550_,
		_w3551_,
		_w3552_
	);
	LUT2 #(
		.INIT('h1)
	) name2045 (
		_w3539_,
		_w3552_,
		_w3553_
	);
	LUT2 #(
		.INIT('h2)
	) name2046 (
		_w1976_,
		_w3553_,
		_w3554_
	);
	LUT2 #(
		.INIT('h1)
	) name2047 (
		_w1714_,
		_w3308_,
		_w3555_
	);
	LUT2 #(
		.INIT('h2)
	) name2048 (
		_w1973_,
		_w3555_,
		_w3556_
	);
	LUT2 #(
		.INIT('h1)
	) name2049 (
		_w3554_,
		_w3556_,
		_w3557_
	);
	LUT2 #(
		.INIT('h2)
	) name2050 (
		_w2023_,
		_w3354_,
		_w3558_
	);
	LUT2 #(
		.INIT('h2)
	) name2051 (
		\TM0_pad ,
		\_2181__reg/NET0131 ,
		_w3559_
	);
	LUT2 #(
		.INIT('h2)
	) name2052 (
		\WX5991_reg/NET0131 ,
		\WX6055_reg/NET0131 ,
		_w3560_
	);
	LUT2 #(
		.INIT('h4)
	) name2053 (
		\WX5991_reg/NET0131 ,
		\WX6055_reg/NET0131 ,
		_w3561_
	);
	LUT2 #(
		.INIT('h1)
	) name2054 (
		_w3560_,
		_w3561_,
		_w3562_
	);
	LUT2 #(
		.INIT('h2)
	) name2055 (
		\WX5863_reg/NET0131 ,
		\WX5927_reg/NET0131 ,
		_w3563_
	);
	LUT2 #(
		.INIT('h4)
	) name2056 (
		\WX5863_reg/NET0131 ,
		\WX5927_reg/NET0131 ,
		_w3564_
	);
	LUT2 #(
		.INIT('h1)
	) name2057 (
		_w3563_,
		_w3564_,
		_w3565_
	);
	LUT2 #(
		.INIT('h4)
	) name2058 (
		_w3562_,
		_w3565_,
		_w3566_
	);
	LUT2 #(
		.INIT('h2)
	) name2059 (
		_w3562_,
		_w3565_,
		_w3567_
	);
	LUT2 #(
		.INIT('h1)
	) name2060 (
		\TM0_pad ,
		_w3566_,
		_w3568_
	);
	LUT2 #(
		.INIT('h4)
	) name2061 (
		_w3567_,
		_w3568_,
		_w3569_
	);
	LUT2 #(
		.INIT('h2)
	) name2062 (
		_w1976_,
		_w3559_,
		_w3570_
	);
	LUT2 #(
		.INIT('h4)
	) name2063 (
		_w3569_,
		_w3570_,
		_w3571_
	);
	LUT2 #(
		.INIT('h1)
	) name2064 (
		_w3558_,
		_w3571_,
		_w3572_
	);
	LUT2 #(
		.INIT('h2)
	) name2065 (
		_w3172_,
		_w3408_,
		_w3573_
	);
	LUT2 #(
		.INIT('h2)
	) name2066 (
		\TM0_pad ,
		\_2214__reg/NET0131 ,
		_w3574_
	);
	LUT2 #(
		.INIT('h2)
	) name2067 (
		\WX7282_reg/NET0131 ,
		\WX7346_reg/NET0131 ,
		_w3575_
	);
	LUT2 #(
		.INIT('h4)
	) name2068 (
		\WX7282_reg/NET0131 ,
		\WX7346_reg/NET0131 ,
		_w3576_
	);
	LUT2 #(
		.INIT('h1)
	) name2069 (
		_w3575_,
		_w3576_,
		_w3577_
	);
	LUT2 #(
		.INIT('h2)
	) name2070 (
		\WX7154_reg/NET0131 ,
		\WX7218_reg/NET0131 ,
		_w3578_
	);
	LUT2 #(
		.INIT('h4)
	) name2071 (
		\WX7154_reg/NET0131 ,
		\WX7218_reg/NET0131 ,
		_w3579_
	);
	LUT2 #(
		.INIT('h1)
	) name2072 (
		_w3578_,
		_w3579_,
		_w3580_
	);
	LUT2 #(
		.INIT('h4)
	) name2073 (
		_w3577_,
		_w3580_,
		_w3581_
	);
	LUT2 #(
		.INIT('h2)
	) name2074 (
		_w3577_,
		_w3580_,
		_w3582_
	);
	LUT2 #(
		.INIT('h1)
	) name2075 (
		\TM0_pad ,
		_w3581_,
		_w3583_
	);
	LUT2 #(
		.INIT('h4)
	) name2076 (
		_w3582_,
		_w3583_,
		_w3584_
	);
	LUT2 #(
		.INIT('h2)
	) name2077 (
		_w1976_,
		_w3574_,
		_w3585_
	);
	LUT2 #(
		.INIT('h4)
	) name2078 (
		_w3584_,
		_w3585_,
		_w3586_
	);
	LUT2 #(
		.INIT('h1)
	) name2079 (
		_w3573_,
		_w3586_,
		_w3587_
	);
	LUT2 #(
		.INIT('h2)
	) name2080 (
		_w3011_,
		_w3423_,
		_w3588_
	);
	LUT2 #(
		.INIT('h2)
	) name2081 (
		\TM0_pad ,
		\_2247__reg/NET0131 ,
		_w3589_
	);
	LUT2 #(
		.INIT('h2)
	) name2082 (
		\WX8573_reg/NET0131 ,
		\WX8637_reg/NET0131 ,
		_w3590_
	);
	LUT2 #(
		.INIT('h4)
	) name2083 (
		\WX8573_reg/NET0131 ,
		\WX8637_reg/NET0131 ,
		_w3591_
	);
	LUT2 #(
		.INIT('h1)
	) name2084 (
		_w3590_,
		_w3591_,
		_w3592_
	);
	LUT2 #(
		.INIT('h2)
	) name2085 (
		\WX8445_reg/NET0131 ,
		\WX8509_reg/NET0131 ,
		_w3593_
	);
	LUT2 #(
		.INIT('h4)
	) name2086 (
		\WX8445_reg/NET0131 ,
		\WX8509_reg/NET0131 ,
		_w3594_
	);
	LUT2 #(
		.INIT('h1)
	) name2087 (
		_w3593_,
		_w3594_,
		_w3595_
	);
	LUT2 #(
		.INIT('h4)
	) name2088 (
		_w3592_,
		_w3595_,
		_w3596_
	);
	LUT2 #(
		.INIT('h2)
	) name2089 (
		_w3592_,
		_w3595_,
		_w3597_
	);
	LUT2 #(
		.INIT('h1)
	) name2090 (
		\TM0_pad ,
		_w3596_,
		_w3598_
	);
	LUT2 #(
		.INIT('h4)
	) name2091 (
		_w3597_,
		_w3598_,
		_w3599_
	);
	LUT2 #(
		.INIT('h2)
	) name2092 (
		_w1976_,
		_w3589_,
		_w3600_
	);
	LUT2 #(
		.INIT('h4)
	) name2093 (
		_w3599_,
		_w3600_,
		_w3601_
	);
	LUT2 #(
		.INIT('h1)
	) name2094 (
		_w3588_,
		_w3601_,
		_w3602_
	);
	LUT2 #(
		.INIT('h1)
	) name2095 (
		\TM0_pad ,
		_w1691_,
		_w3603_
	);
	LUT2 #(
		.INIT('h1)
	) name2096 (
		_w1682_,
		_w3603_,
		_w3604_
	);
	LUT2 #(
		.INIT('h2)
	) name2097 (
		_w1973_,
		_w3604_,
		_w3605_
	);
	LUT2 #(
		.INIT('h8)
	) name2098 (
		\TM0_pad ,
		\_2097__reg/NET0131 ,
		_w3606_
	);
	LUT2 #(
		.INIT('h2)
	) name2099 (
		\WX2088_reg/NET0131 ,
		\WX2152_reg/NET0131 ,
		_w3607_
	);
	LUT2 #(
		.INIT('h4)
	) name2100 (
		\WX2088_reg/NET0131 ,
		\WX2152_reg/NET0131 ,
		_w3608_
	);
	LUT2 #(
		.INIT('h1)
	) name2101 (
		_w3607_,
		_w3608_,
		_w3609_
	);
	LUT2 #(
		.INIT('h2)
	) name2102 (
		\WX2024_reg/NET0131 ,
		_w3609_,
		_w3610_
	);
	LUT2 #(
		.INIT('h4)
	) name2103 (
		\WX2024_reg/NET0131 ,
		_w3609_,
		_w3611_
	);
	LUT2 #(
		.INIT('h1)
	) name2104 (
		_w3610_,
		_w3611_,
		_w3612_
	);
	LUT2 #(
		.INIT('h2)
	) name2105 (
		\TM1_pad ,
		\WX1960_reg/NET0131 ,
		_w3613_
	);
	LUT2 #(
		.INIT('h4)
	) name2106 (
		\TM1_pad ,
		\WX1960_reg/NET0131 ,
		_w3614_
	);
	LUT2 #(
		.INIT('h1)
	) name2107 (
		_w3613_,
		_w3614_,
		_w3615_
	);
	LUT2 #(
		.INIT('h4)
	) name2108 (
		_w3612_,
		_w3615_,
		_w3616_
	);
	LUT2 #(
		.INIT('h2)
	) name2109 (
		_w3612_,
		_w3615_,
		_w3617_
	);
	LUT2 #(
		.INIT('h1)
	) name2110 (
		\TM0_pad ,
		_w3616_,
		_w3618_
	);
	LUT2 #(
		.INIT('h4)
	) name2111 (
		_w3617_,
		_w3618_,
		_w3619_
	);
	LUT2 #(
		.INIT('h1)
	) name2112 (
		_w3606_,
		_w3619_,
		_w3620_
	);
	LUT2 #(
		.INIT('h2)
	) name2113 (
		_w1976_,
		_w3620_,
		_w3621_
	);
	LUT2 #(
		.INIT('h1)
	) name2114 (
		_w3605_,
		_w3621_,
		_w3622_
	);
	LUT2 #(
		.INIT('h2)
	) name2115 (
		\WX11135_reg/NET0131 ,
		\WX11199_reg/NET0131 ,
		_w3623_
	);
	LUT2 #(
		.INIT('h4)
	) name2116 (
		\WX11135_reg/NET0131 ,
		\WX11199_reg/NET0131 ,
		_w3624_
	);
	LUT2 #(
		.INIT('h1)
	) name2117 (
		_w3623_,
		_w3624_,
		_w3625_
	);
	LUT2 #(
		.INIT('h2)
	) name2118 (
		\WX11071_reg/NET0131 ,
		_w3625_,
		_w3626_
	);
	LUT2 #(
		.INIT('h4)
	) name2119 (
		\WX11071_reg/NET0131 ,
		_w3625_,
		_w3627_
	);
	LUT2 #(
		.INIT('h1)
	) name2120 (
		_w3626_,
		_w3627_,
		_w3628_
	);
	LUT2 #(
		.INIT('h2)
	) name2121 (
		\TM1_pad ,
		\WX11007_reg/NET0131 ,
		_w3629_
	);
	LUT2 #(
		.INIT('h4)
	) name2122 (
		\TM1_pad ,
		\WX11007_reg/NET0131 ,
		_w3630_
	);
	LUT2 #(
		.INIT('h1)
	) name2123 (
		_w3629_,
		_w3630_,
		_w3631_
	);
	LUT2 #(
		.INIT('h4)
	) name2124 (
		_w3628_,
		_w3631_,
		_w3632_
	);
	LUT2 #(
		.INIT('h2)
	) name2125 (
		_w3628_,
		_w3631_,
		_w3633_
	);
	LUT2 #(
		.INIT('h1)
	) name2126 (
		\TM0_pad ,
		_w3632_,
		_w3634_
	);
	LUT2 #(
		.INIT('h4)
	) name2127 (
		_w3633_,
		_w3634_,
		_w3635_
	);
	LUT2 #(
		.INIT('h1)
	) name2128 (
		_w1714_,
		_w3635_,
		_w3636_
	);
	LUT2 #(
		.INIT('h2)
	) name2129 (
		_w1973_,
		_w3636_,
		_w3637_
	);
	LUT2 #(
		.INIT('h1)
	) name2130 (
		\DATA_0_22_pad ,
		\TM0_pad ,
		_w3638_
	);
	LUT2 #(
		.INIT('h2)
	) name2131 (
		\TM0_pad ,
		\_2355__reg/NET0131 ,
		_w3639_
	);
	LUT2 #(
		.INIT('h2)
	) name2132 (
		_w1976_,
		_w3638_,
		_w3640_
	);
	LUT2 #(
		.INIT('h4)
	) name2133 (
		_w3639_,
		_w3640_,
		_w3641_
	);
	LUT2 #(
		.INIT('h1)
	) name2134 (
		_w3637_,
		_w3641_,
		_w3642_
	);
	LUT2 #(
		.INIT('h8)
	) name2135 (
		RESET_pad,
		\WX10845_reg/NET0131 ,
		_w3643_
	);
	LUT2 #(
		.INIT('h4)
	) name2136 (
		_w1920_,
		_w1973_,
		_w3644_
	);
	LUT2 #(
		.INIT('h2)
	) name2137 (
		\WX3409_reg/NET0131 ,
		\WX3473_reg/NET0131 ,
		_w3645_
	);
	LUT2 #(
		.INIT('h4)
	) name2138 (
		\WX3409_reg/NET0131 ,
		\WX3473_reg/NET0131 ,
		_w3646_
	);
	LUT2 #(
		.INIT('h1)
	) name2139 (
		_w3645_,
		_w3646_,
		_w3647_
	);
	LUT2 #(
		.INIT('h2)
	) name2140 (
		\WX3281_reg/NET0131 ,
		\WX3345_reg/NET0131 ,
		_w3648_
	);
	LUT2 #(
		.INIT('h4)
	) name2141 (
		\WX3281_reg/NET0131 ,
		\WX3345_reg/NET0131 ,
		_w3649_
	);
	LUT2 #(
		.INIT('h1)
	) name2142 (
		_w3648_,
		_w3649_,
		_w3650_
	);
	LUT2 #(
		.INIT('h4)
	) name2143 (
		_w3647_,
		_w3650_,
		_w3651_
	);
	LUT2 #(
		.INIT('h2)
	) name2144 (
		_w3647_,
		_w3650_,
		_w3652_
	);
	LUT2 #(
		.INIT('h1)
	) name2145 (
		\TM0_pad ,
		_w3651_,
		_w3653_
	);
	LUT2 #(
		.INIT('h4)
	) name2146 (
		_w3652_,
		_w3653_,
		_w3654_
	);
	LUT2 #(
		.INIT('h2)
	) name2147 (
		_w3644_,
		_w3654_,
		_w3655_
	);
	LUT2 #(
		.INIT('h2)
	) name2148 (
		\TM0_pad ,
		\_2147__reg/NET0131 ,
		_w3656_
	);
	LUT2 #(
		.INIT('h2)
	) name2149 (
		\WX4702_reg/NET0131 ,
		\WX4766_reg/NET0131 ,
		_w3657_
	);
	LUT2 #(
		.INIT('h4)
	) name2150 (
		\WX4702_reg/NET0131 ,
		\WX4766_reg/NET0131 ,
		_w3658_
	);
	LUT2 #(
		.INIT('h1)
	) name2151 (
		_w3657_,
		_w3658_,
		_w3659_
	);
	LUT2 #(
		.INIT('h2)
	) name2152 (
		\WX4574_reg/NET0131 ,
		\WX4638_reg/NET0131 ,
		_w3660_
	);
	LUT2 #(
		.INIT('h4)
	) name2153 (
		\WX4574_reg/NET0131 ,
		\WX4638_reg/NET0131 ,
		_w3661_
	);
	LUT2 #(
		.INIT('h1)
	) name2154 (
		_w3660_,
		_w3661_,
		_w3662_
	);
	LUT2 #(
		.INIT('h4)
	) name2155 (
		_w3659_,
		_w3662_,
		_w3663_
	);
	LUT2 #(
		.INIT('h2)
	) name2156 (
		_w3659_,
		_w3662_,
		_w3664_
	);
	LUT2 #(
		.INIT('h1)
	) name2157 (
		\TM0_pad ,
		_w3663_,
		_w3665_
	);
	LUT2 #(
		.INIT('h4)
	) name2158 (
		_w3664_,
		_w3665_,
		_w3666_
	);
	LUT2 #(
		.INIT('h2)
	) name2159 (
		_w1976_,
		_w3656_,
		_w3667_
	);
	LUT2 #(
		.INIT('h4)
	) name2160 (
		_w3666_,
		_w3667_,
		_w3668_
	);
	LUT2 #(
		.INIT('h1)
	) name2161 (
		_w3655_,
		_w3668_,
		_w3669_
	);
	LUT2 #(
		.INIT('h2)
	) name2162 (
		_w3011_,
		_w3599_,
		_w3670_
	);
	LUT2 #(
		.INIT('h2)
	) name2163 (
		\TM0_pad ,
		\_2279__reg/NET0131 ,
		_w3671_
	);
	LUT2 #(
		.INIT('h2)
	) name2164 (
		\WX9866_reg/NET0131 ,
		\WX9930_reg/NET0131 ,
		_w3672_
	);
	LUT2 #(
		.INIT('h4)
	) name2165 (
		\WX9866_reg/NET0131 ,
		\WX9930_reg/NET0131 ,
		_w3673_
	);
	LUT2 #(
		.INIT('h1)
	) name2166 (
		_w3672_,
		_w3673_,
		_w3674_
	);
	LUT2 #(
		.INIT('h2)
	) name2167 (
		\WX9738_reg/NET0131 ,
		\WX9802_reg/NET0131 ,
		_w3675_
	);
	LUT2 #(
		.INIT('h4)
	) name2168 (
		\WX9738_reg/NET0131 ,
		\WX9802_reg/NET0131 ,
		_w3676_
	);
	LUT2 #(
		.INIT('h1)
	) name2169 (
		_w3675_,
		_w3676_,
		_w3677_
	);
	LUT2 #(
		.INIT('h4)
	) name2170 (
		_w3674_,
		_w3677_,
		_w3678_
	);
	LUT2 #(
		.INIT('h2)
	) name2171 (
		_w3674_,
		_w3677_,
		_w3679_
	);
	LUT2 #(
		.INIT('h1)
	) name2172 (
		\TM0_pad ,
		_w3678_,
		_w3680_
	);
	LUT2 #(
		.INIT('h4)
	) name2173 (
		_w3679_,
		_w3680_,
		_w3681_
	);
	LUT2 #(
		.INIT('h2)
	) name2174 (
		_w1976_,
		_w3671_,
		_w3682_
	);
	LUT2 #(
		.INIT('h4)
	) name2175 (
		_w3681_,
		_w3682_,
		_w3683_
	);
	LUT2 #(
		.INIT('h1)
	) name2176 (
		_w3670_,
		_w3683_,
		_w3684_
	);
	LUT2 #(
		.INIT('h2)
	) name2177 (
		_w2846_,
		_w3520_,
		_w3685_
	);
	LUT2 #(
		.INIT('h2)
	) name2178 (
		\TM0_pad ,
		\_2312__reg/NET0131 ,
		_w3686_
	);
	LUT2 #(
		.INIT('h2)
	) name2179 (
		\WX11157_reg/NET0131 ,
		\WX11221_reg/NET0131 ,
		_w3687_
	);
	LUT2 #(
		.INIT('h4)
	) name2180 (
		\WX11157_reg/NET0131 ,
		\WX11221_reg/NET0131 ,
		_w3688_
	);
	LUT2 #(
		.INIT('h1)
	) name2181 (
		_w3687_,
		_w3688_,
		_w3689_
	);
	LUT2 #(
		.INIT('h2)
	) name2182 (
		\WX11029_reg/NET0131 ,
		\WX11093_reg/NET0131 ,
		_w3690_
	);
	LUT2 #(
		.INIT('h4)
	) name2183 (
		\WX11029_reg/NET0131 ,
		\WX11093_reg/NET0131 ,
		_w3691_
	);
	LUT2 #(
		.INIT('h1)
	) name2184 (
		_w3690_,
		_w3691_,
		_w3692_
	);
	LUT2 #(
		.INIT('h4)
	) name2185 (
		_w3689_,
		_w3692_,
		_w3693_
	);
	LUT2 #(
		.INIT('h2)
	) name2186 (
		_w3689_,
		_w3692_,
		_w3694_
	);
	LUT2 #(
		.INIT('h1)
	) name2187 (
		\TM0_pad ,
		_w3693_,
		_w3695_
	);
	LUT2 #(
		.INIT('h4)
	) name2188 (
		_w3694_,
		_w3695_,
		_w3696_
	);
	LUT2 #(
		.INIT('h2)
	) name2189 (
		_w1976_,
		_w3686_,
		_w3697_
	);
	LUT2 #(
		.INIT('h4)
	) name2190 (
		_w3696_,
		_w3697_,
		_w3698_
	);
	LUT2 #(
		.INIT('h1)
	) name2191 (
		_w3685_,
		_w3698_,
		_w3699_
	);
	LUT2 #(
		.INIT('h8)
	) name2192 (
		\TM0_pad ,
		\_2130__reg/NET0131 ,
		_w3700_
	);
	LUT2 #(
		.INIT('h2)
	) name2193 (
		\WX3379_reg/NET0131 ,
		\WX3443_reg/NET0131 ,
		_w3701_
	);
	LUT2 #(
		.INIT('h4)
	) name2194 (
		\WX3379_reg/NET0131 ,
		\WX3443_reg/NET0131 ,
		_w3702_
	);
	LUT2 #(
		.INIT('h1)
	) name2195 (
		_w3701_,
		_w3702_,
		_w3703_
	);
	LUT2 #(
		.INIT('h2)
	) name2196 (
		\WX3315_reg/NET0131 ,
		_w3703_,
		_w3704_
	);
	LUT2 #(
		.INIT('h4)
	) name2197 (
		\WX3315_reg/NET0131 ,
		_w3703_,
		_w3705_
	);
	LUT2 #(
		.INIT('h1)
	) name2198 (
		_w3704_,
		_w3705_,
		_w3706_
	);
	LUT2 #(
		.INIT('h2)
	) name2199 (
		\TM1_pad ,
		\WX3251_reg/NET0131 ,
		_w3707_
	);
	LUT2 #(
		.INIT('h4)
	) name2200 (
		\TM1_pad ,
		\WX3251_reg/NET0131 ,
		_w3708_
	);
	LUT2 #(
		.INIT('h1)
	) name2201 (
		_w3707_,
		_w3708_,
		_w3709_
	);
	LUT2 #(
		.INIT('h4)
	) name2202 (
		_w3706_,
		_w3709_,
		_w3710_
	);
	LUT2 #(
		.INIT('h2)
	) name2203 (
		_w3706_,
		_w3709_,
		_w3711_
	);
	LUT2 #(
		.INIT('h1)
	) name2204 (
		\TM0_pad ,
		_w3710_,
		_w3712_
	);
	LUT2 #(
		.INIT('h4)
	) name2205 (
		_w3711_,
		_w3712_,
		_w3713_
	);
	LUT2 #(
		.INIT('h1)
	) name2206 (
		_w3700_,
		_w3713_,
		_w3714_
	);
	LUT2 #(
		.INIT('h2)
	) name2207 (
		_w1976_,
		_w3714_,
		_w3715_
	);
	LUT2 #(
		.INIT('h1)
	) name2208 (
		_w1698_,
		_w3458_,
		_w3716_
	);
	LUT2 #(
		.INIT('h2)
	) name2209 (
		_w1973_,
		_w3716_,
		_w3717_
	);
	LUT2 #(
		.INIT('h1)
	) name2210 (
		_w3715_,
		_w3717_,
		_w3718_
	);
	LUT2 #(
		.INIT('h2)
	) name2211 (
		_w3483_,
		_w3505_,
		_w3719_
	);
	LUT2 #(
		.INIT('h2)
	) name2212 (
		\TM0_pad ,
		\_2180__reg/NET0131 ,
		_w3720_
	);
	LUT2 #(
		.INIT('h2)
	) name2213 (
		\WX5993_reg/NET0131 ,
		\WX6057_reg/NET0131 ,
		_w3721_
	);
	LUT2 #(
		.INIT('h4)
	) name2214 (
		\WX5993_reg/NET0131 ,
		\WX6057_reg/NET0131 ,
		_w3722_
	);
	LUT2 #(
		.INIT('h1)
	) name2215 (
		_w3721_,
		_w3722_,
		_w3723_
	);
	LUT2 #(
		.INIT('h2)
	) name2216 (
		\WX5865_reg/NET0131 ,
		\WX5929_reg/NET0131 ,
		_w3724_
	);
	LUT2 #(
		.INIT('h4)
	) name2217 (
		\WX5865_reg/NET0131 ,
		\WX5929_reg/NET0131 ,
		_w3725_
	);
	LUT2 #(
		.INIT('h1)
	) name2218 (
		_w3724_,
		_w3725_,
		_w3726_
	);
	LUT2 #(
		.INIT('h4)
	) name2219 (
		_w3723_,
		_w3726_,
		_w3727_
	);
	LUT2 #(
		.INIT('h2)
	) name2220 (
		_w3723_,
		_w3726_,
		_w3728_
	);
	LUT2 #(
		.INIT('h1)
	) name2221 (
		\TM0_pad ,
		_w3727_,
		_w3729_
	);
	LUT2 #(
		.INIT('h4)
	) name2222 (
		_w3728_,
		_w3729_,
		_w3730_
	);
	LUT2 #(
		.INIT('h2)
	) name2223 (
		_w1976_,
		_w3720_,
		_w3731_
	);
	LUT2 #(
		.INIT('h4)
	) name2224 (
		_w3730_,
		_w3731_,
		_w3732_
	);
	LUT2 #(
		.INIT('h1)
	) name2225 (
		_w3719_,
		_w3732_,
		_w3733_
	);
	LUT2 #(
		.INIT('h2)
	) name2226 (
		_w2023_,
		_w3569_,
		_w3734_
	);
	LUT2 #(
		.INIT('h2)
	) name2227 (
		\TM0_pad ,
		\_2213__reg/NET0131 ,
		_w3735_
	);
	LUT2 #(
		.INIT('h2)
	) name2228 (
		\WX7284_reg/NET0131 ,
		\WX7348_reg/NET0131 ,
		_w3736_
	);
	LUT2 #(
		.INIT('h4)
	) name2229 (
		\WX7284_reg/NET0131 ,
		\WX7348_reg/NET0131 ,
		_w3737_
	);
	LUT2 #(
		.INIT('h1)
	) name2230 (
		_w3736_,
		_w3737_,
		_w3738_
	);
	LUT2 #(
		.INIT('h2)
	) name2231 (
		\WX7156_reg/NET0131 ,
		\WX7220_reg/NET0131 ,
		_w3739_
	);
	LUT2 #(
		.INIT('h4)
	) name2232 (
		\WX7156_reg/NET0131 ,
		\WX7220_reg/NET0131 ,
		_w3740_
	);
	LUT2 #(
		.INIT('h1)
	) name2233 (
		_w3739_,
		_w3740_,
		_w3741_
	);
	LUT2 #(
		.INIT('h4)
	) name2234 (
		_w3738_,
		_w3741_,
		_w3742_
	);
	LUT2 #(
		.INIT('h2)
	) name2235 (
		_w3738_,
		_w3741_,
		_w3743_
	);
	LUT2 #(
		.INIT('h1)
	) name2236 (
		\TM0_pad ,
		_w3742_,
		_w3744_
	);
	LUT2 #(
		.INIT('h4)
	) name2237 (
		_w3743_,
		_w3744_,
		_w3745_
	);
	LUT2 #(
		.INIT('h2)
	) name2238 (
		_w1976_,
		_w3735_,
		_w3746_
	);
	LUT2 #(
		.INIT('h4)
	) name2239 (
		_w3745_,
		_w3746_,
		_w3747_
	);
	LUT2 #(
		.INIT('h1)
	) name2240 (
		_w3734_,
		_w3747_,
		_w3748_
	);
	LUT2 #(
		.INIT('h2)
	) name2241 (
		_w3172_,
		_w3584_,
		_w3749_
	);
	LUT2 #(
		.INIT('h2)
	) name2242 (
		\TM0_pad ,
		\_2246__reg/NET0131 ,
		_w3750_
	);
	LUT2 #(
		.INIT('h2)
	) name2243 (
		\WX8575_reg/NET0131 ,
		\WX8639_reg/NET0131 ,
		_w3751_
	);
	LUT2 #(
		.INIT('h4)
	) name2244 (
		\WX8575_reg/NET0131 ,
		\WX8639_reg/NET0131 ,
		_w3752_
	);
	LUT2 #(
		.INIT('h1)
	) name2245 (
		_w3751_,
		_w3752_,
		_w3753_
	);
	LUT2 #(
		.INIT('h2)
	) name2246 (
		\WX8447_reg/NET0131 ,
		\WX8511_reg/NET0131 ,
		_w3754_
	);
	LUT2 #(
		.INIT('h4)
	) name2247 (
		\WX8447_reg/NET0131 ,
		\WX8511_reg/NET0131 ,
		_w3755_
	);
	LUT2 #(
		.INIT('h1)
	) name2248 (
		_w3754_,
		_w3755_,
		_w3756_
	);
	LUT2 #(
		.INIT('h4)
	) name2249 (
		_w3753_,
		_w3756_,
		_w3757_
	);
	LUT2 #(
		.INIT('h2)
	) name2250 (
		_w3753_,
		_w3756_,
		_w3758_
	);
	LUT2 #(
		.INIT('h1)
	) name2251 (
		\TM0_pad ,
		_w3757_,
		_w3759_
	);
	LUT2 #(
		.INIT('h4)
	) name2252 (
		_w3758_,
		_w3759_,
		_w3760_
	);
	LUT2 #(
		.INIT('h2)
	) name2253 (
		_w1976_,
		_w3750_,
		_w3761_
	);
	LUT2 #(
		.INIT('h4)
	) name2254 (
		_w3760_,
		_w3761_,
		_w3762_
	);
	LUT2 #(
		.INIT('h1)
	) name2255 (
		_w3749_,
		_w3762_,
		_w3763_
	);
	LUT2 #(
		.INIT('h1)
	) name2256 (
		\TM0_pad ,
		_w1662_,
		_w3764_
	);
	LUT2 #(
		.INIT('h1)
	) name2257 (
		_w1653_,
		_w3764_,
		_w3765_
	);
	LUT2 #(
		.INIT('h2)
	) name2258 (
		_w1973_,
		_w3765_,
		_w3766_
	);
	LUT2 #(
		.INIT('h8)
	) name2259 (
		\TM0_pad ,
		\_2096__reg/NET0131 ,
		_w3767_
	);
	LUT2 #(
		.INIT('h2)
	) name2260 (
		\WX2090_reg/NET0131 ,
		\WX2154_reg/NET0131 ,
		_w3768_
	);
	LUT2 #(
		.INIT('h4)
	) name2261 (
		\WX2090_reg/NET0131 ,
		\WX2154_reg/NET0131 ,
		_w3769_
	);
	LUT2 #(
		.INIT('h1)
	) name2262 (
		_w3768_,
		_w3769_,
		_w3770_
	);
	LUT2 #(
		.INIT('h2)
	) name2263 (
		\WX2026_reg/NET0131 ,
		_w3770_,
		_w3771_
	);
	LUT2 #(
		.INIT('h4)
	) name2264 (
		\WX2026_reg/NET0131 ,
		_w3770_,
		_w3772_
	);
	LUT2 #(
		.INIT('h1)
	) name2265 (
		_w3771_,
		_w3772_,
		_w3773_
	);
	LUT2 #(
		.INIT('h2)
	) name2266 (
		\TM1_pad ,
		\WX1962_reg/NET0131 ,
		_w3774_
	);
	LUT2 #(
		.INIT('h4)
	) name2267 (
		\TM1_pad ,
		\WX1962_reg/NET0131 ,
		_w3775_
	);
	LUT2 #(
		.INIT('h1)
	) name2268 (
		_w3774_,
		_w3775_,
		_w3776_
	);
	LUT2 #(
		.INIT('h4)
	) name2269 (
		_w3773_,
		_w3776_,
		_w3777_
	);
	LUT2 #(
		.INIT('h2)
	) name2270 (
		_w3773_,
		_w3776_,
		_w3778_
	);
	LUT2 #(
		.INIT('h1)
	) name2271 (
		\TM0_pad ,
		_w3777_,
		_w3779_
	);
	LUT2 #(
		.INIT('h4)
	) name2272 (
		_w3778_,
		_w3779_,
		_w3780_
	);
	LUT2 #(
		.INIT('h1)
	) name2273 (
		_w3767_,
		_w3780_,
		_w3781_
	);
	LUT2 #(
		.INIT('h2)
	) name2274 (
		_w1976_,
		_w3781_,
		_w3782_
	);
	LUT2 #(
		.INIT('h1)
	) name2275 (
		_w3766_,
		_w3782_,
		_w3783_
	);
	LUT2 #(
		.INIT('h2)
	) name2276 (
		\WX11137_reg/NET0131 ,
		\WX11201_reg/NET0131 ,
		_w3784_
	);
	LUT2 #(
		.INIT('h4)
	) name2277 (
		\WX11137_reg/NET0131 ,
		\WX11201_reg/NET0131 ,
		_w3785_
	);
	LUT2 #(
		.INIT('h1)
	) name2278 (
		_w3784_,
		_w3785_,
		_w3786_
	);
	LUT2 #(
		.INIT('h2)
	) name2279 (
		\WX11073_reg/NET0131 ,
		_w3786_,
		_w3787_
	);
	LUT2 #(
		.INIT('h4)
	) name2280 (
		\WX11073_reg/NET0131 ,
		_w3786_,
		_w3788_
	);
	LUT2 #(
		.INIT('h1)
	) name2281 (
		_w3787_,
		_w3788_,
		_w3789_
	);
	LUT2 #(
		.INIT('h2)
	) name2282 (
		\TM1_pad ,
		\WX11009_reg/NET0131 ,
		_w3790_
	);
	LUT2 #(
		.INIT('h4)
	) name2283 (
		\TM1_pad ,
		\WX11009_reg/NET0131 ,
		_w3791_
	);
	LUT2 #(
		.INIT('h1)
	) name2284 (
		_w3790_,
		_w3791_,
		_w3792_
	);
	LUT2 #(
		.INIT('h4)
	) name2285 (
		_w3789_,
		_w3792_,
		_w3793_
	);
	LUT2 #(
		.INIT('h2)
	) name2286 (
		_w3789_,
		_w3792_,
		_w3794_
	);
	LUT2 #(
		.INIT('h1)
	) name2287 (
		\TM0_pad ,
		_w3793_,
		_w3795_
	);
	LUT2 #(
		.INIT('h4)
	) name2288 (
		_w3794_,
		_w3795_,
		_w3796_
	);
	LUT2 #(
		.INIT('h1)
	) name2289 (
		_w1698_,
		_w3796_,
		_w3797_
	);
	LUT2 #(
		.INIT('h2)
	) name2290 (
		_w1973_,
		_w3797_,
		_w3798_
	);
	LUT2 #(
		.INIT('h1)
	) name2291 (
		\DATA_0_21_pad ,
		\TM0_pad ,
		_w3799_
	);
	LUT2 #(
		.INIT('h2)
	) name2292 (
		\TM0_pad ,
		\_2354__reg/NET0131 ,
		_w3800_
	);
	LUT2 #(
		.INIT('h2)
	) name2293 (
		_w1976_,
		_w3799_,
		_w3801_
	);
	LUT2 #(
		.INIT('h4)
	) name2294 (
		_w3800_,
		_w3801_,
		_w3802_
	);
	LUT2 #(
		.INIT('h1)
	) name2295 (
		_w3798_,
		_w3802_,
		_w3803_
	);
	LUT2 #(
		.INIT('h8)
	) name2296 (
		RESET_pad,
		\WX10847_reg/NET0131 ,
		_w3804_
	);
	LUT2 #(
		.INIT('h4)
	) name2297 (
		_w1907_,
		_w1973_,
		_w3805_
	);
	LUT2 #(
		.INIT('h2)
	) name2298 (
		\WX3411_reg/NET0131 ,
		\WX3475_reg/NET0131 ,
		_w3806_
	);
	LUT2 #(
		.INIT('h4)
	) name2299 (
		\WX3411_reg/NET0131 ,
		\WX3475_reg/NET0131 ,
		_w3807_
	);
	LUT2 #(
		.INIT('h1)
	) name2300 (
		_w3806_,
		_w3807_,
		_w3808_
	);
	LUT2 #(
		.INIT('h2)
	) name2301 (
		\WX3283_reg/NET0131 ,
		\WX3347_reg/NET0131 ,
		_w3809_
	);
	LUT2 #(
		.INIT('h4)
	) name2302 (
		\WX3283_reg/NET0131 ,
		\WX3347_reg/NET0131 ,
		_w3810_
	);
	LUT2 #(
		.INIT('h1)
	) name2303 (
		_w3809_,
		_w3810_,
		_w3811_
	);
	LUT2 #(
		.INIT('h4)
	) name2304 (
		_w3808_,
		_w3811_,
		_w3812_
	);
	LUT2 #(
		.INIT('h2)
	) name2305 (
		_w3808_,
		_w3811_,
		_w3813_
	);
	LUT2 #(
		.INIT('h1)
	) name2306 (
		\TM0_pad ,
		_w3812_,
		_w3814_
	);
	LUT2 #(
		.INIT('h4)
	) name2307 (
		_w3813_,
		_w3814_,
		_w3815_
	);
	LUT2 #(
		.INIT('h2)
	) name2308 (
		_w3805_,
		_w3815_,
		_w3816_
	);
	LUT2 #(
		.INIT('h2)
	) name2309 (
		\TM0_pad ,
		\_2146__reg/NET0131 ,
		_w3817_
	);
	LUT2 #(
		.INIT('h2)
	) name2310 (
		\WX4704_reg/NET0131 ,
		\WX4768_reg/NET0131 ,
		_w3818_
	);
	LUT2 #(
		.INIT('h4)
	) name2311 (
		\WX4704_reg/NET0131 ,
		\WX4768_reg/NET0131 ,
		_w3819_
	);
	LUT2 #(
		.INIT('h1)
	) name2312 (
		_w3818_,
		_w3819_,
		_w3820_
	);
	LUT2 #(
		.INIT('h2)
	) name2313 (
		\WX4576_reg/NET0131 ,
		\WX4640_reg/NET0131 ,
		_w3821_
	);
	LUT2 #(
		.INIT('h4)
	) name2314 (
		\WX4576_reg/NET0131 ,
		\WX4640_reg/NET0131 ,
		_w3822_
	);
	LUT2 #(
		.INIT('h1)
	) name2315 (
		_w3821_,
		_w3822_,
		_w3823_
	);
	LUT2 #(
		.INIT('h4)
	) name2316 (
		_w3820_,
		_w3823_,
		_w3824_
	);
	LUT2 #(
		.INIT('h2)
	) name2317 (
		_w3820_,
		_w3823_,
		_w3825_
	);
	LUT2 #(
		.INIT('h1)
	) name2318 (
		\TM0_pad ,
		_w3824_,
		_w3826_
	);
	LUT2 #(
		.INIT('h4)
	) name2319 (
		_w3825_,
		_w3826_,
		_w3827_
	);
	LUT2 #(
		.INIT('h2)
	) name2320 (
		_w1976_,
		_w3817_,
		_w3828_
	);
	LUT2 #(
		.INIT('h4)
	) name2321 (
		_w3827_,
		_w3828_,
		_w3829_
	);
	LUT2 #(
		.INIT('h1)
	) name2322 (
		_w3816_,
		_w3829_,
		_w3830_
	);
	LUT2 #(
		.INIT('h2)
	) name2323 (
		_w3172_,
		_w3760_,
		_w3831_
	);
	LUT2 #(
		.INIT('h2)
	) name2324 (
		\TM0_pad ,
		\_2278__reg/NET0131 ,
		_w3832_
	);
	LUT2 #(
		.INIT('h2)
	) name2325 (
		\WX9868_reg/NET0131 ,
		\WX9932_reg/NET0131 ,
		_w3833_
	);
	LUT2 #(
		.INIT('h4)
	) name2326 (
		\WX9868_reg/NET0131 ,
		\WX9932_reg/NET0131 ,
		_w3834_
	);
	LUT2 #(
		.INIT('h1)
	) name2327 (
		_w3833_,
		_w3834_,
		_w3835_
	);
	LUT2 #(
		.INIT('h2)
	) name2328 (
		\WX9740_reg/NET0131 ,
		\WX9804_reg/NET0131 ,
		_w3836_
	);
	LUT2 #(
		.INIT('h4)
	) name2329 (
		\WX9740_reg/NET0131 ,
		\WX9804_reg/NET0131 ,
		_w3837_
	);
	LUT2 #(
		.INIT('h1)
	) name2330 (
		_w3836_,
		_w3837_,
		_w3838_
	);
	LUT2 #(
		.INIT('h4)
	) name2331 (
		_w3835_,
		_w3838_,
		_w3839_
	);
	LUT2 #(
		.INIT('h2)
	) name2332 (
		_w3835_,
		_w3838_,
		_w3840_
	);
	LUT2 #(
		.INIT('h1)
	) name2333 (
		\TM0_pad ,
		_w3839_,
		_w3841_
	);
	LUT2 #(
		.INIT('h4)
	) name2334 (
		_w3840_,
		_w3841_,
		_w3842_
	);
	LUT2 #(
		.INIT('h2)
	) name2335 (
		_w1976_,
		_w3832_,
		_w3843_
	);
	LUT2 #(
		.INIT('h4)
	) name2336 (
		_w3842_,
		_w3843_,
		_w3844_
	);
	LUT2 #(
		.INIT('h1)
	) name2337 (
		_w3831_,
		_w3844_,
		_w3845_
	);
	LUT2 #(
		.INIT('h2)
	) name2338 (
		_w3011_,
		_w3681_,
		_w3846_
	);
	LUT2 #(
		.INIT('h2)
	) name2339 (
		\TM0_pad ,
		\_2311__reg/NET0131 ,
		_w3847_
	);
	LUT2 #(
		.INIT('h2)
	) name2340 (
		\WX11159_reg/NET0131 ,
		\WX11223_reg/NET0131 ,
		_w3848_
	);
	LUT2 #(
		.INIT('h4)
	) name2341 (
		\WX11159_reg/NET0131 ,
		\WX11223_reg/NET0131 ,
		_w3849_
	);
	LUT2 #(
		.INIT('h1)
	) name2342 (
		_w3848_,
		_w3849_,
		_w3850_
	);
	LUT2 #(
		.INIT('h2)
	) name2343 (
		\WX11031_reg/NET0131 ,
		\WX11095_reg/NET0131 ,
		_w3851_
	);
	LUT2 #(
		.INIT('h4)
	) name2344 (
		\WX11031_reg/NET0131 ,
		\WX11095_reg/NET0131 ,
		_w3852_
	);
	LUT2 #(
		.INIT('h1)
	) name2345 (
		_w3851_,
		_w3852_,
		_w3853_
	);
	LUT2 #(
		.INIT('h4)
	) name2346 (
		_w3850_,
		_w3853_,
		_w3854_
	);
	LUT2 #(
		.INIT('h2)
	) name2347 (
		_w3850_,
		_w3853_,
		_w3855_
	);
	LUT2 #(
		.INIT('h1)
	) name2348 (
		\TM0_pad ,
		_w3854_,
		_w3856_
	);
	LUT2 #(
		.INIT('h4)
	) name2349 (
		_w3855_,
		_w3856_,
		_w3857_
	);
	LUT2 #(
		.INIT('h2)
	) name2350 (
		_w1976_,
		_w3847_,
		_w3858_
	);
	LUT2 #(
		.INIT('h4)
	) name2351 (
		_w3857_,
		_w3858_,
		_w3859_
	);
	LUT2 #(
		.INIT('h1)
	) name2352 (
		_w3846_,
		_w3859_,
		_w3860_
	);
	LUT2 #(
		.INIT('h8)
	) name2353 (
		\TM0_pad ,
		\_2129__reg/NET0131 ,
		_w3861_
	);
	LUT2 #(
		.INIT('h2)
	) name2354 (
		\WX3381_reg/NET0131 ,
		\WX3445_reg/NET0131 ,
		_w3862_
	);
	LUT2 #(
		.INIT('h4)
	) name2355 (
		\WX3381_reg/NET0131 ,
		\WX3445_reg/NET0131 ,
		_w3863_
	);
	LUT2 #(
		.INIT('h1)
	) name2356 (
		_w3862_,
		_w3863_,
		_w3864_
	);
	LUT2 #(
		.INIT('h2)
	) name2357 (
		\WX3317_reg/NET0131 ,
		_w3864_,
		_w3865_
	);
	LUT2 #(
		.INIT('h4)
	) name2358 (
		\WX3317_reg/NET0131 ,
		_w3864_,
		_w3866_
	);
	LUT2 #(
		.INIT('h1)
	) name2359 (
		_w3865_,
		_w3866_,
		_w3867_
	);
	LUT2 #(
		.INIT('h2)
	) name2360 (
		\TM1_pad ,
		\WX3253_reg/NET0131 ,
		_w3868_
	);
	LUT2 #(
		.INIT('h4)
	) name2361 (
		\TM1_pad ,
		\WX3253_reg/NET0131 ,
		_w3869_
	);
	LUT2 #(
		.INIT('h1)
	) name2362 (
		_w3868_,
		_w3869_,
		_w3870_
	);
	LUT2 #(
		.INIT('h4)
	) name2363 (
		_w3867_,
		_w3870_,
		_w3871_
	);
	LUT2 #(
		.INIT('h2)
	) name2364 (
		_w3867_,
		_w3870_,
		_w3872_
	);
	LUT2 #(
		.INIT('h1)
	) name2365 (
		\TM0_pad ,
		_w3871_,
		_w3873_
	);
	LUT2 #(
		.INIT('h4)
	) name2366 (
		_w3872_,
		_w3873_,
		_w3874_
	);
	LUT2 #(
		.INIT('h1)
	) name2367 (
		_w3861_,
		_w3874_,
		_w3875_
	);
	LUT2 #(
		.INIT('h2)
	) name2368 (
		_w1976_,
		_w3875_,
		_w3876_
	);
	LUT2 #(
		.INIT('h1)
	) name2369 (
		_w1682_,
		_w3619_,
		_w3877_
	);
	LUT2 #(
		.INIT('h2)
	) name2370 (
		_w1973_,
		_w3877_,
		_w3878_
	);
	LUT2 #(
		.INIT('h1)
	) name2371 (
		_w3876_,
		_w3878_,
		_w3879_
	);
	LUT2 #(
		.INIT('h2)
	) name2372 (
		_w3644_,
		_w3666_,
		_w3880_
	);
	LUT2 #(
		.INIT('h2)
	) name2373 (
		\TM0_pad ,
		\_2179__reg/NET0131 ,
		_w3881_
	);
	LUT2 #(
		.INIT('h2)
	) name2374 (
		\WX5995_reg/NET0131 ,
		\WX6059_reg/NET0131 ,
		_w3882_
	);
	LUT2 #(
		.INIT('h4)
	) name2375 (
		\WX5995_reg/NET0131 ,
		\WX6059_reg/NET0131 ,
		_w3883_
	);
	LUT2 #(
		.INIT('h1)
	) name2376 (
		_w3882_,
		_w3883_,
		_w3884_
	);
	LUT2 #(
		.INIT('h2)
	) name2377 (
		\WX5867_reg/NET0131 ,
		\WX5931_reg/NET0131 ,
		_w3885_
	);
	LUT2 #(
		.INIT('h4)
	) name2378 (
		\WX5867_reg/NET0131 ,
		\WX5931_reg/NET0131 ,
		_w3886_
	);
	LUT2 #(
		.INIT('h1)
	) name2379 (
		_w3885_,
		_w3886_,
		_w3887_
	);
	LUT2 #(
		.INIT('h4)
	) name2380 (
		_w3884_,
		_w3887_,
		_w3888_
	);
	LUT2 #(
		.INIT('h2)
	) name2381 (
		_w3884_,
		_w3887_,
		_w3889_
	);
	LUT2 #(
		.INIT('h1)
	) name2382 (
		\TM0_pad ,
		_w3888_,
		_w3890_
	);
	LUT2 #(
		.INIT('h4)
	) name2383 (
		_w3889_,
		_w3890_,
		_w3891_
	);
	LUT2 #(
		.INIT('h2)
	) name2384 (
		_w1976_,
		_w3881_,
		_w3892_
	);
	LUT2 #(
		.INIT('h4)
	) name2385 (
		_w3891_,
		_w3892_,
		_w3893_
	);
	LUT2 #(
		.INIT('h1)
	) name2386 (
		_w3880_,
		_w3893_,
		_w3894_
	);
	LUT2 #(
		.INIT('h2)
	) name2387 (
		_w3483_,
		_w3730_,
		_w3895_
	);
	LUT2 #(
		.INIT('h2)
	) name2388 (
		\TM0_pad ,
		\_2212__reg/NET0131 ,
		_w3896_
	);
	LUT2 #(
		.INIT('h2)
	) name2389 (
		\WX7286_reg/NET0131 ,
		\WX7350_reg/NET0131 ,
		_w3897_
	);
	LUT2 #(
		.INIT('h4)
	) name2390 (
		\WX7286_reg/NET0131 ,
		\WX7350_reg/NET0131 ,
		_w3898_
	);
	LUT2 #(
		.INIT('h1)
	) name2391 (
		_w3897_,
		_w3898_,
		_w3899_
	);
	LUT2 #(
		.INIT('h2)
	) name2392 (
		\WX7158_reg/NET0131 ,
		\WX7222_reg/NET0131 ,
		_w3900_
	);
	LUT2 #(
		.INIT('h4)
	) name2393 (
		\WX7158_reg/NET0131 ,
		\WX7222_reg/NET0131 ,
		_w3901_
	);
	LUT2 #(
		.INIT('h1)
	) name2394 (
		_w3900_,
		_w3901_,
		_w3902_
	);
	LUT2 #(
		.INIT('h4)
	) name2395 (
		_w3899_,
		_w3902_,
		_w3903_
	);
	LUT2 #(
		.INIT('h2)
	) name2396 (
		_w3899_,
		_w3902_,
		_w3904_
	);
	LUT2 #(
		.INIT('h1)
	) name2397 (
		\TM0_pad ,
		_w3903_,
		_w3905_
	);
	LUT2 #(
		.INIT('h4)
	) name2398 (
		_w3904_,
		_w3905_,
		_w3906_
	);
	LUT2 #(
		.INIT('h2)
	) name2399 (
		_w1976_,
		_w3896_,
		_w3907_
	);
	LUT2 #(
		.INIT('h4)
	) name2400 (
		_w3906_,
		_w3907_,
		_w3908_
	);
	LUT2 #(
		.INIT('h1)
	) name2401 (
		_w3895_,
		_w3908_,
		_w3909_
	);
	LUT2 #(
		.INIT('h2)
	) name2402 (
		_w2023_,
		_w3745_,
		_w3910_
	);
	LUT2 #(
		.INIT('h2)
	) name2403 (
		\TM0_pad ,
		\_2245__reg/NET0131 ,
		_w3911_
	);
	LUT2 #(
		.INIT('h2)
	) name2404 (
		\WX8577_reg/NET0131 ,
		\WX8641_reg/NET0131 ,
		_w3912_
	);
	LUT2 #(
		.INIT('h4)
	) name2405 (
		\WX8577_reg/NET0131 ,
		\WX8641_reg/NET0131 ,
		_w3913_
	);
	LUT2 #(
		.INIT('h1)
	) name2406 (
		_w3912_,
		_w3913_,
		_w3914_
	);
	LUT2 #(
		.INIT('h2)
	) name2407 (
		\WX8449_reg/NET0131 ,
		\WX8513_reg/NET0131 ,
		_w3915_
	);
	LUT2 #(
		.INIT('h4)
	) name2408 (
		\WX8449_reg/NET0131 ,
		\WX8513_reg/NET0131 ,
		_w3916_
	);
	LUT2 #(
		.INIT('h1)
	) name2409 (
		_w3915_,
		_w3916_,
		_w3917_
	);
	LUT2 #(
		.INIT('h4)
	) name2410 (
		_w3914_,
		_w3917_,
		_w3918_
	);
	LUT2 #(
		.INIT('h2)
	) name2411 (
		_w3914_,
		_w3917_,
		_w3919_
	);
	LUT2 #(
		.INIT('h1)
	) name2412 (
		\TM0_pad ,
		_w3918_,
		_w3920_
	);
	LUT2 #(
		.INIT('h4)
	) name2413 (
		_w3919_,
		_w3920_,
		_w3921_
	);
	LUT2 #(
		.INIT('h2)
	) name2414 (
		_w1976_,
		_w3911_,
		_w3922_
	);
	LUT2 #(
		.INIT('h4)
	) name2415 (
		_w3921_,
		_w3922_,
		_w3923_
	);
	LUT2 #(
		.INIT('h1)
	) name2416 (
		_w3910_,
		_w3923_,
		_w3924_
	);
	LUT2 #(
		.INIT('h1)
	) name2417 (
		\TM0_pad ,
		_w1646_,
		_w3925_
	);
	LUT2 #(
		.INIT('h1)
	) name2418 (
		_w1637_,
		_w3925_,
		_w3926_
	);
	LUT2 #(
		.INIT('h2)
	) name2419 (
		_w1973_,
		_w3926_,
		_w3927_
	);
	LUT2 #(
		.INIT('h8)
	) name2420 (
		\TM0_pad ,
		\_2095__reg/NET0131 ,
		_w3928_
	);
	LUT2 #(
		.INIT('h2)
	) name2421 (
		\WX2092_reg/NET0131 ,
		\WX2156_reg/NET0131 ,
		_w3929_
	);
	LUT2 #(
		.INIT('h4)
	) name2422 (
		\WX2092_reg/NET0131 ,
		\WX2156_reg/NET0131 ,
		_w3930_
	);
	LUT2 #(
		.INIT('h1)
	) name2423 (
		_w3929_,
		_w3930_,
		_w3931_
	);
	LUT2 #(
		.INIT('h2)
	) name2424 (
		\WX2028_reg/NET0131 ,
		_w3931_,
		_w3932_
	);
	LUT2 #(
		.INIT('h4)
	) name2425 (
		\WX2028_reg/NET0131 ,
		_w3931_,
		_w3933_
	);
	LUT2 #(
		.INIT('h1)
	) name2426 (
		_w3932_,
		_w3933_,
		_w3934_
	);
	LUT2 #(
		.INIT('h2)
	) name2427 (
		\TM1_pad ,
		\WX1964_reg/NET0131 ,
		_w3935_
	);
	LUT2 #(
		.INIT('h4)
	) name2428 (
		\TM1_pad ,
		\WX1964_reg/NET0131 ,
		_w3936_
	);
	LUT2 #(
		.INIT('h1)
	) name2429 (
		_w3935_,
		_w3936_,
		_w3937_
	);
	LUT2 #(
		.INIT('h4)
	) name2430 (
		_w3934_,
		_w3937_,
		_w3938_
	);
	LUT2 #(
		.INIT('h2)
	) name2431 (
		_w3934_,
		_w3937_,
		_w3939_
	);
	LUT2 #(
		.INIT('h1)
	) name2432 (
		\TM0_pad ,
		_w3938_,
		_w3940_
	);
	LUT2 #(
		.INIT('h4)
	) name2433 (
		_w3939_,
		_w3940_,
		_w3941_
	);
	LUT2 #(
		.INIT('h1)
	) name2434 (
		_w3928_,
		_w3941_,
		_w3942_
	);
	LUT2 #(
		.INIT('h2)
	) name2435 (
		_w1976_,
		_w3942_,
		_w3943_
	);
	LUT2 #(
		.INIT('h1)
	) name2436 (
		_w3927_,
		_w3943_,
		_w3944_
	);
	LUT2 #(
		.INIT('h1)
	) name2437 (
		_w1682_,
		_w2186_,
		_w3945_
	);
	LUT2 #(
		.INIT('h2)
	) name2438 (
		_w1973_,
		_w3945_,
		_w3946_
	);
	LUT2 #(
		.INIT('h1)
	) name2439 (
		\DATA_0_20_pad ,
		\TM0_pad ,
		_w3947_
	);
	LUT2 #(
		.INIT('h2)
	) name2440 (
		\TM0_pad ,
		\_2353__reg/NET0131 ,
		_w3948_
	);
	LUT2 #(
		.INIT('h2)
	) name2441 (
		_w1976_,
		_w3947_,
		_w3949_
	);
	LUT2 #(
		.INIT('h4)
	) name2442 (
		_w3948_,
		_w3949_,
		_w3950_
	);
	LUT2 #(
		.INIT('h1)
	) name2443 (
		_w3946_,
		_w3950_,
		_w3951_
	);
	LUT2 #(
		.INIT('h8)
	) name2444 (
		RESET_pad,
		\WX10849_reg/NET0131 ,
		_w3952_
	);
	LUT2 #(
		.INIT('h4)
	) name2445 (
		_w1894_,
		_w1973_,
		_w3953_
	);
	LUT2 #(
		.INIT('h2)
	) name2446 (
		\WX3413_reg/NET0131 ,
		\WX3477_reg/NET0131 ,
		_w3954_
	);
	LUT2 #(
		.INIT('h4)
	) name2447 (
		\WX3413_reg/NET0131 ,
		\WX3477_reg/NET0131 ,
		_w3955_
	);
	LUT2 #(
		.INIT('h1)
	) name2448 (
		_w3954_,
		_w3955_,
		_w3956_
	);
	LUT2 #(
		.INIT('h2)
	) name2449 (
		\WX3285_reg/NET0131 ,
		\WX3349_reg/NET0131 ,
		_w3957_
	);
	LUT2 #(
		.INIT('h4)
	) name2450 (
		\WX3285_reg/NET0131 ,
		\WX3349_reg/NET0131 ,
		_w3958_
	);
	LUT2 #(
		.INIT('h1)
	) name2451 (
		_w3957_,
		_w3958_,
		_w3959_
	);
	LUT2 #(
		.INIT('h4)
	) name2452 (
		_w3956_,
		_w3959_,
		_w3960_
	);
	LUT2 #(
		.INIT('h2)
	) name2453 (
		_w3956_,
		_w3959_,
		_w3961_
	);
	LUT2 #(
		.INIT('h1)
	) name2454 (
		\TM0_pad ,
		_w3960_,
		_w3962_
	);
	LUT2 #(
		.INIT('h4)
	) name2455 (
		_w3961_,
		_w3962_,
		_w3963_
	);
	LUT2 #(
		.INIT('h2)
	) name2456 (
		_w3953_,
		_w3963_,
		_w3964_
	);
	LUT2 #(
		.INIT('h2)
	) name2457 (
		\TM0_pad ,
		\_2145__reg/NET0131 ,
		_w3965_
	);
	LUT2 #(
		.INIT('h2)
	) name2458 (
		\WX4706_reg/NET0131 ,
		\WX4770_reg/NET0131 ,
		_w3966_
	);
	LUT2 #(
		.INIT('h4)
	) name2459 (
		\WX4706_reg/NET0131 ,
		\WX4770_reg/NET0131 ,
		_w3967_
	);
	LUT2 #(
		.INIT('h1)
	) name2460 (
		_w3966_,
		_w3967_,
		_w3968_
	);
	LUT2 #(
		.INIT('h2)
	) name2461 (
		\WX4578_reg/NET0131 ,
		\WX4642_reg/NET0131 ,
		_w3969_
	);
	LUT2 #(
		.INIT('h4)
	) name2462 (
		\WX4578_reg/NET0131 ,
		\WX4642_reg/NET0131 ,
		_w3970_
	);
	LUT2 #(
		.INIT('h1)
	) name2463 (
		_w3969_,
		_w3970_,
		_w3971_
	);
	LUT2 #(
		.INIT('h4)
	) name2464 (
		_w3968_,
		_w3971_,
		_w3972_
	);
	LUT2 #(
		.INIT('h2)
	) name2465 (
		_w3968_,
		_w3971_,
		_w3973_
	);
	LUT2 #(
		.INIT('h1)
	) name2466 (
		\TM0_pad ,
		_w3972_,
		_w3974_
	);
	LUT2 #(
		.INIT('h4)
	) name2467 (
		_w3973_,
		_w3974_,
		_w3975_
	);
	LUT2 #(
		.INIT('h2)
	) name2468 (
		_w1976_,
		_w3965_,
		_w3976_
	);
	LUT2 #(
		.INIT('h4)
	) name2469 (
		_w3975_,
		_w3976_,
		_w3977_
	);
	LUT2 #(
		.INIT('h1)
	) name2470 (
		_w3964_,
		_w3977_,
		_w3978_
	);
	LUT2 #(
		.INIT('h2)
	) name2471 (
		_w2023_,
		_w3921_,
		_w3979_
	);
	LUT2 #(
		.INIT('h2)
	) name2472 (
		\TM0_pad ,
		\_2277__reg/NET0131 ,
		_w3980_
	);
	LUT2 #(
		.INIT('h2)
	) name2473 (
		\WX9870_reg/NET0131 ,
		\WX9934_reg/NET0131 ,
		_w3981_
	);
	LUT2 #(
		.INIT('h4)
	) name2474 (
		\WX9870_reg/NET0131 ,
		\WX9934_reg/NET0131 ,
		_w3982_
	);
	LUT2 #(
		.INIT('h1)
	) name2475 (
		_w3981_,
		_w3982_,
		_w3983_
	);
	LUT2 #(
		.INIT('h2)
	) name2476 (
		\WX9742_reg/NET0131 ,
		\WX9806_reg/NET0131 ,
		_w3984_
	);
	LUT2 #(
		.INIT('h4)
	) name2477 (
		\WX9742_reg/NET0131 ,
		\WX9806_reg/NET0131 ,
		_w3985_
	);
	LUT2 #(
		.INIT('h1)
	) name2478 (
		_w3984_,
		_w3985_,
		_w3986_
	);
	LUT2 #(
		.INIT('h4)
	) name2479 (
		_w3983_,
		_w3986_,
		_w3987_
	);
	LUT2 #(
		.INIT('h2)
	) name2480 (
		_w3983_,
		_w3986_,
		_w3988_
	);
	LUT2 #(
		.INIT('h1)
	) name2481 (
		\TM0_pad ,
		_w3987_,
		_w3989_
	);
	LUT2 #(
		.INIT('h4)
	) name2482 (
		_w3988_,
		_w3989_,
		_w3990_
	);
	LUT2 #(
		.INIT('h2)
	) name2483 (
		_w1976_,
		_w3980_,
		_w3991_
	);
	LUT2 #(
		.INIT('h4)
	) name2484 (
		_w3990_,
		_w3991_,
		_w3992_
	);
	LUT2 #(
		.INIT('h1)
	) name2485 (
		_w3979_,
		_w3992_,
		_w3993_
	);
	LUT2 #(
		.INIT('h2)
	) name2486 (
		_w3172_,
		_w3842_,
		_w3994_
	);
	LUT2 #(
		.INIT('h2)
	) name2487 (
		\TM0_pad ,
		\_2310__reg/NET0131 ,
		_w3995_
	);
	LUT2 #(
		.INIT('h2)
	) name2488 (
		\WX11161_reg/NET0131 ,
		\WX11225_reg/NET0131 ,
		_w3996_
	);
	LUT2 #(
		.INIT('h4)
	) name2489 (
		\WX11161_reg/NET0131 ,
		\WX11225_reg/NET0131 ,
		_w3997_
	);
	LUT2 #(
		.INIT('h1)
	) name2490 (
		_w3996_,
		_w3997_,
		_w3998_
	);
	LUT2 #(
		.INIT('h2)
	) name2491 (
		\WX11033_reg/NET0131 ,
		\WX11097_reg/NET0131 ,
		_w3999_
	);
	LUT2 #(
		.INIT('h4)
	) name2492 (
		\WX11033_reg/NET0131 ,
		\WX11097_reg/NET0131 ,
		_w4000_
	);
	LUT2 #(
		.INIT('h1)
	) name2493 (
		_w3999_,
		_w4000_,
		_w4001_
	);
	LUT2 #(
		.INIT('h4)
	) name2494 (
		_w3998_,
		_w4001_,
		_w4002_
	);
	LUT2 #(
		.INIT('h2)
	) name2495 (
		_w3998_,
		_w4001_,
		_w4003_
	);
	LUT2 #(
		.INIT('h1)
	) name2496 (
		\TM0_pad ,
		_w4002_,
		_w4004_
	);
	LUT2 #(
		.INIT('h4)
	) name2497 (
		_w4003_,
		_w4004_,
		_w4005_
	);
	LUT2 #(
		.INIT('h2)
	) name2498 (
		_w1976_,
		_w3995_,
		_w4006_
	);
	LUT2 #(
		.INIT('h4)
	) name2499 (
		_w4005_,
		_w4006_,
		_w4007_
	);
	LUT2 #(
		.INIT('h1)
	) name2500 (
		_w3994_,
		_w4007_,
		_w4008_
	);
	LUT2 #(
		.INIT('h8)
	) name2501 (
		\TM0_pad ,
		\_2128__reg/NET0131 ,
		_w4009_
	);
	LUT2 #(
		.INIT('h2)
	) name2502 (
		\WX3383_reg/NET0131 ,
		\WX3447_reg/NET0131 ,
		_w4010_
	);
	LUT2 #(
		.INIT('h4)
	) name2503 (
		\WX3383_reg/NET0131 ,
		\WX3447_reg/NET0131 ,
		_w4011_
	);
	LUT2 #(
		.INIT('h1)
	) name2504 (
		_w4010_,
		_w4011_,
		_w4012_
	);
	LUT2 #(
		.INIT('h2)
	) name2505 (
		\WX3319_reg/NET0131 ,
		_w4012_,
		_w4013_
	);
	LUT2 #(
		.INIT('h4)
	) name2506 (
		\WX3319_reg/NET0131 ,
		_w4012_,
		_w4014_
	);
	LUT2 #(
		.INIT('h1)
	) name2507 (
		_w4013_,
		_w4014_,
		_w4015_
	);
	LUT2 #(
		.INIT('h2)
	) name2508 (
		\TM1_pad ,
		\WX3255_reg/NET0131 ,
		_w4016_
	);
	LUT2 #(
		.INIT('h4)
	) name2509 (
		\TM1_pad ,
		\WX3255_reg/NET0131 ,
		_w4017_
	);
	LUT2 #(
		.INIT('h1)
	) name2510 (
		_w4016_,
		_w4017_,
		_w4018_
	);
	LUT2 #(
		.INIT('h4)
	) name2511 (
		_w4015_,
		_w4018_,
		_w4019_
	);
	LUT2 #(
		.INIT('h2)
	) name2512 (
		_w4015_,
		_w4018_,
		_w4020_
	);
	LUT2 #(
		.INIT('h1)
	) name2513 (
		\TM0_pad ,
		_w4019_,
		_w4021_
	);
	LUT2 #(
		.INIT('h4)
	) name2514 (
		_w4020_,
		_w4021_,
		_w4022_
	);
	LUT2 #(
		.INIT('h1)
	) name2515 (
		_w4009_,
		_w4022_,
		_w4023_
	);
	LUT2 #(
		.INIT('h2)
	) name2516 (
		_w1976_,
		_w4023_,
		_w4024_
	);
	LUT2 #(
		.INIT('h1)
	) name2517 (
		_w1653_,
		_w3780_,
		_w4025_
	);
	LUT2 #(
		.INIT('h2)
	) name2518 (
		_w1973_,
		_w4025_,
		_w4026_
	);
	LUT2 #(
		.INIT('h1)
	) name2519 (
		_w4024_,
		_w4026_,
		_w4027_
	);
	LUT2 #(
		.INIT('h2)
	) name2520 (
		_w3805_,
		_w3827_,
		_w4028_
	);
	LUT2 #(
		.INIT('h2)
	) name2521 (
		\TM0_pad ,
		\_2178__reg/NET0131 ,
		_w4029_
	);
	LUT2 #(
		.INIT('h2)
	) name2522 (
		\WX5997_reg/NET0131 ,
		\WX6061_reg/NET0131 ,
		_w4030_
	);
	LUT2 #(
		.INIT('h4)
	) name2523 (
		\WX5997_reg/NET0131 ,
		\WX6061_reg/NET0131 ,
		_w4031_
	);
	LUT2 #(
		.INIT('h1)
	) name2524 (
		_w4030_,
		_w4031_,
		_w4032_
	);
	LUT2 #(
		.INIT('h2)
	) name2525 (
		\WX5869_reg/NET0131 ,
		\WX5933_reg/NET0131 ,
		_w4033_
	);
	LUT2 #(
		.INIT('h4)
	) name2526 (
		\WX5869_reg/NET0131 ,
		\WX5933_reg/NET0131 ,
		_w4034_
	);
	LUT2 #(
		.INIT('h1)
	) name2527 (
		_w4033_,
		_w4034_,
		_w4035_
	);
	LUT2 #(
		.INIT('h4)
	) name2528 (
		_w4032_,
		_w4035_,
		_w4036_
	);
	LUT2 #(
		.INIT('h2)
	) name2529 (
		_w4032_,
		_w4035_,
		_w4037_
	);
	LUT2 #(
		.INIT('h1)
	) name2530 (
		\TM0_pad ,
		_w4036_,
		_w4038_
	);
	LUT2 #(
		.INIT('h4)
	) name2531 (
		_w4037_,
		_w4038_,
		_w4039_
	);
	LUT2 #(
		.INIT('h2)
	) name2532 (
		_w1976_,
		_w4029_,
		_w4040_
	);
	LUT2 #(
		.INIT('h4)
	) name2533 (
		_w4039_,
		_w4040_,
		_w4041_
	);
	LUT2 #(
		.INIT('h1)
	) name2534 (
		_w4028_,
		_w4041_,
		_w4042_
	);
	LUT2 #(
		.INIT('h2)
	) name2535 (
		_w3644_,
		_w3891_,
		_w4043_
	);
	LUT2 #(
		.INIT('h2)
	) name2536 (
		\TM0_pad ,
		\_2211__reg/NET0131 ,
		_w4044_
	);
	LUT2 #(
		.INIT('h2)
	) name2537 (
		\WX7288_reg/NET0131 ,
		\WX7352_reg/NET0131 ,
		_w4045_
	);
	LUT2 #(
		.INIT('h4)
	) name2538 (
		\WX7288_reg/NET0131 ,
		\WX7352_reg/NET0131 ,
		_w4046_
	);
	LUT2 #(
		.INIT('h1)
	) name2539 (
		_w4045_,
		_w4046_,
		_w4047_
	);
	LUT2 #(
		.INIT('h2)
	) name2540 (
		\WX7160_reg/NET0131 ,
		\WX7224_reg/NET0131 ,
		_w4048_
	);
	LUT2 #(
		.INIT('h4)
	) name2541 (
		\WX7160_reg/NET0131 ,
		\WX7224_reg/NET0131 ,
		_w4049_
	);
	LUT2 #(
		.INIT('h1)
	) name2542 (
		_w4048_,
		_w4049_,
		_w4050_
	);
	LUT2 #(
		.INIT('h4)
	) name2543 (
		_w4047_,
		_w4050_,
		_w4051_
	);
	LUT2 #(
		.INIT('h2)
	) name2544 (
		_w4047_,
		_w4050_,
		_w4052_
	);
	LUT2 #(
		.INIT('h1)
	) name2545 (
		\TM0_pad ,
		_w4051_,
		_w4053_
	);
	LUT2 #(
		.INIT('h4)
	) name2546 (
		_w4052_,
		_w4053_,
		_w4054_
	);
	LUT2 #(
		.INIT('h2)
	) name2547 (
		_w1976_,
		_w4044_,
		_w4055_
	);
	LUT2 #(
		.INIT('h4)
	) name2548 (
		_w4054_,
		_w4055_,
		_w4056_
	);
	LUT2 #(
		.INIT('h1)
	) name2549 (
		_w4043_,
		_w4056_,
		_w4057_
	);
	LUT2 #(
		.INIT('h2)
	) name2550 (
		_w3483_,
		_w3906_,
		_w4058_
	);
	LUT2 #(
		.INIT('h2)
	) name2551 (
		\TM0_pad ,
		\_2244__reg/NET0131 ,
		_w4059_
	);
	LUT2 #(
		.INIT('h2)
	) name2552 (
		\WX8579_reg/NET0131 ,
		\WX8643_reg/NET0131 ,
		_w4060_
	);
	LUT2 #(
		.INIT('h4)
	) name2553 (
		\WX8579_reg/NET0131 ,
		\WX8643_reg/NET0131 ,
		_w4061_
	);
	LUT2 #(
		.INIT('h1)
	) name2554 (
		_w4060_,
		_w4061_,
		_w4062_
	);
	LUT2 #(
		.INIT('h2)
	) name2555 (
		\WX8451_reg/NET0131 ,
		\WX8515_reg/NET0131 ,
		_w4063_
	);
	LUT2 #(
		.INIT('h4)
	) name2556 (
		\WX8451_reg/NET0131 ,
		\WX8515_reg/NET0131 ,
		_w4064_
	);
	LUT2 #(
		.INIT('h1)
	) name2557 (
		_w4063_,
		_w4064_,
		_w4065_
	);
	LUT2 #(
		.INIT('h4)
	) name2558 (
		_w4062_,
		_w4065_,
		_w4066_
	);
	LUT2 #(
		.INIT('h2)
	) name2559 (
		_w4062_,
		_w4065_,
		_w4067_
	);
	LUT2 #(
		.INIT('h1)
	) name2560 (
		\TM0_pad ,
		_w4066_,
		_w4068_
	);
	LUT2 #(
		.INIT('h4)
	) name2561 (
		_w4067_,
		_w4068_,
		_w4069_
	);
	LUT2 #(
		.INIT('h2)
	) name2562 (
		_w1976_,
		_w4059_,
		_w4070_
	);
	LUT2 #(
		.INIT('h4)
	) name2563 (
		_w4069_,
		_w4070_,
		_w4071_
	);
	LUT2 #(
		.INIT('h1)
	) name2564 (
		_w4058_,
		_w4071_,
		_w4072_
	);
	LUT2 #(
		.INIT('h8)
	) name2565 (
		\TM0_pad ,
		\_2094__reg/NET0131 ,
		_w4073_
	);
	LUT2 #(
		.INIT('h2)
	) name2566 (
		\WX2094_reg/NET0131 ,
		\WX2158_reg/NET0131 ,
		_w4074_
	);
	LUT2 #(
		.INIT('h4)
	) name2567 (
		\WX2094_reg/NET0131 ,
		\WX2158_reg/NET0131 ,
		_w4075_
	);
	LUT2 #(
		.INIT('h1)
	) name2568 (
		_w4074_,
		_w4075_,
		_w4076_
	);
	LUT2 #(
		.INIT('h2)
	) name2569 (
		\WX2030_reg/NET0131 ,
		_w4076_,
		_w4077_
	);
	LUT2 #(
		.INIT('h4)
	) name2570 (
		\WX2030_reg/NET0131 ,
		_w4076_,
		_w4078_
	);
	LUT2 #(
		.INIT('h1)
	) name2571 (
		_w4077_,
		_w4078_,
		_w4079_
	);
	LUT2 #(
		.INIT('h2)
	) name2572 (
		\TM1_pad ,
		\WX1966_reg/NET0131 ,
		_w4080_
	);
	LUT2 #(
		.INIT('h4)
	) name2573 (
		\TM1_pad ,
		\WX1966_reg/NET0131 ,
		_w4081_
	);
	LUT2 #(
		.INIT('h1)
	) name2574 (
		_w4080_,
		_w4081_,
		_w4082_
	);
	LUT2 #(
		.INIT('h4)
	) name2575 (
		_w4079_,
		_w4082_,
		_w4083_
	);
	LUT2 #(
		.INIT('h2)
	) name2576 (
		_w4079_,
		_w4082_,
		_w4084_
	);
	LUT2 #(
		.INIT('h1)
	) name2577 (
		\TM0_pad ,
		_w4083_,
		_w4085_
	);
	LUT2 #(
		.INIT('h4)
	) name2578 (
		_w4084_,
		_w4085_,
		_w4086_
	);
	LUT2 #(
		.INIT('h1)
	) name2579 (
		_w4073_,
		_w4086_,
		_w4087_
	);
	LUT2 #(
		.INIT('h2)
	) name2580 (
		_w1976_,
		_w4087_,
		_w4088_
	);
	LUT2 #(
		.INIT('h1)
	) name2581 (
		\TM0_pad ,
		_w1630_,
		_w4089_
	);
	LUT2 #(
		.INIT('h1)
	) name2582 (
		_w1621_,
		_w4089_,
		_w4090_
	);
	LUT2 #(
		.INIT('h2)
	) name2583 (
		_w1973_,
		_w4090_,
		_w4091_
	);
	LUT2 #(
		.INIT('h1)
	) name2584 (
		_w4088_,
		_w4091_,
		_w4092_
	);
	LUT2 #(
		.INIT('h1)
	) name2585 (
		_w1653_,
		_w2418_,
		_w4093_
	);
	LUT2 #(
		.INIT('h2)
	) name2586 (
		_w1973_,
		_w4093_,
		_w4094_
	);
	LUT2 #(
		.INIT('h1)
	) name2587 (
		\DATA_0_19_pad ,
		\TM0_pad ,
		_w4095_
	);
	LUT2 #(
		.INIT('h2)
	) name2588 (
		\TM0_pad ,
		\_2352__reg/NET0131 ,
		_w4096_
	);
	LUT2 #(
		.INIT('h2)
	) name2589 (
		_w1976_,
		_w4095_,
		_w4097_
	);
	LUT2 #(
		.INIT('h4)
	) name2590 (
		_w4096_,
		_w4097_,
		_w4098_
	);
	LUT2 #(
		.INIT('h1)
	) name2591 (
		_w4094_,
		_w4098_,
		_w4099_
	);
	LUT2 #(
		.INIT('h8)
	) name2592 (
		RESET_pad,
		\WX10851_reg/NET0131 ,
		_w4100_
	);
	LUT2 #(
		.INIT('h4)
	) name2593 (
		_w1881_,
		_w1973_,
		_w4101_
	);
	LUT2 #(
		.INIT('h2)
	) name2594 (
		\WX3415_reg/NET0131 ,
		\WX3479_reg/NET0131 ,
		_w4102_
	);
	LUT2 #(
		.INIT('h4)
	) name2595 (
		\WX3415_reg/NET0131 ,
		\WX3479_reg/NET0131 ,
		_w4103_
	);
	LUT2 #(
		.INIT('h1)
	) name2596 (
		_w4102_,
		_w4103_,
		_w4104_
	);
	LUT2 #(
		.INIT('h2)
	) name2597 (
		\WX3287_reg/NET0131 ,
		\WX3351_reg/NET0131 ,
		_w4105_
	);
	LUT2 #(
		.INIT('h4)
	) name2598 (
		\WX3287_reg/NET0131 ,
		\WX3351_reg/NET0131 ,
		_w4106_
	);
	LUT2 #(
		.INIT('h1)
	) name2599 (
		_w4105_,
		_w4106_,
		_w4107_
	);
	LUT2 #(
		.INIT('h4)
	) name2600 (
		_w4104_,
		_w4107_,
		_w4108_
	);
	LUT2 #(
		.INIT('h2)
	) name2601 (
		_w4104_,
		_w4107_,
		_w4109_
	);
	LUT2 #(
		.INIT('h1)
	) name2602 (
		\TM0_pad ,
		_w4108_,
		_w4110_
	);
	LUT2 #(
		.INIT('h4)
	) name2603 (
		_w4109_,
		_w4110_,
		_w4111_
	);
	LUT2 #(
		.INIT('h2)
	) name2604 (
		_w4101_,
		_w4111_,
		_w4112_
	);
	LUT2 #(
		.INIT('h2)
	) name2605 (
		\TM0_pad ,
		\_2144__reg/NET0131 ,
		_w4113_
	);
	LUT2 #(
		.INIT('h2)
	) name2606 (
		\WX4708_reg/NET0131 ,
		\WX4772_reg/NET0131 ,
		_w4114_
	);
	LUT2 #(
		.INIT('h4)
	) name2607 (
		\WX4708_reg/NET0131 ,
		\WX4772_reg/NET0131 ,
		_w4115_
	);
	LUT2 #(
		.INIT('h1)
	) name2608 (
		_w4114_,
		_w4115_,
		_w4116_
	);
	LUT2 #(
		.INIT('h2)
	) name2609 (
		\WX4580_reg/NET0131 ,
		\WX4644_reg/NET0131 ,
		_w4117_
	);
	LUT2 #(
		.INIT('h4)
	) name2610 (
		\WX4580_reg/NET0131 ,
		\WX4644_reg/NET0131 ,
		_w4118_
	);
	LUT2 #(
		.INIT('h1)
	) name2611 (
		_w4117_,
		_w4118_,
		_w4119_
	);
	LUT2 #(
		.INIT('h4)
	) name2612 (
		_w4116_,
		_w4119_,
		_w4120_
	);
	LUT2 #(
		.INIT('h2)
	) name2613 (
		_w4116_,
		_w4119_,
		_w4121_
	);
	LUT2 #(
		.INIT('h1)
	) name2614 (
		\TM0_pad ,
		_w4120_,
		_w4122_
	);
	LUT2 #(
		.INIT('h4)
	) name2615 (
		_w4121_,
		_w4122_,
		_w4123_
	);
	LUT2 #(
		.INIT('h2)
	) name2616 (
		_w1976_,
		_w4113_,
		_w4124_
	);
	LUT2 #(
		.INIT('h4)
	) name2617 (
		_w4123_,
		_w4124_,
		_w4125_
	);
	LUT2 #(
		.INIT('h1)
	) name2618 (
		_w4112_,
		_w4125_,
		_w4126_
	);
	LUT2 #(
		.INIT('h2)
	) name2619 (
		_w3483_,
		_w4069_,
		_w4127_
	);
	LUT2 #(
		.INIT('h2)
	) name2620 (
		\TM0_pad ,
		\_2276__reg/NET0131 ,
		_w4128_
	);
	LUT2 #(
		.INIT('h2)
	) name2621 (
		\WX9872_reg/NET0131 ,
		\WX9936_reg/NET0131 ,
		_w4129_
	);
	LUT2 #(
		.INIT('h4)
	) name2622 (
		\WX9872_reg/NET0131 ,
		\WX9936_reg/NET0131 ,
		_w4130_
	);
	LUT2 #(
		.INIT('h1)
	) name2623 (
		_w4129_,
		_w4130_,
		_w4131_
	);
	LUT2 #(
		.INIT('h2)
	) name2624 (
		\WX9744_reg/NET0131 ,
		\WX9808_reg/NET0131 ,
		_w4132_
	);
	LUT2 #(
		.INIT('h4)
	) name2625 (
		\WX9744_reg/NET0131 ,
		\WX9808_reg/NET0131 ,
		_w4133_
	);
	LUT2 #(
		.INIT('h1)
	) name2626 (
		_w4132_,
		_w4133_,
		_w4134_
	);
	LUT2 #(
		.INIT('h4)
	) name2627 (
		_w4131_,
		_w4134_,
		_w4135_
	);
	LUT2 #(
		.INIT('h2)
	) name2628 (
		_w4131_,
		_w4134_,
		_w4136_
	);
	LUT2 #(
		.INIT('h1)
	) name2629 (
		\TM0_pad ,
		_w4135_,
		_w4137_
	);
	LUT2 #(
		.INIT('h4)
	) name2630 (
		_w4136_,
		_w4137_,
		_w4138_
	);
	LUT2 #(
		.INIT('h2)
	) name2631 (
		_w1976_,
		_w4128_,
		_w4139_
	);
	LUT2 #(
		.INIT('h4)
	) name2632 (
		_w4138_,
		_w4139_,
		_w4140_
	);
	LUT2 #(
		.INIT('h1)
	) name2633 (
		_w4127_,
		_w4140_,
		_w4141_
	);
	LUT2 #(
		.INIT('h2)
	) name2634 (
		_w2023_,
		_w3990_,
		_w4142_
	);
	LUT2 #(
		.INIT('h2)
	) name2635 (
		\TM0_pad ,
		\_2309__reg/NET0131 ,
		_w4143_
	);
	LUT2 #(
		.INIT('h2)
	) name2636 (
		_w1976_,
		_w4143_,
		_w4144_
	);
	LUT2 #(
		.INIT('h4)
	) name2637 (
		_w2033_,
		_w4144_,
		_w4145_
	);
	LUT2 #(
		.INIT('h1)
	) name2638 (
		_w4142_,
		_w4145_,
		_w4146_
	);
	LUT2 #(
		.INIT('h8)
	) name2639 (
		\TM0_pad ,
		\_2127__reg/NET0131 ,
		_w4147_
	);
	LUT2 #(
		.INIT('h2)
	) name2640 (
		\WX3385_reg/NET0131 ,
		\WX3449_reg/NET0131 ,
		_w4148_
	);
	LUT2 #(
		.INIT('h4)
	) name2641 (
		\WX3385_reg/NET0131 ,
		\WX3449_reg/NET0131 ,
		_w4149_
	);
	LUT2 #(
		.INIT('h1)
	) name2642 (
		_w4148_,
		_w4149_,
		_w4150_
	);
	LUT2 #(
		.INIT('h2)
	) name2643 (
		\WX3321_reg/NET0131 ,
		_w4150_,
		_w4151_
	);
	LUT2 #(
		.INIT('h4)
	) name2644 (
		\WX3321_reg/NET0131 ,
		_w4150_,
		_w4152_
	);
	LUT2 #(
		.INIT('h1)
	) name2645 (
		_w4151_,
		_w4152_,
		_w4153_
	);
	LUT2 #(
		.INIT('h2)
	) name2646 (
		\TM1_pad ,
		\WX3257_reg/NET0131 ,
		_w4154_
	);
	LUT2 #(
		.INIT('h4)
	) name2647 (
		\TM1_pad ,
		\WX3257_reg/NET0131 ,
		_w4155_
	);
	LUT2 #(
		.INIT('h1)
	) name2648 (
		_w4154_,
		_w4155_,
		_w4156_
	);
	LUT2 #(
		.INIT('h4)
	) name2649 (
		_w4153_,
		_w4156_,
		_w4157_
	);
	LUT2 #(
		.INIT('h2)
	) name2650 (
		_w4153_,
		_w4156_,
		_w4158_
	);
	LUT2 #(
		.INIT('h1)
	) name2651 (
		\TM0_pad ,
		_w4157_,
		_w4159_
	);
	LUT2 #(
		.INIT('h4)
	) name2652 (
		_w4158_,
		_w4159_,
		_w4160_
	);
	LUT2 #(
		.INIT('h1)
	) name2653 (
		_w4147_,
		_w4160_,
		_w4161_
	);
	LUT2 #(
		.INIT('h2)
	) name2654 (
		_w1976_,
		_w4161_,
		_w4162_
	);
	LUT2 #(
		.INIT('h1)
	) name2655 (
		_w1637_,
		_w3941_,
		_w4163_
	);
	LUT2 #(
		.INIT('h2)
	) name2656 (
		_w1973_,
		_w4163_,
		_w4164_
	);
	LUT2 #(
		.INIT('h1)
	) name2657 (
		_w4162_,
		_w4164_,
		_w4165_
	);
	LUT2 #(
		.INIT('h2)
	) name2658 (
		_w3953_,
		_w3975_,
		_w4166_
	);
	LUT2 #(
		.INIT('h2)
	) name2659 (
		\TM0_pad ,
		\_2177__reg/NET0131 ,
		_w4167_
	);
	LUT2 #(
		.INIT('h2)
	) name2660 (
		\WX5999_reg/NET0131 ,
		\WX6063_reg/NET0131 ,
		_w4168_
	);
	LUT2 #(
		.INIT('h4)
	) name2661 (
		\WX5999_reg/NET0131 ,
		\WX6063_reg/NET0131 ,
		_w4169_
	);
	LUT2 #(
		.INIT('h1)
	) name2662 (
		_w4168_,
		_w4169_,
		_w4170_
	);
	LUT2 #(
		.INIT('h2)
	) name2663 (
		\WX5871_reg/NET0131 ,
		\WX5935_reg/NET0131 ,
		_w4171_
	);
	LUT2 #(
		.INIT('h4)
	) name2664 (
		\WX5871_reg/NET0131 ,
		\WX5935_reg/NET0131 ,
		_w4172_
	);
	LUT2 #(
		.INIT('h1)
	) name2665 (
		_w4171_,
		_w4172_,
		_w4173_
	);
	LUT2 #(
		.INIT('h4)
	) name2666 (
		_w4170_,
		_w4173_,
		_w4174_
	);
	LUT2 #(
		.INIT('h2)
	) name2667 (
		_w4170_,
		_w4173_,
		_w4175_
	);
	LUT2 #(
		.INIT('h1)
	) name2668 (
		\TM0_pad ,
		_w4174_,
		_w4176_
	);
	LUT2 #(
		.INIT('h4)
	) name2669 (
		_w4175_,
		_w4176_,
		_w4177_
	);
	LUT2 #(
		.INIT('h2)
	) name2670 (
		_w1976_,
		_w4167_,
		_w4178_
	);
	LUT2 #(
		.INIT('h4)
	) name2671 (
		_w4177_,
		_w4178_,
		_w4179_
	);
	LUT2 #(
		.INIT('h1)
	) name2672 (
		_w4166_,
		_w4179_,
		_w4180_
	);
	LUT2 #(
		.INIT('h2)
	) name2673 (
		_w3805_,
		_w4039_,
		_w4181_
	);
	LUT2 #(
		.INIT('h2)
	) name2674 (
		\TM0_pad ,
		\_2210__reg/NET0131 ,
		_w4182_
	);
	LUT2 #(
		.INIT('h2)
	) name2675 (
		\WX7290_reg/NET0131 ,
		\WX7354_reg/NET0131 ,
		_w4183_
	);
	LUT2 #(
		.INIT('h4)
	) name2676 (
		\WX7290_reg/NET0131 ,
		\WX7354_reg/NET0131 ,
		_w4184_
	);
	LUT2 #(
		.INIT('h1)
	) name2677 (
		_w4183_,
		_w4184_,
		_w4185_
	);
	LUT2 #(
		.INIT('h2)
	) name2678 (
		\WX7162_reg/NET0131 ,
		\WX7226_reg/NET0131 ,
		_w4186_
	);
	LUT2 #(
		.INIT('h4)
	) name2679 (
		\WX7162_reg/NET0131 ,
		\WX7226_reg/NET0131 ,
		_w4187_
	);
	LUT2 #(
		.INIT('h1)
	) name2680 (
		_w4186_,
		_w4187_,
		_w4188_
	);
	LUT2 #(
		.INIT('h4)
	) name2681 (
		_w4185_,
		_w4188_,
		_w4189_
	);
	LUT2 #(
		.INIT('h2)
	) name2682 (
		_w4185_,
		_w4188_,
		_w4190_
	);
	LUT2 #(
		.INIT('h1)
	) name2683 (
		\TM0_pad ,
		_w4189_,
		_w4191_
	);
	LUT2 #(
		.INIT('h4)
	) name2684 (
		_w4190_,
		_w4191_,
		_w4192_
	);
	LUT2 #(
		.INIT('h2)
	) name2685 (
		_w1976_,
		_w4182_,
		_w4193_
	);
	LUT2 #(
		.INIT('h4)
	) name2686 (
		_w4192_,
		_w4193_,
		_w4194_
	);
	LUT2 #(
		.INIT('h1)
	) name2687 (
		_w4181_,
		_w4194_,
		_w4195_
	);
	LUT2 #(
		.INIT('h2)
	) name2688 (
		_w3644_,
		_w4054_,
		_w4196_
	);
	LUT2 #(
		.INIT('h2)
	) name2689 (
		\TM0_pad ,
		\_2243__reg/NET0131 ,
		_w4197_
	);
	LUT2 #(
		.INIT('h2)
	) name2690 (
		\WX8581_reg/NET0131 ,
		\WX8645_reg/NET0131 ,
		_w4198_
	);
	LUT2 #(
		.INIT('h4)
	) name2691 (
		\WX8581_reg/NET0131 ,
		\WX8645_reg/NET0131 ,
		_w4199_
	);
	LUT2 #(
		.INIT('h1)
	) name2692 (
		_w4198_,
		_w4199_,
		_w4200_
	);
	LUT2 #(
		.INIT('h2)
	) name2693 (
		\WX8453_reg/NET0131 ,
		\WX8517_reg/NET0131 ,
		_w4201_
	);
	LUT2 #(
		.INIT('h4)
	) name2694 (
		\WX8453_reg/NET0131 ,
		\WX8517_reg/NET0131 ,
		_w4202_
	);
	LUT2 #(
		.INIT('h1)
	) name2695 (
		_w4201_,
		_w4202_,
		_w4203_
	);
	LUT2 #(
		.INIT('h4)
	) name2696 (
		_w4200_,
		_w4203_,
		_w4204_
	);
	LUT2 #(
		.INIT('h2)
	) name2697 (
		_w4200_,
		_w4203_,
		_w4205_
	);
	LUT2 #(
		.INIT('h1)
	) name2698 (
		\TM0_pad ,
		_w4204_,
		_w4206_
	);
	LUT2 #(
		.INIT('h4)
	) name2699 (
		_w4205_,
		_w4206_,
		_w4207_
	);
	LUT2 #(
		.INIT('h2)
	) name2700 (
		_w1976_,
		_w4197_,
		_w4208_
	);
	LUT2 #(
		.INIT('h4)
	) name2701 (
		_w4207_,
		_w4208_,
		_w4209_
	);
	LUT2 #(
		.INIT('h1)
	) name2702 (
		_w4196_,
		_w4209_,
		_w4210_
	);
	LUT2 #(
		.INIT('h1)
	) name2703 (
		\TM0_pad ,
		_w1614_,
		_w4211_
	);
	LUT2 #(
		.INIT('h1)
	) name2704 (
		_w1605_,
		_w4211_,
		_w4212_
	);
	LUT2 #(
		.INIT('h2)
	) name2705 (
		_w1973_,
		_w4212_,
		_w4213_
	);
	LUT2 #(
		.INIT('h8)
	) name2706 (
		\TM0_pad ,
		\_2093__reg/NET0131 ,
		_w4214_
	);
	LUT2 #(
		.INIT('h2)
	) name2707 (
		\WX2096_reg/NET0131 ,
		\WX2160_reg/NET0131 ,
		_w4215_
	);
	LUT2 #(
		.INIT('h4)
	) name2708 (
		\WX2096_reg/NET0131 ,
		\WX2160_reg/NET0131 ,
		_w4216_
	);
	LUT2 #(
		.INIT('h1)
	) name2709 (
		_w4215_,
		_w4216_,
		_w4217_
	);
	LUT2 #(
		.INIT('h2)
	) name2710 (
		\WX2032_reg/NET0131 ,
		_w4217_,
		_w4218_
	);
	LUT2 #(
		.INIT('h4)
	) name2711 (
		\WX2032_reg/NET0131 ,
		_w4217_,
		_w4219_
	);
	LUT2 #(
		.INIT('h1)
	) name2712 (
		_w4218_,
		_w4219_,
		_w4220_
	);
	LUT2 #(
		.INIT('h2)
	) name2713 (
		\TM1_pad ,
		\WX1968_reg/NET0131 ,
		_w4221_
	);
	LUT2 #(
		.INIT('h4)
	) name2714 (
		\TM1_pad ,
		\WX1968_reg/NET0131 ,
		_w4222_
	);
	LUT2 #(
		.INIT('h1)
	) name2715 (
		_w4221_,
		_w4222_,
		_w4223_
	);
	LUT2 #(
		.INIT('h4)
	) name2716 (
		_w4220_,
		_w4223_,
		_w4224_
	);
	LUT2 #(
		.INIT('h2)
	) name2717 (
		_w4220_,
		_w4223_,
		_w4225_
	);
	LUT2 #(
		.INIT('h1)
	) name2718 (
		\TM0_pad ,
		_w4224_,
		_w4226_
	);
	LUT2 #(
		.INIT('h4)
	) name2719 (
		_w4225_,
		_w4226_,
		_w4227_
	);
	LUT2 #(
		.INIT('h1)
	) name2720 (
		_w4214_,
		_w4227_,
		_w4228_
	);
	LUT2 #(
		.INIT('h2)
	) name2721 (
		_w1976_,
		_w4228_,
		_w4229_
	);
	LUT2 #(
		.INIT('h1)
	) name2722 (
		_w4213_,
		_w4229_,
		_w4230_
	);
	LUT2 #(
		.INIT('h1)
	) name2723 (
		_w1637_,
		_w2594_,
		_w4231_
	);
	LUT2 #(
		.INIT('h2)
	) name2724 (
		_w1973_,
		_w4231_,
		_w4232_
	);
	LUT2 #(
		.INIT('h1)
	) name2725 (
		\DATA_0_18_pad ,
		\TM0_pad ,
		_w4233_
	);
	LUT2 #(
		.INIT('h2)
	) name2726 (
		\TM0_pad ,
		\_2351__reg/NET0131 ,
		_w4234_
	);
	LUT2 #(
		.INIT('h2)
	) name2727 (
		_w1976_,
		_w4233_,
		_w4235_
	);
	LUT2 #(
		.INIT('h4)
	) name2728 (
		_w4234_,
		_w4235_,
		_w4236_
	);
	LUT2 #(
		.INIT('h1)
	) name2729 (
		_w4232_,
		_w4236_,
		_w4237_
	);
	LUT2 #(
		.INIT('h8)
	) name2730 (
		RESET_pad,
		\WX10853_reg/NET0131 ,
		_w4238_
	);
	LUT2 #(
		.INIT('h4)
	) name2731 (
		_w1836_,
		_w1973_,
		_w4239_
	);
	LUT2 #(
		.INIT('h2)
	) name2732 (
		\WX3417_reg/NET0131 ,
		\WX3481_reg/NET0131 ,
		_w4240_
	);
	LUT2 #(
		.INIT('h4)
	) name2733 (
		\WX3417_reg/NET0131 ,
		\WX3481_reg/NET0131 ,
		_w4241_
	);
	LUT2 #(
		.INIT('h1)
	) name2734 (
		_w4240_,
		_w4241_,
		_w4242_
	);
	LUT2 #(
		.INIT('h2)
	) name2735 (
		\WX3289_reg/NET0131 ,
		\WX3353_reg/NET0131 ,
		_w4243_
	);
	LUT2 #(
		.INIT('h4)
	) name2736 (
		\WX3289_reg/NET0131 ,
		\WX3353_reg/NET0131 ,
		_w4244_
	);
	LUT2 #(
		.INIT('h1)
	) name2737 (
		_w4243_,
		_w4244_,
		_w4245_
	);
	LUT2 #(
		.INIT('h4)
	) name2738 (
		_w4242_,
		_w4245_,
		_w4246_
	);
	LUT2 #(
		.INIT('h2)
	) name2739 (
		_w4242_,
		_w4245_,
		_w4247_
	);
	LUT2 #(
		.INIT('h1)
	) name2740 (
		\TM0_pad ,
		_w4246_,
		_w4248_
	);
	LUT2 #(
		.INIT('h4)
	) name2741 (
		_w4247_,
		_w4248_,
		_w4249_
	);
	LUT2 #(
		.INIT('h2)
	) name2742 (
		_w4239_,
		_w4249_,
		_w4250_
	);
	LUT2 #(
		.INIT('h2)
	) name2743 (
		\TM0_pad ,
		\_2143__reg/NET0131 ,
		_w4251_
	);
	LUT2 #(
		.INIT('h2)
	) name2744 (
		\WX4710_reg/NET0131 ,
		\WX4774_reg/NET0131 ,
		_w4252_
	);
	LUT2 #(
		.INIT('h4)
	) name2745 (
		\WX4710_reg/NET0131 ,
		\WX4774_reg/NET0131 ,
		_w4253_
	);
	LUT2 #(
		.INIT('h1)
	) name2746 (
		_w4252_,
		_w4253_,
		_w4254_
	);
	LUT2 #(
		.INIT('h2)
	) name2747 (
		\WX4582_reg/NET0131 ,
		\WX4646_reg/NET0131 ,
		_w4255_
	);
	LUT2 #(
		.INIT('h4)
	) name2748 (
		\WX4582_reg/NET0131 ,
		\WX4646_reg/NET0131 ,
		_w4256_
	);
	LUT2 #(
		.INIT('h1)
	) name2749 (
		_w4255_,
		_w4256_,
		_w4257_
	);
	LUT2 #(
		.INIT('h4)
	) name2750 (
		_w4254_,
		_w4257_,
		_w4258_
	);
	LUT2 #(
		.INIT('h2)
	) name2751 (
		_w4254_,
		_w4257_,
		_w4259_
	);
	LUT2 #(
		.INIT('h1)
	) name2752 (
		\TM0_pad ,
		_w4258_,
		_w4260_
	);
	LUT2 #(
		.INIT('h4)
	) name2753 (
		_w4259_,
		_w4260_,
		_w4261_
	);
	LUT2 #(
		.INIT('h2)
	) name2754 (
		_w1976_,
		_w4251_,
		_w4262_
	);
	LUT2 #(
		.INIT('h4)
	) name2755 (
		_w4261_,
		_w4262_,
		_w4263_
	);
	LUT2 #(
		.INIT('h1)
	) name2756 (
		_w4250_,
		_w4263_,
		_w4264_
	);
	LUT2 #(
		.INIT('h2)
	) name2757 (
		_w3644_,
		_w4207_,
		_w4265_
	);
	LUT2 #(
		.INIT('h2)
	) name2758 (
		\TM0_pad ,
		\_2275__reg/NET0131 ,
		_w4266_
	);
	LUT2 #(
		.INIT('h2)
	) name2759 (
		\WX9874_reg/NET0131 ,
		\WX9938_reg/NET0131 ,
		_w4267_
	);
	LUT2 #(
		.INIT('h4)
	) name2760 (
		\WX9874_reg/NET0131 ,
		\WX9938_reg/NET0131 ,
		_w4268_
	);
	LUT2 #(
		.INIT('h1)
	) name2761 (
		_w4267_,
		_w4268_,
		_w4269_
	);
	LUT2 #(
		.INIT('h2)
	) name2762 (
		\WX9746_reg/NET0131 ,
		\WX9810_reg/NET0131 ,
		_w4270_
	);
	LUT2 #(
		.INIT('h4)
	) name2763 (
		\WX9746_reg/NET0131 ,
		\WX9810_reg/NET0131 ,
		_w4271_
	);
	LUT2 #(
		.INIT('h1)
	) name2764 (
		_w4270_,
		_w4271_,
		_w4272_
	);
	LUT2 #(
		.INIT('h4)
	) name2765 (
		_w4269_,
		_w4272_,
		_w4273_
	);
	LUT2 #(
		.INIT('h2)
	) name2766 (
		_w4269_,
		_w4272_,
		_w4274_
	);
	LUT2 #(
		.INIT('h1)
	) name2767 (
		\TM0_pad ,
		_w4273_,
		_w4275_
	);
	LUT2 #(
		.INIT('h4)
	) name2768 (
		_w4274_,
		_w4275_,
		_w4276_
	);
	LUT2 #(
		.INIT('h2)
	) name2769 (
		_w1976_,
		_w4266_,
		_w4277_
	);
	LUT2 #(
		.INIT('h4)
	) name2770 (
		_w4276_,
		_w4277_,
		_w4278_
	);
	LUT2 #(
		.INIT('h1)
	) name2771 (
		_w4265_,
		_w4278_,
		_w4279_
	);
	LUT2 #(
		.INIT('h2)
	) name2772 (
		_w3483_,
		_w4138_,
		_w4280_
	);
	LUT2 #(
		.INIT('h2)
	) name2773 (
		\TM0_pad ,
		\_2308__reg/NET0131 ,
		_w4281_
	);
	LUT2 #(
		.INIT('h2)
	) name2774 (
		\WX11165_reg/NET0131 ,
		\WX11229_reg/NET0131 ,
		_w4282_
	);
	LUT2 #(
		.INIT('h4)
	) name2775 (
		\WX11165_reg/NET0131 ,
		\WX11229_reg/NET0131 ,
		_w4283_
	);
	LUT2 #(
		.INIT('h1)
	) name2776 (
		_w4282_,
		_w4283_,
		_w4284_
	);
	LUT2 #(
		.INIT('h2)
	) name2777 (
		\WX11037_reg/NET0131 ,
		\WX11101_reg/NET0131 ,
		_w4285_
	);
	LUT2 #(
		.INIT('h4)
	) name2778 (
		\WX11037_reg/NET0131 ,
		\WX11101_reg/NET0131 ,
		_w4286_
	);
	LUT2 #(
		.INIT('h1)
	) name2779 (
		_w4285_,
		_w4286_,
		_w4287_
	);
	LUT2 #(
		.INIT('h4)
	) name2780 (
		_w4284_,
		_w4287_,
		_w4288_
	);
	LUT2 #(
		.INIT('h2)
	) name2781 (
		_w4284_,
		_w4287_,
		_w4289_
	);
	LUT2 #(
		.INIT('h1)
	) name2782 (
		\TM0_pad ,
		_w4288_,
		_w4290_
	);
	LUT2 #(
		.INIT('h4)
	) name2783 (
		_w4289_,
		_w4290_,
		_w4291_
	);
	LUT2 #(
		.INIT('h2)
	) name2784 (
		_w1976_,
		_w4281_,
		_w4292_
	);
	LUT2 #(
		.INIT('h4)
	) name2785 (
		_w4291_,
		_w4292_,
		_w4293_
	);
	LUT2 #(
		.INIT('h1)
	) name2786 (
		_w4280_,
		_w4293_,
		_w4294_
	);
	LUT2 #(
		.INIT('h2)
	) name2787 (
		_w4101_,
		_w4123_,
		_w4295_
	);
	LUT2 #(
		.INIT('h2)
	) name2788 (
		\TM0_pad ,
		\_2176__reg/NET0131 ,
		_w4296_
	);
	LUT2 #(
		.INIT('h2)
	) name2789 (
		\WX6001_reg/NET0131 ,
		\WX6065_reg/NET0131 ,
		_w4297_
	);
	LUT2 #(
		.INIT('h4)
	) name2790 (
		\WX6001_reg/NET0131 ,
		\WX6065_reg/NET0131 ,
		_w4298_
	);
	LUT2 #(
		.INIT('h1)
	) name2791 (
		_w4297_,
		_w4298_,
		_w4299_
	);
	LUT2 #(
		.INIT('h2)
	) name2792 (
		\WX5873_reg/NET0131 ,
		\WX5937_reg/NET0131 ,
		_w4300_
	);
	LUT2 #(
		.INIT('h4)
	) name2793 (
		\WX5873_reg/NET0131 ,
		\WX5937_reg/NET0131 ,
		_w4301_
	);
	LUT2 #(
		.INIT('h1)
	) name2794 (
		_w4300_,
		_w4301_,
		_w4302_
	);
	LUT2 #(
		.INIT('h4)
	) name2795 (
		_w4299_,
		_w4302_,
		_w4303_
	);
	LUT2 #(
		.INIT('h2)
	) name2796 (
		_w4299_,
		_w4302_,
		_w4304_
	);
	LUT2 #(
		.INIT('h1)
	) name2797 (
		\TM0_pad ,
		_w4303_,
		_w4305_
	);
	LUT2 #(
		.INIT('h4)
	) name2798 (
		_w4304_,
		_w4305_,
		_w4306_
	);
	LUT2 #(
		.INIT('h2)
	) name2799 (
		_w1976_,
		_w4296_,
		_w4307_
	);
	LUT2 #(
		.INIT('h4)
	) name2800 (
		_w4306_,
		_w4307_,
		_w4308_
	);
	LUT2 #(
		.INIT('h1)
	) name2801 (
		_w4295_,
		_w4308_,
		_w4309_
	);
	LUT2 #(
		.INIT('h8)
	) name2802 (
		\TM0_pad ,
		\_2126__reg/NET0131 ,
		_w4310_
	);
	LUT2 #(
		.INIT('h2)
	) name2803 (
		\WX3387_reg/NET0131 ,
		\WX3451_reg/NET0131 ,
		_w4311_
	);
	LUT2 #(
		.INIT('h4)
	) name2804 (
		\WX3387_reg/NET0131 ,
		\WX3451_reg/NET0131 ,
		_w4312_
	);
	LUT2 #(
		.INIT('h1)
	) name2805 (
		_w4311_,
		_w4312_,
		_w4313_
	);
	LUT2 #(
		.INIT('h2)
	) name2806 (
		\WX3323_reg/NET0131 ,
		_w4313_,
		_w4314_
	);
	LUT2 #(
		.INIT('h4)
	) name2807 (
		\WX3323_reg/NET0131 ,
		_w4313_,
		_w4315_
	);
	LUT2 #(
		.INIT('h1)
	) name2808 (
		_w4314_,
		_w4315_,
		_w4316_
	);
	LUT2 #(
		.INIT('h2)
	) name2809 (
		\TM1_pad ,
		\WX3259_reg/NET0131 ,
		_w4317_
	);
	LUT2 #(
		.INIT('h4)
	) name2810 (
		\TM1_pad ,
		\WX3259_reg/NET0131 ,
		_w4318_
	);
	LUT2 #(
		.INIT('h1)
	) name2811 (
		_w4317_,
		_w4318_,
		_w4319_
	);
	LUT2 #(
		.INIT('h4)
	) name2812 (
		_w4316_,
		_w4319_,
		_w4320_
	);
	LUT2 #(
		.INIT('h2)
	) name2813 (
		_w4316_,
		_w4319_,
		_w4321_
	);
	LUT2 #(
		.INIT('h1)
	) name2814 (
		\TM0_pad ,
		_w4320_,
		_w4322_
	);
	LUT2 #(
		.INIT('h4)
	) name2815 (
		_w4321_,
		_w4322_,
		_w4323_
	);
	LUT2 #(
		.INIT('h1)
	) name2816 (
		_w4310_,
		_w4323_,
		_w4324_
	);
	LUT2 #(
		.INIT('h2)
	) name2817 (
		_w1976_,
		_w4324_,
		_w4325_
	);
	LUT2 #(
		.INIT('h1)
	) name2818 (
		_w1621_,
		_w4086_,
		_w4326_
	);
	LUT2 #(
		.INIT('h2)
	) name2819 (
		_w1973_,
		_w4326_,
		_w4327_
	);
	LUT2 #(
		.INIT('h1)
	) name2820 (
		_w4325_,
		_w4327_,
		_w4328_
	);
	LUT2 #(
		.INIT('h2)
	) name2821 (
		_w3953_,
		_w4177_,
		_w4329_
	);
	LUT2 #(
		.INIT('h2)
	) name2822 (
		\TM0_pad ,
		\_2209__reg/NET0131 ,
		_w4330_
	);
	LUT2 #(
		.INIT('h2)
	) name2823 (
		\WX7292_reg/NET0131 ,
		\WX7356_reg/NET0131 ,
		_w4331_
	);
	LUT2 #(
		.INIT('h4)
	) name2824 (
		\WX7292_reg/NET0131 ,
		\WX7356_reg/NET0131 ,
		_w4332_
	);
	LUT2 #(
		.INIT('h1)
	) name2825 (
		_w4331_,
		_w4332_,
		_w4333_
	);
	LUT2 #(
		.INIT('h2)
	) name2826 (
		\WX7164_reg/NET0131 ,
		\WX7228_reg/NET0131 ,
		_w4334_
	);
	LUT2 #(
		.INIT('h4)
	) name2827 (
		\WX7164_reg/NET0131 ,
		\WX7228_reg/NET0131 ,
		_w4335_
	);
	LUT2 #(
		.INIT('h1)
	) name2828 (
		_w4334_,
		_w4335_,
		_w4336_
	);
	LUT2 #(
		.INIT('h4)
	) name2829 (
		_w4333_,
		_w4336_,
		_w4337_
	);
	LUT2 #(
		.INIT('h2)
	) name2830 (
		_w4333_,
		_w4336_,
		_w4338_
	);
	LUT2 #(
		.INIT('h1)
	) name2831 (
		\TM0_pad ,
		_w4337_,
		_w4339_
	);
	LUT2 #(
		.INIT('h4)
	) name2832 (
		_w4338_,
		_w4339_,
		_w4340_
	);
	LUT2 #(
		.INIT('h2)
	) name2833 (
		_w1976_,
		_w4330_,
		_w4341_
	);
	LUT2 #(
		.INIT('h4)
	) name2834 (
		_w4340_,
		_w4341_,
		_w4342_
	);
	LUT2 #(
		.INIT('h1)
	) name2835 (
		_w4329_,
		_w4342_,
		_w4343_
	);
	LUT2 #(
		.INIT('h2)
	) name2836 (
		_w3805_,
		_w4192_,
		_w4344_
	);
	LUT2 #(
		.INIT('h2)
	) name2837 (
		\TM0_pad ,
		\_2242__reg/NET0131 ,
		_w4345_
	);
	LUT2 #(
		.INIT('h2)
	) name2838 (
		\WX8583_reg/NET0131 ,
		\WX8647_reg/NET0131 ,
		_w4346_
	);
	LUT2 #(
		.INIT('h4)
	) name2839 (
		\WX8583_reg/NET0131 ,
		\WX8647_reg/NET0131 ,
		_w4347_
	);
	LUT2 #(
		.INIT('h1)
	) name2840 (
		_w4346_,
		_w4347_,
		_w4348_
	);
	LUT2 #(
		.INIT('h2)
	) name2841 (
		\WX8455_reg/NET0131 ,
		\WX8519_reg/NET0131 ,
		_w4349_
	);
	LUT2 #(
		.INIT('h4)
	) name2842 (
		\WX8455_reg/NET0131 ,
		\WX8519_reg/NET0131 ,
		_w4350_
	);
	LUT2 #(
		.INIT('h1)
	) name2843 (
		_w4349_,
		_w4350_,
		_w4351_
	);
	LUT2 #(
		.INIT('h4)
	) name2844 (
		_w4348_,
		_w4351_,
		_w4352_
	);
	LUT2 #(
		.INIT('h2)
	) name2845 (
		_w4348_,
		_w4351_,
		_w4353_
	);
	LUT2 #(
		.INIT('h1)
	) name2846 (
		\TM0_pad ,
		_w4352_,
		_w4354_
	);
	LUT2 #(
		.INIT('h4)
	) name2847 (
		_w4353_,
		_w4354_,
		_w4355_
	);
	LUT2 #(
		.INIT('h2)
	) name2848 (
		_w1976_,
		_w4345_,
		_w4356_
	);
	LUT2 #(
		.INIT('h4)
	) name2849 (
		_w4355_,
		_w4356_,
		_w4357_
	);
	LUT2 #(
		.INIT('h1)
	) name2850 (
		_w4344_,
		_w4357_,
		_w4358_
	);
	LUT2 #(
		.INIT('h1)
	) name2851 (
		_w1621_,
		_w2754_,
		_w4359_
	);
	LUT2 #(
		.INIT('h2)
	) name2852 (
		_w1973_,
		_w4359_,
		_w4360_
	);
	LUT2 #(
		.INIT('h1)
	) name2853 (
		\DATA_0_17_pad ,
		\TM0_pad ,
		_w4361_
	);
	LUT2 #(
		.INIT('h2)
	) name2854 (
		\TM0_pad ,
		\_2350__reg/NET0131 ,
		_w4362_
	);
	LUT2 #(
		.INIT('h2)
	) name2855 (
		_w1976_,
		_w4361_,
		_w4363_
	);
	LUT2 #(
		.INIT('h4)
	) name2856 (
		_w4362_,
		_w4363_,
		_w4364_
	);
	LUT2 #(
		.INIT('h1)
	) name2857 (
		_w4360_,
		_w4364_,
		_w4365_
	);
	LUT2 #(
		.INIT('h8)
	) name2858 (
		RESET_pad,
		\WX10855_reg/NET0131 ,
		_w4366_
	);
	LUT2 #(
		.INIT('h2)
	) name2859 (
		_w3953_,
		_w4340_,
		_w4367_
	);
	LUT2 #(
		.INIT('h2)
	) name2860 (
		\TM0_pad ,
		\_2241__reg/NET0131 ,
		_w4368_
	);
	LUT2 #(
		.INIT('h2)
	) name2861 (
		\WX8585_reg/NET0131 ,
		\WX8649_reg/NET0131 ,
		_w4369_
	);
	LUT2 #(
		.INIT('h4)
	) name2862 (
		\WX8585_reg/NET0131 ,
		\WX8649_reg/NET0131 ,
		_w4370_
	);
	LUT2 #(
		.INIT('h1)
	) name2863 (
		_w4369_,
		_w4370_,
		_w4371_
	);
	LUT2 #(
		.INIT('h2)
	) name2864 (
		\WX8457_reg/NET0131 ,
		\WX8521_reg/NET0131 ,
		_w4372_
	);
	LUT2 #(
		.INIT('h4)
	) name2865 (
		\WX8457_reg/NET0131 ,
		\WX8521_reg/NET0131 ,
		_w4373_
	);
	LUT2 #(
		.INIT('h1)
	) name2866 (
		_w4372_,
		_w4373_,
		_w4374_
	);
	LUT2 #(
		.INIT('h4)
	) name2867 (
		_w4371_,
		_w4374_,
		_w4375_
	);
	LUT2 #(
		.INIT('h2)
	) name2868 (
		_w4371_,
		_w4374_,
		_w4376_
	);
	LUT2 #(
		.INIT('h1)
	) name2869 (
		\TM0_pad ,
		_w4375_,
		_w4377_
	);
	LUT2 #(
		.INIT('h4)
	) name2870 (
		_w4376_,
		_w4377_,
		_w4378_
	);
	LUT2 #(
		.INIT('h2)
	) name2871 (
		_w1976_,
		_w4368_,
		_w4379_
	);
	LUT2 #(
		.INIT('h4)
	) name2872 (
		_w4378_,
		_w4379_,
		_w4380_
	);
	LUT2 #(
		.INIT('h1)
	) name2873 (
		_w4367_,
		_w4380_,
		_w4381_
	);
	LUT2 #(
		.INIT('h4)
	) name2874 (
		_w1663_,
		_w1973_,
		_w4382_
	);
	LUT2 #(
		.INIT('h2)
	) name2875 (
		\WX3419_reg/NET0131 ,
		\WX3483_reg/NET0131 ,
		_w4383_
	);
	LUT2 #(
		.INIT('h4)
	) name2876 (
		\WX3419_reg/NET0131 ,
		\WX3483_reg/NET0131 ,
		_w4384_
	);
	LUT2 #(
		.INIT('h1)
	) name2877 (
		_w4383_,
		_w4384_,
		_w4385_
	);
	LUT2 #(
		.INIT('h2)
	) name2878 (
		\WX3291_reg/NET0131 ,
		\WX3355_reg/NET0131 ,
		_w4386_
	);
	LUT2 #(
		.INIT('h4)
	) name2879 (
		\WX3291_reg/NET0131 ,
		\WX3355_reg/NET0131 ,
		_w4387_
	);
	LUT2 #(
		.INIT('h1)
	) name2880 (
		_w4386_,
		_w4387_,
		_w4388_
	);
	LUT2 #(
		.INIT('h4)
	) name2881 (
		_w4385_,
		_w4388_,
		_w4389_
	);
	LUT2 #(
		.INIT('h2)
	) name2882 (
		_w4385_,
		_w4388_,
		_w4390_
	);
	LUT2 #(
		.INIT('h1)
	) name2883 (
		\TM0_pad ,
		_w4389_,
		_w4391_
	);
	LUT2 #(
		.INIT('h4)
	) name2884 (
		_w4390_,
		_w4391_,
		_w4392_
	);
	LUT2 #(
		.INIT('h2)
	) name2885 (
		_w4382_,
		_w4392_,
		_w4393_
	);
	LUT2 #(
		.INIT('h2)
	) name2886 (
		\TM0_pad ,
		\_2142__reg/NET0131 ,
		_w4394_
	);
	LUT2 #(
		.INIT('h2)
	) name2887 (
		\WX4712_reg/NET0131 ,
		\WX4776_reg/NET0131 ,
		_w4395_
	);
	LUT2 #(
		.INIT('h4)
	) name2888 (
		\WX4712_reg/NET0131 ,
		\WX4776_reg/NET0131 ,
		_w4396_
	);
	LUT2 #(
		.INIT('h1)
	) name2889 (
		_w4395_,
		_w4396_,
		_w4397_
	);
	LUT2 #(
		.INIT('h2)
	) name2890 (
		\WX4584_reg/NET0131 ,
		\WX4648_reg/NET0131 ,
		_w4398_
	);
	LUT2 #(
		.INIT('h4)
	) name2891 (
		\WX4584_reg/NET0131 ,
		\WX4648_reg/NET0131 ,
		_w4399_
	);
	LUT2 #(
		.INIT('h1)
	) name2892 (
		_w4398_,
		_w4399_,
		_w4400_
	);
	LUT2 #(
		.INIT('h4)
	) name2893 (
		_w4397_,
		_w4400_,
		_w4401_
	);
	LUT2 #(
		.INIT('h2)
	) name2894 (
		_w4397_,
		_w4400_,
		_w4402_
	);
	LUT2 #(
		.INIT('h1)
	) name2895 (
		\TM0_pad ,
		_w4401_,
		_w4403_
	);
	LUT2 #(
		.INIT('h4)
	) name2896 (
		_w4402_,
		_w4403_,
		_w4404_
	);
	LUT2 #(
		.INIT('h2)
	) name2897 (
		_w1976_,
		_w4394_,
		_w4405_
	);
	LUT2 #(
		.INIT('h4)
	) name2898 (
		_w4404_,
		_w4405_,
		_w4406_
	);
	LUT2 #(
		.INIT('h1)
	) name2899 (
		_w4393_,
		_w4406_,
		_w4407_
	);
	LUT2 #(
		.INIT('h2)
	) name2900 (
		_w3805_,
		_w4355_,
		_w4408_
	);
	LUT2 #(
		.INIT('h2)
	) name2901 (
		\TM0_pad ,
		\_2274__reg/NET0131 ,
		_w4409_
	);
	LUT2 #(
		.INIT('h2)
	) name2902 (
		\WX9876_reg/NET0131 ,
		\WX9940_reg/NET0131 ,
		_w4410_
	);
	LUT2 #(
		.INIT('h4)
	) name2903 (
		\WX9876_reg/NET0131 ,
		\WX9940_reg/NET0131 ,
		_w4411_
	);
	LUT2 #(
		.INIT('h1)
	) name2904 (
		_w4410_,
		_w4411_,
		_w4412_
	);
	LUT2 #(
		.INIT('h2)
	) name2905 (
		\WX9748_reg/NET0131 ,
		\WX9812_reg/NET0131 ,
		_w4413_
	);
	LUT2 #(
		.INIT('h4)
	) name2906 (
		\WX9748_reg/NET0131 ,
		\WX9812_reg/NET0131 ,
		_w4414_
	);
	LUT2 #(
		.INIT('h1)
	) name2907 (
		_w4413_,
		_w4414_,
		_w4415_
	);
	LUT2 #(
		.INIT('h4)
	) name2908 (
		_w4412_,
		_w4415_,
		_w4416_
	);
	LUT2 #(
		.INIT('h2)
	) name2909 (
		_w4412_,
		_w4415_,
		_w4417_
	);
	LUT2 #(
		.INIT('h1)
	) name2910 (
		\TM0_pad ,
		_w4416_,
		_w4418_
	);
	LUT2 #(
		.INIT('h4)
	) name2911 (
		_w4417_,
		_w4418_,
		_w4419_
	);
	LUT2 #(
		.INIT('h2)
	) name2912 (
		_w1976_,
		_w4409_,
		_w4420_
	);
	LUT2 #(
		.INIT('h4)
	) name2913 (
		_w4419_,
		_w4420_,
		_w4421_
	);
	LUT2 #(
		.INIT('h1)
	) name2914 (
		_w4408_,
		_w4421_,
		_w4422_
	);
	LUT2 #(
		.INIT('h2)
	) name2915 (
		_w3644_,
		_w4276_,
		_w4423_
	);
	LUT2 #(
		.INIT('h2)
	) name2916 (
		\TM0_pad ,
		\_2307__reg/NET0131 ,
		_w4424_
	);
	LUT2 #(
		.INIT('h2)
	) name2917 (
		\WX11167_reg/NET0131 ,
		\WX11231_reg/NET0131 ,
		_w4425_
	);
	LUT2 #(
		.INIT('h4)
	) name2918 (
		\WX11167_reg/NET0131 ,
		\WX11231_reg/NET0131 ,
		_w4426_
	);
	LUT2 #(
		.INIT('h1)
	) name2919 (
		_w4425_,
		_w4426_,
		_w4427_
	);
	LUT2 #(
		.INIT('h2)
	) name2920 (
		\WX11039_reg/NET0131 ,
		\WX11103_reg/NET0131 ,
		_w4428_
	);
	LUT2 #(
		.INIT('h4)
	) name2921 (
		\WX11039_reg/NET0131 ,
		\WX11103_reg/NET0131 ,
		_w4429_
	);
	LUT2 #(
		.INIT('h1)
	) name2922 (
		_w4428_,
		_w4429_,
		_w4430_
	);
	LUT2 #(
		.INIT('h4)
	) name2923 (
		_w4427_,
		_w4430_,
		_w4431_
	);
	LUT2 #(
		.INIT('h2)
	) name2924 (
		_w4427_,
		_w4430_,
		_w4432_
	);
	LUT2 #(
		.INIT('h1)
	) name2925 (
		\TM0_pad ,
		_w4431_,
		_w4433_
	);
	LUT2 #(
		.INIT('h4)
	) name2926 (
		_w4432_,
		_w4433_,
		_w4434_
	);
	LUT2 #(
		.INIT('h2)
	) name2927 (
		_w1976_,
		_w4424_,
		_w4435_
	);
	LUT2 #(
		.INIT('h4)
	) name2928 (
		_w4434_,
		_w4435_,
		_w4436_
	);
	LUT2 #(
		.INIT('h1)
	) name2929 (
		_w4423_,
		_w4436_,
		_w4437_
	);
	LUT2 #(
		.INIT('h2)
	) name2930 (
		_w4239_,
		_w4261_,
		_w4438_
	);
	LUT2 #(
		.INIT('h2)
	) name2931 (
		\TM0_pad ,
		\_2175__reg/NET0131 ,
		_w4439_
	);
	LUT2 #(
		.INIT('h2)
	) name2932 (
		\WX6003_reg/NET0131 ,
		\WX6067_reg/NET0131 ,
		_w4440_
	);
	LUT2 #(
		.INIT('h4)
	) name2933 (
		\WX6003_reg/NET0131 ,
		\WX6067_reg/NET0131 ,
		_w4441_
	);
	LUT2 #(
		.INIT('h1)
	) name2934 (
		_w4440_,
		_w4441_,
		_w4442_
	);
	LUT2 #(
		.INIT('h2)
	) name2935 (
		\WX5875_reg/NET0131 ,
		\WX5939_reg/NET0131 ,
		_w4443_
	);
	LUT2 #(
		.INIT('h4)
	) name2936 (
		\WX5875_reg/NET0131 ,
		\WX5939_reg/NET0131 ,
		_w4444_
	);
	LUT2 #(
		.INIT('h1)
	) name2937 (
		_w4443_,
		_w4444_,
		_w4445_
	);
	LUT2 #(
		.INIT('h4)
	) name2938 (
		_w4442_,
		_w4445_,
		_w4446_
	);
	LUT2 #(
		.INIT('h2)
	) name2939 (
		_w4442_,
		_w4445_,
		_w4447_
	);
	LUT2 #(
		.INIT('h1)
	) name2940 (
		\TM0_pad ,
		_w4446_,
		_w4448_
	);
	LUT2 #(
		.INIT('h4)
	) name2941 (
		_w4447_,
		_w4448_,
		_w4449_
	);
	LUT2 #(
		.INIT('h2)
	) name2942 (
		_w1976_,
		_w4439_,
		_w4450_
	);
	LUT2 #(
		.INIT('h4)
	) name2943 (
		_w4449_,
		_w4450_,
		_w4451_
	);
	LUT2 #(
		.INIT('h1)
	) name2944 (
		_w4438_,
		_w4451_,
		_w4452_
	);
	LUT2 #(
		.INIT('h8)
	) name2945 (
		\TM0_pad ,
		\_2125__reg/NET0131 ,
		_w4453_
	);
	LUT2 #(
		.INIT('h2)
	) name2946 (
		\WX3389_reg/NET0131 ,
		\WX3453_reg/NET0131 ,
		_w4454_
	);
	LUT2 #(
		.INIT('h4)
	) name2947 (
		\WX3389_reg/NET0131 ,
		\WX3453_reg/NET0131 ,
		_w4455_
	);
	LUT2 #(
		.INIT('h1)
	) name2948 (
		_w4454_,
		_w4455_,
		_w4456_
	);
	LUT2 #(
		.INIT('h2)
	) name2949 (
		\WX3325_reg/NET0131 ,
		_w4456_,
		_w4457_
	);
	LUT2 #(
		.INIT('h4)
	) name2950 (
		\WX3325_reg/NET0131 ,
		_w4456_,
		_w4458_
	);
	LUT2 #(
		.INIT('h1)
	) name2951 (
		_w4457_,
		_w4458_,
		_w4459_
	);
	LUT2 #(
		.INIT('h2)
	) name2952 (
		\TM1_pad ,
		\WX3261_reg/NET0131 ,
		_w4460_
	);
	LUT2 #(
		.INIT('h4)
	) name2953 (
		\TM1_pad ,
		\WX3261_reg/NET0131 ,
		_w4461_
	);
	LUT2 #(
		.INIT('h1)
	) name2954 (
		_w4460_,
		_w4461_,
		_w4462_
	);
	LUT2 #(
		.INIT('h4)
	) name2955 (
		_w4459_,
		_w4462_,
		_w4463_
	);
	LUT2 #(
		.INIT('h2)
	) name2956 (
		_w4459_,
		_w4462_,
		_w4464_
	);
	LUT2 #(
		.INIT('h1)
	) name2957 (
		\TM0_pad ,
		_w4463_,
		_w4465_
	);
	LUT2 #(
		.INIT('h4)
	) name2958 (
		_w4464_,
		_w4465_,
		_w4466_
	);
	LUT2 #(
		.INIT('h1)
	) name2959 (
		_w4453_,
		_w4466_,
		_w4467_
	);
	LUT2 #(
		.INIT('h2)
	) name2960 (
		_w1976_,
		_w4467_,
		_w4468_
	);
	LUT2 #(
		.INIT('h1)
	) name2961 (
		_w1605_,
		_w4227_,
		_w4469_
	);
	LUT2 #(
		.INIT('h2)
	) name2962 (
		_w1973_,
		_w4469_,
		_w4470_
	);
	LUT2 #(
		.INIT('h1)
	) name2963 (
		_w4468_,
		_w4470_,
		_w4471_
	);
	LUT2 #(
		.INIT('h2)
	) name2964 (
		_w4101_,
		_w4306_,
		_w4472_
	);
	LUT2 #(
		.INIT('h2)
	) name2965 (
		\TM0_pad ,
		\_2208__reg/NET0131 ,
		_w4473_
	);
	LUT2 #(
		.INIT('h2)
	) name2966 (
		\WX7294_reg/NET0131 ,
		\WX7358_reg/NET0131 ,
		_w4474_
	);
	LUT2 #(
		.INIT('h4)
	) name2967 (
		\WX7294_reg/NET0131 ,
		\WX7358_reg/NET0131 ,
		_w4475_
	);
	LUT2 #(
		.INIT('h1)
	) name2968 (
		_w4474_,
		_w4475_,
		_w4476_
	);
	LUT2 #(
		.INIT('h2)
	) name2969 (
		\WX7166_reg/NET0131 ,
		\WX7230_reg/NET0131 ,
		_w4477_
	);
	LUT2 #(
		.INIT('h4)
	) name2970 (
		\WX7166_reg/NET0131 ,
		\WX7230_reg/NET0131 ,
		_w4478_
	);
	LUT2 #(
		.INIT('h1)
	) name2971 (
		_w4477_,
		_w4478_,
		_w4479_
	);
	LUT2 #(
		.INIT('h4)
	) name2972 (
		_w4476_,
		_w4479_,
		_w4480_
	);
	LUT2 #(
		.INIT('h2)
	) name2973 (
		_w4476_,
		_w4479_,
		_w4481_
	);
	LUT2 #(
		.INIT('h1)
	) name2974 (
		\TM0_pad ,
		_w4480_,
		_w4482_
	);
	LUT2 #(
		.INIT('h4)
	) name2975 (
		_w4481_,
		_w4482_,
		_w4483_
	);
	LUT2 #(
		.INIT('h2)
	) name2976 (
		_w1976_,
		_w4473_,
		_w4484_
	);
	LUT2 #(
		.INIT('h4)
	) name2977 (
		_w4483_,
		_w4484_,
		_w4485_
	);
	LUT2 #(
		.INIT('h1)
	) name2978 (
		_w4472_,
		_w4485_,
		_w4486_
	);
	LUT2 #(
		.INIT('h1)
	) name2979 (
		_w1605_,
		_w2919_,
		_w4487_
	);
	LUT2 #(
		.INIT('h2)
	) name2980 (
		_w1973_,
		_w4487_,
		_w4488_
	);
	LUT2 #(
		.INIT('h1)
	) name2981 (
		\DATA_0_16_pad ,
		\TM0_pad ,
		_w4489_
	);
	LUT2 #(
		.INIT('h2)
	) name2982 (
		\TM0_pad ,
		\_2349__reg/NET0131 ,
		_w4490_
	);
	LUT2 #(
		.INIT('h2)
	) name2983 (
		_w1976_,
		_w4489_,
		_w4491_
	);
	LUT2 #(
		.INIT('h4)
	) name2984 (
		_w4490_,
		_w4491_,
		_w4492_
	);
	LUT2 #(
		.INIT('h1)
	) name2985 (
		_w4488_,
		_w4492_,
		_w4493_
	);
	LUT2 #(
		.INIT('h8)
	) name2986 (
		RESET_pad,
		\WX10857_reg/NET0131 ,
		_w4494_
	);
	LUT2 #(
		.INIT('h2)
	) name2987 (
		_w4101_,
		_w4483_,
		_w4495_
	);
	LUT2 #(
		.INIT('h2)
	) name2988 (
		\TM0_pad ,
		\_2240__reg/NET0131 ,
		_w4496_
	);
	LUT2 #(
		.INIT('h2)
	) name2989 (
		\WX8587_reg/NET0131 ,
		\WX8651_reg/NET0131 ,
		_w4497_
	);
	LUT2 #(
		.INIT('h4)
	) name2990 (
		\WX8587_reg/NET0131 ,
		\WX8651_reg/NET0131 ,
		_w4498_
	);
	LUT2 #(
		.INIT('h1)
	) name2991 (
		_w4497_,
		_w4498_,
		_w4499_
	);
	LUT2 #(
		.INIT('h2)
	) name2992 (
		\WX8459_reg/NET0131 ,
		\WX8523_reg/NET0131 ,
		_w4500_
	);
	LUT2 #(
		.INIT('h4)
	) name2993 (
		\WX8459_reg/NET0131 ,
		\WX8523_reg/NET0131 ,
		_w4501_
	);
	LUT2 #(
		.INIT('h1)
	) name2994 (
		_w4500_,
		_w4501_,
		_w4502_
	);
	LUT2 #(
		.INIT('h4)
	) name2995 (
		_w4499_,
		_w4502_,
		_w4503_
	);
	LUT2 #(
		.INIT('h2)
	) name2996 (
		_w4499_,
		_w4502_,
		_w4504_
	);
	LUT2 #(
		.INIT('h1)
	) name2997 (
		\TM0_pad ,
		_w4503_,
		_w4505_
	);
	LUT2 #(
		.INIT('h4)
	) name2998 (
		_w4504_,
		_w4505_,
		_w4506_
	);
	LUT2 #(
		.INIT('h2)
	) name2999 (
		_w1976_,
		_w4496_,
		_w4507_
	);
	LUT2 #(
		.INIT('h4)
	) name3000 (
		_w4506_,
		_w4507_,
		_w4508_
	);
	LUT2 #(
		.INIT('h1)
	) name3001 (
		_w4495_,
		_w4508_,
		_w4509_
	);
	LUT2 #(
		.INIT('h4)
	) name3002 (
		_w1508_,
		_w1973_,
		_w4510_
	);
	LUT2 #(
		.INIT('h2)
	) name3003 (
		\WX3421_reg/NET0131 ,
		\WX3485_reg/NET0131 ,
		_w4511_
	);
	LUT2 #(
		.INIT('h4)
	) name3004 (
		\WX3421_reg/NET0131 ,
		\WX3485_reg/NET0131 ,
		_w4512_
	);
	LUT2 #(
		.INIT('h1)
	) name3005 (
		_w4511_,
		_w4512_,
		_w4513_
	);
	LUT2 #(
		.INIT('h2)
	) name3006 (
		\WX3293_reg/NET0131 ,
		\WX3357_reg/NET0131 ,
		_w4514_
	);
	LUT2 #(
		.INIT('h4)
	) name3007 (
		\WX3293_reg/NET0131 ,
		\WX3357_reg/NET0131 ,
		_w4515_
	);
	LUT2 #(
		.INIT('h1)
	) name3008 (
		_w4514_,
		_w4515_,
		_w4516_
	);
	LUT2 #(
		.INIT('h4)
	) name3009 (
		_w4513_,
		_w4516_,
		_w4517_
	);
	LUT2 #(
		.INIT('h2)
	) name3010 (
		_w4513_,
		_w4516_,
		_w4518_
	);
	LUT2 #(
		.INIT('h1)
	) name3011 (
		\TM0_pad ,
		_w4517_,
		_w4519_
	);
	LUT2 #(
		.INIT('h4)
	) name3012 (
		_w4518_,
		_w4519_,
		_w4520_
	);
	LUT2 #(
		.INIT('h2)
	) name3013 (
		_w4510_,
		_w4520_,
		_w4521_
	);
	LUT2 #(
		.INIT('h2)
	) name3014 (
		\TM0_pad ,
		\_2141__reg/NET0131 ,
		_w4522_
	);
	LUT2 #(
		.INIT('h2)
	) name3015 (
		\WX4714_reg/NET0131 ,
		\WX4778_reg/NET0131 ,
		_w4523_
	);
	LUT2 #(
		.INIT('h4)
	) name3016 (
		\WX4714_reg/NET0131 ,
		\WX4778_reg/NET0131 ,
		_w4524_
	);
	LUT2 #(
		.INIT('h1)
	) name3017 (
		_w4523_,
		_w4524_,
		_w4525_
	);
	LUT2 #(
		.INIT('h2)
	) name3018 (
		\WX4586_reg/NET0131 ,
		\WX4650_reg/NET0131 ,
		_w4526_
	);
	LUT2 #(
		.INIT('h4)
	) name3019 (
		\WX4586_reg/NET0131 ,
		\WX4650_reg/NET0131 ,
		_w4527_
	);
	LUT2 #(
		.INIT('h1)
	) name3020 (
		_w4526_,
		_w4527_,
		_w4528_
	);
	LUT2 #(
		.INIT('h4)
	) name3021 (
		_w4525_,
		_w4528_,
		_w4529_
	);
	LUT2 #(
		.INIT('h2)
	) name3022 (
		_w4525_,
		_w4528_,
		_w4530_
	);
	LUT2 #(
		.INIT('h1)
	) name3023 (
		\TM0_pad ,
		_w4529_,
		_w4531_
	);
	LUT2 #(
		.INIT('h4)
	) name3024 (
		_w4530_,
		_w4531_,
		_w4532_
	);
	LUT2 #(
		.INIT('h2)
	) name3025 (
		_w1976_,
		_w4522_,
		_w4533_
	);
	LUT2 #(
		.INIT('h4)
	) name3026 (
		_w4532_,
		_w4533_,
		_w4534_
	);
	LUT2 #(
		.INIT('h1)
	) name3027 (
		_w4521_,
		_w4534_,
		_w4535_
	);
	LUT2 #(
		.INIT('h2)
	) name3028 (
		_w3953_,
		_w4378_,
		_w4536_
	);
	LUT2 #(
		.INIT('h2)
	) name3029 (
		\TM0_pad ,
		\_2273__reg/NET0131 ,
		_w4537_
	);
	LUT2 #(
		.INIT('h2)
	) name3030 (
		\WX9878_reg/NET0131 ,
		\WX9942_reg/NET0131 ,
		_w4538_
	);
	LUT2 #(
		.INIT('h4)
	) name3031 (
		\WX9878_reg/NET0131 ,
		\WX9942_reg/NET0131 ,
		_w4539_
	);
	LUT2 #(
		.INIT('h1)
	) name3032 (
		_w4538_,
		_w4539_,
		_w4540_
	);
	LUT2 #(
		.INIT('h2)
	) name3033 (
		\WX9750_reg/NET0131 ,
		\WX9814_reg/NET0131 ,
		_w4541_
	);
	LUT2 #(
		.INIT('h4)
	) name3034 (
		\WX9750_reg/NET0131 ,
		\WX9814_reg/NET0131 ,
		_w4542_
	);
	LUT2 #(
		.INIT('h1)
	) name3035 (
		_w4541_,
		_w4542_,
		_w4543_
	);
	LUT2 #(
		.INIT('h4)
	) name3036 (
		_w4540_,
		_w4543_,
		_w4544_
	);
	LUT2 #(
		.INIT('h2)
	) name3037 (
		_w4540_,
		_w4543_,
		_w4545_
	);
	LUT2 #(
		.INIT('h1)
	) name3038 (
		\TM0_pad ,
		_w4544_,
		_w4546_
	);
	LUT2 #(
		.INIT('h4)
	) name3039 (
		_w4545_,
		_w4546_,
		_w4547_
	);
	LUT2 #(
		.INIT('h2)
	) name3040 (
		_w1976_,
		_w4537_,
		_w4548_
	);
	LUT2 #(
		.INIT('h4)
	) name3041 (
		_w4547_,
		_w4548_,
		_w4549_
	);
	LUT2 #(
		.INIT('h1)
	) name3042 (
		_w4536_,
		_w4549_,
		_w4550_
	);
	LUT2 #(
		.INIT('h2)
	) name3043 (
		_w3805_,
		_w4419_,
		_w4551_
	);
	LUT2 #(
		.INIT('h2)
	) name3044 (
		\TM0_pad ,
		\_2306__reg/NET0131 ,
		_w4552_
	);
	LUT2 #(
		.INIT('h2)
	) name3045 (
		\WX11169_reg/NET0131 ,
		\WX11233_reg/NET0131 ,
		_w4553_
	);
	LUT2 #(
		.INIT('h4)
	) name3046 (
		\WX11169_reg/NET0131 ,
		\WX11233_reg/NET0131 ,
		_w4554_
	);
	LUT2 #(
		.INIT('h1)
	) name3047 (
		_w4553_,
		_w4554_,
		_w4555_
	);
	LUT2 #(
		.INIT('h2)
	) name3048 (
		\WX11041_reg/NET0131 ,
		\WX11105_reg/NET0131 ,
		_w4556_
	);
	LUT2 #(
		.INIT('h4)
	) name3049 (
		\WX11041_reg/NET0131 ,
		\WX11105_reg/NET0131 ,
		_w4557_
	);
	LUT2 #(
		.INIT('h1)
	) name3050 (
		_w4556_,
		_w4557_,
		_w4558_
	);
	LUT2 #(
		.INIT('h4)
	) name3051 (
		_w4555_,
		_w4558_,
		_w4559_
	);
	LUT2 #(
		.INIT('h2)
	) name3052 (
		_w4555_,
		_w4558_,
		_w4560_
	);
	LUT2 #(
		.INIT('h1)
	) name3053 (
		\TM0_pad ,
		_w4559_,
		_w4561_
	);
	LUT2 #(
		.INIT('h4)
	) name3054 (
		_w4560_,
		_w4561_,
		_w4562_
	);
	LUT2 #(
		.INIT('h2)
	) name3055 (
		_w1976_,
		_w4552_,
		_w4563_
	);
	LUT2 #(
		.INIT('h4)
	) name3056 (
		_w4562_,
		_w4563_,
		_w4564_
	);
	LUT2 #(
		.INIT('h1)
	) name3057 (
		_w4551_,
		_w4564_,
		_w4565_
	);
	LUT2 #(
		.INIT('h2)
	) name3058 (
		_w4382_,
		_w4404_,
		_w4566_
	);
	LUT2 #(
		.INIT('h2)
	) name3059 (
		\TM0_pad ,
		\_2174__reg/NET0131 ,
		_w4567_
	);
	LUT2 #(
		.INIT('h2)
	) name3060 (
		\WX6005_reg/NET0131 ,
		\WX6069_reg/NET0131 ,
		_w4568_
	);
	LUT2 #(
		.INIT('h4)
	) name3061 (
		\WX6005_reg/NET0131 ,
		\WX6069_reg/NET0131 ,
		_w4569_
	);
	LUT2 #(
		.INIT('h1)
	) name3062 (
		_w4568_,
		_w4569_,
		_w4570_
	);
	LUT2 #(
		.INIT('h2)
	) name3063 (
		\WX5877_reg/NET0131 ,
		\WX5941_reg/NET0131 ,
		_w4571_
	);
	LUT2 #(
		.INIT('h4)
	) name3064 (
		\WX5877_reg/NET0131 ,
		\WX5941_reg/NET0131 ,
		_w4572_
	);
	LUT2 #(
		.INIT('h1)
	) name3065 (
		_w4571_,
		_w4572_,
		_w4573_
	);
	LUT2 #(
		.INIT('h4)
	) name3066 (
		_w4570_,
		_w4573_,
		_w4574_
	);
	LUT2 #(
		.INIT('h2)
	) name3067 (
		_w4570_,
		_w4573_,
		_w4575_
	);
	LUT2 #(
		.INIT('h1)
	) name3068 (
		\TM0_pad ,
		_w4574_,
		_w4576_
	);
	LUT2 #(
		.INIT('h4)
	) name3069 (
		_w4575_,
		_w4576_,
		_w4577_
	);
	LUT2 #(
		.INIT('h2)
	) name3070 (
		_w1976_,
		_w4567_,
		_w4578_
	);
	LUT2 #(
		.INIT('h4)
	) name3071 (
		_w4577_,
		_w4578_,
		_w4579_
	);
	LUT2 #(
		.INIT('h1)
	) name3072 (
		_w4566_,
		_w4579_,
		_w4580_
	);
	LUT2 #(
		.INIT('h2)
	) name3073 (
		_w1974_,
		_w1987_,
		_w4581_
	);
	LUT2 #(
		.INIT('h2)
	) name3074 (
		\TM0_pad ,
		\_2124__reg/NET0131 ,
		_w4582_
	);
	LUT2 #(
		.INIT('h2)
	) name3075 (
		_w1976_,
		_w4582_,
		_w4583_
	);
	LUT2 #(
		.INIT('h4)
	) name3076 (
		_w2106_,
		_w4583_,
		_w4584_
	);
	LUT2 #(
		.INIT('h1)
	) name3077 (
		_w4581_,
		_w4584_,
		_w4585_
	);
	LUT2 #(
		.INIT('h2)
	) name3078 (
		_w4239_,
		_w4449_,
		_w4586_
	);
	LUT2 #(
		.INIT('h2)
	) name3079 (
		\TM0_pad ,
		\_2207__reg/NET0131 ,
		_w4587_
	);
	LUT2 #(
		.INIT('h2)
	) name3080 (
		\WX7296_reg/NET0131 ,
		\WX7360_reg/NET0131 ,
		_w4588_
	);
	LUT2 #(
		.INIT('h4)
	) name3081 (
		\WX7296_reg/NET0131 ,
		\WX7360_reg/NET0131 ,
		_w4589_
	);
	LUT2 #(
		.INIT('h1)
	) name3082 (
		_w4588_,
		_w4589_,
		_w4590_
	);
	LUT2 #(
		.INIT('h2)
	) name3083 (
		\WX7168_reg/NET0131 ,
		\WX7232_reg/NET0131 ,
		_w4591_
	);
	LUT2 #(
		.INIT('h4)
	) name3084 (
		\WX7168_reg/NET0131 ,
		\WX7232_reg/NET0131 ,
		_w4592_
	);
	LUT2 #(
		.INIT('h1)
	) name3085 (
		_w4591_,
		_w4592_,
		_w4593_
	);
	LUT2 #(
		.INIT('h4)
	) name3086 (
		_w4590_,
		_w4593_,
		_w4594_
	);
	LUT2 #(
		.INIT('h2)
	) name3087 (
		_w4590_,
		_w4593_,
		_w4595_
	);
	LUT2 #(
		.INIT('h1)
	) name3088 (
		\TM0_pad ,
		_w4594_,
		_w4596_
	);
	LUT2 #(
		.INIT('h4)
	) name3089 (
		_w4595_,
		_w4596_,
		_w4597_
	);
	LUT2 #(
		.INIT('h2)
	) name3090 (
		_w1976_,
		_w4587_,
		_w4598_
	);
	LUT2 #(
		.INIT('h4)
	) name3091 (
		_w4597_,
		_w4598_,
		_w4599_
	);
	LUT2 #(
		.INIT('h1)
	) name3092 (
		_w4586_,
		_w4599_,
		_w4600_
	);
	LUT2 #(
		.INIT('h1)
	) name3093 (
		\TM0_pad ,
		_w1569_,
		_w4601_
	);
	LUT2 #(
		.INIT('h2)
	) name3094 (
		_w2040_,
		_w4601_,
		_w4602_
	);
	LUT2 #(
		.INIT('h2)
	) name3095 (
		\TM0_pad ,
		\_2090__reg/NET0131 ,
		_w4603_
	);
	LUT2 #(
		.INIT('h2)
	) name3096 (
		\WX2102_reg/NET0131 ,
		\WX2166_reg/NET0131 ,
		_w4604_
	);
	LUT2 #(
		.INIT('h4)
	) name3097 (
		\WX2102_reg/NET0131 ,
		\WX2166_reg/NET0131 ,
		_w4605_
	);
	LUT2 #(
		.INIT('h1)
	) name3098 (
		_w4604_,
		_w4605_,
		_w4606_
	);
	LUT2 #(
		.INIT('h2)
	) name3099 (
		\WX1974_reg/NET0131 ,
		\WX2038_reg/NET0131 ,
		_w4607_
	);
	LUT2 #(
		.INIT('h4)
	) name3100 (
		\WX1974_reg/NET0131 ,
		\WX2038_reg/NET0131 ,
		_w4608_
	);
	LUT2 #(
		.INIT('h1)
	) name3101 (
		_w4607_,
		_w4608_,
		_w4609_
	);
	LUT2 #(
		.INIT('h4)
	) name3102 (
		_w4606_,
		_w4609_,
		_w4610_
	);
	LUT2 #(
		.INIT('h2)
	) name3103 (
		_w4606_,
		_w4609_,
		_w4611_
	);
	LUT2 #(
		.INIT('h1)
	) name3104 (
		\TM0_pad ,
		_w4610_,
		_w4612_
	);
	LUT2 #(
		.INIT('h4)
	) name3105 (
		_w4611_,
		_w4612_,
		_w4613_
	);
	LUT2 #(
		.INIT('h2)
	) name3106 (
		_w1976_,
		_w4603_,
		_w4614_
	);
	LUT2 #(
		.INIT('h4)
	) name3107 (
		_w4613_,
		_w4614_,
		_w4615_
	);
	LUT2 #(
		.INIT('h1)
	) name3108 (
		_w4602_,
		_w4615_,
		_w4616_
	);
	LUT2 #(
		.INIT('h8)
	) name3109 (
		RESET_pad,
		\WX10859_reg/NET0131 ,
		_w4617_
	);
	LUT2 #(
		.INIT('h2)
	) name3110 (
		_w4239_,
		_w4597_,
		_w4618_
	);
	LUT2 #(
		.INIT('h2)
	) name3111 (
		\TM0_pad ,
		\_2239__reg/NET0131 ,
		_w4619_
	);
	LUT2 #(
		.INIT('h2)
	) name3112 (
		\WX8589_reg/NET0131 ,
		\WX8653_reg/NET0131 ,
		_w4620_
	);
	LUT2 #(
		.INIT('h4)
	) name3113 (
		\WX8589_reg/NET0131 ,
		\WX8653_reg/NET0131 ,
		_w4621_
	);
	LUT2 #(
		.INIT('h1)
	) name3114 (
		_w4620_,
		_w4621_,
		_w4622_
	);
	LUT2 #(
		.INIT('h2)
	) name3115 (
		\WX8461_reg/NET0131 ,
		\WX8525_reg/NET0131 ,
		_w4623_
	);
	LUT2 #(
		.INIT('h4)
	) name3116 (
		\WX8461_reg/NET0131 ,
		\WX8525_reg/NET0131 ,
		_w4624_
	);
	LUT2 #(
		.INIT('h1)
	) name3117 (
		_w4623_,
		_w4624_,
		_w4625_
	);
	LUT2 #(
		.INIT('h4)
	) name3118 (
		_w4622_,
		_w4625_,
		_w4626_
	);
	LUT2 #(
		.INIT('h2)
	) name3119 (
		_w4622_,
		_w4625_,
		_w4627_
	);
	LUT2 #(
		.INIT('h1)
	) name3120 (
		\TM0_pad ,
		_w4626_,
		_w4628_
	);
	LUT2 #(
		.INIT('h4)
	) name3121 (
		_w4627_,
		_w4628_,
		_w4629_
	);
	LUT2 #(
		.INIT('h2)
	) name3122 (
		_w1976_,
		_w4619_,
		_w4630_
	);
	LUT2 #(
		.INIT('h4)
	) name3123 (
		_w4629_,
		_w4630_,
		_w4631_
	);
	LUT2 #(
		.INIT('h1)
	) name3124 (
		_w4618_,
		_w4631_,
		_w4632_
	);
	LUT2 #(
		.INIT('h2)
	) name3125 (
		_w4101_,
		_w4506_,
		_w4633_
	);
	LUT2 #(
		.INIT('h2)
	) name3126 (
		\TM0_pad ,
		\_2272__reg/NET0131 ,
		_w4634_
	);
	LUT2 #(
		.INIT('h2)
	) name3127 (
		\WX9880_reg/NET0131 ,
		\WX9944_reg/NET0131 ,
		_w4635_
	);
	LUT2 #(
		.INIT('h4)
	) name3128 (
		\WX9880_reg/NET0131 ,
		\WX9944_reg/NET0131 ,
		_w4636_
	);
	LUT2 #(
		.INIT('h1)
	) name3129 (
		_w4635_,
		_w4636_,
		_w4637_
	);
	LUT2 #(
		.INIT('h2)
	) name3130 (
		\WX9752_reg/NET0131 ,
		\WX9816_reg/NET0131 ,
		_w4638_
	);
	LUT2 #(
		.INIT('h4)
	) name3131 (
		\WX9752_reg/NET0131 ,
		\WX9816_reg/NET0131 ,
		_w4639_
	);
	LUT2 #(
		.INIT('h1)
	) name3132 (
		_w4638_,
		_w4639_,
		_w4640_
	);
	LUT2 #(
		.INIT('h4)
	) name3133 (
		_w4637_,
		_w4640_,
		_w4641_
	);
	LUT2 #(
		.INIT('h2)
	) name3134 (
		_w4637_,
		_w4640_,
		_w4642_
	);
	LUT2 #(
		.INIT('h1)
	) name3135 (
		\TM0_pad ,
		_w4641_,
		_w4643_
	);
	LUT2 #(
		.INIT('h4)
	) name3136 (
		_w4642_,
		_w4643_,
		_w4644_
	);
	LUT2 #(
		.INIT('h2)
	) name3137 (
		_w1976_,
		_w4634_,
		_w4645_
	);
	LUT2 #(
		.INIT('h4)
	) name3138 (
		_w4644_,
		_w4645_,
		_w4646_
	);
	LUT2 #(
		.INIT('h1)
	) name3139 (
		_w4633_,
		_w4646_,
		_w4647_
	);
	LUT2 #(
		.INIT('h2)
	) name3140 (
		_w3953_,
		_w4547_,
		_w4648_
	);
	LUT2 #(
		.INIT('h2)
	) name3141 (
		\TM0_pad ,
		\_2305__reg/NET0131 ,
		_w4649_
	);
	LUT2 #(
		.INIT('h2)
	) name3142 (
		\WX11171_reg/NET0131 ,
		\WX11235_reg/NET0131 ,
		_w4650_
	);
	LUT2 #(
		.INIT('h4)
	) name3143 (
		\WX11171_reg/NET0131 ,
		\WX11235_reg/NET0131 ,
		_w4651_
	);
	LUT2 #(
		.INIT('h1)
	) name3144 (
		_w4650_,
		_w4651_,
		_w4652_
	);
	LUT2 #(
		.INIT('h2)
	) name3145 (
		\WX11043_reg/NET0131 ,
		\WX11107_reg/NET0131 ,
		_w4653_
	);
	LUT2 #(
		.INIT('h4)
	) name3146 (
		\WX11043_reg/NET0131 ,
		\WX11107_reg/NET0131 ,
		_w4654_
	);
	LUT2 #(
		.INIT('h1)
	) name3147 (
		_w4653_,
		_w4654_,
		_w4655_
	);
	LUT2 #(
		.INIT('h4)
	) name3148 (
		_w4652_,
		_w4655_,
		_w4656_
	);
	LUT2 #(
		.INIT('h2)
	) name3149 (
		_w4652_,
		_w4655_,
		_w4657_
	);
	LUT2 #(
		.INIT('h1)
	) name3150 (
		\TM0_pad ,
		_w4656_,
		_w4658_
	);
	LUT2 #(
		.INIT('h4)
	) name3151 (
		_w4657_,
		_w4658_,
		_w4659_
	);
	LUT2 #(
		.INIT('h2)
	) name3152 (
		_w1976_,
		_w4649_,
		_w4660_
	);
	LUT2 #(
		.INIT('h4)
	) name3153 (
		_w4659_,
		_w4660_,
		_w4661_
	);
	LUT2 #(
		.INIT('h1)
	) name3154 (
		_w4648_,
		_w4661_,
		_w4662_
	);
	LUT2 #(
		.INIT('h2)
	) name3155 (
		_w4510_,
		_w4532_,
		_w4663_
	);
	LUT2 #(
		.INIT('h2)
	) name3156 (
		\TM0_pad ,
		\_2173__reg/NET0131 ,
		_w4664_
	);
	LUT2 #(
		.INIT('h2)
	) name3157 (
		\WX6007_reg/NET0131 ,
		\WX6071_reg/NET0131 ,
		_w4665_
	);
	LUT2 #(
		.INIT('h4)
	) name3158 (
		\WX6007_reg/NET0131 ,
		\WX6071_reg/NET0131 ,
		_w4666_
	);
	LUT2 #(
		.INIT('h1)
	) name3159 (
		_w4665_,
		_w4666_,
		_w4667_
	);
	LUT2 #(
		.INIT('h2)
	) name3160 (
		\WX5879_reg/NET0131 ,
		\WX5943_reg/NET0131 ,
		_w4668_
	);
	LUT2 #(
		.INIT('h4)
	) name3161 (
		\WX5879_reg/NET0131 ,
		\WX5943_reg/NET0131 ,
		_w4669_
	);
	LUT2 #(
		.INIT('h1)
	) name3162 (
		_w4668_,
		_w4669_,
		_w4670_
	);
	LUT2 #(
		.INIT('h4)
	) name3163 (
		_w4667_,
		_w4670_,
		_w4671_
	);
	LUT2 #(
		.INIT('h2)
	) name3164 (
		_w4667_,
		_w4670_,
		_w4672_
	);
	LUT2 #(
		.INIT('h1)
	) name3165 (
		\TM0_pad ,
		_w4671_,
		_w4673_
	);
	LUT2 #(
		.INIT('h4)
	) name3166 (
		_w4672_,
		_w4673_,
		_w4674_
	);
	LUT2 #(
		.INIT('h2)
	) name3167 (
		_w1976_,
		_w4664_,
		_w4675_
	);
	LUT2 #(
		.INIT('h4)
	) name3168 (
		_w4674_,
		_w4675_,
		_w4676_
	);
	LUT2 #(
		.INIT('h1)
	) name3169 (
		_w4663_,
		_w4676_,
		_w4677_
	);
	LUT2 #(
		.INIT('h2)
	) name3170 (
		\WX2100_reg/NET0131 ,
		\WX2164_reg/NET0131 ,
		_w4678_
	);
	LUT2 #(
		.INIT('h4)
	) name3171 (
		\WX2100_reg/NET0131 ,
		\WX2164_reg/NET0131 ,
		_w4679_
	);
	LUT2 #(
		.INIT('h1)
	) name3172 (
		_w4678_,
		_w4679_,
		_w4680_
	);
	LUT2 #(
		.INIT('h2)
	) name3173 (
		\WX1972_reg/NET0131 ,
		\WX2036_reg/NET0131 ,
		_w4681_
	);
	LUT2 #(
		.INIT('h4)
	) name3174 (
		\WX1972_reg/NET0131 ,
		\WX2036_reg/NET0131 ,
		_w4682_
	);
	LUT2 #(
		.INIT('h1)
	) name3175 (
		_w4681_,
		_w4682_,
		_w4683_
	);
	LUT2 #(
		.INIT('h4)
	) name3176 (
		_w4680_,
		_w4683_,
		_w4684_
	);
	LUT2 #(
		.INIT('h2)
	) name3177 (
		_w4680_,
		_w4683_,
		_w4685_
	);
	LUT2 #(
		.INIT('h1)
	) name3178 (
		\TM0_pad ,
		_w4684_,
		_w4686_
	);
	LUT2 #(
		.INIT('h4)
	) name3179 (
		_w4685_,
		_w4686_,
		_w4687_
	);
	LUT2 #(
		.INIT('h2)
	) name3180 (
		_w2341_,
		_w4687_,
		_w4688_
	);
	LUT2 #(
		.INIT('h2)
	) name3181 (
		\TM0_pad ,
		\_2123__reg/NET0131 ,
		_w4689_
	);
	LUT2 #(
		.INIT('h2)
	) name3182 (
		_w1976_,
		_w4689_,
		_w4690_
	);
	LUT2 #(
		.INIT('h4)
	) name3183 (
		_w2351_,
		_w4690_,
		_w4691_
	);
	LUT2 #(
		.INIT('h1)
	) name3184 (
		_w4688_,
		_w4691_,
		_w4692_
	);
	LUT2 #(
		.INIT('h2)
	) name3185 (
		_w4382_,
		_w4577_,
		_w4693_
	);
	LUT2 #(
		.INIT('h2)
	) name3186 (
		\TM0_pad ,
		\_2206__reg/NET0131 ,
		_w4694_
	);
	LUT2 #(
		.INIT('h2)
	) name3187 (
		\WX7298_reg/NET0131 ,
		\WX7362_reg/NET0131 ,
		_w4695_
	);
	LUT2 #(
		.INIT('h4)
	) name3188 (
		\WX7298_reg/NET0131 ,
		\WX7362_reg/NET0131 ,
		_w4696_
	);
	LUT2 #(
		.INIT('h1)
	) name3189 (
		_w4695_,
		_w4696_,
		_w4697_
	);
	LUT2 #(
		.INIT('h2)
	) name3190 (
		\WX7170_reg/NET0131 ,
		\WX7234_reg/NET0131 ,
		_w4698_
	);
	LUT2 #(
		.INIT('h4)
	) name3191 (
		\WX7170_reg/NET0131 ,
		\WX7234_reg/NET0131 ,
		_w4699_
	);
	LUT2 #(
		.INIT('h1)
	) name3192 (
		_w4698_,
		_w4699_,
		_w4700_
	);
	LUT2 #(
		.INIT('h4)
	) name3193 (
		_w4697_,
		_w4700_,
		_w4701_
	);
	LUT2 #(
		.INIT('h2)
	) name3194 (
		_w4697_,
		_w4700_,
		_w4702_
	);
	LUT2 #(
		.INIT('h1)
	) name3195 (
		\TM0_pad ,
		_w4701_,
		_w4703_
	);
	LUT2 #(
		.INIT('h4)
	) name3196 (
		_w4702_,
		_w4703_,
		_w4704_
	);
	LUT2 #(
		.INIT('h2)
	) name3197 (
		_w1976_,
		_w4694_,
		_w4705_
	);
	LUT2 #(
		.INIT('h4)
	) name3198 (
		_w4704_,
		_w4705_,
		_w4706_
	);
	LUT2 #(
		.INIT('h1)
	) name3199 (
		_w4693_,
		_w4706_,
		_w4707_
	);
	LUT2 #(
		.INIT('h8)
	) name3200 (
		\TM0_pad ,
		\_2172__reg/NET0131 ,
		_w4708_
	);
	LUT2 #(
		.INIT('h2)
	) name3201 (
		\WX4652_reg/NET0131 ,
		\WX4716_reg/NET0131 ,
		_w4709_
	);
	LUT2 #(
		.INIT('h4)
	) name3202 (
		\WX4652_reg/NET0131 ,
		\WX4716_reg/NET0131 ,
		_w4710_
	);
	LUT2 #(
		.INIT('h1)
	) name3203 (
		_w4709_,
		_w4710_,
		_w4711_
	);
	LUT2 #(
		.INIT('h2)
	) name3204 (
		\WX4588_reg/NET0131 ,
		_w4711_,
		_w4712_
	);
	LUT2 #(
		.INIT('h4)
	) name3205 (
		\WX4588_reg/NET0131 ,
		_w4711_,
		_w4713_
	);
	LUT2 #(
		.INIT('h1)
	) name3206 (
		_w4712_,
		_w4713_,
		_w4714_
	);
	LUT2 #(
		.INIT('h2)
	) name3207 (
		\TM1_pad ,
		\WX4524_reg/NET0131 ,
		_w4715_
	);
	LUT2 #(
		.INIT('h4)
	) name3208 (
		\TM1_pad ,
		\WX4524_reg/NET0131 ,
		_w4716_
	);
	LUT2 #(
		.INIT('h1)
	) name3209 (
		_w4715_,
		_w4716_,
		_w4717_
	);
	LUT2 #(
		.INIT('h4)
	) name3210 (
		_w4714_,
		_w4717_,
		_w4718_
	);
	LUT2 #(
		.INIT('h2)
	) name3211 (
		_w4714_,
		_w4717_,
		_w4719_
	);
	LUT2 #(
		.INIT('h1)
	) name3212 (
		\TM0_pad ,
		_w4718_,
		_w4720_
	);
	LUT2 #(
		.INIT('h4)
	) name3213 (
		_w4719_,
		_w4720_,
		_w4721_
	);
	LUT2 #(
		.INIT('h1)
	) name3214 (
		_w4708_,
		_w4721_,
		_w4722_
	);
	LUT2 #(
		.INIT('h2)
	) name3215 (
		_w1976_,
		_w4722_,
		_w4723_
	);
	LUT2 #(
		.INIT('h2)
	) name3216 (
		\WX3359_reg/NET0131 ,
		\WX3423_reg/NET0131 ,
		_w4724_
	);
	LUT2 #(
		.INIT('h4)
	) name3217 (
		\WX3359_reg/NET0131 ,
		\WX3423_reg/NET0131 ,
		_w4725_
	);
	LUT2 #(
		.INIT('h1)
	) name3218 (
		_w4724_,
		_w4725_,
		_w4726_
	);
	LUT2 #(
		.INIT('h2)
	) name3219 (
		\WX3295_reg/NET0131 ,
		_w4726_,
		_w4727_
	);
	LUT2 #(
		.INIT('h4)
	) name3220 (
		\WX3295_reg/NET0131 ,
		_w4726_,
		_w4728_
	);
	LUT2 #(
		.INIT('h1)
	) name3221 (
		_w4727_,
		_w4728_,
		_w4729_
	);
	LUT2 #(
		.INIT('h2)
	) name3222 (
		\TM1_pad ,
		\WX3231_reg/NET0131 ,
		_w4730_
	);
	LUT2 #(
		.INIT('h4)
	) name3223 (
		\TM1_pad ,
		\WX3231_reg/NET0131 ,
		_w4731_
	);
	LUT2 #(
		.INIT('h1)
	) name3224 (
		_w4730_,
		_w4731_,
		_w4732_
	);
	LUT2 #(
		.INIT('h4)
	) name3225 (
		_w4729_,
		_w4732_,
		_w4733_
	);
	LUT2 #(
		.INIT('h2)
	) name3226 (
		_w4729_,
		_w4732_,
		_w4734_
	);
	LUT2 #(
		.INIT('h1)
	) name3227 (
		\TM0_pad ,
		_w4733_,
		_w4735_
	);
	LUT2 #(
		.INIT('h4)
	) name3228 (
		_w4734_,
		_w4735_,
		_w4736_
	);
	LUT2 #(
		.INIT('h1)
	) name3229 (
		_w1871_,
		_w4736_,
		_w4737_
	);
	LUT2 #(
		.INIT('h2)
	) name3230 (
		_w1973_,
		_w4737_,
		_w4738_
	);
	LUT2 #(
		.INIT('h1)
	) name3231 (
		_w4723_,
		_w4738_,
		_w4739_
	);
	LUT2 #(
		.INIT('h1)
	) name3232 (
		\TM0_pad ,
		_w1556_,
		_w4740_
	);
	LUT2 #(
		.INIT('h2)
	) name3233 (
		_w2677_,
		_w4740_,
		_w4741_
	);
	LUT2 #(
		.INIT('h2)
	) name3234 (
		\TM0_pad ,
		\_2089__reg/NET0131 ,
		_w4742_
	);
	LUT2 #(
		.INIT('h2)
	) name3235 (
		\WX2104_reg/NET0131 ,
		\WX2168_reg/NET0131 ,
		_w4743_
	);
	LUT2 #(
		.INIT('h4)
	) name3236 (
		\WX2104_reg/NET0131 ,
		\WX2168_reg/NET0131 ,
		_w4744_
	);
	LUT2 #(
		.INIT('h1)
	) name3237 (
		_w4743_,
		_w4744_,
		_w4745_
	);
	LUT2 #(
		.INIT('h2)
	) name3238 (
		\WX1976_reg/NET0131 ,
		\WX2040_reg/NET0131 ,
		_w4746_
	);
	LUT2 #(
		.INIT('h4)
	) name3239 (
		\WX1976_reg/NET0131 ,
		\WX2040_reg/NET0131 ,
		_w4747_
	);
	LUT2 #(
		.INIT('h1)
	) name3240 (
		_w4746_,
		_w4747_,
		_w4748_
	);
	LUT2 #(
		.INIT('h4)
	) name3241 (
		_w4745_,
		_w4748_,
		_w4749_
	);
	LUT2 #(
		.INIT('h2)
	) name3242 (
		_w4745_,
		_w4748_,
		_w4750_
	);
	LUT2 #(
		.INIT('h1)
	) name3243 (
		\TM0_pad ,
		_w4749_,
		_w4751_
	);
	LUT2 #(
		.INIT('h4)
	) name3244 (
		_w4750_,
		_w4751_,
		_w4752_
	);
	LUT2 #(
		.INIT('h2)
	) name3245 (
		_w1976_,
		_w4742_,
		_w4753_
	);
	LUT2 #(
		.INIT('h4)
	) name3246 (
		_w4752_,
		_w4753_,
		_w4754_
	);
	LUT2 #(
		.INIT('h1)
	) name3247 (
		_w4741_,
		_w4754_,
		_w4755_
	);
	LUT2 #(
		.INIT('h2)
	) name3248 (
		_w2341_,
		_w3224_,
		_w4756_
	);
	LUT2 #(
		.INIT('h1)
	) name3249 (
		\DATA_0_14_pad ,
		\TM0_pad ,
		_w4757_
	);
	LUT2 #(
		.INIT('h2)
	) name3250 (
		\TM0_pad ,
		\_2347__reg/NET0131 ,
		_w4758_
	);
	LUT2 #(
		.INIT('h2)
	) name3251 (
		_w1976_,
		_w4757_,
		_w4759_
	);
	LUT2 #(
		.INIT('h4)
	) name3252 (
		_w4758_,
		_w4759_,
		_w4760_
	);
	LUT2 #(
		.INIT('h1)
	) name3253 (
		_w4756_,
		_w4760_,
		_w4761_
	);
	LUT2 #(
		.INIT('h8)
	) name3254 (
		RESET_pad,
		\WX10861_reg/NET0131 ,
		_w4762_
	);
	LUT2 #(
		.INIT('h2)
	) name3255 (
		_w4382_,
		_w4704_,
		_w4763_
	);
	LUT2 #(
		.INIT('h2)
	) name3256 (
		\TM0_pad ,
		\_2238__reg/NET0131 ,
		_w4764_
	);
	LUT2 #(
		.INIT('h2)
	) name3257 (
		\WX8591_reg/NET0131 ,
		\WX8655_reg/NET0131 ,
		_w4765_
	);
	LUT2 #(
		.INIT('h4)
	) name3258 (
		\WX8591_reg/NET0131 ,
		\WX8655_reg/NET0131 ,
		_w4766_
	);
	LUT2 #(
		.INIT('h1)
	) name3259 (
		_w4765_,
		_w4766_,
		_w4767_
	);
	LUT2 #(
		.INIT('h2)
	) name3260 (
		\WX8463_reg/NET0131 ,
		\WX8527_reg/NET0131 ,
		_w4768_
	);
	LUT2 #(
		.INIT('h4)
	) name3261 (
		\WX8463_reg/NET0131 ,
		\WX8527_reg/NET0131 ,
		_w4769_
	);
	LUT2 #(
		.INIT('h1)
	) name3262 (
		_w4768_,
		_w4769_,
		_w4770_
	);
	LUT2 #(
		.INIT('h4)
	) name3263 (
		_w4767_,
		_w4770_,
		_w4771_
	);
	LUT2 #(
		.INIT('h2)
	) name3264 (
		_w4767_,
		_w4770_,
		_w4772_
	);
	LUT2 #(
		.INIT('h1)
	) name3265 (
		\TM0_pad ,
		_w4771_,
		_w4773_
	);
	LUT2 #(
		.INIT('h4)
	) name3266 (
		_w4772_,
		_w4773_,
		_w4774_
	);
	LUT2 #(
		.INIT('h2)
	) name3267 (
		_w1976_,
		_w4764_,
		_w4775_
	);
	LUT2 #(
		.INIT('h4)
	) name3268 (
		_w4774_,
		_w4775_,
		_w4776_
	);
	LUT2 #(
		.INIT('h1)
	) name3269 (
		_w4763_,
		_w4776_,
		_w4777_
	);
	LUT2 #(
		.INIT('h2)
	) name3270 (
		_w4239_,
		_w4629_,
		_w4778_
	);
	LUT2 #(
		.INIT('h2)
	) name3271 (
		\TM0_pad ,
		\_2271__reg/NET0131 ,
		_w4779_
	);
	LUT2 #(
		.INIT('h2)
	) name3272 (
		\WX9882_reg/NET0131 ,
		\WX9946_reg/NET0131 ,
		_w4780_
	);
	LUT2 #(
		.INIT('h4)
	) name3273 (
		\WX9882_reg/NET0131 ,
		\WX9946_reg/NET0131 ,
		_w4781_
	);
	LUT2 #(
		.INIT('h1)
	) name3274 (
		_w4780_,
		_w4781_,
		_w4782_
	);
	LUT2 #(
		.INIT('h2)
	) name3275 (
		\WX9754_reg/NET0131 ,
		\WX9818_reg/NET0131 ,
		_w4783_
	);
	LUT2 #(
		.INIT('h4)
	) name3276 (
		\WX9754_reg/NET0131 ,
		\WX9818_reg/NET0131 ,
		_w4784_
	);
	LUT2 #(
		.INIT('h1)
	) name3277 (
		_w4783_,
		_w4784_,
		_w4785_
	);
	LUT2 #(
		.INIT('h4)
	) name3278 (
		_w4782_,
		_w4785_,
		_w4786_
	);
	LUT2 #(
		.INIT('h2)
	) name3279 (
		_w4782_,
		_w4785_,
		_w4787_
	);
	LUT2 #(
		.INIT('h1)
	) name3280 (
		\TM0_pad ,
		_w4786_,
		_w4788_
	);
	LUT2 #(
		.INIT('h4)
	) name3281 (
		_w4787_,
		_w4788_,
		_w4789_
	);
	LUT2 #(
		.INIT('h2)
	) name3282 (
		_w1976_,
		_w4779_,
		_w4790_
	);
	LUT2 #(
		.INIT('h4)
	) name3283 (
		_w4789_,
		_w4790_,
		_w4791_
	);
	LUT2 #(
		.INIT('h1)
	) name3284 (
		_w4778_,
		_w4791_,
		_w4792_
	);
	LUT2 #(
		.INIT('h8)
	) name3285 (
		\TM0_pad ,
		\_2204__reg/NET0131 ,
		_w4793_
	);
	LUT2 #(
		.INIT('h2)
	) name3286 (
		\WX5945_reg/NET0131 ,
		\WX6009_reg/NET0131 ,
		_w4794_
	);
	LUT2 #(
		.INIT('h4)
	) name3287 (
		\WX5945_reg/NET0131 ,
		\WX6009_reg/NET0131 ,
		_w4795_
	);
	LUT2 #(
		.INIT('h1)
	) name3288 (
		_w4794_,
		_w4795_,
		_w4796_
	);
	LUT2 #(
		.INIT('h2)
	) name3289 (
		\WX5881_reg/NET0131 ,
		_w4796_,
		_w4797_
	);
	LUT2 #(
		.INIT('h4)
	) name3290 (
		\WX5881_reg/NET0131 ,
		_w4796_,
		_w4798_
	);
	LUT2 #(
		.INIT('h1)
	) name3291 (
		_w4797_,
		_w4798_,
		_w4799_
	);
	LUT2 #(
		.INIT('h2)
	) name3292 (
		\TM1_pad ,
		\WX5817_reg/NET0131 ,
		_w4800_
	);
	LUT2 #(
		.INIT('h4)
	) name3293 (
		\TM1_pad ,
		\WX5817_reg/NET0131 ,
		_w4801_
	);
	LUT2 #(
		.INIT('h1)
	) name3294 (
		_w4800_,
		_w4801_,
		_w4802_
	);
	LUT2 #(
		.INIT('h4)
	) name3295 (
		_w4799_,
		_w4802_,
		_w4803_
	);
	LUT2 #(
		.INIT('h2)
	) name3296 (
		_w4799_,
		_w4802_,
		_w4804_
	);
	LUT2 #(
		.INIT('h1)
	) name3297 (
		\TM0_pad ,
		_w4803_,
		_w4805_
	);
	LUT2 #(
		.INIT('h4)
	) name3298 (
		_w4804_,
		_w4805_,
		_w4806_
	);
	LUT2 #(
		.INIT('h1)
	) name3299 (
		_w4793_,
		_w4806_,
		_w4807_
	);
	LUT2 #(
		.INIT('h2)
	) name3300 (
		_w1976_,
		_w4807_,
		_w4808_
	);
	LUT2 #(
		.INIT('h1)
	) name3301 (
		_w1871_,
		_w4721_,
		_w4809_
	);
	LUT2 #(
		.INIT('h2)
	) name3302 (
		_w1973_,
		_w4809_,
		_w4810_
	);
	LUT2 #(
		.INIT('h1)
	) name3303 (
		_w4808_,
		_w4810_,
		_w4811_
	);
	LUT2 #(
		.INIT('h2)
	) name3304 (
		_w4101_,
		_w4644_,
		_w4812_
	);
	LUT2 #(
		.INIT('h2)
	) name3305 (
		\TM0_pad ,
		\_2304__reg/NET0131 ,
		_w4813_
	);
	LUT2 #(
		.INIT('h2)
	) name3306 (
		\WX11173_reg/NET0131 ,
		\WX11237_reg/NET0131 ,
		_w4814_
	);
	LUT2 #(
		.INIT('h4)
	) name3307 (
		\WX11173_reg/NET0131 ,
		\WX11237_reg/NET0131 ,
		_w4815_
	);
	LUT2 #(
		.INIT('h1)
	) name3308 (
		_w4814_,
		_w4815_,
		_w4816_
	);
	LUT2 #(
		.INIT('h2)
	) name3309 (
		\WX11045_reg/NET0131 ,
		\WX11109_reg/NET0131 ,
		_w4817_
	);
	LUT2 #(
		.INIT('h4)
	) name3310 (
		\WX11045_reg/NET0131 ,
		\WX11109_reg/NET0131 ,
		_w4818_
	);
	LUT2 #(
		.INIT('h1)
	) name3311 (
		_w4817_,
		_w4818_,
		_w4819_
	);
	LUT2 #(
		.INIT('h4)
	) name3312 (
		_w4816_,
		_w4819_,
		_w4820_
	);
	LUT2 #(
		.INIT('h2)
	) name3313 (
		_w4816_,
		_w4819_,
		_w4821_
	);
	LUT2 #(
		.INIT('h1)
	) name3314 (
		\TM0_pad ,
		_w4820_,
		_w4822_
	);
	LUT2 #(
		.INIT('h4)
	) name3315 (
		_w4821_,
		_w4822_,
		_w4823_
	);
	LUT2 #(
		.INIT('h2)
	) name3316 (
		_w1976_,
		_w4813_,
		_w4824_
	);
	LUT2 #(
		.INIT('h4)
	) name3317 (
		_w4823_,
		_w4824_,
		_w4825_
	);
	LUT2 #(
		.INIT('h1)
	) name3318 (
		_w4812_,
		_w4825_,
		_w4826_
	);
	LUT2 #(
		.INIT('h2)
	) name3319 (
		_w2040_,
		_w4613_,
		_w4827_
	);
	LUT2 #(
		.INIT('h2)
	) name3320 (
		\TM0_pad ,
		\_2122__reg/NET0131 ,
		_w4828_
	);
	LUT2 #(
		.INIT('h2)
	) name3321 (
		_w1976_,
		_w4828_,
		_w4829_
	);
	LUT2 #(
		.INIT('h4)
	) name3322 (
		_w2527_,
		_w4829_,
		_w4830_
	);
	LUT2 #(
		.INIT('h1)
	) name3323 (
		_w4827_,
		_w4830_,
		_w4831_
	);
	LUT2 #(
		.INIT('h2)
	) name3324 (
		_w4510_,
		_w4674_,
		_w4832_
	);
	LUT2 #(
		.INIT('h2)
	) name3325 (
		\TM0_pad ,
		\_2205__reg/NET0131 ,
		_w4833_
	);
	LUT2 #(
		.INIT('h2)
	) name3326 (
		\WX7300_reg/NET0131 ,
		\WX7364_reg/NET0131 ,
		_w4834_
	);
	LUT2 #(
		.INIT('h4)
	) name3327 (
		\WX7300_reg/NET0131 ,
		\WX7364_reg/NET0131 ,
		_w4835_
	);
	LUT2 #(
		.INIT('h1)
	) name3328 (
		_w4834_,
		_w4835_,
		_w4836_
	);
	LUT2 #(
		.INIT('h2)
	) name3329 (
		\WX7172_reg/NET0131 ,
		\WX7236_reg/NET0131 ,
		_w4837_
	);
	LUT2 #(
		.INIT('h4)
	) name3330 (
		\WX7172_reg/NET0131 ,
		\WX7236_reg/NET0131 ,
		_w4838_
	);
	LUT2 #(
		.INIT('h1)
	) name3331 (
		_w4837_,
		_w4838_,
		_w4839_
	);
	LUT2 #(
		.INIT('h4)
	) name3332 (
		_w4836_,
		_w4839_,
		_w4840_
	);
	LUT2 #(
		.INIT('h2)
	) name3333 (
		_w4836_,
		_w4839_,
		_w4841_
	);
	LUT2 #(
		.INIT('h1)
	) name3334 (
		\TM0_pad ,
		_w4840_,
		_w4842_
	);
	LUT2 #(
		.INIT('h4)
	) name3335 (
		_w4841_,
		_w4842_,
		_w4843_
	);
	LUT2 #(
		.INIT('h2)
	) name3336 (
		_w1976_,
		_w4833_,
		_w4844_
	);
	LUT2 #(
		.INIT('h4)
	) name3337 (
		_w4843_,
		_w4844_,
		_w4845_
	);
	LUT2 #(
		.INIT('h1)
	) name3338 (
		_w4832_,
		_w4845_,
		_w4846_
	);
	LUT2 #(
		.INIT('h8)
	) name3339 (
		\TM0_pad ,
		\_2171__reg/NET0131 ,
		_w4847_
	);
	LUT2 #(
		.INIT('h2)
	) name3340 (
		\WX4654_reg/NET0131 ,
		\WX4718_reg/NET0131 ,
		_w4848_
	);
	LUT2 #(
		.INIT('h4)
	) name3341 (
		\WX4654_reg/NET0131 ,
		\WX4718_reg/NET0131 ,
		_w4849_
	);
	LUT2 #(
		.INIT('h1)
	) name3342 (
		_w4848_,
		_w4849_,
		_w4850_
	);
	LUT2 #(
		.INIT('h2)
	) name3343 (
		\WX4590_reg/NET0131 ,
		_w4850_,
		_w4851_
	);
	LUT2 #(
		.INIT('h4)
	) name3344 (
		\WX4590_reg/NET0131 ,
		_w4850_,
		_w4852_
	);
	LUT2 #(
		.INIT('h1)
	) name3345 (
		_w4851_,
		_w4852_,
		_w4853_
	);
	LUT2 #(
		.INIT('h2)
	) name3346 (
		\TM1_pad ,
		\WX4526_reg/NET0131 ,
		_w4854_
	);
	LUT2 #(
		.INIT('h4)
	) name3347 (
		\TM1_pad ,
		\WX4526_reg/NET0131 ,
		_w4855_
	);
	LUT2 #(
		.INIT('h1)
	) name3348 (
		_w4854_,
		_w4855_,
		_w4856_
	);
	LUT2 #(
		.INIT('h4)
	) name3349 (
		_w4853_,
		_w4856_,
		_w4857_
	);
	LUT2 #(
		.INIT('h2)
	) name3350 (
		_w4853_,
		_w4856_,
		_w4858_
	);
	LUT2 #(
		.INIT('h1)
	) name3351 (
		\TM0_pad ,
		_w4857_,
		_w4859_
	);
	LUT2 #(
		.INIT('h4)
	) name3352 (
		_w4858_,
		_w4859_,
		_w4860_
	);
	LUT2 #(
		.INIT('h1)
	) name3353 (
		_w4847_,
		_w4860_,
		_w4861_
	);
	LUT2 #(
		.INIT('h2)
	) name3354 (
		_w1976_,
		_w4861_,
		_w4862_
	);
	LUT2 #(
		.INIT('h1)
	) name3355 (
		_w1855_,
		_w2135_,
		_w4863_
	);
	LUT2 #(
		.INIT('h2)
	) name3356 (
		_w1973_,
		_w4863_,
		_w4864_
	);
	LUT2 #(
		.INIT('h1)
	) name3357 (
		_w4862_,
		_w4864_,
		_w4865_
	);
	LUT2 #(
		.INIT('h8)
	) name3358 (
		RESET_pad,
		\WX10863_reg/NET0131 ,
		_w4866_
	);
	LUT2 #(
		.INIT('h2)
	) name3359 (
		_w4510_,
		_w4843_,
		_w4867_
	);
	LUT2 #(
		.INIT('h2)
	) name3360 (
		\TM0_pad ,
		\_2237__reg/NET0131 ,
		_w4868_
	);
	LUT2 #(
		.INIT('h2)
	) name3361 (
		\WX8593_reg/NET0131 ,
		\WX8657_reg/NET0131 ,
		_w4869_
	);
	LUT2 #(
		.INIT('h4)
	) name3362 (
		\WX8593_reg/NET0131 ,
		\WX8657_reg/NET0131 ,
		_w4870_
	);
	LUT2 #(
		.INIT('h1)
	) name3363 (
		_w4869_,
		_w4870_,
		_w4871_
	);
	LUT2 #(
		.INIT('h2)
	) name3364 (
		\WX8465_reg/NET0131 ,
		\WX8529_reg/NET0131 ,
		_w4872_
	);
	LUT2 #(
		.INIT('h4)
	) name3365 (
		\WX8465_reg/NET0131 ,
		\WX8529_reg/NET0131 ,
		_w4873_
	);
	LUT2 #(
		.INIT('h1)
	) name3366 (
		_w4872_,
		_w4873_,
		_w4874_
	);
	LUT2 #(
		.INIT('h4)
	) name3367 (
		_w4871_,
		_w4874_,
		_w4875_
	);
	LUT2 #(
		.INIT('h2)
	) name3368 (
		_w4871_,
		_w4874_,
		_w4876_
	);
	LUT2 #(
		.INIT('h1)
	) name3369 (
		\TM0_pad ,
		_w4875_,
		_w4877_
	);
	LUT2 #(
		.INIT('h4)
	) name3370 (
		_w4876_,
		_w4877_,
		_w4878_
	);
	LUT2 #(
		.INIT('h2)
	) name3371 (
		_w1976_,
		_w4868_,
		_w4879_
	);
	LUT2 #(
		.INIT('h4)
	) name3372 (
		_w4878_,
		_w4879_,
		_w4880_
	);
	LUT2 #(
		.INIT('h1)
	) name3373 (
		_w4867_,
		_w4880_,
		_w4881_
	);
	LUT2 #(
		.INIT('h2)
	) name3374 (
		_w4382_,
		_w4774_,
		_w4882_
	);
	LUT2 #(
		.INIT('h2)
	) name3375 (
		\TM0_pad ,
		\_2270__reg/NET0131 ,
		_w4883_
	);
	LUT2 #(
		.INIT('h2)
	) name3376 (
		\WX9884_reg/NET0131 ,
		\WX9948_reg/NET0131 ,
		_w4884_
	);
	LUT2 #(
		.INIT('h4)
	) name3377 (
		\WX9884_reg/NET0131 ,
		\WX9948_reg/NET0131 ,
		_w4885_
	);
	LUT2 #(
		.INIT('h1)
	) name3378 (
		_w4884_,
		_w4885_,
		_w4886_
	);
	LUT2 #(
		.INIT('h2)
	) name3379 (
		\WX9756_reg/NET0131 ,
		\WX9820_reg/NET0131 ,
		_w4887_
	);
	LUT2 #(
		.INIT('h4)
	) name3380 (
		\WX9756_reg/NET0131 ,
		\WX9820_reg/NET0131 ,
		_w4888_
	);
	LUT2 #(
		.INIT('h1)
	) name3381 (
		_w4887_,
		_w4888_,
		_w4889_
	);
	LUT2 #(
		.INIT('h4)
	) name3382 (
		_w4886_,
		_w4889_,
		_w4890_
	);
	LUT2 #(
		.INIT('h2)
	) name3383 (
		_w4886_,
		_w4889_,
		_w4891_
	);
	LUT2 #(
		.INIT('h1)
	) name3384 (
		\TM0_pad ,
		_w4890_,
		_w4892_
	);
	LUT2 #(
		.INIT('h4)
	) name3385 (
		_w4891_,
		_w4892_,
		_w4893_
	);
	LUT2 #(
		.INIT('h2)
	) name3386 (
		_w1976_,
		_w4883_,
		_w4894_
	);
	LUT2 #(
		.INIT('h4)
	) name3387 (
		_w4893_,
		_w4894_,
		_w4895_
	);
	LUT2 #(
		.INIT('h1)
	) name3388 (
		_w4882_,
		_w4895_,
		_w4896_
	);
	LUT2 #(
		.INIT('h8)
	) name3389 (
		\TM0_pad ,
		\_2203__reg/NET0131 ,
		_w4897_
	);
	LUT2 #(
		.INIT('h2)
	) name3390 (
		\WX5947_reg/NET0131 ,
		\WX6011_reg/NET0131 ,
		_w4898_
	);
	LUT2 #(
		.INIT('h4)
	) name3391 (
		\WX5947_reg/NET0131 ,
		\WX6011_reg/NET0131 ,
		_w4899_
	);
	LUT2 #(
		.INIT('h1)
	) name3392 (
		_w4898_,
		_w4899_,
		_w4900_
	);
	LUT2 #(
		.INIT('h2)
	) name3393 (
		\WX5883_reg/NET0131 ,
		_w4900_,
		_w4901_
	);
	LUT2 #(
		.INIT('h4)
	) name3394 (
		\WX5883_reg/NET0131 ,
		_w4900_,
		_w4902_
	);
	LUT2 #(
		.INIT('h1)
	) name3395 (
		_w4901_,
		_w4902_,
		_w4903_
	);
	LUT2 #(
		.INIT('h2)
	) name3396 (
		\TM1_pad ,
		\WX5819_reg/NET0131 ,
		_w4904_
	);
	LUT2 #(
		.INIT('h4)
	) name3397 (
		\TM1_pad ,
		\WX5819_reg/NET0131 ,
		_w4905_
	);
	LUT2 #(
		.INIT('h1)
	) name3398 (
		_w4904_,
		_w4905_,
		_w4906_
	);
	LUT2 #(
		.INIT('h4)
	) name3399 (
		_w4903_,
		_w4906_,
		_w4907_
	);
	LUT2 #(
		.INIT('h2)
	) name3400 (
		_w4903_,
		_w4906_,
		_w4908_
	);
	LUT2 #(
		.INIT('h1)
	) name3401 (
		\TM0_pad ,
		_w4907_,
		_w4909_
	);
	LUT2 #(
		.INIT('h4)
	) name3402 (
		_w4908_,
		_w4909_,
		_w4910_
	);
	LUT2 #(
		.INIT('h1)
	) name3403 (
		_w4897_,
		_w4910_,
		_w4911_
	);
	LUT2 #(
		.INIT('h2)
	) name3404 (
		_w1976_,
		_w4911_,
		_w4912_
	);
	LUT2 #(
		.INIT('h1)
	) name3405 (
		_w1855_,
		_w4860_,
		_w4913_
	);
	LUT2 #(
		.INIT('h2)
	) name3406 (
		_w1973_,
		_w4913_,
		_w4914_
	);
	LUT2 #(
		.INIT('h1)
	) name3407 (
		_w4912_,
		_w4914_,
		_w4915_
	);
	LUT2 #(
		.INIT('h2)
	) name3408 (
		_w4239_,
		_w4789_,
		_w4916_
	);
	LUT2 #(
		.INIT('h2)
	) name3409 (
		\TM0_pad ,
		\_2303__reg/NET0131 ,
		_w4917_
	);
	LUT2 #(
		.INIT('h2)
	) name3410 (
		\WX11175_reg/NET0131 ,
		\WX11239_reg/NET0131 ,
		_w4918_
	);
	LUT2 #(
		.INIT('h4)
	) name3411 (
		\WX11175_reg/NET0131 ,
		\WX11239_reg/NET0131 ,
		_w4919_
	);
	LUT2 #(
		.INIT('h1)
	) name3412 (
		_w4918_,
		_w4919_,
		_w4920_
	);
	LUT2 #(
		.INIT('h2)
	) name3413 (
		\WX11047_reg/NET0131 ,
		\WX11111_reg/NET0131 ,
		_w4921_
	);
	LUT2 #(
		.INIT('h4)
	) name3414 (
		\WX11047_reg/NET0131 ,
		\WX11111_reg/NET0131 ,
		_w4922_
	);
	LUT2 #(
		.INIT('h1)
	) name3415 (
		_w4921_,
		_w4922_,
		_w4923_
	);
	LUT2 #(
		.INIT('h4)
	) name3416 (
		_w4920_,
		_w4923_,
		_w4924_
	);
	LUT2 #(
		.INIT('h2)
	) name3417 (
		_w4920_,
		_w4923_,
		_w4925_
	);
	LUT2 #(
		.INIT('h1)
	) name3418 (
		\TM0_pad ,
		_w4924_,
		_w4926_
	);
	LUT2 #(
		.INIT('h4)
	) name3419 (
		_w4925_,
		_w4926_,
		_w4927_
	);
	LUT2 #(
		.INIT('h2)
	) name3420 (
		_w1976_,
		_w4917_,
		_w4928_
	);
	LUT2 #(
		.INIT('h4)
	) name3421 (
		_w4927_,
		_w4928_,
		_w4929_
	);
	LUT2 #(
		.INIT('h1)
	) name3422 (
		_w4916_,
		_w4929_,
		_w4930_
	);
	LUT2 #(
		.INIT('h8)
	) name3423 (
		\TM0_pad ,
		\_2236__reg/NET0131 ,
		_w4931_
	);
	LUT2 #(
		.INIT('h2)
	) name3424 (
		\WX7238_reg/NET0131 ,
		\WX7302_reg/NET0131 ,
		_w4932_
	);
	LUT2 #(
		.INIT('h4)
	) name3425 (
		\WX7238_reg/NET0131 ,
		\WX7302_reg/NET0131 ,
		_w4933_
	);
	LUT2 #(
		.INIT('h1)
	) name3426 (
		_w4932_,
		_w4933_,
		_w4934_
	);
	LUT2 #(
		.INIT('h2)
	) name3427 (
		\WX7174_reg/NET0131 ,
		_w4934_,
		_w4935_
	);
	LUT2 #(
		.INIT('h4)
	) name3428 (
		\WX7174_reg/NET0131 ,
		_w4934_,
		_w4936_
	);
	LUT2 #(
		.INIT('h1)
	) name3429 (
		_w4935_,
		_w4936_,
		_w4937_
	);
	LUT2 #(
		.INIT('h2)
	) name3430 (
		\TM1_pad ,
		\WX7110_reg/NET0131 ,
		_w4938_
	);
	LUT2 #(
		.INIT('h4)
	) name3431 (
		\TM1_pad ,
		\WX7110_reg/NET0131 ,
		_w4939_
	);
	LUT2 #(
		.INIT('h1)
	) name3432 (
		_w4938_,
		_w4939_,
		_w4940_
	);
	LUT2 #(
		.INIT('h4)
	) name3433 (
		_w4937_,
		_w4940_,
		_w4941_
	);
	LUT2 #(
		.INIT('h2)
	) name3434 (
		_w4937_,
		_w4940_,
		_w4942_
	);
	LUT2 #(
		.INIT('h1)
	) name3435 (
		\TM0_pad ,
		_w4941_,
		_w4943_
	);
	LUT2 #(
		.INIT('h4)
	) name3436 (
		_w4942_,
		_w4943_,
		_w4944_
	);
	LUT2 #(
		.INIT('h1)
	) name3437 (
		_w4931_,
		_w4944_,
		_w4945_
	);
	LUT2 #(
		.INIT('h2)
	) name3438 (
		_w1976_,
		_w4945_,
		_w4946_
	);
	LUT2 #(
		.INIT('h1)
	) name3439 (
		_w1871_,
		_w4806_,
		_w4947_
	);
	LUT2 #(
		.INIT('h2)
	) name3440 (
		_w1973_,
		_w4947_,
		_w4948_
	);
	LUT2 #(
		.INIT('h1)
	) name3441 (
		_w4946_,
		_w4948_,
		_w4949_
	);
	LUT2 #(
		.INIT('h2)
	) name3442 (
		_w2677_,
		_w4752_,
		_w4950_
	);
	LUT2 #(
		.INIT('h2)
	) name3443 (
		\TM0_pad ,
		\_2121__reg/NET0131 ,
		_w4951_
	);
	LUT2 #(
		.INIT('h2)
	) name3444 (
		_w1976_,
		_w4951_,
		_w4952_
	);
	LUT2 #(
		.INIT('h4)
	) name3445 (
		_w2687_,
		_w4952_,
		_w4953_
	);
	LUT2 #(
		.INIT('h1)
	) name3446 (
		_w4950_,
		_w4953_,
		_w4954_
	);
	LUT2 #(
		.INIT('h8)
	) name3447 (
		\TM0_pad ,
		\_2170__reg/NET0131 ,
		_w4955_
	);
	LUT2 #(
		.INIT('h2)
	) name3448 (
		\WX4656_reg/NET0131 ,
		\WX4720_reg/NET0131 ,
		_w4956_
	);
	LUT2 #(
		.INIT('h4)
	) name3449 (
		\WX4656_reg/NET0131 ,
		\WX4720_reg/NET0131 ,
		_w4957_
	);
	LUT2 #(
		.INIT('h1)
	) name3450 (
		_w4956_,
		_w4957_,
		_w4958_
	);
	LUT2 #(
		.INIT('h2)
	) name3451 (
		\WX4592_reg/NET0131 ,
		_w4958_,
		_w4959_
	);
	LUT2 #(
		.INIT('h4)
	) name3452 (
		\WX4592_reg/NET0131 ,
		_w4958_,
		_w4960_
	);
	LUT2 #(
		.INIT('h1)
	) name3453 (
		_w4959_,
		_w4960_,
		_w4961_
	);
	LUT2 #(
		.INIT('h2)
	) name3454 (
		\TM1_pad ,
		\WX4528_reg/NET0131 ,
		_w4962_
	);
	LUT2 #(
		.INIT('h4)
	) name3455 (
		\TM1_pad ,
		\WX4528_reg/NET0131 ,
		_w4963_
	);
	LUT2 #(
		.INIT('h1)
	) name3456 (
		_w4962_,
		_w4963_,
		_w4964_
	);
	LUT2 #(
		.INIT('h4)
	) name3457 (
		_w4961_,
		_w4964_,
		_w4965_
	);
	LUT2 #(
		.INIT('h2)
	) name3458 (
		_w4961_,
		_w4964_,
		_w4966_
	);
	LUT2 #(
		.INIT('h1)
	) name3459 (
		\TM0_pad ,
		_w4965_,
		_w4967_
	);
	LUT2 #(
		.INIT('h4)
	) name3460 (
		_w4966_,
		_w4967_,
		_w4968_
	);
	LUT2 #(
		.INIT('h1)
	) name3461 (
		_w4955_,
		_w4968_,
		_w4969_
	);
	LUT2 #(
		.INIT('h2)
	) name3462 (
		_w1976_,
		_w4969_,
		_w4970_
	);
	LUT2 #(
		.INIT('h1)
	) name3463 (
		_w1826_,
		_w2399_,
		_w4971_
	);
	LUT2 #(
		.INIT('h2)
	) name3464 (
		_w1973_,
		_w4971_,
		_w4972_
	);
	LUT2 #(
		.INIT('h1)
	) name3465 (
		_w4970_,
		_w4972_,
		_w4973_
	);
	LUT2 #(
		.INIT('h1)
	) name3466 (
		\TM0_pad ,
		_w1530_,
		_w4974_
	);
	LUT2 #(
		.INIT('h2)
	) name3467 (
		_w3011_,
		_w4974_,
		_w4975_
	);
	LUT2 #(
		.INIT('h2)
	) name3468 (
		\TM0_pad ,
		\_2087__reg/NET0131 ,
		_w4976_
	);
	LUT2 #(
		.INIT('h2)
	) name3469 (
		\WX2108_reg/NET0131 ,
		\WX2172_reg/NET0131 ,
		_w4977_
	);
	LUT2 #(
		.INIT('h4)
	) name3470 (
		\WX2108_reg/NET0131 ,
		\WX2172_reg/NET0131 ,
		_w4978_
	);
	LUT2 #(
		.INIT('h1)
	) name3471 (
		_w4977_,
		_w4978_,
		_w4979_
	);
	LUT2 #(
		.INIT('h2)
	) name3472 (
		\WX1980_reg/NET0131 ,
		\WX2044_reg/NET0131 ,
		_w4980_
	);
	LUT2 #(
		.INIT('h4)
	) name3473 (
		\WX1980_reg/NET0131 ,
		\WX2044_reg/NET0131 ,
		_w4981_
	);
	LUT2 #(
		.INIT('h1)
	) name3474 (
		_w4980_,
		_w4981_,
		_w4982_
	);
	LUT2 #(
		.INIT('h4)
	) name3475 (
		_w4979_,
		_w4982_,
		_w4983_
	);
	LUT2 #(
		.INIT('h2)
	) name3476 (
		_w4979_,
		_w4982_,
		_w4984_
	);
	LUT2 #(
		.INIT('h1)
	) name3477 (
		\TM0_pad ,
		_w4983_,
		_w4985_
	);
	LUT2 #(
		.INIT('h4)
	) name3478 (
		_w4984_,
		_w4985_,
		_w4986_
	);
	LUT2 #(
		.INIT('h2)
	) name3479 (
		_w1976_,
		_w4976_,
		_w4987_
	);
	LUT2 #(
		.INIT('h4)
	) name3480 (
		_w4986_,
		_w4987_,
		_w4988_
	);
	LUT2 #(
		.INIT('h1)
	) name3481 (
		_w4975_,
		_w4988_,
		_w4989_
	);
	LUT2 #(
		.INIT('h2)
	) name3482 (
		_w2677_,
		_w3535_,
		_w4990_
	);
	LUT2 #(
		.INIT('h1)
	) name3483 (
		\DATA_0_12_pad ,
		\TM0_pad ,
		_w4991_
	);
	LUT2 #(
		.INIT('h2)
	) name3484 (
		\TM0_pad ,
		\_2345__reg/NET0131 ,
		_w4992_
	);
	LUT2 #(
		.INIT('h2)
	) name3485 (
		_w1976_,
		_w4991_,
		_w4993_
	);
	LUT2 #(
		.INIT('h4)
	) name3486 (
		_w4992_,
		_w4993_,
		_w4994_
	);
	LUT2 #(
		.INIT('h1)
	) name3487 (
		_w4990_,
		_w4994_,
		_w4995_
	);
	LUT2 #(
		.INIT('h8)
	) name3488 (
		RESET_pad,
		\WX10865_reg/NET0131 ,
		_w4996_
	);
	LUT2 #(
		.INIT('h2)
	) name3489 (
		_w4510_,
		_w4878_,
		_w4997_
	);
	LUT2 #(
		.INIT('h2)
	) name3490 (
		\TM0_pad ,
		\_2269__reg/NET0131 ,
		_w4998_
	);
	LUT2 #(
		.INIT('h2)
	) name3491 (
		\WX9886_reg/NET0131 ,
		\WX9950_reg/NET0131 ,
		_w4999_
	);
	LUT2 #(
		.INIT('h4)
	) name3492 (
		\WX9886_reg/NET0131 ,
		\WX9950_reg/NET0131 ,
		_w5000_
	);
	LUT2 #(
		.INIT('h1)
	) name3493 (
		_w4999_,
		_w5000_,
		_w5001_
	);
	LUT2 #(
		.INIT('h2)
	) name3494 (
		\WX9758_reg/NET0131 ,
		\WX9822_reg/NET0131 ,
		_w5002_
	);
	LUT2 #(
		.INIT('h4)
	) name3495 (
		\WX9758_reg/NET0131 ,
		\WX9822_reg/NET0131 ,
		_w5003_
	);
	LUT2 #(
		.INIT('h1)
	) name3496 (
		_w5002_,
		_w5003_,
		_w5004_
	);
	LUT2 #(
		.INIT('h4)
	) name3497 (
		_w5001_,
		_w5004_,
		_w5005_
	);
	LUT2 #(
		.INIT('h2)
	) name3498 (
		_w5001_,
		_w5004_,
		_w5006_
	);
	LUT2 #(
		.INIT('h1)
	) name3499 (
		\TM0_pad ,
		_w5005_,
		_w5007_
	);
	LUT2 #(
		.INIT('h4)
	) name3500 (
		_w5006_,
		_w5007_,
		_w5008_
	);
	LUT2 #(
		.INIT('h2)
	) name3501 (
		_w1976_,
		_w4998_,
		_w5009_
	);
	LUT2 #(
		.INIT('h4)
	) name3502 (
		_w5008_,
		_w5009_,
		_w5010_
	);
	LUT2 #(
		.INIT('h1)
	) name3503 (
		_w4997_,
		_w5010_,
		_w5011_
	);
	LUT2 #(
		.INIT('h8)
	) name3504 (
		\TM0_pad ,
		\_2202__reg/NET0131 ,
		_w5012_
	);
	LUT2 #(
		.INIT('h2)
	) name3505 (
		\WX5949_reg/NET0131 ,
		\WX6013_reg/NET0131 ,
		_w5013_
	);
	LUT2 #(
		.INIT('h4)
	) name3506 (
		\WX5949_reg/NET0131 ,
		\WX6013_reg/NET0131 ,
		_w5014_
	);
	LUT2 #(
		.INIT('h1)
	) name3507 (
		_w5013_,
		_w5014_,
		_w5015_
	);
	LUT2 #(
		.INIT('h2)
	) name3508 (
		\WX5885_reg/NET0131 ,
		_w5015_,
		_w5016_
	);
	LUT2 #(
		.INIT('h4)
	) name3509 (
		\WX5885_reg/NET0131 ,
		_w5015_,
		_w5017_
	);
	LUT2 #(
		.INIT('h1)
	) name3510 (
		_w5016_,
		_w5017_,
		_w5018_
	);
	LUT2 #(
		.INIT('h2)
	) name3511 (
		\TM1_pad ,
		\WX5821_reg/NET0131 ,
		_w5019_
	);
	LUT2 #(
		.INIT('h4)
	) name3512 (
		\TM1_pad ,
		\WX5821_reg/NET0131 ,
		_w5020_
	);
	LUT2 #(
		.INIT('h1)
	) name3513 (
		_w5019_,
		_w5020_,
		_w5021_
	);
	LUT2 #(
		.INIT('h4)
	) name3514 (
		_w5018_,
		_w5021_,
		_w5022_
	);
	LUT2 #(
		.INIT('h2)
	) name3515 (
		_w5018_,
		_w5021_,
		_w5023_
	);
	LUT2 #(
		.INIT('h1)
	) name3516 (
		\TM0_pad ,
		_w5022_,
		_w5024_
	);
	LUT2 #(
		.INIT('h4)
	) name3517 (
		_w5023_,
		_w5024_,
		_w5025_
	);
	LUT2 #(
		.INIT('h1)
	) name3518 (
		_w5012_,
		_w5025_,
		_w5026_
	);
	LUT2 #(
		.INIT('h2)
	) name3519 (
		_w1976_,
		_w5026_,
		_w5027_
	);
	LUT2 #(
		.INIT('h1)
	) name3520 (
		_w1826_,
		_w4968_,
		_w5028_
	);
	LUT2 #(
		.INIT('h2)
	) name3521 (
		_w1973_,
		_w5028_,
		_w5029_
	);
	LUT2 #(
		.INIT('h1)
	) name3522 (
		_w5027_,
		_w5029_,
		_w5030_
	);
	LUT2 #(
		.INIT('h2)
	) name3523 (
		_w4382_,
		_w4893_,
		_w5031_
	);
	LUT2 #(
		.INIT('h2)
	) name3524 (
		\TM0_pad ,
		\_2302__reg/NET0131 ,
		_w5032_
	);
	LUT2 #(
		.INIT('h2)
	) name3525 (
		\WX11177_reg/NET0131 ,
		\WX11241_reg/NET0131 ,
		_w5033_
	);
	LUT2 #(
		.INIT('h4)
	) name3526 (
		\WX11177_reg/NET0131 ,
		\WX11241_reg/NET0131 ,
		_w5034_
	);
	LUT2 #(
		.INIT('h1)
	) name3527 (
		_w5033_,
		_w5034_,
		_w5035_
	);
	LUT2 #(
		.INIT('h2)
	) name3528 (
		\WX11049_reg/NET0131 ,
		\WX11113_reg/NET0131 ,
		_w5036_
	);
	LUT2 #(
		.INIT('h4)
	) name3529 (
		\WX11049_reg/NET0131 ,
		\WX11113_reg/NET0131 ,
		_w5037_
	);
	LUT2 #(
		.INIT('h1)
	) name3530 (
		_w5036_,
		_w5037_,
		_w5038_
	);
	LUT2 #(
		.INIT('h4)
	) name3531 (
		_w5035_,
		_w5038_,
		_w5039_
	);
	LUT2 #(
		.INIT('h2)
	) name3532 (
		_w5035_,
		_w5038_,
		_w5040_
	);
	LUT2 #(
		.INIT('h1)
	) name3533 (
		\TM0_pad ,
		_w5039_,
		_w5041_
	);
	LUT2 #(
		.INIT('h4)
	) name3534 (
		_w5040_,
		_w5041_,
		_w5042_
	);
	LUT2 #(
		.INIT('h2)
	) name3535 (
		_w1976_,
		_w5032_,
		_w5043_
	);
	LUT2 #(
		.INIT('h4)
	) name3536 (
		_w5042_,
		_w5043_,
		_w5044_
	);
	LUT2 #(
		.INIT('h1)
	) name3537 (
		_w5031_,
		_w5044_,
		_w5045_
	);
	LUT2 #(
		.INIT('h8)
	) name3538 (
		\TM0_pad ,
		\_2235__reg/NET0131 ,
		_w5046_
	);
	LUT2 #(
		.INIT('h2)
	) name3539 (
		\TM1_pad ,
		\WX7112_reg/NET0131 ,
		_w5047_
	);
	LUT2 #(
		.INIT('h4)
	) name3540 (
		\TM1_pad ,
		\WX7112_reg/NET0131 ,
		_w5048_
	);
	LUT2 #(
		.INIT('h1)
	) name3541 (
		_w5047_,
		_w5048_,
		_w5049_
	);
	LUT2 #(
		.INIT('h1)
	) name3542 (
		\WX7176_reg/NET0131 ,
		_w5049_,
		_w5050_
	);
	LUT2 #(
		.INIT('h8)
	) name3543 (
		\WX7176_reg/NET0131 ,
		_w5049_,
		_w5051_
	);
	LUT2 #(
		.INIT('h1)
	) name3544 (
		_w5050_,
		_w5051_,
		_w5052_
	);
	LUT2 #(
		.INIT('h2)
	) name3545 (
		\WX7240_reg/NET0131 ,
		\WX7304_reg/NET0131 ,
		_w5053_
	);
	LUT2 #(
		.INIT('h4)
	) name3546 (
		\WX7240_reg/NET0131 ,
		\WX7304_reg/NET0131 ,
		_w5054_
	);
	LUT2 #(
		.INIT('h1)
	) name3547 (
		_w5053_,
		_w5054_,
		_w5055_
	);
	LUT2 #(
		.INIT('h1)
	) name3548 (
		_w5052_,
		_w5055_,
		_w5056_
	);
	LUT2 #(
		.INIT('h8)
	) name3549 (
		_w5052_,
		_w5055_,
		_w5057_
	);
	LUT2 #(
		.INIT('h1)
	) name3550 (
		\TM0_pad ,
		_w5056_,
		_w5058_
	);
	LUT2 #(
		.INIT('h4)
	) name3551 (
		_w5057_,
		_w5058_,
		_w5059_
	);
	LUT2 #(
		.INIT('h1)
	) name3552 (
		_w5046_,
		_w5059_,
		_w5060_
	);
	LUT2 #(
		.INIT('h2)
	) name3553 (
		_w1976_,
		_w5060_,
		_w5061_
	);
	LUT2 #(
		.INIT('h1)
	) name3554 (
		_w1855_,
		_w4910_,
		_w5062_
	);
	LUT2 #(
		.INIT('h2)
	) name3555 (
		_w1973_,
		_w5062_,
		_w5063_
	);
	LUT2 #(
		.INIT('h1)
	) name3556 (
		_w5061_,
		_w5063_,
		_w5064_
	);
	LUT2 #(
		.INIT('h2)
	) name3557 (
		\WX2106_reg/NET0131 ,
		\WX2170_reg/NET0131 ,
		_w5065_
	);
	LUT2 #(
		.INIT('h4)
	) name3558 (
		\WX2106_reg/NET0131 ,
		\WX2170_reg/NET0131 ,
		_w5066_
	);
	LUT2 #(
		.INIT('h1)
	) name3559 (
		_w5065_,
		_w5066_,
		_w5067_
	);
	LUT2 #(
		.INIT('h2)
	) name3560 (
		\WX1978_reg/NET0131 ,
		\WX2042_reg/NET0131 ,
		_w5068_
	);
	LUT2 #(
		.INIT('h4)
	) name3561 (
		\WX1978_reg/NET0131 ,
		\WX2042_reg/NET0131 ,
		_w5069_
	);
	LUT2 #(
		.INIT('h1)
	) name3562 (
		_w5068_,
		_w5069_,
		_w5070_
	);
	LUT2 #(
		.INIT('h4)
	) name3563 (
		_w5067_,
		_w5070_,
		_w5071_
	);
	LUT2 #(
		.INIT('h2)
	) name3564 (
		_w5067_,
		_w5070_,
		_w5072_
	);
	LUT2 #(
		.INIT('h1)
	) name3565 (
		\TM0_pad ,
		_w5071_,
		_w5073_
	);
	LUT2 #(
		.INIT('h4)
	) name3566 (
		_w5072_,
		_w5073_,
		_w5074_
	);
	LUT2 #(
		.INIT('h2)
	) name3567 (
		_w2846_,
		_w5074_,
		_w5075_
	);
	LUT2 #(
		.INIT('h2)
	) name3568 (
		\TM0_pad ,
		\_2120__reg/NET0131 ,
		_w5076_
	);
	LUT2 #(
		.INIT('h2)
	) name3569 (
		_w1976_,
		_w5076_,
		_w5077_
	);
	LUT2 #(
		.INIT('h4)
	) name3570 (
		_w2856_,
		_w5077_,
		_w5078_
	);
	LUT2 #(
		.INIT('h1)
	) name3571 (
		_w5075_,
		_w5078_,
		_w5079_
	);
	LUT2 #(
		.INIT('h8)
	) name3572 (
		\TM0_pad ,
		\_2268__reg/NET0131 ,
		_w5080_
	);
	LUT2 #(
		.INIT('h2)
	) name3573 (
		\WX8531_reg/NET0131 ,
		\WX8595_reg/NET0131 ,
		_w5081_
	);
	LUT2 #(
		.INIT('h4)
	) name3574 (
		\WX8531_reg/NET0131 ,
		\WX8595_reg/NET0131 ,
		_w5082_
	);
	LUT2 #(
		.INIT('h1)
	) name3575 (
		_w5081_,
		_w5082_,
		_w5083_
	);
	LUT2 #(
		.INIT('h2)
	) name3576 (
		\WX8467_reg/NET0131 ,
		_w5083_,
		_w5084_
	);
	LUT2 #(
		.INIT('h4)
	) name3577 (
		\WX8467_reg/NET0131 ,
		_w5083_,
		_w5085_
	);
	LUT2 #(
		.INIT('h1)
	) name3578 (
		_w5084_,
		_w5085_,
		_w5086_
	);
	LUT2 #(
		.INIT('h2)
	) name3579 (
		\TM1_pad ,
		\WX8403_reg/NET0131 ,
		_w5087_
	);
	LUT2 #(
		.INIT('h4)
	) name3580 (
		\TM1_pad ,
		\WX8403_reg/NET0131 ,
		_w5088_
	);
	LUT2 #(
		.INIT('h1)
	) name3581 (
		_w5087_,
		_w5088_,
		_w5089_
	);
	LUT2 #(
		.INIT('h4)
	) name3582 (
		_w5086_,
		_w5089_,
		_w5090_
	);
	LUT2 #(
		.INIT('h2)
	) name3583 (
		_w5086_,
		_w5089_,
		_w5091_
	);
	LUT2 #(
		.INIT('h1)
	) name3584 (
		\TM0_pad ,
		_w5090_,
		_w5092_
	);
	LUT2 #(
		.INIT('h4)
	) name3585 (
		_w5091_,
		_w5092_,
		_w5093_
	);
	LUT2 #(
		.INIT('h1)
	) name3586 (
		_w5080_,
		_w5093_,
		_w5094_
	);
	LUT2 #(
		.INIT('h2)
	) name3587 (
		_w1976_,
		_w5094_,
		_w5095_
	);
	LUT2 #(
		.INIT('h1)
	) name3588 (
		_w1871_,
		_w4944_,
		_w5096_
	);
	LUT2 #(
		.INIT('h2)
	) name3589 (
		_w1973_,
		_w5096_,
		_w5097_
	);
	LUT2 #(
		.INIT('h1)
	) name3590 (
		_w5095_,
		_w5097_,
		_w5098_
	);
	LUT2 #(
		.INIT('h8)
	) name3591 (
		\TM0_pad ,
		\_2169__reg/NET0131 ,
		_w5099_
	);
	LUT2 #(
		.INIT('h2)
	) name3592 (
		\WX4658_reg/NET0131 ,
		\WX4722_reg/NET0131 ,
		_w5100_
	);
	LUT2 #(
		.INIT('h4)
	) name3593 (
		\WX4658_reg/NET0131 ,
		\WX4722_reg/NET0131 ,
		_w5101_
	);
	LUT2 #(
		.INIT('h1)
	) name3594 (
		_w5100_,
		_w5101_,
		_w5102_
	);
	LUT2 #(
		.INIT('h2)
	) name3595 (
		\WX4594_reg/NET0131 ,
		_w5102_,
		_w5103_
	);
	LUT2 #(
		.INIT('h4)
	) name3596 (
		\WX4594_reg/NET0131 ,
		_w5102_,
		_w5104_
	);
	LUT2 #(
		.INIT('h1)
	) name3597 (
		_w5103_,
		_w5104_,
		_w5105_
	);
	LUT2 #(
		.INIT('h2)
	) name3598 (
		\TM1_pad ,
		\WX4530_reg/NET0131 ,
		_w5106_
	);
	LUT2 #(
		.INIT('h4)
	) name3599 (
		\TM1_pad ,
		\WX4530_reg/NET0131 ,
		_w5107_
	);
	LUT2 #(
		.INIT('h1)
	) name3600 (
		_w5106_,
		_w5107_,
		_w5108_
	);
	LUT2 #(
		.INIT('h4)
	) name3601 (
		_w5105_,
		_w5108_,
		_w5109_
	);
	LUT2 #(
		.INIT('h2)
	) name3602 (
		_w5105_,
		_w5108_,
		_w5110_
	);
	LUT2 #(
		.INIT('h1)
	) name3603 (
		\TM0_pad ,
		_w5109_,
		_w5111_
	);
	LUT2 #(
		.INIT('h4)
	) name3604 (
		_w5110_,
		_w5111_,
		_w5112_
	);
	LUT2 #(
		.INIT('h1)
	) name3605 (
		_w5099_,
		_w5112_,
		_w5113_
	);
	LUT2 #(
		.INIT('h2)
	) name3606 (
		_w1976_,
		_w5113_,
		_w5114_
	);
	LUT2 #(
		.INIT('h1)
	) name3607 (
		_w1810_,
		_w2575_,
		_w5115_
	);
	LUT2 #(
		.INIT('h2)
	) name3608 (
		_w1973_,
		_w5115_,
		_w5116_
	);
	LUT2 #(
		.INIT('h1)
	) name3609 (
		_w5114_,
		_w5116_,
		_w5117_
	);
	LUT2 #(
		.INIT('h2)
	) name3610 (
		_w2846_,
		_w3696_,
		_w5118_
	);
	LUT2 #(
		.INIT('h1)
	) name3611 (
		\DATA_0_11_pad ,
		\TM0_pad ,
		_w5119_
	);
	LUT2 #(
		.INIT('h2)
	) name3612 (
		\TM0_pad ,
		\_2344__reg/NET0131 ,
		_w5120_
	);
	LUT2 #(
		.INIT('h2)
	) name3613 (
		_w1976_,
		_w5119_,
		_w5121_
	);
	LUT2 #(
		.INIT('h4)
	) name3614 (
		_w5120_,
		_w5121_,
		_w5122_
	);
	LUT2 #(
		.INIT('h1)
	) name3615 (
		_w5118_,
		_w5122_,
		_w5123_
	);
	LUT2 #(
		.INIT('h8)
	) name3616 (
		RESET_pad,
		\WX10867_reg/NET0131 ,
		_w5124_
	);
	LUT2 #(
		.INIT('h8)
	) name3617 (
		\TM0_pad ,
		\_2300__reg/NET0131 ,
		_w5125_
	);
	LUT2 #(
		.INIT('h2)
	) name3618 (
		\WX9824_reg/NET0131 ,
		\WX9888_reg/NET0131 ,
		_w5126_
	);
	LUT2 #(
		.INIT('h4)
	) name3619 (
		\WX9824_reg/NET0131 ,
		\WX9888_reg/NET0131 ,
		_w5127_
	);
	LUT2 #(
		.INIT('h1)
	) name3620 (
		_w5126_,
		_w5127_,
		_w5128_
	);
	LUT2 #(
		.INIT('h2)
	) name3621 (
		\WX9760_reg/NET0131 ,
		_w5128_,
		_w5129_
	);
	LUT2 #(
		.INIT('h4)
	) name3622 (
		\WX9760_reg/NET0131 ,
		_w5128_,
		_w5130_
	);
	LUT2 #(
		.INIT('h1)
	) name3623 (
		_w5129_,
		_w5130_,
		_w5131_
	);
	LUT2 #(
		.INIT('h2)
	) name3624 (
		\TM1_pad ,
		\WX9696_reg/NET0131 ,
		_w5132_
	);
	LUT2 #(
		.INIT('h4)
	) name3625 (
		\TM1_pad ,
		\WX9696_reg/NET0131 ,
		_w5133_
	);
	LUT2 #(
		.INIT('h1)
	) name3626 (
		_w5132_,
		_w5133_,
		_w5134_
	);
	LUT2 #(
		.INIT('h4)
	) name3627 (
		_w5131_,
		_w5134_,
		_w5135_
	);
	LUT2 #(
		.INIT('h2)
	) name3628 (
		_w5131_,
		_w5134_,
		_w5136_
	);
	LUT2 #(
		.INIT('h1)
	) name3629 (
		\TM0_pad ,
		_w5135_,
		_w5137_
	);
	LUT2 #(
		.INIT('h4)
	) name3630 (
		_w5136_,
		_w5137_,
		_w5138_
	);
	LUT2 #(
		.INIT('h1)
	) name3631 (
		_w5125_,
		_w5138_,
		_w5139_
	);
	LUT2 #(
		.INIT('h2)
	) name3632 (
		_w1976_,
		_w5139_,
		_w5140_
	);
	LUT2 #(
		.INIT('h1)
	) name3633 (
		_w1871_,
		_w5093_,
		_w5141_
	);
	LUT2 #(
		.INIT('h2)
	) name3634 (
		_w1973_,
		_w5141_,
		_w5142_
	);
	LUT2 #(
		.INIT('h1)
	) name3635 (
		_w5140_,
		_w5142_,
		_w5143_
	);
	LUT2 #(
		.INIT('h8)
	) name3636 (
		\TM0_pad ,
		\_2201__reg/NET0131 ,
		_w5144_
	);
	LUT2 #(
		.INIT('h2)
	) name3637 (
		\WX5951_reg/NET0131 ,
		\WX6015_reg/NET0131 ,
		_w5145_
	);
	LUT2 #(
		.INIT('h4)
	) name3638 (
		\WX5951_reg/NET0131 ,
		\WX6015_reg/NET0131 ,
		_w5146_
	);
	LUT2 #(
		.INIT('h1)
	) name3639 (
		_w5145_,
		_w5146_,
		_w5147_
	);
	LUT2 #(
		.INIT('h2)
	) name3640 (
		\WX5887_reg/NET0131 ,
		_w5147_,
		_w5148_
	);
	LUT2 #(
		.INIT('h4)
	) name3641 (
		\WX5887_reg/NET0131 ,
		_w5147_,
		_w5149_
	);
	LUT2 #(
		.INIT('h1)
	) name3642 (
		_w5148_,
		_w5149_,
		_w5150_
	);
	LUT2 #(
		.INIT('h2)
	) name3643 (
		\TM1_pad ,
		\WX5823_reg/NET0131 ,
		_w5151_
	);
	LUT2 #(
		.INIT('h4)
	) name3644 (
		\TM1_pad ,
		\WX5823_reg/NET0131 ,
		_w5152_
	);
	LUT2 #(
		.INIT('h1)
	) name3645 (
		_w5151_,
		_w5152_,
		_w5153_
	);
	LUT2 #(
		.INIT('h4)
	) name3646 (
		_w5150_,
		_w5153_,
		_w5154_
	);
	LUT2 #(
		.INIT('h2)
	) name3647 (
		_w5150_,
		_w5153_,
		_w5155_
	);
	LUT2 #(
		.INIT('h1)
	) name3648 (
		\TM0_pad ,
		_w5154_,
		_w5156_
	);
	LUT2 #(
		.INIT('h4)
	) name3649 (
		_w5155_,
		_w5156_,
		_w5157_
	);
	LUT2 #(
		.INIT('h1)
	) name3650 (
		_w5144_,
		_w5157_,
		_w5158_
	);
	LUT2 #(
		.INIT('h2)
	) name3651 (
		_w1976_,
		_w5158_,
		_w5159_
	);
	LUT2 #(
		.INIT('h1)
	) name3652 (
		_w1810_,
		_w5112_,
		_w5160_
	);
	LUT2 #(
		.INIT('h2)
	) name3653 (
		_w1973_,
		_w5160_,
		_w5161_
	);
	LUT2 #(
		.INIT('h1)
	) name3654 (
		_w5159_,
		_w5161_,
		_w5162_
	);
	LUT2 #(
		.INIT('h2)
	) name3655 (
		_w4510_,
		_w5008_,
		_w5163_
	);
	LUT2 #(
		.INIT('h2)
	) name3656 (
		\TM0_pad ,
		\_2301__reg/NET0131 ,
		_w5164_
	);
	LUT2 #(
		.INIT('h2)
	) name3657 (
		\WX11179_reg/NET0131 ,
		\WX11243_reg/NET0131 ,
		_w5165_
	);
	LUT2 #(
		.INIT('h4)
	) name3658 (
		\WX11179_reg/NET0131 ,
		\WX11243_reg/NET0131 ,
		_w5166_
	);
	LUT2 #(
		.INIT('h1)
	) name3659 (
		_w5165_,
		_w5166_,
		_w5167_
	);
	LUT2 #(
		.INIT('h2)
	) name3660 (
		\WX11051_reg/NET0131 ,
		\WX11115_reg/NET0131 ,
		_w5168_
	);
	LUT2 #(
		.INIT('h4)
	) name3661 (
		\WX11051_reg/NET0131 ,
		\WX11115_reg/NET0131 ,
		_w5169_
	);
	LUT2 #(
		.INIT('h1)
	) name3662 (
		_w5168_,
		_w5169_,
		_w5170_
	);
	LUT2 #(
		.INIT('h4)
	) name3663 (
		_w5167_,
		_w5170_,
		_w5171_
	);
	LUT2 #(
		.INIT('h2)
	) name3664 (
		_w5167_,
		_w5170_,
		_w5172_
	);
	LUT2 #(
		.INIT('h1)
	) name3665 (
		\TM0_pad ,
		_w5171_,
		_w5173_
	);
	LUT2 #(
		.INIT('h4)
	) name3666 (
		_w5172_,
		_w5173_,
		_w5174_
	);
	LUT2 #(
		.INIT('h2)
	) name3667 (
		_w1976_,
		_w5164_,
		_w5175_
	);
	LUT2 #(
		.INIT('h4)
	) name3668 (
		_w5174_,
		_w5175_,
		_w5176_
	);
	LUT2 #(
		.INIT('h1)
	) name3669 (
		_w5163_,
		_w5176_,
		_w5177_
	);
	LUT2 #(
		.INIT('h8)
	) name3670 (
		\TM0_pad ,
		\_2234__reg/NET0131 ,
		_w5178_
	);
	LUT2 #(
		.INIT('h2)
	) name3671 (
		\WX7242_reg/NET0131 ,
		\WX7306_reg/NET0131 ,
		_w5179_
	);
	LUT2 #(
		.INIT('h4)
	) name3672 (
		\WX7242_reg/NET0131 ,
		\WX7306_reg/NET0131 ,
		_w5180_
	);
	LUT2 #(
		.INIT('h1)
	) name3673 (
		_w5179_,
		_w5180_,
		_w5181_
	);
	LUT2 #(
		.INIT('h2)
	) name3674 (
		\WX7178_reg/NET0131 ,
		_w5181_,
		_w5182_
	);
	LUT2 #(
		.INIT('h4)
	) name3675 (
		\WX7178_reg/NET0131 ,
		_w5181_,
		_w5183_
	);
	LUT2 #(
		.INIT('h1)
	) name3676 (
		_w5182_,
		_w5183_,
		_w5184_
	);
	LUT2 #(
		.INIT('h2)
	) name3677 (
		\TM1_pad ,
		\WX7114_reg/NET0131 ,
		_w5185_
	);
	LUT2 #(
		.INIT('h4)
	) name3678 (
		\TM1_pad ,
		\WX7114_reg/NET0131 ,
		_w5186_
	);
	LUT2 #(
		.INIT('h1)
	) name3679 (
		_w5185_,
		_w5186_,
		_w5187_
	);
	LUT2 #(
		.INIT('h4)
	) name3680 (
		_w5184_,
		_w5187_,
		_w5188_
	);
	LUT2 #(
		.INIT('h2)
	) name3681 (
		_w5184_,
		_w5187_,
		_w5189_
	);
	LUT2 #(
		.INIT('h1)
	) name3682 (
		\TM0_pad ,
		_w5188_,
		_w5190_
	);
	LUT2 #(
		.INIT('h4)
	) name3683 (
		_w5189_,
		_w5190_,
		_w5191_
	);
	LUT2 #(
		.INIT('h1)
	) name3684 (
		_w5178_,
		_w5191_,
		_w5192_
	);
	LUT2 #(
		.INIT('h2)
	) name3685 (
		_w1976_,
		_w5192_,
		_w5193_
	);
	LUT2 #(
		.INIT('h1)
	) name3686 (
		_w1826_,
		_w5025_,
		_w5194_
	);
	LUT2 #(
		.INIT('h2)
	) name3687 (
		_w1973_,
		_w5194_,
		_w5195_
	);
	LUT2 #(
		.INIT('h1)
	) name3688 (
		_w5193_,
		_w5195_,
		_w5196_
	);
	LUT2 #(
		.INIT('h2)
	) name3689 (
		_w3011_,
		_w4986_,
		_w5197_
	);
	LUT2 #(
		.INIT('h2)
	) name3690 (
		\TM0_pad ,
		\_2119__reg/NET0131 ,
		_w5198_
	);
	LUT2 #(
		.INIT('h2)
	) name3691 (
		_w1976_,
		_w5198_,
		_w5199_
	);
	LUT2 #(
		.INIT('h4)
	) name3692 (
		_w3021_,
		_w5199_,
		_w5200_
	);
	LUT2 #(
		.INIT('h1)
	) name3693 (
		_w5197_,
		_w5200_,
		_w5201_
	);
	LUT2 #(
		.INIT('h8)
	) name3694 (
		\TM0_pad ,
		\_2267__reg/NET0131 ,
		_w5202_
	);
	LUT2 #(
		.INIT('h2)
	) name3695 (
		\WX8533_reg/NET0131 ,
		\WX8597_reg/NET0131 ,
		_w5203_
	);
	LUT2 #(
		.INIT('h4)
	) name3696 (
		\WX8533_reg/NET0131 ,
		\WX8597_reg/NET0131 ,
		_w5204_
	);
	LUT2 #(
		.INIT('h1)
	) name3697 (
		_w5203_,
		_w5204_,
		_w5205_
	);
	LUT2 #(
		.INIT('h2)
	) name3698 (
		\WX8469_reg/NET0131 ,
		_w5205_,
		_w5206_
	);
	LUT2 #(
		.INIT('h4)
	) name3699 (
		\WX8469_reg/NET0131 ,
		_w5205_,
		_w5207_
	);
	LUT2 #(
		.INIT('h1)
	) name3700 (
		_w5206_,
		_w5207_,
		_w5208_
	);
	LUT2 #(
		.INIT('h2)
	) name3701 (
		\TM1_pad ,
		\WX8405_reg/NET0131 ,
		_w5209_
	);
	LUT2 #(
		.INIT('h4)
	) name3702 (
		\TM1_pad ,
		\WX8405_reg/NET0131 ,
		_w5210_
	);
	LUT2 #(
		.INIT('h1)
	) name3703 (
		_w5209_,
		_w5210_,
		_w5211_
	);
	LUT2 #(
		.INIT('h4)
	) name3704 (
		_w5208_,
		_w5211_,
		_w5212_
	);
	LUT2 #(
		.INIT('h2)
	) name3705 (
		_w5208_,
		_w5211_,
		_w5213_
	);
	LUT2 #(
		.INIT('h1)
	) name3706 (
		\TM0_pad ,
		_w5212_,
		_w5214_
	);
	LUT2 #(
		.INIT('h4)
	) name3707 (
		_w5213_,
		_w5214_,
		_w5215_
	);
	LUT2 #(
		.INIT('h1)
	) name3708 (
		_w5202_,
		_w5215_,
		_w5216_
	);
	LUT2 #(
		.INIT('h2)
	) name3709 (
		_w1976_,
		_w5216_,
		_w5217_
	);
	LUT2 #(
		.INIT('h1)
	) name3710 (
		_w1855_,
		_w5059_,
		_w5218_
	);
	LUT2 #(
		.INIT('h2)
	) name3711 (
		_w1973_,
		_w5218_,
		_w5219_
	);
	LUT2 #(
		.INIT('h1)
	) name3712 (
		_w5217_,
		_w5219_,
		_w5220_
	);
	LUT2 #(
		.INIT('h8)
	) name3713 (
		\TM0_pad ,
		\_2168__reg/NET0131 ,
		_w5221_
	);
	LUT2 #(
		.INIT('h2)
	) name3714 (
		\WX4660_reg/NET0131 ,
		\WX4724_reg/NET0131 ,
		_w5222_
	);
	LUT2 #(
		.INIT('h4)
	) name3715 (
		\WX4660_reg/NET0131 ,
		\WX4724_reg/NET0131 ,
		_w5223_
	);
	LUT2 #(
		.INIT('h1)
	) name3716 (
		_w5222_,
		_w5223_,
		_w5224_
	);
	LUT2 #(
		.INIT('h2)
	) name3717 (
		\WX4596_reg/NET0131 ,
		_w5224_,
		_w5225_
	);
	LUT2 #(
		.INIT('h4)
	) name3718 (
		\WX4596_reg/NET0131 ,
		_w5224_,
		_w5226_
	);
	LUT2 #(
		.INIT('h1)
	) name3719 (
		_w5225_,
		_w5226_,
		_w5227_
	);
	LUT2 #(
		.INIT('h2)
	) name3720 (
		\TM1_pad ,
		\WX4532_reg/NET0131 ,
		_w5228_
	);
	LUT2 #(
		.INIT('h4)
	) name3721 (
		\TM1_pad ,
		\WX4532_reg/NET0131 ,
		_w5229_
	);
	LUT2 #(
		.INIT('h1)
	) name3722 (
		_w5228_,
		_w5229_,
		_w5230_
	);
	LUT2 #(
		.INIT('h4)
	) name3723 (
		_w5227_,
		_w5230_,
		_w5231_
	);
	LUT2 #(
		.INIT('h2)
	) name3724 (
		_w5227_,
		_w5230_,
		_w5232_
	);
	LUT2 #(
		.INIT('h1)
	) name3725 (
		\TM0_pad ,
		_w5231_,
		_w5233_
	);
	LUT2 #(
		.INIT('h4)
	) name3726 (
		_w5232_,
		_w5233_,
		_w5234_
	);
	LUT2 #(
		.INIT('h1)
	) name3727 (
		_w5221_,
		_w5234_,
		_w5235_
	);
	LUT2 #(
		.INIT('h2)
	) name3728 (
		_w1976_,
		_w5235_,
		_w5236_
	);
	LUT2 #(
		.INIT('h1)
	) name3729 (
		_w1794_,
		_w2735_,
		_w5237_
	);
	LUT2 #(
		.INIT('h2)
	) name3730 (
		_w1973_,
		_w5237_,
		_w5238_
	);
	LUT2 #(
		.INIT('h1)
	) name3731 (
		_w5236_,
		_w5238_,
		_w5239_
	);
	LUT2 #(
		.INIT('h2)
	) name3732 (
		_w3011_,
		_w3857_,
		_w5240_
	);
	LUT2 #(
		.INIT('h1)
	) name3733 (
		\DATA_0_10_pad ,
		\TM0_pad ,
		_w5241_
	);
	LUT2 #(
		.INIT('h2)
	) name3734 (
		\TM0_pad ,
		\_2343__reg/NET0131 ,
		_w5242_
	);
	LUT2 #(
		.INIT('h2)
	) name3735 (
		_w1976_,
		_w5241_,
		_w5243_
	);
	LUT2 #(
		.INIT('h4)
	) name3736 (
		_w5242_,
		_w5243_,
		_w5244_
	);
	LUT2 #(
		.INIT('h1)
	) name3737 (
		_w5240_,
		_w5244_,
		_w5245_
	);
	LUT2 #(
		.INIT('h8)
	) name3738 (
		RESET_pad,
		\WX10869_reg/NET0131 ,
		_w5246_
	);
	LUT2 #(
		.INIT('h8)
	) name3739 (
		\TM0_pad ,
		\_2299__reg/NET0131 ,
		_w5247_
	);
	LUT2 #(
		.INIT('h2)
	) name3740 (
		\WX9826_reg/NET0131 ,
		\WX9890_reg/NET0131 ,
		_w5248_
	);
	LUT2 #(
		.INIT('h4)
	) name3741 (
		\WX9826_reg/NET0131 ,
		\WX9890_reg/NET0131 ,
		_w5249_
	);
	LUT2 #(
		.INIT('h1)
	) name3742 (
		_w5248_,
		_w5249_,
		_w5250_
	);
	LUT2 #(
		.INIT('h2)
	) name3743 (
		\WX9762_reg/NET0131 ,
		_w5250_,
		_w5251_
	);
	LUT2 #(
		.INIT('h4)
	) name3744 (
		\WX9762_reg/NET0131 ,
		_w5250_,
		_w5252_
	);
	LUT2 #(
		.INIT('h1)
	) name3745 (
		_w5251_,
		_w5252_,
		_w5253_
	);
	LUT2 #(
		.INIT('h2)
	) name3746 (
		\TM1_pad ,
		\WX9698_reg/NET0131 ,
		_w5254_
	);
	LUT2 #(
		.INIT('h4)
	) name3747 (
		\TM1_pad ,
		\WX9698_reg/NET0131 ,
		_w5255_
	);
	LUT2 #(
		.INIT('h1)
	) name3748 (
		_w5254_,
		_w5255_,
		_w5256_
	);
	LUT2 #(
		.INIT('h4)
	) name3749 (
		_w5253_,
		_w5256_,
		_w5257_
	);
	LUT2 #(
		.INIT('h2)
	) name3750 (
		_w5253_,
		_w5256_,
		_w5258_
	);
	LUT2 #(
		.INIT('h1)
	) name3751 (
		\TM0_pad ,
		_w5257_,
		_w5259_
	);
	LUT2 #(
		.INIT('h4)
	) name3752 (
		_w5258_,
		_w5259_,
		_w5260_
	);
	LUT2 #(
		.INIT('h1)
	) name3753 (
		_w5247_,
		_w5260_,
		_w5261_
	);
	LUT2 #(
		.INIT('h2)
	) name3754 (
		_w1976_,
		_w5261_,
		_w5262_
	);
	LUT2 #(
		.INIT('h1)
	) name3755 (
		_w1855_,
		_w5215_,
		_w5263_
	);
	LUT2 #(
		.INIT('h2)
	) name3756 (
		_w1973_,
		_w5263_,
		_w5264_
	);
	LUT2 #(
		.INIT('h1)
	) name3757 (
		_w5262_,
		_w5264_,
		_w5265_
	);
	LUT2 #(
		.INIT('h8)
	) name3758 (
		\TM0_pad ,
		\_2332__reg/NET0131 ,
		_w5266_
	);
	LUT2 #(
		.INIT('h2)
	) name3759 (
		\TM1_pad ,
		\WX10989_reg/NET0131 ,
		_w5267_
	);
	LUT2 #(
		.INIT('h4)
	) name3760 (
		\TM1_pad ,
		\WX10989_reg/NET0131 ,
		_w5268_
	);
	LUT2 #(
		.INIT('h1)
	) name3761 (
		_w5267_,
		_w5268_,
		_w5269_
	);
	LUT2 #(
		.INIT('h1)
	) name3762 (
		\WX11053_reg/NET0131 ,
		_w5269_,
		_w5270_
	);
	LUT2 #(
		.INIT('h8)
	) name3763 (
		\WX11053_reg/NET0131 ,
		_w5269_,
		_w5271_
	);
	LUT2 #(
		.INIT('h1)
	) name3764 (
		_w5270_,
		_w5271_,
		_w5272_
	);
	LUT2 #(
		.INIT('h2)
	) name3765 (
		\WX11117_reg/NET0131 ,
		\WX11181_reg/NET0131 ,
		_w5273_
	);
	LUT2 #(
		.INIT('h4)
	) name3766 (
		\WX11117_reg/NET0131 ,
		\WX11181_reg/NET0131 ,
		_w5274_
	);
	LUT2 #(
		.INIT('h1)
	) name3767 (
		_w5273_,
		_w5274_,
		_w5275_
	);
	LUT2 #(
		.INIT('h8)
	) name3768 (
		_w5272_,
		_w5275_,
		_w5276_
	);
	LUT2 #(
		.INIT('h1)
	) name3769 (
		_w5272_,
		_w5275_,
		_w5277_
	);
	LUT2 #(
		.INIT('h1)
	) name3770 (
		\TM0_pad ,
		_w5276_,
		_w5278_
	);
	LUT2 #(
		.INIT('h4)
	) name3771 (
		_w5277_,
		_w5278_,
		_w5279_
	);
	LUT2 #(
		.INIT('h1)
	) name3772 (
		_w5266_,
		_w5279_,
		_w5280_
	);
	LUT2 #(
		.INIT('h2)
	) name3773 (
		_w1976_,
		_w5280_,
		_w5281_
	);
	LUT2 #(
		.INIT('h1)
	) name3774 (
		_w1871_,
		_w5138_,
		_w5282_
	);
	LUT2 #(
		.INIT('h2)
	) name3775 (
		_w1973_,
		_w5282_,
		_w5283_
	);
	LUT2 #(
		.INIT('h1)
	) name3776 (
		_w5281_,
		_w5283_,
		_w5284_
	);
	LUT2 #(
		.INIT('h8)
	) name3777 (
		\TM0_pad ,
		\_2200__reg/NET0131 ,
		_w5285_
	);
	LUT2 #(
		.INIT('h2)
	) name3778 (
		\WX5953_reg/NET0131 ,
		\WX6017_reg/NET0131 ,
		_w5286_
	);
	LUT2 #(
		.INIT('h4)
	) name3779 (
		\WX5953_reg/NET0131 ,
		\WX6017_reg/NET0131 ,
		_w5287_
	);
	LUT2 #(
		.INIT('h1)
	) name3780 (
		_w5286_,
		_w5287_,
		_w5288_
	);
	LUT2 #(
		.INIT('h2)
	) name3781 (
		\WX5889_reg/NET0131 ,
		_w5288_,
		_w5289_
	);
	LUT2 #(
		.INIT('h4)
	) name3782 (
		\WX5889_reg/NET0131 ,
		_w5288_,
		_w5290_
	);
	LUT2 #(
		.INIT('h1)
	) name3783 (
		_w5289_,
		_w5290_,
		_w5291_
	);
	LUT2 #(
		.INIT('h2)
	) name3784 (
		\TM1_pad ,
		\WX5825_reg/NET0131 ,
		_w5292_
	);
	LUT2 #(
		.INIT('h4)
	) name3785 (
		\TM1_pad ,
		\WX5825_reg/NET0131 ,
		_w5293_
	);
	LUT2 #(
		.INIT('h1)
	) name3786 (
		_w5292_,
		_w5293_,
		_w5294_
	);
	LUT2 #(
		.INIT('h4)
	) name3787 (
		_w5291_,
		_w5294_,
		_w5295_
	);
	LUT2 #(
		.INIT('h2)
	) name3788 (
		_w5291_,
		_w5294_,
		_w5296_
	);
	LUT2 #(
		.INIT('h1)
	) name3789 (
		\TM0_pad ,
		_w5295_,
		_w5297_
	);
	LUT2 #(
		.INIT('h4)
	) name3790 (
		_w5296_,
		_w5297_,
		_w5298_
	);
	LUT2 #(
		.INIT('h1)
	) name3791 (
		_w5285_,
		_w5298_,
		_w5299_
	);
	LUT2 #(
		.INIT('h2)
	) name3792 (
		_w1976_,
		_w5299_,
		_w5300_
	);
	LUT2 #(
		.INIT('h1)
	) name3793 (
		_w1794_,
		_w5234_,
		_w5301_
	);
	LUT2 #(
		.INIT('h2)
	) name3794 (
		_w1973_,
		_w5301_,
		_w5302_
	);
	LUT2 #(
		.INIT('h1)
	) name3795 (
		_w5300_,
		_w5302_,
		_w5303_
	);
	LUT2 #(
		.INIT('h8)
	) name3796 (
		\TM0_pad ,
		\_2233__reg/NET0131 ,
		_w5304_
	);
	LUT2 #(
		.INIT('h2)
	) name3797 (
		\WX7244_reg/NET0131 ,
		\WX7308_reg/NET0131 ,
		_w5305_
	);
	LUT2 #(
		.INIT('h4)
	) name3798 (
		\WX7244_reg/NET0131 ,
		\WX7308_reg/NET0131 ,
		_w5306_
	);
	LUT2 #(
		.INIT('h1)
	) name3799 (
		_w5305_,
		_w5306_,
		_w5307_
	);
	LUT2 #(
		.INIT('h2)
	) name3800 (
		\WX7180_reg/NET0131 ,
		_w5307_,
		_w5308_
	);
	LUT2 #(
		.INIT('h4)
	) name3801 (
		\WX7180_reg/NET0131 ,
		_w5307_,
		_w5309_
	);
	LUT2 #(
		.INIT('h1)
	) name3802 (
		_w5308_,
		_w5309_,
		_w5310_
	);
	LUT2 #(
		.INIT('h2)
	) name3803 (
		\TM1_pad ,
		\WX7116_reg/NET0131 ,
		_w5311_
	);
	LUT2 #(
		.INIT('h4)
	) name3804 (
		\TM1_pad ,
		\WX7116_reg/NET0131 ,
		_w5312_
	);
	LUT2 #(
		.INIT('h1)
	) name3805 (
		_w5311_,
		_w5312_,
		_w5313_
	);
	LUT2 #(
		.INIT('h4)
	) name3806 (
		_w5310_,
		_w5313_,
		_w5314_
	);
	LUT2 #(
		.INIT('h2)
	) name3807 (
		_w5310_,
		_w5313_,
		_w5315_
	);
	LUT2 #(
		.INIT('h1)
	) name3808 (
		\TM0_pad ,
		_w5314_,
		_w5316_
	);
	LUT2 #(
		.INIT('h4)
	) name3809 (
		_w5315_,
		_w5316_,
		_w5317_
	);
	LUT2 #(
		.INIT('h1)
	) name3810 (
		_w5304_,
		_w5317_,
		_w5318_
	);
	LUT2 #(
		.INIT('h2)
	) name3811 (
		_w1976_,
		_w5318_,
		_w5319_
	);
	LUT2 #(
		.INIT('h1)
	) name3812 (
		_w1810_,
		_w5157_,
		_w5320_
	);
	LUT2 #(
		.INIT('h2)
	) name3813 (
		_w1973_,
		_w5320_,
		_w5321_
	);
	LUT2 #(
		.INIT('h1)
	) name3814 (
		_w5319_,
		_w5321_,
		_w5322_
	);
	LUT2 #(
		.INIT('h2)
	) name3815 (
		\WX2110_reg/NET0131 ,
		\WX2174_reg/NET0131 ,
		_w5323_
	);
	LUT2 #(
		.INIT('h4)
	) name3816 (
		\WX2110_reg/NET0131 ,
		\WX2174_reg/NET0131 ,
		_w5324_
	);
	LUT2 #(
		.INIT('h1)
	) name3817 (
		_w5323_,
		_w5324_,
		_w5325_
	);
	LUT2 #(
		.INIT('h2)
	) name3818 (
		\WX1982_reg/NET0131 ,
		\WX2046_reg/NET0131 ,
		_w5326_
	);
	LUT2 #(
		.INIT('h4)
	) name3819 (
		\WX1982_reg/NET0131 ,
		\WX2046_reg/NET0131 ,
		_w5327_
	);
	LUT2 #(
		.INIT('h1)
	) name3820 (
		_w5326_,
		_w5327_,
		_w5328_
	);
	LUT2 #(
		.INIT('h4)
	) name3821 (
		_w5325_,
		_w5328_,
		_w5329_
	);
	LUT2 #(
		.INIT('h2)
	) name3822 (
		_w5325_,
		_w5328_,
		_w5330_
	);
	LUT2 #(
		.INIT('h1)
	) name3823 (
		\TM0_pad ,
		_w5329_,
		_w5331_
	);
	LUT2 #(
		.INIT('h4)
	) name3824 (
		_w5330_,
		_w5331_,
		_w5332_
	);
	LUT2 #(
		.INIT('h2)
	) name3825 (
		_w3172_,
		_w5332_,
		_w5333_
	);
	LUT2 #(
		.INIT('h2)
	) name3826 (
		\TM0_pad ,
		\_2118__reg/NET0131 ,
		_w5334_
	);
	LUT2 #(
		.INIT('h2)
	) name3827 (
		_w1976_,
		_w5334_,
		_w5335_
	);
	LUT2 #(
		.INIT('h4)
	) name3828 (
		_w3182_,
		_w5335_,
		_w5336_
	);
	LUT2 #(
		.INIT('h1)
	) name3829 (
		_w5333_,
		_w5336_,
		_w5337_
	);
	LUT2 #(
		.INIT('h8)
	) name3830 (
		\TM0_pad ,
		\_2266__reg/NET0131 ,
		_w5338_
	);
	LUT2 #(
		.INIT('h2)
	) name3831 (
		\WX8535_reg/NET0131 ,
		\WX8599_reg/NET0131 ,
		_w5339_
	);
	LUT2 #(
		.INIT('h4)
	) name3832 (
		\WX8535_reg/NET0131 ,
		\WX8599_reg/NET0131 ,
		_w5340_
	);
	LUT2 #(
		.INIT('h1)
	) name3833 (
		_w5339_,
		_w5340_,
		_w5341_
	);
	LUT2 #(
		.INIT('h2)
	) name3834 (
		\WX8471_reg/NET0131 ,
		_w5341_,
		_w5342_
	);
	LUT2 #(
		.INIT('h4)
	) name3835 (
		\WX8471_reg/NET0131 ,
		_w5341_,
		_w5343_
	);
	LUT2 #(
		.INIT('h1)
	) name3836 (
		_w5342_,
		_w5343_,
		_w5344_
	);
	LUT2 #(
		.INIT('h2)
	) name3837 (
		\TM1_pad ,
		\WX8407_reg/NET0131 ,
		_w5345_
	);
	LUT2 #(
		.INIT('h4)
	) name3838 (
		\TM1_pad ,
		\WX8407_reg/NET0131 ,
		_w5346_
	);
	LUT2 #(
		.INIT('h1)
	) name3839 (
		_w5345_,
		_w5346_,
		_w5347_
	);
	LUT2 #(
		.INIT('h4)
	) name3840 (
		_w5344_,
		_w5347_,
		_w5348_
	);
	LUT2 #(
		.INIT('h2)
	) name3841 (
		_w5344_,
		_w5347_,
		_w5349_
	);
	LUT2 #(
		.INIT('h1)
	) name3842 (
		\TM0_pad ,
		_w5348_,
		_w5350_
	);
	LUT2 #(
		.INIT('h4)
	) name3843 (
		_w5349_,
		_w5350_,
		_w5351_
	);
	LUT2 #(
		.INIT('h1)
	) name3844 (
		_w5338_,
		_w5351_,
		_w5352_
	);
	LUT2 #(
		.INIT('h2)
	) name3845 (
		_w1976_,
		_w5352_,
		_w5353_
	);
	LUT2 #(
		.INIT('h1)
	) name3846 (
		_w1826_,
		_w5191_,
		_w5354_
	);
	LUT2 #(
		.INIT('h2)
	) name3847 (
		_w1973_,
		_w5354_,
		_w5355_
	);
	LUT2 #(
		.INIT('h1)
	) name3848 (
		_w5353_,
		_w5355_,
		_w5356_
	);
	LUT2 #(
		.INIT('h8)
	) name3849 (
		\TM0_pad ,
		\_2167__reg/NET0131 ,
		_w5357_
	);
	LUT2 #(
		.INIT('h2)
	) name3850 (
		\WX4662_reg/NET0131 ,
		\WX4726_reg/NET0131 ,
		_w5358_
	);
	LUT2 #(
		.INIT('h4)
	) name3851 (
		\WX4662_reg/NET0131 ,
		\WX4726_reg/NET0131 ,
		_w5359_
	);
	LUT2 #(
		.INIT('h1)
	) name3852 (
		_w5358_,
		_w5359_,
		_w5360_
	);
	LUT2 #(
		.INIT('h2)
	) name3853 (
		\WX4598_reg/NET0131 ,
		_w5360_,
		_w5361_
	);
	LUT2 #(
		.INIT('h4)
	) name3854 (
		\WX4598_reg/NET0131 ,
		_w5360_,
		_w5362_
	);
	LUT2 #(
		.INIT('h1)
	) name3855 (
		_w5361_,
		_w5362_,
		_w5363_
	);
	LUT2 #(
		.INIT('h2)
	) name3856 (
		\TM1_pad ,
		\WX4534_reg/NET0131 ,
		_w5364_
	);
	LUT2 #(
		.INIT('h4)
	) name3857 (
		\TM1_pad ,
		\WX4534_reg/NET0131 ,
		_w5365_
	);
	LUT2 #(
		.INIT('h1)
	) name3858 (
		_w5364_,
		_w5365_,
		_w5366_
	);
	LUT2 #(
		.INIT('h4)
	) name3859 (
		_w5363_,
		_w5366_,
		_w5367_
	);
	LUT2 #(
		.INIT('h2)
	) name3860 (
		_w5363_,
		_w5366_,
		_w5368_
	);
	LUT2 #(
		.INIT('h1)
	) name3861 (
		\TM0_pad ,
		_w5367_,
		_w5369_
	);
	LUT2 #(
		.INIT('h4)
	) name3862 (
		_w5368_,
		_w5369_,
		_w5370_
	);
	LUT2 #(
		.INIT('h1)
	) name3863 (
		_w5357_,
		_w5370_,
		_w5371_
	);
	LUT2 #(
		.INIT('h2)
	) name3864 (
		_w1976_,
		_w5371_,
		_w5372_
	);
	LUT2 #(
		.INIT('h1)
	) name3865 (
		_w1778_,
		_w2900_,
		_w5373_
	);
	LUT2 #(
		.INIT('h2)
	) name3866 (
		_w1973_,
		_w5373_,
		_w5374_
	);
	LUT2 #(
		.INIT('h1)
	) name3867 (
		_w5372_,
		_w5374_,
		_w5375_
	);
	LUT2 #(
		.INIT('h2)
	) name3868 (
		_w3172_,
		_w4005_,
		_w5376_
	);
	LUT2 #(
		.INIT('h1)
	) name3869 (
		\DATA_0_9_pad ,
		\TM0_pad ,
		_w5377_
	);
	LUT2 #(
		.INIT('h2)
	) name3870 (
		\TM0_pad ,
		\_2342__reg/NET0131 ,
		_w5378_
	);
	LUT2 #(
		.INIT('h2)
	) name3871 (
		_w1976_,
		_w5377_,
		_w5379_
	);
	LUT2 #(
		.INIT('h4)
	) name3872 (
		_w5378_,
		_w5379_,
		_w5380_
	);
	LUT2 #(
		.INIT('h1)
	) name3873 (
		_w5376_,
		_w5380_,
		_w5381_
	);
	LUT2 #(
		.INIT('h8)
	) name3874 (
		RESET_pad,
		\WX10871_reg/NET0131 ,
		_w5382_
	);
	LUT2 #(
		.INIT('h8)
	) name3875 (
		\TM0_pad ,
		\_2298__reg/NET0131 ,
		_w5383_
	);
	LUT2 #(
		.INIT('h2)
	) name3876 (
		\WX9828_reg/NET0131 ,
		\WX9892_reg/NET0131 ,
		_w5384_
	);
	LUT2 #(
		.INIT('h4)
	) name3877 (
		\WX9828_reg/NET0131 ,
		\WX9892_reg/NET0131 ,
		_w5385_
	);
	LUT2 #(
		.INIT('h1)
	) name3878 (
		_w5384_,
		_w5385_,
		_w5386_
	);
	LUT2 #(
		.INIT('h2)
	) name3879 (
		\WX9764_reg/NET0131 ,
		_w5386_,
		_w5387_
	);
	LUT2 #(
		.INIT('h4)
	) name3880 (
		\WX9764_reg/NET0131 ,
		_w5386_,
		_w5388_
	);
	LUT2 #(
		.INIT('h1)
	) name3881 (
		_w5387_,
		_w5388_,
		_w5389_
	);
	LUT2 #(
		.INIT('h2)
	) name3882 (
		\TM1_pad ,
		\WX9700_reg/NET0131 ,
		_w5390_
	);
	LUT2 #(
		.INIT('h4)
	) name3883 (
		\TM1_pad ,
		\WX9700_reg/NET0131 ,
		_w5391_
	);
	LUT2 #(
		.INIT('h1)
	) name3884 (
		_w5390_,
		_w5391_,
		_w5392_
	);
	LUT2 #(
		.INIT('h4)
	) name3885 (
		_w5389_,
		_w5392_,
		_w5393_
	);
	LUT2 #(
		.INIT('h2)
	) name3886 (
		_w5389_,
		_w5392_,
		_w5394_
	);
	LUT2 #(
		.INIT('h1)
	) name3887 (
		\TM0_pad ,
		_w5393_,
		_w5395_
	);
	LUT2 #(
		.INIT('h4)
	) name3888 (
		_w5394_,
		_w5395_,
		_w5396_
	);
	LUT2 #(
		.INIT('h1)
	) name3889 (
		_w5383_,
		_w5396_,
		_w5397_
	);
	LUT2 #(
		.INIT('h2)
	) name3890 (
		_w1976_,
		_w5397_,
		_w5398_
	);
	LUT2 #(
		.INIT('h1)
	) name3891 (
		_w1826_,
		_w5351_,
		_w5399_
	);
	LUT2 #(
		.INIT('h2)
	) name3892 (
		_w1973_,
		_w5399_,
		_w5400_
	);
	LUT2 #(
		.INIT('h1)
	) name3893 (
		_w5398_,
		_w5400_,
		_w5401_
	);
	LUT2 #(
		.INIT('h8)
	) name3894 (
		\TM0_pad ,
		\_2331__reg/NET0131 ,
		_w5402_
	);
	LUT2 #(
		.INIT('h1)
	) name3895 (
		_w2333_,
		_w5402_,
		_w5403_
	);
	LUT2 #(
		.INIT('h2)
	) name3896 (
		_w1976_,
		_w5403_,
		_w5404_
	);
	LUT2 #(
		.INIT('h1)
	) name3897 (
		_w1855_,
		_w5260_,
		_w5405_
	);
	LUT2 #(
		.INIT('h2)
	) name3898 (
		_w1973_,
		_w5405_,
		_w5406_
	);
	LUT2 #(
		.INIT('h1)
	) name3899 (
		_w5404_,
		_w5406_,
		_w5407_
	);
	LUT2 #(
		.INIT('h8)
	) name3900 (
		\TM0_pad ,
		\_2199__reg/NET0131 ,
		_w5408_
	);
	LUT2 #(
		.INIT('h2)
	) name3901 (
		\WX5955_reg/NET0131 ,
		\WX6019_reg/NET0131 ,
		_w5409_
	);
	LUT2 #(
		.INIT('h4)
	) name3902 (
		\WX5955_reg/NET0131 ,
		\WX6019_reg/NET0131 ,
		_w5410_
	);
	LUT2 #(
		.INIT('h1)
	) name3903 (
		_w5409_,
		_w5410_,
		_w5411_
	);
	LUT2 #(
		.INIT('h2)
	) name3904 (
		\WX5891_reg/NET0131 ,
		_w5411_,
		_w5412_
	);
	LUT2 #(
		.INIT('h4)
	) name3905 (
		\WX5891_reg/NET0131 ,
		_w5411_,
		_w5413_
	);
	LUT2 #(
		.INIT('h1)
	) name3906 (
		_w5412_,
		_w5413_,
		_w5414_
	);
	LUT2 #(
		.INIT('h2)
	) name3907 (
		\TM1_pad ,
		\WX5827_reg/NET0131 ,
		_w5415_
	);
	LUT2 #(
		.INIT('h4)
	) name3908 (
		\TM1_pad ,
		\WX5827_reg/NET0131 ,
		_w5416_
	);
	LUT2 #(
		.INIT('h1)
	) name3909 (
		_w5415_,
		_w5416_,
		_w5417_
	);
	LUT2 #(
		.INIT('h4)
	) name3910 (
		_w5414_,
		_w5417_,
		_w5418_
	);
	LUT2 #(
		.INIT('h2)
	) name3911 (
		_w5414_,
		_w5417_,
		_w5419_
	);
	LUT2 #(
		.INIT('h1)
	) name3912 (
		\TM0_pad ,
		_w5418_,
		_w5420_
	);
	LUT2 #(
		.INIT('h4)
	) name3913 (
		_w5419_,
		_w5420_,
		_w5421_
	);
	LUT2 #(
		.INIT('h1)
	) name3914 (
		_w5408_,
		_w5421_,
		_w5422_
	);
	LUT2 #(
		.INIT('h2)
	) name3915 (
		_w1976_,
		_w5422_,
		_w5423_
	);
	LUT2 #(
		.INIT('h1)
	) name3916 (
		_w1778_,
		_w5370_,
		_w5424_
	);
	LUT2 #(
		.INIT('h2)
	) name3917 (
		_w1973_,
		_w5424_,
		_w5425_
	);
	LUT2 #(
		.INIT('h1)
	) name3918 (
		_w5423_,
		_w5425_,
		_w5426_
	);
	LUT2 #(
		.INIT('h8)
	) name3919 (
		\TM0_pad ,
		\_2232__reg/NET0131 ,
		_w5427_
	);
	LUT2 #(
		.INIT('h2)
	) name3920 (
		\WX7246_reg/NET0131 ,
		\WX7310_reg/NET0131 ,
		_w5428_
	);
	LUT2 #(
		.INIT('h4)
	) name3921 (
		\WX7246_reg/NET0131 ,
		\WX7310_reg/NET0131 ,
		_w5429_
	);
	LUT2 #(
		.INIT('h1)
	) name3922 (
		_w5428_,
		_w5429_,
		_w5430_
	);
	LUT2 #(
		.INIT('h2)
	) name3923 (
		\WX7182_reg/NET0131 ,
		_w5430_,
		_w5431_
	);
	LUT2 #(
		.INIT('h4)
	) name3924 (
		\WX7182_reg/NET0131 ,
		_w5430_,
		_w5432_
	);
	LUT2 #(
		.INIT('h1)
	) name3925 (
		_w5431_,
		_w5432_,
		_w5433_
	);
	LUT2 #(
		.INIT('h2)
	) name3926 (
		\TM1_pad ,
		\WX7118_reg/NET0131 ,
		_w5434_
	);
	LUT2 #(
		.INIT('h4)
	) name3927 (
		\TM1_pad ,
		\WX7118_reg/NET0131 ,
		_w5435_
	);
	LUT2 #(
		.INIT('h1)
	) name3928 (
		_w5434_,
		_w5435_,
		_w5436_
	);
	LUT2 #(
		.INIT('h4)
	) name3929 (
		_w5433_,
		_w5436_,
		_w5437_
	);
	LUT2 #(
		.INIT('h2)
	) name3930 (
		_w5433_,
		_w5436_,
		_w5438_
	);
	LUT2 #(
		.INIT('h1)
	) name3931 (
		\TM0_pad ,
		_w5437_,
		_w5439_
	);
	LUT2 #(
		.INIT('h4)
	) name3932 (
		_w5438_,
		_w5439_,
		_w5440_
	);
	LUT2 #(
		.INIT('h1)
	) name3933 (
		_w5427_,
		_w5440_,
		_w5441_
	);
	LUT2 #(
		.INIT('h2)
	) name3934 (
		_w1976_,
		_w5441_,
		_w5442_
	);
	LUT2 #(
		.INIT('h1)
	) name3935 (
		_w1794_,
		_w5298_,
		_w5443_
	);
	LUT2 #(
		.INIT('h2)
	) name3936 (
		_w1973_,
		_w5443_,
		_w5444_
	);
	LUT2 #(
		.INIT('h1)
	) name3937 (
		_w5442_,
		_w5444_,
		_w5445_
	);
	LUT2 #(
		.INIT('h2)
	) name3938 (
		\WX2112_reg/NET0131 ,
		\WX2176_reg/NET0131 ,
		_w5446_
	);
	LUT2 #(
		.INIT('h4)
	) name3939 (
		\WX2112_reg/NET0131 ,
		\WX2176_reg/NET0131 ,
		_w5447_
	);
	LUT2 #(
		.INIT('h1)
	) name3940 (
		_w5446_,
		_w5447_,
		_w5448_
	);
	LUT2 #(
		.INIT('h2)
	) name3941 (
		\WX1984_reg/NET0131 ,
		\WX2048_reg/NET0131 ,
		_w5449_
	);
	LUT2 #(
		.INIT('h4)
	) name3942 (
		\WX1984_reg/NET0131 ,
		\WX2048_reg/NET0131 ,
		_w5450_
	);
	LUT2 #(
		.INIT('h1)
	) name3943 (
		_w5449_,
		_w5450_,
		_w5451_
	);
	LUT2 #(
		.INIT('h4)
	) name3944 (
		_w5448_,
		_w5451_,
		_w5452_
	);
	LUT2 #(
		.INIT('h2)
	) name3945 (
		_w5448_,
		_w5451_,
		_w5453_
	);
	LUT2 #(
		.INIT('h1)
	) name3946 (
		\TM0_pad ,
		_w5452_,
		_w5454_
	);
	LUT2 #(
		.INIT('h4)
	) name3947 (
		_w5453_,
		_w5454_,
		_w5455_
	);
	LUT2 #(
		.INIT('h2)
	) name3948 (
		_w2023_,
		_w5455_,
		_w5456_
	);
	LUT2 #(
		.INIT('h2)
	) name3949 (
		\TM0_pad ,
		\_2117__reg/NET0131 ,
		_w5457_
	);
	LUT2 #(
		.INIT('h2)
	) name3950 (
		_w1976_,
		_w5457_,
		_w5458_
	);
	LUT2 #(
		.INIT('h4)
	) name3951 (
		_w3342_,
		_w5458_,
		_w5459_
	);
	LUT2 #(
		.INIT('h1)
	) name3952 (
		_w5456_,
		_w5459_,
		_w5460_
	);
	LUT2 #(
		.INIT('h8)
	) name3953 (
		\TM0_pad ,
		\_2265__reg/NET0131 ,
		_w5461_
	);
	LUT2 #(
		.INIT('h2)
	) name3954 (
		\WX8537_reg/NET0131 ,
		\WX8601_reg/NET0131 ,
		_w5462_
	);
	LUT2 #(
		.INIT('h4)
	) name3955 (
		\WX8537_reg/NET0131 ,
		\WX8601_reg/NET0131 ,
		_w5463_
	);
	LUT2 #(
		.INIT('h1)
	) name3956 (
		_w5462_,
		_w5463_,
		_w5464_
	);
	LUT2 #(
		.INIT('h2)
	) name3957 (
		\WX8473_reg/NET0131 ,
		_w5464_,
		_w5465_
	);
	LUT2 #(
		.INIT('h4)
	) name3958 (
		\WX8473_reg/NET0131 ,
		_w5464_,
		_w5466_
	);
	LUT2 #(
		.INIT('h1)
	) name3959 (
		_w5465_,
		_w5466_,
		_w5467_
	);
	LUT2 #(
		.INIT('h2)
	) name3960 (
		\TM1_pad ,
		\WX8409_reg/NET0131 ,
		_w5468_
	);
	LUT2 #(
		.INIT('h4)
	) name3961 (
		\TM1_pad ,
		\WX8409_reg/NET0131 ,
		_w5469_
	);
	LUT2 #(
		.INIT('h1)
	) name3962 (
		_w5468_,
		_w5469_,
		_w5470_
	);
	LUT2 #(
		.INIT('h4)
	) name3963 (
		_w5467_,
		_w5470_,
		_w5471_
	);
	LUT2 #(
		.INIT('h2)
	) name3964 (
		_w5467_,
		_w5470_,
		_w5472_
	);
	LUT2 #(
		.INIT('h1)
	) name3965 (
		\TM0_pad ,
		_w5471_,
		_w5473_
	);
	LUT2 #(
		.INIT('h4)
	) name3966 (
		_w5472_,
		_w5473_,
		_w5474_
	);
	LUT2 #(
		.INIT('h1)
	) name3967 (
		_w5461_,
		_w5474_,
		_w5475_
	);
	LUT2 #(
		.INIT('h2)
	) name3968 (
		_w1976_,
		_w5475_,
		_w5476_
	);
	LUT2 #(
		.INIT('h1)
	) name3969 (
		_w1810_,
		_w5317_,
		_w5477_
	);
	LUT2 #(
		.INIT('h2)
	) name3970 (
		_w1973_,
		_w5477_,
		_w5478_
	);
	LUT2 #(
		.INIT('h1)
	) name3971 (
		_w5476_,
		_w5478_,
		_w5479_
	);
	LUT2 #(
		.INIT('h8)
	) name3972 (
		\TM0_pad ,
		\_2166__reg/NET0131 ,
		_w5480_
	);
	LUT2 #(
		.INIT('h2)
	) name3973 (
		\WX4664_reg/NET0131 ,
		\WX4728_reg/NET0131 ,
		_w5481_
	);
	LUT2 #(
		.INIT('h4)
	) name3974 (
		\WX4664_reg/NET0131 ,
		\WX4728_reg/NET0131 ,
		_w5482_
	);
	LUT2 #(
		.INIT('h1)
	) name3975 (
		_w5481_,
		_w5482_,
		_w5483_
	);
	LUT2 #(
		.INIT('h2)
	) name3976 (
		\WX4600_reg/NET0131 ,
		_w5483_,
		_w5484_
	);
	LUT2 #(
		.INIT('h4)
	) name3977 (
		\WX4600_reg/NET0131 ,
		_w5483_,
		_w5485_
	);
	LUT2 #(
		.INIT('h1)
	) name3978 (
		_w5484_,
		_w5485_,
		_w5486_
	);
	LUT2 #(
		.INIT('h2)
	) name3979 (
		\TM1_pad ,
		\WX4536_reg/NET0131 ,
		_w5487_
	);
	LUT2 #(
		.INIT('h4)
	) name3980 (
		\TM1_pad ,
		\WX4536_reg/NET0131 ,
		_w5488_
	);
	LUT2 #(
		.INIT('h1)
	) name3981 (
		_w5487_,
		_w5488_,
		_w5489_
	);
	LUT2 #(
		.INIT('h4)
	) name3982 (
		_w5486_,
		_w5489_,
		_w5490_
	);
	LUT2 #(
		.INIT('h2)
	) name3983 (
		_w5486_,
		_w5489_,
		_w5491_
	);
	LUT2 #(
		.INIT('h1)
	) name3984 (
		\TM0_pad ,
		_w5490_,
		_w5492_
	);
	LUT2 #(
		.INIT('h4)
	) name3985 (
		_w5491_,
		_w5492_,
		_w5493_
	);
	LUT2 #(
		.INIT('h1)
	) name3986 (
		_w5480_,
		_w5493_,
		_w5494_
	);
	LUT2 #(
		.INIT('h2)
	) name3987 (
		_w1976_,
		_w5494_,
		_w5495_
	);
	LUT2 #(
		.INIT('h1)
	) name3988 (
		_w1762_,
		_w3065_,
		_w5496_
	);
	LUT2 #(
		.INIT('h2)
	) name3989 (
		_w1973_,
		_w5496_,
		_w5497_
	);
	LUT2 #(
		.INIT('h1)
	) name3990 (
		_w5495_,
		_w5497_,
		_w5498_
	);
	LUT2 #(
		.INIT('h1)
	) name3991 (
		\TM0_pad ,
		_w1929_,
		_w5499_
	);
	LUT2 #(
		.INIT('h2)
	) name3992 (
		_w3644_,
		_w5499_,
		_w5500_
	);
	LUT2 #(
		.INIT('h2)
	) name3993 (
		\TM0_pad ,
		\_2083__reg/NET0131 ,
		_w5501_
	);
	LUT2 #(
		.INIT('h2)
	) name3994 (
		\WX2116_reg/NET0131 ,
		\WX2180_reg/NET0131 ,
		_w5502_
	);
	LUT2 #(
		.INIT('h4)
	) name3995 (
		\WX2116_reg/NET0131 ,
		\WX2180_reg/NET0131 ,
		_w5503_
	);
	LUT2 #(
		.INIT('h1)
	) name3996 (
		_w5502_,
		_w5503_,
		_w5504_
	);
	LUT2 #(
		.INIT('h2)
	) name3997 (
		\WX1988_reg/NET0131 ,
		\WX2052_reg/NET0131 ,
		_w5505_
	);
	LUT2 #(
		.INIT('h4)
	) name3998 (
		\WX1988_reg/NET0131 ,
		\WX2052_reg/NET0131 ,
		_w5506_
	);
	LUT2 #(
		.INIT('h1)
	) name3999 (
		_w5505_,
		_w5506_,
		_w5507_
	);
	LUT2 #(
		.INIT('h4)
	) name4000 (
		_w5504_,
		_w5507_,
		_w5508_
	);
	LUT2 #(
		.INIT('h2)
	) name4001 (
		_w5504_,
		_w5507_,
		_w5509_
	);
	LUT2 #(
		.INIT('h1)
	) name4002 (
		\TM0_pad ,
		_w5508_,
		_w5510_
	);
	LUT2 #(
		.INIT('h4)
	) name4003 (
		_w5509_,
		_w5510_,
		_w5511_
	);
	LUT2 #(
		.INIT('h2)
	) name4004 (
		_w1976_,
		_w5501_,
		_w5512_
	);
	LUT2 #(
		.INIT('h4)
	) name4005 (
		_w5511_,
		_w5512_,
		_w5513_
	);
	LUT2 #(
		.INIT('h1)
	) name4006 (
		_w5500_,
		_w5513_,
		_w5514_
	);
	LUT2 #(
		.INIT('h8)
	) name4007 (
		RESET_pad,
		\WX10873_reg/NET0131 ,
		_w5515_
	);
	LUT2 #(
		.INIT('h8)
	) name4008 (
		\TM0_pad ,
		\_2297__reg/NET0131 ,
		_w5516_
	);
	LUT2 #(
		.INIT('h1)
	) name4009 (
		_w2003_,
		_w5516_,
		_w5517_
	);
	LUT2 #(
		.INIT('h2)
	) name4010 (
		_w1976_,
		_w5517_,
		_w5518_
	);
	LUT2 #(
		.INIT('h1)
	) name4011 (
		_w1810_,
		_w5474_,
		_w5519_
	);
	LUT2 #(
		.INIT('h2)
	) name4012 (
		_w1973_,
		_w5519_,
		_w5520_
	);
	LUT2 #(
		.INIT('h1)
	) name4013 (
		_w5518_,
		_w5520_,
		_w5521_
	);
	LUT2 #(
		.INIT('h8)
	) name4014 (
		\TM0_pad ,
		\_2330__reg/NET0131 ,
		_w5522_
	);
	LUT2 #(
		.INIT('h1)
	) name4015 (
		_w2509_,
		_w5522_,
		_w5523_
	);
	LUT2 #(
		.INIT('h2)
	) name4016 (
		_w1976_,
		_w5523_,
		_w5524_
	);
	LUT2 #(
		.INIT('h1)
	) name4017 (
		_w1826_,
		_w5396_,
		_w5525_
	);
	LUT2 #(
		.INIT('h2)
	) name4018 (
		_w1973_,
		_w5525_,
		_w5526_
	);
	LUT2 #(
		.INIT('h1)
	) name4019 (
		_w5524_,
		_w5526_,
		_w5527_
	);
	LUT2 #(
		.INIT('h8)
	) name4020 (
		\TM0_pad ,
		\_2198__reg/NET0131 ,
		_w5528_
	);
	LUT2 #(
		.INIT('h2)
	) name4021 (
		\WX5957_reg/NET0131 ,
		\WX6021_reg/NET0131 ,
		_w5529_
	);
	LUT2 #(
		.INIT('h4)
	) name4022 (
		\WX5957_reg/NET0131 ,
		\WX6021_reg/NET0131 ,
		_w5530_
	);
	LUT2 #(
		.INIT('h1)
	) name4023 (
		_w5529_,
		_w5530_,
		_w5531_
	);
	LUT2 #(
		.INIT('h2)
	) name4024 (
		\WX5893_reg/NET0131 ,
		_w5531_,
		_w5532_
	);
	LUT2 #(
		.INIT('h4)
	) name4025 (
		\WX5893_reg/NET0131 ,
		_w5531_,
		_w5533_
	);
	LUT2 #(
		.INIT('h1)
	) name4026 (
		_w5532_,
		_w5533_,
		_w5534_
	);
	LUT2 #(
		.INIT('h2)
	) name4027 (
		\TM1_pad ,
		\WX5829_reg/NET0131 ,
		_w5535_
	);
	LUT2 #(
		.INIT('h4)
	) name4028 (
		\TM1_pad ,
		\WX5829_reg/NET0131 ,
		_w5536_
	);
	LUT2 #(
		.INIT('h1)
	) name4029 (
		_w5535_,
		_w5536_,
		_w5537_
	);
	LUT2 #(
		.INIT('h4)
	) name4030 (
		_w5534_,
		_w5537_,
		_w5538_
	);
	LUT2 #(
		.INIT('h2)
	) name4031 (
		_w5534_,
		_w5537_,
		_w5539_
	);
	LUT2 #(
		.INIT('h1)
	) name4032 (
		\TM0_pad ,
		_w5538_,
		_w5540_
	);
	LUT2 #(
		.INIT('h4)
	) name4033 (
		_w5539_,
		_w5540_,
		_w5541_
	);
	LUT2 #(
		.INIT('h1)
	) name4034 (
		_w5528_,
		_w5541_,
		_w5542_
	);
	LUT2 #(
		.INIT('h2)
	) name4035 (
		_w1976_,
		_w5542_,
		_w5543_
	);
	LUT2 #(
		.INIT('h1)
	) name4036 (
		_w1762_,
		_w5493_,
		_w5544_
	);
	LUT2 #(
		.INIT('h2)
	) name4037 (
		_w1973_,
		_w5544_,
		_w5545_
	);
	LUT2 #(
		.INIT('h1)
	) name4038 (
		_w5543_,
		_w5545_,
		_w5546_
	);
	LUT2 #(
		.INIT('h8)
	) name4039 (
		\TM0_pad ,
		\_2231__reg/NET0131 ,
		_w5547_
	);
	LUT2 #(
		.INIT('h2)
	) name4040 (
		\WX7248_reg/NET0131 ,
		\WX7312_reg/NET0131 ,
		_w5548_
	);
	LUT2 #(
		.INIT('h4)
	) name4041 (
		\WX7248_reg/NET0131 ,
		\WX7312_reg/NET0131 ,
		_w5549_
	);
	LUT2 #(
		.INIT('h1)
	) name4042 (
		_w5548_,
		_w5549_,
		_w5550_
	);
	LUT2 #(
		.INIT('h2)
	) name4043 (
		\WX7184_reg/NET0131 ,
		_w5550_,
		_w5551_
	);
	LUT2 #(
		.INIT('h4)
	) name4044 (
		\WX7184_reg/NET0131 ,
		_w5550_,
		_w5552_
	);
	LUT2 #(
		.INIT('h1)
	) name4045 (
		_w5551_,
		_w5552_,
		_w5553_
	);
	LUT2 #(
		.INIT('h2)
	) name4046 (
		\TM1_pad ,
		\WX7120_reg/NET0131 ,
		_w5554_
	);
	LUT2 #(
		.INIT('h4)
	) name4047 (
		\TM1_pad ,
		\WX7120_reg/NET0131 ,
		_w5555_
	);
	LUT2 #(
		.INIT('h1)
	) name4048 (
		_w5554_,
		_w5555_,
		_w5556_
	);
	LUT2 #(
		.INIT('h4)
	) name4049 (
		_w5553_,
		_w5556_,
		_w5557_
	);
	LUT2 #(
		.INIT('h2)
	) name4050 (
		_w5553_,
		_w5556_,
		_w5558_
	);
	LUT2 #(
		.INIT('h1)
	) name4051 (
		\TM0_pad ,
		_w5557_,
		_w5559_
	);
	LUT2 #(
		.INIT('h4)
	) name4052 (
		_w5558_,
		_w5559_,
		_w5560_
	);
	LUT2 #(
		.INIT('h1)
	) name4053 (
		_w5547_,
		_w5560_,
		_w5561_
	);
	LUT2 #(
		.INIT('h2)
	) name4054 (
		_w1976_,
		_w5561_,
		_w5562_
	);
	LUT2 #(
		.INIT('h1)
	) name4055 (
		_w1778_,
		_w5421_,
		_w5563_
	);
	LUT2 #(
		.INIT('h2)
	) name4056 (
		_w1973_,
		_w5563_,
		_w5564_
	);
	LUT2 #(
		.INIT('h1)
	) name4057 (
		_w5562_,
		_w5564_,
		_w5565_
	);
	LUT2 #(
		.INIT('h2)
	) name4058 (
		\WX2114_reg/NET0131 ,
		\WX2178_reg/NET0131 ,
		_w5566_
	);
	LUT2 #(
		.INIT('h4)
	) name4059 (
		\WX2114_reg/NET0131 ,
		\WX2178_reg/NET0131 ,
		_w5567_
	);
	LUT2 #(
		.INIT('h1)
	) name4060 (
		_w5566_,
		_w5567_,
		_w5568_
	);
	LUT2 #(
		.INIT('h2)
	) name4061 (
		\WX1986_reg/NET0131 ,
		\WX2050_reg/NET0131 ,
		_w5569_
	);
	LUT2 #(
		.INIT('h4)
	) name4062 (
		\WX1986_reg/NET0131 ,
		\WX2050_reg/NET0131 ,
		_w5570_
	);
	LUT2 #(
		.INIT('h1)
	) name4063 (
		_w5569_,
		_w5570_,
		_w5571_
	);
	LUT2 #(
		.INIT('h4)
	) name4064 (
		_w5568_,
		_w5571_,
		_w5572_
	);
	LUT2 #(
		.INIT('h2)
	) name4065 (
		_w5568_,
		_w5571_,
		_w5573_
	);
	LUT2 #(
		.INIT('h1)
	) name4066 (
		\TM0_pad ,
		_w5572_,
		_w5574_
	);
	LUT2 #(
		.INIT('h4)
	) name4067 (
		_w5573_,
		_w5574_,
		_w5575_
	);
	LUT2 #(
		.INIT('h2)
	) name4068 (
		_w3483_,
		_w5575_,
		_w5576_
	);
	LUT2 #(
		.INIT('h2)
	) name4069 (
		\TM0_pad ,
		\_2116__reg/NET0131 ,
		_w5577_
	);
	LUT2 #(
		.INIT('h2)
	) name4070 (
		_w1976_,
		_w5577_,
		_w5578_
	);
	LUT2 #(
		.INIT('h4)
	) name4071 (
		_w3493_,
		_w5578_,
		_w5579_
	);
	LUT2 #(
		.INIT('h1)
	) name4072 (
		_w5576_,
		_w5579_,
		_w5580_
	);
	LUT2 #(
		.INIT('h8)
	) name4073 (
		\TM0_pad ,
		\_2264__reg/NET0131 ,
		_w5581_
	);
	LUT2 #(
		.INIT('h2)
	) name4074 (
		\WX8539_reg/NET0131 ,
		\WX8603_reg/NET0131 ,
		_w5582_
	);
	LUT2 #(
		.INIT('h4)
	) name4075 (
		\WX8539_reg/NET0131 ,
		\WX8603_reg/NET0131 ,
		_w5583_
	);
	LUT2 #(
		.INIT('h1)
	) name4076 (
		_w5582_,
		_w5583_,
		_w5584_
	);
	LUT2 #(
		.INIT('h2)
	) name4077 (
		\WX8475_reg/NET0131 ,
		_w5584_,
		_w5585_
	);
	LUT2 #(
		.INIT('h4)
	) name4078 (
		\WX8475_reg/NET0131 ,
		_w5584_,
		_w5586_
	);
	LUT2 #(
		.INIT('h1)
	) name4079 (
		_w5585_,
		_w5586_,
		_w5587_
	);
	LUT2 #(
		.INIT('h2)
	) name4080 (
		\TM1_pad ,
		\WX8411_reg/NET0131 ,
		_w5588_
	);
	LUT2 #(
		.INIT('h4)
	) name4081 (
		\TM1_pad ,
		\WX8411_reg/NET0131 ,
		_w5589_
	);
	LUT2 #(
		.INIT('h1)
	) name4082 (
		_w5588_,
		_w5589_,
		_w5590_
	);
	LUT2 #(
		.INIT('h4)
	) name4083 (
		_w5587_,
		_w5590_,
		_w5591_
	);
	LUT2 #(
		.INIT('h2)
	) name4084 (
		_w5587_,
		_w5590_,
		_w5592_
	);
	LUT2 #(
		.INIT('h1)
	) name4085 (
		\TM0_pad ,
		_w5591_,
		_w5593_
	);
	LUT2 #(
		.INIT('h4)
	) name4086 (
		_w5592_,
		_w5593_,
		_w5594_
	);
	LUT2 #(
		.INIT('h1)
	) name4087 (
		_w5581_,
		_w5594_,
		_w5595_
	);
	LUT2 #(
		.INIT('h2)
	) name4088 (
		_w1976_,
		_w5595_,
		_w5596_
	);
	LUT2 #(
		.INIT('h1)
	) name4089 (
		_w1794_,
		_w5440_,
		_w5597_
	);
	LUT2 #(
		.INIT('h2)
	) name4090 (
		_w1973_,
		_w5597_,
		_w5598_
	);
	LUT2 #(
		.INIT('h1)
	) name4091 (
		_w5596_,
		_w5598_,
		_w5599_
	);
	LUT2 #(
		.INIT('h8)
	) name4092 (
		\TM0_pad ,
		\_2165__reg/NET0131 ,
		_w5600_
	);
	LUT2 #(
		.INIT('h2)
	) name4093 (
		\WX4666_reg/NET0131 ,
		\WX4730_reg/NET0131 ,
		_w5601_
	);
	LUT2 #(
		.INIT('h4)
	) name4094 (
		\WX4666_reg/NET0131 ,
		\WX4730_reg/NET0131 ,
		_w5602_
	);
	LUT2 #(
		.INIT('h1)
	) name4095 (
		_w5601_,
		_w5602_,
		_w5603_
	);
	LUT2 #(
		.INIT('h2)
	) name4096 (
		\WX4602_reg/NET0131 ,
		_w5603_,
		_w5604_
	);
	LUT2 #(
		.INIT('h4)
	) name4097 (
		\WX4602_reg/NET0131 ,
		_w5603_,
		_w5605_
	);
	LUT2 #(
		.INIT('h1)
	) name4098 (
		_w5604_,
		_w5605_,
		_w5606_
	);
	LUT2 #(
		.INIT('h2)
	) name4099 (
		\TM1_pad ,
		\WX4538_reg/NET0131 ,
		_w5607_
	);
	LUT2 #(
		.INIT('h4)
	) name4100 (
		\TM1_pad ,
		\WX4538_reg/NET0131 ,
		_w5608_
	);
	LUT2 #(
		.INIT('h1)
	) name4101 (
		_w5607_,
		_w5608_,
		_w5609_
	);
	LUT2 #(
		.INIT('h4)
	) name4102 (
		_w5606_,
		_w5609_,
		_w5610_
	);
	LUT2 #(
		.INIT('h2)
	) name4103 (
		_w5606_,
		_w5609_,
		_w5611_
	);
	LUT2 #(
		.INIT('h1)
	) name4104 (
		\TM0_pad ,
		_w5610_,
		_w5612_
	);
	LUT2 #(
		.INIT('h4)
	) name4105 (
		_w5611_,
		_w5612_,
		_w5613_
	);
	LUT2 #(
		.INIT('h1)
	) name4106 (
		_w5600_,
		_w5613_,
		_w5614_
	);
	LUT2 #(
		.INIT('h2)
	) name4107 (
		_w1976_,
		_w5614_,
		_w5615_
	);
	LUT2 #(
		.INIT('h1)
	) name4108 (
		_w1746_,
		_w3241_,
		_w5616_
	);
	LUT2 #(
		.INIT('h2)
	) name4109 (
		_w1973_,
		_w5616_,
		_w5617_
	);
	LUT2 #(
		.INIT('h1)
	) name4110 (
		_w5615_,
		_w5617_,
		_w5618_
	);
	LUT2 #(
		.INIT('h1)
	) name4111 (
		\TM0_pad ,
		_w1916_,
		_w5619_
	);
	LUT2 #(
		.INIT('h2)
	) name4112 (
		_w3805_,
		_w5619_,
		_w5620_
	);
	LUT2 #(
		.INIT('h2)
	) name4113 (
		\TM0_pad ,
		\_2082__reg/NET0131 ,
		_w5621_
	);
	LUT2 #(
		.INIT('h2)
	) name4114 (
		\WX2118_reg/NET0131 ,
		\WX2182_reg/NET0131 ,
		_w5622_
	);
	LUT2 #(
		.INIT('h4)
	) name4115 (
		\WX2118_reg/NET0131 ,
		\WX2182_reg/NET0131 ,
		_w5623_
	);
	LUT2 #(
		.INIT('h1)
	) name4116 (
		_w5622_,
		_w5623_,
		_w5624_
	);
	LUT2 #(
		.INIT('h2)
	) name4117 (
		\WX1990_reg/NET0131 ,
		\WX2054_reg/NET0131 ,
		_w5625_
	);
	LUT2 #(
		.INIT('h4)
	) name4118 (
		\WX1990_reg/NET0131 ,
		\WX2054_reg/NET0131 ,
		_w5626_
	);
	LUT2 #(
		.INIT('h1)
	) name4119 (
		_w5625_,
		_w5626_,
		_w5627_
	);
	LUT2 #(
		.INIT('h4)
	) name4120 (
		_w5624_,
		_w5627_,
		_w5628_
	);
	LUT2 #(
		.INIT('h2)
	) name4121 (
		_w5624_,
		_w5627_,
		_w5629_
	);
	LUT2 #(
		.INIT('h1)
	) name4122 (
		\TM0_pad ,
		_w5628_,
		_w5630_
	);
	LUT2 #(
		.INIT('h4)
	) name4123 (
		_w5629_,
		_w5630_,
		_w5631_
	);
	LUT2 #(
		.INIT('h2)
	) name4124 (
		_w1976_,
		_w5621_,
		_w5632_
	);
	LUT2 #(
		.INIT('h4)
	) name4125 (
		_w5631_,
		_w5632_,
		_w5633_
	);
	LUT2 #(
		.INIT('h1)
	) name4126 (
		_w5620_,
		_w5633_,
		_w5634_
	);
	LUT2 #(
		.INIT('h2)
	) name4127 (
		_w3483_,
		_w4291_,
		_w5635_
	);
	LUT2 #(
		.INIT('h1)
	) name4128 (
		\DATA_0_7_pad ,
		\TM0_pad ,
		_w5636_
	);
	LUT2 #(
		.INIT('h2)
	) name4129 (
		\TM0_pad ,
		\_2340__reg/NET0131 ,
		_w5637_
	);
	LUT2 #(
		.INIT('h2)
	) name4130 (
		_w1976_,
		_w5636_,
		_w5638_
	);
	LUT2 #(
		.INIT('h4)
	) name4131 (
		_w5637_,
		_w5638_,
		_w5639_
	);
	LUT2 #(
		.INIT('h1)
	) name4132 (
		_w5635_,
		_w5639_,
		_w5640_
	);
	LUT2 #(
		.INIT('h8)
	) name4133 (
		RESET_pad,
		\WX10875_reg/NET0131 ,
		_w5641_
	);
	LUT2 #(
		.INIT('h8)
	) name4134 (
		\TM0_pad ,
		\_2296__reg/NET0131 ,
		_w5642_
	);
	LUT2 #(
		.INIT('h2)
	) name4135 (
		\WX9832_reg/NET0131 ,
		\WX9896_reg/NET0131 ,
		_w5643_
	);
	LUT2 #(
		.INIT('h4)
	) name4136 (
		\WX9832_reg/NET0131 ,
		\WX9896_reg/NET0131 ,
		_w5644_
	);
	LUT2 #(
		.INIT('h1)
	) name4137 (
		_w5643_,
		_w5644_,
		_w5645_
	);
	LUT2 #(
		.INIT('h2)
	) name4138 (
		\WX9768_reg/NET0131 ,
		_w5645_,
		_w5646_
	);
	LUT2 #(
		.INIT('h4)
	) name4139 (
		\WX9768_reg/NET0131 ,
		_w5645_,
		_w5647_
	);
	LUT2 #(
		.INIT('h1)
	) name4140 (
		_w5646_,
		_w5647_,
		_w5648_
	);
	LUT2 #(
		.INIT('h2)
	) name4141 (
		\TM1_pad ,
		\WX9704_reg/NET0131 ,
		_w5649_
	);
	LUT2 #(
		.INIT('h4)
	) name4142 (
		\TM1_pad ,
		\WX9704_reg/NET0131 ,
		_w5650_
	);
	LUT2 #(
		.INIT('h1)
	) name4143 (
		_w5649_,
		_w5650_,
		_w5651_
	);
	LUT2 #(
		.INIT('h4)
	) name4144 (
		_w5648_,
		_w5651_,
		_w5652_
	);
	LUT2 #(
		.INIT('h2)
	) name4145 (
		_w5648_,
		_w5651_,
		_w5653_
	);
	LUT2 #(
		.INIT('h1)
	) name4146 (
		\TM0_pad ,
		_w5652_,
		_w5654_
	);
	LUT2 #(
		.INIT('h4)
	) name4147 (
		_w5653_,
		_w5654_,
		_w5655_
	);
	LUT2 #(
		.INIT('h1)
	) name4148 (
		_w5642_,
		_w5655_,
		_w5656_
	);
	LUT2 #(
		.INIT('h2)
	) name4149 (
		_w1976_,
		_w5656_,
		_w5657_
	);
	LUT2 #(
		.INIT('h1)
	) name4150 (
		_w1794_,
		_w5594_,
		_w5658_
	);
	LUT2 #(
		.INIT('h2)
	) name4151 (
		_w1973_,
		_w5658_,
		_w5659_
	);
	LUT2 #(
		.INIT('h1)
	) name4152 (
		_w5657_,
		_w5659_,
		_w5660_
	);
	LUT2 #(
		.INIT('h8)
	) name4153 (
		\TM0_pad ,
		\_2197__reg/NET0131 ,
		_w5661_
	);
	LUT2 #(
		.INIT('h2)
	) name4154 (
		\WX5959_reg/NET0131 ,
		\WX6023_reg/NET0131 ,
		_w5662_
	);
	LUT2 #(
		.INIT('h4)
	) name4155 (
		\WX5959_reg/NET0131 ,
		\WX6023_reg/NET0131 ,
		_w5663_
	);
	LUT2 #(
		.INIT('h1)
	) name4156 (
		_w5662_,
		_w5663_,
		_w5664_
	);
	LUT2 #(
		.INIT('h2)
	) name4157 (
		\WX5895_reg/NET0131 ,
		_w5664_,
		_w5665_
	);
	LUT2 #(
		.INIT('h4)
	) name4158 (
		\WX5895_reg/NET0131 ,
		_w5664_,
		_w5666_
	);
	LUT2 #(
		.INIT('h1)
	) name4159 (
		_w5665_,
		_w5666_,
		_w5667_
	);
	LUT2 #(
		.INIT('h2)
	) name4160 (
		\TM1_pad ,
		\WX5831_reg/NET0131 ,
		_w5668_
	);
	LUT2 #(
		.INIT('h4)
	) name4161 (
		\TM1_pad ,
		\WX5831_reg/NET0131 ,
		_w5669_
	);
	LUT2 #(
		.INIT('h1)
	) name4162 (
		_w5668_,
		_w5669_,
		_w5670_
	);
	LUT2 #(
		.INIT('h4)
	) name4163 (
		_w5667_,
		_w5670_,
		_w5671_
	);
	LUT2 #(
		.INIT('h2)
	) name4164 (
		_w5667_,
		_w5670_,
		_w5672_
	);
	LUT2 #(
		.INIT('h1)
	) name4165 (
		\TM0_pad ,
		_w5671_,
		_w5673_
	);
	LUT2 #(
		.INIT('h4)
	) name4166 (
		_w5672_,
		_w5673_,
		_w5674_
	);
	LUT2 #(
		.INIT('h1)
	) name4167 (
		_w5661_,
		_w5674_,
		_w5675_
	);
	LUT2 #(
		.INIT('h2)
	) name4168 (
		_w1976_,
		_w5675_,
		_w5676_
	);
	LUT2 #(
		.INIT('h1)
	) name4169 (
		_w1746_,
		_w5613_,
		_w5677_
	);
	LUT2 #(
		.INIT('h2)
	) name4170 (
		_w1973_,
		_w5677_,
		_w5678_
	);
	LUT2 #(
		.INIT('h1)
	) name4171 (
		_w5676_,
		_w5678_,
		_w5679_
	);
	LUT2 #(
		.INIT('h8)
	) name4172 (
		\TM0_pad ,
		\_2230__reg/NET0131 ,
		_w5680_
	);
	LUT2 #(
		.INIT('h2)
	) name4173 (
		\WX7250_reg/NET0131 ,
		\WX7314_reg/NET0131 ,
		_w5681_
	);
	LUT2 #(
		.INIT('h4)
	) name4174 (
		\WX7250_reg/NET0131 ,
		\WX7314_reg/NET0131 ,
		_w5682_
	);
	LUT2 #(
		.INIT('h1)
	) name4175 (
		_w5681_,
		_w5682_,
		_w5683_
	);
	LUT2 #(
		.INIT('h2)
	) name4176 (
		\WX7186_reg/NET0131 ,
		_w5683_,
		_w5684_
	);
	LUT2 #(
		.INIT('h4)
	) name4177 (
		\WX7186_reg/NET0131 ,
		_w5683_,
		_w5685_
	);
	LUT2 #(
		.INIT('h1)
	) name4178 (
		_w5684_,
		_w5685_,
		_w5686_
	);
	LUT2 #(
		.INIT('h2)
	) name4179 (
		\TM1_pad ,
		\WX7122_reg/NET0131 ,
		_w5687_
	);
	LUT2 #(
		.INIT('h4)
	) name4180 (
		\TM1_pad ,
		\WX7122_reg/NET0131 ,
		_w5688_
	);
	LUT2 #(
		.INIT('h1)
	) name4181 (
		_w5687_,
		_w5688_,
		_w5689_
	);
	LUT2 #(
		.INIT('h4)
	) name4182 (
		_w5686_,
		_w5689_,
		_w5690_
	);
	LUT2 #(
		.INIT('h2)
	) name4183 (
		_w5686_,
		_w5689_,
		_w5691_
	);
	LUT2 #(
		.INIT('h1)
	) name4184 (
		\TM0_pad ,
		_w5690_,
		_w5692_
	);
	LUT2 #(
		.INIT('h4)
	) name4185 (
		_w5691_,
		_w5692_,
		_w5693_
	);
	LUT2 #(
		.INIT('h1)
	) name4186 (
		_w5680_,
		_w5693_,
		_w5694_
	);
	LUT2 #(
		.INIT('h2)
	) name4187 (
		_w1976_,
		_w5694_,
		_w5695_
	);
	LUT2 #(
		.INIT('h1)
	) name4188 (
		_w1762_,
		_w5541_,
		_w5696_
	);
	LUT2 #(
		.INIT('h2)
	) name4189 (
		_w1973_,
		_w5696_,
		_w5697_
	);
	LUT2 #(
		.INIT('h1)
	) name4190 (
		_w5695_,
		_w5697_,
		_w5698_
	);
	LUT2 #(
		.INIT('h2)
	) name4191 (
		_w3644_,
		_w5511_,
		_w5699_
	);
	LUT2 #(
		.INIT('h2)
	) name4192 (
		\TM0_pad ,
		\_2115__reg/NET0131 ,
		_w5700_
	);
	LUT2 #(
		.INIT('h2)
	) name4193 (
		_w1976_,
		_w5700_,
		_w5701_
	);
	LUT2 #(
		.INIT('h4)
	) name4194 (
		_w3654_,
		_w5701_,
		_w5702_
	);
	LUT2 #(
		.INIT('h1)
	) name4195 (
		_w5699_,
		_w5702_,
		_w5703_
	);
	LUT2 #(
		.INIT('h8)
	) name4196 (
		\TM0_pad ,
		\_2263__reg/NET0131 ,
		_w5704_
	);
	LUT2 #(
		.INIT('h2)
	) name4197 (
		\WX8541_reg/NET0131 ,
		\WX8605_reg/NET0131 ,
		_w5705_
	);
	LUT2 #(
		.INIT('h4)
	) name4198 (
		\WX8541_reg/NET0131 ,
		\WX8605_reg/NET0131 ,
		_w5706_
	);
	LUT2 #(
		.INIT('h1)
	) name4199 (
		_w5705_,
		_w5706_,
		_w5707_
	);
	LUT2 #(
		.INIT('h2)
	) name4200 (
		\WX8477_reg/NET0131 ,
		_w5707_,
		_w5708_
	);
	LUT2 #(
		.INIT('h4)
	) name4201 (
		\WX8477_reg/NET0131 ,
		_w5707_,
		_w5709_
	);
	LUT2 #(
		.INIT('h1)
	) name4202 (
		_w5708_,
		_w5709_,
		_w5710_
	);
	LUT2 #(
		.INIT('h2)
	) name4203 (
		\TM1_pad ,
		\WX8413_reg/NET0131 ,
		_w5711_
	);
	LUT2 #(
		.INIT('h4)
	) name4204 (
		\TM1_pad ,
		\WX8413_reg/NET0131 ,
		_w5712_
	);
	LUT2 #(
		.INIT('h1)
	) name4205 (
		_w5711_,
		_w5712_,
		_w5713_
	);
	LUT2 #(
		.INIT('h4)
	) name4206 (
		_w5710_,
		_w5713_,
		_w5714_
	);
	LUT2 #(
		.INIT('h2)
	) name4207 (
		_w5710_,
		_w5713_,
		_w5715_
	);
	LUT2 #(
		.INIT('h1)
	) name4208 (
		\TM0_pad ,
		_w5714_,
		_w5716_
	);
	LUT2 #(
		.INIT('h4)
	) name4209 (
		_w5715_,
		_w5716_,
		_w5717_
	);
	LUT2 #(
		.INIT('h1)
	) name4210 (
		_w5704_,
		_w5717_,
		_w5718_
	);
	LUT2 #(
		.INIT('h2)
	) name4211 (
		_w1976_,
		_w5718_,
		_w5719_
	);
	LUT2 #(
		.INIT('h1)
	) name4212 (
		_w1778_,
		_w5560_,
		_w5720_
	);
	LUT2 #(
		.INIT('h2)
	) name4213 (
		_w1973_,
		_w5720_,
		_w5721_
	);
	LUT2 #(
		.INIT('h1)
	) name4214 (
		_w5719_,
		_w5721_,
		_w5722_
	);
	LUT2 #(
		.INIT('h8)
	) name4215 (
		\TM0_pad ,
		\_2164__reg/NET0131 ,
		_w5723_
	);
	LUT2 #(
		.INIT('h2)
	) name4216 (
		\WX4668_reg/NET0131 ,
		\WX4732_reg/NET0131 ,
		_w5724_
	);
	LUT2 #(
		.INIT('h4)
	) name4217 (
		\WX4668_reg/NET0131 ,
		\WX4732_reg/NET0131 ,
		_w5725_
	);
	LUT2 #(
		.INIT('h1)
	) name4218 (
		_w5724_,
		_w5725_,
		_w5726_
	);
	LUT2 #(
		.INIT('h2)
	) name4219 (
		\WX4604_reg/NET0131 ,
		_w5726_,
		_w5727_
	);
	LUT2 #(
		.INIT('h4)
	) name4220 (
		\WX4604_reg/NET0131 ,
		_w5726_,
		_w5728_
	);
	LUT2 #(
		.INIT('h1)
	) name4221 (
		_w5727_,
		_w5728_,
		_w5729_
	);
	LUT2 #(
		.INIT('h2)
	) name4222 (
		\TM1_pad ,
		\WX4540_reg/NET0131 ,
		_w5730_
	);
	LUT2 #(
		.INIT('h4)
	) name4223 (
		\TM1_pad ,
		\WX4540_reg/NET0131 ,
		_w5731_
	);
	LUT2 #(
		.INIT('h1)
	) name4224 (
		_w5730_,
		_w5731_,
		_w5732_
	);
	LUT2 #(
		.INIT('h4)
	) name4225 (
		_w5729_,
		_w5732_,
		_w5733_
	);
	LUT2 #(
		.INIT('h2)
	) name4226 (
		_w5729_,
		_w5732_,
		_w5734_
	);
	LUT2 #(
		.INIT('h1)
	) name4227 (
		\TM0_pad ,
		_w5733_,
		_w5735_
	);
	LUT2 #(
		.INIT('h4)
	) name4228 (
		_w5734_,
		_w5735_,
		_w5736_
	);
	LUT2 #(
		.INIT('h1)
	) name4229 (
		_w5723_,
		_w5736_,
		_w5737_
	);
	LUT2 #(
		.INIT('h2)
	) name4230 (
		_w1976_,
		_w5737_,
		_w5738_
	);
	LUT2 #(
		.INIT('h1)
	) name4231 (
		_w1730_,
		_w3391_,
		_w5739_
	);
	LUT2 #(
		.INIT('h2)
	) name4232 (
		_w1973_,
		_w5739_,
		_w5740_
	);
	LUT2 #(
		.INIT('h1)
	) name4233 (
		_w5738_,
		_w5740_,
		_w5741_
	);
	LUT2 #(
		.INIT('h1)
	) name4234 (
		\TM0_pad ,
		_w1880_,
		_w5742_
	);
	LUT2 #(
		.INIT('h1)
	) name4235 (
		_w1871_,
		_w5742_,
		_w5743_
	);
	LUT2 #(
		.INIT('h2)
	) name4236 (
		_w1973_,
		_w5743_,
		_w5744_
	);
	LUT2 #(
		.INIT('h8)
	) name4237 (
		\TM0_pad ,
		\_2108__reg/NET0131 ,
		_w5745_
	);
	LUT2 #(
		.INIT('h2)
	) name4238 (
		\TM1_pad ,
		\WX1938_reg/NET0131 ,
		_w5746_
	);
	LUT2 #(
		.INIT('h4)
	) name4239 (
		\TM1_pad ,
		\WX1938_reg/NET0131 ,
		_w5747_
	);
	LUT2 #(
		.INIT('h1)
	) name4240 (
		_w5746_,
		_w5747_,
		_w5748_
	);
	LUT2 #(
		.INIT('h1)
	) name4241 (
		\WX2002_reg/NET0131 ,
		_w5748_,
		_w5749_
	);
	LUT2 #(
		.INIT('h8)
	) name4242 (
		\WX2002_reg/NET0131 ,
		_w5748_,
		_w5750_
	);
	LUT2 #(
		.INIT('h1)
	) name4243 (
		_w5749_,
		_w5750_,
		_w5751_
	);
	LUT2 #(
		.INIT('h2)
	) name4244 (
		\WX2066_reg/NET0131 ,
		\WX2130_reg/NET0131 ,
		_w5752_
	);
	LUT2 #(
		.INIT('h4)
	) name4245 (
		\WX2066_reg/NET0131 ,
		\WX2130_reg/NET0131 ,
		_w5753_
	);
	LUT2 #(
		.INIT('h1)
	) name4246 (
		_w5752_,
		_w5753_,
		_w5754_
	);
	LUT2 #(
		.INIT('h8)
	) name4247 (
		_w5751_,
		_w5754_,
		_w5755_
	);
	LUT2 #(
		.INIT('h1)
	) name4248 (
		_w5751_,
		_w5754_,
		_w5756_
	);
	LUT2 #(
		.INIT('h1)
	) name4249 (
		\TM0_pad ,
		_w5755_,
		_w5757_
	);
	LUT2 #(
		.INIT('h4)
	) name4250 (
		_w5756_,
		_w5757_,
		_w5758_
	);
	LUT2 #(
		.INIT('h1)
	) name4251 (
		_w5745_,
		_w5758_,
		_w5759_
	);
	LUT2 #(
		.INIT('h2)
	) name4252 (
		_w1976_,
		_w5759_,
		_w5760_
	);
	LUT2 #(
		.INIT('h1)
	) name4253 (
		_w5744_,
		_w5760_,
		_w5761_
	);
	LUT2 #(
		.INIT('h2)
	) name4254 (
		_w3644_,
		_w4434_,
		_w5762_
	);
	LUT2 #(
		.INIT('h1)
	) name4255 (
		\DATA_0_6_pad ,
		\TM0_pad ,
		_w5763_
	);
	LUT2 #(
		.INIT('h2)
	) name4256 (
		\TM0_pad ,
		\_2339__reg/NET0131 ,
		_w5764_
	);
	LUT2 #(
		.INIT('h2)
	) name4257 (
		_w1976_,
		_w5763_,
		_w5765_
	);
	LUT2 #(
		.INIT('h4)
	) name4258 (
		_w5764_,
		_w5765_,
		_w5766_
	);
	LUT2 #(
		.INIT('h1)
	) name4259 (
		_w5762_,
		_w5766_,
		_w5767_
	);
	LUT2 #(
		.INIT('h8)
	) name4260 (
		RESET_pad,
		\WX10877_reg/NET0131 ,
		_w5768_
	);
	LUT2 #(
		.INIT('h8)
	) name4261 (
		\TM0_pad ,
		\_2163__reg/NET0131 ,
		_w5769_
	);
	LUT2 #(
		.INIT('h2)
	) name4262 (
		\WX4670_reg/NET0131 ,
		\WX4734_reg/NET0131 ,
		_w5770_
	);
	LUT2 #(
		.INIT('h4)
	) name4263 (
		\WX4670_reg/NET0131 ,
		\WX4734_reg/NET0131 ,
		_w5771_
	);
	LUT2 #(
		.INIT('h1)
	) name4264 (
		_w5770_,
		_w5771_,
		_w5772_
	);
	LUT2 #(
		.INIT('h2)
	) name4265 (
		\WX4606_reg/NET0131 ,
		_w5772_,
		_w5773_
	);
	LUT2 #(
		.INIT('h4)
	) name4266 (
		\WX4606_reg/NET0131 ,
		_w5772_,
		_w5774_
	);
	LUT2 #(
		.INIT('h1)
	) name4267 (
		_w5773_,
		_w5774_,
		_w5775_
	);
	LUT2 #(
		.INIT('h2)
	) name4268 (
		\TM1_pad ,
		\WX4542_reg/NET0131 ,
		_w5776_
	);
	LUT2 #(
		.INIT('h4)
	) name4269 (
		\TM1_pad ,
		\WX4542_reg/NET0131 ,
		_w5777_
	);
	LUT2 #(
		.INIT('h1)
	) name4270 (
		_w5776_,
		_w5777_,
		_w5778_
	);
	LUT2 #(
		.INIT('h4)
	) name4271 (
		_w5775_,
		_w5778_,
		_w5779_
	);
	LUT2 #(
		.INIT('h2)
	) name4272 (
		_w5775_,
		_w5778_,
		_w5780_
	);
	LUT2 #(
		.INIT('h1)
	) name4273 (
		\TM0_pad ,
		_w5779_,
		_w5781_
	);
	LUT2 #(
		.INIT('h4)
	) name4274 (
		_w5780_,
		_w5781_,
		_w5782_
	);
	LUT2 #(
		.INIT('h1)
	) name4275 (
		_w5769_,
		_w5782_,
		_w5783_
	);
	LUT2 #(
		.INIT('h2)
	) name4276 (
		_w1976_,
		_w5783_,
		_w5784_
	);
	LUT2 #(
		.INIT('h1)
	) name4277 (
		_w1714_,
		_w3552_,
		_w5785_
	);
	LUT2 #(
		.INIT('h2)
	) name4278 (
		_w1973_,
		_w5785_,
		_w5786_
	);
	LUT2 #(
		.INIT('h1)
	) name4279 (
		_w5784_,
		_w5786_,
		_w5787_
	);
	LUT2 #(
		.INIT('h8)
	) name4280 (
		\TM0_pad ,
		\_2295__reg/NET0131 ,
		_w5788_
	);
	LUT2 #(
		.INIT('h2)
	) name4281 (
		\WX9834_reg/NET0131 ,
		\WX9898_reg/NET0131 ,
		_w5789_
	);
	LUT2 #(
		.INIT('h4)
	) name4282 (
		\WX9834_reg/NET0131 ,
		\WX9898_reg/NET0131 ,
		_w5790_
	);
	LUT2 #(
		.INIT('h1)
	) name4283 (
		_w5789_,
		_w5790_,
		_w5791_
	);
	LUT2 #(
		.INIT('h2)
	) name4284 (
		\WX9770_reg/NET0131 ,
		_w5791_,
		_w5792_
	);
	LUT2 #(
		.INIT('h4)
	) name4285 (
		\WX9770_reg/NET0131 ,
		_w5791_,
		_w5793_
	);
	LUT2 #(
		.INIT('h1)
	) name4286 (
		_w5792_,
		_w5793_,
		_w5794_
	);
	LUT2 #(
		.INIT('h2)
	) name4287 (
		\TM1_pad ,
		\WX9706_reg/NET0131 ,
		_w5795_
	);
	LUT2 #(
		.INIT('h4)
	) name4288 (
		\TM1_pad ,
		\WX9706_reg/NET0131 ,
		_w5796_
	);
	LUT2 #(
		.INIT('h1)
	) name4289 (
		_w5795_,
		_w5796_,
		_w5797_
	);
	LUT2 #(
		.INIT('h4)
	) name4290 (
		_w5794_,
		_w5797_,
		_w5798_
	);
	LUT2 #(
		.INIT('h2)
	) name4291 (
		_w5794_,
		_w5797_,
		_w5799_
	);
	LUT2 #(
		.INIT('h1)
	) name4292 (
		\TM0_pad ,
		_w5798_,
		_w5800_
	);
	LUT2 #(
		.INIT('h4)
	) name4293 (
		_w5799_,
		_w5800_,
		_w5801_
	);
	LUT2 #(
		.INIT('h1)
	) name4294 (
		_w5788_,
		_w5801_,
		_w5802_
	);
	LUT2 #(
		.INIT('h2)
	) name4295 (
		_w1976_,
		_w5802_,
		_w5803_
	);
	LUT2 #(
		.INIT('h1)
	) name4296 (
		_w1778_,
		_w5717_,
		_w5804_
	);
	LUT2 #(
		.INIT('h2)
	) name4297 (
		_w1973_,
		_w5804_,
		_w5805_
	);
	LUT2 #(
		.INIT('h1)
	) name4298 (
		_w5803_,
		_w5805_,
		_w5806_
	);
	LUT2 #(
		.INIT('h8)
	) name4299 (
		\TM0_pad ,
		\_2328__reg/NET0131 ,
		_w5807_
	);
	LUT2 #(
		.INIT('h1)
	) name4300 (
		_w2837_,
		_w5807_,
		_w5808_
	);
	LUT2 #(
		.INIT('h2)
	) name4301 (
		_w1976_,
		_w5808_,
		_w5809_
	);
	LUT2 #(
		.INIT('h1)
	) name4302 (
		_w1794_,
		_w5655_,
		_w5810_
	);
	LUT2 #(
		.INIT('h2)
	) name4303 (
		_w1973_,
		_w5810_,
		_w5811_
	);
	LUT2 #(
		.INIT('h1)
	) name4304 (
		_w5809_,
		_w5811_,
		_w5812_
	);
	LUT2 #(
		.INIT('h8)
	) name4305 (
		\TM0_pad ,
		\_2196__reg/NET0131 ,
		_w5813_
	);
	LUT2 #(
		.INIT('h2)
	) name4306 (
		\WX5961_reg/NET0131 ,
		\WX6025_reg/NET0131 ,
		_w5814_
	);
	LUT2 #(
		.INIT('h4)
	) name4307 (
		\WX5961_reg/NET0131 ,
		\WX6025_reg/NET0131 ,
		_w5815_
	);
	LUT2 #(
		.INIT('h1)
	) name4308 (
		_w5814_,
		_w5815_,
		_w5816_
	);
	LUT2 #(
		.INIT('h2)
	) name4309 (
		\WX5897_reg/NET0131 ,
		_w5816_,
		_w5817_
	);
	LUT2 #(
		.INIT('h4)
	) name4310 (
		\WX5897_reg/NET0131 ,
		_w5816_,
		_w5818_
	);
	LUT2 #(
		.INIT('h1)
	) name4311 (
		_w5817_,
		_w5818_,
		_w5819_
	);
	LUT2 #(
		.INIT('h2)
	) name4312 (
		\TM1_pad ,
		\WX5833_reg/NET0131 ,
		_w5820_
	);
	LUT2 #(
		.INIT('h4)
	) name4313 (
		\TM1_pad ,
		\WX5833_reg/NET0131 ,
		_w5821_
	);
	LUT2 #(
		.INIT('h1)
	) name4314 (
		_w5820_,
		_w5821_,
		_w5822_
	);
	LUT2 #(
		.INIT('h4)
	) name4315 (
		_w5819_,
		_w5822_,
		_w5823_
	);
	LUT2 #(
		.INIT('h2)
	) name4316 (
		_w5819_,
		_w5822_,
		_w5824_
	);
	LUT2 #(
		.INIT('h1)
	) name4317 (
		\TM0_pad ,
		_w5823_,
		_w5825_
	);
	LUT2 #(
		.INIT('h4)
	) name4318 (
		_w5824_,
		_w5825_,
		_w5826_
	);
	LUT2 #(
		.INIT('h1)
	) name4319 (
		_w5813_,
		_w5826_,
		_w5827_
	);
	LUT2 #(
		.INIT('h2)
	) name4320 (
		_w1976_,
		_w5827_,
		_w5828_
	);
	LUT2 #(
		.INIT('h1)
	) name4321 (
		_w1730_,
		_w5736_,
		_w5829_
	);
	LUT2 #(
		.INIT('h2)
	) name4322 (
		_w1973_,
		_w5829_,
		_w5830_
	);
	LUT2 #(
		.INIT('h1)
	) name4323 (
		_w5828_,
		_w5830_,
		_w5831_
	);
	LUT2 #(
		.INIT('h8)
	) name4324 (
		\TM0_pad ,
		\_2229__reg/NET0131 ,
		_w5832_
	);
	LUT2 #(
		.INIT('h2)
	) name4325 (
		\WX7252_reg/NET0131 ,
		\WX7316_reg/NET0131 ,
		_w5833_
	);
	LUT2 #(
		.INIT('h4)
	) name4326 (
		\WX7252_reg/NET0131 ,
		\WX7316_reg/NET0131 ,
		_w5834_
	);
	LUT2 #(
		.INIT('h1)
	) name4327 (
		_w5833_,
		_w5834_,
		_w5835_
	);
	LUT2 #(
		.INIT('h2)
	) name4328 (
		\WX7188_reg/NET0131 ,
		_w5835_,
		_w5836_
	);
	LUT2 #(
		.INIT('h4)
	) name4329 (
		\WX7188_reg/NET0131 ,
		_w5835_,
		_w5837_
	);
	LUT2 #(
		.INIT('h1)
	) name4330 (
		_w5836_,
		_w5837_,
		_w5838_
	);
	LUT2 #(
		.INIT('h2)
	) name4331 (
		\TM1_pad ,
		\WX7124_reg/NET0131 ,
		_w5839_
	);
	LUT2 #(
		.INIT('h4)
	) name4332 (
		\TM1_pad ,
		\WX7124_reg/NET0131 ,
		_w5840_
	);
	LUT2 #(
		.INIT('h1)
	) name4333 (
		_w5839_,
		_w5840_,
		_w5841_
	);
	LUT2 #(
		.INIT('h4)
	) name4334 (
		_w5838_,
		_w5841_,
		_w5842_
	);
	LUT2 #(
		.INIT('h2)
	) name4335 (
		_w5838_,
		_w5841_,
		_w5843_
	);
	LUT2 #(
		.INIT('h1)
	) name4336 (
		\TM0_pad ,
		_w5842_,
		_w5844_
	);
	LUT2 #(
		.INIT('h4)
	) name4337 (
		_w5843_,
		_w5844_,
		_w5845_
	);
	LUT2 #(
		.INIT('h1)
	) name4338 (
		_w5832_,
		_w5845_,
		_w5846_
	);
	LUT2 #(
		.INIT('h2)
	) name4339 (
		_w1976_,
		_w5846_,
		_w5847_
	);
	LUT2 #(
		.INIT('h1)
	) name4340 (
		_w1746_,
		_w5674_,
		_w5848_
	);
	LUT2 #(
		.INIT('h2)
	) name4341 (
		_w1973_,
		_w5848_,
		_w5849_
	);
	LUT2 #(
		.INIT('h1)
	) name4342 (
		_w5847_,
		_w5849_,
		_w5850_
	);
	LUT2 #(
		.INIT('h2)
	) name4343 (
		_w3805_,
		_w5631_,
		_w5851_
	);
	LUT2 #(
		.INIT('h2)
	) name4344 (
		\TM0_pad ,
		\_2114__reg/NET0131 ,
		_w5852_
	);
	LUT2 #(
		.INIT('h2)
	) name4345 (
		_w1976_,
		_w5852_,
		_w5853_
	);
	LUT2 #(
		.INIT('h4)
	) name4346 (
		_w3815_,
		_w5853_,
		_w5854_
	);
	LUT2 #(
		.INIT('h1)
	) name4347 (
		_w5851_,
		_w5854_,
		_w5855_
	);
	LUT2 #(
		.INIT('h8)
	) name4348 (
		\TM0_pad ,
		\_2262__reg/NET0131 ,
		_w5856_
	);
	LUT2 #(
		.INIT('h2)
	) name4349 (
		\WX8543_reg/NET0131 ,
		\WX8607_reg/NET0131 ,
		_w5857_
	);
	LUT2 #(
		.INIT('h4)
	) name4350 (
		\WX8543_reg/NET0131 ,
		\WX8607_reg/NET0131 ,
		_w5858_
	);
	LUT2 #(
		.INIT('h1)
	) name4351 (
		_w5857_,
		_w5858_,
		_w5859_
	);
	LUT2 #(
		.INIT('h2)
	) name4352 (
		\WX8479_reg/NET0131 ,
		_w5859_,
		_w5860_
	);
	LUT2 #(
		.INIT('h4)
	) name4353 (
		\WX8479_reg/NET0131 ,
		_w5859_,
		_w5861_
	);
	LUT2 #(
		.INIT('h1)
	) name4354 (
		_w5860_,
		_w5861_,
		_w5862_
	);
	LUT2 #(
		.INIT('h2)
	) name4355 (
		\TM1_pad ,
		\WX8415_reg/NET0131 ,
		_w5863_
	);
	LUT2 #(
		.INIT('h4)
	) name4356 (
		\TM1_pad ,
		\WX8415_reg/NET0131 ,
		_w5864_
	);
	LUT2 #(
		.INIT('h1)
	) name4357 (
		_w5863_,
		_w5864_,
		_w5865_
	);
	LUT2 #(
		.INIT('h4)
	) name4358 (
		_w5862_,
		_w5865_,
		_w5866_
	);
	LUT2 #(
		.INIT('h2)
	) name4359 (
		_w5862_,
		_w5865_,
		_w5867_
	);
	LUT2 #(
		.INIT('h1)
	) name4360 (
		\TM0_pad ,
		_w5866_,
		_w5868_
	);
	LUT2 #(
		.INIT('h4)
	) name4361 (
		_w5867_,
		_w5868_,
		_w5869_
	);
	LUT2 #(
		.INIT('h1)
	) name4362 (
		_w5856_,
		_w5869_,
		_w5870_
	);
	LUT2 #(
		.INIT('h2)
	) name4363 (
		_w1976_,
		_w5870_,
		_w5871_
	);
	LUT2 #(
		.INIT('h1)
	) name4364 (
		_w1762_,
		_w5693_,
		_w5872_
	);
	LUT2 #(
		.INIT('h2)
	) name4365 (
		_w1973_,
		_w5872_,
		_w5873_
	);
	LUT2 #(
		.INIT('h1)
	) name4366 (
		_w5871_,
		_w5873_,
		_w5874_
	);
	LUT2 #(
		.INIT('h1)
	) name4367 (
		\TM0_pad ,
		_w1890_,
		_w5875_
	);
	LUT2 #(
		.INIT('h2)
	) name4368 (
		_w4101_,
		_w5875_,
		_w5876_
	);
	LUT2 #(
		.INIT('h2)
	) name4369 (
		\TM0_pad ,
		\_2080__reg/NET0131 ,
		_w5877_
	);
	LUT2 #(
		.INIT('h2)
	) name4370 (
		\WX2122_reg/NET0131 ,
		\WX2186_reg/NET0131 ,
		_w5878_
	);
	LUT2 #(
		.INIT('h4)
	) name4371 (
		\WX2122_reg/NET0131 ,
		\WX2186_reg/NET0131 ,
		_w5879_
	);
	LUT2 #(
		.INIT('h1)
	) name4372 (
		_w5878_,
		_w5879_,
		_w5880_
	);
	LUT2 #(
		.INIT('h2)
	) name4373 (
		\WX1994_reg/NET0131 ,
		\WX2058_reg/NET0131 ,
		_w5881_
	);
	LUT2 #(
		.INIT('h4)
	) name4374 (
		\WX1994_reg/NET0131 ,
		\WX2058_reg/NET0131 ,
		_w5882_
	);
	LUT2 #(
		.INIT('h1)
	) name4375 (
		_w5881_,
		_w5882_,
		_w5883_
	);
	LUT2 #(
		.INIT('h4)
	) name4376 (
		_w5880_,
		_w5883_,
		_w5884_
	);
	LUT2 #(
		.INIT('h2)
	) name4377 (
		_w5880_,
		_w5883_,
		_w5885_
	);
	LUT2 #(
		.INIT('h1)
	) name4378 (
		\TM0_pad ,
		_w5884_,
		_w5886_
	);
	LUT2 #(
		.INIT('h4)
	) name4379 (
		_w5885_,
		_w5886_,
		_w5887_
	);
	LUT2 #(
		.INIT('h2)
	) name4380 (
		_w1976_,
		_w5877_,
		_w5888_
	);
	LUT2 #(
		.INIT('h4)
	) name4381 (
		_w5887_,
		_w5888_,
		_w5889_
	);
	LUT2 #(
		.INIT('h1)
	) name4382 (
		_w5876_,
		_w5889_,
		_w5890_
	);
	LUT2 #(
		.INIT('h2)
	) name4383 (
		_w3805_,
		_w4562_,
		_w5891_
	);
	LUT2 #(
		.INIT('h1)
	) name4384 (
		\DATA_0_5_pad ,
		\TM0_pad ,
		_w5892_
	);
	LUT2 #(
		.INIT('h2)
	) name4385 (
		\TM0_pad ,
		\_2338__reg/NET0131 ,
		_w5893_
	);
	LUT2 #(
		.INIT('h2)
	) name4386 (
		_w1976_,
		_w5892_,
		_w5894_
	);
	LUT2 #(
		.INIT('h4)
	) name4387 (
		_w5893_,
		_w5894_,
		_w5895_
	);
	LUT2 #(
		.INIT('h1)
	) name4388 (
		_w5891_,
		_w5895_,
		_w5896_
	);
	LUT2 #(
		.INIT('h8)
	) name4389 (
		RESET_pad,
		\WX10879_reg/NET0131 ,
		_w5897_
	);
	LUT2 #(
		.INIT('h8)
	) name4390 (
		\TM0_pad ,
		\_2162__reg/NET0131 ,
		_w5898_
	);
	LUT2 #(
		.INIT('h2)
	) name4391 (
		\WX4672_reg/NET0131 ,
		\WX4736_reg/NET0131 ,
		_w5899_
	);
	LUT2 #(
		.INIT('h4)
	) name4392 (
		\WX4672_reg/NET0131 ,
		\WX4736_reg/NET0131 ,
		_w5900_
	);
	LUT2 #(
		.INIT('h1)
	) name4393 (
		_w5899_,
		_w5900_,
		_w5901_
	);
	LUT2 #(
		.INIT('h2)
	) name4394 (
		\WX4608_reg/NET0131 ,
		_w5901_,
		_w5902_
	);
	LUT2 #(
		.INIT('h4)
	) name4395 (
		\WX4608_reg/NET0131 ,
		_w5901_,
		_w5903_
	);
	LUT2 #(
		.INIT('h1)
	) name4396 (
		_w5902_,
		_w5903_,
		_w5904_
	);
	LUT2 #(
		.INIT('h2)
	) name4397 (
		\TM1_pad ,
		\WX4544_reg/NET0131 ,
		_w5905_
	);
	LUT2 #(
		.INIT('h4)
	) name4398 (
		\TM1_pad ,
		\WX4544_reg/NET0131 ,
		_w5906_
	);
	LUT2 #(
		.INIT('h1)
	) name4399 (
		_w5905_,
		_w5906_,
		_w5907_
	);
	LUT2 #(
		.INIT('h4)
	) name4400 (
		_w5904_,
		_w5907_,
		_w5908_
	);
	LUT2 #(
		.INIT('h2)
	) name4401 (
		_w5904_,
		_w5907_,
		_w5909_
	);
	LUT2 #(
		.INIT('h1)
	) name4402 (
		\TM0_pad ,
		_w5908_,
		_w5910_
	);
	LUT2 #(
		.INIT('h4)
	) name4403 (
		_w5909_,
		_w5910_,
		_w5911_
	);
	LUT2 #(
		.INIT('h1)
	) name4404 (
		_w5898_,
		_w5911_,
		_w5912_
	);
	LUT2 #(
		.INIT('h2)
	) name4405 (
		_w1976_,
		_w5912_,
		_w5913_
	);
	LUT2 #(
		.INIT('h1)
	) name4406 (
		_w1698_,
		_w3713_,
		_w5914_
	);
	LUT2 #(
		.INIT('h2)
	) name4407 (
		_w1973_,
		_w5914_,
		_w5915_
	);
	LUT2 #(
		.INIT('h1)
	) name4408 (
		_w5913_,
		_w5915_,
		_w5916_
	);
	LUT2 #(
		.INIT('h8)
	) name4409 (
		\TM0_pad ,
		\_2294__reg/NET0131 ,
		_w5917_
	);
	LUT2 #(
		.INIT('h2)
	) name4410 (
		\WX9836_reg/NET0131 ,
		\WX9900_reg/NET0131 ,
		_w5918_
	);
	LUT2 #(
		.INIT('h4)
	) name4411 (
		\WX9836_reg/NET0131 ,
		\WX9900_reg/NET0131 ,
		_w5919_
	);
	LUT2 #(
		.INIT('h1)
	) name4412 (
		_w5918_,
		_w5919_,
		_w5920_
	);
	LUT2 #(
		.INIT('h2)
	) name4413 (
		\WX9772_reg/NET0131 ,
		_w5920_,
		_w5921_
	);
	LUT2 #(
		.INIT('h4)
	) name4414 (
		\WX9772_reg/NET0131 ,
		_w5920_,
		_w5922_
	);
	LUT2 #(
		.INIT('h1)
	) name4415 (
		_w5921_,
		_w5922_,
		_w5923_
	);
	LUT2 #(
		.INIT('h2)
	) name4416 (
		\TM1_pad ,
		\WX9708_reg/NET0131 ,
		_w5924_
	);
	LUT2 #(
		.INIT('h4)
	) name4417 (
		\TM1_pad ,
		\WX9708_reg/NET0131 ,
		_w5925_
	);
	LUT2 #(
		.INIT('h1)
	) name4418 (
		_w5924_,
		_w5925_,
		_w5926_
	);
	LUT2 #(
		.INIT('h4)
	) name4419 (
		_w5923_,
		_w5926_,
		_w5927_
	);
	LUT2 #(
		.INIT('h2)
	) name4420 (
		_w5923_,
		_w5926_,
		_w5928_
	);
	LUT2 #(
		.INIT('h1)
	) name4421 (
		\TM0_pad ,
		_w5927_,
		_w5929_
	);
	LUT2 #(
		.INIT('h4)
	) name4422 (
		_w5928_,
		_w5929_,
		_w5930_
	);
	LUT2 #(
		.INIT('h1)
	) name4423 (
		_w5917_,
		_w5930_,
		_w5931_
	);
	LUT2 #(
		.INIT('h2)
	) name4424 (
		_w1976_,
		_w5931_,
		_w5932_
	);
	LUT2 #(
		.INIT('h1)
	) name4425 (
		_w1762_,
		_w5869_,
		_w5933_
	);
	LUT2 #(
		.INIT('h2)
	) name4426 (
		_w1973_,
		_w5933_,
		_w5934_
	);
	LUT2 #(
		.INIT('h1)
	) name4427 (
		_w5932_,
		_w5934_,
		_w5935_
	);
	LUT2 #(
		.INIT('h8)
	) name4428 (
		\TM0_pad ,
		\_2140__reg/NET0131 ,
		_w5936_
	);
	LUT2 #(
		.INIT('h1)
	) name4429 (
		_w4736_,
		_w5936_,
		_w5937_
	);
	LUT2 #(
		.INIT('h2)
	) name4430 (
		_w1976_,
		_w5937_,
		_w5938_
	);
	LUT2 #(
		.INIT('h1)
	) name4431 (
		_w1871_,
		_w5758_,
		_w5939_
	);
	LUT2 #(
		.INIT('h2)
	) name4432 (
		_w1973_,
		_w5939_,
		_w5940_
	);
	LUT2 #(
		.INIT('h1)
	) name4433 (
		_w5938_,
		_w5940_,
		_w5941_
	);
	LUT2 #(
		.INIT('h8)
	) name4434 (
		\TM0_pad ,
		\_2327__reg/NET0131 ,
		_w5942_
	);
	LUT2 #(
		.INIT('h1)
	) name4435 (
		_w3002_,
		_w5942_,
		_w5943_
	);
	LUT2 #(
		.INIT('h2)
	) name4436 (
		_w1976_,
		_w5943_,
		_w5944_
	);
	LUT2 #(
		.INIT('h1)
	) name4437 (
		_w1778_,
		_w5801_,
		_w5945_
	);
	LUT2 #(
		.INIT('h2)
	) name4438 (
		_w1973_,
		_w5945_,
		_w5946_
	);
	LUT2 #(
		.INIT('h1)
	) name4439 (
		_w5944_,
		_w5946_,
		_w5947_
	);
	LUT2 #(
		.INIT('h8)
	) name4440 (
		\TM0_pad ,
		\_2195__reg/NET0131 ,
		_w5948_
	);
	LUT2 #(
		.INIT('h2)
	) name4441 (
		\WX5963_reg/NET0131 ,
		\WX6027_reg/NET0131 ,
		_w5949_
	);
	LUT2 #(
		.INIT('h4)
	) name4442 (
		\WX5963_reg/NET0131 ,
		\WX6027_reg/NET0131 ,
		_w5950_
	);
	LUT2 #(
		.INIT('h1)
	) name4443 (
		_w5949_,
		_w5950_,
		_w5951_
	);
	LUT2 #(
		.INIT('h2)
	) name4444 (
		\WX5899_reg/NET0131 ,
		_w5951_,
		_w5952_
	);
	LUT2 #(
		.INIT('h4)
	) name4445 (
		\WX5899_reg/NET0131 ,
		_w5951_,
		_w5953_
	);
	LUT2 #(
		.INIT('h1)
	) name4446 (
		_w5952_,
		_w5953_,
		_w5954_
	);
	LUT2 #(
		.INIT('h2)
	) name4447 (
		\TM1_pad ,
		\WX5835_reg/NET0131 ,
		_w5955_
	);
	LUT2 #(
		.INIT('h4)
	) name4448 (
		\TM1_pad ,
		\WX5835_reg/NET0131 ,
		_w5956_
	);
	LUT2 #(
		.INIT('h1)
	) name4449 (
		_w5955_,
		_w5956_,
		_w5957_
	);
	LUT2 #(
		.INIT('h4)
	) name4450 (
		_w5954_,
		_w5957_,
		_w5958_
	);
	LUT2 #(
		.INIT('h2)
	) name4451 (
		_w5954_,
		_w5957_,
		_w5959_
	);
	LUT2 #(
		.INIT('h1)
	) name4452 (
		\TM0_pad ,
		_w5958_,
		_w5960_
	);
	LUT2 #(
		.INIT('h4)
	) name4453 (
		_w5959_,
		_w5960_,
		_w5961_
	);
	LUT2 #(
		.INIT('h1)
	) name4454 (
		_w5948_,
		_w5961_,
		_w5962_
	);
	LUT2 #(
		.INIT('h2)
	) name4455 (
		_w1976_,
		_w5962_,
		_w5963_
	);
	LUT2 #(
		.INIT('h1)
	) name4456 (
		_w1714_,
		_w5782_,
		_w5964_
	);
	LUT2 #(
		.INIT('h2)
	) name4457 (
		_w1973_,
		_w5964_,
		_w5965_
	);
	LUT2 #(
		.INIT('h1)
	) name4458 (
		_w5963_,
		_w5965_,
		_w5966_
	);
	LUT2 #(
		.INIT('h8)
	) name4459 (
		\TM0_pad ,
		\_2228__reg/NET0131 ,
		_w5967_
	);
	LUT2 #(
		.INIT('h2)
	) name4460 (
		\WX7254_reg/NET0131 ,
		\WX7318_reg/NET0131 ,
		_w5968_
	);
	LUT2 #(
		.INIT('h4)
	) name4461 (
		\WX7254_reg/NET0131 ,
		\WX7318_reg/NET0131 ,
		_w5969_
	);
	LUT2 #(
		.INIT('h1)
	) name4462 (
		_w5968_,
		_w5969_,
		_w5970_
	);
	LUT2 #(
		.INIT('h2)
	) name4463 (
		\WX7190_reg/NET0131 ,
		_w5970_,
		_w5971_
	);
	LUT2 #(
		.INIT('h4)
	) name4464 (
		\WX7190_reg/NET0131 ,
		_w5970_,
		_w5972_
	);
	LUT2 #(
		.INIT('h1)
	) name4465 (
		_w5971_,
		_w5972_,
		_w5973_
	);
	LUT2 #(
		.INIT('h2)
	) name4466 (
		\TM1_pad ,
		\WX7126_reg/NET0131 ,
		_w5974_
	);
	LUT2 #(
		.INIT('h4)
	) name4467 (
		\TM1_pad ,
		\WX7126_reg/NET0131 ,
		_w5975_
	);
	LUT2 #(
		.INIT('h1)
	) name4468 (
		_w5974_,
		_w5975_,
		_w5976_
	);
	LUT2 #(
		.INIT('h4)
	) name4469 (
		_w5973_,
		_w5976_,
		_w5977_
	);
	LUT2 #(
		.INIT('h2)
	) name4470 (
		_w5973_,
		_w5976_,
		_w5978_
	);
	LUT2 #(
		.INIT('h1)
	) name4471 (
		\TM0_pad ,
		_w5977_,
		_w5979_
	);
	LUT2 #(
		.INIT('h4)
	) name4472 (
		_w5978_,
		_w5979_,
		_w5980_
	);
	LUT2 #(
		.INIT('h1)
	) name4473 (
		_w5967_,
		_w5980_,
		_w5981_
	);
	LUT2 #(
		.INIT('h2)
	) name4474 (
		_w1976_,
		_w5981_,
		_w5982_
	);
	LUT2 #(
		.INIT('h1)
	) name4475 (
		_w1730_,
		_w5826_,
		_w5983_
	);
	LUT2 #(
		.INIT('h2)
	) name4476 (
		_w1973_,
		_w5983_,
		_w5984_
	);
	LUT2 #(
		.INIT('h1)
	) name4477 (
		_w5982_,
		_w5984_,
		_w5985_
	);
	LUT2 #(
		.INIT('h2)
	) name4478 (
		\WX2120_reg/NET0131 ,
		\WX2184_reg/NET0131 ,
		_w5986_
	);
	LUT2 #(
		.INIT('h4)
	) name4479 (
		\WX2120_reg/NET0131 ,
		\WX2184_reg/NET0131 ,
		_w5987_
	);
	LUT2 #(
		.INIT('h1)
	) name4480 (
		_w5986_,
		_w5987_,
		_w5988_
	);
	LUT2 #(
		.INIT('h2)
	) name4481 (
		\WX1992_reg/NET0131 ,
		\WX2056_reg/NET0131 ,
		_w5989_
	);
	LUT2 #(
		.INIT('h4)
	) name4482 (
		\WX1992_reg/NET0131 ,
		\WX2056_reg/NET0131 ,
		_w5990_
	);
	LUT2 #(
		.INIT('h1)
	) name4483 (
		_w5989_,
		_w5990_,
		_w5991_
	);
	LUT2 #(
		.INIT('h4)
	) name4484 (
		_w5988_,
		_w5991_,
		_w5992_
	);
	LUT2 #(
		.INIT('h2)
	) name4485 (
		_w5988_,
		_w5991_,
		_w5993_
	);
	LUT2 #(
		.INIT('h1)
	) name4486 (
		\TM0_pad ,
		_w5992_,
		_w5994_
	);
	LUT2 #(
		.INIT('h4)
	) name4487 (
		_w5993_,
		_w5994_,
		_w5995_
	);
	LUT2 #(
		.INIT('h2)
	) name4488 (
		_w3953_,
		_w5995_,
		_w5996_
	);
	LUT2 #(
		.INIT('h2)
	) name4489 (
		\TM0_pad ,
		\_2113__reg/NET0131 ,
		_w5997_
	);
	LUT2 #(
		.INIT('h2)
	) name4490 (
		_w1976_,
		_w5997_,
		_w5998_
	);
	LUT2 #(
		.INIT('h4)
	) name4491 (
		_w3963_,
		_w5998_,
		_w5999_
	);
	LUT2 #(
		.INIT('h1)
	) name4492 (
		_w5996_,
		_w5999_,
		_w6000_
	);
	LUT2 #(
		.INIT('h8)
	) name4493 (
		\TM0_pad ,
		\_2261__reg/NET0131 ,
		_w6001_
	);
	LUT2 #(
		.INIT('h2)
	) name4494 (
		\WX8545_reg/NET0131 ,
		\WX8609_reg/NET0131 ,
		_w6002_
	);
	LUT2 #(
		.INIT('h4)
	) name4495 (
		\WX8545_reg/NET0131 ,
		\WX8609_reg/NET0131 ,
		_w6003_
	);
	LUT2 #(
		.INIT('h1)
	) name4496 (
		_w6002_,
		_w6003_,
		_w6004_
	);
	LUT2 #(
		.INIT('h2)
	) name4497 (
		\WX8481_reg/NET0131 ,
		_w6004_,
		_w6005_
	);
	LUT2 #(
		.INIT('h4)
	) name4498 (
		\WX8481_reg/NET0131 ,
		_w6004_,
		_w6006_
	);
	LUT2 #(
		.INIT('h1)
	) name4499 (
		_w6005_,
		_w6006_,
		_w6007_
	);
	LUT2 #(
		.INIT('h2)
	) name4500 (
		\TM1_pad ,
		\WX8417_reg/NET0131 ,
		_w6008_
	);
	LUT2 #(
		.INIT('h4)
	) name4501 (
		\TM1_pad ,
		\WX8417_reg/NET0131 ,
		_w6009_
	);
	LUT2 #(
		.INIT('h1)
	) name4502 (
		_w6008_,
		_w6009_,
		_w6010_
	);
	LUT2 #(
		.INIT('h4)
	) name4503 (
		_w6007_,
		_w6010_,
		_w6011_
	);
	LUT2 #(
		.INIT('h2)
	) name4504 (
		_w6007_,
		_w6010_,
		_w6012_
	);
	LUT2 #(
		.INIT('h1)
	) name4505 (
		\TM0_pad ,
		_w6011_,
		_w6013_
	);
	LUT2 #(
		.INIT('h4)
	) name4506 (
		_w6012_,
		_w6013_,
		_w6014_
	);
	LUT2 #(
		.INIT('h1)
	) name4507 (
		_w6001_,
		_w6014_,
		_w6015_
	);
	LUT2 #(
		.INIT('h2)
	) name4508 (
		_w1976_,
		_w6015_,
		_w6016_
	);
	LUT2 #(
		.INIT('h1)
	) name4509 (
		_w1746_,
		_w5845_,
		_w6017_
	);
	LUT2 #(
		.INIT('h2)
	) name4510 (
		_w1973_,
		_w6017_,
		_w6018_
	);
	LUT2 #(
		.INIT('h1)
	) name4511 (
		_w6016_,
		_w6018_,
		_w6019_
	);
	LUT2 #(
		.INIT('h1)
	) name4512 (
		\TM0_pad ,
		_w1845_,
		_w6020_
	);
	LUT2 #(
		.INIT('h2)
	) name4513 (
		_w4239_,
		_w6020_,
		_w6021_
	);
	LUT2 #(
		.INIT('h2)
	) name4514 (
		\TM0_pad ,
		\_2079__reg/NET0131 ,
		_w6022_
	);
	LUT2 #(
		.INIT('h2)
	) name4515 (
		\WX2124_reg/NET0131 ,
		\WX2188_reg/NET0131 ,
		_w6023_
	);
	LUT2 #(
		.INIT('h4)
	) name4516 (
		\WX2124_reg/NET0131 ,
		\WX2188_reg/NET0131 ,
		_w6024_
	);
	LUT2 #(
		.INIT('h1)
	) name4517 (
		_w6023_,
		_w6024_,
		_w6025_
	);
	LUT2 #(
		.INIT('h2)
	) name4518 (
		\WX1996_reg/NET0131 ,
		\WX2060_reg/NET0131 ,
		_w6026_
	);
	LUT2 #(
		.INIT('h4)
	) name4519 (
		\WX1996_reg/NET0131 ,
		\WX2060_reg/NET0131 ,
		_w6027_
	);
	LUT2 #(
		.INIT('h1)
	) name4520 (
		_w6026_,
		_w6027_,
		_w6028_
	);
	LUT2 #(
		.INIT('h4)
	) name4521 (
		_w6025_,
		_w6028_,
		_w6029_
	);
	LUT2 #(
		.INIT('h2)
	) name4522 (
		_w6025_,
		_w6028_,
		_w6030_
	);
	LUT2 #(
		.INIT('h1)
	) name4523 (
		\TM0_pad ,
		_w6029_,
		_w6031_
	);
	LUT2 #(
		.INIT('h4)
	) name4524 (
		_w6030_,
		_w6031_,
		_w6032_
	);
	LUT2 #(
		.INIT('h2)
	) name4525 (
		_w1976_,
		_w6022_,
		_w6033_
	);
	LUT2 #(
		.INIT('h4)
	) name4526 (
		_w6032_,
		_w6033_,
		_w6034_
	);
	LUT2 #(
		.INIT('h1)
	) name4527 (
		_w6021_,
		_w6034_,
		_w6035_
	);
	LUT2 #(
		.INIT('h1)
	) name4528 (
		\TM0_pad ,
		_w1517_,
		_w6036_
	);
	LUT2 #(
		.INIT('h2)
	) name4529 (
		_w4510_,
		_w6036_,
		_w6037_
	);
	LUT2 #(
		.INIT('h2)
	) name4530 (
		\TM0_pad ,
		\_2077__reg/NET0131 ,
		_w6038_
	);
	LUT2 #(
		.INIT('h2)
	) name4531 (
		\WX2128_reg/NET0131 ,
		\WX2192_reg/NET0131 ,
		_w6039_
	);
	LUT2 #(
		.INIT('h4)
	) name4532 (
		\WX2128_reg/NET0131 ,
		\WX2192_reg/NET0131 ,
		_w6040_
	);
	LUT2 #(
		.INIT('h1)
	) name4533 (
		_w6039_,
		_w6040_,
		_w6041_
	);
	LUT2 #(
		.INIT('h2)
	) name4534 (
		\WX2000_reg/NET0131 ,
		\WX2064_reg/NET0131 ,
		_w6042_
	);
	LUT2 #(
		.INIT('h4)
	) name4535 (
		\WX2000_reg/NET0131 ,
		\WX2064_reg/NET0131 ,
		_w6043_
	);
	LUT2 #(
		.INIT('h1)
	) name4536 (
		_w6042_,
		_w6043_,
		_w6044_
	);
	LUT2 #(
		.INIT('h4)
	) name4537 (
		_w6041_,
		_w6044_,
		_w6045_
	);
	LUT2 #(
		.INIT('h2)
	) name4538 (
		_w6041_,
		_w6044_,
		_w6046_
	);
	LUT2 #(
		.INIT('h1)
	) name4539 (
		\TM0_pad ,
		_w6045_,
		_w6047_
	);
	LUT2 #(
		.INIT('h4)
	) name4540 (
		_w6046_,
		_w6047_,
		_w6048_
	);
	LUT2 #(
		.INIT('h2)
	) name4541 (
		_w1976_,
		_w6038_,
		_w6049_
	);
	LUT2 #(
		.INIT('h4)
	) name4542 (
		_w6048_,
		_w6049_,
		_w6050_
	);
	LUT2 #(
		.INIT('h1)
	) name4543 (
		_w6037_,
		_w6050_,
		_w6051_
	);
	LUT2 #(
		.INIT('h1)
	) name4544 (
		_w1871_,
		_w5279_,
		_w6052_
	);
	LUT2 #(
		.INIT('h2)
	) name4545 (
		_w1973_,
		_w6052_,
		_w6053_
	);
	LUT2 #(
		.INIT('h1)
	) name4546 (
		\DATA_0_31_pad ,
		\TM0_pad ,
		_w6054_
	);
	LUT2 #(
		.INIT('h2)
	) name4547 (
		\TM0_pad ,
		\_2364__reg/NET0131 ,
		_w6055_
	);
	LUT2 #(
		.INIT('h2)
	) name4548 (
		_w1976_,
		_w6054_,
		_w6056_
	);
	LUT2 #(
		.INIT('h4)
	) name4549 (
		_w6055_,
		_w6056_,
		_w6057_
	);
	LUT2 #(
		.INIT('h1)
	) name4550 (
		_w6053_,
		_w6057_,
		_w6058_
	);
	LUT2 #(
		.INIT('h2)
	) name4551 (
		_w3953_,
		_w4659_,
		_w6059_
	);
	LUT2 #(
		.INIT('h1)
	) name4552 (
		\DATA_0_4_pad ,
		\TM0_pad ,
		_w6060_
	);
	LUT2 #(
		.INIT('h2)
	) name4553 (
		\TM0_pad ,
		\_2337__reg/NET0131 ,
		_w6061_
	);
	LUT2 #(
		.INIT('h2)
	) name4554 (
		_w1976_,
		_w6060_,
		_w6062_
	);
	LUT2 #(
		.INIT('h4)
	) name4555 (
		_w6061_,
		_w6062_,
		_w6063_
	);
	LUT2 #(
		.INIT('h1)
	) name4556 (
		_w6059_,
		_w6063_,
		_w6064_
	);
	LUT2 #(
		.INIT('h8)
	) name4557 (
		RESET_pad,
		\WX10881_reg/NET0131 ,
		_w6065_
	);
	LUT2 #(
		.INIT('h8)
	) name4558 (
		\TM0_pad ,
		\_2161__reg/NET0131 ,
		_w6066_
	);
	LUT2 #(
		.INIT('h2)
	) name4559 (
		\WX4674_reg/NET0131 ,
		\WX4738_reg/NET0131 ,
		_w6067_
	);
	LUT2 #(
		.INIT('h4)
	) name4560 (
		\WX4674_reg/NET0131 ,
		\WX4738_reg/NET0131 ,
		_w6068_
	);
	LUT2 #(
		.INIT('h1)
	) name4561 (
		_w6067_,
		_w6068_,
		_w6069_
	);
	LUT2 #(
		.INIT('h2)
	) name4562 (
		\WX4610_reg/NET0131 ,
		_w6069_,
		_w6070_
	);
	LUT2 #(
		.INIT('h4)
	) name4563 (
		\WX4610_reg/NET0131 ,
		_w6069_,
		_w6071_
	);
	LUT2 #(
		.INIT('h1)
	) name4564 (
		_w6070_,
		_w6071_,
		_w6072_
	);
	LUT2 #(
		.INIT('h2)
	) name4565 (
		\TM1_pad ,
		\WX4546_reg/NET0131 ,
		_w6073_
	);
	LUT2 #(
		.INIT('h4)
	) name4566 (
		\TM1_pad ,
		\WX4546_reg/NET0131 ,
		_w6074_
	);
	LUT2 #(
		.INIT('h1)
	) name4567 (
		_w6073_,
		_w6074_,
		_w6075_
	);
	LUT2 #(
		.INIT('h4)
	) name4568 (
		_w6072_,
		_w6075_,
		_w6076_
	);
	LUT2 #(
		.INIT('h2)
	) name4569 (
		_w6072_,
		_w6075_,
		_w6077_
	);
	LUT2 #(
		.INIT('h1)
	) name4570 (
		\TM0_pad ,
		_w6076_,
		_w6078_
	);
	LUT2 #(
		.INIT('h4)
	) name4571 (
		_w6077_,
		_w6078_,
		_w6079_
	);
	LUT2 #(
		.INIT('h1)
	) name4572 (
		_w6066_,
		_w6079_,
		_w6080_
	);
	LUT2 #(
		.INIT('h2)
	) name4573 (
		_w1976_,
		_w6080_,
		_w6081_
	);
	LUT2 #(
		.INIT('h1)
	) name4574 (
		_w1682_,
		_w3874_,
		_w6082_
	);
	LUT2 #(
		.INIT('h2)
	) name4575 (
		_w1973_,
		_w6082_,
		_w6083_
	);
	LUT2 #(
		.INIT('h1)
	) name4576 (
		_w6081_,
		_w6083_,
		_w6084_
	);
	LUT2 #(
		.INIT('h8)
	) name4577 (
		\TM0_pad ,
		\_2293__reg/NET0131 ,
		_w6085_
	);
	LUT2 #(
		.INIT('h2)
	) name4578 (
		\WX9838_reg/NET0131 ,
		\WX9902_reg/NET0131 ,
		_w6086_
	);
	LUT2 #(
		.INIT('h4)
	) name4579 (
		\WX9838_reg/NET0131 ,
		\WX9902_reg/NET0131 ,
		_w6087_
	);
	LUT2 #(
		.INIT('h1)
	) name4580 (
		_w6086_,
		_w6087_,
		_w6088_
	);
	LUT2 #(
		.INIT('h2)
	) name4581 (
		\WX9774_reg/NET0131 ,
		_w6088_,
		_w6089_
	);
	LUT2 #(
		.INIT('h4)
	) name4582 (
		\WX9774_reg/NET0131 ,
		_w6088_,
		_w6090_
	);
	LUT2 #(
		.INIT('h1)
	) name4583 (
		_w6089_,
		_w6090_,
		_w6091_
	);
	LUT2 #(
		.INIT('h2)
	) name4584 (
		\TM1_pad ,
		\WX9710_reg/NET0131 ,
		_w6092_
	);
	LUT2 #(
		.INIT('h4)
	) name4585 (
		\TM1_pad ,
		\WX9710_reg/NET0131 ,
		_w6093_
	);
	LUT2 #(
		.INIT('h1)
	) name4586 (
		_w6092_,
		_w6093_,
		_w6094_
	);
	LUT2 #(
		.INIT('h4)
	) name4587 (
		_w6091_,
		_w6094_,
		_w6095_
	);
	LUT2 #(
		.INIT('h2)
	) name4588 (
		_w6091_,
		_w6094_,
		_w6096_
	);
	LUT2 #(
		.INIT('h1)
	) name4589 (
		\TM0_pad ,
		_w6095_,
		_w6097_
	);
	LUT2 #(
		.INIT('h4)
	) name4590 (
		_w6096_,
		_w6097_,
		_w6098_
	);
	LUT2 #(
		.INIT('h1)
	) name4591 (
		_w6085_,
		_w6098_,
		_w6099_
	);
	LUT2 #(
		.INIT('h2)
	) name4592 (
		_w1976_,
		_w6099_,
		_w6100_
	);
	LUT2 #(
		.INIT('h1)
	) name4593 (
		_w1746_,
		_w6014_,
		_w6101_
	);
	LUT2 #(
		.INIT('h2)
	) name4594 (
		_w1973_,
		_w6101_,
		_w6102_
	);
	LUT2 #(
		.INIT('h1)
	) name4595 (
		_w6100_,
		_w6102_,
		_w6103_
	);
	LUT2 #(
		.INIT('h8)
	) name4596 (
		\TM0_pad ,
		\_2326__reg/NET0131 ,
		_w6104_
	);
	LUT2 #(
		.INIT('h1)
	) name4597 (
		_w3163_,
		_w6104_,
		_w6105_
	);
	LUT2 #(
		.INIT('h2)
	) name4598 (
		_w1976_,
		_w6105_,
		_w6106_
	);
	LUT2 #(
		.INIT('h1)
	) name4599 (
		_w1762_,
		_w5930_,
		_w6107_
	);
	LUT2 #(
		.INIT('h2)
	) name4600 (
		_w1973_,
		_w6107_,
		_w6108_
	);
	LUT2 #(
		.INIT('h1)
	) name4601 (
		_w6106_,
		_w6108_,
		_w6109_
	);
	LUT2 #(
		.INIT('h8)
	) name4602 (
		\TM0_pad ,
		\_2194__reg/NET0131 ,
		_w6110_
	);
	LUT2 #(
		.INIT('h2)
	) name4603 (
		\WX5965_reg/NET0131 ,
		\WX6029_reg/NET0131 ,
		_w6111_
	);
	LUT2 #(
		.INIT('h4)
	) name4604 (
		\WX5965_reg/NET0131 ,
		\WX6029_reg/NET0131 ,
		_w6112_
	);
	LUT2 #(
		.INIT('h1)
	) name4605 (
		_w6111_,
		_w6112_,
		_w6113_
	);
	LUT2 #(
		.INIT('h2)
	) name4606 (
		\WX5901_reg/NET0131 ,
		_w6113_,
		_w6114_
	);
	LUT2 #(
		.INIT('h4)
	) name4607 (
		\WX5901_reg/NET0131 ,
		_w6113_,
		_w6115_
	);
	LUT2 #(
		.INIT('h1)
	) name4608 (
		_w6114_,
		_w6115_,
		_w6116_
	);
	LUT2 #(
		.INIT('h2)
	) name4609 (
		\TM1_pad ,
		\WX5837_reg/NET0131 ,
		_w6117_
	);
	LUT2 #(
		.INIT('h4)
	) name4610 (
		\TM1_pad ,
		\WX5837_reg/NET0131 ,
		_w6118_
	);
	LUT2 #(
		.INIT('h1)
	) name4611 (
		_w6117_,
		_w6118_,
		_w6119_
	);
	LUT2 #(
		.INIT('h4)
	) name4612 (
		_w6116_,
		_w6119_,
		_w6120_
	);
	LUT2 #(
		.INIT('h2)
	) name4613 (
		_w6116_,
		_w6119_,
		_w6121_
	);
	LUT2 #(
		.INIT('h1)
	) name4614 (
		\TM0_pad ,
		_w6120_,
		_w6122_
	);
	LUT2 #(
		.INIT('h4)
	) name4615 (
		_w6121_,
		_w6122_,
		_w6123_
	);
	LUT2 #(
		.INIT('h1)
	) name4616 (
		_w6110_,
		_w6123_,
		_w6124_
	);
	LUT2 #(
		.INIT('h2)
	) name4617 (
		_w1976_,
		_w6124_,
		_w6125_
	);
	LUT2 #(
		.INIT('h1)
	) name4618 (
		_w1698_,
		_w5911_,
		_w6126_
	);
	LUT2 #(
		.INIT('h2)
	) name4619 (
		_w1973_,
		_w6126_,
		_w6127_
	);
	LUT2 #(
		.INIT('h1)
	) name4620 (
		_w6125_,
		_w6127_,
		_w6128_
	);
	LUT2 #(
		.INIT('h8)
	) name4621 (
		\TM0_pad ,
		\_2227__reg/NET0131 ,
		_w6129_
	);
	LUT2 #(
		.INIT('h2)
	) name4622 (
		\WX7256_reg/NET0131 ,
		\WX7320_reg/NET0131 ,
		_w6130_
	);
	LUT2 #(
		.INIT('h4)
	) name4623 (
		\WX7256_reg/NET0131 ,
		\WX7320_reg/NET0131 ,
		_w6131_
	);
	LUT2 #(
		.INIT('h1)
	) name4624 (
		_w6130_,
		_w6131_,
		_w6132_
	);
	LUT2 #(
		.INIT('h2)
	) name4625 (
		\WX7192_reg/NET0131 ,
		_w6132_,
		_w6133_
	);
	LUT2 #(
		.INIT('h4)
	) name4626 (
		\WX7192_reg/NET0131 ,
		_w6132_,
		_w6134_
	);
	LUT2 #(
		.INIT('h1)
	) name4627 (
		_w6133_,
		_w6134_,
		_w6135_
	);
	LUT2 #(
		.INIT('h2)
	) name4628 (
		\TM1_pad ,
		\WX7128_reg/NET0131 ,
		_w6136_
	);
	LUT2 #(
		.INIT('h4)
	) name4629 (
		\TM1_pad ,
		\WX7128_reg/NET0131 ,
		_w6137_
	);
	LUT2 #(
		.INIT('h1)
	) name4630 (
		_w6136_,
		_w6137_,
		_w6138_
	);
	LUT2 #(
		.INIT('h4)
	) name4631 (
		_w6135_,
		_w6138_,
		_w6139_
	);
	LUT2 #(
		.INIT('h2)
	) name4632 (
		_w6135_,
		_w6138_,
		_w6140_
	);
	LUT2 #(
		.INIT('h1)
	) name4633 (
		\TM0_pad ,
		_w6139_,
		_w6141_
	);
	LUT2 #(
		.INIT('h4)
	) name4634 (
		_w6140_,
		_w6141_,
		_w6142_
	);
	LUT2 #(
		.INIT('h1)
	) name4635 (
		_w6129_,
		_w6142_,
		_w6143_
	);
	LUT2 #(
		.INIT('h2)
	) name4636 (
		_w1976_,
		_w6143_,
		_w6144_
	);
	LUT2 #(
		.INIT('h1)
	) name4637 (
		_w1714_,
		_w5961_,
		_w6145_
	);
	LUT2 #(
		.INIT('h2)
	) name4638 (
		_w1973_,
		_w6145_,
		_w6146_
	);
	LUT2 #(
		.INIT('h1)
	) name4639 (
		_w6144_,
		_w6146_,
		_w6147_
	);
	LUT2 #(
		.INIT('h2)
	) name4640 (
		_w4101_,
		_w5887_,
		_w6148_
	);
	LUT2 #(
		.INIT('h2)
	) name4641 (
		\TM0_pad ,
		\_2112__reg/NET0131 ,
		_w6149_
	);
	LUT2 #(
		.INIT('h2)
	) name4642 (
		_w1976_,
		_w6149_,
		_w6150_
	);
	LUT2 #(
		.INIT('h4)
	) name4643 (
		_w4111_,
		_w6150_,
		_w6151_
	);
	LUT2 #(
		.INIT('h1)
	) name4644 (
		_w6148_,
		_w6151_,
		_w6152_
	);
	LUT2 #(
		.INIT('h8)
	) name4645 (
		\TM0_pad ,
		\_2260__reg/NET0131 ,
		_w6153_
	);
	LUT2 #(
		.INIT('h2)
	) name4646 (
		\WX8547_reg/NET0131 ,
		\WX8611_reg/NET0131 ,
		_w6154_
	);
	LUT2 #(
		.INIT('h4)
	) name4647 (
		\WX8547_reg/NET0131 ,
		\WX8611_reg/NET0131 ,
		_w6155_
	);
	LUT2 #(
		.INIT('h1)
	) name4648 (
		_w6154_,
		_w6155_,
		_w6156_
	);
	LUT2 #(
		.INIT('h2)
	) name4649 (
		\WX8483_reg/NET0131 ,
		_w6156_,
		_w6157_
	);
	LUT2 #(
		.INIT('h4)
	) name4650 (
		\WX8483_reg/NET0131 ,
		_w6156_,
		_w6158_
	);
	LUT2 #(
		.INIT('h1)
	) name4651 (
		_w6157_,
		_w6158_,
		_w6159_
	);
	LUT2 #(
		.INIT('h2)
	) name4652 (
		\TM1_pad ,
		\WX8419_reg/NET0131 ,
		_w6160_
	);
	LUT2 #(
		.INIT('h4)
	) name4653 (
		\TM1_pad ,
		\WX8419_reg/NET0131 ,
		_w6161_
	);
	LUT2 #(
		.INIT('h1)
	) name4654 (
		_w6160_,
		_w6161_,
		_w6162_
	);
	LUT2 #(
		.INIT('h4)
	) name4655 (
		_w6159_,
		_w6162_,
		_w6163_
	);
	LUT2 #(
		.INIT('h2)
	) name4656 (
		_w6159_,
		_w6162_,
		_w6164_
	);
	LUT2 #(
		.INIT('h1)
	) name4657 (
		\TM0_pad ,
		_w6163_,
		_w6165_
	);
	LUT2 #(
		.INIT('h4)
	) name4658 (
		_w6164_,
		_w6165_,
		_w6166_
	);
	LUT2 #(
		.INIT('h1)
	) name4659 (
		_w6153_,
		_w6166_,
		_w6167_
	);
	LUT2 #(
		.INIT('h2)
	) name4660 (
		_w1976_,
		_w6167_,
		_w6168_
	);
	LUT2 #(
		.INIT('h1)
	) name4661 (
		_w1730_,
		_w5980_,
		_w6169_
	);
	LUT2 #(
		.INIT('h2)
	) name4662 (
		_w1973_,
		_w6169_,
		_w6170_
	);
	LUT2 #(
		.INIT('h1)
	) name4663 (
		_w6168_,
		_w6170_,
		_w6171_
	);
	LUT2 #(
		.INIT('h2)
	) name4664 (
		_w4101_,
		_w4823_,
		_w6172_
	);
	LUT2 #(
		.INIT('h1)
	) name4665 (
		\DATA_0_3_pad ,
		\TM0_pad ,
		_w6173_
	);
	LUT2 #(
		.INIT('h2)
	) name4666 (
		\TM0_pad ,
		\_2336__reg/NET0131 ,
		_w6174_
	);
	LUT2 #(
		.INIT('h2)
	) name4667 (
		_w1976_,
		_w6173_,
		_w6175_
	);
	LUT2 #(
		.INIT('h4)
	) name4668 (
		_w6174_,
		_w6175_,
		_w6176_
	);
	LUT2 #(
		.INIT('h1)
	) name4669 (
		_w6172_,
		_w6176_,
		_w6177_
	);
	LUT2 #(
		.INIT('h8)
	) name4670 (
		RESET_pad,
		\WX10883_reg/NET0131 ,
		_w6178_
	);
	LUT2 #(
		.INIT('h8)
	) name4671 (
		\TM0_pad ,
		\_2160__reg/NET0131 ,
		_w6179_
	);
	LUT2 #(
		.INIT('h2)
	) name4672 (
		\TM1_pad ,
		\WX4548_reg/NET0131 ,
		_w6180_
	);
	LUT2 #(
		.INIT('h4)
	) name4673 (
		\TM1_pad ,
		\WX4548_reg/NET0131 ,
		_w6181_
	);
	LUT2 #(
		.INIT('h1)
	) name4674 (
		_w6180_,
		_w6181_,
		_w6182_
	);
	LUT2 #(
		.INIT('h1)
	) name4675 (
		\WX4612_reg/NET0131 ,
		_w6182_,
		_w6183_
	);
	LUT2 #(
		.INIT('h8)
	) name4676 (
		\WX4612_reg/NET0131 ,
		_w6182_,
		_w6184_
	);
	LUT2 #(
		.INIT('h1)
	) name4677 (
		_w6183_,
		_w6184_,
		_w6185_
	);
	LUT2 #(
		.INIT('h2)
	) name4678 (
		\WX4676_reg/NET0131 ,
		\WX4740_reg/NET0131 ,
		_w6186_
	);
	LUT2 #(
		.INIT('h4)
	) name4679 (
		\WX4676_reg/NET0131 ,
		\WX4740_reg/NET0131 ,
		_w6187_
	);
	LUT2 #(
		.INIT('h1)
	) name4680 (
		_w6186_,
		_w6187_,
		_w6188_
	);
	LUT2 #(
		.INIT('h1)
	) name4681 (
		_w6185_,
		_w6188_,
		_w6189_
	);
	LUT2 #(
		.INIT('h8)
	) name4682 (
		_w6185_,
		_w6188_,
		_w6190_
	);
	LUT2 #(
		.INIT('h1)
	) name4683 (
		\TM0_pad ,
		_w6189_,
		_w6191_
	);
	LUT2 #(
		.INIT('h4)
	) name4684 (
		_w6190_,
		_w6191_,
		_w6192_
	);
	LUT2 #(
		.INIT('h1)
	) name4685 (
		_w6179_,
		_w6192_,
		_w6193_
	);
	LUT2 #(
		.INIT('h2)
	) name4686 (
		_w1976_,
		_w6193_,
		_w6194_
	);
	LUT2 #(
		.INIT('h1)
	) name4687 (
		_w1653_,
		_w4022_,
		_w6195_
	);
	LUT2 #(
		.INIT('h2)
	) name4688 (
		_w1973_,
		_w6195_,
		_w6196_
	);
	LUT2 #(
		.INIT('h1)
	) name4689 (
		_w6194_,
		_w6196_,
		_w6197_
	);
	LUT2 #(
		.INIT('h8)
	) name4690 (
		\TM0_pad ,
		\_2159__reg/NET0131 ,
		_w6198_
	);
	LUT2 #(
		.INIT('h2)
	) name4691 (
		\WX4678_reg/NET0131 ,
		\WX4742_reg/NET0131 ,
		_w6199_
	);
	LUT2 #(
		.INIT('h4)
	) name4692 (
		\WX4678_reg/NET0131 ,
		\WX4742_reg/NET0131 ,
		_w6200_
	);
	LUT2 #(
		.INIT('h1)
	) name4693 (
		_w6199_,
		_w6200_,
		_w6201_
	);
	LUT2 #(
		.INIT('h2)
	) name4694 (
		\WX4614_reg/NET0131 ,
		_w6201_,
		_w6202_
	);
	LUT2 #(
		.INIT('h4)
	) name4695 (
		\WX4614_reg/NET0131 ,
		_w6201_,
		_w6203_
	);
	LUT2 #(
		.INIT('h1)
	) name4696 (
		_w6202_,
		_w6203_,
		_w6204_
	);
	LUT2 #(
		.INIT('h2)
	) name4697 (
		\TM1_pad ,
		\WX4550_reg/NET0131 ,
		_w6205_
	);
	LUT2 #(
		.INIT('h4)
	) name4698 (
		\TM1_pad ,
		\WX4550_reg/NET0131 ,
		_w6206_
	);
	LUT2 #(
		.INIT('h1)
	) name4699 (
		_w6205_,
		_w6206_,
		_w6207_
	);
	LUT2 #(
		.INIT('h4)
	) name4700 (
		_w6204_,
		_w6207_,
		_w6208_
	);
	LUT2 #(
		.INIT('h2)
	) name4701 (
		_w6204_,
		_w6207_,
		_w6209_
	);
	LUT2 #(
		.INIT('h1)
	) name4702 (
		\TM0_pad ,
		_w6208_,
		_w6210_
	);
	LUT2 #(
		.INIT('h4)
	) name4703 (
		_w6209_,
		_w6210_,
		_w6211_
	);
	LUT2 #(
		.INIT('h1)
	) name4704 (
		_w6198_,
		_w6211_,
		_w6212_
	);
	LUT2 #(
		.INIT('h2)
	) name4705 (
		_w1976_,
		_w6212_,
		_w6213_
	);
	LUT2 #(
		.INIT('h1)
	) name4706 (
		_w1637_,
		_w4160_,
		_w6214_
	);
	LUT2 #(
		.INIT('h2)
	) name4707 (
		_w1973_,
		_w6214_,
		_w6215_
	);
	LUT2 #(
		.INIT('h1)
	) name4708 (
		_w6213_,
		_w6215_,
		_w6216_
	);
	LUT2 #(
		.INIT('h8)
	) name4709 (
		\TM0_pad ,
		\_2158__reg/NET0131 ,
		_w6217_
	);
	LUT2 #(
		.INIT('h2)
	) name4710 (
		\WX4680_reg/NET0131 ,
		\WX4744_reg/NET0131 ,
		_w6218_
	);
	LUT2 #(
		.INIT('h4)
	) name4711 (
		\WX4680_reg/NET0131 ,
		\WX4744_reg/NET0131 ,
		_w6219_
	);
	LUT2 #(
		.INIT('h1)
	) name4712 (
		_w6218_,
		_w6219_,
		_w6220_
	);
	LUT2 #(
		.INIT('h2)
	) name4713 (
		\WX4616_reg/NET0131 ,
		_w6220_,
		_w6221_
	);
	LUT2 #(
		.INIT('h4)
	) name4714 (
		\WX4616_reg/NET0131 ,
		_w6220_,
		_w6222_
	);
	LUT2 #(
		.INIT('h1)
	) name4715 (
		_w6221_,
		_w6222_,
		_w6223_
	);
	LUT2 #(
		.INIT('h2)
	) name4716 (
		\TM1_pad ,
		\WX4552_reg/NET0131 ,
		_w6224_
	);
	LUT2 #(
		.INIT('h4)
	) name4717 (
		\TM1_pad ,
		\WX4552_reg/NET0131 ,
		_w6225_
	);
	LUT2 #(
		.INIT('h1)
	) name4718 (
		_w6224_,
		_w6225_,
		_w6226_
	);
	LUT2 #(
		.INIT('h4)
	) name4719 (
		_w6223_,
		_w6226_,
		_w6227_
	);
	LUT2 #(
		.INIT('h2)
	) name4720 (
		_w6223_,
		_w6226_,
		_w6228_
	);
	LUT2 #(
		.INIT('h1)
	) name4721 (
		\TM0_pad ,
		_w6227_,
		_w6229_
	);
	LUT2 #(
		.INIT('h4)
	) name4722 (
		_w6228_,
		_w6229_,
		_w6230_
	);
	LUT2 #(
		.INIT('h1)
	) name4723 (
		_w6217_,
		_w6230_,
		_w6231_
	);
	LUT2 #(
		.INIT('h2)
	) name4724 (
		_w1976_,
		_w6231_,
		_w6232_
	);
	LUT2 #(
		.INIT('h1)
	) name4725 (
		_w1621_,
		_w4323_,
		_w6233_
	);
	LUT2 #(
		.INIT('h2)
	) name4726 (
		_w1973_,
		_w6233_,
		_w6234_
	);
	LUT2 #(
		.INIT('h1)
	) name4727 (
		_w6232_,
		_w6234_,
		_w6235_
	);
	LUT2 #(
		.INIT('h8)
	) name4728 (
		\TM0_pad ,
		\_2157__reg/NET0131 ,
		_w6236_
	);
	LUT2 #(
		.INIT('h1)
	) name4729 (
		_w2233_,
		_w6236_,
		_w6237_
	);
	LUT2 #(
		.INIT('h2)
	) name4730 (
		_w1976_,
		_w6237_,
		_w6238_
	);
	LUT2 #(
		.INIT('h1)
	) name4731 (
		_w1605_,
		_w4466_,
		_w6239_
	);
	LUT2 #(
		.INIT('h2)
	) name4732 (
		_w1973_,
		_w6239_,
		_w6240_
	);
	LUT2 #(
		.INIT('h1)
	) name4733 (
		_w6238_,
		_w6240_,
		_w6241_
	);
	LUT2 #(
		.INIT('h8)
	) name4734 (
		\TM0_pad ,
		\_2292__reg/NET0131 ,
		_w6242_
	);
	LUT2 #(
		.INIT('h2)
	) name4735 (
		\WX9840_reg/NET0131 ,
		\WX9904_reg/NET0131 ,
		_w6243_
	);
	LUT2 #(
		.INIT('h4)
	) name4736 (
		\WX9840_reg/NET0131 ,
		\WX9904_reg/NET0131 ,
		_w6244_
	);
	LUT2 #(
		.INIT('h1)
	) name4737 (
		_w6243_,
		_w6244_,
		_w6245_
	);
	LUT2 #(
		.INIT('h2)
	) name4738 (
		\WX9776_reg/NET0131 ,
		_w6245_,
		_w6246_
	);
	LUT2 #(
		.INIT('h4)
	) name4739 (
		\WX9776_reg/NET0131 ,
		_w6245_,
		_w6247_
	);
	LUT2 #(
		.INIT('h1)
	) name4740 (
		_w6246_,
		_w6247_,
		_w6248_
	);
	LUT2 #(
		.INIT('h2)
	) name4741 (
		\TM1_pad ,
		\WX9712_reg/NET0131 ,
		_w6249_
	);
	LUT2 #(
		.INIT('h4)
	) name4742 (
		\TM1_pad ,
		\WX9712_reg/NET0131 ,
		_w6250_
	);
	LUT2 #(
		.INIT('h1)
	) name4743 (
		_w6249_,
		_w6250_,
		_w6251_
	);
	LUT2 #(
		.INIT('h4)
	) name4744 (
		_w6248_,
		_w6251_,
		_w6252_
	);
	LUT2 #(
		.INIT('h2)
	) name4745 (
		_w6248_,
		_w6251_,
		_w6253_
	);
	LUT2 #(
		.INIT('h1)
	) name4746 (
		\TM0_pad ,
		_w6252_,
		_w6254_
	);
	LUT2 #(
		.INIT('h4)
	) name4747 (
		_w6253_,
		_w6254_,
		_w6255_
	);
	LUT2 #(
		.INIT('h1)
	) name4748 (
		_w6242_,
		_w6255_,
		_w6256_
	);
	LUT2 #(
		.INIT('h2)
	) name4749 (
		_w1976_,
		_w6256_,
		_w6257_
	);
	LUT2 #(
		.INIT('h1)
	) name4750 (
		_w1730_,
		_w6166_,
		_w6258_
	);
	LUT2 #(
		.INIT('h2)
	) name4751 (
		_w1973_,
		_w6258_,
		_w6259_
	);
	LUT2 #(
		.INIT('h1)
	) name4752 (
		_w6257_,
		_w6259_,
		_w6260_
	);
	LUT2 #(
		.INIT('h8)
	) name4753 (
		\TM0_pad ,
		\_2291__reg/NET0131 ,
		_w6261_
	);
	LUT2 #(
		.INIT('h2)
	) name4754 (
		\WX9842_reg/NET0131 ,
		\WX9906_reg/NET0131 ,
		_w6262_
	);
	LUT2 #(
		.INIT('h4)
	) name4755 (
		\WX9842_reg/NET0131 ,
		\WX9906_reg/NET0131 ,
		_w6263_
	);
	LUT2 #(
		.INIT('h1)
	) name4756 (
		_w6262_,
		_w6263_,
		_w6264_
	);
	LUT2 #(
		.INIT('h2)
	) name4757 (
		\WX9778_reg/NET0131 ,
		_w6264_,
		_w6265_
	);
	LUT2 #(
		.INIT('h4)
	) name4758 (
		\WX9778_reg/NET0131 ,
		_w6264_,
		_w6266_
	);
	LUT2 #(
		.INIT('h1)
	) name4759 (
		_w6265_,
		_w6266_,
		_w6267_
	);
	LUT2 #(
		.INIT('h2)
	) name4760 (
		\TM1_pad ,
		\WX9714_reg/NET0131 ,
		_w6268_
	);
	LUT2 #(
		.INIT('h4)
	) name4761 (
		\TM1_pad ,
		\WX9714_reg/NET0131 ,
		_w6269_
	);
	LUT2 #(
		.INIT('h1)
	) name4762 (
		_w6268_,
		_w6269_,
		_w6270_
	);
	LUT2 #(
		.INIT('h4)
	) name4763 (
		_w6267_,
		_w6270_,
		_w6271_
	);
	LUT2 #(
		.INIT('h2)
	) name4764 (
		_w6267_,
		_w6270_,
		_w6272_
	);
	LUT2 #(
		.INIT('h1)
	) name4765 (
		\TM0_pad ,
		_w6271_,
		_w6273_
	);
	LUT2 #(
		.INIT('h4)
	) name4766 (
		_w6272_,
		_w6273_,
		_w6274_
	);
	LUT2 #(
		.INIT('h1)
	) name4767 (
		_w6261_,
		_w6274_,
		_w6275_
	);
	LUT2 #(
		.INIT('h2)
	) name4768 (
		_w1976_,
		_w6275_,
		_w6276_
	);
	LUT2 #(
		.INIT('h2)
	) name4769 (
		\WX8549_reg/NET0131 ,
		\WX8613_reg/NET0131 ,
		_w6277_
	);
	LUT2 #(
		.INIT('h4)
	) name4770 (
		\WX8549_reg/NET0131 ,
		\WX8613_reg/NET0131 ,
		_w6278_
	);
	LUT2 #(
		.INIT('h1)
	) name4771 (
		_w6277_,
		_w6278_,
		_w6279_
	);
	LUT2 #(
		.INIT('h2)
	) name4772 (
		\WX8485_reg/NET0131 ,
		_w6279_,
		_w6280_
	);
	LUT2 #(
		.INIT('h4)
	) name4773 (
		\WX8485_reg/NET0131 ,
		_w6279_,
		_w6281_
	);
	LUT2 #(
		.INIT('h1)
	) name4774 (
		_w6280_,
		_w6281_,
		_w6282_
	);
	LUT2 #(
		.INIT('h2)
	) name4775 (
		\TM1_pad ,
		\WX8421_reg/NET0131 ,
		_w6283_
	);
	LUT2 #(
		.INIT('h4)
	) name4776 (
		\TM1_pad ,
		\WX8421_reg/NET0131 ,
		_w6284_
	);
	LUT2 #(
		.INIT('h1)
	) name4777 (
		_w6283_,
		_w6284_,
		_w6285_
	);
	LUT2 #(
		.INIT('h4)
	) name4778 (
		_w6282_,
		_w6285_,
		_w6286_
	);
	LUT2 #(
		.INIT('h2)
	) name4779 (
		_w6282_,
		_w6285_,
		_w6287_
	);
	LUT2 #(
		.INIT('h1)
	) name4780 (
		\TM0_pad ,
		_w6286_,
		_w6288_
	);
	LUT2 #(
		.INIT('h4)
	) name4781 (
		_w6287_,
		_w6288_,
		_w6289_
	);
	LUT2 #(
		.INIT('h1)
	) name4782 (
		_w1714_,
		_w6289_,
		_w6290_
	);
	LUT2 #(
		.INIT('h2)
	) name4783 (
		_w1973_,
		_w6290_,
		_w6291_
	);
	LUT2 #(
		.INIT('h1)
	) name4784 (
		_w6276_,
		_w6291_,
		_w6292_
	);
	LUT2 #(
		.INIT('h8)
	) name4785 (
		\TM0_pad ,
		\_2290__reg/NET0131 ,
		_w6293_
	);
	LUT2 #(
		.INIT('h2)
	) name4786 (
		\WX9844_reg/NET0131 ,
		\WX9908_reg/NET0131 ,
		_w6294_
	);
	LUT2 #(
		.INIT('h4)
	) name4787 (
		\WX9844_reg/NET0131 ,
		\WX9908_reg/NET0131 ,
		_w6295_
	);
	LUT2 #(
		.INIT('h1)
	) name4788 (
		_w6294_,
		_w6295_,
		_w6296_
	);
	LUT2 #(
		.INIT('h2)
	) name4789 (
		\WX9780_reg/NET0131 ,
		_w6296_,
		_w6297_
	);
	LUT2 #(
		.INIT('h4)
	) name4790 (
		\WX9780_reg/NET0131 ,
		_w6296_,
		_w6298_
	);
	LUT2 #(
		.INIT('h1)
	) name4791 (
		_w6297_,
		_w6298_,
		_w6299_
	);
	LUT2 #(
		.INIT('h2)
	) name4792 (
		\TM1_pad ,
		\WX9716_reg/NET0131 ,
		_w6300_
	);
	LUT2 #(
		.INIT('h4)
	) name4793 (
		\TM1_pad ,
		\WX9716_reg/NET0131 ,
		_w6301_
	);
	LUT2 #(
		.INIT('h1)
	) name4794 (
		_w6300_,
		_w6301_,
		_w6302_
	);
	LUT2 #(
		.INIT('h4)
	) name4795 (
		_w6299_,
		_w6302_,
		_w6303_
	);
	LUT2 #(
		.INIT('h2)
	) name4796 (
		_w6299_,
		_w6302_,
		_w6304_
	);
	LUT2 #(
		.INIT('h1)
	) name4797 (
		\TM0_pad ,
		_w6303_,
		_w6305_
	);
	LUT2 #(
		.INIT('h4)
	) name4798 (
		_w6304_,
		_w6305_,
		_w6306_
	);
	LUT2 #(
		.INIT('h1)
	) name4799 (
		_w6293_,
		_w6306_,
		_w6307_
	);
	LUT2 #(
		.INIT('h2)
	) name4800 (
		_w1976_,
		_w6307_,
		_w6308_
	);
	LUT2 #(
		.INIT('h2)
	) name4801 (
		\WX8551_reg/NET0131 ,
		\WX8615_reg/NET0131 ,
		_w6309_
	);
	LUT2 #(
		.INIT('h4)
	) name4802 (
		\WX8551_reg/NET0131 ,
		\WX8615_reg/NET0131 ,
		_w6310_
	);
	LUT2 #(
		.INIT('h1)
	) name4803 (
		_w6309_,
		_w6310_,
		_w6311_
	);
	LUT2 #(
		.INIT('h2)
	) name4804 (
		\WX8487_reg/NET0131 ,
		_w6311_,
		_w6312_
	);
	LUT2 #(
		.INIT('h4)
	) name4805 (
		\WX8487_reg/NET0131 ,
		_w6311_,
		_w6313_
	);
	LUT2 #(
		.INIT('h1)
	) name4806 (
		_w6312_,
		_w6313_,
		_w6314_
	);
	LUT2 #(
		.INIT('h2)
	) name4807 (
		\TM1_pad ,
		\WX8423_reg/NET0131 ,
		_w6315_
	);
	LUT2 #(
		.INIT('h4)
	) name4808 (
		\TM1_pad ,
		\WX8423_reg/NET0131 ,
		_w6316_
	);
	LUT2 #(
		.INIT('h1)
	) name4809 (
		_w6315_,
		_w6316_,
		_w6317_
	);
	LUT2 #(
		.INIT('h4)
	) name4810 (
		_w6314_,
		_w6317_,
		_w6318_
	);
	LUT2 #(
		.INIT('h2)
	) name4811 (
		_w6314_,
		_w6317_,
		_w6319_
	);
	LUT2 #(
		.INIT('h1)
	) name4812 (
		\TM0_pad ,
		_w6318_,
		_w6320_
	);
	LUT2 #(
		.INIT('h4)
	) name4813 (
		_w6319_,
		_w6320_,
		_w6321_
	);
	LUT2 #(
		.INIT('h1)
	) name4814 (
		_w1698_,
		_w6321_,
		_w6322_
	);
	LUT2 #(
		.INIT('h2)
	) name4815 (
		_w1973_,
		_w6322_,
		_w6323_
	);
	LUT2 #(
		.INIT('h1)
	) name4816 (
		_w6308_,
		_w6323_,
		_w6324_
	);
	LUT2 #(
		.INIT('h8)
	) name4817 (
		\TM0_pad ,
		\_2289__reg/NET0131 ,
		_w6325_
	);
	LUT2 #(
		.INIT('h1)
	) name4818 (
		_w2201_,
		_w6325_,
		_w6326_
	);
	LUT2 #(
		.INIT('h2)
	) name4819 (
		_w1976_,
		_w6326_,
		_w6327_
	);
	LUT2 #(
		.INIT('h2)
	) name4820 (
		\WX8553_reg/NET0131 ,
		\WX8617_reg/NET0131 ,
		_w6328_
	);
	LUT2 #(
		.INIT('h4)
	) name4821 (
		\WX8553_reg/NET0131 ,
		\WX8617_reg/NET0131 ,
		_w6329_
	);
	LUT2 #(
		.INIT('h1)
	) name4822 (
		_w6328_,
		_w6329_,
		_w6330_
	);
	LUT2 #(
		.INIT('h2)
	) name4823 (
		\WX8489_reg/NET0131 ,
		_w6330_,
		_w6331_
	);
	LUT2 #(
		.INIT('h4)
	) name4824 (
		\WX8489_reg/NET0131 ,
		_w6330_,
		_w6332_
	);
	LUT2 #(
		.INIT('h1)
	) name4825 (
		_w6331_,
		_w6332_,
		_w6333_
	);
	LUT2 #(
		.INIT('h2)
	) name4826 (
		\TM1_pad ,
		\WX8425_reg/NET0131 ,
		_w6334_
	);
	LUT2 #(
		.INIT('h4)
	) name4827 (
		\TM1_pad ,
		\WX8425_reg/NET0131 ,
		_w6335_
	);
	LUT2 #(
		.INIT('h1)
	) name4828 (
		_w6334_,
		_w6335_,
		_w6336_
	);
	LUT2 #(
		.INIT('h4)
	) name4829 (
		_w6333_,
		_w6336_,
		_w6337_
	);
	LUT2 #(
		.INIT('h2)
	) name4830 (
		_w6333_,
		_w6336_,
		_w6338_
	);
	LUT2 #(
		.INIT('h1)
	) name4831 (
		\TM0_pad ,
		_w6337_,
		_w6339_
	);
	LUT2 #(
		.INIT('h4)
	) name4832 (
		_w6338_,
		_w6339_,
		_w6340_
	);
	LUT2 #(
		.INIT('h1)
	) name4833 (
		_w1682_,
		_w6340_,
		_w6341_
	);
	LUT2 #(
		.INIT('h2)
	) name4834 (
		_w1973_,
		_w6341_,
		_w6342_
	);
	LUT2 #(
		.INIT('h1)
	) name4835 (
		_w6327_,
		_w6342_,
		_w6343_
	);
	LUT2 #(
		.INIT('h8)
	) name4836 (
		\TM0_pad ,
		\_2325__reg/NET0131 ,
		_w6344_
	);
	LUT2 #(
		.INIT('h1)
	) name4837 (
		_w3324_,
		_w6344_,
		_w6345_
	);
	LUT2 #(
		.INIT('h2)
	) name4838 (
		_w1976_,
		_w6345_,
		_w6346_
	);
	LUT2 #(
		.INIT('h1)
	) name4839 (
		_w1746_,
		_w6098_,
		_w6347_
	);
	LUT2 #(
		.INIT('h2)
	) name4840 (
		_w1973_,
		_w6347_,
		_w6348_
	);
	LUT2 #(
		.INIT('h1)
	) name4841 (
		_w6346_,
		_w6348_,
		_w6349_
	);
	LUT2 #(
		.INIT('h8)
	) name4842 (
		\TM0_pad ,
		\_2324__reg/NET0131 ,
		_w6350_
	);
	LUT2 #(
		.INIT('h1)
	) name4843 (
		_w3474_,
		_w6350_,
		_w6351_
	);
	LUT2 #(
		.INIT('h2)
	) name4844 (
		_w1976_,
		_w6351_,
		_w6352_
	);
	LUT2 #(
		.INIT('h1)
	) name4845 (
		_w1730_,
		_w6255_,
		_w6353_
	);
	LUT2 #(
		.INIT('h2)
	) name4846 (
		_w1973_,
		_w6353_,
		_w6354_
	);
	LUT2 #(
		.INIT('h1)
	) name4847 (
		_w6352_,
		_w6354_,
		_w6355_
	);
	LUT2 #(
		.INIT('h8)
	) name4848 (
		\TM0_pad ,
		\_2323__reg/NET0131 ,
		_w6356_
	);
	LUT2 #(
		.INIT('h1)
	) name4849 (
		_w3635_,
		_w6356_,
		_w6357_
	);
	LUT2 #(
		.INIT('h2)
	) name4850 (
		_w1976_,
		_w6357_,
		_w6358_
	);
	LUT2 #(
		.INIT('h1)
	) name4851 (
		_w1714_,
		_w6274_,
		_w6359_
	);
	LUT2 #(
		.INIT('h2)
	) name4852 (
		_w1973_,
		_w6359_,
		_w6360_
	);
	LUT2 #(
		.INIT('h1)
	) name4853 (
		_w6358_,
		_w6360_,
		_w6361_
	);
	LUT2 #(
		.INIT('h8)
	) name4854 (
		\TM0_pad ,
		\_2322__reg/NET0131 ,
		_w6362_
	);
	LUT2 #(
		.INIT('h1)
	) name4855 (
		_w3796_,
		_w6362_,
		_w6363_
	);
	LUT2 #(
		.INIT('h2)
	) name4856 (
		_w1976_,
		_w6363_,
		_w6364_
	);
	LUT2 #(
		.INIT('h1)
	) name4857 (
		_w1698_,
		_w6306_,
		_w6365_
	);
	LUT2 #(
		.INIT('h2)
	) name4858 (
		_w1973_,
		_w6365_,
		_w6366_
	);
	LUT2 #(
		.INIT('h1)
	) name4859 (
		_w6364_,
		_w6366_,
		_w6367_
	);
	LUT2 #(
		.INIT('h8)
	) name4860 (
		\TM0_pad ,
		\_2193__reg/NET0131 ,
		_w6368_
	);
	LUT2 #(
		.INIT('h2)
	) name4861 (
		\WX5967_reg/NET0131 ,
		\WX6031_reg/NET0131 ,
		_w6369_
	);
	LUT2 #(
		.INIT('h4)
	) name4862 (
		\WX5967_reg/NET0131 ,
		\WX6031_reg/NET0131 ,
		_w6370_
	);
	LUT2 #(
		.INIT('h1)
	) name4863 (
		_w6369_,
		_w6370_,
		_w6371_
	);
	LUT2 #(
		.INIT('h2)
	) name4864 (
		\WX5903_reg/NET0131 ,
		_w6371_,
		_w6372_
	);
	LUT2 #(
		.INIT('h4)
	) name4865 (
		\WX5903_reg/NET0131 ,
		_w6371_,
		_w6373_
	);
	LUT2 #(
		.INIT('h1)
	) name4866 (
		_w6372_,
		_w6373_,
		_w6374_
	);
	LUT2 #(
		.INIT('h2)
	) name4867 (
		\TM1_pad ,
		\WX5839_reg/NET0131 ,
		_w6375_
	);
	LUT2 #(
		.INIT('h4)
	) name4868 (
		\TM1_pad ,
		\WX5839_reg/NET0131 ,
		_w6376_
	);
	LUT2 #(
		.INIT('h1)
	) name4869 (
		_w6375_,
		_w6376_,
		_w6377_
	);
	LUT2 #(
		.INIT('h4)
	) name4870 (
		_w6374_,
		_w6377_,
		_w6378_
	);
	LUT2 #(
		.INIT('h2)
	) name4871 (
		_w6374_,
		_w6377_,
		_w6379_
	);
	LUT2 #(
		.INIT('h1)
	) name4872 (
		\TM0_pad ,
		_w6378_,
		_w6380_
	);
	LUT2 #(
		.INIT('h4)
	) name4873 (
		_w6379_,
		_w6380_,
		_w6381_
	);
	LUT2 #(
		.INIT('h1)
	) name4874 (
		_w6368_,
		_w6381_,
		_w6382_
	);
	LUT2 #(
		.INIT('h2)
	) name4875 (
		_w1976_,
		_w6382_,
		_w6383_
	);
	LUT2 #(
		.INIT('h1)
	) name4876 (
		_w1682_,
		_w6079_,
		_w6384_
	);
	LUT2 #(
		.INIT('h2)
	) name4877 (
		_w1973_,
		_w6384_,
		_w6385_
	);
	LUT2 #(
		.INIT('h1)
	) name4878 (
		_w6383_,
		_w6385_,
		_w6386_
	);
	LUT2 #(
		.INIT('h8)
	) name4879 (
		\TM0_pad ,
		\_2192__reg/NET0131 ,
		_w6387_
	);
	LUT2 #(
		.INIT('h2)
	) name4880 (
		\WX5969_reg/NET0131 ,
		\WX6033_reg/NET0131 ,
		_w6388_
	);
	LUT2 #(
		.INIT('h4)
	) name4881 (
		\WX5969_reg/NET0131 ,
		\WX6033_reg/NET0131 ,
		_w6389_
	);
	LUT2 #(
		.INIT('h1)
	) name4882 (
		_w6388_,
		_w6389_,
		_w6390_
	);
	LUT2 #(
		.INIT('h2)
	) name4883 (
		\WX5905_reg/NET0131 ,
		_w6390_,
		_w6391_
	);
	LUT2 #(
		.INIT('h4)
	) name4884 (
		\WX5905_reg/NET0131 ,
		_w6390_,
		_w6392_
	);
	LUT2 #(
		.INIT('h1)
	) name4885 (
		_w6391_,
		_w6392_,
		_w6393_
	);
	LUT2 #(
		.INIT('h2)
	) name4886 (
		\TM1_pad ,
		\WX5841_reg/NET0131 ,
		_w6394_
	);
	LUT2 #(
		.INIT('h4)
	) name4887 (
		\TM1_pad ,
		\WX5841_reg/NET0131 ,
		_w6395_
	);
	LUT2 #(
		.INIT('h1)
	) name4888 (
		_w6394_,
		_w6395_,
		_w6396_
	);
	LUT2 #(
		.INIT('h4)
	) name4889 (
		_w6393_,
		_w6396_,
		_w6397_
	);
	LUT2 #(
		.INIT('h2)
	) name4890 (
		_w6393_,
		_w6396_,
		_w6398_
	);
	LUT2 #(
		.INIT('h1)
	) name4891 (
		\TM0_pad ,
		_w6397_,
		_w6399_
	);
	LUT2 #(
		.INIT('h4)
	) name4892 (
		_w6398_,
		_w6399_,
		_w6400_
	);
	LUT2 #(
		.INIT('h1)
	) name4893 (
		_w6387_,
		_w6400_,
		_w6401_
	);
	LUT2 #(
		.INIT('h2)
	) name4894 (
		_w1976_,
		_w6401_,
		_w6402_
	);
	LUT2 #(
		.INIT('h1)
	) name4895 (
		_w1653_,
		_w6192_,
		_w6403_
	);
	LUT2 #(
		.INIT('h2)
	) name4896 (
		_w1973_,
		_w6403_,
		_w6404_
	);
	LUT2 #(
		.INIT('h1)
	) name4897 (
		_w6402_,
		_w6404_,
		_w6405_
	);
	LUT2 #(
		.INIT('h8)
	) name4898 (
		\TM0_pad ,
		\_2191__reg/NET0131 ,
		_w6406_
	);
	LUT2 #(
		.INIT('h2)
	) name4899 (
		\WX5971_reg/NET0131 ,
		\WX6035_reg/NET0131 ,
		_w6407_
	);
	LUT2 #(
		.INIT('h4)
	) name4900 (
		\WX5971_reg/NET0131 ,
		\WX6035_reg/NET0131 ,
		_w6408_
	);
	LUT2 #(
		.INIT('h1)
	) name4901 (
		_w6407_,
		_w6408_,
		_w6409_
	);
	LUT2 #(
		.INIT('h2)
	) name4902 (
		\WX5907_reg/NET0131 ,
		_w6409_,
		_w6410_
	);
	LUT2 #(
		.INIT('h4)
	) name4903 (
		\WX5907_reg/NET0131 ,
		_w6409_,
		_w6411_
	);
	LUT2 #(
		.INIT('h1)
	) name4904 (
		_w6410_,
		_w6411_,
		_w6412_
	);
	LUT2 #(
		.INIT('h2)
	) name4905 (
		\TM1_pad ,
		\WX5843_reg/NET0131 ,
		_w6413_
	);
	LUT2 #(
		.INIT('h4)
	) name4906 (
		\TM1_pad ,
		\WX5843_reg/NET0131 ,
		_w6414_
	);
	LUT2 #(
		.INIT('h1)
	) name4907 (
		_w6413_,
		_w6414_,
		_w6415_
	);
	LUT2 #(
		.INIT('h4)
	) name4908 (
		_w6412_,
		_w6415_,
		_w6416_
	);
	LUT2 #(
		.INIT('h2)
	) name4909 (
		_w6412_,
		_w6415_,
		_w6417_
	);
	LUT2 #(
		.INIT('h1)
	) name4910 (
		\TM0_pad ,
		_w6416_,
		_w6418_
	);
	LUT2 #(
		.INIT('h4)
	) name4911 (
		_w6417_,
		_w6418_,
		_w6419_
	);
	LUT2 #(
		.INIT('h1)
	) name4912 (
		_w6406_,
		_w6419_,
		_w6420_
	);
	LUT2 #(
		.INIT('h2)
	) name4913 (
		_w1976_,
		_w6420_,
		_w6421_
	);
	LUT2 #(
		.INIT('h1)
	) name4914 (
		_w1637_,
		_w6211_,
		_w6422_
	);
	LUT2 #(
		.INIT('h2)
	) name4915 (
		_w1973_,
		_w6422_,
		_w6423_
	);
	LUT2 #(
		.INIT('h1)
	) name4916 (
		_w6421_,
		_w6423_,
		_w6424_
	);
	LUT2 #(
		.INIT('h8)
	) name4917 (
		\TM0_pad ,
		\_2190__reg/NET0131 ,
		_w6425_
	);
	LUT2 #(
		.INIT('h1)
	) name4918 (
		_w2265_,
		_w6425_,
		_w6426_
	);
	LUT2 #(
		.INIT('h2)
	) name4919 (
		_w1976_,
		_w6426_,
		_w6427_
	);
	LUT2 #(
		.INIT('h1)
	) name4920 (
		_w1621_,
		_w6230_,
		_w6428_
	);
	LUT2 #(
		.INIT('h2)
	) name4921 (
		_w1973_,
		_w6428_,
		_w6429_
	);
	LUT2 #(
		.INIT('h1)
	) name4922 (
		_w6427_,
		_w6429_,
		_w6430_
	);
	LUT2 #(
		.INIT('h8)
	) name4923 (
		\TM0_pad ,
		\_2226__reg/NET0131 ,
		_w6431_
	);
	LUT2 #(
		.INIT('h2)
	) name4924 (
		\WX7258_reg/NET0131 ,
		\WX7322_reg/NET0131 ,
		_w6432_
	);
	LUT2 #(
		.INIT('h4)
	) name4925 (
		\WX7258_reg/NET0131 ,
		\WX7322_reg/NET0131 ,
		_w6433_
	);
	LUT2 #(
		.INIT('h1)
	) name4926 (
		_w6432_,
		_w6433_,
		_w6434_
	);
	LUT2 #(
		.INIT('h2)
	) name4927 (
		\WX7194_reg/NET0131 ,
		_w6434_,
		_w6435_
	);
	LUT2 #(
		.INIT('h4)
	) name4928 (
		\WX7194_reg/NET0131 ,
		_w6434_,
		_w6436_
	);
	LUT2 #(
		.INIT('h1)
	) name4929 (
		_w6435_,
		_w6436_,
		_w6437_
	);
	LUT2 #(
		.INIT('h2)
	) name4930 (
		\TM1_pad ,
		\WX7130_reg/NET0131 ,
		_w6438_
	);
	LUT2 #(
		.INIT('h4)
	) name4931 (
		\TM1_pad ,
		\WX7130_reg/NET0131 ,
		_w6439_
	);
	LUT2 #(
		.INIT('h1)
	) name4932 (
		_w6438_,
		_w6439_,
		_w6440_
	);
	LUT2 #(
		.INIT('h4)
	) name4933 (
		_w6437_,
		_w6440_,
		_w6441_
	);
	LUT2 #(
		.INIT('h2)
	) name4934 (
		_w6437_,
		_w6440_,
		_w6442_
	);
	LUT2 #(
		.INIT('h1)
	) name4935 (
		\TM0_pad ,
		_w6441_,
		_w6443_
	);
	LUT2 #(
		.INIT('h4)
	) name4936 (
		_w6442_,
		_w6443_,
		_w6444_
	);
	LUT2 #(
		.INIT('h1)
	) name4937 (
		_w6431_,
		_w6444_,
		_w6445_
	);
	LUT2 #(
		.INIT('h2)
	) name4938 (
		_w1976_,
		_w6445_,
		_w6446_
	);
	LUT2 #(
		.INIT('h1)
	) name4939 (
		_w1698_,
		_w6123_,
		_w6447_
	);
	LUT2 #(
		.INIT('h2)
	) name4940 (
		_w1973_,
		_w6447_,
		_w6448_
	);
	LUT2 #(
		.INIT('h1)
	) name4941 (
		_w6446_,
		_w6448_,
		_w6449_
	);
	LUT2 #(
		.INIT('h8)
	) name4942 (
		\TM0_pad ,
		\_2225__reg/NET0131 ,
		_w6450_
	);
	LUT2 #(
		.INIT('h2)
	) name4943 (
		\WX7260_reg/NET0131 ,
		\WX7324_reg/NET0131 ,
		_w6451_
	);
	LUT2 #(
		.INIT('h4)
	) name4944 (
		\WX7260_reg/NET0131 ,
		\WX7324_reg/NET0131 ,
		_w6452_
	);
	LUT2 #(
		.INIT('h1)
	) name4945 (
		_w6451_,
		_w6452_,
		_w6453_
	);
	LUT2 #(
		.INIT('h2)
	) name4946 (
		\WX7196_reg/NET0131 ,
		_w6453_,
		_w6454_
	);
	LUT2 #(
		.INIT('h4)
	) name4947 (
		\WX7196_reg/NET0131 ,
		_w6453_,
		_w6455_
	);
	LUT2 #(
		.INIT('h1)
	) name4948 (
		_w6454_,
		_w6455_,
		_w6456_
	);
	LUT2 #(
		.INIT('h2)
	) name4949 (
		\TM1_pad ,
		\WX7132_reg/NET0131 ,
		_w6457_
	);
	LUT2 #(
		.INIT('h4)
	) name4950 (
		\TM1_pad ,
		\WX7132_reg/NET0131 ,
		_w6458_
	);
	LUT2 #(
		.INIT('h1)
	) name4951 (
		_w6457_,
		_w6458_,
		_w6459_
	);
	LUT2 #(
		.INIT('h4)
	) name4952 (
		_w6456_,
		_w6459_,
		_w6460_
	);
	LUT2 #(
		.INIT('h2)
	) name4953 (
		_w6456_,
		_w6459_,
		_w6461_
	);
	LUT2 #(
		.INIT('h1)
	) name4954 (
		\TM0_pad ,
		_w6460_,
		_w6462_
	);
	LUT2 #(
		.INIT('h4)
	) name4955 (
		_w6461_,
		_w6462_,
		_w6463_
	);
	LUT2 #(
		.INIT('h1)
	) name4956 (
		_w6450_,
		_w6463_,
		_w6464_
	);
	LUT2 #(
		.INIT('h2)
	) name4957 (
		_w1976_,
		_w6464_,
		_w6465_
	);
	LUT2 #(
		.INIT('h1)
	) name4958 (
		_w1682_,
		_w6381_,
		_w6466_
	);
	LUT2 #(
		.INIT('h2)
	) name4959 (
		_w1973_,
		_w6466_,
		_w6467_
	);
	LUT2 #(
		.INIT('h1)
	) name4960 (
		_w6465_,
		_w6467_,
		_w6468_
	);
	LUT2 #(
		.INIT('h8)
	) name4961 (
		\TM0_pad ,
		\_2224__reg/NET0131 ,
		_w6469_
	);
	LUT2 #(
		.INIT('h2)
	) name4962 (
		\WX7262_reg/NET0131 ,
		\WX7326_reg/NET0131 ,
		_w6470_
	);
	LUT2 #(
		.INIT('h4)
	) name4963 (
		\WX7262_reg/NET0131 ,
		\WX7326_reg/NET0131 ,
		_w6471_
	);
	LUT2 #(
		.INIT('h1)
	) name4964 (
		_w6470_,
		_w6471_,
		_w6472_
	);
	LUT2 #(
		.INIT('h2)
	) name4965 (
		\WX7198_reg/NET0131 ,
		_w6472_,
		_w6473_
	);
	LUT2 #(
		.INIT('h4)
	) name4966 (
		\WX7198_reg/NET0131 ,
		_w6472_,
		_w6474_
	);
	LUT2 #(
		.INIT('h1)
	) name4967 (
		_w6473_,
		_w6474_,
		_w6475_
	);
	LUT2 #(
		.INIT('h2)
	) name4968 (
		\TM1_pad ,
		\WX7134_reg/NET0131 ,
		_w6476_
	);
	LUT2 #(
		.INIT('h4)
	) name4969 (
		\TM1_pad ,
		\WX7134_reg/NET0131 ,
		_w6477_
	);
	LUT2 #(
		.INIT('h1)
	) name4970 (
		_w6476_,
		_w6477_,
		_w6478_
	);
	LUT2 #(
		.INIT('h4)
	) name4971 (
		_w6475_,
		_w6478_,
		_w6479_
	);
	LUT2 #(
		.INIT('h2)
	) name4972 (
		_w6475_,
		_w6478_,
		_w6480_
	);
	LUT2 #(
		.INIT('h1)
	) name4973 (
		\TM0_pad ,
		_w6479_,
		_w6481_
	);
	LUT2 #(
		.INIT('h4)
	) name4974 (
		_w6480_,
		_w6481_,
		_w6482_
	);
	LUT2 #(
		.INIT('h1)
	) name4975 (
		_w6469_,
		_w6482_,
		_w6483_
	);
	LUT2 #(
		.INIT('h2)
	) name4976 (
		_w1976_,
		_w6483_,
		_w6484_
	);
	LUT2 #(
		.INIT('h1)
	) name4977 (
		_w1653_,
		_w6400_,
		_w6485_
	);
	LUT2 #(
		.INIT('h2)
	) name4978 (
		_w1973_,
		_w6485_,
		_w6486_
	);
	LUT2 #(
		.INIT('h1)
	) name4979 (
		_w6484_,
		_w6486_,
		_w6487_
	);
	LUT2 #(
		.INIT('h8)
	) name4980 (
		\TM0_pad ,
		\_2223__reg/NET0131 ,
		_w6488_
	);
	LUT2 #(
		.INIT('h1)
	) name4981 (
		_w2297_,
		_w6488_,
		_w6489_
	);
	LUT2 #(
		.INIT('h2)
	) name4982 (
		_w1976_,
		_w6489_,
		_w6490_
	);
	LUT2 #(
		.INIT('h1)
	) name4983 (
		_w1637_,
		_w6419_,
		_w6491_
	);
	LUT2 #(
		.INIT('h2)
	) name4984 (
		_w1973_,
		_w6491_,
		_w6492_
	);
	LUT2 #(
		.INIT('h1)
	) name4985 (
		_w6490_,
		_w6492_,
		_w6493_
	);
	LUT2 #(
		.INIT('h2)
	) name4986 (
		_w4239_,
		_w6032_,
		_w6494_
	);
	LUT2 #(
		.INIT('h2)
	) name4987 (
		\TM0_pad ,
		\_2111__reg/NET0131 ,
		_w6495_
	);
	LUT2 #(
		.INIT('h2)
	) name4988 (
		_w1976_,
		_w6495_,
		_w6496_
	);
	LUT2 #(
		.INIT('h4)
	) name4989 (
		_w4249_,
		_w6496_,
		_w6497_
	);
	LUT2 #(
		.INIT('h1)
	) name4990 (
		_w6494_,
		_w6497_,
		_w6498_
	);
	LUT2 #(
		.INIT('h2)
	) name4991 (
		\WX2126_reg/NET0131 ,
		\WX2190_reg/NET0131 ,
		_w6499_
	);
	LUT2 #(
		.INIT('h4)
	) name4992 (
		\WX2126_reg/NET0131 ,
		\WX2190_reg/NET0131 ,
		_w6500_
	);
	LUT2 #(
		.INIT('h1)
	) name4993 (
		_w6499_,
		_w6500_,
		_w6501_
	);
	LUT2 #(
		.INIT('h2)
	) name4994 (
		\WX1998_reg/NET0131 ,
		\WX2062_reg/NET0131 ,
		_w6502_
	);
	LUT2 #(
		.INIT('h4)
	) name4995 (
		\WX1998_reg/NET0131 ,
		\WX2062_reg/NET0131 ,
		_w6503_
	);
	LUT2 #(
		.INIT('h1)
	) name4996 (
		_w6502_,
		_w6503_,
		_w6504_
	);
	LUT2 #(
		.INIT('h4)
	) name4997 (
		_w6501_,
		_w6504_,
		_w6505_
	);
	LUT2 #(
		.INIT('h2)
	) name4998 (
		_w6501_,
		_w6504_,
		_w6506_
	);
	LUT2 #(
		.INIT('h1)
	) name4999 (
		\TM0_pad ,
		_w6505_,
		_w6507_
	);
	LUT2 #(
		.INIT('h4)
	) name5000 (
		_w6506_,
		_w6507_,
		_w6508_
	);
	LUT2 #(
		.INIT('h2)
	) name5001 (
		_w4382_,
		_w6508_,
		_w6509_
	);
	LUT2 #(
		.INIT('h2)
	) name5002 (
		\TM0_pad ,
		\_2110__reg/NET0131 ,
		_w6510_
	);
	LUT2 #(
		.INIT('h2)
	) name5003 (
		_w1976_,
		_w6510_,
		_w6511_
	);
	LUT2 #(
		.INIT('h4)
	) name5004 (
		_w4392_,
		_w6511_,
		_w6512_
	);
	LUT2 #(
		.INIT('h1)
	) name5005 (
		_w6509_,
		_w6512_,
		_w6513_
	);
	LUT2 #(
		.INIT('h2)
	) name5006 (
		_w4510_,
		_w6048_,
		_w6514_
	);
	LUT2 #(
		.INIT('h2)
	) name5007 (
		\TM0_pad ,
		\_2109__reg/NET0131 ,
		_w6515_
	);
	LUT2 #(
		.INIT('h2)
	) name5008 (
		_w1976_,
		_w6515_,
		_w6516_
	);
	LUT2 #(
		.INIT('h4)
	) name5009 (
		_w4520_,
		_w6516_,
		_w6517_
	);
	LUT2 #(
		.INIT('h1)
	) name5010 (
		_w6514_,
		_w6517_,
		_w6518_
	);
	LUT2 #(
		.INIT('h8)
	) name5011 (
		\TM0_pad ,
		\_2259__reg/NET0131 ,
		_w6519_
	);
	LUT2 #(
		.INIT('h1)
	) name5012 (
		_w6289_,
		_w6519_,
		_w6520_
	);
	LUT2 #(
		.INIT('h2)
	) name5013 (
		_w1976_,
		_w6520_,
		_w6521_
	);
	LUT2 #(
		.INIT('h1)
	) name5014 (
		_w1714_,
		_w6142_,
		_w6522_
	);
	LUT2 #(
		.INIT('h2)
	) name5015 (
		_w1973_,
		_w6522_,
		_w6523_
	);
	LUT2 #(
		.INIT('h1)
	) name5016 (
		_w6521_,
		_w6523_,
		_w6524_
	);
	LUT2 #(
		.INIT('h8)
	) name5017 (
		\TM0_pad ,
		\_2258__reg/NET0131 ,
		_w6525_
	);
	LUT2 #(
		.INIT('h1)
	) name5018 (
		_w6321_,
		_w6525_,
		_w6526_
	);
	LUT2 #(
		.INIT('h2)
	) name5019 (
		_w1976_,
		_w6526_,
		_w6527_
	);
	LUT2 #(
		.INIT('h1)
	) name5020 (
		_w1698_,
		_w6444_,
		_w6528_
	);
	LUT2 #(
		.INIT('h2)
	) name5021 (
		_w1973_,
		_w6528_,
		_w6529_
	);
	LUT2 #(
		.INIT('h1)
	) name5022 (
		_w6527_,
		_w6529_,
		_w6530_
	);
	LUT2 #(
		.INIT('h8)
	) name5023 (
		\TM0_pad ,
		\_2257__reg/NET0131 ,
		_w6531_
	);
	LUT2 #(
		.INIT('h1)
	) name5024 (
		_w6340_,
		_w6531_,
		_w6532_
	);
	LUT2 #(
		.INIT('h2)
	) name5025 (
		_w1976_,
		_w6532_,
		_w6533_
	);
	LUT2 #(
		.INIT('h1)
	) name5026 (
		_w1682_,
		_w6463_,
		_w6534_
	);
	LUT2 #(
		.INIT('h2)
	) name5027 (
		_w1973_,
		_w6534_,
		_w6535_
	);
	LUT2 #(
		.INIT('h1)
	) name5028 (
		_w6533_,
		_w6535_,
		_w6536_
	);
	LUT2 #(
		.INIT('h8)
	) name5029 (
		\TM0_pad ,
		\_2256__reg/NET0131 ,
		_w6537_
	);
	LUT2 #(
		.INIT('h1)
	) name5030 (
		_w2169_,
		_w6537_,
		_w6538_
	);
	LUT2 #(
		.INIT('h2)
	) name5031 (
		_w1976_,
		_w6538_,
		_w6539_
	);
	LUT2 #(
		.INIT('h1)
	) name5032 (
		_w1653_,
		_w6482_,
		_w6540_
	);
	LUT2 #(
		.INIT('h2)
	) name5033 (
		_w1973_,
		_w6540_,
		_w6541_
	);
	LUT2 #(
		.INIT('h1)
	) name5034 (
		_w6539_,
		_w6541_,
		_w6542_
	);
	LUT2 #(
		.INIT('h2)
	) name5035 (
		_w4239_,
		_w4927_,
		_w6543_
	);
	LUT2 #(
		.INIT('h1)
	) name5036 (
		\DATA_0_2_pad ,
		\TM0_pad ,
		_w6544_
	);
	LUT2 #(
		.INIT('h2)
	) name5037 (
		\TM0_pad ,
		\_2335__reg/NET0131 ,
		_w6545_
	);
	LUT2 #(
		.INIT('h2)
	) name5038 (
		_w1976_,
		_w6544_,
		_w6546_
	);
	LUT2 #(
		.INIT('h4)
	) name5039 (
		_w6545_,
		_w6546_,
		_w6547_
	);
	LUT2 #(
		.INIT('h1)
	) name5040 (
		_w6543_,
		_w6547_,
		_w6548_
	);
	LUT2 #(
		.INIT('h2)
	) name5041 (
		_w4382_,
		_w5042_,
		_w6549_
	);
	LUT2 #(
		.INIT('h1)
	) name5042 (
		\DATA_0_1_pad ,
		\TM0_pad ,
		_w6550_
	);
	LUT2 #(
		.INIT('h2)
	) name5043 (
		\TM0_pad ,
		\_2334__reg/NET0131 ,
		_w6551_
	);
	LUT2 #(
		.INIT('h2)
	) name5044 (
		_w1976_,
		_w6550_,
		_w6552_
	);
	LUT2 #(
		.INIT('h4)
	) name5045 (
		_w6551_,
		_w6552_,
		_w6553_
	);
	LUT2 #(
		.INIT('h1)
	) name5046 (
		_w6549_,
		_w6553_,
		_w6554_
	);
	LUT2 #(
		.INIT('h2)
	) name5047 (
		_w4510_,
		_w5174_,
		_w6555_
	);
	LUT2 #(
		.INIT('h1)
	) name5048 (
		\DATA_0_0_pad ,
		\TM0_pad ,
		_w6556_
	);
	LUT2 #(
		.INIT('h2)
	) name5049 (
		\TM0_pad ,
		\_2333__reg/NET0131 ,
		_w6557_
	);
	LUT2 #(
		.INIT('h2)
	) name5050 (
		_w1976_,
		_w6556_,
		_w6558_
	);
	LUT2 #(
		.INIT('h4)
	) name5051 (
		_w6557_,
		_w6558_,
		_w6559_
	);
	LUT2 #(
		.INIT('h1)
	) name5052 (
		_w6555_,
		_w6559_,
		_w6560_
	);
	LUT2 #(
		.INIT('h8)
	) name5053 (
		RESET_pad,
		\WX10885_reg/NET0131 ,
		_w6561_
	);
	LUT2 #(
		.INIT('h1)
	) name5054 (
		\WX837_reg/NET0131 ,
		\_2107__reg/NET0131 ,
		_w6562_
	);
	LUT2 #(
		.INIT('h8)
	) name5055 (
		\WX837_reg/NET0131 ,
		\_2107__reg/NET0131 ,
		_w6563_
	);
	LUT2 #(
		.INIT('h1)
	) name5056 (
		_w6562_,
		_w6563_,
		_w6564_
	);
	LUT2 #(
		.INIT('h2)
	) name5057 (
		RESET_pad,
		_w6564_,
		_w6565_
	);
	LUT2 #(
		.INIT('h1)
	) name5058 (
		\WX2130_reg/NET0131 ,
		\_2139__reg/NET0131 ,
		_w6566_
	);
	LUT2 #(
		.INIT('h8)
	) name5059 (
		\WX2130_reg/NET0131 ,
		\_2139__reg/NET0131 ,
		_w6567_
	);
	LUT2 #(
		.INIT('h1)
	) name5060 (
		_w6566_,
		_w6567_,
		_w6568_
	);
	LUT2 #(
		.INIT('h2)
	) name5061 (
		RESET_pad,
		_w6568_,
		_w6569_
	);
	LUT2 #(
		.INIT('h1)
	) name5062 (
		\WX11181_reg/NET0131 ,
		\_2363__reg/NET0131 ,
		_w6570_
	);
	LUT2 #(
		.INIT('h8)
	) name5063 (
		\WX11181_reg/NET0131 ,
		\_2363__reg/NET0131 ,
		_w6571_
	);
	LUT2 #(
		.INIT('h1)
	) name5064 (
		_w6570_,
		_w6571_,
		_w6572_
	);
	LUT2 #(
		.INIT('h2)
	) name5065 (
		RESET_pad,
		_w6572_,
		_w6573_
	);
	LUT2 #(
		.INIT('h8)
	) name5066 (
		RESET_pad,
		\WX10887_reg/NET0131 ,
		_w6574_
	);
	LUT2 #(
		.INIT('h1)
	) name5067 (
		\WX891_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w6575_
	);
	LUT2 #(
		.INIT('h8)
	) name5068 (
		\WX891_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w6576_
	);
	LUT2 #(
		.INIT('h1)
	) name5069 (
		_w6575_,
		_w6576_,
		_w6577_
	);
	LUT2 #(
		.INIT('h2)
	) name5070 (
		\_2080__reg/NET0131 ,
		_w6577_,
		_w6578_
	);
	LUT2 #(
		.INIT('h4)
	) name5071 (
		\_2080__reg/NET0131 ,
		_w6577_,
		_w6579_
	);
	LUT2 #(
		.INIT('h2)
	) name5072 (
		RESET_pad,
		_w6578_,
		_w6580_
	);
	LUT2 #(
		.INIT('h4)
	) name5073 (
		_w6579_,
		_w6580_,
		_w6581_
	);
	LUT2 #(
		.INIT('h1)
	) name5074 (
		\WX877_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w6582_
	);
	LUT2 #(
		.INIT('h8)
	) name5075 (
		\WX877_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w6583_
	);
	LUT2 #(
		.INIT('h1)
	) name5076 (
		_w6582_,
		_w6583_,
		_w6584_
	);
	LUT2 #(
		.INIT('h2)
	) name5077 (
		\_2087__reg/NET0131 ,
		_w6584_,
		_w6585_
	);
	LUT2 #(
		.INIT('h4)
	) name5078 (
		\_2087__reg/NET0131 ,
		_w6584_,
		_w6586_
	);
	LUT2 #(
		.INIT('h2)
	) name5079 (
		RESET_pad,
		_w6585_,
		_w6587_
	);
	LUT2 #(
		.INIT('h4)
	) name5080 (
		_w6586_,
		_w6587_,
		_w6588_
	);
	LUT2 #(
		.INIT('h1)
	) name5081 (
		\WX867_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w6589_
	);
	LUT2 #(
		.INIT('h8)
	) name5082 (
		\WX867_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w6590_
	);
	LUT2 #(
		.INIT('h1)
	) name5083 (
		_w6589_,
		_w6590_,
		_w6591_
	);
	LUT2 #(
		.INIT('h2)
	) name5084 (
		\_2092__reg/NET0131 ,
		_w6591_,
		_w6592_
	);
	LUT2 #(
		.INIT('h4)
	) name5085 (
		\_2092__reg/NET0131 ,
		_w6591_,
		_w6593_
	);
	LUT2 #(
		.INIT('h2)
	) name5086 (
		RESET_pad,
		_w6592_,
		_w6594_
	);
	LUT2 #(
		.INIT('h4)
	) name5087 (
		_w6593_,
		_w6594_,
		_w6595_
	);
	LUT2 #(
		.INIT('h1)
	) name5088 (
		\WX2184_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w6596_
	);
	LUT2 #(
		.INIT('h8)
	) name5089 (
		\WX2184_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w6597_
	);
	LUT2 #(
		.INIT('h1)
	) name5090 (
		_w6596_,
		_w6597_,
		_w6598_
	);
	LUT2 #(
		.INIT('h2)
	) name5091 (
		\_2112__reg/NET0131 ,
		_w6598_,
		_w6599_
	);
	LUT2 #(
		.INIT('h4)
	) name5092 (
		\_2112__reg/NET0131 ,
		_w6598_,
		_w6600_
	);
	LUT2 #(
		.INIT('h2)
	) name5093 (
		RESET_pad,
		_w6599_,
		_w6601_
	);
	LUT2 #(
		.INIT('h4)
	) name5094 (
		_w6600_,
		_w6601_,
		_w6602_
	);
	LUT2 #(
		.INIT('h1)
	) name5095 (
		\WX2170_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w6603_
	);
	LUT2 #(
		.INIT('h8)
	) name5096 (
		\WX2170_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w6604_
	);
	LUT2 #(
		.INIT('h1)
	) name5097 (
		_w6603_,
		_w6604_,
		_w6605_
	);
	LUT2 #(
		.INIT('h2)
	) name5098 (
		\_2119__reg/NET0131 ,
		_w6605_,
		_w6606_
	);
	LUT2 #(
		.INIT('h4)
	) name5099 (
		\_2119__reg/NET0131 ,
		_w6605_,
		_w6607_
	);
	LUT2 #(
		.INIT('h2)
	) name5100 (
		RESET_pad,
		_w6606_,
		_w6608_
	);
	LUT2 #(
		.INIT('h4)
	) name5101 (
		_w6607_,
		_w6608_,
		_w6609_
	);
	LUT2 #(
		.INIT('h1)
	) name5102 (
		\WX2160_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w6610_
	);
	LUT2 #(
		.INIT('h8)
	) name5103 (
		\WX2160_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w6611_
	);
	LUT2 #(
		.INIT('h1)
	) name5104 (
		_w6610_,
		_w6611_,
		_w6612_
	);
	LUT2 #(
		.INIT('h2)
	) name5105 (
		\_2124__reg/NET0131 ,
		_w6612_,
		_w6613_
	);
	LUT2 #(
		.INIT('h4)
	) name5106 (
		\_2124__reg/NET0131 ,
		_w6612_,
		_w6614_
	);
	LUT2 #(
		.INIT('h2)
	) name5107 (
		RESET_pad,
		_w6613_,
		_w6615_
	);
	LUT2 #(
		.INIT('h4)
	) name5108 (
		_w6614_,
		_w6615_,
		_w6616_
	);
	LUT2 #(
		.INIT('h1)
	) name5109 (
		\WX3477_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w6617_
	);
	LUT2 #(
		.INIT('h8)
	) name5110 (
		\WX3477_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w6618_
	);
	LUT2 #(
		.INIT('h1)
	) name5111 (
		_w6617_,
		_w6618_,
		_w6619_
	);
	LUT2 #(
		.INIT('h2)
	) name5112 (
		\_2144__reg/NET0131 ,
		_w6619_,
		_w6620_
	);
	LUT2 #(
		.INIT('h4)
	) name5113 (
		\_2144__reg/NET0131 ,
		_w6619_,
		_w6621_
	);
	LUT2 #(
		.INIT('h2)
	) name5114 (
		RESET_pad,
		_w6620_,
		_w6622_
	);
	LUT2 #(
		.INIT('h4)
	) name5115 (
		_w6621_,
		_w6622_,
		_w6623_
	);
	LUT2 #(
		.INIT('h1)
	) name5116 (
		\WX3463_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w6624_
	);
	LUT2 #(
		.INIT('h8)
	) name5117 (
		\WX3463_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w6625_
	);
	LUT2 #(
		.INIT('h1)
	) name5118 (
		_w6624_,
		_w6625_,
		_w6626_
	);
	LUT2 #(
		.INIT('h2)
	) name5119 (
		\_2151__reg/NET0131 ,
		_w6626_,
		_w6627_
	);
	LUT2 #(
		.INIT('h4)
	) name5120 (
		\_2151__reg/NET0131 ,
		_w6626_,
		_w6628_
	);
	LUT2 #(
		.INIT('h2)
	) name5121 (
		RESET_pad,
		_w6627_,
		_w6629_
	);
	LUT2 #(
		.INIT('h4)
	) name5122 (
		_w6628_,
		_w6629_,
		_w6630_
	);
	LUT2 #(
		.INIT('h1)
	) name5123 (
		\WX3453_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w6631_
	);
	LUT2 #(
		.INIT('h8)
	) name5124 (
		\WX3453_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w6632_
	);
	LUT2 #(
		.INIT('h1)
	) name5125 (
		_w6631_,
		_w6632_,
		_w6633_
	);
	LUT2 #(
		.INIT('h2)
	) name5126 (
		\_2156__reg/NET0131 ,
		_w6633_,
		_w6634_
	);
	LUT2 #(
		.INIT('h4)
	) name5127 (
		\_2156__reg/NET0131 ,
		_w6633_,
		_w6635_
	);
	LUT2 #(
		.INIT('h2)
	) name5128 (
		RESET_pad,
		_w6634_,
		_w6636_
	);
	LUT2 #(
		.INIT('h4)
	) name5129 (
		_w6635_,
		_w6636_,
		_w6637_
	);
	LUT2 #(
		.INIT('h1)
	) name5130 (
		\WX4770_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w6638_
	);
	LUT2 #(
		.INIT('h8)
	) name5131 (
		\WX4770_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w6639_
	);
	LUT2 #(
		.INIT('h1)
	) name5132 (
		_w6638_,
		_w6639_,
		_w6640_
	);
	LUT2 #(
		.INIT('h2)
	) name5133 (
		\_2176__reg/NET0131 ,
		_w6640_,
		_w6641_
	);
	LUT2 #(
		.INIT('h4)
	) name5134 (
		\_2176__reg/NET0131 ,
		_w6640_,
		_w6642_
	);
	LUT2 #(
		.INIT('h2)
	) name5135 (
		RESET_pad,
		_w6641_,
		_w6643_
	);
	LUT2 #(
		.INIT('h4)
	) name5136 (
		_w6642_,
		_w6643_,
		_w6644_
	);
	LUT2 #(
		.INIT('h1)
	) name5137 (
		\WX4756_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w6645_
	);
	LUT2 #(
		.INIT('h8)
	) name5138 (
		\WX4756_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w6646_
	);
	LUT2 #(
		.INIT('h1)
	) name5139 (
		_w6645_,
		_w6646_,
		_w6647_
	);
	LUT2 #(
		.INIT('h2)
	) name5140 (
		\_2183__reg/NET0131 ,
		_w6647_,
		_w6648_
	);
	LUT2 #(
		.INIT('h4)
	) name5141 (
		\_2183__reg/NET0131 ,
		_w6647_,
		_w6649_
	);
	LUT2 #(
		.INIT('h2)
	) name5142 (
		RESET_pad,
		_w6648_,
		_w6650_
	);
	LUT2 #(
		.INIT('h4)
	) name5143 (
		_w6649_,
		_w6650_,
		_w6651_
	);
	LUT2 #(
		.INIT('h1)
	) name5144 (
		\WX4746_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w6652_
	);
	LUT2 #(
		.INIT('h8)
	) name5145 (
		\WX4746_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w6653_
	);
	LUT2 #(
		.INIT('h1)
	) name5146 (
		_w6652_,
		_w6653_,
		_w6654_
	);
	LUT2 #(
		.INIT('h2)
	) name5147 (
		\_2188__reg/NET0131 ,
		_w6654_,
		_w6655_
	);
	LUT2 #(
		.INIT('h4)
	) name5148 (
		\_2188__reg/NET0131 ,
		_w6654_,
		_w6656_
	);
	LUT2 #(
		.INIT('h2)
	) name5149 (
		RESET_pad,
		_w6655_,
		_w6657_
	);
	LUT2 #(
		.INIT('h4)
	) name5150 (
		_w6656_,
		_w6657_,
		_w6658_
	);
	LUT2 #(
		.INIT('h1)
	) name5151 (
		\WX6063_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w6659_
	);
	LUT2 #(
		.INIT('h8)
	) name5152 (
		\WX6063_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w6660_
	);
	LUT2 #(
		.INIT('h1)
	) name5153 (
		_w6659_,
		_w6660_,
		_w6661_
	);
	LUT2 #(
		.INIT('h2)
	) name5154 (
		\_2208__reg/NET0131 ,
		_w6661_,
		_w6662_
	);
	LUT2 #(
		.INIT('h4)
	) name5155 (
		\_2208__reg/NET0131 ,
		_w6661_,
		_w6663_
	);
	LUT2 #(
		.INIT('h2)
	) name5156 (
		RESET_pad,
		_w6662_,
		_w6664_
	);
	LUT2 #(
		.INIT('h4)
	) name5157 (
		_w6663_,
		_w6664_,
		_w6665_
	);
	LUT2 #(
		.INIT('h1)
	) name5158 (
		\WX6049_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w6666_
	);
	LUT2 #(
		.INIT('h8)
	) name5159 (
		\WX6049_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w6667_
	);
	LUT2 #(
		.INIT('h1)
	) name5160 (
		_w6666_,
		_w6667_,
		_w6668_
	);
	LUT2 #(
		.INIT('h2)
	) name5161 (
		\_2215__reg/NET0131 ,
		_w6668_,
		_w6669_
	);
	LUT2 #(
		.INIT('h4)
	) name5162 (
		\_2215__reg/NET0131 ,
		_w6668_,
		_w6670_
	);
	LUT2 #(
		.INIT('h2)
	) name5163 (
		RESET_pad,
		_w6669_,
		_w6671_
	);
	LUT2 #(
		.INIT('h4)
	) name5164 (
		_w6670_,
		_w6671_,
		_w6672_
	);
	LUT2 #(
		.INIT('h1)
	) name5165 (
		\WX6039_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w6673_
	);
	LUT2 #(
		.INIT('h8)
	) name5166 (
		\WX6039_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w6674_
	);
	LUT2 #(
		.INIT('h1)
	) name5167 (
		_w6673_,
		_w6674_,
		_w6675_
	);
	LUT2 #(
		.INIT('h2)
	) name5168 (
		\_2220__reg/NET0131 ,
		_w6675_,
		_w6676_
	);
	LUT2 #(
		.INIT('h4)
	) name5169 (
		\_2220__reg/NET0131 ,
		_w6675_,
		_w6677_
	);
	LUT2 #(
		.INIT('h2)
	) name5170 (
		RESET_pad,
		_w6676_,
		_w6678_
	);
	LUT2 #(
		.INIT('h4)
	) name5171 (
		_w6677_,
		_w6678_,
		_w6679_
	);
	LUT2 #(
		.INIT('h1)
	) name5172 (
		\WX7356_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w6680_
	);
	LUT2 #(
		.INIT('h8)
	) name5173 (
		\WX7356_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w6681_
	);
	LUT2 #(
		.INIT('h1)
	) name5174 (
		_w6680_,
		_w6681_,
		_w6682_
	);
	LUT2 #(
		.INIT('h2)
	) name5175 (
		\_2240__reg/NET0131 ,
		_w6682_,
		_w6683_
	);
	LUT2 #(
		.INIT('h4)
	) name5176 (
		\_2240__reg/NET0131 ,
		_w6682_,
		_w6684_
	);
	LUT2 #(
		.INIT('h2)
	) name5177 (
		RESET_pad,
		_w6683_,
		_w6685_
	);
	LUT2 #(
		.INIT('h4)
	) name5178 (
		_w6684_,
		_w6685_,
		_w6686_
	);
	LUT2 #(
		.INIT('h1)
	) name5179 (
		\WX7342_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w6687_
	);
	LUT2 #(
		.INIT('h8)
	) name5180 (
		\WX7342_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w6688_
	);
	LUT2 #(
		.INIT('h1)
	) name5181 (
		_w6687_,
		_w6688_,
		_w6689_
	);
	LUT2 #(
		.INIT('h2)
	) name5182 (
		\_2247__reg/NET0131 ,
		_w6689_,
		_w6690_
	);
	LUT2 #(
		.INIT('h4)
	) name5183 (
		\_2247__reg/NET0131 ,
		_w6689_,
		_w6691_
	);
	LUT2 #(
		.INIT('h2)
	) name5184 (
		RESET_pad,
		_w6690_,
		_w6692_
	);
	LUT2 #(
		.INIT('h4)
	) name5185 (
		_w6691_,
		_w6692_,
		_w6693_
	);
	LUT2 #(
		.INIT('h1)
	) name5186 (
		\WX7332_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w6694_
	);
	LUT2 #(
		.INIT('h8)
	) name5187 (
		\WX7332_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w6695_
	);
	LUT2 #(
		.INIT('h1)
	) name5188 (
		_w6694_,
		_w6695_,
		_w6696_
	);
	LUT2 #(
		.INIT('h2)
	) name5189 (
		\_2252__reg/NET0131 ,
		_w6696_,
		_w6697_
	);
	LUT2 #(
		.INIT('h4)
	) name5190 (
		\_2252__reg/NET0131 ,
		_w6696_,
		_w6698_
	);
	LUT2 #(
		.INIT('h2)
	) name5191 (
		RESET_pad,
		_w6697_,
		_w6699_
	);
	LUT2 #(
		.INIT('h4)
	) name5192 (
		_w6698_,
		_w6699_,
		_w6700_
	);
	LUT2 #(
		.INIT('h1)
	) name5193 (
		\WX8649_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w6701_
	);
	LUT2 #(
		.INIT('h8)
	) name5194 (
		\WX8649_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w6702_
	);
	LUT2 #(
		.INIT('h1)
	) name5195 (
		_w6701_,
		_w6702_,
		_w6703_
	);
	LUT2 #(
		.INIT('h2)
	) name5196 (
		\_2272__reg/NET0131 ,
		_w6703_,
		_w6704_
	);
	LUT2 #(
		.INIT('h4)
	) name5197 (
		\_2272__reg/NET0131 ,
		_w6703_,
		_w6705_
	);
	LUT2 #(
		.INIT('h2)
	) name5198 (
		RESET_pad,
		_w6704_,
		_w6706_
	);
	LUT2 #(
		.INIT('h4)
	) name5199 (
		_w6705_,
		_w6706_,
		_w6707_
	);
	LUT2 #(
		.INIT('h1)
	) name5200 (
		\WX8635_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w6708_
	);
	LUT2 #(
		.INIT('h8)
	) name5201 (
		\WX8635_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w6709_
	);
	LUT2 #(
		.INIT('h1)
	) name5202 (
		_w6708_,
		_w6709_,
		_w6710_
	);
	LUT2 #(
		.INIT('h2)
	) name5203 (
		\_2279__reg/NET0131 ,
		_w6710_,
		_w6711_
	);
	LUT2 #(
		.INIT('h4)
	) name5204 (
		\_2279__reg/NET0131 ,
		_w6710_,
		_w6712_
	);
	LUT2 #(
		.INIT('h2)
	) name5205 (
		RESET_pad,
		_w6711_,
		_w6713_
	);
	LUT2 #(
		.INIT('h4)
	) name5206 (
		_w6712_,
		_w6713_,
		_w6714_
	);
	LUT2 #(
		.INIT('h1)
	) name5207 (
		\WX8625_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w6715_
	);
	LUT2 #(
		.INIT('h8)
	) name5208 (
		\WX8625_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w6716_
	);
	LUT2 #(
		.INIT('h1)
	) name5209 (
		_w6715_,
		_w6716_,
		_w6717_
	);
	LUT2 #(
		.INIT('h2)
	) name5210 (
		\_2284__reg/NET0131 ,
		_w6717_,
		_w6718_
	);
	LUT2 #(
		.INIT('h4)
	) name5211 (
		\_2284__reg/NET0131 ,
		_w6717_,
		_w6719_
	);
	LUT2 #(
		.INIT('h2)
	) name5212 (
		RESET_pad,
		_w6718_,
		_w6720_
	);
	LUT2 #(
		.INIT('h4)
	) name5213 (
		_w6719_,
		_w6720_,
		_w6721_
	);
	LUT2 #(
		.INIT('h1)
	) name5214 (
		\WX9942_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w6722_
	);
	LUT2 #(
		.INIT('h8)
	) name5215 (
		\WX9942_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w6723_
	);
	LUT2 #(
		.INIT('h1)
	) name5216 (
		_w6722_,
		_w6723_,
		_w6724_
	);
	LUT2 #(
		.INIT('h2)
	) name5217 (
		\_2304__reg/NET0131 ,
		_w6724_,
		_w6725_
	);
	LUT2 #(
		.INIT('h4)
	) name5218 (
		\_2304__reg/NET0131 ,
		_w6724_,
		_w6726_
	);
	LUT2 #(
		.INIT('h2)
	) name5219 (
		RESET_pad,
		_w6725_,
		_w6727_
	);
	LUT2 #(
		.INIT('h4)
	) name5220 (
		_w6726_,
		_w6727_,
		_w6728_
	);
	LUT2 #(
		.INIT('h1)
	) name5221 (
		\WX9928_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w6729_
	);
	LUT2 #(
		.INIT('h8)
	) name5222 (
		\WX9928_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w6730_
	);
	LUT2 #(
		.INIT('h1)
	) name5223 (
		_w6729_,
		_w6730_,
		_w6731_
	);
	LUT2 #(
		.INIT('h2)
	) name5224 (
		\_2311__reg/NET0131 ,
		_w6731_,
		_w6732_
	);
	LUT2 #(
		.INIT('h4)
	) name5225 (
		\_2311__reg/NET0131 ,
		_w6731_,
		_w6733_
	);
	LUT2 #(
		.INIT('h2)
	) name5226 (
		RESET_pad,
		_w6732_,
		_w6734_
	);
	LUT2 #(
		.INIT('h4)
	) name5227 (
		_w6733_,
		_w6734_,
		_w6735_
	);
	LUT2 #(
		.INIT('h1)
	) name5228 (
		\WX9918_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w6736_
	);
	LUT2 #(
		.INIT('h8)
	) name5229 (
		\WX9918_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w6737_
	);
	LUT2 #(
		.INIT('h1)
	) name5230 (
		_w6736_,
		_w6737_,
		_w6738_
	);
	LUT2 #(
		.INIT('h2)
	) name5231 (
		\_2316__reg/NET0131 ,
		_w6738_,
		_w6739_
	);
	LUT2 #(
		.INIT('h4)
	) name5232 (
		\_2316__reg/NET0131 ,
		_w6738_,
		_w6740_
	);
	LUT2 #(
		.INIT('h2)
	) name5233 (
		RESET_pad,
		_w6739_,
		_w6741_
	);
	LUT2 #(
		.INIT('h4)
	) name5234 (
		_w6740_,
		_w6741_,
		_w6742_
	);
	LUT2 #(
		.INIT('h1)
	) name5235 (
		\WX11235_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w6743_
	);
	LUT2 #(
		.INIT('h8)
	) name5236 (
		\WX11235_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w6744_
	);
	LUT2 #(
		.INIT('h1)
	) name5237 (
		_w6743_,
		_w6744_,
		_w6745_
	);
	LUT2 #(
		.INIT('h2)
	) name5238 (
		\_2336__reg/NET0131 ,
		_w6745_,
		_w6746_
	);
	LUT2 #(
		.INIT('h4)
	) name5239 (
		\_2336__reg/NET0131 ,
		_w6745_,
		_w6747_
	);
	LUT2 #(
		.INIT('h2)
	) name5240 (
		RESET_pad,
		_w6746_,
		_w6748_
	);
	LUT2 #(
		.INIT('h4)
	) name5241 (
		_w6747_,
		_w6748_,
		_w6749_
	);
	LUT2 #(
		.INIT('h1)
	) name5242 (
		\WX11221_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w6750_
	);
	LUT2 #(
		.INIT('h8)
	) name5243 (
		\WX11221_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w6751_
	);
	LUT2 #(
		.INIT('h1)
	) name5244 (
		_w6750_,
		_w6751_,
		_w6752_
	);
	LUT2 #(
		.INIT('h2)
	) name5245 (
		\_2343__reg/NET0131 ,
		_w6752_,
		_w6753_
	);
	LUT2 #(
		.INIT('h4)
	) name5246 (
		\_2343__reg/NET0131 ,
		_w6752_,
		_w6754_
	);
	LUT2 #(
		.INIT('h2)
	) name5247 (
		RESET_pad,
		_w6753_,
		_w6755_
	);
	LUT2 #(
		.INIT('h4)
	) name5248 (
		_w6754_,
		_w6755_,
		_w6756_
	);
	LUT2 #(
		.INIT('h1)
	) name5249 (
		\WX11211_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w6757_
	);
	LUT2 #(
		.INIT('h8)
	) name5250 (
		\WX11211_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w6758_
	);
	LUT2 #(
		.INIT('h1)
	) name5251 (
		_w6757_,
		_w6758_,
		_w6759_
	);
	LUT2 #(
		.INIT('h2)
	) name5252 (
		\_2348__reg/NET0131 ,
		_w6759_,
		_w6760_
	);
	LUT2 #(
		.INIT('h4)
	) name5253 (
		\_2348__reg/NET0131 ,
		_w6759_,
		_w6761_
	);
	LUT2 #(
		.INIT('h2)
	) name5254 (
		RESET_pad,
		_w6760_,
		_w6762_
	);
	LUT2 #(
		.INIT('h4)
	) name5255 (
		_w6761_,
		_w6762_,
		_w6763_
	);
	LUT2 #(
		.INIT('h8)
	) name5256 (
		RESET_pad,
		\WX11117_reg/NET0131 ,
		_w6764_
	);
	LUT2 #(
		.INIT('h8)
	) name5257 (
		RESET_pad,
		\WX773_reg/NET0131 ,
		_w6765_
	);
	LUT2 #(
		.INIT('h8)
	) name5258 (
		RESET_pad,
		\WX10889_reg/NET0131 ,
		_w6766_
	);
	LUT2 #(
		.INIT('h8)
	) name5259 (
		RESET_pad,
		\WX2066_reg/NET0131 ,
		_w6767_
	);
	LUT2 #(
		.INIT('h1)
	) name5260 (
		\WX3475_reg/NET0131 ,
		\_2145__reg/NET0131 ,
		_w6768_
	);
	LUT2 #(
		.INIT('h8)
	) name5261 (
		\WX3475_reg/NET0131 ,
		\_2145__reg/NET0131 ,
		_w6769_
	);
	LUT2 #(
		.INIT('h1)
	) name5262 (
		_w6768_,
		_w6769_,
		_w6770_
	);
	LUT2 #(
		.INIT('h2)
	) name5263 (
		RESET_pad,
		_w6770_,
		_w6771_
	);
	LUT2 #(
		.INIT('h1)
	) name5264 (
		\WX3427_reg/NET0131 ,
		\_2169__reg/NET0131 ,
		_w6772_
	);
	LUT2 #(
		.INIT('h8)
	) name5265 (
		\WX3427_reg/NET0131 ,
		\_2169__reg/NET0131 ,
		_w6773_
	);
	LUT2 #(
		.INIT('h1)
	) name5266 (
		_w6772_,
		_w6773_,
		_w6774_
	);
	LUT2 #(
		.INIT('h2)
	) name5267 (
		RESET_pad,
		_w6774_,
		_w6775_
	);
	LUT2 #(
		.INIT('h1)
	) name5268 (
		\WX2132_reg/NET0131 ,
		\_2138__reg/NET0131 ,
		_w6776_
	);
	LUT2 #(
		.INIT('h8)
	) name5269 (
		\WX2132_reg/NET0131 ,
		\_2138__reg/NET0131 ,
		_w6777_
	);
	LUT2 #(
		.INIT('h1)
	) name5270 (
		_w6776_,
		_w6777_,
		_w6778_
	);
	LUT2 #(
		.INIT('h2)
	) name5271 (
		RESET_pad,
		_w6778_,
		_w6779_
	);
	LUT2 #(
		.INIT('h1)
	) name5272 (
		\WX11215_reg/NET0131 ,
		\_2346__reg/NET0131 ,
		_w6780_
	);
	LUT2 #(
		.INIT('h8)
	) name5273 (
		\WX11215_reg/NET0131 ,
		\_2346__reg/NET0131 ,
		_w6781_
	);
	LUT2 #(
		.INIT('h1)
	) name5274 (
		_w6780_,
		_w6781_,
		_w6782_
	);
	LUT2 #(
		.INIT('h2)
	) name5275 (
		RESET_pad,
		_w6782_,
		_w6783_
	);
	LUT2 #(
		.INIT('h1)
	) name5276 (
		\WX8599_reg/NET0131 ,
		\_2297__reg/NET0131 ,
		_w6784_
	);
	LUT2 #(
		.INIT('h8)
	) name5277 (
		\WX8599_reg/NET0131 ,
		\_2297__reg/NET0131 ,
		_w6785_
	);
	LUT2 #(
		.INIT('h1)
	) name5278 (
		_w6784_,
		_w6785_,
		_w6786_
	);
	LUT2 #(
		.INIT('h2)
	) name5279 (
		RESET_pad,
		_w6786_,
		_w6787_
	);
	LUT2 #(
		.INIT('h1)
	) name5280 (
		\WX6043_reg/NET0131 ,
		\_2218__reg/NET0131 ,
		_w6788_
	);
	LUT2 #(
		.INIT('h8)
	) name5281 (
		\WX6043_reg/NET0131 ,
		\_2218__reg/NET0131 ,
		_w6789_
	);
	LUT2 #(
		.INIT('h1)
	) name5282 (
		_w6788_,
		_w6789_,
		_w6790_
	);
	LUT2 #(
		.INIT('h2)
	) name5283 (
		RESET_pad,
		_w6790_,
		_w6791_
	);
	LUT2 #(
		.INIT('h1)
	) name5284 (
		\WX3461_reg/NET0131 ,
		\_2152__reg/NET0131 ,
		_w6792_
	);
	LUT2 #(
		.INIT('h8)
	) name5285 (
		\WX3461_reg/NET0131 ,
		\_2152__reg/NET0131 ,
		_w6793_
	);
	LUT2 #(
		.INIT('h1)
	) name5286 (
		_w6792_,
		_w6793_,
		_w6794_
	);
	LUT2 #(
		.INIT('h2)
	) name5287 (
		RESET_pad,
		_w6794_,
		_w6795_
	);
	LUT2 #(
		.INIT('h1)
	) name5288 (
		\WX857_reg/NET0131 ,
		\_2097__reg/NET0131 ,
		_w6796_
	);
	LUT2 #(
		.INIT('h8)
	) name5289 (
		\WX857_reg/NET0131 ,
		\_2097__reg/NET0131 ,
		_w6797_
	);
	LUT2 #(
		.INIT('h1)
	) name5290 (
		_w6796_,
		_w6797_,
		_w6798_
	);
	LUT2 #(
		.INIT('h2)
	) name5291 (
		RESET_pad,
		_w6798_,
		_w6799_
	);
	LUT2 #(
		.INIT('h1)
	) name5292 (
		\WX9934_reg/NET0131 ,
		\_2308__reg/NET0131 ,
		_w6800_
	);
	LUT2 #(
		.INIT('h8)
	) name5293 (
		\WX9934_reg/NET0131 ,
		\_2308__reg/NET0131 ,
		_w6801_
	);
	LUT2 #(
		.INIT('h1)
	) name5294 (
		_w6800_,
		_w6801_,
		_w6802_
	);
	LUT2 #(
		.INIT('h2)
	) name5295 (
		RESET_pad,
		_w6802_,
		_w6803_
	);
	LUT2 #(
		.INIT('h1)
	) name5296 (
		\WX7312_reg/NET0131 ,
		\_2262__reg/NET0131 ,
		_w6804_
	);
	LUT2 #(
		.INIT('h8)
	) name5297 (
		\WX7312_reg/NET0131 ,
		\_2262__reg/NET0131 ,
		_w6805_
	);
	LUT2 #(
		.INIT('h1)
	) name5298 (
		_w6804_,
		_w6805_,
		_w6806_
	);
	LUT2 #(
		.INIT('h2)
	) name5299 (
		RESET_pad,
		_w6806_,
		_w6807_
	);
	LUT2 #(
		.INIT('h1)
	) name5300 (
		\WX7338_reg/NET0131 ,
		\_2249__reg/NET0131 ,
		_w6808_
	);
	LUT2 #(
		.INIT('h8)
	) name5301 (
		\WX7338_reg/NET0131 ,
		\_2249__reg/NET0131 ,
		_w6809_
	);
	LUT2 #(
		.INIT('h1)
	) name5302 (
		_w6808_,
		_w6809_,
		_w6810_
	);
	LUT2 #(
		.INIT('h2)
	) name5303 (
		RESET_pad,
		_w6810_,
		_w6811_
	);
	LUT2 #(
		.INIT('h1)
	) name5304 (
		\WX8605_reg/NET0131 ,
		\_2294__reg/NET0131 ,
		_w6812_
	);
	LUT2 #(
		.INIT('h8)
	) name5305 (
		\WX8605_reg/NET0131 ,
		\_2294__reg/NET0131 ,
		_w6813_
	);
	LUT2 #(
		.INIT('h1)
	) name5306 (
		_w6812_,
		_w6813_,
		_w6814_
	);
	LUT2 #(
		.INIT('h2)
	) name5307 (
		RESET_pad,
		_w6814_,
		_w6815_
	);
	LUT2 #(
		.INIT('h1)
	) name5308 (
		\WX8601_reg/NET0131 ,
		\_2296__reg/NET0131 ,
		_w6816_
	);
	LUT2 #(
		.INIT('h8)
	) name5309 (
		\WX8601_reg/NET0131 ,
		\_2296__reg/NET0131 ,
		_w6817_
	);
	LUT2 #(
		.INIT('h1)
	) name5310 (
		_w6816_,
		_w6817_,
		_w6818_
	);
	LUT2 #(
		.INIT('h2)
	) name5311 (
		RESET_pad,
		_w6818_,
		_w6819_
	);
	LUT2 #(
		.INIT('h1)
	) name5312 (
		\WX8603_reg/NET0131 ,
		\_2295__reg/NET0131 ,
		_w6820_
	);
	LUT2 #(
		.INIT('h8)
	) name5313 (
		\WX8603_reg/NET0131 ,
		\_2295__reg/NET0131 ,
		_w6821_
	);
	LUT2 #(
		.INIT('h1)
	) name5314 (
		_w6820_,
		_w6821_,
		_w6822_
	);
	LUT2 #(
		.INIT('h2)
	) name5315 (
		RESET_pad,
		_w6822_,
		_w6823_
	);
	LUT2 #(
		.INIT('h1)
	) name5316 (
		\WX6037_reg/NET0131 ,
		\_2221__reg/NET0131 ,
		_w6824_
	);
	LUT2 #(
		.INIT('h8)
	) name5317 (
		\WX6037_reg/NET0131 ,
		\_2221__reg/NET0131 ,
		_w6825_
	);
	LUT2 #(
		.INIT('h1)
	) name5318 (
		_w6824_,
		_w6825_,
		_w6826_
	);
	LUT2 #(
		.INIT('h2)
	) name5319 (
		RESET_pad,
		_w6826_,
		_w6827_
	);
	LUT2 #(
		.INIT('h1)
	) name5320 (
		\WX8619_reg/NET0131 ,
		\_2287__reg/NET0131 ,
		_w6828_
	);
	LUT2 #(
		.INIT('h8)
	) name5321 (
		\WX8619_reg/NET0131 ,
		\_2287__reg/NET0131 ,
		_w6829_
	);
	LUT2 #(
		.INIT('h1)
	) name5322 (
		_w6828_,
		_w6829_,
		_w6830_
	);
	LUT2 #(
		.INIT('h2)
	) name5323 (
		RESET_pad,
		_w6830_,
		_w6831_
	);
	LUT2 #(
		.INIT('h1)
	) name5324 (
		\WX7362_reg/NET0131 ,
		\_2237__reg/NET0131 ,
		_w6832_
	);
	LUT2 #(
		.INIT('h8)
	) name5325 (
		\WX7362_reg/NET0131 ,
		\_2237__reg/NET0131 ,
		_w6833_
	);
	LUT2 #(
		.INIT('h1)
	) name5326 (
		_w6832_,
		_w6833_,
		_w6834_
	);
	LUT2 #(
		.INIT('h2)
	) name5327 (
		RESET_pad,
		_w6834_,
		_w6835_
	);
	LUT2 #(
		.INIT('h1)
	) name5328 (
		\WX3425_reg/NET0131 ,
		\_2170__reg/NET0131 ,
		_w6836_
	);
	LUT2 #(
		.INIT('h8)
	) name5329 (
		\WX3425_reg/NET0131 ,
		\_2170__reg/NET0131 ,
		_w6837_
	);
	LUT2 #(
		.INIT('h1)
	) name5330 (
		_w6836_,
		_w6837_,
		_w6838_
	);
	LUT2 #(
		.INIT('h2)
	) name5331 (
		RESET_pad,
		_w6838_,
		_w6839_
	);
	LUT2 #(
		.INIT('h1)
	) name5332 (
		\WX4728_reg/NET0131 ,
		\_2197__reg/NET0131 ,
		_w6840_
	);
	LUT2 #(
		.INIT('h8)
	) name5333 (
		\WX4728_reg/NET0131 ,
		\_2197__reg/NET0131 ,
		_w6841_
	);
	LUT2 #(
		.INIT('h1)
	) name5334 (
		_w6840_,
		_w6841_,
		_w6842_
	);
	LUT2 #(
		.INIT('h2)
	) name5335 (
		RESET_pad,
		_w6842_,
		_w6843_
	);
	LUT2 #(
		.INIT('h1)
	) name5336 (
		\WX3485_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w6844_
	);
	LUT2 #(
		.INIT('h8)
	) name5337 (
		\WX3485_reg/NET0131 ,
		\_2172__reg/NET0131 ,
		_w6845_
	);
	LUT2 #(
		.INIT('h1)
	) name5338 (
		_w6844_,
		_w6845_,
		_w6846_
	);
	LUT2 #(
		.INIT('h2)
	) name5339 (
		RESET_pad,
		_w6846_,
		_w6847_
	);
	LUT2 #(
		.INIT('h1)
	) name5340 (
		\WX7328_reg/NET0131 ,
		\_2254__reg/NET0131 ,
		_w6848_
	);
	LUT2 #(
		.INIT('h8)
	) name5341 (
		\WX7328_reg/NET0131 ,
		\_2254__reg/NET0131 ,
		_w6849_
	);
	LUT2 #(
		.INIT('h1)
	) name5342 (
		_w6848_,
		_w6849_,
		_w6850_
	);
	LUT2 #(
		.INIT('h2)
	) name5343 (
		RESET_pad,
		_w6850_,
		_w6851_
	);
	LUT2 #(
		.INIT('h1)
	) name5344 (
		\WX9930_reg/NET0131 ,
		\_2310__reg/NET0131 ,
		_w6852_
	);
	LUT2 #(
		.INIT('h8)
	) name5345 (
		\WX9930_reg/NET0131 ,
		\_2310__reg/NET0131 ,
		_w6853_
	);
	LUT2 #(
		.INIT('h1)
	) name5346 (
		_w6852_,
		_w6853_,
		_w6854_
	);
	LUT2 #(
		.INIT('h2)
	) name5347 (
		RESET_pad,
		_w6854_,
		_w6855_
	);
	LUT2 #(
		.INIT('h1)
	) name5348 (
		\WX2148_reg/NET0131 ,
		\_2130__reg/NET0131 ,
		_w6856_
	);
	LUT2 #(
		.INIT('h8)
	) name5349 (
		\WX2148_reg/NET0131 ,
		\_2130__reg/NET0131 ,
		_w6857_
	);
	LUT2 #(
		.INIT('h1)
	) name5350 (
		_w6856_,
		_w6857_,
		_w6858_
	);
	LUT2 #(
		.INIT('h2)
	) name5351 (
		RESET_pad,
		_w6858_,
		_w6859_
	);
	LUT2 #(
		.INIT('h1)
	) name5352 (
		\WX7340_reg/NET0131 ,
		\_2248__reg/NET0131 ,
		_w6860_
	);
	LUT2 #(
		.INIT('h8)
	) name5353 (
		\WX7340_reg/NET0131 ,
		\_2248__reg/NET0131 ,
		_w6861_
	);
	LUT2 #(
		.INIT('h1)
	) name5354 (
		_w6860_,
		_w6861_,
		_w6862_
	);
	LUT2 #(
		.INIT('h2)
	) name5355 (
		RESET_pad,
		_w6862_,
		_w6863_
	);
	LUT2 #(
		.INIT('h1)
	) name5356 (
		\WX6061_reg/NET0131 ,
		\_2209__reg/NET0131 ,
		_w6864_
	);
	LUT2 #(
		.INIT('h8)
	) name5357 (
		\WX6061_reg/NET0131 ,
		\_2209__reg/NET0131 ,
		_w6865_
	);
	LUT2 #(
		.INIT('h1)
	) name5358 (
		_w6864_,
		_w6865_,
		_w6866_
	);
	LUT2 #(
		.INIT('h2)
	) name5359 (
		RESET_pad,
		_w6866_,
		_w6867_
	);
	LUT2 #(
		.INIT('h1)
	) name5360 (
		\WX8657_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w6868_
	);
	LUT2 #(
		.INIT('h8)
	) name5361 (
		\WX8657_reg/NET0131 ,
		\_2300__reg/NET0131 ,
		_w6869_
	);
	LUT2 #(
		.INIT('h1)
	) name5362 (
		_w6868_,
		_w6869_,
		_w6870_
	);
	LUT2 #(
		.INIT('h2)
	) name5363 (
		RESET_pad,
		_w6870_,
		_w6871_
	);
	LUT2 #(
		.INIT('h1)
	) name5364 (
		\WX2172_reg/NET0131 ,
		\_2118__reg/NET0131 ,
		_w6872_
	);
	LUT2 #(
		.INIT('h8)
	) name5365 (
		\WX2172_reg/NET0131 ,
		\_2118__reg/NET0131 ,
		_w6873_
	);
	LUT2 #(
		.INIT('h1)
	) name5366 (
		_w6872_,
		_w6873_,
		_w6874_
	);
	LUT2 #(
		.INIT('h2)
	) name5367 (
		RESET_pad,
		_w6874_,
		_w6875_
	);
	LUT2 #(
		.INIT('h1)
	) name5368 (
		\WX8607_reg/NET0131 ,
		\_2293__reg/NET0131 ,
		_w6876_
	);
	LUT2 #(
		.INIT('h8)
	) name5369 (
		\WX8607_reg/NET0131 ,
		\_2293__reg/NET0131 ,
		_w6877_
	);
	LUT2 #(
		.INIT('h1)
	) name5370 (
		_w6876_,
		_w6877_,
		_w6878_
	);
	LUT2 #(
		.INIT('h2)
	) name5371 (
		RESET_pad,
		_w6878_,
		_w6879_
	);
	LUT2 #(
		.INIT('h1)
	) name5372 (
		\WX899_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w6880_
	);
	LUT2 #(
		.INIT('h8)
	) name5373 (
		\WX899_reg/NET0131 ,
		\_2108__reg/NET0131 ,
		_w6881_
	);
	LUT2 #(
		.INIT('h1)
	) name5374 (
		_w6880_,
		_w6881_,
		_w6882_
	);
	LUT2 #(
		.INIT('h2)
	) name5375 (
		RESET_pad,
		_w6882_,
		_w6883_
	);
	LUT2 #(
		.INIT('h1)
	) name5376 (
		\WX897_reg/NET0131 ,
		\_2077__reg/NET0131 ,
		_w6884_
	);
	LUT2 #(
		.INIT('h8)
	) name5377 (
		\WX897_reg/NET0131 ,
		\_2077__reg/NET0131 ,
		_w6885_
	);
	LUT2 #(
		.INIT('h1)
	) name5378 (
		_w6884_,
		_w6885_,
		_w6886_
	);
	LUT2 #(
		.INIT('h2)
	) name5379 (
		RESET_pad,
		_w6886_,
		_w6887_
	);
	LUT2 #(
		.INIT('h1)
	) name5380 (
		\WX895_reg/NET0131 ,
		\_2078__reg/NET0131 ,
		_w6888_
	);
	LUT2 #(
		.INIT('h8)
	) name5381 (
		\WX895_reg/NET0131 ,
		\_2078__reg/NET0131 ,
		_w6889_
	);
	LUT2 #(
		.INIT('h1)
	) name5382 (
		_w6888_,
		_w6889_,
		_w6890_
	);
	LUT2 #(
		.INIT('h2)
	) name5383 (
		RESET_pad,
		_w6890_,
		_w6891_
	);
	LUT2 #(
		.INIT('h1)
	) name5384 (
		\WX893_reg/NET0131 ,
		\_2079__reg/NET0131 ,
		_w6892_
	);
	LUT2 #(
		.INIT('h8)
	) name5385 (
		\WX893_reg/NET0131 ,
		\_2079__reg/NET0131 ,
		_w6893_
	);
	LUT2 #(
		.INIT('h1)
	) name5386 (
		_w6892_,
		_w6893_,
		_w6894_
	);
	LUT2 #(
		.INIT('h2)
	) name5387 (
		RESET_pad,
		_w6894_,
		_w6895_
	);
	LUT2 #(
		.INIT('h1)
	) name5388 (
		\WX889_reg/NET0131 ,
		\_2081__reg/NET0131 ,
		_w6896_
	);
	LUT2 #(
		.INIT('h8)
	) name5389 (
		\WX889_reg/NET0131 ,
		\_2081__reg/NET0131 ,
		_w6897_
	);
	LUT2 #(
		.INIT('h1)
	) name5390 (
		_w6896_,
		_w6897_,
		_w6898_
	);
	LUT2 #(
		.INIT('h2)
	) name5391 (
		RESET_pad,
		_w6898_,
		_w6899_
	);
	LUT2 #(
		.INIT('h1)
	) name5392 (
		\WX887_reg/NET0131 ,
		\_2082__reg/NET0131 ,
		_w6900_
	);
	LUT2 #(
		.INIT('h8)
	) name5393 (
		\WX887_reg/NET0131 ,
		\_2082__reg/NET0131 ,
		_w6901_
	);
	LUT2 #(
		.INIT('h1)
	) name5394 (
		_w6900_,
		_w6901_,
		_w6902_
	);
	LUT2 #(
		.INIT('h2)
	) name5395 (
		RESET_pad,
		_w6902_,
		_w6903_
	);
	LUT2 #(
		.INIT('h1)
	) name5396 (
		\WX883_reg/NET0131 ,
		\_2084__reg/NET0131 ,
		_w6904_
	);
	LUT2 #(
		.INIT('h8)
	) name5397 (
		\WX883_reg/NET0131 ,
		\_2084__reg/NET0131 ,
		_w6905_
	);
	LUT2 #(
		.INIT('h1)
	) name5398 (
		_w6904_,
		_w6905_,
		_w6906_
	);
	LUT2 #(
		.INIT('h2)
	) name5399 (
		RESET_pad,
		_w6906_,
		_w6907_
	);
	LUT2 #(
		.INIT('h1)
	) name5400 (
		\WX881_reg/NET0131 ,
		\_2085__reg/NET0131 ,
		_w6908_
	);
	LUT2 #(
		.INIT('h8)
	) name5401 (
		\WX881_reg/NET0131 ,
		\_2085__reg/NET0131 ,
		_w6909_
	);
	LUT2 #(
		.INIT('h1)
	) name5402 (
		_w6908_,
		_w6909_,
		_w6910_
	);
	LUT2 #(
		.INIT('h2)
	) name5403 (
		RESET_pad,
		_w6910_,
		_w6911_
	);
	LUT2 #(
		.INIT('h1)
	) name5404 (
		\WX875_reg/NET0131 ,
		\_2088__reg/NET0131 ,
		_w6912_
	);
	LUT2 #(
		.INIT('h8)
	) name5405 (
		\WX875_reg/NET0131 ,
		\_2088__reg/NET0131 ,
		_w6913_
	);
	LUT2 #(
		.INIT('h1)
	) name5406 (
		_w6912_,
		_w6913_,
		_w6914_
	);
	LUT2 #(
		.INIT('h2)
	) name5407 (
		RESET_pad,
		_w6914_,
		_w6915_
	);
	LUT2 #(
		.INIT('h1)
	) name5408 (
		\WX873_reg/NET0131 ,
		\_2089__reg/NET0131 ,
		_w6916_
	);
	LUT2 #(
		.INIT('h8)
	) name5409 (
		\WX873_reg/NET0131 ,
		\_2089__reg/NET0131 ,
		_w6917_
	);
	LUT2 #(
		.INIT('h1)
	) name5410 (
		_w6916_,
		_w6917_,
		_w6918_
	);
	LUT2 #(
		.INIT('h2)
	) name5411 (
		RESET_pad,
		_w6918_,
		_w6919_
	);
	LUT2 #(
		.INIT('h1)
	) name5412 (
		\WX869_reg/NET0131 ,
		\_2091__reg/NET0131 ,
		_w6920_
	);
	LUT2 #(
		.INIT('h8)
	) name5413 (
		\WX869_reg/NET0131 ,
		\_2091__reg/NET0131 ,
		_w6921_
	);
	LUT2 #(
		.INIT('h1)
	) name5414 (
		_w6920_,
		_w6921_,
		_w6922_
	);
	LUT2 #(
		.INIT('h2)
	) name5415 (
		RESET_pad,
		_w6922_,
		_w6923_
	);
	LUT2 #(
		.INIT('h1)
	) name5416 (
		\WX865_reg/NET0131 ,
		\_2093__reg/NET0131 ,
		_w6924_
	);
	LUT2 #(
		.INIT('h8)
	) name5417 (
		\WX865_reg/NET0131 ,
		\_2093__reg/NET0131 ,
		_w6925_
	);
	LUT2 #(
		.INIT('h1)
	) name5418 (
		_w6924_,
		_w6925_,
		_w6926_
	);
	LUT2 #(
		.INIT('h2)
	) name5419 (
		RESET_pad,
		_w6926_,
		_w6927_
	);
	LUT2 #(
		.INIT('h1)
	) name5420 (
		\WX863_reg/NET0131 ,
		\_2094__reg/NET0131 ,
		_w6928_
	);
	LUT2 #(
		.INIT('h8)
	) name5421 (
		\WX863_reg/NET0131 ,
		\_2094__reg/NET0131 ,
		_w6929_
	);
	LUT2 #(
		.INIT('h1)
	) name5422 (
		_w6928_,
		_w6929_,
		_w6930_
	);
	LUT2 #(
		.INIT('h2)
	) name5423 (
		RESET_pad,
		_w6930_,
		_w6931_
	);
	LUT2 #(
		.INIT('h1)
	) name5424 (
		\WX855_reg/NET0131 ,
		\_2098__reg/NET0131 ,
		_w6932_
	);
	LUT2 #(
		.INIT('h8)
	) name5425 (
		\WX855_reg/NET0131 ,
		\_2098__reg/NET0131 ,
		_w6933_
	);
	LUT2 #(
		.INIT('h1)
	) name5426 (
		_w6932_,
		_w6933_,
		_w6934_
	);
	LUT2 #(
		.INIT('h2)
	) name5427 (
		RESET_pad,
		_w6934_,
		_w6935_
	);
	LUT2 #(
		.INIT('h1)
	) name5428 (
		\WX851_reg/NET0131 ,
		\_2100__reg/NET0131 ,
		_w6936_
	);
	LUT2 #(
		.INIT('h8)
	) name5429 (
		\WX851_reg/NET0131 ,
		\_2100__reg/NET0131 ,
		_w6937_
	);
	LUT2 #(
		.INIT('h1)
	) name5430 (
		_w6936_,
		_w6937_,
		_w6938_
	);
	LUT2 #(
		.INIT('h2)
	) name5431 (
		RESET_pad,
		_w6938_,
		_w6939_
	);
	LUT2 #(
		.INIT('h1)
	) name5432 (
		\WX845_reg/NET0131 ,
		\_2103__reg/NET0131 ,
		_w6940_
	);
	LUT2 #(
		.INIT('h8)
	) name5433 (
		\WX845_reg/NET0131 ,
		\_2103__reg/NET0131 ,
		_w6941_
	);
	LUT2 #(
		.INIT('h1)
	) name5434 (
		_w6940_,
		_w6941_,
		_w6942_
	);
	LUT2 #(
		.INIT('h2)
	) name5435 (
		RESET_pad,
		_w6942_,
		_w6943_
	);
	LUT2 #(
		.INIT('h1)
	) name5436 (
		\WX843_reg/NET0131 ,
		\_2104__reg/NET0131 ,
		_w6944_
	);
	LUT2 #(
		.INIT('h8)
	) name5437 (
		\WX843_reg/NET0131 ,
		\_2104__reg/NET0131 ,
		_w6945_
	);
	LUT2 #(
		.INIT('h1)
	) name5438 (
		_w6944_,
		_w6945_,
		_w6946_
	);
	LUT2 #(
		.INIT('h2)
	) name5439 (
		RESET_pad,
		_w6946_,
		_w6947_
	);
	LUT2 #(
		.INIT('h1)
	) name5440 (
		\WX841_reg/NET0131 ,
		\_2105__reg/NET0131 ,
		_w6948_
	);
	LUT2 #(
		.INIT('h8)
	) name5441 (
		\WX841_reg/NET0131 ,
		\_2105__reg/NET0131 ,
		_w6949_
	);
	LUT2 #(
		.INIT('h1)
	) name5442 (
		_w6948_,
		_w6949_,
		_w6950_
	);
	LUT2 #(
		.INIT('h2)
	) name5443 (
		RESET_pad,
		_w6950_,
		_w6951_
	);
	LUT2 #(
		.INIT('h1)
	) name5444 (
		\WX839_reg/NET0131 ,
		\_2106__reg/NET0131 ,
		_w6952_
	);
	LUT2 #(
		.INIT('h8)
	) name5445 (
		\WX839_reg/NET0131 ,
		\_2106__reg/NET0131 ,
		_w6953_
	);
	LUT2 #(
		.INIT('h1)
	) name5446 (
		_w6952_,
		_w6953_,
		_w6954_
	);
	LUT2 #(
		.INIT('h2)
	) name5447 (
		RESET_pad,
		_w6954_,
		_w6955_
	);
	LUT2 #(
		.INIT('h1)
	) name5448 (
		\WX2192_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w6956_
	);
	LUT2 #(
		.INIT('h8)
	) name5449 (
		\WX2192_reg/NET0131 ,
		\_2140__reg/NET0131 ,
		_w6957_
	);
	LUT2 #(
		.INIT('h1)
	) name5450 (
		_w6956_,
		_w6957_,
		_w6958_
	);
	LUT2 #(
		.INIT('h2)
	) name5451 (
		RESET_pad,
		_w6958_,
		_w6959_
	);
	LUT2 #(
		.INIT('h1)
	) name5452 (
		\WX2190_reg/NET0131 ,
		\_2109__reg/NET0131 ,
		_w6960_
	);
	LUT2 #(
		.INIT('h8)
	) name5453 (
		\WX2190_reg/NET0131 ,
		\_2109__reg/NET0131 ,
		_w6961_
	);
	LUT2 #(
		.INIT('h1)
	) name5454 (
		_w6960_,
		_w6961_,
		_w6962_
	);
	LUT2 #(
		.INIT('h2)
	) name5455 (
		RESET_pad,
		_w6962_,
		_w6963_
	);
	LUT2 #(
		.INIT('h1)
	) name5456 (
		\WX2188_reg/NET0131 ,
		\_2110__reg/NET0131 ,
		_w6964_
	);
	LUT2 #(
		.INIT('h8)
	) name5457 (
		\WX2188_reg/NET0131 ,
		\_2110__reg/NET0131 ,
		_w6965_
	);
	LUT2 #(
		.INIT('h1)
	) name5458 (
		_w6964_,
		_w6965_,
		_w6966_
	);
	LUT2 #(
		.INIT('h2)
	) name5459 (
		RESET_pad,
		_w6966_,
		_w6967_
	);
	LUT2 #(
		.INIT('h1)
	) name5460 (
		\WX2186_reg/NET0131 ,
		\_2111__reg/NET0131 ,
		_w6968_
	);
	LUT2 #(
		.INIT('h8)
	) name5461 (
		\WX2186_reg/NET0131 ,
		\_2111__reg/NET0131 ,
		_w6969_
	);
	LUT2 #(
		.INIT('h1)
	) name5462 (
		_w6968_,
		_w6969_,
		_w6970_
	);
	LUT2 #(
		.INIT('h2)
	) name5463 (
		RESET_pad,
		_w6970_,
		_w6971_
	);
	LUT2 #(
		.INIT('h1)
	) name5464 (
		\WX2182_reg/NET0131 ,
		\_2113__reg/NET0131 ,
		_w6972_
	);
	LUT2 #(
		.INIT('h8)
	) name5465 (
		\WX2182_reg/NET0131 ,
		\_2113__reg/NET0131 ,
		_w6973_
	);
	LUT2 #(
		.INIT('h1)
	) name5466 (
		_w6972_,
		_w6973_,
		_w6974_
	);
	LUT2 #(
		.INIT('h2)
	) name5467 (
		RESET_pad,
		_w6974_,
		_w6975_
	);
	LUT2 #(
		.INIT('h1)
	) name5468 (
		\WX2180_reg/NET0131 ,
		\_2114__reg/NET0131 ,
		_w6976_
	);
	LUT2 #(
		.INIT('h8)
	) name5469 (
		\WX2180_reg/NET0131 ,
		\_2114__reg/NET0131 ,
		_w6977_
	);
	LUT2 #(
		.INIT('h1)
	) name5470 (
		_w6976_,
		_w6977_,
		_w6978_
	);
	LUT2 #(
		.INIT('h2)
	) name5471 (
		RESET_pad,
		_w6978_,
		_w6979_
	);
	LUT2 #(
		.INIT('h1)
	) name5472 (
		\WX2174_reg/NET0131 ,
		\_2117__reg/NET0131 ,
		_w6980_
	);
	LUT2 #(
		.INIT('h8)
	) name5473 (
		\WX2174_reg/NET0131 ,
		\_2117__reg/NET0131 ,
		_w6981_
	);
	LUT2 #(
		.INIT('h1)
	) name5474 (
		_w6980_,
		_w6981_,
		_w6982_
	);
	LUT2 #(
		.INIT('h2)
	) name5475 (
		RESET_pad,
		_w6982_,
		_w6983_
	);
	LUT2 #(
		.INIT('h1)
	) name5476 (
		\WX2168_reg/NET0131 ,
		\_2120__reg/NET0131 ,
		_w6984_
	);
	LUT2 #(
		.INIT('h8)
	) name5477 (
		\WX2168_reg/NET0131 ,
		\_2120__reg/NET0131 ,
		_w6985_
	);
	LUT2 #(
		.INIT('h1)
	) name5478 (
		_w6984_,
		_w6985_,
		_w6986_
	);
	LUT2 #(
		.INIT('h2)
	) name5479 (
		RESET_pad,
		_w6986_,
		_w6987_
	);
	LUT2 #(
		.INIT('h1)
	) name5480 (
		\WX2166_reg/NET0131 ,
		\_2121__reg/NET0131 ,
		_w6988_
	);
	LUT2 #(
		.INIT('h8)
	) name5481 (
		\WX2166_reg/NET0131 ,
		\_2121__reg/NET0131 ,
		_w6989_
	);
	LUT2 #(
		.INIT('h1)
	) name5482 (
		_w6988_,
		_w6989_,
		_w6990_
	);
	LUT2 #(
		.INIT('h2)
	) name5483 (
		RESET_pad,
		_w6990_,
		_w6991_
	);
	LUT2 #(
		.INIT('h1)
	) name5484 (
		\WX2164_reg/NET0131 ,
		\_2122__reg/NET0131 ,
		_w6992_
	);
	LUT2 #(
		.INIT('h8)
	) name5485 (
		\WX2164_reg/NET0131 ,
		\_2122__reg/NET0131 ,
		_w6993_
	);
	LUT2 #(
		.INIT('h1)
	) name5486 (
		_w6992_,
		_w6993_,
		_w6994_
	);
	LUT2 #(
		.INIT('h2)
	) name5487 (
		RESET_pad,
		_w6994_,
		_w6995_
	);
	LUT2 #(
		.INIT('h1)
	) name5488 (
		\WX2162_reg/NET0131 ,
		\_2123__reg/NET0131 ,
		_w6996_
	);
	LUT2 #(
		.INIT('h8)
	) name5489 (
		\WX2162_reg/NET0131 ,
		\_2123__reg/NET0131 ,
		_w6997_
	);
	LUT2 #(
		.INIT('h1)
	) name5490 (
		_w6996_,
		_w6997_,
		_w6998_
	);
	LUT2 #(
		.INIT('h2)
	) name5491 (
		RESET_pad,
		_w6998_,
		_w6999_
	);
	LUT2 #(
		.INIT('h1)
	) name5492 (
		\WX2158_reg/NET0131 ,
		\_2125__reg/NET0131 ,
		_w7000_
	);
	LUT2 #(
		.INIT('h8)
	) name5493 (
		\WX2158_reg/NET0131 ,
		\_2125__reg/NET0131 ,
		_w7001_
	);
	LUT2 #(
		.INIT('h1)
	) name5494 (
		_w7000_,
		_w7001_,
		_w7002_
	);
	LUT2 #(
		.INIT('h2)
	) name5495 (
		RESET_pad,
		_w7002_,
		_w7003_
	);
	LUT2 #(
		.INIT('h1)
	) name5496 (
		\WX2156_reg/NET0131 ,
		\_2126__reg/NET0131 ,
		_w7004_
	);
	LUT2 #(
		.INIT('h8)
	) name5497 (
		\WX2156_reg/NET0131 ,
		\_2126__reg/NET0131 ,
		_w7005_
	);
	LUT2 #(
		.INIT('h1)
	) name5498 (
		_w7004_,
		_w7005_,
		_w7006_
	);
	LUT2 #(
		.INIT('h2)
	) name5499 (
		RESET_pad,
		_w7006_,
		_w7007_
	);
	LUT2 #(
		.INIT('h1)
	) name5500 (
		\WX2154_reg/NET0131 ,
		\_2127__reg/NET0131 ,
		_w7008_
	);
	LUT2 #(
		.INIT('h8)
	) name5501 (
		\WX2154_reg/NET0131 ,
		\_2127__reg/NET0131 ,
		_w7009_
	);
	LUT2 #(
		.INIT('h1)
	) name5502 (
		_w7008_,
		_w7009_,
		_w7010_
	);
	LUT2 #(
		.INIT('h2)
	) name5503 (
		RESET_pad,
		_w7010_,
		_w7011_
	);
	LUT2 #(
		.INIT('h1)
	) name5504 (
		\WX2146_reg/NET0131 ,
		\_2131__reg/NET0131 ,
		_w7012_
	);
	LUT2 #(
		.INIT('h8)
	) name5505 (
		\WX2146_reg/NET0131 ,
		\_2131__reg/NET0131 ,
		_w7013_
	);
	LUT2 #(
		.INIT('h1)
	) name5506 (
		_w7012_,
		_w7013_,
		_w7014_
	);
	LUT2 #(
		.INIT('h2)
	) name5507 (
		RESET_pad,
		_w7014_,
		_w7015_
	);
	LUT2 #(
		.INIT('h1)
	) name5508 (
		\WX2144_reg/NET0131 ,
		\_2132__reg/NET0131 ,
		_w7016_
	);
	LUT2 #(
		.INIT('h8)
	) name5509 (
		\WX2144_reg/NET0131 ,
		\_2132__reg/NET0131 ,
		_w7017_
	);
	LUT2 #(
		.INIT('h1)
	) name5510 (
		_w7016_,
		_w7017_,
		_w7018_
	);
	LUT2 #(
		.INIT('h2)
	) name5511 (
		RESET_pad,
		_w7018_,
		_w7019_
	);
	LUT2 #(
		.INIT('h1)
	) name5512 (
		\WX2142_reg/NET0131 ,
		\_2133__reg/NET0131 ,
		_w7020_
	);
	LUT2 #(
		.INIT('h8)
	) name5513 (
		\WX2142_reg/NET0131 ,
		\_2133__reg/NET0131 ,
		_w7021_
	);
	LUT2 #(
		.INIT('h1)
	) name5514 (
		_w7020_,
		_w7021_,
		_w7022_
	);
	LUT2 #(
		.INIT('h2)
	) name5515 (
		RESET_pad,
		_w7022_,
		_w7023_
	);
	LUT2 #(
		.INIT('h1)
	) name5516 (
		\WX2138_reg/NET0131 ,
		\_2135__reg/NET0131 ,
		_w7024_
	);
	LUT2 #(
		.INIT('h8)
	) name5517 (
		\WX2138_reg/NET0131 ,
		\_2135__reg/NET0131 ,
		_w7025_
	);
	LUT2 #(
		.INIT('h1)
	) name5518 (
		_w7024_,
		_w7025_,
		_w7026_
	);
	LUT2 #(
		.INIT('h2)
	) name5519 (
		RESET_pad,
		_w7026_,
		_w7027_
	);
	LUT2 #(
		.INIT('h1)
	) name5520 (
		\WX2134_reg/NET0131 ,
		\_2137__reg/NET0131 ,
		_w7028_
	);
	LUT2 #(
		.INIT('h8)
	) name5521 (
		\WX2134_reg/NET0131 ,
		\_2137__reg/NET0131 ,
		_w7029_
	);
	LUT2 #(
		.INIT('h1)
	) name5522 (
		_w7028_,
		_w7029_,
		_w7030_
	);
	LUT2 #(
		.INIT('h2)
	) name5523 (
		RESET_pad,
		_w7030_,
		_w7031_
	);
	LUT2 #(
		.INIT('h1)
	) name5524 (
		\WX7348_reg/NET0131 ,
		\_2244__reg/NET0131 ,
		_w7032_
	);
	LUT2 #(
		.INIT('h8)
	) name5525 (
		\WX7348_reg/NET0131 ,
		\_2244__reg/NET0131 ,
		_w7033_
	);
	LUT2 #(
		.INIT('h1)
	) name5526 (
		_w7032_,
		_w7033_,
		_w7034_
	);
	LUT2 #(
		.INIT('h2)
	) name5527 (
		RESET_pad,
		_w7034_,
		_w7035_
	);
	LUT2 #(
		.INIT('h1)
	) name5528 (
		\WX3483_reg/NET0131 ,
		\_2141__reg/NET0131 ,
		_w7036_
	);
	LUT2 #(
		.INIT('h8)
	) name5529 (
		\WX3483_reg/NET0131 ,
		\_2141__reg/NET0131 ,
		_w7037_
	);
	LUT2 #(
		.INIT('h1)
	) name5530 (
		_w7036_,
		_w7037_,
		_w7038_
	);
	LUT2 #(
		.INIT('h2)
	) name5531 (
		RESET_pad,
		_w7038_,
		_w7039_
	);
	LUT2 #(
		.INIT('h1)
	) name5532 (
		\WX3481_reg/NET0131 ,
		\_2142__reg/NET0131 ,
		_w7040_
	);
	LUT2 #(
		.INIT('h8)
	) name5533 (
		\WX3481_reg/NET0131 ,
		\_2142__reg/NET0131 ,
		_w7041_
	);
	LUT2 #(
		.INIT('h1)
	) name5534 (
		_w7040_,
		_w7041_,
		_w7042_
	);
	LUT2 #(
		.INIT('h2)
	) name5535 (
		RESET_pad,
		_w7042_,
		_w7043_
	);
	LUT2 #(
		.INIT('h1)
	) name5536 (
		\WX3479_reg/NET0131 ,
		\_2143__reg/NET0131 ,
		_w7044_
	);
	LUT2 #(
		.INIT('h8)
	) name5537 (
		\WX3479_reg/NET0131 ,
		\_2143__reg/NET0131 ,
		_w7045_
	);
	LUT2 #(
		.INIT('h1)
	) name5538 (
		_w7044_,
		_w7045_,
		_w7046_
	);
	LUT2 #(
		.INIT('h2)
	) name5539 (
		RESET_pad,
		_w7046_,
		_w7047_
	);
	LUT2 #(
		.INIT('h1)
	) name5540 (
		\WX3473_reg/NET0131 ,
		\_2146__reg/NET0131 ,
		_w7048_
	);
	LUT2 #(
		.INIT('h8)
	) name5541 (
		\WX3473_reg/NET0131 ,
		\_2146__reg/NET0131 ,
		_w7049_
	);
	LUT2 #(
		.INIT('h1)
	) name5542 (
		_w7048_,
		_w7049_,
		_w7050_
	);
	LUT2 #(
		.INIT('h2)
	) name5543 (
		RESET_pad,
		_w7050_,
		_w7051_
	);
	LUT2 #(
		.INIT('h1)
	) name5544 (
		\WX3471_reg/NET0131 ,
		\_2147__reg/NET0131 ,
		_w7052_
	);
	LUT2 #(
		.INIT('h8)
	) name5545 (
		\WX3471_reg/NET0131 ,
		\_2147__reg/NET0131 ,
		_w7053_
	);
	LUT2 #(
		.INIT('h1)
	) name5546 (
		_w7052_,
		_w7053_,
		_w7054_
	);
	LUT2 #(
		.INIT('h2)
	) name5547 (
		RESET_pad,
		_w7054_,
		_w7055_
	);
	LUT2 #(
		.INIT('h1)
	) name5548 (
		\WX3469_reg/NET0131 ,
		\_2148__reg/NET0131 ,
		_w7056_
	);
	LUT2 #(
		.INIT('h8)
	) name5549 (
		\WX3469_reg/NET0131 ,
		\_2148__reg/NET0131 ,
		_w7057_
	);
	LUT2 #(
		.INIT('h1)
	) name5550 (
		_w7056_,
		_w7057_,
		_w7058_
	);
	LUT2 #(
		.INIT('h2)
	) name5551 (
		RESET_pad,
		_w7058_,
		_w7059_
	);
	LUT2 #(
		.INIT('h1)
	) name5552 (
		\WX3465_reg/NET0131 ,
		\_2150__reg/NET0131 ,
		_w7060_
	);
	LUT2 #(
		.INIT('h8)
	) name5553 (
		\WX3465_reg/NET0131 ,
		\_2150__reg/NET0131 ,
		_w7061_
	);
	LUT2 #(
		.INIT('h1)
	) name5554 (
		_w7060_,
		_w7061_,
		_w7062_
	);
	LUT2 #(
		.INIT('h2)
	) name5555 (
		RESET_pad,
		_w7062_,
		_w7063_
	);
	LUT2 #(
		.INIT('h1)
	) name5556 (
		\WX3459_reg/NET0131 ,
		\_2153__reg/NET0131 ,
		_w7064_
	);
	LUT2 #(
		.INIT('h8)
	) name5557 (
		\WX3459_reg/NET0131 ,
		\_2153__reg/NET0131 ,
		_w7065_
	);
	LUT2 #(
		.INIT('h1)
	) name5558 (
		_w7064_,
		_w7065_,
		_w7066_
	);
	LUT2 #(
		.INIT('h2)
	) name5559 (
		RESET_pad,
		_w7066_,
		_w7067_
	);
	LUT2 #(
		.INIT('h1)
	) name5560 (
		\WX3457_reg/NET0131 ,
		\_2154__reg/NET0131 ,
		_w7068_
	);
	LUT2 #(
		.INIT('h8)
	) name5561 (
		\WX3457_reg/NET0131 ,
		\_2154__reg/NET0131 ,
		_w7069_
	);
	LUT2 #(
		.INIT('h1)
	) name5562 (
		_w7068_,
		_w7069_,
		_w7070_
	);
	LUT2 #(
		.INIT('h2)
	) name5563 (
		RESET_pad,
		_w7070_,
		_w7071_
	);
	LUT2 #(
		.INIT('h1)
	) name5564 (
		\WX3455_reg/NET0131 ,
		\_2155__reg/NET0131 ,
		_w7072_
	);
	LUT2 #(
		.INIT('h8)
	) name5565 (
		\WX3455_reg/NET0131 ,
		\_2155__reg/NET0131 ,
		_w7073_
	);
	LUT2 #(
		.INIT('h1)
	) name5566 (
		_w7072_,
		_w7073_,
		_w7074_
	);
	LUT2 #(
		.INIT('h2)
	) name5567 (
		RESET_pad,
		_w7074_,
		_w7075_
	);
	LUT2 #(
		.INIT('h1)
	) name5568 (
		\WX3451_reg/NET0131 ,
		\_2157__reg/NET0131 ,
		_w7076_
	);
	LUT2 #(
		.INIT('h8)
	) name5569 (
		\WX3451_reg/NET0131 ,
		\_2157__reg/NET0131 ,
		_w7077_
	);
	LUT2 #(
		.INIT('h1)
	) name5570 (
		_w7076_,
		_w7077_,
		_w7078_
	);
	LUT2 #(
		.INIT('h2)
	) name5571 (
		RESET_pad,
		_w7078_,
		_w7079_
	);
	LUT2 #(
		.INIT('h1)
	) name5572 (
		\WX3449_reg/NET0131 ,
		\_2158__reg/NET0131 ,
		_w7080_
	);
	LUT2 #(
		.INIT('h8)
	) name5573 (
		\WX3449_reg/NET0131 ,
		\_2158__reg/NET0131 ,
		_w7081_
	);
	LUT2 #(
		.INIT('h1)
	) name5574 (
		_w7080_,
		_w7081_,
		_w7082_
	);
	LUT2 #(
		.INIT('h2)
	) name5575 (
		RESET_pad,
		_w7082_,
		_w7083_
	);
	LUT2 #(
		.INIT('h1)
	) name5576 (
		\WX3445_reg/NET0131 ,
		\_2160__reg/NET0131 ,
		_w7084_
	);
	LUT2 #(
		.INIT('h8)
	) name5577 (
		\WX3445_reg/NET0131 ,
		\_2160__reg/NET0131 ,
		_w7085_
	);
	LUT2 #(
		.INIT('h1)
	) name5578 (
		_w7084_,
		_w7085_,
		_w7086_
	);
	LUT2 #(
		.INIT('h2)
	) name5579 (
		RESET_pad,
		_w7086_,
		_w7087_
	);
	LUT2 #(
		.INIT('h1)
	) name5580 (
		\WX3443_reg/NET0131 ,
		\_2161__reg/NET0131 ,
		_w7088_
	);
	LUT2 #(
		.INIT('h8)
	) name5581 (
		\WX3443_reg/NET0131 ,
		\_2161__reg/NET0131 ,
		_w7089_
	);
	LUT2 #(
		.INIT('h1)
	) name5582 (
		_w7088_,
		_w7089_,
		_w7090_
	);
	LUT2 #(
		.INIT('h2)
	) name5583 (
		RESET_pad,
		_w7090_,
		_w7091_
	);
	LUT2 #(
		.INIT('h1)
	) name5584 (
		\WX3441_reg/NET0131 ,
		\_2162__reg/NET0131 ,
		_w7092_
	);
	LUT2 #(
		.INIT('h8)
	) name5585 (
		\WX3441_reg/NET0131 ,
		\_2162__reg/NET0131 ,
		_w7093_
	);
	LUT2 #(
		.INIT('h1)
	) name5586 (
		_w7092_,
		_w7093_,
		_w7094_
	);
	LUT2 #(
		.INIT('h2)
	) name5587 (
		RESET_pad,
		_w7094_,
		_w7095_
	);
	LUT2 #(
		.INIT('h1)
	) name5588 (
		\WX3439_reg/NET0131 ,
		\_2163__reg/NET0131 ,
		_w7096_
	);
	LUT2 #(
		.INIT('h8)
	) name5589 (
		\WX3439_reg/NET0131 ,
		\_2163__reg/NET0131 ,
		_w7097_
	);
	LUT2 #(
		.INIT('h1)
	) name5590 (
		_w7096_,
		_w7097_,
		_w7098_
	);
	LUT2 #(
		.INIT('h2)
	) name5591 (
		RESET_pad,
		_w7098_,
		_w7099_
	);
	LUT2 #(
		.INIT('h1)
	) name5592 (
		\WX3437_reg/NET0131 ,
		\_2164__reg/NET0131 ,
		_w7100_
	);
	LUT2 #(
		.INIT('h8)
	) name5593 (
		\WX3437_reg/NET0131 ,
		\_2164__reg/NET0131 ,
		_w7101_
	);
	LUT2 #(
		.INIT('h1)
	) name5594 (
		_w7100_,
		_w7101_,
		_w7102_
	);
	LUT2 #(
		.INIT('h2)
	) name5595 (
		RESET_pad,
		_w7102_,
		_w7103_
	);
	LUT2 #(
		.INIT('h1)
	) name5596 (
		\WX3435_reg/NET0131 ,
		\_2165__reg/NET0131 ,
		_w7104_
	);
	LUT2 #(
		.INIT('h8)
	) name5597 (
		\WX3435_reg/NET0131 ,
		\_2165__reg/NET0131 ,
		_w7105_
	);
	LUT2 #(
		.INIT('h1)
	) name5598 (
		_w7104_,
		_w7105_,
		_w7106_
	);
	LUT2 #(
		.INIT('h2)
	) name5599 (
		RESET_pad,
		_w7106_,
		_w7107_
	);
	LUT2 #(
		.INIT('h1)
	) name5600 (
		\WX3433_reg/NET0131 ,
		\_2166__reg/NET0131 ,
		_w7108_
	);
	LUT2 #(
		.INIT('h8)
	) name5601 (
		\WX3433_reg/NET0131 ,
		\_2166__reg/NET0131 ,
		_w7109_
	);
	LUT2 #(
		.INIT('h1)
	) name5602 (
		_w7108_,
		_w7109_,
		_w7110_
	);
	LUT2 #(
		.INIT('h2)
	) name5603 (
		RESET_pad,
		_w7110_,
		_w7111_
	);
	LUT2 #(
		.INIT('h1)
	) name5604 (
		\WX3431_reg/NET0131 ,
		\_2167__reg/NET0131 ,
		_w7112_
	);
	LUT2 #(
		.INIT('h8)
	) name5605 (
		\WX3431_reg/NET0131 ,
		\_2167__reg/NET0131 ,
		_w7113_
	);
	LUT2 #(
		.INIT('h1)
	) name5606 (
		_w7112_,
		_w7113_,
		_w7114_
	);
	LUT2 #(
		.INIT('h2)
	) name5607 (
		RESET_pad,
		_w7114_,
		_w7115_
	);
	LUT2 #(
		.INIT('h1)
	) name5608 (
		\WX3429_reg/NET0131 ,
		\_2168__reg/NET0131 ,
		_w7116_
	);
	LUT2 #(
		.INIT('h8)
	) name5609 (
		\WX3429_reg/NET0131 ,
		\_2168__reg/NET0131 ,
		_w7117_
	);
	LUT2 #(
		.INIT('h1)
	) name5610 (
		_w7116_,
		_w7117_,
		_w7118_
	);
	LUT2 #(
		.INIT('h2)
	) name5611 (
		RESET_pad,
		_w7118_,
		_w7119_
	);
	LUT2 #(
		.INIT('h1)
	) name5612 (
		\WX3423_reg/NET0131 ,
		\_2171__reg/NET0131 ,
		_w7120_
	);
	LUT2 #(
		.INIT('h8)
	) name5613 (
		\WX3423_reg/NET0131 ,
		\_2171__reg/NET0131 ,
		_w7121_
	);
	LUT2 #(
		.INIT('h1)
	) name5614 (
		_w7120_,
		_w7121_,
		_w7122_
	);
	LUT2 #(
		.INIT('h2)
	) name5615 (
		RESET_pad,
		_w7122_,
		_w7123_
	);
	LUT2 #(
		.INIT('h1)
	) name5616 (
		\WX4778_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w7124_
	);
	LUT2 #(
		.INIT('h8)
	) name5617 (
		\WX4778_reg/NET0131 ,
		\_2204__reg/NET0131 ,
		_w7125_
	);
	LUT2 #(
		.INIT('h1)
	) name5618 (
		_w7124_,
		_w7125_,
		_w7126_
	);
	LUT2 #(
		.INIT('h2)
	) name5619 (
		RESET_pad,
		_w7126_,
		_w7127_
	);
	LUT2 #(
		.INIT('h1)
	) name5620 (
		\WX4776_reg/NET0131 ,
		\_2173__reg/NET0131 ,
		_w7128_
	);
	LUT2 #(
		.INIT('h8)
	) name5621 (
		\WX4776_reg/NET0131 ,
		\_2173__reg/NET0131 ,
		_w7129_
	);
	LUT2 #(
		.INIT('h1)
	) name5622 (
		_w7128_,
		_w7129_,
		_w7130_
	);
	LUT2 #(
		.INIT('h2)
	) name5623 (
		RESET_pad,
		_w7130_,
		_w7131_
	);
	LUT2 #(
		.INIT('h1)
	) name5624 (
		\WX4774_reg/NET0131 ,
		\_2174__reg/NET0131 ,
		_w7132_
	);
	LUT2 #(
		.INIT('h8)
	) name5625 (
		\WX4774_reg/NET0131 ,
		\_2174__reg/NET0131 ,
		_w7133_
	);
	LUT2 #(
		.INIT('h1)
	) name5626 (
		_w7132_,
		_w7133_,
		_w7134_
	);
	LUT2 #(
		.INIT('h2)
	) name5627 (
		RESET_pad,
		_w7134_,
		_w7135_
	);
	LUT2 #(
		.INIT('h1)
	) name5628 (
		\WX4772_reg/NET0131 ,
		\_2175__reg/NET0131 ,
		_w7136_
	);
	LUT2 #(
		.INIT('h8)
	) name5629 (
		\WX4772_reg/NET0131 ,
		\_2175__reg/NET0131 ,
		_w7137_
	);
	LUT2 #(
		.INIT('h1)
	) name5630 (
		_w7136_,
		_w7137_,
		_w7138_
	);
	LUT2 #(
		.INIT('h2)
	) name5631 (
		RESET_pad,
		_w7138_,
		_w7139_
	);
	LUT2 #(
		.INIT('h1)
	) name5632 (
		\WX7316_reg/NET0131 ,
		\_2260__reg/NET0131 ,
		_w7140_
	);
	LUT2 #(
		.INIT('h8)
	) name5633 (
		\WX7316_reg/NET0131 ,
		\_2260__reg/NET0131 ,
		_w7141_
	);
	LUT2 #(
		.INIT('h1)
	) name5634 (
		_w7140_,
		_w7141_,
		_w7142_
	);
	LUT2 #(
		.INIT('h2)
	) name5635 (
		RESET_pad,
		_w7142_,
		_w7143_
	);
	LUT2 #(
		.INIT('h1)
	) name5636 (
		\WX4768_reg/NET0131 ,
		\_2177__reg/NET0131 ,
		_w7144_
	);
	LUT2 #(
		.INIT('h8)
	) name5637 (
		\WX4768_reg/NET0131 ,
		\_2177__reg/NET0131 ,
		_w7145_
	);
	LUT2 #(
		.INIT('h1)
	) name5638 (
		_w7144_,
		_w7145_,
		_w7146_
	);
	LUT2 #(
		.INIT('h2)
	) name5639 (
		RESET_pad,
		_w7146_,
		_w7147_
	);
	LUT2 #(
		.INIT('h1)
	) name5640 (
		\WX4766_reg/NET0131 ,
		\_2178__reg/NET0131 ,
		_w7148_
	);
	LUT2 #(
		.INIT('h8)
	) name5641 (
		\WX4766_reg/NET0131 ,
		\_2178__reg/NET0131 ,
		_w7149_
	);
	LUT2 #(
		.INIT('h1)
	) name5642 (
		_w7148_,
		_w7149_,
		_w7150_
	);
	LUT2 #(
		.INIT('h2)
	) name5643 (
		RESET_pad,
		_w7150_,
		_w7151_
	);
	LUT2 #(
		.INIT('h1)
	) name5644 (
		\WX4764_reg/NET0131 ,
		\_2179__reg/NET0131 ,
		_w7152_
	);
	LUT2 #(
		.INIT('h8)
	) name5645 (
		\WX4764_reg/NET0131 ,
		\_2179__reg/NET0131 ,
		_w7153_
	);
	LUT2 #(
		.INIT('h1)
	) name5646 (
		_w7152_,
		_w7153_,
		_w7154_
	);
	LUT2 #(
		.INIT('h2)
	) name5647 (
		RESET_pad,
		_w7154_,
		_w7155_
	);
	LUT2 #(
		.INIT('h1)
	) name5648 (
		\WX4760_reg/NET0131 ,
		\_2181__reg/NET0131 ,
		_w7156_
	);
	LUT2 #(
		.INIT('h8)
	) name5649 (
		\WX4760_reg/NET0131 ,
		\_2181__reg/NET0131 ,
		_w7157_
	);
	LUT2 #(
		.INIT('h1)
	) name5650 (
		_w7156_,
		_w7157_,
		_w7158_
	);
	LUT2 #(
		.INIT('h2)
	) name5651 (
		RESET_pad,
		_w7158_,
		_w7159_
	);
	LUT2 #(
		.INIT('h1)
	) name5652 (
		\WX4758_reg/NET0131 ,
		\_2182__reg/NET0131 ,
		_w7160_
	);
	LUT2 #(
		.INIT('h8)
	) name5653 (
		\WX4758_reg/NET0131 ,
		\_2182__reg/NET0131 ,
		_w7161_
	);
	LUT2 #(
		.INIT('h1)
	) name5654 (
		_w7160_,
		_w7161_,
		_w7162_
	);
	LUT2 #(
		.INIT('h2)
	) name5655 (
		RESET_pad,
		_w7162_,
		_w7163_
	);
	LUT2 #(
		.INIT('h1)
	) name5656 (
		\WX4754_reg/NET0131 ,
		\_2184__reg/NET0131 ,
		_w7164_
	);
	LUT2 #(
		.INIT('h8)
	) name5657 (
		\WX4754_reg/NET0131 ,
		\_2184__reg/NET0131 ,
		_w7165_
	);
	LUT2 #(
		.INIT('h1)
	) name5658 (
		_w7164_,
		_w7165_,
		_w7166_
	);
	LUT2 #(
		.INIT('h2)
	) name5659 (
		RESET_pad,
		_w7166_,
		_w7167_
	);
	LUT2 #(
		.INIT('h1)
	) name5660 (
		\WX4752_reg/NET0131 ,
		\_2185__reg/NET0131 ,
		_w7168_
	);
	LUT2 #(
		.INIT('h8)
	) name5661 (
		\WX4752_reg/NET0131 ,
		\_2185__reg/NET0131 ,
		_w7169_
	);
	LUT2 #(
		.INIT('h1)
	) name5662 (
		_w7168_,
		_w7169_,
		_w7170_
	);
	LUT2 #(
		.INIT('h2)
	) name5663 (
		RESET_pad,
		_w7170_,
		_w7171_
	);
	LUT2 #(
		.INIT('h1)
	) name5664 (
		\WX4750_reg/NET0131 ,
		\_2186__reg/NET0131 ,
		_w7172_
	);
	LUT2 #(
		.INIT('h8)
	) name5665 (
		\WX4750_reg/NET0131 ,
		\_2186__reg/NET0131 ,
		_w7173_
	);
	LUT2 #(
		.INIT('h1)
	) name5666 (
		_w7172_,
		_w7173_,
		_w7174_
	);
	LUT2 #(
		.INIT('h2)
	) name5667 (
		RESET_pad,
		_w7174_,
		_w7175_
	);
	LUT2 #(
		.INIT('h1)
	) name5668 (
		\WX4748_reg/NET0131 ,
		\_2187__reg/NET0131 ,
		_w7176_
	);
	LUT2 #(
		.INIT('h8)
	) name5669 (
		\WX4748_reg/NET0131 ,
		\_2187__reg/NET0131 ,
		_w7177_
	);
	LUT2 #(
		.INIT('h1)
	) name5670 (
		_w7176_,
		_w7177_,
		_w7178_
	);
	LUT2 #(
		.INIT('h2)
	) name5671 (
		RESET_pad,
		_w7178_,
		_w7179_
	);
	LUT2 #(
		.INIT('h1)
	) name5672 (
		\WX4744_reg/NET0131 ,
		\_2189__reg/NET0131 ,
		_w7180_
	);
	LUT2 #(
		.INIT('h8)
	) name5673 (
		\WX4744_reg/NET0131 ,
		\_2189__reg/NET0131 ,
		_w7181_
	);
	LUT2 #(
		.INIT('h1)
	) name5674 (
		_w7180_,
		_w7181_,
		_w7182_
	);
	LUT2 #(
		.INIT('h2)
	) name5675 (
		RESET_pad,
		_w7182_,
		_w7183_
	);
	LUT2 #(
		.INIT('h1)
	) name5676 (
		\WX4742_reg/NET0131 ,
		\_2190__reg/NET0131 ,
		_w7184_
	);
	LUT2 #(
		.INIT('h8)
	) name5677 (
		\WX4742_reg/NET0131 ,
		\_2190__reg/NET0131 ,
		_w7185_
	);
	LUT2 #(
		.INIT('h1)
	) name5678 (
		_w7184_,
		_w7185_,
		_w7186_
	);
	LUT2 #(
		.INIT('h2)
	) name5679 (
		RESET_pad,
		_w7186_,
		_w7187_
	);
	LUT2 #(
		.INIT('h1)
	) name5680 (
		\WX4740_reg/NET0131 ,
		\_2191__reg/NET0131 ,
		_w7188_
	);
	LUT2 #(
		.INIT('h8)
	) name5681 (
		\WX4740_reg/NET0131 ,
		\_2191__reg/NET0131 ,
		_w7189_
	);
	LUT2 #(
		.INIT('h1)
	) name5682 (
		_w7188_,
		_w7189_,
		_w7190_
	);
	LUT2 #(
		.INIT('h2)
	) name5683 (
		RESET_pad,
		_w7190_,
		_w7191_
	);
	LUT2 #(
		.INIT('h1)
	) name5684 (
		\WX4738_reg/NET0131 ,
		\_2192__reg/NET0131 ,
		_w7192_
	);
	LUT2 #(
		.INIT('h8)
	) name5685 (
		\WX4738_reg/NET0131 ,
		\_2192__reg/NET0131 ,
		_w7193_
	);
	LUT2 #(
		.INIT('h1)
	) name5686 (
		_w7192_,
		_w7193_,
		_w7194_
	);
	LUT2 #(
		.INIT('h2)
	) name5687 (
		RESET_pad,
		_w7194_,
		_w7195_
	);
	LUT2 #(
		.INIT('h1)
	) name5688 (
		\WX4736_reg/NET0131 ,
		\_2193__reg/NET0131 ,
		_w7196_
	);
	LUT2 #(
		.INIT('h8)
	) name5689 (
		\WX4736_reg/NET0131 ,
		\_2193__reg/NET0131 ,
		_w7197_
	);
	LUT2 #(
		.INIT('h1)
	) name5690 (
		_w7196_,
		_w7197_,
		_w7198_
	);
	LUT2 #(
		.INIT('h2)
	) name5691 (
		RESET_pad,
		_w7198_,
		_w7199_
	);
	LUT2 #(
		.INIT('h1)
	) name5692 (
		\WX4734_reg/NET0131 ,
		\_2194__reg/NET0131 ,
		_w7200_
	);
	LUT2 #(
		.INIT('h8)
	) name5693 (
		\WX4734_reg/NET0131 ,
		\_2194__reg/NET0131 ,
		_w7201_
	);
	LUT2 #(
		.INIT('h1)
	) name5694 (
		_w7200_,
		_w7201_,
		_w7202_
	);
	LUT2 #(
		.INIT('h2)
	) name5695 (
		RESET_pad,
		_w7202_,
		_w7203_
	);
	LUT2 #(
		.INIT('h1)
	) name5696 (
		\WX4732_reg/NET0131 ,
		\_2195__reg/NET0131 ,
		_w7204_
	);
	LUT2 #(
		.INIT('h8)
	) name5697 (
		\WX4732_reg/NET0131 ,
		\_2195__reg/NET0131 ,
		_w7205_
	);
	LUT2 #(
		.INIT('h1)
	) name5698 (
		_w7204_,
		_w7205_,
		_w7206_
	);
	LUT2 #(
		.INIT('h2)
	) name5699 (
		RESET_pad,
		_w7206_,
		_w7207_
	);
	LUT2 #(
		.INIT('h1)
	) name5700 (
		\WX4730_reg/NET0131 ,
		\_2196__reg/NET0131 ,
		_w7208_
	);
	LUT2 #(
		.INIT('h8)
	) name5701 (
		\WX4730_reg/NET0131 ,
		\_2196__reg/NET0131 ,
		_w7209_
	);
	LUT2 #(
		.INIT('h1)
	) name5702 (
		_w7208_,
		_w7209_,
		_w7210_
	);
	LUT2 #(
		.INIT('h2)
	) name5703 (
		RESET_pad,
		_w7210_,
		_w7211_
	);
	LUT2 #(
		.INIT('h1)
	) name5704 (
		\WX4724_reg/NET0131 ,
		\_2199__reg/NET0131 ,
		_w7212_
	);
	LUT2 #(
		.INIT('h8)
	) name5705 (
		\WX4724_reg/NET0131 ,
		\_2199__reg/NET0131 ,
		_w7213_
	);
	LUT2 #(
		.INIT('h1)
	) name5706 (
		_w7212_,
		_w7213_,
		_w7214_
	);
	LUT2 #(
		.INIT('h2)
	) name5707 (
		RESET_pad,
		_w7214_,
		_w7215_
	);
	LUT2 #(
		.INIT('h1)
	) name5708 (
		\WX4722_reg/NET0131 ,
		\_2200__reg/NET0131 ,
		_w7216_
	);
	LUT2 #(
		.INIT('h8)
	) name5709 (
		\WX4722_reg/NET0131 ,
		\_2200__reg/NET0131 ,
		_w7217_
	);
	LUT2 #(
		.INIT('h1)
	) name5710 (
		_w7216_,
		_w7217_,
		_w7218_
	);
	LUT2 #(
		.INIT('h2)
	) name5711 (
		RESET_pad,
		_w7218_,
		_w7219_
	);
	LUT2 #(
		.INIT('h1)
	) name5712 (
		\WX4720_reg/NET0131 ,
		\_2201__reg/NET0131 ,
		_w7220_
	);
	LUT2 #(
		.INIT('h8)
	) name5713 (
		\WX4720_reg/NET0131 ,
		\_2201__reg/NET0131 ,
		_w7221_
	);
	LUT2 #(
		.INIT('h1)
	) name5714 (
		_w7220_,
		_w7221_,
		_w7222_
	);
	LUT2 #(
		.INIT('h2)
	) name5715 (
		RESET_pad,
		_w7222_,
		_w7223_
	);
	LUT2 #(
		.INIT('h1)
	) name5716 (
		\WX4718_reg/NET0131 ,
		\_2202__reg/NET0131 ,
		_w7224_
	);
	LUT2 #(
		.INIT('h8)
	) name5717 (
		\WX4718_reg/NET0131 ,
		\_2202__reg/NET0131 ,
		_w7225_
	);
	LUT2 #(
		.INIT('h1)
	) name5718 (
		_w7224_,
		_w7225_,
		_w7226_
	);
	LUT2 #(
		.INIT('h2)
	) name5719 (
		RESET_pad,
		_w7226_,
		_w7227_
	);
	LUT2 #(
		.INIT('h1)
	) name5720 (
		\WX4716_reg/NET0131 ,
		\_2203__reg/NET0131 ,
		_w7228_
	);
	LUT2 #(
		.INIT('h8)
	) name5721 (
		\WX4716_reg/NET0131 ,
		\_2203__reg/NET0131 ,
		_w7229_
	);
	LUT2 #(
		.INIT('h1)
	) name5722 (
		_w7228_,
		_w7229_,
		_w7230_
	);
	LUT2 #(
		.INIT('h2)
	) name5723 (
		RESET_pad,
		_w7230_,
		_w7231_
	);
	LUT2 #(
		.INIT('h1)
	) name5724 (
		\WX6071_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w7232_
	);
	LUT2 #(
		.INIT('h8)
	) name5725 (
		\WX6071_reg/NET0131 ,
		\_2236__reg/NET0131 ,
		_w7233_
	);
	LUT2 #(
		.INIT('h1)
	) name5726 (
		_w7232_,
		_w7233_,
		_w7234_
	);
	LUT2 #(
		.INIT('h2)
	) name5727 (
		RESET_pad,
		_w7234_,
		_w7235_
	);
	LUT2 #(
		.INIT('h1)
	) name5728 (
		\WX6067_reg/NET0131 ,
		\_2206__reg/NET0131 ,
		_w7236_
	);
	LUT2 #(
		.INIT('h8)
	) name5729 (
		\WX6067_reg/NET0131 ,
		\_2206__reg/NET0131 ,
		_w7237_
	);
	LUT2 #(
		.INIT('h1)
	) name5730 (
		_w7236_,
		_w7237_,
		_w7238_
	);
	LUT2 #(
		.INIT('h2)
	) name5731 (
		RESET_pad,
		_w7238_,
		_w7239_
	);
	LUT2 #(
		.INIT('h1)
	) name5732 (
		\WX6065_reg/NET0131 ,
		\_2207__reg/NET0131 ,
		_w7240_
	);
	LUT2 #(
		.INIT('h8)
	) name5733 (
		\WX6065_reg/NET0131 ,
		\_2207__reg/NET0131 ,
		_w7241_
	);
	LUT2 #(
		.INIT('h1)
	) name5734 (
		_w7240_,
		_w7241_,
		_w7242_
	);
	LUT2 #(
		.INIT('h2)
	) name5735 (
		RESET_pad,
		_w7242_,
		_w7243_
	);
	LUT2 #(
		.INIT('h1)
	) name5736 (
		\WX6059_reg/NET0131 ,
		\_2210__reg/NET0131 ,
		_w7244_
	);
	LUT2 #(
		.INIT('h8)
	) name5737 (
		\WX6059_reg/NET0131 ,
		\_2210__reg/NET0131 ,
		_w7245_
	);
	LUT2 #(
		.INIT('h1)
	) name5738 (
		_w7244_,
		_w7245_,
		_w7246_
	);
	LUT2 #(
		.INIT('h2)
	) name5739 (
		RESET_pad,
		_w7246_,
		_w7247_
	);
	LUT2 #(
		.INIT('h1)
	) name5740 (
		\WX6057_reg/NET0131 ,
		\_2211__reg/NET0131 ,
		_w7248_
	);
	LUT2 #(
		.INIT('h8)
	) name5741 (
		\WX6057_reg/NET0131 ,
		\_2211__reg/NET0131 ,
		_w7249_
	);
	LUT2 #(
		.INIT('h1)
	) name5742 (
		_w7248_,
		_w7249_,
		_w7250_
	);
	LUT2 #(
		.INIT('h2)
	) name5743 (
		RESET_pad,
		_w7250_,
		_w7251_
	);
	LUT2 #(
		.INIT('h1)
	) name5744 (
		\WX6055_reg/NET0131 ,
		\_2212__reg/NET0131 ,
		_w7252_
	);
	LUT2 #(
		.INIT('h8)
	) name5745 (
		\WX6055_reg/NET0131 ,
		\_2212__reg/NET0131 ,
		_w7253_
	);
	LUT2 #(
		.INIT('h1)
	) name5746 (
		_w7252_,
		_w7253_,
		_w7254_
	);
	LUT2 #(
		.INIT('h2)
	) name5747 (
		RESET_pad,
		_w7254_,
		_w7255_
	);
	LUT2 #(
		.INIT('h1)
	) name5748 (
		\WX6053_reg/NET0131 ,
		\_2213__reg/NET0131 ,
		_w7256_
	);
	LUT2 #(
		.INIT('h8)
	) name5749 (
		\WX6053_reg/NET0131 ,
		\_2213__reg/NET0131 ,
		_w7257_
	);
	LUT2 #(
		.INIT('h1)
	) name5750 (
		_w7256_,
		_w7257_,
		_w7258_
	);
	LUT2 #(
		.INIT('h2)
	) name5751 (
		RESET_pad,
		_w7258_,
		_w7259_
	);
	LUT2 #(
		.INIT('h1)
	) name5752 (
		\WX6051_reg/NET0131 ,
		\_2214__reg/NET0131 ,
		_w7260_
	);
	LUT2 #(
		.INIT('h8)
	) name5753 (
		\WX6051_reg/NET0131 ,
		\_2214__reg/NET0131 ,
		_w7261_
	);
	LUT2 #(
		.INIT('h1)
	) name5754 (
		_w7260_,
		_w7261_,
		_w7262_
	);
	LUT2 #(
		.INIT('h2)
	) name5755 (
		RESET_pad,
		_w7262_,
		_w7263_
	);
	LUT2 #(
		.INIT('h1)
	) name5756 (
		\WX6047_reg/NET0131 ,
		\_2216__reg/NET0131 ,
		_w7264_
	);
	LUT2 #(
		.INIT('h8)
	) name5757 (
		\WX6047_reg/NET0131 ,
		\_2216__reg/NET0131 ,
		_w7265_
	);
	LUT2 #(
		.INIT('h1)
	) name5758 (
		_w7264_,
		_w7265_,
		_w7266_
	);
	LUT2 #(
		.INIT('h2)
	) name5759 (
		RESET_pad,
		_w7266_,
		_w7267_
	);
	LUT2 #(
		.INIT('h1)
	) name5760 (
		\WX6045_reg/NET0131 ,
		\_2217__reg/NET0131 ,
		_w7268_
	);
	LUT2 #(
		.INIT('h8)
	) name5761 (
		\WX6045_reg/NET0131 ,
		\_2217__reg/NET0131 ,
		_w7269_
	);
	LUT2 #(
		.INIT('h1)
	) name5762 (
		_w7268_,
		_w7269_,
		_w7270_
	);
	LUT2 #(
		.INIT('h2)
	) name5763 (
		RESET_pad,
		_w7270_,
		_w7271_
	);
	LUT2 #(
		.INIT('h1)
	) name5764 (
		\WX6035_reg/NET0131 ,
		\_2222__reg/NET0131 ,
		_w7272_
	);
	LUT2 #(
		.INIT('h8)
	) name5765 (
		\WX6035_reg/NET0131 ,
		\_2222__reg/NET0131 ,
		_w7273_
	);
	LUT2 #(
		.INIT('h1)
	) name5766 (
		_w7272_,
		_w7273_,
		_w7274_
	);
	LUT2 #(
		.INIT('h2)
	) name5767 (
		RESET_pad,
		_w7274_,
		_w7275_
	);
	LUT2 #(
		.INIT('h1)
	) name5768 (
		\WX6033_reg/NET0131 ,
		\_2223__reg/NET0131 ,
		_w7276_
	);
	LUT2 #(
		.INIT('h8)
	) name5769 (
		\WX6033_reg/NET0131 ,
		\_2223__reg/NET0131 ,
		_w7277_
	);
	LUT2 #(
		.INIT('h1)
	) name5770 (
		_w7276_,
		_w7277_,
		_w7278_
	);
	LUT2 #(
		.INIT('h2)
	) name5771 (
		RESET_pad,
		_w7278_,
		_w7279_
	);
	LUT2 #(
		.INIT('h1)
	) name5772 (
		\WX6031_reg/NET0131 ,
		\_2224__reg/NET0131 ,
		_w7280_
	);
	LUT2 #(
		.INIT('h8)
	) name5773 (
		\WX6031_reg/NET0131 ,
		\_2224__reg/NET0131 ,
		_w7281_
	);
	LUT2 #(
		.INIT('h1)
	) name5774 (
		_w7280_,
		_w7281_,
		_w7282_
	);
	LUT2 #(
		.INIT('h2)
	) name5775 (
		RESET_pad,
		_w7282_,
		_w7283_
	);
	LUT2 #(
		.INIT('h1)
	) name5776 (
		\WX6029_reg/NET0131 ,
		\_2225__reg/NET0131 ,
		_w7284_
	);
	LUT2 #(
		.INIT('h8)
	) name5777 (
		\WX6029_reg/NET0131 ,
		\_2225__reg/NET0131 ,
		_w7285_
	);
	LUT2 #(
		.INIT('h1)
	) name5778 (
		_w7284_,
		_w7285_,
		_w7286_
	);
	LUT2 #(
		.INIT('h2)
	) name5779 (
		RESET_pad,
		_w7286_,
		_w7287_
	);
	LUT2 #(
		.INIT('h1)
	) name5780 (
		\WX6023_reg/NET0131 ,
		\_2228__reg/NET0131 ,
		_w7288_
	);
	LUT2 #(
		.INIT('h8)
	) name5781 (
		\WX6023_reg/NET0131 ,
		\_2228__reg/NET0131 ,
		_w7289_
	);
	LUT2 #(
		.INIT('h1)
	) name5782 (
		_w7288_,
		_w7289_,
		_w7290_
	);
	LUT2 #(
		.INIT('h2)
	) name5783 (
		RESET_pad,
		_w7290_,
		_w7291_
	);
	LUT2 #(
		.INIT('h1)
	) name5784 (
		\WX6021_reg/NET0131 ,
		\_2229__reg/NET0131 ,
		_w7292_
	);
	LUT2 #(
		.INIT('h8)
	) name5785 (
		\WX6021_reg/NET0131 ,
		\_2229__reg/NET0131 ,
		_w7293_
	);
	LUT2 #(
		.INIT('h1)
	) name5786 (
		_w7292_,
		_w7293_,
		_w7294_
	);
	LUT2 #(
		.INIT('h2)
	) name5787 (
		RESET_pad,
		_w7294_,
		_w7295_
	);
	LUT2 #(
		.INIT('h1)
	) name5788 (
		\WX6019_reg/NET0131 ,
		\_2230__reg/NET0131 ,
		_w7296_
	);
	LUT2 #(
		.INIT('h8)
	) name5789 (
		\WX6019_reg/NET0131 ,
		\_2230__reg/NET0131 ,
		_w7297_
	);
	LUT2 #(
		.INIT('h1)
	) name5790 (
		_w7296_,
		_w7297_,
		_w7298_
	);
	LUT2 #(
		.INIT('h2)
	) name5791 (
		RESET_pad,
		_w7298_,
		_w7299_
	);
	LUT2 #(
		.INIT('h1)
	) name5792 (
		\WX6015_reg/NET0131 ,
		\_2232__reg/NET0131 ,
		_w7300_
	);
	LUT2 #(
		.INIT('h8)
	) name5793 (
		\WX6015_reg/NET0131 ,
		\_2232__reg/NET0131 ,
		_w7301_
	);
	LUT2 #(
		.INIT('h1)
	) name5794 (
		_w7300_,
		_w7301_,
		_w7302_
	);
	LUT2 #(
		.INIT('h2)
	) name5795 (
		RESET_pad,
		_w7302_,
		_w7303_
	);
	LUT2 #(
		.INIT('h1)
	) name5796 (
		\WX6011_reg/NET0131 ,
		\_2234__reg/NET0131 ,
		_w7304_
	);
	LUT2 #(
		.INIT('h8)
	) name5797 (
		\WX6011_reg/NET0131 ,
		\_2234__reg/NET0131 ,
		_w7305_
	);
	LUT2 #(
		.INIT('h1)
	) name5798 (
		_w7304_,
		_w7305_,
		_w7306_
	);
	LUT2 #(
		.INIT('h2)
	) name5799 (
		RESET_pad,
		_w7306_,
		_w7307_
	);
	LUT2 #(
		.INIT('h1)
	) name5800 (
		\WX6009_reg/NET0131 ,
		\_2235__reg/NET0131 ,
		_w7308_
	);
	LUT2 #(
		.INIT('h8)
	) name5801 (
		\WX6009_reg/NET0131 ,
		\_2235__reg/NET0131 ,
		_w7309_
	);
	LUT2 #(
		.INIT('h1)
	) name5802 (
		_w7308_,
		_w7309_,
		_w7310_
	);
	LUT2 #(
		.INIT('h2)
	) name5803 (
		RESET_pad,
		_w7310_,
		_w7311_
	);
	LUT2 #(
		.INIT('h1)
	) name5804 (
		\WX7364_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w7312_
	);
	LUT2 #(
		.INIT('h8)
	) name5805 (
		\WX7364_reg/NET0131 ,
		\_2268__reg/NET0131 ,
		_w7313_
	);
	LUT2 #(
		.INIT('h1)
	) name5806 (
		_w7312_,
		_w7313_,
		_w7314_
	);
	LUT2 #(
		.INIT('h2)
	) name5807 (
		RESET_pad,
		_w7314_,
		_w7315_
	);
	LUT2 #(
		.INIT('h1)
	) name5808 (
		\WX7360_reg/NET0131 ,
		\_2238__reg/NET0131 ,
		_w7316_
	);
	LUT2 #(
		.INIT('h8)
	) name5809 (
		\WX7360_reg/NET0131 ,
		\_2238__reg/NET0131 ,
		_w7317_
	);
	LUT2 #(
		.INIT('h1)
	) name5810 (
		_w7316_,
		_w7317_,
		_w7318_
	);
	LUT2 #(
		.INIT('h2)
	) name5811 (
		RESET_pad,
		_w7318_,
		_w7319_
	);
	LUT2 #(
		.INIT('h1)
	) name5812 (
		\WX7358_reg/NET0131 ,
		\_2239__reg/NET0131 ,
		_w7320_
	);
	LUT2 #(
		.INIT('h8)
	) name5813 (
		\WX7358_reg/NET0131 ,
		\_2239__reg/NET0131 ,
		_w7321_
	);
	LUT2 #(
		.INIT('h1)
	) name5814 (
		_w7320_,
		_w7321_,
		_w7322_
	);
	LUT2 #(
		.INIT('h2)
	) name5815 (
		RESET_pad,
		_w7322_,
		_w7323_
	);
	LUT2 #(
		.INIT('h1)
	) name5816 (
		\WX7354_reg/NET0131 ,
		\_2241__reg/NET0131 ,
		_w7324_
	);
	LUT2 #(
		.INIT('h8)
	) name5817 (
		\WX7354_reg/NET0131 ,
		\_2241__reg/NET0131 ,
		_w7325_
	);
	LUT2 #(
		.INIT('h1)
	) name5818 (
		_w7324_,
		_w7325_,
		_w7326_
	);
	LUT2 #(
		.INIT('h2)
	) name5819 (
		RESET_pad,
		_w7326_,
		_w7327_
	);
	LUT2 #(
		.INIT('h1)
	) name5820 (
		\WX7352_reg/NET0131 ,
		\_2242__reg/NET0131 ,
		_w7328_
	);
	LUT2 #(
		.INIT('h8)
	) name5821 (
		\WX7352_reg/NET0131 ,
		\_2242__reg/NET0131 ,
		_w7329_
	);
	LUT2 #(
		.INIT('h1)
	) name5822 (
		_w7328_,
		_w7329_,
		_w7330_
	);
	LUT2 #(
		.INIT('h2)
	) name5823 (
		RESET_pad,
		_w7330_,
		_w7331_
	);
	LUT2 #(
		.INIT('h1)
	) name5824 (
		\WX6025_reg/NET0131 ,
		\_2227__reg/NET0131 ,
		_w7332_
	);
	LUT2 #(
		.INIT('h8)
	) name5825 (
		\WX6025_reg/NET0131 ,
		\_2227__reg/NET0131 ,
		_w7333_
	);
	LUT2 #(
		.INIT('h1)
	) name5826 (
		_w7332_,
		_w7333_,
		_w7334_
	);
	LUT2 #(
		.INIT('h2)
	) name5827 (
		RESET_pad,
		_w7334_,
		_w7335_
	);
	LUT2 #(
		.INIT('h1)
	) name5828 (
		\WX8647_reg/NET0131 ,
		\_2273__reg/NET0131 ,
		_w7336_
	);
	LUT2 #(
		.INIT('h8)
	) name5829 (
		\WX8647_reg/NET0131 ,
		\_2273__reg/NET0131 ,
		_w7337_
	);
	LUT2 #(
		.INIT('h1)
	) name5830 (
		_w7336_,
		_w7337_,
		_w7338_
	);
	LUT2 #(
		.INIT('h2)
	) name5831 (
		RESET_pad,
		_w7338_,
		_w7339_
	);
	LUT2 #(
		.INIT('h1)
	) name5832 (
		\WX7336_reg/NET0131 ,
		\_2250__reg/NET0131 ,
		_w7340_
	);
	LUT2 #(
		.INIT('h8)
	) name5833 (
		\WX7336_reg/NET0131 ,
		\_2250__reg/NET0131 ,
		_w7341_
	);
	LUT2 #(
		.INIT('h1)
	) name5834 (
		_w7340_,
		_w7341_,
		_w7342_
	);
	LUT2 #(
		.INIT('h2)
	) name5835 (
		RESET_pad,
		_w7342_,
		_w7343_
	);
	LUT2 #(
		.INIT('h1)
	) name5836 (
		\WX7330_reg/NET0131 ,
		\_2253__reg/NET0131 ,
		_w7344_
	);
	LUT2 #(
		.INIT('h8)
	) name5837 (
		\WX7330_reg/NET0131 ,
		\_2253__reg/NET0131 ,
		_w7345_
	);
	LUT2 #(
		.INIT('h1)
	) name5838 (
		_w7344_,
		_w7345_,
		_w7346_
	);
	LUT2 #(
		.INIT('h2)
	) name5839 (
		RESET_pad,
		_w7346_,
		_w7347_
	);
	LUT2 #(
		.INIT('h1)
	) name5840 (
		\WX7326_reg/NET0131 ,
		\_2255__reg/NET0131 ,
		_w7348_
	);
	LUT2 #(
		.INIT('h8)
	) name5841 (
		\WX7326_reg/NET0131 ,
		\_2255__reg/NET0131 ,
		_w7349_
	);
	LUT2 #(
		.INIT('h1)
	) name5842 (
		_w7348_,
		_w7349_,
		_w7350_
	);
	LUT2 #(
		.INIT('h2)
	) name5843 (
		RESET_pad,
		_w7350_,
		_w7351_
	);
	LUT2 #(
		.INIT('h1)
	) name5844 (
		\WX7322_reg/NET0131 ,
		\_2257__reg/NET0131 ,
		_w7352_
	);
	LUT2 #(
		.INIT('h8)
	) name5845 (
		\WX7322_reg/NET0131 ,
		\_2257__reg/NET0131 ,
		_w7353_
	);
	LUT2 #(
		.INIT('h1)
	) name5846 (
		_w7352_,
		_w7353_,
		_w7354_
	);
	LUT2 #(
		.INIT('h2)
	) name5847 (
		RESET_pad,
		_w7354_,
		_w7355_
	);
	LUT2 #(
		.INIT('h1)
	) name5848 (
		\WX7320_reg/NET0131 ,
		\_2258__reg/NET0131 ,
		_w7356_
	);
	LUT2 #(
		.INIT('h8)
	) name5849 (
		\WX7320_reg/NET0131 ,
		\_2258__reg/NET0131 ,
		_w7357_
	);
	LUT2 #(
		.INIT('h1)
	) name5850 (
		_w7356_,
		_w7357_,
		_w7358_
	);
	LUT2 #(
		.INIT('h2)
	) name5851 (
		RESET_pad,
		_w7358_,
		_w7359_
	);
	LUT2 #(
		.INIT('h1)
	) name5852 (
		\WX7318_reg/NET0131 ,
		\_2259__reg/NET0131 ,
		_w7360_
	);
	LUT2 #(
		.INIT('h8)
	) name5853 (
		\WX7318_reg/NET0131 ,
		\_2259__reg/NET0131 ,
		_w7361_
	);
	LUT2 #(
		.INIT('h1)
	) name5854 (
		_w7360_,
		_w7361_,
		_w7362_
	);
	LUT2 #(
		.INIT('h2)
	) name5855 (
		RESET_pad,
		_w7362_,
		_w7363_
	);
	LUT2 #(
		.INIT('h1)
	) name5856 (
		\WX6069_reg/NET0131 ,
		\_2205__reg/NET0131 ,
		_w7364_
	);
	LUT2 #(
		.INIT('h8)
	) name5857 (
		\WX6069_reg/NET0131 ,
		\_2205__reg/NET0131 ,
		_w7365_
	);
	LUT2 #(
		.INIT('h1)
	) name5858 (
		_w7364_,
		_w7365_,
		_w7366_
	);
	LUT2 #(
		.INIT('h2)
	) name5859 (
		RESET_pad,
		_w7366_,
		_w7367_
	);
	LUT2 #(
		.INIT('h1)
	) name5860 (
		\WX7314_reg/NET0131 ,
		\_2261__reg/NET0131 ,
		_w7368_
	);
	LUT2 #(
		.INIT('h8)
	) name5861 (
		\WX7314_reg/NET0131 ,
		\_2261__reg/NET0131 ,
		_w7369_
	);
	LUT2 #(
		.INIT('h1)
	) name5862 (
		_w7368_,
		_w7369_,
		_w7370_
	);
	LUT2 #(
		.INIT('h2)
	) name5863 (
		RESET_pad,
		_w7370_,
		_w7371_
	);
	LUT2 #(
		.INIT('h1)
	) name5864 (
		\WX6017_reg/NET0131 ,
		\_2231__reg/NET0131 ,
		_w7372_
	);
	LUT2 #(
		.INIT('h8)
	) name5865 (
		\WX6017_reg/NET0131 ,
		\_2231__reg/NET0131 ,
		_w7373_
	);
	LUT2 #(
		.INIT('h1)
	) name5866 (
		_w7372_,
		_w7373_,
		_w7374_
	);
	LUT2 #(
		.INIT('h2)
	) name5867 (
		RESET_pad,
		_w7374_,
		_w7375_
	);
	LUT2 #(
		.INIT('h1)
	) name5868 (
		\WX6027_reg/NET0131 ,
		\_2226__reg/NET0131 ,
		_w7376_
	);
	LUT2 #(
		.INIT('h8)
	) name5869 (
		\WX6027_reg/NET0131 ,
		\_2226__reg/NET0131 ,
		_w7377_
	);
	LUT2 #(
		.INIT('h1)
	) name5870 (
		_w7376_,
		_w7377_,
		_w7378_
	);
	LUT2 #(
		.INIT('h2)
	) name5871 (
		RESET_pad,
		_w7378_,
		_w7379_
	);
	LUT2 #(
		.INIT('h1)
	) name5872 (
		\WX7306_reg/NET0131 ,
		\_2265__reg/NET0131 ,
		_w7380_
	);
	LUT2 #(
		.INIT('h8)
	) name5873 (
		\WX7306_reg/NET0131 ,
		\_2265__reg/NET0131 ,
		_w7381_
	);
	LUT2 #(
		.INIT('h1)
	) name5874 (
		_w7380_,
		_w7381_,
		_w7382_
	);
	LUT2 #(
		.INIT('h2)
	) name5875 (
		RESET_pad,
		_w7382_,
		_w7383_
	);
	LUT2 #(
		.INIT('h1)
	) name5876 (
		\WX7302_reg/NET0131 ,
		\_2267__reg/NET0131 ,
		_w7384_
	);
	LUT2 #(
		.INIT('h8)
	) name5877 (
		\WX7302_reg/NET0131 ,
		\_2267__reg/NET0131 ,
		_w7385_
	);
	LUT2 #(
		.INIT('h1)
	) name5878 (
		_w7384_,
		_w7385_,
		_w7386_
	);
	LUT2 #(
		.INIT('h2)
	) name5879 (
		RESET_pad,
		_w7386_,
		_w7387_
	);
	LUT2 #(
		.INIT('h1)
	) name5880 (
		\WX8655_reg/NET0131 ,
		\_2269__reg/NET0131 ,
		_w7388_
	);
	LUT2 #(
		.INIT('h8)
	) name5881 (
		\WX8655_reg/NET0131 ,
		\_2269__reg/NET0131 ,
		_w7389_
	);
	LUT2 #(
		.INIT('h1)
	) name5882 (
		_w7388_,
		_w7389_,
		_w7390_
	);
	LUT2 #(
		.INIT('h2)
	) name5883 (
		RESET_pad,
		_w7390_,
		_w7391_
	);
	LUT2 #(
		.INIT('h1)
	) name5884 (
		\WX8653_reg/NET0131 ,
		\_2270__reg/NET0131 ,
		_w7392_
	);
	LUT2 #(
		.INIT('h8)
	) name5885 (
		\WX8653_reg/NET0131 ,
		\_2270__reg/NET0131 ,
		_w7393_
	);
	LUT2 #(
		.INIT('h1)
	) name5886 (
		_w7392_,
		_w7393_,
		_w7394_
	);
	LUT2 #(
		.INIT('h2)
	) name5887 (
		RESET_pad,
		_w7394_,
		_w7395_
	);
	LUT2 #(
		.INIT('h1)
	) name5888 (
		\WX8651_reg/NET0131 ,
		\_2271__reg/NET0131 ,
		_w7396_
	);
	LUT2 #(
		.INIT('h8)
	) name5889 (
		\WX8651_reg/NET0131 ,
		\_2271__reg/NET0131 ,
		_w7397_
	);
	LUT2 #(
		.INIT('h1)
	) name5890 (
		_w7396_,
		_w7397_,
		_w7398_
	);
	LUT2 #(
		.INIT('h2)
	) name5891 (
		RESET_pad,
		_w7398_,
		_w7399_
	);
	LUT2 #(
		.INIT('h1)
	) name5892 (
		\WX8645_reg/NET0131 ,
		\_2274__reg/NET0131 ,
		_w7400_
	);
	LUT2 #(
		.INIT('h8)
	) name5893 (
		\WX8645_reg/NET0131 ,
		\_2274__reg/NET0131 ,
		_w7401_
	);
	LUT2 #(
		.INIT('h1)
	) name5894 (
		_w7400_,
		_w7401_,
		_w7402_
	);
	LUT2 #(
		.INIT('h2)
	) name5895 (
		RESET_pad,
		_w7402_,
		_w7403_
	);
	LUT2 #(
		.INIT('h1)
	) name5896 (
		\WX8641_reg/NET0131 ,
		\_2276__reg/NET0131 ,
		_w7404_
	);
	LUT2 #(
		.INIT('h8)
	) name5897 (
		\WX8641_reg/NET0131 ,
		\_2276__reg/NET0131 ,
		_w7405_
	);
	LUT2 #(
		.INIT('h1)
	) name5898 (
		_w7404_,
		_w7405_,
		_w7406_
	);
	LUT2 #(
		.INIT('h2)
	) name5899 (
		RESET_pad,
		_w7406_,
		_w7407_
	);
	LUT2 #(
		.INIT('h1)
	) name5900 (
		\WX8637_reg/NET0131 ,
		\_2278__reg/NET0131 ,
		_w7408_
	);
	LUT2 #(
		.INIT('h8)
	) name5901 (
		\WX8637_reg/NET0131 ,
		\_2278__reg/NET0131 ,
		_w7409_
	);
	LUT2 #(
		.INIT('h1)
	) name5902 (
		_w7408_,
		_w7409_,
		_w7410_
	);
	LUT2 #(
		.INIT('h2)
	) name5903 (
		RESET_pad,
		_w7410_,
		_w7411_
	);
	LUT2 #(
		.INIT('h1)
	) name5904 (
		\WX8631_reg/NET0131 ,
		\_2281__reg/NET0131 ,
		_w7412_
	);
	LUT2 #(
		.INIT('h8)
	) name5905 (
		\WX8631_reg/NET0131 ,
		\_2281__reg/NET0131 ,
		_w7413_
	);
	LUT2 #(
		.INIT('h1)
	) name5906 (
		_w7412_,
		_w7413_,
		_w7414_
	);
	LUT2 #(
		.INIT('h2)
	) name5907 (
		RESET_pad,
		_w7414_,
		_w7415_
	);
	LUT2 #(
		.INIT('h1)
	) name5908 (
		\WX8629_reg/NET0131 ,
		\_2282__reg/NET0131 ,
		_w7416_
	);
	LUT2 #(
		.INIT('h8)
	) name5909 (
		\WX8629_reg/NET0131 ,
		\_2282__reg/NET0131 ,
		_w7417_
	);
	LUT2 #(
		.INIT('h1)
	) name5910 (
		_w7416_,
		_w7417_,
		_w7418_
	);
	LUT2 #(
		.INIT('h2)
	) name5911 (
		RESET_pad,
		_w7418_,
		_w7419_
	);
	LUT2 #(
		.INIT('h1)
	) name5912 (
		\WX8627_reg/NET0131 ,
		\_2283__reg/NET0131 ,
		_w7420_
	);
	LUT2 #(
		.INIT('h8)
	) name5913 (
		\WX8627_reg/NET0131 ,
		\_2283__reg/NET0131 ,
		_w7421_
	);
	LUT2 #(
		.INIT('h1)
	) name5914 (
		_w7420_,
		_w7421_,
		_w7422_
	);
	LUT2 #(
		.INIT('h2)
	) name5915 (
		RESET_pad,
		_w7422_,
		_w7423_
	);
	LUT2 #(
		.INIT('h1)
	) name5916 (
		\WX8621_reg/NET0131 ,
		\_2286__reg/NET0131 ,
		_w7424_
	);
	LUT2 #(
		.INIT('h8)
	) name5917 (
		\WX8621_reg/NET0131 ,
		\_2286__reg/NET0131 ,
		_w7425_
	);
	LUT2 #(
		.INIT('h1)
	) name5918 (
		_w7424_,
		_w7425_,
		_w7426_
	);
	LUT2 #(
		.INIT('h2)
	) name5919 (
		RESET_pad,
		_w7426_,
		_w7427_
	);
	LUT2 #(
		.INIT('h1)
	) name5920 (
		\WX8617_reg/NET0131 ,
		\_2288__reg/NET0131 ,
		_w7428_
	);
	LUT2 #(
		.INIT('h8)
	) name5921 (
		\WX8617_reg/NET0131 ,
		\_2288__reg/NET0131 ,
		_w7429_
	);
	LUT2 #(
		.INIT('h1)
	) name5922 (
		_w7428_,
		_w7429_,
		_w7430_
	);
	LUT2 #(
		.INIT('h2)
	) name5923 (
		RESET_pad,
		_w7430_,
		_w7431_
	);
	LUT2 #(
		.INIT('h1)
	) name5924 (
		\WX8615_reg/NET0131 ,
		\_2289__reg/NET0131 ,
		_w7432_
	);
	LUT2 #(
		.INIT('h8)
	) name5925 (
		\WX8615_reg/NET0131 ,
		\_2289__reg/NET0131 ,
		_w7433_
	);
	LUT2 #(
		.INIT('h1)
	) name5926 (
		_w7432_,
		_w7433_,
		_w7434_
	);
	LUT2 #(
		.INIT('h2)
	) name5927 (
		RESET_pad,
		_w7434_,
		_w7435_
	);
	LUT2 #(
		.INIT('h1)
	) name5928 (
		\WX8613_reg/NET0131 ,
		\_2290__reg/NET0131 ,
		_w7436_
	);
	LUT2 #(
		.INIT('h8)
	) name5929 (
		\WX8613_reg/NET0131 ,
		\_2290__reg/NET0131 ,
		_w7437_
	);
	LUT2 #(
		.INIT('h1)
	) name5930 (
		_w7436_,
		_w7437_,
		_w7438_
	);
	LUT2 #(
		.INIT('h2)
	) name5931 (
		RESET_pad,
		_w7438_,
		_w7439_
	);
	LUT2 #(
		.INIT('h1)
	) name5932 (
		\WX8611_reg/NET0131 ,
		\_2291__reg/NET0131 ,
		_w7440_
	);
	LUT2 #(
		.INIT('h8)
	) name5933 (
		\WX8611_reg/NET0131 ,
		\_2291__reg/NET0131 ,
		_w7441_
	);
	LUT2 #(
		.INIT('h1)
	) name5934 (
		_w7440_,
		_w7441_,
		_w7442_
	);
	LUT2 #(
		.INIT('h2)
	) name5935 (
		RESET_pad,
		_w7442_,
		_w7443_
	);
	LUT2 #(
		.INIT('h1)
	) name5936 (
		\WX8609_reg/NET0131 ,
		\_2292__reg/NET0131 ,
		_w7444_
	);
	LUT2 #(
		.INIT('h8)
	) name5937 (
		\WX8609_reg/NET0131 ,
		\_2292__reg/NET0131 ,
		_w7445_
	);
	LUT2 #(
		.INIT('h1)
	) name5938 (
		_w7444_,
		_w7445_,
		_w7446_
	);
	LUT2 #(
		.INIT('h2)
	) name5939 (
		RESET_pad,
		_w7446_,
		_w7447_
	);
	LUT2 #(
		.INIT('h1)
	) name5940 (
		\WX8597_reg/NET0131 ,
		\_2298__reg/NET0131 ,
		_w7448_
	);
	LUT2 #(
		.INIT('h8)
	) name5941 (
		\WX8597_reg/NET0131 ,
		\_2298__reg/NET0131 ,
		_w7449_
	);
	LUT2 #(
		.INIT('h1)
	) name5942 (
		_w7448_,
		_w7449_,
		_w7450_
	);
	LUT2 #(
		.INIT('h2)
	) name5943 (
		RESET_pad,
		_w7450_,
		_w7451_
	);
	LUT2 #(
		.INIT('h1)
	) name5944 (
		\WX8595_reg/NET0131 ,
		\_2299__reg/NET0131 ,
		_w7452_
	);
	LUT2 #(
		.INIT('h8)
	) name5945 (
		\WX8595_reg/NET0131 ,
		\_2299__reg/NET0131 ,
		_w7453_
	);
	LUT2 #(
		.INIT('h1)
	) name5946 (
		_w7452_,
		_w7453_,
		_w7454_
	);
	LUT2 #(
		.INIT('h2)
	) name5947 (
		RESET_pad,
		_w7454_,
		_w7455_
	);
	LUT2 #(
		.INIT('h1)
	) name5948 (
		\WX9950_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w7456_
	);
	LUT2 #(
		.INIT('h8)
	) name5949 (
		\WX9950_reg/NET0131 ,
		\_2332__reg/NET0131 ,
		_w7457_
	);
	LUT2 #(
		.INIT('h1)
	) name5950 (
		_w7456_,
		_w7457_,
		_w7458_
	);
	LUT2 #(
		.INIT('h2)
	) name5951 (
		RESET_pad,
		_w7458_,
		_w7459_
	);
	LUT2 #(
		.INIT('h1)
	) name5952 (
		\WX9948_reg/NET0131 ,
		\_2301__reg/NET0131 ,
		_w7460_
	);
	LUT2 #(
		.INIT('h8)
	) name5953 (
		\WX9948_reg/NET0131 ,
		\_2301__reg/NET0131 ,
		_w7461_
	);
	LUT2 #(
		.INIT('h1)
	) name5954 (
		_w7460_,
		_w7461_,
		_w7462_
	);
	LUT2 #(
		.INIT('h2)
	) name5955 (
		RESET_pad,
		_w7462_,
		_w7463_
	);
	LUT2 #(
		.INIT('h1)
	) name5956 (
		\WX9946_reg/NET0131 ,
		\_2302__reg/NET0131 ,
		_w7464_
	);
	LUT2 #(
		.INIT('h8)
	) name5957 (
		\WX9946_reg/NET0131 ,
		\_2302__reg/NET0131 ,
		_w7465_
	);
	LUT2 #(
		.INIT('h1)
	) name5958 (
		_w7464_,
		_w7465_,
		_w7466_
	);
	LUT2 #(
		.INIT('h2)
	) name5959 (
		RESET_pad,
		_w7466_,
		_w7467_
	);
	LUT2 #(
		.INIT('h1)
	) name5960 (
		\WX9940_reg/NET0131 ,
		\_2305__reg/NET0131 ,
		_w7468_
	);
	LUT2 #(
		.INIT('h8)
	) name5961 (
		\WX9940_reg/NET0131 ,
		\_2305__reg/NET0131 ,
		_w7469_
	);
	LUT2 #(
		.INIT('h1)
	) name5962 (
		_w7468_,
		_w7469_,
		_w7470_
	);
	LUT2 #(
		.INIT('h2)
	) name5963 (
		RESET_pad,
		_w7470_,
		_w7471_
	);
	LUT2 #(
		.INIT('h1)
	) name5964 (
		\WX9938_reg/NET0131 ,
		\_2306__reg/NET0131 ,
		_w7472_
	);
	LUT2 #(
		.INIT('h8)
	) name5965 (
		\WX9938_reg/NET0131 ,
		\_2306__reg/NET0131 ,
		_w7473_
	);
	LUT2 #(
		.INIT('h1)
	) name5966 (
		_w7472_,
		_w7473_,
		_w7474_
	);
	LUT2 #(
		.INIT('h2)
	) name5967 (
		RESET_pad,
		_w7474_,
		_w7475_
	);
	LUT2 #(
		.INIT('h1)
	) name5968 (
		\WX9932_reg/NET0131 ,
		\_2309__reg/NET0131 ,
		_w7476_
	);
	LUT2 #(
		.INIT('h8)
	) name5969 (
		\WX9932_reg/NET0131 ,
		\_2309__reg/NET0131 ,
		_w7477_
	);
	LUT2 #(
		.INIT('h1)
	) name5970 (
		_w7476_,
		_w7477_,
		_w7478_
	);
	LUT2 #(
		.INIT('h2)
	) name5971 (
		RESET_pad,
		_w7478_,
		_w7479_
	);
	LUT2 #(
		.INIT('h1)
	) name5972 (
		\WX9926_reg/NET0131 ,
		\_2312__reg/NET0131 ,
		_w7480_
	);
	LUT2 #(
		.INIT('h8)
	) name5973 (
		\WX9926_reg/NET0131 ,
		\_2312__reg/NET0131 ,
		_w7481_
	);
	LUT2 #(
		.INIT('h1)
	) name5974 (
		_w7480_,
		_w7481_,
		_w7482_
	);
	LUT2 #(
		.INIT('h2)
	) name5975 (
		RESET_pad,
		_w7482_,
		_w7483_
	);
	LUT2 #(
		.INIT('h1)
	) name5976 (
		\WX9922_reg/NET0131 ,
		\_2314__reg/NET0131 ,
		_w7484_
	);
	LUT2 #(
		.INIT('h8)
	) name5977 (
		\WX9922_reg/NET0131 ,
		\_2314__reg/NET0131 ,
		_w7485_
	);
	LUT2 #(
		.INIT('h1)
	) name5978 (
		_w7484_,
		_w7485_,
		_w7486_
	);
	LUT2 #(
		.INIT('h2)
	) name5979 (
		RESET_pad,
		_w7486_,
		_w7487_
	);
	LUT2 #(
		.INIT('h1)
	) name5980 (
		\WX9920_reg/NET0131 ,
		\_2315__reg/NET0131 ,
		_w7488_
	);
	LUT2 #(
		.INIT('h8)
	) name5981 (
		\WX9920_reg/NET0131 ,
		\_2315__reg/NET0131 ,
		_w7489_
	);
	LUT2 #(
		.INIT('h1)
	) name5982 (
		_w7488_,
		_w7489_,
		_w7490_
	);
	LUT2 #(
		.INIT('h2)
	) name5983 (
		RESET_pad,
		_w7490_,
		_w7491_
	);
	LUT2 #(
		.INIT('h1)
	) name5984 (
		\WX9916_reg/NET0131 ,
		\_2317__reg/NET0131 ,
		_w7492_
	);
	LUT2 #(
		.INIT('h8)
	) name5985 (
		\WX9916_reg/NET0131 ,
		\_2317__reg/NET0131 ,
		_w7493_
	);
	LUT2 #(
		.INIT('h1)
	) name5986 (
		_w7492_,
		_w7493_,
		_w7494_
	);
	LUT2 #(
		.INIT('h2)
	) name5987 (
		RESET_pad,
		_w7494_,
		_w7495_
	);
	LUT2 #(
		.INIT('h1)
	) name5988 (
		\WX9914_reg/NET0131 ,
		\_2318__reg/NET0131 ,
		_w7496_
	);
	LUT2 #(
		.INIT('h8)
	) name5989 (
		\WX9914_reg/NET0131 ,
		\_2318__reg/NET0131 ,
		_w7497_
	);
	LUT2 #(
		.INIT('h1)
	) name5990 (
		_w7496_,
		_w7497_,
		_w7498_
	);
	LUT2 #(
		.INIT('h2)
	) name5991 (
		RESET_pad,
		_w7498_,
		_w7499_
	);
	LUT2 #(
		.INIT('h1)
	) name5992 (
		\WX9912_reg/NET0131 ,
		\_2319__reg/NET0131 ,
		_w7500_
	);
	LUT2 #(
		.INIT('h8)
	) name5993 (
		\WX9912_reg/NET0131 ,
		\_2319__reg/NET0131 ,
		_w7501_
	);
	LUT2 #(
		.INIT('h1)
	) name5994 (
		_w7500_,
		_w7501_,
		_w7502_
	);
	LUT2 #(
		.INIT('h2)
	) name5995 (
		RESET_pad,
		_w7502_,
		_w7503_
	);
	LUT2 #(
		.INIT('h1)
	) name5996 (
		\WX9910_reg/NET0131 ,
		\_2320__reg/NET0131 ,
		_w7504_
	);
	LUT2 #(
		.INIT('h8)
	) name5997 (
		\WX9910_reg/NET0131 ,
		\_2320__reg/NET0131 ,
		_w7505_
	);
	LUT2 #(
		.INIT('h1)
	) name5998 (
		_w7504_,
		_w7505_,
		_w7506_
	);
	LUT2 #(
		.INIT('h2)
	) name5999 (
		RESET_pad,
		_w7506_,
		_w7507_
	);
	LUT2 #(
		.INIT('h1)
	) name6000 (
		\WX9908_reg/NET0131 ,
		\_2321__reg/NET0131 ,
		_w7508_
	);
	LUT2 #(
		.INIT('h8)
	) name6001 (
		\WX9908_reg/NET0131 ,
		\_2321__reg/NET0131 ,
		_w7509_
	);
	LUT2 #(
		.INIT('h1)
	) name6002 (
		_w7508_,
		_w7509_,
		_w7510_
	);
	LUT2 #(
		.INIT('h2)
	) name6003 (
		RESET_pad,
		_w7510_,
		_w7511_
	);
	LUT2 #(
		.INIT('h1)
	) name6004 (
		\WX9906_reg/NET0131 ,
		\_2322__reg/NET0131 ,
		_w7512_
	);
	LUT2 #(
		.INIT('h8)
	) name6005 (
		\WX9906_reg/NET0131 ,
		\_2322__reg/NET0131 ,
		_w7513_
	);
	LUT2 #(
		.INIT('h1)
	) name6006 (
		_w7512_,
		_w7513_,
		_w7514_
	);
	LUT2 #(
		.INIT('h2)
	) name6007 (
		RESET_pad,
		_w7514_,
		_w7515_
	);
	LUT2 #(
		.INIT('h1)
	) name6008 (
		\WX9904_reg/NET0131 ,
		\_2323__reg/NET0131 ,
		_w7516_
	);
	LUT2 #(
		.INIT('h8)
	) name6009 (
		\WX9904_reg/NET0131 ,
		\_2323__reg/NET0131 ,
		_w7517_
	);
	LUT2 #(
		.INIT('h1)
	) name6010 (
		_w7516_,
		_w7517_,
		_w7518_
	);
	LUT2 #(
		.INIT('h2)
	) name6011 (
		RESET_pad,
		_w7518_,
		_w7519_
	);
	LUT2 #(
		.INIT('h1)
	) name6012 (
		\WX9902_reg/NET0131 ,
		\_2324__reg/NET0131 ,
		_w7520_
	);
	LUT2 #(
		.INIT('h8)
	) name6013 (
		\WX9902_reg/NET0131 ,
		\_2324__reg/NET0131 ,
		_w7521_
	);
	LUT2 #(
		.INIT('h1)
	) name6014 (
		_w7520_,
		_w7521_,
		_w7522_
	);
	LUT2 #(
		.INIT('h2)
	) name6015 (
		RESET_pad,
		_w7522_,
		_w7523_
	);
	LUT2 #(
		.INIT('h1)
	) name6016 (
		\WX9900_reg/NET0131 ,
		\_2325__reg/NET0131 ,
		_w7524_
	);
	LUT2 #(
		.INIT('h8)
	) name6017 (
		\WX9900_reg/NET0131 ,
		\_2325__reg/NET0131 ,
		_w7525_
	);
	LUT2 #(
		.INIT('h1)
	) name6018 (
		_w7524_,
		_w7525_,
		_w7526_
	);
	LUT2 #(
		.INIT('h2)
	) name6019 (
		RESET_pad,
		_w7526_,
		_w7527_
	);
	LUT2 #(
		.INIT('h1)
	) name6020 (
		\WX9898_reg/NET0131 ,
		\_2326__reg/NET0131 ,
		_w7528_
	);
	LUT2 #(
		.INIT('h8)
	) name6021 (
		\WX9898_reg/NET0131 ,
		\_2326__reg/NET0131 ,
		_w7529_
	);
	LUT2 #(
		.INIT('h1)
	) name6022 (
		_w7528_,
		_w7529_,
		_w7530_
	);
	LUT2 #(
		.INIT('h2)
	) name6023 (
		RESET_pad,
		_w7530_,
		_w7531_
	);
	LUT2 #(
		.INIT('h1)
	) name6024 (
		\WX9896_reg/NET0131 ,
		\_2327__reg/NET0131 ,
		_w7532_
	);
	LUT2 #(
		.INIT('h8)
	) name6025 (
		\WX9896_reg/NET0131 ,
		\_2327__reg/NET0131 ,
		_w7533_
	);
	LUT2 #(
		.INIT('h1)
	) name6026 (
		_w7532_,
		_w7533_,
		_w7534_
	);
	LUT2 #(
		.INIT('h2)
	) name6027 (
		RESET_pad,
		_w7534_,
		_w7535_
	);
	LUT2 #(
		.INIT('h1)
	) name6028 (
		\WX9894_reg/NET0131 ,
		\_2328__reg/NET0131 ,
		_w7536_
	);
	LUT2 #(
		.INIT('h8)
	) name6029 (
		\WX9894_reg/NET0131 ,
		\_2328__reg/NET0131 ,
		_w7537_
	);
	LUT2 #(
		.INIT('h1)
	) name6030 (
		_w7536_,
		_w7537_,
		_w7538_
	);
	LUT2 #(
		.INIT('h2)
	) name6031 (
		RESET_pad,
		_w7538_,
		_w7539_
	);
	LUT2 #(
		.INIT('h1)
	) name6032 (
		\WX9892_reg/NET0131 ,
		\_2329__reg/NET0131 ,
		_w7540_
	);
	LUT2 #(
		.INIT('h8)
	) name6033 (
		\WX9892_reg/NET0131 ,
		\_2329__reg/NET0131 ,
		_w7541_
	);
	LUT2 #(
		.INIT('h1)
	) name6034 (
		_w7540_,
		_w7541_,
		_w7542_
	);
	LUT2 #(
		.INIT('h2)
	) name6035 (
		RESET_pad,
		_w7542_,
		_w7543_
	);
	LUT2 #(
		.INIT('h1)
	) name6036 (
		\WX9888_reg/NET0131 ,
		\_2331__reg/NET0131 ,
		_w7544_
	);
	LUT2 #(
		.INIT('h8)
	) name6037 (
		\WX9888_reg/NET0131 ,
		\_2331__reg/NET0131 ,
		_w7545_
	);
	LUT2 #(
		.INIT('h1)
	) name6038 (
		_w7544_,
		_w7545_,
		_w7546_
	);
	LUT2 #(
		.INIT('h2)
	) name6039 (
		RESET_pad,
		_w7546_,
		_w7547_
	);
	LUT2 #(
		.INIT('h1)
	) name6040 (
		\WX11243_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w7548_
	);
	LUT2 #(
		.INIT('h8)
	) name6041 (
		\WX11243_reg/NET0131 ,
		\_2364__reg/NET0131 ,
		_w7549_
	);
	LUT2 #(
		.INIT('h1)
	) name6042 (
		_w7548_,
		_w7549_,
		_w7550_
	);
	LUT2 #(
		.INIT('h2)
	) name6043 (
		RESET_pad,
		_w7550_,
		_w7551_
	);
	LUT2 #(
		.INIT('h1)
	) name6044 (
		\WX11241_reg/NET0131 ,
		\_2333__reg/NET0131 ,
		_w7552_
	);
	LUT2 #(
		.INIT('h8)
	) name6045 (
		\WX11241_reg/NET0131 ,
		\_2333__reg/NET0131 ,
		_w7553_
	);
	LUT2 #(
		.INIT('h1)
	) name6046 (
		_w7552_,
		_w7553_,
		_w7554_
	);
	LUT2 #(
		.INIT('h2)
	) name6047 (
		RESET_pad,
		_w7554_,
		_w7555_
	);
	LUT2 #(
		.INIT('h1)
	) name6048 (
		\WX11239_reg/NET0131 ,
		\_2334__reg/NET0131 ,
		_w7556_
	);
	LUT2 #(
		.INIT('h8)
	) name6049 (
		\WX11239_reg/NET0131 ,
		\_2334__reg/NET0131 ,
		_w7557_
	);
	LUT2 #(
		.INIT('h1)
	) name6050 (
		_w7556_,
		_w7557_,
		_w7558_
	);
	LUT2 #(
		.INIT('h2)
	) name6051 (
		RESET_pad,
		_w7558_,
		_w7559_
	);
	LUT2 #(
		.INIT('h1)
	) name6052 (
		\WX11237_reg/NET0131 ,
		\_2335__reg/NET0131 ,
		_w7560_
	);
	LUT2 #(
		.INIT('h8)
	) name6053 (
		\WX11237_reg/NET0131 ,
		\_2335__reg/NET0131 ,
		_w7561_
	);
	LUT2 #(
		.INIT('h1)
	) name6054 (
		_w7560_,
		_w7561_,
		_w7562_
	);
	LUT2 #(
		.INIT('h2)
	) name6055 (
		RESET_pad,
		_w7562_,
		_w7563_
	);
	LUT2 #(
		.INIT('h1)
	) name6056 (
		\WX11233_reg/NET0131 ,
		\_2337__reg/NET0131 ,
		_w7564_
	);
	LUT2 #(
		.INIT('h8)
	) name6057 (
		\WX11233_reg/NET0131 ,
		\_2337__reg/NET0131 ,
		_w7565_
	);
	LUT2 #(
		.INIT('h1)
	) name6058 (
		_w7564_,
		_w7565_,
		_w7566_
	);
	LUT2 #(
		.INIT('h2)
	) name6059 (
		RESET_pad,
		_w7566_,
		_w7567_
	);
	LUT2 #(
		.INIT('h1)
	) name6060 (
		\WX11231_reg/NET0131 ,
		\_2338__reg/NET0131 ,
		_w7568_
	);
	LUT2 #(
		.INIT('h8)
	) name6061 (
		\WX11231_reg/NET0131 ,
		\_2338__reg/NET0131 ,
		_w7569_
	);
	LUT2 #(
		.INIT('h1)
	) name6062 (
		_w7568_,
		_w7569_,
		_w7570_
	);
	LUT2 #(
		.INIT('h2)
	) name6063 (
		RESET_pad,
		_w7570_,
		_w7571_
	);
	LUT2 #(
		.INIT('h1)
	) name6064 (
		\WX11229_reg/NET0131 ,
		\_2339__reg/NET0131 ,
		_w7572_
	);
	LUT2 #(
		.INIT('h8)
	) name6065 (
		\WX11229_reg/NET0131 ,
		\_2339__reg/NET0131 ,
		_w7573_
	);
	LUT2 #(
		.INIT('h1)
	) name6066 (
		_w7572_,
		_w7573_,
		_w7574_
	);
	LUT2 #(
		.INIT('h2)
	) name6067 (
		RESET_pad,
		_w7574_,
		_w7575_
	);
	LUT2 #(
		.INIT('h1)
	) name6068 (
		\WX11227_reg/NET0131 ,
		\_2340__reg/NET0131 ,
		_w7576_
	);
	LUT2 #(
		.INIT('h8)
	) name6069 (
		\WX11227_reg/NET0131 ,
		\_2340__reg/NET0131 ,
		_w7577_
	);
	LUT2 #(
		.INIT('h1)
	) name6070 (
		_w7576_,
		_w7577_,
		_w7578_
	);
	LUT2 #(
		.INIT('h2)
	) name6071 (
		RESET_pad,
		_w7578_,
		_w7579_
	);
	LUT2 #(
		.INIT('h1)
	) name6072 (
		\WX11225_reg/NET0131 ,
		\_2341__reg/NET0131 ,
		_w7580_
	);
	LUT2 #(
		.INIT('h8)
	) name6073 (
		\WX11225_reg/NET0131 ,
		\_2341__reg/NET0131 ,
		_w7581_
	);
	LUT2 #(
		.INIT('h1)
	) name6074 (
		_w7580_,
		_w7581_,
		_w7582_
	);
	LUT2 #(
		.INIT('h2)
	) name6075 (
		RESET_pad,
		_w7582_,
		_w7583_
	);
	LUT2 #(
		.INIT('h1)
	) name6076 (
		\WX11223_reg/NET0131 ,
		\_2342__reg/NET0131 ,
		_w7584_
	);
	LUT2 #(
		.INIT('h8)
	) name6077 (
		\WX11223_reg/NET0131 ,
		\_2342__reg/NET0131 ,
		_w7585_
	);
	LUT2 #(
		.INIT('h1)
	) name6078 (
		_w7584_,
		_w7585_,
		_w7586_
	);
	LUT2 #(
		.INIT('h2)
	) name6079 (
		RESET_pad,
		_w7586_,
		_w7587_
	);
	LUT2 #(
		.INIT('h1)
	) name6080 (
		\WX11219_reg/NET0131 ,
		\_2344__reg/NET0131 ,
		_w7588_
	);
	LUT2 #(
		.INIT('h8)
	) name6081 (
		\WX11219_reg/NET0131 ,
		\_2344__reg/NET0131 ,
		_w7589_
	);
	LUT2 #(
		.INIT('h1)
	) name6082 (
		_w7588_,
		_w7589_,
		_w7590_
	);
	LUT2 #(
		.INIT('h2)
	) name6083 (
		RESET_pad,
		_w7590_,
		_w7591_
	);
	LUT2 #(
		.INIT('h1)
	) name6084 (
		\WX11217_reg/NET0131 ,
		\_2345__reg/NET0131 ,
		_w7592_
	);
	LUT2 #(
		.INIT('h8)
	) name6085 (
		\WX11217_reg/NET0131 ,
		\_2345__reg/NET0131 ,
		_w7593_
	);
	LUT2 #(
		.INIT('h1)
	) name6086 (
		_w7592_,
		_w7593_,
		_w7594_
	);
	LUT2 #(
		.INIT('h2)
	) name6087 (
		RESET_pad,
		_w7594_,
		_w7595_
	);
	LUT2 #(
		.INIT('h1)
	) name6088 (
		\WX11213_reg/NET0131 ,
		\_2347__reg/NET0131 ,
		_w7596_
	);
	LUT2 #(
		.INIT('h8)
	) name6089 (
		\WX11213_reg/NET0131 ,
		\_2347__reg/NET0131 ,
		_w7597_
	);
	LUT2 #(
		.INIT('h1)
	) name6090 (
		_w7596_,
		_w7597_,
		_w7598_
	);
	LUT2 #(
		.INIT('h2)
	) name6091 (
		RESET_pad,
		_w7598_,
		_w7599_
	);
	LUT2 #(
		.INIT('h1)
	) name6092 (
		\WX11209_reg/NET0131 ,
		\_2349__reg/NET0131 ,
		_w7600_
	);
	LUT2 #(
		.INIT('h8)
	) name6093 (
		\WX11209_reg/NET0131 ,
		\_2349__reg/NET0131 ,
		_w7601_
	);
	LUT2 #(
		.INIT('h1)
	) name6094 (
		_w7600_,
		_w7601_,
		_w7602_
	);
	LUT2 #(
		.INIT('h2)
	) name6095 (
		RESET_pad,
		_w7602_,
		_w7603_
	);
	LUT2 #(
		.INIT('h1)
	) name6096 (
		\WX11207_reg/NET0131 ,
		\_2350__reg/NET0131 ,
		_w7604_
	);
	LUT2 #(
		.INIT('h8)
	) name6097 (
		\WX11207_reg/NET0131 ,
		\_2350__reg/NET0131 ,
		_w7605_
	);
	LUT2 #(
		.INIT('h1)
	) name6098 (
		_w7604_,
		_w7605_,
		_w7606_
	);
	LUT2 #(
		.INIT('h2)
	) name6099 (
		RESET_pad,
		_w7606_,
		_w7607_
	);
	LUT2 #(
		.INIT('h1)
	) name6100 (
		\WX11205_reg/NET0131 ,
		\_2351__reg/NET0131 ,
		_w7608_
	);
	LUT2 #(
		.INIT('h8)
	) name6101 (
		\WX11205_reg/NET0131 ,
		\_2351__reg/NET0131 ,
		_w7609_
	);
	LUT2 #(
		.INIT('h1)
	) name6102 (
		_w7608_,
		_w7609_,
		_w7610_
	);
	LUT2 #(
		.INIT('h2)
	) name6103 (
		RESET_pad,
		_w7610_,
		_w7611_
	);
	LUT2 #(
		.INIT('h1)
	) name6104 (
		\WX11203_reg/NET0131 ,
		\_2352__reg/NET0131 ,
		_w7612_
	);
	LUT2 #(
		.INIT('h8)
	) name6105 (
		\WX11203_reg/NET0131 ,
		\_2352__reg/NET0131 ,
		_w7613_
	);
	LUT2 #(
		.INIT('h1)
	) name6106 (
		_w7612_,
		_w7613_,
		_w7614_
	);
	LUT2 #(
		.INIT('h2)
	) name6107 (
		RESET_pad,
		_w7614_,
		_w7615_
	);
	LUT2 #(
		.INIT('h1)
	) name6108 (
		\WX11201_reg/NET0131 ,
		\_2353__reg/NET0131 ,
		_w7616_
	);
	LUT2 #(
		.INIT('h8)
	) name6109 (
		\WX11201_reg/NET0131 ,
		\_2353__reg/NET0131 ,
		_w7617_
	);
	LUT2 #(
		.INIT('h1)
	) name6110 (
		_w7616_,
		_w7617_,
		_w7618_
	);
	LUT2 #(
		.INIT('h2)
	) name6111 (
		RESET_pad,
		_w7618_,
		_w7619_
	);
	LUT2 #(
		.INIT('h1)
	) name6112 (
		\WX11199_reg/NET0131 ,
		\_2354__reg/NET0131 ,
		_w7620_
	);
	LUT2 #(
		.INIT('h8)
	) name6113 (
		\WX11199_reg/NET0131 ,
		\_2354__reg/NET0131 ,
		_w7621_
	);
	LUT2 #(
		.INIT('h1)
	) name6114 (
		_w7620_,
		_w7621_,
		_w7622_
	);
	LUT2 #(
		.INIT('h2)
	) name6115 (
		RESET_pad,
		_w7622_,
		_w7623_
	);
	LUT2 #(
		.INIT('h1)
	) name6116 (
		\WX11197_reg/NET0131 ,
		\_2355__reg/NET0131 ,
		_w7624_
	);
	LUT2 #(
		.INIT('h8)
	) name6117 (
		\WX11197_reg/NET0131 ,
		\_2355__reg/NET0131 ,
		_w7625_
	);
	LUT2 #(
		.INIT('h1)
	) name6118 (
		_w7624_,
		_w7625_,
		_w7626_
	);
	LUT2 #(
		.INIT('h2)
	) name6119 (
		RESET_pad,
		_w7626_,
		_w7627_
	);
	LUT2 #(
		.INIT('h1)
	) name6120 (
		\WX11195_reg/NET0131 ,
		\_2356__reg/NET0131 ,
		_w7628_
	);
	LUT2 #(
		.INIT('h8)
	) name6121 (
		\WX11195_reg/NET0131 ,
		\_2356__reg/NET0131 ,
		_w7629_
	);
	LUT2 #(
		.INIT('h1)
	) name6122 (
		_w7628_,
		_w7629_,
		_w7630_
	);
	LUT2 #(
		.INIT('h2)
	) name6123 (
		RESET_pad,
		_w7630_,
		_w7631_
	);
	LUT2 #(
		.INIT('h1)
	) name6124 (
		\WX11193_reg/NET0131 ,
		\_2357__reg/NET0131 ,
		_w7632_
	);
	LUT2 #(
		.INIT('h8)
	) name6125 (
		\WX11193_reg/NET0131 ,
		\_2357__reg/NET0131 ,
		_w7633_
	);
	LUT2 #(
		.INIT('h1)
	) name6126 (
		_w7632_,
		_w7633_,
		_w7634_
	);
	LUT2 #(
		.INIT('h2)
	) name6127 (
		RESET_pad,
		_w7634_,
		_w7635_
	);
	LUT2 #(
		.INIT('h1)
	) name6128 (
		\WX11191_reg/NET0131 ,
		\_2358__reg/NET0131 ,
		_w7636_
	);
	LUT2 #(
		.INIT('h8)
	) name6129 (
		\WX11191_reg/NET0131 ,
		\_2358__reg/NET0131 ,
		_w7637_
	);
	LUT2 #(
		.INIT('h1)
	) name6130 (
		_w7636_,
		_w7637_,
		_w7638_
	);
	LUT2 #(
		.INIT('h2)
	) name6131 (
		RESET_pad,
		_w7638_,
		_w7639_
	);
	LUT2 #(
		.INIT('h1)
	) name6132 (
		\WX11189_reg/NET0131 ,
		\_2359__reg/NET0131 ,
		_w7640_
	);
	LUT2 #(
		.INIT('h8)
	) name6133 (
		\WX11189_reg/NET0131 ,
		\_2359__reg/NET0131 ,
		_w7641_
	);
	LUT2 #(
		.INIT('h1)
	) name6134 (
		_w7640_,
		_w7641_,
		_w7642_
	);
	LUT2 #(
		.INIT('h2)
	) name6135 (
		RESET_pad,
		_w7642_,
		_w7643_
	);
	LUT2 #(
		.INIT('h1)
	) name6136 (
		\WX11187_reg/NET0131 ,
		\_2360__reg/NET0131 ,
		_w7644_
	);
	LUT2 #(
		.INIT('h8)
	) name6137 (
		\WX11187_reg/NET0131 ,
		\_2360__reg/NET0131 ,
		_w7645_
	);
	LUT2 #(
		.INIT('h1)
	) name6138 (
		_w7644_,
		_w7645_,
		_w7646_
	);
	LUT2 #(
		.INIT('h2)
	) name6139 (
		RESET_pad,
		_w7646_,
		_w7647_
	);
	LUT2 #(
		.INIT('h1)
	) name6140 (
		\WX11183_reg/NET0131 ,
		\_2362__reg/NET0131 ,
		_w7648_
	);
	LUT2 #(
		.INIT('h8)
	) name6141 (
		\WX11183_reg/NET0131 ,
		\_2362__reg/NET0131 ,
		_w7649_
	);
	LUT2 #(
		.INIT('h1)
	) name6142 (
		_w7648_,
		_w7649_,
		_w7650_
	);
	LUT2 #(
		.INIT('h2)
	) name6143 (
		RESET_pad,
		_w7650_,
		_w7651_
	);
	LUT2 #(
		.INIT('h1)
	) name6144 (
		\WX2150_reg/NET0131 ,
		\_2129__reg/NET0131 ,
		_w7652_
	);
	LUT2 #(
		.INIT('h8)
	) name6145 (
		\WX2150_reg/NET0131 ,
		\_2129__reg/NET0131 ,
		_w7653_
	);
	LUT2 #(
		.INIT('h1)
	) name6146 (
		_w7652_,
		_w7653_,
		_w7654_
	);
	LUT2 #(
		.INIT('h2)
	) name6147 (
		RESET_pad,
		_w7654_,
		_w7655_
	);
	LUT2 #(
		.INIT('h1)
	) name6148 (
		\WX7304_reg/NET0131 ,
		\_2266__reg/NET0131 ,
		_w7656_
	);
	LUT2 #(
		.INIT('h8)
	) name6149 (
		\WX7304_reg/NET0131 ,
		\_2266__reg/NET0131 ,
		_w7657_
	);
	LUT2 #(
		.INIT('h1)
	) name6150 (
		_w7656_,
		_w7657_,
		_w7658_
	);
	LUT2 #(
		.INIT('h2)
	) name6151 (
		RESET_pad,
		_w7658_,
		_w7659_
	);
	LUT2 #(
		.INIT('h1)
	) name6152 (
		\WX2136_reg/NET0131 ,
		\_2136__reg/NET0131 ,
		_w7660_
	);
	LUT2 #(
		.INIT('h8)
	) name6153 (
		\WX2136_reg/NET0131 ,
		\_2136__reg/NET0131 ,
		_w7661_
	);
	LUT2 #(
		.INIT('h1)
	) name6154 (
		_w7660_,
		_w7661_,
		_w7662_
	);
	LUT2 #(
		.INIT('h2)
	) name6155 (
		RESET_pad,
		_w7662_,
		_w7663_
	);
	LUT2 #(
		.INIT('h1)
	) name6156 (
		\WX3467_reg/NET0131 ,
		\_2149__reg/NET0131 ,
		_w7664_
	);
	LUT2 #(
		.INIT('h8)
	) name6157 (
		\WX3467_reg/NET0131 ,
		\_2149__reg/NET0131 ,
		_w7665_
	);
	LUT2 #(
		.INIT('h1)
	) name6158 (
		_w7664_,
		_w7665_,
		_w7666_
	);
	LUT2 #(
		.INIT('h2)
	) name6159 (
		RESET_pad,
		_w7666_,
		_w7667_
	);
	LUT2 #(
		.INIT('h1)
	) name6160 (
		\WX8633_reg/NET0131 ,
		\_2280__reg/NET0131 ,
		_w7668_
	);
	LUT2 #(
		.INIT('h8)
	) name6161 (
		\WX8633_reg/NET0131 ,
		\_2280__reg/NET0131 ,
		_w7669_
	);
	LUT2 #(
		.INIT('h1)
	) name6162 (
		_w7668_,
		_w7669_,
		_w7670_
	);
	LUT2 #(
		.INIT('h2)
	) name6163 (
		RESET_pad,
		_w7670_,
		_w7671_
	);
	LUT2 #(
		.INIT('h1)
	) name6164 (
		\WX853_reg/NET0131 ,
		\_2099__reg/NET0131 ,
		_w7672_
	);
	LUT2 #(
		.INIT('h8)
	) name6165 (
		\WX853_reg/NET0131 ,
		\_2099__reg/NET0131 ,
		_w7673_
	);
	LUT2 #(
		.INIT('h1)
	) name6166 (
		_w7672_,
		_w7673_,
		_w7674_
	);
	LUT2 #(
		.INIT('h2)
	) name6167 (
		RESET_pad,
		_w7674_,
		_w7675_
	);
	LUT2 #(
		.INIT('h1)
	) name6168 (
		\WX859_reg/NET0131 ,
		\_2096__reg/NET0131 ,
		_w7676_
	);
	LUT2 #(
		.INIT('h8)
	) name6169 (
		\WX859_reg/NET0131 ,
		\_2096__reg/NET0131 ,
		_w7677_
	);
	LUT2 #(
		.INIT('h1)
	) name6170 (
		_w7676_,
		_w7677_,
		_w7678_
	);
	LUT2 #(
		.INIT('h2)
	) name6171 (
		RESET_pad,
		_w7678_,
		_w7679_
	);
	LUT2 #(
		.INIT('h1)
	) name6172 (
		\WX7310_reg/NET0131 ,
		\_2263__reg/NET0131 ,
		_w7680_
	);
	LUT2 #(
		.INIT('h8)
	) name6173 (
		\WX7310_reg/NET0131 ,
		\_2263__reg/NET0131 ,
		_w7681_
	);
	LUT2 #(
		.INIT('h1)
	) name6174 (
		_w7680_,
		_w7681_,
		_w7682_
	);
	LUT2 #(
		.INIT('h2)
	) name6175 (
		RESET_pad,
		_w7682_,
		_w7683_
	);
	LUT2 #(
		.INIT('h1)
	) name6176 (
		\WX9936_reg/NET0131 ,
		\_2307__reg/NET0131 ,
		_w7684_
	);
	LUT2 #(
		.INIT('h8)
	) name6177 (
		\WX9936_reg/NET0131 ,
		\_2307__reg/NET0131 ,
		_w7685_
	);
	LUT2 #(
		.INIT('h1)
	) name6178 (
		_w7684_,
		_w7685_,
		_w7686_
	);
	LUT2 #(
		.INIT('h2)
	) name6179 (
		RESET_pad,
		_w7686_,
		_w7687_
	);
	LUT2 #(
		.INIT('h1)
	) name6180 (
		\WX849_reg/NET0131 ,
		\_2101__reg/NET0131 ,
		_w7688_
	);
	LUT2 #(
		.INIT('h8)
	) name6181 (
		\WX849_reg/NET0131 ,
		\_2101__reg/NET0131 ,
		_w7689_
	);
	LUT2 #(
		.INIT('h1)
	) name6182 (
		_w7688_,
		_w7689_,
		_w7690_
	);
	LUT2 #(
		.INIT('h2)
	) name6183 (
		RESET_pad,
		_w7690_,
		_w7691_
	);
	LUT2 #(
		.INIT('h1)
	) name6184 (
		\WX2140_reg/NET0131 ,
		\_2134__reg/NET0131 ,
		_w7692_
	);
	LUT2 #(
		.INIT('h8)
	) name6185 (
		\WX2140_reg/NET0131 ,
		\_2134__reg/NET0131 ,
		_w7693_
	);
	LUT2 #(
		.INIT('h1)
	) name6186 (
		_w7692_,
		_w7693_,
		_w7694_
	);
	LUT2 #(
		.INIT('h2)
	) name6187 (
		RESET_pad,
		_w7694_,
		_w7695_
	);
	LUT2 #(
		.INIT('h1)
	) name6188 (
		\WX2178_reg/NET0131 ,
		\_2115__reg/NET0131 ,
		_w7696_
	);
	LUT2 #(
		.INIT('h8)
	) name6189 (
		\WX2178_reg/NET0131 ,
		\_2115__reg/NET0131 ,
		_w7697_
	);
	LUT2 #(
		.INIT('h1)
	) name6190 (
		_w7696_,
		_w7697_,
		_w7698_
	);
	LUT2 #(
		.INIT('h2)
	) name6191 (
		RESET_pad,
		_w7698_,
		_w7699_
	);
	LUT2 #(
		.INIT('h1)
	) name6192 (
		\WX8623_reg/NET0131 ,
		\_2285__reg/NET0131 ,
		_w7700_
	);
	LUT2 #(
		.INIT('h8)
	) name6193 (
		\WX8623_reg/NET0131 ,
		\_2285__reg/NET0131 ,
		_w7701_
	);
	LUT2 #(
		.INIT('h1)
	) name6194 (
		_w7700_,
		_w7701_,
		_w7702_
	);
	LUT2 #(
		.INIT('h2)
	) name6195 (
		RESET_pad,
		_w7702_,
		_w7703_
	);
	LUT2 #(
		.INIT('h1)
	) name6196 (
		\WX2176_reg/NET0131 ,
		\_2116__reg/NET0131 ,
		_w7704_
	);
	LUT2 #(
		.INIT('h8)
	) name6197 (
		\WX2176_reg/NET0131 ,
		\_2116__reg/NET0131 ,
		_w7705_
	);
	LUT2 #(
		.INIT('h1)
	) name6198 (
		_w7704_,
		_w7705_,
		_w7706_
	);
	LUT2 #(
		.INIT('h2)
	) name6199 (
		RESET_pad,
		_w7706_,
		_w7707_
	);
	LUT2 #(
		.INIT('h1)
	) name6200 (
		\WX7346_reg/NET0131 ,
		\_2245__reg/NET0131 ,
		_w7708_
	);
	LUT2 #(
		.INIT('h8)
	) name6201 (
		\WX7346_reg/NET0131 ,
		\_2245__reg/NET0131 ,
		_w7709_
	);
	LUT2 #(
		.INIT('h1)
	) name6202 (
		_w7708_,
		_w7709_,
		_w7710_
	);
	LUT2 #(
		.INIT('h2)
	) name6203 (
		RESET_pad,
		_w7710_,
		_w7711_
	);
	LUT2 #(
		.INIT('h1)
	) name6204 (
		\WX6041_reg/NET0131 ,
		\_2219__reg/NET0131 ,
		_w7712_
	);
	LUT2 #(
		.INIT('h8)
	) name6205 (
		\WX6041_reg/NET0131 ,
		\_2219__reg/NET0131 ,
		_w7713_
	);
	LUT2 #(
		.INIT('h1)
	) name6206 (
		_w7712_,
		_w7713_,
		_w7714_
	);
	LUT2 #(
		.INIT('h2)
	) name6207 (
		RESET_pad,
		_w7714_,
		_w7715_
	);
	LUT2 #(
		.INIT('h1)
	) name6208 (
		\WX7350_reg/NET0131 ,
		\_2243__reg/NET0131 ,
		_w7716_
	);
	LUT2 #(
		.INIT('h8)
	) name6209 (
		\WX7350_reg/NET0131 ,
		\_2243__reg/NET0131 ,
		_w7717_
	);
	LUT2 #(
		.INIT('h1)
	) name6210 (
		_w7716_,
		_w7717_,
		_w7718_
	);
	LUT2 #(
		.INIT('h2)
	) name6211 (
		RESET_pad,
		_w7718_,
		_w7719_
	);
	LUT2 #(
		.INIT('h1)
	) name6212 (
		\WX4762_reg/NET0131 ,
		\_2180__reg/NET0131 ,
		_w7720_
	);
	LUT2 #(
		.INIT('h8)
	) name6213 (
		\WX4762_reg/NET0131 ,
		\_2180__reg/NET0131 ,
		_w7721_
	);
	LUT2 #(
		.INIT('h1)
	) name6214 (
		_w7720_,
		_w7721_,
		_w7722_
	);
	LUT2 #(
		.INIT('h2)
	) name6215 (
		RESET_pad,
		_w7722_,
		_w7723_
	);
	LUT2 #(
		.INIT('h1)
	) name6216 (
		\WX871_reg/NET0131 ,
		\_2090__reg/NET0131 ,
		_w7724_
	);
	LUT2 #(
		.INIT('h8)
	) name6217 (
		\WX871_reg/NET0131 ,
		\_2090__reg/NET0131 ,
		_w7725_
	);
	LUT2 #(
		.INIT('h1)
	) name6218 (
		_w7724_,
		_w7725_,
		_w7726_
	);
	LUT2 #(
		.INIT('h2)
	) name6219 (
		RESET_pad,
		_w7726_,
		_w7727_
	);
	LUT2 #(
		.INIT('h1)
	) name6220 (
		\WX885_reg/NET0131 ,
		\_2083__reg/NET0131 ,
		_w7728_
	);
	LUT2 #(
		.INIT('h8)
	) name6221 (
		\WX885_reg/NET0131 ,
		\_2083__reg/NET0131 ,
		_w7729_
	);
	LUT2 #(
		.INIT('h1)
	) name6222 (
		_w7728_,
		_w7729_,
		_w7730_
	);
	LUT2 #(
		.INIT('h2)
	) name6223 (
		RESET_pad,
		_w7730_,
		_w7731_
	);
	LUT2 #(
		.INIT('h1)
	) name6224 (
		\WX11185_reg/NET0131 ,
		\_2361__reg/NET0131 ,
		_w7732_
	);
	LUT2 #(
		.INIT('h8)
	) name6225 (
		\WX11185_reg/NET0131 ,
		\_2361__reg/NET0131 ,
		_w7733_
	);
	LUT2 #(
		.INIT('h1)
	) name6226 (
		_w7732_,
		_w7733_,
		_w7734_
	);
	LUT2 #(
		.INIT('h2)
	) name6227 (
		RESET_pad,
		_w7734_,
		_w7735_
	);
	LUT2 #(
		.INIT('h1)
	) name6228 (
		\WX9890_reg/NET0131 ,
		\_2330__reg/NET0131 ,
		_w7736_
	);
	LUT2 #(
		.INIT('h8)
	) name6229 (
		\WX9890_reg/NET0131 ,
		\_2330__reg/NET0131 ,
		_w7737_
	);
	LUT2 #(
		.INIT('h1)
	) name6230 (
		_w7736_,
		_w7737_,
		_w7738_
	);
	LUT2 #(
		.INIT('h2)
	) name6231 (
		RESET_pad,
		_w7738_,
		_w7739_
	);
	LUT2 #(
		.INIT('h1)
	) name6232 (
		\WX9944_reg/NET0131 ,
		\_2303__reg/NET0131 ,
		_w7740_
	);
	LUT2 #(
		.INIT('h8)
	) name6233 (
		\WX9944_reg/NET0131 ,
		\_2303__reg/NET0131 ,
		_w7741_
	);
	LUT2 #(
		.INIT('h1)
	) name6234 (
		_w7740_,
		_w7741_,
		_w7742_
	);
	LUT2 #(
		.INIT('h2)
	) name6235 (
		RESET_pad,
		_w7742_,
		_w7743_
	);
	LUT2 #(
		.INIT('h1)
	) name6236 (
		\WX7344_reg/NET0131 ,
		\_2246__reg/NET0131 ,
		_w7744_
	);
	LUT2 #(
		.INIT('h8)
	) name6237 (
		\WX7344_reg/NET0131 ,
		\_2246__reg/NET0131 ,
		_w7745_
	);
	LUT2 #(
		.INIT('h1)
	) name6238 (
		_w7744_,
		_w7745_,
		_w7746_
	);
	LUT2 #(
		.INIT('h2)
	) name6239 (
		RESET_pad,
		_w7746_,
		_w7747_
	);
	LUT2 #(
		.INIT('h1)
	) name6240 (
		\WX7324_reg/NET0131 ,
		\_2256__reg/NET0131 ,
		_w7748_
	);
	LUT2 #(
		.INIT('h8)
	) name6241 (
		\WX7324_reg/NET0131 ,
		\_2256__reg/NET0131 ,
		_w7749_
	);
	LUT2 #(
		.INIT('h1)
	) name6242 (
		_w7748_,
		_w7749_,
		_w7750_
	);
	LUT2 #(
		.INIT('h2)
	) name6243 (
		RESET_pad,
		_w7750_,
		_w7751_
	);
	LUT2 #(
		.INIT('h1)
	) name6244 (
		\WX6013_reg/NET0131 ,
		\_2233__reg/NET0131 ,
		_w7752_
	);
	LUT2 #(
		.INIT('h8)
	) name6245 (
		\WX6013_reg/NET0131 ,
		\_2233__reg/NET0131 ,
		_w7753_
	);
	LUT2 #(
		.INIT('h1)
	) name6246 (
		_w7752_,
		_w7753_,
		_w7754_
	);
	LUT2 #(
		.INIT('h2)
	) name6247 (
		RESET_pad,
		_w7754_,
		_w7755_
	);
	LUT2 #(
		.INIT('h1)
	) name6248 (
		\WX2152_reg/NET0131 ,
		\_2128__reg/NET0131 ,
		_w7756_
	);
	LUT2 #(
		.INIT('h8)
	) name6249 (
		\WX2152_reg/NET0131 ,
		\_2128__reg/NET0131 ,
		_w7757_
	);
	LUT2 #(
		.INIT('h1)
	) name6250 (
		_w7756_,
		_w7757_,
		_w7758_
	);
	LUT2 #(
		.INIT('h2)
	) name6251 (
		RESET_pad,
		_w7758_,
		_w7759_
	);
	LUT2 #(
		.INIT('h1)
	) name6252 (
		\WX847_reg/NET0131 ,
		\_2102__reg/NET0131 ,
		_w7760_
	);
	LUT2 #(
		.INIT('h8)
	) name6253 (
		\WX847_reg/NET0131 ,
		\_2102__reg/NET0131 ,
		_w7761_
	);
	LUT2 #(
		.INIT('h1)
	) name6254 (
		_w7760_,
		_w7761_,
		_w7762_
	);
	LUT2 #(
		.INIT('h2)
	) name6255 (
		RESET_pad,
		_w7762_,
		_w7763_
	);
	LUT2 #(
		.INIT('h1)
	) name6256 (
		\WX3447_reg/NET0131 ,
		\_2159__reg/NET0131 ,
		_w7764_
	);
	LUT2 #(
		.INIT('h8)
	) name6257 (
		\WX3447_reg/NET0131 ,
		\_2159__reg/NET0131 ,
		_w7765_
	);
	LUT2 #(
		.INIT('h1)
	) name6258 (
		_w7764_,
		_w7765_,
		_w7766_
	);
	LUT2 #(
		.INIT('h2)
	) name6259 (
		RESET_pad,
		_w7766_,
		_w7767_
	);
	LUT2 #(
		.INIT('h1)
	) name6260 (
		\WX9924_reg/NET0131 ,
		\_2313__reg/NET0131 ,
		_w7768_
	);
	LUT2 #(
		.INIT('h8)
	) name6261 (
		\WX9924_reg/NET0131 ,
		\_2313__reg/NET0131 ,
		_w7769_
	);
	LUT2 #(
		.INIT('h1)
	) name6262 (
		_w7768_,
		_w7769_,
		_w7770_
	);
	LUT2 #(
		.INIT('h2)
	) name6263 (
		RESET_pad,
		_w7770_,
		_w7771_
	);
	LUT2 #(
		.INIT('h1)
	) name6264 (
		\WX861_reg/NET0131 ,
		\_2095__reg/NET0131 ,
		_w7772_
	);
	LUT2 #(
		.INIT('h8)
	) name6265 (
		\WX861_reg/NET0131 ,
		\_2095__reg/NET0131 ,
		_w7773_
	);
	LUT2 #(
		.INIT('h1)
	) name6266 (
		_w7772_,
		_w7773_,
		_w7774_
	);
	LUT2 #(
		.INIT('h2)
	) name6267 (
		RESET_pad,
		_w7774_,
		_w7775_
	);
	LUT2 #(
		.INIT('h1)
	) name6268 (
		\WX8639_reg/NET0131 ,
		\_2277__reg/NET0131 ,
		_w7776_
	);
	LUT2 #(
		.INIT('h8)
	) name6269 (
		\WX8639_reg/NET0131 ,
		\_2277__reg/NET0131 ,
		_w7777_
	);
	LUT2 #(
		.INIT('h1)
	) name6270 (
		_w7776_,
		_w7777_,
		_w7778_
	);
	LUT2 #(
		.INIT('h2)
	) name6271 (
		RESET_pad,
		_w7778_,
		_w7779_
	);
	LUT2 #(
		.INIT('h1)
	) name6272 (
		\WX7308_reg/NET0131 ,
		\_2264__reg/NET0131 ,
		_w7780_
	);
	LUT2 #(
		.INIT('h8)
	) name6273 (
		\WX7308_reg/NET0131 ,
		\_2264__reg/NET0131 ,
		_w7781_
	);
	LUT2 #(
		.INIT('h1)
	) name6274 (
		_w7780_,
		_w7781_,
		_w7782_
	);
	LUT2 #(
		.INIT('h2)
	) name6275 (
		RESET_pad,
		_w7782_,
		_w7783_
	);
	LUT2 #(
		.INIT('h1)
	) name6276 (
		\WX879_reg/NET0131 ,
		\_2086__reg/NET0131 ,
		_w7784_
	);
	LUT2 #(
		.INIT('h8)
	) name6277 (
		\WX879_reg/NET0131 ,
		\_2086__reg/NET0131 ,
		_w7785_
	);
	LUT2 #(
		.INIT('h1)
	) name6278 (
		_w7784_,
		_w7785_,
		_w7786_
	);
	LUT2 #(
		.INIT('h2)
	) name6279 (
		RESET_pad,
		_w7786_,
		_w7787_
	);
	LUT2 #(
		.INIT('h1)
	) name6280 (
		\WX7334_reg/NET0131 ,
		\_2251__reg/NET0131 ,
		_w7788_
	);
	LUT2 #(
		.INIT('h8)
	) name6281 (
		\WX7334_reg/NET0131 ,
		\_2251__reg/NET0131 ,
		_w7789_
	);
	LUT2 #(
		.INIT('h1)
	) name6282 (
		_w7788_,
		_w7789_,
		_w7790_
	);
	LUT2 #(
		.INIT('h2)
	) name6283 (
		RESET_pad,
		_w7790_,
		_w7791_
	);
	LUT2 #(
		.INIT('h1)
	) name6284 (
		\WX8643_reg/NET0131 ,
		\_2275__reg/NET0131 ,
		_w7792_
	);
	LUT2 #(
		.INIT('h8)
	) name6285 (
		\WX8643_reg/NET0131 ,
		\_2275__reg/NET0131 ,
		_w7793_
	);
	LUT2 #(
		.INIT('h1)
	) name6286 (
		_w7792_,
		_w7793_,
		_w7794_
	);
	LUT2 #(
		.INIT('h2)
	) name6287 (
		RESET_pad,
		_w7794_,
		_w7795_
	);
	LUT2 #(
		.INIT('h1)
	) name6288 (
		\WX4726_reg/NET0131 ,
		\_2198__reg/NET0131 ,
		_w7796_
	);
	LUT2 #(
		.INIT('h8)
	) name6289 (
		\WX4726_reg/NET0131 ,
		\_2198__reg/NET0131 ,
		_w7797_
	);
	LUT2 #(
		.INIT('h1)
	) name6290 (
		_w7796_,
		_w7797_,
		_w7798_
	);
	LUT2 #(
		.INIT('h2)
	) name6291 (
		RESET_pad,
		_w7798_,
		_w7799_
	);
	LUT2 #(
		.INIT('h8)
	) name6292 (
		RESET_pad,
		\WX11053_reg/NET0131 ,
		_w7800_
	);
	LUT2 #(
		.INIT('h8)
	) name6293 (
		RESET_pad,
		\WX709_reg/NET0131 ,
		_w7801_
	);
	LUT2 #(
		.INIT('h8)
	) name6294 (
		RESET_pad,
		\WX10891_reg/NET0131 ,
		_w7802_
	);
	LUT2 #(
		.INIT('h8)
	) name6295 (
		RESET_pad,
		\WX2002_reg/NET0131 ,
		_w7803_
	);
	LUT2 #(
		.INIT('h2)
	) name6296 (
		RESET_pad,
		\WX10829_reg/NET0131 ,
		_w7804_
	);
	LUT2 #(
		.INIT('h8)
	) name6297 (
		RESET_pad,
		\WX11059_reg/NET0131 ,
		_w7805_
	);
	LUT2 #(
		.INIT('h8)
	) name6298 (
		RESET_pad,
		\WX3271_reg/NET0131 ,
		_w7806_
	);
	LUT2 #(
		.INIT('h8)
	) name6299 (
		RESET_pad,
		\WX11033_reg/NET0131 ,
		_w7807_
	);
	LUT2 #(
		.INIT('h8)
	) name6300 (
		RESET_pad,
		\WX7252_reg/NET0131 ,
		_w7808_
	);
	LUT2 #(
		.INIT('h8)
	) name6301 (
		RESET_pad,
		\WX3257_reg/NET0131 ,
		_w7809_
	);
	LUT2 #(
		.INIT('h8)
	) name6302 (
		RESET_pad,
		\WX3403_reg/NET0131 ,
		_w7810_
	);
	LUT2 #(
		.INIT('h8)
	) name6303 (
		RESET_pad,
		\WX11115_reg/NET0131 ,
		_w7811_
	);
	LUT2 #(
		.INIT('h8)
	) name6304 (
		RESET_pad,
		\WX11049_reg/NET0131 ,
		_w7812_
	);
	LUT2 #(
		.INIT('h8)
	) name6305 (
		RESET_pad,
		\WX9714_reg/NET0131 ,
		_w7813_
	);
	LUT2 #(
		.INIT('h8)
	) name6306 (
		RESET_pad,
		\WX2004_reg/NET0131 ,
		_w7814_
	);
	LUT2 #(
		.INIT('h8)
	) name6307 (
		RESET_pad,
		\WX11037_reg/NET0131 ,
		_w7815_
	);
	LUT2 #(
		.INIT('h8)
	) name6308 (
		RESET_pad,
		\WX9852_reg/NET0131 ,
		_w7816_
	);
	LUT2 #(
		.INIT('h8)
	) name6309 (
		RESET_pad,
		\WX9702_reg/NET0131 ,
		_w7817_
	);
	LUT2 #(
		.INIT('h8)
	) name6310 (
		RESET_pad,
		\WX9876_reg/NET0131 ,
		_w7818_
	);
	LUT2 #(
		.INIT('h8)
	) name6311 (
		RESET_pad,
		\WX11121_reg/NET0131 ,
		_w7819_
	);
	LUT2 #(
		.INIT('h8)
	) name6312 (
		RESET_pad,
		\WX7114_reg/NET0131 ,
		_w7820_
	);
	LUT2 #(
		.INIT('h8)
	) name6313 (
		RESET_pad,
		\WX1986_reg/NET0131 ,
		_w7821_
	);
	LUT2 #(
		.INIT('h8)
	) name6314 (
		RESET_pad,
		\WX9802_reg/NET0131 ,
		_w7822_
	);
	LUT2 #(
		.INIT('h8)
	) name6315 (
		RESET_pad,
		\WX9824_reg/NET0131 ,
		_w7823_
	);
	LUT2 #(
		.INIT('h8)
	) name6316 (
		RESET_pad,
		\WX7220_reg/NET0131 ,
		_w7824_
	);
	LUT2 #(
		.INIT('h8)
	) name6317 (
		RESET_pad,
		\WX9806_reg/NET0131 ,
		_w7825_
	);
	LUT2 #(
		.INIT('h8)
	) name6318 (
		RESET_pad,
		\WX11073_reg/NET0131 ,
		_w7826_
	);
	LUT2 #(
		.INIT('h8)
	) name6319 (
		RESET_pad,
		\WX9878_reg/NET0131 ,
		_w7827_
	);
	LUT2 #(
		.INIT('h8)
	) name6320 (
		RESET_pad,
		\WX11111_reg/NET0131 ,
		_w7828_
	);
	LUT2 #(
		.INIT('h8)
	) name6321 (
		RESET_pad,
		\WX11169_reg/NET0131 ,
		_w7829_
	);
	LUT2 #(
		.INIT('h8)
	) name6322 (
		RESET_pad,
		\WX1998_reg/NET0131 ,
		_w7830_
	);
	LUT2 #(
		.INIT('h8)
	) name6323 (
		RESET_pad,
		\WX9850_reg/NET0131 ,
		_w7831_
	);
	LUT2 #(
		.INIT('h8)
	) name6324 (
		RESET_pad,
		\WX11079_reg/NET0131 ,
		_w7832_
	);
	LUT2 #(
		.INIT('h8)
	) name6325 (
		RESET_pad,
		\WX7110_reg/NET0131 ,
		_w7833_
	);
	LUT2 #(
		.INIT('h8)
	) name6326 (
		RESET_pad,
		\WX7240_reg/NET0131 ,
		_w7834_
	);
	LUT2 #(
		.INIT('h8)
	) name6327 (
		RESET_pad,
		\WX1954_reg/NET0131 ,
		_w7835_
	);
	LUT2 #(
		.INIT('h8)
	) name6328 (
		RESET_pad,
		\WX11081_reg/NET0131 ,
		_w7836_
	);
	LUT2 #(
		.INIT('h8)
	) name6329 (
		RESET_pad,
		\WX11083_reg/NET0131 ,
		_w7837_
	);
	LUT2 #(
		.INIT('h8)
	) name6330 (
		RESET_pad,
		\WX3339_reg/NET0131 ,
		_w7838_
	);
	LUT2 #(
		.INIT('h8)
	) name6331 (
		RESET_pad,
		\WX8491_reg/NET0131 ,
		_w7839_
	);
	LUT2 #(
		.INIT('h8)
	) name6332 (
		RESET_pad,
		\WX11175_reg/NET0131 ,
		_w7840_
	);
	LUT2 #(
		.INIT('h8)
	) name6333 (
		RESET_pad,
		\WX11089_reg/NET0131 ,
		_w7841_
	);
	LUT2 #(
		.INIT('h8)
	) name6334 (
		RESET_pad,
		\WX9770_reg/NET0131 ,
		_w7842_
	);
	LUT2 #(
		.INIT('h8)
	) name6335 (
		RESET_pad,
		\WX2068_reg/NET0131 ,
		_w7843_
	);
	LUT2 #(
		.INIT('h8)
	) name6336 (
		RESET_pad,
		\WX823_reg/NET0131 ,
		_w7844_
	);
	LUT2 #(
		.INIT('h8)
	) name6337 (
		RESET_pad,
		\WX5941_reg/NET0131 ,
		_w7845_
	);
	LUT2 #(
		.INIT('h8)
	) name6338 (
		RESET_pad,
		\WX11093_reg/NET0131 ,
		_w7846_
	);
	LUT2 #(
		.INIT('h8)
	) name6339 (
		RESET_pad,
		\WX5919_reg/NET0131 ,
		_w7847_
	);
	LUT2 #(
		.INIT('h8)
	) name6340 (
		RESET_pad,
		\WX7160_reg/NET0131 ,
		_w7848_
	);
	LUT2 #(
		.INIT('h8)
	) name6341 (
		RESET_pad,
		\WX791_reg/NET0131 ,
		_w7849_
	);
	LUT2 #(
		.INIT('h8)
	) name6342 (
		RESET_pad,
		\WX11095_reg/NET0131 ,
		_w7850_
	);
	LUT2 #(
		.INIT('h8)
	) name6343 (
		RESET_pad,
		\WX3349_reg/NET0131 ,
		_w7851_
	);
	LUT2 #(
		.INIT('h8)
	) name6344 (
		RESET_pad,
		\WX9708_reg/NET0131 ,
		_w7852_
	);
	LUT2 #(
		.INIT('h8)
	) name6345 (
		RESET_pad,
		\WX769_reg/NET0131 ,
		_w7853_
	);
	LUT2 #(
		.INIT('h8)
	) name6346 (
		RESET_pad,
		\WX11153_reg/NET0131 ,
		_w7854_
	);
	LUT2 #(
		.INIT('h8)
	) name6347 (
		RESET_pad,
		\WX7182_reg/NET0131 ,
		_w7855_
	);
	LUT2 #(
		.INIT('h8)
	) name6348 (
		RESET_pad,
		\WX7238_reg/NET0131 ,
		_w7856_
	);
	LUT2 #(
		.INIT('h8)
	) name6349 (
		RESET_pad,
		\WX11103_reg/NET0131 ,
		_w7857_
	);
	LUT2 #(
		.INIT('h8)
	) name6350 (
		RESET_pad,
		\WX5925_reg/NET0131 ,
		_w7858_
	);
	LUT2 #(
		.INIT('h8)
	) name6351 (
		RESET_pad,
		\WX7196_reg/NET0131 ,
		_w7859_
	);
	LUT2 #(
		.INIT('h8)
	) name6352 (
		RESET_pad,
		\WX7204_reg/NET0131 ,
		_w7860_
	);
	LUT2 #(
		.INIT('h8)
	) name6353 (
		RESET_pad,
		\WX3279_reg/NET0131 ,
		_w7861_
	);
	LUT2 #(
		.INIT('h8)
	) name6354 (
		RESET_pad,
		\WX5953_reg/NET0131 ,
		_w7862_
	);
	LUT2 #(
		.INIT('h8)
	) name6355 (
		RESET_pad,
		\WX3285_reg/NET0131 ,
		_w7863_
	);
	LUT2 #(
		.INIT('h8)
	) name6356 (
		RESET_pad,
		\WX4594_reg/NET0131 ,
		_w7864_
	);
	LUT2 #(
		.INIT('h8)
	) name6357 (
		RESET_pad,
		\WX777_reg/NET0131 ,
		_w7865_
	);
	LUT2 #(
		.INIT('h8)
	) name6358 (
		RESET_pad,
		\WX7164_reg/NET0131 ,
		_w7866_
	);
	LUT2 #(
		.INIT('h8)
	) name6359 (
		RESET_pad,
		\WX11167_reg/NET0131 ,
		_w7867_
	);
	LUT2 #(
		.INIT('h8)
	) name6360 (
		RESET_pad,
		\WX719_reg/NET0131 ,
		_w7868_
	);
	LUT2 #(
		.INIT('h8)
	) name6361 (
		RESET_pad,
		\WX707_reg/NET0131 ,
		_w7869_
	);
	LUT2 #(
		.INIT('h8)
	) name6362 (
		RESET_pad,
		\WX7294_reg/NET0131 ,
		_w7870_
	);
	LUT2 #(
		.INIT('h8)
	) name6363 (
		RESET_pad,
		\WX11113_reg/NET0131 ,
		_w7871_
	);
	LUT2 #(
		.INIT('h8)
	) name6364 (
		RESET_pad,
		\WX1988_reg/NET0131 ,
		_w7872_
	);
	LUT2 #(
		.INIT('h8)
	) name6365 (
		RESET_pad,
		\WX7234_reg/NET0131 ,
		_w7873_
	);
	LUT2 #(
		.INIT('h8)
	) name6366 (
		RESET_pad,
		\WX9712_reg/NET0131 ,
		_w7874_
	);
	LUT2 #(
		.INIT('h8)
	) name6367 (
		RESET_pad,
		\WX5929_reg/NET0131 ,
		_w7875_
	);
	LUT2 #(
		.INIT('h8)
	) name6368 (
		RESET_pad,
		\WX7244_reg/NET0131 ,
		_w7876_
	);
	LUT2 #(
		.INIT('h8)
	) name6369 (
		RESET_pad,
		\WX7248_reg/NET0131 ,
		_w7877_
	);
	LUT2 #(
		.INIT('h8)
	) name6370 (
		RESET_pad,
		\WX9882_reg/NET0131 ,
		_w7878_
	);
	LUT2 #(
		.INIT('h8)
	) name6371 (
		RESET_pad,
		\WX4550_reg/NET0131 ,
		_w7879_
	);
	LUT2 #(
		.INIT('h8)
	) name6372 (
		RESET_pad,
		\WX665_reg/NET0131 ,
		_w7880_
	);
	LUT2 #(
		.INIT('h8)
	) name6373 (
		RESET_pad,
		\WX7232_reg/NET0131 ,
		_w7881_
	);
	LUT2 #(
		.INIT('h8)
	) name6374 (
		RESET_pad,
		\WX705_reg/NET0131 ,
		_w7882_
	);
	LUT2 #(
		.INIT('h8)
	) name6375 (
		RESET_pad,
		\WX2064_reg/NET0131 ,
		_w7883_
	);
	LUT2 #(
		.INIT('h8)
	) name6376 (
		RESET_pad,
		\WX5927_reg/NET0131 ,
		_w7884_
	);
	LUT2 #(
		.INIT('h8)
	) name6377 (
		RESET_pad,
		\WX9822_reg/NET0131 ,
		_w7885_
	);
	LUT2 #(
		.INIT('h8)
	) name6378 (
		RESET_pad,
		\WX7276_reg/NET0131 ,
		_w7886_
	);
	LUT2 #(
		.INIT('h8)
	) name6379 (
		RESET_pad,
		\WX3277_reg/NET0131 ,
		_w7887_
	);
	LUT2 #(
		.INIT('h8)
	) name6380 (
		RESET_pad,
		\WX7284_reg/NET0131 ,
		_w7888_
	);
	LUT2 #(
		.INIT('h8)
	) name6381 (
		RESET_pad,
		\WX11177_reg/NET0131 ,
		_w7889_
	);
	LUT2 #(
		.INIT('h8)
	) name6382 (
		RESET_pad,
		\WX645_reg/NET0131 ,
		_w7890_
	);
	LUT2 #(
		.INIT('h8)
	) name6383 (
		RESET_pad,
		\WX11133_reg/NET0131 ,
		_w7891_
	);
	LUT2 #(
		.INIT('h8)
	) name6384 (
		RESET_pad,
		\WX1992_reg/NET0131 ,
		_w7892_
	);
	LUT2 #(
		.INIT('h8)
	) name6385 (
		RESET_pad,
		\WX11135_reg/NET0131 ,
		_w7893_
	);
	LUT2 #(
		.INIT('h8)
	) name6386 (
		RESET_pad,
		\WX11137_reg/NET0131 ,
		_w7894_
	);
	LUT2 #(
		.INIT('h8)
	) name6387 (
		RESET_pad,
		\WX2072_reg/NET0131 ,
		_w7895_
	);
	LUT2 #(
		.INIT('h8)
	) name6388 (
		RESET_pad,
		\WX11161_reg/NET0131 ,
		_w7896_
	);
	LUT2 #(
		.INIT('h8)
	) name6389 (
		RESET_pad,
		\WX5933_reg/NET0131 ,
		_w7897_
	);
	LUT2 #(
		.INIT('h8)
	) name6390 (
		RESET_pad,
		\WX3379_reg/NET0131 ,
		_w7898_
	);
	LUT2 #(
		.INIT('h8)
	) name6391 (
		RESET_pad,
		\WX4556_reg/NET0131 ,
		_w7899_
	);
	LUT2 #(
		.INIT('h8)
	) name6392 (
		RESET_pad,
		\WX11143_reg/NET0131 ,
		_w7900_
	);
	LUT2 #(
		.INIT('h8)
	) name6393 (
		RESET_pad,
		\WX9750_reg/NET0131 ,
		_w7901_
	);
	LUT2 #(
		.INIT('h8)
	) name6394 (
		RESET_pad,
		\WX9786_reg/NET0131 ,
		_w7902_
	);
	LUT2 #(
		.INIT('h8)
	) name6395 (
		RESET_pad,
		\WX7230_reg/NET0131 ,
		_w7903_
	);
	LUT2 #(
		.INIT('h8)
	) name6396 (
		RESET_pad,
		\WX3237_reg/NET0131 ,
		_w7904_
	);
	LUT2 #(
		.INIT('h8)
	) name6397 (
		RESET_pad,
		\WX11041_reg/NET0131 ,
		_w7905_
	);
	LUT2 #(
		.INIT('h8)
	) name6398 (
		RESET_pad,
		\WX5939_reg/NET0131 ,
		_w7906_
	);
	LUT2 #(
		.INIT('h8)
	) name6399 (
		RESET_pad,
		\WX9716_reg/NET0131 ,
		_w7907_
	);
	LUT2 #(
		.INIT('h8)
	) name6400 (
		RESET_pad,
		\WX5871_reg/NET0131 ,
		_w7908_
	);
	LUT2 #(
		.INIT('h8)
	) name6401 (
		RESET_pad,
		\WX757_reg/NET0131 ,
		_w7909_
	);
	LUT2 #(
		.INIT('h8)
	) name6402 (
		RESET_pad,
		\WX11045_reg/NET0131 ,
		_w7910_
	);
	LUT2 #(
		.INIT('h8)
	) name6403 (
		RESET_pad,
		\WX9744_reg/NET0131 ,
		_w7911_
	);
	LUT2 #(
		.INIT('h8)
	) name6404 (
		RESET_pad,
		\WX9762_reg/NET0131 ,
		_w7912_
	);
	LUT2 #(
		.INIT('h8)
	) name6405 (
		RESET_pad,
		\WX4558_reg/NET0131 ,
		_w7913_
	);
	LUT2 #(
		.INIT('h8)
	) name6406 (
		RESET_pad,
		\WX3273_reg/NET0131 ,
		_w7914_
	);
	LUT2 #(
		.INIT('h8)
	) name6407 (
		RESET_pad,
		\WX5945_reg/NET0131 ,
		_w7915_
	);
	LUT2 #(
		.INIT('h8)
	) name6408 (
		RESET_pad,
		\WX9860_reg/NET0131 ,
		_w7916_
	);
	LUT2 #(
		.INIT('h8)
	) name6409 (
		RESET_pad,
		\WX7228_reg/NET0131 ,
		_w7917_
	);
	LUT2 #(
		.INIT('h8)
	) name6410 (
		RESET_pad,
		\WX7226_reg/NET0131 ,
		_w7918_
	);
	LUT2 #(
		.INIT('h8)
	) name6411 (
		RESET_pad,
		\WX4542_reg/NET0131 ,
		_w7919_
	);
	LUT2 #(
		.INIT('h8)
	) name6412 (
		RESET_pad,
		\WX9808_reg/NET0131 ,
		_w7920_
	);
	LUT2 #(
		.INIT('h8)
	) name6413 (
		RESET_pad,
		\WX11109_reg/NET0131 ,
		_w7921_
	);
	LUT2 #(
		.INIT('h8)
	) name6414 (
		RESET_pad,
		\WX8423_reg/NET0131 ,
		_w7922_
	);
	LUT2 #(
		.INIT('h8)
	) name6415 (
		RESET_pad,
		\WX3327_reg/NET0131 ,
		_w7923_
	);
	LUT2 #(
		.INIT('h8)
	) name6416 (
		RESET_pad,
		\WX807_reg/NET0131 ,
		_w7924_
	);
	LUT2 #(
		.INIT('h8)
	) name6417 (
		RESET_pad,
		\WX8533_reg/NET0131 ,
		_w7925_
	);
	LUT2 #(
		.INIT('h8)
	) name6418 (
		RESET_pad,
		\WX7222_reg/NET0131 ,
		_w7926_
	);
	LUT2 #(
		.INIT('h8)
	) name6419 (
		RESET_pad,
		\WX9856_reg/NET0131 ,
		_w7927_
	);
	LUT2 #(
		.INIT('h8)
	) name6420 (
		RESET_pad,
		\WX1984_reg/NET0131 ,
		_w7928_
	);
	LUT2 #(
		.INIT('h8)
	) name6421 (
		RESET_pad,
		\WX7118_reg/NET0131 ,
		_w7929_
	);
	LUT2 #(
		.INIT('h8)
	) name6422 (
		RESET_pad,
		\WX7218_reg/NET0131 ,
		_w7930_
	);
	LUT2 #(
		.INIT('h8)
	) name6423 (
		RESET_pad,
		\WX7224_reg/NET0131 ,
		_w7931_
	);
	LUT2 #(
		.INIT('h8)
	) name6424 (
		RESET_pad,
		\WX4544_reg/NET0131 ,
		_w7932_
	);
	LUT2 #(
		.INIT('h8)
	) name6425 (
		RESET_pad,
		\WX4560_reg/NET0131 ,
		_w7933_
	);
	LUT2 #(
		.INIT('h8)
	) name6426 (
		RESET_pad,
		\WX667_reg/NET0131 ,
		_w7934_
	);
	LUT2 #(
		.INIT('h8)
	) name6427 (
		RESET_pad,
		\WX7214_reg/NET0131 ,
		_w7935_
	);
	LUT2 #(
		.INIT('h8)
	) name6428 (
		RESET_pad,
		\WX3319_reg/NET0131 ,
		_w7936_
	);
	LUT2 #(
		.INIT('h8)
	) name6429 (
		RESET_pad,
		\WX663_reg/NET0131 ,
		_w7937_
	);
	LUT2 #(
		.INIT('h8)
	) name6430 (
		RESET_pad,
		\WX4598_reg/NET0131 ,
		_w7938_
	);
	LUT2 #(
		.INIT('h8)
	) name6431 (
		RESET_pad,
		\WX9820_reg/NET0131 ,
		_w7939_
	);
	LUT2 #(
		.INIT('h8)
	) name6432 (
		RESET_pad,
		\WX5979_reg/NET0131 ,
		_w7940_
	);
	LUT2 #(
		.INIT('h8)
	) name6433 (
		RESET_pad,
		\WX11107_reg/NET0131 ,
		_w7941_
	);
	LUT2 #(
		.INIT('h8)
	) name6434 (
		RESET_pad,
		\WX9698_reg/NET0131 ,
		_w7942_
	);
	LUT2 #(
		.INIT('h8)
	) name6435 (
		RESET_pad,
		\WX7198_reg/NET0131 ,
		_w7943_
	);
	LUT2 #(
		.INIT('h8)
	) name6436 (
		RESET_pad,
		\WX3365_reg/NET0131 ,
		_w7944_
	);
	LUT2 #(
		.INIT('h8)
	) name6437 (
		RESET_pad,
		\WX11131_reg/NET0131 ,
		_w7945_
	);
	LUT2 #(
		.INIT('h8)
	) name6438 (
		RESET_pad,
		\WX3361_reg/NET0131 ,
		_w7946_
	);
	LUT2 #(
		.INIT('h8)
	) name6439 (
		RESET_pad,
		\WX11163_reg/NET0131 ,
		_w7947_
	);
	LUT2 #(
		.INIT('h8)
	) name6440 (
		RESET_pad,
		\WX8517_reg/NET0131 ,
		_w7948_
	);
	LUT2 #(
		.INIT('h8)
	) name6441 (
		RESET_pad,
		\WX9772_reg/NET0131 ,
		_w7949_
	);
	LUT2 #(
		.INIT('h8)
	) name6442 (
		RESET_pad,
		\WX11105_reg/NET0131 ,
		_w7950_
	);
	LUT2 #(
		.INIT('h8)
	) name6443 (
		RESET_pad,
		\WX11123_reg/NET0131 ,
		_w7951_
	);
	LUT2 #(
		.INIT('h8)
	) name6444 (
		RESET_pad,
		\WX3351_reg/NET0131 ,
		_w7952_
	);
	LUT2 #(
		.INIT('h8)
	) name6445 (
		RESET_pad,
		\WX4562_reg/NET0131 ,
		_w7953_
	);
	LUT2 #(
		.INIT('h8)
	) name6446 (
		RESET_pad,
		\WX4540_reg/NET0131 ,
		_w7954_
	);
	LUT2 #(
		.INIT('h8)
	) name6447 (
		RESET_pad,
		\WX5879_reg/NET0131 ,
		_w7955_
	);
	LUT2 #(
		.INIT('h8)
	) name6448 (
		RESET_pad,
		\WX5875_reg/NET0131 ,
		_w7956_
	);
	LUT2 #(
		.INIT('h8)
	) name6449 (
		RESET_pad,
		\WX5991_reg/NET0131 ,
		_w7957_
	);
	LUT2 #(
		.INIT('h8)
	) name6450 (
		RESET_pad,
		\WX2056_reg/NET0131 ,
		_w7958_
	);
	LUT2 #(
		.INIT('h8)
	) name6451 (
		RESET_pad,
		\WX3263_reg/NET0131 ,
		_w7959_
	);
	LUT2 #(
		.INIT('h8)
	) name6452 (
		RESET_pad,
		\WX7166_reg/NET0131 ,
		_w7960_
	);
	LUT2 #(
		.INIT('h8)
	) name6453 (
		RESET_pad,
		\WX7190_reg/NET0131 ,
		_w7961_
	);
	LUT2 #(
		.INIT('h8)
	) name6454 (
		RESET_pad,
		\WX1972_reg/NET0131 ,
		_w7962_
	);
	LUT2 #(
		.INIT('h8)
	) name6455 (
		RESET_pad,
		\WX661_reg/NET0131 ,
		_w7963_
	);
	LUT2 #(
		.INIT('h8)
	) name6456 (
		RESET_pad,
		\WX9774_reg/NET0131 ,
		_w7964_
	);
	LUT2 #(
		.INIT('h8)
	) name6457 (
		RESET_pad,
		\WX1994_reg/NET0131 ,
		_w7965_
	);
	LUT2 #(
		.INIT('h8)
	) name6458 (
		RESET_pad,
		\WX7256_reg/NET0131 ,
		_w7966_
	);
	LUT2 #(
		.INIT('h8)
	) name6459 (
		RESET_pad,
		\WX5985_reg/NET0131 ,
		_w7967_
	);
	LUT2 #(
		.INIT('h8)
	) name6460 (
		RESET_pad,
		\WX7192_reg/NET0131 ,
		_w7968_
	);
	LUT2 #(
		.INIT('h8)
	) name6461 (
		RESET_pad,
		\WX7194_reg/NET0131 ,
		_w7969_
	);
	LUT2 #(
		.INIT('h8)
	) name6462 (
		RESET_pad,
		\WX8445_reg/NET0131 ,
		_w7970_
	);
	LUT2 #(
		.INIT('h8)
	) name6463 (
		RESET_pad,
		\WX5999_reg/NET0131 ,
		_w7971_
	);
	LUT2 #(
		.INIT('h8)
	) name6464 (
		RESET_pad,
		\WX1966_reg/NET0131 ,
		_w7972_
	);
	LUT2 #(
		.INIT('h8)
	) name6465 (
		RESET_pad,
		\WX9726_reg/NET0131 ,
		_w7973_
	);
	LUT2 #(
		.INIT('h8)
	) name6466 (
		RESET_pad,
		\WX9704_reg/NET0131 ,
		_w7974_
	);
	LUT2 #(
		.INIT('h8)
	) name6467 (
		RESET_pad,
		\WX7186_reg/NET0131 ,
		_w7975_
	);
	LUT2 #(
		.INIT('h8)
	) name6468 (
		RESET_pad,
		\WX8441_reg/NET0131 ,
		_w7976_
	);
	LUT2 #(
		.INIT('h8)
	) name6469 (
		RESET_pad,
		\WX5923_reg/NET0131 ,
		_w7977_
	);
	LUT2 #(
		.INIT('h8)
	) name6470 (
		RESET_pad,
		\WX2128_reg/NET0131 ,
		_w7978_
	);
	LUT2 #(
		.INIT('h8)
	) name6471 (
		RESET_pad,
		\WX2126_reg/NET0131 ,
		_w7979_
	);
	LUT2 #(
		.INIT('h8)
	) name6472 (
		RESET_pad,
		\WX7180_reg/NET0131 ,
		_w7980_
	);
	LUT2 #(
		.INIT('h8)
	) name6473 (
		RESET_pad,
		\WX721_reg/NET0131 ,
		_w7981_
	);
	LUT2 #(
		.INIT('h8)
	) name6474 (
		RESET_pad,
		\WX7278_reg/NET0131 ,
		_w7982_
	);
	LUT2 #(
		.INIT('h8)
	) name6475 (
		RESET_pad,
		\WX835_reg/NET0131 ,
		_w7983_
	);
	LUT2 #(
		.INIT('h8)
	) name6476 (
		RESET_pad,
		\WX5997_reg/NET0131 ,
		_w7984_
	);
	LUT2 #(
		.INIT('h8)
	) name6477 (
		RESET_pad,
		\WX3363_reg/NET0131 ,
		_w7985_
	);
	LUT2 #(
		.INIT('h8)
	) name6478 (
		RESET_pad,
		\WX5921_reg/NET0131 ,
		_w7986_
	);
	LUT2 #(
		.INIT('h8)
	) name6479 (
		RESET_pad,
		\WX659_reg/NET0131 ,
		_w7987_
	);
	LUT2 #(
		.INIT('h8)
	) name6480 (
		RESET_pad,
		\WX3259_reg/NET0131 ,
		_w7988_
	);
	LUT2 #(
		.INIT('h8)
	) name6481 (
		RESET_pad,
		\WX9780_reg/NET0131 ,
		_w7989_
	);
	LUT2 #(
		.INIT('h8)
	) name6482 (
		RESET_pad,
		\WX1956_reg/NET0131 ,
		_w7990_
	);
	LUT2 #(
		.INIT('h8)
	) name6483 (
		RESET_pad,
		\WX11099_reg/NET0131 ,
		_w7991_
	);
	LUT2 #(
		.INIT('h8)
	) name6484 (
		RESET_pad,
		\WX2088_reg/NET0131 ,
		_w7992_
	);
	LUT2 #(
		.INIT('h8)
	) name6485 (
		RESET_pad,
		\WX9800_reg/NET0131 ,
		_w7993_
	);
	LUT2 #(
		.INIT('h8)
	) name6486 (
		RESET_pad,
		\WX767_reg/NET0131 ,
		_w7994_
	);
	LUT2 #(
		.INIT('h8)
	) name6487 (
		RESET_pad,
		\WX7280_reg/NET0131 ,
		_w7995_
	);
	LUT2 #(
		.INIT('h8)
	) name6488 (
		RESET_pad,
		\WX8519_reg/NET0131 ,
		_w7996_
	);
	LUT2 #(
		.INIT('h8)
	) name6489 (
		RESET_pad,
		\WX771_reg/NET0131 ,
		_w7997_
	);
	LUT2 #(
		.INIT('h8)
	) name6490 (
		RESET_pad,
		\WX781_reg/NET0131 ,
		_w7998_
	);
	LUT2 #(
		.INIT('h8)
	) name6491 (
		RESET_pad,
		\WX1958_reg/NET0131 ,
		_w7999_
	);
	LUT2 #(
		.INIT('h8)
	) name6492 (
		RESET_pad,
		\WX3289_reg/NET0131 ,
		_w8000_
	);
	LUT2 #(
		.INIT('h8)
	) name6493 (
		RESET_pad,
		\WX4638_reg/NET0131 ,
		_w8001_
	);
	LUT2 #(
		.INIT('h8)
	) name6494 (
		RESET_pad,
		\WX687_reg/NET0131 ,
		_w8002_
	);
	LUT2 #(
		.INIT('h8)
	) name6495 (
		RESET_pad,
		\WX2112_reg/NET0131 ,
		_w8003_
	);
	LUT2 #(
		.INIT('h8)
	) name6496 (
		RESET_pad,
		\WX9730_reg/NET0131 ,
		_w8004_
	);
	LUT2 #(
		.INIT('h8)
	) name6497 (
		RESET_pad,
		\WX9754_reg/NET0131 ,
		_w8005_
	);
	LUT2 #(
		.INIT('h8)
	) name6498 (
		RESET_pad,
		\WX787_reg/NET0131 ,
		_w8006_
	);
	LUT2 #(
		.INIT('h8)
	) name6499 (
		RESET_pad,
		\WX731_reg/NET0131 ,
		_w8007_
	);
	LUT2 #(
		.INIT('h8)
	) name6500 (
		RESET_pad,
		\WX3415_reg/NET0131 ,
		_w8008_
	);
	LUT2 #(
		.INIT('h8)
	) name6501 (
		RESET_pad,
		\WX3255_reg/NET0131 ,
		_w8009_
	);
	LUT2 #(
		.INIT('h8)
	) name6502 (
		RESET_pad,
		\WX2122_reg/NET0131 ,
		_w8010_
	);
	LUT2 #(
		.INIT('h8)
	) name6503 (
		RESET_pad,
		\WX8529_reg/NET0131 ,
		_w8011_
	);
	LUT2 #(
		.INIT('h8)
	) name6504 (
		RESET_pad,
		\WX9832_reg/NET0131 ,
		_w8012_
	);
	LUT2 #(
		.INIT('h8)
	) name6505 (
		RESET_pad,
		\WX8449_reg/NET0131 ,
		_w8013_
	);
	LUT2 #(
		.INIT('h8)
	) name6506 (
		RESET_pad,
		\WX727_reg/NET0131 ,
		_w8014_
	);
	LUT2 #(
		.INIT('h8)
	) name6507 (
		RESET_pad,
		\WX7158_reg/NET0131 ,
		_w8015_
	);
	LUT2 #(
		.INIT('h8)
	) name6508 (
		RESET_pad,
		\WX11011_reg/NET0131 ,
		_w8016_
	);
	LUT2 #(
		.INIT('h8)
	) name6509 (
		RESET_pad,
		\WX7152_reg/NET0131 ,
		_w8017_
	);
	LUT2 #(
		.INIT('h8)
	) name6510 (
		RESET_pad,
		\WX4676_reg/NET0131 ,
		_w8018_
	);
	LUT2 #(
		.INIT('h8)
	) name6511 (
		RESET_pad,
		\WX7156_reg/NET0131 ,
		_w8019_
	);
	LUT2 #(
		.INIT('h8)
	) name6512 (
		RESET_pad,
		\WX7154_reg/NET0131 ,
		_w8020_
	);
	LUT2 #(
		.INIT('h8)
	) name6513 (
		RESET_pad,
		\WX657_reg/NET0131 ,
		_w8021_
	);
	LUT2 #(
		.INIT('h8)
	) name6514 (
		RESET_pad,
		\WX9816_reg/NET0131 ,
		_w8022_
	);
	LUT2 #(
		.INIT('h8)
	) name6515 (
		RESET_pad,
		\WX831_reg/NET0131 ,
		_w8023_
	);
	LUT2 #(
		.INIT('h8)
	) name6516 (
		RESET_pad,
		\WX7134_reg/NET0131 ,
		_w8024_
	);
	LUT2 #(
		.INIT('h8)
	) name6517 (
		RESET_pad,
		\WX7246_reg/NET0131 ,
		_w8025_
	);
	LUT2 #(
		.INIT('h8)
	) name6518 (
		RESET_pad,
		\WX7144_reg/NET0131 ,
		_w8026_
	);
	LUT2 #(
		.INIT('h8)
	) name6519 (
		RESET_pad,
		\WX9736_reg/NET0131 ,
		_w8027_
	);
	LUT2 #(
		.INIT('h8)
	) name6520 (
		RESET_pad,
		\WX1946_reg/NET0131 ,
		_w8028_
	);
	LUT2 #(
		.INIT('h8)
	) name6521 (
		RESET_pad,
		\WX7150_reg/NET0131 ,
		_w8029_
	);
	LUT2 #(
		.INIT('h8)
	) name6522 (
		RESET_pad,
		\WX2000_reg/NET0131 ,
		_w8030_
	);
	LUT2 #(
		.INIT('h8)
	) name6523 (
		RESET_pad,
		\WX761_reg/NET0131 ,
		_w8031_
	);
	LUT2 #(
		.INIT('h8)
	) name6524 (
		RESET_pad,
		\WX9842_reg/NET0131 ,
		_w8032_
	);
	LUT2 #(
		.INIT('h8)
	) name6525 (
		RESET_pad,
		\WX819_reg/NET0131 ,
		_w8033_
	);
	LUT2 #(
		.INIT('h8)
	) name6526 (
		RESET_pad,
		\WX7148_reg/NET0131 ,
		_w8034_
	);
	LUT2 #(
		.INIT('h8)
	) name6527 (
		RESET_pad,
		\WX3321_reg/NET0131 ,
		_w8035_
	);
	LUT2 #(
		.INIT('h8)
	) name6528 (
		RESET_pad,
		\WX4634_reg/NET0131 ,
		_w8036_
	);
	LUT2 #(
		.INIT('h8)
	) name6529 (
		RESET_pad,
		\WX11087_reg/NET0131 ,
		_w8037_
	);
	LUT2 #(
		.INIT('h8)
	) name6530 (
		RESET_pad,
		\WX7124_reg/NET0131 ,
		_w8038_
	);
	LUT2 #(
		.INIT('h8)
	) name6531 (
		RESET_pad,
		\WX3301_reg/NET0131 ,
		_w8039_
	);
	LUT2 #(
		.INIT('h8)
	) name6532 (
		RESET_pad,
		\WX3409_reg/NET0131 ,
		_w8040_
	);
	LUT2 #(
		.INIT('h8)
	) name6533 (
		RESET_pad,
		\WX9778_reg/NET0131 ,
		_w8041_
	);
	LUT2 #(
		.INIT('h8)
	) name6534 (
		RESET_pad,
		\WX7272_reg/NET0131 ,
		_w8042_
	);
	LUT2 #(
		.INIT('h8)
	) name6535 (
		RESET_pad,
		\WX7138_reg/NET0131 ,
		_w8043_
	);
	LUT2 #(
		.INIT('h8)
	) name6536 (
		RESET_pad,
		\WX2118_reg/NET0131 ,
		_w8044_
	);
	LUT2 #(
		.INIT('h8)
	) name6537 (
		RESET_pad,
		\WX4626_reg/NET0131 ,
		_w8045_
	);
	LUT2 #(
		.INIT('h8)
	) name6538 (
		RESET_pad,
		\WX5949_reg/NET0131 ,
		_w8046_
	);
	LUT2 #(
		.INIT('h8)
	) name6539 (
		RESET_pad,
		\WX693_reg/NET0131 ,
		_w8047_
	);
	LUT2 #(
		.INIT('h8)
	) name6540 (
		RESET_pad,
		\WX3265_reg/NET0131 ,
		_w8048_
	);
	LUT2 #(
		.INIT('h8)
	) name6541 (
		RESET_pad,
		\WX11141_reg/NET0131 ,
		_w8049_
	);
	LUT2 #(
		.INIT('h8)
	) name6542 (
		RESET_pad,
		\WX5947_reg/NET0131 ,
		_w8050_
	);
	LUT2 #(
		.INIT('h8)
	) name6543 (
		RESET_pad,
		\WX2114_reg/NET0131 ,
		_w8051_
	);
	LUT2 #(
		.INIT('h8)
	) name6544 (
		RESET_pad,
		\WX4584_reg/NET0131 ,
		_w8052_
	);
	LUT2 #(
		.INIT('h8)
	) name6545 (
		RESET_pad,
		\WX735_reg/NET0131 ,
		_w8053_
	);
	LUT2 #(
		.INIT('h8)
	) name6546 (
		RESET_pad,
		\WX3267_reg/NET0131 ,
		_w8054_
	);
	LUT2 #(
		.INIT('h8)
	) name6547 (
		RESET_pad,
		\WX7120_reg/NET0131 ,
		_w8055_
	);
	LUT2 #(
		.INIT('h8)
	) name6548 (
		RESET_pad,
		\WX7132_reg/NET0131 ,
		_w8056_
	);
	LUT2 #(
		.INIT('h8)
	) name6549 (
		RESET_pad,
		\WX3357_reg/NET0131 ,
		_w8057_
	);
	LUT2 #(
		.INIT('h8)
	) name6550 (
		RESET_pad,
		\WX3281_reg/NET0131 ,
		_w8058_
	);
	LUT2 #(
		.INIT('h8)
	) name6551 (
		RESET_pad,
		\WX3247_reg/NET0131 ,
		_w8059_
	);
	LUT2 #(
		.INIT('h8)
	) name6552 (
		RESET_pad,
		\WX9798_reg/NET0131 ,
		_w8060_
	);
	LUT2 #(
		.INIT('h8)
	) name6553 (
		RESET_pad,
		\WX11119_reg/NET0131 ,
		_w8061_
	);
	LUT2 #(
		.INIT('h8)
	) name6554 (
		RESET_pad,
		\WX7126_reg/NET0131 ,
		_w8062_
	);
	LUT2 #(
		.INIT('h8)
	) name6555 (
		RESET_pad,
		\WX5937_reg/NET0131 ,
		_w8063_
	);
	LUT2 #(
		.INIT('h8)
	) name6556 (
		RESET_pad,
		\WX7128_reg/NET0131 ,
		_w8064_
	);
	LUT2 #(
		.INIT('h8)
	) name6557 (
		RESET_pad,
		\WX3347_reg/NET0131 ,
		_w8065_
	);
	LUT2 #(
		.INIT('h8)
	) name6558 (
		RESET_pad,
		\WX2060_reg/NET0131 ,
		_w8066_
	);
	LUT2 #(
		.INIT('h8)
	) name6559 (
		RESET_pad,
		\WX7130_reg/NET0131 ,
		_w8067_
	);
	LUT2 #(
		.INIT('h8)
	) name6560 (
		RESET_pad,
		\WX9742_reg/NET0131 ,
		_w8068_
	);
	LUT2 #(
		.INIT('h8)
	) name6561 (
		RESET_pad,
		\WX11085_reg/NET0131 ,
		_w8069_
	);
	LUT2 #(
		.INIT('h8)
	) name6562 (
		RESET_pad,
		\WX11043_reg/NET0131 ,
		_w8070_
	);
	LUT2 #(
		.INIT('h8)
	) name6563 (
		RESET_pad,
		\WX3283_reg/NET0131 ,
		_w8071_
	);
	LUT2 #(
		.INIT('h8)
	) name6564 (
		RESET_pad,
		\WX755_reg/NET0131 ,
		_w8072_
	);
	LUT2 #(
		.INIT('h8)
	) name6565 (
		RESET_pad,
		\WX8447_reg/NET0131 ,
		_w8073_
	);
	LUT2 #(
		.INIT('h8)
	) name6566 (
		RESET_pad,
		\WX669_reg/NET0131 ,
		_w8074_
	);
	LUT2 #(
		.INIT('h8)
	) name6567 (
		RESET_pad,
		\WX4564_reg/NET0131 ,
		_w8075_
	);
	LUT2 #(
		.INIT('h8)
	) name6568 (
		RESET_pad,
		\WX685_reg/NET0131 ,
		_w8076_
	);
	LUT2 #(
		.INIT('h8)
	) name6569 (
		RESET_pad,
		\WX11067_reg/NET0131 ,
		_w8077_
	);
	LUT2 #(
		.INIT('h8)
	) name6570 (
		RESET_pad,
		\WX8453_reg/NET0131 ,
		_w8078_
	);
	LUT2 #(
		.INIT('h8)
	) name6571 (
		RESET_pad,
		\WX4538_reg/NET0131 ,
		_w8079_
	);
	LUT2 #(
		.INIT('h8)
	) name6572 (
		RESET_pad,
		\WX5959_reg/NET0131 ,
		_w8080_
	);
	LUT2 #(
		.INIT('h8)
	) name6573 (
		RESET_pad,
		\WX3355_reg/NET0131 ,
		_w8081_
	);
	LUT2 #(
		.INIT('h8)
	) name6574 (
		RESET_pad,
		\WX4588_reg/NET0131 ,
		_w8082_
	);
	LUT2 #(
		.INIT('h8)
	) name6575 (
		RESET_pad,
		\WX9724_reg/NET0131 ,
		_w8083_
	);
	LUT2 #(
		.INIT('h8)
	) name6576 (
		RESET_pad,
		\WX5965_reg/NET0131 ,
		_w8084_
	);
	LUT2 #(
		.INIT('h8)
	) name6577 (
		RESET_pad,
		\WX11147_reg/NET0131 ,
		_w8085_
	);
	LUT2 #(
		.INIT('h8)
	) name6578 (
		RESET_pad,
		\WX7122_reg/NET0131 ,
		_w8086_
	);
	LUT2 #(
		.INIT('h8)
	) name6579 (
		RESET_pad,
		\WX695_reg/NET0131 ,
		_w8087_
	);
	LUT2 #(
		.INIT('h8)
	) name6580 (
		RESET_pad,
		\WX4636_reg/NET0131 ,
		_w8088_
	);
	LUT2 #(
		.INIT('h8)
	) name6581 (
		RESET_pad,
		\WX4628_reg/NET0131 ,
		_w8089_
	);
	LUT2 #(
		.INIT('h8)
	) name6582 (
		RESET_pad,
		\WX8551_reg/NET0131 ,
		_w8090_
	);
	LUT2 #(
		.INIT('h8)
	) name6583 (
		RESET_pad,
		\WX9872_reg/NET0131 ,
		_w8091_
	);
	LUT2 #(
		.INIT('h8)
	) name6584 (
		RESET_pad,
		\WX5861_reg/NET0131 ,
		_w8092_
	);
	LUT2 #(
		.INIT('h8)
	) name6585 (
		RESET_pad,
		\WX8407_reg/NET0131 ,
		_w8093_
	);
	LUT2 #(
		.INIT('h8)
	) name6586 (
		RESET_pad,
		\WX8547_reg/NET0131 ,
		_w8094_
	);
	LUT2 #(
		.INIT('h8)
	) name6587 (
		RESET_pad,
		\WX9862_reg/NET0131 ,
		_w8095_
	);
	LUT2 #(
		.INIT('h8)
	) name6588 (
		RESET_pad,
		\WX4570_reg/NET0131 ,
		_w8096_
	);
	LUT2 #(
		.INIT('h8)
	) name6589 (
		RESET_pad,
		\WX11027_reg/NET0131 ,
		_w8097_
	);
	LUT2 #(
		.INIT('h8)
	) name6590 (
		RESET_pad,
		\WX11139_reg/NET0131 ,
		_w8098_
	);
	LUT2 #(
		.INIT('h8)
	) name6591 (
		RESET_pad,
		\WX4652_reg/NET0131 ,
		_w8099_
	);
	LUT2 #(
		.INIT('h8)
	) name6592 (
		RESET_pad,
		\WX729_reg/NET0131 ,
		_w8100_
	);
	LUT2 #(
		.INIT('h8)
	) name6593 (
		RESET_pad,
		\WX5957_reg/NET0131 ,
		_w8101_
	);
	LUT2 #(
		.INIT('h8)
	) name6594 (
		RESET_pad,
		\WX3287_reg/NET0131 ,
		_w8102_
	);
	LUT2 #(
		.INIT('h8)
	) name6595 (
		RESET_pad,
		\WX801_reg/NET0131 ,
		_w8103_
	);
	LUT2 #(
		.INIT('h8)
	) name6596 (
		RESET_pad,
		\WX805_reg/NET0131 ,
		_w8104_
	);
	LUT2 #(
		.INIT('h8)
	) name6597 (
		RESET_pad,
		\WX11149_reg/NET0131 ,
		_w8105_
	);
	LUT2 #(
		.INIT('h8)
	) name6598 (
		RESET_pad,
		\WX691_reg/NET0131 ,
		_w8106_
	);
	LUT2 #(
		.INIT('h8)
	) name6599 (
		RESET_pad,
		\WX8557_reg/NET0131 ,
		_w8107_
	);
	LUT2 #(
		.INIT('h8)
	) name6600 (
		RESET_pad,
		\WX9722_reg/NET0131 ,
		_w8108_
	);
	LUT2 #(
		.INIT('h8)
	) name6601 (
		RESET_pad,
		\WX9840_reg/NET0131 ,
		_w8109_
	);
	LUT2 #(
		.INIT('h8)
	) name6602 (
		RESET_pad,
		\WX9764_reg/NET0131 ,
		_w8110_
	);
	LUT2 #(
		.INIT('h8)
	) name6603 (
		RESET_pad,
		\WX2076_reg/NET0131 ,
		_w8111_
	);
	LUT2 #(
		.INIT('h8)
	) name6604 (
		RESET_pad,
		\WX7116_reg/NET0131 ,
		_w8112_
	);
	LUT2 #(
		.INIT('h8)
	) name6605 (
		RESET_pad,
		\WX9796_reg/NET0131 ,
		_w8113_
	);
	LUT2 #(
		.INIT('h8)
	) name6606 (
		RESET_pad,
		\WX9776_reg/NET0131 ,
		_w8114_
	);
	LUT2 #(
		.INIT('h8)
	) name6607 (
		RESET_pad,
		\WX11071_reg/NET0131 ,
		_w8115_
	);
	LUT2 #(
		.INIT('h8)
	) name6608 (
		RESET_pad,
		\WX9760_reg/NET0131 ,
		_w8116_
	);
	LUT2 #(
		.INIT('h8)
	) name6609 (
		RESET_pad,
		\WX4576_reg/NET0131 ,
		_w8117_
	);
	LUT2 #(
		.INIT('h8)
	) name6610 (
		RESET_pad,
		\WX803_reg/NET0131 ,
		_w8118_
	);
	LUT2 #(
		.INIT('h8)
	) name6611 (
		RESET_pad,
		\WX3395_reg/NET0131 ,
		_w8119_
	);
	LUT2 #(
		.INIT('h8)
	) name6612 (
		RESET_pad,
		\WX4526_reg/NET0131 ,
		_w8120_
	);
	LUT2 #(
		.INIT('h8)
	) name6613 (
		RESET_pad,
		\WX9790_reg/NET0131 ,
		_w8121_
	);
	LUT2 #(
		.INIT('h8)
	) name6614 (
		RESET_pad,
		\WX9768_reg/NET0131 ,
		_w8122_
	);
	LUT2 #(
		.INIT('h8)
	) name6615 (
		RESET_pad,
		\WX653_reg/NET0131 ,
		_w8123_
	);
	LUT2 #(
		.INIT('h8)
	) name6616 (
		RESET_pad,
		\WX4662_reg/NET0131 ,
		_w8124_
	);
	LUT2 #(
		.INIT('h8)
	) name6617 (
		RESET_pad,
		\WX4580_reg/NET0131 ,
		_w8125_
	);
	LUT2 #(
		.INIT('h8)
	) name6618 (
		RESET_pad,
		\WX9728_reg/NET0131 ,
		_w8126_
	);
	LUT2 #(
		.INIT('h8)
	) name6619 (
		RESET_pad,
		\WX9718_reg/NET0131 ,
		_w8127_
	);
	LUT2 #(
		.INIT('h8)
	) name6620 (
		RESET_pad,
		\WX3405_reg/NET0131 ,
		_w8128_
	);
	LUT2 #(
		.INIT('h8)
	) name6621 (
		RESET_pad,
		\WX3245_reg/NET0131 ,
		_w8129_
	);
	LUT2 #(
		.INIT('h8)
	) name6622 (
		RESET_pad,
		\WX2010_reg/NET0131 ,
		_w8130_
	);
	LUT2 #(
		.INIT('h8)
	) name6623 (
		RESET_pad,
		\WX4682_reg/NET0131 ,
		_w8131_
	);
	LUT2 #(
		.INIT('h8)
	) name6624 (
		RESET_pad,
		\WX8589_reg/NET0131 ,
		_w8132_
	);
	LUT2 #(
		.INIT('h8)
	) name6625 (
		RESET_pad,
		\WX4688_reg/NET0131 ,
		_w8133_
	);
	LUT2 #(
		.INIT('h8)
	) name6626 (
		RESET_pad,
		\WX9706_reg/NET0131 ,
		_w8134_
	);
	LUT2 #(
		.INIT('h8)
	) name6627 (
		RESET_pad,
		\WX4690_reg/NET0131 ,
		_w8135_
	);
	LUT2 #(
		.INIT('h8)
	) name6628 (
		RESET_pad,
		\WX3243_reg/NET0131 ,
		_w8136_
	);
	LUT2 #(
		.INIT('h8)
	) name6629 (
		RESET_pad,
		\WX3241_reg/NET0131 ,
		_w8137_
	);
	LUT2 #(
		.INIT('h8)
	) name6630 (
		RESET_pad,
		\WX4698_reg/NET0131 ,
		_w8138_
	);
	LUT2 #(
		.INIT('h8)
	) name6631 (
		RESET_pad,
		\WX8591_reg/NET0131 ,
		_w8139_
	);
	LUT2 #(
		.INIT('h8)
	) name6632 (
		RESET_pad,
		\WX3239_reg/NET0131 ,
		_w8140_
	);
	LUT2 #(
		.INIT('h8)
	) name6633 (
		RESET_pad,
		\WX4704_reg/NET0131 ,
		_w8141_
	);
	LUT2 #(
		.INIT('h8)
	) name6634 (
		RESET_pad,
		\WX8583_reg/NET0131 ,
		_w8142_
	);
	LUT2 #(
		.INIT('h8)
	) name6635 (
		RESET_pad,
		\WX11029_reg/NET0131 ,
		_w8143_
	);
	LUT2 #(
		.INIT('h8)
	) name6636 (
		RESET_pad,
		\WX4712_reg/NET0131 ,
		_w8144_
	);
	LUT2 #(
		.INIT('h8)
	) name6637 (
		RESET_pad,
		\WX743_reg/NET0131 ,
		_w8145_
	);
	LUT2 #(
		.INIT('h8)
	) name6638 (
		RESET_pad,
		\WX8565_reg/NET0131 ,
		_w8146_
	);
	LUT2 #(
		.INIT('h8)
	) name6639 (
		RESET_pad,
		\WX8579_reg/NET0131 ,
		_w8147_
	);
	LUT2 #(
		.INIT('h8)
	) name6640 (
		RESET_pad,
		\WX3383_reg/NET0131 ,
		_w8148_
	);
	LUT2 #(
		.INIT('h8)
	) name6641 (
		RESET_pad,
		\WX8559_reg/NET0131 ,
		_w8149_
	);
	LUT2 #(
		.INIT('h8)
	) name6642 (
		RESET_pad,
		\WX2104_reg/NET0131 ,
		_w8150_
	);
	LUT2 #(
		.INIT('h8)
	) name6643 (
		RESET_pad,
		\WX4678_reg/NET0131 ,
		_w8151_
	);
	LUT2 #(
		.INIT('h8)
	) name6644 (
		RESET_pad,
		\WX689_reg/NET0131 ,
		_w8152_
	);
	LUT2 #(
		.INIT('h8)
	) name6645 (
		RESET_pad,
		\WX3233_reg/NET0131 ,
		_w8153_
	);
	LUT2 #(
		.INIT('h8)
	) name6646 (
		RESET_pad,
		\WX3393_reg/NET0131 ,
		_w8154_
	);
	LUT2 #(
		.INIT('h8)
	) name6647 (
		RESET_pad,
		\WX8455_reg/NET0131 ,
		_w8155_
	);
	LUT2 #(
		.INIT('h8)
	) name6648 (
		RESET_pad,
		\WX3235_reg/NET0131 ,
		_w8156_
	);
	LUT2 #(
		.INIT('h8)
	) name6649 (
		RESET_pad,
		\WX739_reg/NET0131 ,
		_w8157_
	);
	LUT2 #(
		.INIT('h8)
	) name6650 (
		RESET_pad,
		\WX8567_reg/NET0131 ,
		_w8158_
	);
	LUT2 #(
		.INIT('h8)
	) name6651 (
		RESET_pad,
		\WX8573_reg/NET0131 ,
		_w8159_
	);
	LUT2 #(
		.INIT('h8)
	) name6652 (
		RESET_pad,
		\WX3391_reg/NET0131 ,
		_w8160_
	);
	LUT2 #(
		.INIT('h8)
	) name6653 (
		RESET_pad,
		\WX10995_reg/NET0131 ,
		_w8161_
	);
	LUT2 #(
		.INIT('h8)
	) name6654 (
		RESET_pad,
		\WX8571_reg/NET0131 ,
		_w8162_
	);
	LUT2 #(
		.INIT('h8)
	) name6655 (
		RESET_pad,
		\WX2108_reg/NET0131 ,
		_w8163_
	);
	LUT2 #(
		.INIT('h8)
	) name6656 (
		RESET_pad,
		\WX2008_reg/NET0131 ,
		_w8164_
	);
	LUT2 #(
		.INIT('h8)
	) name6657 (
		RESET_pad,
		\WX7242_reg/NET0131 ,
		_w8165_
	);
	LUT2 #(
		.INIT('h8)
	) name6658 (
		RESET_pad,
		\WX11015_reg/NET0131 ,
		_w8166_
	);
	LUT2 #(
		.INIT('h8)
	) name6659 (
		RESET_pad,
		\WX9864_reg/NET0131 ,
		_w8167_
	);
	LUT2 #(
		.INIT('h8)
	) name6660 (
		RESET_pad,
		\WX3385_reg/NET0131 ,
		_w8168_
	);
	LUT2 #(
		.INIT('h8)
	) name6661 (
		RESET_pad,
		\WX4710_reg/NET0131 ,
		_w8169_
	);
	LUT2 #(
		.INIT('h8)
	) name6662 (
		RESET_pad,
		\WX779_reg/NET0131 ,
		_w8170_
	);
	LUT2 #(
		.INIT('h8)
	) name6663 (
		RESET_pad,
		\WX753_reg/NET0131 ,
		_w8171_
	);
	LUT2 #(
		.INIT('h8)
	) name6664 (
		RESET_pad,
		\WX733_reg/NET0131 ,
		_w8172_
	);
	LUT2 #(
		.INIT('h8)
	) name6665 (
		RESET_pad,
		\WX2012_reg/NET0131 ,
		_w8173_
	);
	LUT2 #(
		.INIT('h8)
	) name6666 (
		RESET_pad,
		\WX2086_reg/NET0131 ,
		_w8174_
	);
	LUT2 #(
		.INIT('h8)
	) name6667 (
		RESET_pad,
		\WX4680_reg/NET0131 ,
		_w8175_
	);
	LUT2 #(
		.INIT('h8)
	) name6668 (
		RESET_pad,
		\WX4696_reg/NET0131 ,
		_w8176_
	);
	LUT2 #(
		.INIT('h8)
	) name6669 (
		RESET_pad,
		\WX8561_reg/NET0131 ,
		_w8177_
	);
	LUT2 #(
		.INIT('h8)
	) name6670 (
		RESET_pad,
		\WX11077_reg/NET0131 ,
		_w8178_
	);
	LUT2 #(
		.INIT('h8)
	) name6671 (
		RESET_pad,
		\WX2106_reg/NET0131 ,
		_w8179_
	);
	LUT2 #(
		.INIT('h8)
	) name6672 (
		RESET_pad,
		\WX4686_reg/NET0131 ,
		_w8180_
	);
	LUT2 #(
		.INIT('h8)
	) name6673 (
		RESET_pad,
		\WX3335_reg/NET0131 ,
		_w8181_
	);
	LUT2 #(
		.INIT('h8)
	) name6674 (
		RESET_pad,
		\WX4666_reg/NET0131 ,
		_w8182_
	);
	LUT2 #(
		.INIT('h8)
	) name6675 (
		RESET_pad,
		\WX9830_reg/NET0131 ,
		_w8183_
	);
	LUT2 #(
		.INIT('h8)
	) name6676 (
		RESET_pad,
		\WX9788_reg/NET0131 ,
		_w8184_
	);
	LUT2 #(
		.INIT('h8)
	) name6677 (
		RESET_pad,
		\WX4674_reg/NET0131 ,
		_w8185_
	);
	LUT2 #(
		.INIT('h8)
	) name6678 (
		RESET_pad,
		\WX9838_reg/NET0131 ,
		_w8186_
	);
	LUT2 #(
		.INIT('h8)
	) name6679 (
		RESET_pad,
		\WX4670_reg/NET0131 ,
		_w8187_
	);
	LUT2 #(
		.INIT('h8)
	) name6680 (
		RESET_pad,
		\WX3253_reg/NET0131 ,
		_w8188_
	);
	LUT2 #(
		.INIT('h8)
	) name6681 (
		RESET_pad,
		\WX4664_reg/NET0131 ,
		_w8189_
	);
	LUT2 #(
		.INIT('h8)
	) name6682 (
		RESET_pad,
		\WX7296_reg/NET0131 ,
		_w8190_
	);
	LUT2 #(
		.INIT('h8)
	) name6683 (
		RESET_pad,
		\WX4660_reg/NET0131 ,
		_w8191_
	);
	LUT2 #(
		.INIT('h8)
	) name6684 (
		RESET_pad,
		\WX9696_reg/NET0131 ,
		_w8192_
	);
	LUT2 #(
		.INIT('h8)
	) name6685 (
		RESET_pad,
		\WX4566_reg/NET0131 ,
		_w8193_
	);
	LUT2 #(
		.INIT('h8)
	) name6686 (
		RESET_pad,
		\WX11001_reg/NET0131 ,
		_w8194_
	);
	LUT2 #(
		.INIT('h8)
	) name6687 (
		RESET_pad,
		\WX9812_reg/NET0131 ,
		_w8195_
	);
	LUT2 #(
		.INIT('h8)
	) name6688 (
		RESET_pad,
		\WX4620_reg/NET0131 ,
		_w8196_
	);
	LUT2 #(
		.INIT('h8)
	) name6689 (
		RESET_pad,
		\WX3407_reg/NET0131 ,
		_w8197_
	);
	LUT2 #(
		.INIT('h8)
	) name6690 (
		RESET_pad,
		\WX821_reg/NET0131 ,
		_w8198_
	);
	LUT2 #(
		.INIT('h8)
	) name6691 (
		RESET_pad,
		\WX8531_reg/NET0131 ,
		_w8199_
	);
	LUT2 #(
		.INIT('h8)
	) name6692 (
		RESET_pad,
		\WX2102_reg/NET0131 ,
		_w8200_
	);
	LUT2 #(
		.INIT('h8)
	) name6693 (
		RESET_pad,
		\WX649_reg/NET0131 ,
		_w8201_
	);
	LUT2 #(
		.INIT('h8)
	) name6694 (
		RESET_pad,
		\WX829_reg/NET0131 ,
		_w8202_
	);
	LUT2 #(
		.INIT('h8)
	) name6695 (
		RESET_pad,
		\WX8555_reg/NET0131 ,
		_w8203_
	);
	LUT2 #(
		.INIT('h8)
	) name6696 (
		RESET_pad,
		\WX3295_reg/NET0131 ,
		_w8204_
	);
	LUT2 #(
		.INIT('h8)
	) name6697 (
		RESET_pad,
		\WX2100_reg/NET0131 ,
		_w8205_
	);
	LUT2 #(
		.INIT('h8)
	) name6698 (
		RESET_pad,
		\WX825_reg/NET0131 ,
		_w8206_
	);
	LUT2 #(
		.INIT('h8)
	) name6699 (
		RESET_pad,
		\WX11017_reg/NET0131 ,
		_w8207_
	);
	LUT2 #(
		.INIT('h8)
	) name6700 (
		RESET_pad,
		\WX5951_reg/NET0131 ,
		_w8208_
	);
	LUT2 #(
		.INIT('h8)
	) name6701 (
		RESET_pad,
		\WX2098_reg/NET0131 ,
		_w8209_
	);
	LUT2 #(
		.INIT('h8)
	) name6702 (
		RESET_pad,
		\WX3297_reg/NET0131 ,
		_w8210_
	);
	LUT2 #(
		.INIT('h8)
	) name6703 (
		RESET_pad,
		\WX5849_reg/NET0131 ,
		_w8211_
	);
	LUT2 #(
		.INIT('h8)
	) name6704 (
		RESET_pad,
		\WX8553_reg/NET0131 ,
		_w8212_
	);
	LUT2 #(
		.INIT('h8)
	) name6705 (
		RESET_pad,
		\WX2016_reg/NET0131 ,
		_w8213_
	);
	LUT2 #(
		.INIT('h8)
	) name6706 (
		RESET_pad,
		\WX11063_reg/NET0131 ,
		_w8214_
	);
	LUT2 #(
		.INIT('h8)
	) name6707 (
		RESET_pad,
		\WX9700_reg/NET0131 ,
		_w8215_
	);
	LUT2 #(
		.INIT('h8)
	) name6708 (
		RESET_pad,
		\WX8463_reg/NET0131 ,
		_w8216_
	);
	LUT2 #(
		.INIT('h8)
	) name6709 (
		RESET_pad,
		\WX2096_reg/NET0131 ,
		_w8217_
	);
	LUT2 #(
		.INIT('h8)
	) name6710 (
		RESET_pad,
		\WX3331_reg/NET0131 ,
		_w8218_
	);
	LUT2 #(
		.INIT('h8)
	) name6711 (
		RESET_pad,
		\WX3299_reg/NET0131 ,
		_w8219_
	);
	LUT2 #(
		.INIT('h8)
	) name6712 (
		RESET_pad,
		\WX8549_reg/NET0131 ,
		_w8220_
	);
	LUT2 #(
		.INIT('h8)
	) name6713 (
		RESET_pad,
		\WX795_reg/NET0131 ,
		_w8221_
	);
	LUT2 #(
		.INIT('h8)
	) name6714 (
		RESET_pad,
		\WX3375_reg/NET0131 ,
		_w8222_
	);
	LUT2 #(
		.INIT('h8)
	) name6715 (
		RESET_pad,
		\WX5859_reg/NET0131 ,
		_w8223_
	);
	LUT2 #(
		.INIT('h8)
	) name6716 (
		RESET_pad,
		\WX4548_reg/NET0131 ,
		_w8224_
	);
	LUT2 #(
		.INIT('h8)
	) name6717 (
		RESET_pad,
		\WX3419_reg/NET0131 ,
		_w8225_
	);
	LUT2 #(
		.INIT('h8)
	) name6718 (
		RESET_pad,
		\WX8545_reg/NET0131 ,
		_w8226_
	);
	LUT2 #(
		.INIT('h8)
	) name6719 (
		RESET_pad,
		\WX4622_reg/NET0131 ,
		_w8227_
	);
	LUT2 #(
		.INIT('h8)
	) name6720 (
		RESET_pad,
		\WX8539_reg/NET0131 ,
		_w8228_
	);
	LUT2 #(
		.INIT('h8)
	) name6721 (
		RESET_pad,
		\WX2094_reg/NET0131 ,
		_w8229_
	);
	LUT2 #(
		.INIT('h8)
	) name6722 (
		RESET_pad,
		\WX2048_reg/NET0131 ,
		_w8230_
	);
	LUT2 #(
		.INIT('h8)
	) name6723 (
		RESET_pad,
		\WX723_reg/NET0131 ,
		_w8231_
	);
	LUT2 #(
		.INIT('h8)
	) name6724 (
		RESET_pad,
		\WX4600_reg/NET0131 ,
		_w8232_
	);
	LUT2 #(
		.INIT('h8)
	) name6725 (
		RESET_pad,
		\WX4602_reg/NET0131 ,
		_w8233_
	);
	LUT2 #(
		.INIT('h8)
	) name6726 (
		RESET_pad,
		\WX8405_reg/NET0131 ,
		_w8234_
	);
	LUT2 #(
		.INIT('h8)
	) name6727 (
		RESET_pad,
		\WX4650_reg/NET0131 ,
		_w8235_
	);
	LUT2 #(
		.INIT('h8)
	) name6728 (
		RESET_pad,
		\WX8543_reg/NET0131 ,
		_w8236_
	);
	LUT2 #(
		.INIT('h8)
	) name6729 (
		RESET_pad,
		\WX10997_reg/NET0131 ,
		_w8237_
	);
	LUT2 #(
		.INIT('h8)
	) name6730 (
		RESET_pad,
		\WX7282_reg/NET0131 ,
		_w8238_
	);
	LUT2 #(
		.INIT('h8)
	) name6731 (
		RESET_pad,
		\WX9884_reg/NET0131 ,
		_w8239_
	);
	LUT2 #(
		.INIT('h8)
	) name6732 (
		RESET_pad,
		\WX5899_reg/NET0131 ,
		_w8240_
	);
	LUT2 #(
		.INIT('h8)
	) name6733 (
		RESET_pad,
		\WX3369_reg/NET0131 ,
		_w8241_
	);
	LUT2 #(
		.INIT('h8)
	) name6734 (
		RESET_pad,
		\WX4616_reg/NET0131 ,
		_w8242_
	);
	LUT2 #(
		.INIT('h8)
	) name6735 (
		RESET_pad,
		\WX8457_reg/NET0131 ,
		_w8243_
	);
	LUT2 #(
		.INIT('h8)
	) name6736 (
		RESET_pad,
		\WX5855_reg/NET0131 ,
		_w8244_
	);
	LUT2 #(
		.INIT('h8)
	) name6737 (
		RESET_pad,
		\WX8435_reg/NET0131 ,
		_w8245_
	);
	LUT2 #(
		.INIT('h8)
	) name6738 (
		RESET_pad,
		\WX759_reg/NET0131 ,
		_w8246_
	);
	LUT2 #(
		.INIT('h8)
	) name6739 (
		RESET_pad,
		\WX8537_reg/NET0131 ,
		_w8247_
	);
	LUT2 #(
		.INIT('h8)
	) name6740 (
		RESET_pad,
		\WX9854_reg/NET0131 ,
		_w8248_
	);
	LUT2 #(
		.INIT('h8)
	) name6741 (
		RESET_pad,
		\WX10999_reg/NET0131 ,
		_w8249_
	);
	LUT2 #(
		.INIT('h8)
	) name6742 (
		RESET_pad,
		\WX7250_reg/NET0131 ,
		_w8250_
	);
	LUT2 #(
		.INIT('h8)
	) name6743 (
		RESET_pad,
		\WX1978_reg/NET0131 ,
		_w8251_
	);
	LUT2 #(
		.INIT('h8)
	) name6744 (
		RESET_pad,
		\WX651_reg/NET0131 ,
		_w8252_
	);
	LUT2 #(
		.INIT('h8)
	) name6745 (
		RESET_pad,
		\WX3387_reg/NET0131 ,
		_w8253_
	);
	LUT2 #(
		.INIT('h8)
	) name6746 (
		RESET_pad,
		\WX681_reg/NET0131 ,
		_w8254_
	);
	LUT2 #(
		.INIT('h8)
	) name6747 (
		RESET_pad,
		\WX8535_reg/NET0131 ,
		_w8255_
	);
	LUT2 #(
		.INIT('h8)
	) name6748 (
		RESET_pad,
		\WX7212_reg/NET0131 ,
		_w8256_
	);
	LUT2 #(
		.INIT('h8)
	) name6749 (
		RESET_pad,
		\WX5981_reg/NET0131 ,
		_w8257_
	);
	LUT2 #(
		.INIT('h8)
	) name6750 (
		RESET_pad,
		\WX4586_reg/NET0131 ,
		_w8258_
	);
	LUT2 #(
		.INIT('h8)
	) name6751 (
		RESET_pad,
		\WX4656_reg/NET0131 ,
		_w8259_
	);
	LUT2 #(
		.INIT('h8)
	) name6752 (
		RESET_pad,
		\WX3333_reg/NET0131 ,
		_w8260_
	);
	LUT2 #(
		.INIT('h8)
	) name6753 (
		RESET_pad,
		\WX9826_reg/NET0131 ,
		_w8261_
	);
	LUT2 #(
		.INIT('h8)
	) name6754 (
		RESET_pad,
		\WX2092_reg/NET0131 ,
		_w8262_
	);
	LUT2 #(
		.INIT('h8)
	) name6755 (
		RESET_pad,
		\WX4624_reg/NET0131 ,
		_w8263_
	);
	LUT2 #(
		.INIT('h8)
	) name6756 (
		RESET_pad,
		\WX7136_reg/NET0131 ,
		_w8264_
	);
	LUT2 #(
		.INIT('h8)
	) name6757 (
		RESET_pad,
		\WX7268_reg/NET0131 ,
		_w8265_
	);
	LUT2 #(
		.INIT('h8)
	) name6758 (
		RESET_pad,
		\WX4642_reg/NET0131 ,
		_w8266_
	);
	LUT2 #(
		.INIT('h8)
	) name6759 (
		RESET_pad,
		\WX8409_reg/NET0131 ,
		_w8267_
	);
	LUT2 #(
		.INIT('h8)
	) name6760 (
		RESET_pad,
		\WX4618_reg/NET0131 ,
		_w8268_
	);
	LUT2 #(
		.INIT('h8)
	) name6761 (
		RESET_pad,
		\WX4612_reg/NET0131 ,
		_w8269_
	);
	LUT2 #(
		.INIT('h8)
	) name6762 (
		RESET_pad,
		\WX7292_reg/NET0131 ,
		_w8270_
	);
	LUT2 #(
		.INIT('h8)
	) name6763 (
		RESET_pad,
		\WX3231_reg/NET0131 ,
		_w8271_
	);
	LUT2 #(
		.INIT('h8)
	) name6764 (
		RESET_pad,
		\WX8489_reg/NET0131 ,
		_w8272_
	);
	LUT2 #(
		.INIT('h8)
	) name6765 (
		RESET_pad,
		\WX3305_reg/NET0131 ,
		_w8273_
	);
	LUT2 #(
		.INIT('h8)
	) name6766 (
		RESET_pad,
		\WX8525_reg/NET0131 ,
		_w8274_
	);
	LUT2 #(
		.INIT('h8)
	) name6767 (
		RESET_pad,
		\WX11159_reg/NET0131 ,
		_w8275_
	);
	LUT2 #(
		.INIT('h8)
	) name6768 (
		RESET_pad,
		\WX3367_reg/NET0131 ,
		_w8276_
	);
	LUT2 #(
		.INIT('h8)
	) name6769 (
		RESET_pad,
		\WX11061_reg/NET0131 ,
		_w8277_
	);
	LUT2 #(
		.INIT('h8)
	) name6770 (
		RESET_pad,
		\WX8569_reg/NET0131 ,
		_w8278_
	);
	LUT2 #(
		.INIT('h8)
	) name6771 (
		RESET_pad,
		\WX11125_reg/NET0131 ,
		_w8279_
	);
	LUT2 #(
		.INIT('h8)
	) name6772 (
		RESET_pad,
		\WX809_reg/NET0131 ,
		_w8280_
	);
	LUT2 #(
		.INIT('h8)
	) name6773 (
		RESET_pad,
		\WX683_reg/NET0131 ,
		_w8281_
	);
	LUT2 #(
		.INIT('h8)
	) name6774 (
		RESET_pad,
		\WX8413_reg/NET0131 ,
		_w8282_
	);
	LUT2 #(
		.INIT('h8)
	) name6775 (
		RESET_pad,
		\WX2062_reg/NET0131 ,
		_w8283_
	);
	LUT2 #(
		.INIT('h8)
	) name6776 (
		RESET_pad,
		\WX9758_reg/NET0131 ,
		_w8284_
	);
	LUT2 #(
		.INIT('h8)
	) name6777 (
		RESET_pad,
		\WX3397_reg/NET0131 ,
		_w8285_
	);
	LUT2 #(
		.INIT('h8)
	) name6778 (
		RESET_pad,
		\WX7300_reg/NET0131 ,
		_w8286_
	);
	LUT2 #(
		.INIT('h8)
	) name6779 (
		RESET_pad,
		\WX6003_reg/NET0131 ,
		_w8287_
	);
	LUT2 #(
		.INIT('h8)
	) name6780 (
		RESET_pad,
		\WX4646_reg/NET0131 ,
		_w8288_
	);
	LUT2 #(
		.INIT('h8)
	) name6781 (
		RESET_pad,
		\WX9880_reg/NET0131 ,
		_w8289_
	);
	LUT2 #(
		.INIT('h8)
	) name6782 (
		RESET_pad,
		\WX7258_reg/NET0131 ,
		_w8290_
	);
	LUT2 #(
		.INIT('h8)
	) name6783 (
		RESET_pad,
		\WX8593_reg/NET0131 ,
		_w8291_
	);
	LUT2 #(
		.INIT('h8)
	) name6784 (
		RESET_pad,
		\WX11057_reg/NET0131 ,
		_w8292_
	);
	LUT2 #(
		.INIT('h8)
	) name6785 (
		RESET_pad,
		\WX675_reg/NET0131 ,
		_w8293_
	);
	LUT2 #(
		.INIT('h8)
	) name6786 (
		RESET_pad,
		\WX3371_reg/NET0131 ,
		_w8294_
	);
	LUT2 #(
		.INIT('h8)
	) name6787 (
		RESET_pad,
		\WX783_reg/NET0131 ,
		_w8295_
	);
	LUT2 #(
		.INIT('h8)
	) name6788 (
		RESET_pad,
		\WX8411_reg/NET0131 ,
		_w8296_
	);
	LUT2 #(
		.INIT('h8)
	) name6789 (
		RESET_pad,
		\WX9836_reg/NET0131 ,
		_w8297_
	);
	LUT2 #(
		.INIT('h8)
	) name6790 (
		RESET_pad,
		\WX11055_reg/NET0131 ,
		_w8298_
	);
	LUT2 #(
		.INIT('h8)
	) name6791 (
		RESET_pad,
		\WX8467_reg/NET0131 ,
		_w8299_
	);
	LUT2 #(
		.INIT('h8)
	) name6792 (
		RESET_pad,
		\WX817_reg/NET0131 ,
		_w8300_
	);
	LUT2 #(
		.INIT('h8)
	) name6793 (
		RESET_pad,
		\WX9870_reg/NET0131 ,
		_w8301_
	);
	LUT2 #(
		.INIT('h8)
	) name6794 (
		RESET_pad,
		\WX7262_reg/NET0131 ,
		_w8302_
	);
	LUT2 #(
		.INIT('h8)
	) name6795 (
		RESET_pad,
		\WX7264_reg/NET0131 ,
		_w8303_
	);
	LUT2 #(
		.INIT('h8)
	) name6796 (
		RESET_pad,
		\WX4604_reg/NET0131 ,
		_w8304_
	);
	LUT2 #(
		.INIT('h8)
	) name6797 (
		RESET_pad,
		\WX9804_reg/NET0131 ,
		_w8305_
	);
	LUT2 #(
		.INIT('h8)
	) name6798 (
		RESET_pad,
		\WX8429_reg/NET0131 ,
		_w8306_
	);
	LUT2 #(
		.INIT('h8)
	) name6799 (
		RESET_pad,
		\WX815_reg/NET0131 ,
		_w8307_
	);
	LUT2 #(
		.INIT('h8)
	) name6800 (
		RESET_pad,
		\WX5877_reg/NET0131 ,
		_w8308_
	);
	LUT2 #(
		.INIT('h8)
	) name6801 (
		RESET_pad,
		\WX6001_reg/NET0131 ,
		_w8309_
	);
	LUT2 #(
		.INIT('h8)
	) name6802 (
		RESET_pad,
		\WX8521_reg/NET0131 ,
		_w8310_
	);
	LUT2 #(
		.INIT('h8)
	) name6803 (
		RESET_pad,
		\WX7270_reg/NET0131 ,
		_w8311_
	);
	LUT2 #(
		.INIT('h8)
	) name6804 (
		RESET_pad,
		\WX677_reg/NET0131 ,
		_w8312_
	);
	LUT2 #(
		.INIT('h8)
	) name6805 (
		RESET_pad,
		\WX5989_reg/NET0131 ,
		_w8313_
	);
	LUT2 #(
		.INIT('h8)
	) name6806 (
		RESET_pad,
		\WX5993_reg/NET0131 ,
		_w8314_
	);
	LUT2 #(
		.INIT('h8)
	) name6807 (
		RESET_pad,
		\WX3303_reg/NET0131 ,
		_w8315_
	);
	LUT2 #(
		.INIT('h8)
	) name6808 (
		RESET_pad,
		\WX7142_reg/NET0131 ,
		_w8316_
	);
	LUT2 #(
		.INIT('h8)
	) name6809 (
		RESET_pad,
		\WX793_reg/NET0131 ,
		_w8317_
	);
	LUT2 #(
		.INIT('h8)
	) name6810 (
		RESET_pad,
		\WX9756_reg/NET0131 ,
		_w8318_
	);
	LUT2 #(
		.INIT('h8)
	) name6811 (
		RESET_pad,
		\WX7260_reg/NET0131 ,
		_w8319_
	);
	LUT2 #(
		.INIT('h8)
	) name6812 (
		RESET_pad,
		\WX5903_reg/NET0131 ,
		_w8320_
	);
	LUT2 #(
		.INIT('h8)
	) name6813 (
		RESET_pad,
		\WX11065_reg/NET0131 ,
		_w8321_
	);
	LUT2 #(
		.INIT('h8)
	) name6814 (
		RESET_pad,
		\WX4534_reg/NET0131 ,
		_w8322_
	);
	LUT2 #(
		.INIT('h8)
	) name6815 (
		RESET_pad,
		\WX4546_reg/NET0131 ,
		_w8323_
	);
	LUT2 #(
		.INIT('h8)
	) name6816 (
		RESET_pad,
		\WX2074_reg/NET0131 ,
		_w8324_
	);
	LUT2 #(
		.INIT('h8)
	) name6817 (
		RESET_pad,
		\WX8483_reg/NET0131 ,
		_w8325_
	);
	LUT2 #(
		.INIT('h8)
	) name6818 (
		RESET_pad,
		\WX3307_reg/NET0131 ,
		_w8326_
	);
	LUT2 #(
		.INIT('h8)
	) name6819 (
		RESET_pad,
		\WX9866_reg/NET0131 ,
		_w8327_
	);
	LUT2 #(
		.INIT('h8)
	) name6820 (
		RESET_pad,
		\WX4610_reg/NET0131 ,
		_w8328_
	);
	LUT2 #(
		.INIT('h8)
	) name6821 (
		RESET_pad,
		\WX4582_reg/NET0131 ,
		_w8329_
	);
	LUT2 #(
		.INIT('h8)
	) name6822 (
		RESET_pad,
		\WX5987_reg/NET0131 ,
		_w8330_
	);
	LUT2 #(
		.INIT('h8)
	) name6823 (
		RESET_pad,
		\WX11051_reg/NET0131 ,
		_w8331_
	);
	LUT2 #(
		.INIT('h8)
	) name6824 (
		RESET_pad,
		\WX4640_reg/NET0131 ,
		_w8332_
	);
	LUT2 #(
		.INIT('h8)
	) name6825 (
		RESET_pad,
		\WX655_reg/NET0131 ,
		_w8333_
	);
	LUT2 #(
		.INIT('h8)
	) name6826 (
		RESET_pad,
		\WX4596_reg/NET0131 ,
		_w8334_
	);
	LUT2 #(
		.INIT('h8)
	) name6827 (
		RESET_pad,
		\WX673_reg/NET0131 ,
		_w8335_
	);
	LUT2 #(
		.INIT('h8)
	) name6828 (
		RESET_pad,
		\WX4592_reg/NET0131 ,
		_w8336_
	);
	LUT2 #(
		.INIT('h8)
	) name6829 (
		RESET_pad,
		\WX7298_reg/NET0131 ,
		_w8337_
	);
	LUT2 #(
		.INIT('h8)
	) name6830 (
		RESET_pad,
		\WX2078_reg/NET0131 ,
		_w8338_
	);
	LUT2 #(
		.INIT('h8)
	) name6831 (
		RESET_pad,
		\WX2038_reg/NET0131 ,
		_w8339_
	);
	LUT2 #(
		.INIT('h8)
	) name6832 (
		RESET_pad,
		\WX11003_reg/NET0131 ,
		_w8340_
	);
	LUT2 #(
		.INIT('h8)
	) name6833 (
		RESET_pad,
		\WX5881_reg/NET0131 ,
		_w8341_
	);
	LUT2 #(
		.INIT('h8)
	) name6834 (
		RESET_pad,
		\WX4644_reg/NET0131 ,
		_w8342_
	);
	LUT2 #(
		.INIT('h8)
	) name6835 (
		RESET_pad,
		\WX2120_reg/NET0131 ,
		_w8343_
	);
	LUT2 #(
		.INIT('h8)
	) name6836 (
		RESET_pad,
		\WX4654_reg/NET0131 ,
		_w8344_
	);
	LUT2 #(
		.INIT('h8)
	) name6837 (
		RESET_pad,
		\WX3353_reg/NET0131 ,
		_w8345_
	);
	LUT2 #(
		.INIT('h8)
	) name6838 (
		RESET_pad,
		\WX5983_reg/NET0131 ,
		_w8346_
	);
	LUT2 #(
		.INIT('h8)
	) name6839 (
		RESET_pad,
		\WX4572_reg/NET0131 ,
		_w8347_
	);
	LUT2 #(
		.INIT('h8)
	) name6840 (
		RESET_pad,
		\WX8427_reg/NET0131 ,
		_w8348_
	);
	LUT2 #(
		.INIT('h8)
	) name6841 (
		RESET_pad,
		\WX4684_reg/NET0131 ,
		_w8349_
	);
	LUT2 #(
		.INIT('h8)
	) name6842 (
		RESET_pad,
		\WX4694_reg/NET0131 ,
		_w8350_
	);
	LUT2 #(
		.INIT('h8)
	) name6843 (
		RESET_pad,
		\WX833_reg/NET0131 ,
		_w8351_
	);
	LUT2 #(
		.INIT('h8)
	) name6844 (
		RESET_pad,
		\WX9886_reg/NET0131 ,
		_w8352_
	);
	LUT2 #(
		.INIT('h8)
	) name6845 (
		RESET_pad,
		\WX4552_reg/NET0131 ,
		_w8353_
	);
	LUT2 #(
		.INIT('h8)
	) name6846 (
		RESET_pad,
		\WX4606_reg/NET0131 ,
		_w8354_
	);
	LUT2 #(
		.INIT('h8)
	) name6847 (
		RESET_pad,
		\WX4536_reg/NET0131 ,
		_w8355_
	);
	LUT2 #(
		.INIT('h8)
	) name6848 (
		RESET_pad,
		\WX7140_reg/NET0131 ,
		_w8356_
	);
	LUT2 #(
		.INIT('h8)
	) name6849 (
		RESET_pad,
		\WX5975_reg/NET0131 ,
		_w8357_
	);
	LUT2 #(
		.INIT('h8)
	) name6850 (
		RESET_pad,
		\WX2110_reg/NET0131 ,
		_w8358_
	);
	LUT2 #(
		.INIT('h8)
	) name6851 (
		RESET_pad,
		\WX7274_reg/NET0131 ,
		_w8359_
	);
	LUT2 #(
		.INIT('h8)
	) name6852 (
		RESET_pad,
		\WX5977_reg/NET0131 ,
		_w8360_
	);
	LUT2 #(
		.INIT('h8)
	) name6853 (
		RESET_pad,
		\WX3417_reg/NET0131 ,
		_w8361_
	);
	LUT2 #(
		.INIT('h8)
	) name6854 (
		RESET_pad,
		\WX8507_reg/NET0131 ,
		_w8362_
	);
	LUT2 #(
		.INIT('h8)
	) name6855 (
		RESET_pad,
		\WX9720_reg/NET0131 ,
		_w8363_
	);
	LUT2 #(
		.INIT('h8)
	) name6856 (
		RESET_pad,
		\WX5971_reg/NET0131 ,
		_w8364_
	);
	LUT2 #(
		.INIT('h8)
	) name6857 (
		RESET_pad,
		\WX5967_reg/NET0131 ,
		_w8365_
	);
	LUT2 #(
		.INIT('h8)
	) name6858 (
		RESET_pad,
		\WX7146_reg/NET0131 ,
		_w8366_
	);
	LUT2 #(
		.INIT('h8)
	) name6859 (
		RESET_pad,
		\WX8541_reg/NET0131 ,
		_w8367_
	);
	LUT2 #(
		.INIT('h8)
	) name6860 (
		RESET_pad,
		\WX5969_reg/NET0131 ,
		_w8368_
	);
	LUT2 #(
		.INIT('h8)
	) name6861 (
		RESET_pad,
		\WX3373_reg/NET0131 ,
		_w8369_
	);
	LUT2 #(
		.INIT('h8)
	) name6862 (
		RESET_pad,
		\WX5963_reg/NET0131 ,
		_w8370_
	);
	LUT2 #(
		.INIT('h8)
	) name6863 (
		RESET_pad,
		\WX8513_reg/NET0131 ,
		_w8371_
	);
	LUT2 #(
		.INIT('h8)
	) name6864 (
		RESET_pad,
		\WX8509_reg/NET0131 ,
		_w8372_
	);
	LUT2 #(
		.INIT('h8)
	) name6865 (
		RESET_pad,
		\WX8433_reg/NET0131 ,
		_w8373_
	);
	LUT2 #(
		.INIT('h8)
	) name6866 (
		RESET_pad,
		\WX11047_reg/NET0131 ,
		_w8374_
	);
	LUT2 #(
		.INIT('h8)
	) name6867 (
		RESET_pad,
		\WX1942_reg/NET0131 ,
		_w8375_
	);
	LUT2 #(
		.INIT('h8)
	) name6868 (
		RESET_pad,
		\WX5961_reg/NET0131 ,
		_w8376_
	);
	LUT2 #(
		.INIT('h8)
	) name6869 (
		RESET_pad,
		\WX8511_reg/NET0131 ,
		_w8377_
	);
	LUT2 #(
		.INIT('h8)
	) name6870 (
		RESET_pad,
		\WX8431_reg/NET0131 ,
		_w8378_
	);
	LUT2 #(
		.INIT('h8)
	) name6871 (
		RESET_pad,
		\WX7286_reg/NET0131 ,
		_w8379_
	);
	LUT2 #(
		.INIT('h8)
	) name6872 (
		RESET_pad,
		\WX7288_reg/NET0131 ,
		_w8380_
	);
	LUT2 #(
		.INIT('h8)
	) name6873 (
		RESET_pad,
		\WX3343_reg/NET0131 ,
		_w8381_
	);
	LUT2 #(
		.INIT('h8)
	) name6874 (
		RESET_pad,
		\WX7112_reg/NET0131 ,
		_w8382_
	);
	LUT2 #(
		.INIT('h8)
	) name6875 (
		RESET_pad,
		\WX9766_reg/NET0131 ,
		_w8383_
	);
	LUT2 #(
		.INIT('h8)
	) name6876 (
		RESET_pad,
		\WX3315_reg/NET0131 ,
		_w8384_
	);
	LUT2 #(
		.INIT('h8)
	) name6877 (
		RESET_pad,
		\WX2070_reg/NET0131 ,
		_w8385_
	);
	LUT2 #(
		.INIT('h8)
	) name6878 (
		RESET_pad,
		\WX11091_reg/NET0131 ,
		_w8386_
	);
	LUT2 #(
		.INIT('h8)
	) name6879 (
		RESET_pad,
		\WX3377_reg/NET0131 ,
		_w8387_
	);
	LUT2 #(
		.INIT('h8)
	) name6880 (
		RESET_pad,
		\WX5943_reg/NET0131 ,
		_w8388_
	);
	LUT2 #(
		.INIT('h8)
	) name6881 (
		RESET_pad,
		\WX8479_reg/NET0131 ,
		_w8389_
	);
	LUT2 #(
		.INIT('h8)
	) name6882 (
		RESET_pad,
		\WX1948_reg/NET0131 ,
		_w8390_
	);
	LUT2 #(
		.INIT('h8)
	) name6883 (
		RESET_pad,
		\WX747_reg/NET0131 ,
		_w8391_
	);
	LUT2 #(
		.INIT('h8)
	) name6884 (
		RESET_pad,
		\WX8439_reg/NET0131 ,
		_w8392_
	);
	LUT2 #(
		.INIT('h8)
	) name6885 (
		RESET_pad,
		\WX9738_reg/NET0131 ,
		_w8393_
	);
	LUT2 #(
		.INIT('h8)
	) name6886 (
		RESET_pad,
		\WX9858_reg/NET0131 ,
		_w8394_
	);
	LUT2 #(
		.INIT('h8)
	) name6887 (
		RESET_pad,
		\WX7216_reg/NET0131 ,
		_w8395_
	);
	LUT2 #(
		.INIT('h8)
	) name6888 (
		RESET_pad,
		\WX2022_reg/NET0131 ,
		_w8396_
	);
	LUT2 #(
		.INIT('h8)
	) name6889 (
		RESET_pad,
		\WX4702_reg/NET0131 ,
		_w8397_
	);
	LUT2 #(
		.INIT('h8)
	) name6890 (
		RESET_pad,
		\WX4524_reg/NET0131 ,
		_w8398_
	);
	LUT2 #(
		.INIT('h8)
	) name6891 (
		RESET_pad,
		\WX5853_reg/NET0131 ,
		_w8399_
	);
	LUT2 #(
		.INIT('h8)
	) name6892 (
		RESET_pad,
		\WX5889_reg/NET0131 ,
		_w8400_
	);
	LUT2 #(
		.INIT('h8)
	) name6893 (
		RESET_pad,
		\WX8477_reg/NET0131 ,
		_w8401_
	);
	LUT2 #(
		.INIT('h8)
	) name6894 (
		RESET_pad,
		\WX4608_reg/NET0131 ,
		_w8402_
	);
	LUT2 #(
		.INIT('h8)
	) name6895 (
		RESET_pad,
		\WX5915_reg/NET0131 ,
		_w8403_
	);
	LUT2 #(
		.INIT('h8)
	) name6896 (
		RESET_pad,
		\WX8495_reg/NET0131 ,
		_w8404_
	);
	LUT2 #(
		.INIT('h8)
	) name6897 (
		RESET_pad,
		\WX3313_reg/NET0131 ,
		_w8405_
	);
	LUT2 #(
		.INIT('h8)
	) name6898 (
		RESET_pad,
		\WX8437_reg/NET0131 ,
		_w8406_
	);
	LUT2 #(
		.INIT('h8)
	) name6899 (
		RESET_pad,
		\WX5935_reg/NET0131 ,
		_w8407_
	);
	LUT2 #(
		.INIT('h8)
	) name6900 (
		RESET_pad,
		\WX715_reg/NET0131 ,
		_w8408_
	);
	LUT2 #(
		.INIT('h8)
	) name6901 (
		RESET_pad,
		\WX8501_reg/NET0131 ,
		_w8409_
	);
	LUT2 #(
		.INIT('h8)
	) name6902 (
		RESET_pad,
		\WX11009_reg/NET0131 ,
		_w8410_
	);
	LUT2 #(
		.INIT('h8)
	) name6903 (
		RESET_pad,
		\WX5931_reg/NET0131 ,
		_w8411_
	);
	LUT2 #(
		.INIT('h8)
	) name6904 (
		RESET_pad,
		\WX4590_reg/NET0131 ,
		_w8412_
	);
	LUT2 #(
		.INIT('h8)
	) name6905 (
		RESET_pad,
		\WX2124_reg/NET0131 ,
		_w8413_
	);
	LUT2 #(
		.INIT('h8)
	) name6906 (
		RESET_pad,
		\WX775_reg/NET0131 ,
		_w8414_
	);
	LUT2 #(
		.INIT('h8)
	) name6907 (
		RESET_pad,
		\WX9792_reg/NET0131 ,
		_w8415_
	);
	LUT2 #(
		.INIT('h8)
	) name6908 (
		RESET_pad,
		\WX811_reg/NET0131 ,
		_w8416_
	);
	LUT2 #(
		.INIT('h8)
	) name6909 (
		RESET_pad,
		\WX8499_reg/NET0131 ,
		_w8417_
	);
	LUT2 #(
		.INIT('h8)
	) name6910 (
		RESET_pad,
		\WX10991_reg/NET0131 ,
		_w8418_
	);
	LUT2 #(
		.INIT('h8)
	) name6911 (
		RESET_pad,
		\WX7162_reg/NET0131 ,
		_w8419_
	);
	LUT2 #(
		.INIT('h8)
	) name6912 (
		RESET_pad,
		\WX3411_reg/NET0131 ,
		_w8420_
	);
	LUT2 #(
		.INIT('h8)
	) name6913 (
		RESET_pad,
		\WX8497_reg/NET0131 ,
		_w8421_
	);
	LUT2 #(
		.INIT('h8)
	) name6914 (
		RESET_pad,
		\WX703_reg/NET0131 ,
		_w8422_
	);
	LUT2 #(
		.INIT('h8)
	) name6915 (
		RESET_pad,
		\WX5917_reg/NET0131 ,
		_w8423_
	);
	LUT2 #(
		.INIT('h8)
	) name6916 (
		RESET_pad,
		\WX11157_reg/NET0131 ,
		_w8424_
	);
	LUT2 #(
		.INIT('h8)
	) name6917 (
		RESET_pad,
		\WX1970_reg/NET0131 ,
		_w8425_
	);
	LUT2 #(
		.INIT('h8)
	) name6918 (
		RESET_pad,
		\WX1974_reg/NET0131 ,
		_w8426_
	);
	LUT2 #(
		.INIT('h8)
	) name6919 (
		RESET_pad,
		\WX8493_reg/NET0131 ,
		_w8427_
	);
	LUT2 #(
		.INIT('h8)
	) name6920 (
		RESET_pad,
		\WX9828_reg/NET0131 ,
		_w8428_
	);
	LUT2 #(
		.INIT('h8)
	) name6921 (
		RESET_pad,
		\WX5911_reg/NET0131 ,
		_w8429_
	);
	LUT2 #(
		.INIT('h8)
	) name6922 (
		RESET_pad,
		\WX797_reg/NET0131 ,
		_w8430_
	);
	LUT2 #(
		.INIT('h8)
	) name6923 (
		RESET_pad,
		\WX1962_reg/NET0131 ,
		_w8431_
	);
	LUT2 #(
		.INIT('h8)
	) name6924 (
		RESET_pad,
		\WX2040_reg/NET0131 ,
		_w8432_
	);
	LUT2 #(
		.INIT('h8)
	) name6925 (
		RESET_pad,
		\WX827_reg/NET0131 ,
		_w8433_
	);
	LUT2 #(
		.INIT('h8)
	) name6926 (
		RESET_pad,
		\WX8487_reg/NET0131 ,
		_w8434_
	);
	LUT2 #(
		.INIT('h8)
	) name6927 (
		RESET_pad,
		\WX5913_reg/NET0131 ,
		_w8435_
	);
	LUT2 #(
		.INIT('h8)
	) name6928 (
		RESET_pad,
		\WX1952_reg/NET0131 ,
		_w8436_
	);
	LUT2 #(
		.INIT('h8)
	) name6929 (
		RESET_pad,
		\WX5905_reg/NET0131 ,
		_w8437_
	);
	LUT2 #(
		.INIT('h8)
	) name6930 (
		RESET_pad,
		\WX3345_reg/NET0131 ,
		_w8438_
	);
	LUT2 #(
		.INIT('h8)
	) name6931 (
		RESET_pad,
		\WX9748_reg/NET0131 ,
		_w8439_
	);
	LUT2 #(
		.INIT('h8)
	) name6932 (
		RESET_pad,
		\WX2058_reg/NET0131 ,
		_w8440_
	);
	LUT2 #(
		.INIT('h8)
	) name6933 (
		RESET_pad,
		\WX5907_reg/NET0131 ,
		_w8441_
	);
	LUT2 #(
		.INIT('h8)
	) name6934 (
		RESET_pad,
		\WX3249_reg/NET0131 ,
		_w8442_
	);
	LUT2 #(
		.INIT('h8)
	) name6935 (
		RESET_pad,
		\WX1944_reg/NET0131 ,
		_w8443_
	);
	LUT2 #(
		.INIT('h8)
	) name6936 (
		RESET_pad,
		\WX4630_reg/NET0131 ,
		_w8444_
	);
	LUT2 #(
		.INIT('h8)
	) name6937 (
		RESET_pad,
		\WX5895_reg/NET0131 ,
		_w8445_
	);
	LUT2 #(
		.INIT('h8)
	) name6938 (
		RESET_pad,
		\WX5887_reg/NET0131 ,
		_w8446_
	);
	LUT2 #(
		.INIT('h8)
	) name6939 (
		RESET_pad,
		\WX1938_reg/NET0131 ,
		_w8447_
	);
	LUT2 #(
		.INIT('h8)
	) name6940 (
		RESET_pad,
		\WX1940_reg/NET0131 ,
		_w8448_
	);
	LUT2 #(
		.INIT('h8)
	) name6941 (
		RESET_pad,
		\WX8403_reg/NET0131 ,
		_w8449_
	);
	LUT2 #(
		.INIT('h8)
	) name6942 (
		RESET_pad,
		\WX725_reg/NET0131 ,
		_w8450_
	);
	LUT2 #(
		.INIT('h8)
	) name6943 (
		RESET_pad,
		\WX5897_reg/NET0131 ,
		_w8451_
	);
	LUT2 #(
		.INIT('h8)
	) name6944 (
		RESET_pad,
		\WX11173_reg/NET0131 ,
		_w8452_
	);
	LUT2 #(
		.INIT('h8)
	) name6945 (
		RESET_pad,
		\WX8425_reg/NET0131 ,
		_w8453_
	);
	LUT2 #(
		.INIT('h8)
	) name6946 (
		RESET_pad,
		\WX7170_reg/NET0131 ,
		_w8454_
	);
	LUT2 #(
		.INIT('h8)
	) name6947 (
		RESET_pad,
		\WX8465_reg/NET0131 ,
		_w8455_
	);
	LUT2 #(
		.INIT('h8)
	) name6948 (
		RESET_pad,
		\WX4530_reg/NET0131 ,
		_w8456_
	);
	LUT2 #(
		.INIT('h8)
	) name6949 (
		RESET_pad,
		\WX7172_reg/NET0131 ,
		_w8457_
	);
	LUT2 #(
		.INIT('h8)
	) name6950 (
		RESET_pad,
		\WX5893_reg/NET0131 ,
		_w8458_
	);
	LUT2 #(
		.INIT('h8)
	) name6951 (
		RESET_pad,
		\WX785_reg/NET0131 ,
		_w8459_
	);
	LUT2 #(
		.INIT('h8)
	) name6952 (
		RESET_pad,
		\WX2050_reg/NET0131 ,
		_w8460_
	);
	LUT2 #(
		.INIT('h8)
	) name6953 (
		RESET_pad,
		\WX8585_reg/NET0131 ,
		_w8461_
	);
	LUT2 #(
		.INIT('h8)
	) name6954 (
		RESET_pad,
		\WX8587_reg/NET0131 ,
		_w8462_
	);
	LUT2 #(
		.INIT('h8)
	) name6955 (
		RESET_pad,
		\WX5891_reg/NET0131 ,
		_w8463_
	);
	LUT2 #(
		.INIT('h8)
	) name6956 (
		RESET_pad,
		\WX671_reg/NET0131 ,
		_w8464_
	);
	LUT2 #(
		.INIT('h8)
	) name6957 (
		RESET_pad,
		\WX2028_reg/NET0131 ,
		_w8465_
	);
	LUT2 #(
		.INIT('h8)
	) name6958 (
		RESET_pad,
		\WX11097_reg/NET0131 ,
		_w8466_
	);
	LUT2 #(
		.INIT('h8)
	) name6959 (
		RESET_pad,
		\WX2116_reg/NET0131 ,
		_w8467_
	);
	LUT2 #(
		.INIT('h8)
	) name6960 (
		RESET_pad,
		\WX11151_reg/NET0131 ,
		_w8468_
	);
	LUT2 #(
		.INIT('h8)
	) name6961 (
		RESET_pad,
		\WX679_reg/NET0131 ,
		_w8469_
	);
	LUT2 #(
		.INIT('h8)
	) name6962 (
		RESET_pad,
		\WX2024_reg/NET0131 ,
		_w8470_
	);
	LUT2 #(
		.INIT('h8)
	) name6963 (
		RESET_pad,
		\WX4706_reg/NET0131 ,
		_w8471_
	);
	LUT2 #(
		.INIT('h8)
	) name6964 (
		RESET_pad,
		\WX7168_reg/NET0131 ,
		_w8472_
	);
	LUT2 #(
		.INIT('h8)
	) name6965 (
		RESET_pad,
		\WX4554_reg/NET0131 ,
		_w8473_
	);
	LUT2 #(
		.INIT('h8)
	) name6966 (
		RESET_pad,
		\WX8421_reg/NET0131 ,
		_w8474_
	);
	LUT2 #(
		.INIT('h8)
	) name6967 (
		RESET_pad,
		\WX2090_reg/NET0131 ,
		_w8475_
	);
	LUT2 #(
		.INIT('h8)
	) name6968 (
		RESET_pad,
		\WX9784_reg/NET0131 ,
		_w8476_
	);
	LUT2 #(
		.INIT('h8)
	) name6969 (
		RESET_pad,
		\WX4714_reg/NET0131 ,
		_w8477_
	);
	LUT2 #(
		.INIT('h8)
	) name6970 (
		RESET_pad,
		\WX11013_reg/NET0131 ,
		_w8478_
	);
	LUT2 #(
		.INIT('h8)
	) name6971 (
		RESET_pad,
		\WX2052_reg/NET0131 ,
		_w8479_
	);
	LUT2 #(
		.INIT('h8)
	) name6972 (
		RESET_pad,
		\WX8417_reg/NET0131 ,
		_w8480_
	);
	LUT2 #(
		.INIT('h8)
	) name6973 (
		RESET_pad,
		\WX3341_reg/NET0131 ,
		_w8481_
	);
	LUT2 #(
		.INIT('h8)
	) name6974 (
		RESET_pad,
		\WX5883_reg/NET0131 ,
		_w8482_
	);
	LUT2 #(
		.INIT('h8)
	) name6975 (
		RESET_pad,
		\WX3323_reg/NET0131 ,
		_w8483_
	);
	LUT2 #(
		.INIT('h8)
	) name6976 (
		RESET_pad,
		\WX9868_reg/NET0131 ,
		_w8484_
	);
	LUT2 #(
		.INIT('h8)
	) name6977 (
		RESET_pad,
		\WX8461_reg/NET0131 ,
		_w8485_
	);
	LUT2 #(
		.INIT('h8)
	) name6978 (
		RESET_pad,
		\WX3329_reg/NET0131 ,
		_w8486_
	);
	LUT2 #(
		.INIT('h8)
	) name6979 (
		RESET_pad,
		\WX11171_reg/NET0131 ,
		_w8487_
	);
	LUT2 #(
		.INIT('h8)
	) name6980 (
		RESET_pad,
		\WX9734_reg/NET0131 ,
		_w8488_
	);
	LUT2 #(
		.INIT('h8)
	) name6981 (
		RESET_pad,
		\WX7176_reg/NET0131 ,
		_w8489_
	);
	LUT2 #(
		.INIT('h8)
	) name6982 (
		RESET_pad,
		\WX2018_reg/NET0131 ,
		_w8490_
	);
	LUT2 #(
		.INIT('h8)
	) name6983 (
		RESET_pad,
		\WX9834_reg/NET0131 ,
		_w8491_
	);
	LUT2 #(
		.INIT('h8)
	) name6984 (
		RESET_pad,
		\WX3401_reg/NET0131 ,
		_w8492_
	);
	LUT2 #(
		.INIT('h8)
	) name6985 (
		RESET_pad,
		\WX2006_reg/NET0131 ,
		_w8493_
	);
	LUT2 #(
		.INIT('h8)
	) name6986 (
		RESET_pad,
		\WX3337_reg/NET0131 ,
		_w8494_
	);
	LUT2 #(
		.INIT('h8)
	) name6987 (
		RESET_pad,
		\WX8503_reg/NET0131 ,
		_w8495_
	);
	LUT2 #(
		.INIT('h8)
	) name6988 (
		RESET_pad,
		\WX5867_reg/NET0131 ,
		_w8496_
	);
	LUT2 #(
		.INIT('h8)
	) name6989 (
		RESET_pad,
		\WX6005_reg/NET0131 ,
		_w8497_
	);
	LUT2 #(
		.INIT('h8)
	) name6990 (
		RESET_pad,
		\WX11025_reg/NET0131 ,
		_w8498_
	);
	LUT2 #(
		.INIT('h8)
	) name6991 (
		RESET_pad,
		\WX1990_reg/NET0131 ,
		_w8499_
	);
	LUT2 #(
		.INIT('h8)
	) name6992 (
		RESET_pad,
		\WX5831_reg/NET0131 ,
		_w8500_
	);
	LUT2 #(
		.INIT('h8)
	) name6993 (
		RESET_pad,
		\WX5955_reg/NET0131 ,
		_w8501_
	);
	LUT2 #(
		.INIT('h8)
	) name6994 (
		RESET_pad,
		\WX8523_reg/NET0131 ,
		_w8502_
	);
	LUT2 #(
		.INIT('h8)
	) name6995 (
		RESET_pad,
		\WX2084_reg/NET0131 ,
		_w8503_
	);
	LUT2 #(
		.INIT('h8)
	) name6996 (
		RESET_pad,
		\WX789_reg/NET0131 ,
		_w8504_
	);
	LUT2 #(
		.INIT('h8)
	) name6997 (
		RESET_pad,
		\WX3381_reg/NET0131 ,
		_w8505_
	);
	LUT2 #(
		.INIT('h8)
	) name6998 (
		RESET_pad,
		\WX5865_reg/NET0131 ,
		_w8506_
	);
	LUT2 #(
		.INIT('h8)
	) name6999 (
		RESET_pad,
		\WX5885_reg/NET0131 ,
		_w8507_
	);
	LUT2 #(
		.INIT('h8)
	) name7000 (
		RESET_pad,
		\WX9794_reg/NET0131 ,
		_w8508_
	);
	LUT2 #(
		.INIT('h8)
	) name7001 (
		RESET_pad,
		\WX5819_reg/NET0131 ,
		_w8509_
	);
	LUT2 #(
		.INIT('h8)
	) name7002 (
		RESET_pad,
		\WX5863_reg/NET0131 ,
		_w8510_
	);
	LUT2 #(
		.INIT('h8)
	) name7003 (
		RESET_pad,
		\WX2042_reg/NET0131 ,
		_w8511_
	);
	LUT2 #(
		.INIT('h8)
	) name7004 (
		RESET_pad,
		\WX7178_reg/NET0131 ,
		_w8512_
	);
	LUT2 #(
		.INIT('h8)
	) name7005 (
		RESET_pad,
		\WX813_reg/NET0131 ,
		_w8513_
	);
	LUT2 #(
		.INIT('h8)
	) name7006 (
		RESET_pad,
		\WX5821_reg/NET0131 ,
		_w8514_
	);
	LUT2 #(
		.INIT('h8)
	) name7007 (
		RESET_pad,
		\WX5851_reg/NET0131 ,
		_w8515_
	);
	LUT2 #(
		.INIT('h8)
	) name7008 (
		RESET_pad,
		\WX8473_reg/NET0131 ,
		_w8516_
	);
	LUT2 #(
		.INIT('h8)
	) name7009 (
		RESET_pad,
		\WX4578_reg/NET0131 ,
		_w8517_
	);
	LUT2 #(
		.INIT('h8)
	) name7010 (
		RESET_pad,
		\WX3421_reg/NET0131 ,
		_w8518_
	);
	LUT2 #(
		.INIT('h8)
	) name7011 (
		RESET_pad,
		\WX9732_reg/NET0131 ,
		_w8519_
	);
	LUT2 #(
		.INIT('h8)
	) name7012 (
		RESET_pad,
		\WX11127_reg/NET0131 ,
		_w8520_
	);
	LUT2 #(
		.INIT('h8)
	) name7013 (
		RESET_pad,
		\WX5847_reg/NET0131 ,
		_w8521_
	);
	LUT2 #(
		.INIT('h8)
	) name7014 (
		RESET_pad,
		\WX8469_reg/NET0131 ,
		_w8522_
	);
	LUT2 #(
		.INIT('h8)
	) name7015 (
		RESET_pad,
		\WX763_reg/NET0131 ,
		_w8523_
	);
	LUT2 #(
		.INIT('h8)
	) name7016 (
		RESET_pad,
		\WX2036_reg/NET0131 ,
		_w8524_
	);
	LUT2 #(
		.INIT('h8)
	) name7017 (
		RESET_pad,
		\WX8475_reg/NET0131 ,
		_w8525_
	);
	LUT2 #(
		.INIT('h8)
	) name7018 (
		RESET_pad,
		\WX11021_reg/NET0131 ,
		_w8526_
	);
	LUT2 #(
		.INIT('h8)
	) name7019 (
		RESET_pad,
		\WX5901_reg/NET0131 ,
		_w8527_
	);
	LUT2 #(
		.INIT('h8)
	) name7020 (
		RESET_pad,
		\WX11005_reg/NET0131 ,
		_w8528_
	);
	LUT2 #(
		.INIT('h8)
	) name7021 (
		RESET_pad,
		\WX3275_reg/NET0131 ,
		_w8529_
	);
	LUT2 #(
		.INIT('h8)
	) name7022 (
		RESET_pad,
		\WX4632_reg/NET0131 ,
		_w8530_
	);
	LUT2 #(
		.INIT('h8)
	) name7023 (
		RESET_pad,
		\WX5841_reg/NET0131 ,
		_w8531_
	);
	LUT2 #(
		.INIT('h8)
	) name7024 (
		RESET_pad,
		\WX5973_reg/NET0131 ,
		_w8532_
	);
	LUT2 #(
		.INIT('h8)
	) name7025 (
		RESET_pad,
		\WX11019_reg/NET0131 ,
		_w8533_
	);
	LUT2 #(
		.INIT('h8)
	) name7026 (
		RESET_pad,
		\WX5829_reg/NET0131 ,
		_w8534_
	);
	LUT2 #(
		.INIT('h8)
	) name7027 (
		RESET_pad,
		\WX647_reg/NET0131 ,
		_w8535_
	);
	LUT2 #(
		.INIT('h8)
	) name7028 (
		RESET_pad,
		\WX5833_reg/NET0131 ,
		_w8536_
	);
	LUT2 #(
		.INIT('h8)
	) name7029 (
		RESET_pad,
		\WX5995_reg/NET0131 ,
		_w8537_
	);
	LUT2 #(
		.INIT('h8)
	) name7030 (
		RESET_pad,
		\WX3261_reg/NET0131 ,
		_w8538_
	);
	LUT2 #(
		.INIT('h8)
	) name7031 (
		RESET_pad,
		\WX7184_reg/NET0131 ,
		_w8539_
	);
	LUT2 #(
		.INIT('h8)
	) name7032 (
		RESET_pad,
		\WX11165_reg/NET0131 ,
		_w8540_
	);
	LUT2 #(
		.INIT('h8)
	) name7033 (
		RESET_pad,
		\WX8419_reg/NET0131 ,
		_w8541_
	);
	LUT2 #(
		.INIT('h8)
	) name7034 (
		RESET_pad,
		\WX697_reg/NET0131 ,
		_w8542_
	);
	LUT2 #(
		.INIT('h8)
	) name7035 (
		RESET_pad,
		\WX5823_reg/NET0131 ,
		_w8543_
	);
	LUT2 #(
		.INIT('h8)
	) name7036 (
		RESET_pad,
		\WX5857_reg/NET0131 ,
		_w8544_
	);
	LUT2 #(
		.INIT('h8)
	) name7037 (
		RESET_pad,
		\WX717_reg/NET0131 ,
		_w8545_
	);
	LUT2 #(
		.INIT('h8)
	) name7038 (
		RESET_pad,
		\WX4528_reg/NET0131 ,
		_w8546_
	);
	LUT2 #(
		.INIT('h8)
	) name7039 (
		RESET_pad,
		\WX5843_reg/NET0131 ,
		_w8547_
	);
	LUT2 #(
		.INIT('h8)
	) name7040 (
		RESET_pad,
		\WX5827_reg/NET0131 ,
		_w8548_
	);
	LUT2 #(
		.INIT('h8)
	) name7041 (
		RESET_pad,
		\WX7254_reg/NET0131 ,
		_w8549_
	);
	LUT2 #(
		.INIT('h8)
	) name7042 (
		RESET_pad,
		\WX5835_reg/NET0131 ,
		_w8550_
	);
	LUT2 #(
		.INIT('h8)
	) name7043 (
		RESET_pad,
		\WX737_reg/NET0131 ,
		_w8551_
	);
	LUT2 #(
		.INIT('h8)
	) name7044 (
		RESET_pad,
		\WX3293_reg/NET0131 ,
		_w8552_
	);
	LUT2 #(
		.INIT('h8)
	) name7045 (
		RESET_pad,
		\WX9846_reg/NET0131 ,
		_w8553_
	);
	LUT2 #(
		.INIT('h8)
	) name7046 (
		RESET_pad,
		\WX1964_reg/NET0131 ,
		_w8554_
	);
	LUT2 #(
		.INIT('h8)
	) name7047 (
		RESET_pad,
		\WX9814_reg/NET0131 ,
		_w8555_
	);
	LUT2 #(
		.INIT('h8)
	) name7048 (
		RESET_pad,
		\WX8505_reg/NET0131 ,
		_w8556_
	);
	LUT2 #(
		.INIT('h8)
	) name7049 (
		RESET_pad,
		\WX4658_reg/NET0131 ,
		_w8557_
	);
	LUT2 #(
		.INIT('h8)
	) name7050 (
		RESET_pad,
		\WX5825_reg/NET0131 ,
		_w8558_
	);
	LUT2 #(
		.INIT('h8)
	) name7051 (
		RESET_pad,
		\WX7188_reg/NET0131 ,
		_w8559_
	);
	LUT2 #(
		.INIT('h8)
	) name7052 (
		RESET_pad,
		\WX3399_reg/NET0131 ,
		_w8560_
	);
	LUT2 #(
		.INIT('h8)
	) name7053 (
		RESET_pad,
		\WX2034_reg/NET0131 ,
		_w8561_
	);
	LUT2 #(
		.INIT('h8)
	) name7054 (
		RESET_pad,
		\WX8471_reg/NET0131 ,
		_w8562_
	);
	LUT2 #(
		.INIT('h8)
	) name7055 (
		RESET_pad,
		\WX1968_reg/NET0131 ,
		_w8563_
	);
	LUT2 #(
		.INIT('h8)
	) name7056 (
		RESET_pad,
		\WX7290_reg/NET0131 ,
		_w8564_
	);
	LUT2 #(
		.INIT('h8)
	) name7057 (
		RESET_pad,
		\WX11101_reg/NET0131 ,
		_w8565_
	);
	LUT2 #(
		.INIT('h8)
	) name7058 (
		RESET_pad,
		\WX5837_reg/NET0131 ,
		_w8566_
	);
	LUT2 #(
		.INIT('h8)
	) name7059 (
		RESET_pad,
		\WX8459_reg/NET0131 ,
		_w8567_
	);
	LUT2 #(
		.INIT('h8)
	) name7060 (
		RESET_pad,
		\WX5817_reg/NET0131 ,
		_w8568_
	);
	LUT2 #(
		.INIT('h8)
	) name7061 (
		RESET_pad,
		\WX4668_reg/NET0131 ,
		_w8569_
	);
	LUT2 #(
		.INIT('h8)
	) name7062 (
		RESET_pad,
		\WX4614_reg/NET0131 ,
		_w8570_
	);
	LUT2 #(
		.INIT('h8)
	) name7063 (
		RESET_pad,
		\WX4672_reg/NET0131 ,
		_w8571_
	);
	LUT2 #(
		.INIT('h8)
	) name7064 (
		RESET_pad,
		\WX9844_reg/NET0131 ,
		_w8572_
	);
	LUT2 #(
		.INIT('h8)
	) name7065 (
		RESET_pad,
		\WX4648_reg/NET0131 ,
		_w8573_
	);
	LUT2 #(
		.INIT('h8)
	) name7066 (
		RESET_pad,
		\WX3325_reg/NET0131 ,
		_w8574_
	);
	LUT2 #(
		.INIT('h8)
	) name7067 (
		RESET_pad,
		\WX713_reg/NET0131 ,
		_w8575_
	);
	LUT2 #(
		.INIT('h8)
	) name7068 (
		RESET_pad,
		\WX11069_reg/NET0131 ,
		_w8576_
	);
	LUT2 #(
		.INIT('h8)
	) name7069 (
		RESET_pad,
		\WX9746_reg/NET0131 ,
		_w8577_
	);
	LUT2 #(
		.INIT('h8)
	) name7070 (
		RESET_pad,
		\WX9874_reg/NET0131 ,
		_w8578_
	);
	LUT2 #(
		.INIT('h8)
	) name7071 (
		RESET_pad,
		\WX8451_reg/NET0131 ,
		_w8579_
	);
	LUT2 #(
		.INIT('h8)
	) name7072 (
		RESET_pad,
		\WX1950_reg/NET0131 ,
		_w8580_
	);
	LUT2 #(
		.INIT('h8)
	) name7073 (
		RESET_pad,
		\WX5909_reg/NET0131 ,
		_w8581_
	);
	LUT2 #(
		.INIT('h8)
	) name7074 (
		RESET_pad,
		\WX8515_reg/NET0131 ,
		_w8582_
	);
	LUT2 #(
		.INIT('h8)
	) name7075 (
		RESET_pad,
		\WX1960_reg/NET0131 ,
		_w8583_
	);
	LUT2 #(
		.INIT('h8)
	) name7076 (
		RESET_pad,
		\WX7236_reg/NET0131 ,
		_w8584_
	);
	LUT2 #(
		.INIT('h8)
	) name7077 (
		RESET_pad,
		\WX4700_reg/NET0131 ,
		_w8585_
	);
	LUT2 #(
		.INIT('h8)
	) name7078 (
		RESET_pad,
		\WX4692_reg/NET0131 ,
		_w8586_
	);
	LUT2 #(
		.INIT('h8)
	) name7079 (
		RESET_pad,
		\WX1976_reg/NET0131 ,
		_w8587_
	);
	LUT2 #(
		.INIT('h8)
	) name7080 (
		RESET_pad,
		\WX1980_reg/NET0131 ,
		_w8588_
	);
	LUT2 #(
		.INIT('h8)
	) name7081 (
		RESET_pad,
		\WX8443_reg/NET0131 ,
		_w8589_
	);
	LUT2 #(
		.INIT('h8)
	) name7082 (
		RESET_pad,
		\WX1996_reg/NET0131 ,
		_w8590_
	);
	LUT2 #(
		.INIT('h8)
	) name7083 (
		RESET_pad,
		\WX2032_reg/NET0131 ,
		_w8591_
	);
	LUT2 #(
		.INIT('h8)
	) name7084 (
		RESET_pad,
		\WX9848_reg/NET0131 ,
		_w8592_
	);
	LUT2 #(
		.INIT('h8)
	) name7085 (
		RESET_pad,
		\WX11023_reg/NET0131 ,
		_w8593_
	);
	LUT2 #(
		.INIT('h8)
	) name7086 (
		RESET_pad,
		\WX3317_reg/NET0131 ,
		_w8594_
	);
	LUT2 #(
		.INIT('h8)
	) name7087 (
		RESET_pad,
		\WX9740_reg/NET0131 ,
		_w8595_
	);
	LUT2 #(
		.INIT('h8)
	) name7088 (
		RESET_pad,
		\WX2014_reg/NET0131 ,
		_w8596_
	);
	LUT2 #(
		.INIT('h8)
	) name7089 (
		RESET_pad,
		\WX11155_reg/NET0131 ,
		_w8597_
	);
	LUT2 #(
		.INIT('h8)
	) name7090 (
		RESET_pad,
		\WX2020_reg/NET0131 ,
		_w8598_
	);
	LUT2 #(
		.INIT('h8)
	) name7091 (
		RESET_pad,
		\WX6007_reg/NET0131 ,
		_w8599_
	);
	LUT2 #(
		.INIT('h8)
	) name7092 (
		RESET_pad,
		\WX4708_reg/NET0131 ,
		_w8600_
	);
	LUT2 #(
		.INIT('h8)
	) name7093 (
		RESET_pad,
		\WX2044_reg/NET0131 ,
		_w8601_
	);
	LUT2 #(
		.INIT('h8)
	) name7094 (
		RESET_pad,
		\WX2046_reg/NET0131 ,
		_w8602_
	);
	LUT2 #(
		.INIT('h8)
	) name7095 (
		RESET_pad,
		\WX3359_reg/NET0131 ,
		_w8603_
	);
	LUT2 #(
		.INIT('h8)
	) name7096 (
		RESET_pad,
		\WX2054_reg/NET0131 ,
		_w8604_
	);
	LUT2 #(
		.INIT('h8)
	) name7097 (
		RESET_pad,
		\WX5869_reg/NET0131 ,
		_w8605_
	);
	LUT2 #(
		.INIT('h8)
	) name7098 (
		RESET_pad,
		\WX11179_reg/NET0131 ,
		_w8606_
	);
	LUT2 #(
		.INIT('h8)
	) name7099 (
		RESET_pad,
		\WX11129_reg/NET0131 ,
		_w8607_
	);
	LUT2 #(
		.INIT('h8)
	) name7100 (
		RESET_pad,
		\WX11145_reg/NET0131 ,
		_w8608_
	);
	LUT2 #(
		.INIT('h8)
	) name7101 (
		RESET_pad,
		\WX699_reg/NET0131 ,
		_w8609_
	);
	LUT2 #(
		.INIT('h8)
	) name7102 (
		RESET_pad,
		\WX2080_reg/NET0131 ,
		_w8610_
	);
	LUT2 #(
		.INIT('h8)
	) name7103 (
		RESET_pad,
		\WX2082_reg/NET0131 ,
		_w8611_
	);
	LUT2 #(
		.INIT('h8)
	) name7104 (
		RESET_pad,
		\WX2030_reg/NET0131 ,
		_w8612_
	);
	LUT2 #(
		.INIT('h8)
	) name7105 (
		RESET_pad,
		\WX11075_reg/NET0131 ,
		_w8613_
	);
	LUT2 #(
		.INIT('h8)
	) name7106 (
		RESET_pad,
		\WX3311_reg/NET0131 ,
		_w8614_
	);
	LUT2 #(
		.INIT('h8)
	) name7107 (
		RESET_pad,
		\WX9818_reg/NET0131 ,
		_w8615_
	);
	LUT2 #(
		.INIT('h8)
	) name7108 (
		RESET_pad,
		\WX701_reg/NET0131 ,
		_w8616_
	);
	LUT2 #(
		.INIT('h8)
	) name7109 (
		RESET_pad,
		\WX2026_reg/NET0131 ,
		_w8617_
	);
	LUT2 #(
		.INIT('h8)
	) name7110 (
		RESET_pad,
		\WX5839_reg/NET0131 ,
		_w8618_
	);
	LUT2 #(
		.INIT('h8)
	) name7111 (
		RESET_pad,
		\WX11007_reg/NET0131 ,
		_w8619_
	);
	LUT2 #(
		.INIT('h8)
	) name7112 (
		RESET_pad,
		\WX8563_reg/NET0131 ,
		_w8620_
	);
	LUT2 #(
		.INIT('h8)
	) name7113 (
		RESET_pad,
		\WX3309_reg/NET0131 ,
		_w8621_
	);
	LUT2 #(
		.INIT('h8)
	) name7114 (
		RESET_pad,
		\WX9710_reg/NET0131 ,
		_w8622_
	);
	LUT2 #(
		.INIT('h8)
	) name7115 (
		RESET_pad,
		\WX4574_reg/NET0131 ,
		_w8623_
	);
	LUT2 #(
		.INIT('h8)
	) name7116 (
		RESET_pad,
		\WX7202_reg/NET0131 ,
		_w8624_
	);
	LUT2 #(
		.INIT('h8)
	) name7117 (
		RESET_pad,
		\WX8415_reg/NET0131 ,
		_w8625_
	);
	LUT2 #(
		.INIT('h8)
	) name7118 (
		RESET_pad,
		\WX9810_reg/NET0131 ,
		_w8626_
	);
	LUT2 #(
		.INIT('h8)
	) name7119 (
		RESET_pad,
		\WX3269_reg/NET0131 ,
		_w8627_
	);
	LUT2 #(
		.INIT('h8)
	) name7120 (
		RESET_pad,
		\WX7200_reg/NET0131 ,
		_w8628_
	);
	LUT2 #(
		.INIT('h8)
	) name7121 (
		RESET_pad,
		\WX9752_reg/NET0131 ,
		_w8629_
	);
	LUT2 #(
		.INIT('h8)
	) name7122 (
		RESET_pad,
		\WX7174_reg/NET0131 ,
		_w8630_
	);
	LUT2 #(
		.INIT('h8)
	) name7123 (
		RESET_pad,
		\WX3389_reg/NET0131 ,
		_w8631_
	);
	LUT2 #(
		.INIT('h8)
	) name7124 (
		RESET_pad,
		\WX8581_reg/NET0131 ,
		_w8632_
	);
	LUT2 #(
		.INIT('h8)
	) name7125 (
		RESET_pad,
		\WX5845_reg/NET0131 ,
		_w8633_
	);
	LUT2 #(
		.INIT('h8)
	) name7126 (
		RESET_pad,
		\WX5873_reg/NET0131 ,
		_w8634_
	);
	LUT2 #(
		.INIT('h8)
	) name7127 (
		RESET_pad,
		\WX9782_reg/NET0131 ,
		_w8635_
	);
	LUT2 #(
		.INIT('h8)
	) name7128 (
		RESET_pad,
		\WX7208_reg/NET0131 ,
		_w8636_
	);
	LUT2 #(
		.INIT('h8)
	) name7129 (
		RESET_pad,
		\WX8485_reg/NET0131 ,
		_w8637_
	);
	LUT2 #(
		.INIT('h8)
	) name7130 (
		RESET_pad,
		\WX8575_reg/NET0131 ,
		_w8638_
	);
	LUT2 #(
		.INIT('h8)
	) name7131 (
		RESET_pad,
		\WX8481_reg/NET0131 ,
		_w8639_
	);
	LUT2 #(
		.INIT('h8)
	) name7132 (
		RESET_pad,
		\WX4532_reg/NET0131 ,
		_w8640_
	);
	LUT2 #(
		.INIT('h8)
	) name7133 (
		RESET_pad,
		\WX11031_reg/NET0131 ,
		_w8641_
	);
	LUT2 #(
		.INIT('h8)
	) name7134 (
		RESET_pad,
		\WX7210_reg/NET0131 ,
		_w8642_
	);
	LUT2 #(
		.INIT('h8)
	) name7135 (
		RESET_pad,
		\WX7206_reg/NET0131 ,
		_w8643_
	);
	LUT2 #(
		.INIT('h8)
	) name7136 (
		RESET_pad,
		\WX10989_reg/NET0131 ,
		_w8644_
	);
	LUT2 #(
		.INIT('h8)
	) name7137 (
		RESET_pad,
		\WX765_reg/NET0131 ,
		_w8645_
	);
	LUT2 #(
		.INIT('h8)
	) name7138 (
		RESET_pad,
		\WX799_reg/NET0131 ,
		_w8646_
	);
	LUT2 #(
		.INIT('h8)
	) name7139 (
		RESET_pad,
		\WX711_reg/NET0131 ,
		_w8647_
	);
	LUT2 #(
		.INIT('h8)
	) name7140 (
		RESET_pad,
		\WX751_reg/NET0131 ,
		_w8648_
	);
	LUT2 #(
		.INIT('h8)
	) name7141 (
		RESET_pad,
		\WX10993_reg/NET0131 ,
		_w8649_
	);
	LUT2 #(
		.INIT('h8)
	) name7142 (
		RESET_pad,
		\WX3413_reg/NET0131 ,
		_w8650_
	);
	LUT2 #(
		.INIT('h8)
	) name7143 (
		RESET_pad,
		\WX8577_reg/NET0131 ,
		_w8651_
	);
	LUT2 #(
		.INIT('h8)
	) name7144 (
		RESET_pad,
		\WX3291_reg/NET0131 ,
		_w8652_
	);
	LUT2 #(
		.INIT('h8)
	) name7145 (
		RESET_pad,
		\WX741_reg/NET0131 ,
		_w8653_
	);
	LUT2 #(
		.INIT('h8)
	) name7146 (
		RESET_pad,
		\WX749_reg/NET0131 ,
		_w8654_
	);
	LUT2 #(
		.INIT('h8)
	) name7147 (
		RESET_pad,
		\WX7266_reg/NET0131 ,
		_w8655_
	);
	LUT2 #(
		.INIT('h8)
	) name7148 (
		RESET_pad,
		\WX4568_reg/NET0131 ,
		_w8656_
	);
	LUT2 #(
		.INIT('h8)
	) name7149 (
		RESET_pad,
		\WX8527_reg/NET0131 ,
		_w8657_
	);
	LUT2 #(
		.INIT('h8)
	) name7150 (
		RESET_pad,
		\WX1982_reg/NET0131 ,
		_w8658_
	);
	LUT2 #(
		.INIT('h8)
	) name7151 (
		RESET_pad,
		\WX11035_reg/NET0131 ,
		_w8659_
	);
	LUT2 #(
		.INIT('h8)
	) name7152 (
		RESET_pad,
		\WX11039_reg/NET0131 ,
		_w8660_
	);
	LUT2 #(
		.INIT('h8)
	) name7153 (
		RESET_pad,
		\WX3251_reg/NET0131 ,
		_w8661_
	);
	LUT2 #(
		.INIT('h8)
	) name7154 (
		RESET_pad,
		\WX745_reg/NET0131 ,
		_w8662_
	);
	LUT2 #(
		.INIT('h1)
	) name7155 (
		\TM0_pad ,
		_w1543_,
		_w8663_
	);
	LUT2 #(
		.INIT('h2)
	) name7156 (
		_w2846_,
		_w8663_,
		_w8664_
	);
	LUT2 #(
		.INIT('h2)
	) name7157 (
		\TM0_pad ,
		\_2088__reg/NET0131 ,
		_w8665_
	);
	LUT2 #(
		.INIT('h2)
	) name7158 (
		_w1976_,
		_w8665_,
		_w8666_
	);
	LUT2 #(
		.INIT('h4)
	) name7159 (
		_w5074_,
		_w8666_,
		_w8667_
	);
	LUT2 #(
		.INIT('h1)
	) name7160 (
		_w8664_,
		_w8667_,
		_w8668_
	);
	LUT2 #(
		.INIT('h1)
	) name7161 (
		\TM0_pad ,
		_w1955_,
		_w8669_
	);
	LUT2 #(
		.INIT('h2)
	) name7162 (
		_w2023_,
		_w8669_,
		_w8670_
	);
	LUT2 #(
		.INIT('h2)
	) name7163 (
		\TM0_pad ,
		\_2085__reg/NET0131 ,
		_w8671_
	);
	LUT2 #(
		.INIT('h2)
	) name7164 (
		_w1976_,
		_w8671_,
		_w8672_
	);
	LUT2 #(
		.INIT('h4)
	) name7165 (
		_w5455_,
		_w8672_,
		_w8673_
	);
	LUT2 #(
		.INIT('h1)
	) name7166 (
		_w8670_,
		_w8673_,
		_w8674_
	);
	LUT2 #(
		.INIT('h1)
	) name7167 (
		\TM0_pad ,
		_w1903_,
		_w8675_
	);
	LUT2 #(
		.INIT('h2)
	) name7168 (
		_w3953_,
		_w8675_,
		_w8676_
	);
	LUT2 #(
		.INIT('h2)
	) name7169 (
		\TM0_pad ,
		\_2081__reg/NET0131 ,
		_w8677_
	);
	LUT2 #(
		.INIT('h2)
	) name7170 (
		_w1976_,
		_w8677_,
		_w8678_
	);
	LUT2 #(
		.INIT('h4)
	) name7171 (
		_w5995_,
		_w8678_,
		_w8679_
	);
	LUT2 #(
		.INIT('h1)
	) name7172 (
		_w8676_,
		_w8679_,
		_w8680_
	);
	LUT2 #(
		.INIT('h1)
	) name7173 (
		\TM0_pad ,
		_w1582_,
		_w8681_
	);
	LUT2 #(
		.INIT('h2)
	) name7174 (
		_w2341_,
		_w8681_,
		_w8682_
	);
	LUT2 #(
		.INIT('h2)
	) name7175 (
		\TM0_pad ,
		\_2091__reg/NET0131 ,
		_w8683_
	);
	LUT2 #(
		.INIT('h2)
	) name7176 (
		_w1976_,
		_w8683_,
		_w8684_
	);
	LUT2 #(
		.INIT('h4)
	) name7177 (
		_w4687_,
		_w8684_,
		_w8685_
	);
	LUT2 #(
		.INIT('h1)
	) name7178 (
		_w8682_,
		_w8685_,
		_w8686_
	);
	LUT2 #(
		.INIT('h1)
	) name7179 (
		\TM0_pad ,
		_w1968_,
		_w8687_
	);
	LUT2 #(
		.INIT('h2)
	) name7180 (
		_w3172_,
		_w8687_,
		_w8688_
	);
	LUT2 #(
		.INIT('h2)
	) name7181 (
		\TM0_pad ,
		\_2086__reg/NET0131 ,
		_w8689_
	);
	LUT2 #(
		.INIT('h2)
	) name7182 (
		_w1976_,
		_w8689_,
		_w8690_
	);
	LUT2 #(
		.INIT('h4)
	) name7183 (
		_w5332_,
		_w8690_,
		_w8691_
	);
	LUT2 #(
		.INIT('h1)
	) name7184 (
		_w8688_,
		_w8691_,
		_w8692_
	);
	LUT2 #(
		.INIT('h1)
	) name7185 (
		\TM0_pad ,
		_w1942_,
		_w8693_
	);
	LUT2 #(
		.INIT('h2)
	) name7186 (
		_w3483_,
		_w8693_,
		_w8694_
	);
	LUT2 #(
		.INIT('h2)
	) name7187 (
		\TM0_pad ,
		\_2084__reg/NET0131 ,
		_w8695_
	);
	LUT2 #(
		.INIT('h2)
	) name7188 (
		_w1976_,
		_w8695_,
		_w8696_
	);
	LUT2 #(
		.INIT('h4)
	) name7189 (
		_w5575_,
		_w8696_,
		_w8697_
	);
	LUT2 #(
		.INIT('h1)
	) name7190 (
		_w8694_,
		_w8697_,
		_w8698_
	);
	LUT2 #(
		.INIT('h1)
	) name7191 (
		\TM0_pad ,
		_w1672_,
		_w8699_
	);
	LUT2 #(
		.INIT('h2)
	) name7192 (
		_w4382_,
		_w8699_,
		_w8700_
	);
	LUT2 #(
		.INIT('h2)
	) name7193 (
		\TM0_pad ,
		\_2078__reg/NET0131 ,
		_w8701_
	);
	LUT2 #(
		.INIT('h2)
	) name7194 (
		_w1976_,
		_w8701_,
		_w8702_
	);
	LUT2 #(
		.INIT('h4)
	) name7195 (
		_w6508_,
		_w8702_,
		_w8703_
	);
	LUT2 #(
		.INIT('h1)
	) name7196 (
		_w8700_,
		_w8703_,
		_w8704_
	);
	LUT2 #(
		.INIT('h2)
	) name7197 (
		_w1974_,
		_w3082_,
		_w8705_
	);
	LUT2 #(
		.INIT('h1)
	) name7198 (
		\DATA_0_15_pad ,
		\TM0_pad ,
		_w8706_
	);
	LUT2 #(
		.INIT('h2)
	) name7199 (
		\TM0_pad ,
		\_2348__reg/NET0131 ,
		_w8707_
	);
	LUT2 #(
		.INIT('h2)
	) name7200 (
		_w1976_,
		_w8706_,
		_w8708_
	);
	LUT2 #(
		.INIT('h4)
	) name7201 (
		_w8707_,
		_w8708_,
		_w8709_
	);
	LUT2 #(
		.INIT('h1)
	) name7202 (
		_w8705_,
		_w8709_,
		_w8710_
	);
	assign \DATA_9_0_pad  = _w1520_ ;
	assign \DATA_9_10_pad  = _w1533_ ;
	assign \DATA_9_11_pad  = _w1546_ ;
	assign \DATA_9_12_pad  = _w1559_ ;
	assign \DATA_9_13_pad  = _w1572_ ;
	assign \DATA_9_14_pad  = _w1585_ ;
	assign \DATA_9_15_pad  = _w1598_ ;
	assign \DATA_9_16_pad  = _w1614_ ;
	assign \DATA_9_17_pad  = _w1630_ ;
	assign \DATA_9_18_pad  = _w1646_ ;
	assign \DATA_9_19_pad  = _w1662_ ;
	assign \DATA_9_1_pad  = _w1675_ ;
	assign \DATA_9_20_pad  = _w1691_ ;
	assign \DATA_9_21_pad  = _w1707_ ;
	assign \DATA_9_22_pad  = _w1723_ ;
	assign \DATA_9_23_pad  = _w1739_ ;
	assign \DATA_9_24_pad  = _w1755_ ;
	assign \DATA_9_25_pad  = _w1771_ ;
	assign \DATA_9_26_pad  = _w1787_ ;
	assign \DATA_9_27_pad  = _w1803_ ;
	assign \DATA_9_28_pad  = _w1819_ ;
	assign \DATA_9_29_pad  = _w1835_ ;
	assign \DATA_9_2_pad  = _w1848_ ;
	assign \DATA_9_30_pad  = _w1864_ ;
	assign \DATA_9_31_pad  = _w1880_ ;
	assign \DATA_9_3_pad  = _w1893_ ;
	assign \DATA_9_4_pad  = _w1906_ ;
	assign \DATA_9_5_pad  = _w1919_ ;
	assign \DATA_9_6_pad  = _w1932_ ;
	assign \DATA_9_7_pad  = _w1945_ ;
	assign \DATA_9_8_pad  = _w1958_ ;
	assign \DATA_9_9_pad  = _w1971_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b0;
	assign \g19/_0_  = _w1990_ ;
	assign \g35/_0_  = _w2022_ ;
	assign \g36/_0_  = _w2039_ ;
	assign \g40/_0_  = _w2056_ ;
	assign \g55780/_0_  = _w2076_ ;
	assign \g55783/_0_  = _w2096_ ;
	assign \g55795/_0_  = _w2121_ ;
	assign \g55796/_0_  = _w2140_ ;
	assign \g55797/_0_  = _w2172_ ;
	assign \g55798/_0_  = _w2204_ ;
	assign \g55799/_0_  = _w2236_ ;
	assign \g55800/_0_  = _w2268_ ;
	assign \g55801/_0_  = _w2300_ ;
	assign \g55802/_0_  = _w2320_ ;
	assign \g55803/_0_  = _w2340_ ;
	assign \g55834/_0_  = _w2366_ ;
	assign \g55835/_0_  = _w2385_ ;
	assign \g55836/_0_  = _w2404_ ;
	assign \g55837/_0_  = _w2423_ ;
	assign \g55838/_0_  = _w2438_ ;
	assign \g55839/_0_  = _w2457_ ;
	assign \g55840/_0_  = _w2476_ ;
	assign \g55841/_0_  = _w2496_ ;
	assign \g55842/_0_  = _w2516_ ;
	assign \g55856/_0_  = _w2517_ ;
	assign \g55894/_0_  = _w2542_ ;
	assign \g55895/_0_  = _w2561_ ;
	assign \g55896/_0_  = _w2580_ ;
	assign \g55897/_0_  = _w2599_ ;
	assign \g55898/_0_  = _w2614_ ;
	assign \g55899/_0_  = _w2629_ ;
	assign \g55900/_0_  = _w2648_ ;
	assign \g55901/_0_  = _w2668_ ;
	assign \g55902/_0_  = _w2675_ ;
	assign \g55916/_0_  = _w2676_ ;
	assign \g55953/_0_  = _w2702_ ;
	assign \g55954/_0_  = _w2721_ ;
	assign \g55955/_0_  = _w2740_ ;
	assign \g55956/_0_  = _w2759_ ;
	assign \g55957/_0_  = _w2774_ ;
	assign \g55958/_0_  = _w2789_ ;
	assign \g55959/_0_  = _w2804_ ;
	assign \g55960/_0_  = _w2824_ ;
	assign \g55961/_0_  = _w2844_ ;
	assign \g55975/_0_  = _w2845_ ;
	assign \g56012/_0_  = _w2871_ ;
	assign \g56013/_0_  = _w2886_ ;
	assign \g56014/_0_  = _w2905_ ;
	assign \g56015/_0_  = _w2924_ ;
	assign \g56016/_0_  = _w2939_ ;
	assign \g56017/_0_  = _w2954_ ;
	assign \g56018/_0_  = _w2969_ ;
	assign \g56019/_0_  = _w2989_ ;
	assign \g56020/_0_  = _w3009_ ;
	assign \g56034/_0_  = _w3010_ ;
	assign \g56071/_0_  = _w3036_ ;
	assign \g56072/_0_  = _w3051_ ;
	assign \g56073/_0_  = _w3070_ ;
	assign \g56074/_0_  = _w3085_ ;
	assign \g56075/_0_  = _w3100_ ;
	assign \g56076/_0_  = _w3115_ ;
	assign \g56077/_0_  = _w3130_ ;
	assign \g56078/_0_  = _w3150_ ;
	assign \g56079/_0_  = _w3170_ ;
	assign \g56093/_0_  = _w3171_ ;
	assign \g56130/_0_  = _w3197_ ;
	assign \g56131/_0_  = _w3212_ ;
	assign \g56132/_0_  = _w3227_ ;
	assign \g56133/_0_  = _w3246_ ;
	assign \g56134/_0_  = _w3261_ ;
	assign \g56135/_0_  = _w3276_ ;
	assign \g56136/_0_  = _w3291_ ;
	assign \g56137/_0_  = _w3311_ ;
	assign \g56138/_0_  = _w3331_ ;
	assign \g56152/_0_  = _w3332_ ;
	assign \g56189/_0_  = _w3357_ ;
	assign \g56190/_0_  = _w3372_ ;
	assign \g56191/_0_  = _w3377_ ;
	assign \g56192/_0_  = _w3396_ ;
	assign \g56193/_0_  = _w3411_ ;
	assign \g56194/_0_  = _w3426_ ;
	assign \g56195/_0_  = _w3441_ ;
	assign \g56196/_0_  = _w3461_ ;
	assign \g56197/_0_  = _w3481_ ;
	assign \g56211/_0_  = _w3482_ ;
	assign \g56248/_0_  = _w3508_ ;
	assign \g56249/_0_  = _w3523_ ;
	assign \g56250/_0_  = _w3538_ ;
	assign \g56251/_0_  = _w3557_ ;
	assign \g56252/_0_  = _w3572_ ;
	assign \g56253/_0_  = _w3587_ ;
	assign \g56254/_0_  = _w3602_ ;
	assign \g56255/_0_  = _w3622_ ;
	assign \g56256/_0_  = _w3642_ ;
	assign \g56270/_0_  = _w3643_ ;
	assign \g56307/_0_  = _w3669_ ;
	assign \g56308/_0_  = _w3684_ ;
	assign \g56309/_0_  = _w3699_ ;
	assign \g56310/_0_  = _w3718_ ;
	assign \g56311/_0_  = _w3733_ ;
	assign \g56312/_0_  = _w3748_ ;
	assign \g56313/_0_  = _w3763_ ;
	assign \g56314/_0_  = _w3783_ ;
	assign \g56315/_0_  = _w3803_ ;
	assign \g56329/_0_  = _w3804_ ;
	assign \g56366/_0_  = _w3830_ ;
	assign \g56367/_0_  = _w3845_ ;
	assign \g56368/_0_  = _w3860_ ;
	assign \g56369/_0_  = _w3879_ ;
	assign \g56370/_0_  = _w3894_ ;
	assign \g56371/_0_  = _w3909_ ;
	assign \g56372/_0_  = _w3924_ ;
	assign \g56373/_0_  = _w3944_ ;
	assign \g56374/_0_  = _w3951_ ;
	assign \g56388/_0_  = _w3952_ ;
	assign \g56425/_0_  = _w3978_ ;
	assign \g56426/_0_  = _w3993_ ;
	assign \g56427/_0_  = _w4008_ ;
	assign \g56428/_0_  = _w4027_ ;
	assign \g56429/_0_  = _w4042_ ;
	assign \g56430/_0_  = _w4057_ ;
	assign \g56431/_0_  = _w4072_ ;
	assign \g56432/_0_  = _w4092_ ;
	assign \g56433/_0_  = _w4099_ ;
	assign \g56447/_0_  = _w4100_ ;
	assign \g56484/_0_  = _w4126_ ;
	assign \g56485/_0_  = _w4141_ ;
	assign \g56486/_0_  = _w4146_ ;
	assign \g56487/_0_  = _w4165_ ;
	assign \g56488/_0_  = _w4180_ ;
	assign \g56489/_0_  = _w4195_ ;
	assign \g56490/_0_  = _w4210_ ;
	assign \g56491/_0_  = _w4230_ ;
	assign \g56492/_0_  = _w4237_ ;
	assign \g56507/_0_  = _w4238_ ;
	assign \g56543/_0_  = _w4264_ ;
	assign \g56544/_0_  = _w4279_ ;
	assign \g56545/_0_  = _w4294_ ;
	assign \g56546/_0_  = _w4309_ ;
	assign \g56547/_0_  = _w4328_ ;
	assign \g56548/_0_  = _w4343_ ;
	assign \g56549/_0_  = _w4358_ ;
	assign \g56551/_0_  = _w4365_ ;
	assign \g56567/_0_  = _w4366_ ;
	assign \g56602/_0_  = _w4381_ ;
	assign \g56603/_0_  = _w4407_ ;
	assign \g56604/_0_  = _w4422_ ;
	assign \g56605/_0_  = _w4437_ ;
	assign \g56606/_0_  = _w4452_ ;
	assign \g56607/_0_  = _w4471_ ;
	assign \g56608/_0_  = _w4486_ ;
	assign \g56610/_0_  = _w4493_ ;
	assign \g56627/_0_  = _w4494_ ;
	assign \g56661/_0_  = _w4509_ ;
	assign \g56662/_0_  = _w4535_ ;
	assign \g56663/_0_  = _w4550_ ;
	assign \g56664/_0_  = _w4565_ ;
	assign \g56665/_0_  = _w4580_ ;
	assign \g56666/_0_  = _w4585_ ;
	assign \g56667/_0_  = _w4600_ ;
	assign \g56668/_0_  = _w4616_ ;
	assign \g56686/_0_  = _w4617_ ;
	assign \g56720/_0_  = _w4632_ ;
	assign \g56721/_0_  = _w4647_ ;
	assign \g56722/_0_  = _w4662_ ;
	assign \g56723/_0_  = _w4677_ ;
	assign \g56724/_0_  = _w4692_ ;
	assign \g56725/_0_  = _w4707_ ;
	assign \g56726/_0_  = _w4739_ ;
	assign \g56727/_0_  = _w4755_ ;
	assign \g56728/_0_  = _w4761_ ;
	assign \g56745/_0_  = _w4762_ ;
	assign \g56779/_0_  = _w4777_ ;
	assign \g56780/_0_  = _w4792_ ;
	assign \g56781/_0_  = _w4811_ ;
	assign \g56782/_0_  = _w4826_ ;
	assign \g56783/_0_  = _w4831_ ;
	assign \g56784/_0_  = _w4846_ ;
	assign \g56785/_0_  = _w4865_ ;
	assign \g56804/_0_  = _w4866_ ;
	assign \g56838/_0_  = _w4881_ ;
	assign \g56839/_0_  = _w4896_ ;
	assign \g56840/_0_  = _w4915_ ;
	assign \g56841/_0_  = _w4930_ ;
	assign \g56842/_0_  = _w4949_ ;
	assign \g56843/_0_  = _w4954_ ;
	assign \g56844/_0_  = _w4973_ ;
	assign \g56845/_0_  = _w4989_ ;
	assign \g56846/_0_  = _w4995_ ;
	assign \g56863/_0_  = _w4996_ ;
	assign \g56897/_0_  = _w5011_ ;
	assign \g56898/_0_  = _w5030_ ;
	assign \g56899/_0_  = _w5045_ ;
	assign \g56900/_0_  = _w5064_ ;
	assign \g56901/_0_  = _w5079_ ;
	assign \g56902/_0_  = _w5098_ ;
	assign \g56903/_0_  = _w5117_ ;
	assign \g56905/_0_  = _w5123_ ;
	assign \g56921/_0_  = _w5124_ ;
	assign \g56956/_0_  = _w5143_ ;
	assign \g56957/_0_  = _w5162_ ;
	assign \g56958/_0_  = _w5177_ ;
	assign \g56959/_0_  = _w5196_ ;
	assign \g56960/_0_  = _w5201_ ;
	assign \g56961/_0_  = _w5220_ ;
	assign \g56962/_0_  = _w5239_ ;
	assign \g56964/_0_  = _w5245_ ;
	assign \g56980/_0_  = _w5246_ ;
	assign \g57015/_0_  = _w5265_ ;
	assign \g57016/_0_  = _w5284_ ;
	assign \g57017/_0_  = _w5303_ ;
	assign \g57018/_0_  = _w5322_ ;
	assign \g57019/_0_  = _w5337_ ;
	assign \g57020/_0_  = _w5356_ ;
	assign \g57021/_0_  = _w5375_ ;
	assign \g57023/_0_  = _w5381_ ;
	assign \g57040/_0_  = _w5382_ ;
	assign \g57074/_0_  = _w5401_ ;
	assign \g57075/_0_  = _w5407_ ;
	assign \g57076/_0_  = _w5426_ ;
	assign \g57077/_0_  = _w5445_ ;
	assign \g57078/_0_  = _w5460_ ;
	assign \g57079/_0_  = _w5479_ ;
	assign \g57080/_0_  = _w5498_ ;
	assign \g57081/_0_  = _w5514_ ;
	assign \g57099/_0_  = _w5515_ ;
	assign \g57133/_0_  = _w5521_ ;
	assign \g57134/_0_  = _w5527_ ;
	assign \g57135/_0_  = _w5546_ ;
	assign \g57136/_0_  = _w5565_ ;
	assign \g57137/_0_  = _w5580_ ;
	assign \g57138/_0_  = _w5599_ ;
	assign \g57139/_0_  = _w5618_ ;
	assign \g57140/_0_  = _w5634_ ;
	assign \g57141/_0_  = _w5640_ ;
	assign \g57159/_0_  = _w5641_ ;
	assign \g57193/_0_  = _w5660_ ;
	assign \g57195/_0_  = _w5679_ ;
	assign \g57196/_0_  = _w5698_ ;
	assign \g57197/_0_  = _w5703_ ;
	assign \g57198/_0_  = _w5722_ ;
	assign \g57199/_0_  = _w5741_ ;
	assign \g57200/_0_  = _w5761_ ;
	assign \g57202/_0_  = _w5767_ ;
	assign \g57219/_0_  = _w5768_ ;
	assign \g57254/_0_  = _w5787_ ;
	assign \g57255/_0_  = _w5806_ ;
	assign \g57256/_0_  = _w5812_ ;
	assign \g57257/_0_  = _w5831_ ;
	assign \g57258/_0_  = _w5850_ ;
	assign \g57259/_0_  = _w5855_ ;
	assign \g57260/_0_  = _w5874_ ;
	assign \g57262/_0_  = _w5890_ ;
	assign \g57263/_0_  = _w5896_ ;
	assign \g57285/_0_  = _w5897_ ;
	assign \g57318/_0_  = _w5916_ ;
	assign \g57319/_0_  = _w5935_ ;
	assign \g57320/_0_  = _w5941_ ;
	assign \g57321/_0_  = _w5947_ ;
	assign \g57322/_0_  = _w5966_ ;
	assign \g57323/_0_  = _w5985_ ;
	assign \g57324/_0_  = _w6000_ ;
	assign \g57325/_0_  = _w6019_ ;
	assign \g57326/_0_  = _w6035_ ;
	assign \g57328/_0_  = _w6051_ ;
	assign \g57329/_0_  = _w6058_ ;
	assign \g57330/_0_  = _w6064_ ;
	assign \g57350/_0_  = _w6065_ ;
	assign \g57387/_0_  = _w6084_ ;
	assign \g57388/_0_  = _w6103_ ;
	assign \g57390/_0_  = _w6109_ ;
	assign \g57391/_0_  = _w6128_ ;
	assign \g57392/_0_  = _w6147_ ;
	assign \g57393/_0_  = _w6152_ ;
	assign \g57395/_0_  = _w6171_ ;
	assign \g57396/_0_  = _w6177_ ;
	assign \g57439/_0_  = _w6178_ ;
	assign \g57476/_0_  = _w6197_ ;
	assign \g57477/_0_  = _w6216_ ;
	assign \g57478/_0_  = _w6235_ ;
	assign \g57479/_0_  = _w6241_ ;
	assign \g57480/_0_  = _w6260_ ;
	assign \g57481/_0_  = _w6292_ ;
	assign \g57482/_0_  = _w6324_ ;
	assign \g57483/_0_  = _w6343_ ;
	assign \g57484/_0_  = _w6349_ ;
	assign \g57485/_0_  = _w6355_ ;
	assign \g57486/_0_  = _w6361_ ;
	assign \g57487/_0_  = _w6367_ ;
	assign \g57488/_0_  = _w6386_ ;
	assign \g57489/_0_  = _w6405_ ;
	assign \g57490/_0_  = _w6424_ ;
	assign \g57491/_0_  = _w6430_ ;
	assign \g57492/_0_  = _w6449_ ;
	assign \g57493/_0_  = _w6468_ ;
	assign \g57494/_0_  = _w6487_ ;
	assign \g57495/_0_  = _w6493_ ;
	assign \g57496/_0_  = _w6498_ ;
	assign \g57497/_0_  = _w6513_ ;
	assign \g57498/_0_  = _w6518_ ;
	assign \g57499/_0_  = _w6524_ ;
	assign \g57500/_0_  = _w6530_ ;
	assign \g57501/_0_  = _w6536_ ;
	assign \g57502/_0_  = _w6542_ ;
	assign \g57503/_0_  = _w6548_ ;
	assign \g57504/_0_  = _w6554_ ;
	assign \g57505/_0_  = _w6560_ ;
	assign \g57524/_0_  = _w6561_ ;
	assign \g57537/_0_  = _w6565_ ;
	assign \g57541/_0_  = _w6569_ ;
	assign \g57543/_0_  = _w6573_ ;
	assign \g58163/_0_  = _w6574_ ;
	assign \g58572/_0_  = _w6581_ ;
	assign \g58573/_0_  = _w6588_ ;
	assign \g58574/_0_  = _w6595_ ;
	assign \g58575/_0_  = _w6602_ ;
	assign \g58576/_0_  = _w6609_ ;
	assign \g58577/_0_  = _w6616_ ;
	assign \g58578/_0_  = _w6623_ ;
	assign \g58579/_0_  = _w6630_ ;
	assign \g58580/_0_  = _w6637_ ;
	assign \g58581/_0_  = _w6644_ ;
	assign \g58582/_0_  = _w6651_ ;
	assign \g58583/_0_  = _w6658_ ;
	assign \g58584/_0_  = _w6665_ ;
	assign \g58585/_0_  = _w6672_ ;
	assign \g58586/_0_  = _w6679_ ;
	assign \g58587/_0_  = _w6686_ ;
	assign \g58588/_0_  = _w6693_ ;
	assign \g58589/_0_  = _w6700_ ;
	assign \g58590/_0_  = _w6707_ ;
	assign \g58591/_0_  = _w6714_ ;
	assign \g58592/_0_  = _w6721_ ;
	assign \g58593/_0_  = _w6728_ ;
	assign \g58594/_0_  = _w6735_ ;
	assign \g58595/_0_  = _w6742_ ;
	assign \g58596/_0_  = _w6749_ ;
	assign \g58597/_0_  = _w6756_ ;
	assign \g58598/_0_  = _w6763_ ;
	assign \g58600/_0_  = _w6764_ ;
	assign \g58602/_0_  = _w6765_ ;
	assign \g58604/_0_  = _w6766_ ;
	assign \g58615/_0_  = _w6767_ ;
	assign \g59240/_0_  = _w6771_ ;
	assign \g59241/_0_  = _w6775_ ;
	assign \g59242/_0_  = _w6779_ ;
	assign \g59243/_0_  = _w6783_ ;
	assign \g59244/_0_  = _w6787_ ;
	assign \g59245/_0_  = _w6791_ ;
	assign \g59246/_0_  = _w6795_ ;
	assign \g59247/_0_  = _w6799_ ;
	assign \g59248/_0_  = _w6803_ ;
	assign \g59249/_0_  = _w6807_ ;
	assign \g59250/_0_  = _w6811_ ;
	assign \g59251/_0_  = _w6815_ ;
	assign \g59252/_0_  = _w6819_ ;
	assign \g59253/_0_  = _w6823_ ;
	assign \g59254/_0_  = _w6827_ ;
	assign \g59255/_0_  = _w6831_ ;
	assign \g59256/_0_  = _w6835_ ;
	assign \g59257/_0_  = _w6839_ ;
	assign \g59258/_0_  = _w6843_ ;
	assign \g59259/_0_  = _w6847_ ;
	assign \g59260/_0_  = _w6851_ ;
	assign \g59261/_0_  = _w6855_ ;
	assign \g59262/_0_  = _w6859_ ;
	assign \g59263/_0_  = _w6863_ ;
	assign \g59264/_0_  = _w6867_ ;
	assign \g59265/_0_  = _w6871_ ;
	assign \g59266/_0_  = _w6875_ ;
	assign \g59267/_0_  = _w6879_ ;
	assign \g59268/_0_  = _w6883_ ;
	assign \g59269/_0_  = _w6887_ ;
	assign \g59270/_0_  = _w6891_ ;
	assign \g59271/_0_  = _w6895_ ;
	assign \g59272/_0_  = _w6899_ ;
	assign \g59273/_0_  = _w6903_ ;
	assign \g59274/_0_  = _w6907_ ;
	assign \g59275/_0_  = _w6911_ ;
	assign \g59276/_0_  = _w6915_ ;
	assign \g59277/_0_  = _w6919_ ;
	assign \g59278/_0_  = _w6923_ ;
	assign \g59279/_0_  = _w6927_ ;
	assign \g59280/_0_  = _w6931_ ;
	assign \g59281/_0_  = _w6935_ ;
	assign \g59282/_0_  = _w6939_ ;
	assign \g59283/_0_  = _w6943_ ;
	assign \g59284/_0_  = _w6947_ ;
	assign \g59285/_0_  = _w6951_ ;
	assign \g59286/_0_  = _w6955_ ;
	assign \g59287/_0_  = _w6959_ ;
	assign \g59288/_0_  = _w6963_ ;
	assign \g59289/_0_  = _w6967_ ;
	assign \g59290/_0_  = _w6971_ ;
	assign \g59291/_0_  = _w6975_ ;
	assign \g59292/_0_  = _w6979_ ;
	assign \g59293/_0_  = _w6983_ ;
	assign \g59294/_0_  = _w6987_ ;
	assign \g59295/_0_  = _w6991_ ;
	assign \g59296/_0_  = _w6995_ ;
	assign \g59297/_0_  = _w6999_ ;
	assign \g59298/_0_  = _w7003_ ;
	assign \g59299/_0_  = _w7007_ ;
	assign \g59300/_0_  = _w7011_ ;
	assign \g59301/_0_  = _w7015_ ;
	assign \g59302/_0_  = _w7019_ ;
	assign \g59303/_0_  = _w7023_ ;
	assign \g59304/_0_  = _w7027_ ;
	assign \g59305/_0_  = _w7031_ ;
	assign \g59306/_0_  = _w7035_ ;
	assign \g59307/_0_  = _w7039_ ;
	assign \g59308/_0_  = _w7043_ ;
	assign \g59309/_0_  = _w7047_ ;
	assign \g59310/_0_  = _w7051_ ;
	assign \g59311/_0_  = _w7055_ ;
	assign \g59312/_0_  = _w7059_ ;
	assign \g59313/_0_  = _w7063_ ;
	assign \g59314/_0_  = _w7067_ ;
	assign \g59315/_0_  = _w7071_ ;
	assign \g59316/_0_  = _w7075_ ;
	assign \g59317/_0_  = _w7079_ ;
	assign \g59318/_0_  = _w7083_ ;
	assign \g59319/_0_  = _w7087_ ;
	assign \g59320/_0_  = _w7091_ ;
	assign \g59321/_0_  = _w7095_ ;
	assign \g59322/_0_  = _w7099_ ;
	assign \g59323/_0_  = _w7103_ ;
	assign \g59324/_0_  = _w7107_ ;
	assign \g59325/_0_  = _w7111_ ;
	assign \g59326/_0_  = _w7115_ ;
	assign \g59327/_0_  = _w7119_ ;
	assign \g59328/_0_  = _w7123_ ;
	assign \g59329/_0_  = _w7127_ ;
	assign \g59330/_0_  = _w7131_ ;
	assign \g59331/_0_  = _w7135_ ;
	assign \g59332/_0_  = _w7139_ ;
	assign \g59333/_0_  = _w7143_ ;
	assign \g59334/_0_  = _w7147_ ;
	assign \g59335/_0_  = _w7151_ ;
	assign \g59336/_0_  = _w7155_ ;
	assign \g59337/_0_  = _w7159_ ;
	assign \g59338/_0_  = _w7163_ ;
	assign \g59339/_0_  = _w7167_ ;
	assign \g59340/_0_  = _w7171_ ;
	assign \g59341/_0_  = _w7175_ ;
	assign \g59342/_0_  = _w7179_ ;
	assign \g59343/_0_  = _w7183_ ;
	assign \g59344/_0_  = _w7187_ ;
	assign \g59345/_0_  = _w7191_ ;
	assign \g59346/_0_  = _w7195_ ;
	assign \g59347/_0_  = _w7199_ ;
	assign \g59348/_0_  = _w7203_ ;
	assign \g59349/_0_  = _w7207_ ;
	assign \g59350/_0_  = _w7211_ ;
	assign \g59351/_0_  = _w7215_ ;
	assign \g59352/_0_  = _w7219_ ;
	assign \g59353/_0_  = _w7223_ ;
	assign \g59354/_0_  = _w7227_ ;
	assign \g59355/_0_  = _w7231_ ;
	assign \g59356/_0_  = _w7235_ ;
	assign \g59357/_0_  = _w7239_ ;
	assign \g59358/_0_  = _w7243_ ;
	assign \g59359/_0_  = _w7247_ ;
	assign \g59360/_0_  = _w7251_ ;
	assign \g59361/_0_  = _w7255_ ;
	assign \g59362/_0_  = _w7259_ ;
	assign \g59363/_0_  = _w7263_ ;
	assign \g59364/_0_  = _w7267_ ;
	assign \g59365/_0_  = _w7271_ ;
	assign \g59366/_0_  = _w7275_ ;
	assign \g59367/_0_  = _w7279_ ;
	assign \g59368/_0_  = _w7283_ ;
	assign \g59369/_0_  = _w7287_ ;
	assign \g59370/_0_  = _w7291_ ;
	assign \g59371/_0_  = _w7295_ ;
	assign \g59372/_0_  = _w7299_ ;
	assign \g59373/_0_  = _w7303_ ;
	assign \g59374/_0_  = _w7307_ ;
	assign \g59375/_0_  = _w7311_ ;
	assign \g59376/_0_  = _w7315_ ;
	assign \g59377/_0_  = _w7319_ ;
	assign \g59378/_0_  = _w7323_ ;
	assign \g59379/_0_  = _w7327_ ;
	assign \g59380/_0_  = _w7331_ ;
	assign \g59381/_0_  = _w7335_ ;
	assign \g59382/_0_  = _w7339_ ;
	assign \g59383/_0_  = _w7343_ ;
	assign \g59384/_0_  = _w7347_ ;
	assign \g59385/_0_  = _w7351_ ;
	assign \g59386/_0_  = _w7355_ ;
	assign \g59387/_0_  = _w7359_ ;
	assign \g59388/_0_  = _w7363_ ;
	assign \g59389/_0_  = _w7367_ ;
	assign \g59390/_0_  = _w7371_ ;
	assign \g59391/_0_  = _w7375_ ;
	assign \g59392/_0_  = _w7379_ ;
	assign \g59393/_0_  = _w7383_ ;
	assign \g59394/_0_  = _w7387_ ;
	assign \g59395/_0_  = _w7391_ ;
	assign \g59396/_0_  = _w7395_ ;
	assign \g59397/_0_  = _w7399_ ;
	assign \g59398/_0_  = _w7403_ ;
	assign \g59399/_0_  = _w7407_ ;
	assign \g59400/_0_  = _w7411_ ;
	assign \g59401/_0_  = _w7415_ ;
	assign \g59402/_0_  = _w7419_ ;
	assign \g59403/_0_  = _w7423_ ;
	assign \g59404/_0_  = _w7427_ ;
	assign \g59405/_0_  = _w7431_ ;
	assign \g59406/_0_  = _w7435_ ;
	assign \g59407/_0_  = _w7439_ ;
	assign \g59408/_0_  = _w7443_ ;
	assign \g59409/_0_  = _w7447_ ;
	assign \g59410/_0_  = _w7451_ ;
	assign \g59411/_0_  = _w7455_ ;
	assign \g59412/_0_  = _w7459_ ;
	assign \g59413/_0_  = _w7463_ ;
	assign \g59414/_0_  = _w7467_ ;
	assign \g59415/_0_  = _w7471_ ;
	assign \g59416/_0_  = _w7475_ ;
	assign \g59417/_0_  = _w7479_ ;
	assign \g59418/_0_  = _w7483_ ;
	assign \g59419/_0_  = _w7487_ ;
	assign \g59420/_0_  = _w7491_ ;
	assign \g59421/_0_  = _w7495_ ;
	assign \g59422/_0_  = _w7499_ ;
	assign \g59423/_0_  = _w7503_ ;
	assign \g59424/_0_  = _w7507_ ;
	assign \g59425/_0_  = _w7511_ ;
	assign \g59426/_0_  = _w7515_ ;
	assign \g59427/_0_  = _w7519_ ;
	assign \g59428/_0_  = _w7523_ ;
	assign \g59429/_0_  = _w7527_ ;
	assign \g59430/_0_  = _w7531_ ;
	assign \g59431/_0_  = _w7535_ ;
	assign \g59432/_0_  = _w7539_ ;
	assign \g59433/_0_  = _w7543_ ;
	assign \g59434/_0_  = _w7547_ ;
	assign \g59435/_0_  = _w7551_ ;
	assign \g59436/_0_  = _w7555_ ;
	assign \g59437/_0_  = _w7559_ ;
	assign \g59438/_0_  = _w7563_ ;
	assign \g59439/_0_  = _w7567_ ;
	assign \g59440/_0_  = _w7571_ ;
	assign \g59441/_0_  = _w7575_ ;
	assign \g59442/_0_  = _w7579_ ;
	assign \g59443/_0_  = _w7583_ ;
	assign \g59444/_0_  = _w7587_ ;
	assign \g59445/_0_  = _w7591_ ;
	assign \g59446/_0_  = _w7595_ ;
	assign \g59447/_0_  = _w7599_ ;
	assign \g59448/_0_  = _w7603_ ;
	assign \g59449/_0_  = _w7607_ ;
	assign \g59450/_0_  = _w7611_ ;
	assign \g59451/_0_  = _w7615_ ;
	assign \g59452/_0_  = _w7619_ ;
	assign \g59453/_0_  = _w7623_ ;
	assign \g59454/_0_  = _w7627_ ;
	assign \g59455/_0_  = _w7631_ ;
	assign \g59456/_0_  = _w7635_ ;
	assign \g59457/_0_  = _w7639_ ;
	assign \g59458/_0_  = _w7643_ ;
	assign \g59459/_0_  = _w7647_ ;
	assign \g59460/_0_  = _w7651_ ;
	assign \g59461/_0_  = _w7655_ ;
	assign \g59462/_0_  = _w7659_ ;
	assign \g59463/_0_  = _w7663_ ;
	assign \g59464/_0_  = _w7667_ ;
	assign \g59465/_0_  = _w7671_ ;
	assign \g59466/_0_  = _w7675_ ;
	assign \g59467/_0_  = _w7679_ ;
	assign \g59468/_0_  = _w7683_ ;
	assign \g59469/_0_  = _w7687_ ;
	assign \g59470/_0_  = _w7691_ ;
	assign \g59471/_0_  = _w7695_ ;
	assign \g59472/_0_  = _w7699_ ;
	assign \g59473/_0_  = _w7703_ ;
	assign \g59474/_0_  = _w7707_ ;
	assign \g59475/_0_  = _w7711_ ;
	assign \g59476/_0_  = _w7715_ ;
	assign \g59477/_0_  = _w7719_ ;
	assign \g59478/_0_  = _w7723_ ;
	assign \g59479/_0_  = _w7727_ ;
	assign \g59480/_0_  = _w7731_ ;
	assign \g59481/_0_  = _w7735_ ;
	assign \g59482/_0_  = _w7739_ ;
	assign \g59483/_0_  = _w7743_ ;
	assign \g59484/_0_  = _w7747_ ;
	assign \g59485/_0_  = _w7751_ ;
	assign \g59486/_0_  = _w7755_ ;
	assign \g59487/_0_  = _w7759_ ;
	assign \g59488/_0_  = _w7763_ ;
	assign \g59489/_0_  = _w7767_ ;
	assign \g59490/_0_  = _w7771_ ;
	assign \g59491/_0_  = _w7775_ ;
	assign \g59492/_0_  = _w7779_ ;
	assign \g59493/_0_  = _w7783_ ;
	assign \g59494/_0_  = _w7787_ ;
	assign \g59495/_0_  = _w7791_ ;
	assign \g59496/_0_  = _w7795_ ;
	assign \g59497/_0_  = _w7799_ ;
	assign \g59498/_0_  = _w7800_ ;
	assign \g59500/_0_  = _w7801_ ;
	assign \g59503/_0_  = _w7802_ ;
	assign \g59512/_0_  = _w7803_ ;
	assign \g61336/_0_  = _w7804_ ;
	assign \g61521/_0_  = _w7805_ ;
	assign \g61523/_0_  = _w7806_ ;
	assign \g61524/_0_  = _w7807_ ;
	assign \g61526/_0_  = _w7808_ ;
	assign \g61527/_0_  = _w7809_ ;
	assign \g61528/_0_  = _w7810_ ;
	assign \g61529/_0_  = _w7811_ ;
	assign \g61530/_0_  = _w7812_ ;
	assign \g61531/_0_  = _w7813_ ;
	assign \g61532/_0_  = _w7814_ ;
	assign \g61533/_0_  = _w7815_ ;
	assign \g61535/_0_  = _w7816_ ;
	assign \g61537/_0_  = _w7817_ ;
	assign \g61539/_0_  = _w7818_ ;
	assign \g61540/_0_  = _w7819_ ;
	assign \g61541/_0_  = _w7820_ ;
	assign \g61542/_0_  = _w7821_ ;
	assign \g61546/_0_  = _w7822_ ;
	assign \g61550/_0_  = _w7823_ ;
	assign \g61551/_0_  = _w7824_ ;
	assign \g61552/_0_  = _w7825_ ;
	assign \g61554/_0_  = _w7826_ ;
	assign \g61555/_0_  = _w7827_ ;
	assign \g61556/_0_  = _w7828_ ;
	assign \g61558/_0_  = _w7829_ ;
	assign \g61559/_0_  = _w7830_ ;
	assign \g61561/_0_  = _w7831_ ;
	assign \g61562/_0_  = _w7832_ ;
	assign \g61563/_0_  = _w7833_ ;
	assign \g61564/_0_  = _w7834_ ;
	assign \g61565/_0_  = _w7835_ ;
	assign \g61566/_0_  = _w7836_ ;
	assign \g61568/_0_  = _w7837_ ;
	assign \g61570/_0_  = _w7838_ ;
	assign \g61571/_0_  = _w7839_ ;
	assign \g61572/_0_  = _w7840_ ;
	assign \g61573/_0_  = _w7841_ ;
	assign \g61577/_0_  = _w7842_ ;
	assign \g61578/_0_  = _w7843_ ;
	assign \g61579/_0_  = _w7844_ ;
	assign \g61580/_0_  = _w7845_ ;
	assign \g61581/_0_  = _w7846_ ;
	assign \g61582/_0_  = _w7847_ ;
	assign \g61583/_0_  = _w7848_ ;
	assign \g61584/_0_  = _w7849_ ;
	assign \g61585/_0_  = _w7850_ ;
	assign \g61586/_0_  = _w7851_ ;
	assign \g61587/_0_  = _w7852_ ;
	assign \g61588/_0_  = _w7853_ ;
	assign \g61589/_0_  = _w7854_ ;
	assign \g61591/_0_  = _w7855_ ;
	assign \g61592/_0_  = _w7856_ ;
	assign \g61594/_0_  = _w7857_ ;
	assign \g61595/_0_  = _w7858_ ;
	assign \g61596/_0_  = _w7859_ ;
	assign \g61597/_0_  = _w7860_ ;
	assign \g61598/_0_  = _w7861_ ;
	assign \g61599/_0_  = _w7862_ ;
	assign \g61600/_0_  = _w7863_ ;
	assign \g61601/_0_  = _w7864_ ;
	assign \g61605/_0_  = _w7865_ ;
	assign \g61606/_0_  = _w7866_ ;
	assign \g61607/_0_  = _w7867_ ;
	assign \g61608/_0_  = _w7868_ ;
	assign \g61609/_0_  = _w7869_ ;
	assign \g61610/_0_  = _w7870_ ;
	assign \g61611/_0_  = _w7871_ ;
	assign \g61612/_0_  = _w7872_ ;
	assign \g61613/_0_  = _w7873_ ;
	assign \g61615/_0_  = _w7874_ ;
	assign \g61616/_0_  = _w7875_ ;
	assign \g61617/_0_  = _w7876_ ;
	assign \g61618/_0_  = _w7877_ ;
	assign \g61619/_0_  = _w7878_ ;
	assign \g61620/_0_  = _w7879_ ;
	assign \g61621/_0_  = _w7880_ ;
	assign \g61623/_0_  = _w7881_ ;
	assign \g61624/_0_  = _w7882_ ;
	assign \g61625/_0_  = _w7883_ ;
	assign \g61626/_0_  = _w7884_ ;
	assign \g61627/_0_  = _w7885_ ;
	assign \g61629/_0_  = _w7886_ ;
	assign \g61630/_0_  = _w7887_ ;
	assign \g61631/_0_  = _w7888_ ;
	assign \g61632/_0_  = _w7889_ ;
	assign \g61633/_0_  = _w7890_ ;
	assign \g61634/_0_  = _w7891_ ;
	assign \g61636/_0_  = _w7892_ ;
	assign \g61638/_0_  = _w7893_ ;
	assign \g61639/_0_  = _w7894_ ;
	assign \g61640/_0_  = _w7895_ ;
	assign \g61641/_0_  = _w7896_ ;
	assign \g61642/_0_  = _w7897_ ;
	assign \g61644/_0_  = _w7898_ ;
	assign \g61647/_0_  = _w7899_ ;
	assign \g61648/_0_  = _w7900_ ;
	assign \g61649/_0_  = _w7901_ ;
	assign \g61650/_0_  = _w7902_ ;
	assign \g61653/_0_  = _w7903_ ;
	assign \g61654/_0_  = _w7904_ ;
	assign \g61655/_0_  = _w7905_ ;
	assign \g61656/_0_  = _w7906_ ;
	assign \g61658/_0_  = _w7907_ ;
	assign \g61661/_0_  = _w7908_ ;
	assign \g61662/_0_  = _w7909_ ;
	assign \g61663/_0_  = _w7910_ ;
	assign \g61664/_0_  = _w7911_ ;
	assign \g61666/_0_  = _w7912_ ;
	assign \g61667/_0_  = _w7913_ ;
	assign \g61668/_0_  = _w7914_ ;
	assign \g61670/_0_  = _w7915_ ;
	assign \g61671/_0_  = _w7916_ ;
	assign \g61672/_0_  = _w7917_ ;
	assign \g61673/_0_  = _w7918_ ;
	assign \g61675/_0_  = _w7919_ ;
	assign \g61676/_0_  = _w7920_ ;
	assign \g61680/_0_  = _w7921_ ;
	assign \g61681/_0_  = _w7922_ ;
	assign \g61682/_0_  = _w7923_ ;
	assign \g61683/_0_  = _w7924_ ;
	assign \g61684/_0_  = _w7925_ ;
	assign \g61686/_0_  = _w7926_ ;
	assign \g61687/_0_  = _w7927_ ;
	assign \g61688/_0_  = _w7928_ ;
	assign \g61689/_0_  = _w7929_ ;
	assign \g61690/_0_  = _w7930_ ;
	assign \g61691/_0_  = _w7931_ ;
	assign \g61693/_0_  = _w7932_ ;
	assign \g61694/_0_  = _w7933_ ;
	assign \g61696/_0_  = _w7934_ ;
	assign \g61697/_0_  = _w7935_ ;
	assign \g61698/_0_  = _w7936_ ;
	assign \g61699/_0_  = _w7937_ ;
	assign \g61700/_0_  = _w7938_ ;
	assign \g61701/_0_  = _w7939_ ;
	assign \g61702/_0_  = _w7940_ ;
	assign \g61703/_0_  = _w7941_ ;
	assign \g61704/_0_  = _w7942_ ;
	assign \g61705/_0_  = _w7943_ ;
	assign \g61706/_0_  = _w7944_ ;
	assign \g61707/_0_  = _w7945_ ;
	assign \g61708/_0_  = _w7946_ ;
	assign \g61711/_0_  = _w7947_ ;
	assign \g61712/_0_  = _w7948_ ;
	assign \g61714/_0_  = _w7949_ ;
	assign \g61716/_0_  = _w7950_ ;
	assign \g61717/_0_  = _w7951_ ;
	assign \g61719/_0_  = _w7952_ ;
	assign \g61720/_0_  = _w7953_ ;
	assign \g61721/_0_  = _w7954_ ;
	assign \g61724/_0_  = _w7955_ ;
	assign \g61725/_0_  = _w7956_ ;
	assign \g61728/_0_  = _w7957_ ;
	assign \g61729/_0_  = _w7958_ ;
	assign \g61731/_0_  = _w7959_ ;
	assign \g61732/_0_  = _w7960_ ;
	assign \g61733/_0_  = _w7961_ ;
	assign \g61736/_0_  = _w7962_ ;
	assign \g61737/_0_  = _w7963_ ;
	assign \g61739/_0_  = _w7964_ ;
	assign \g61740/_0_  = _w7965_ ;
	assign \g61741/_0_  = _w7966_ ;
	assign \g61743/_0_  = _w7967_ ;
	assign \g61744/_0_  = _w7968_ ;
	assign \g61745/_0_  = _w7969_ ;
	assign \g61746/_0_  = _w7970_ ;
	assign \g61747/_0_  = _w7971_ ;
	assign \g61748/_0_  = _w7972_ ;
	assign \g61749/_0_  = _w7973_ ;
	assign \g61750/_0_  = _w7974_ ;
	assign \g61751/_0_  = _w7975_ ;
	assign \g61752/_0_  = _w7976_ ;
	assign \g61753/_0_  = _w7977_ ;
	assign \g61754/_0_  = _w7978_ ;
	assign \g61755/_0_  = _w7979_ ;
	assign \g61757/_0_  = _w7980_ ;
	assign \g61758/_0_  = _w7981_ ;
	assign \g61759/_0_  = _w7982_ ;
	assign \g61760/_0_  = _w7983_ ;
	assign \g61761/_0_  = _w7984_ ;
	assign \g61762/_0_  = _w7985_ ;
	assign \g61763/_0_  = _w7986_ ;
	assign \g61764/_0_  = _w7987_ ;
	assign \g61765/_0_  = _w7988_ ;
	assign \g61766/_0_  = _w7989_ ;
	assign \g61767/_0_  = _w7990_ ;
	assign \g61768/_0_  = _w7991_ ;
	assign \g61769/_0_  = _w7992_ ;
	assign \g61770/_0_  = _w7993_ ;
	assign \g61771/_0_  = _w7994_ ;
	assign \g61772/_0_  = _w7995_ ;
	assign \g61773/_0_  = _w7996_ ;
	assign \g61774/_0_  = _w7997_ ;
	assign \g61775/_0_  = _w7998_ ;
	assign \g61776/_0_  = _w7999_ ;
	assign \g61777/_0_  = _w8000_ ;
	assign \g61778/_0_  = _w8001_ ;
	assign \g61780/_0_  = _w8002_ ;
	assign \g61781/_0_  = _w8003_ ;
	assign \g61783/_0_  = _w8004_ ;
	assign \g61784/_0_  = _w8005_ ;
	assign \g61786/_0_  = _w8006_ ;
	assign \g61787/_0_  = _w8007_ ;
	assign \g61790/_0_  = _w8008_ ;
	assign \g61791/_0_  = _w8009_ ;
	assign \g61794/_0_  = _w8010_ ;
	assign \g61795/_0_  = _w8011_ ;
	assign \g61796/_0_  = _w8012_ ;
	assign \g61797/_0_  = _w8013_ ;
	assign \g61798/_0_  = _w8014_ ;
	assign \g61799/_0_  = _w8015_ ;
	assign \g61800/_0_  = _w8016_ ;
	assign \g61801/_0_  = _w8017_ ;
	assign \g61802/_0_  = _w8018_ ;
	assign \g61803/_0_  = _w8019_ ;
	assign \g61805/_0_  = _w8020_ ;
	assign \g61806/_0_  = _w8021_ ;
	assign \g61807/_0_  = _w8022_ ;
	assign \g61808/_0_  = _w8023_ ;
	assign \g61809/_0_  = _w8024_ ;
	assign \g61810/_0_  = _w8025_ ;
	assign \g61811/_0_  = _w8026_ ;
	assign \g61812/_0_  = _w8027_ ;
	assign \g61813/_0_  = _w8028_ ;
	assign \g61816/_0_  = _w8029_ ;
	assign \g61817/_0_  = _w8030_ ;
	assign \g61818/_0_  = _w8031_ ;
	assign \g61820/_0_  = _w8032_ ;
	assign \g61822/_0_  = _w8033_ ;
	assign \g61823/_0_  = _w8034_ ;
	assign \g61825/_0_  = _w8035_ ;
	assign \g61826/_0_  = _w8036_ ;
	assign \g61827/_0_  = _w8037_ ;
	assign \g61828/_0_  = _w8038_ ;
	assign \g61829/_0_  = _w8039_ ;
	assign \g61832/_0_  = _w8040_ ;
	assign \g61834/_0_  = _w8041_ ;
	assign \g61835/_0_  = _w8042_ ;
	assign \g61837/_0_  = _w8043_ ;
	assign \g61838/_0_  = _w8044_ ;
	assign \g61839/_0_  = _w8045_ ;
	assign \g61840/_0_  = _w8046_ ;
	assign \g61844/_0_  = _w8047_ ;
	assign \g61847/_0_  = _w8048_ ;
	assign \g61848/_0_  = _w8049_ ;
	assign \g61849/_0_  = _w8050_ ;
	assign \g61850/_0_  = _w8051_ ;
	assign \g61851/_0_  = _w8052_ ;
	assign \g61853/_0_  = _w8053_ ;
	assign \g61854/_0_  = _w8054_ ;
	assign \g61855/_0_  = _w8055_ ;
	assign \g61856/_0_  = _w8056_ ;
	assign \g61858/_0_  = _w8057_ ;
	assign \g61859/_0_  = _w8058_ ;
	assign \g61861/_0_  = _w8059_ ;
	assign \g61862/_0_  = _w8060_ ;
	assign \g61863/_0_  = _w8061_ ;
	assign \g61864/_0_  = _w8062_ ;
	assign \g61865/_0_  = _w8063_ ;
	assign \g61866/_0_  = _w8064_ ;
	assign \g61867/_0_  = _w8065_ ;
	assign \g61868/_0_  = _w8066_ ;
	assign \g61869/_0_  = _w8067_ ;
	assign \g61870/_0_  = _w8068_ ;
	assign \g61871/_0_  = _w8069_ ;
	assign \g61873/_0_  = _w8070_ ;
	assign \g61874/_0_  = _w8071_ ;
	assign \g61875/_0_  = _w8072_ ;
	assign \g61877/_0_  = _w8073_ ;
	assign \g61878/_0_  = _w8074_ ;
	assign \g61879/_0_  = _w8075_ ;
	assign \g61880/_0_  = _w8076_ ;
	assign \g61881/_0_  = _w8077_ ;
	assign \g61883/_0_  = _w8078_ ;
	assign \g61884/_0_  = _w8079_ ;
	assign \g61886/_0_  = _w8080_ ;
	assign \g61887/_0_  = _w8081_ ;
	assign \g61890/_0_  = _w8082_ ;
	assign \g61891/_0_  = _w8083_ ;
	assign \g61892/_0_  = _w8084_ ;
	assign \g61893/_0_  = _w8085_ ;
	assign \g61894/_0_  = _w8086_ ;
	assign \g61895/_0_  = _w8087_ ;
	assign \g61900/_0_  = _w8088_ ;
	assign \g61901/_0_  = _w8089_ ;
	assign \g61902/_0_  = _w8090_ ;
	assign \g61904/_0_  = _w8091_ ;
	assign \g61905/_0_  = _w8092_ ;
	assign \g61906/_0_  = _w8093_ ;
	assign \g61907/_0_  = _w8094_ ;
	assign \g61914/_0_  = _w8095_ ;
	assign \g61915/_0_  = _w8096_ ;
	assign \g61917/_0_  = _w8097_ ;
	assign \g61919/_0_  = _w8098_ ;
	assign \g61921/_0_  = _w8099_ ;
	assign \g61924/_0_  = _w8100_ ;
	assign \g61925/_0_  = _w8101_ ;
	assign \g61926/_0_  = _w8102_ ;
	assign \g61927/_0_  = _w8103_ ;
	assign \g61928/_0_  = _w8104_ ;
	assign \g61929/_0_  = _w8105_ ;
	assign \g61930/_0_  = _w8106_ ;
	assign \g61931/_0_  = _w8107_ ;
	assign \g61932/_0_  = _w8108_ ;
	assign \g61933/_0_  = _w8109_ ;
	assign \g61934/_0_  = _w8110_ ;
	assign \g61935/_0_  = _w8111_ ;
	assign \g61936/_0_  = _w8112_ ;
	assign \g61937/_0_  = _w8113_ ;
	assign \g61938/_0_  = _w8114_ ;
	assign \g61939/_0_  = _w8115_ ;
	assign \g61943/_0_  = _w8116_ ;
	assign \g61944/_0_  = _w8117_ ;
	assign \g61945/_0_  = _w8118_ ;
	assign \g61947/_0_  = _w8119_ ;
	assign \g61948/_0_  = _w8120_ ;
	assign \g61949/_0_  = _w8121_ ;
	assign \g61950/_0_  = _w8122_ ;
	assign \g61951/_0_  = _w8123_ ;
	assign \g61952/_0_  = _w8124_ ;
	assign \g61953/_0_  = _w8125_ ;
	assign \g61955/_0_  = _w8126_ ;
	assign \g61956/_0_  = _w8127_ ;
	assign \g61957/_0_  = _w8128_ ;
	assign \g61958/_0_  = _w8129_ ;
	assign \g61959/_0_  = _w8130_ ;
	assign \g61960/_0_  = _w8131_ ;
	assign \g61961/_0_  = _w8132_ ;
	assign \g61962/_0_  = _w8133_ ;
	assign \g61963/_0_  = _w8134_ ;
	assign \g61964/_0_  = _w8135_ ;
	assign \g61965/_0_  = _w8136_ ;
	assign \g61966/_0_  = _w8137_ ;
	assign \g61967/_0_  = _w8138_ ;
	assign \g61968/_0_  = _w8139_ ;
	assign \g61969/_0_  = _w8140_ ;
	assign \g61970/_0_  = _w8141_ ;
	assign \g61971/_0_  = _w8142_ ;
	assign \g61972/_0_  = _w8143_ ;
	assign \g61973/_0_  = _w8144_ ;
	assign \g61974/_0_  = _w8145_ ;
	assign \g61976/_0_  = _w8146_ ;
	assign \g61978/_0_  = _w8147_ ;
	assign \g61980/_0_  = _w8148_ ;
	assign \g61981/_0_  = _w8149_ ;
	assign \g61982/_0_  = _w8150_ ;
	assign \g61983/_0_  = _w8151_ ;
	assign \g61984/_0_  = _w8152_ ;
	assign \g61985/_0_  = _w8153_ ;
	assign \g61986/_0_  = _w8154_ ;
	assign \g61987/_0_  = _w8155_ ;
	assign \g61988/_0_  = _w8156_ ;
	assign \g61989/_0_  = _w8157_ ;
	assign \g61990/_0_  = _w8158_ ;
	assign \g61992/_0_  = _w8159_ ;
	assign \g61994/_0_  = _w8160_ ;
	assign \g61995/_0_  = _w8161_ ;
	assign \g61996/_0_  = _w8162_ ;
	assign \g61997/_0_  = _w8163_ ;
	assign \g61998/_0_  = _w8164_ ;
	assign \g62000/_0_  = _w8165_ ;
	assign \g62001/_0_  = _w8166_ ;
	assign \g62002/_0_  = _w8167_ ;
	assign \g62003/_0_  = _w8168_ ;
	assign \g62004/_0_  = _w8169_ ;
	assign \g62005/_0_  = _w8170_ ;
	assign \g62007/_0_  = _w8171_ ;
	assign \g62008/_0_  = _w8172_ ;
	assign \g62009/_0_  = _w8173_ ;
	assign \g62010/_0_  = _w8174_ ;
	assign \g62011/_0_  = _w8175_ ;
	assign \g62012/_0_  = _w8176_ ;
	assign \g62013/_0_  = _w8177_ ;
	assign \g62014/_0_  = _w8178_ ;
	assign \g62015/_0_  = _w8179_ ;
	assign \g62016/_0_  = _w8180_ ;
	assign \g62017/_0_  = _w8181_ ;
	assign \g62018/_0_  = _w8182_ ;
	assign \g62019/_0_  = _w8183_ ;
	assign \g62020/_0_  = _w8184_ ;
	assign \g62021/_0_  = _w8185_ ;
	assign \g62022/_0_  = _w8186_ ;
	assign \g62023/_0_  = _w8187_ ;
	assign \g62024/_0_  = _w8188_ ;
	assign \g62025/_0_  = _w8189_ ;
	assign \g62026/_0_  = _w8190_ ;
	assign \g62027/_0_  = _w8191_ ;
	assign \g62030/_0_  = _w8192_ ;
	assign \g62033/_0_  = _w8193_ ;
	assign \g62034/_0_  = _w8194_ ;
	assign \g62036/_0_  = _w8195_ ;
	assign \g62038/_0_  = _w8196_ ;
	assign \g62041/_0_  = _w8197_ ;
	assign \g62042/_0_  = _w8198_ ;
	assign \g62043/_0_  = _w8199_ ;
	assign \g62044/_0_  = _w8200_ ;
	assign \g62045/_0_  = _w8201_ ;
	assign \g62046/_0_  = _w8202_ ;
	assign \g62047/_0_  = _w8203_ ;
	assign \g62048/_0_  = _w8204_ ;
	assign \g62050/_0_  = _w8205_ ;
	assign \g62051/_0_  = _w8206_ ;
	assign \g62052/_0_  = _w8207_ ;
	assign \g62055/_0_  = _w8208_ ;
	assign \g62057/_0_  = _w8209_ ;
	assign \g62058/_0_  = _w8210_ ;
	assign \g62059/_0_  = _w8211_ ;
	assign \g62060/_0_  = _w8212_ ;
	assign \g62061/_0_  = _w8213_ ;
	assign \g62062/_0_  = _w8214_ ;
	assign \g62064/_0_  = _w8215_ ;
	assign \g62065/_0_  = _w8216_ ;
	assign \g62066/_0_  = _w8217_ ;
	assign \g62067/_0_  = _w8218_ ;
	assign \g62068/_0_  = _w8219_ ;
	assign \g62072/_0_  = _w8220_ ;
	assign \g62073/_0_  = _w8221_ ;
	assign \g62074/_0_  = _w8222_ ;
	assign \g62075/_0_  = _w8223_ ;
	assign \g62076/_0_  = _w8224_ ;
	assign \g62077/_0_  = _w8225_ ;
	assign \g62078/_0_  = _w8226_ ;
	assign \g62080/_0_  = _w8227_ ;
	assign \g62081/_0_  = _w8228_ ;
	assign \g62082/_0_  = _w8229_ ;
	assign \g62084/_0_  = _w8230_ ;
	assign \g62085/_0_  = _w8231_ ;
	assign \g62086/_0_  = _w8232_ ;
	assign \g62087/_0_  = _w8233_ ;
	assign \g62088/_0_  = _w8234_ ;
	assign \g62089/_0_  = _w8235_ ;
	assign \g62090/_0_  = _w8236_ ;
	assign \g62091/_0_  = _w8237_ ;
	assign \g62092/_0_  = _w8238_ ;
	assign \g62094/_0_  = _w8239_ ;
	assign \g62096/_0_  = _w8240_ ;
	assign \g62097/_0_  = _w8241_ ;
	assign \g62098/_0_  = _w8242_ ;
	assign \g62099/_0_  = _w8243_ ;
	assign \g62100/_0_  = _w8244_ ;
	assign \g62101/_0_  = _w8245_ ;
	assign \g62102/_0_  = _w8246_ ;
	assign \g62104/_0_  = _w8247_ ;
	assign \g62106/_0_  = _w8248_ ;
	assign \g62107/_0_  = _w8249_ ;
	assign \g62108/_0_  = _w8250_ ;
	assign \g62110/_0_  = _w8251_ ;
	assign \g62112/_0_  = _w8252_ ;
	assign \g62113/_0_  = _w8253_ ;
	assign \g62114/_0_  = _w8254_ ;
	assign \g62116/_0_  = _w8255_ ;
	assign \g62117/_0_  = _w8256_ ;
	assign \g62118/_0_  = _w8257_ ;
	assign \g62119/_0_  = _w8258_ ;
	assign \g62120/_0_  = _w8259_ ;
	assign \g62121/_0_  = _w8260_ ;
	assign \g62122/_0_  = _w8261_ ;
	assign \g62124/_0_  = _w8262_ ;
	assign \g62126/_0_  = _w8263_ ;
	assign \g62127/_0_  = _w8264_ ;
	assign \g62128/_0_  = _w8265_ ;
	assign \g62129/_0_  = _w8266_ ;
	assign \g62130/_0_  = _w8267_ ;
	assign \g62131/_0_  = _w8268_ ;
	assign \g62132/_0_  = _w8269_ ;
	assign \g62133/_0_  = _w8270_ ;
	assign \g62135/_0_  = _w8271_ ;
	assign \g62136/_0_  = _w8272_ ;
	assign \g62137/_0_  = _w8273_ ;
	assign \g62138/_0_  = _w8274_ ;
	assign \g62140/_0_  = _w8275_ ;
	assign \g62143/_0_  = _w8276_ ;
	assign \g62144/_0_  = _w8277_ ;
	assign \g62149/_0_  = _w8278_ ;
	assign \g62150/_0_  = _w8279_ ;
	assign \g62151/_0_  = _w8280_ ;
	assign \g62153/_0_  = _w8281_ ;
	assign \g62155/_0_  = _w8282_ ;
	assign \g62156/_0_  = _w8283_ ;
	assign \g62158/_0_  = _w8284_ ;
	assign \g62160/_0_  = _w8285_ ;
	assign \g62161/_0_  = _w8286_ ;
	assign \g62162/_0_  = _w8287_ ;
	assign \g62164/_0_  = _w8288_ ;
	assign \g62165/_0_  = _w8289_ ;
	assign \g62166/_0_  = _w8290_ ;
	assign \g62167/_0_  = _w8291_ ;
	assign \g62168/_0_  = _w8292_ ;
	assign \g62169/_0_  = _w8293_ ;
	assign \g62172/_0_  = _w8294_ ;
	assign \g62173/_0_  = _w8295_ ;
	assign \g62175/_0_  = _w8296_ ;
	assign \g62176/_0_  = _w8297_ ;
	assign \g62177/_0_  = _w8298_ ;
	assign \g62178/_0_  = _w8299_ ;
	assign \g62179/_0_  = _w8300_ ;
	assign \g62180/_0_  = _w8301_ ;
	assign \g62181/_0_  = _w8302_ ;
	assign \g62182/_0_  = _w8303_ ;
	assign \g62183/_0_  = _w8304_ ;
	assign \g62184/_0_  = _w8305_ ;
	assign \g62185/_0_  = _w8306_ ;
	assign \g62186/_0_  = _w8307_ ;
	assign \g62188/_0_  = _w8308_ ;
	assign \g62189/_0_  = _w8309_ ;
	assign \g62190/_0_  = _w8310_ ;
	assign \g62191/_0_  = _w8311_ ;
	assign \g62193/_0_  = _w8312_ ;
	assign \g62194/_0_  = _w8313_ ;
	assign \g62195/_0_  = _w8314_ ;
	assign \g62196/_0_  = _w8315_ ;
	assign \g62197/_0_  = _w8316_ ;
	assign \g62200/_0_  = _w8317_ ;
	assign \g62201/_0_  = _w8318_ ;
	assign \g62202/_0_  = _w8319_ ;
	assign \g62203/_0_  = _w8320_ ;
	assign \g62205/_0_  = _w8321_ ;
	assign \g62206/_0_  = _w8322_ ;
	assign \g62207/_0_  = _w8323_ ;
	assign \g62208/_0_  = _w8324_ ;
	assign \g62209/_0_  = _w8325_ ;
	assign \g62210/_0_  = _w8326_ ;
	assign \g62211/_0_  = _w8327_ ;
	assign \g62215/_0_  = _w8328_ ;
	assign \g62218/_0_  = _w8329_ ;
	assign \g62219/_0_  = _w8330_ ;
	assign \g62221/_0_  = _w8331_ ;
	assign \g62222/_0_  = _w8332_ ;
	assign \g62223/_0_  = _w8333_ ;
	assign \g62224/_0_  = _w8334_ ;
	assign \g62225/_0_  = _w8335_ ;
	assign \g62226/_0_  = _w8336_ ;
	assign \g62229/_0_  = _w8337_ ;
	assign \g62230/_0_  = _w8338_ ;
	assign \g62231/_0_  = _w8339_ ;
	assign \g62233/_0_  = _w8340_ ;
	assign \g62236/_0_  = _w8341_ ;
	assign \g62237/_0_  = _w8342_ ;
	assign \g62238/_0_  = _w8343_ ;
	assign \g62240/_0_  = _w8344_ ;
	assign \g62241/_0_  = _w8345_ ;
	assign \g62243/_0_  = _w8346_ ;
	assign \g62244/_0_  = _w8347_ ;
	assign \g62245/_0_  = _w8348_ ;
	assign \g62247/_0_  = _w8349_ ;
	assign \g62248/_0_  = _w8350_ ;
	assign \g62250/_0_  = _w8351_ ;
	assign \g62252/_0_  = _w8352_ ;
	assign \g62253/_0_  = _w8353_ ;
	assign \g62255/_0_  = _w8354_ ;
	assign \g62256/_0_  = _w8355_ ;
	assign \g62257/_0_  = _w8356_ ;
	assign \g62258/_0_  = _w8357_ ;
	assign \g62259/_0_  = _w8358_ ;
	assign \g62260/_0_  = _w8359_ ;
	assign \g62261/_0_  = _w8360_ ;
	assign \g62262/_0_  = _w8361_ ;
	assign \g62263/_0_  = _w8362_ ;
	assign \g62264/_0_  = _w8363_ ;
	assign \g62265/_0_  = _w8364_ ;
	assign \g62267/_0_  = _w8365_ ;
	assign \g62269/_0_  = _w8366_ ;
	assign \g62270/_0_  = _w8367_ ;
	assign \g62272/_0_  = _w8368_ ;
	assign \g62274/_0_  = _w8369_ ;
	assign \g62277/_0_  = _w8370_ ;
	assign \g62279/_0_  = _w8371_ ;
	assign \g62280/_0_  = _w8372_ ;
	assign \g62281/_0_  = _w8373_ ;
	assign \g62283/_0_  = _w8374_ ;
	assign \g62284/_0_  = _w8375_ ;
	assign \g62285/_0_  = _w8376_ ;
	assign \g62286/_0_  = _w8377_ ;
	assign \g62288/_0_  = _w8378_ ;
	assign \g62289/_0_  = _w8379_ ;
	assign \g62290/_0_  = _w8380_ ;
	assign \g62294/_0_  = _w8381_ ;
	assign \g62295/_0_  = _w8382_ ;
	assign \g62296/_0_  = _w8383_ ;
	assign \g62297/_0_  = _w8384_ ;
	assign \g62298/_0_  = _w8385_ ;
	assign \g62299/_0_  = _w8386_ ;
	assign \g62303/_0_  = _w8387_ ;
	assign \g62305/_0_  = _w8388_ ;
	assign \g62306/_0_  = _w8389_ ;
	assign \g62307/_0_  = _w8390_ ;
	assign \g62309/_0_  = _w8391_ ;
	assign \g62311/_0_  = _w8392_ ;
	assign \g62312/_0_  = _w8393_ ;
	assign \g62313/_0_  = _w8394_ ;
	assign \g62314/_0_  = _w8395_ ;
	assign \g62315/_0_  = _w8396_ ;
	assign \g62316/_0_  = _w8397_ ;
	assign \g62317/_0_  = _w8398_ ;
	assign \g62318/_0_  = _w8399_ ;
	assign \g62319/_0_  = _w8400_ ;
	assign \g62320/_0_  = _w8401_ ;
	assign \g62322/_0_  = _w8402_ ;
	assign \g62324/_0_  = _w8403_ ;
	assign \g62325/_0_  = _w8404_ ;
	assign \g62326/_0_  = _w8405_ ;
	assign \g62327/_0_  = _w8406_ ;
	assign \g62329/_0_  = _w8407_ ;
	assign \g62330/_0_  = _w8408_ ;
	assign \g62331/_0_  = _w8409_ ;
	assign \g62332/_0_  = _w8410_ ;
	assign \g62333/_0_  = _w8411_ ;
	assign \g62335/_0_  = _w8412_ ;
	assign \g62336/_0_  = _w8413_ ;
	assign \g62338/_0_  = _w8414_ ;
	assign \g62341/_0_  = _w8415_ ;
	assign \g62342/_0_  = _w8416_ ;
	assign \g62344/_0_  = _w8417_ ;
	assign \g62345/_0_  = _w8418_ ;
	assign \g62348/_0_  = _w8419_ ;
	assign \g62349/_0_  = _w8420_ ;
	assign \g62350/_0_  = _w8421_ ;
	assign \g62353/_0_  = _w8422_ ;
	assign \g62354/_0_  = _w8423_ ;
	assign \g62355/_0_  = _w8424_ ;
	assign \g62356/_0_  = _w8425_ ;
	assign \g62359/_0_  = _w8426_ ;
	assign \g62362/_0_  = _w8427_ ;
	assign \g62363/_0_  = _w8428_ ;
	assign \g62364/_0_  = _w8429_ ;
	assign \g62365/_0_  = _w8430_ ;
	assign \g62366/_0_  = _w8431_ ;
	assign \g62367/_0_  = _w8432_ ;
	assign \g62368/_0_  = _w8433_ ;
	assign \g62369/_0_  = _w8434_ ;
	assign \g62370/_0_  = _w8435_ ;
	assign \g62371/_0_  = _w8436_ ;
	assign \g62372/_0_  = _w8437_ ;
	assign \g62373/_0_  = _w8438_ ;
	assign \g62374/_0_  = _w8439_ ;
	assign \g62376/_0_  = _w8440_ ;
	assign \g62467/_0_  = _w8441_ ;
	assign \g62468/_0_  = _w8442_ ;
	assign \g62469/_0_  = _w8443_ ;
	assign \g62470/_0_  = _w8444_ ;
	assign \g62471/_0_  = _w8445_ ;
	assign \g62472/_0_  = _w8446_ ;
	assign \g62473/_0_  = _w8447_ ;
	assign \g62474/_0_  = _w8448_ ;
	assign \g62475/_0_  = _w8449_ ;
	assign \g62478/_0_  = _w8450_ ;
	assign \g62480/_0_  = _w8451_ ;
	assign \g62481/_0_  = _w8452_ ;
	assign \g62482/_0_  = _w8453_ ;
	assign \g62483/_0_  = _w8454_ ;
	assign \g62484/_0_  = _w8455_ ;
	assign \g62485/_0_  = _w8456_ ;
	assign \g62486/_0_  = _w8457_ ;
	assign \g62487/_0_  = _w8458_ ;
	assign \g62488/_0_  = _w8459_ ;
	assign \g62489/_0_  = _w8460_ ;
	assign \g62490/_0_  = _w8461_ ;
	assign \g62491/_0_  = _w8462_ ;
	assign \g62492/_0_  = _w8463_ ;
	assign \g62493/_0_  = _w8464_ ;
	assign \g62494/_0_  = _w8465_ ;
	assign \g62495/_0_  = _w8466_ ;
	assign \g62496/_0_  = _w8467_ ;
	assign \g62497/_0_  = _w8468_ ;
	assign \g62498/_0_  = _w8469_ ;
	assign \g62499/_0_  = _w8470_ ;
	assign \g62500/_0_  = _w8471_ ;
	assign \g62501/_0_  = _w8472_ ;
	assign \g62502/_0_  = _w8473_ ;
	assign \g62503/_0_  = _w8474_ ;
	assign \g62504/_0_  = _w8475_ ;
	assign \g62509/_0_  = _w8476_ ;
	assign \g62510/_0_  = _w8477_ ;
	assign \g62511/_0_  = _w8478_ ;
	assign \g62512/_0_  = _w8479_ ;
	assign \g62513/_0_  = _w8480_ ;
	assign \g62514/_0_  = _w8481_ ;
	assign \g62515/_0_  = _w8482_ ;
	assign \g62516/_0_  = _w8483_ ;
	assign \g62517/_0_  = _w8484_ ;
	assign \g62518/_0_  = _w8485_ ;
	assign \g62519/_0_  = _w8486_ ;
	assign \g62520/_0_  = _w8487_ ;
	assign \g62521/_0_  = _w8488_ ;
	assign \g62523/_0_  = _w8489_ ;
	assign \g62526/_0_  = _w8490_ ;
	assign \g62528/_0_  = _w8491_ ;
	assign \g62529/_0_  = _w8492_ ;
	assign \g62531/_0_  = _w8493_ ;
	assign \g62532/_0_  = _w8494_ ;
	assign \g62533/_0_  = _w8495_ ;
	assign \g62534/_0_  = _w8496_ ;
	assign \g62535/_0_  = _w8497_ ;
	assign \g62536/_0_  = _w8498_ ;
	assign \g62537/_0_  = _w8499_ ;
	assign \g62539/_0_  = _w8500_ ;
	assign \g62540/_0_  = _w8501_ ;
	assign \g62541/_0_  = _w8502_ ;
	assign \g62542/_0_  = _w8503_ ;
	assign \g62543/_0_  = _w8504_ ;
	assign \g62544/_0_  = _w8505_ ;
	assign \g62545/_0_  = _w8506_ ;
	assign \g62547/_0_  = _w8507_ ;
	assign \g62548/_0_  = _w8508_ ;
	assign \g62549/_0_  = _w8509_ ;
	assign \g62550/_0_  = _w8510_ ;
	assign \g62551/_0_  = _w8511_ ;
	assign \g62552/_0_  = _w8512_ ;
	assign \g62553/_0_  = _w8513_ ;
	assign \g62554/_0_  = _w8514_ ;
	assign \g62555/_0_  = _w8515_ ;
	assign \g62556/_0_  = _w8516_ ;
	assign \g62557/_0_  = _w8517_ ;
	assign \g62560/_0_  = _w8518_ ;
	assign \g62562/_0_  = _w8519_ ;
	assign \g62563/_0_  = _w8520_ ;
	assign \g62564/_0_  = _w8521_ ;
	assign \g62565/_0_  = _w8522_ ;
	assign \g62566/_0_  = _w8523_ ;
	assign \g62567/_0_  = _w8524_ ;
	assign \g62569/_0_  = _w8525_ ;
	assign \g62570/_0_  = _w8526_ ;
	assign \g62571/_0_  = _w8527_ ;
	assign \g62572/_0_  = _w8528_ ;
	assign \g62573/_0_  = _w8529_ ;
	assign \g62574/_0_  = _w8530_ ;
	assign \g62576/_0_  = _w8531_ ;
	assign \g62577/_0_  = _w8532_ ;
	assign \g62581/_0_  = _w8533_ ;
	assign \g62582/_0_  = _w8534_ ;
	assign \g62584/_0_  = _w8535_ ;
	assign \g62585/_0_  = _w8536_ ;
	assign \g62586/_0_  = _w8537_ ;
	assign \g62588/_0_  = _w8538_ ;
	assign \g62589/_0_  = _w8539_ ;
	assign \g62593/_0_  = _w8540_ ;
	assign \g62594/_0_  = _w8541_ ;
	assign \g62595/_0_  = _w8542_ ;
	assign \g62596/_0_  = _w8543_ ;
	assign \g62597/_0_  = _w8544_ ;
	assign \g62598/_0_  = _w8545_ ;
	assign \g62599/_0_  = _w8546_ ;
	assign \g62600/_0_  = _w8547_ ;
	assign \g62601/_0_  = _w8548_ ;
	assign \g62602/_0_  = _w8549_ ;
	assign \g62603/_0_  = _w8550_ ;
	assign \g62604/_0_  = _w8551_ ;
	assign \g62605/_0_  = _w8552_ ;
	assign \g62606/_0_  = _w8553_ ;
	assign \g62607/_0_  = _w8554_ ;
	assign \g62608/_0_  = _w8555_ ;
	assign \g62609/_0_  = _w8556_ ;
	assign \g62610/_0_  = _w8557_ ;
	assign \g62612/_0_  = _w8558_ ;
	assign \g62613/_0_  = _w8559_ ;
	assign \g62614/_0_  = _w8560_ ;
	assign \g62615/_0_  = _w8561_ ;
	assign \g62617/_0_  = _w8562_ ;
	assign \g62618/_0_  = _w8563_ ;
	assign \g62620/_0_  = _w8564_ ;
	assign \g62621/_0_  = _w8565_ ;
	assign \g62622/_0_  = _w8566_ ;
	assign \g62624/_0_  = _w8567_ ;
	assign \g62625/_0_  = _w8568_ ;
	assign \g62626/_0_  = _w8569_ ;
	assign \g62627/_0_  = _w8570_ ;
	assign \g62629/_0_  = _w8571_ ;
	assign \g62630/_0_  = _w8572_ ;
	assign \g62632/_0_  = _w8573_ ;
	assign \g62633/_0_  = _w8574_ ;
	assign \g62635/_0_  = _w8575_ ;
	assign \g62636/_0_  = _w8576_ ;
	assign \g62637/_0_  = _w8577_ ;
	assign \g62638/_0_  = _w8578_ ;
	assign \g62640/_0_  = _w8579_ ;
	assign \g62641/_0_  = _w8580_ ;
	assign \g62642/_0_  = _w8581_ ;
	assign \g62643/_0_  = _w8582_ ;
	assign \g62644/_0_  = _w8583_ ;
	assign \g62646/_0_  = _w8584_ ;
	assign \g62647/_0_  = _w8585_ ;
	assign \g62649/_0_  = _w8586_ ;
	assign \g62650/_0_  = _w8587_ ;
	assign \g62651/_0_  = _w8588_ ;
	assign \g62653/_0_  = _w8589_ ;
	assign \g62655/_0_  = _w8590_ ;
	assign \g62656/_0_  = _w8591_ ;
	assign \g62657/_0_  = _w8592_ ;
	assign \g62658/_0_  = _w8593_ ;
	assign \g62660/_0_  = _w8594_ ;
	assign \g62661/_0_  = _w8595_ ;
	assign \g62662/_0_  = _w8596_ ;
	assign \g62663/_0_  = _w8597_ ;
	assign \g62664/_0_  = _w8598_ ;
	assign \g62665/_0_  = _w8599_ ;
	assign \g62667/_0_  = _w8600_ ;
	assign \g62669/_0_  = _w8601_ ;
	assign \g62670/_0_  = _w8602_ ;
	assign \g62671/_0_  = _w8603_ ;
	assign \g62672/_0_  = _w8604_ ;
	assign \g62674/_0_  = _w8605_ ;
	assign \g62675/_0_  = _w8606_ ;
	assign \g62676/_0_  = _w8607_ ;
	assign \g62677/_0_  = _w8608_ ;
	assign \g62678/_0_  = _w8609_ ;
	assign \g62679/_0_  = _w8610_ ;
	assign \g62680/_0_  = _w8611_ ;
	assign \g62681/_0_  = _w8612_ ;
	assign \g62682/_0_  = _w8613_ ;
	assign \g62684/_0_  = _w8614_ ;
	assign \g62685/_0_  = _w8615_ ;
	assign \g62686/_0_  = _w8616_ ;
	assign \g62687/_0_  = _w8617_ ;
	assign \g62690/_0_  = _w8618_ ;
	assign \g62693/_0_  = _w8619_ ;
	assign \g62698/_0_  = _w8620_ ;
	assign \g62699/_0_  = _w8621_ ;
	assign \g62700/_0_  = _w8622_ ;
	assign \g62701/_0_  = _w8623_ ;
	assign \g62702/_0_  = _w8624_ ;
	assign \g62703/_0_  = _w8625_ ;
	assign \g62704/_0_  = _w8626_ ;
	assign \g62709/_0_  = _w8627_ ;
	assign \g62710/_0_  = _w8628_ ;
	assign \g62711/_0_  = _w8629_ ;
	assign \g62714/_0_  = _w8630_ ;
	assign \g62715/_0_  = _w8631_ ;
	assign \g62717/_0_  = _w8632_ ;
	assign \g62718/_0_  = _w8633_ ;
	assign \g62719/_0_  = _w8634_ ;
	assign \g62720/_0_  = _w8635_ ;
	assign \g62721/_0_  = _w8636_ ;
	assign \g62723/_0_  = _w8637_ ;
	assign \g62725/_0_  = _w8638_ ;
	assign \g62726/_0_  = _w8639_ ;
	assign \g62729/_0_  = _w8640_ ;
	assign \g62731/_0_  = _w8641_ ;
	assign \g62733/_0_  = _w8642_ ;
	assign \g62738/_0_  = _w8643_ ;
	assign \g62741/_0_  = _w8644_ ;
	assign \g62742/_0_  = _w8645_ ;
	assign \g62744/_0_  = _w8646_ ;
	assign \g62745/_0_  = _w8647_ ;
	assign \g62746/_0_  = _w8648_ ;
	assign \g62747/_0_  = _w8649_ ;
	assign \g62748/_0_  = _w8650_ ;
	assign \g62749/_0_  = _w8651_ ;
	assign \g62753/_0_  = _w8652_ ;
	assign \g62755/_0_  = _w8653_ ;
	assign \g62756/_0_  = _w8654_ ;
	assign \g62758/_0_  = _w8655_ ;
	assign \g62759/_0_  = _w8656_ ;
	assign \g62760/_0_  = _w8657_ ;
	assign \g62761/_0_  = _w8658_ ;
	assign \g62763/_0_  = _w8659_ ;
	assign \g62766/_0_  = _w8660_ ;
	assign \g62767/_0_  = _w8661_ ;
	assign \g62768/_0_  = _w8662_ ;
	assign \g65554/_0_  = _w8668_ ;
	assign \g65561/_0_  = _w8674_ ;
	assign \g65569/_0_  = _w8680_ ;
	assign \g65580/_0_  = _w8686_ ;
	assign \g65599/_0_  = _w8692_ ;
	assign \g65606/_0_  = _w8698_ ;
	assign \g65636/_0_  = _w8704_ ;
	assign \g65864/_0_  = _w8710_ ;
endmodule;