module top( \g1000_reg/NET0131  , \g1001_reg/NET0131  , \g1002_reg/NET0131  , \g1003_reg/NET0131  , \g1004_reg/NET0131  , \g1005_reg/NET0131  , \g1006_reg/NET0131  , \g1007_reg/NET0131  , \g1008_reg/NET0131  , \g1009_reg/NET0131  , \g1010_reg/NET0131  , \g1011_reg/NET0131  , \g1018_reg/NET0131  , \g101_reg/NET0131  , \g1024_reg/NET0131  , \g1030_reg/NET0131  , \g1033_reg/NET0131  , \g1036_reg/NET0131  , \g1038_reg/NET0131  , \g1040_reg/NET0131  , \g1041_reg/NET0131  , \g1045_reg/NET0131  , \g1048_reg/NET0131  , \g1051_reg/NET0131  , \g1053_reg/NET0131  , \g1055_reg/NET0131  , \g1056_reg/NET0131  , \g105_reg/NET0131  , \g1060_reg/NET0131  , \g1063_reg/NET0131  , \g1066_reg/NET0131  , \g1068_reg/NET0131  , \g1070_reg/NET0131  , \g1071_reg/NET0131  , \g1075_reg/NET0131  , \g1078_reg/NET0131  , \g1081_reg/NET0131  , \g1083_reg/NET0131  , \g1085_reg/NET0131  , \g1088_reg/NET0131  , \g1089_reg/NET0131  , \g1090_reg/NET0131  , \g1091_reg/NET0131  , \g1092_reg/NET0131  , \g1095_reg/NET0131  , \g1098_reg/NET0131  , \g109_reg/NET0131  , \g1101_reg/NET0131  , \g1104_reg/NET0131  , \g1107_reg/NET0131  , \g1110_reg/NET0131  , \g1113_reg/NET0131  , \g1114_reg/NET0131  , \g1115_reg/NET0131  , \g1116_reg/NET0131  , \g1119_reg/NET0131  , \g1122_reg/NET0131  , \g1125_reg/NET0131  , \g1128_reg/NET0131  , \g1131_reg/NET0131  , \g1134_reg/NET0131  , \g1135_reg/NET0131  , \g1136_reg/NET0131  , \g1138_reg/NET0131  , \g113_reg/NET0131  , \g1140_reg/NET0131  , \g1151_reg/NET0131  , \g1164_reg/NET0131  , \g1165_reg/NET0131  , \g1166_reg/NET0131  , \g1167_reg/NET0131  , \g1171_reg/NET0131  , \g1173_reg/NET0131  , \g1174_reg/NET0131  , \g1175_reg/NET0131  , \g1176_reg/NET0131  , \g1177_reg/NET0131  , \g117_reg/NET0131  , \g1180_reg/NET0131  , \g1183_reg/NET0131  , \g1186_reg/NET0131  , \g1192_reg/NET0131  , \g1193_reg/NET0131  , \g1196_reg/NET0131  , \g1210_reg/NET0131  , \g1211_reg/NET0131  , \g1215_reg/NET0131  , \g1216_reg/NET0131  , \g1217_reg/NET0131  , \g1218_reg/NET0131  , \g1219_reg/NET0131  , \g121_reg/NET0131  , \g1220_reg/NET0131  , \g1222_reg/NET0131  , \g1223_reg/NET0131  , \g1224_reg/NET0131  , \g1227_reg/NET0131  , \g1228_reg/NET0131  , \g1230_reg/NET0131  , \g1234_reg/NET0131  , \g1240_reg/NET0131  , \g1243_reg/NET0131  , \g1245_reg/NET0131  , \g1249_pad  , \g1251_reg/NET0131  , \g1253_reg/NET0131  , \g1255_reg/NET0131  , \g1257_reg/NET0131  , \g1259_reg/NET0131  , \g125_reg/NET0131  , \g1261_reg/NET0131  , \g1262_reg/NET0131  , \g1263_reg/NET0131  , \g1264_reg/NET0131  , \g1265_reg/NET0131  , \g1266_reg/NET0131  , \g1267_reg/NET0131  , \g1268_reg/NET0131  , \g1269_reg/NET0131  , \g1270_reg/NET0131  , \g1271_reg/NET0131  , \g1272_reg/NET0131  , \g1273_reg/NET0131  , \g1276_reg/NET0131  , \g1279_reg/NET0131  , \g1282_reg/NET0131  , \g1285_reg/NET0131  , \g1288_reg/NET0131  , \g1291_reg/NET0131  , \g1294_reg/NET0131  , \g1297_reg/NET0131  , \g129_reg/NET0131  , \g1300_reg/NET0131  , \g1303_reg/NET0131  , \g1306_reg/NET0131  , \g130_reg/NET0131  , \g1316_reg/NET0131  , \g1319_reg/NET0131  , \g131_reg/NET0131  , \g1326_reg/NET0131  , \g132_reg/NET0131  , \g1332_reg/NET0131  , \g1339_reg/NET0131  , \g133_reg/NET0131  , \g1345_reg/NET0131  , \g1346_reg/NET0131  , \g134_reg/NET0131  , \g1352_reg/NET0131  , \g1358_reg/NET0131  , \g1365_reg/NET0131  , \g1372_reg/NET0131  , \g1378_reg/NET0131  , \g1384_reg/NET0131  , \g1385_reg/NET0131  , \g1386_reg/NET0131  , \g1387_reg/NET0131  , \g1388_reg/NET0131  , \g1389_reg/NET0131  , \g1390_reg/NET0131  , \g1391_reg/NET0131  , \g1392_reg/NET0131  , \g1393_reg/NET0131  , \g1394_reg/NET0131  , \g1395_reg/NET0131  , \g1396_reg/NET0131  , \g1397_reg/NET0131  , \g1398_reg/NET0131  , \g1399_reg/NET0131  , \g1400_reg/NET0131  , \g1401_reg/NET0131  , \g1402_reg/NET0131  , \g1403_reg/NET0131  , \g1404_reg/NET0131  , \g1405_reg/NET0131  , \g1406_reg/NET0131  , \g1407_reg/NET0131  , \g1408_reg/NET0131  , \g1409_reg/NET0131  , \g1410_reg/NET0131  , \g1411_reg/NET0131  , \g1412_reg/NET0131  , \g1413_reg/NET0131  , \g1414_reg/NET0131  , \g1415_reg/NET0131  , \g1416_reg/NET0131  , \g1417_reg/NET0131  , \g1418_reg/NET0131  , \g1419_reg/NET0131  , \g141_reg/NET0131  , \g1420_reg/NET0131  , \g1421_reg/NET0131  , \g1422_reg/NET0131  , \g1423_reg/NET0131  , \g1424_reg/NET0131  , \g1425_reg/NET0131  , \g1426_reg/NET0131  , \g142_reg/NET0131  , \g1430_reg/NET0131  , \g1435_reg/NET0131  , \g1439_reg/NET0131  , \g143_reg/NET0131  , \g1444_reg/NET0131  , \g1448_reg/NET0131  , \g144_reg/NET0131  , \g1453_reg/NET0131  , \g1457_reg/NET0131  , \g145_reg/NET0131  , \g1462_reg/NET0131  , \g1466_reg/NET0131  , \g146_reg/NET0131  , \g1471_reg/NET0131  , \g1476_reg/NET0131  , \g147_reg/NET0131  , \g1481_reg/NET0131  , \g1486_reg/NET0131  , \g148_reg/NET0131  , \g1491_reg/NET0131  , \g1496_reg/NET0131  , \g149_reg/NET0131  , \g1501_reg/NET0131  , \g1506_reg/NET0131  , \g150_reg/NET0131  , \g1511_reg/NET0131  , \g1512_reg/NET0131  , \g1513_reg/NET0131  , \g1514_reg/NET0131  , \g1515_reg/NET0131  , \g1516_reg/NET0131  , \g151_reg/NET0131  , \g1523_reg/NET0131  , \g1524_reg/NET0131  , \g1525_reg/NET0131  , \g1526_reg/NET0131  , \g1527_reg/NET0131  , \g1528_reg/NET0131  , \g1529_reg/NET0131  , \g152_reg/NET0131  , \g1530_reg/NET0131  , \g1531_reg/NET0131  , \g1532_reg/NET0131  , \g1533_reg/NET0131  , \g1534_reg/NET0131  , \g1535_reg/NET0131  , \g1536_reg/NET0131  , \g1537_reg/NET0131  , \g1538_reg/NET0131  , \g1539_reg/NET0131  , \g153_reg/NET0131  , \g1540_reg/NET0131  , \g1541_reg/NET0131  , \g1542_reg/NET0131  , \g1543_reg/NET0131  , \g1544_reg/NET0131  , \g1545_reg/NET0131  , \g1546_reg/NET0131  , \g154_reg/NET0131  , \g1550_reg/NET0131  , \g1551_reg/NET0131  , \g1552_reg/NET0131  , \g1553_reg/NET0131  , \g1554_reg/NET0131  , \g1555_reg/NET0131  , \g1556_reg/NET0131  , \g1557_reg/NET0131  , \g1558_reg/NET0131  , \g1559_reg/NET0131  , \g155_reg/NET0131  , \g1560_reg/NET0131  , \g1561_reg/NET0131  , \g1563_reg/NET0131  , \g1567_reg/NET0131  , \g156_reg/NET0131  , \g1570_reg/NET0131  , \g1573_reg/NET0131  , \g1576_reg/NET0131  , \g1579_reg/NET0131  , \g157_reg/NET0131  , \g1582_reg/NET0131  , \g1585_reg/NET0131  , \g1588_reg/NET0131  , \g158_reg/NET0131  , \g1591_reg/NET0131  , \g1594_reg/NET0131  , \g1597_reg/NET0131  , \g159_reg/NET0131  , \g1600_reg/NET0131  , \g1603_reg/NET0131  , \g1606_reg/NET0131  , \g1609_reg/NET0131  , \g160_reg/NET0131  , \g1612_reg/NET0131  , \g1615_reg/NET0131  , \g1618_reg/NET0131  , \g161_reg/NET0131  , \g1621_reg/NET0131  , \g1624_reg/NET0131  , \g1627_reg/NET0131  , \g16297_pad  , \g162_reg/NET0131  , \g1630_reg/NET0131  , \g1633_reg/NET0131  , \g16355_pad  , \g1636_reg/NET0131  , \g16399_pad  , \g1639_reg/NET0131  , \g163_reg/NET0131  , \g1642_reg/NET0131  , \g16437_pad  , \g1645_reg/NET0131  , \g1648_reg/NET0131  , \g164_reg/NET0131  , \g1651_reg/NET0131  , \g1654_reg/NET0131  , \g1660_reg/NET0131  , \g1662_reg/NET0131  , \g1664_reg/NET0131  , \g1666_reg/NET0131  , \g1668_reg/NET0131  , \g1670_reg/NET0131  , \g1672_reg/NET0131  , \g1679_reg/NET0131  , \g1680_reg/NET0131  , \g1686_reg/NET0131  , \g168_reg/NET0131  , \g1693_reg/NET0131  , \g1694_reg/NET0131  , \g1695_reg/NET0131  , \g1696_reg/NET0131  , \g1697_reg/NET0131  , \g1698_reg/NET0131  , \g1699_reg/NET0131  , \g169_reg/NET0131  , \g1700_reg/NET0131  , \g1701_reg/NET0131  , \g1702_reg/NET0131  , \g1703_reg/NET0131  , \g1704_reg/NET0131  , \g1705_reg/NET0131  , \g170_reg/NET0131  , \g171_reg/NET0131  , \g1724_reg/NET0131  , \g1727_reg/NET0131  , \g172_reg/NET0131  , \g1730_reg/NET0131  , \g1732_reg/NET0131  , \g1734_reg/NET0131  , \g1735_reg/NET0131  , \g1739_reg/NET0131  , \g173_reg/NET0131  , \g1742_reg/NET0131  , \g1745_reg/NET0131  , \g1747_reg/NET0131  , \g1749_reg/NET0131  , \g174_reg/NET0131  , \g1750_reg/NET0131  , \g1754_reg/NET0131  , \g1757_reg/NET0131  , \g175_reg/NET0131  , \g1760_reg/NET0131  , \g1762_reg/NET0131  , \g1764_reg/NET0131  , \g1765_reg/NET0131  , \g1769_reg/NET0131  , \g176_reg/NET0131  , \g1772_reg/NET0131  , \g1775_reg/NET0131  , \g1777_reg/NET0131  , \g1779_reg/NET0131  , \g177_reg/NET0131  , \g1783_reg/NET0131  , \g1784_reg/NET0131  , \g1785_reg/NET0131  , \g1789_reg/NET0131  , \g178_reg/NET0131  , \g1792_reg/NET0131  , \g1795_reg/NET0131  , \g1798_reg/NET0131  , \g179_reg/NET0131  , \g1801_reg/NET0131  , \g1804_reg/NET0131  , \g1807_reg/NET0131  , \g1808_reg/NET0131  , \g1809_reg/NET0131  , \g1810_reg/NET0131  , \g1813_reg/NET0131  , \g1816_reg/NET0131  , \g1819_reg/NET0131  , \g1822_reg/NET0131  , \g1825_reg/NET0131  , \g1828_reg/NET0131  , \g1829_reg/NET0131  , \g1830_reg/NET0131  , \g1832_reg/NET0131  , \g1834_reg/NET0131  , \g1845_reg/NET0131  , \g1846_reg/NET0131  , \g1849_reg/NET0131  , \g1852_reg/NET0131  , \g1858_reg/NET0131  , \g1859_reg/NET0131  , \g185_reg/NET0131  , \g1860_reg/NET0131  , \g1861_reg/NET0131  , \g1865_reg/NET0131  , \g1867_reg/NET0131  , \g1868_reg/NET0131  , \g1869_reg/NET0131  , \g186_reg/NET0131  , \g1870_reg/NET0131  , \g1871_reg/NET0131  , \g1874_reg/NET0131  , \g1877_reg/NET0131  , \g1880_reg/NET0131  , \g1886_reg/NET0131  , \g1887_reg/NET0131  , \g189_reg/NET0131  , \g1904_reg/NET0131  , \g1905_reg/NET0131  , \g1909_reg/NET0131  , \g1910_reg/NET0131  , \g1911_reg/NET0131  , \g1912_reg/NET0131  , \g1913_reg/NET0131  , \g1914_reg/NET0131  , \g1916_reg/NET0131  , \g1917_reg/NET0131  , \g1918_reg/NET0131  , \g1921_reg/NET0131  , \g1922_reg/NET0131  , \g1924_reg/NET0131  , \g1928_reg/NET0131  , \g192_reg/NET0131  , \g1939_reg/NET0131  , \g1943_pad  , \g1945_reg/NET0131  , \g1947_reg/NET0131  , \g1949_reg/NET0131  , \g1951_reg/NET0131  , \g1953_reg/NET0131  , \g1955_reg/NET0131  , \g1956_reg/NET0131  , \g1957_reg/NET0131  , \g1958_reg/NET0131  , \g1959_reg/NET0131  , \g195_reg/NET0131  , \g1960_reg/NET0131  , \g1961_reg/NET0131  , \g1962_reg/NET0131  , \g1963_reg/NET0131  , \g1964_reg/NET0131  , \g1965_reg/NET0131  , \g1966_reg/NET0131  , \g1967_reg/NET0131  , \g1970_reg/NET0131  , \g1973_reg/NET0131  , \g1976_reg/NET0131  , \g1979_reg/NET0131  , \g1982_reg/NET0131  , \g1985_reg/NET0131  , \g1988_reg/NET0131  , \g198_reg/NET0131  , \g1991_reg/NET0131  , \g1994_reg/NET0131  , \g1997_reg/NET0131  , \g2000_reg/NET0131  , \g201_reg/NET0131  , \g204_reg/NET0131  , \g2078_reg/NET0131  , \g2079_reg/NET0131  , \g207_reg/NET0131  , \g2080_reg/NET0131  , \g2081_reg/NET0131  , \g2082_reg/NET0131  , \g2083_reg/NET0131  , \g2084_reg/NET0131  , \g2085_reg/NET0131  , \g2086_reg/NET0131  , \g2087_reg/NET0131  , \g2088_reg/NET0131  , \g2089_reg/NET0131  , \g2090_reg/NET0131  , \g2091_reg/NET0131  , \g2092_reg/NET0131  , \g2093_reg/NET0131  , \g2094_reg/NET0131  , \g2095_reg/NET0131  , \g2096_reg/NET0131  , \g2097_reg/NET0131  , \g2098_reg/NET0131  , \g2099_reg/NET0131  , \g2100_reg/NET0131  , \g2101_reg/NET0131  , \g2102_reg/NET0131  , \g2103_reg/NET0131  , \g2104_reg/NET0131  , \g2105_reg/NET0131  , \g2106_reg/NET0131  , \g2107_reg/NET0131  , \g2108_reg/NET0131  , \g2109_reg/NET0131  , \g210_reg/NET0131  , \g2110_reg/NET0131  , \g2111_reg/NET0131  , \g2112_reg/NET0131  , \g2113_reg/NET0131  , \g2114_reg/NET0131  , \g2115_reg/NET0131  , \g2116_reg/NET0131  , \g2117_reg/NET0131  , \g2118_reg/NET0131  , \g2119_reg/NET0131  , \g213_reg/NET0131  , \g2165_reg/NET0131  , \g216_reg/NET0131  , \g2170_reg/NET0131  , \g2175_reg/NET0131  , \g2180_reg/NET0131  , \g2185_reg/NET0131  , \g2190_reg/NET0131  , \g2195_reg/NET0131  , \g219_reg/NET0131  , \g2200_reg/NET0131  , \g2205_reg/NET0131  , \g2206_reg/NET0131  , \g2207_reg/NET0131  , \g2208_reg/NET0131  , \g2209_reg/NET0131  , \g2210_reg/NET0131  , \g2217_reg/NET0131  , \g2218_reg/NET0131  , \g2219_reg/NET0131  , \g2220_reg/NET0131  , \g2221_reg/NET0131  , \g2222_reg/NET0131  , \g2223_reg/NET0131  , \g2224_reg/NET0131  , \g2225_reg/NET0131  , \g2226_reg/NET0131  , \g2227_reg/NET0131  , \g2228_reg/NET0131  , \g2229_reg/NET0131  , \g222_reg/NET0131  , \g2230_reg/NET0131  , \g2231_reg/NET0131  , \g2232_reg/NET0131  , \g2233_reg/NET0131  , \g2234_reg/NET0131  , \g2235_reg/NET0131  , \g2236_reg/NET0131  , \g2237_reg/NET0131  , \g2238_reg/NET0131  , \g2239_reg/NET0131  , \g2240_reg/NET0131  , \g2244_reg/NET0131  , \g2245_reg/NET0131  , \g2246_reg/NET0131  , \g2247_reg/NET0131  , \g2248_reg/NET0131  , \g2249_reg/NET0131  , \g2250_reg/NET0131  , \g2251_reg/NET0131  , \g2252_reg/NET0131  , \g2253_reg/NET0131  , \g2254_reg/NET0131  , \g2255_reg/NET0131  , \g225_reg/NET0131  , \g2261_reg/NET0131  , \g2264_reg/NET0131  , \g2267_reg/NET0131  , \g2270_reg/NET0131  , \g2273_reg/NET0131  , \g2276_reg/NET0131  , \g2279_reg/NET0131  , \g2282_reg/NET0131  , \g2285_reg/NET0131  , \g2288_reg/NET0131  , \g228_reg/NET0131  , \g2291_reg/NET0131  , \g2294_reg/NET0131  , \g2297_reg/NET0131  , \g2300_reg/NET0131  , \g2303_reg/NET0131  , \g2306_reg/NET0131  , \g2309_reg/NET0131  , \g2312_reg/NET0131  , \g2315_reg/NET0131  , \g2318_reg/NET0131  , \g231_reg/NET0131  , \g2321_reg/NET0131  , \g2324_reg/NET0131  , \g2327_reg/NET0131  , \g2330_reg/NET0131  , \g2333_reg/NET0131  , \g2336_reg/NET0131  , \g2339_reg/NET0131  , \g2342_reg/NET0131  , \g2345_reg/NET0131  , \g2348_reg/NET0131  , \g234_reg/NET0131  , \g2354_reg/NET0131  , \g2356_reg/NET0131  , \g2358_reg/NET0131  , \g2360_reg/NET0131  , \g2362_reg/NET0131  , \g2364_reg/NET0131  , \g2366_reg/NET0131  , \g2373_reg/NET0131  , \g2374_reg/NET0131  , \g237_reg/NET0131  , \g2380_reg/NET0131  , \g2387_reg/NET0131  , \g2388_reg/NET0131  , \g2389_reg/NET0131  , \g2390_reg/NET0131  , \g2391_reg/NET0131  , \g2392_reg/NET0131  , \g2393_reg/NET0131  , \g2394_reg/NET0131  , \g2395_reg/NET0131  , \g2396_reg/NET0131  , \g2397_reg/NET0131  , \g2398_reg/NET0131  , \g2399_reg/NET0131  , \g240_reg/NET0131  , \g2418_reg/NET0131  , \g2421_reg/NET0131  , \g2424_reg/NET0131  , \g2426_reg/NET0131  , \g2428_reg/NET0131  , \g2429_reg/NET0131  , \g2433_reg/NET0131  , \g2436_reg/NET0131  , \g2439_reg/NET0131  , \g243_reg/NET0131  , \g2441_reg/NET0131  , \g2443_reg/NET0131  , \g2444_reg/NET0131  , \g2448_reg/NET0131  , \g2451_reg/NET0131  , \g2454_reg/NET0131  , \g2456_reg/NET0131  , \g2458_reg/NET0131  , \g2459_reg/NET0131  , \g2463_reg/NET0131  , \g2466_reg/NET0131  , \g2469_reg/NET0131  , \g246_reg/NET0131  , \g2471_reg/NET0131  , \g2473_reg/NET0131  , \g2477_reg/NET0131  , \g2478_reg/NET0131  , \g2479_reg/NET0131  , \g2483_reg/NET0131  , \g2486_reg/NET0131  , \g2489_reg/NET0131  , \g2492_reg/NET0131  , \g2495_reg/NET0131  , \g2498_reg/NET0131  , \g249_reg/NET0131  , \g2501_reg/NET0131  , \g2502_reg/NET0131  , \g2503_reg/NET0131  , \g2504_reg/NET0131  , \g2507_reg/NET0131  , \g2510_reg/NET0131  , \g2513_reg/NET0131  , \g2516_reg/NET0131  , \g2519_reg/NET0131  , \g2522_reg/NET0131  , \g2523_reg/NET0131  , \g2524_reg/NET0131  , \g2526_reg/NET0131  , \g2528_reg/NET0131  , \g252_reg/NET0131  , \g2539_reg/NET0131  , \g2540_reg/NET0131  , \g2543_reg/NET0131  , \g2546_reg/NET0131  , \g2552_reg/NET0131  , \g2553_reg/NET0131  , \g2554_reg/NET0131  , \g2555_reg/NET0131  , \g2559_reg/NET0131  , \g255_reg/NET0131  , \g2561_reg/NET0131  , \g2562_reg/NET0131  , \g2563_reg/NET0131  , \g2564_reg/NET0131  , \g2565_reg/NET0131  , \g2568_reg/NET0131  , \g2571_reg/NET0131  , \g2574_reg/NET0131  , \g2580_reg/NET0131  , \g2581_reg/NET0131  , \g258_reg/NET0131  , \g2598_reg/NET0131  , \g2599_reg/NET0131  , \g2603_reg/NET0131  , \g2604_reg/NET0131  , \g2605_reg/NET0131  , \g2606_reg/NET0131  , \g2607_reg/NET0131  , \g2608_reg/NET0131  , \g2610_reg/NET0131  , \g2611_reg/NET0131  , \g2612_reg/NET0131  , \g2615_reg/NET0131  , \g2616_reg/NET0131  , \g2618_reg/NET0131  , \g261_reg/NET0131  , \g2622_reg/NET0131  , \g2633_reg/NET0131  , \g2637_pad  , \g2639_reg/NET0131  , \g2641_reg/NET0131  , \g2643_reg/NET0131  , \g2645_reg/NET0131  , \g2647_reg/NET0131  , \g2649_reg/NET0131  , \g264_reg/NET0131  , \g2650_reg/NET0131  , \g2651_reg/NET0131  , \g2652_reg/NET0131  , \g2653_reg/NET0131  , \g2654_reg/NET0131  , \g2655_reg/NET0131  , \g2656_reg/NET0131  , \g2657_reg/NET0131  , \g2658_reg/NET0131  , \g2659_reg/NET0131  , \g2660_reg/NET0131  , \g2661_reg/NET0131  , \g2664_reg/NET0131  , \g2667_reg/NET0131  , \g2670_reg/NET0131  , \g2673_reg/NET0131  , \g2676_reg/NET0131  , \g2679_reg/NET0131  , \g267_reg/NET0131  , \g2682_reg/NET0131  , \g2685_reg/NET0131  , \g2688_reg/NET0131  , \g2691_reg/NET0131  , \g2694_reg/NET0131  , \g270_reg/NET0131  , \g273_reg/NET0131  , \g2772_reg/NET0131  , \g2773_reg/NET0131  , \g2774_reg/NET0131  , \g2775_reg/NET0131  , \g2776_reg/NET0131  , \g2777_reg/NET0131  , \g2778_reg/NET0131  , \g2779_reg/NET0131  , \g2780_reg/NET0131  , \g2781_reg/NET0131  , \g2782_reg/NET0131  , \g2783_reg/NET0131  , \g2784_reg/NET0131  , \g2785_reg/NET0131  , \g2786_reg/NET0131  , \g2787_reg/NET0131  , \g2788_reg/NET0131  , \g2789_reg/NET0131  , \g2790_reg/NET0131  , \g2791_reg/NET0131  , \g2792_reg/NET0131  , \g2793_reg/NET0131  , \g2794_reg/NET0131  , \g2795_reg/NET0131  , \g2796_reg/NET0131  , \g2797_reg/NET0131  , \g2798_reg/NET0131  , \g2799_reg/NET0131  , \g279_reg/NET0131  , \g2800_reg/NET0131  , \g2801_reg/NET0131  , \g2802_reg/NET0131  , \g2803_reg/NET0131  , \g2804_reg/NET0131  , \g2805_reg/NET0131  , \g2806_reg/NET0131  , \g2807_reg/NET0131  , \g2808_reg/NET0131  , \g2809_reg/NET0131  , \g2810_reg/NET0131  , \g2811_reg/NET0131  , \g2812_reg/NET0131  , \g2813_reg/NET0131  , \g2814_reg/NET0131  , \g2817_reg/NET0131  , \g281_reg/NET0131  , \g283_reg/NET0131  , \g285_reg/NET0131  , \g2874_reg/NET0131  , \g2879_reg/NET0131  , \g287_reg/NET0131  , \g2883_reg/NET0131  , \g2888_reg/NET0131  , \g2892_reg/NET0131  , \g2896_reg/NET0131  , \g289_reg/NET0131  , \g2900_reg/NET0131  , \g2903_reg/NET0131  , \g2908_reg/NET0131  , \g2912_reg/NET0131  , \g2917_reg/NET0131  , \g291_reg/NET0131  , \g2920_reg/NET0131  , \g2924_reg/NET0131  , \g2929_reg/NET0131  , \g2933_reg/NET0131  , \g2934_reg/NET0131  , \g2935_reg/NET0131  , \g2938_reg/NET0131  , \g2941_reg/NET0131  , \g2944_reg/NET0131  , \g2947_reg/NET0131  , \g2950_reg/NET0131  , \g2953_reg/NET0131  , \g2956_reg/NET0131  , \g2959_reg/NET0131  , \g2962_reg/NET0131  , \g2963_reg/NET0131  , \g2966_reg/NET0131  , \g2969_reg/NET0131  , \g2972_reg/NET0131  , \g2975_reg/NET0131  , \g2978_reg/NET0131  , \g2981_reg/NET0131  , \g2984_reg/NET0131  , \g2985_reg/NET0131  , \g2986_reg/NET0131  , \g2987_reg/NET0131  , \g298_reg/NET0131  , \g2990_reg/NET0131  , \g2991_reg/NET0131  , \g2992_reg/NET0131  , \g2993_reg/NET0131  , \g2997_reg/NET0131  , \g2998_reg/NET0131  , \g299_reg/NET0131  , \g3002_reg/NET0131  , \g3006_reg/NET0131  , \g3010_reg/NET0131  , \g3013_reg/NET0131  , \g3018_reg/NET0131  , \g3024_reg/NET0131  , \g3028_reg/NET0131  , \g3032_reg/NET0131  , \g3036_reg/NET0131  , \g3043_reg/NET0131  , \g3044_reg/NET0131  , \g3045_reg/NET0131  , \g3046_reg/NET0131  , \g3047_reg/NET0131  , \g3048_reg/NET0131  , \g3049_reg/NET0131  , \g3050_reg/NET0131  , \g3051_reg/NET0131  , \g3052_reg/NET0131  , \g3053_reg/NET0131  , \g3054_reg/NET0131  , \g3055_reg/NET0131  , \g3056_reg/NET0131  , \g3057_reg/NET0131  , \g3058_reg/NET0131  , \g3059_reg/NET0131  , \g305_reg/NET0131  , \g3060_reg/NET0131  , \g3061_reg/NET0131  , \g3062_reg/NET0131  , \g3063_reg/NET0131  , \g3064_reg/NET0131  , \g3065_reg/NET0131  , \g3066_reg/NET0131  , \g3067_reg/NET0131  , \g3068_reg/NET0131  , \g3069_reg/NET0131  , \g3070_reg/NET0131  , \g3071_reg/NET0131  , \g3072_reg/NET0131  , \g3073_reg/NET0131  , \g3074_reg/NET0131  , \g3075_reg/NET0131  , \g3076_reg/NET0131  , \g3077_reg/NET0131  , \g3078_reg/NET0131  , \g3079_reg/NET0131  , \g3080_reg/NET0131  , \g3083_reg/NET0131  , \g3097_reg/NET0131  , \g3110_reg/NET0131  , \g3114_reg/NET0131  , \g3120_reg/NET0131  , \g312_reg/NET0131  , \g3139_reg/NET0131  , \g313_reg/NET0131  , \g314_reg/NET0131  , \g315_reg/NET0131  , \g316_reg/NET0131  , \g317_reg/NET0131  , \g318_reg/NET0131  , \g319_reg/NET0131  , \g320_reg/NET0131  , \g321_reg/NET0131  , \g3229_pad  , \g322_reg/NET0131  , \g3230_pad  , \g3231_pad  , \g3233_pad  , \g3234_pad  , \g323_reg/NET0131  , \g324_reg/NET0131  , \g343_reg/NET0131  , \g346_reg/NET0131  , \g349_reg/NET0131  , \g351_reg/NET0131  , \g353_reg/NET0131  , \g354_reg/NET0131  , \g358_reg/NET0131  , \g361_reg/NET0131  , \g364_reg/NET0131  , \g366_reg/NET0131  , \g368_reg/NET0131  , \g369_reg/NET0131  , \g373_reg/NET0131  , \g376_reg/NET0131  , \g379_reg/NET0131  , \g381_reg/NET0131  , \g383_reg/NET0131  , \g384_reg/NET0131  , \g388_reg/NET0131  , \g391_reg/NET0131  , \g394_reg/NET0131  , \g396_reg/NET0131  , \g398_reg/NET0131  , \g402_reg/NET0131  , \g403_reg/NET0131  , \g404_reg/NET0131  , \g408_reg/NET0131  , \g411_reg/NET0131  , \g414_reg/NET0131  , \g417_reg/NET0131  , \g420_reg/NET0131  , \g423_reg/NET0131  , \g426_reg/NET0131  , \g427_reg/NET0131  , \g428_reg/NET0131  , \g429_reg/NET0131  , \g432_reg/NET0131  , \g435_reg/NET0131  , \g438_reg/NET0131  , \g441_reg/NET0131  , \g444_reg/NET0131  , \g447_reg/NET0131  , \g448_reg/NET0131  , \g449_reg/NET0131  , \g451_reg/NET0131  , \g453_reg/NET0131  , \g464_reg/NET0131  , \g465_reg/NET0131  , \g468_reg/NET0131  , \g471_reg/NET0131  , \g477_reg/NET0131  , \g478_reg/NET0131  , \g479_reg/NET0131  , \g480_reg/NET0131  , \g484_reg/NET0131  , \g486_reg/NET0131  , \g487_reg/NET0131  , \g488_reg/NET0131  , \g489_reg/NET0131  , \g490_reg/NET0131  , \g493_reg/NET0131  , \g496_reg/NET0131  , \g499_reg/NET0131  , \g506_reg/NET0131  , \g507_reg/NET0131  , \g51_pad  , \g524_reg/NET0131  , \g525_reg/NET0131  , \g529_reg/NET0131  , \g530_reg/NET0131  , \g531_reg/NET0131  , \g532_reg/NET0131  , \g533_reg/NET0131  , \g534_reg/NET0131  , \g536_reg/NET0131  , \g537_reg/NET0131  , \g5388_pad  , \g538_reg/NET0131  , \g541_reg/NET0131  , \g542_reg/NET0131  , \g544_reg/NET0131  , \g548_reg/NET0131  , \g559_reg/NET0131  , \g563_pad  , \g5657_pad  , \g565_reg/NET0131  , \g567_reg/NET0131  , \g569_reg/NET0131  , \g571_reg/NET0131  , \g573_reg/NET0131  , \g575_reg/NET0131  , \g576_reg/NET0131  , \g577_reg/NET0131  , \g578_reg/NET0131  , \g579_reg/NET0131  , \g580_reg/NET0131  , \g581_reg/NET0131  , \g582_reg/NET0131  , \g583_reg/NET0131  , \g584_reg/NET0131  , \g585_reg/NET0131  , \g586_reg/NET0131  , \g587_reg/NET0131  , \g590_reg/NET0131  , \g593_reg/NET0131  , \g596_reg/NET0131  , \g599_reg/NET0131  , \g602_reg/NET0131  , \g605_reg/NET0131  , \g608_reg/NET0131  , \g611_reg/NET0131  , \g614_reg/NET0131  , \g617_reg/NET0131  , \g620_reg/NET0131  , \g698_reg/NET0131  , \g699_reg/NET0131  , \g700_reg/NET0131  , \g701_reg/NET0131  , \g702_reg/NET0131  , \g703_reg/NET0131  , \g704_reg/NET0131  , \g705_reg/NET0131  , \g706_reg/NET0131  , \g707_reg/NET0131  , \g708_reg/NET0131  , \g709_reg/NET0131  , \g710_reg/NET0131  , \g711_reg/NET0131  , \g712_reg/NET0131  , \g713_reg/NET0131  , \g714_reg/NET0131  , \g715_reg/NET0131  , \g716_reg/NET0131  , \g717_reg/NET0131  , \g718_reg/NET0131  , \g719_reg/NET0131  , \g720_reg/NET0131  , \g721_reg/NET0131  , \g722_reg/NET0131  , \g723_reg/NET0131  , \g724_reg/NET0131  , \g725_reg/NET0131  , \g726_reg/NET0131  , \g727_reg/NET0131  , \g728_reg/NET0131  , \g729_reg/NET0131  , \g730_reg/NET0131  , \g731_reg/NET0131  , \g732_reg/NET0131  , \g733_reg/NET0131  , \g734_reg/NET0131  , \g735_reg/NET0131  , \g736_reg/NET0131  , \g737_reg/NET0131  , \g738_reg/NET0131  , \g739_reg/NET0131  , \g785_reg/NET0131  , \g789_reg/NET0131  , \g793_reg/NET0131  , \g7961_pad  , \g797_reg/NET0131  , \g801_reg/NET0131  , \g805_reg/NET0131  , \g809_reg/NET0131  , \g813_reg/NET0131  , \g817_reg/NET0131  , \g818_reg/NET0131  , \g819_reg/NET0131  , \g820_reg/NET0131  , \g821_reg/NET0131  , \g822_reg/NET0131  , \g8259_pad  , \g8260_pad  , \g8261_pad  , \g8262_pad  , \g8263_pad  , \g8264_pad  , \g8265_pad  , \g8266_pad  , \g8268_pad  , \g8269_pad  , \g8270_pad  , \g8271_pad  , \g8272_pad  , \g8273_pad  , \g8274_pad  , \g8275_pad  , \g829_reg/NET0131  , \g830_reg/NET0131  , \g831_reg/NET0131  , \g832_reg/NET0131  , \g833_reg/NET0131  , \g834_reg/NET0131  , \g835_reg/NET0131  , \g836_reg/NET0131  , \g837_reg/NET0131  , \g838_reg/NET0131  , \g839_reg/NET0131  , \g840_reg/NET0131  , \g841_reg/NET0131  , \g842_reg/NET0131  , \g843_reg/NET0131  , \g844_reg/NET0131  , \g845_reg/NET0131  , \g846_reg/NET0131  , \g847_reg/NET0131  , \g848_reg/NET0131  , \g849_reg/NET0131  , \g850_reg/NET0131  , \g851_reg/NET0131  , \g852_reg/NET0131  , \g856_reg/NET0131  , \g857_reg/NET0131  , \g858_reg/NET0131  , \g859_reg/NET0131  , \g860_reg/NET0131  , \g861_reg/NET0131  , \g862_reg/NET0131  , \g863_reg/NET0131  , \g864_reg/NET0131  , \g865_reg/NET0131  , \g866_reg/NET0131  , \g867_reg/NET0131  , \g873_reg/NET0131  , \g876_reg/NET0131  , \g879_reg/NET0131  , \g882_reg/NET0131  , \g885_reg/NET0131  , \g888_reg/NET0131  , \g891_reg/NET0131  , \g894_reg/NET0131  , \g897_reg/NET0131  , \g900_reg/NET0131  , \g903_reg/NET0131  , \g906_reg/NET0131  , \g909_reg/NET0131  , \g912_reg/NET0131  , \g915_reg/NET0131  , \g918_reg/NET0131  , \g921_reg/NET0131  , \g924_reg/NET0131  , \g927_reg/NET0131  , \g930_reg/NET0131  , \g933_reg/NET0131  , \g936_reg/NET0131  , \g939_reg/NET0131  , \g942_reg/NET0131  , \g945_reg/NET0131  , \g948_reg/NET0131  , \g951_reg/NET0131  , \g954_reg/NET0131  , \g957_reg/NET0131  , \g960_reg/NET0131  , \g966_reg/NET0131  , \g968_reg/NET0131  , \g970_reg/NET0131  , \g972_reg/NET0131  , \g974_reg/NET0131  , \g976_reg/NET0131  , \g978_reg/NET0131  , \g97_reg/NET0131  , \g985_reg/NET0131  , \g986_reg/NET0131  , \g992_reg/NET0131  , \g999_reg/NET0131  , \_al_n0  , \_al_n1  , \g101_reg/P0001  , \g105_reg/P0001  , \g109_reg/P0001  , \g1138_reg/P0001  , \g113_reg/P0001  , \g1140_reg/P0001  , \g117_reg/P0001  , \g121_reg/P0001  , \g125_reg/P0001  , \g1471_reg/P0001  , \g1476_reg/P0001  , \g1481_reg/P0001  , \g1486_reg/P0001  , \g1491_reg/P0001  , \g1496_reg/P0001  , \g1501_reg/P0001  , \g1506_reg/P0001  , \g16496_pad  , \g1660_reg/P0001  , \g1662_reg/P0001  , \g1664_reg/P0001  , \g1666_reg/P0001  , \g1668_reg/P0001  , \g1670_reg/P0001  , \g1672_reg/P0001  , \g18/_0_  , \g1832_reg/P0001  , \g1834_reg/P0001  , \g2165_reg/P0001  , \g2170_reg/P0001  , \g2175_reg/P0001  , \g2180_reg/P0001  , \g2185_reg/P0001  , \g2190_reg/P0001  , \g2195_reg/P0001  , \g2200_reg/P0001  , \g2354_reg/P0001  , \g2356_reg/P0001  , \g2358_reg/P0001  , \g2360_reg/P0001  , \g2362_reg/P0001  , \g2364_reg/P0001  , \g2366_reg/P0001  , \g2526_reg/P0001  , \g2528_reg/P0001  , \g25489_pad  , \g279_reg/P0001  , \g281_reg/P0001  , \g283_reg/P0001  , \g285_reg/P0001  , \g2879_reg/NET0131_syn_2  , \g287_reg/P0001  , \g289_reg/P0001  , \g291_reg/P0001  , \g451_reg/P0001  , \g453_reg/P0001  , \g59421/_3_  , \g59425/_1_  , \g59435/_0_  , \g59436/_0_  , \g59441/_3_  , \g59442/_0_  , \g59445/_0_  , \g59453/_0_  , \g59462/_3_  , \g59466/_3_  , \g59467/_3_  , \g59468/_3_  , \g59469/_3_  , \g59470/_3_  , \g59471/_3_  , \g59472/_3_  , \g59473/_3_  , \g59489/_0_  , \g59498/_0_  , \g59499/_0_  , \g59500/_0_  , \g59502/_2_  , \g59503/_0_  , \g59505/_2_  , \g59507/_0_  , \g59508/_0_  , \g59533/_3_  , \g59534/_3_  , \g59535/_3_  , \g59536/_3_  , \g59537/_3_  , \g59538/_3_  , \g59539/_3_  , \g59540/_3_  , \g59548/_0_  , \g59550/_0_  , \g59551/_0_  , \g59552/_0_  , \g59554/_0_  , \g59555/_0_  , \g59556/_0_  , \g59557/_0_  , \g59558/_0_  , \g59559/_0_  , \g59560/_0_  , \g59561/_0_  , \g59639/_0_  , \g59694/_2_  , \g59695/_0_  , \g59697/_2_  , \g59698/_0_  , \g59699/_0_  , \g59700/_0_  , \g59705/_0_  , \g59706/_0_  , \g59707/_0_  , \g59708/_0_  , \g59709/_0_  , \g59710/_0_  , \g59711/_0_  , \g59712/_0_  , \g59713/_0_  , \g59714/_0_  , \g59715/_0_  , \g59716/_0_  , \g59717/_0_  , \g59718/_0_  , \g59719/_0_  , \g59720/_0_  , \g59721/_0_  , \g59722/_0_  , \g59723/_0_  , \g59724/_0_  , \g59725/_0_  , \g59726/_0_  , \g59727/_0_  , \g59728/_0_  , \g59729/_0_  , \g59730/_0_  , \g59731/_0_  , \g59732/_0_  , \g59733/_0_  , \g59734/_0_  , \g59735/_0_  , \g59736/_0_  , \g59737/_0_  , \g59738/_0_  , \g59739/_0_  , \g59740/_0_  , \g59741/_0_  , \g59742/_0_  , \g59743/_0_  , \g59744/_0_  , \g59745/_0_  , \g59747/_0_  , \g59748/_0_  , \g59749/_0_  , \g59750/_0_  , \g59751/_0_  , \g59752/_0_  , \g59753/_0_  , \g59754/_0_  , \g59755/_0_  , \g59756/_0_  , \g59757/_0_  , \g59758/_0_  , \g59759/_0_  , \g59760/_0_  , \g59761/_0_  , \g59762/_0_  , \g59763/_0_  , \g59764/_0_  , \g59765/_0_  , \g59766/_0_  , \g59915/_0_  , \g59952/_2_  , \g60046/_0_  , \g60048/_0_  , \g60049/_0_  , \g60051/_0_  , \g60063/_0_  , \g60103/_0_  , \g60104/_0_  , \g60105/_0_  , \g60107/_2_  , \g60108/_0_  , \g60109/_0_  , \g60110/_0_  , \g60112/_2_  , \g60119/_0_  , \g60120/_0_  , \g60121/_0_  , \g60122/_0_  , \g60123/_0_  , \g60124/_0_  , \g60126/_0_  , \g60127/_0_  , \g60128/_0_  , \g60129/_0_  , \g60130/_0_  , \g60135/_0_  , \g60136/_0_  , \g60137/_0_  , \g60138/_0_  , \g60139/_0_  , \g60143/_3_  , \g60144/_0_  , \g60145/_0_  , \g60339/_0_  , \g60404/_0_  , \g60427/_0_  , \g60428/_0_  , \g60429/_0_  , \g60434/_0_  , \g60435/_0_  , \g60437/_0_  , \g60438/_0_  , \g60439/_0_  , \g60440/_0_  , \g60441/_0_  , \g60448/_0_  , \g60451/_0_  , \g60452/_0_  , \g60453/_0_  , \g60459/_0_  , \g60460/_0_  , \g60523/_0_  , \g60534/_0_  , \g60535/_0_  , \g60536/_0_  , \g60585/_0_  , \g60586/_0_  , \g60587/_0_  , \g60588/_0_  , \g60591/_0_  , \g60592/_0_  , \g60599/_0_  , \g60601/_0_  , \g60602/_0_  , \g60603/_0_  , \g60604/_0_  , \g60605/_0_  , \g60606/_0_  , \g60607/_0_  , \g60608/_0_  , \g60609/_0_  , \g60613/_0_  , \g60614/_0_  , \g60615/_0_  , \g60694/_0_  , \g60708/_0_  , \g60709/_0_  , \g60710/_0_  , \g60785/_0_  , \g60787/_0_  , \g60788/_0_  , \g60799/_0_  , \g60801/_0_  , \g60802/_0_  , \g60803/_1__syn_2  , \g60805/_1__syn_2  , \g60806/_1__syn_2  , \g60808/_0_  , \g60810/_0_  , \g60811/_0_  , \g60825/_3_  , \g60896/_0_  , \g60980/_0_  , \g60981/_0_  , \g60985/_0_  , \g60986/_0_  , \g61012/_0_  , \g61013/_0_  , \g61015/_0_  , \g61017/_0_  , \g61122/_0_  , \g61123/_0_  , \g61124/_0_  , \g61125/_0_  , \g61222/_0_  , \g61223/_0_  , \g61224/_0_  , \g61225/_0_  , \g61228/_0_  , \g61229/_0_  , \g61230/_0_  , \g61231/_0_  , \g61281/_0_  , \g61293/_1_  , \g61307/_0__syn_2  , \g61309/_0__syn_2  , \g61310/_0__syn_2  , \g61311/_1_  , \g61312/_1_  , \g61313/_1_  , \g61324/_1_  , \g61325/_1_  , \g61326/_1_  , \g61328/_1_  , \g61329/_1_  , \g61330/_1_  , \g61332/_1_  , \g61333/_1_  , \g61334/_1_  , \g61335/_1_  , \g61336/_0_  , \g61338/_0_  , \g61339/_0_  , \g61340/_0_  , \g61377/_1_  , \g61378/_1_  , \g61379/_1_  , \g61388/_1_  , \g61391/_0_  , \g61394/_1_  , \g61395/_1_  , \g61396/_1_  , \g61398/_1_  , \g61399/_1_  , \g61421/_1_  , \g61422/_1_  , \g61423/_1_  , \g61524/_0_  , \g61525/_0_  , \g61526/_0_  , \g61527/_0_  , \g61528/_0_  , \g61529/_0_  , \g61530/_0_  , \g61531/_0_  , \g61532/_0_  , \g61533/_0_  , \g61534/_0_  , \g61535/_0_  , \g61536/_0_  , \g61537/_0_  , \g61538/_0_  , \g61539/_0_  , \g61540/_0_  , \g61541/_0_  , \g61542/_0_  , \g61543/_0_  , \g61544/_0_  , \g61545/_0_  , \g61546/_0_  , \g61547/_0_  , \g61548/_0_  , \g61549/_0_  , \g61550/_0_  , \g61551/_0_  , \g61552/_0_  , \g61553/_0_  , \g61554/_0_  , \g61555/_0_  , \g61556/_0_  , \g61557/_0_  , \g61558/_0_  , \g61559/_0_  , \g61560/_0_  , \g61561/_0_  , \g61562/_0_  , \g61563/_0_  , \g61564/_0_  , \g61565/_0_  , \g61566/_0_  , \g61620/_0_  , \g61621/_0_  , \g61622/_0_  , \g61623/_0_  , \g61753/_0_  , \g61764/_0_  , \g61786/_0_  , \g61795/_0_  , \g61801/_0_  , \g61803/_0_  , \g61808/_0_  , \g61848/_0_  , \g61850/_0_  , \g61851/_0_  , \g62097/_0_  , \g62102/_0_  , \g62115/_0_  , \g62119/_0_  , \g62130/_1_  , \g62131/_0_  , \g62132/_0_  , \g62139/_1_  , \g62140/_1_  , \g62141/_1_  , \g62144/_0_  , \g62145/_0_  , \g62146/_0_  , \g62147/_0_  , \g62150/_0_  , \g62151/_1_  , \g62152/_0_  , \g62153/_1_  , \g62156/_1_  , \g62157/_0_  , \g62159/_0_  , \g62161/_0_  , \g62187/_1_  , \g62190/_1_  , \g62191/_1_  , \g62192/_1_  , \g62194/_1_  , \g62195/_1_  , \g62196/_1_  , \g62203/_0_  , \g62204/_1_  , \g62207/_0__syn_2  , \g62208/_1_  , \g62209/_1_  , \g62210/_1_  , \g62211/_1_  , \g62212/_1_  , \g62217/_0_  , \g62286/_0_  , \g62287/_0_  , \g62288/_0_  , \g62289/_0_  , \g62290/_0_  , \g62291/_0_  , \g62292/_0_  , \g62435/_0_  , \g62436/_0_  , \g62439/_0_  , \g62456/_0_  , \g62486/_1_  , \g62492/_1_  , \g62494/_0_  , \g62495/_1_  , \g62497/_0_  , \g62537/_0_  , \g62544/_0_  , \g62546/_0_  , \g62547/_0_  , \g62549/_3_  , \g62552/_0_  , \g62554/_0_  , \g62555/_0_  , \g62556/_0_  , \g62558/_0_  , \g62559/_0_  , \g62561/_0_  , \g62562/_0_  , \g62566/_0_  , \g62567/_0_  , \g62568/_0_  , \g62569/_0_  , \g62570/_0_  , \g62571/_0_  , \g62572/_0_  , \g62573/_0_  , \g62574/_0_  , \g62575/_0_  , \g62576/_0_  , \g62577/_0_  , \g62578/_0_  , \g62579/_0_  , \g62580/_0_  , \g62581/_0_  , \g62582/_0_  , \g62583/_0_  , \g62584/_0_  , \g62585/_0_  , \g62586/_0_  , \g62587/_0_  , \g62588/_0_  , \g62589/_0_  , \g62590/_0_  , \g62591/_0_  , \g62592/_0_  , \g62593/_0_  , \g62594/_0_  , \g62595/_0_  , \g62596/_0_  , \g62597/_0_  , \g62602/_0_  , \g62607/_0_  , \g62608/_0_  , \g62609/_0_  , \g62619/_0_  , \g62620/_0_  , \g62621/_0_  , \g62622/_0_  , \g62623/_0_  , \g62624/_0_  , \g62626/_0_  , \g62627/_0_  , \g62628/_0_  , \g62629/_0_  , \g62630/_0_  , \g62631/_0_  , \g62632/_0_  , \g62633/_0_  , \g62634/_0_  , \g62635/_0_  , \g62636/_0_  , \g62637/_0_  , \g62638/_0_  , \g62639/_0_  , \g62640/_0_  , \g62641/_0_  , \g62642/_0_  , \g62643/_0_  , \g62644/_0_  , \g62645/_0_  , \g62646/_0_  , \g62647/_0_  , \g62648/_0_  , \g62649/_0_  , \g62650/_0_  , \g62651/_0_  , \g62652/_0_  , \g62653/_0_  , \g62654/_0_  , \g62655/_0_  , \g62656/_0_  , \g62657/_0_  , \g62658/_0_  , \g62659/_0_  , \g62660/_0_  , \g62661/_0_  , \g62674/_0_  , \g62682/_0_  , \g62683/_0_  , \g62689/_0_  , \g62690/_0_  , \g62691/_0_  , \g62694/_0_  , \g62695/_0_  , \g62696/_0_  , \g62698/_0_  , \g62699/_0_  , \g62700/_0_  , \g62723/_0_  , \g62724/_0_  , \g62725/_0_  , \g62726/_0_  , \g62727/_0_  , \g62728/_0_  , \g62735/_0_  , \g62736/_0_  , \g62737/_0_  , \g62738/_0_  , \g62739/_0_  , \g62740/_0_  , \g62754/_0_  , \g62762/_0_  , \g62763/_0_  , \g62764/_0_  , \g62780/_0_  , \g62781/_0_  , \g62785/_0_  , \g62786/_0_  , \g62787/_0_  , \g62791/_0_  , \g62792/_0_  , \g62794/_0_  , \g62804/_0_  , \g62806/_0_  , \g62807/_0_  , \g62811/_0_  , \g62968/_0_  , \g63005/_0_  , \g63041/_0_  , \g63116/_0_  , \g63157/_0_  , \g63164/_0_  , \g63170/_0_  , \g63189/_0_  , \g63202/_0_  , \g63206/_0_  , \g63207/_0_  , \g63265/_0_  , \g63266/_0_  , \g63269/_0_  , \g63271/_0_  , \g63272/_0_  , \g63273/_0_  , \g63274/_0_  , \g63275/_0_  , \g63276/_0_  , \g63277/_0_  , \g63278/_0_  , \g63280/_0_  , \g63281/_0_  , \g63282/_0_  , \g63283/_0_  , \g63284/_0_  , \g63285/_0_  , \g63286/_0_  , \g63287/_0_  , \g63288/_0_  , \g63289/_0_  , \g63290/_0_  , \g63292/_0_  , \g63293/_0_  , \g63294/_0_  , \g63295/_0_  , \g63296/_0_  , \g63297/_0_  , \g63298/_0_  , \g63299/_0_  , \g63302/_0_  , \g63303/_0_  , \g63304/_0_  , \g63305/_0_  , \g63306/_0_  , \g63307/_0_  , \g63308/_0_  , \g63309/_0_  , \g63310/_0_  , \g63311/_0_  , \g63312/_0_  , \g63313/_0_  , \g63314/_0_  , \g63315/_0_  , \g63316/_0_  , \g63317/_0_  , \g63318/_0_  , \g63319/_0_  , \g63320/_0_  , \g63321/_0_  , \g63322/_0_  , \g63323/_0_  , \g63324/_0_  , \g63325/_0_  , \g63326/_0_  , \g63327/_0_  , \g63328/_0_  , \g63329/_0_  , \g63330/_0_  , \g63331/_0_  , \g63339/_0_  , \g63505/_0_  , \g63525/_0_  , \g63543/_1_  , \g63602/_0_  , \g63653/_0_  , \g63663/_1_  , \g63677/_0_  , \g63694/_0_  , \g63729/_0_  , \g63766/_0_  , \g63771/_1_  , \g63773/_1_  , \g63784/_1_  , \g63964/_0_  , \g63965/_0_  , \g63966/_0_  , \g63967/_0_  , \g64257/_1_  , \g64266/_0_  , \g64275/_0_  , \g64400/_0_  , \g64416/_0_  , \g64470/_3_  , \g64473/_0_  , \g64474/_0_  , \g64475/_0_  , \g64479/_0_  , \g64480/_0_  , \g64481/_0_  , \g64483/_0_  , \g64484/_0_  , \g64485/_0_  , \g64486/_0_  , \g64493/_0_  , \g64494/_0_  , \g64495/_0_  , \g64496/_0_  , \g64505/_3_  , \g64507/_0_  , \g64508/_0_  , \g64510/_0_  , \g64511/_0_  , \g64544/_0_  , \g64545/_0_  , \g64546/_0_  , \g64639/_0_  , \g64641/_0_  , \g64642/_0_  , \g64645/_0_  , \g64650/_0_  , \g64737/_0_  , \g64738/_0_  , \g65066/_0_  , \g65070/_0_  , \g65090/_0_  , \g65102/_0_  , \g65102/_3_  , \g65126/_3_  , \g65147/_3_  , \g65163/_0_  , \g65176/_3_  , \g65178/_0_  , \g65182/_0_  , \g65190/_1_  , \g65191/_0_  , \g65196/_0_  , \g65268/_0_  , \g65275/_0_  , \g65290/_0_  , \g65290/_3_  , \g65291/_0_  , \g65292/_0_  , \g65298/_0_  , \g65298/_3_  , \g65314/_0_  , \g65314/_3_  , \g65319/_3_  , \g65335/_0_  , \g65342/_0_  , \g65348/_0_  , \g65422/_0_  , \g65465/_1_  , \g65469/_1_  , \g65478/_1_  , \g65507/_0_  , \g65548/_0_  , \g65699/_1_  , \g65713/_1_  , \g65835/_0_  , \g65860/_0_  , \g65863/_0_  , \g66094/_1_  , \g66102/_0_  , \g66107/_0_  , \g66130/_3_  , \g66131/_3_  , \g66228/_1_  , \g66348/_1_  , \g66543/_0_  , \g66549/_1_  , \g66640/_3_  , \g66641/_3_  , \g66950/_1_  , \g67111/_0_  , \g67219/_0_  , \g67263/_0_  , \g67909/_1_  , \g68049/_0_  , \g68220/_0_  , \g68413/_0_  , \g68511/_0_  , \g68536/_0_  , \g68543/_1_  , \g68554/_0_  , \g68559/_0_  , \g70915/_0_  , \g71108/_1_  , \g71115/_2_  , \g71244_dup/_0_  , \g71368/_0_  , \g71581/_0_  , \g71720/_0_  , \g785_reg/P0001  , \g789_reg/P0001  , \g797_reg/P0001  , \g809_reg/P0001  , \g813_reg/P0001  , \g966_reg/P0001  , \g968_reg/P0001  , \g970_reg/P0001  , \g972_reg/P0001  , \g974_reg/P0001  , \g976_reg/P0001  , \g978_reg/P0001  );
  input \g1000_reg/NET0131  ;
  input \g1001_reg/NET0131  ;
  input \g1002_reg/NET0131  ;
  input \g1003_reg/NET0131  ;
  input \g1004_reg/NET0131  ;
  input \g1005_reg/NET0131  ;
  input \g1006_reg/NET0131  ;
  input \g1007_reg/NET0131  ;
  input \g1008_reg/NET0131  ;
  input \g1009_reg/NET0131  ;
  input \g1010_reg/NET0131  ;
  input \g1011_reg/NET0131  ;
  input \g1018_reg/NET0131  ;
  input \g101_reg/NET0131  ;
  input \g1024_reg/NET0131  ;
  input \g1030_reg/NET0131  ;
  input \g1033_reg/NET0131  ;
  input \g1036_reg/NET0131  ;
  input \g1038_reg/NET0131  ;
  input \g1040_reg/NET0131  ;
  input \g1041_reg/NET0131  ;
  input \g1045_reg/NET0131  ;
  input \g1048_reg/NET0131  ;
  input \g1051_reg/NET0131  ;
  input \g1053_reg/NET0131  ;
  input \g1055_reg/NET0131  ;
  input \g1056_reg/NET0131  ;
  input \g105_reg/NET0131  ;
  input \g1060_reg/NET0131  ;
  input \g1063_reg/NET0131  ;
  input \g1066_reg/NET0131  ;
  input \g1068_reg/NET0131  ;
  input \g1070_reg/NET0131  ;
  input \g1071_reg/NET0131  ;
  input \g1075_reg/NET0131  ;
  input \g1078_reg/NET0131  ;
  input \g1081_reg/NET0131  ;
  input \g1083_reg/NET0131  ;
  input \g1085_reg/NET0131  ;
  input \g1088_reg/NET0131  ;
  input \g1089_reg/NET0131  ;
  input \g1090_reg/NET0131  ;
  input \g1091_reg/NET0131  ;
  input \g1092_reg/NET0131  ;
  input \g1095_reg/NET0131  ;
  input \g1098_reg/NET0131  ;
  input \g109_reg/NET0131  ;
  input \g1101_reg/NET0131  ;
  input \g1104_reg/NET0131  ;
  input \g1107_reg/NET0131  ;
  input \g1110_reg/NET0131  ;
  input \g1113_reg/NET0131  ;
  input \g1114_reg/NET0131  ;
  input \g1115_reg/NET0131  ;
  input \g1116_reg/NET0131  ;
  input \g1119_reg/NET0131  ;
  input \g1122_reg/NET0131  ;
  input \g1125_reg/NET0131  ;
  input \g1128_reg/NET0131  ;
  input \g1131_reg/NET0131  ;
  input \g1134_reg/NET0131  ;
  input \g1135_reg/NET0131  ;
  input \g1136_reg/NET0131  ;
  input \g1138_reg/NET0131  ;
  input \g113_reg/NET0131  ;
  input \g1140_reg/NET0131  ;
  input \g1151_reg/NET0131  ;
  input \g1164_reg/NET0131  ;
  input \g1165_reg/NET0131  ;
  input \g1166_reg/NET0131  ;
  input \g1167_reg/NET0131  ;
  input \g1171_reg/NET0131  ;
  input \g1173_reg/NET0131  ;
  input \g1174_reg/NET0131  ;
  input \g1175_reg/NET0131  ;
  input \g1176_reg/NET0131  ;
  input \g1177_reg/NET0131  ;
  input \g117_reg/NET0131  ;
  input \g1180_reg/NET0131  ;
  input \g1183_reg/NET0131  ;
  input \g1186_reg/NET0131  ;
  input \g1192_reg/NET0131  ;
  input \g1193_reg/NET0131  ;
  input \g1196_reg/NET0131  ;
  input \g1210_reg/NET0131  ;
  input \g1211_reg/NET0131  ;
  input \g1215_reg/NET0131  ;
  input \g1216_reg/NET0131  ;
  input \g1217_reg/NET0131  ;
  input \g1218_reg/NET0131  ;
  input \g1219_reg/NET0131  ;
  input \g121_reg/NET0131  ;
  input \g1220_reg/NET0131  ;
  input \g1222_reg/NET0131  ;
  input \g1223_reg/NET0131  ;
  input \g1224_reg/NET0131  ;
  input \g1227_reg/NET0131  ;
  input \g1228_reg/NET0131  ;
  input \g1230_reg/NET0131  ;
  input \g1234_reg/NET0131  ;
  input \g1240_reg/NET0131  ;
  input \g1243_reg/NET0131  ;
  input \g1245_reg/NET0131  ;
  input \g1249_pad  ;
  input \g1251_reg/NET0131  ;
  input \g1253_reg/NET0131  ;
  input \g1255_reg/NET0131  ;
  input \g1257_reg/NET0131  ;
  input \g1259_reg/NET0131  ;
  input \g125_reg/NET0131  ;
  input \g1261_reg/NET0131  ;
  input \g1262_reg/NET0131  ;
  input \g1263_reg/NET0131  ;
  input \g1264_reg/NET0131  ;
  input \g1265_reg/NET0131  ;
  input \g1266_reg/NET0131  ;
  input \g1267_reg/NET0131  ;
  input \g1268_reg/NET0131  ;
  input \g1269_reg/NET0131  ;
  input \g1270_reg/NET0131  ;
  input \g1271_reg/NET0131  ;
  input \g1272_reg/NET0131  ;
  input \g1273_reg/NET0131  ;
  input \g1276_reg/NET0131  ;
  input \g1279_reg/NET0131  ;
  input \g1282_reg/NET0131  ;
  input \g1285_reg/NET0131  ;
  input \g1288_reg/NET0131  ;
  input \g1291_reg/NET0131  ;
  input \g1294_reg/NET0131  ;
  input \g1297_reg/NET0131  ;
  input \g129_reg/NET0131  ;
  input \g1300_reg/NET0131  ;
  input \g1303_reg/NET0131  ;
  input \g1306_reg/NET0131  ;
  input \g130_reg/NET0131  ;
  input \g1316_reg/NET0131  ;
  input \g1319_reg/NET0131  ;
  input \g131_reg/NET0131  ;
  input \g1326_reg/NET0131  ;
  input \g132_reg/NET0131  ;
  input \g1332_reg/NET0131  ;
  input \g1339_reg/NET0131  ;
  input \g133_reg/NET0131  ;
  input \g1345_reg/NET0131  ;
  input \g1346_reg/NET0131  ;
  input \g134_reg/NET0131  ;
  input \g1352_reg/NET0131  ;
  input \g1358_reg/NET0131  ;
  input \g1365_reg/NET0131  ;
  input \g1372_reg/NET0131  ;
  input \g1378_reg/NET0131  ;
  input \g1384_reg/NET0131  ;
  input \g1385_reg/NET0131  ;
  input \g1386_reg/NET0131  ;
  input \g1387_reg/NET0131  ;
  input \g1388_reg/NET0131  ;
  input \g1389_reg/NET0131  ;
  input \g1390_reg/NET0131  ;
  input \g1391_reg/NET0131  ;
  input \g1392_reg/NET0131  ;
  input \g1393_reg/NET0131  ;
  input \g1394_reg/NET0131  ;
  input \g1395_reg/NET0131  ;
  input \g1396_reg/NET0131  ;
  input \g1397_reg/NET0131  ;
  input \g1398_reg/NET0131  ;
  input \g1399_reg/NET0131  ;
  input \g1400_reg/NET0131  ;
  input \g1401_reg/NET0131  ;
  input \g1402_reg/NET0131  ;
  input \g1403_reg/NET0131  ;
  input \g1404_reg/NET0131  ;
  input \g1405_reg/NET0131  ;
  input \g1406_reg/NET0131  ;
  input \g1407_reg/NET0131  ;
  input \g1408_reg/NET0131  ;
  input \g1409_reg/NET0131  ;
  input \g1410_reg/NET0131  ;
  input \g1411_reg/NET0131  ;
  input \g1412_reg/NET0131  ;
  input \g1413_reg/NET0131  ;
  input \g1414_reg/NET0131  ;
  input \g1415_reg/NET0131  ;
  input \g1416_reg/NET0131  ;
  input \g1417_reg/NET0131  ;
  input \g1418_reg/NET0131  ;
  input \g1419_reg/NET0131  ;
  input \g141_reg/NET0131  ;
  input \g1420_reg/NET0131  ;
  input \g1421_reg/NET0131  ;
  input \g1422_reg/NET0131  ;
  input \g1423_reg/NET0131  ;
  input \g1424_reg/NET0131  ;
  input \g1425_reg/NET0131  ;
  input \g1426_reg/NET0131  ;
  input \g142_reg/NET0131  ;
  input \g1430_reg/NET0131  ;
  input \g1435_reg/NET0131  ;
  input \g1439_reg/NET0131  ;
  input \g143_reg/NET0131  ;
  input \g1444_reg/NET0131  ;
  input \g1448_reg/NET0131  ;
  input \g144_reg/NET0131  ;
  input \g1453_reg/NET0131  ;
  input \g1457_reg/NET0131  ;
  input \g145_reg/NET0131  ;
  input \g1462_reg/NET0131  ;
  input \g1466_reg/NET0131  ;
  input \g146_reg/NET0131  ;
  input \g1471_reg/NET0131  ;
  input \g1476_reg/NET0131  ;
  input \g147_reg/NET0131  ;
  input \g1481_reg/NET0131  ;
  input \g1486_reg/NET0131  ;
  input \g148_reg/NET0131  ;
  input \g1491_reg/NET0131  ;
  input \g1496_reg/NET0131  ;
  input \g149_reg/NET0131  ;
  input \g1501_reg/NET0131  ;
  input \g1506_reg/NET0131  ;
  input \g150_reg/NET0131  ;
  input \g1511_reg/NET0131  ;
  input \g1512_reg/NET0131  ;
  input \g1513_reg/NET0131  ;
  input \g1514_reg/NET0131  ;
  input \g1515_reg/NET0131  ;
  input \g1516_reg/NET0131  ;
  input \g151_reg/NET0131  ;
  input \g1523_reg/NET0131  ;
  input \g1524_reg/NET0131  ;
  input \g1525_reg/NET0131  ;
  input \g1526_reg/NET0131  ;
  input \g1527_reg/NET0131  ;
  input \g1528_reg/NET0131  ;
  input \g1529_reg/NET0131  ;
  input \g152_reg/NET0131  ;
  input \g1530_reg/NET0131  ;
  input \g1531_reg/NET0131  ;
  input \g1532_reg/NET0131  ;
  input \g1533_reg/NET0131  ;
  input \g1534_reg/NET0131  ;
  input \g1535_reg/NET0131  ;
  input \g1536_reg/NET0131  ;
  input \g1537_reg/NET0131  ;
  input \g1538_reg/NET0131  ;
  input \g1539_reg/NET0131  ;
  input \g153_reg/NET0131  ;
  input \g1540_reg/NET0131  ;
  input \g1541_reg/NET0131  ;
  input \g1542_reg/NET0131  ;
  input \g1543_reg/NET0131  ;
  input \g1544_reg/NET0131  ;
  input \g1545_reg/NET0131  ;
  input \g1546_reg/NET0131  ;
  input \g154_reg/NET0131  ;
  input \g1550_reg/NET0131  ;
  input \g1551_reg/NET0131  ;
  input \g1552_reg/NET0131  ;
  input \g1553_reg/NET0131  ;
  input \g1554_reg/NET0131  ;
  input \g1555_reg/NET0131  ;
  input \g1556_reg/NET0131  ;
  input \g1557_reg/NET0131  ;
  input \g1558_reg/NET0131  ;
  input \g1559_reg/NET0131  ;
  input \g155_reg/NET0131  ;
  input \g1560_reg/NET0131  ;
  input \g1561_reg/NET0131  ;
  input \g1563_reg/NET0131  ;
  input \g1567_reg/NET0131  ;
  input \g156_reg/NET0131  ;
  input \g1570_reg/NET0131  ;
  input \g1573_reg/NET0131  ;
  input \g1576_reg/NET0131  ;
  input \g1579_reg/NET0131  ;
  input \g157_reg/NET0131  ;
  input \g1582_reg/NET0131  ;
  input \g1585_reg/NET0131  ;
  input \g1588_reg/NET0131  ;
  input \g158_reg/NET0131  ;
  input \g1591_reg/NET0131  ;
  input \g1594_reg/NET0131  ;
  input \g1597_reg/NET0131  ;
  input \g159_reg/NET0131  ;
  input \g1600_reg/NET0131  ;
  input \g1603_reg/NET0131  ;
  input \g1606_reg/NET0131  ;
  input \g1609_reg/NET0131  ;
  input \g160_reg/NET0131  ;
  input \g1612_reg/NET0131  ;
  input \g1615_reg/NET0131  ;
  input \g1618_reg/NET0131  ;
  input \g161_reg/NET0131  ;
  input \g1621_reg/NET0131  ;
  input \g1624_reg/NET0131  ;
  input \g1627_reg/NET0131  ;
  input \g16297_pad  ;
  input \g162_reg/NET0131  ;
  input \g1630_reg/NET0131  ;
  input \g1633_reg/NET0131  ;
  input \g16355_pad  ;
  input \g1636_reg/NET0131  ;
  input \g16399_pad  ;
  input \g1639_reg/NET0131  ;
  input \g163_reg/NET0131  ;
  input \g1642_reg/NET0131  ;
  input \g16437_pad  ;
  input \g1645_reg/NET0131  ;
  input \g1648_reg/NET0131  ;
  input \g164_reg/NET0131  ;
  input \g1651_reg/NET0131  ;
  input \g1654_reg/NET0131  ;
  input \g1660_reg/NET0131  ;
  input \g1662_reg/NET0131  ;
  input \g1664_reg/NET0131  ;
  input \g1666_reg/NET0131  ;
  input \g1668_reg/NET0131  ;
  input \g1670_reg/NET0131  ;
  input \g1672_reg/NET0131  ;
  input \g1679_reg/NET0131  ;
  input \g1680_reg/NET0131  ;
  input \g1686_reg/NET0131  ;
  input \g168_reg/NET0131  ;
  input \g1693_reg/NET0131  ;
  input \g1694_reg/NET0131  ;
  input \g1695_reg/NET0131  ;
  input \g1696_reg/NET0131  ;
  input \g1697_reg/NET0131  ;
  input \g1698_reg/NET0131  ;
  input \g1699_reg/NET0131  ;
  input \g169_reg/NET0131  ;
  input \g1700_reg/NET0131  ;
  input \g1701_reg/NET0131  ;
  input \g1702_reg/NET0131  ;
  input \g1703_reg/NET0131  ;
  input \g1704_reg/NET0131  ;
  input \g1705_reg/NET0131  ;
  input \g170_reg/NET0131  ;
  input \g171_reg/NET0131  ;
  input \g1724_reg/NET0131  ;
  input \g1727_reg/NET0131  ;
  input \g172_reg/NET0131  ;
  input \g1730_reg/NET0131  ;
  input \g1732_reg/NET0131  ;
  input \g1734_reg/NET0131  ;
  input \g1735_reg/NET0131  ;
  input \g1739_reg/NET0131  ;
  input \g173_reg/NET0131  ;
  input \g1742_reg/NET0131  ;
  input \g1745_reg/NET0131  ;
  input \g1747_reg/NET0131  ;
  input \g1749_reg/NET0131  ;
  input \g174_reg/NET0131  ;
  input \g1750_reg/NET0131  ;
  input \g1754_reg/NET0131  ;
  input \g1757_reg/NET0131  ;
  input \g175_reg/NET0131  ;
  input \g1760_reg/NET0131  ;
  input \g1762_reg/NET0131  ;
  input \g1764_reg/NET0131  ;
  input \g1765_reg/NET0131  ;
  input \g1769_reg/NET0131  ;
  input \g176_reg/NET0131  ;
  input \g1772_reg/NET0131  ;
  input \g1775_reg/NET0131  ;
  input \g1777_reg/NET0131  ;
  input \g1779_reg/NET0131  ;
  input \g177_reg/NET0131  ;
  input \g1783_reg/NET0131  ;
  input \g1784_reg/NET0131  ;
  input \g1785_reg/NET0131  ;
  input \g1789_reg/NET0131  ;
  input \g178_reg/NET0131  ;
  input \g1792_reg/NET0131  ;
  input \g1795_reg/NET0131  ;
  input \g1798_reg/NET0131  ;
  input \g179_reg/NET0131  ;
  input \g1801_reg/NET0131  ;
  input \g1804_reg/NET0131  ;
  input \g1807_reg/NET0131  ;
  input \g1808_reg/NET0131  ;
  input \g1809_reg/NET0131  ;
  input \g1810_reg/NET0131  ;
  input \g1813_reg/NET0131  ;
  input \g1816_reg/NET0131  ;
  input \g1819_reg/NET0131  ;
  input \g1822_reg/NET0131  ;
  input \g1825_reg/NET0131  ;
  input \g1828_reg/NET0131  ;
  input \g1829_reg/NET0131  ;
  input \g1830_reg/NET0131  ;
  input \g1832_reg/NET0131  ;
  input \g1834_reg/NET0131  ;
  input \g1845_reg/NET0131  ;
  input \g1846_reg/NET0131  ;
  input \g1849_reg/NET0131  ;
  input \g1852_reg/NET0131  ;
  input \g1858_reg/NET0131  ;
  input \g1859_reg/NET0131  ;
  input \g185_reg/NET0131  ;
  input \g1860_reg/NET0131  ;
  input \g1861_reg/NET0131  ;
  input \g1865_reg/NET0131  ;
  input \g1867_reg/NET0131  ;
  input \g1868_reg/NET0131  ;
  input \g1869_reg/NET0131  ;
  input \g186_reg/NET0131  ;
  input \g1870_reg/NET0131  ;
  input \g1871_reg/NET0131  ;
  input \g1874_reg/NET0131  ;
  input \g1877_reg/NET0131  ;
  input \g1880_reg/NET0131  ;
  input \g1886_reg/NET0131  ;
  input \g1887_reg/NET0131  ;
  input \g189_reg/NET0131  ;
  input \g1904_reg/NET0131  ;
  input \g1905_reg/NET0131  ;
  input \g1909_reg/NET0131  ;
  input \g1910_reg/NET0131  ;
  input \g1911_reg/NET0131  ;
  input \g1912_reg/NET0131  ;
  input \g1913_reg/NET0131  ;
  input \g1914_reg/NET0131  ;
  input \g1916_reg/NET0131  ;
  input \g1917_reg/NET0131  ;
  input \g1918_reg/NET0131  ;
  input \g1921_reg/NET0131  ;
  input \g1922_reg/NET0131  ;
  input \g1924_reg/NET0131  ;
  input \g1928_reg/NET0131  ;
  input \g192_reg/NET0131  ;
  input \g1939_reg/NET0131  ;
  input \g1943_pad  ;
  input \g1945_reg/NET0131  ;
  input \g1947_reg/NET0131  ;
  input \g1949_reg/NET0131  ;
  input \g1951_reg/NET0131  ;
  input \g1953_reg/NET0131  ;
  input \g1955_reg/NET0131  ;
  input \g1956_reg/NET0131  ;
  input \g1957_reg/NET0131  ;
  input \g1958_reg/NET0131  ;
  input \g1959_reg/NET0131  ;
  input \g195_reg/NET0131  ;
  input \g1960_reg/NET0131  ;
  input \g1961_reg/NET0131  ;
  input \g1962_reg/NET0131  ;
  input \g1963_reg/NET0131  ;
  input \g1964_reg/NET0131  ;
  input \g1965_reg/NET0131  ;
  input \g1966_reg/NET0131  ;
  input \g1967_reg/NET0131  ;
  input \g1970_reg/NET0131  ;
  input \g1973_reg/NET0131  ;
  input \g1976_reg/NET0131  ;
  input \g1979_reg/NET0131  ;
  input \g1982_reg/NET0131  ;
  input \g1985_reg/NET0131  ;
  input \g1988_reg/NET0131  ;
  input \g198_reg/NET0131  ;
  input \g1991_reg/NET0131  ;
  input \g1994_reg/NET0131  ;
  input \g1997_reg/NET0131  ;
  input \g2000_reg/NET0131  ;
  input \g201_reg/NET0131  ;
  input \g204_reg/NET0131  ;
  input \g2078_reg/NET0131  ;
  input \g2079_reg/NET0131  ;
  input \g207_reg/NET0131  ;
  input \g2080_reg/NET0131  ;
  input \g2081_reg/NET0131  ;
  input \g2082_reg/NET0131  ;
  input \g2083_reg/NET0131  ;
  input \g2084_reg/NET0131  ;
  input \g2085_reg/NET0131  ;
  input \g2086_reg/NET0131  ;
  input \g2087_reg/NET0131  ;
  input \g2088_reg/NET0131  ;
  input \g2089_reg/NET0131  ;
  input \g2090_reg/NET0131  ;
  input \g2091_reg/NET0131  ;
  input \g2092_reg/NET0131  ;
  input \g2093_reg/NET0131  ;
  input \g2094_reg/NET0131  ;
  input \g2095_reg/NET0131  ;
  input \g2096_reg/NET0131  ;
  input \g2097_reg/NET0131  ;
  input \g2098_reg/NET0131  ;
  input \g2099_reg/NET0131  ;
  input \g2100_reg/NET0131  ;
  input \g2101_reg/NET0131  ;
  input \g2102_reg/NET0131  ;
  input \g2103_reg/NET0131  ;
  input \g2104_reg/NET0131  ;
  input \g2105_reg/NET0131  ;
  input \g2106_reg/NET0131  ;
  input \g2107_reg/NET0131  ;
  input \g2108_reg/NET0131  ;
  input \g2109_reg/NET0131  ;
  input \g210_reg/NET0131  ;
  input \g2110_reg/NET0131  ;
  input \g2111_reg/NET0131  ;
  input \g2112_reg/NET0131  ;
  input \g2113_reg/NET0131  ;
  input \g2114_reg/NET0131  ;
  input \g2115_reg/NET0131  ;
  input \g2116_reg/NET0131  ;
  input \g2117_reg/NET0131  ;
  input \g2118_reg/NET0131  ;
  input \g2119_reg/NET0131  ;
  input \g213_reg/NET0131  ;
  input \g2165_reg/NET0131  ;
  input \g216_reg/NET0131  ;
  input \g2170_reg/NET0131  ;
  input \g2175_reg/NET0131  ;
  input \g2180_reg/NET0131  ;
  input \g2185_reg/NET0131  ;
  input \g2190_reg/NET0131  ;
  input \g2195_reg/NET0131  ;
  input \g219_reg/NET0131  ;
  input \g2200_reg/NET0131  ;
  input \g2205_reg/NET0131  ;
  input \g2206_reg/NET0131  ;
  input \g2207_reg/NET0131  ;
  input \g2208_reg/NET0131  ;
  input \g2209_reg/NET0131  ;
  input \g2210_reg/NET0131  ;
  input \g2217_reg/NET0131  ;
  input \g2218_reg/NET0131  ;
  input \g2219_reg/NET0131  ;
  input \g2220_reg/NET0131  ;
  input \g2221_reg/NET0131  ;
  input \g2222_reg/NET0131  ;
  input \g2223_reg/NET0131  ;
  input \g2224_reg/NET0131  ;
  input \g2225_reg/NET0131  ;
  input \g2226_reg/NET0131  ;
  input \g2227_reg/NET0131  ;
  input \g2228_reg/NET0131  ;
  input \g2229_reg/NET0131  ;
  input \g222_reg/NET0131  ;
  input \g2230_reg/NET0131  ;
  input \g2231_reg/NET0131  ;
  input \g2232_reg/NET0131  ;
  input \g2233_reg/NET0131  ;
  input \g2234_reg/NET0131  ;
  input \g2235_reg/NET0131  ;
  input \g2236_reg/NET0131  ;
  input \g2237_reg/NET0131  ;
  input \g2238_reg/NET0131  ;
  input \g2239_reg/NET0131  ;
  input \g2240_reg/NET0131  ;
  input \g2244_reg/NET0131  ;
  input \g2245_reg/NET0131  ;
  input \g2246_reg/NET0131  ;
  input \g2247_reg/NET0131  ;
  input \g2248_reg/NET0131  ;
  input \g2249_reg/NET0131  ;
  input \g2250_reg/NET0131  ;
  input \g2251_reg/NET0131  ;
  input \g2252_reg/NET0131  ;
  input \g2253_reg/NET0131  ;
  input \g2254_reg/NET0131  ;
  input \g2255_reg/NET0131  ;
  input \g225_reg/NET0131  ;
  input \g2261_reg/NET0131  ;
  input \g2264_reg/NET0131  ;
  input \g2267_reg/NET0131  ;
  input \g2270_reg/NET0131  ;
  input \g2273_reg/NET0131  ;
  input \g2276_reg/NET0131  ;
  input \g2279_reg/NET0131  ;
  input \g2282_reg/NET0131  ;
  input \g2285_reg/NET0131  ;
  input \g2288_reg/NET0131  ;
  input \g228_reg/NET0131  ;
  input \g2291_reg/NET0131  ;
  input \g2294_reg/NET0131  ;
  input \g2297_reg/NET0131  ;
  input \g2300_reg/NET0131  ;
  input \g2303_reg/NET0131  ;
  input \g2306_reg/NET0131  ;
  input \g2309_reg/NET0131  ;
  input \g2312_reg/NET0131  ;
  input \g2315_reg/NET0131  ;
  input \g2318_reg/NET0131  ;
  input \g231_reg/NET0131  ;
  input \g2321_reg/NET0131  ;
  input \g2324_reg/NET0131  ;
  input \g2327_reg/NET0131  ;
  input \g2330_reg/NET0131  ;
  input \g2333_reg/NET0131  ;
  input \g2336_reg/NET0131  ;
  input \g2339_reg/NET0131  ;
  input \g2342_reg/NET0131  ;
  input \g2345_reg/NET0131  ;
  input \g2348_reg/NET0131  ;
  input \g234_reg/NET0131  ;
  input \g2354_reg/NET0131  ;
  input \g2356_reg/NET0131  ;
  input \g2358_reg/NET0131  ;
  input \g2360_reg/NET0131  ;
  input \g2362_reg/NET0131  ;
  input \g2364_reg/NET0131  ;
  input \g2366_reg/NET0131  ;
  input \g2373_reg/NET0131  ;
  input \g2374_reg/NET0131  ;
  input \g237_reg/NET0131  ;
  input \g2380_reg/NET0131  ;
  input \g2387_reg/NET0131  ;
  input \g2388_reg/NET0131  ;
  input \g2389_reg/NET0131  ;
  input \g2390_reg/NET0131  ;
  input \g2391_reg/NET0131  ;
  input \g2392_reg/NET0131  ;
  input \g2393_reg/NET0131  ;
  input \g2394_reg/NET0131  ;
  input \g2395_reg/NET0131  ;
  input \g2396_reg/NET0131  ;
  input \g2397_reg/NET0131  ;
  input \g2398_reg/NET0131  ;
  input \g2399_reg/NET0131  ;
  input \g240_reg/NET0131  ;
  input \g2418_reg/NET0131  ;
  input \g2421_reg/NET0131  ;
  input \g2424_reg/NET0131  ;
  input \g2426_reg/NET0131  ;
  input \g2428_reg/NET0131  ;
  input \g2429_reg/NET0131  ;
  input \g2433_reg/NET0131  ;
  input \g2436_reg/NET0131  ;
  input \g2439_reg/NET0131  ;
  input \g243_reg/NET0131  ;
  input \g2441_reg/NET0131  ;
  input \g2443_reg/NET0131  ;
  input \g2444_reg/NET0131  ;
  input \g2448_reg/NET0131  ;
  input \g2451_reg/NET0131  ;
  input \g2454_reg/NET0131  ;
  input \g2456_reg/NET0131  ;
  input \g2458_reg/NET0131  ;
  input \g2459_reg/NET0131  ;
  input \g2463_reg/NET0131  ;
  input \g2466_reg/NET0131  ;
  input \g2469_reg/NET0131  ;
  input \g246_reg/NET0131  ;
  input \g2471_reg/NET0131  ;
  input \g2473_reg/NET0131  ;
  input \g2477_reg/NET0131  ;
  input \g2478_reg/NET0131  ;
  input \g2479_reg/NET0131  ;
  input \g2483_reg/NET0131  ;
  input \g2486_reg/NET0131  ;
  input \g2489_reg/NET0131  ;
  input \g2492_reg/NET0131  ;
  input \g2495_reg/NET0131  ;
  input \g2498_reg/NET0131  ;
  input \g249_reg/NET0131  ;
  input \g2501_reg/NET0131  ;
  input \g2502_reg/NET0131  ;
  input \g2503_reg/NET0131  ;
  input \g2504_reg/NET0131  ;
  input \g2507_reg/NET0131  ;
  input \g2510_reg/NET0131  ;
  input \g2513_reg/NET0131  ;
  input \g2516_reg/NET0131  ;
  input \g2519_reg/NET0131  ;
  input \g2522_reg/NET0131  ;
  input \g2523_reg/NET0131  ;
  input \g2524_reg/NET0131  ;
  input \g2526_reg/NET0131  ;
  input \g2528_reg/NET0131  ;
  input \g252_reg/NET0131  ;
  input \g2539_reg/NET0131  ;
  input \g2540_reg/NET0131  ;
  input \g2543_reg/NET0131  ;
  input \g2546_reg/NET0131  ;
  input \g2552_reg/NET0131  ;
  input \g2553_reg/NET0131  ;
  input \g2554_reg/NET0131  ;
  input \g2555_reg/NET0131  ;
  input \g2559_reg/NET0131  ;
  input \g255_reg/NET0131  ;
  input \g2561_reg/NET0131  ;
  input \g2562_reg/NET0131  ;
  input \g2563_reg/NET0131  ;
  input \g2564_reg/NET0131  ;
  input \g2565_reg/NET0131  ;
  input \g2568_reg/NET0131  ;
  input \g2571_reg/NET0131  ;
  input \g2574_reg/NET0131  ;
  input \g2580_reg/NET0131  ;
  input \g2581_reg/NET0131  ;
  input \g258_reg/NET0131  ;
  input \g2598_reg/NET0131  ;
  input \g2599_reg/NET0131  ;
  input \g2603_reg/NET0131  ;
  input \g2604_reg/NET0131  ;
  input \g2605_reg/NET0131  ;
  input \g2606_reg/NET0131  ;
  input \g2607_reg/NET0131  ;
  input \g2608_reg/NET0131  ;
  input \g2610_reg/NET0131  ;
  input \g2611_reg/NET0131  ;
  input \g2612_reg/NET0131  ;
  input \g2615_reg/NET0131  ;
  input \g2616_reg/NET0131  ;
  input \g2618_reg/NET0131  ;
  input \g261_reg/NET0131  ;
  input \g2622_reg/NET0131  ;
  input \g2633_reg/NET0131  ;
  input \g2637_pad  ;
  input \g2639_reg/NET0131  ;
  input \g2641_reg/NET0131  ;
  input \g2643_reg/NET0131  ;
  input \g2645_reg/NET0131  ;
  input \g2647_reg/NET0131  ;
  input \g2649_reg/NET0131  ;
  input \g264_reg/NET0131  ;
  input \g2650_reg/NET0131  ;
  input \g2651_reg/NET0131  ;
  input \g2652_reg/NET0131  ;
  input \g2653_reg/NET0131  ;
  input \g2654_reg/NET0131  ;
  input \g2655_reg/NET0131  ;
  input \g2656_reg/NET0131  ;
  input \g2657_reg/NET0131  ;
  input \g2658_reg/NET0131  ;
  input \g2659_reg/NET0131  ;
  input \g2660_reg/NET0131  ;
  input \g2661_reg/NET0131  ;
  input \g2664_reg/NET0131  ;
  input \g2667_reg/NET0131  ;
  input \g2670_reg/NET0131  ;
  input \g2673_reg/NET0131  ;
  input \g2676_reg/NET0131  ;
  input \g2679_reg/NET0131  ;
  input \g267_reg/NET0131  ;
  input \g2682_reg/NET0131  ;
  input \g2685_reg/NET0131  ;
  input \g2688_reg/NET0131  ;
  input \g2691_reg/NET0131  ;
  input \g2694_reg/NET0131  ;
  input \g270_reg/NET0131  ;
  input \g273_reg/NET0131  ;
  input \g2772_reg/NET0131  ;
  input \g2773_reg/NET0131  ;
  input \g2774_reg/NET0131  ;
  input \g2775_reg/NET0131  ;
  input \g2776_reg/NET0131  ;
  input \g2777_reg/NET0131  ;
  input \g2778_reg/NET0131  ;
  input \g2779_reg/NET0131  ;
  input \g2780_reg/NET0131  ;
  input \g2781_reg/NET0131  ;
  input \g2782_reg/NET0131  ;
  input \g2783_reg/NET0131  ;
  input \g2784_reg/NET0131  ;
  input \g2785_reg/NET0131  ;
  input \g2786_reg/NET0131  ;
  input \g2787_reg/NET0131  ;
  input \g2788_reg/NET0131  ;
  input \g2789_reg/NET0131  ;
  input \g2790_reg/NET0131  ;
  input \g2791_reg/NET0131  ;
  input \g2792_reg/NET0131  ;
  input \g2793_reg/NET0131  ;
  input \g2794_reg/NET0131  ;
  input \g2795_reg/NET0131  ;
  input \g2796_reg/NET0131  ;
  input \g2797_reg/NET0131  ;
  input \g2798_reg/NET0131  ;
  input \g2799_reg/NET0131  ;
  input \g279_reg/NET0131  ;
  input \g2800_reg/NET0131  ;
  input \g2801_reg/NET0131  ;
  input \g2802_reg/NET0131  ;
  input \g2803_reg/NET0131  ;
  input \g2804_reg/NET0131  ;
  input \g2805_reg/NET0131  ;
  input \g2806_reg/NET0131  ;
  input \g2807_reg/NET0131  ;
  input \g2808_reg/NET0131  ;
  input \g2809_reg/NET0131  ;
  input \g2810_reg/NET0131  ;
  input \g2811_reg/NET0131  ;
  input \g2812_reg/NET0131  ;
  input \g2813_reg/NET0131  ;
  input \g2814_reg/NET0131  ;
  input \g2817_reg/NET0131  ;
  input \g281_reg/NET0131  ;
  input \g283_reg/NET0131  ;
  input \g285_reg/NET0131  ;
  input \g2874_reg/NET0131  ;
  input \g2879_reg/NET0131  ;
  input \g287_reg/NET0131  ;
  input \g2883_reg/NET0131  ;
  input \g2888_reg/NET0131  ;
  input \g2892_reg/NET0131  ;
  input \g2896_reg/NET0131  ;
  input \g289_reg/NET0131  ;
  input \g2900_reg/NET0131  ;
  input \g2903_reg/NET0131  ;
  input \g2908_reg/NET0131  ;
  input \g2912_reg/NET0131  ;
  input \g2917_reg/NET0131  ;
  input \g291_reg/NET0131  ;
  input \g2920_reg/NET0131  ;
  input \g2924_reg/NET0131  ;
  input \g2929_reg/NET0131  ;
  input \g2933_reg/NET0131  ;
  input \g2934_reg/NET0131  ;
  input \g2935_reg/NET0131  ;
  input \g2938_reg/NET0131  ;
  input \g2941_reg/NET0131  ;
  input \g2944_reg/NET0131  ;
  input \g2947_reg/NET0131  ;
  input \g2950_reg/NET0131  ;
  input \g2953_reg/NET0131  ;
  input \g2956_reg/NET0131  ;
  input \g2959_reg/NET0131  ;
  input \g2962_reg/NET0131  ;
  input \g2963_reg/NET0131  ;
  input \g2966_reg/NET0131  ;
  input \g2969_reg/NET0131  ;
  input \g2972_reg/NET0131  ;
  input \g2975_reg/NET0131  ;
  input \g2978_reg/NET0131  ;
  input \g2981_reg/NET0131  ;
  input \g2984_reg/NET0131  ;
  input \g2985_reg/NET0131  ;
  input \g2986_reg/NET0131  ;
  input \g2987_reg/NET0131  ;
  input \g298_reg/NET0131  ;
  input \g2990_reg/NET0131  ;
  input \g2991_reg/NET0131  ;
  input \g2992_reg/NET0131  ;
  input \g2993_reg/NET0131  ;
  input \g2997_reg/NET0131  ;
  input \g2998_reg/NET0131  ;
  input \g299_reg/NET0131  ;
  input \g3002_reg/NET0131  ;
  input \g3006_reg/NET0131  ;
  input \g3010_reg/NET0131  ;
  input \g3013_reg/NET0131  ;
  input \g3018_reg/NET0131  ;
  input \g3024_reg/NET0131  ;
  input \g3028_reg/NET0131  ;
  input \g3032_reg/NET0131  ;
  input \g3036_reg/NET0131  ;
  input \g3043_reg/NET0131  ;
  input \g3044_reg/NET0131  ;
  input \g3045_reg/NET0131  ;
  input \g3046_reg/NET0131  ;
  input \g3047_reg/NET0131  ;
  input \g3048_reg/NET0131  ;
  input \g3049_reg/NET0131  ;
  input \g3050_reg/NET0131  ;
  input \g3051_reg/NET0131  ;
  input \g3052_reg/NET0131  ;
  input \g3053_reg/NET0131  ;
  input \g3054_reg/NET0131  ;
  input \g3055_reg/NET0131  ;
  input \g3056_reg/NET0131  ;
  input \g3057_reg/NET0131  ;
  input \g3058_reg/NET0131  ;
  input \g3059_reg/NET0131  ;
  input \g305_reg/NET0131  ;
  input \g3060_reg/NET0131  ;
  input \g3061_reg/NET0131  ;
  input \g3062_reg/NET0131  ;
  input \g3063_reg/NET0131  ;
  input \g3064_reg/NET0131  ;
  input \g3065_reg/NET0131  ;
  input \g3066_reg/NET0131  ;
  input \g3067_reg/NET0131  ;
  input \g3068_reg/NET0131  ;
  input \g3069_reg/NET0131  ;
  input \g3070_reg/NET0131  ;
  input \g3071_reg/NET0131  ;
  input \g3072_reg/NET0131  ;
  input \g3073_reg/NET0131  ;
  input \g3074_reg/NET0131  ;
  input \g3075_reg/NET0131  ;
  input \g3076_reg/NET0131  ;
  input \g3077_reg/NET0131  ;
  input \g3078_reg/NET0131  ;
  input \g3079_reg/NET0131  ;
  input \g3080_reg/NET0131  ;
  input \g3083_reg/NET0131  ;
  input \g3097_reg/NET0131  ;
  input \g3110_reg/NET0131  ;
  input \g3114_reg/NET0131  ;
  input \g3120_reg/NET0131  ;
  input \g312_reg/NET0131  ;
  input \g3139_reg/NET0131  ;
  input \g313_reg/NET0131  ;
  input \g314_reg/NET0131  ;
  input \g315_reg/NET0131  ;
  input \g316_reg/NET0131  ;
  input \g317_reg/NET0131  ;
  input \g318_reg/NET0131  ;
  input \g319_reg/NET0131  ;
  input \g320_reg/NET0131  ;
  input \g321_reg/NET0131  ;
  input \g3229_pad  ;
  input \g322_reg/NET0131  ;
  input \g3230_pad  ;
  input \g3231_pad  ;
  input \g3233_pad  ;
  input \g3234_pad  ;
  input \g323_reg/NET0131  ;
  input \g324_reg/NET0131  ;
  input \g343_reg/NET0131  ;
  input \g346_reg/NET0131  ;
  input \g349_reg/NET0131  ;
  input \g351_reg/NET0131  ;
  input \g353_reg/NET0131  ;
  input \g354_reg/NET0131  ;
  input \g358_reg/NET0131  ;
  input \g361_reg/NET0131  ;
  input \g364_reg/NET0131  ;
  input \g366_reg/NET0131  ;
  input \g368_reg/NET0131  ;
  input \g369_reg/NET0131  ;
  input \g373_reg/NET0131  ;
  input \g376_reg/NET0131  ;
  input \g379_reg/NET0131  ;
  input \g381_reg/NET0131  ;
  input \g383_reg/NET0131  ;
  input \g384_reg/NET0131  ;
  input \g388_reg/NET0131  ;
  input \g391_reg/NET0131  ;
  input \g394_reg/NET0131  ;
  input \g396_reg/NET0131  ;
  input \g398_reg/NET0131  ;
  input \g402_reg/NET0131  ;
  input \g403_reg/NET0131  ;
  input \g404_reg/NET0131  ;
  input \g408_reg/NET0131  ;
  input \g411_reg/NET0131  ;
  input \g414_reg/NET0131  ;
  input \g417_reg/NET0131  ;
  input \g420_reg/NET0131  ;
  input \g423_reg/NET0131  ;
  input \g426_reg/NET0131  ;
  input \g427_reg/NET0131  ;
  input \g428_reg/NET0131  ;
  input \g429_reg/NET0131  ;
  input \g432_reg/NET0131  ;
  input \g435_reg/NET0131  ;
  input \g438_reg/NET0131  ;
  input \g441_reg/NET0131  ;
  input \g444_reg/NET0131  ;
  input \g447_reg/NET0131  ;
  input \g448_reg/NET0131  ;
  input \g449_reg/NET0131  ;
  input \g451_reg/NET0131  ;
  input \g453_reg/NET0131  ;
  input \g464_reg/NET0131  ;
  input \g465_reg/NET0131  ;
  input \g468_reg/NET0131  ;
  input \g471_reg/NET0131  ;
  input \g477_reg/NET0131  ;
  input \g478_reg/NET0131  ;
  input \g479_reg/NET0131  ;
  input \g480_reg/NET0131  ;
  input \g484_reg/NET0131  ;
  input \g486_reg/NET0131  ;
  input \g487_reg/NET0131  ;
  input \g488_reg/NET0131  ;
  input \g489_reg/NET0131  ;
  input \g490_reg/NET0131  ;
  input \g493_reg/NET0131  ;
  input \g496_reg/NET0131  ;
  input \g499_reg/NET0131  ;
  input \g506_reg/NET0131  ;
  input \g507_reg/NET0131  ;
  input \g51_pad  ;
  input \g524_reg/NET0131  ;
  input \g525_reg/NET0131  ;
  input \g529_reg/NET0131  ;
  input \g530_reg/NET0131  ;
  input \g531_reg/NET0131  ;
  input \g532_reg/NET0131  ;
  input \g533_reg/NET0131  ;
  input \g534_reg/NET0131  ;
  input \g536_reg/NET0131  ;
  input \g537_reg/NET0131  ;
  input \g5388_pad  ;
  input \g538_reg/NET0131  ;
  input \g541_reg/NET0131  ;
  input \g542_reg/NET0131  ;
  input \g544_reg/NET0131  ;
  input \g548_reg/NET0131  ;
  input \g559_reg/NET0131  ;
  input \g563_pad  ;
  input \g5657_pad  ;
  input \g565_reg/NET0131  ;
  input \g567_reg/NET0131  ;
  input \g569_reg/NET0131  ;
  input \g571_reg/NET0131  ;
  input \g573_reg/NET0131  ;
  input \g575_reg/NET0131  ;
  input \g576_reg/NET0131  ;
  input \g577_reg/NET0131  ;
  input \g578_reg/NET0131  ;
  input \g579_reg/NET0131  ;
  input \g580_reg/NET0131  ;
  input \g581_reg/NET0131  ;
  input \g582_reg/NET0131  ;
  input \g583_reg/NET0131  ;
  input \g584_reg/NET0131  ;
  input \g585_reg/NET0131  ;
  input \g586_reg/NET0131  ;
  input \g587_reg/NET0131  ;
  input \g590_reg/NET0131  ;
  input \g593_reg/NET0131  ;
  input \g596_reg/NET0131  ;
  input \g599_reg/NET0131  ;
  input \g602_reg/NET0131  ;
  input \g605_reg/NET0131  ;
  input \g608_reg/NET0131  ;
  input \g611_reg/NET0131  ;
  input \g614_reg/NET0131  ;
  input \g617_reg/NET0131  ;
  input \g620_reg/NET0131  ;
  input \g698_reg/NET0131  ;
  input \g699_reg/NET0131  ;
  input \g700_reg/NET0131  ;
  input \g701_reg/NET0131  ;
  input \g702_reg/NET0131  ;
  input \g703_reg/NET0131  ;
  input \g704_reg/NET0131  ;
  input \g705_reg/NET0131  ;
  input \g706_reg/NET0131  ;
  input \g707_reg/NET0131  ;
  input \g708_reg/NET0131  ;
  input \g709_reg/NET0131  ;
  input \g710_reg/NET0131  ;
  input \g711_reg/NET0131  ;
  input \g712_reg/NET0131  ;
  input \g713_reg/NET0131  ;
  input \g714_reg/NET0131  ;
  input \g715_reg/NET0131  ;
  input \g716_reg/NET0131  ;
  input \g717_reg/NET0131  ;
  input \g718_reg/NET0131  ;
  input \g719_reg/NET0131  ;
  input \g720_reg/NET0131  ;
  input \g721_reg/NET0131  ;
  input \g722_reg/NET0131  ;
  input \g723_reg/NET0131  ;
  input \g724_reg/NET0131  ;
  input \g725_reg/NET0131  ;
  input \g726_reg/NET0131  ;
  input \g727_reg/NET0131  ;
  input \g728_reg/NET0131  ;
  input \g729_reg/NET0131  ;
  input \g730_reg/NET0131  ;
  input \g731_reg/NET0131  ;
  input \g732_reg/NET0131  ;
  input \g733_reg/NET0131  ;
  input \g734_reg/NET0131  ;
  input \g735_reg/NET0131  ;
  input \g736_reg/NET0131  ;
  input \g737_reg/NET0131  ;
  input \g738_reg/NET0131  ;
  input \g739_reg/NET0131  ;
  input \g785_reg/NET0131  ;
  input \g789_reg/NET0131  ;
  input \g793_reg/NET0131  ;
  input \g7961_pad  ;
  input \g797_reg/NET0131  ;
  input \g801_reg/NET0131  ;
  input \g805_reg/NET0131  ;
  input \g809_reg/NET0131  ;
  input \g813_reg/NET0131  ;
  input \g817_reg/NET0131  ;
  input \g818_reg/NET0131  ;
  input \g819_reg/NET0131  ;
  input \g820_reg/NET0131  ;
  input \g821_reg/NET0131  ;
  input \g822_reg/NET0131  ;
  input \g8259_pad  ;
  input \g8260_pad  ;
  input \g8261_pad  ;
  input \g8262_pad  ;
  input \g8263_pad  ;
  input \g8264_pad  ;
  input \g8265_pad  ;
  input \g8266_pad  ;
  input \g8268_pad  ;
  input \g8269_pad  ;
  input \g8270_pad  ;
  input \g8271_pad  ;
  input \g8272_pad  ;
  input \g8273_pad  ;
  input \g8274_pad  ;
  input \g8275_pad  ;
  input \g829_reg/NET0131  ;
  input \g830_reg/NET0131  ;
  input \g831_reg/NET0131  ;
  input \g832_reg/NET0131  ;
  input \g833_reg/NET0131  ;
  input \g834_reg/NET0131  ;
  input \g835_reg/NET0131  ;
  input \g836_reg/NET0131  ;
  input \g837_reg/NET0131  ;
  input \g838_reg/NET0131  ;
  input \g839_reg/NET0131  ;
  input \g840_reg/NET0131  ;
  input \g841_reg/NET0131  ;
  input \g842_reg/NET0131  ;
  input \g843_reg/NET0131  ;
  input \g844_reg/NET0131  ;
  input \g845_reg/NET0131  ;
  input \g846_reg/NET0131  ;
  input \g847_reg/NET0131  ;
  input \g848_reg/NET0131  ;
  input \g849_reg/NET0131  ;
  input \g850_reg/NET0131  ;
  input \g851_reg/NET0131  ;
  input \g852_reg/NET0131  ;
  input \g856_reg/NET0131  ;
  input \g857_reg/NET0131  ;
  input \g858_reg/NET0131  ;
  input \g859_reg/NET0131  ;
  input \g860_reg/NET0131  ;
  input \g861_reg/NET0131  ;
  input \g862_reg/NET0131  ;
  input \g863_reg/NET0131  ;
  input \g864_reg/NET0131  ;
  input \g865_reg/NET0131  ;
  input \g866_reg/NET0131  ;
  input \g867_reg/NET0131  ;
  input \g873_reg/NET0131  ;
  input \g876_reg/NET0131  ;
  input \g879_reg/NET0131  ;
  input \g882_reg/NET0131  ;
  input \g885_reg/NET0131  ;
  input \g888_reg/NET0131  ;
  input \g891_reg/NET0131  ;
  input \g894_reg/NET0131  ;
  input \g897_reg/NET0131  ;
  input \g900_reg/NET0131  ;
  input \g903_reg/NET0131  ;
  input \g906_reg/NET0131  ;
  input \g909_reg/NET0131  ;
  input \g912_reg/NET0131  ;
  input \g915_reg/NET0131  ;
  input \g918_reg/NET0131  ;
  input \g921_reg/NET0131  ;
  input \g924_reg/NET0131  ;
  input \g927_reg/NET0131  ;
  input \g930_reg/NET0131  ;
  input \g933_reg/NET0131  ;
  input \g936_reg/NET0131  ;
  input \g939_reg/NET0131  ;
  input \g942_reg/NET0131  ;
  input \g945_reg/NET0131  ;
  input \g948_reg/NET0131  ;
  input \g951_reg/NET0131  ;
  input \g954_reg/NET0131  ;
  input \g957_reg/NET0131  ;
  input \g960_reg/NET0131  ;
  input \g966_reg/NET0131  ;
  input \g968_reg/NET0131  ;
  input \g970_reg/NET0131  ;
  input \g972_reg/NET0131  ;
  input \g974_reg/NET0131  ;
  input \g976_reg/NET0131  ;
  input \g978_reg/NET0131  ;
  input \g97_reg/NET0131  ;
  input \g985_reg/NET0131  ;
  input \g986_reg/NET0131  ;
  input \g992_reg/NET0131  ;
  input \g999_reg/NET0131  ;
  output \_al_n0  ;
  output \_al_n1  ;
  output \g101_reg/P0001  ;
  output \g105_reg/P0001  ;
  output \g109_reg/P0001  ;
  output \g1138_reg/P0001  ;
  output \g113_reg/P0001  ;
  output \g1140_reg/P0001  ;
  output \g117_reg/P0001  ;
  output \g121_reg/P0001  ;
  output \g125_reg/P0001  ;
  output \g1471_reg/P0001  ;
  output \g1476_reg/P0001  ;
  output \g1481_reg/P0001  ;
  output \g1486_reg/P0001  ;
  output \g1491_reg/P0001  ;
  output \g1496_reg/P0001  ;
  output \g1501_reg/P0001  ;
  output \g1506_reg/P0001  ;
  output \g16496_pad  ;
  output \g1660_reg/P0001  ;
  output \g1662_reg/P0001  ;
  output \g1664_reg/P0001  ;
  output \g1666_reg/P0001  ;
  output \g1668_reg/P0001  ;
  output \g1670_reg/P0001  ;
  output \g1672_reg/P0001  ;
  output \g18/_0_  ;
  output \g1832_reg/P0001  ;
  output \g1834_reg/P0001  ;
  output \g2165_reg/P0001  ;
  output \g2170_reg/P0001  ;
  output \g2175_reg/P0001  ;
  output \g2180_reg/P0001  ;
  output \g2185_reg/P0001  ;
  output \g2190_reg/P0001  ;
  output \g2195_reg/P0001  ;
  output \g2200_reg/P0001  ;
  output \g2354_reg/P0001  ;
  output \g2356_reg/P0001  ;
  output \g2358_reg/P0001  ;
  output \g2360_reg/P0001  ;
  output \g2362_reg/P0001  ;
  output \g2364_reg/P0001  ;
  output \g2366_reg/P0001  ;
  output \g2526_reg/P0001  ;
  output \g2528_reg/P0001  ;
  output \g25489_pad  ;
  output \g279_reg/P0001  ;
  output \g281_reg/P0001  ;
  output \g283_reg/P0001  ;
  output \g285_reg/P0001  ;
  output \g2879_reg/NET0131_syn_2  ;
  output \g287_reg/P0001  ;
  output \g289_reg/P0001  ;
  output \g291_reg/P0001  ;
  output \g451_reg/P0001  ;
  output \g453_reg/P0001  ;
  output \g59421/_3_  ;
  output \g59425/_1_  ;
  output \g59435/_0_  ;
  output \g59436/_0_  ;
  output \g59441/_3_  ;
  output \g59442/_0_  ;
  output \g59445/_0_  ;
  output \g59453/_0_  ;
  output \g59462/_3_  ;
  output \g59466/_3_  ;
  output \g59467/_3_  ;
  output \g59468/_3_  ;
  output \g59469/_3_  ;
  output \g59470/_3_  ;
  output \g59471/_3_  ;
  output \g59472/_3_  ;
  output \g59473/_3_  ;
  output \g59489/_0_  ;
  output \g59498/_0_  ;
  output \g59499/_0_  ;
  output \g59500/_0_  ;
  output \g59502/_2_  ;
  output \g59503/_0_  ;
  output \g59505/_2_  ;
  output \g59507/_0_  ;
  output \g59508/_0_  ;
  output \g59533/_3_  ;
  output \g59534/_3_  ;
  output \g59535/_3_  ;
  output \g59536/_3_  ;
  output \g59537/_3_  ;
  output \g59538/_3_  ;
  output \g59539/_3_  ;
  output \g59540/_3_  ;
  output \g59548/_0_  ;
  output \g59550/_0_  ;
  output \g59551/_0_  ;
  output \g59552/_0_  ;
  output \g59554/_0_  ;
  output \g59555/_0_  ;
  output \g59556/_0_  ;
  output \g59557/_0_  ;
  output \g59558/_0_  ;
  output \g59559/_0_  ;
  output \g59560/_0_  ;
  output \g59561/_0_  ;
  output \g59639/_0_  ;
  output \g59694/_2_  ;
  output \g59695/_0_  ;
  output \g59697/_2_  ;
  output \g59698/_0_  ;
  output \g59699/_0_  ;
  output \g59700/_0_  ;
  output \g59705/_0_  ;
  output \g59706/_0_  ;
  output \g59707/_0_  ;
  output \g59708/_0_  ;
  output \g59709/_0_  ;
  output \g59710/_0_  ;
  output \g59711/_0_  ;
  output \g59712/_0_  ;
  output \g59713/_0_  ;
  output \g59714/_0_  ;
  output \g59715/_0_  ;
  output \g59716/_0_  ;
  output \g59717/_0_  ;
  output \g59718/_0_  ;
  output \g59719/_0_  ;
  output \g59720/_0_  ;
  output \g59721/_0_  ;
  output \g59722/_0_  ;
  output \g59723/_0_  ;
  output \g59724/_0_  ;
  output \g59725/_0_  ;
  output \g59726/_0_  ;
  output \g59727/_0_  ;
  output \g59728/_0_  ;
  output \g59729/_0_  ;
  output \g59730/_0_  ;
  output \g59731/_0_  ;
  output \g59732/_0_  ;
  output \g59733/_0_  ;
  output \g59734/_0_  ;
  output \g59735/_0_  ;
  output \g59736/_0_  ;
  output \g59737/_0_  ;
  output \g59738/_0_  ;
  output \g59739/_0_  ;
  output \g59740/_0_  ;
  output \g59741/_0_  ;
  output \g59742/_0_  ;
  output \g59743/_0_  ;
  output \g59744/_0_  ;
  output \g59745/_0_  ;
  output \g59747/_0_  ;
  output \g59748/_0_  ;
  output \g59749/_0_  ;
  output \g59750/_0_  ;
  output \g59751/_0_  ;
  output \g59752/_0_  ;
  output \g59753/_0_  ;
  output \g59754/_0_  ;
  output \g59755/_0_  ;
  output \g59756/_0_  ;
  output \g59757/_0_  ;
  output \g59758/_0_  ;
  output \g59759/_0_  ;
  output \g59760/_0_  ;
  output \g59761/_0_  ;
  output \g59762/_0_  ;
  output \g59763/_0_  ;
  output \g59764/_0_  ;
  output \g59765/_0_  ;
  output \g59766/_0_  ;
  output \g59915/_0_  ;
  output \g59952/_2_  ;
  output \g60046/_0_  ;
  output \g60048/_0_  ;
  output \g60049/_0_  ;
  output \g60051/_0_  ;
  output \g60063/_0_  ;
  output \g60103/_0_  ;
  output \g60104/_0_  ;
  output \g60105/_0_  ;
  output \g60107/_2_  ;
  output \g60108/_0_  ;
  output \g60109/_0_  ;
  output \g60110/_0_  ;
  output \g60112/_2_  ;
  output \g60119/_0_  ;
  output \g60120/_0_  ;
  output \g60121/_0_  ;
  output \g60122/_0_  ;
  output \g60123/_0_  ;
  output \g60124/_0_  ;
  output \g60126/_0_  ;
  output \g60127/_0_  ;
  output \g60128/_0_  ;
  output \g60129/_0_  ;
  output \g60130/_0_  ;
  output \g60135/_0_  ;
  output \g60136/_0_  ;
  output \g60137/_0_  ;
  output \g60138/_0_  ;
  output \g60139/_0_  ;
  output \g60143/_3_  ;
  output \g60144/_0_  ;
  output \g60145/_0_  ;
  output \g60339/_0_  ;
  output \g60404/_0_  ;
  output \g60427/_0_  ;
  output \g60428/_0_  ;
  output \g60429/_0_  ;
  output \g60434/_0_  ;
  output \g60435/_0_  ;
  output \g60437/_0_  ;
  output \g60438/_0_  ;
  output \g60439/_0_  ;
  output \g60440/_0_  ;
  output \g60441/_0_  ;
  output \g60448/_0_  ;
  output \g60451/_0_  ;
  output \g60452/_0_  ;
  output \g60453/_0_  ;
  output \g60459/_0_  ;
  output \g60460/_0_  ;
  output \g60523/_0_  ;
  output \g60534/_0_  ;
  output \g60535/_0_  ;
  output \g60536/_0_  ;
  output \g60585/_0_  ;
  output \g60586/_0_  ;
  output \g60587/_0_  ;
  output \g60588/_0_  ;
  output \g60591/_0_  ;
  output \g60592/_0_  ;
  output \g60599/_0_  ;
  output \g60601/_0_  ;
  output \g60602/_0_  ;
  output \g60603/_0_  ;
  output \g60604/_0_  ;
  output \g60605/_0_  ;
  output \g60606/_0_  ;
  output \g60607/_0_  ;
  output \g60608/_0_  ;
  output \g60609/_0_  ;
  output \g60613/_0_  ;
  output \g60614/_0_  ;
  output \g60615/_0_  ;
  output \g60694/_0_  ;
  output \g60708/_0_  ;
  output \g60709/_0_  ;
  output \g60710/_0_  ;
  output \g60785/_0_  ;
  output \g60787/_0_  ;
  output \g60788/_0_  ;
  output \g60799/_0_  ;
  output \g60801/_0_  ;
  output \g60802/_0_  ;
  output \g60803/_1__syn_2  ;
  output \g60805/_1__syn_2  ;
  output \g60806/_1__syn_2  ;
  output \g60808/_0_  ;
  output \g60810/_0_  ;
  output \g60811/_0_  ;
  output \g60825/_3_  ;
  output \g60896/_0_  ;
  output \g60980/_0_  ;
  output \g60981/_0_  ;
  output \g60985/_0_  ;
  output \g60986/_0_  ;
  output \g61012/_0_  ;
  output \g61013/_0_  ;
  output \g61015/_0_  ;
  output \g61017/_0_  ;
  output \g61122/_0_  ;
  output \g61123/_0_  ;
  output \g61124/_0_  ;
  output \g61125/_0_  ;
  output \g61222/_0_  ;
  output \g61223/_0_  ;
  output \g61224/_0_  ;
  output \g61225/_0_  ;
  output \g61228/_0_  ;
  output \g61229/_0_  ;
  output \g61230/_0_  ;
  output \g61231/_0_  ;
  output \g61281/_0_  ;
  output \g61293/_1_  ;
  output \g61307/_0__syn_2  ;
  output \g61309/_0__syn_2  ;
  output \g61310/_0__syn_2  ;
  output \g61311/_1_  ;
  output \g61312/_1_  ;
  output \g61313/_1_  ;
  output \g61324/_1_  ;
  output \g61325/_1_  ;
  output \g61326/_1_  ;
  output \g61328/_1_  ;
  output \g61329/_1_  ;
  output \g61330/_1_  ;
  output \g61332/_1_  ;
  output \g61333/_1_  ;
  output \g61334/_1_  ;
  output \g61335/_1_  ;
  output \g61336/_0_  ;
  output \g61338/_0_  ;
  output \g61339/_0_  ;
  output \g61340/_0_  ;
  output \g61377/_1_  ;
  output \g61378/_1_  ;
  output \g61379/_1_  ;
  output \g61388/_1_  ;
  output \g61391/_0_  ;
  output \g61394/_1_  ;
  output \g61395/_1_  ;
  output \g61396/_1_  ;
  output \g61398/_1_  ;
  output \g61399/_1_  ;
  output \g61421/_1_  ;
  output \g61422/_1_  ;
  output \g61423/_1_  ;
  output \g61524/_0_  ;
  output \g61525/_0_  ;
  output \g61526/_0_  ;
  output \g61527/_0_  ;
  output \g61528/_0_  ;
  output \g61529/_0_  ;
  output \g61530/_0_  ;
  output \g61531/_0_  ;
  output \g61532/_0_  ;
  output \g61533/_0_  ;
  output \g61534/_0_  ;
  output \g61535/_0_  ;
  output \g61536/_0_  ;
  output \g61537/_0_  ;
  output \g61538/_0_  ;
  output \g61539/_0_  ;
  output \g61540/_0_  ;
  output \g61541/_0_  ;
  output \g61542/_0_  ;
  output \g61543/_0_  ;
  output \g61544/_0_  ;
  output \g61545/_0_  ;
  output \g61546/_0_  ;
  output \g61547/_0_  ;
  output \g61548/_0_  ;
  output \g61549/_0_  ;
  output \g61550/_0_  ;
  output \g61551/_0_  ;
  output \g61552/_0_  ;
  output \g61553/_0_  ;
  output \g61554/_0_  ;
  output \g61555/_0_  ;
  output \g61556/_0_  ;
  output \g61557/_0_  ;
  output \g61558/_0_  ;
  output \g61559/_0_  ;
  output \g61560/_0_  ;
  output \g61561/_0_  ;
  output \g61562/_0_  ;
  output \g61563/_0_  ;
  output \g61564/_0_  ;
  output \g61565/_0_  ;
  output \g61566/_0_  ;
  output \g61620/_0_  ;
  output \g61621/_0_  ;
  output \g61622/_0_  ;
  output \g61623/_0_  ;
  output \g61753/_0_  ;
  output \g61764/_0_  ;
  output \g61786/_0_  ;
  output \g61795/_0_  ;
  output \g61801/_0_  ;
  output \g61803/_0_  ;
  output \g61808/_0_  ;
  output \g61848/_0_  ;
  output \g61850/_0_  ;
  output \g61851/_0_  ;
  output \g62097/_0_  ;
  output \g62102/_0_  ;
  output \g62115/_0_  ;
  output \g62119/_0_  ;
  output \g62130/_1_  ;
  output \g62131/_0_  ;
  output \g62132/_0_  ;
  output \g62139/_1_  ;
  output \g62140/_1_  ;
  output \g62141/_1_  ;
  output \g62144/_0_  ;
  output \g62145/_0_  ;
  output \g62146/_0_  ;
  output \g62147/_0_  ;
  output \g62150/_0_  ;
  output \g62151/_1_  ;
  output \g62152/_0_  ;
  output \g62153/_1_  ;
  output \g62156/_1_  ;
  output \g62157/_0_  ;
  output \g62159/_0_  ;
  output \g62161/_0_  ;
  output \g62187/_1_  ;
  output \g62190/_1_  ;
  output \g62191/_1_  ;
  output \g62192/_1_  ;
  output \g62194/_1_  ;
  output \g62195/_1_  ;
  output \g62196/_1_  ;
  output \g62203/_0_  ;
  output \g62204/_1_  ;
  output \g62207/_0__syn_2  ;
  output \g62208/_1_  ;
  output \g62209/_1_  ;
  output \g62210/_1_  ;
  output \g62211/_1_  ;
  output \g62212/_1_  ;
  output \g62217/_0_  ;
  output \g62286/_0_  ;
  output \g62287/_0_  ;
  output \g62288/_0_  ;
  output \g62289/_0_  ;
  output \g62290/_0_  ;
  output \g62291/_0_  ;
  output \g62292/_0_  ;
  output \g62435/_0_  ;
  output \g62436/_0_  ;
  output \g62439/_0_  ;
  output \g62456/_0_  ;
  output \g62486/_1_  ;
  output \g62492/_1_  ;
  output \g62494/_0_  ;
  output \g62495/_1_  ;
  output \g62497/_0_  ;
  output \g62537/_0_  ;
  output \g62544/_0_  ;
  output \g62546/_0_  ;
  output \g62547/_0_  ;
  output \g62549/_3_  ;
  output \g62552/_0_  ;
  output \g62554/_0_  ;
  output \g62555/_0_  ;
  output \g62556/_0_  ;
  output \g62558/_0_  ;
  output \g62559/_0_  ;
  output \g62561/_0_  ;
  output \g62562/_0_  ;
  output \g62566/_0_  ;
  output \g62567/_0_  ;
  output \g62568/_0_  ;
  output \g62569/_0_  ;
  output \g62570/_0_  ;
  output \g62571/_0_  ;
  output \g62572/_0_  ;
  output \g62573/_0_  ;
  output \g62574/_0_  ;
  output \g62575/_0_  ;
  output \g62576/_0_  ;
  output \g62577/_0_  ;
  output \g62578/_0_  ;
  output \g62579/_0_  ;
  output \g62580/_0_  ;
  output \g62581/_0_  ;
  output \g62582/_0_  ;
  output \g62583/_0_  ;
  output \g62584/_0_  ;
  output \g62585/_0_  ;
  output \g62586/_0_  ;
  output \g62587/_0_  ;
  output \g62588/_0_  ;
  output \g62589/_0_  ;
  output \g62590/_0_  ;
  output \g62591/_0_  ;
  output \g62592/_0_  ;
  output \g62593/_0_  ;
  output \g62594/_0_  ;
  output \g62595/_0_  ;
  output \g62596/_0_  ;
  output \g62597/_0_  ;
  output \g62602/_0_  ;
  output \g62607/_0_  ;
  output \g62608/_0_  ;
  output \g62609/_0_  ;
  output \g62619/_0_  ;
  output \g62620/_0_  ;
  output \g62621/_0_  ;
  output \g62622/_0_  ;
  output \g62623/_0_  ;
  output \g62624/_0_  ;
  output \g62626/_0_  ;
  output \g62627/_0_  ;
  output \g62628/_0_  ;
  output \g62629/_0_  ;
  output \g62630/_0_  ;
  output \g62631/_0_  ;
  output \g62632/_0_  ;
  output \g62633/_0_  ;
  output \g62634/_0_  ;
  output \g62635/_0_  ;
  output \g62636/_0_  ;
  output \g62637/_0_  ;
  output \g62638/_0_  ;
  output \g62639/_0_  ;
  output \g62640/_0_  ;
  output \g62641/_0_  ;
  output \g62642/_0_  ;
  output \g62643/_0_  ;
  output \g62644/_0_  ;
  output \g62645/_0_  ;
  output \g62646/_0_  ;
  output \g62647/_0_  ;
  output \g62648/_0_  ;
  output \g62649/_0_  ;
  output \g62650/_0_  ;
  output \g62651/_0_  ;
  output \g62652/_0_  ;
  output \g62653/_0_  ;
  output \g62654/_0_  ;
  output \g62655/_0_  ;
  output \g62656/_0_  ;
  output \g62657/_0_  ;
  output \g62658/_0_  ;
  output \g62659/_0_  ;
  output \g62660/_0_  ;
  output \g62661/_0_  ;
  output \g62674/_0_  ;
  output \g62682/_0_  ;
  output \g62683/_0_  ;
  output \g62689/_0_  ;
  output \g62690/_0_  ;
  output \g62691/_0_  ;
  output \g62694/_0_  ;
  output \g62695/_0_  ;
  output \g62696/_0_  ;
  output \g62698/_0_  ;
  output \g62699/_0_  ;
  output \g62700/_0_  ;
  output \g62723/_0_  ;
  output \g62724/_0_  ;
  output \g62725/_0_  ;
  output \g62726/_0_  ;
  output \g62727/_0_  ;
  output \g62728/_0_  ;
  output \g62735/_0_  ;
  output \g62736/_0_  ;
  output \g62737/_0_  ;
  output \g62738/_0_  ;
  output \g62739/_0_  ;
  output \g62740/_0_  ;
  output \g62754/_0_  ;
  output \g62762/_0_  ;
  output \g62763/_0_  ;
  output \g62764/_0_  ;
  output \g62780/_0_  ;
  output \g62781/_0_  ;
  output \g62785/_0_  ;
  output \g62786/_0_  ;
  output \g62787/_0_  ;
  output \g62791/_0_  ;
  output \g62792/_0_  ;
  output \g62794/_0_  ;
  output \g62804/_0_  ;
  output \g62806/_0_  ;
  output \g62807/_0_  ;
  output \g62811/_0_  ;
  output \g62968/_0_  ;
  output \g63005/_0_  ;
  output \g63041/_0_  ;
  output \g63116/_0_  ;
  output \g63157/_0_  ;
  output \g63164/_0_  ;
  output \g63170/_0_  ;
  output \g63189/_0_  ;
  output \g63202/_0_  ;
  output \g63206/_0_  ;
  output \g63207/_0_  ;
  output \g63265/_0_  ;
  output \g63266/_0_  ;
  output \g63269/_0_  ;
  output \g63271/_0_  ;
  output \g63272/_0_  ;
  output \g63273/_0_  ;
  output \g63274/_0_  ;
  output \g63275/_0_  ;
  output \g63276/_0_  ;
  output \g63277/_0_  ;
  output \g63278/_0_  ;
  output \g63280/_0_  ;
  output \g63281/_0_  ;
  output \g63282/_0_  ;
  output \g63283/_0_  ;
  output \g63284/_0_  ;
  output \g63285/_0_  ;
  output \g63286/_0_  ;
  output \g63287/_0_  ;
  output \g63288/_0_  ;
  output \g63289/_0_  ;
  output \g63290/_0_  ;
  output \g63292/_0_  ;
  output \g63293/_0_  ;
  output \g63294/_0_  ;
  output \g63295/_0_  ;
  output \g63296/_0_  ;
  output \g63297/_0_  ;
  output \g63298/_0_  ;
  output \g63299/_0_  ;
  output \g63302/_0_  ;
  output \g63303/_0_  ;
  output \g63304/_0_  ;
  output \g63305/_0_  ;
  output \g63306/_0_  ;
  output \g63307/_0_  ;
  output \g63308/_0_  ;
  output \g63309/_0_  ;
  output \g63310/_0_  ;
  output \g63311/_0_  ;
  output \g63312/_0_  ;
  output \g63313/_0_  ;
  output \g63314/_0_  ;
  output \g63315/_0_  ;
  output \g63316/_0_  ;
  output \g63317/_0_  ;
  output \g63318/_0_  ;
  output \g63319/_0_  ;
  output \g63320/_0_  ;
  output \g63321/_0_  ;
  output \g63322/_0_  ;
  output \g63323/_0_  ;
  output \g63324/_0_  ;
  output \g63325/_0_  ;
  output \g63326/_0_  ;
  output \g63327/_0_  ;
  output \g63328/_0_  ;
  output \g63329/_0_  ;
  output \g63330/_0_  ;
  output \g63331/_0_  ;
  output \g63339/_0_  ;
  output \g63505/_0_  ;
  output \g63525/_0_  ;
  output \g63543/_1_  ;
  output \g63602/_0_  ;
  output \g63653/_0_  ;
  output \g63663/_1_  ;
  output \g63677/_0_  ;
  output \g63694/_0_  ;
  output \g63729/_0_  ;
  output \g63766/_0_  ;
  output \g63771/_1_  ;
  output \g63773/_1_  ;
  output \g63784/_1_  ;
  output \g63964/_0_  ;
  output \g63965/_0_  ;
  output \g63966/_0_  ;
  output \g63967/_0_  ;
  output \g64257/_1_  ;
  output \g64266/_0_  ;
  output \g64275/_0_  ;
  output \g64400/_0_  ;
  output \g64416/_0_  ;
  output \g64470/_3_  ;
  output \g64473/_0_  ;
  output \g64474/_0_  ;
  output \g64475/_0_  ;
  output \g64479/_0_  ;
  output \g64480/_0_  ;
  output \g64481/_0_  ;
  output \g64483/_0_  ;
  output \g64484/_0_  ;
  output \g64485/_0_  ;
  output \g64486/_0_  ;
  output \g64493/_0_  ;
  output \g64494/_0_  ;
  output \g64495/_0_  ;
  output \g64496/_0_  ;
  output \g64505/_3_  ;
  output \g64507/_0_  ;
  output \g64508/_0_  ;
  output \g64510/_0_  ;
  output \g64511/_0_  ;
  output \g64544/_0_  ;
  output \g64545/_0_  ;
  output \g64546/_0_  ;
  output \g64639/_0_  ;
  output \g64641/_0_  ;
  output \g64642/_0_  ;
  output \g64645/_0_  ;
  output \g64650/_0_  ;
  output \g64737/_0_  ;
  output \g64738/_0_  ;
  output \g65066/_0_  ;
  output \g65070/_0_  ;
  output \g65090/_0_  ;
  output \g65102/_0_  ;
  output \g65102/_3_  ;
  output \g65126/_3_  ;
  output \g65147/_3_  ;
  output \g65163/_0_  ;
  output \g65176/_3_  ;
  output \g65178/_0_  ;
  output \g65182/_0_  ;
  output \g65190/_1_  ;
  output \g65191/_0_  ;
  output \g65196/_0_  ;
  output \g65268/_0_  ;
  output \g65275/_0_  ;
  output \g65290/_0_  ;
  output \g65290/_3_  ;
  output \g65291/_0_  ;
  output \g65292/_0_  ;
  output \g65298/_0_  ;
  output \g65298/_3_  ;
  output \g65314/_0_  ;
  output \g65314/_3_  ;
  output \g65319/_3_  ;
  output \g65335/_0_  ;
  output \g65342/_0_  ;
  output \g65348/_0_  ;
  output \g65422/_0_  ;
  output \g65465/_1_  ;
  output \g65469/_1_  ;
  output \g65478/_1_  ;
  output \g65507/_0_  ;
  output \g65548/_0_  ;
  output \g65699/_1_  ;
  output \g65713/_1_  ;
  output \g65835/_0_  ;
  output \g65860/_0_  ;
  output \g65863/_0_  ;
  output \g66094/_1_  ;
  output \g66102/_0_  ;
  output \g66107/_0_  ;
  output \g66130/_3_  ;
  output \g66131/_3_  ;
  output \g66228/_1_  ;
  output \g66348/_1_  ;
  output \g66543/_0_  ;
  output \g66549/_1_  ;
  output \g66640/_3_  ;
  output \g66641/_3_  ;
  output \g66950/_1_  ;
  output \g67111/_0_  ;
  output \g67219/_0_  ;
  output \g67263/_0_  ;
  output \g67909/_1_  ;
  output \g68049/_0_  ;
  output \g68220/_0_  ;
  output \g68413/_0_  ;
  output \g68511/_0_  ;
  output \g68536/_0_  ;
  output \g68543/_1_  ;
  output \g68554/_0_  ;
  output \g68559/_0_  ;
  output \g70915/_0_  ;
  output \g71108/_1_  ;
  output \g71115/_2_  ;
  output \g71244_dup/_0_  ;
  output \g71368/_0_  ;
  output \g71581/_0_  ;
  output \g71720/_0_  ;
  output \g785_reg/P0001  ;
  output \g789_reg/P0001  ;
  output \g797_reg/P0001  ;
  output \g809_reg/P0001  ;
  output \g813_reg/P0001  ;
  output \g966_reg/P0001  ;
  output \g968_reg/P0001  ;
  output \g970_reg/P0001  ;
  output \g972_reg/P0001  ;
  output \g974_reg/P0001  ;
  output \g976_reg/P0001  ;
  output \g978_reg/P0001  ;
  wire n1180 , n1181 , n1182 , n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 , n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 , n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 , n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 , n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 , n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 , n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 , n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 , n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 , n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 , n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 , n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 , n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 , n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 , n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 , n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 , n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 , n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 , n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 , n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 , n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 , n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 , n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 , n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 , n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 , n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 , n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 , n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 , n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 , n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 , n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 , n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 , n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 , n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 , n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 , n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 , n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 , n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 , n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 , n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 , n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 , n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 , n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 , n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 , n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 , n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 , n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 , n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 , n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 , n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 , n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 , n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 , n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 , n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 , n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 , n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 , n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 , n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 , n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 , n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 , n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 , n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 , n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 , n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 , n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 , n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 , n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 , n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 , n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 , n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 , n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 , n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 , n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 , n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 , n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 , n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 , n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 , n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 , n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 , n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 , n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 , n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 , n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 , n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 , n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 , n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 , n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 , n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 , n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 , n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 , n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 , n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 , n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 , n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 , n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 , n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 , n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 , n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 , n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 , n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 , n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 , n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 , n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 , n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 , n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 , n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 , n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 , n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 , n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 , n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 , n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 , n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 , n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 , n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 , n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 , n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 , n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 , n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 , n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 , n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 , n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 , n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 , n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 , n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 , n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 , n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 , n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 , n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 , n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 , n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 , n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 , n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 , n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 , n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 , n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 , n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 , n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 , n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 , n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 , n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 , n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 , n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 , n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 , n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 , n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 , n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 , n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 , n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 , n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 , n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 , n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 , n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 , n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 , n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 , n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 , n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 , n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 , n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 , n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 , n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 , n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 , n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 , n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 , n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 , n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 , n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 , n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 , n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 , n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 , n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 , n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 , n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 , n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 , n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 , n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 , n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 , n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 , n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 , n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 , n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 , n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 , n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 , n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 , n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 , n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 , n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 , n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 , n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 , n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 , n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 , n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 , n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 , n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 , n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 , n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 , n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 , n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 , n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 , n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 , n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 , n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 , n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 , n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 , n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 , n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 , n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 , n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 , n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 , n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 , n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 , n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 , n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 , n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 , n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 , n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 , n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 , n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 , n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 , n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 , n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 , n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 , n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 , n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 , n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 , n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 , n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 , n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 , n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 , n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 , n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 , n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 , n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 , n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 , n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 , n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 , n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 , n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 , n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 , n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 , n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 , n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 , n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 , n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 , n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 , n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 , n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 , n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 , n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 , n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 , n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 , n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 , n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 , n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 , n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 , n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 , n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 , n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 , n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 , n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 , n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 , n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 , n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 , n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 , n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 , n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 , n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 , n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 , n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 , n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 , n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 , n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 , n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 , n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 , n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 , n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 , n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 , n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 , n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 , n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 , n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 , n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 , n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 , n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 , n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 , n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 , n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 , n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 , n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 , n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 , n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 , n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 , n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 , n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 , n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 , n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 , n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 , n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 , n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 , n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 , n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 , n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 , n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 , n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 , n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 , n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 , n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 , n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 , n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 , n8363 , n8364 , n8365 ;
  assign n1180 = ~\g2986_reg/NET0131  & \g5388_pad  ;
  assign n1181 = \g2987_reg/NET0131  & ~n1180 ;
  assign n1182 = \g1092_reg/NET0131  & ~\g2394_reg/NET0131  ;
  assign n1183 = ~\g2393_reg/NET0131  & \g7961_pad  ;
  assign n1184 = \g1088_reg/NET0131  & ~\g2395_reg/NET0131  ;
  assign n1185 = ~n1183 & ~n1184 ;
  assign n1186 = ~n1182 & n1185 ;
  assign n1187 = \g1092_reg/NET0131  & \g2336_reg/NET0131  ;
  assign n1188 = \g2333_reg/NET0131  & \g7961_pad  ;
  assign n1189 = \g1088_reg/NET0131  & \g2339_reg/NET0131  ;
  assign n1190 = ~n1188 & ~n1189 ;
  assign n1191 = ~n1187 & n1190 ;
  assign n1192 = ~\g2200_reg/NET0131  & ~n1191 ;
  assign n1193 = \g2200_reg/NET0131  & ~n1187 ;
  assign n1194 = n1190 & n1193 ;
  assign n1195 = ~n1192 & ~n1194 ;
  assign n1196 = \g2306_reg/NET0131  & \g7961_pad  ;
  assign n1197 = \g1088_reg/NET0131  & \g2312_reg/NET0131  ;
  assign n1198 = \g1092_reg/NET0131  & \g2309_reg/NET0131  ;
  assign n1199 = ~n1197 & ~n1198 ;
  assign n1200 = ~n1196 & n1199 ;
  assign n1201 = ~\g2170_reg/NET0131  & ~n1200 ;
  assign n1202 = \g2170_reg/NET0131  & ~n1196 ;
  assign n1203 = n1199 & n1202 ;
  assign n1204 = ~n1201 & ~n1203 ;
  assign n1205 = n1195 & n1204 ;
  assign n1206 = \g2324_reg/NET0131  & \g7961_pad  ;
  assign n1207 = \g1088_reg/NET0131  & \g2330_reg/NET0131  ;
  assign n1208 = ~n1206 & ~n1207 ;
  assign n1209 = \g1092_reg/NET0131  & \g2327_reg/NET0131  ;
  assign n1210 = \g2190_reg/NET0131  & ~n1209 ;
  assign n1211 = n1208 & n1210 ;
  assign n1212 = n1208 & ~n1209 ;
  assign n1213 = ~\g2190_reg/NET0131  & ~n1212 ;
  assign n1214 = ~n1211 & ~n1213 ;
  assign n1215 = \g1088_reg/NET0131  & ~\g2247_reg/NET0131  ;
  assign n1216 = \g1092_reg/NET0131  & ~\g2249_reg/NET0131  ;
  assign n1217 = ~\g2248_reg/NET0131  & \g7961_pad  ;
  assign n1218 = ~n1216 & ~n1217 ;
  assign n1219 = ~n1215 & n1218 ;
  assign n1220 = \g2342_reg/NET0131  & \g7961_pad  ;
  assign n1221 = \g1088_reg/NET0131  & \g2348_reg/NET0131  ;
  assign n1222 = \g1092_reg/NET0131  & \g2345_reg/NET0131  ;
  assign n1223 = ~n1221 & ~n1222 ;
  assign n1224 = ~n1220 & n1223 ;
  assign n1225 = ~n1219 & ~n1224 ;
  assign n1226 = n1219 & n1224 ;
  assign n1227 = ~n1225 & ~n1226 ;
  assign n1228 = \g1092_reg/NET0131  & \g2318_reg/NET0131  ;
  assign n1229 = \g1088_reg/NET0131  & \g2321_reg/NET0131  ;
  assign n1230 = ~n1228 & ~n1229 ;
  assign n1231 = \g2315_reg/NET0131  & \g7961_pad  ;
  assign n1232 = \g2180_reg/NET0131  & ~n1231 ;
  assign n1233 = n1230 & n1232 ;
  assign n1234 = n1230 & ~n1231 ;
  assign n1235 = ~\g2180_reg/NET0131  & ~n1234 ;
  assign n1236 = ~n1233 & ~n1235 ;
  assign n1237 = ~n1227 & n1236 ;
  assign n1238 = ~n1214 & ~n1237 ;
  assign n1239 = ~n1205 & n1238 ;
  assign n1240 = n1204 & n1236 ;
  assign n1241 = n1195 & n1214 ;
  assign n1242 = ~n1240 & ~n1241 ;
  assign n1243 = n1227 & n1242 ;
  assign n1244 = n1195 & ~n1227 ;
  assign n1245 = n1214 & n1236 ;
  assign n1246 = ~n1204 & ~n1245 ;
  assign n1247 = ~n1244 & n1246 ;
  assign n1248 = ~n1243 & ~n1247 ;
  assign n1249 = ~n1239 & n1248 ;
  assign n1250 = \g1088_reg/NET0131  & \g2285_reg/NET0131  ;
  assign n1251 = \g2279_reg/NET0131  & \g7961_pad  ;
  assign n1252 = \g1092_reg/NET0131  & \g2282_reg/NET0131  ;
  assign n1253 = ~n1251 & ~n1252 ;
  assign n1254 = ~n1250 & n1253 ;
  assign n1255 = ~\g2185_reg/NET0131  & ~n1254 ;
  assign n1256 = \g2185_reg/NET0131  & ~n1250 ;
  assign n1257 = n1253 & n1256 ;
  assign n1258 = ~n1255 & ~n1257 ;
  assign n1259 = ~n1227 & n1258 ;
  assign n1260 = n1245 & n1259 ;
  assign n1261 = \g1092_reg/NET0131  & \g2291_reg/NET0131  ;
  assign n1262 = \g2288_reg/NET0131  & \g7961_pad  ;
  assign n1263 = \g1088_reg/NET0131  & \g2294_reg/NET0131  ;
  assign n1264 = ~n1262 & ~n1263 ;
  assign n1265 = ~n1261 & n1264 ;
  assign n1266 = ~\g2195_reg/NET0131  & ~n1265 ;
  assign n1267 = \g2195_reg/NET0131  & ~n1261 ;
  assign n1268 = n1264 & n1267 ;
  assign n1269 = ~n1266 & ~n1268 ;
  assign n1270 = \g1088_reg/NET0131  & ~\g2250_reg/NET0131  ;
  assign n1271 = \g1092_reg/NET0131  & ~\g2252_reg/NET0131  ;
  assign n1272 = ~\g2251_reg/NET0131  & \g7961_pad  ;
  assign n1273 = ~n1271 & ~n1272 ;
  assign n1274 = ~n1270 & n1273 ;
  assign n1275 = \g2297_reg/NET0131  & \g7961_pad  ;
  assign n1276 = \g1088_reg/NET0131  & \g2303_reg/NET0131  ;
  assign n1277 = \g1092_reg/NET0131  & \g2300_reg/NET0131  ;
  assign n1278 = ~n1276 & ~n1277 ;
  assign n1279 = ~n1275 & n1278 ;
  assign n1280 = ~n1274 & ~n1279 ;
  assign n1281 = n1274 & n1279 ;
  assign n1282 = ~n1280 & ~n1281 ;
  assign n1283 = n1269 & ~n1282 ;
  assign n1284 = \g2261_reg/NET0131  & \g7961_pad  ;
  assign n1285 = \g1088_reg/NET0131  & \g2267_reg/NET0131  ;
  assign n1286 = ~n1284 & ~n1285 ;
  assign n1287 = \g1092_reg/NET0131  & \g2264_reg/NET0131  ;
  assign n1288 = \g2165_reg/NET0131  & ~n1287 ;
  assign n1289 = n1286 & n1288 ;
  assign n1290 = n1286 & ~n1287 ;
  assign n1291 = ~\g2165_reg/NET0131  & ~n1290 ;
  assign n1292 = ~n1289 & ~n1291 ;
  assign n1293 = \g2270_reg/NET0131  & \g7961_pad  ;
  assign n1294 = \g1088_reg/NET0131  & \g2276_reg/NET0131  ;
  assign n1295 = \g1092_reg/NET0131  & \g2273_reg/NET0131  ;
  assign n1296 = ~n1294 & ~n1295 ;
  assign n1297 = ~n1293 & n1296 ;
  assign n1298 = ~\g2175_reg/NET0131  & ~n1297 ;
  assign n1299 = \g2175_reg/NET0131  & ~n1293 ;
  assign n1300 = n1296 & n1299 ;
  assign n1301 = ~n1298 & ~n1300 ;
  assign n1302 = n1292 & n1301 ;
  assign n1303 = n1205 & n1302 ;
  assign n1304 = n1283 & n1303 ;
  assign n1305 = n1260 & n1304 ;
  assign n1306 = n1249 & ~n1305 ;
  assign n1307 = n1186 & ~n1306 ;
  assign n1308 = \g1092_reg/NET0131  & ~\g2246_reg/NET0131  ;
  assign n1309 = \g1088_reg/NET0131  & ~\g2244_reg/NET0131  ;
  assign n1310 = ~\g2245_reg/NET0131  & \g7961_pad  ;
  assign n1311 = ~n1309 & ~n1310 ;
  assign n1312 = ~n1308 & n1311 ;
  assign n1313 = ~\g2230_reg/NET0131  & \g7961_pad  ;
  assign n1314 = \g1088_reg/NET0131  & ~\g2229_reg/NET0131  ;
  assign n1315 = ~n1313 & ~n1314 ;
  assign n1316 = \g1092_reg/NET0131  & ~\g2231_reg/NET0131  ;
  assign n1317 = \g2195_reg/NET0131  & ~n1316 ;
  assign n1318 = n1315 & n1317 ;
  assign n1319 = n1315 & ~n1316 ;
  assign n1320 = ~\g2195_reg/NET0131  & ~n1319 ;
  assign n1321 = ~n1318 & ~n1320 ;
  assign n1322 = \g1092_reg/NET0131  & ~\g2237_reg/NET0131  ;
  assign n1323 = ~\g2236_reg/NET0131  & \g7961_pad  ;
  assign n1324 = \g1088_reg/NET0131  & ~\g2235_reg/NET0131  ;
  assign n1325 = ~n1323 & ~n1324 ;
  assign n1326 = ~n1322 & n1325 ;
  assign n1327 = ~n1274 & ~n1326 ;
  assign n1328 = n1274 & n1326 ;
  assign n1329 = ~n1327 & ~n1328 ;
  assign n1330 = n1321 & ~n1329 ;
  assign n1331 = ~\g2224_reg/NET0131  & \g7961_pad  ;
  assign n1332 = \g1088_reg/NET0131  & ~\g2223_reg/NET0131  ;
  assign n1333 = ~n1331 & ~n1332 ;
  assign n1334 = \g1092_reg/NET0131  & ~\g2225_reg/NET0131  ;
  assign n1335 = \g2185_reg/NET0131  & ~n1334 ;
  assign n1336 = n1333 & n1335 ;
  assign n1337 = n1333 & ~n1334 ;
  assign n1338 = ~\g2185_reg/NET0131  & ~n1337 ;
  assign n1339 = ~n1336 & ~n1338 ;
  assign n1340 = \g1092_reg/NET0131  & ~\g2207_reg/NET0131  ;
  assign n1341 = \g1088_reg/NET0131  & ~\g2205_reg/NET0131  ;
  assign n1342 = ~n1340 & ~n1341 ;
  assign n1343 = ~\g2206_reg/NET0131  & \g7961_pad  ;
  assign n1344 = \g2165_reg/NET0131  & ~n1343 ;
  assign n1345 = n1342 & n1344 ;
  assign n1346 = n1342 & ~n1343 ;
  assign n1347 = ~\g2165_reg/NET0131  & ~n1346 ;
  assign n1348 = ~n1345 & ~n1347 ;
  assign n1349 = n1339 & n1348 ;
  assign n1350 = n1330 & n1349 ;
  assign n1351 = ~\g2233_reg/NET0131  & \g7961_pad  ;
  assign n1352 = \g1088_reg/NET0131  & ~\g2232_reg/NET0131  ;
  assign n1353 = ~n1351 & ~n1352 ;
  assign n1354 = \g1092_reg/NET0131  & ~\g2234_reg/NET0131  ;
  assign n1355 = \g2200_reg/NET0131  & ~n1354 ;
  assign n1356 = n1353 & n1355 ;
  assign n1357 = n1353 & ~n1354 ;
  assign n1358 = ~\g2200_reg/NET0131  & ~n1357 ;
  assign n1359 = ~n1356 & ~n1358 ;
  assign n1360 = \g1088_reg/NET0131  & ~\g2208_reg/NET0131  ;
  assign n1361 = \g1092_reg/NET0131  & ~\g2210_reg/NET0131  ;
  assign n1362 = ~n1360 & ~n1361 ;
  assign n1363 = ~\g2209_reg/NET0131  & \g7961_pad  ;
  assign n1364 = \g2170_reg/NET0131  & ~n1363 ;
  assign n1365 = n1362 & n1364 ;
  assign n1366 = n1362 & ~n1363 ;
  assign n1367 = ~\g2170_reg/NET0131  & ~n1366 ;
  assign n1368 = ~n1365 & ~n1367 ;
  assign n1369 = n1359 & n1368 ;
  assign n1370 = \g1563_reg/NET0131  & ~n1312 ;
  assign n1371 = \g1088_reg/NET0131  & ~\g2220_reg/NET0131  ;
  assign n1372 = \g1092_reg/NET0131  & ~\g2222_reg/NET0131  ;
  assign n1373 = ~n1371 & ~n1372 ;
  assign n1374 = ~\g2221_reg/NET0131  & \g7961_pad  ;
  assign n1375 = \g2180_reg/NET0131  & ~n1374 ;
  assign n1376 = n1373 & n1375 ;
  assign n1377 = n1373 & ~n1374 ;
  assign n1378 = ~\g2180_reg/NET0131  & ~n1377 ;
  assign n1379 = ~n1376 & ~n1378 ;
  assign n1380 = n1370 & n1379 ;
  assign n1381 = n1369 & n1380 ;
  assign n1382 = n1350 & n1381 ;
  assign n1383 = n1258 & n1269 ;
  assign n1384 = n1282 & ~n1302 ;
  assign n1385 = ~n1383 & n1384 ;
  assign n1386 = ~n1282 & n1301 ;
  assign n1387 = n1269 & n1292 ;
  assign n1388 = ~n1258 & ~n1387 ;
  assign n1389 = ~n1386 & n1388 ;
  assign n1390 = ~n1385 & ~n1389 ;
  assign n1391 = n1258 & n1301 ;
  assign n1392 = ~n1283 & ~n1391 ;
  assign n1393 = ~n1292 & n1392 ;
  assign n1394 = \g1092_reg/NET0131  & ~\g2219_reg/NET0131  ;
  assign n1395 = \g1088_reg/NET0131  & ~\g2217_reg/NET0131  ;
  assign n1396 = ~n1394 & ~n1395 ;
  assign n1397 = ~\g2218_reg/NET0131  & \g7961_pad  ;
  assign n1398 = \g2175_reg/NET0131  & ~n1397 ;
  assign n1399 = n1396 & n1398 ;
  assign n1400 = n1396 & ~n1397 ;
  assign n1401 = ~\g2175_reg/NET0131  & ~n1400 ;
  assign n1402 = ~n1399 & ~n1401 ;
  assign n1403 = \g1088_reg/NET0131  & ~\g2226_reg/NET0131  ;
  assign n1404 = ~\g2227_reg/NET0131  & \g7961_pad  ;
  assign n1405 = ~n1403 & ~n1404 ;
  assign n1406 = \g1092_reg/NET0131  & ~\g2228_reg/NET0131  ;
  assign n1407 = \g2190_reg/NET0131  & ~n1406 ;
  assign n1408 = n1405 & n1407 ;
  assign n1409 = n1405 & ~n1406 ;
  assign n1410 = ~\g2190_reg/NET0131  & ~n1409 ;
  assign n1411 = ~n1408 & ~n1410 ;
  assign n1412 = n1402 & n1411 ;
  assign n1413 = \g1092_reg/NET0131  & ~\g2240_reg/NET0131  ;
  assign n1414 = \g1088_reg/NET0131  & ~\g2238_reg/NET0131  ;
  assign n1415 = ~\g2239_reg/NET0131  & \g7961_pad  ;
  assign n1416 = ~n1414 & ~n1415 ;
  assign n1417 = ~n1413 & n1416 ;
  assign n1418 = ~n1219 & n1417 ;
  assign n1419 = n1219 & ~n1417 ;
  assign n1420 = ~n1418 & ~n1419 ;
  assign n1421 = \g1092_reg/NET0131  & ~\g2398_reg/NET0131  ;
  assign n1422 = ~\g2397_reg/NET0131  & \g7961_pad  ;
  assign n1423 = \g1088_reg/NET0131  & ~\g2396_reg/NET0131  ;
  assign n1424 = ~n1422 & ~n1423 ;
  assign n1425 = ~n1421 & n1424 ;
  assign n1426 = n1420 & ~n1425 ;
  assign n1427 = n1412 & n1426 ;
  assign n1428 = ~n1393 & n1427 ;
  assign n1429 = n1390 & n1428 ;
  assign n1430 = n1382 & n1429 ;
  assign n1431 = ~n1312 & ~n1430 ;
  assign n1432 = ~n1307 & n1431 ;
  assign n1433 = \g1088_reg/NET0131  & ~\g2389_reg/NET0131  ;
  assign n1434 = ~\g2387_reg/NET0131  & \g7961_pad  ;
  assign n1435 = \g1092_reg/NET0131  & ~\g2388_reg/NET0131  ;
  assign n1436 = ~n1434 & ~n1435 ;
  assign n1437 = ~n1433 & n1436 ;
  assign n1438 = \g1563_reg/NET0131  & ~n1437 ;
  assign n1439 = ~n1432 & n1438 ;
  assign n1440 = \g1092_reg/NET0131  & ~\g2391_reg/NET0131  ;
  assign n1441 = ~\g2390_reg/NET0131  & \g7961_pad  ;
  assign n1442 = \g1088_reg/NET0131  & ~\g2392_reg/NET0131  ;
  assign n1443 = ~n1441 & ~n1442 ;
  assign n1444 = ~n1440 & n1443 ;
  assign n1445 = n1186 & n1437 ;
  assign n1446 = n1444 & n1445 ;
  assign n1447 = \g1088_reg/NET0131  & ~\g2477_reg/NET0131  ;
  assign n1448 = ~\g2478_reg/NET0131  & \g7961_pad  ;
  assign n1449 = \g1092_reg/NET0131  & ~\g2479_reg/NET0131  ;
  assign n1450 = ~n1448 & ~n1449 ;
  assign n1451 = ~n1447 & n1450 ;
  assign n1452 = n1420 & ~n1451 ;
  assign n1453 = n1412 & n1452 ;
  assign n1454 = n1382 & n1453 ;
  assign n1455 = ~n1446 & ~n1454 ;
  assign n1456 = ~n1186 & ~n1425 ;
  assign n1457 = ~n1437 & n1456 ;
  assign n1458 = n1420 & n1457 ;
  assign n1459 = n1412 & n1458 ;
  assign n1460 = n1382 & n1459 ;
  assign n1461 = n1444 & ~n1460 ;
  assign n1462 = n1455 & n1461 ;
  assign n1463 = ~n1439 & n1462 ;
  assign n1464 = n1390 & ~n1393 ;
  assign n1465 = n1186 & ~n1305 ;
  assign n1466 = n1249 & n1465 ;
  assign n1467 = n1464 & ~n1466 ;
  assign n1468 = ~n1437 & ~n1444 ;
  assign n1469 = n1370 & n1468 ;
  assign n1470 = ~n1454 & n1469 ;
  assign n1471 = ~n1467 & n1470 ;
  assign n1472 = ~n1446 & n1471 ;
  assign n1473 = \g7961_pad  & ~n1472 ;
  assign n1474 = ~n1463 & n1473 ;
  assign n1475 = ~\g2390_reg/NET0131  & ~\g7961_pad  ;
  assign n1476 = ~n1474 & ~n1475 ;
  assign n1477 = ~\g2991_reg/NET0131  & ~\g2992_reg/NET0131  ;
  assign n1478 = ~\g3114_reg/NET0131  & \g3120_reg/NET0131  ;
  assign n1479 = n1477 & n1478 ;
  assign n1480 = ~\g2984_reg/NET0131  & ~\g2985_reg/NET0131  ;
  assign n1481 = ~\g3120_reg/NET0131  & ~n1480 ;
  assign n1482 = ~\g3114_reg/NET0131  & \g3139_reg/NET0131  ;
  assign n1483 = ~n1481 & n1482 ;
  assign n1484 = ~n1479 & ~n1483 ;
  assign n1485 = \g3097_reg/NET0131  & \g3120_reg/NET0131  ;
  assign n1486 = \g3139_reg/NET0131  & n1485 ;
  assign n1487 = \g3114_reg/NET0131  & ~n1486 ;
  assign n1488 = n1484 & ~n1487 ;
  assign n1489 = ~\g3230_pad  & \g3233_pad  ;
  assign n1490 = ~\g3110_reg/NET0131  & ~\g3120_reg/NET0131  ;
  assign n1491 = ~\g3114_reg/NET0131  & ~\g3139_reg/NET0131  ;
  assign n1492 = n1490 & n1491 ;
  assign n1493 = n1489 & ~n1492 ;
  assign n1494 = ~\g3139_reg/NET0131  & n1490 ;
  assign n1495 = ~\g3114_reg/NET0131  & n1477 ;
  assign n1496 = n1494 & ~n1495 ;
  assign n1497 = n1489 & ~n1496 ;
  assign n1498 = ~\g8260_pad  & ~\g8263_pad  ;
  assign n1499 = \g8260_pad  & \g8263_pad  ;
  assign n1500 = ~n1498 & ~n1499 ;
  assign n1501 = \g8266_pad  & n1500 ;
  assign n1502 = ~\g8266_pad  & ~n1500 ;
  assign n1503 = ~n1501 & ~n1502 ;
  assign n1504 = \g8259_pad  & ~\g8261_pad  ;
  assign n1505 = ~\g8259_pad  & \g8261_pad  ;
  assign n1506 = ~n1504 & ~n1505 ;
  assign n1507 = \g8265_pad  & n1506 ;
  assign n1508 = ~\g8265_pad  & ~n1506 ;
  assign n1509 = ~n1507 & ~n1508 ;
  assign n1510 = n1503 & n1509 ;
  assign n1511 = ~n1503 & ~n1509 ;
  assign n1512 = ~n1510 & ~n1511 ;
  assign n1513 = \g8262_pad  & ~\g8264_pad  ;
  assign n1514 = ~\g8262_pad  & \g8264_pad  ;
  assign n1515 = ~n1513 & ~n1514 ;
  assign n1516 = \g2990_reg/NET0131  & n1515 ;
  assign n1517 = n1512 & n1516 ;
  assign n1518 = \g2990_reg/NET0131  & ~n1515 ;
  assign n1519 = ~n1512 & n1518 ;
  assign n1520 = ~n1517 & ~n1519 ;
  assign n1521 = ~\g2990_reg/NET0131  & ~n1515 ;
  assign n1522 = n1512 & n1521 ;
  assign n1523 = ~\g2990_reg/NET0131  & n1515 ;
  assign n1524 = ~n1512 & n1523 ;
  assign n1525 = ~n1522 & ~n1524 ;
  assign n1526 = n1520 & n1525 ;
  assign n1527 = \g3120_reg/NET0131  & ~\g3231_pad  ;
  assign n1528 = ~n1515 & ~n1527 ;
  assign n1529 = ~n1512 & n1528 ;
  assign n1530 = n1515 & ~n1527 ;
  assign n1531 = n1512 & n1530 ;
  assign n1532 = ~n1529 & ~n1531 ;
  assign n1533 = ~n1515 & n1527 ;
  assign n1534 = n1512 & n1533 ;
  assign n1535 = n1515 & n1527 ;
  assign n1536 = ~n1512 & n1535 ;
  assign n1537 = ~n1534 & ~n1536 ;
  assign n1538 = n1532 & n1537 ;
  assign n1539 = \g2987_reg/NET0131  & \g2997_reg/NET0131  ;
  assign n1540 = ~\g2987_reg/NET0131  & \g3061_reg/NET0131  ;
  assign n1541 = ~n1539 & ~n1540 ;
  assign n1542 = ~\g8270_pad  & ~\g8271_pad  ;
  assign n1543 = \g8270_pad  & \g8271_pad  ;
  assign n1544 = ~n1542 & ~n1543 ;
  assign n1545 = \g8273_pad  & n1544 ;
  assign n1546 = ~\g8273_pad  & ~n1544 ;
  assign n1547 = ~n1545 & ~n1546 ;
  assign n1548 = \g8268_pad  & ~\g8269_pad  ;
  assign n1549 = ~\g8268_pad  & \g8269_pad  ;
  assign n1550 = ~n1548 & ~n1549 ;
  assign n1551 = \g8272_pad  & n1550 ;
  assign n1552 = ~\g8272_pad  & ~n1550 ;
  assign n1553 = ~n1551 & ~n1552 ;
  assign n1554 = n1547 & n1553 ;
  assign n1555 = ~n1547 & ~n1553 ;
  assign n1556 = ~n1554 & ~n1555 ;
  assign n1557 = \g8274_pad  & ~\g8275_pad  ;
  assign n1558 = ~\g8274_pad  & \g8275_pad  ;
  assign n1559 = ~n1557 & ~n1558 ;
  assign n1560 = \g3083_reg/NET0131  & n1559 ;
  assign n1561 = n1556 & n1560 ;
  assign n1562 = \g3083_reg/NET0131  & ~n1559 ;
  assign n1563 = ~n1556 & n1562 ;
  assign n1564 = ~n1561 & ~n1563 ;
  assign n1565 = ~\g3083_reg/NET0131  & ~n1559 ;
  assign n1566 = n1556 & n1565 ;
  assign n1567 = ~\g3083_reg/NET0131  & n1559 ;
  assign n1568 = ~n1556 & n1567 ;
  assign n1569 = ~n1566 & ~n1568 ;
  assign n1570 = n1564 & n1569 ;
  assign n1571 = n1527 & n1559 ;
  assign n1572 = n1556 & n1571 ;
  assign n1573 = n1527 & ~n1559 ;
  assign n1574 = ~n1556 & n1573 ;
  assign n1575 = ~n1572 & ~n1574 ;
  assign n1576 = ~n1527 & ~n1559 ;
  assign n1577 = n1556 & n1576 ;
  assign n1578 = ~n1527 & n1559 ;
  assign n1579 = ~n1556 & n1578 ;
  assign n1580 = ~n1577 & ~n1579 ;
  assign n1581 = n1575 & n1580 ;
  assign n1582 = ~\g2633_reg/NET0131  & ~\g2637_pad  ;
  assign n1583 = \g2574_reg/NET0131  & ~\g2618_reg/NET0131  ;
  assign n1584 = n1582 & n1583 ;
  assign n1585 = \g2688_reg/NET0131  & \g5657_pad  ;
  assign n1586 = \g1024_reg/NET0131  & \g2694_reg/NET0131  ;
  assign n1587 = \g1018_reg/NET0131  & \g2691_reg/NET0131  ;
  assign n1588 = ~n1586 & ~n1587 ;
  assign n1589 = ~n1585 & n1588 ;
  assign n1590 = ~\g2797_reg/NET0131  & \g5657_pad  ;
  assign n1591 = \g1018_reg/NET0131  & ~\g2798_reg/NET0131  ;
  assign n1592 = \g1024_reg/NET0131  & ~\g2796_reg/NET0131  ;
  assign n1593 = ~n1591 & ~n1592 ;
  assign n1594 = ~n1590 & n1593 ;
  assign n1595 = ~n1589 & n1594 ;
  assign n1596 = ~\g2779_reg/NET0131  & \g5657_pad  ;
  assign n1597 = \g1018_reg/NET0131  & ~\g2780_reg/NET0131  ;
  assign n1598 = \g1024_reg/NET0131  & ~\g2778_reg/NET0131  ;
  assign n1599 = ~n1597 & ~n1598 ;
  assign n1600 = ~n1596 & n1599 ;
  assign n1601 = ~\g2791_reg/NET0131  & \g5657_pad  ;
  assign n1602 = \g1024_reg/NET0131  & ~\g2790_reg/NET0131  ;
  assign n1603 = \g1018_reg/NET0131  & ~\g2792_reg/NET0131  ;
  assign n1604 = ~n1602 & ~n1603 ;
  assign n1605 = ~n1601 & n1604 ;
  assign n1606 = ~n1600 & n1605 ;
  assign n1607 = ~\g2788_reg/NET0131  & \g5657_pad  ;
  assign n1608 = \g1024_reg/NET0131  & ~\g2787_reg/NET0131  ;
  assign n1609 = \g1018_reg/NET0131  & ~\g2789_reg/NET0131  ;
  assign n1610 = ~n1608 & ~n1609 ;
  assign n1611 = ~n1607 & n1610 ;
  assign n1612 = ~\g2785_reg/NET0131  & \g5657_pad  ;
  assign n1613 = \g1024_reg/NET0131  & ~\g2784_reg/NET0131  ;
  assign n1614 = \g1018_reg/NET0131  & ~\g2786_reg/NET0131  ;
  assign n1615 = ~n1613 & ~n1614 ;
  assign n1616 = ~n1612 & n1615 ;
  assign n1617 = n1611 & n1616 ;
  assign n1618 = n1606 & n1617 ;
  assign n1619 = ~\g2794_reg/NET0131  & \g5657_pad  ;
  assign n1620 = \g1024_reg/NET0131  & ~\g2793_reg/NET0131  ;
  assign n1621 = \g1018_reg/NET0131  & ~\g2795_reg/NET0131  ;
  assign n1622 = ~n1620 & ~n1621 ;
  assign n1623 = ~n1619 & n1622 ;
  assign n1624 = ~n1594 & n1623 ;
  assign n1625 = ~\g2782_reg/NET0131  & \g5657_pad  ;
  assign n1626 = \g1018_reg/NET0131  & ~\g2783_reg/NET0131  ;
  assign n1627 = \g1024_reg/NET0131  & ~\g2781_reg/NET0131  ;
  assign n1628 = ~n1626 & ~n1627 ;
  assign n1629 = ~n1625 & n1628 ;
  assign n1630 = ~\g2773_reg/NET0131  & \g5657_pad  ;
  assign n1631 = \g1024_reg/NET0131  & ~\g2772_reg/NET0131  ;
  assign n1632 = \g1018_reg/NET0131  & ~\g2774_reg/NET0131  ;
  assign n1633 = ~n1631 & ~n1632 ;
  assign n1634 = ~n1630 & n1633 ;
  assign n1635 = ~n1629 & n1634 ;
  assign n1636 = n1624 & n1635 ;
  assign n1637 = n1618 & n1636 ;
  assign n1638 = \g1018_reg/NET0131  & ~\g2813_reg/NET0131  ;
  assign n1639 = ~\g2812_reg/NET0131  & \g5657_pad  ;
  assign n1640 = \g1024_reg/NET0131  & ~\g2811_reg/NET0131  ;
  assign n1641 = ~n1639 & ~n1640 ;
  assign n1642 = ~n1638 & n1641 ;
  assign n1643 = \g1024_reg/NET0131  & ~\g2805_reg/NET0131  ;
  assign n1644 = ~\g2806_reg/NET0131  & \g5657_pad  ;
  assign n1645 = \g1018_reg/NET0131  & ~\g2807_reg/NET0131  ;
  assign n1646 = ~n1644 & ~n1645 ;
  assign n1647 = ~n1643 & n1646 ;
  assign n1648 = ~n1642 & ~n1647 ;
  assign n1649 = ~\g2776_reg/NET0131  & \g5657_pad  ;
  assign n1650 = \g1024_reg/NET0131  & ~\g2775_reg/NET0131  ;
  assign n1651 = \g1018_reg/NET0131  & ~\g2777_reg/NET0131  ;
  assign n1652 = ~n1650 & ~n1651 ;
  assign n1653 = ~n1649 & n1652 ;
  assign n1654 = ~\g2800_reg/NET0131  & \g5657_pad  ;
  assign n1655 = \g1018_reg/NET0131  & ~\g2801_reg/NET0131  ;
  assign n1656 = \g1024_reg/NET0131  & ~\g2799_reg/NET0131  ;
  assign n1657 = ~n1655 & ~n1656 ;
  assign n1658 = ~n1654 & n1657 ;
  assign n1659 = ~n1653 & ~n1658 ;
  assign n1660 = n1648 & n1659 ;
  assign n1661 = ~n1589 & n1660 ;
  assign n1662 = n1637 & n1661 ;
  assign n1663 = ~n1595 & ~n1662 ;
  assign n1664 = n1637 & n1660 ;
  assign n1665 = n1589 & ~n1594 ;
  assign n1666 = ~n1664 & n1665 ;
  assign n1667 = n1663 & ~n1666 ;
  assign n1668 = n1584 & n1667 ;
  assign n1669 = \g2679_reg/NET0131  & \g5657_pad  ;
  assign n1670 = \g1024_reg/NET0131  & \g2685_reg/NET0131  ;
  assign n1671 = \g1018_reg/NET0131  & \g2682_reg/NET0131  ;
  assign n1672 = ~n1670 & ~n1671 ;
  assign n1673 = ~n1669 & n1672 ;
  assign n1674 = n1658 & ~n1673 ;
  assign n1675 = n1660 & ~n1673 ;
  assign n1676 = n1637 & n1675 ;
  assign n1677 = ~n1674 & ~n1676 ;
  assign n1678 = ~n1658 & n1673 ;
  assign n1679 = ~n1664 & n1678 ;
  assign n1680 = n1677 & ~n1679 ;
  assign n1681 = n1668 & n1680 ;
  assign n1682 = \g1243_reg/NET0131  & n1584 ;
  assign n1683 = ~n1667 & ~n1680 ;
  assign n1684 = n1682 & ~n1683 ;
  assign n1685 = ~n1681 & n1684 ;
  assign n1686 = n1589 & ~n1600 ;
  assign n1687 = ~n1664 & n1686 ;
  assign n1688 = ~n1589 & n1600 ;
  assign n1689 = ~n1662 & ~n1688 ;
  assign n1690 = ~n1687 & n1689 ;
  assign n1691 = n1584 & n1690 ;
  assign n1692 = ~n1629 & n1673 ;
  assign n1693 = ~n1664 & n1692 ;
  assign n1694 = n1629 & ~n1673 ;
  assign n1695 = ~n1676 & ~n1694 ;
  assign n1696 = ~n1693 & n1695 ;
  assign n1697 = n1691 & ~n1696 ;
  assign n1698 = n1584 & n1696 ;
  assign n1699 = ~n1690 & n1698 ;
  assign n1700 = ~n1697 & ~n1699 ;
  assign n1701 = ~n1589 & ~n1634 ;
  assign n1702 = n1589 & n1634 ;
  assign n1703 = ~n1701 & ~n1702 ;
  assign n1704 = n1584 & ~n1703 ;
  assign n1705 = n1700 & ~n1704 ;
  assign n1706 = ~n1696 & n1704 ;
  assign n1707 = n1690 & n1706 ;
  assign n1708 = n1653 & ~n1673 ;
  assign n1709 = ~n1676 & ~n1708 ;
  assign n1710 = ~n1653 & n1673 ;
  assign n1711 = ~n1664 & n1710 ;
  assign n1712 = n1709 & ~n1711 ;
  assign n1713 = n1584 & n1712 ;
  assign n1714 = ~n1690 & n1704 ;
  assign n1715 = n1698 & n1714 ;
  assign n1716 = n1713 & ~n1715 ;
  assign n1717 = ~n1707 & n1716 ;
  assign n1718 = ~n1705 & n1717 ;
  assign n1719 = ~n1704 & ~n1713 ;
  assign n1720 = n1700 & n1719 ;
  assign n1721 = n1704 & ~n1712 ;
  assign n1722 = ~n1700 & n1721 ;
  assign n1723 = ~n1720 & ~n1722 ;
  assign n1724 = ~n1718 & n1723 ;
  assign n1725 = ~n1623 & ~n1673 ;
  assign n1726 = n1623 & n1673 ;
  assign n1727 = ~n1725 & ~n1726 ;
  assign n1728 = ~n1589 & ~n1616 ;
  assign n1729 = n1589 & n1616 ;
  assign n1730 = ~n1728 & ~n1729 ;
  assign n1731 = ~n1727 & ~n1730 ;
  assign n1732 = n1727 & n1730 ;
  assign n1733 = ~n1731 & ~n1732 ;
  assign n1734 = n1611 & n1673 ;
  assign n1735 = ~n1611 & ~n1673 ;
  assign n1736 = ~n1734 & ~n1735 ;
  assign n1737 = n1584 & ~n1736 ;
  assign n1738 = n1584 & ~n1737 ;
  assign n1739 = n1733 & n1738 ;
  assign n1740 = ~n1733 & n1737 ;
  assign n1741 = ~n1739 & ~n1740 ;
  assign n1742 = n1589 & n1605 ;
  assign n1743 = ~n1589 & ~n1605 ;
  assign n1744 = ~n1742 & ~n1743 ;
  assign n1745 = \g1880_reg/NET0131  & \g1924_reg/NET0131  ;
  assign n1746 = \g5657_pad  & ~n1745 ;
  assign n1747 = ~\g2622_reg/NET0131  & ~\g5657_pad  ;
  assign n1748 = ~\g2574_reg/NET0131  & ~n1747 ;
  assign n1749 = ~n1746 & n1748 ;
  assign n1750 = \g1186_reg/NET0131  & ~\g1230_reg/NET0131  ;
  assign n1751 = \g5657_pad  & n1750 ;
  assign n1752 = \g499_reg/NET0131  & \g544_reg/NET0131  ;
  assign n1753 = ~\g1186_reg/NET0131  & \g5657_pad  ;
  assign n1754 = ~n1752 & n1753 ;
  assign n1755 = ~n1751 & ~n1754 ;
  assign n1756 = ~\g1928_reg/NET0131  & ~\g5657_pad  ;
  assign n1757 = ~\g1880_reg/NET0131  & ~n1756 ;
  assign n1758 = n1748 & n1757 ;
  assign n1759 = n1755 & n1758 ;
  assign n1760 = ~n1749 & ~n1759 ;
  assign n1761 = n1584 & n1760 ;
  assign n1762 = ~n1744 & n1761 ;
  assign n1763 = \g1196_reg/NET0131  & ~n1762 ;
  assign n1764 = n1741 & n1763 ;
  assign n1765 = \g1196_reg/NET0131  & n1762 ;
  assign n1766 = ~n1741 & n1765 ;
  assign n1767 = ~n1764 & ~n1766 ;
  assign n1768 = ~\g1196_reg/NET0131  & ~\g1243_reg/NET0131  ;
  assign n1769 = \g2599_reg/NET0131  & n1768 ;
  assign n1770 = ~\g2612_reg/NET0131  & \g3229_pad  ;
  assign n1771 = n1769 & ~n1770 ;
  assign n1772 = \g2574_reg/NET0131  & \g2618_reg/NET0131  ;
  assign n1773 = n1582 & ~n1772 ;
  assign n1774 = ~\g2615_reg/NET0131  & ~\g3229_pad  ;
  assign n1775 = n1773 & ~n1774 ;
  assign n1776 = n1771 & n1775 ;
  assign n1777 = n1760 & n1776 ;
  assign n1778 = n1767 & ~n1777 ;
  assign n1779 = n1724 & n1778 ;
  assign n1780 = ~n1741 & n1763 ;
  assign n1781 = n1741 & n1765 ;
  assign n1782 = ~n1780 & ~n1781 ;
  assign n1783 = ~n1777 & n1782 ;
  assign n1784 = ~n1724 & n1783 ;
  assign n1785 = ~n1779 & ~n1784 ;
  assign n1786 = ~n1685 & ~n1785 ;
  assign n1787 = \g2987_reg/NET0131  & \g3070_reg/NET0131  ;
  assign n1788 = ~\g2987_reg/NET0131  & \g3051_reg/NET0131  ;
  assign n1789 = ~n1787 & ~n1788 ;
  assign n1790 = \g2987_reg/NET0131  & \g3078_reg/NET0131  ;
  assign n1791 = ~\g2987_reg/NET0131  & \g3060_reg/NET0131  ;
  assign n1792 = ~n1790 & ~n1791 ;
  assign n1793 = \g2987_reg/NET0131  & \g3075_reg/NET0131  ;
  assign n1794 = ~\g2987_reg/NET0131  & \g3057_reg/NET0131  ;
  assign n1795 = ~n1793 & ~n1794 ;
  assign n1796 = \g2987_reg/NET0131  & \g3076_reg/NET0131  ;
  assign n1797 = ~\g2987_reg/NET0131  & \g3058_reg/NET0131  ;
  assign n1798 = ~n1796 & ~n1797 ;
  assign n1799 = \g2987_reg/NET0131  & \g3072_reg/NET0131  ;
  assign n1800 = ~\g2987_reg/NET0131  & \g3053_reg/NET0131  ;
  assign n1801 = ~n1799 & ~n1800 ;
  assign n1802 = \g2987_reg/NET0131  & \g3077_reg/NET0131  ;
  assign n1803 = ~\g2987_reg/NET0131  & \g3059_reg/NET0131  ;
  assign n1804 = ~n1802 & ~n1803 ;
  assign n1805 = \g2987_reg/NET0131  & \g3074_reg/NET0131  ;
  assign n1806 = ~\g2987_reg/NET0131  & \g3056_reg/NET0131  ;
  assign n1807 = ~n1805 & ~n1806 ;
  assign n1808 = \g2987_reg/NET0131  & \g3071_reg/NET0131  ;
  assign n1809 = ~\g2987_reg/NET0131  & \g3052_reg/NET0131  ;
  assign n1810 = ~n1808 & ~n1809 ;
  assign n1811 = \g2987_reg/NET0131  & \g3073_reg/NET0131  ;
  assign n1812 = ~\g2987_reg/NET0131  & \g3055_reg/NET0131  ;
  assign n1813 = ~n1811 & ~n1812 ;
  assign n1814 = ~\g1939_reg/NET0131  & ~\g1943_pad  ;
  assign n1815 = \g1880_reg/NET0131  & ~\g1924_reg/NET0131  ;
  assign n1816 = n1814 & n1815 ;
  assign n1817 = ~\g2100_reg/NET0131  & \g5657_pad  ;
  assign n1818 = \g1024_reg/NET0131  & ~\g2099_reg/NET0131  ;
  assign n1819 = \g1018_reg/NET0131  & ~\g2101_reg/NET0131  ;
  assign n1820 = ~n1818 & ~n1819 ;
  assign n1821 = ~n1817 & n1820 ;
  assign n1822 = \g1024_reg/NET0131  & ~\g2111_reg/NET0131  ;
  assign n1823 = ~\g2112_reg/NET0131  & \g5657_pad  ;
  assign n1824 = \g1018_reg/NET0131  & ~\g2113_reg/NET0131  ;
  assign n1825 = ~n1823 & ~n1824 ;
  assign n1826 = ~n1822 & n1825 ;
  assign n1827 = n1821 & ~n1826 ;
  assign n1828 = ~\g2097_reg/NET0131  & \g5657_pad  ;
  assign n1829 = \g1018_reg/NET0131  & ~\g2098_reg/NET0131  ;
  assign n1830 = \g1024_reg/NET0131  & ~\g2096_reg/NET0131  ;
  assign n1831 = ~n1829 & ~n1830 ;
  assign n1832 = ~n1828 & n1831 ;
  assign n1833 = \g1018_reg/NET0131  & ~\g2119_reg/NET0131  ;
  assign n1834 = \g1024_reg/NET0131  & ~\g2117_reg/NET0131  ;
  assign n1835 = ~\g2118_reg/NET0131  & \g5657_pad  ;
  assign n1836 = ~n1834 & ~n1835 ;
  assign n1837 = ~n1833 & n1836 ;
  assign n1838 = n1832 & ~n1837 ;
  assign n1839 = n1827 & n1838 ;
  assign n1840 = ~\g2103_reg/NET0131  & \g5657_pad  ;
  assign n1841 = \g1024_reg/NET0131  & ~\g2102_reg/NET0131  ;
  assign n1842 = \g1018_reg/NET0131  & ~\g2104_reg/NET0131  ;
  assign n1843 = ~n1841 & ~n1842 ;
  assign n1844 = ~n1840 & n1843 ;
  assign n1845 = ~\g2094_reg/NET0131  & \g5657_pad  ;
  assign n1846 = \g1018_reg/NET0131  & ~\g2095_reg/NET0131  ;
  assign n1847 = \g1024_reg/NET0131  & ~\g2093_reg/NET0131  ;
  assign n1848 = ~n1846 & ~n1847 ;
  assign n1849 = ~n1845 & n1848 ;
  assign n1850 = ~n1844 & n1849 ;
  assign n1851 = ~\g2079_reg/NET0131  & \g5657_pad  ;
  assign n1852 = \g1024_reg/NET0131  & ~\g2078_reg/NET0131  ;
  assign n1853 = \g1018_reg/NET0131  & ~\g2080_reg/NET0131  ;
  assign n1854 = ~n1852 & ~n1853 ;
  assign n1855 = ~n1851 & n1854 ;
  assign n1856 = ~\g2091_reg/NET0131  & \g5657_pad  ;
  assign n1857 = \g1018_reg/NET0131  & ~\g2092_reg/NET0131  ;
  assign n1858 = \g1024_reg/NET0131  & ~\g2090_reg/NET0131  ;
  assign n1859 = ~n1857 & ~n1858 ;
  assign n1860 = ~n1856 & n1859 ;
  assign n1861 = n1855 & n1860 ;
  assign n1862 = n1850 & n1861 ;
  assign n1863 = ~\g2088_reg/NET0131  & \g5657_pad  ;
  assign n1864 = \g1024_reg/NET0131  & ~\g2087_reg/NET0131  ;
  assign n1865 = \g1018_reg/NET0131  & ~\g2089_reg/NET0131  ;
  assign n1866 = ~n1864 & ~n1865 ;
  assign n1867 = ~n1863 & n1866 ;
  assign n1868 = ~\g2082_reg/NET0131  & \g5657_pad  ;
  assign n1869 = \g1018_reg/NET0131  & ~\g2083_reg/NET0131  ;
  assign n1870 = \g1024_reg/NET0131  & ~\g2081_reg/NET0131  ;
  assign n1871 = ~n1869 & ~n1870 ;
  assign n1872 = ~n1868 & n1871 ;
  assign n1873 = ~n1867 & ~n1872 ;
  assign n1874 = ~\g2085_reg/NET0131  & \g5657_pad  ;
  assign n1875 = \g1018_reg/NET0131  & ~\g2086_reg/NET0131  ;
  assign n1876 = \g1024_reg/NET0131  & ~\g2084_reg/NET0131  ;
  assign n1877 = ~n1875 & ~n1876 ;
  assign n1878 = ~n1874 & n1877 ;
  assign n1879 = ~\g2106_reg/NET0131  & \g5657_pad  ;
  assign n1880 = \g1018_reg/NET0131  & ~\g2107_reg/NET0131  ;
  assign n1881 = \g1024_reg/NET0131  & ~\g2105_reg/NET0131  ;
  assign n1882 = ~n1880 & ~n1881 ;
  assign n1883 = ~n1879 & n1882 ;
  assign n1884 = ~n1878 & ~n1883 ;
  assign n1885 = n1873 & n1884 ;
  assign n1886 = n1862 & n1885 ;
  assign n1887 = n1839 & n1886 ;
  assign n1888 = \g1018_reg/NET0131  & \g1988_reg/NET0131  ;
  assign n1889 = \g1985_reg/NET0131  & \g5657_pad  ;
  assign n1890 = \g1024_reg/NET0131  & \g1991_reg/NET0131  ;
  assign n1891 = ~n1889 & ~n1890 ;
  assign n1892 = ~n1888 & n1891 ;
  assign n1893 = ~n1867 & n1892 ;
  assign n1894 = ~n1887 & n1893 ;
  assign n1895 = n1867 & ~n1892 ;
  assign n1896 = n1839 & ~n1892 ;
  assign n1897 = n1886 & n1896 ;
  assign n1898 = ~n1895 & ~n1897 ;
  assign n1899 = ~n1894 & n1898 ;
  assign n1900 = n1816 & n1899 ;
  assign n1901 = \g1024_reg/NET0131  & \g2000_reg/NET0131  ;
  assign n1902 = \g1994_reg/NET0131  & \g5657_pad  ;
  assign n1903 = \g1018_reg/NET0131  & \g1997_reg/NET0131  ;
  assign n1904 = ~n1902 & ~n1903 ;
  assign n1905 = ~n1901 & n1904 ;
  assign n1906 = ~n1878 & n1905 ;
  assign n1907 = ~n1887 & n1906 ;
  assign n1908 = n1878 & ~n1905 ;
  assign n1909 = n1839 & ~n1905 ;
  assign n1910 = n1886 & n1909 ;
  assign n1911 = ~n1908 & ~n1910 ;
  assign n1912 = ~n1907 & n1911 ;
  assign n1913 = n1900 & ~n1912 ;
  assign n1914 = n1816 & n1912 ;
  assign n1915 = ~n1899 & n1914 ;
  assign n1916 = ~n1913 & ~n1915 ;
  assign n1917 = ~n1855 & ~n1905 ;
  assign n1918 = n1855 & n1905 ;
  assign n1919 = ~n1917 & ~n1918 ;
  assign n1920 = n1816 & ~n1919 ;
  assign n1921 = n1916 & ~n1920 ;
  assign n1922 = n1899 & ~n1912 ;
  assign n1923 = ~n1899 & n1912 ;
  assign n1924 = ~n1922 & ~n1923 ;
  assign n1925 = n1920 & ~n1924 ;
  assign n1926 = ~n1921 & ~n1925 ;
  assign n1927 = ~n1872 & n1892 ;
  assign n1928 = ~n1887 & n1927 ;
  assign n1929 = n1872 & ~n1892 ;
  assign n1930 = ~n1897 & ~n1929 ;
  assign n1931 = ~n1928 & n1930 ;
  assign n1932 = ~n1832 & ~n1905 ;
  assign n1933 = n1832 & n1905 ;
  assign n1934 = ~n1932 & ~n1933 ;
  assign n1935 = n1816 & n1934 ;
  assign n1936 = n1931 & n1935 ;
  assign n1937 = n1816 & ~n1934 ;
  assign n1938 = ~n1931 & n1937 ;
  assign n1939 = ~n1936 & ~n1938 ;
  assign n1940 = ~n1860 & ~n1905 ;
  assign n1941 = n1860 & n1905 ;
  assign n1942 = ~n1940 & ~n1941 ;
  assign n1943 = ~n1849 & ~n1892 ;
  assign n1944 = n1849 & n1892 ;
  assign n1945 = ~n1943 & ~n1944 ;
  assign n1946 = ~n1942 & ~n1945 ;
  assign n1947 = n1942 & n1945 ;
  assign n1948 = ~n1946 & ~n1947 ;
  assign n1949 = ~n1821 & ~n1892 ;
  assign n1950 = n1821 & n1892 ;
  assign n1951 = ~n1949 & ~n1950 ;
  assign n1952 = n1816 & ~n1951 ;
  assign n1953 = ~n1948 & n1952 ;
  assign n1954 = n1816 & n1951 ;
  assign n1955 = n1948 & n1954 ;
  assign n1956 = ~n1953 & ~n1955 ;
  assign n1957 = n1939 & ~n1956 ;
  assign n1958 = ~n1939 & n1956 ;
  assign n1959 = ~n1957 & ~n1958 ;
  assign n1960 = ~n1926 & n1959 ;
  assign n1961 = \g1196_reg/NET0131  & n1956 ;
  assign n1962 = n1939 & n1961 ;
  assign n1963 = \g1196_reg/NET0131  & ~n1956 ;
  assign n1964 = ~n1939 & n1963 ;
  assign n1965 = ~n1962 & ~n1964 ;
  assign n1966 = \g1196_reg/NET0131  & ~n1920 ;
  assign n1967 = n1916 & n1966 ;
  assign n1968 = \g1196_reg/NET0131  & n1816 ;
  assign n1969 = ~n1919 & n1968 ;
  assign n1970 = n1816 & n1969 ;
  assign n1971 = ~n1912 & n1970 ;
  assign n1972 = n1899 & n1971 ;
  assign n1973 = n1912 & n1970 ;
  assign n1974 = ~n1899 & n1973 ;
  assign n1975 = ~n1972 & ~n1974 ;
  assign n1976 = ~n1967 & n1975 ;
  assign n1977 = n1965 & n1976 ;
  assign n1978 = ~n1960 & ~n1977 ;
  assign n1979 = ~n1883 & n1892 ;
  assign n1980 = ~n1887 & n1979 ;
  assign n1981 = n1883 & ~n1892 ;
  assign n1982 = ~n1897 & ~n1981 ;
  assign n1983 = ~n1980 & n1982 ;
  assign n1984 = ~n1844 & n1905 ;
  assign n1985 = ~n1887 & n1984 ;
  assign n1986 = n1844 & ~n1905 ;
  assign n1987 = ~n1910 & ~n1986 ;
  assign n1988 = ~n1985 & n1987 ;
  assign n1989 = ~n1983 & n1988 ;
  assign n1990 = n1983 & ~n1988 ;
  assign n1991 = ~n1989 & ~n1990 ;
  assign n1992 = \g1243_reg/NET0131  & n1816 ;
  assign n1993 = ~n1991 & n1992 ;
  assign n1994 = n1755 & n1757 ;
  assign n1995 = \g1905_reg/NET0131  & n1768 ;
  assign n1996 = ~\g1918_reg/NET0131  & \g3229_pad  ;
  assign n1997 = n1995 & ~n1996 ;
  assign n1998 = ~n1745 & n1814 ;
  assign n1999 = ~\g1921_reg/NET0131  & ~\g3229_pad  ;
  assign n2000 = n1998 & ~n1999 ;
  assign n2001 = n1997 & n2000 ;
  assign n2002 = ~n1994 & n2001 ;
  assign n2003 = ~n1993 & ~n2002 ;
  assign n2004 = ~n1978 & n2003 ;
  assign n2005 = ~\g1196_reg/NET0131  & \g1243_reg/NET0131  ;
  assign n2006 = n1760 & n1773 ;
  assign n2007 = n2005 & ~n2006 ;
  assign n2008 = \g2574_reg/NET0131  & n1660 ;
  assign n2009 = n1637 & n2008 ;
  assign n2010 = ~\g2809_reg/NET0131  & \g5657_pad  ;
  assign n2011 = \g1018_reg/NET0131  & ~\g2810_reg/NET0131  ;
  assign n2012 = \g1024_reg/NET0131  & ~\g2808_reg/NET0131  ;
  assign n2013 = ~n2011 & ~n2012 ;
  assign n2014 = ~n2010 & n2013 ;
  assign n2015 = \g2574_reg/NET0131  & ~n2014 ;
  assign n2016 = n2005 & ~n2015 ;
  assign n2017 = ~n2009 & n2016 ;
  assign n2018 = ~n2007 & ~n2017 ;
  assign n2019 = n1584 & ~n1769 ;
  assign n2020 = ~n1727 & n2019 ;
  assign n2021 = ~\g1196_reg/NET0131  & ~\g2599_reg/NET0131  ;
  assign n2022 = ~\g1243_reg/NET0131  & ~n2021 ;
  assign n2023 = ~\g1243_reg/NET0131  & ~\g2599_reg/NET0131  ;
  assign n2024 = ~\g1196_reg/NET0131  & ~\g2603_reg/NET0131  ;
  assign n2025 = ~n2023 & n2024 ;
  assign n2026 = n1773 & n2025 ;
  assign n2027 = n1760 & n2026 ;
  assign n2028 = n2022 & ~n2027 ;
  assign n2029 = ~n2020 & n2028 ;
  assign n2030 = n2018 & ~n2029 ;
  assign n2031 = ~n1730 & n2019 ;
  assign n2032 = ~\g1196_reg/NET0131  & ~\g2606_reg/NET0131  ;
  assign n2033 = ~n2023 & n2032 ;
  assign n2034 = n1773 & n2033 ;
  assign n2035 = n1760 & n2034 ;
  assign n2036 = ~n2031 & ~n2035 ;
  assign n2037 = n2022 & n2036 ;
  assign n2038 = n2018 & ~n2037 ;
  assign n2039 = ~\g1196_reg/NET0131  & ~n2023 ;
  assign n2040 = n1584 & ~n2039 ;
  assign n2041 = n1696 & n2040 ;
  assign n2042 = ~\g1196_reg/NET0131  & ~\g2607_reg/NET0131  ;
  assign n2043 = ~n2023 & n2042 ;
  assign n2044 = n1773 & n2043 ;
  assign n2045 = n1760 & n2044 ;
  assign n2046 = n2022 & ~n2045 ;
  assign n2047 = ~n2041 & n2046 ;
  assign n2048 = ~n2007 & ~n2047 ;
  assign n2049 = n2006 & ~n2015 ;
  assign n2050 = ~n2009 & n2049 ;
  assign n2051 = n2005 & ~n2050 ;
  assign n2052 = ~n1736 & n2019 ;
  assign n2053 = ~\g1196_reg/NET0131  & ~\g2605_reg/NET0131  ;
  assign n2054 = ~n2023 & n2053 ;
  assign n2055 = n1773 & n2054 ;
  assign n2056 = n1760 & n2055 ;
  assign n2057 = ~n2052 & ~n2056 ;
  assign n2058 = n2022 & n2057 ;
  assign n2059 = ~n2051 & ~n2058 ;
  assign n2060 = n1690 & n2040 ;
  assign n2061 = ~\g1196_reg/NET0131  & ~\g2608_reg/NET0131  ;
  assign n2062 = ~n2023 & n2061 ;
  assign n2063 = n1773 & n2062 ;
  assign n2064 = n1760 & n2063 ;
  assign n2065 = n2022 & ~n2064 ;
  assign n2066 = ~n2060 & n2065 ;
  assign n2067 = ~n2007 & ~n2066 ;
  assign n2068 = ~n1744 & n2019 ;
  assign n2069 = ~\g1196_reg/NET0131  & ~\g2604_reg/NET0131  ;
  assign n2070 = ~n2023 & n2069 ;
  assign n2071 = n1773 & n2070 ;
  assign n2072 = n1760 & n2071 ;
  assign n2073 = ~n2068 & ~n2072 ;
  assign n2074 = n2022 & n2073 ;
  assign n2075 = ~n2051 & ~n2074 ;
  assign n2076 = n1584 & n1680 ;
  assign n2077 = n2005 & ~n2076 ;
  assign n2078 = n1712 & n2019 ;
  assign n2079 = ~\g1196_reg/NET0131  & ~\g2610_reg/NET0131  ;
  assign n2080 = ~n2023 & n2079 ;
  assign n2081 = n1773 & n2080 ;
  assign n2082 = n1760 & n2081 ;
  assign n2083 = n2022 & ~n2082 ;
  assign n2084 = ~n2078 & n2083 ;
  assign n2085 = ~n2077 & ~n2084 ;
  assign n2086 = ~n1703 & n2019 ;
  assign n2087 = ~\g1196_reg/NET0131  & ~\g2611_reg/NET0131  ;
  assign n2088 = ~n2023 & n2087 ;
  assign n2089 = n1773 & n2088 ;
  assign n2090 = n1760 & n2089 ;
  assign n2091 = ~n2086 & ~n2090 ;
  assign n2092 = n2022 & n2091 ;
  assign n2093 = ~n2005 & ~n2092 ;
  assign n2094 = n1584 & ~n2092 ;
  assign n2095 = n1667 & n2094 ;
  assign n2096 = ~n2093 & ~n2095 ;
  assign n2097 = \g2987_reg/NET0131  & \g3067_reg/NET0131  ;
  assign n2098 = ~\g2987_reg/NET0131  & \g3048_reg/NET0131  ;
  assign n2099 = ~n2097 & ~n2098 ;
  assign n2100 = \g2987_reg/NET0131  & \g3068_reg/NET0131  ;
  assign n2101 = ~\g2987_reg/NET0131  & \g3049_reg/NET0131  ;
  assign n2102 = ~n2100 & ~n2101 ;
  assign n2103 = \g2987_reg/NET0131  & \g3069_reg/NET0131  ;
  assign n2104 = ~\g2987_reg/NET0131  & \g3050_reg/NET0131  ;
  assign n2105 = ~n2103 & ~n2104 ;
  assign n2106 = \g2987_reg/NET0131  & \g3065_reg/NET0131  ;
  assign n2107 = ~\g2987_reg/NET0131  & \g3046_reg/NET0131  ;
  assign n2108 = ~n2106 & ~n2107 ;
  assign n2109 = \g2987_reg/NET0131  & \g3064_reg/NET0131  ;
  assign n2110 = ~\g2987_reg/NET0131  & \g3045_reg/NET0131  ;
  assign n2111 = ~n2109 & ~n2110 ;
  assign n2112 = \g2987_reg/NET0131  & \g3063_reg/NET0131  ;
  assign n2113 = ~\g2987_reg/NET0131  & \g3044_reg/NET0131  ;
  assign n2114 = ~n2112 & ~n2113 ;
  assign n2115 = \g2987_reg/NET0131  & \g3062_reg/NET0131  ;
  assign n2116 = ~\g2987_reg/NET0131  & \g3043_reg/NET0131  ;
  assign n2117 = ~n2115 & ~n2116 ;
  assign n2118 = \g2987_reg/NET0131  & \g3066_reg/NET0131  ;
  assign n2119 = ~\g2987_reg/NET0131  & \g3047_reg/NET0131  ;
  assign n2120 = ~n2118 & ~n2119 ;
  assign n2121 = ~\g2373_reg/NET0131  & ~\g2374_reg/NET0131  ;
  assign n2122 = ~\g1092_reg/NET0131  & ~\g1686_reg/NET0131  ;
  assign n2123 = \g1680_reg/NET0131  & ~n2122 ;
  assign n2124 = ~\g1679_reg/NET0131  & ~\g1680_reg/NET0131  ;
  assign n2125 = \g1092_reg/NET0131  & ~n2124 ;
  assign n2126 = ~n2123 & n2125 ;
  assign n2127 = ~\g298_reg/NET0131  & ~\g299_reg/NET0131  ;
  assign n2128 = \g1092_reg/NET0131  & ~n2127 ;
  assign n2129 = ~\g1092_reg/NET0131  & ~\g992_reg/NET0131  ;
  assign n2130 = \g986_reg/NET0131  & ~n2129 ;
  assign n2131 = ~n2128 & n2130 ;
  assign n2132 = ~\g985_reg/NET0131  & ~\g986_reg/NET0131  ;
  assign n2133 = \g1092_reg/NET0131  & ~n2132 ;
  assign n2134 = n2125 & n2133 ;
  assign n2135 = ~n2131 & n2134 ;
  assign n2136 = ~n2126 & ~n2135 ;
  assign n2137 = ~\g1092_reg/NET0131  & ~\g2380_reg/NET0131  ;
  assign n2138 = \g2374_reg/NET0131  & ~n2137 ;
  assign n2139 = n2136 & n2138 ;
  assign n2140 = ~n2121 & ~n2139 ;
  assign n2141 = \g315_reg/NET0131  & ~\g7961_pad  ;
  assign n2142 = ~\g315_reg/NET0131  & \g7961_pad  ;
  assign n2143 = \g1088_reg/NET0131  & ~\g317_reg/NET0131  ;
  assign n2144 = \g1092_reg/NET0131  & ~\g316_reg/NET0131  ;
  assign n2145 = ~n2143 & ~n2144 ;
  assign n2146 = ~n2142 & n2145 ;
  assign n2147 = \g1088_reg/NET0131  & ~\g314_reg/NET0131  ;
  assign n2148 = ~\g312_reg/NET0131  & \g7961_pad  ;
  assign n2149 = \g1092_reg/NET0131  & ~\g313_reg/NET0131  ;
  assign n2150 = ~n2148 & ~n2149 ;
  assign n2151 = ~n2147 & n2150 ;
  assign n2152 = n2146 & ~n2151 ;
  assign n2153 = \g1092_reg/NET0131  & ~\g146_reg/NET0131  ;
  assign n2154 = ~\g145_reg/NET0131  & \g7961_pad  ;
  assign n2155 = ~n2153 & ~n2154 ;
  assign n2156 = \g1088_reg/NET0131  & ~\g144_reg/NET0131  ;
  assign n2157 = \g109_reg/NET0131  & ~n2156 ;
  assign n2158 = n2155 & n2157 ;
  assign n2159 = n2155 & ~n2156 ;
  assign n2160 = ~\g109_reg/NET0131  & ~n2159 ;
  assign n2161 = ~n2158 & ~n2160 ;
  assign n2162 = \g1092_reg/NET0131  & ~\g158_reg/NET0131  ;
  assign n2163 = ~\g157_reg/NET0131  & \g7961_pad  ;
  assign n2164 = ~n2162 & ~n2163 ;
  assign n2165 = \g1088_reg/NET0131  & ~\g156_reg/NET0131  ;
  assign n2166 = \g125_reg/NET0131  & ~n2165 ;
  assign n2167 = n2164 & n2166 ;
  assign n2168 = n2164 & ~n2165 ;
  assign n2169 = ~\g125_reg/NET0131  & ~n2168 ;
  assign n2170 = ~n2167 & ~n2169 ;
  assign n2171 = \g1092_reg/NET0131  & ~\g134_reg/NET0131  ;
  assign n2172 = \g1088_reg/NET0131  & ~\g132_reg/NET0131  ;
  assign n2173 = ~n2171 & ~n2172 ;
  assign n2174 = ~\g133_reg/NET0131  & \g7961_pad  ;
  assign n2175 = \g101_reg/NET0131  & ~n2174 ;
  assign n2176 = n2173 & n2175 ;
  assign n2177 = n2173 & ~n2174 ;
  assign n2178 = ~\g101_reg/NET0131  & ~n2177 ;
  assign n2179 = ~n2176 & ~n2178 ;
  assign n2180 = n2170 & n2179 ;
  assign n2181 = n2161 & n2180 ;
  assign n2182 = \g1088_reg/NET0131  & ~\g150_reg/NET0131  ;
  assign n2183 = ~\g151_reg/NET0131  & \g7961_pad  ;
  assign n2184 = ~n2182 & ~n2183 ;
  assign n2185 = \g1092_reg/NET0131  & ~\g152_reg/NET0131  ;
  assign n2186 = \g117_reg/NET0131  & ~n2185 ;
  assign n2187 = n2184 & n2186 ;
  assign n2188 = n2184 & ~n2185 ;
  assign n2189 = ~\g117_reg/NET0131  & ~n2188 ;
  assign n2190 = ~n2187 & ~n2189 ;
  assign n2191 = \g1092_reg/NET0131  & ~\g143_reg/NET0131  ;
  assign n2192 = \g1088_reg/NET0131  & ~\g141_reg/NET0131  ;
  assign n2193 = ~n2191 & ~n2192 ;
  assign n2194 = ~\g142_reg/NET0131  & \g7961_pad  ;
  assign n2195 = \g105_reg/NET0131  & ~n2194 ;
  assign n2196 = n2193 & n2195 ;
  assign n2197 = n2193 & ~n2194 ;
  assign n2198 = ~\g105_reg/NET0131  & ~n2197 ;
  assign n2199 = ~n2196 & ~n2198 ;
  assign n2200 = n2190 & n2199 ;
  assign n2201 = \g1088_reg/NET0131  & ~\g147_reg/NET0131  ;
  assign n2202 = \g1092_reg/NET0131  & ~\g149_reg/NET0131  ;
  assign n2203 = ~n2201 & ~n2202 ;
  assign n2204 = ~\g148_reg/NET0131  & \g7961_pad  ;
  assign n2205 = \g113_reg/NET0131  & ~n2204 ;
  assign n2206 = n2203 & n2205 ;
  assign n2207 = n2203 & ~n2204 ;
  assign n2208 = ~\g113_reg/NET0131  & ~n2207 ;
  assign n2209 = ~n2206 & ~n2208 ;
  assign n2210 = \g1088_reg/NET0131  & ~\g153_reg/NET0131  ;
  assign n2211 = ~\g154_reg/NET0131  & \g7961_pad  ;
  assign n2212 = ~n2210 & ~n2211 ;
  assign n2213 = \g1092_reg/NET0131  & ~\g155_reg/NET0131  ;
  assign n2214 = \g121_reg/NET0131  & ~n2213 ;
  assign n2215 = n2212 & n2214 ;
  assign n2216 = n2212 & ~n2213 ;
  assign n2217 = ~\g121_reg/NET0131  & ~n2216 ;
  assign n2218 = ~n2215 & ~n2217 ;
  assign n2219 = n2209 & n2218 ;
  assign n2220 = n2200 & n2219 ;
  assign n2221 = \g1092_reg/NET0131  & ~\g131_reg/NET0131  ;
  assign n2222 = \g1088_reg/NET0131  & ~\g129_reg/NET0131  ;
  assign n2223 = ~n2221 & ~n2222 ;
  assign n2224 = ~\g130_reg/NET0131  & \g7961_pad  ;
  assign n2225 = \g97_reg/NET0131  & ~n2224 ;
  assign n2226 = n2223 & n2225 ;
  assign n2227 = n2223 & ~n2224 ;
  assign n2228 = ~\g97_reg/NET0131  & ~n2227 ;
  assign n2229 = ~n2226 & ~n2228 ;
  assign n2230 = n2220 & n2229 ;
  assign n2231 = \g1088_reg/NET0131  & ~\g171_reg/NET0131  ;
  assign n2232 = \g1092_reg/NET0131  & ~\g173_reg/NET0131  ;
  assign n2233 = ~\g172_reg/NET0131  & \g7961_pad  ;
  assign n2234 = ~n2232 & ~n2233 ;
  assign n2235 = ~n2231 & n2234 ;
  assign n2236 = ~\g163_reg/NET0131  & \g7961_pad  ;
  assign n2237 = \g1092_reg/NET0131  & ~\g164_reg/NET0131  ;
  assign n2238 = \g1088_reg/NET0131  & ~\g162_reg/NET0131  ;
  assign n2239 = ~n2237 & ~n2238 ;
  assign n2240 = ~n2236 & n2239 ;
  assign n2241 = ~n2235 & ~n2240 ;
  assign n2242 = n2235 & n2240 ;
  assign n2243 = ~n2241 & ~n2242 ;
  assign n2244 = \g1088_reg/NET0131  & ~\g168_reg/NET0131  ;
  assign n2245 = \g1092_reg/NET0131  & ~\g170_reg/NET0131  ;
  assign n2246 = ~\g169_reg/NET0131  & \g7961_pad  ;
  assign n2247 = ~n2245 & ~n2246 ;
  assign n2248 = ~n2244 & n2247 ;
  assign n2249 = \g1563_reg/NET0131  & ~n2248 ;
  assign n2250 = ~n2243 & n2249 ;
  assign n2251 = \g1088_reg/NET0131  & ~\g174_reg/NET0131  ;
  assign n2252 = \g1092_reg/NET0131  & ~\g176_reg/NET0131  ;
  assign n2253 = ~\g175_reg/NET0131  & \g7961_pad  ;
  assign n2254 = ~n2252 & ~n2253 ;
  assign n2255 = ~n2251 & n2254 ;
  assign n2256 = \g1092_reg/NET0131  & ~\g161_reg/NET0131  ;
  assign n2257 = \g1088_reg/NET0131  & ~\g159_reg/NET0131  ;
  assign n2258 = ~\g160_reg/NET0131  & \g7961_pad  ;
  assign n2259 = ~n2257 & ~n2258 ;
  assign n2260 = ~n2256 & n2259 ;
  assign n2261 = ~n2255 & ~n2260 ;
  assign n2262 = n2255 & n2260 ;
  assign n2263 = ~n2261 & ~n2262 ;
  assign n2264 = n2250 & ~n2263 ;
  assign n2265 = \g1088_reg/NET0131  & ~\g320_reg/NET0131  ;
  assign n2266 = ~\g318_reg/NET0131  & \g7961_pad  ;
  assign n2267 = \g1092_reg/NET0131  & ~\g319_reg/NET0131  ;
  assign n2268 = ~n2266 & ~n2267 ;
  assign n2269 = ~n2265 & n2268 ;
  assign n2270 = \g1088_reg/NET0131  & ~\g321_reg/NET0131  ;
  assign n2271 = \g1092_reg/NET0131  & ~\g323_reg/NET0131  ;
  assign n2272 = ~\g322_reg/NET0131  & \g7961_pad  ;
  assign n2273 = ~n2271 & ~n2272 ;
  assign n2274 = ~n2270 & n2273 ;
  assign n2275 = ~n2269 & ~n2274 ;
  assign n2276 = n2264 & n2275 ;
  assign n2277 = n2230 & n2276 ;
  assign n2278 = n2181 & n2277 ;
  assign n2279 = n2152 & n2278 ;
  assign n2280 = \g267_reg/NET0131  & \g7961_pad  ;
  assign n2281 = \g1088_reg/NET0131  & \g273_reg/NET0131  ;
  assign n2282 = \g1092_reg/NET0131  & \g270_reg/NET0131  ;
  assign n2283 = ~n2281 & ~n2282 ;
  assign n2284 = ~n2280 & n2283 ;
  assign n2285 = ~n2235 & ~n2284 ;
  assign n2286 = n2235 & n2284 ;
  assign n2287 = ~n2285 & ~n2286 ;
  assign n2288 = \g1092_reg/NET0131  & \g261_reg/NET0131  ;
  assign n2289 = \g1088_reg/NET0131  & \g264_reg/NET0131  ;
  assign n2290 = ~n2288 & ~n2289 ;
  assign n2291 = \g258_reg/NET0131  & \g7961_pad  ;
  assign n2292 = \g125_reg/NET0131  & ~n2291 ;
  assign n2293 = n2290 & n2292 ;
  assign n2294 = n2290 & ~n2291 ;
  assign n2295 = ~\g125_reg/NET0131  & ~n2294 ;
  assign n2296 = ~n2293 & ~n2295 ;
  assign n2297 = ~n2287 & n2296 ;
  assign n2298 = \g222_reg/NET0131  & \g7961_pad  ;
  assign n2299 = \g1088_reg/NET0131  & \g228_reg/NET0131  ;
  assign n2300 = \g1092_reg/NET0131  & \g225_reg/NET0131  ;
  assign n2301 = ~n2299 & ~n2300 ;
  assign n2302 = ~n2298 & n2301 ;
  assign n2303 = n2255 & n2302 ;
  assign n2304 = ~n2255 & ~n2302 ;
  assign n2305 = ~n2303 & ~n2304 ;
  assign n2306 = \g231_reg/NET0131  & \g7961_pad  ;
  assign n2307 = \g1088_reg/NET0131  & \g237_reg/NET0131  ;
  assign n2308 = ~n2306 & ~n2307 ;
  assign n2309 = \g1092_reg/NET0131  & \g234_reg/NET0131  ;
  assign n2310 = \g101_reg/NET0131  & ~n2309 ;
  assign n2311 = n2308 & n2310 ;
  assign n2312 = n2308 & ~n2309 ;
  assign n2313 = ~\g101_reg/NET0131  & ~n2312 ;
  assign n2314 = ~n2311 & ~n2313 ;
  assign n2315 = ~n2305 & n2314 ;
  assign n2316 = n2297 & n2315 ;
  assign n2317 = \g249_reg/NET0131  & \g7961_pad  ;
  assign n2318 = \g1088_reg/NET0131  & \g255_reg/NET0131  ;
  assign n2319 = ~n2317 & ~n2318 ;
  assign n2320 = \g1092_reg/NET0131  & \g252_reg/NET0131  ;
  assign n2321 = \g117_reg/NET0131  & ~n2320 ;
  assign n2322 = n2319 & n2321 ;
  assign n2323 = n2319 & ~n2320 ;
  assign n2324 = ~\g117_reg/NET0131  & ~n2323 ;
  assign n2325 = ~n2322 & ~n2324 ;
  assign n2326 = \g1088_reg/NET0131  & \g246_reg/NET0131  ;
  assign n2327 = \g1092_reg/NET0131  & \g243_reg/NET0131  ;
  assign n2328 = ~n2326 & ~n2327 ;
  assign n2329 = \g240_reg/NET0131  & \g7961_pad  ;
  assign n2330 = \g109_reg/NET0131  & ~n2329 ;
  assign n2331 = n2328 & n2330 ;
  assign n2332 = n2328 & ~n2329 ;
  assign n2333 = ~\g109_reg/NET0131  & ~n2332 ;
  assign n2334 = ~n2331 & ~n2333 ;
  assign n2335 = n2325 & n2334 ;
  assign n2336 = \g186_reg/NET0131  & \g7961_pad  ;
  assign n2337 = \g1092_reg/NET0131  & \g189_reg/NET0131  ;
  assign n2338 = ~n2336 & ~n2337 ;
  assign n2339 = \g1088_reg/NET0131  & \g192_reg/NET0131  ;
  assign n2340 = \g97_reg/NET0131  & ~n2339 ;
  assign n2341 = n2338 & n2340 ;
  assign n2342 = n2338 & ~n2339 ;
  assign n2343 = ~\g97_reg/NET0131  & ~n2342 ;
  assign n2344 = ~n2341 & ~n2343 ;
  assign n2345 = \g213_reg/NET0131  & \g7961_pad  ;
  assign n2346 = \g1092_reg/NET0131  & \g216_reg/NET0131  ;
  assign n2347 = \g1088_reg/NET0131  & \g219_reg/NET0131  ;
  assign n2348 = ~n2346 & ~n2347 ;
  assign n2349 = ~n2345 & n2348 ;
  assign n2350 = ~\g121_reg/NET0131  & ~n2349 ;
  assign n2351 = \g121_reg/NET0131  & ~n2345 ;
  assign n2352 = n2348 & n2351 ;
  assign n2353 = ~n2350 & ~n2352 ;
  assign n2354 = n2344 & n2353 ;
  assign n2355 = \g1088_reg/NET0131  & \g201_reg/NET0131  ;
  assign n2356 = \g1092_reg/NET0131  & \g198_reg/NET0131  ;
  assign n2357 = ~n2355 & ~n2356 ;
  assign n2358 = \g195_reg/NET0131  & \g7961_pad  ;
  assign n2359 = \g105_reg/NET0131  & ~n2358 ;
  assign n2360 = n2357 & n2359 ;
  assign n2361 = n2357 & ~n2358 ;
  assign n2362 = ~\g105_reg/NET0131  & ~n2361 ;
  assign n2363 = ~n2360 & ~n2362 ;
  assign n2364 = \g1088_reg/NET0131  & \g210_reg/NET0131  ;
  assign n2365 = \g204_reg/NET0131  & \g7961_pad  ;
  assign n2366 = \g1092_reg/NET0131  & \g207_reg/NET0131  ;
  assign n2367 = ~n2365 & ~n2366 ;
  assign n2368 = ~n2364 & n2367 ;
  assign n2369 = ~\g113_reg/NET0131  & ~n2368 ;
  assign n2370 = \g113_reg/NET0131  & ~n2364 ;
  assign n2371 = n2367 & n2370 ;
  assign n2372 = ~n2369 & ~n2371 ;
  assign n2373 = n2363 & n2372 ;
  assign n2374 = n2354 & n2373 ;
  assign n2375 = n2335 & n2374 ;
  assign n2376 = n2316 & n2375 ;
  assign n2377 = n2296 & n2314 ;
  assign n2378 = ~n2325 & ~n2377 ;
  assign n2379 = n2314 & n2334 ;
  assign n2380 = ~n2378 & n2379 ;
  assign n2381 = n2296 & n2325 ;
  assign n2382 = n2287 & ~n2381 ;
  assign n2383 = ~n2380 & n2382 ;
  assign n2384 = ~n2325 & ~n2334 ;
  assign n2385 = ~n2377 & n2384 ;
  assign n2386 = ~n2297 & ~n2314 ;
  assign n2387 = ~n2335 & n2386 ;
  assign n2388 = ~n2385 & ~n2387 ;
  assign n2389 = ~n2383 & n2388 ;
  assign n2390 = ~n2376 & n2389 ;
  assign n2391 = n2269 & ~n2390 ;
  assign n2392 = ~n2305 & n2363 ;
  assign n2393 = ~n2354 & ~n2392 ;
  assign n2394 = ~n2372 & n2393 ;
  assign n2395 = ~n2305 & n2353 ;
  assign n2396 = ~n2344 & ~n2373 ;
  assign n2397 = ~n2395 & n2396 ;
  assign n2398 = ~n2394 & ~n2397 ;
  assign n2399 = n2264 & ~n2274 ;
  assign n2400 = n2230 & n2399 ;
  assign n2401 = n2344 & n2363 ;
  assign n2402 = n2353 & n2372 ;
  assign n2403 = n2305 & ~n2402 ;
  assign n2404 = ~n2401 & n2403 ;
  assign n2405 = n2181 & ~n2404 ;
  assign n2406 = n2400 & n2405 ;
  assign n2407 = n2398 & n2406 ;
  assign n2408 = ~n2248 & ~n2407 ;
  assign n2409 = ~n2391 & n2408 ;
  assign n2410 = \g1563_reg/NET0131  & n2152 ;
  assign n2411 = ~n2409 & n2410 ;
  assign n2412 = ~n2279 & ~n2411 ;
  assign n2413 = n2269 & ~n2376 ;
  assign n2414 = n2389 & n2413 ;
  assign n2415 = n2151 & n2269 ;
  assign n2416 = n2146 & ~n2415 ;
  assign n2417 = ~n2404 & ~n2416 ;
  assign n2418 = n2398 & n2417 ;
  assign n2419 = ~n2414 & n2418 ;
  assign n2420 = ~\g315_reg/NET0131  & ~\g7961_pad  ;
  assign n2421 = \g1092_reg/NET0131  & ~\g404_reg/NET0131  ;
  assign n2422 = ~\g403_reg/NET0131  & \g7961_pad  ;
  assign n2423 = \g1088_reg/NET0131  & ~\g402_reg/NET0131  ;
  assign n2424 = ~n2422 & ~n2423 ;
  assign n2425 = ~n2421 & n2424 ;
  assign n2426 = n2264 & ~n2425 ;
  assign n2427 = n2230 & n2426 ;
  assign n2428 = n2181 & n2427 ;
  assign n2429 = ~n2151 & n2249 ;
  assign n2430 = ~n2416 & ~n2429 ;
  assign n2431 = ~n2428 & ~n2430 ;
  assign n2432 = ~n2420 & n2431 ;
  assign n2433 = ~n2419 & n2432 ;
  assign n2434 = n2412 & n2433 ;
  assign n2435 = ~n2141 & ~n2434 ;
  assign n2436 = ~\g1092_reg/NET0131  & \g316_reg/NET0131  ;
  assign n2437 = ~\g1092_reg/NET0131  & ~\g316_reg/NET0131  ;
  assign n2438 = n2431 & ~n2437 ;
  assign n2439 = ~n2419 & n2438 ;
  assign n2440 = n2412 & n2439 ;
  assign n2441 = ~n2436 & ~n2440 ;
  assign n2442 = ~\g1088_reg/NET0131  & \g317_reg/NET0131  ;
  assign n2443 = ~\g1088_reg/NET0131  & ~\g317_reg/NET0131  ;
  assign n2444 = n2431 & ~n2443 ;
  assign n2445 = ~n2419 & n2444 ;
  assign n2446 = n2412 & n2445 ;
  assign n2447 = ~n2442 & ~n2446 ;
  assign n2448 = \g1003_reg/NET0131  & ~\g1092_reg/NET0131  ;
  assign n2449 = ~\g1003_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n2450 = ~\g1004_reg/NET0131  & \g1088_reg/NET0131  ;
  assign n2451 = ~\g1002_reg/NET0131  & \g7961_pad  ;
  assign n2452 = ~n2450 & ~n2451 ;
  assign n2453 = ~n2449 & n2452 ;
  assign n2454 = ~\g1007_reg/NET0131  & \g1088_reg/NET0131  ;
  assign n2455 = ~\g1006_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n2456 = ~\g1005_reg/NET0131  & \g7961_pad  ;
  assign n2457 = ~n2455 & ~n2456 ;
  assign n2458 = ~n2454 & n2457 ;
  assign n2459 = \g1088_reg/NET0131  & ~\g856_reg/NET0131  ;
  assign n2460 = \g1092_reg/NET0131  & ~\g858_reg/NET0131  ;
  assign n2461 = ~n2459 & ~n2460 ;
  assign n2462 = \g7961_pad  & ~\g857_reg/NET0131  ;
  assign n2463 = \g1563_reg/NET0131  & ~n2462 ;
  assign n2464 = n2461 & n2463 ;
  assign n2465 = ~n2458 & ~n2464 ;
  assign n2466 = ~\g1001_reg/NET0131  & \g1088_reg/NET0131  ;
  assign n2467 = ~\g1000_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n2468 = \g7961_pad  & ~\g999_reg/NET0131  ;
  assign n2469 = ~n2467 & ~n2468 ;
  assign n2470 = ~n2466 & n2469 ;
  assign n2471 = ~n2465 & ~n2470 ;
  assign n2472 = \g7961_pad  & ~\g830_reg/NET0131  ;
  assign n2473 = \g1092_reg/NET0131  & ~\g831_reg/NET0131  ;
  assign n2474 = ~n2472 & ~n2473 ;
  assign n2475 = \g1088_reg/NET0131  & ~\g829_reg/NET0131  ;
  assign n2476 = \g793_reg/NET0131  & ~n2475 ;
  assign n2477 = n2474 & n2476 ;
  assign n2478 = n2474 & ~n2475 ;
  assign n2479 = ~\g793_reg/NET0131  & ~n2478 ;
  assign n2480 = ~n2477 & ~n2479 ;
  assign n2481 = \g7961_pad  & ~\g833_reg/NET0131  ;
  assign n2482 = \g1088_reg/NET0131  & ~\g832_reg/NET0131  ;
  assign n2483 = ~n2481 & ~n2482 ;
  assign n2484 = \g1092_reg/NET0131  & ~\g834_reg/NET0131  ;
  assign n2485 = \g797_reg/NET0131  & ~n2484 ;
  assign n2486 = n2483 & n2485 ;
  assign n2487 = n2483 & ~n2484 ;
  assign n2488 = ~\g797_reg/NET0131  & ~n2487 ;
  assign n2489 = ~n2486 & ~n2488 ;
  assign n2490 = n2480 & n2489 ;
  assign n2491 = \g7961_pad  & ~\g818_reg/NET0131  ;
  assign n2492 = \g1088_reg/NET0131  & ~\g817_reg/NET0131  ;
  assign n2493 = ~n2491 & ~n2492 ;
  assign n2494 = \g1092_reg/NET0131  & ~\g819_reg/NET0131  ;
  assign n2495 = \g785_reg/NET0131  & ~n2494 ;
  assign n2496 = n2493 & n2495 ;
  assign n2497 = n2493 & ~n2494 ;
  assign n2498 = ~\g785_reg/NET0131  & ~n2497 ;
  assign n2499 = ~n2496 & ~n2498 ;
  assign n2500 = \g7961_pad  & ~\g842_reg/NET0131  ;
  assign n2501 = \g1092_reg/NET0131  & ~\g843_reg/NET0131  ;
  assign n2502 = ~n2500 & ~n2501 ;
  assign n2503 = \g1088_reg/NET0131  & ~\g841_reg/NET0131  ;
  assign n2504 = \g809_reg/NET0131  & ~n2503 ;
  assign n2505 = n2502 & n2504 ;
  assign n2506 = n2502 & ~n2503 ;
  assign n2507 = ~\g809_reg/NET0131  & ~n2506 ;
  assign n2508 = ~n2505 & ~n2507 ;
  assign n2509 = n2499 & n2508 ;
  assign n2510 = n2490 & n2509 ;
  assign n2511 = \g1088_reg/NET0131  & ~\g859_reg/NET0131  ;
  assign n2512 = \g7961_pad  & ~\g860_reg/NET0131  ;
  assign n2513 = \g1092_reg/NET0131  & ~\g861_reg/NET0131  ;
  assign n2514 = ~n2512 & ~n2513 ;
  assign n2515 = ~n2511 & n2514 ;
  assign n2516 = \g7961_pad  & ~\g851_reg/NET0131  ;
  assign n2517 = \g1088_reg/NET0131  & ~\g850_reg/NET0131  ;
  assign n2518 = \g1092_reg/NET0131  & ~\g852_reg/NET0131  ;
  assign n2519 = ~n2517 & ~n2518 ;
  assign n2520 = ~n2516 & n2519 ;
  assign n2521 = ~n2515 & ~n2520 ;
  assign n2522 = n2515 & n2520 ;
  assign n2523 = ~n2521 & ~n2522 ;
  assign n2524 = \g1088_reg/NET0131  & ~\g838_reg/NET0131  ;
  assign n2525 = \g1092_reg/NET0131  & ~\g840_reg/NET0131  ;
  assign n2526 = ~n2524 & ~n2525 ;
  assign n2527 = \g7961_pad  & ~\g839_reg/NET0131  ;
  assign n2528 = \g805_reg/NET0131  & ~n2527 ;
  assign n2529 = n2526 & n2528 ;
  assign n2530 = \g7961_pad  & ~\g821_reg/NET0131  ;
  assign n2531 = \g1092_reg/NET0131  & ~\g822_reg/NET0131  ;
  assign n2532 = ~n2530 & ~n2531 ;
  assign n2533 = \g1088_reg/NET0131  & ~\g820_reg/NET0131  ;
  assign n2534 = n2532 & ~n2533 ;
  assign n2535 = ~\g789_reg/NET0131  & ~n2534 ;
  assign n2536 = ~n2529 & ~n2535 ;
  assign n2537 = ~n2523 & n2536 ;
  assign n2538 = \g789_reg/NET0131  & ~n2533 ;
  assign n2539 = n2532 & n2538 ;
  assign n2540 = n2461 & ~n2462 ;
  assign n2541 = \g1563_reg/NET0131  & ~n2540 ;
  assign n2542 = n2526 & ~n2527 ;
  assign n2543 = ~\g805_reg/NET0131  & ~n2542 ;
  assign n2544 = n2541 & ~n2543 ;
  assign n2545 = ~n2539 & n2544 ;
  assign n2546 = n2537 & n2545 ;
  assign n2547 = n2510 & n2546 ;
  assign n2548 = \g7961_pad  & ~\g836_reg/NET0131  ;
  assign n2549 = \g1092_reg/NET0131  & ~\g837_reg/NET0131  ;
  assign n2550 = ~n2548 & ~n2549 ;
  assign n2551 = \g1088_reg/NET0131  & ~\g835_reg/NET0131  ;
  assign n2552 = \g801_reg/NET0131  & ~n2551 ;
  assign n2553 = n2550 & n2552 ;
  assign n2554 = n2550 & ~n2551 ;
  assign n2555 = ~\g801_reg/NET0131  & ~n2554 ;
  assign n2556 = ~n2553 & ~n2555 ;
  assign n2557 = \g1088_reg/NET0131  & ~\g862_reg/NET0131  ;
  assign n2558 = \g7961_pad  & ~\g863_reg/NET0131  ;
  assign n2559 = \g1092_reg/NET0131  & ~\g864_reg/NET0131  ;
  assign n2560 = ~n2558 & ~n2559 ;
  assign n2561 = ~n2557 & n2560 ;
  assign n2562 = \g7961_pad  & ~\g848_reg/NET0131  ;
  assign n2563 = \g1092_reg/NET0131  & ~\g849_reg/NET0131  ;
  assign n2564 = \g1088_reg/NET0131  & ~\g847_reg/NET0131  ;
  assign n2565 = ~n2563 & ~n2564 ;
  assign n2566 = ~n2562 & n2565 ;
  assign n2567 = ~n2561 & ~n2566 ;
  assign n2568 = n2561 & n2566 ;
  assign n2569 = ~n2567 & ~n2568 ;
  assign n2570 = n2556 & ~n2569 ;
  assign n2571 = ~\g1009_reg/NET0131  & \g7961_pad  ;
  assign n2572 = ~\g1010_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n2573 = ~\g1008_reg/NET0131  & \g1088_reg/NET0131  ;
  assign n2574 = ~n2572 & ~n2573 ;
  assign n2575 = ~n2571 & n2574 ;
  assign n2576 = \g1088_reg/NET0131  & ~\g844_reg/NET0131  ;
  assign n2577 = \g1092_reg/NET0131  & ~\g846_reg/NET0131  ;
  assign n2578 = ~n2576 & ~n2577 ;
  assign n2579 = \g7961_pad  & ~\g845_reg/NET0131  ;
  assign n2580 = \g813_reg/NET0131  & ~n2579 ;
  assign n2581 = n2578 & n2580 ;
  assign n2582 = n2578 & ~n2579 ;
  assign n2583 = ~\g813_reg/NET0131  & ~n2582 ;
  assign n2584 = ~n2581 & ~n2583 ;
  assign n2585 = ~n2575 & n2584 ;
  assign n2586 = n2570 & n2585 ;
  assign n2587 = ~n2470 & n2586 ;
  assign n2588 = n2547 & n2587 ;
  assign n2589 = ~n2471 & ~n2588 ;
  assign n2590 = n2453 & ~n2589 ;
  assign n2591 = n2570 & n2584 ;
  assign n2592 = ~\g1090_reg/NET0131  & \g7961_pad  ;
  assign n2593 = ~\g1091_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n2594 = \g1088_reg/NET0131  & ~\g1089_reg/NET0131  ;
  assign n2595 = ~n2593 & ~n2594 ;
  assign n2596 = ~n2592 & n2595 ;
  assign n2597 = n2591 & ~n2596 ;
  assign n2598 = n2547 & n2597 ;
  assign n2599 = n2458 & n2470 ;
  assign n2600 = n2453 & n2599 ;
  assign n2601 = ~n2598 & ~n2600 ;
  assign n2602 = ~n2590 & n2601 ;
  assign n2603 = \g1088_reg/NET0131  & \g897_reg/NET0131  ;
  assign n2604 = \g7961_pad  & \g891_reg/NET0131  ;
  assign n2605 = \g1092_reg/NET0131  & \g894_reg/NET0131  ;
  assign n2606 = ~n2604 & ~n2605 ;
  assign n2607 = ~n2603 & n2606 ;
  assign n2608 = ~\g801_reg/NET0131  & ~n2607 ;
  assign n2609 = \g801_reg/NET0131  & ~n2603 ;
  assign n2610 = n2606 & n2609 ;
  assign n2611 = ~n2608 & ~n2610 ;
  assign n2612 = \g7961_pad  & \g909_reg/NET0131  ;
  assign n2613 = \g1088_reg/NET0131  & \g915_reg/NET0131  ;
  assign n2614 = \g1092_reg/NET0131  & \g912_reg/NET0131  ;
  assign n2615 = ~n2613 & ~n2614 ;
  assign n2616 = ~n2612 & n2615 ;
  assign n2617 = ~n2561 & ~n2616 ;
  assign n2618 = n2561 & n2616 ;
  assign n2619 = ~n2617 & ~n2618 ;
  assign n2620 = \g7961_pad  & \g882_reg/NET0131  ;
  assign n2621 = \g1088_reg/NET0131  & \g888_reg/NET0131  ;
  assign n2622 = \g1092_reg/NET0131  & \g885_reg/NET0131  ;
  assign n2623 = ~n2621 & ~n2622 ;
  assign n2624 = ~n2620 & n2623 ;
  assign n2625 = ~\g793_reg/NET0131  & ~n2624 ;
  assign n2626 = \g793_reg/NET0131  & ~n2620 ;
  assign n2627 = n2623 & n2626 ;
  assign n2628 = ~n2625 & ~n2627 ;
  assign n2629 = ~n2619 & n2628 ;
  assign n2630 = ~n2611 & ~n2629 ;
  assign n2631 = \g7961_pad  & \g900_reg/NET0131  ;
  assign n2632 = \g1092_reg/NET0131  & \g903_reg/NET0131  ;
  assign n2633 = \g1088_reg/NET0131  & \g906_reg/NET0131  ;
  assign n2634 = ~n2632 & ~n2633 ;
  assign n2635 = ~n2631 & n2634 ;
  assign n2636 = ~\g809_reg/NET0131  & ~n2635 ;
  assign n2637 = \g809_reg/NET0131  & ~n2631 ;
  assign n2638 = n2634 & n2637 ;
  assign n2639 = ~n2636 & ~n2638 ;
  assign n2640 = ~n2619 & n2639 ;
  assign n2641 = ~n2630 & n2640 ;
  assign n2642 = \g7961_pad  & \g873_reg/NET0131  ;
  assign n2643 = \g1092_reg/NET0131  & \g876_reg/NET0131  ;
  assign n2644 = ~n2642 & ~n2643 ;
  assign n2645 = \g1088_reg/NET0131  & \g879_reg/NET0131  ;
  assign n2646 = \g785_reg/NET0131  & ~n2645 ;
  assign n2647 = n2644 & n2646 ;
  assign n2648 = n2644 & ~n2645 ;
  assign n2649 = ~\g785_reg/NET0131  & ~n2648 ;
  assign n2650 = ~n2647 & ~n2649 ;
  assign n2651 = n2611 & n2628 ;
  assign n2652 = ~n2650 & ~n2651 ;
  assign n2653 = ~n2641 & n2652 ;
  assign n2654 = ~n2611 & ~n2639 ;
  assign n2655 = ~n2629 & n2654 ;
  assign n2656 = n2611 & n2639 ;
  assign n2657 = n2628 & n2650 ;
  assign n2658 = ~n2656 & ~n2657 ;
  assign n2659 = n2619 & n2658 ;
  assign n2660 = ~n2655 & ~n2659 ;
  assign n2661 = ~n2653 & n2660 ;
  assign n2662 = n2541 & ~n2661 ;
  assign n2663 = \g1563_reg/NET0131  & n2586 ;
  assign n2664 = n2547 & n2663 ;
  assign n2665 = ~n2662 & n2664 ;
  assign n2666 = \g7961_pad  & \g927_reg/NET0131  ;
  assign n2667 = \g1088_reg/NET0131  & \g933_reg/NET0131  ;
  assign n2668 = \g1092_reg/NET0131  & \g930_reg/NET0131  ;
  assign n2669 = ~n2667 & ~n2668 ;
  assign n2670 = ~n2666 & n2669 ;
  assign n2671 = ~\g797_reg/NET0131  & ~n2670 ;
  assign n2672 = \g797_reg/NET0131  & ~n2666 ;
  assign n2673 = n2669 & n2672 ;
  assign n2674 = ~n2671 & ~n2673 ;
  assign n2675 = \g7961_pad  & \g954_reg/NET0131  ;
  assign n2676 = \g1088_reg/NET0131  & \g960_reg/NET0131  ;
  assign n2677 = \g1092_reg/NET0131  & \g957_reg/NET0131  ;
  assign n2678 = ~n2676 & ~n2677 ;
  assign n2679 = ~n2675 & n2678 ;
  assign n2680 = ~n2515 & ~n2679 ;
  assign n2681 = n2515 & n2679 ;
  assign n2682 = ~n2680 & ~n2681 ;
  assign n2683 = n2674 & ~n2682 ;
  assign n2684 = \g7961_pad  & \g918_reg/NET0131  ;
  assign n2685 = \g1088_reg/NET0131  & \g924_reg/NET0131  ;
  assign n2686 = \g1092_reg/NET0131  & \g921_reg/NET0131  ;
  assign n2687 = ~n2685 & ~n2686 ;
  assign n2688 = ~n2684 & n2687 ;
  assign n2689 = ~\g789_reg/NET0131  & ~n2688 ;
  assign n2690 = \g789_reg/NET0131  & ~n2684 ;
  assign n2691 = n2687 & n2690 ;
  assign n2692 = ~n2689 & ~n2691 ;
  assign n2693 = n2674 & n2692 ;
  assign n2694 = n2682 & ~n2693 ;
  assign n2695 = \g1092_reg/NET0131  & \g948_reg/NET0131  ;
  assign n2696 = \g7961_pad  & \g945_reg/NET0131  ;
  assign n2697 = \g1088_reg/NET0131  & \g951_reg/NET0131  ;
  assign n2698 = ~n2696 & ~n2697 ;
  assign n2699 = ~n2695 & n2698 ;
  assign n2700 = ~\g813_reg/NET0131  & ~n2699 ;
  assign n2701 = \g813_reg/NET0131  & ~n2695 ;
  assign n2702 = n2698 & n2701 ;
  assign n2703 = ~n2700 & ~n2702 ;
  assign n2704 = n2692 & n2703 ;
  assign n2705 = ~n2694 & n2704 ;
  assign n2706 = ~n2683 & ~n2705 ;
  assign n2707 = \g1088_reg/NET0131  & \g942_reg/NET0131  ;
  assign n2708 = \g7961_pad  & \g936_reg/NET0131  ;
  assign n2709 = \g1092_reg/NET0131  & \g939_reg/NET0131  ;
  assign n2710 = ~n2708 & ~n2709 ;
  assign n2711 = ~n2707 & n2710 ;
  assign n2712 = ~\g805_reg/NET0131  & ~n2711 ;
  assign n2713 = \g805_reg/NET0131  & ~n2707 ;
  assign n2714 = n2710 & n2713 ;
  assign n2715 = ~n2712 & ~n2714 ;
  assign n2716 = n2682 & ~n2703 ;
  assign n2717 = ~n2693 & n2716 ;
  assign n2718 = n2715 & ~n2717 ;
  assign n2719 = n2541 & ~n2718 ;
  assign n2720 = n2706 & n2719 ;
  assign n2721 = n2674 & n2715 ;
  assign n2722 = ~n2682 & n2703 ;
  assign n2723 = ~n2721 & ~n2722 ;
  assign n2724 = n2541 & ~n2692 ;
  assign n2725 = n2723 & n2724 ;
  assign n2726 = ~n2600 & ~n2725 ;
  assign n2727 = ~n2598 & n2726 ;
  assign n2728 = ~n2720 & n2727 ;
  assign n2729 = \g1563_reg/NET0131  & n2540 ;
  assign n2730 = n2657 & n2722 ;
  assign n2731 = n2656 & n2730 ;
  assign n2732 = ~n2619 & n2692 ;
  assign n2733 = n2721 & n2732 ;
  assign n2734 = \g1563_reg/NET0131  & n2733 ;
  assign n2735 = n2731 & n2734 ;
  assign n2736 = ~n2729 & ~n2735 ;
  assign n2737 = n2458 & n2736 ;
  assign n2738 = n2728 & n2737 ;
  assign n2739 = ~n2665 & n2738 ;
  assign n2740 = ~n2602 & ~n2739 ;
  assign n2741 = ~\g1003_reg/NET0131  & ~\g1092_reg/NET0131  ;
  assign n2742 = n2731 & n2733 ;
  assign n2743 = ~n2470 & ~n2742 ;
  assign n2744 = n2706 & ~n2718 ;
  assign n2745 = ~n2692 & n2723 ;
  assign n2746 = n2458 & n2541 ;
  assign n2747 = ~n2745 & n2746 ;
  assign n2748 = ~n2744 & n2747 ;
  assign n2749 = n2743 & n2748 ;
  assign n2750 = ~n2470 & n2541 ;
  assign n2751 = ~n2661 & n2750 ;
  assign n2752 = ~n2453 & ~n2751 ;
  assign n2753 = ~n2749 & n2752 ;
  assign n2754 = ~n2741 & ~n2753 ;
  assign n2755 = ~n2740 & n2754 ;
  assign n2756 = ~n2448 & ~n2755 ;
  assign n2757 = \g1092_reg/NET0131  & ~n1472 ;
  assign n2758 = ~n1463 & n2757 ;
  assign n2759 = ~\g1092_reg/NET0131  & ~\g2391_reg/NET0131  ;
  assign n2760 = ~n2758 & ~n2759 ;
  assign n2761 = \g1088_reg/NET0131  & ~n1472 ;
  assign n2762 = ~n1463 & n2761 ;
  assign n2763 = ~\g1088_reg/NET0131  & ~\g2392_reg/NET0131  ;
  assign n2764 = ~n2762 & ~n2763 ;
  assign n2765 = \g1004_reg/NET0131  & ~\g1088_reg/NET0131  ;
  assign n2766 = ~\g1004_reg/NET0131  & ~\g1088_reg/NET0131  ;
  assign n2767 = ~n2753 & ~n2766 ;
  assign n2768 = ~n2740 & n2767 ;
  assign n2769 = ~n2765 & ~n2768 ;
  assign n2770 = \g1002_reg/NET0131  & ~\g7961_pad  ;
  assign n2771 = ~\g1002_reg/NET0131  & ~\g7961_pad  ;
  assign n2772 = ~n2753 & ~n2771 ;
  assign n2773 = ~n2740 & n2772 ;
  assign n2774 = ~n2770 & ~n2773 ;
  assign n2775 = \g1088_reg/NET0131  & ~\g1550_reg/NET0131  ;
  assign n2776 = \g1092_reg/NET0131  & ~\g1552_reg/NET0131  ;
  assign n2777 = ~\g1551_reg/NET0131  & \g7961_pad  ;
  assign n2778 = ~n2776 & ~n2777 ;
  assign n2779 = ~n2775 & n2778 ;
  assign n2780 = \g1563_reg/NET0131  & ~n2779 ;
  assign n2781 = \g1088_reg/NET0131  & ~\g1556_reg/NET0131  ;
  assign n2782 = \g1092_reg/NET0131  & ~\g1558_reg/NET0131  ;
  assign n2783 = ~\g1557_reg/NET0131  & \g7961_pad  ;
  assign n2784 = ~n2782 & ~n2783 ;
  assign n2785 = ~n2781 & n2784 ;
  assign n2786 = \g1603_reg/NET0131  & \g7961_pad  ;
  assign n2787 = \g1088_reg/NET0131  & \g1609_reg/NET0131  ;
  assign n2788 = \g1092_reg/NET0131  & \g1606_reg/NET0131  ;
  assign n2789 = ~n2787 & ~n2788 ;
  assign n2790 = ~n2786 & n2789 ;
  assign n2791 = ~n2785 & ~n2790 ;
  assign n2792 = n2785 & n2790 ;
  assign n2793 = ~n2791 & ~n2792 ;
  assign n2794 = \g1594_reg/NET0131  & \g7961_pad  ;
  assign n2795 = \g1092_reg/NET0131  & \g1597_reg/NET0131  ;
  assign n2796 = \g1088_reg/NET0131  & \g1600_reg/NET0131  ;
  assign n2797 = ~n2795 & ~n2796 ;
  assign n2798 = ~n2794 & n2797 ;
  assign n2799 = ~\g1501_reg/NET0131  & ~n2798 ;
  assign n2800 = \g1501_reg/NET0131  & ~n2794 ;
  assign n2801 = n2797 & n2800 ;
  assign n2802 = ~n2799 & ~n2801 ;
  assign n2803 = \g1088_reg/NET0131  & \g1591_reg/NET0131  ;
  assign n2804 = \g1585_reg/NET0131  & \g7961_pad  ;
  assign n2805 = \g1092_reg/NET0131  & \g1588_reg/NET0131  ;
  assign n2806 = ~n2804 & ~n2805 ;
  assign n2807 = ~n2803 & n2806 ;
  assign n2808 = ~\g1491_reg/NET0131  & ~n2807 ;
  assign n2809 = \g1491_reg/NET0131  & ~n2803 ;
  assign n2810 = n2806 & n2809 ;
  assign n2811 = ~n2808 & ~n2810 ;
  assign n2812 = n2802 & n2811 ;
  assign n2813 = \g1567_reg/NET0131  & \g7961_pad  ;
  assign n2814 = \g1088_reg/NET0131  & \g1573_reg/NET0131  ;
  assign n2815 = ~n2813 & ~n2814 ;
  assign n2816 = \g1092_reg/NET0131  & \g1570_reg/NET0131  ;
  assign n2817 = \g1471_reg/NET0131  & ~n2816 ;
  assign n2818 = n2815 & n2817 ;
  assign n2819 = n2815 & ~n2816 ;
  assign n2820 = ~\g1471_reg/NET0131  & ~n2819 ;
  assign n2821 = ~n2818 & ~n2820 ;
  assign n2822 = \g1576_reg/NET0131  & \g7961_pad  ;
  assign n2823 = \g1088_reg/NET0131  & \g1582_reg/NET0131  ;
  assign n2824 = \g1092_reg/NET0131  & \g1579_reg/NET0131  ;
  assign n2825 = ~n2823 & ~n2824 ;
  assign n2826 = ~n2822 & n2825 ;
  assign n2827 = ~\g1481_reg/NET0131  & ~n2826 ;
  assign n2828 = \g1481_reg/NET0131  & ~n2822 ;
  assign n2829 = n2825 & n2828 ;
  assign n2830 = ~n2827 & ~n2829 ;
  assign n2831 = n2821 & n2830 ;
  assign n2832 = ~n2812 & ~n2831 ;
  assign n2833 = n2793 & n2832 ;
  assign n2834 = ~n2793 & n2830 ;
  assign n2835 = n2802 & n2821 ;
  assign n2836 = ~n2811 & ~n2835 ;
  assign n2837 = ~n2834 & n2836 ;
  assign n2838 = ~n2793 & n2802 ;
  assign n2839 = n2811 & n2830 ;
  assign n2840 = ~n2821 & ~n2839 ;
  assign n2841 = ~n2838 & n2840 ;
  assign n2842 = ~n2837 & ~n2841 ;
  assign n2843 = ~n2833 & n2842 ;
  assign n2844 = n2780 & ~n2843 ;
  assign n2845 = \g1088_reg/NET0131  & ~\g1529_reg/NET0131  ;
  assign n2846 = \g1092_reg/NET0131  & ~\g1531_reg/NET0131  ;
  assign n2847 = ~n2845 & ~n2846 ;
  assign n2848 = ~\g1530_reg/NET0131  & \g7961_pad  ;
  assign n2849 = \g1491_reg/NET0131  & ~n2848 ;
  assign n2850 = n2847 & n2849 ;
  assign n2851 = n2847 & ~n2848 ;
  assign n2852 = ~\g1491_reg/NET0131  & ~n2851 ;
  assign n2853 = ~n2850 & ~n2852 ;
  assign n2854 = ~\g1515_reg/NET0131  & \g7961_pad  ;
  assign n2855 = \g1088_reg/NET0131  & ~\g1514_reg/NET0131  ;
  assign n2856 = ~n2854 & ~n2855 ;
  assign n2857 = \g1092_reg/NET0131  & ~\g1516_reg/NET0131  ;
  assign n2858 = \g1476_reg/NET0131  & ~n2857 ;
  assign n2859 = n2856 & n2858 ;
  assign n2860 = n2856 & ~n2857 ;
  assign n2861 = ~\g1476_reg/NET0131  & ~n2860 ;
  assign n2862 = ~n2859 & ~n2861 ;
  assign n2863 = n2853 & n2862 ;
  assign n2864 = \g1092_reg/NET0131  & ~\g1537_reg/NET0131  ;
  assign n2865 = \g1088_reg/NET0131  & ~\g1535_reg/NET0131  ;
  assign n2866 = ~n2864 & ~n2865 ;
  assign n2867 = ~\g1536_reg/NET0131  & \g7961_pad  ;
  assign n2868 = \g1501_reg/NET0131  & ~n2867 ;
  assign n2869 = n2866 & n2868 ;
  assign n2870 = n2866 & ~n2867 ;
  assign n2871 = ~\g1501_reg/NET0131  & ~n2870 ;
  assign n2872 = ~n2869 & ~n2871 ;
  assign n2873 = ~\g1539_reg/NET0131  & \g7961_pad  ;
  assign n2874 = \g1088_reg/NET0131  & ~\g1538_reg/NET0131  ;
  assign n2875 = ~n2873 & ~n2874 ;
  assign n2876 = \g1092_reg/NET0131  & ~\g1540_reg/NET0131  ;
  assign n2877 = \g1506_reg/NET0131  & ~n2876 ;
  assign n2878 = n2875 & n2877 ;
  assign n2879 = n2875 & ~n2876 ;
  assign n2880 = ~\g1506_reg/NET0131  & ~n2879 ;
  assign n2881 = ~n2878 & ~n2880 ;
  assign n2882 = n2872 & n2881 ;
  assign n2883 = n2863 & n2882 ;
  assign n2884 = ~\g1527_reg/NET0131  & \g7961_pad  ;
  assign n2885 = \g1088_reg/NET0131  & ~\g1526_reg/NET0131  ;
  assign n2886 = ~n2884 & ~n2885 ;
  assign n2887 = \g1092_reg/NET0131  & ~\g1528_reg/NET0131  ;
  assign n2888 = \g1486_reg/NET0131  & ~n2887 ;
  assign n2889 = n2886 & n2888 ;
  assign n2890 = n2886 & ~n2887 ;
  assign n2891 = ~\g1486_reg/NET0131  & ~n2890 ;
  assign n2892 = ~n2889 & ~n2891 ;
  assign n2893 = ~\g1512_reg/NET0131  & \g7961_pad  ;
  assign n2894 = \g1088_reg/NET0131  & ~\g1511_reg/NET0131  ;
  assign n2895 = ~n2893 & ~n2894 ;
  assign n2896 = \g1092_reg/NET0131  & ~\g1513_reg/NET0131  ;
  assign n2897 = \g1471_reg/NET0131  & ~n2896 ;
  assign n2898 = n2895 & n2897 ;
  assign n2899 = n2895 & ~n2896 ;
  assign n2900 = ~\g1471_reg/NET0131  & ~n2899 ;
  assign n2901 = ~n2898 & ~n2900 ;
  assign n2902 = n2892 & n2901 ;
  assign n2903 = \g1092_reg/NET0131  & ~\g1525_reg/NET0131  ;
  assign n2904 = ~\g1524_reg/NET0131  & \g7961_pad  ;
  assign n2905 = ~n2903 & ~n2904 ;
  assign n2906 = \g1088_reg/NET0131  & ~\g1523_reg/NET0131  ;
  assign n2907 = \g1481_reg/NET0131  & ~n2906 ;
  assign n2908 = n2905 & n2907 ;
  assign n2909 = n2905 & ~n2906 ;
  assign n2910 = ~\g1481_reg/NET0131  & ~n2909 ;
  assign n2911 = ~n2908 & ~n2910 ;
  assign n2912 = n2780 & n2911 ;
  assign n2913 = n2902 & n2912 ;
  assign n2914 = n2883 & n2913 ;
  assign n2915 = \g1092_reg/NET0131  & ~\g1534_reg/NET0131  ;
  assign n2916 = \g1088_reg/NET0131  & ~\g1532_reg/NET0131  ;
  assign n2917 = ~n2915 & ~n2916 ;
  assign n2918 = ~\g1533_reg/NET0131  & \g7961_pad  ;
  assign n2919 = \g1496_reg/NET0131  & ~n2918 ;
  assign n2920 = n2917 & n2919 ;
  assign n2921 = n2917 & ~n2918 ;
  assign n2922 = ~\g1496_reg/NET0131  & ~n2921 ;
  assign n2923 = ~n2920 & ~n2922 ;
  assign n2924 = \g1088_reg/NET0131  & ~\g1553_reg/NET0131  ;
  assign n2925 = \g1092_reg/NET0131  & ~\g1555_reg/NET0131  ;
  assign n2926 = ~\g1554_reg/NET0131  & \g7961_pad  ;
  assign n2927 = ~n2925 & ~n2926 ;
  assign n2928 = ~n2924 & n2927 ;
  assign n2929 = ~\g1545_reg/NET0131  & \g7961_pad  ;
  assign n2930 = \g1092_reg/NET0131  & ~\g1546_reg/NET0131  ;
  assign n2931 = \g1088_reg/NET0131  & ~\g1544_reg/NET0131  ;
  assign n2932 = ~n2930 & ~n2931 ;
  assign n2933 = ~n2929 & n2932 ;
  assign n2934 = ~n2928 & ~n2933 ;
  assign n2935 = n2928 & n2933 ;
  assign n2936 = ~n2934 & ~n2935 ;
  assign n2937 = n2923 & ~n2936 ;
  assign n2938 = ~\g1542_reg/NET0131  & \g7961_pad  ;
  assign n2939 = \g1092_reg/NET0131  & ~\g1543_reg/NET0131  ;
  assign n2940 = \g1088_reg/NET0131  & ~\g1541_reg/NET0131  ;
  assign n2941 = ~n2939 & ~n2940 ;
  assign n2942 = ~n2938 & n2941 ;
  assign n2943 = ~n2785 & ~n2942 ;
  assign n2944 = n2785 & n2942 ;
  assign n2945 = ~n2943 & ~n2944 ;
  assign n2946 = \g1088_reg/NET0131  & ~\g1702_reg/NET0131  ;
  assign n2947 = ~\g1703_reg/NET0131  & \g7961_pad  ;
  assign n2948 = \g1092_reg/NET0131  & ~\g1704_reg/NET0131  ;
  assign n2949 = ~n2947 & ~n2948 ;
  assign n2950 = ~n2946 & n2949 ;
  assign n2951 = ~n2945 & ~n2950 ;
  assign n2952 = n2937 & n2951 ;
  assign n2953 = \g1563_reg/NET0131  & n2952 ;
  assign n2954 = n2914 & n2953 ;
  assign n2955 = ~n2844 & n2954 ;
  assign n2956 = \g1630_reg/NET0131  & \g7961_pad  ;
  assign n2957 = \g1088_reg/NET0131  & \g1636_reg/NET0131  ;
  assign n2958 = ~n2956 & ~n2957 ;
  assign n2959 = \g1092_reg/NET0131  & \g1633_reg/NET0131  ;
  assign n2960 = \g1496_reg/NET0131  & ~n2959 ;
  assign n2961 = n2958 & n2960 ;
  assign n2962 = n2958 & ~n2959 ;
  assign n2963 = ~\g1496_reg/NET0131  & ~n2962 ;
  assign n2964 = ~n2961 & ~n2963 ;
  assign n2965 = \g1612_reg/NET0131  & \g7961_pad  ;
  assign n2966 = \g1088_reg/NET0131  & \g1618_reg/NET0131  ;
  assign n2967 = \g1092_reg/NET0131  & \g1615_reg/NET0131  ;
  assign n2968 = ~n2966 & ~n2967 ;
  assign n2969 = ~n2965 & n2968 ;
  assign n2970 = ~\g1476_reg/NET0131  & ~n2969 ;
  assign n2971 = \g1476_reg/NET0131  & ~n2965 ;
  assign n2972 = n2968 & n2971 ;
  assign n2973 = ~n2970 & ~n2972 ;
  assign n2974 = \g1639_reg/NET0131  & \g7961_pad  ;
  assign n2975 = \g1092_reg/NET0131  & \g1642_reg/NET0131  ;
  assign n2976 = \g1088_reg/NET0131  & \g1645_reg/NET0131  ;
  assign n2977 = ~n2975 & ~n2976 ;
  assign n2978 = ~n2974 & n2977 ;
  assign n2979 = ~\g1506_reg/NET0131  & ~n2978 ;
  assign n2980 = \g1506_reg/NET0131  & ~n2974 ;
  assign n2981 = n2977 & n2980 ;
  assign n2982 = ~n2979 & ~n2981 ;
  assign n2983 = n2973 & n2982 ;
  assign n2984 = ~n2964 & ~n2983 ;
  assign n2985 = \g1092_reg/NET0131  & \g1624_reg/NET0131  ;
  assign n2986 = \g1088_reg/NET0131  & \g1627_reg/NET0131  ;
  assign n2987 = ~n2985 & ~n2986 ;
  assign n2988 = \g1621_reg/NET0131  & \g7961_pad  ;
  assign n2989 = \g1486_reg/NET0131  & ~n2988 ;
  assign n2990 = n2987 & n2989 ;
  assign n2991 = n2987 & ~n2988 ;
  assign n2992 = ~\g1486_reg/NET0131  & ~n2991 ;
  assign n2993 = ~n2990 & ~n2992 ;
  assign n2994 = n2973 & n2993 ;
  assign n2995 = ~n2984 & n2994 ;
  assign n2996 = \g1648_reg/NET0131  & \g7961_pad  ;
  assign n2997 = \g1088_reg/NET0131  & \g1654_reg/NET0131  ;
  assign n2998 = \g1092_reg/NET0131  & \g1651_reg/NET0131  ;
  assign n2999 = ~n2997 & ~n2998 ;
  assign n3000 = ~n2996 & n2999 ;
  assign n3001 = ~n2928 & ~n3000 ;
  assign n3002 = n2928 & n3000 ;
  assign n3003 = ~n3001 & ~n3002 ;
  assign n3004 = n2964 & n2982 ;
  assign n3005 = n3003 & ~n3004 ;
  assign n3006 = ~n2995 & n3005 ;
  assign n3007 = ~n2964 & ~n2993 ;
  assign n3008 = ~n2983 & n3007 ;
  assign n3009 = n2982 & ~n3003 ;
  assign n3010 = n2964 & n2993 ;
  assign n3011 = ~n2973 & ~n3010 ;
  assign n3012 = ~n3009 & n3011 ;
  assign n3013 = ~n3008 & ~n3012 ;
  assign n3014 = ~n3006 & n3013 ;
  assign n3015 = n2780 & ~n3014 ;
  assign n3016 = \g1092_reg/NET0131  & ~\g1700_reg/NET0131  ;
  assign n3017 = ~\g1699_reg/NET0131  & \g7961_pad  ;
  assign n3018 = \g1088_reg/NET0131  & ~\g1701_reg/NET0131  ;
  assign n3019 = ~n3017 & ~n3018 ;
  assign n3020 = ~n3016 & n3019 ;
  assign n3021 = \g1563_reg/NET0131  & n2779 ;
  assign n3022 = n2834 & n3010 ;
  assign n3023 = n3009 & n3022 ;
  assign n3024 = n2821 & n2973 ;
  assign n3025 = n2812 & n3024 ;
  assign n3026 = \g1563_reg/NET0131  & n3025 ;
  assign n3027 = n3023 & n3026 ;
  assign n3028 = ~n3021 & ~n3027 ;
  assign n3029 = n3020 & n3028 ;
  assign n3030 = ~n3015 & n3029 ;
  assign n3031 = ~n2955 & n3030 ;
  assign n3032 = \g1088_reg/NET0131  & ~\g1695_reg/NET0131  ;
  assign n3033 = ~\g1693_reg/NET0131  & \g7961_pad  ;
  assign n3034 = \g1092_reg/NET0131  & ~\g1694_reg/NET0131  ;
  assign n3035 = ~n3033 & ~n3034 ;
  assign n3036 = ~n3032 & n3035 ;
  assign n3037 = \g1563_reg/NET0131  & ~n2775 ;
  assign n3038 = n2778 & n3037 ;
  assign n3039 = ~n3020 & ~n3038 ;
  assign n3040 = ~n3036 & ~n3039 ;
  assign n3041 = n2952 & ~n3036 ;
  assign n3042 = n2914 & n3041 ;
  assign n3043 = ~n3040 & ~n3042 ;
  assign n3044 = ~\g1696_reg/NET0131  & \g7961_pad  ;
  assign n3045 = \g1088_reg/NET0131  & ~\g1698_reg/NET0131  ;
  assign n3046 = \g1092_reg/NET0131  & ~\g1697_reg/NET0131  ;
  assign n3047 = ~n3045 & ~n3046 ;
  assign n3048 = ~n3044 & n3047 ;
  assign n3049 = \g7961_pad  & n3048 ;
  assign n3050 = ~n3043 & n3049 ;
  assign n3051 = ~n3031 & n3050 ;
  assign n3052 = ~n3006 & ~n3012 ;
  assign n3053 = n3023 & n3025 ;
  assign n3054 = ~n3008 & n3020 ;
  assign n3055 = n2780 & n3054 ;
  assign n3056 = ~n3053 & n3055 ;
  assign n3057 = n3052 & n3056 ;
  assign n3058 = ~n2844 & ~n3057 ;
  assign n3059 = \g1088_reg/NET0131  & ~\g1783_reg/NET0131  ;
  assign n3060 = ~\g1784_reg/NET0131  & \g7961_pad  ;
  assign n3061 = \g1092_reg/NET0131  & ~\g1785_reg/NET0131  ;
  assign n3062 = ~n3060 & ~n3061 ;
  assign n3063 = ~n3059 & n3062 ;
  assign n3064 = ~n2945 & ~n3063 ;
  assign n3065 = n2937 & n3064 ;
  assign n3066 = n2914 & n3065 ;
  assign n3067 = ~n3036 & ~n3066 ;
  assign n3068 = ~n3058 & n3067 ;
  assign n3069 = n3020 & n3036 ;
  assign n3070 = n3048 & ~n3069 ;
  assign n3071 = ~n3066 & n3070 ;
  assign n3072 = \g7961_pad  & ~n3071 ;
  assign n3073 = ~n3068 & n3072 ;
  assign n3074 = ~\g1696_reg/NET0131  & ~\g7961_pad  ;
  assign n3075 = ~n3073 & ~n3074 ;
  assign n3076 = ~n3051 & n3075 ;
  assign n3077 = \g1092_reg/NET0131  & n3048 ;
  assign n3078 = ~n3043 & n3077 ;
  assign n3079 = ~n3031 & n3078 ;
  assign n3080 = \g1092_reg/NET0131  & ~n3071 ;
  assign n3081 = ~n3068 & n3080 ;
  assign n3082 = ~\g1092_reg/NET0131  & ~\g1697_reg/NET0131  ;
  assign n3083 = ~n3081 & ~n3082 ;
  assign n3084 = ~n3079 & n3083 ;
  assign n3085 = \g1088_reg/NET0131  & n3048 ;
  assign n3086 = ~n3043 & n3085 ;
  assign n3087 = ~n3031 & n3086 ;
  assign n3088 = \g1088_reg/NET0131  & ~n3071 ;
  assign n3089 = ~n3068 & n3088 ;
  assign n3090 = ~\g1088_reg/NET0131  & ~\g1698_reg/NET0131  ;
  assign n3091 = ~n3089 & ~n3090 ;
  assign n3092 = ~n3087 & n3091 ;
  assign n3093 = \g1234_reg/NET0131  & ~\g5657_pad  ;
  assign n3094 = ~\g1186_reg/NET0131  & ~n3093 ;
  assign n3095 = \g5657_pad  & n1752 ;
  assign n3096 = n3094 & ~n3095 ;
  assign n3097 = ~n1750 & ~n3096 ;
  assign n3098 = ~\g1245_reg/NET0131  & ~\g1249_pad  ;
  assign n3099 = \g1186_reg/NET0131  & n3098 ;
  assign n3100 = ~n3097 & n3099 ;
  assign n3101 = \g1018_reg/NET0131  & ~\g1425_reg/NET0131  ;
  assign n3102 = ~\g1424_reg/NET0131  & \g5657_pad  ;
  assign n3103 = \g1024_reg/NET0131  & ~\g1423_reg/NET0131  ;
  assign n3104 = ~n3102 & ~n3103 ;
  assign n3105 = ~n3101 & n3104 ;
  assign n3106 = \g1024_reg/NET0131  & ~\g1417_reg/NET0131  ;
  assign n3107 = ~\g1418_reg/NET0131  & \g5657_pad  ;
  assign n3108 = \g1018_reg/NET0131  & ~\g1419_reg/NET0131  ;
  assign n3109 = ~n3107 & ~n3108 ;
  assign n3110 = ~n3106 & n3109 ;
  assign n3111 = ~n3105 & ~n3110 ;
  assign n3112 = ~\g1391_reg/NET0131  & \g5657_pad  ;
  assign n3113 = \g1018_reg/NET0131  & ~\g1392_reg/NET0131  ;
  assign n3114 = \g1024_reg/NET0131  & ~\g1390_reg/NET0131  ;
  assign n3115 = ~n3113 & ~n3114 ;
  assign n3116 = ~n3112 & n3115 ;
  assign n3117 = ~\g1400_reg/NET0131  & \g5657_pad  ;
  assign n3118 = \g1018_reg/NET0131  & ~\g1401_reg/NET0131  ;
  assign n3119 = \g1024_reg/NET0131  & ~\g1399_reg/NET0131  ;
  assign n3120 = ~n3118 & ~n3119 ;
  assign n3121 = ~n3117 & n3120 ;
  assign n3122 = ~n3116 & n3121 ;
  assign n3123 = n3111 & n3122 ;
  assign n3124 = ~\g1409_reg/NET0131  & \g5657_pad  ;
  assign n3125 = \g1018_reg/NET0131  & ~\g1410_reg/NET0131  ;
  assign n3126 = \g1024_reg/NET0131  & ~\g1408_reg/NET0131  ;
  assign n3127 = ~n3125 & ~n3126 ;
  assign n3128 = ~n3124 & n3127 ;
  assign n3129 = ~\g1397_reg/NET0131  & \g5657_pad  ;
  assign n3130 = \g1024_reg/NET0131  & ~\g1396_reg/NET0131  ;
  assign n3131 = \g1018_reg/NET0131  & ~\g1398_reg/NET0131  ;
  assign n3132 = ~n3130 & ~n3131 ;
  assign n3133 = ~n3129 & n3132 ;
  assign n3134 = ~n3128 & n3133 ;
  assign n3135 = ~\g1385_reg/NET0131  & \g5657_pad  ;
  assign n3136 = \g1024_reg/NET0131  & ~\g1384_reg/NET0131  ;
  assign n3137 = \g1018_reg/NET0131  & ~\g1386_reg/NET0131  ;
  assign n3138 = ~n3136 & ~n3137 ;
  assign n3139 = ~n3135 & n3138 ;
  assign n3140 = ~\g1388_reg/NET0131  & \g5657_pad  ;
  assign n3141 = \g1018_reg/NET0131  & ~\g1389_reg/NET0131  ;
  assign n3142 = \g1024_reg/NET0131  & ~\g1387_reg/NET0131  ;
  assign n3143 = ~n3141 & ~n3142 ;
  assign n3144 = ~n3140 & n3143 ;
  assign n3145 = n3139 & ~n3144 ;
  assign n3146 = n3134 & n3145 ;
  assign n3147 = ~\g1403_reg/NET0131  & \g5657_pad  ;
  assign n3148 = \g1018_reg/NET0131  & ~\g1404_reg/NET0131  ;
  assign n3149 = \g1024_reg/NET0131  & ~\g1402_reg/NET0131  ;
  assign n3150 = ~n3148 & ~n3149 ;
  assign n3151 = ~n3147 & n3150 ;
  assign n3152 = ~\g1394_reg/NET0131  & \g5657_pad  ;
  assign n3153 = \g1018_reg/NET0131  & ~\g1395_reg/NET0131  ;
  assign n3154 = \g1024_reg/NET0131  & ~\g1393_reg/NET0131  ;
  assign n3155 = ~n3153 & ~n3154 ;
  assign n3156 = ~n3152 & n3155 ;
  assign n3157 = n3151 & ~n3156 ;
  assign n3158 = ~\g1412_reg/NET0131  & \g5657_pad  ;
  assign n3159 = \g1024_reg/NET0131  & ~\g1411_reg/NET0131  ;
  assign n3160 = \g1018_reg/NET0131  & ~\g1413_reg/NET0131  ;
  assign n3161 = ~n3159 & ~n3160 ;
  assign n3162 = ~n3158 & n3161 ;
  assign n3163 = ~\g1406_reg/NET0131  & \g5657_pad  ;
  assign n3164 = \g1018_reg/NET0131  & ~\g1407_reg/NET0131  ;
  assign n3165 = \g1024_reg/NET0131  & ~\g1405_reg/NET0131  ;
  assign n3166 = ~n3164 & ~n3165 ;
  assign n3167 = ~n3163 & n3166 ;
  assign n3168 = ~n3162 & n3167 ;
  assign n3169 = n3157 & n3168 ;
  assign n3170 = n3146 & n3169 ;
  assign n3171 = n3123 & n3170 ;
  assign n3172 = \g1300_reg/NET0131  & \g5657_pad  ;
  assign n3173 = \g1018_reg/NET0131  & \g1303_reg/NET0131  ;
  assign n3174 = \g1024_reg/NET0131  & \g1306_reg/NET0131  ;
  assign n3175 = ~n3173 & ~n3174 ;
  assign n3176 = ~n3172 & n3175 ;
  assign n3177 = ~n3116 & n3176 ;
  assign n3178 = ~n3171 & n3177 ;
  assign n3179 = n3116 & ~n3176 ;
  assign n3180 = n3123 & ~n3176 ;
  assign n3181 = n3170 & n3180 ;
  assign n3182 = ~n3179 & ~n3181 ;
  assign n3183 = ~n3178 & n3182 ;
  assign n3184 = \g1018_reg/NET0131  & \g1294_reg/NET0131  ;
  assign n3185 = \g1291_reg/NET0131  & \g5657_pad  ;
  assign n3186 = \g1024_reg/NET0131  & \g1297_reg/NET0131  ;
  assign n3187 = ~n3185 & ~n3186 ;
  assign n3188 = ~n3184 & n3187 ;
  assign n3189 = ~n3156 & n3188 ;
  assign n3190 = ~n3171 & n3189 ;
  assign n3191 = n3156 & ~n3188 ;
  assign n3192 = n3123 & ~n3188 ;
  assign n3193 = n3170 & n3192 ;
  assign n3194 = ~n3191 & ~n3193 ;
  assign n3195 = ~n3190 & n3194 ;
  assign n3196 = ~n3183 & n3195 ;
  assign n3197 = n3183 & ~n3195 ;
  assign n3198 = ~n3196 & ~n3197 ;
  assign n3199 = n3100 & ~n3198 ;
  assign n3200 = n3139 & n3176 ;
  assign n3201 = ~n3139 & ~n3176 ;
  assign n3202 = ~n3200 & ~n3201 ;
  assign n3203 = n3100 & ~n3202 ;
  assign n3204 = ~n3144 & n3188 ;
  assign n3205 = ~n3171 & n3204 ;
  assign n3206 = n3144 & ~n3188 ;
  assign n3207 = ~n3193 & ~n3206 ;
  assign n3208 = n3100 & n3207 ;
  assign n3209 = ~n3205 & n3208 ;
  assign n3210 = ~n3203 & ~n3209 ;
  assign n3211 = ~n3151 & ~n3176 ;
  assign n3212 = n3151 & n3176 ;
  assign n3213 = ~n3211 & ~n3212 ;
  assign n3214 = n3100 & ~n3213 ;
  assign n3215 = n3167 & n3188 ;
  assign n3216 = ~n3167 & ~n3188 ;
  assign n3217 = ~n3215 & ~n3216 ;
  assign n3218 = n3214 & n3217 ;
  assign n3219 = n3100 & ~n3217 ;
  assign n3220 = n3213 & n3219 ;
  assign n3221 = ~n3218 & ~n3220 ;
  assign n3222 = n3121 & n3188 ;
  assign n3223 = ~n3121 & ~n3188 ;
  assign n3224 = ~n3222 & ~n3223 ;
  assign n3225 = n3100 & ~n3224 ;
  assign n3226 = ~n3133 & ~n3176 ;
  assign n3227 = n3133 & n3176 ;
  assign n3228 = ~n3226 & ~n3227 ;
  assign n3229 = n3100 & ~n3228 ;
  assign n3230 = n3225 & ~n3229 ;
  assign n3231 = ~n3221 & n3230 ;
  assign n3232 = n3225 & n3229 ;
  assign n3233 = n3221 & n3232 ;
  assign n3234 = ~n3231 & ~n3233 ;
  assign n3235 = ~n3225 & ~n3229 ;
  assign n3236 = n3221 & n3235 ;
  assign n3237 = ~n3225 & n3229 ;
  assign n3238 = ~n3221 & n3237 ;
  assign n3239 = ~n3236 & ~n3238 ;
  assign n3240 = n3234 & n3239 ;
  assign n3241 = n3210 & ~n3240 ;
  assign n3242 = ~n3199 & n3241 ;
  assign n3243 = n3203 & n3209 ;
  assign n3244 = ~n3240 & n3243 ;
  assign n3245 = ~n3199 & n3244 ;
  assign n3246 = ~n3242 & ~n3245 ;
  assign n3247 = n3203 & ~n3209 ;
  assign n3248 = ~n3240 & n3247 ;
  assign n3249 = n3199 & n3248 ;
  assign n3250 = ~n3203 & n3209 ;
  assign n3251 = ~n3240 & n3250 ;
  assign n3252 = n3199 & n3251 ;
  assign n3253 = ~n3249 & ~n3252 ;
  assign n3254 = n3246 & n3253 ;
  assign n3255 = n3240 & n3247 ;
  assign n3256 = ~n3199 & n3255 ;
  assign n3257 = n3240 & n3250 ;
  assign n3258 = ~n3199 & n3257 ;
  assign n3259 = ~n3256 & ~n3258 ;
  assign n3260 = n3210 & n3240 ;
  assign n3261 = n3199 & n3260 ;
  assign n3262 = n3240 & n3243 ;
  assign n3263 = n3199 & n3262 ;
  assign n3264 = ~n3261 & ~n3263 ;
  assign n3265 = n3259 & n3264 ;
  assign n3266 = n3254 & n3265 ;
  assign n3267 = \g1196_reg/NET0131  & n3266 ;
  assign n3268 = ~n3162 & n3188 ;
  assign n3269 = ~n3171 & n3268 ;
  assign n3270 = n3162 & ~n3188 ;
  assign n3271 = ~n3193 & ~n3270 ;
  assign n3272 = ~n3269 & n3271 ;
  assign n3273 = ~n3128 & n3176 ;
  assign n3274 = ~n3171 & n3273 ;
  assign n3275 = n3128 & ~n3176 ;
  assign n3276 = ~n3181 & ~n3275 ;
  assign n3277 = ~n3274 & n3276 ;
  assign n3278 = ~n3272 & n3277 ;
  assign n3279 = n3272 & ~n3277 ;
  assign n3280 = ~n3278 & ~n3279 ;
  assign n3281 = \g1243_reg/NET0131  & n3100 ;
  assign n3282 = ~n3280 & n3281 ;
  assign n3283 = \g1211_reg/NET0131  & n1768 ;
  assign n3284 = ~\g1224_reg/NET0131  & \g3229_pad  ;
  assign n3285 = n3283 & ~n3284 ;
  assign n3286 = ~\g1227_reg/NET0131  & ~\g3229_pad  ;
  assign n3287 = n3098 & ~n3286 ;
  assign n3288 = n3285 & n3287 ;
  assign n3289 = ~n3097 & n3288 ;
  assign n3290 = ~n3282 & ~n3289 ;
  assign n3291 = ~n3267 & n3290 ;
  assign n3292 = n1816 & ~n1995 ;
  assign n3293 = ~n1934 & n3292 ;
  assign n3294 = ~\g1196_reg/NET0131  & ~\g1905_reg/NET0131  ;
  assign n3295 = ~\g1243_reg/NET0131  & ~n3294 ;
  assign n3296 = ~\g1243_reg/NET0131  & ~\g1905_reg/NET0131  ;
  assign n3297 = ~\g1196_reg/NET0131  & ~\g1910_reg/NET0131  ;
  assign n3298 = ~n3296 & n3297 ;
  assign n3299 = n1998 & n3298 ;
  assign n3300 = n3295 & ~n3299 ;
  assign n3301 = n1757 & n3295 ;
  assign n3302 = n1755 & n3301 ;
  assign n3303 = ~n3300 & ~n3302 ;
  assign n3304 = ~n3293 & ~n3303 ;
  assign n3305 = ~n2005 & ~n3304 ;
  assign n3306 = ~\g2115_reg/NET0131  & \g5657_pad  ;
  assign n3307 = \g1018_reg/NET0131  & ~\g2116_reg/NET0131  ;
  assign n3308 = \g1024_reg/NET0131  & ~\g2114_reg/NET0131  ;
  assign n3309 = ~n3307 & ~n3308 ;
  assign n3310 = ~n3306 & n3309 ;
  assign n3311 = \g1880_reg/NET0131  & ~n3310 ;
  assign n3312 = \g1880_reg/NET0131  & n1839 ;
  assign n3313 = n1886 & n3312 ;
  assign n3314 = ~n3311 & ~n3313 ;
  assign n3315 = ~n1994 & n1998 ;
  assign n3316 = ~n3304 & n3315 ;
  assign n3317 = n3314 & n3316 ;
  assign n3318 = ~n3305 & ~n3317 ;
  assign n3319 = ~n1951 & n3292 ;
  assign n3320 = ~\g1196_reg/NET0131  & ~\g1909_reg/NET0131  ;
  assign n3321 = ~n3296 & n3320 ;
  assign n3322 = n1998 & n3321 ;
  assign n3323 = ~n1994 & n3322 ;
  assign n3324 = n3295 & ~n3323 ;
  assign n3325 = ~n3319 & n3324 ;
  assign n3326 = ~n2005 & ~n3325 ;
  assign n3327 = n3315 & ~n3325 ;
  assign n3328 = ~n3314 & n3327 ;
  assign n3329 = ~n3326 & ~n3328 ;
  assign n3330 = ~n1945 & n3292 ;
  assign n3331 = ~\g1196_reg/NET0131  & ~\g1911_reg/NET0131  ;
  assign n3332 = ~n3296 & n3331 ;
  assign n3333 = n1998 & n3332 ;
  assign n3334 = ~n1994 & n3333 ;
  assign n3335 = n3295 & ~n3334 ;
  assign n3336 = ~n3330 & n3335 ;
  assign n3337 = ~n2005 & ~n3336 ;
  assign n3338 = n3315 & ~n3336 ;
  assign n3339 = n3314 & n3338 ;
  assign n3340 = ~n3337 & ~n3339 ;
  assign n3341 = ~n1942 & n3292 ;
  assign n3342 = ~\g1196_reg/NET0131  & ~\g1912_reg/NET0131  ;
  assign n3343 = ~n3296 & n3342 ;
  assign n3344 = n1998 & n3343 ;
  assign n3345 = ~n1994 & n3344 ;
  assign n3346 = n3295 & ~n3345 ;
  assign n3347 = ~n3341 & n3346 ;
  assign n3348 = ~n2005 & ~n3347 ;
  assign n3349 = n3315 & ~n3347 ;
  assign n3350 = ~n3314 & n3349 ;
  assign n3351 = ~n3348 & ~n3350 ;
  assign n3352 = ~n1998 & n2005 ;
  assign n3353 = n1757 & n2005 ;
  assign n3354 = n1755 & n3353 ;
  assign n3355 = ~n3352 & ~n3354 ;
  assign n3356 = ~\g1196_reg/NET0131  & ~n3296 ;
  assign n3357 = n1816 & ~n3356 ;
  assign n3358 = n1899 & n3357 ;
  assign n3359 = ~\g1196_reg/NET0131  & ~\g1913_reg/NET0131  ;
  assign n3360 = ~n3296 & n3359 ;
  assign n3361 = n1998 & n3360 ;
  assign n3362 = ~n1994 & n3361 ;
  assign n3363 = n3295 & ~n3362 ;
  assign n3364 = ~n3358 & n3363 ;
  assign n3365 = n3355 & ~n3364 ;
  assign n3366 = n1912 & n3357 ;
  assign n3367 = ~\g1196_reg/NET0131  & ~\g1914_reg/NET0131  ;
  assign n3368 = ~n3296 & n3367 ;
  assign n3369 = n1998 & n3368 ;
  assign n3370 = ~n1994 & n3369 ;
  assign n3371 = n3295 & ~n3370 ;
  assign n3372 = ~n3366 & n3371 ;
  assign n3373 = n3355 & ~n3372 ;
  assign n3374 = \g1563_reg/NET0131  & ~n2244 ;
  assign n3375 = n2247 & n3374 ;
  assign n3376 = ~n2151 & n3375 ;
  assign n3377 = n2146 & ~n2269 ;
  assign n3378 = ~n2274 & n3377 ;
  assign n3379 = n2264 & n3378 ;
  assign n3380 = n2230 & n3379 ;
  assign n3381 = ~n2151 & n2181 ;
  assign n3382 = n3380 & n3381 ;
  assign n3383 = ~n3376 & ~n3382 ;
  assign n3384 = ~n2146 & ~n2361 ;
  assign n3385 = n2415 & n3384 ;
  assign n3386 = ~n2284 & ~n2302 ;
  assign n3387 = ~n2312 & ~n2332 ;
  assign n3388 = n3386 & n3387 ;
  assign n3389 = n3385 & n3388 ;
  assign n3390 = n2323 & n2349 ;
  assign n3391 = n2342 & n2368 ;
  assign n3392 = n2294 & n3391 ;
  assign n3393 = n3390 & n3392 ;
  assign n3394 = n3389 & n3393 ;
  assign n3395 = ~n2428 & ~n3394 ;
  assign n3396 = n3383 & n3395 ;
  assign n3397 = ~\g105_reg/NET0131  & ~n3396 ;
  assign n3398 = n2398 & ~n2404 ;
  assign n3399 = n2389 & n3398 ;
  assign n3400 = n2249 & ~n3399 ;
  assign n3401 = ~n2151 & n2269 ;
  assign n3402 = n2146 & ~n2274 ;
  assign n3403 = n3401 & n3402 ;
  assign n3404 = n2264 & n3403 ;
  assign n3405 = n2230 & n3404 ;
  assign n3406 = n2181 & n3405 ;
  assign n3407 = ~\g105_reg/NET0131  & n3406 ;
  assign n3408 = ~n3400 & n3407 ;
  assign n3409 = ~n3397 & ~n3408 ;
  assign n3410 = ~n3400 & n3406 ;
  assign n3411 = ~n2428 & n3383 ;
  assign n3412 = n2284 & n2302 ;
  assign n3413 = n2146 & n2312 ;
  assign n3414 = n2332 & n2361 ;
  assign n3415 = n3413 & n3414 ;
  assign n3416 = n3412 & n3415 ;
  assign n3417 = n3393 & n3416 ;
  assign n3418 = ~n3394 & ~n3417 ;
  assign n3419 = ~n2146 & n2415 ;
  assign n3420 = ~n3418 & n3419 ;
  assign n3421 = n2146 & ~n2342 ;
  assign n3422 = ~n2146 & n2342 ;
  assign n3423 = n2415 & ~n3422 ;
  assign n3424 = ~n3421 & n3423 ;
  assign n3425 = ~n2146 & ~n2312 ;
  assign n3426 = ~n3413 & ~n3425 ;
  assign n3427 = n2361 & ~n3426 ;
  assign n3428 = n3424 & n3427 ;
  assign n3429 = ~n3420 & n3428 ;
  assign n3430 = n2415 & ~n3418 ;
  assign n3431 = n3424 & ~n3426 ;
  assign n3432 = ~n2361 & ~n3431 ;
  assign n3433 = ~n3430 & ~n3432 ;
  assign n3434 = ~n3420 & ~n3433 ;
  assign n3435 = ~n3429 & ~n3434 ;
  assign n3436 = n3411 & n3435 ;
  assign n3437 = ~n3410 & n3436 ;
  assign n3438 = n3409 & ~n3437 ;
  assign n3439 = \g7961_pad  & ~n3438 ;
  assign n3440 = ~\g195_reg/NET0131  & ~\g7961_pad  ;
  assign n3441 = ~n3439 & ~n3440 ;
  assign n3442 = \g1092_reg/NET0131  & ~n3438 ;
  assign n3443 = ~\g1092_reg/NET0131  & ~\g198_reg/NET0131  ;
  assign n3444 = ~n3442 & ~n3443 ;
  assign n3445 = \g1088_reg/NET0131  & ~n3438 ;
  assign n3446 = ~\g1088_reg/NET0131  & ~\g201_reg/NET0131  ;
  assign n3447 = ~n3445 & ~n3446 ;
  assign n3448 = n2453 & ~n2470 ;
  assign n3449 = n2458 & ~n2575 ;
  assign n3450 = n3448 & n3449 ;
  assign n3451 = n2591 & n3450 ;
  assign n3452 = n2547 & n3451 ;
  assign n3453 = ~n2725 & n3452 ;
  assign n3454 = ~n2720 & n3453 ;
  assign n3455 = ~n2662 & n3454 ;
  assign n3456 = n2453 & ~n2458 ;
  assign n3457 = ~n2464 & ~n3456 ;
  assign n3458 = ~n2470 & ~n3457 ;
  assign n3459 = n2464 & n3458 ;
  assign n3460 = n2586 & n3458 ;
  assign n3461 = n2547 & n3460 ;
  assign n3462 = ~n3459 & ~n3461 ;
  assign n3463 = ~n2598 & n3462 ;
  assign n3464 = ~n2453 & n2599 ;
  assign n3465 = n2635 & n2711 ;
  assign n3466 = n2607 & n2699 ;
  assign n3467 = n2648 & n3466 ;
  assign n3468 = n3465 & n3467 ;
  assign n3469 = n2670 & n2679 ;
  assign n3470 = n2616 & n3469 ;
  assign n3471 = n2453 & n2688 ;
  assign n3472 = n2624 & n3471 ;
  assign n3473 = n3470 & n3472 ;
  assign n3474 = n3468 & n3473 ;
  assign n3475 = ~n2453 & ~n2624 ;
  assign n3476 = n2599 & n3475 ;
  assign n3477 = ~n2670 & ~n2679 ;
  assign n3478 = ~n2616 & ~n2688 ;
  assign n3479 = n3477 & n3478 ;
  assign n3480 = n3476 & n3479 ;
  assign n3481 = n3468 & n3480 ;
  assign n3482 = ~n3474 & ~n3481 ;
  assign n3483 = n3464 & ~n3482 ;
  assign n3484 = n2599 & ~n3482 ;
  assign n3485 = n2453 & ~n2648 ;
  assign n3486 = n2599 & ~n3485 ;
  assign n3487 = ~n2648 & ~n2688 ;
  assign n3488 = ~n3471 & ~n3487 ;
  assign n3489 = n3486 & ~n3488 ;
  assign n3490 = ~n2624 & ~n3489 ;
  assign n3491 = n2624 & n3489 ;
  assign n3492 = ~n3490 & ~n3491 ;
  assign n3493 = ~n3484 & n3492 ;
  assign n3494 = ~n3483 & ~n3493 ;
  assign n3495 = n3463 & ~n3494 ;
  assign n3496 = ~n3455 & n3495 ;
  assign n3497 = \g7961_pad  & n3496 ;
  assign n3498 = ~n3455 & n3463 ;
  assign n3499 = ~\g793_reg/NET0131  & \g7961_pad  ;
  assign n3500 = ~n3498 & n3499 ;
  assign n3501 = ~n3497 & ~n3500 ;
  assign n3502 = ~\g7961_pad  & ~\g882_reg/NET0131  ;
  assign n3503 = n3501 & ~n3502 ;
  assign n3504 = \g1092_reg/NET0131  & n3496 ;
  assign n3505 = \g1092_reg/NET0131  & ~\g793_reg/NET0131  ;
  assign n3506 = ~n3498 & n3505 ;
  assign n3507 = ~n3504 & ~n3506 ;
  assign n3508 = ~\g1092_reg/NET0131  & ~\g885_reg/NET0131  ;
  assign n3509 = n3507 & ~n3508 ;
  assign n3510 = \g1088_reg/NET0131  & n3496 ;
  assign n3511 = \g1088_reg/NET0131  & ~\g793_reg/NET0131  ;
  assign n3512 = ~n3498 & n3511 ;
  assign n3513 = ~n3510 & ~n3512 ;
  assign n3514 = ~\g1088_reg/NET0131  & ~\g888_reg/NET0131  ;
  assign n3515 = n3513 & ~n3514 ;
  assign n3516 = ~n2453 & n2648 ;
  assign n3517 = n2599 & n3516 ;
  assign n3518 = n3486 & ~n3517 ;
  assign n3519 = ~n2688 & ~n3518 ;
  assign n3520 = n2688 & ~n3485 ;
  assign n3521 = n2599 & ~n3516 ;
  assign n3522 = n3520 & n3521 ;
  assign n3523 = ~n3519 & ~n3522 ;
  assign n3524 = ~n3484 & n3523 ;
  assign n3525 = ~n3483 & ~n3524 ;
  assign n3526 = n3463 & ~n3525 ;
  assign n3527 = ~n3455 & n3526 ;
  assign n3528 = \g7961_pad  & n3527 ;
  assign n3529 = ~\g789_reg/NET0131  & \g7961_pad  ;
  assign n3530 = ~n3498 & n3529 ;
  assign n3531 = ~n3528 & ~n3530 ;
  assign n3532 = ~\g7961_pad  & ~\g918_reg/NET0131  ;
  assign n3533 = n3531 & ~n3532 ;
  assign n3534 = \g1092_reg/NET0131  & n3527 ;
  assign n3535 = \g1092_reg/NET0131  & ~\g789_reg/NET0131  ;
  assign n3536 = ~n3498 & n3535 ;
  assign n3537 = ~n3534 & ~n3536 ;
  assign n3538 = ~\g1092_reg/NET0131  & ~\g921_reg/NET0131  ;
  assign n3539 = n3537 & ~n3538 ;
  assign n3540 = \g1088_reg/NET0131  & n3527 ;
  assign n3541 = \g1088_reg/NET0131  & ~\g789_reg/NET0131  ;
  assign n3542 = ~n3498 & n3541 ;
  assign n3543 = ~n3540 & ~n3542 ;
  assign n3544 = ~\g1088_reg/NET0131  & ~\g924_reg/NET0131  ;
  assign n3545 = n3543 & ~n3544 ;
  assign n3546 = ~n2670 & ~n3489 ;
  assign n3547 = n2624 & ~n3464 ;
  assign n3548 = ~n2670 & ~n3476 ;
  assign n3549 = ~n3547 & n3548 ;
  assign n3550 = ~n3546 & ~n3549 ;
  assign n3551 = ~n3476 & ~n3547 ;
  assign n3552 = n2670 & n3489 ;
  assign n3553 = ~n3551 & n3552 ;
  assign n3554 = n3550 & ~n3553 ;
  assign n3555 = ~n3484 & n3554 ;
  assign n3556 = ~n3483 & ~n3555 ;
  assign n3557 = n3463 & ~n3556 ;
  assign n3558 = ~n3455 & n3557 ;
  assign n3559 = \g7961_pad  & n3558 ;
  assign n3560 = \g7961_pad  & ~\g797_reg/NET0131  ;
  assign n3561 = ~n3498 & n3560 ;
  assign n3562 = ~n3559 & ~n3561 ;
  assign n3563 = ~\g7961_pad  & ~\g927_reg/NET0131  ;
  assign n3564 = n3562 & ~n3563 ;
  assign n3565 = \g1088_reg/NET0131  & n3558 ;
  assign n3566 = \g1088_reg/NET0131  & ~\g797_reg/NET0131  ;
  assign n3567 = ~n3498 & n3566 ;
  assign n3568 = ~n3565 & ~n3567 ;
  assign n3569 = ~\g1088_reg/NET0131  & ~\g933_reg/NET0131  ;
  assign n3570 = n3568 & ~n3569 ;
  assign n3571 = \g1092_reg/NET0131  & n3558 ;
  assign n3572 = \g1092_reg/NET0131  & ~\g797_reg/NET0131  ;
  assign n3573 = ~n3498 & n3572 ;
  assign n3574 = ~n3571 & ~n3573 ;
  assign n3575 = ~\g1092_reg/NET0131  & ~\g930_reg/NET0131  ;
  assign n3576 = n3574 & ~n3575 ;
  assign n3577 = ~\g7961_pad  & \g954_reg/NET0131  ;
  assign n3578 = n3463 & n3483 ;
  assign n3579 = ~n3455 & n3578 ;
  assign n3580 = n2515 & ~n3498 ;
  assign n3581 = ~n3579 & ~n3580 ;
  assign n3582 = ~\g7961_pad  & ~\g954_reg/NET0131  ;
  assign n3583 = ~n2598 & ~n3484 ;
  assign n3584 = n3462 & n3583 ;
  assign n3585 = n3489 & ~n3551 ;
  assign n3586 = ~n2670 & ~n3464 ;
  assign n3587 = ~n2453 & n2670 ;
  assign n3588 = n2599 & n3587 ;
  assign n3589 = ~n3586 & ~n3588 ;
  assign n3590 = ~n2607 & ~n3464 ;
  assign n3591 = ~n2453 & n2607 ;
  assign n3592 = n2599 & n3591 ;
  assign n3593 = ~n3590 & ~n3592 ;
  assign n3594 = n3589 & n3593 ;
  assign n3595 = n3585 & n3594 ;
  assign n3596 = ~n2453 & ~n2635 ;
  assign n3597 = n2599 & n3596 ;
  assign n3598 = ~n3465 & ~n3597 ;
  assign n3599 = ~n2607 & n2711 ;
  assign n3600 = ~n3598 & ~n3599 ;
  assign n3601 = ~n2699 & ~n3464 ;
  assign n3602 = ~n2453 & n2699 ;
  assign n3603 = n2599 & n3602 ;
  assign n3604 = ~n3601 & ~n3603 ;
  assign n3605 = n3600 & n3604 ;
  assign n3606 = ~n2616 & ~n3464 ;
  assign n3607 = ~n2453 & n2616 ;
  assign n3608 = n2599 & n3607 ;
  assign n3609 = ~n3606 & ~n3608 ;
  assign n3610 = n3605 & n3609 ;
  assign n3611 = n3595 & n3610 ;
  assign n3612 = ~n2679 & n3611 ;
  assign n3613 = n2679 & ~n3611 ;
  assign n3614 = ~n3612 & ~n3613 ;
  assign n3615 = ~n3455 & ~n3614 ;
  assign n3616 = n3584 & n3615 ;
  assign n3617 = ~n3582 & ~n3616 ;
  assign n3618 = n3581 & n3617 ;
  assign n3619 = ~n3577 & ~n3618 ;
  assign n3620 = ~\g1092_reg/NET0131  & \g957_reg/NET0131  ;
  assign n3621 = ~\g1092_reg/NET0131  & ~\g957_reg/NET0131  ;
  assign n3622 = ~n3616 & ~n3621 ;
  assign n3623 = n3581 & n3622 ;
  assign n3624 = ~n3620 & ~n3623 ;
  assign n3625 = ~\g1088_reg/NET0131  & \g960_reg/NET0131  ;
  assign n3626 = ~\g1088_reg/NET0131  & ~\g960_reg/NET0131  ;
  assign n3627 = ~n3616 & ~n3626 ;
  assign n3628 = n3581 & n3627 ;
  assign n3629 = ~n3625 & ~n3628 ;
  assign n3630 = ~n2844 & ~n3015 ;
  assign n3631 = ~n2950 & n3048 ;
  assign n3632 = n2937 & ~n2945 ;
  assign n3633 = n3020 & ~n3036 ;
  assign n3634 = n3632 & n3633 ;
  assign n3635 = n2914 & n3634 ;
  assign n3636 = n3631 & n3635 ;
  assign n3637 = n3630 & n3636 ;
  assign n3638 = ~n3020 & n3048 ;
  assign n3639 = ~n3038 & ~n3638 ;
  assign n3640 = ~n3036 & ~n3639 ;
  assign n3641 = n3038 & n3640 ;
  assign n3642 = n2952 & n3640 ;
  assign n3643 = n2914 & n3642 ;
  assign n3644 = ~n3641 & ~n3643 ;
  assign n3645 = ~n3066 & n3644 ;
  assign n3646 = ~n3048 & n3069 ;
  assign n3647 = n2798 & n2962 ;
  assign n3648 = n2819 & n2978 ;
  assign n3649 = n2807 & n3648 ;
  assign n3650 = n3647 & n3649 ;
  assign n3651 = n2969 & n3048 ;
  assign n3652 = n2826 & n2991 ;
  assign n3653 = n2790 & n3000 ;
  assign n3654 = n3652 & n3653 ;
  assign n3655 = n3651 & n3654 ;
  assign n3656 = n3650 & n3655 ;
  assign n3657 = ~n2790 & ~n3048 ;
  assign n3658 = n3069 & n3657 ;
  assign n3659 = ~n2826 & ~n2991 ;
  assign n3660 = ~n2969 & ~n3000 ;
  assign n3661 = n3659 & n3660 ;
  assign n3662 = n3658 & n3661 ;
  assign n3663 = n3650 & n3662 ;
  assign n3664 = ~n3656 & ~n3663 ;
  assign n3665 = n3646 & ~n3664 ;
  assign n3666 = n3069 & ~n3664 ;
  assign n3667 = ~n2819 & n3048 ;
  assign n3668 = n3069 & ~n3667 ;
  assign n3669 = ~n2819 & ~n2969 ;
  assign n3670 = ~n3651 & ~n3669 ;
  assign n3671 = n3668 & ~n3670 ;
  assign n3672 = ~n2826 & n3671 ;
  assign n3673 = n2826 & ~n3671 ;
  assign n3674 = ~n3672 & ~n3673 ;
  assign n3675 = ~n3666 & ~n3674 ;
  assign n3676 = ~n3665 & ~n3675 ;
  assign n3677 = n3645 & ~n3676 ;
  assign n3678 = ~n3637 & n3677 ;
  assign n3679 = \g7961_pad  & n3678 ;
  assign n3680 = ~n3637 & n3645 ;
  assign n3681 = ~\g1481_reg/NET0131  & \g7961_pad  ;
  assign n3682 = ~n3680 & n3681 ;
  assign n3683 = ~n3679 & ~n3682 ;
  assign n3684 = ~\g1576_reg/NET0131  & ~\g7961_pad  ;
  assign n3685 = n3683 & ~n3684 ;
  assign n3686 = n1249 & n1464 ;
  assign n3687 = n1370 & ~n3686 ;
  assign n3688 = ~n1425 & n1444 ;
  assign n3689 = n1412 & n1420 ;
  assign n3690 = n1186 & ~n1437 ;
  assign n3691 = n3689 & n3690 ;
  assign n3692 = n1382 & n3691 ;
  assign n3693 = n3688 & n3692 ;
  assign n3694 = ~n3687 & n3693 ;
  assign n3695 = ~n1186 & n1444 ;
  assign n3696 = ~n1425 & ~n1437 ;
  assign n3697 = n3695 & n3696 ;
  assign n3698 = n3689 & n3697 ;
  assign n3699 = n1382 & n3698 ;
  assign n3700 = \g1563_reg/NET0131  & ~n1308 ;
  assign n3701 = n1311 & n3700 ;
  assign n3702 = ~n1437 & n3701 ;
  assign n3703 = ~n1454 & ~n3702 ;
  assign n3704 = ~n3699 & n3703 ;
  assign n3705 = ~n1444 & n1445 ;
  assign n3706 = n1191 & n1265 ;
  assign n3707 = n1212 & n1254 ;
  assign n3708 = n1290 & n3707 ;
  assign n3709 = n3706 & n3708 ;
  assign n3710 = n1224 & n1234 ;
  assign n3711 = n1279 & n3710 ;
  assign n3712 = n1200 & n1444 ;
  assign n3713 = n1297 & n3712 ;
  assign n3714 = n3711 & n3713 ;
  assign n3715 = n3709 & n3714 ;
  assign n3716 = ~n1279 & ~n1444 ;
  assign n3717 = n1445 & n3716 ;
  assign n3718 = ~n1224 & ~n1234 ;
  assign n3719 = ~n1200 & ~n1297 ;
  assign n3720 = n3718 & n3719 ;
  assign n3721 = n3717 & n3720 ;
  assign n3722 = n3709 & n3721 ;
  assign n3723 = ~n3715 & ~n3722 ;
  assign n3724 = n3705 & ~n3723 ;
  assign n3725 = n1445 & ~n3723 ;
  assign n3726 = ~n1290 & n1444 ;
  assign n3727 = n1445 & ~n3726 ;
  assign n3728 = ~n1200 & ~n1290 ;
  assign n3729 = ~n3712 & ~n3728 ;
  assign n3730 = n3727 & ~n3729 ;
  assign n3731 = ~n1297 & n3730 ;
  assign n3732 = n1297 & ~n3730 ;
  assign n3733 = ~n3731 & ~n3732 ;
  assign n3734 = ~n3725 & ~n3733 ;
  assign n3735 = ~n3724 & ~n3734 ;
  assign n3736 = n3704 & ~n3735 ;
  assign n3737 = ~n3694 & n3736 ;
  assign n3738 = \g7961_pad  & n3737 ;
  assign n3739 = ~n3694 & n3704 ;
  assign n3740 = ~\g2175_reg/NET0131  & \g7961_pad  ;
  assign n3741 = ~n3739 & n3740 ;
  assign n3742 = ~n3738 & ~n3741 ;
  assign n3743 = ~\g2270_reg/NET0131  & ~\g7961_pad  ;
  assign n3744 = n3742 & ~n3743 ;
  assign n3745 = \g1088_reg/NET0131  & n3737 ;
  assign n3746 = \g1088_reg/NET0131  & ~\g2175_reg/NET0131  ;
  assign n3747 = ~n3739 & n3746 ;
  assign n3748 = ~n3745 & ~n3747 ;
  assign n3749 = ~\g1088_reg/NET0131  & ~\g2276_reg/NET0131  ;
  assign n3750 = n3748 & ~n3749 ;
  assign n3751 = \g1092_reg/NET0131  & n3737 ;
  assign n3752 = \g1092_reg/NET0131  & ~\g2175_reg/NET0131  ;
  assign n3753 = ~n3739 & n3752 ;
  assign n3754 = ~n3751 & ~n3753 ;
  assign n3755 = ~\g1092_reg/NET0131  & ~\g2273_reg/NET0131  ;
  assign n3756 = n3754 & ~n3755 ;
  assign n3757 = \g1092_reg/NET0131  & n3678 ;
  assign n3758 = \g1092_reg/NET0131  & ~\g1481_reg/NET0131  ;
  assign n3759 = ~n3680 & n3758 ;
  assign n3760 = ~n3757 & ~n3759 ;
  assign n3761 = ~\g1092_reg/NET0131  & ~\g1579_reg/NET0131  ;
  assign n3762 = n3760 & ~n3761 ;
  assign n3763 = ~n1290 & ~n1444 ;
  assign n3764 = n1445 & n3763 ;
  assign n3765 = n1290 & n1444 ;
  assign n3766 = n1445 & n3765 ;
  assign n3767 = ~n3764 & ~n3766 ;
  assign n3768 = n1200 & n3767 ;
  assign n3769 = ~n1200 & ~n3767 ;
  assign n3770 = ~n3768 & ~n3769 ;
  assign n3771 = ~n3725 & ~n3770 ;
  assign n3772 = ~n3724 & ~n3771 ;
  assign n3773 = n3704 & ~n3772 ;
  assign n3774 = ~n3694 & n3773 ;
  assign n3775 = \g7961_pad  & n3774 ;
  assign n3776 = ~\g2170_reg/NET0131  & \g7961_pad  ;
  assign n3777 = ~n3739 & n3776 ;
  assign n3778 = ~n3775 & ~n3777 ;
  assign n3779 = ~\g2306_reg/NET0131  & ~\g7961_pad  ;
  assign n3780 = n3778 & ~n3779 ;
  assign n3781 = \g1088_reg/NET0131  & n3678 ;
  assign n3782 = \g1088_reg/NET0131  & ~\g1481_reg/NET0131  ;
  assign n3783 = ~n3680 & n3782 ;
  assign n3784 = ~n3781 & ~n3783 ;
  assign n3785 = ~\g1088_reg/NET0131  & ~\g1582_reg/NET0131  ;
  assign n3786 = n3784 & ~n3785 ;
  assign n3787 = \g1092_reg/NET0131  & n3774 ;
  assign n3788 = \g1092_reg/NET0131  & ~\g2170_reg/NET0131  ;
  assign n3789 = ~n3739 & n3788 ;
  assign n3790 = ~n3787 & ~n3789 ;
  assign n3791 = ~\g1092_reg/NET0131  & ~\g2309_reg/NET0131  ;
  assign n3792 = n3790 & ~n3791 ;
  assign n3793 = \g1088_reg/NET0131  & n3774 ;
  assign n3794 = \g1088_reg/NET0131  & ~\g2170_reg/NET0131  ;
  assign n3795 = ~n3739 & n3794 ;
  assign n3796 = ~n3793 & ~n3795 ;
  assign n3797 = ~\g1088_reg/NET0131  & ~\g2312_reg/NET0131  ;
  assign n3798 = n3796 & ~n3797 ;
  assign n3799 = ~n1234 & ~n3730 ;
  assign n3800 = ~n1234 & n1297 ;
  assign n3801 = n3705 & n3800 ;
  assign n3802 = ~n1234 & ~n1297 ;
  assign n3803 = ~n3705 & n3802 ;
  assign n3804 = ~n3801 & ~n3803 ;
  assign n3805 = ~n3799 & n3804 ;
  assign n3806 = ~n1297 & ~n3705 ;
  assign n3807 = n3730 & ~n3806 ;
  assign n3808 = n1297 & ~n1444 ;
  assign n3809 = n1445 & n3808 ;
  assign n3810 = n1234 & ~n3809 ;
  assign n3811 = n3807 & n3810 ;
  assign n3812 = n3805 & ~n3811 ;
  assign n3813 = ~n3725 & n3812 ;
  assign n3814 = ~n3724 & ~n3813 ;
  assign n3815 = n3704 & ~n3814 ;
  assign n3816 = ~n3694 & n3815 ;
  assign n3817 = \g7961_pad  & n3816 ;
  assign n3818 = ~\g2180_reg/NET0131  & \g7961_pad  ;
  assign n3819 = ~n3739 & n3818 ;
  assign n3820 = ~n3817 & ~n3819 ;
  assign n3821 = ~\g2315_reg/NET0131  & ~\g7961_pad  ;
  assign n3822 = n3820 & ~n3821 ;
  assign n3823 = \g1092_reg/NET0131  & n3816 ;
  assign n3824 = \g1092_reg/NET0131  & ~\g2180_reg/NET0131  ;
  assign n3825 = ~n3739 & n3824 ;
  assign n3826 = ~n3823 & ~n3825 ;
  assign n3827 = ~\g1092_reg/NET0131  & ~\g2318_reg/NET0131  ;
  assign n3828 = n3826 & ~n3827 ;
  assign n3829 = ~\g101_reg/NET0131  & ~n3396 ;
  assign n3830 = ~\g101_reg/NET0131  & n3406 ;
  assign n3831 = ~n3400 & n3830 ;
  assign n3832 = ~n3829 & ~n3831 ;
  assign n3833 = n2312 & ~n3421 ;
  assign n3834 = n3423 & n3833 ;
  assign n3835 = ~n3420 & n3834 ;
  assign n3836 = ~n2312 & ~n3424 ;
  assign n3837 = ~n3430 & ~n3836 ;
  assign n3838 = ~n3420 & ~n3837 ;
  assign n3839 = ~n3835 & ~n3838 ;
  assign n3840 = n3411 & n3839 ;
  assign n3841 = ~n3410 & n3840 ;
  assign n3842 = n3832 & ~n3841 ;
  assign n3843 = \g7961_pad  & ~n3842 ;
  assign n3844 = ~\g231_reg/NET0131  & ~\g7961_pad  ;
  assign n3845 = ~n3843 & ~n3844 ;
  assign n3846 = \g1088_reg/NET0131  & n3816 ;
  assign n3847 = \g1088_reg/NET0131  & ~\g2180_reg/NET0131  ;
  assign n3848 = ~n3739 & n3847 ;
  assign n3849 = ~n3846 & ~n3848 ;
  assign n3850 = ~\g1088_reg/NET0131  & ~\g2321_reg/NET0131  ;
  assign n3851 = n3849 & ~n3850 ;
  assign n3852 = \g2342_reg/NET0131  & ~\g7961_pad  ;
  assign n3853 = n3704 & n3724 ;
  assign n3854 = ~n3694 & n3853 ;
  assign n3855 = n1219 & ~n3739 ;
  assign n3856 = ~n3854 & ~n3855 ;
  assign n3857 = ~\g2342_reg/NET0131  & ~\g7961_pad  ;
  assign n3858 = ~n3699 & ~n3725 ;
  assign n3859 = n3703 & n3858 ;
  assign n3860 = ~n1234 & ~n1444 ;
  assign n3861 = n1445 & n3860 ;
  assign n3862 = ~n1254 & ~n3861 ;
  assign n3863 = ~n1234 & n1254 ;
  assign n3864 = n1254 & ~n1444 ;
  assign n3865 = n1445 & n3864 ;
  assign n3866 = ~n3863 & ~n3865 ;
  assign n3867 = ~n3862 & n3866 ;
  assign n3868 = ~n1212 & ~n3705 ;
  assign n3869 = n1212 & ~n1444 ;
  assign n3870 = n1445 & n3869 ;
  assign n3871 = ~n3809 & ~n3870 ;
  assign n3872 = ~n3868 & n3871 ;
  assign n3873 = n3867 & n3872 ;
  assign n3874 = ~n1265 & ~n3705 ;
  assign n3875 = ~n1191 & ~n1265 ;
  assign n3876 = ~n3706 & ~n3875 ;
  assign n3877 = n1265 & ~n1444 ;
  assign n3878 = n1445 & n3877 ;
  assign n3879 = ~n3876 & ~n3878 ;
  assign n3880 = ~n3874 & n3879 ;
  assign n3881 = n3807 & n3880 ;
  assign n3882 = n3873 & n3881 ;
  assign n3883 = n1279 & ~n3705 ;
  assign n3884 = ~n3717 & ~n3883 ;
  assign n3885 = ~n1224 & ~n3884 ;
  assign n3886 = n3882 & n3885 ;
  assign n3887 = n3882 & ~n3884 ;
  assign n3888 = n1224 & ~n3887 ;
  assign n3889 = ~n3886 & ~n3888 ;
  assign n3890 = n3859 & ~n3889 ;
  assign n3891 = ~n3694 & n3890 ;
  assign n3892 = ~n3857 & ~n3891 ;
  assign n3893 = n3856 & n3892 ;
  assign n3894 = ~n3852 & ~n3893 ;
  assign n3895 = ~\g1092_reg/NET0131  & \g2345_reg/NET0131  ;
  assign n3896 = ~\g1092_reg/NET0131  & ~\g2345_reg/NET0131  ;
  assign n3897 = ~n3891 & ~n3896 ;
  assign n3898 = n3856 & n3897 ;
  assign n3899 = ~n3895 & ~n3898 ;
  assign n3900 = ~\g1088_reg/NET0131  & \g2348_reg/NET0131  ;
  assign n3901 = ~\g1088_reg/NET0131  & ~\g2348_reg/NET0131  ;
  assign n3902 = ~n3891 & ~n3901 ;
  assign n3903 = n3856 & n3902 ;
  assign n3904 = ~n3900 & ~n3903 ;
  assign n3905 = \g1092_reg/NET0131  & ~n3842 ;
  assign n3906 = ~\g1092_reg/NET0131  & ~\g234_reg/NET0131  ;
  assign n3907 = ~n3905 & ~n3906 ;
  assign n3908 = \g1088_reg/NET0131  & ~n3842 ;
  assign n3909 = ~\g1088_reg/NET0131  & ~\g237_reg/NET0131  ;
  assign n3910 = ~n3908 & ~n3909 ;
  assign n3911 = n2819 & ~n3048 ;
  assign n3912 = n3069 & n3911 ;
  assign n3913 = n3668 & ~n3912 ;
  assign n3914 = ~n2969 & ~n3913 ;
  assign n3915 = n2969 & n3913 ;
  assign n3916 = ~n3914 & ~n3915 ;
  assign n3917 = ~n3666 & n3916 ;
  assign n3918 = ~n3665 & ~n3917 ;
  assign n3919 = n3645 & ~n3918 ;
  assign n3920 = ~n3637 & n3919 ;
  assign n3921 = \g7961_pad  & n3920 ;
  assign n3922 = ~\g1476_reg/NET0131  & \g7961_pad  ;
  assign n3923 = ~n3680 & n3922 ;
  assign n3924 = ~n3921 & ~n3923 ;
  assign n3925 = ~\g1612_reg/NET0131  & ~\g7961_pad  ;
  assign n3926 = n3924 & ~n3925 ;
  assign n3927 = \g1092_reg/NET0131  & n3920 ;
  assign n3928 = \g1092_reg/NET0131  & ~\g1476_reg/NET0131  ;
  assign n3929 = ~n3680 & n3928 ;
  assign n3930 = ~n3927 & ~n3929 ;
  assign n3931 = ~\g1092_reg/NET0131  & ~\g1615_reg/NET0131  ;
  assign n3932 = n3930 & ~n3931 ;
  assign n3933 = \g1088_reg/NET0131  & n3920 ;
  assign n3934 = \g1088_reg/NET0131  & ~\g1476_reg/NET0131  ;
  assign n3935 = ~n3680 & n3934 ;
  assign n3936 = ~n3933 & ~n3935 ;
  assign n3937 = ~\g1088_reg/NET0131  & ~\g1618_reg/NET0131  ;
  assign n3938 = n3936 & ~n3937 ;
  assign n3939 = ~n2991 & ~n3671 ;
  assign n3940 = n2826 & ~n2991 ;
  assign n3941 = n3646 & n3940 ;
  assign n3942 = ~n3646 & n3659 ;
  assign n3943 = ~n3941 & ~n3942 ;
  assign n3944 = ~n3939 & n3943 ;
  assign n3945 = n2826 & ~n3048 ;
  assign n3946 = n3069 & n3945 ;
  assign n3947 = n3671 & ~n3946 ;
  assign n3948 = n2991 & ~n3048 ;
  assign n3949 = n3069 & n3948 ;
  assign n3950 = ~n3652 & ~n3949 ;
  assign n3951 = n3947 & ~n3950 ;
  assign n3952 = n3944 & ~n3951 ;
  assign n3953 = ~n3666 & n3952 ;
  assign n3954 = ~n3665 & ~n3953 ;
  assign n3955 = n3645 & ~n3954 ;
  assign n3956 = ~n3637 & n3955 ;
  assign n3957 = \g7961_pad  & n3956 ;
  assign n3958 = ~\g1486_reg/NET0131  & \g7961_pad  ;
  assign n3959 = ~n3680 & n3958 ;
  assign n3960 = ~n3957 & ~n3959 ;
  assign n3961 = ~\g1621_reg/NET0131  & ~\g7961_pad  ;
  assign n3962 = n3960 & ~n3961 ;
  assign n3963 = \g1092_reg/NET0131  & n3956 ;
  assign n3964 = \g1092_reg/NET0131  & ~\g1486_reg/NET0131  ;
  assign n3965 = ~n3680 & n3964 ;
  assign n3966 = ~n3963 & ~n3965 ;
  assign n3967 = ~\g1092_reg/NET0131  & ~\g1624_reg/NET0131  ;
  assign n3968 = n3966 & ~n3967 ;
  assign n3969 = ~n2428 & ~n3430 ;
  assign n3970 = n3383 & n3969 ;
  assign n3971 = ~\g109_reg/NET0131  & ~n3970 ;
  assign n3972 = ~\g109_reg/NET0131  & n3406 ;
  assign n3973 = ~n3400 & n3972 ;
  assign n3974 = ~n3971 & ~n3973 ;
  assign n3975 = n2146 & ~n2428 ;
  assign n3976 = n3383 & n3975 ;
  assign n3977 = \g7961_pad  & ~n3976 ;
  assign n3978 = \g7961_pad  & n3406 ;
  assign n3979 = ~n3400 & n3978 ;
  assign n3980 = ~n3977 & ~n3979 ;
  assign n3981 = ~n3974 & ~n3980 ;
  assign n3982 = n2332 & n3385 ;
  assign n3983 = n3414 & ~n3419 ;
  assign n3984 = ~n3982 & ~n3983 ;
  assign n3985 = n3431 & ~n3984 ;
  assign n3986 = ~n3420 & n3985 ;
  assign n3987 = n2361 & ~n3419 ;
  assign n3988 = ~n3385 & ~n3987 ;
  assign n3989 = n3431 & ~n3988 ;
  assign n3990 = ~n2332 & ~n3989 ;
  assign n3991 = ~n3430 & ~n3990 ;
  assign n3992 = ~n3420 & ~n3991 ;
  assign n3993 = ~n3986 & ~n3992 ;
  assign n3994 = n3411 & n3993 ;
  assign n3995 = ~n3410 & n3994 ;
  assign n3996 = \g7961_pad  & n3995 ;
  assign n3997 = ~\g240_reg/NET0131  & ~\g7961_pad  ;
  assign n3998 = ~n3996 & ~n3997 ;
  assign n3999 = ~n3981 & n3998 ;
  assign n4000 = \g1088_reg/NET0131  & n3956 ;
  assign n4001 = \g1088_reg/NET0131  & ~\g1486_reg/NET0131  ;
  assign n4002 = ~n3680 & n4001 ;
  assign n4003 = ~n4000 & ~n4002 ;
  assign n4004 = ~\g1088_reg/NET0131  & ~\g1627_reg/NET0131  ;
  assign n4005 = n4003 & ~n4004 ;
  assign n4006 = \g1092_reg/NET0131  & ~n3976 ;
  assign n4007 = \g1092_reg/NET0131  & n3406 ;
  assign n4008 = ~n3400 & n4007 ;
  assign n4009 = ~n4006 & ~n4008 ;
  assign n4010 = ~n3974 & ~n4009 ;
  assign n4011 = \g1092_reg/NET0131  & n3995 ;
  assign n4012 = ~\g1092_reg/NET0131  & ~\g243_reg/NET0131  ;
  assign n4013 = ~n4011 & ~n4012 ;
  assign n4014 = ~n4010 & n4013 ;
  assign n4015 = ~\g1092_reg/NET0131  & \g1651_reg/NET0131  ;
  assign n4016 = n3645 & n3665 ;
  assign n4017 = ~n3637 & n4016 ;
  assign n4018 = n2928 & ~n3680 ;
  assign n4019 = ~n4017 & ~n4018 ;
  assign n4020 = ~\g1092_reg/NET0131  & ~\g1651_reg/NET0131  ;
  assign n4021 = ~n3066 & ~n3666 ;
  assign n4022 = n3644 & n4021 ;
  assign n4023 = ~n2991 & ~n3048 ;
  assign n4024 = n3069 & n4023 ;
  assign n4025 = ~n3652 & ~n4024 ;
  assign n4026 = n3947 & ~n4025 ;
  assign n4027 = ~n2807 & ~n3646 ;
  assign n4028 = ~n2798 & ~n3048 ;
  assign n4029 = n3069 & n4028 ;
  assign n4030 = ~n3647 & ~n4029 ;
  assign n4031 = n2807 & ~n3048 ;
  assign n4032 = n3069 & n4031 ;
  assign n4033 = n2962 & ~n3048 ;
  assign n4034 = n3069 & n4033 ;
  assign n4035 = ~n4032 & ~n4034 ;
  assign n4036 = ~n4030 & n4035 ;
  assign n4037 = ~n4027 & n4036 ;
  assign n4038 = n4026 & n4037 ;
  assign n4039 = n2790 & ~n3646 ;
  assign n4040 = ~n3658 & ~n4039 ;
  assign n4041 = ~n2978 & ~n3646 ;
  assign n4042 = n2978 & ~n3048 ;
  assign n4043 = n3069 & n4042 ;
  assign n4044 = ~n4041 & ~n4043 ;
  assign n4045 = ~n4040 & n4044 ;
  assign n4046 = n4038 & n4045 ;
  assign n4047 = ~n3000 & ~n4046 ;
  assign n4048 = n3000 & n4045 ;
  assign n4049 = n4038 & n4048 ;
  assign n4050 = ~n4047 & ~n4049 ;
  assign n4051 = n4022 & n4050 ;
  assign n4052 = ~n3637 & n4051 ;
  assign n4053 = ~n4020 & ~n4052 ;
  assign n4054 = n4019 & n4053 ;
  assign n4055 = ~n4015 & ~n4054 ;
  assign n4056 = \g1648_reg/NET0131  & ~\g7961_pad  ;
  assign n4057 = ~\g1648_reg/NET0131  & ~\g7961_pad  ;
  assign n4058 = ~n4052 & ~n4057 ;
  assign n4059 = n4019 & n4058 ;
  assign n4060 = ~n4056 & ~n4059 ;
  assign n4061 = ~\g1088_reg/NET0131  & \g1654_reg/NET0131  ;
  assign n4062 = ~\g1088_reg/NET0131  & ~\g1654_reg/NET0131  ;
  assign n4063 = ~n4052 & ~n4062 ;
  assign n4064 = n4019 & n4063 ;
  assign n4065 = ~n4061 & ~n4064 ;
  assign n4066 = \g267_reg/NET0131  & ~\g7961_pad  ;
  assign n4067 = ~n2428 & n3420 ;
  assign n4068 = n3383 & n4067 ;
  assign n4069 = ~n3410 & n4068 ;
  assign n4070 = n2235 & ~n3396 ;
  assign n4071 = n2235 & n3406 ;
  assign n4072 = ~n3400 & n4071 ;
  assign n4073 = ~n4070 & ~n4072 ;
  assign n4074 = ~n4069 & n4073 ;
  assign n4075 = ~\g267_reg/NET0131  & ~\g7961_pad  ;
  assign n4076 = n2332 & n2368 ;
  assign n4077 = ~n3419 & n4076 ;
  assign n4078 = ~n2332 & ~n2368 ;
  assign n4079 = n3419 & n4078 ;
  assign n4080 = ~n4077 & ~n4079 ;
  assign n4081 = ~n2323 & ~n3419 ;
  assign n4082 = ~n2323 & ~n2349 ;
  assign n4083 = ~n3390 & ~n4082 ;
  assign n4084 = ~n2146 & n2323 ;
  assign n4085 = n2415 & n4084 ;
  assign n4086 = ~n4083 & ~n4085 ;
  assign n4087 = ~n4081 & n4086 ;
  assign n4088 = ~n4080 & n4087 ;
  assign n4089 = n3989 & n4088 ;
  assign n4090 = ~n2294 & ~n3419 ;
  assign n4091 = ~n2146 & n2294 ;
  assign n4092 = n2415 & n4091 ;
  assign n4093 = ~n4090 & ~n4092 ;
  assign n4094 = ~n2302 & ~n3419 ;
  assign n4095 = ~n2146 & n2302 ;
  assign n4096 = n2415 & n4095 ;
  assign n4097 = ~n4094 & ~n4096 ;
  assign n4098 = n4093 & n4097 ;
  assign n4099 = ~n2284 & n4098 ;
  assign n4100 = n4089 & n4099 ;
  assign n4101 = n4089 & n4098 ;
  assign n4102 = n2284 & ~n4101 ;
  assign n4103 = ~n4100 & ~n4102 ;
  assign n4104 = n3970 & ~n4103 ;
  assign n4105 = ~n3410 & n4104 ;
  assign n4106 = ~n4075 & ~n4105 ;
  assign n4107 = n4074 & n4106 ;
  assign n4108 = ~n4066 & ~n4107 ;
  assign n4109 = ~\g1092_reg/NET0131  & \g270_reg/NET0131  ;
  assign n4110 = ~\g1092_reg/NET0131  & ~\g270_reg/NET0131  ;
  assign n4111 = ~n4105 & ~n4110 ;
  assign n4112 = n4074 & n4111 ;
  assign n4113 = ~n4109 & ~n4112 ;
  assign n4114 = ~\g1088_reg/NET0131  & \g273_reg/NET0131  ;
  assign n4115 = ~\g1088_reg/NET0131  & ~\g273_reg/NET0131  ;
  assign n4116 = ~n4105 & ~n4115 ;
  assign n4117 = n4074 & n4116 ;
  assign n4118 = ~n4114 & ~n4117 ;
  assign n4119 = n1816 & n1983 ;
  assign n4120 = n2005 & ~n4119 ;
  assign n4121 = n1931 & n3292 ;
  assign n4122 = ~\g1196_reg/NET0131  & ~\g1916_reg/NET0131  ;
  assign n4123 = ~n3296 & n4122 ;
  assign n4124 = n1998 & n4123 ;
  assign n4125 = ~n1994 & n4124 ;
  assign n4126 = n3295 & ~n4125 ;
  assign n4127 = ~n4121 & n4126 ;
  assign n4128 = ~n4120 & ~n4127 ;
  assign n4129 = ~n1919 & n3292 ;
  assign n4130 = ~\g1196_reg/NET0131  & ~\g1917_reg/NET0131  ;
  assign n4131 = ~n3296 & n4130 ;
  assign n4132 = n1998 & n4131 ;
  assign n4133 = n3295 & ~n4132 ;
  assign n4134 = ~n3302 & ~n4133 ;
  assign n4135 = ~n4129 & ~n4134 ;
  assign n4136 = ~n2005 & ~n4135 ;
  assign n4137 = n1816 & ~n4135 ;
  assign n4138 = n1988 & n4137 ;
  assign n4139 = ~n4136 & ~n4138 ;
  assign n4140 = ~\g1088_reg/NET0131  & \g915_reg/NET0131  ;
  assign n4141 = n2561 & ~n3498 ;
  assign n4142 = ~n3579 & ~n4141 ;
  assign n4143 = ~\g1088_reg/NET0131  & ~\g915_reg/NET0131  ;
  assign n4144 = n3595 & n3605 ;
  assign n4145 = ~n2616 & ~n4144 ;
  assign n4146 = n2616 & n3600 ;
  assign n4147 = n3604 & n4146 ;
  assign n4148 = n3595 & n4147 ;
  assign n4149 = ~n3484 & ~n4148 ;
  assign n4150 = ~n4145 & n4149 ;
  assign n4151 = n3498 & n4150 ;
  assign n4152 = ~n4143 & ~n4151 ;
  assign n4153 = n4142 & n4152 ;
  assign n4154 = ~n4140 & ~n4153 ;
  assign n4155 = ~\g7961_pad  & \g909_reg/NET0131  ;
  assign n4156 = ~\g7961_pad  & ~\g909_reg/NET0131  ;
  assign n4157 = ~n4151 & ~n4156 ;
  assign n4158 = n4142 & n4157 ;
  assign n4159 = ~n4155 & ~n4158 ;
  assign n4160 = ~\g1092_reg/NET0131  & \g912_reg/NET0131  ;
  assign n4161 = ~\g1092_reg/NET0131  & ~\g912_reg/NET0131  ;
  assign n4162 = ~n4151 & ~n4161 ;
  assign n4163 = n4142 & n4162 ;
  assign n4164 = ~n4160 & ~n4163 ;
  assign n4165 = \g222_reg/NET0131  & ~\g7961_pad  ;
  assign n4166 = n2255 & ~n3396 ;
  assign n4167 = n2255 & n3406 ;
  assign n4168 = ~n3400 & n4167 ;
  assign n4169 = ~n4166 & ~n4168 ;
  assign n4170 = ~n4069 & n4169 ;
  assign n4171 = ~\g222_reg/NET0131  & ~\g7961_pad  ;
  assign n4172 = n2302 & n4093 ;
  assign n4173 = n4089 & n4172 ;
  assign n4174 = n4089 & n4093 ;
  assign n4175 = ~n2302 & ~n4174 ;
  assign n4176 = ~n4173 & ~n4175 ;
  assign n4177 = n3970 & n4176 ;
  assign n4178 = ~n3410 & n4177 ;
  assign n4179 = ~n4171 & ~n4178 ;
  assign n4180 = n4170 & n4179 ;
  assign n4181 = ~n4165 & ~n4180 ;
  assign n4182 = ~\g1092_reg/NET0131  & \g225_reg/NET0131  ;
  assign n4183 = ~\g1092_reg/NET0131  & ~\g225_reg/NET0131  ;
  assign n4184 = ~n4178 & ~n4183 ;
  assign n4185 = n4170 & n4184 ;
  assign n4186 = ~n4182 & ~n4185 ;
  assign n4187 = ~\g1088_reg/NET0131  & \g228_reg/NET0131  ;
  assign n4188 = ~\g1088_reg/NET0131  & ~\g228_reg/NET0131  ;
  assign n4189 = ~n4178 & ~n4188 ;
  assign n4190 = n4170 & n4189 ;
  assign n4191 = ~n4187 & ~n4190 ;
  assign n4192 = n1274 & ~n3739 ;
  assign n4193 = ~n1279 & ~n3882 ;
  assign n4194 = n1279 & n3882 ;
  assign n4195 = ~n4193 & ~n4194 ;
  assign n4196 = n3859 & n4195 ;
  assign n4197 = ~n3694 & n4196 ;
  assign n4198 = ~n3854 & ~n4197 ;
  assign n4199 = ~n4192 & n4198 ;
  assign n4200 = \g7961_pad  & ~n4199 ;
  assign n4201 = ~\g2297_reg/NET0131  & ~\g7961_pad  ;
  assign n4202 = ~n4200 & ~n4201 ;
  assign n4203 = \g1092_reg/NET0131  & ~n4199 ;
  assign n4204 = ~\g1092_reg/NET0131  & ~\g2300_reg/NET0131  ;
  assign n4205 = ~n4203 & ~n4204 ;
  assign n4206 = \g1088_reg/NET0131  & ~n4199 ;
  assign n4207 = ~\g1088_reg/NET0131  & ~\g2303_reg/NET0131  ;
  assign n4208 = ~n4206 & ~n4207 ;
  assign n4209 = \g1603_reg/NET0131  & ~\g7961_pad  ;
  assign n4210 = n2785 & ~n3680 ;
  assign n4211 = ~n4017 & ~n4210 ;
  assign n4212 = ~\g1603_reg/NET0131  & ~\g7961_pad  ;
  assign n4213 = n4038 & n4044 ;
  assign n4214 = ~n2790 & ~n4213 ;
  assign n4215 = n2790 & n4044 ;
  assign n4216 = n4038 & n4215 ;
  assign n4217 = ~n3666 & ~n4216 ;
  assign n4218 = ~n4214 & n4217 ;
  assign n4219 = n3645 & n4218 ;
  assign n4220 = ~n3637 & n4219 ;
  assign n4221 = ~n4212 & ~n4220 ;
  assign n4222 = n4211 & n4221 ;
  assign n4223 = ~n4209 & ~n4222 ;
  assign n4224 = ~\g1092_reg/NET0131  & \g1606_reg/NET0131  ;
  assign n4225 = ~\g1092_reg/NET0131  & ~\g1606_reg/NET0131  ;
  assign n4226 = ~n4220 & ~n4225 ;
  assign n4227 = n4211 & n4226 ;
  assign n4228 = ~n4224 & ~n4227 ;
  assign n4229 = ~\g1088_reg/NET0131  & \g1609_reg/NET0131  ;
  assign n4230 = ~\g1088_reg/NET0131  & ~\g1609_reg/NET0131  ;
  assign n4231 = ~n4220 & ~n4230 ;
  assign n4232 = n4211 & n4231 ;
  assign n4233 = ~n4229 & ~n4232 ;
  assign n4234 = ~\g559_reg/NET0131  & ~\g563_pad  ;
  assign n4235 = \g499_reg/NET0131  & ~\g544_reg/NET0131  ;
  assign n4236 = n4234 & n4235 ;
  assign n4237 = \g5657_pad  & ~\g705_reg/NET0131  ;
  assign n4238 = \g1024_reg/NET0131  & ~\g704_reg/NET0131  ;
  assign n4239 = \g1018_reg/NET0131  & ~\g706_reg/NET0131  ;
  assign n4240 = ~n4238 & ~n4239 ;
  assign n4241 = ~n4237 & n4240 ;
  assign n4242 = \g5657_pad  & ~\g714_reg/NET0131  ;
  assign n4243 = \g1024_reg/NET0131  & ~\g713_reg/NET0131  ;
  assign n4244 = \g1018_reg/NET0131  & ~\g715_reg/NET0131  ;
  assign n4245 = ~n4243 & ~n4244 ;
  assign n4246 = ~n4242 & n4245 ;
  assign n4247 = ~n4241 & n4246 ;
  assign n4248 = \g5657_pad  & ~\g720_reg/NET0131  ;
  assign n4249 = \g1024_reg/NET0131  & ~\g719_reg/NET0131  ;
  assign n4250 = \g1018_reg/NET0131  & ~\g721_reg/NET0131  ;
  assign n4251 = ~n4249 & ~n4250 ;
  assign n4252 = ~n4248 & n4251 ;
  assign n4253 = \g5657_pad  & ~\g738_reg/NET0131  ;
  assign n4254 = \g1018_reg/NET0131  & ~\g739_reg/NET0131  ;
  assign n4255 = \g1024_reg/NET0131  & ~\g737_reg/NET0131  ;
  assign n4256 = ~n4254 & ~n4255 ;
  assign n4257 = ~n4253 & n4256 ;
  assign n4258 = n4252 & ~n4257 ;
  assign n4259 = n4247 & n4258 ;
  assign n4260 = \g5657_pad  & ~\g723_reg/NET0131  ;
  assign n4261 = \g1018_reg/NET0131  & ~\g724_reg/NET0131  ;
  assign n4262 = \g1024_reg/NET0131  & ~\g722_reg/NET0131  ;
  assign n4263 = ~n4261 & ~n4262 ;
  assign n4264 = ~n4260 & n4263 ;
  assign n4265 = \g5657_pad  & ~\g702_reg/NET0131  ;
  assign n4266 = \g1024_reg/NET0131  & ~\g701_reg/NET0131  ;
  assign n4267 = \g1018_reg/NET0131  & ~\g703_reg/NET0131  ;
  assign n4268 = ~n4266 & ~n4267 ;
  assign n4269 = ~n4265 & n4268 ;
  assign n4270 = ~n4264 & ~n4269 ;
  assign n4271 = \g5657_pad  & ~\g708_reg/NET0131  ;
  assign n4272 = \g1018_reg/NET0131  & ~\g709_reg/NET0131  ;
  assign n4273 = \g1024_reg/NET0131  & ~\g707_reg/NET0131  ;
  assign n4274 = ~n4272 & ~n4273 ;
  assign n4275 = ~n4271 & n4274 ;
  assign n4276 = \g5657_pad  & ~\g699_reg/NET0131  ;
  assign n4277 = \g1024_reg/NET0131  & ~\g698_reg/NET0131  ;
  assign n4278 = \g1018_reg/NET0131  & ~\g700_reg/NET0131  ;
  assign n4279 = ~n4277 & ~n4278 ;
  assign n4280 = ~n4276 & n4279 ;
  assign n4281 = ~n4275 & n4280 ;
  assign n4282 = n4270 & n4281 ;
  assign n4283 = \g5657_pad  & ~\g726_reg/NET0131  ;
  assign n4284 = \g1024_reg/NET0131  & ~\g725_reg/NET0131  ;
  assign n4285 = \g1018_reg/NET0131  & ~\g727_reg/NET0131  ;
  assign n4286 = ~n4284 & ~n4285 ;
  assign n4287 = ~n4283 & n4286 ;
  assign n4288 = \g1024_reg/NET0131  & ~\g731_reg/NET0131  ;
  assign n4289 = \g5657_pad  & ~\g732_reg/NET0131  ;
  assign n4290 = \g1018_reg/NET0131  & ~\g733_reg/NET0131  ;
  assign n4291 = ~n4289 & ~n4290 ;
  assign n4292 = ~n4288 & n4291 ;
  assign n4293 = ~n4287 & ~n4292 ;
  assign n4294 = \g5657_pad  & ~\g711_reg/NET0131  ;
  assign n4295 = \g1018_reg/NET0131  & ~\g712_reg/NET0131  ;
  assign n4296 = \g1024_reg/NET0131  & ~\g710_reg/NET0131  ;
  assign n4297 = ~n4295 & ~n4296 ;
  assign n4298 = ~n4294 & n4297 ;
  assign n4299 = \g5657_pad  & ~\g717_reg/NET0131  ;
  assign n4300 = \g1024_reg/NET0131  & ~\g716_reg/NET0131  ;
  assign n4301 = \g1018_reg/NET0131  & ~\g718_reg/NET0131  ;
  assign n4302 = ~n4300 & ~n4301 ;
  assign n4303 = ~n4299 & n4302 ;
  assign n4304 = n4298 & n4303 ;
  assign n4305 = n4293 & n4304 ;
  assign n4306 = n4282 & n4305 ;
  assign n4307 = n4259 & n4306 ;
  assign n4308 = \g1024_reg/NET0131  & \g611_reg/NET0131  ;
  assign n4309 = \g5657_pad  & \g605_reg/NET0131  ;
  assign n4310 = \g1018_reg/NET0131  & \g608_reg/NET0131  ;
  assign n4311 = ~n4309 & ~n4310 ;
  assign n4312 = ~n4308 & n4311 ;
  assign n4313 = ~n4275 & n4312 ;
  assign n4314 = ~n4307 & n4313 ;
  assign n4315 = n4275 & ~n4312 ;
  assign n4316 = n4259 & ~n4312 ;
  assign n4317 = n4306 & n4316 ;
  assign n4318 = ~n4315 & ~n4317 ;
  assign n4319 = ~n4314 & n4318 ;
  assign n4320 = n4236 & n4319 ;
  assign n4321 = \g1018_reg/NET0131  & \g617_reg/NET0131  ;
  assign n4322 = \g5657_pad  & \g614_reg/NET0131  ;
  assign n4323 = \g1024_reg/NET0131  & \g620_reg/NET0131  ;
  assign n4324 = ~n4322 & ~n4323 ;
  assign n4325 = ~n4321 & n4324 ;
  assign n4326 = ~n4241 & n4325 ;
  assign n4327 = ~n4307 & n4326 ;
  assign n4328 = n4241 & ~n4325 ;
  assign n4329 = n4259 & ~n4325 ;
  assign n4330 = n4306 & n4329 ;
  assign n4331 = ~n4328 & ~n4330 ;
  assign n4332 = ~n4327 & n4331 ;
  assign n4333 = n4320 & ~n4332 ;
  assign n4334 = n4236 & n4332 ;
  assign n4335 = ~n4319 & n4334 ;
  assign n4336 = ~n4333 & ~n4335 ;
  assign n4337 = ~n4280 & ~n4325 ;
  assign n4338 = n4280 & n4325 ;
  assign n4339 = ~n4337 & ~n4338 ;
  assign n4340 = n4236 & ~n4339 ;
  assign n4341 = ~n4269 & n4312 ;
  assign n4342 = ~n4307 & n4341 ;
  assign n4343 = n4269 & ~n4312 ;
  assign n4344 = ~n4317 & ~n4343 ;
  assign n4345 = ~n4342 & n4344 ;
  assign n4346 = n4340 & ~n4345 ;
  assign n4347 = n4236 & n4339 ;
  assign n4348 = n4345 & n4347 ;
  assign n4349 = ~n4346 & ~n4348 ;
  assign n4350 = ~n4298 & ~n4325 ;
  assign n4351 = n4298 & n4325 ;
  assign n4352 = ~n4350 & ~n4351 ;
  assign n4353 = n4236 & ~n4352 ;
  assign n4354 = n4246 & n4312 ;
  assign n4355 = ~n4246 & ~n4312 ;
  assign n4356 = ~n4354 & ~n4355 ;
  assign n4357 = n4353 & n4356 ;
  assign n4358 = n4236 & ~n4356 ;
  assign n4359 = n4352 & n4358 ;
  assign n4360 = ~n4357 & ~n4359 ;
  assign n4361 = n4252 & n4312 ;
  assign n4362 = ~n4252 & ~n4312 ;
  assign n4363 = ~n4361 & ~n4362 ;
  assign n4364 = n4236 & ~n4363 ;
  assign n4365 = ~n4303 & ~n4325 ;
  assign n4366 = n4303 & n4325 ;
  assign n4367 = ~n4365 & ~n4366 ;
  assign n4368 = n4364 & n4367 ;
  assign n4369 = n4236 & ~n4367 ;
  assign n4370 = n4363 & n4369 ;
  assign n4371 = ~n4368 & ~n4370 ;
  assign n4372 = ~n4360 & ~n4371 ;
  assign n4373 = ~n4349 & n4372 ;
  assign n4374 = ~n4336 & n4373 ;
  assign n4375 = ~n4360 & n4371 ;
  assign n4376 = ~n4349 & n4375 ;
  assign n4377 = n4336 & n4376 ;
  assign n4378 = ~n4374 & ~n4377 ;
  assign n4379 = n4236 & ~n4332 ;
  assign n4380 = n4319 & n4375 ;
  assign n4381 = n4379 & n4380 ;
  assign n4382 = ~n4319 & n4375 ;
  assign n4383 = n4334 & n4382 ;
  assign n4384 = ~n4381 & ~n4383 ;
  assign n4385 = n4349 & ~n4384 ;
  assign n4386 = n4349 & n4372 ;
  assign n4387 = n4336 & n4386 ;
  assign n4388 = ~n4385 & ~n4387 ;
  assign n4389 = n4378 & n4388 ;
  assign n4390 = n4360 & n4371 ;
  assign n4391 = ~n4349 & n4390 ;
  assign n4392 = ~n4336 & n4391 ;
  assign n4393 = n4360 & ~n4371 ;
  assign n4394 = ~n4349 & n4393 ;
  assign n4395 = n4336 & n4394 ;
  assign n4396 = ~n4392 & ~n4395 ;
  assign n4397 = n4319 & n4393 ;
  assign n4398 = n4379 & n4397 ;
  assign n4399 = ~n4319 & n4393 ;
  assign n4400 = n4334 & n4399 ;
  assign n4401 = ~n4398 & ~n4400 ;
  assign n4402 = n4349 & ~n4401 ;
  assign n4403 = n4349 & n4390 ;
  assign n4404 = n4336 & n4403 ;
  assign n4405 = ~n4402 & ~n4404 ;
  assign n4406 = \g1196_reg/NET0131  & n4405 ;
  assign n4407 = n4396 & n4406 ;
  assign n4408 = n4389 & n4407 ;
  assign n4409 = ~n4264 & n4325 ;
  assign n4410 = ~n4307 & n4409 ;
  assign n4411 = n4264 & ~n4325 ;
  assign n4412 = ~n4330 & ~n4411 ;
  assign n4413 = ~n4410 & n4412 ;
  assign n4414 = ~n4287 & n4312 ;
  assign n4415 = ~n4307 & n4414 ;
  assign n4416 = n4287 & ~n4312 ;
  assign n4417 = ~n4317 & ~n4416 ;
  assign n4418 = ~n4415 & n4417 ;
  assign n4419 = ~n4413 & n4418 ;
  assign n4420 = n4413 & ~n4418 ;
  assign n4421 = ~n4419 & ~n4420 ;
  assign n4422 = \g1243_reg/NET0131  & n4236 ;
  assign n4423 = ~n4421 & n4422 ;
  assign n4424 = ~\g499_reg/NET0131  & \g548_reg/NET0131  ;
  assign n4425 = ~\g5657_pad  & n4424 ;
  assign n4426 = ~n1752 & n4234 ;
  assign n4427 = ~n4425 & n4426 ;
  assign n4428 = ~\g499_reg/NET0131  & \g5657_pad  ;
  assign n4429 = n4427 & ~n4428 ;
  assign n4430 = \g525_reg/NET0131  & n1768 ;
  assign n4431 = ~\g3229_pad  & ~\g541_reg/NET0131  ;
  assign n4432 = \g3229_pad  & ~\g538_reg/NET0131  ;
  assign n4433 = ~n4431 & ~n4432 ;
  assign n4434 = n4430 & n4433 ;
  assign n4435 = n4429 & n4434 ;
  assign n4436 = ~n4423 & ~n4435 ;
  assign n4437 = ~n4408 & n4436 ;
  assign n4438 = ~n2123 & ~n2124 ;
  assign n4439 = ~n2124 & n2133 ;
  assign n4440 = ~n2131 & n4439 ;
  assign n4441 = ~n4438 & ~n4440 ;
  assign n4442 = n2146 & ~n2248 ;
  assign n4443 = ~n3399 & n4442 ;
  assign n4444 = \g1563_reg/NET0131  & ~n4443 ;
  assign n4445 = n2269 & ~n4444 ;
  assign n4446 = n2249 & ~n2269 ;
  assign n4447 = ~n3399 & n4446 ;
  assign n4448 = n2249 & ~n2376 ;
  assign n4449 = ~n4447 & ~n4448 ;
  assign n4450 = ~n2146 & ~n4449 ;
  assign n4451 = ~n4445 & ~n4450 ;
  assign n4452 = ~n2151 & ~n2428 ;
  assign n4453 = ~n4451 & n4452 ;
  assign n4454 = n1370 & n1444 ;
  assign n4455 = ~n3686 & n4454 ;
  assign n4456 = n1370 & ~n1444 ;
  assign n4457 = \g1563_reg/NET0131  & ~n4456 ;
  assign n4458 = \g1563_reg/NET0131  & n1260 ;
  assign n4459 = n1304 & n4458 ;
  assign n4460 = ~n4457 & ~n4459 ;
  assign n4461 = ~n4455 & ~n4460 ;
  assign n4462 = ~n1186 & ~n4456 ;
  assign n4463 = ~n1186 & n1260 ;
  assign n4464 = n1304 & n4463 ;
  assign n4465 = ~n4462 & ~n4464 ;
  assign n4466 = ~n1437 & ~n1454 ;
  assign n4467 = n4465 & n4466 ;
  assign n4468 = ~n4461 & n4467 ;
  assign n4469 = ~n2720 & ~n2725 ;
  assign n4470 = ~n2662 & n4469 ;
  assign n4471 = n2453 & n2458 ;
  assign n4472 = ~n4470 & n4471 ;
  assign n4473 = ~\g1563_reg/NET0131  & ~n2454 ;
  assign n4474 = n2457 & n4473 ;
  assign n4475 = ~n2453 & ~n2540 ;
  assign n4476 = \g1563_reg/NET0131  & n4475 ;
  assign n4477 = ~n2742 & n4476 ;
  assign n4478 = ~n4474 & ~n4477 ;
  assign n4479 = ~n4472 & n4478 ;
  assign n4480 = ~n2470 & ~n2598 ;
  assign n4481 = ~n4479 & n4480 ;
  assign n4482 = \g1563_reg/NET0131  & ~n3044 ;
  assign n4483 = n3047 & n4482 ;
  assign n4484 = ~n2779 & n4483 ;
  assign n4485 = ~n3014 & n4484 ;
  assign n4486 = ~n2843 & n4484 ;
  assign n4487 = ~n4485 & ~n4486 ;
  assign n4488 = n2780 & ~n3048 ;
  assign n4489 = \g1563_reg/NET0131  & ~n4488 ;
  assign n4490 = ~n3027 & ~n4489 ;
  assign n4491 = n4487 & ~n4490 ;
  assign n4492 = ~n3020 & ~n4488 ;
  assign n4493 = ~n3020 & n3025 ;
  assign n4494 = n3023 & n4493 ;
  assign n4495 = ~n4492 & ~n4494 ;
  assign n4496 = n3067 & n4495 ;
  assign n4497 = ~n4491 & n4496 ;
  assign n4498 = \g2580_reg/NET0131  & \g2581_reg/NET0131  ;
  assign n4499 = \g1192_reg/NET0131  & ~\g1193_reg/NET0131  ;
  assign n4500 = \g1018_reg/NET0131  & n4499 ;
  assign n4501 = \g506_reg/NET0131  & ~\g507_reg/NET0131  ;
  assign n4502 = \g1018_reg/NET0131  & ~\g1192_reg/NET0131  ;
  assign n4503 = n4501 & n4502 ;
  assign n4504 = ~n4500 & ~n4503 ;
  assign n4505 = ~\g1018_reg/NET0131  & ~\g16399_pad  ;
  assign n4506 = ~\g1886_reg/NET0131  & ~n4505 ;
  assign n4507 = n4504 & n4506 ;
  assign n4508 = \g1886_reg/NET0131  & \g1887_reg/NET0131  ;
  assign n4509 = \g1018_reg/NET0131  & ~n4508 ;
  assign n4510 = ~n4507 & n4509 ;
  assign n4511 = ~\g1018_reg/NET0131  & ~\g16437_pad  ;
  assign n4512 = ~\g2580_reg/NET0131  & ~n4511 ;
  assign n4513 = ~n4510 & n4512 ;
  assign n4514 = ~n4498 & ~n4513 ;
  assign n4515 = \g805_reg/NET0131  & ~n3498 ;
  assign n4516 = n2711 & ~n3595 ;
  assign n4517 = ~n2711 & n3595 ;
  assign n4518 = ~n4516 & ~n4517 ;
  assign n4519 = ~n3484 & n4518 ;
  assign n4520 = n3498 & n4519 ;
  assign n4521 = ~n4515 & ~n4520 ;
  assign n4522 = ~\g117_reg/NET0131  & ~n3411 ;
  assign n4523 = ~\g117_reg/NET0131  & n3406 ;
  assign n4524 = ~n3400 & n4523 ;
  assign n4525 = ~n4522 & ~n4524 ;
  assign n4526 = n3989 & ~n4080 ;
  assign n4527 = ~n2323 & ~n4526 ;
  assign n4528 = n2323 & ~n4080 ;
  assign n4529 = n3989 & n4528 ;
  assign n4530 = ~n4527 & ~n4529 ;
  assign n4531 = ~n3430 & ~n4530 ;
  assign n4532 = n3411 & ~n4531 ;
  assign n4533 = ~n3410 & n4532 ;
  assign n4534 = n4525 & ~n4533 ;
  assign n4535 = n3100 & n3123 ;
  assign n4536 = n3170 & n4535 ;
  assign n4537 = \g1018_reg/NET0131  & ~\g1422_reg/NET0131  ;
  assign n4538 = ~\g1421_reg/NET0131  & \g5657_pad  ;
  assign n4539 = \g1024_reg/NET0131  & ~\g1420_reg/NET0131  ;
  assign n4540 = ~n4538 & ~n4539 ;
  assign n4541 = ~n4537 & n4540 ;
  assign n4542 = n3099 & ~n4541 ;
  assign n4543 = ~n3097 & n4542 ;
  assign n4544 = n2005 & ~n4543 ;
  assign n4545 = ~n4536 & n4544 ;
  assign n4546 = ~\g1211_reg/NET0131  & ~\g1243_reg/NET0131  ;
  assign n4547 = ~\g1196_reg/NET0131  & ~n4546 ;
  assign n4548 = n3099 & ~n4547 ;
  assign n4549 = ~n3097 & n4548 ;
  assign n4550 = ~n3217 & n4549 ;
  assign n4551 = ~\g1196_reg/NET0131  & ~\g1211_reg/NET0131  ;
  assign n4552 = ~\g1243_reg/NET0131  & ~n4551 ;
  assign n4553 = ~\g1215_reg/NET0131  & n3098 ;
  assign n4554 = n4547 & n4553 ;
  assign n4555 = n4552 & ~n4554 ;
  assign n4556 = ~n1750 & n4552 ;
  assign n4557 = ~n3096 & n4556 ;
  assign n4558 = ~n4555 & ~n4557 ;
  assign n4559 = ~n4550 & ~n4558 ;
  assign n4560 = ~n4545 & ~n4559 ;
  assign n4561 = \g1186_reg/NET0131  & n3123 ;
  assign n4562 = n3170 & n4561 ;
  assign n4563 = ~n3097 & n3098 ;
  assign n4564 = \g1186_reg/NET0131  & ~n4541 ;
  assign n4565 = n4563 & ~n4564 ;
  assign n4566 = ~n4562 & n4565 ;
  assign n4567 = n2005 & ~n4566 ;
  assign n4568 = n3099 & ~n3283 ;
  assign n4569 = ~n3097 & n4568 ;
  assign n4570 = ~n3224 & n4569 ;
  assign n4571 = ~\g1217_reg/NET0131  & n3098 ;
  assign n4572 = n4547 & n4571 ;
  assign n4573 = ~n3097 & n4572 ;
  assign n4574 = n4552 & ~n4573 ;
  assign n4575 = ~n4570 & n4574 ;
  assign n4576 = ~n4567 & ~n4575 ;
  assign n4577 = ~n3228 & n4569 ;
  assign n4578 = ~\g1218_reg/NET0131  & n3098 ;
  assign n4579 = n4547 & n4578 ;
  assign n4580 = ~n3097 & n4579 ;
  assign n4581 = n4552 & ~n4580 ;
  assign n4582 = ~n4577 & n4581 ;
  assign n4583 = ~n4545 & ~n4582 ;
  assign n4584 = n2005 & ~n3098 ;
  assign n4585 = ~n1750 & n2005 ;
  assign n4586 = ~n3096 & n4585 ;
  assign n4587 = ~n4584 & ~n4586 ;
  assign n4588 = ~\g1219_reg/NET0131  & n3098 ;
  assign n4589 = n4547 & n4588 ;
  assign n4590 = n4552 & ~n4589 ;
  assign n4591 = ~n4557 & ~n4590 ;
  assign n4592 = n4587 & n4591 ;
  assign n4593 = n4549 & n4587 ;
  assign n4594 = n3195 & n4593 ;
  assign n4595 = ~n4592 & ~n4594 ;
  assign n4596 = ~\g1220_reg/NET0131  & n3098 ;
  assign n4597 = n4547 & n4596 ;
  assign n4598 = n4552 & ~n4597 ;
  assign n4599 = ~n4557 & ~n4598 ;
  assign n4600 = n4587 & n4599 ;
  assign n4601 = n3183 & n4593 ;
  assign n4602 = ~n4600 & ~n4601 ;
  assign n4603 = ~n3213 & n4549 ;
  assign n4604 = ~\g1216_reg/NET0131  & n3098 ;
  assign n4605 = n4547 & n4604 ;
  assign n4606 = ~n3097 & n4605 ;
  assign n4607 = n4552 & ~n4606 ;
  assign n4608 = ~n4603 & n4607 ;
  assign n4609 = ~n4567 & ~n4608 ;
  assign n4610 = \g1496_reg/NET0131  & ~n3680 ;
  assign n4611 = ~n4027 & ~n4032 ;
  assign n4612 = n4026 & n4611 ;
  assign n4613 = n2962 & ~n4612 ;
  assign n4614 = ~n2962 & n4611 ;
  assign n4615 = n4026 & n4614 ;
  assign n4616 = ~n4613 & ~n4615 ;
  assign n4617 = n4022 & n4616 ;
  assign n4618 = ~n3637 & n4617 ;
  assign n4619 = ~n4610 & ~n4618 ;
  assign n4620 = n3411 & n3430 ;
  assign n4621 = ~n3410 & n4620 ;
  assign n4622 = ~\g97_reg/NET0131  & ~n3411 ;
  assign n4623 = ~\g97_reg/NET0131  & n3406 ;
  assign n4624 = ~n3400 & n4623 ;
  assign n4625 = ~n4622 & ~n4624 ;
  assign n4626 = ~n2342 & ~n2415 ;
  assign n4627 = n2342 & n2415 ;
  assign n4628 = ~n4626 & ~n4627 ;
  assign n4629 = ~n3430 & n4628 ;
  assign n4630 = ~n2428 & n4629 ;
  assign n4631 = n3383 & n4630 ;
  assign n4632 = ~n3410 & n4631 ;
  assign n4633 = n4625 & ~n4632 ;
  assign n4634 = ~n4621 & n4633 ;
  assign n4635 = ~\g113_reg/NET0131  & ~n3411 ;
  assign n4636 = ~\g113_reg/NET0131  & n3406 ;
  assign n4637 = ~n3400 & n4636 ;
  assign n4638 = ~n4635 & ~n4637 ;
  assign n4639 = ~n2146 & n2332 ;
  assign n4640 = n2415 & n4639 ;
  assign n4641 = ~n2332 & ~n3419 ;
  assign n4642 = ~n4640 & ~n4641 ;
  assign n4643 = n2368 & n4642 ;
  assign n4644 = n3989 & n4643 ;
  assign n4645 = n3989 & n4642 ;
  assign n4646 = ~n2368 & ~n4645 ;
  assign n4647 = ~n4644 & ~n4646 ;
  assign n4648 = n3970 & n4647 ;
  assign n4649 = ~n3410 & n4648 ;
  assign n4650 = n4638 & ~n4649 ;
  assign n4651 = ~n4621 & n4650 ;
  assign n4652 = \g785_reg/NET0131  & ~n3498 ;
  assign n4653 = n2599 & n2648 ;
  assign n4654 = ~n2599 & ~n2648 ;
  assign n4655 = ~n4653 & ~n4654 ;
  assign n4656 = ~n3484 & ~n4655 ;
  assign n4657 = n3463 & n4656 ;
  assign n4658 = ~n3455 & n4657 ;
  assign n4659 = ~n4652 & ~n4658 ;
  assign n4660 = \g1471_reg/NET0131  & ~n3680 ;
  assign n4661 = n2819 & n3069 ;
  assign n4662 = ~n2819 & ~n3069 ;
  assign n4663 = ~n4661 & ~n4662 ;
  assign n4664 = n4022 & ~n4663 ;
  assign n4665 = ~n3637 & n4664 ;
  assign n4666 = ~n4660 & ~n4665 ;
  assign n4667 = \g801_reg/NET0131  & ~n3498 ;
  assign n4668 = n3585 & n3589 ;
  assign n4669 = n2607 & ~n4668 ;
  assign n4670 = ~n2607 & n3589 ;
  assign n4671 = n3585 & n4670 ;
  assign n4672 = ~n3484 & ~n4671 ;
  assign n4673 = ~n4669 & n4672 ;
  assign n4674 = n3463 & n4673 ;
  assign n4675 = ~n3455 & n4674 ;
  assign n4676 = ~n4667 & ~n4675 ;
  assign n4677 = \g2165_reg/NET0131  & ~n3739 ;
  assign n4678 = ~n1290 & n1445 ;
  assign n4679 = n1290 & ~n1445 ;
  assign n4680 = ~n4678 & ~n4679 ;
  assign n4681 = ~n3725 & n4680 ;
  assign n4682 = n3704 & n4681 ;
  assign n4683 = ~n3694 & n4682 ;
  assign n4684 = ~n4677 & ~n4683 ;
  assign n4685 = ~n3694 & n3859 ;
  assign n4686 = \g2185_reg/NET0131  & ~n3739 ;
  assign n4687 = ~n4685 & ~n4686 ;
  assign n4688 = n1234 & n1297 ;
  assign n4689 = ~n3705 & n4688 ;
  assign n4690 = n3730 & n4689 ;
  assign n4691 = ~n1297 & n3861 ;
  assign n4692 = n3730 & n4691 ;
  assign n4693 = ~n4690 & ~n4692 ;
  assign n4694 = ~n1254 & ~n4693 ;
  assign n4695 = n1254 & n4693 ;
  assign n4696 = ~n4694 & ~n4695 ;
  assign n4697 = ~n3725 & ~n4696 ;
  assign n4698 = n3704 & n4697 ;
  assign n4699 = ~n3694 & n4698 ;
  assign n4700 = ~n4687 & ~n4699 ;
  assign n4701 = \g2195_reg/NET0131  & ~n3739 ;
  assign n4702 = n3807 & n3873 ;
  assign n4703 = n1265 & ~n4702 ;
  assign n4704 = ~n1265 & n3807 ;
  assign n4705 = n3873 & n4704 ;
  assign n4706 = ~n4703 & ~n4705 ;
  assign n4707 = n3859 & n4706 ;
  assign n4708 = ~n3694 & n4707 ;
  assign n4709 = ~n4701 & ~n4708 ;
  assign n4710 = \g1491_reg/NET0131  & ~n3680 ;
  assign n4711 = n2807 & ~n4026 ;
  assign n4712 = ~n2807 & ~n4025 ;
  assign n4713 = n3947 & n4712 ;
  assign n4714 = ~n4711 & ~n4713 ;
  assign n4715 = n4022 & n4714 ;
  assign n4716 = ~n3637 & n4715 ;
  assign n4717 = ~n4710 & ~n4716 ;
  assign n4718 = \g1501_reg/NET0131  & ~n3680 ;
  assign n4719 = ~n2807 & ~n2962 ;
  assign n4720 = n3646 & n4719 ;
  assign n4721 = n2807 & n2962 ;
  assign n4722 = ~n3646 & n4721 ;
  assign n4723 = ~n4720 & ~n4722 ;
  assign n4724 = n4026 & ~n4723 ;
  assign n4725 = ~n2798 & ~n4724 ;
  assign n4726 = n2798 & ~n4723 ;
  assign n4727 = n4026 & n4726 ;
  assign n4728 = ~n4725 & ~n4727 ;
  assign n4729 = n4022 & ~n4728 ;
  assign n4730 = ~n3637 & n4729 ;
  assign n4731 = ~n4718 & ~n4730 ;
  assign n4732 = ~n3455 & n3584 ;
  assign n4733 = \g809_reg/NET0131  & ~n3498 ;
  assign n4734 = ~n4732 & ~n4733 ;
  assign n4735 = ~n2711 & ~n3464 ;
  assign n4736 = ~n3599 & ~n4735 ;
  assign n4737 = ~n2635 & n4736 ;
  assign n4738 = n3595 & n4737 ;
  assign n4739 = n3595 & n4736 ;
  assign n4740 = n2635 & ~n4739 ;
  assign n4741 = ~n4738 & ~n4740 ;
  assign n4742 = n4732 & ~n4741 ;
  assign n4743 = ~n4734 & ~n4742 ;
  assign n4744 = \g2200_reg/NET0131  & ~n3739 ;
  assign n4745 = ~n3874 & ~n3878 ;
  assign n4746 = n3807 & n4745 ;
  assign n4747 = n3873 & n4746 ;
  assign n4748 = ~n1191 & ~n4747 ;
  assign n4749 = n1191 & n4747 ;
  assign n4750 = ~n4748 & ~n4749 ;
  assign n4751 = n3859 & ~n4750 ;
  assign n4752 = ~n3694 & n4751 ;
  assign n4753 = ~n4744 & ~n4752 ;
  assign n4754 = \g1506_reg/NET0131  & ~n3680 ;
  assign n4755 = n2978 & ~n4038 ;
  assign n4756 = ~n2978 & ~n4027 ;
  assign n4757 = n4036 & n4756 ;
  assign n4758 = n4026 & n4757 ;
  assign n4759 = ~n4755 & ~n4758 ;
  assign n4760 = n4022 & n4759 ;
  assign n4761 = ~n3637 & n4760 ;
  assign n4762 = ~n4754 & ~n4761 ;
  assign n4763 = \g813_reg/NET0131  & ~n3498 ;
  assign n4764 = n3595 & n3600 ;
  assign n4765 = n2699 & ~n4764 ;
  assign n4766 = ~n2699 & ~n3599 ;
  assign n4767 = ~n3598 & n4766 ;
  assign n4768 = n3595 & n4767 ;
  assign n4769 = ~n4765 & ~n4768 ;
  assign n4770 = n4732 & n4769 ;
  assign n4771 = ~n4763 & ~n4770 ;
  assign n4772 = \g125_reg/NET0131  & ~n3411 ;
  assign n4773 = \g125_reg/NET0131  & n3406 ;
  assign n4774 = ~n3400 & n4773 ;
  assign n4775 = ~n4772 & ~n4774 ;
  assign n4776 = ~n2294 & ~n4085 ;
  assign n4777 = ~n4081 & n4776 ;
  assign n4778 = ~n4083 & n4777 ;
  assign n4779 = n4526 & n4778 ;
  assign n4780 = n2294 & ~n4089 ;
  assign n4781 = ~n4779 & ~n4780 ;
  assign n4782 = n3970 & n4781 ;
  assign n4783 = ~n3410 & n4782 ;
  assign n4784 = n4775 & ~n4783 ;
  assign n4785 = n1760 & ~n1772 ;
  assign n4786 = n3100 & n3272 ;
  assign n4787 = n2005 & ~n4786 ;
  assign n4788 = ~n3204 & ~n3283 ;
  assign n4789 = n3123 & ~n3283 ;
  assign n4790 = n3170 & n4789 ;
  assign n4791 = ~n4788 & ~n4790 ;
  assign n4792 = n3208 & ~n4791 ;
  assign n4793 = ~\g1222_reg/NET0131  & n3098 ;
  assign n4794 = n4547 & n4793 ;
  assign n4795 = ~n3097 & n4794 ;
  assign n4796 = n4552 & ~n4795 ;
  assign n4797 = ~n4792 & n4796 ;
  assign n4798 = ~n4787 & ~n4797 ;
  assign n4799 = ~n3202 & n4569 ;
  assign n4800 = ~\g1223_reg/NET0131  & n3098 ;
  assign n4801 = n4547 & n4800 ;
  assign n4802 = ~n3097 & n4801 ;
  assign n4803 = n4552 & ~n4802 ;
  assign n4804 = ~n4799 & n4803 ;
  assign n4805 = ~n2005 & ~n4804 ;
  assign n4806 = n3100 & ~n4804 ;
  assign n4807 = n3277 & n4806 ;
  assign n4808 = ~n4805 & ~n4807 ;
  assign n4809 = ~n2131 & ~n2132 ;
  assign n4810 = ~n2151 & ~n3377 ;
  assign n4811 = n2249 & n4810 ;
  assign n4812 = ~n3399 & n4811 ;
  assign n4813 = ~n3419 & ~n4812 ;
  assign n4814 = ~n2428 & ~n4813 ;
  assign n4815 = ~n2598 & n3464 ;
  assign n4816 = ~n2470 & ~n3456 ;
  assign n4817 = ~n2598 & n4816 ;
  assign n4818 = ~n4470 & n4817 ;
  assign n4819 = ~n4815 & ~n4818 ;
  assign n4820 = ~n1454 & n3705 ;
  assign n4821 = n1370 & ~n1437 ;
  assign n4822 = ~n3695 & n4821 ;
  assign n4823 = ~n1454 & n4822 ;
  assign n4824 = ~n3686 & n4823 ;
  assign n4825 = ~n4820 & ~n4824 ;
  assign n4826 = ~n3036 & ~n3638 ;
  assign n4827 = n2780 & n4826 ;
  assign n4828 = ~n3014 & n4827 ;
  assign n4829 = ~n2843 & n4827 ;
  assign n4830 = ~n4828 & ~n4829 ;
  assign n4831 = ~n3646 & n4830 ;
  assign n4832 = ~n3066 & ~n4831 ;
  assign n4833 = ~\g1243_reg/NET0131  & ~\g525_reg/NET0131  ;
  assign n4834 = ~\g1196_reg/NET0131  & ~n4833 ;
  assign n4835 = n4236 & ~n4834 ;
  assign n4836 = ~n4367 & n4835 ;
  assign n4837 = ~\g1196_reg/NET0131  & ~\g525_reg/NET0131  ;
  assign n4838 = ~\g1243_reg/NET0131  & ~n4837 ;
  assign n4839 = ~\g530_reg/NET0131  & ~n4428 ;
  assign n4840 = n4834 & n4839 ;
  assign n4841 = n4427 & n4840 ;
  assign n4842 = n4838 & ~n4841 ;
  assign n4843 = ~n4836 & n4842 ;
  assign n4844 = ~n2005 & ~n4843 ;
  assign n4845 = \g5657_pad  & ~\g735_reg/NET0131  ;
  assign n4846 = \g1018_reg/NET0131  & ~\g736_reg/NET0131  ;
  assign n4847 = \g1024_reg/NET0131  & ~\g734_reg/NET0131  ;
  assign n4848 = ~n4846 & ~n4847 ;
  assign n4849 = ~n4845 & n4848 ;
  assign n4850 = \g499_reg/NET0131  & ~n4849 ;
  assign n4851 = \g499_reg/NET0131  & n4259 ;
  assign n4852 = n4306 & n4851 ;
  assign n4853 = ~n4850 & ~n4852 ;
  assign n4854 = n4429 & ~n4843 ;
  assign n4855 = n4853 & n4854 ;
  assign n4856 = ~n4844 & ~n4855 ;
  assign n4857 = ~n4356 & n4835 ;
  assign n4858 = ~\g531_reg/NET0131  & ~n4428 ;
  assign n4859 = n4834 & n4858 ;
  assign n4860 = n4427 & n4859 ;
  assign n4861 = n4838 & ~n4860 ;
  assign n4862 = ~n4857 & n4861 ;
  assign n4863 = ~n2005 & ~n4862 ;
  assign n4864 = n4429 & ~n4862 ;
  assign n4865 = n4853 & n4864 ;
  assign n4866 = ~n4863 & ~n4865 ;
  assign n4867 = ~n4363 & n4835 ;
  assign n4868 = ~\g529_reg/NET0131  & ~n4428 ;
  assign n4869 = n4834 & n4868 ;
  assign n4870 = n4427 & n4869 ;
  assign n4871 = n4838 & ~n4870 ;
  assign n4872 = ~n4867 & n4871 ;
  assign n4873 = ~n2005 & ~n4872 ;
  assign n4874 = n4427 & ~n4872 ;
  assign n4875 = ~n4853 & n4874 ;
  assign n4876 = ~n4873 & ~n4875 ;
  assign n4877 = ~n4352 & n4835 ;
  assign n4878 = ~\g532_reg/NET0131  & ~n4428 ;
  assign n4879 = n4834 & n4878 ;
  assign n4880 = n4427 & n4879 ;
  assign n4881 = n4838 & ~n4880 ;
  assign n4882 = ~n4877 & n4881 ;
  assign n4883 = ~n2005 & ~n4882 ;
  assign n4884 = n4427 & ~n4882 ;
  assign n4885 = ~n4853 & n4884 ;
  assign n4886 = ~n4883 & ~n4885 ;
  assign n4887 = n2005 & ~n4429 ;
  assign n4888 = ~\g533_reg/NET0131  & ~n4428 ;
  assign n4889 = n4834 & n4888 ;
  assign n4890 = n4427 & n4889 ;
  assign n4891 = n4838 & ~n4890 ;
  assign n4892 = ~n4887 & ~n4891 ;
  assign n4893 = n4835 & ~n4887 ;
  assign n4894 = n4319 & n4893 ;
  assign n4895 = ~n4892 & ~n4894 ;
  assign n4896 = ~\g534_reg/NET0131  & ~n4428 ;
  assign n4897 = n4834 & n4896 ;
  assign n4898 = n4427 & n4897 ;
  assign n4899 = n4838 & ~n4898 ;
  assign n4900 = ~n4887 & ~n4899 ;
  assign n4901 = n4332 & n4893 ;
  assign n4902 = ~n4900 & ~n4901 ;
  assign n4903 = ~n4507 & ~n4508 ;
  assign n4904 = \g1018_reg/NET0131  & \g1038_reg/NET0131  ;
  assign n4905 = \g1036_reg/NET0131  & \g5657_pad  ;
  assign n4906 = \g1024_reg/NET0131  & \g1040_reg/NET0131  ;
  assign n4907 = ~n4905 & ~n4906 ;
  assign n4908 = ~n4904 & n4907 ;
  assign n4909 = \g1024_reg/NET0131  & \g1055_reg/NET0131  ;
  assign n4910 = \g1051_reg/NET0131  & \g5657_pad  ;
  assign n4911 = \g1018_reg/NET0131  & \g1053_reg/NET0131  ;
  assign n4912 = ~n4910 & ~n4911 ;
  assign n4913 = ~n4909 & n4912 ;
  assign n4914 = n4908 & n4913 ;
  assign n4915 = ~\g1262_reg/NET0131  & \g5657_pad  ;
  assign n4916 = \g1024_reg/NET0131  & ~\g1261_reg/NET0131  ;
  assign n4917 = \g1018_reg/NET0131  & ~\g1263_reg/NET0131  ;
  assign n4918 = ~n4916 & ~n4917 ;
  assign n4919 = ~n4915 & n4918 ;
  assign n4920 = \g1024_reg/NET0131  & ~\g1264_reg/NET0131  ;
  assign n4921 = \g1018_reg/NET0131  & ~\g1266_reg/NET0131  ;
  assign n4922 = ~\g1265_reg/NET0131  & \g5657_pad  ;
  assign n4923 = ~n4921 & ~n4922 ;
  assign n4924 = ~n4920 & n4923 ;
  assign n4925 = ~n4919 & n4924 ;
  assign n4926 = n4914 & n4925 ;
  assign n4927 = \g1024_reg/NET0131  & \g1070_reg/NET0131  ;
  assign n4928 = \g1066_reg/NET0131  & \g5657_pad  ;
  assign n4929 = \g1018_reg/NET0131  & \g1068_reg/NET0131  ;
  assign n4930 = ~n4928 & ~n4929 ;
  assign n4931 = ~n4927 & n4930 ;
  assign n4932 = ~n4913 & ~n4931 ;
  assign n4933 = ~n4908 & n4932 ;
  assign n4934 = \g1018_reg/NET0131  & ~\g1269_reg/NET0131  ;
  assign n4935 = ~\g1268_reg/NET0131  & \g5657_pad  ;
  assign n4936 = \g1024_reg/NET0131  & ~\g1267_reg/NET0131  ;
  assign n4937 = ~n4935 & ~n4936 ;
  assign n4938 = ~n4934 & n4937 ;
  assign n4939 = n4919 & ~n4938 ;
  assign n4940 = n4933 & n4939 ;
  assign n4941 = ~n4926 & ~n4940 ;
  assign n4942 = n4908 & n4931 ;
  assign n4943 = n4913 & ~n4938 ;
  assign n4944 = ~n4919 & n4943 ;
  assign n4945 = ~n4942 & n4944 ;
  assign n4946 = n4941 & ~n4945 ;
  assign n4947 = n4908 & n4924 ;
  assign n4948 = n4932 & n4947 ;
  assign n4949 = n4919 & n4948 ;
  assign n4950 = \g1024_reg/NET0131  & ~\g1270_reg/NET0131  ;
  assign n4951 = \g1018_reg/NET0131  & ~\g1272_reg/NET0131  ;
  assign n4952 = ~\g1271_reg/NET0131  & \g5657_pad  ;
  assign n4953 = ~n4951 & ~n4952 ;
  assign n4954 = ~n4950 & n4953 ;
  assign n4955 = ~n4908 & n4954 ;
  assign n4956 = n4938 & ~n4955 ;
  assign n4957 = \g1011_reg/NET0131  & \g1024_reg/NET0131  ;
  assign n4958 = \g1081_reg/NET0131  & \g5657_pad  ;
  assign n4959 = \g1018_reg/NET0131  & \g1083_reg/NET0131  ;
  assign n4960 = ~n4958 & ~n4959 ;
  assign n4961 = ~n4957 & n4960 ;
  assign n4962 = n4919 & n4961 ;
  assign n4963 = ~n4956 & n4962 ;
  assign n4964 = ~n4949 & ~n4963 ;
  assign n4965 = ~n4908 & n4931 ;
  assign n4966 = ~n4924 & ~n4943 ;
  assign n4967 = n4965 & n4966 ;
  assign n4968 = n4964 & ~n4967 ;
  assign n4969 = n4946 & n4968 ;
  assign n4970 = \g1018_reg/NET0131  & \g1253_reg/NET0131  ;
  assign n4971 = \g1251_reg/NET0131  & \g5657_pad  ;
  assign n4972 = \g1024_reg/NET0131  & \g1176_reg/NET0131  ;
  assign n4973 = ~n4971 & ~n4972 ;
  assign n4974 = ~n4970 & n4973 ;
  assign n4975 = \g1228_reg/NET0131  & \g185_reg/NET0131  ;
  assign n4976 = ~n4974 & n4975 ;
  assign n4977 = \g1018_reg/NET0131  & \g1285_reg/NET0131  ;
  assign n4978 = \g1282_reg/NET0131  & \g5657_pad  ;
  assign n4979 = \g1024_reg/NET0131  & \g1288_reg/NET0131  ;
  assign n4980 = ~n4978 & ~n4979 ;
  assign n4981 = ~n4977 & n4980 ;
  assign n4982 = ~n4976 & n4981 ;
  assign n4983 = n4931 & ~n4954 ;
  assign n4984 = n4924 & n4938 ;
  assign n4985 = ~n4913 & n4931 ;
  assign n4986 = n4984 & n4985 ;
  assign n4987 = ~n4983 & ~n4986 ;
  assign n4988 = ~n4919 & ~n4954 ;
  assign n4989 = ~n4961 & n4988 ;
  assign n4990 = n4908 & ~n4989 ;
  assign n4991 = n4987 & n4990 ;
  assign n4992 = n4913 & ~n4931 ;
  assign n4993 = ~n4919 & n4954 ;
  assign n4994 = n4992 & n4993 ;
  assign n4995 = ~n4913 & ~n4961 ;
  assign n4996 = ~n4924 & n4938 ;
  assign n4997 = n4995 & n4996 ;
  assign n4998 = ~n4994 & ~n4997 ;
  assign n4999 = ~n4908 & n4998 ;
  assign n5000 = ~n4991 & ~n4999 ;
  assign n5001 = n4982 & ~n5000 ;
  assign n5002 = n4969 & n5001 ;
  assign n5003 = ~n4924 & n4942 ;
  assign n5004 = n4961 & n4984 ;
  assign n5005 = ~n5003 & ~n5004 ;
  assign n5006 = ~n4919 & ~n5005 ;
  assign n5007 = n4919 & ~n4924 ;
  assign n5008 = n4992 & n5007 ;
  assign n5009 = ~n5006 & ~n5008 ;
  assign n5010 = ~n4908 & ~n4984 ;
  assign n5011 = ~n4908 & n4919 ;
  assign n5012 = ~n4919 & ~n4938 ;
  assign n5013 = ~n5011 & ~n5012 ;
  assign n5014 = ~n5010 & ~n5013 ;
  assign n5015 = n4995 & n5014 ;
  assign n5016 = n4943 & n5011 ;
  assign n5017 = n4914 & n4996 ;
  assign n5018 = ~n5016 & ~n5017 ;
  assign n5019 = ~n5015 & n5018 ;
  assign n5020 = n5009 & n5019 ;
  assign n5021 = n4948 & n4993 ;
  assign n5022 = n4919 & n4924 ;
  assign n5023 = n4965 & n5022 ;
  assign n5024 = n4954 & n5023 ;
  assign n5025 = ~n5021 & ~n5024 ;
  assign n5026 = ~n4908 & ~n4954 ;
  assign n5027 = n4932 & n5026 ;
  assign n5028 = \g1255_reg/NET0131  & \g5657_pad  ;
  assign n5029 = \g1018_reg/NET0131  & \g1257_reg/NET0131  ;
  assign n5030 = \g1024_reg/NET0131  & \g1259_reg/NET0131  ;
  assign n5031 = ~n5029 & ~n5030 ;
  assign n5032 = ~n5028 & n5031 ;
  assign n5033 = \g1210_reg/NET0131  & \g185_reg/NET0131  ;
  assign n5034 = ~n5032 & n5033 ;
  assign n5035 = \g1024_reg/NET0131  & \g1279_reg/NET0131  ;
  assign n5036 = \g1273_reg/NET0131  & \g5657_pad  ;
  assign n5037 = \g1018_reg/NET0131  & \g1276_reg/NET0131  ;
  assign n5038 = ~n5036 & ~n5037 ;
  assign n5039 = ~n5035 & n5038 ;
  assign n5040 = ~n5034 & n5039 ;
  assign n5041 = ~n4982 & ~n5040 ;
  assign n5042 = ~n5027 & ~n5041 ;
  assign n5043 = n5025 & n5042 ;
  assign n5044 = n5020 & n5043 ;
  assign n5045 = ~n5002 & n5044 ;
  assign n5046 = ~\g3010_reg/NET0131  & \g3013_reg/NET0131  ;
  assign n5047 = \g3024_reg/NET0131  & n5046 ;
  assign n5048 = \g3002_reg/NET0131  & ~\g3006_reg/NET0131  ;
  assign n5049 = ~\g2993_reg/NET0131  & \g2998_reg/NET0131  ;
  assign n5050 = n5048 & n5049 ;
  assign n5051 = n5047 & n5050 ;
  assign n5052 = ~\g3032_reg/NET0131  & ~\g3036_reg/NET0131  ;
  assign n5053 = \g3018_reg/NET0131  & \g3028_reg/NET0131  ;
  assign n5054 = \g1024_reg/NET0131  & n5053 ;
  assign n5055 = n5052 & n5054 ;
  assign n5056 = n5051 & n5055 ;
  assign n5057 = ~n5045 & n5056 ;
  assign n5058 = n5052 & n5053 ;
  assign n5059 = n5051 & n5058 ;
  assign n5060 = \g1024_reg/NET0131  & n3176 ;
  assign n5061 = ~n5059 & n5060 ;
  assign n5062 = ~\g1024_reg/NET0131  & ~\g1306_reg/NET0131  ;
  assign n5063 = ~n5061 & ~n5062 ;
  assign n5064 = ~n5057 & n5063 ;
  assign n5065 = \g1018_reg/NET0131  & \g2426_reg/NET0131  ;
  assign n5066 = \g2424_reg/NET0131  & \g5657_pad  ;
  assign n5067 = \g1024_reg/NET0131  & \g2428_reg/NET0131  ;
  assign n5068 = ~n5066 & ~n5067 ;
  assign n5069 = ~n5065 & n5068 ;
  assign n5070 = \g1018_reg/NET0131  & \g2441_reg/NET0131  ;
  assign n5071 = \g2439_reg/NET0131  & \g5657_pad  ;
  assign n5072 = \g1024_reg/NET0131  & \g2443_reg/NET0131  ;
  assign n5073 = ~n5071 & ~n5072 ;
  assign n5074 = ~n5070 & n5073 ;
  assign n5075 = n5069 & n5074 ;
  assign n5076 = ~\g2653_reg/NET0131  & \g5657_pad  ;
  assign n5077 = \g1018_reg/NET0131  & ~\g2654_reg/NET0131  ;
  assign n5078 = \g1024_reg/NET0131  & ~\g2652_reg/NET0131  ;
  assign n5079 = ~n5077 & ~n5078 ;
  assign n5080 = ~n5076 & n5079 ;
  assign n5081 = ~\g2650_reg/NET0131  & \g5657_pad  ;
  assign n5082 = \g1024_reg/NET0131  & ~\g2649_reg/NET0131  ;
  assign n5083 = \g1018_reg/NET0131  & ~\g2651_reg/NET0131  ;
  assign n5084 = ~n5082 & ~n5083 ;
  assign n5085 = ~n5081 & n5084 ;
  assign n5086 = n5080 & ~n5085 ;
  assign n5087 = n5075 & n5086 ;
  assign n5088 = ~n5069 & n5074 ;
  assign n5089 = \g1018_reg/NET0131  & ~\g2657_reg/NET0131  ;
  assign n5090 = \g1024_reg/NET0131  & ~\g2655_reg/NET0131  ;
  assign n5091 = ~\g2656_reg/NET0131  & \g5657_pad  ;
  assign n5092 = ~n5090 & ~n5091 ;
  assign n5093 = ~n5089 & n5092 ;
  assign n5094 = ~n5085 & ~n5093 ;
  assign n5095 = n5088 & n5094 ;
  assign n5096 = ~n5087 & ~n5095 ;
  assign n5097 = \g1018_reg/NET0131  & \g2456_reg/NET0131  ;
  assign n5098 = \g2454_reg/NET0131  & \g5657_pad  ;
  assign n5099 = \g1024_reg/NET0131  & \g2458_reg/NET0131  ;
  assign n5100 = ~n5098 & ~n5099 ;
  assign n5101 = ~n5097 & n5100 ;
  assign n5102 = ~n5069 & n5101 ;
  assign n5103 = ~n5074 & ~n5080 ;
  assign n5104 = n5102 & n5103 ;
  assign n5105 = n5096 & ~n5104 ;
  assign n5106 = n5069 & n5101 ;
  assign n5107 = ~\g2659_reg/NET0131  & \g5657_pad  ;
  assign n5108 = \g1018_reg/NET0131  & ~\g2660_reg/NET0131  ;
  assign n5109 = \g1024_reg/NET0131  & ~\g2658_reg/NET0131  ;
  assign n5110 = ~n5108 & ~n5109 ;
  assign n5111 = ~n5107 & n5110 ;
  assign n5112 = n5106 & ~n5111 ;
  assign n5113 = n5069 & ~n5085 ;
  assign n5114 = \g1018_reg/NET0131  & \g2471_reg/NET0131  ;
  assign n5115 = \g2469_reg/NET0131  & \g5657_pad  ;
  assign n5116 = \g1024_reg/NET0131  & \g2399_reg/NET0131  ;
  assign n5117 = ~n5115 & ~n5116 ;
  assign n5118 = ~n5114 & n5117 ;
  assign n5119 = ~n5111 & ~n5118 ;
  assign n5120 = n5113 & n5119 ;
  assign n5121 = ~n5112 & ~n5120 ;
  assign n5122 = ~n5069 & n5085 ;
  assign n5123 = n5111 & n5118 ;
  assign n5124 = n5122 & n5123 ;
  assign n5125 = n5121 & ~n5124 ;
  assign n5126 = n5105 & n5125 ;
  assign n5127 = n5074 & ~n5101 ;
  assign n5128 = ~n5085 & n5111 ;
  assign n5129 = ~n5069 & n5128 ;
  assign n5130 = ~n5094 & ~n5129 ;
  assign n5131 = n5127 & ~n5130 ;
  assign n5132 = n5085 & ~n5093 ;
  assign n5133 = ~n5074 & ~n5101 ;
  assign n5134 = ~n5069 & n5133 ;
  assign n5135 = ~n5118 & ~n5134 ;
  assign n5136 = n5132 & ~n5135 ;
  assign n5137 = ~n5131 & ~n5136 ;
  assign n5138 = n5126 & n5137 ;
  assign n5139 = ~n5074 & ~n5118 ;
  assign n5140 = ~n5101 & ~n5139 ;
  assign n5141 = ~n5080 & n5093 ;
  assign n5142 = ~n5069 & n5141 ;
  assign n5143 = ~n5140 & n5142 ;
  assign n5144 = n5080 & n5093 ;
  assign n5145 = ~n5074 & n5106 ;
  assign n5146 = n5144 & n5145 ;
  assign n5147 = ~n5143 & ~n5146 ;
  assign n5148 = \g1024_reg/NET0131  & \g2564_reg/NET0131  ;
  assign n5149 = \g2639_reg/NET0131  & \g5657_pad  ;
  assign n5150 = \g1018_reg/NET0131  & \g2641_reg/NET0131  ;
  assign n5151 = ~n5149 & ~n5150 ;
  assign n5152 = ~n5148 & n5151 ;
  assign n5153 = \g185_reg/NET0131  & \g2616_reg/NET0131  ;
  assign n5154 = ~n5152 & n5153 ;
  assign n5155 = \g1024_reg/NET0131  & \g2676_reg/NET0131  ;
  assign n5156 = \g2670_reg/NET0131  & \g5657_pad  ;
  assign n5157 = \g1018_reg/NET0131  & \g2673_reg/NET0131  ;
  assign n5158 = ~n5156 & ~n5157 ;
  assign n5159 = ~n5155 & n5158 ;
  assign n5160 = ~n5154 & n5159 ;
  assign n5161 = n5069 & n5133 ;
  assign n5162 = n5080 & n5085 ;
  assign n5163 = n5161 & n5162 ;
  assign n5164 = n5160 & ~n5163 ;
  assign n5165 = n5147 & n5164 ;
  assign n5166 = n5138 & n5165 ;
  assign n5167 = n5075 & ~n5080 ;
  assign n5168 = n5086 & n5118 ;
  assign n5169 = ~n5167 & ~n5168 ;
  assign n5170 = n5093 & ~n5169 ;
  assign n5171 = n5122 & n5144 ;
  assign n5172 = ~n5093 & n5113 ;
  assign n5173 = ~n5171 & ~n5172 ;
  assign n5174 = n5139 & ~n5173 ;
  assign n5175 = ~n5080 & n5085 ;
  assign n5176 = n5127 & n5175 ;
  assign n5177 = ~n5080 & ~n5085 ;
  assign n5178 = n5106 & n5177 ;
  assign n5179 = ~n5176 & ~n5178 ;
  assign n5180 = n5088 & n5132 ;
  assign n5181 = n5179 & ~n5180 ;
  assign n5182 = ~n5174 & n5181 ;
  assign n5183 = ~n5170 & n5182 ;
  assign n5184 = ~n5069 & ~n5111 ;
  assign n5185 = n5133 & n5184 ;
  assign n5186 = n5086 & n5111 ;
  assign n5187 = n5161 & n5186 ;
  assign n5188 = ~n5185 & ~n5187 ;
  assign n5189 = n5102 & n5162 ;
  assign n5190 = n5111 & n5189 ;
  assign n5191 = \g2643_reg/NET0131  & \g5657_pad  ;
  assign n5192 = \g1018_reg/NET0131  & \g2645_reg/NET0131  ;
  assign n5193 = \g1024_reg/NET0131  & \g2647_reg/NET0131  ;
  assign n5194 = ~n5192 & ~n5193 ;
  assign n5195 = ~n5191 & n5194 ;
  assign n5196 = \g185_reg/NET0131  & \g2598_reg/NET0131  ;
  assign n5197 = ~n5195 & n5196 ;
  assign n5198 = \g1024_reg/NET0131  & \g2667_reg/NET0131  ;
  assign n5199 = \g2661_reg/NET0131  & \g5657_pad  ;
  assign n5200 = \g1018_reg/NET0131  & \g2664_reg/NET0131  ;
  assign n5201 = ~n5199 & ~n5200 ;
  assign n5202 = ~n5198 & n5201 ;
  assign n5203 = ~n5197 & n5202 ;
  assign n5204 = ~n5160 & ~n5203 ;
  assign n5205 = ~n5190 & ~n5204 ;
  assign n5206 = n5188 & n5205 ;
  assign n5207 = n5183 & n5206 ;
  assign n5208 = ~n5166 & n5207 ;
  assign n5209 = \g5657_pad  & n5053 ;
  assign n5210 = n5052 & n5209 ;
  assign n5211 = n5051 & n5210 ;
  assign n5212 = ~n5208 & n5211 ;
  assign n5213 = \g5657_pad  & n1589 ;
  assign n5214 = ~n5059 & n5213 ;
  assign n5215 = ~\g2688_reg/NET0131  & ~\g5657_pad  ;
  assign n5216 = ~n5214 & ~n5215 ;
  assign n5217 = ~n5212 & n5216 ;
  assign n5218 = \g1018_reg/NET0131  & n5053 ;
  assign n5219 = n5052 & n5218 ;
  assign n5220 = n5051 & n5219 ;
  assign n5221 = ~n5208 & n5220 ;
  assign n5222 = \g1018_reg/NET0131  & n1589 ;
  assign n5223 = ~n5059 & n5222 ;
  assign n5224 = ~\g1018_reg/NET0131  & ~\g2691_reg/NET0131  ;
  assign n5225 = ~n5223 & ~n5224 ;
  assign n5226 = ~n5221 & n5225 ;
  assign n5227 = n5056 & ~n5208 ;
  assign n5228 = \g1024_reg/NET0131  & n1589 ;
  assign n5229 = ~n5059 & n5228 ;
  assign n5230 = ~\g1024_reg/NET0131  & ~\g2694_reg/NET0131  ;
  assign n5231 = ~n5229 & ~n5230 ;
  assign n5232 = ~n5227 & n5231 ;
  assign n5233 = n4236 & n4418 ;
  assign n5234 = n2005 & ~n5233 ;
  assign n5235 = n4345 & n4835 ;
  assign n5236 = ~\g536_reg/NET0131  & ~n4428 ;
  assign n5237 = n4834 & n5236 ;
  assign n5238 = n4427 & n5237 ;
  assign n5239 = n4838 & ~n5238 ;
  assign n5240 = ~n5235 & n5239 ;
  assign n5241 = ~n5234 & ~n5240 ;
  assign n5242 = ~n4339 & n4835 ;
  assign n5243 = ~\g537_reg/NET0131  & ~n4428 ;
  assign n5244 = n4834 & n5243 ;
  assign n5245 = n4427 & n5244 ;
  assign n5246 = n4838 & ~n5245 ;
  assign n5247 = ~n5242 & n5246 ;
  assign n5248 = ~n2005 & ~n5247 ;
  assign n5249 = n4236 & ~n5247 ;
  assign n5250 = n4413 & n5249 ;
  assign n5251 = ~n5248 & ~n5250 ;
  assign n5252 = ~n1745 & ~n1994 ;
  assign n5253 = ~\g2679_reg/NET0131  & ~\g5657_pad  ;
  assign n5254 = n5188 & ~n5190 ;
  assign n5255 = ~n5170 & n5203 ;
  assign n5256 = n5182 & n5255 ;
  assign n5257 = n5254 & n5256 ;
  assign n5258 = n5147 & ~n5163 ;
  assign n5259 = n5059 & ~n5204 ;
  assign n5260 = n5258 & n5259 ;
  assign n5261 = n5138 & n5260 ;
  assign n5262 = ~n5257 & n5261 ;
  assign n5263 = \g2679_reg/NET0131  & ~\g5657_pad  ;
  assign n5264 = ~n1673 & ~n5059 ;
  assign n5265 = ~n5263 & ~n5264 ;
  assign n5266 = ~n5262 & n5265 ;
  assign n5267 = ~n5253 & ~n5266 ;
  assign n5268 = ~\g1018_reg/NET0131  & ~\g2682_reg/NET0131  ;
  assign n5269 = ~\g1018_reg/NET0131  & \g2682_reg/NET0131  ;
  assign n5270 = ~n5264 & ~n5269 ;
  assign n5271 = ~n5262 & n5270 ;
  assign n5272 = ~n5268 & ~n5271 ;
  assign n5273 = ~\g1024_reg/NET0131  & ~\g2685_reg/NET0131  ;
  assign n5274 = ~\g1024_reg/NET0131  & \g2685_reg/NET0131  ;
  assign n5275 = ~n5264 & ~n5274 ;
  assign n5276 = ~n5262 & n5275 ;
  assign n5277 = ~n5273 & ~n5276 ;
  assign n5278 = ~n2151 & n3377 ;
  assign n5279 = n2249 & ~n5278 ;
  assign n5280 = ~n3399 & n5279 ;
  assign n5281 = n2181 & n2264 ;
  assign n5282 = n2230 & n5281 ;
  assign n5283 = ~n2146 & ~n2269 ;
  assign n5284 = ~n2151 & ~n5283 ;
  assign n5285 = n5282 & n5284 ;
  assign n5286 = ~n5280 & n5285 ;
  assign n5287 = ~n1437 & n3695 ;
  assign n5288 = n1420 & n5287 ;
  assign n5289 = n1412 & n5288 ;
  assign n5290 = n1382 & n5289 ;
  assign n5291 = ~n3692 & ~n5290 ;
  assign n5292 = n1370 & ~n5290 ;
  assign n5293 = ~n3686 & n5292 ;
  assign n5294 = ~n5291 & ~n5293 ;
  assign n5295 = ~n2470 & n2584 ;
  assign n5296 = n2570 & n5295 ;
  assign n5297 = n3456 & n5296 ;
  assign n5298 = n2547 & n5297 ;
  assign n5299 = n2547 & n5296 ;
  assign n5300 = ~n2725 & n5299 ;
  assign n5301 = ~n2720 & n5300 ;
  assign n5302 = ~n2662 & n5301 ;
  assign n5303 = n2458 & n5302 ;
  assign n5304 = ~n5298 & ~n5303 ;
  assign n5305 = n3630 & n3635 ;
  assign n5306 = ~n3036 & n3638 ;
  assign n5307 = n3632 & n5306 ;
  assign n5308 = n2914 & n5307 ;
  assign n5309 = ~n5305 & ~n5308 ;
  assign n5310 = ~\g1345_reg/NET0131  & \g2599_reg/NET0131  ;
  assign n5311 = \g2612_reg/NET0131  & \g5657_pad  ;
  assign n5312 = n5310 & n5311 ;
  assign n5313 = \g2809_reg/NET0131  & ~n5312 ;
  assign n5314 = \g1024_reg/NET0131  & ~\g2802_reg/NET0131  ;
  assign n5315 = \g1018_reg/NET0131  & ~\g2804_reg/NET0131  ;
  assign n5316 = ~\g2803_reg/NET0131  & \g5657_pad  ;
  assign n5317 = ~n5315 & ~n5316 ;
  assign n5318 = ~n5314 & n5317 ;
  assign n5319 = n1647 & n5318 ;
  assign n5320 = n5312 & n5319 ;
  assign n5321 = ~n5313 & ~n5320 ;
  assign n5322 = ~\g1319_reg/NET0131  & ~n1653 ;
  assign n5323 = \g1339_reg/NET0131  & ~n1596 ;
  assign n5324 = n1599 & n5323 ;
  assign n5325 = ~n5322 & ~n5324 ;
  assign n5326 = ~\g1378_reg/NET0131  & ~n1658 ;
  assign n5327 = ~\g1332_reg/NET0131  & ~n1629 ;
  assign n5328 = ~n5326 & ~n5327 ;
  assign n5329 = n5325 & n5328 ;
  assign n5330 = ~\g1346_reg/NET0131  & ~n1616 ;
  assign n5331 = ~\g1352_reg/NET0131  & ~n1605 ;
  assign n5332 = ~n5330 & ~n5331 ;
  assign n5333 = \g1352_reg/NET0131  & ~n1601 ;
  assign n5334 = n1604 & n5333 ;
  assign n5335 = ~\g1372_reg/NET0131  & ~n1594 ;
  assign n5336 = ~n5334 & ~n5335 ;
  assign n5337 = n5332 & n5336 ;
  assign n5338 = n5329 & n5337 ;
  assign n5339 = ~\g1339_reg/NET0131  & ~n1600 ;
  assign n5340 = \g1365_reg/NET0131  & ~n1619 ;
  assign n5341 = n1622 & n5340 ;
  assign n5342 = ~n5339 & ~n5341 ;
  assign n5343 = \g1372_reg/NET0131  & ~n1590 ;
  assign n5344 = n1593 & n5343 ;
  assign n5345 = \g1378_reg/NET0131  & ~n1654 ;
  assign n5346 = n1657 & n5345 ;
  assign n5347 = ~n5344 & ~n5346 ;
  assign n5348 = ~\g1326_reg/NET0131  & ~n1634 ;
  assign n5349 = n5347 & ~n5348 ;
  assign n5350 = n5342 & n5349 ;
  assign n5351 = ~\g1365_reg/NET0131  & ~n1623 ;
  assign n5352 = ~\g1358_reg/NET0131  & ~n1611 ;
  assign n5353 = ~n5351 & ~n5352 ;
  assign n5354 = \g1319_reg/NET0131  & ~n1649 ;
  assign n5355 = n1652 & n5354 ;
  assign n5356 = \g1332_reg/NET0131  & ~n1625 ;
  assign n5357 = n1628 & n5356 ;
  assign n5358 = ~n5355 & ~n5357 ;
  assign n5359 = \g1346_reg/NET0131  & ~n1612 ;
  assign n5360 = n1615 & n5359 ;
  assign n5361 = n5358 & ~n5360 ;
  assign n5362 = n5353 & n5361 ;
  assign n5363 = n5350 & n5362 ;
  assign n5364 = n5338 & n5363 ;
  assign n5365 = \g1358_reg/NET0131  & ~n1607 ;
  assign n5366 = n1610 & n5365 ;
  assign n5367 = \g1326_reg/NET0131  & ~n1630 ;
  assign n5368 = n1633 & n5367 ;
  assign n5369 = ~n5366 & ~n5368 ;
  assign n5370 = ~n5313 & n5369 ;
  assign n5371 = n5364 & n5370 ;
  assign n5372 = ~n5321 & ~n5371 ;
  assign n5373 = \g1018_reg/NET0131  & \g2612_reg/NET0131  ;
  assign n5374 = n5310 & n5373 ;
  assign n5375 = \g2810_reg/NET0131  & ~n5374 ;
  assign n5376 = n5319 & n5374 ;
  assign n5377 = ~n5375 & ~n5376 ;
  assign n5378 = n5369 & ~n5375 ;
  assign n5379 = n5364 & n5378 ;
  assign n5380 = ~n5377 & ~n5379 ;
  assign n5381 = \g1211_reg/NET0131  & \g1224_reg/NET0131  ;
  assign n5382 = \g1024_reg/NET0131  & ~\g1345_reg/NET0131  ;
  assign n5383 = n5381 & n5382 ;
  assign n5384 = \g1420_reg/NET0131  & ~n5383 ;
  assign n5385 = \g1024_reg/NET0131  & ~\g1414_reg/NET0131  ;
  assign n5386 = \g1018_reg/NET0131  & ~\g1416_reg/NET0131  ;
  assign n5387 = ~\g1415_reg/NET0131  & \g5657_pad  ;
  assign n5388 = ~n5386 & ~n5387 ;
  assign n5389 = ~n5385 & n5388 ;
  assign n5390 = n3110 & n5389 ;
  assign n5391 = n5383 & n5390 ;
  assign n5392 = ~n5384 & ~n5391 ;
  assign n5393 = ~\g1346_reg/NET0131  & ~n3133 ;
  assign n5394 = \g1319_reg/NET0131  & ~n3140 ;
  assign n5395 = n3143 & n5394 ;
  assign n5396 = ~n5393 & ~n5395 ;
  assign n5397 = ~\g1332_reg/NET0131  & ~n3156 ;
  assign n5398 = ~\g1358_reg/NET0131  & ~n3121 ;
  assign n5399 = ~n5397 & ~n5398 ;
  assign n5400 = n5396 & n5399 ;
  assign n5401 = ~\g1339_reg/NET0131  & ~n3116 ;
  assign n5402 = ~\g1372_reg/NET0131  & ~n3128 ;
  assign n5403 = ~n5401 & ~n5402 ;
  assign n5404 = \g1372_reg/NET0131  & ~n3124 ;
  assign n5405 = n3127 & n5404 ;
  assign n5406 = ~\g1365_reg/NET0131  & ~n3167 ;
  assign n5407 = ~n5405 & ~n5406 ;
  assign n5408 = n5403 & n5407 ;
  assign n5409 = n5400 & n5408 ;
  assign n5410 = ~\g1319_reg/NET0131  & ~n3144 ;
  assign n5411 = \g1378_reg/NET0131  & ~n3158 ;
  assign n5412 = n3161 & n5411 ;
  assign n5413 = ~n5410 & ~n5412 ;
  assign n5414 = \g1365_reg/NET0131  & ~n3163 ;
  assign n5415 = n3166 & n5414 ;
  assign n5416 = \g1332_reg/NET0131  & ~n3152 ;
  assign n5417 = n3155 & n5416 ;
  assign n5418 = ~n5415 & ~n5417 ;
  assign n5419 = ~\g1326_reg/NET0131  & ~n3139 ;
  assign n5420 = n5418 & ~n5419 ;
  assign n5421 = n5413 & n5420 ;
  assign n5422 = ~\g1378_reg/NET0131  & ~n3162 ;
  assign n5423 = ~\g1352_reg/NET0131  & ~n3151 ;
  assign n5424 = ~n5422 & ~n5423 ;
  assign n5425 = \g1346_reg/NET0131  & ~n3129 ;
  assign n5426 = n3132 & n5425 ;
  assign n5427 = \g1358_reg/NET0131  & ~n3117 ;
  assign n5428 = n3120 & n5427 ;
  assign n5429 = ~n5426 & ~n5428 ;
  assign n5430 = \g1339_reg/NET0131  & ~n3112 ;
  assign n5431 = n3115 & n5430 ;
  assign n5432 = n5429 & ~n5431 ;
  assign n5433 = n5424 & n5432 ;
  assign n5434 = n5421 & n5433 ;
  assign n5435 = n5409 & n5434 ;
  assign n5436 = \g1352_reg/NET0131  & ~n3147 ;
  assign n5437 = n3150 & n5436 ;
  assign n5438 = \g1326_reg/NET0131  & ~n3135 ;
  assign n5439 = n3138 & n5438 ;
  assign n5440 = ~n5437 & ~n5439 ;
  assign n5441 = ~n5384 & n5440 ;
  assign n5442 = n5435 & n5441 ;
  assign n5443 = ~n5392 & ~n5442 ;
  assign n5444 = \g1018_reg/NET0131  & ~\g1345_reg/NET0131  ;
  assign n5445 = n5381 & n5444 ;
  assign n5446 = \g1422_reg/NET0131  & ~n5445 ;
  assign n5447 = n5390 & n5445 ;
  assign n5448 = ~n5446 & ~n5447 ;
  assign n5449 = n5440 & ~n5446 ;
  assign n5450 = n5435 & n5449 ;
  assign n5451 = ~n5448 & ~n5450 ;
  assign n5452 = ~\g1345_reg/NET0131  & \g5657_pad  ;
  assign n5453 = n5381 & n5452 ;
  assign n5454 = \g1421_reg/NET0131  & ~n5453 ;
  assign n5455 = n5390 & n5453 ;
  assign n5456 = ~n5454 & ~n5455 ;
  assign n5457 = n5440 & ~n5454 ;
  assign n5458 = n5435 & n5457 ;
  assign n5459 = ~n5456 & ~n5458 ;
  assign n5460 = ~\g1345_reg/NET0131  & \g1905_reg/NET0131  ;
  assign n5461 = \g1024_reg/NET0131  & \g1918_reg/NET0131  ;
  assign n5462 = n5460 & n5461 ;
  assign n5463 = \g2114_reg/NET0131  & ~n5462 ;
  assign n5464 = \g1024_reg/NET0131  & ~\g2108_reg/NET0131  ;
  assign n5465 = \g1018_reg/NET0131  & ~\g2110_reg/NET0131  ;
  assign n5466 = ~\g2109_reg/NET0131  & \g5657_pad  ;
  assign n5467 = ~n5465 & ~n5466 ;
  assign n5468 = ~n5464 & n5467 ;
  assign n5469 = n1826 & n5468 ;
  assign n5470 = n5462 & n5469 ;
  assign n5471 = ~n5463 & ~n5470 ;
  assign n5472 = ~\g1346_reg/NET0131  & ~n1860 ;
  assign n5473 = \g1319_reg/NET0131  & ~n1868 ;
  assign n5474 = n1871 & n5473 ;
  assign n5475 = ~n5472 & ~n5474 ;
  assign n5476 = ~\g1358_reg/NET0131  & ~n1849 ;
  assign n5477 = ~\g1332_reg/NET0131  & ~n1867 ;
  assign n5478 = ~n5476 & ~n5477 ;
  assign n5479 = n5475 & n5478 ;
  assign n5480 = ~\g1339_reg/NET0131  & ~n1878 ;
  assign n5481 = ~\g1378_reg/NET0131  & ~n1883 ;
  assign n5482 = ~n5480 & ~n5481 ;
  assign n5483 = \g1378_reg/NET0131  & ~n1879 ;
  assign n5484 = n1882 & n5483 ;
  assign n5485 = ~\g1372_reg/NET0131  & ~n1844 ;
  assign n5486 = ~n5484 & ~n5485 ;
  assign n5487 = n5482 & n5486 ;
  assign n5488 = n5479 & n5487 ;
  assign n5489 = ~\g1319_reg/NET0131  & ~n1872 ;
  assign n5490 = \g1352_reg/NET0131  & ~n1828 ;
  assign n5491 = n1831 & n5490 ;
  assign n5492 = ~n5489 & ~n5491 ;
  assign n5493 = \g1372_reg/NET0131  & ~n1840 ;
  assign n5494 = n1843 & n5493 ;
  assign n5495 = \g1358_reg/NET0131  & ~n1845 ;
  assign n5496 = n1848 & n5495 ;
  assign n5497 = ~n5494 & ~n5496 ;
  assign n5498 = ~\g1326_reg/NET0131  & ~n1855 ;
  assign n5499 = n5497 & ~n5498 ;
  assign n5500 = n5492 & n5499 ;
  assign n5501 = ~\g1352_reg/NET0131  & ~n1832 ;
  assign n5502 = ~\g1365_reg/NET0131  & ~n1821 ;
  assign n5503 = ~n5501 & ~n5502 ;
  assign n5504 = \g1346_reg/NET0131  & ~n1856 ;
  assign n5505 = n1859 & n5504 ;
  assign n5506 = \g1332_reg/NET0131  & ~n1863 ;
  assign n5507 = n1866 & n5506 ;
  assign n5508 = ~n5505 & ~n5507 ;
  assign n5509 = \g1339_reg/NET0131  & ~n1874 ;
  assign n5510 = n1877 & n5509 ;
  assign n5511 = n5508 & ~n5510 ;
  assign n5512 = n5503 & n5511 ;
  assign n5513 = n5500 & n5512 ;
  assign n5514 = n5488 & n5513 ;
  assign n5515 = \g1365_reg/NET0131  & ~n1817 ;
  assign n5516 = n1820 & n5515 ;
  assign n5517 = \g1326_reg/NET0131  & ~n1851 ;
  assign n5518 = n1854 & n5517 ;
  assign n5519 = ~n5516 & ~n5518 ;
  assign n5520 = ~n5463 & n5519 ;
  assign n5521 = n5514 & n5520 ;
  assign n5522 = ~n5471 & ~n5521 ;
  assign n5523 = ~\g1345_reg/NET0131  & \g525_reg/NET0131  ;
  assign n5524 = \g1024_reg/NET0131  & \g538_reg/NET0131  ;
  assign n5525 = n5523 & n5524 ;
  assign n5526 = \g734_reg/NET0131  & ~n5525 ;
  assign n5527 = \g1024_reg/NET0131  & ~\g728_reg/NET0131  ;
  assign n5528 = \g1018_reg/NET0131  & ~\g730_reg/NET0131  ;
  assign n5529 = \g5657_pad  & ~\g729_reg/NET0131  ;
  assign n5530 = ~n5528 & ~n5529 ;
  assign n5531 = ~n5527 & n5530 ;
  assign n5532 = n4292 & n5531 ;
  assign n5533 = n5525 & n5532 ;
  assign n5534 = ~n5526 & ~n5533 ;
  assign n5535 = ~\g1326_reg/NET0131  & ~n4280 ;
  assign n5536 = \g1319_reg/NET0131  & ~n4265 ;
  assign n5537 = n4268 & n5536 ;
  assign n5538 = ~n5535 & ~n5537 ;
  assign n5539 = ~\g1358_reg/NET0131  & ~n4246 ;
  assign n5540 = ~\g1352_reg/NET0131  & ~n4303 ;
  assign n5541 = ~n5539 & ~n5540 ;
  assign n5542 = n5538 & n5541 ;
  assign n5543 = ~\g1339_reg/NET0131  & ~n4241 ;
  assign n5544 = ~\g1378_reg/NET0131  & ~n4287 ;
  assign n5545 = ~n5543 & ~n5544 ;
  assign n5546 = \g1378_reg/NET0131  & ~n4283 ;
  assign n5547 = n4286 & n5546 ;
  assign n5548 = ~\g1372_reg/NET0131  & ~n4264 ;
  assign n5549 = ~n5547 & ~n5548 ;
  assign n5550 = n5545 & n5549 ;
  assign n5551 = n5542 & n5550 ;
  assign n5552 = ~\g1319_reg/NET0131  & ~n4269 ;
  assign n5553 = \g1332_reg/NET0131  & ~n4271 ;
  assign n5554 = n4274 & n5553 ;
  assign n5555 = ~n5552 & ~n5554 ;
  assign n5556 = \g1372_reg/NET0131  & ~n4260 ;
  assign n5557 = n4263 & n5556 ;
  assign n5558 = \g1358_reg/NET0131  & ~n4242 ;
  assign n5559 = n4245 & n5558 ;
  assign n5560 = ~n5557 & ~n5559 ;
  assign n5561 = ~\g1346_reg/NET0131  & ~n4298 ;
  assign n5562 = n5560 & ~n5561 ;
  assign n5563 = n5555 & n5562 ;
  assign n5564 = ~\g1332_reg/NET0131  & ~n4275 ;
  assign n5565 = ~\g1365_reg/NET0131  & ~n4252 ;
  assign n5566 = ~n5564 & ~n5565 ;
  assign n5567 = \g1326_reg/NET0131  & ~n4276 ;
  assign n5568 = n4279 & n5567 ;
  assign n5569 = \g1352_reg/NET0131  & ~n4299 ;
  assign n5570 = n4302 & n5569 ;
  assign n5571 = ~n5568 & ~n5570 ;
  assign n5572 = \g1339_reg/NET0131  & ~n4237 ;
  assign n5573 = n4240 & n5572 ;
  assign n5574 = n5571 & ~n5573 ;
  assign n5575 = n5566 & n5574 ;
  assign n5576 = n5563 & n5575 ;
  assign n5577 = n5551 & n5576 ;
  assign n5578 = \g1365_reg/NET0131  & ~n4248 ;
  assign n5579 = n4251 & n5578 ;
  assign n5580 = \g1346_reg/NET0131  & ~n4294 ;
  assign n5581 = n4297 & n5580 ;
  assign n5582 = ~n5579 & ~n5581 ;
  assign n5583 = ~n5526 & n5582 ;
  assign n5584 = n5577 & n5583 ;
  assign n5585 = ~n5534 & ~n5584 ;
  assign n5586 = \g525_reg/NET0131  & \g538_reg/NET0131  ;
  assign n5587 = n5452 & n5586 ;
  assign n5588 = \g735_reg/NET0131  & ~n5587 ;
  assign n5589 = n5532 & n5587 ;
  assign n5590 = ~n5588 & ~n5589 ;
  assign n5591 = n5582 & ~n5588 ;
  assign n5592 = n5577 & n5591 ;
  assign n5593 = ~n5590 & ~n5592 ;
  assign n5594 = \g1018_reg/NET0131  & \g538_reg/NET0131  ;
  assign n5595 = n5523 & n5594 ;
  assign n5596 = \g736_reg/NET0131  & ~n5595 ;
  assign n5597 = n5532 & n5595 ;
  assign n5598 = ~n5596 & ~n5597 ;
  assign n5599 = n5582 & ~n5596 ;
  assign n5600 = n5577 & n5599 ;
  assign n5601 = ~n5598 & ~n5600 ;
  assign n5602 = \g1018_reg/NET0131  & \g1918_reg/NET0131  ;
  assign n5603 = n5460 & n5602 ;
  assign n5604 = \g2116_reg/NET0131  & ~n5603 ;
  assign n5605 = n5469 & n5603 ;
  assign n5606 = ~n5604 & ~n5605 ;
  assign n5607 = n5519 & ~n5604 ;
  assign n5608 = n5514 & n5607 ;
  assign n5609 = ~n5606 & ~n5608 ;
  assign n5610 = \g1905_reg/NET0131  & \g1918_reg/NET0131  ;
  assign n5611 = n5452 & n5610 ;
  assign n5612 = \g2115_reg/NET0131  & ~n5611 ;
  assign n5613 = n5469 & n5611 ;
  assign n5614 = ~n5612 & ~n5613 ;
  assign n5615 = n5519 & ~n5612 ;
  assign n5616 = n5514 & n5615 ;
  assign n5617 = ~n5614 & ~n5616 ;
  assign n5618 = \g1024_reg/NET0131  & \g2612_reg/NET0131  ;
  assign n5619 = n5310 & n5618 ;
  assign n5620 = \g2808_reg/NET0131  & ~n5619 ;
  assign n5621 = n5319 & n5619 ;
  assign n5622 = ~n5620 & ~n5621 ;
  assign n5623 = n5369 & ~n5620 ;
  assign n5624 = n5364 & n5623 ;
  assign n5625 = ~n5622 & ~n5624 ;
  assign n5626 = ~n1905 & ~n5059 ;
  assign n5627 = \g1018_reg/NET0131  & \g1747_reg/NET0131  ;
  assign n5628 = \g1745_reg/NET0131  & \g5657_pad  ;
  assign n5629 = \g1024_reg/NET0131  & \g1749_reg/NET0131  ;
  assign n5630 = ~n5628 & ~n5629 ;
  assign n5631 = ~n5627 & n5630 ;
  assign n5632 = \g1018_reg/NET0131  & \g1762_reg/NET0131  ;
  assign n5633 = \g1760_reg/NET0131  & \g5657_pad  ;
  assign n5634 = \g1024_reg/NET0131  & \g1764_reg/NET0131  ;
  assign n5635 = ~n5633 & ~n5634 ;
  assign n5636 = ~n5632 & n5635 ;
  assign n5637 = \g1018_reg/NET0131  & \g1732_reg/NET0131  ;
  assign n5638 = \g1730_reg/NET0131  & \g5657_pad  ;
  assign n5639 = \g1024_reg/NET0131  & \g1734_reg/NET0131  ;
  assign n5640 = ~n5638 & ~n5639 ;
  assign n5641 = ~n5637 & n5640 ;
  assign n5642 = n5636 & n5641 ;
  assign n5643 = ~\g1959_reg/NET0131  & \g5657_pad  ;
  assign n5644 = \g1018_reg/NET0131  & ~\g1960_reg/NET0131  ;
  assign n5645 = \g1024_reg/NET0131  & ~\g1958_reg/NET0131  ;
  assign n5646 = ~n5644 & ~n5645 ;
  assign n5647 = ~n5643 & n5646 ;
  assign n5648 = \g1024_reg/NET0131  & ~\g1961_reg/NET0131  ;
  assign n5649 = \g1018_reg/NET0131  & ~\g1963_reg/NET0131  ;
  assign n5650 = ~\g1962_reg/NET0131  & \g5657_pad  ;
  assign n5651 = ~n5649 & ~n5650 ;
  assign n5652 = ~n5648 & n5651 ;
  assign n5653 = n5647 & n5652 ;
  assign n5654 = n5642 & n5653 ;
  assign n5655 = n5636 & ~n5641 ;
  assign n5656 = ~n5647 & n5655 ;
  assign n5657 = ~\g1956_reg/NET0131  & \g5657_pad  ;
  assign n5658 = \g1018_reg/NET0131  & ~\g1957_reg/NET0131  ;
  assign n5659 = \g1024_reg/NET0131  & ~\g1955_reg/NET0131  ;
  assign n5660 = ~n5658 & ~n5659 ;
  assign n5661 = ~n5657 & n5660 ;
  assign n5662 = ~n5652 & n5661 ;
  assign n5663 = ~n5636 & ~n5641 ;
  assign n5664 = n5662 & n5663 ;
  assign n5665 = ~n5656 & ~n5664 ;
  assign n5666 = ~n5654 & n5665 ;
  assign n5667 = ~n5631 & ~n5666 ;
  assign n5668 = n5647 & n5661 ;
  assign n5669 = ~n5631 & ~n5636 ;
  assign n5670 = n5641 & n5669 ;
  assign n5671 = n5668 & n5670 ;
  assign n5672 = \g1018_reg/NET0131  & \g1777_reg/NET0131  ;
  assign n5673 = \g1775_reg/NET0131  & \g5657_pad  ;
  assign n5674 = \g1024_reg/NET0131  & \g1705_reg/NET0131  ;
  assign n5675 = ~n5673 & ~n5674 ;
  assign n5676 = ~n5672 & n5675 ;
  assign n5677 = ~n5631 & ~n5676 ;
  assign n5678 = ~n5636 & ~n5677 ;
  assign n5679 = ~n5647 & n5652 ;
  assign n5680 = ~n5641 & n5679 ;
  assign n5681 = ~n5678 & n5680 ;
  assign n5682 = ~n5671 & ~n5681 ;
  assign n5683 = n5662 & n5676 ;
  assign n5684 = ~n5641 & n5661 ;
  assign n5685 = \g1024_reg/NET0131  & ~\g1964_reg/NET0131  ;
  assign n5686 = \g1018_reg/NET0131  & ~\g1966_reg/NET0131  ;
  assign n5687 = ~\g1965_reg/NET0131  & \g5657_pad  ;
  assign n5688 = ~n5686 & ~n5687 ;
  assign n5689 = ~n5685 & n5688 ;
  assign n5690 = n5676 & n5689 ;
  assign n5691 = n5684 & n5690 ;
  assign n5692 = ~n5683 & ~n5691 ;
  assign n5693 = n5642 & ~n5689 ;
  assign n5694 = n5631 & n5641 ;
  assign n5695 = n5647 & ~n5661 ;
  assign n5696 = n5694 & n5695 ;
  assign n5697 = ~n5693 & ~n5696 ;
  assign n5698 = n5692 & n5697 ;
  assign n5699 = n5682 & n5698 ;
  assign n5700 = ~n5667 & n5699 ;
  assign n5701 = ~n5642 & ~n5652 ;
  assign n5702 = n5663 & n5689 ;
  assign n5703 = ~n5701 & ~n5702 ;
  assign n5704 = n5631 & ~n5661 ;
  assign n5705 = ~n5703 & n5704 ;
  assign n5706 = ~n5676 & ~n5689 ;
  assign n5707 = n5641 & ~n5661 ;
  assign n5708 = n5706 & n5707 ;
  assign n5709 = \g1018_reg/NET0131  & \g1947_reg/NET0131  ;
  assign n5710 = \g1945_reg/NET0131  & \g5657_pad  ;
  assign n5711 = \g1024_reg/NET0131  & \g1870_reg/NET0131  ;
  assign n5712 = ~n5710 & ~n5711 ;
  assign n5713 = ~n5709 & n5712 ;
  assign n5714 = \g185_reg/NET0131  & \g1922_reg/NET0131  ;
  assign n5715 = ~n5713 & n5714 ;
  assign n5716 = \g1018_reg/NET0131  & \g1979_reg/NET0131  ;
  assign n5717 = \g1976_reg/NET0131  & \g5657_pad  ;
  assign n5718 = \g1024_reg/NET0131  & \g1982_reg/NET0131  ;
  assign n5719 = ~n5717 & ~n5718 ;
  assign n5720 = ~n5716 & n5719 ;
  assign n5721 = ~n5715 & n5720 ;
  assign n5722 = ~n5708 & n5721 ;
  assign n5723 = ~n5705 & n5722 ;
  assign n5724 = n5700 & n5723 ;
  assign n5725 = n5689 & n5695 ;
  assign n5726 = n5670 & n5725 ;
  assign n5727 = n5655 & n5689 ;
  assign n5728 = n5668 & n5727 ;
  assign n5729 = n5652 & n5676 ;
  assign n5730 = n5695 & n5729 ;
  assign n5731 = ~n5647 & ~n5661 ;
  assign n5732 = n5642 & n5731 ;
  assign n5733 = ~n5730 & ~n5732 ;
  assign n5734 = ~n5728 & n5733 ;
  assign n5735 = ~n5726 & n5734 ;
  assign n5736 = ~n5652 & ~n5661 ;
  assign n5737 = ~n5684 & ~n5736 ;
  assign n5738 = ~n5641 & ~n5653 ;
  assign n5739 = ~n5737 & ~n5738 ;
  assign n5740 = n5677 & n5739 ;
  assign n5741 = n5679 & n5694 ;
  assign n5742 = n5631 & ~n5641 ;
  assign n5743 = n5662 & n5742 ;
  assign n5744 = ~n5741 & ~n5743 ;
  assign n5745 = ~n5647 & n5661 ;
  assign n5746 = n5631 & ~n5636 ;
  assign n5747 = n5745 & n5746 ;
  assign n5748 = ~n5641 & ~n5689 ;
  assign n5749 = n5669 & n5748 ;
  assign n5750 = ~n5747 & ~n5749 ;
  assign n5751 = n5744 & n5750 ;
  assign n5752 = ~n5740 & n5751 ;
  assign n5753 = n5735 & n5752 ;
  assign n5754 = \g1949_reg/NET0131  & \g5657_pad  ;
  assign n5755 = \g1018_reg/NET0131  & \g1951_reg/NET0131  ;
  assign n5756 = \g1024_reg/NET0131  & \g1953_reg/NET0131  ;
  assign n5757 = ~n5755 & ~n5756 ;
  assign n5758 = ~n5754 & n5757 ;
  assign n5759 = \g185_reg/NET0131  & \g1904_reg/NET0131  ;
  assign n5760 = ~n5758 & n5759 ;
  assign n5761 = \g1024_reg/NET0131  & \g1973_reg/NET0131  ;
  assign n5762 = \g1967_reg/NET0131  & \g5657_pad  ;
  assign n5763 = \g1018_reg/NET0131  & \g1970_reg/NET0131  ;
  assign n5764 = ~n5762 & ~n5763 ;
  assign n5765 = ~n5761 & n5764 ;
  assign n5766 = ~n5760 & n5765 ;
  assign n5767 = ~n5721 & ~n5766 ;
  assign n5768 = n5059 & ~n5767 ;
  assign n5769 = n5753 & n5768 ;
  assign n5770 = ~n5724 & n5769 ;
  assign n5771 = ~n5626 & ~n5770 ;
  assign n5772 = ~n4325 & ~n5059 ;
  assign n5773 = \g5657_pad  & ~\g576_reg/NET0131  ;
  assign n5774 = \g1024_reg/NET0131  & ~\g575_reg/NET0131  ;
  assign n5775 = \g1018_reg/NET0131  & ~\g577_reg/NET0131  ;
  assign n5776 = ~n5774 & ~n5775 ;
  assign n5777 = ~n5773 & n5776 ;
  assign n5778 = \g1024_reg/NET0131  & ~\g578_reg/NET0131  ;
  assign n5779 = \g1018_reg/NET0131  & ~\g580_reg/NET0131  ;
  assign n5780 = \g5657_pad  & ~\g579_reg/NET0131  ;
  assign n5781 = ~n5779 & ~n5780 ;
  assign n5782 = ~n5778 & n5781 ;
  assign n5783 = ~n5777 & n5782 ;
  assign n5784 = \g1018_reg/NET0131  & \g366_reg/NET0131  ;
  assign n5785 = \g364_reg/NET0131  & \g5657_pad  ;
  assign n5786 = \g1024_reg/NET0131  & \g368_reg/NET0131  ;
  assign n5787 = ~n5785 & ~n5786 ;
  assign n5788 = ~n5784 & n5787 ;
  assign n5789 = \g1018_reg/NET0131  & \g351_reg/NET0131  ;
  assign n5790 = \g349_reg/NET0131  & \g5657_pad  ;
  assign n5791 = \g1024_reg/NET0131  & \g353_reg/NET0131  ;
  assign n5792 = ~n5790 & ~n5791 ;
  assign n5793 = ~n5789 & n5792 ;
  assign n5794 = n5788 & n5793 ;
  assign n5795 = n5783 & n5794 ;
  assign n5796 = n5788 & ~n5793 ;
  assign n5797 = \g1024_reg/NET0131  & ~\g581_reg/NET0131  ;
  assign n5798 = \g1018_reg/NET0131  & ~\g583_reg/NET0131  ;
  assign n5799 = \g5657_pad  & ~\g582_reg/NET0131  ;
  assign n5800 = ~n5798 & ~n5799 ;
  assign n5801 = ~n5797 & n5800 ;
  assign n5802 = ~n5777 & ~n5801 ;
  assign n5803 = n5796 & n5802 ;
  assign n5804 = ~n5795 & ~n5803 ;
  assign n5805 = \g1018_reg/NET0131  & \g381_reg/NET0131  ;
  assign n5806 = \g379_reg/NET0131  & \g5657_pad  ;
  assign n5807 = \g1024_reg/NET0131  & \g383_reg/NET0131  ;
  assign n5808 = ~n5806 & ~n5807 ;
  assign n5809 = ~n5805 & n5808 ;
  assign n5810 = ~n5782 & n5809 ;
  assign n5811 = ~n5788 & ~n5793 ;
  assign n5812 = n5810 & n5811 ;
  assign n5813 = \g5657_pad  & ~\g585_reg/NET0131  ;
  assign n5814 = \g1018_reg/NET0131  & ~\g586_reg/NET0131  ;
  assign n5815 = \g1024_reg/NET0131  & ~\g584_reg/NET0131  ;
  assign n5816 = ~n5814 & ~n5815 ;
  assign n5817 = ~n5813 & n5816 ;
  assign n5818 = ~n5793 & n5817 ;
  assign n5819 = \g1018_reg/NET0131  & \g396_reg/NET0131  ;
  assign n5820 = \g394_reg/NET0131  & \g5657_pad  ;
  assign n5821 = \g1024_reg/NET0131  & \g324_reg/NET0131  ;
  assign n5822 = ~n5820 & ~n5821 ;
  assign n5823 = ~n5819 & n5822 ;
  assign n5824 = n5777 & n5823 ;
  assign n5825 = n5818 & n5824 ;
  assign n5826 = ~n5812 & ~n5825 ;
  assign n5827 = n5804 & n5826 ;
  assign n5828 = n5801 & ~n5818 ;
  assign n5829 = n5788 & ~n5809 ;
  assign n5830 = ~n5777 & n5829 ;
  assign n5831 = ~n5828 & n5830 ;
  assign n5832 = n5777 & n5782 ;
  assign n5833 = ~n5788 & n5793 ;
  assign n5834 = ~n5809 & n5833 ;
  assign n5835 = n5832 & n5834 ;
  assign n5836 = ~n5831 & ~n5835 ;
  assign n5837 = n5827 & n5836 ;
  assign n5838 = n5777 & ~n5801 ;
  assign n5839 = ~n5809 & n5811 ;
  assign n5840 = ~n5823 & ~n5839 ;
  assign n5841 = n5838 & ~n5840 ;
  assign n5842 = ~n5782 & n5801 ;
  assign n5843 = ~n5793 & n5809 ;
  assign n5844 = n5811 & ~n5823 ;
  assign n5845 = ~n5843 & ~n5844 ;
  assign n5846 = n5842 & ~n5845 ;
  assign n5847 = ~n5841 & ~n5846 ;
  assign n5848 = n5837 & n5847 ;
  assign n5849 = \g1018_reg/NET0131  & \g567_reg/NET0131  ;
  assign n5850 = \g5657_pad  & \g565_reg/NET0131  ;
  assign n5851 = \g1024_reg/NET0131  & \g489_reg/NET0131  ;
  assign n5852 = ~n5850 & ~n5851 ;
  assign n5853 = ~n5849 & n5852 ;
  assign n5854 = \g185_reg/NET0131  & \g542_reg/NET0131  ;
  assign n5855 = ~n5853 & n5854 ;
  assign n5856 = \g1024_reg/NET0131  & \g602_reg/NET0131  ;
  assign n5857 = \g5657_pad  & \g596_reg/NET0131  ;
  assign n5858 = \g1018_reg/NET0131  & \g599_reg/NET0131  ;
  assign n5859 = ~n5857 & ~n5858 ;
  assign n5860 = ~n5856 & n5859 ;
  assign n5861 = ~n5855 & n5860 ;
  assign n5862 = ~n5788 & n5809 ;
  assign n5863 = n5782 & n5801 ;
  assign n5864 = n5862 & n5863 ;
  assign n5865 = n5793 & n5864 ;
  assign n5866 = ~n5777 & ~n5823 ;
  assign n5867 = ~n5809 & ~n5866 ;
  assign n5868 = n5793 & ~n5817 ;
  assign n5869 = ~n5867 & n5868 ;
  assign n5870 = ~n5865 & ~n5869 ;
  assign n5871 = n5861 & n5870 ;
  assign n5872 = n5848 & n5871 ;
  assign n5873 = n5796 & n5838 ;
  assign n5874 = n5777 & ~n5782 ;
  assign n5875 = n5829 & n5874 ;
  assign n5876 = ~n5873 & ~n5875 ;
  assign n5877 = ~n5809 & n5817 ;
  assign n5878 = n5833 & n5877 ;
  assign n5879 = n5783 & n5878 ;
  assign n5880 = n5802 & ~n5823 ;
  assign n5881 = n5833 & n5880 ;
  assign n5882 = ~n5879 & ~n5881 ;
  assign n5883 = n5832 & n5843 ;
  assign n5884 = n5817 & n5883 ;
  assign n5885 = ~n5777 & n5793 ;
  assign n5886 = n5810 & n5885 ;
  assign n5887 = ~n5809 & ~n5817 ;
  assign n5888 = n5811 & n5887 ;
  assign n5889 = ~n5886 & ~n5888 ;
  assign n5890 = ~n5884 & n5889 ;
  assign n5891 = n5882 & n5890 ;
  assign n5892 = n5876 & n5891 ;
  assign n5893 = n5832 & n5844 ;
  assign n5894 = ~n5782 & n5794 ;
  assign n5895 = n5783 & n5823 ;
  assign n5896 = ~n5894 & ~n5895 ;
  assign n5897 = ~n5893 & n5896 ;
  assign n5898 = n5801 & ~n5897 ;
  assign n5899 = \g5657_pad  & \g569_reg/NET0131  ;
  assign n5900 = \g1018_reg/NET0131  & \g571_reg/NET0131  ;
  assign n5901 = \g1024_reg/NET0131  & \g573_reg/NET0131  ;
  assign n5902 = ~n5900 & ~n5901 ;
  assign n5903 = ~n5899 & n5902 ;
  assign n5904 = \g185_reg/NET0131  & \g524_reg/NET0131  ;
  assign n5905 = ~n5903 & n5904 ;
  assign n5906 = \g1018_reg/NET0131  & \g590_reg/NET0131  ;
  assign n5907 = \g5657_pad  & \g587_reg/NET0131  ;
  assign n5908 = \g1024_reg/NET0131  & \g593_reg/NET0131  ;
  assign n5909 = ~n5907 & ~n5908 ;
  assign n5910 = ~n5906 & n5909 ;
  assign n5911 = ~n5905 & n5910 ;
  assign n5912 = ~n5861 & ~n5911 ;
  assign n5913 = n5059 & ~n5912 ;
  assign n5914 = ~n5898 & n5913 ;
  assign n5915 = n5892 & n5914 ;
  assign n5916 = ~n5872 & n5915 ;
  assign n5917 = ~n5772 & ~n5916 ;
  assign n5918 = n3176 & ~n5059 ;
  assign n5919 = ~n5045 & n5059 ;
  assign n5920 = ~n5918 & ~n5919 ;
  assign n5921 = ~\g1092_reg/NET0131  & \g299_reg/NET0131  ;
  assign n5922 = \g305_reg/NET0131  & n5921 ;
  assign n5923 = ~n2127 & ~n5922 ;
  assign n5924 = ~n1892 & ~n5059 ;
  assign n5925 = ~n5726 & n5766 ;
  assign n5926 = n5734 & n5925 ;
  assign n5927 = n5752 & n5926 ;
  assign n5928 = n5059 & ~n5708 ;
  assign n5929 = ~n5767 & n5928 ;
  assign n5930 = ~n5705 & n5929 ;
  assign n5931 = n5700 & n5930 ;
  assign n5932 = ~n5927 & n5931 ;
  assign n5933 = ~n5924 & ~n5932 ;
  assign n5934 = ~n3188 & ~n5059 ;
  assign n5935 = n5025 & ~n5027 ;
  assign n5936 = ~n5008 & n5040 ;
  assign n5937 = ~n5006 & n5936 ;
  assign n5938 = n5019 & n5937 ;
  assign n5939 = n5935 & n5938 ;
  assign n5940 = ~n5041 & n5059 ;
  assign n5941 = ~n5000 & n5940 ;
  assign n5942 = n4969 & n5941 ;
  assign n5943 = ~n5939 & n5942 ;
  assign n5944 = ~n5934 & ~n5943 ;
  assign n5945 = ~n4312 & ~n5059 ;
  assign n5946 = ~n5898 & n5911 ;
  assign n5947 = n5892 & n5946 ;
  assign n5948 = n5870 & n5913 ;
  assign n5949 = n5848 & n5948 ;
  assign n5950 = ~n5947 & n5949 ;
  assign n5951 = ~n5945 & ~n5950 ;
  assign n5952 = \g1088_reg/NET0131  & \g1563_reg/NET0131  ;
  assign n5953 = n2248 & ~n5278 ;
  assign n5954 = n2316 & ~n5278 ;
  assign n5955 = n2375 & n5954 ;
  assign n5956 = ~n5953 & ~n5955 ;
  assign n5957 = n5952 & n5956 ;
  assign n5958 = \g1563_reg/NET0131  & \g7961_pad  ;
  assign n5959 = n5956 & n5958 ;
  assign n5960 = \g1092_reg/NET0131  & \g1563_reg/NET0131  ;
  assign n5961 = n5956 & n5960 ;
  assign n5962 = n1260 & ~n5287 ;
  assign n5963 = n1304 & n5962 ;
  assign n5964 = n1312 & ~n5287 ;
  assign n5965 = n5952 & ~n5964 ;
  assign n5966 = ~n5963 & n5965 ;
  assign n5967 = n5958 & ~n5964 ;
  assign n5968 = ~n5963 & n5967 ;
  assign n5969 = n5960 & ~n5964 ;
  assign n5970 = ~n5963 & n5969 ;
  assign n5971 = ~n2470 & n3456 ;
  assign n5972 = n2656 & ~n5971 ;
  assign n5973 = n2730 & n5972 ;
  assign n5974 = n2733 & n5973 ;
  assign n5975 = n2540 & ~n5971 ;
  assign n5976 = n5952 & ~n5975 ;
  assign n5977 = ~n5974 & n5976 ;
  assign n5978 = n5958 & ~n5975 ;
  assign n5979 = ~n5974 & n5978 ;
  assign n5980 = n5960 & ~n5975 ;
  assign n5981 = ~n5974 & n5980 ;
  assign n5982 = n2779 & ~n5306 ;
  assign n5983 = n3025 & ~n5306 ;
  assign n5984 = n3023 & n5983 ;
  assign n5985 = ~n5982 & ~n5984 ;
  assign n5986 = n5952 & n5985 ;
  assign n5987 = n5958 & n5985 ;
  assign n5988 = n5960 & n5985 ;
  assign n5989 = ~\g1018_reg/NET0131  & \g16355_pad  ;
  assign n5990 = ~\g1192_reg/NET0131  & ~n5989 ;
  assign n5991 = \g1018_reg/NET0131  & ~n4501 ;
  assign n5992 = n5990 & ~n5991 ;
  assign n5993 = ~n4499 & ~n5992 ;
  assign n5994 = \g1332_reg/NET0131  & \g1346_reg/NET0131  ;
  assign n5995 = \g1339_reg/NET0131  & n5994 ;
  assign n5996 = \g1319_reg/NET0131  & \g1326_reg/NET0131  ;
  assign n5997 = n5382 & n5996 ;
  assign n5998 = n5995 & n5997 ;
  assign n5999 = \g1352_reg/NET0131  & \g1365_reg/NET0131  ;
  assign n6000 = \g1358_reg/NET0131  & n5999 ;
  assign n6001 = \g1372_reg/NET0131  & \g1378_reg/NET0131  ;
  assign n6002 = n6000 & n6001 ;
  assign n6003 = n5998 & n6002 ;
  assign n6004 = \g1018_reg/NET0131  & \g1316_reg/NET0131  ;
  assign n6005 = \g1378_reg/NET0131  & ~n6004 ;
  assign n6006 = \g1372_reg/NET0131  & ~n6004 ;
  assign n6007 = n6000 & n6006 ;
  assign n6008 = n5998 & n6007 ;
  assign n6009 = ~n6005 & ~n6008 ;
  assign n6010 = ~n6003 & ~n6009 ;
  assign n6011 = \g1092_reg/NET0131  & \g1098_reg/NET0131  ;
  assign n6012 = \g1095_reg/NET0131  & \g7961_pad  ;
  assign n6013 = \g1088_reg/NET0131  & \g1101_reg/NET0131  ;
  assign n6014 = ~n6012 & ~n6013 ;
  assign n6015 = ~n6011 & n6014 ;
  assign n6016 = \g1088_reg/NET0131  & ~\g1113_reg/NET0131  ;
  assign n6017 = ~\g1114_reg/NET0131  & \g7961_pad  ;
  assign n6018 = \g1092_reg/NET0131  & ~\g1115_reg/NET0131  ;
  assign n6019 = ~n6017 & ~n6018 ;
  assign n6020 = ~n6016 & n6019 ;
  assign n6021 = ~n6015 & ~n6020 ;
  assign n6022 = \g1563_reg/NET0131  & n6021 ;
  assign n6023 = \g1092_reg/NET0131  & \g1107_reg/NET0131  ;
  assign n6024 = \g1104_reg/NET0131  & \g7961_pad  ;
  assign n6025 = \g1088_reg/NET0131  & \g1110_reg/NET0131  ;
  assign n6026 = ~n6024 & ~n6025 ;
  assign n6027 = ~n6023 & n6026 ;
  assign n6028 = ~n6022 & ~n6027 ;
  assign n6029 = ~n2540 & ~n6021 ;
  assign n6030 = ~n2515 & ~n2561 ;
  assign n6031 = \g805_reg/NET0131  & \g809_reg/NET0131  ;
  assign n6032 = \g793_reg/NET0131  & \g797_reg/NET0131  ;
  assign n6033 = n6031 & n6032 ;
  assign n6034 = \g801_reg/NET0131  & \g813_reg/NET0131  ;
  assign n6035 = \g785_reg/NET0131  & \g789_reg/NET0131  ;
  assign n6036 = n6034 & n6035 ;
  assign n6037 = n6033 & n6036 ;
  assign n6038 = \g1563_reg/NET0131  & n6037 ;
  assign n6039 = n6030 & n6038 ;
  assign n6040 = ~n6029 & n6039 ;
  assign n6041 = ~n6028 & ~n6040 ;
  assign n6042 = \g1092_reg/NET0131  & \g411_reg/NET0131  ;
  assign n6043 = \g408_reg/NET0131  & \g7961_pad  ;
  assign n6044 = \g1088_reg/NET0131  & \g414_reg/NET0131  ;
  assign n6045 = ~n6043 & ~n6044 ;
  assign n6046 = ~n6042 & n6045 ;
  assign n6047 = \g1088_reg/NET0131  & ~\g426_reg/NET0131  ;
  assign n6048 = ~\g427_reg/NET0131  & \g7961_pad  ;
  assign n6049 = \g1092_reg/NET0131  & ~\g428_reg/NET0131  ;
  assign n6050 = ~n6048 & ~n6049 ;
  assign n6051 = ~n6047 & n6050 ;
  assign n6052 = ~n6046 & ~n6051 ;
  assign n6053 = \g1563_reg/NET0131  & n6052 ;
  assign n6054 = \g1092_reg/NET0131  & \g420_reg/NET0131  ;
  assign n6055 = \g417_reg/NET0131  & \g7961_pad  ;
  assign n6056 = \g1088_reg/NET0131  & \g423_reg/NET0131  ;
  assign n6057 = ~n6055 & ~n6056 ;
  assign n6058 = ~n6054 & n6057 ;
  assign n6059 = ~n6053 & ~n6058 ;
  assign n6060 = ~n2248 & ~n6052 ;
  assign n6061 = ~n2235 & ~n2255 ;
  assign n6062 = \g121_reg/NET0131  & \g97_reg/NET0131  ;
  assign n6063 = \g109_reg/NET0131  & \g117_reg/NET0131  ;
  assign n6064 = n6062 & n6063 ;
  assign n6065 = \g113_reg/NET0131  & \g125_reg/NET0131  ;
  assign n6066 = \g101_reg/NET0131  & \g105_reg/NET0131  ;
  assign n6067 = n6065 & n6066 ;
  assign n6068 = n6064 & n6067 ;
  assign n6069 = \g1563_reg/NET0131  & n6068 ;
  assign n6070 = n6061 & n6069 ;
  assign n6071 = ~n6060 & n6070 ;
  assign n6072 = ~n6059 & ~n6071 ;
  assign n6073 = \g1092_reg/NET0131  & \g2486_reg/NET0131  ;
  assign n6074 = \g2483_reg/NET0131  & \g7961_pad  ;
  assign n6075 = \g1088_reg/NET0131  & \g2489_reg/NET0131  ;
  assign n6076 = ~n6074 & ~n6075 ;
  assign n6077 = ~n6073 & n6076 ;
  assign n6078 = \g1088_reg/NET0131  & ~\g2501_reg/NET0131  ;
  assign n6079 = ~\g2502_reg/NET0131  & \g7961_pad  ;
  assign n6080 = \g1092_reg/NET0131  & ~\g2503_reg/NET0131  ;
  assign n6081 = ~n6079 & ~n6080 ;
  assign n6082 = ~n6078 & n6081 ;
  assign n6083 = ~n6077 & ~n6082 ;
  assign n6084 = \g1563_reg/NET0131  & n6083 ;
  assign n6085 = \g1092_reg/NET0131  & \g2495_reg/NET0131  ;
  assign n6086 = \g2492_reg/NET0131  & \g7961_pad  ;
  assign n6087 = \g1088_reg/NET0131  & \g2498_reg/NET0131  ;
  assign n6088 = ~n6086 & ~n6087 ;
  assign n6089 = ~n6085 & n6088 ;
  assign n6090 = ~n6084 & ~n6089 ;
  assign n6091 = ~n1312 & ~n6083 ;
  assign n6092 = ~n1219 & ~n1274 ;
  assign n6093 = \g2190_reg/NET0131  & \g2195_reg/NET0131  ;
  assign n6094 = \g2175_reg/NET0131  & \g2180_reg/NET0131  ;
  assign n6095 = n6093 & n6094 ;
  assign n6096 = \g2185_reg/NET0131  & \g2200_reg/NET0131  ;
  assign n6097 = \g2165_reg/NET0131  & \g2170_reg/NET0131  ;
  assign n6098 = n6096 & n6097 ;
  assign n6099 = n6095 & n6098 ;
  assign n6100 = \g1563_reg/NET0131  & n6099 ;
  assign n6101 = n6092 & n6100 ;
  assign n6102 = ~n6091 & n6101 ;
  assign n6103 = ~n6090 & ~n6102 ;
  assign n6104 = \g1088_reg/NET0131  & ~\g1807_reg/NET0131  ;
  assign n6105 = ~\g1808_reg/NET0131  & \g7961_pad  ;
  assign n6106 = \g1092_reg/NET0131  & ~\g1809_reg/NET0131  ;
  assign n6107 = ~n6105 & ~n6106 ;
  assign n6108 = ~n6104 & n6107 ;
  assign n6109 = \g1092_reg/NET0131  & \g1792_reg/NET0131  ;
  assign n6110 = \g1789_reg/NET0131  & \g7961_pad  ;
  assign n6111 = \g1088_reg/NET0131  & \g1795_reg/NET0131  ;
  assign n6112 = ~n6110 & ~n6111 ;
  assign n6113 = ~n6109 & n6112 ;
  assign n6114 = ~n6108 & ~n6113 ;
  assign n6115 = \g1563_reg/NET0131  & n6114 ;
  assign n6116 = \g1092_reg/NET0131  & \g1801_reg/NET0131  ;
  assign n6117 = \g1798_reg/NET0131  & \g7961_pad  ;
  assign n6118 = \g1088_reg/NET0131  & \g1804_reg/NET0131  ;
  assign n6119 = ~n6117 & ~n6118 ;
  assign n6120 = ~n6116 & n6119 ;
  assign n6121 = ~n6115 & ~n6120 ;
  assign n6122 = ~n2779 & ~n6114 ;
  assign n6123 = ~n2785 & ~n2928 ;
  assign n6124 = \g1496_reg/NET0131  & \g1501_reg/NET0131  ;
  assign n6125 = \g1481_reg/NET0131  & \g1486_reg/NET0131  ;
  assign n6126 = n6124 & n6125 ;
  assign n6127 = \g1491_reg/NET0131  & \g1506_reg/NET0131  ;
  assign n6128 = \g1471_reg/NET0131  & \g1476_reg/NET0131  ;
  assign n6129 = n6127 & n6128 ;
  assign n6130 = n6126 & n6129 ;
  assign n6131 = \g1563_reg/NET0131  & n6130 ;
  assign n6132 = n6123 & n6131 ;
  assign n6133 = ~n6122 & n6132 ;
  assign n6134 = ~n6121 & ~n6133 ;
  assign n6135 = n2584 & n2596 ;
  assign n6136 = n2570 & n6135 ;
  assign n6137 = n2547 & n6136 ;
  assign n6138 = n2425 & n5282 ;
  assign n6139 = n1420 & n1451 ;
  assign n6140 = n1412 & n6139 ;
  assign n6141 = n1382 & n6140 ;
  assign n6142 = n3063 & n3632 ;
  assign n6143 = n2914 & n6142 ;
  assign n6144 = ~\g1563_reg/NET0131  & ~n6015 ;
  assign n6145 = n6030 & n6037 ;
  assign n6146 = ~n2540 & n6027 ;
  assign n6147 = n6145 & ~n6146 ;
  assign n6148 = \g1563_reg/NET0131  & ~n6027 ;
  assign n6149 = ~n6039 & ~n6148 ;
  assign n6150 = ~n6147 & ~n6149 ;
  assign n6151 = ~n6021 & n6150 ;
  assign n6152 = ~n6144 & ~n6151 ;
  assign n6153 = ~\g1563_reg/NET0131  & ~n6046 ;
  assign n6154 = n6061 & n6068 ;
  assign n6155 = ~n2248 & n6058 ;
  assign n6156 = n6154 & ~n6155 ;
  assign n6157 = \g1563_reg/NET0131  & ~n6058 ;
  assign n6158 = ~n6070 & ~n6157 ;
  assign n6159 = ~n6156 & ~n6158 ;
  assign n6160 = ~n6052 & n6159 ;
  assign n6161 = ~n6153 & ~n6160 ;
  assign n6162 = ~\g1563_reg/NET0131  & ~n6077 ;
  assign n6163 = n6092 & n6099 ;
  assign n6164 = ~n1312 & n6089 ;
  assign n6165 = n6163 & ~n6164 ;
  assign n6166 = \g1563_reg/NET0131  & ~n6089 ;
  assign n6167 = ~n6101 & ~n6166 ;
  assign n6168 = ~n6165 & ~n6167 ;
  assign n6169 = ~n6083 & n6168 ;
  assign n6170 = ~n6162 & ~n6169 ;
  assign n6171 = ~\g1563_reg/NET0131  & ~n6113 ;
  assign n6172 = n6123 & n6130 ;
  assign n6173 = ~n2779 & n6120 ;
  assign n6174 = n6172 & ~n6173 ;
  assign n6175 = \g1563_reg/NET0131  & ~n6120 ;
  assign n6176 = ~n6132 & ~n6175 ;
  assign n6177 = ~n6174 & ~n6176 ;
  assign n6178 = ~n6114 & n6177 ;
  assign n6179 = ~n6171 & ~n6178 ;
  assign n6180 = ~n5059 & ~n5766 ;
  assign n6181 = ~n5059 & ~n5721 ;
  assign n6182 = ~n5059 & ~n5911 ;
  assign n6183 = ~n5059 & ~n5861 ;
  assign n6184 = ~n5040 & ~n5059 ;
  assign n6185 = ~n4982 & ~n5059 ;
  assign n6186 = ~n5059 & ~n5203 ;
  assign n6187 = ~n5059 & ~n5160 ;
  assign n6188 = n5998 & n6000 ;
  assign n6189 = n6006 & ~n6188 ;
  assign n6190 = ~\g1372_reg/NET0131  & ~n6004 ;
  assign n6191 = n6000 & n6190 ;
  assign n6192 = n5998 & n6191 ;
  assign n6193 = ~n6189 & ~n6192 ;
  assign n6194 = ~n1480 & n1492 ;
  assign n6195 = n1489 & ~n6194 ;
  assign n6196 = \g1088_reg/NET0131  & ~n6021 ;
  assign n6197 = n6150 & n6196 ;
  assign n6198 = \g7961_pad  & ~n6021 ;
  assign n6199 = n6150 & n6198 ;
  assign n6200 = \g1092_reg/NET0131  & ~n6021 ;
  assign n6201 = n6150 & n6200 ;
  assign n6202 = \g1088_reg/NET0131  & ~n6052 ;
  assign n6203 = n6159 & n6202 ;
  assign n6204 = \g7961_pad  & ~n6052 ;
  assign n6205 = n6159 & n6204 ;
  assign n6206 = \g1092_reg/NET0131  & ~n6052 ;
  assign n6207 = n6159 & n6206 ;
  assign n6208 = \g1088_reg/NET0131  & ~n6083 ;
  assign n6209 = n6168 & n6208 ;
  assign n6210 = \g7961_pad  & ~n6083 ;
  assign n6211 = n6168 & n6210 ;
  assign n6212 = \g1092_reg/NET0131  & ~n6083 ;
  assign n6213 = n6168 & n6212 ;
  assign n6214 = \g1088_reg/NET0131  & ~n6114 ;
  assign n6215 = n6177 & n6214 ;
  assign n6216 = \g7961_pad  & ~n6114 ;
  assign n6217 = n6177 & n6216 ;
  assign n6218 = \g1092_reg/NET0131  & ~n6114 ;
  assign n6219 = n6177 & n6218 ;
  assign n6220 = \g1426_reg/NET0131  & ~n2280 ;
  assign n6221 = n2283 & n6220 ;
  assign n6222 = ~\g1457_reg/NET0131  & ~n2361 ;
  assign n6223 = ~n6221 & ~n6222 ;
  assign n6224 = \g1457_reg/NET0131  & ~n2358 ;
  assign n6225 = n2357 & n6224 ;
  assign n6226 = \g1448_reg/NET0131  & ~n2364 ;
  assign n6227 = n2367 & n6226 ;
  assign n6228 = ~n6225 & ~n6227 ;
  assign n6229 = n6223 & n6228 ;
  assign n6230 = \g1435_reg/NET0131  & ~n2291 ;
  assign n6231 = n2290 & n6230 ;
  assign n6232 = \g1466_reg/NET0131  & ~n2339 ;
  assign n6233 = n2338 & n6232 ;
  assign n6234 = ~n6231 & ~n6233 ;
  assign n6235 = ~\g1435_reg/NET0131  & ~n2294 ;
  assign n6236 = ~\g1426_reg/NET0131  & ~n2284 ;
  assign n6237 = ~n6235 & ~n6236 ;
  assign n6238 = n6234 & n6237 ;
  assign n6239 = n6229 & n6238 ;
  assign n6240 = ~\g2896_reg/NET0131  & ~\g2900_reg/NET0131  ;
  assign n6241 = ~\g2892_reg/NET0131  & ~\g2903_reg/NET0131  ;
  assign n6242 = ~\g2908_reg/NET0131  & n6241 ;
  assign n6243 = n6240 & n6242 ;
  assign n6244 = ~n2146 & n2151 ;
  assign n6245 = ~n2269 & n6244 ;
  assign n6246 = ~n6243 & ~n6245 ;
  assign n6247 = \g1453_reg/NET0131  & ~n2329 ;
  assign n6248 = n2328 & n6247 ;
  assign n6249 = \g1439_reg/NET0131  & ~n2345 ;
  assign n6250 = n2348 & n6249 ;
  assign n6251 = ~n6248 & ~n6250 ;
  assign n6252 = ~\g1439_reg/NET0131  & ~n2349 ;
  assign n6253 = ~\g1453_reg/NET0131  & ~n2332 ;
  assign n6254 = ~n6252 & ~n6253 ;
  assign n6255 = n6251 & n6254 ;
  assign n6256 = n6246 & n6255 ;
  assign n6257 = n6239 & n6256 ;
  assign n6258 = \g1462_reg/NET0131  & ~n2312 ;
  assign n6259 = ~\g1462_reg/NET0131  & ~n2309 ;
  assign n6260 = n2308 & n6259 ;
  assign n6261 = ~n6258 & ~n6260 ;
  assign n6262 = \g1430_reg/NET0131  & ~n2302 ;
  assign n6263 = ~\g1430_reg/NET0131  & ~n2298 ;
  assign n6264 = n2301 & n6263 ;
  assign n6265 = ~n6262 & ~n6264 ;
  assign n6266 = ~n6261 & ~n6265 ;
  assign n6267 = ~\g1448_reg/NET0131  & ~n2368 ;
  assign n6268 = ~\g1466_reg/NET0131  & ~n2342 ;
  assign n6269 = ~n6267 & ~n6268 ;
  assign n6270 = \g1444_reg/NET0131  & ~n2323 ;
  assign n6271 = ~\g1444_reg/NET0131  & ~n2320 ;
  assign n6272 = n2319 & n6271 ;
  assign n6273 = ~n6270 & ~n6272 ;
  assign n6274 = n6269 & ~n6273 ;
  assign n6275 = n6266 & n6274 ;
  assign n6276 = n6257 & n6275 ;
  assign n6277 = n2415 & n3390 ;
  assign n6278 = n3392 & n6277 ;
  assign n6279 = n3412 & n3414 ;
  assign n6280 = n3413 & n6279 ;
  assign n6281 = n6278 & n6280 ;
  assign n6282 = ~n6276 & ~n6281 ;
  assign n6283 = \g1444_reg/NET0131  & ~n2707 ;
  assign n6284 = n2710 & n6283 ;
  assign n6285 = ~\g1426_reg/NET0131  & ~n2679 ;
  assign n6286 = ~n6284 & ~n6285 ;
  assign n6287 = ~\g1430_reg/NET0131  & ~n2616 ;
  assign n6288 = ~\g1457_reg/NET0131  & ~n2624 ;
  assign n6289 = ~n6287 & ~n6288 ;
  assign n6290 = n6286 & n6289 ;
  assign n6291 = \g1426_reg/NET0131  & ~n2675 ;
  assign n6292 = n2678 & n6291 ;
  assign n6293 = \g1453_reg/NET0131  & ~n2666 ;
  assign n6294 = n2669 & n6293 ;
  assign n6295 = ~n6292 & ~n6294 ;
  assign n6296 = ~\g1439_reg/NET0131  & ~n2635 ;
  assign n6297 = ~\g1448_reg/NET0131  & ~n2607 ;
  assign n6298 = ~n6296 & ~n6297 ;
  assign n6299 = n6295 & n6298 ;
  assign n6300 = n6290 & n6299 ;
  assign n6301 = \g1448_reg/NET0131  & ~n2603 ;
  assign n6302 = n2606 & n6301 ;
  assign n6303 = ~\g1435_reg/NET0131  & ~n2699 ;
  assign n6304 = \g1435_reg/NET0131  & ~n2695 ;
  assign n6305 = n2698 & n6304 ;
  assign n6306 = \g1430_reg/NET0131  & ~n2612 ;
  assign n6307 = n2615 & n6306 ;
  assign n6308 = ~n6305 & ~n6307 ;
  assign n6309 = ~n6303 & n6308 ;
  assign n6310 = ~n6302 & n6309 ;
  assign n6311 = ~\g1453_reg/NET0131  & ~n2670 ;
  assign n6312 = ~\g1444_reg/NET0131  & ~n2711 ;
  assign n6313 = ~n6311 & ~n6312 ;
  assign n6314 = ~\g1462_reg/NET0131  & ~n2688 ;
  assign n6315 = ~\g1466_reg/NET0131  & ~n2648 ;
  assign n6316 = ~n6314 & ~n6315 ;
  assign n6317 = n6313 & n6316 ;
  assign n6318 = n6310 & n6317 ;
  assign n6319 = ~n2453 & ~n2458 ;
  assign n6320 = n2470 & n6319 ;
  assign n6321 = ~n6243 & ~n6320 ;
  assign n6322 = \g1439_reg/NET0131  & ~n2631 ;
  assign n6323 = n2634 & n6322 ;
  assign n6324 = \g1457_reg/NET0131  & ~n2620 ;
  assign n6325 = n2623 & n6324 ;
  assign n6326 = ~n6323 & ~n6325 ;
  assign n6327 = \g1462_reg/NET0131  & ~n2684 ;
  assign n6328 = n2687 & n6327 ;
  assign n6329 = \g1466_reg/NET0131  & ~n2645 ;
  assign n6330 = n2644 & n6329 ;
  assign n6331 = ~n6328 & ~n6330 ;
  assign n6332 = n6326 & n6331 ;
  assign n6333 = n6321 & n6332 ;
  assign n6334 = n6318 & n6333 ;
  assign n6335 = n6300 & n6334 ;
  assign n6336 = n2599 & n3465 ;
  assign n6337 = n3467 & n6336 ;
  assign n6338 = n3473 & n6337 ;
  assign n6339 = ~n6335 & ~n6338 ;
  assign n6340 = \g1439_reg/NET0131  & ~n1261 ;
  assign n6341 = n1264 & n6340 ;
  assign n6342 = ~\g1426_reg/NET0131  & ~n1224 ;
  assign n6343 = ~n6341 & ~n6342 ;
  assign n6344 = ~\g1439_reg/NET0131  & ~n1265 ;
  assign n6345 = \g1430_reg/NET0131  & ~n1275 ;
  assign n6346 = n1278 & n6345 ;
  assign n6347 = ~n6344 & ~n6346 ;
  assign n6348 = n6343 & n6347 ;
  assign n6349 = \g1457_reg/NET0131  & ~n1293 ;
  assign n6350 = n1296 & n6349 ;
  assign n6351 = \g1426_reg/NET0131  & ~n1220 ;
  assign n6352 = n1223 & n6351 ;
  assign n6353 = ~n6350 & ~n6352 ;
  assign n6354 = ~\g1457_reg/NET0131  & ~n1297 ;
  assign n6355 = ~\g1444_reg/NET0131  & ~n1212 ;
  assign n6356 = ~n6354 & ~n6355 ;
  assign n6357 = n6353 & n6356 ;
  assign n6358 = n6348 & n6357 ;
  assign n6359 = ~\g1462_reg/NET0131  & ~n1200 ;
  assign n6360 = ~\g1435_reg/NET0131  & ~n1191 ;
  assign n6361 = ~n6359 & ~n6360 ;
  assign n6362 = \g1444_reg/NET0131  & ~n1209 ;
  assign n6363 = n1208 & n6362 ;
  assign n6364 = n6361 & ~n6363 ;
  assign n6365 = ~\g1466_reg/NET0131  & ~n1290 ;
  assign n6366 = ~\g1430_reg/NET0131  & ~n1279 ;
  assign n6367 = ~n6365 & ~n6366 ;
  assign n6368 = \g1435_reg/NET0131  & ~n1187 ;
  assign n6369 = n1190 & n6368 ;
  assign n6370 = \g1453_reg/NET0131  & ~n1231 ;
  assign n6371 = n1230 & n6370 ;
  assign n6372 = ~n6369 & ~n6371 ;
  assign n6373 = ~\g1453_reg/NET0131  & ~n1234 ;
  assign n6374 = n6372 & ~n6373 ;
  assign n6375 = n6367 & n6374 ;
  assign n6376 = n6364 & n6375 ;
  assign n6377 = ~n1186 & n1437 ;
  assign n6378 = ~n1444 & n6377 ;
  assign n6379 = ~n6243 & ~n6378 ;
  assign n6380 = \g1462_reg/NET0131  & ~n1196 ;
  assign n6381 = n1199 & n6380 ;
  assign n6382 = \g1466_reg/NET0131  & ~n1287 ;
  assign n6383 = n1286 & n6382 ;
  assign n6384 = ~n6381 & ~n6383 ;
  assign n6385 = ~\g1448_reg/NET0131  & ~n1254 ;
  assign n6386 = \g1448_reg/NET0131  & ~n1250 ;
  assign n6387 = n1253 & n6386 ;
  assign n6388 = ~n6385 & ~n6387 ;
  assign n6389 = n6384 & n6388 ;
  assign n6390 = n6379 & n6389 ;
  assign n6391 = n6376 & n6390 ;
  assign n6392 = n6358 & n6391 ;
  assign n6393 = n1445 & n3706 ;
  assign n6394 = n3708 & n6393 ;
  assign n6395 = n3714 & n6394 ;
  assign n6396 = ~n6392 & ~n6395 ;
  assign n6397 = \g1448_reg/NET0131  & ~n2803 ;
  assign n6398 = n2806 & n6397 ;
  assign n6399 = \g1430_reg/NET0131  & ~n2786 ;
  assign n6400 = n2789 & n6399 ;
  assign n6401 = ~n6398 & ~n6400 ;
  assign n6402 = ~\g1439_reg/NET0131  & ~n2798 ;
  assign n6403 = ~\g1426_reg/NET0131  & ~n3000 ;
  assign n6404 = ~n6402 & ~n6403 ;
  assign n6405 = n6401 & n6404 ;
  assign n6406 = \g1439_reg/NET0131  & ~n2794 ;
  assign n6407 = n2797 & n6406 ;
  assign n6408 = \g1462_reg/NET0131  & ~n2965 ;
  assign n6409 = n2968 & n6408 ;
  assign n6410 = ~n6407 & ~n6409 ;
  assign n6411 = \g1457_reg/NET0131  & ~n2822 ;
  assign n6412 = n2825 & n6411 ;
  assign n6413 = n6410 & ~n6412 ;
  assign n6414 = ~n3020 & n3036 ;
  assign n6415 = ~n3048 & n6414 ;
  assign n6416 = \g1444_reg/NET0131  & ~n2959 ;
  assign n6417 = n2958 & n6416 ;
  assign n6418 = ~n6243 & ~n6417 ;
  assign n6419 = ~n6415 & n6418 ;
  assign n6420 = n6413 & n6419 ;
  assign n6421 = n6405 & n6420 ;
  assign n6422 = \g1466_reg/NET0131  & ~n2816 ;
  assign n6423 = n2815 & n6422 ;
  assign n6424 = ~\g1448_reg/NET0131  & ~n2807 ;
  assign n6425 = ~n6423 & ~n6424 ;
  assign n6426 = ~\g1453_reg/NET0131  & ~n2991 ;
  assign n6427 = ~\g1462_reg/NET0131  & ~n2969 ;
  assign n6428 = ~n6426 & ~n6427 ;
  assign n6429 = n6425 & n6428 ;
  assign n6430 = ~\g1435_reg/NET0131  & ~n2974 ;
  assign n6431 = n2977 & n6430 ;
  assign n6432 = \g1435_reg/NET0131  & ~n2978 ;
  assign n6433 = ~n6431 & ~n6432 ;
  assign n6434 = \g1453_reg/NET0131  & ~n2988 ;
  assign n6435 = n2987 & n6434 ;
  assign n6436 = \g1426_reg/NET0131  & ~n2996 ;
  assign n6437 = n2999 & n6436 ;
  assign n6438 = ~n6435 & ~n6437 ;
  assign n6439 = ~n6433 & n6438 ;
  assign n6440 = ~\g1430_reg/NET0131  & ~n2790 ;
  assign n6441 = ~\g1466_reg/NET0131  & ~n2819 ;
  assign n6442 = ~n6440 & ~n6441 ;
  assign n6443 = ~\g1457_reg/NET0131  & ~n2826 ;
  assign n6444 = ~\g1444_reg/NET0131  & ~n2962 ;
  assign n6445 = ~n6443 & ~n6444 ;
  assign n6446 = n6442 & n6445 ;
  assign n6447 = n6439 & n6446 ;
  assign n6448 = n6429 & n6447 ;
  assign n6449 = n6421 & n6448 ;
  assign n6450 = n3069 & n3647 ;
  assign n6451 = n3649 & n6450 ;
  assign n6452 = n3655 & n6451 ;
  assign n6453 = ~n6449 & ~n6452 ;
  assign n6454 = \g1092_reg/NET0131  & ~\g1561_reg/NET0131  ;
  assign n6455 = \g1088_reg/NET0131  & ~\g1559_reg/NET0131  ;
  assign n6456 = ~\g1560_reg/NET0131  & \g7961_pad  ;
  assign n6457 = ~n6455 & ~n6456 ;
  assign n6458 = ~n6454 & n6457 ;
  assign n6459 = n6130 & ~n6458 ;
  assign n6460 = n5960 & ~n6459 ;
  assign n6461 = \g1810_reg/NET0131  & \g7961_pad  ;
  assign n6462 = ~\g1563_reg/NET0131  & ~n6461 ;
  assign n6463 = \g1088_reg/NET0131  & \g1816_reg/NET0131  ;
  assign n6464 = \g1092_reg/NET0131  & ~\g1813_reg/NET0131  ;
  assign n6465 = ~n6463 & n6464 ;
  assign n6466 = n6462 & n6465 ;
  assign n6467 = ~\g1092_reg/NET0131  & ~\g1813_reg/NET0131  ;
  assign n6468 = ~n6466 & ~n6467 ;
  assign n6469 = ~n6460 & n6468 ;
  assign n6470 = \g1092_reg/NET0131  & ~\g867_reg/NET0131  ;
  assign n6471 = \g1088_reg/NET0131  & ~\g865_reg/NET0131  ;
  assign n6472 = \g7961_pad  & ~\g866_reg/NET0131  ;
  assign n6473 = ~n6471 & ~n6472 ;
  assign n6474 = ~n6470 & n6473 ;
  assign n6475 = n6037 & ~n6474 ;
  assign n6476 = n5958 & ~n6475 ;
  assign n6477 = \g1092_reg/NET0131  & \g1119_reg/NET0131  ;
  assign n6478 = \g1088_reg/NET0131  & \g1122_reg/NET0131  ;
  assign n6479 = ~n6477 & ~n6478 ;
  assign n6480 = ~\g1116_reg/NET0131  & \g7961_pad  ;
  assign n6481 = ~\g1563_reg/NET0131  & n6480 ;
  assign n6482 = n6479 & n6481 ;
  assign n6483 = ~\g1116_reg/NET0131  & ~\g7961_pad  ;
  assign n6484 = ~n6482 & ~n6483 ;
  assign n6485 = ~n6476 & n6484 ;
  assign n6486 = n5960 & ~n6475 ;
  assign n6487 = \g1116_reg/NET0131  & \g7961_pad  ;
  assign n6488 = ~\g1563_reg/NET0131  & ~n6487 ;
  assign n6489 = \g1092_reg/NET0131  & ~\g1119_reg/NET0131  ;
  assign n6490 = ~n6478 & n6489 ;
  assign n6491 = n6488 & n6490 ;
  assign n6492 = ~\g1092_reg/NET0131  & ~\g1119_reg/NET0131  ;
  assign n6493 = ~n6491 & ~n6492 ;
  assign n6494 = ~n6486 & n6493 ;
  assign n6495 = n5952 & ~n6475 ;
  assign n6496 = \g1088_reg/NET0131  & ~\g1122_reg/NET0131  ;
  assign n6497 = ~n6477 & n6496 ;
  assign n6498 = n6488 & n6497 ;
  assign n6499 = ~\g1088_reg/NET0131  & ~\g1122_reg/NET0131  ;
  assign n6500 = ~n6498 & ~n6499 ;
  assign n6501 = ~n6495 & n6500 ;
  assign n6502 = \g1088_reg/NET0131  & ~\g1828_reg/NET0131  ;
  assign n6503 = ~\g1829_reg/NET0131  & \g7961_pad  ;
  assign n6504 = \g1092_reg/NET0131  & ~\g1830_reg/NET0131  ;
  assign n6505 = ~n6503 & ~n6504 ;
  assign n6506 = ~n6502 & n6505 ;
  assign n6507 = \g1092_reg/NET0131  & \g1822_reg/NET0131  ;
  assign n6508 = \g1819_reg/NET0131  & \g7961_pad  ;
  assign n6509 = \g1088_reg/NET0131  & \g1825_reg/NET0131  ;
  assign n6510 = ~n6508 & ~n6509 ;
  assign n6511 = ~n6507 & n6510 ;
  assign n6512 = \g1092_reg/NET0131  & \g1813_reg/NET0131  ;
  assign n6513 = ~n6463 & ~n6512 ;
  assign n6514 = ~n6461 & n6513 ;
  assign n6515 = n6511 & n6514 ;
  assign n6516 = n6506 & ~n6515 ;
  assign n6517 = \g1563_reg/NET0131  & n6514 ;
  assign n6518 = ~n6459 & n6517 ;
  assign n6519 = \g1563_reg/NET0131  & n6511 ;
  assign n6520 = n6459 & n6519 ;
  assign n6521 = ~n6518 & ~n6520 ;
  assign n6522 = n6516 & ~n6521 ;
  assign n6523 = ~n6459 & ~n6514 ;
  assign n6524 = ~n6515 & ~n6523 ;
  assign n6525 = ~n6459 & n6511 ;
  assign n6526 = \g1563_reg/NET0131  & ~n6525 ;
  assign n6527 = ~n6524 & n6526 ;
  assign n6528 = ~n6522 & ~n6527 ;
  assign n6529 = \g1088_reg/NET0131  & ~n6528 ;
  assign n6530 = \g7961_pad  & ~n6528 ;
  assign n6531 = \g1092_reg/NET0131  & ~n6528 ;
  assign n6532 = \g1092_reg/NET0131  & \g432_reg/NET0131  ;
  assign n6533 = \g429_reg/NET0131  & \g7961_pad  ;
  assign n6534 = \g1088_reg/NET0131  & \g435_reg/NET0131  ;
  assign n6535 = ~n6533 & ~n6534 ;
  assign n6536 = ~n6532 & n6535 ;
  assign n6537 = \g1092_reg/NET0131  & \g441_reg/NET0131  ;
  assign n6538 = \g438_reg/NET0131  & \g7961_pad  ;
  assign n6539 = \g1088_reg/NET0131  & \g444_reg/NET0131  ;
  assign n6540 = ~n6538 & ~n6539 ;
  assign n6541 = ~n6537 & n6540 ;
  assign n6542 = ~n6536 & n6541 ;
  assign n6543 = \g1092_reg/NET0131  & ~\g179_reg/NET0131  ;
  assign n6544 = \g1088_reg/NET0131  & ~\g177_reg/NET0131  ;
  assign n6545 = ~\g178_reg/NET0131  & \g7961_pad  ;
  assign n6546 = ~n6544 & ~n6545 ;
  assign n6547 = ~n6543 & n6546 ;
  assign n6548 = n6068 & ~n6547 ;
  assign n6549 = ~n6541 & ~n6548 ;
  assign n6550 = ~n6542 & ~n6549 ;
  assign n6551 = ~n6536 & ~n6548 ;
  assign n6552 = ~\g448_reg/NET0131  & \g7961_pad  ;
  assign n6553 = \g1092_reg/NET0131  & ~\g449_reg/NET0131  ;
  assign n6554 = ~n6552 & ~n6553 ;
  assign n6555 = \g1088_reg/NET0131  & ~\g447_reg/NET0131  ;
  assign n6556 = \g1563_reg/NET0131  & ~n6555 ;
  assign n6557 = n6554 & n6556 ;
  assign n6558 = ~n6551 & n6557 ;
  assign n6559 = ~n6550 & n6558 ;
  assign n6560 = n6541 & n6548 ;
  assign n6561 = ~n6551 & ~n6560 ;
  assign n6562 = \g1563_reg/NET0131  & ~n6542 ;
  assign n6563 = ~n6561 & n6562 ;
  assign n6564 = ~n6559 & ~n6563 ;
  assign n6565 = \g7961_pad  & ~n6564 ;
  assign n6566 = \g1088_reg/NET0131  & \g1466_reg/NET0131  ;
  assign n6567 = \g1462_reg/NET0131  & n6566 ;
  assign n6568 = \g1448_reg/NET0131  & \g1457_reg/NET0131  ;
  assign n6569 = \g1453_reg/NET0131  & n6568 ;
  assign n6570 = n6567 & n6569 ;
  assign n6571 = ~n6243 & n6570 ;
  assign n6572 = \g1435_reg/NET0131  & \g1444_reg/NET0131  ;
  assign n6573 = \g1439_reg/NET0131  & n6572 ;
  assign n6574 = \g1426_reg/NET0131  & \g1430_reg/NET0131  ;
  assign n6575 = n6573 & n6574 ;
  assign n6576 = n6571 & n6575 ;
  assign n6577 = n5952 & n6240 ;
  assign n6578 = n6242 & n6577 ;
  assign n6579 = \g1426_reg/NET0131  & ~n6578 ;
  assign n6580 = \g1430_reg/NET0131  & n6573 ;
  assign n6581 = ~n6578 & n6580 ;
  assign n6582 = n6571 & n6581 ;
  assign n6583 = ~n6579 & ~n6582 ;
  assign n6584 = ~n6576 & ~n6583 ;
  assign n6585 = \g1088_reg/NET0131  & ~n6564 ;
  assign n6586 = \g1092_reg/NET0131  & ~n6564 ;
  assign n6587 = \g1088_reg/NET0131  & ~\g1134_reg/NET0131  ;
  assign n6588 = ~\g1135_reg/NET0131  & \g7961_pad  ;
  assign n6589 = \g1092_reg/NET0131  & ~\g1136_reg/NET0131  ;
  assign n6590 = ~n6588 & ~n6589 ;
  assign n6591 = ~n6587 & n6590 ;
  assign n6592 = \g1092_reg/NET0131  & \g1128_reg/NET0131  ;
  assign n6593 = \g1125_reg/NET0131  & \g7961_pad  ;
  assign n6594 = \g1088_reg/NET0131  & \g1131_reg/NET0131  ;
  assign n6595 = ~n6593 & ~n6594 ;
  assign n6596 = ~n6592 & n6595 ;
  assign n6597 = n6479 & ~n6487 ;
  assign n6598 = n6596 & n6597 ;
  assign n6599 = n6591 & ~n6598 ;
  assign n6600 = \g1563_reg/NET0131  & n6597 ;
  assign n6601 = ~n6475 & n6600 ;
  assign n6602 = \g1563_reg/NET0131  & n6596 ;
  assign n6603 = n6475 & n6602 ;
  assign n6604 = ~n6601 & ~n6603 ;
  assign n6605 = n6599 & ~n6604 ;
  assign n6606 = ~n6475 & ~n6597 ;
  assign n6607 = ~n6598 & ~n6606 ;
  assign n6608 = ~n6475 & n6596 ;
  assign n6609 = \g1563_reg/NET0131  & ~n6608 ;
  assign n6610 = ~n6607 & n6609 ;
  assign n6611 = ~n6605 & ~n6610 ;
  assign n6612 = \g1088_reg/NET0131  & ~n6611 ;
  assign n6613 = \g7961_pad  & ~n6611 ;
  assign n6614 = \g1092_reg/NET0131  & ~n6611 ;
  assign n6615 = \g1092_reg/NET0131  & \g2507_reg/NET0131  ;
  assign n6616 = \g2504_reg/NET0131  & \g7961_pad  ;
  assign n6617 = \g1088_reg/NET0131  & \g2510_reg/NET0131  ;
  assign n6618 = ~n6616 & ~n6617 ;
  assign n6619 = ~n6615 & n6618 ;
  assign n6620 = \g1092_reg/NET0131  & \g2516_reg/NET0131  ;
  assign n6621 = \g2513_reg/NET0131  & \g7961_pad  ;
  assign n6622 = \g1088_reg/NET0131  & \g2519_reg/NET0131  ;
  assign n6623 = ~n6621 & ~n6622 ;
  assign n6624 = ~n6620 & n6623 ;
  assign n6625 = ~n6619 & n6624 ;
  assign n6626 = ~\g2254_reg/NET0131  & \g7961_pad  ;
  assign n6627 = \g1092_reg/NET0131  & ~\g2255_reg/NET0131  ;
  assign n6628 = \g1088_reg/NET0131  & ~\g2253_reg/NET0131  ;
  assign n6629 = ~n6627 & ~n6628 ;
  assign n6630 = ~n6626 & n6629 ;
  assign n6631 = n6099 & ~n6630 ;
  assign n6632 = ~n6624 & ~n6631 ;
  assign n6633 = ~n6625 & ~n6632 ;
  assign n6634 = ~n6619 & ~n6631 ;
  assign n6635 = ~\g2523_reg/NET0131  & \g7961_pad  ;
  assign n6636 = \g1092_reg/NET0131  & ~\g2524_reg/NET0131  ;
  assign n6637 = ~n6635 & ~n6636 ;
  assign n6638 = \g1088_reg/NET0131  & ~\g2522_reg/NET0131  ;
  assign n6639 = \g1563_reg/NET0131  & ~n6638 ;
  assign n6640 = n6637 & n6639 ;
  assign n6641 = ~n6634 & n6640 ;
  assign n6642 = ~n6633 & n6641 ;
  assign n6643 = n6624 & n6631 ;
  assign n6644 = ~n6634 & ~n6643 ;
  assign n6645 = \g1563_reg/NET0131  & ~n6625 ;
  assign n6646 = ~n6644 & n6645 ;
  assign n6647 = ~n6642 & ~n6646 ;
  assign n6648 = \g1088_reg/NET0131  & ~n6647 ;
  assign n6649 = \g7961_pad  & ~n6647 ;
  assign n6650 = \g1092_reg/NET0131  & ~n6647 ;
  assign n6651 = \g1092_reg/NET0131  & n2600 ;
  assign n6652 = \g1092_reg/NET0131  & ~n6243 ;
  assign n6653 = ~n6320 & n6652 ;
  assign n6654 = ~n6651 & ~n6653 ;
  assign n6655 = ~\g1056_reg/NET0131  & \g7961_pad  ;
  assign n6656 = ~\g1045_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n6657 = ~\g1048_reg/NET0131  & \g1088_reg/NET0131  ;
  assign n6658 = ~n6656 & ~n6657 ;
  assign n6659 = ~n6655 & n6658 ;
  assign n6660 = ~\g1085_reg/NET0131  & \g7961_pad  ;
  assign n6661 = ~\g1075_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n6662 = ~\g1078_reg/NET0131  & \g1088_reg/NET0131  ;
  assign n6663 = ~n6661 & ~n6662 ;
  assign n6664 = ~n6660 & n6663 ;
  assign n6665 = n6659 & n6664 ;
  assign n6666 = ~\g1041_reg/NET0131  & \g7961_pad  ;
  assign n6667 = ~\g1030_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n6668 = ~\g1033_reg/NET0131  & \g1088_reg/NET0131  ;
  assign n6669 = ~n6667 & ~n6668 ;
  assign n6670 = ~n6666 & n6669 ;
  assign n6671 = \g3229_pad  & ~n6670 ;
  assign n6672 = ~\g3229_pad  & ~n6666 ;
  assign n6673 = n6669 & n6672 ;
  assign n6674 = ~n6671 & ~n6673 ;
  assign n6675 = ~n6665 & ~n6674 ;
  assign n6676 = n6659 & ~n6673 ;
  assign n6677 = ~n6671 & n6676 ;
  assign n6678 = ~n6675 & ~n6677 ;
  assign n6679 = ~n6654 & ~n6678 ;
  assign n6680 = \g1060_reg/NET0131  & n6654 ;
  assign n6681 = ~n6679 & ~n6680 ;
  assign n6682 = \g1088_reg/NET0131  & n2600 ;
  assign n6683 = \g1088_reg/NET0131  & ~n6243 ;
  assign n6684 = ~n6320 & n6683 ;
  assign n6685 = ~n6682 & ~n6684 ;
  assign n6686 = ~n6678 & ~n6685 ;
  assign n6687 = \g1063_reg/NET0131  & n6685 ;
  assign n6688 = ~n6686 & ~n6687 ;
  assign n6689 = \g7961_pad  & n2600 ;
  assign n6690 = \g7961_pad  & ~n6243 ;
  assign n6691 = ~n6320 & n6690 ;
  assign n6692 = ~n6689 & ~n6691 ;
  assign n6693 = ~n6678 & ~n6692 ;
  assign n6694 = \g1071_reg/NET0131  & n6692 ;
  assign n6695 = ~n6693 & ~n6694 ;
  assign n6696 = \g1871_reg/NET0131  & \g5657_pad  ;
  assign n6697 = \g1024_reg/NET0131  & \g1877_reg/NET0131  ;
  assign n6698 = ~n6696 & ~n6697 ;
  assign n6699 = \g1018_reg/NET0131  & \g1874_reg/NET0131  ;
  assign n6700 = \g1196_reg/NET0131  & ~n6699 ;
  assign n6701 = n6698 & n6700 ;
  assign n6702 = ~n1905 & n6701 ;
  assign n6703 = \g1024_reg/NET0131  & n6702 ;
  assign n6704 = n6698 & ~n6699 ;
  assign n6705 = ~n1892 & ~n6704 ;
  assign n6706 = ~\g3002_reg/NET0131  & ~\g3006_reg/NET0131  ;
  assign n6707 = ~\g3010_reg/NET0131  & ~\g3013_reg/NET0131  ;
  assign n6708 = ~\g3024_reg/NET0131  & n6707 ;
  assign n6709 = n6706 & n6708 ;
  assign n6710 = \g1024_reg/NET0131  & ~n6709 ;
  assign n6711 = ~n6705 & n6710 ;
  assign n6712 = ~n6703 & ~n6711 ;
  assign n6713 = \g1955_reg/NET0131  & n6712 ;
  assign n6714 = ~n5661 & n5689 ;
  assign n6715 = ~\g3229_pad  & ~n5679 ;
  assign n6716 = ~n6714 & n6715 ;
  assign n6717 = n5689 & ~n5736 ;
  assign n6718 = \g3229_pad  & ~n5695 ;
  assign n6719 = n6717 & n6718 ;
  assign n6720 = ~n6716 & ~n6719 ;
  assign n6721 = ~n6712 & ~n6720 ;
  assign n6722 = ~n6713 & ~n6721 ;
  assign n6723 = \g5657_pad  & n6702 ;
  assign n6724 = \g5657_pad  & ~n6709 ;
  assign n6725 = ~n6705 & n6724 ;
  assign n6726 = ~n6723 & ~n6725 ;
  assign n6727 = \g1956_reg/NET0131  & n6726 ;
  assign n6728 = ~n6720 & ~n6726 ;
  assign n6729 = ~n6727 & ~n6728 ;
  assign n6730 = \g1018_reg/NET0131  & n6702 ;
  assign n6731 = \g1018_reg/NET0131  & ~n6709 ;
  assign n6732 = ~n6705 & n6731 ;
  assign n6733 = ~n6730 & ~n6732 ;
  assign n6734 = \g1957_reg/NET0131  & n6733 ;
  assign n6735 = ~n6720 & ~n6733 ;
  assign n6736 = ~n6734 & ~n6735 ;
  assign n6737 = n2146 & n2415 ;
  assign n6738 = \g1092_reg/NET0131  & n6737 ;
  assign n6739 = ~n6245 & n6652 ;
  assign n6740 = ~n6738 & ~n6739 ;
  assign n6741 = \g343_reg/NET0131  & n6740 ;
  assign n6742 = ~\g398_reg/NET0131  & \g7961_pad  ;
  assign n6743 = \g1092_reg/NET0131  & ~\g388_reg/NET0131  ;
  assign n6744 = \g1088_reg/NET0131  & ~\g391_reg/NET0131  ;
  assign n6745 = ~n6743 & ~n6744 ;
  assign n6746 = ~n6742 & n6745 ;
  assign n6747 = ~\g354_reg/NET0131  & \g7961_pad  ;
  assign n6748 = \g1088_reg/NET0131  & ~\g346_reg/NET0131  ;
  assign n6749 = \g1092_reg/NET0131  & ~\g343_reg/NET0131  ;
  assign n6750 = ~n6748 & ~n6749 ;
  assign n6751 = ~n6747 & n6750 ;
  assign n6752 = n6746 & ~n6751 ;
  assign n6753 = ~\g369_reg/NET0131  & \g7961_pad  ;
  assign n6754 = \g1092_reg/NET0131  & ~\g358_reg/NET0131  ;
  assign n6755 = \g1088_reg/NET0131  & ~\g361_reg/NET0131  ;
  assign n6756 = ~n6754 & ~n6755 ;
  assign n6757 = ~n6753 & n6756 ;
  assign n6758 = \g1092_reg/NET0131  & ~\g373_reg/NET0131  ;
  assign n6759 = \g1088_reg/NET0131  & ~\g376_reg/NET0131  ;
  assign n6760 = ~\g384_reg/NET0131  & \g7961_pad  ;
  assign n6761 = ~n6759 & ~n6760 ;
  assign n6762 = ~n6758 & n6761 ;
  assign n6763 = ~n6757 & n6762 ;
  assign n6764 = ~n6752 & ~n6763 ;
  assign n6765 = ~\g3229_pad  & ~n6764 ;
  assign n6766 = \g3229_pad  & ~n6746 ;
  assign n6767 = \g3229_pad  & ~n6751 ;
  assign n6768 = ~n6763 & n6767 ;
  assign n6769 = ~n6766 & ~n6768 ;
  assign n6770 = ~n6765 & n6769 ;
  assign n6771 = ~n6740 & n6770 ;
  assign n6772 = ~n6741 & ~n6771 ;
  assign n6773 = \g1088_reg/NET0131  & n6737 ;
  assign n6774 = ~n6245 & n6683 ;
  assign n6775 = ~n6773 & ~n6774 ;
  assign n6776 = \g346_reg/NET0131  & n6775 ;
  assign n6777 = n6770 & ~n6775 ;
  assign n6778 = ~n6776 & ~n6777 ;
  assign n6779 = \g7961_pad  & n6737 ;
  assign n6780 = ~n6245 & n6690 ;
  assign n6781 = ~n6779 & ~n6780 ;
  assign n6782 = \g354_reg/NET0131  & n6781 ;
  assign n6783 = n6770 & ~n6781 ;
  assign n6784 = ~n6782 & ~n6783 ;
  assign n6785 = ~\g3229_pad  & ~n6747 ;
  assign n6786 = n6750 & n6785 ;
  assign n6787 = n6757 & ~n6786 ;
  assign n6788 = ~n6767 & n6787 ;
  assign n6789 = ~n6767 & ~n6786 ;
  assign n6790 = n6746 & n6757 ;
  assign n6791 = ~n6789 & ~n6790 ;
  assign n6792 = ~n6788 & ~n6791 ;
  assign n6793 = ~n6740 & ~n6792 ;
  assign n6794 = \g373_reg/NET0131  & n6740 ;
  assign n6795 = ~n6793 & ~n6794 ;
  assign n6796 = ~n6775 & ~n6792 ;
  assign n6797 = \g376_reg/NET0131  & n6775 ;
  assign n6798 = ~n6796 & ~n6797 ;
  assign n6799 = ~n6781 & ~n6792 ;
  assign n6800 = \g384_reg/NET0131  & n6781 ;
  assign n6801 = ~n6799 & ~n6800 ;
  assign n6802 = \g490_reg/NET0131  & \g5657_pad  ;
  assign n6803 = \g1024_reg/NET0131  & \g496_reg/NET0131  ;
  assign n6804 = ~n6802 & ~n6803 ;
  assign n6805 = \g1018_reg/NET0131  & \g493_reg/NET0131  ;
  assign n6806 = \g1196_reg/NET0131  & ~n6805 ;
  assign n6807 = n6804 & n6806 ;
  assign n6808 = ~n4325 & n6807 ;
  assign n6809 = \g1024_reg/NET0131  & n6808 ;
  assign n6810 = n6804 & ~n6805 ;
  assign n6811 = ~n4312 & ~n6810 ;
  assign n6812 = n6710 & ~n6811 ;
  assign n6813 = ~n6809 & ~n6812 ;
  assign n6814 = \g575_reg/NET0131  & n6813 ;
  assign n6815 = ~n5777 & n5817 ;
  assign n6816 = ~\g3229_pad  & ~n6815 ;
  assign n6817 = ~n5842 & n6816 ;
  assign n6818 = ~n5783 & n5817 ;
  assign n6819 = \g3229_pad  & ~n5802 ;
  assign n6820 = n6818 & n6819 ;
  assign n6821 = ~n6817 & ~n6820 ;
  assign n6822 = ~n6813 & ~n6821 ;
  assign n6823 = ~n6814 & ~n6822 ;
  assign n6824 = \g5657_pad  & n6808 ;
  assign n6825 = n6724 & ~n6811 ;
  assign n6826 = ~n6824 & ~n6825 ;
  assign n6827 = \g576_reg/NET0131  & n6826 ;
  assign n6828 = ~n6821 & ~n6826 ;
  assign n6829 = ~n6827 & ~n6828 ;
  assign n6830 = \g1018_reg/NET0131  & n6808 ;
  assign n6831 = n6731 & ~n6811 ;
  assign n6832 = ~n6830 & ~n6831 ;
  assign n6833 = \g577_reg/NET0131  & n6832 ;
  assign n6834 = ~n6821 & ~n6832 ;
  assign n6835 = ~n6833 & ~n6834 ;
  assign n6836 = ~\g1018_reg/NET0131  & ~\g16297_pad  ;
  assign n6837 = ~\g506_reg/NET0131  & n6836 ;
  assign n6838 = ~n4501 & ~n6837 ;
  assign n6839 = \g1177_reg/NET0131  & \g5657_pad  ;
  assign n6840 = \g1024_reg/NET0131  & \g1183_reg/NET0131  ;
  assign n6841 = ~n6839 & ~n6840 ;
  assign n6842 = \g1018_reg/NET0131  & \g1180_reg/NET0131  ;
  assign n6843 = \g1196_reg/NET0131  & ~n6842 ;
  assign n6844 = n6841 & n6843 ;
  assign n6845 = ~n3176 & n6844 ;
  assign n6846 = \g1024_reg/NET0131  & n6845 ;
  assign n6847 = n6841 & ~n6842 ;
  assign n6848 = ~n3188 & ~n6847 ;
  assign n6849 = n6710 & ~n6848 ;
  assign n6850 = ~n6846 & ~n6849 ;
  assign n6851 = \g1261_reg/NET0131  & n6850 ;
  assign n6852 = ~n4993 & ~n4996 ;
  assign n6853 = ~\g3229_pad  & n6852 ;
  assign n6854 = ~n4925 & ~n5012 ;
  assign n6855 = \g3229_pad  & n4954 ;
  assign n6856 = n6854 & n6855 ;
  assign n6857 = ~n6853 & ~n6856 ;
  assign n6858 = ~n6850 & ~n6857 ;
  assign n6859 = ~n6851 & ~n6858 ;
  assign n6860 = \g5657_pad  & n6845 ;
  assign n6861 = n6724 & ~n6848 ;
  assign n6862 = ~n6860 & ~n6861 ;
  assign n6863 = \g1262_reg/NET0131  & n6862 ;
  assign n6864 = ~n6857 & ~n6862 ;
  assign n6865 = ~n6863 & ~n6864 ;
  assign n6866 = \g1018_reg/NET0131  & n6845 ;
  assign n6867 = n6731 & ~n6848 ;
  assign n6868 = ~n6866 & ~n6867 ;
  assign n6869 = \g1263_reg/NET0131  & n6868 ;
  assign n6870 = ~n6857 & ~n6868 ;
  assign n6871 = ~n6869 & ~n6870 ;
  assign n6872 = ~n4925 & ~n5007 ;
  assign n6873 = n4924 & ~n4954 ;
  assign n6874 = \g3229_pad  & ~n6873 ;
  assign n6875 = ~n6872 & n6874 ;
  assign n6876 = ~\g3229_pad  & ~n6873 ;
  assign n6877 = n6872 & n6876 ;
  assign n6878 = ~n6875 & ~n6877 ;
  assign n6879 = ~n6850 & n6878 ;
  assign n6880 = \g1267_reg/NET0131  & n6850 ;
  assign n6881 = ~n6879 & ~n6880 ;
  assign n6882 = \g1092_reg/NET0131  & n1446 ;
  assign n6883 = ~n6378 & n6652 ;
  assign n6884 = ~n6882 & ~n6883 ;
  assign n6885 = \g2418_reg/NET0131  & n6884 ;
  assign n6886 = ~\g2473_reg/NET0131  & \g7961_pad  ;
  assign n6887 = \g1092_reg/NET0131  & ~\g2463_reg/NET0131  ;
  assign n6888 = \g1088_reg/NET0131  & ~\g2466_reg/NET0131  ;
  assign n6889 = ~n6887 & ~n6888 ;
  assign n6890 = ~n6886 & n6889 ;
  assign n6891 = ~\g2429_reg/NET0131  & \g7961_pad  ;
  assign n6892 = \g1088_reg/NET0131  & ~\g2421_reg/NET0131  ;
  assign n6893 = \g1092_reg/NET0131  & ~\g2418_reg/NET0131  ;
  assign n6894 = ~n6892 & ~n6893 ;
  assign n6895 = ~n6891 & n6894 ;
  assign n6896 = n6890 & ~n6895 ;
  assign n6897 = ~\g2444_reg/NET0131  & \g7961_pad  ;
  assign n6898 = \g1092_reg/NET0131  & ~\g2433_reg/NET0131  ;
  assign n6899 = \g1088_reg/NET0131  & ~\g2436_reg/NET0131  ;
  assign n6900 = ~n6898 & ~n6899 ;
  assign n6901 = ~n6897 & n6900 ;
  assign n6902 = \g1092_reg/NET0131  & ~\g2448_reg/NET0131  ;
  assign n6903 = \g1088_reg/NET0131  & ~\g2451_reg/NET0131  ;
  assign n6904 = ~\g2459_reg/NET0131  & \g7961_pad  ;
  assign n6905 = ~n6903 & ~n6904 ;
  assign n6906 = ~n6902 & n6905 ;
  assign n6907 = ~n6901 & n6906 ;
  assign n6908 = ~n6896 & ~n6907 ;
  assign n6909 = ~\g3229_pad  & ~n6908 ;
  assign n6910 = \g3229_pad  & ~n6890 ;
  assign n6911 = \g3229_pad  & ~n6895 ;
  assign n6912 = ~n6907 & n6911 ;
  assign n6913 = ~n6910 & ~n6912 ;
  assign n6914 = ~n6909 & n6913 ;
  assign n6915 = ~n6884 & n6914 ;
  assign n6916 = ~n6885 & ~n6915 ;
  assign n6917 = ~n6862 & n6878 ;
  assign n6918 = \g1268_reg/NET0131  & n6862 ;
  assign n6919 = ~n6917 & ~n6918 ;
  assign n6920 = ~n6868 & n6878 ;
  assign n6921 = \g1269_reg/NET0131  & n6868 ;
  assign n6922 = ~n6920 & ~n6921 ;
  assign n6923 = \g1088_reg/NET0131  & n1446 ;
  assign n6924 = ~n6378 & n6683 ;
  assign n6925 = ~n6923 & ~n6924 ;
  assign n6926 = \g2421_reg/NET0131  & n6925 ;
  assign n6927 = n6914 & ~n6925 ;
  assign n6928 = ~n6926 & ~n6927 ;
  assign n6929 = \g7961_pad  & n1446 ;
  assign n6930 = ~n6378 & n6690 ;
  assign n6931 = ~n6929 & ~n6930 ;
  assign n6932 = \g2429_reg/NET0131  & n6931 ;
  assign n6933 = n6914 & ~n6931 ;
  assign n6934 = ~n6932 & ~n6933 ;
  assign n6935 = ~\g3229_pad  & ~n6891 ;
  assign n6936 = n6894 & n6935 ;
  assign n6937 = n6901 & ~n6936 ;
  assign n6938 = ~n6911 & n6937 ;
  assign n6939 = ~n6911 & ~n6936 ;
  assign n6940 = n6890 & n6901 ;
  assign n6941 = ~n6939 & ~n6940 ;
  assign n6942 = ~n6938 & ~n6941 ;
  assign n6943 = ~n6884 & ~n6942 ;
  assign n6944 = \g2448_reg/NET0131  & n6884 ;
  assign n6945 = ~n6943 & ~n6944 ;
  assign n6946 = ~n6925 & ~n6942 ;
  assign n6947 = \g2451_reg/NET0131  & n6925 ;
  assign n6948 = ~n6946 & ~n6947 ;
  assign n6949 = ~n6931 & ~n6942 ;
  assign n6950 = \g2459_reg/NET0131  & n6931 ;
  assign n6951 = ~n6949 & ~n6950 ;
  assign n6952 = \g1030_reg/NET0131  & n6654 ;
  assign n6953 = ~\g1060_reg/NET0131  & \g1092_reg/NET0131  ;
  assign n6954 = ~\g1063_reg/NET0131  & \g1088_reg/NET0131  ;
  assign n6955 = ~\g1071_reg/NET0131  & \g7961_pad  ;
  assign n6956 = ~n6954 & ~n6955 ;
  assign n6957 = ~n6953 & n6956 ;
  assign n6958 = ~n6659 & n6957 ;
  assign n6959 = n6664 & ~n6670 ;
  assign n6960 = ~n6958 & ~n6959 ;
  assign n6961 = ~\g3229_pad  & ~n6960 ;
  assign n6962 = \g3229_pad  & ~n6664 ;
  assign n6963 = n6671 & ~n6958 ;
  assign n6964 = ~n6962 & ~n6963 ;
  assign n6965 = ~n6961 & n6964 ;
  assign n6966 = ~n6654 & n6965 ;
  assign n6967 = ~n6952 & ~n6966 ;
  assign n6968 = \g2565_reg/NET0131  & \g5657_pad  ;
  assign n6969 = \g1024_reg/NET0131  & \g2571_reg/NET0131  ;
  assign n6970 = ~n6968 & ~n6969 ;
  assign n6971 = \g1018_reg/NET0131  & \g2568_reg/NET0131  ;
  assign n6972 = \g1196_reg/NET0131  & ~n6971 ;
  assign n6973 = n6970 & n6972 ;
  assign n6974 = ~n1589 & n6973 ;
  assign n6975 = \g1024_reg/NET0131  & n6974 ;
  assign n6976 = n6970 & ~n6971 ;
  assign n6977 = ~n1673 & ~n6976 ;
  assign n6978 = n6710 & ~n6977 ;
  assign n6979 = ~n6975 & ~n6978 ;
  assign n6980 = \g2649_reg/NET0131  & n6979 ;
  assign n6981 = ~\g3229_pad  & ~n5128 ;
  assign n6982 = ~n5141 & n6981 ;
  assign n6983 = ~n5086 & n5111 ;
  assign n6984 = \g3229_pad  & ~n5094 ;
  assign n6985 = n6983 & n6984 ;
  assign n6986 = ~n6982 & ~n6985 ;
  assign n6987 = ~n6979 & ~n6986 ;
  assign n6988 = ~n6980 & ~n6987 ;
  assign n6989 = n3048 & n3069 ;
  assign n6990 = \g1092_reg/NET0131  & n6989 ;
  assign n6991 = ~n6415 & n6652 ;
  assign n6992 = ~n6990 & ~n6991 ;
  assign n6993 = \g1724_reg/NET0131  & n6992 ;
  assign n6994 = ~\g1779_reg/NET0131  & \g7961_pad  ;
  assign n6995 = \g1092_reg/NET0131  & ~\g1769_reg/NET0131  ;
  assign n6996 = \g1088_reg/NET0131  & ~\g1772_reg/NET0131  ;
  assign n6997 = ~n6995 & ~n6996 ;
  assign n6998 = ~n6994 & n6997 ;
  assign n6999 = ~\g1735_reg/NET0131  & \g7961_pad  ;
  assign n7000 = \g1088_reg/NET0131  & ~\g1727_reg/NET0131  ;
  assign n7001 = \g1092_reg/NET0131  & ~\g1724_reg/NET0131  ;
  assign n7002 = ~n7000 & ~n7001 ;
  assign n7003 = ~n6999 & n7002 ;
  assign n7004 = n6998 & ~n7003 ;
  assign n7005 = ~\g1750_reg/NET0131  & \g7961_pad  ;
  assign n7006 = \g1092_reg/NET0131  & ~\g1739_reg/NET0131  ;
  assign n7007 = \g1088_reg/NET0131  & ~\g1742_reg/NET0131  ;
  assign n7008 = ~n7006 & ~n7007 ;
  assign n7009 = ~n7005 & n7008 ;
  assign n7010 = \g1092_reg/NET0131  & ~\g1754_reg/NET0131  ;
  assign n7011 = \g1088_reg/NET0131  & ~\g1757_reg/NET0131  ;
  assign n7012 = ~\g1765_reg/NET0131  & \g7961_pad  ;
  assign n7013 = ~n7011 & ~n7012 ;
  assign n7014 = ~n7010 & n7013 ;
  assign n7015 = ~n7009 & n7014 ;
  assign n7016 = ~n7004 & ~n7015 ;
  assign n7017 = ~\g3229_pad  & ~n7016 ;
  assign n7018 = \g3229_pad  & ~n6998 ;
  assign n7019 = \g3229_pad  & ~n7003 ;
  assign n7020 = ~n7015 & n7019 ;
  assign n7021 = ~n7018 & ~n7020 ;
  assign n7022 = ~n7017 & n7021 ;
  assign n7023 = ~n6992 & n7022 ;
  assign n7024 = ~n6993 & ~n7023 ;
  assign n7025 = \g5657_pad  & n6974 ;
  assign n7026 = n6724 & ~n6977 ;
  assign n7027 = ~n7025 & ~n7026 ;
  assign n7028 = \g2650_reg/NET0131  & n7027 ;
  assign n7029 = ~n6986 & ~n7027 ;
  assign n7030 = ~n7028 & ~n7029 ;
  assign n7031 = \g1018_reg/NET0131  & n6974 ;
  assign n7032 = n6731 & ~n6977 ;
  assign n7033 = ~n7031 & ~n7032 ;
  assign n7034 = \g2651_reg/NET0131  & n7033 ;
  assign n7035 = ~n6986 & ~n7033 ;
  assign n7036 = ~n7034 & ~n7035 ;
  assign n7037 = \g2655_reg/NET0131  & n6979 ;
  assign n7038 = ~\g3229_pad  & n5177 ;
  assign n7039 = ~\g3229_pad  & ~n5107 ;
  assign n7040 = n5110 & n7039 ;
  assign n7041 = n5162 & n7040 ;
  assign n7042 = ~n7038 & ~n7041 ;
  assign n7043 = \g3229_pad  & ~n5081 ;
  assign n7044 = n5084 & n7043 ;
  assign n7045 = ~n5080 & n7044 ;
  assign n7046 = \g3229_pad  & ~n5107 ;
  assign n7047 = n5110 & n7046 ;
  assign n7048 = n5086 & n7047 ;
  assign n7049 = ~n7045 & ~n7048 ;
  assign n7050 = n7042 & n7049 ;
  assign n7051 = ~n6979 & n7050 ;
  assign n7052 = ~n7037 & ~n7051 ;
  assign n7053 = \g2656_reg/NET0131  & n7027 ;
  assign n7054 = ~n7027 & n7050 ;
  assign n7055 = ~n7053 & ~n7054 ;
  assign n7056 = \g2657_reg/NET0131  & n7033 ;
  assign n7057 = ~n7033 & n7050 ;
  assign n7058 = ~n7056 & ~n7057 ;
  assign n7059 = \g1088_reg/NET0131  & n6989 ;
  assign n7060 = ~n6415 & n6683 ;
  assign n7061 = ~n7059 & ~n7060 ;
  assign n7062 = \g1727_reg/NET0131  & n7061 ;
  assign n7063 = n7022 & ~n7061 ;
  assign n7064 = ~n7062 & ~n7063 ;
  assign n7065 = \g7961_pad  & n6989 ;
  assign n7066 = ~n6415 & n6690 ;
  assign n7067 = ~n7065 & ~n7066 ;
  assign n7068 = \g1735_reg/NET0131  & n7067 ;
  assign n7069 = n7022 & ~n7067 ;
  assign n7070 = ~n7068 & ~n7069 ;
  assign n7071 = ~\g3229_pad  & ~n6999 ;
  assign n7072 = n7002 & n7071 ;
  assign n7073 = n7009 & ~n7072 ;
  assign n7074 = ~n7019 & n7073 ;
  assign n7075 = ~n7019 & ~n7072 ;
  assign n7076 = n6998 & n7009 ;
  assign n7077 = ~n7075 & ~n7076 ;
  assign n7078 = ~n7074 & ~n7077 ;
  assign n7079 = ~n6992 & ~n7078 ;
  assign n7080 = \g1754_reg/NET0131  & n6992 ;
  assign n7081 = ~n7079 & ~n7080 ;
  assign n7082 = ~n7061 & ~n7078 ;
  assign n7083 = \g1757_reg/NET0131  & n7061 ;
  assign n7084 = ~n7082 & ~n7083 ;
  assign n7085 = ~n7067 & ~n7078 ;
  assign n7086 = \g1765_reg/NET0131  & n7067 ;
  assign n7087 = ~n7085 & ~n7086 ;
  assign n7088 = \g1033_reg/NET0131  & n6685 ;
  assign n7089 = ~n6685 & n6965 ;
  assign n7090 = ~n7088 & ~n7089 ;
  assign n7091 = \g1041_reg/NET0131  & n6692 ;
  assign n7092 = ~n6692 & n6965 ;
  assign n7093 = ~n7091 & ~n7092 ;
  assign n7094 = ~n6506 & ~n6515 ;
  assign n7095 = n6511 & n7094 ;
  assign n7096 = ~n6521 & n7095 ;
  assign n7097 = ~n6521 & n7094 ;
  assign n7098 = ~n6511 & ~n7097 ;
  assign n7099 = ~n7096 & ~n7098 ;
  assign n7100 = ~n6591 & ~n6598 ;
  assign n7101 = n6596 & n7100 ;
  assign n7102 = ~n6604 & n7101 ;
  assign n7103 = ~n6604 & n7100 ;
  assign n7104 = ~n6596 & ~n7103 ;
  assign n7105 = ~n7102 & ~n7104 ;
  assign n7106 = n6554 & ~n6555 ;
  assign n7107 = \g1563_reg/NET0131  & ~n7106 ;
  assign n7108 = ~n6551 & n7107 ;
  assign n7109 = ~n6550 & n7108 ;
  assign n7110 = n6541 & ~n7109 ;
  assign n7111 = ~n6541 & n6549 ;
  assign n7112 = n7108 & n7111 ;
  assign n7113 = ~n7110 & ~n7112 ;
  assign n7114 = n6637 & ~n6638 ;
  assign n7115 = \g1563_reg/NET0131  & ~n7114 ;
  assign n7116 = ~n6634 & n7115 ;
  assign n7117 = ~n6633 & n7116 ;
  assign n7118 = n6624 & ~n7117 ;
  assign n7119 = ~n6624 & n6632 ;
  assign n7120 = n7116 & n7119 ;
  assign n7121 = ~n7118 & ~n7120 ;
  assign n7122 = ~n6015 & n6020 ;
  assign n7123 = n6150 & n7122 ;
  assign n7124 = ~n6046 & n6051 ;
  assign n7125 = n6159 & n7124 ;
  assign n7126 = ~n6077 & n6082 ;
  assign n7127 = n6168 & n7126 ;
  assign n7128 = n6108 & ~n6113 ;
  assign n7129 = n6177 & n7128 ;
  assign n7130 = \g3024_reg/NET0131  & \g3080_reg/NET0131  ;
  assign n7131 = n5046 & n7130 ;
  assign n7132 = n5050 & n7131 ;
  assign n7133 = ~\g3028_reg/NET0131  & \g3032_reg/NET0131  ;
  assign n7134 = ~\g3036_reg/NET0131  & n7133 ;
  assign n7135 = ~\g3028_reg/NET0131  & ~\g3234_pad  ;
  assign n7136 = \g3018_reg/NET0131  & n7135 ;
  assign n7137 = ~n7134 & n7136 ;
  assign n7138 = n7132 & n7137 ;
  assign n7139 = \g3018_reg/NET0131  & n7132 ;
  assign n7140 = \g3028_reg/NET0131  & ~\g3234_pad  ;
  assign n7141 = ~n7139 & n7140 ;
  assign n7142 = ~n7138 & ~n7141 ;
  assign n7143 = ~\g1425_reg/NET0131  & ~n5445 ;
  assign n7144 = ~n6004 & ~n7143 ;
  assign n7145 = ~\g739_reg/NET0131  & ~n5595 ;
  assign n7146 = ~n6004 & ~n7145 ;
  assign n7147 = \g1563_reg/NET0131  & ~n6548 ;
  assign n7148 = ~\g1563_reg/NET0131  & ~n6532 ;
  assign n7149 = n6535 & n7148 ;
  assign n7150 = ~n7147 & ~n7149 ;
  assign n7151 = \g1563_reg/NET0131  & ~n6631 ;
  assign n7152 = ~\g1563_reg/NET0131  & ~n6615 ;
  assign n7153 = n6618 & n7152 ;
  assign n7154 = ~n7151 & ~n7153 ;
  assign n7155 = n6462 & n6513 ;
  assign n7156 = \g1563_reg/NET0131  & ~n6459 ;
  assign n7157 = ~n7155 & ~n7156 ;
  assign n7158 = \g3018_reg/NET0131  & \g3036_reg/NET0131  ;
  assign n7159 = \g3028_reg/NET0131  & n7158 ;
  assign n7160 = n7132 & n7159 ;
  assign n7161 = \g3018_reg/NET0131  & n7134 ;
  assign n7162 = n7132 & n7161 ;
  assign n7163 = ~\g3234_pad  & ~n7162 ;
  assign n7164 = n5053 & n7132 ;
  assign n7165 = ~\g3036_reg/NET0131  & ~n7164 ;
  assign n7166 = n7163 & ~n7165 ;
  assign n7167 = ~n7160 & n7166 ;
  assign n7168 = \g3032_reg/NET0131  & n7160 ;
  assign n7169 = ~\g3032_reg/NET0131  & ~n7160 ;
  assign n7170 = ~n7168 & ~n7169 ;
  assign n7171 = n7163 & n7170 ;
  assign n7172 = \g1352_reg/NET0131  & \g1358_reg/NET0131  ;
  assign n7173 = n5998 & n7172 ;
  assign n7174 = ~\g1365_reg/NET0131  & ~n7173 ;
  assign n7175 = ~n6004 & ~n6188 ;
  assign n7176 = ~n7174 & n7175 ;
  assign n7177 = \g3018_reg/NET0131  & ~\g3234_pad  ;
  assign n7178 = ~n7134 & n7177 ;
  assign n7179 = n7132 & n7178 ;
  assign n7180 = ~\g3018_reg/NET0131  & ~\g3234_pad  ;
  assign n7181 = ~n7132 & n7180 ;
  assign n7182 = ~n7179 & ~n7181 ;
  assign n7183 = ~\g3234_pad  & ~n7132 ;
  assign n7184 = \g2993_reg/NET0131  & \g2998_reg/NET0131  ;
  assign n7185 = \g3006_reg/NET0131  & \g3080_reg/NET0131  ;
  assign n7186 = n7184 & n7185 ;
  assign n7187 = \g3002_reg/NET0131  & \g3013_reg/NET0131  ;
  assign n7188 = \g3010_reg/NET0131  & \g3024_reg/NET0131  ;
  assign n7189 = n7187 & n7188 ;
  assign n7190 = n7186 & n7189 ;
  assign n7191 = \g3010_reg/NET0131  & n7187 ;
  assign n7192 = n7186 & n7191 ;
  assign n7193 = ~\g3024_reg/NET0131  & ~n7192 ;
  assign n7194 = ~n7190 & ~n7193 ;
  assign n7195 = n7183 & n7194 ;
  assign n7196 = ~\g3229_pad  & n5731 ;
  assign n7197 = ~\g3229_pad  & ~n5685 ;
  assign n7198 = n5688 & n7197 ;
  assign n7199 = n5668 & n7198 ;
  assign n7200 = ~n7196 & ~n7199 ;
  assign n7201 = \g3229_pad  & ~n5657 ;
  assign n7202 = n5660 & n7201 ;
  assign n7203 = ~n5647 & n7202 ;
  assign n7204 = \g3229_pad  & ~n5685 ;
  assign n7205 = n5688 & n7204 ;
  assign n7206 = n5695 & n7205 ;
  assign n7207 = ~n7203 & ~n7206 ;
  assign n7208 = n7200 & n7207 ;
  assign n7209 = n6571 & n6573 ;
  assign n7210 = \g1430_reg/NET0131  & ~n6578 ;
  assign n7211 = ~n7209 & n7210 ;
  assign n7212 = ~\g1430_reg/NET0131  & n6573 ;
  assign n7213 = ~n6578 & n7212 ;
  assign n7214 = n6571 & n7213 ;
  assign n7215 = ~n7211 & ~n7214 ;
  assign n7216 = \g1439_reg/NET0131  & \g1444_reg/NET0131  ;
  assign n7217 = n6571 & n7216 ;
  assign n7218 = ~\g1435_reg/NET0131  & ~n7217 ;
  assign n7219 = ~n6578 & ~n7209 ;
  assign n7220 = ~n7218 & n7219 ;
  assign n7221 = \g1444_reg/NET0131  & ~n6578 ;
  assign n7222 = ~n6571 & n7221 ;
  assign n7223 = ~\g1444_reg/NET0131  & ~n6578 ;
  assign n7224 = n6571 & n7223 ;
  assign n7225 = ~n7222 & ~n7224 ;
  assign n7226 = \g1457_reg/NET0131  & n6567 ;
  assign n7227 = ~n6243 & n7226 ;
  assign n7228 = ~\g1453_reg/NET0131  & ~n7227 ;
  assign n7229 = \g1453_reg/NET0131  & \g1457_reg/NET0131  ;
  assign n7230 = n6567 & n7229 ;
  assign n7231 = ~n6243 & n7230 ;
  assign n7232 = ~n6578 & ~n7231 ;
  assign n7233 = ~n7228 & n7232 ;
  assign n7234 = ~n6243 & n6567 ;
  assign n7235 = ~\g1462_reg/NET0131  & ~n6566 ;
  assign n7236 = ~\g1462_reg/NET0131  & n6240 ;
  assign n7237 = n6242 & n7236 ;
  assign n7238 = ~n7235 & ~n7237 ;
  assign n7239 = ~n7234 & n7238 ;
  assign n7240 = ~n6578 & n7239 ;
  assign n7241 = \g3229_pad  & ~n5773 ;
  assign n7242 = n5776 & n7241 ;
  assign n7243 = ~n5782 & n7242 ;
  assign n7244 = \g3229_pad  & ~n5813 ;
  assign n7245 = n5816 & n7244 ;
  assign n7246 = n5783 & n7245 ;
  assign n7247 = ~n7243 & ~n7246 ;
  assign n7248 = ~\g3229_pad  & ~n5813 ;
  assign n7249 = n5816 & n7248 ;
  assign n7250 = n5832 & n7249 ;
  assign n7251 = ~n5777 & ~n5782 ;
  assign n7252 = ~\g3229_pad  & n7251 ;
  assign n7253 = ~n7250 & ~n7252 ;
  assign n7254 = n7247 & n7253 ;
  assign n7255 = \g1358_reg/NET0131  & n5998 ;
  assign n7256 = ~\g1352_reg/NET0131  & ~n7255 ;
  assign n7257 = ~n6004 & ~n7173 ;
  assign n7258 = ~n7256 & n7257 ;
  assign n7259 = ~\g2883_reg/NET0131  & \g2888_reg/NET0131  ;
  assign n7260 = n6240 & n7259 ;
  assign n7261 = \g2892_reg/NET0131  & \g2903_reg/NET0131  ;
  assign n7262 = \g2908_reg/NET0131  & \g2950_reg/NET0131  ;
  assign n7263 = n7261 & n7262 ;
  assign n7264 = n7260 & n7263 ;
  assign n7265 = ~\g2917_reg/NET0131  & \g2920_reg/NET0131  ;
  assign n7266 = ~\g2924_reg/NET0131  & n7265 ;
  assign n7267 = \g2912_reg/NET0131  & n7266 ;
  assign n7268 = n7264 & n7267 ;
  assign n7269 = ~\g2814_reg/NET0131  & ~n7268 ;
  assign n7270 = n7260 & n7262 ;
  assign n7271 = \g2912_reg/NET0131  & \g2924_reg/NET0131  ;
  assign n7272 = \g2917_reg/NET0131  & n7271 ;
  assign n7273 = n7261 & n7272 ;
  assign n7274 = n7270 & n7273 ;
  assign n7275 = ~\g2920_reg/NET0131  & ~n7274 ;
  assign n7276 = n7269 & ~n7275 ;
  assign n7277 = \g2920_reg/NET0131  & n7272 ;
  assign n7278 = n7264 & n7277 ;
  assign n7279 = n7276 & ~n7278 ;
  assign n7280 = ~\g2813_reg/NET0131  & ~n5374 ;
  assign n7281 = ~n6004 & ~n7280 ;
  assign n7282 = \g1024_reg/NET0131  & \g1316_reg/NET0131  ;
  assign n7283 = ~\g1423_reg/NET0131  & ~n5383 ;
  assign n7284 = ~n7282 & ~n7283 ;
  assign n7285 = \g1316_reg/NET0131  & \g5657_pad  ;
  assign n7286 = ~\g1424_reg/NET0131  & ~n5453 ;
  assign n7287 = ~n7285 & ~n7286 ;
  assign n7288 = ~\g737_reg/NET0131  & ~n5525 ;
  assign n7289 = ~n7282 & ~n7288 ;
  assign n7290 = ~\g2119_reg/NET0131  & ~n5603 ;
  assign n7291 = ~n6004 & ~n7290 ;
  assign n7292 = ~\g738_reg/NET0131  & ~n5587 ;
  assign n7293 = ~n7285 & ~n7292 ;
  assign n7294 = \g1444_reg/NET0131  & n6571 ;
  assign n7295 = ~\g1439_reg/NET0131  & ~n7294 ;
  assign n7296 = ~n6578 & ~n7217 ;
  assign n7297 = ~n7295 & n7296 ;
  assign n7298 = ~\g1448_reg/NET0131  & ~n7231 ;
  assign n7299 = ~n6571 & ~n6578 ;
  assign n7300 = ~n7298 & n7299 ;
  assign n7301 = ~n6243 & n6566 ;
  assign n7302 = ~\g1088_reg/NET0131  & ~\g1466_reg/NET0131  ;
  assign n7303 = ~\g1466_reg/NET0131  & n6240 ;
  assign n7304 = n6242 & n7303 ;
  assign n7305 = ~n7302 & ~n7304 ;
  assign n7306 = ~n7301 & n7305 ;
  assign n7307 = ~n6578 & n7306 ;
  assign n7308 = \g1457_reg/NET0131  & ~n6567 ;
  assign n7309 = \g1457_reg/NET0131  & n6240 ;
  assign n7310 = n6242 & n7309 ;
  assign n7311 = ~n7308 & ~n7310 ;
  assign n7312 = ~n6578 & ~n7311 ;
  assign n7313 = ~\g1457_reg/NET0131  & n6567 ;
  assign n7314 = ~n6243 & n7313 ;
  assign n7315 = ~n7312 & ~n7314 ;
  assign n7316 = \g1332_reg/NET0131  & \g1339_reg/NET0131  ;
  assign n7317 = n5997 & n7316 ;
  assign n7318 = ~\g1346_reg/NET0131  & ~n7317 ;
  assign n7319 = ~n5998 & ~n6004 ;
  assign n7320 = ~n7318 & n7319 ;
  assign n7321 = \g1358_reg/NET0131  & ~n6004 ;
  assign n7322 = ~n5998 & n7321 ;
  assign n7323 = ~\g1358_reg/NET0131  & ~n6004 ;
  assign n7324 = n5998 & n7323 ;
  assign n7325 = ~n7322 & ~n7324 ;
  assign n7326 = ~\g3229_pad  & ~n5081 ;
  assign n7327 = n5084 & n7326 ;
  assign n7328 = ~n5093 & n7327 ;
  assign n7329 = ~n5141 & ~n7328 ;
  assign n7330 = \g3229_pad  & ~n5085 ;
  assign n7331 = ~n5093 & n7330 ;
  assign n7332 = n7329 & ~n7331 ;
  assign n7333 = ~n6705 & ~n6709 ;
  assign n7334 = ~n6702 & ~n7333 ;
  assign n7335 = ~n6709 & ~n6811 ;
  assign n7336 = ~n6808 & ~n7335 ;
  assign n7337 = ~n6709 & ~n6848 ;
  assign n7338 = ~n6845 & ~n7337 ;
  assign n7339 = ~n6709 & ~n6977 ;
  assign n7340 = ~n6974 & ~n7339 ;
  assign n7341 = n6677 & n6957 ;
  assign n7342 = ~\g3229_pad  & ~n5648 ;
  assign n7343 = n5651 & n7342 ;
  assign n7344 = n5695 & n7343 ;
  assign n7345 = \g3229_pad  & ~n5648 ;
  assign n7346 = n5651 & n7345 ;
  assign n7347 = n5668 & n7346 ;
  assign n7348 = ~n7344 & ~n7347 ;
  assign n7349 = n6762 & n6788 ;
  assign n7350 = ~\g3229_pad  & ~n5797 ;
  assign n7351 = n5800 & n7350 ;
  assign n7352 = n5783 & n7351 ;
  assign n7353 = \g3229_pad  & ~n5797 ;
  assign n7354 = n5800 & n7353 ;
  assign n7355 = n5832 & n7354 ;
  assign n7356 = ~n7352 & ~n7355 ;
  assign n7357 = ~\g3229_pad  & ~n4934 ;
  assign n7358 = n4937 & n7357 ;
  assign n7359 = n4925 & n7358 ;
  assign n7360 = \g3229_pad  & ~n4934 ;
  assign n7361 = n4937 & n7360 ;
  assign n7362 = n5022 & n7361 ;
  assign n7363 = ~n7359 & ~n7362 ;
  assign n7364 = n6906 & n6938 ;
  assign n7365 = \g3229_pad  & ~n5089 ;
  assign n7366 = n5092 & n7365 ;
  assign n7367 = n5162 & n7366 ;
  assign n7368 = ~\g3229_pad  & ~n5089 ;
  assign n7369 = n5092 & n7368 ;
  assign n7370 = n5086 & n7369 ;
  assign n7371 = ~n7367 & ~n7370 ;
  assign n7372 = n7014 & n7074 ;
  assign n7373 = ~\g1384_reg/NET0131  & ~n5383 ;
  assign n7374 = \g1326_reg/NET0131  & n5382 ;
  assign n7375 = n5381 & n7374 ;
  assign n7376 = ~n7373 & ~n7375 ;
  assign n7377 = \g1385_reg/NET0131  & ~n5453 ;
  assign n7378 = ~\g1326_reg/NET0131  & n5453 ;
  assign n7379 = ~n7377 & ~n7378 ;
  assign n7380 = ~\g2811_reg/NET0131  & ~n5619 ;
  assign n7381 = ~n7282 & ~n7380 ;
  assign n7382 = \g1386_reg/NET0131  & ~n5445 ;
  assign n7383 = ~\g1326_reg/NET0131  & n5445 ;
  assign n7384 = ~n7382 & ~n7383 ;
  assign n7385 = ~\g2812_reg/NET0131  & ~n5312 ;
  assign n7386 = ~n7285 & ~n7385 ;
  assign n7387 = \g1387_reg/NET0131  & ~n5383 ;
  assign n7388 = ~\g1319_reg/NET0131  & n5383 ;
  assign n7389 = ~n7387 & ~n7388 ;
  assign n7390 = \g1388_reg/NET0131  & ~n5453 ;
  assign n7391 = ~\g1319_reg/NET0131  & n5453 ;
  assign n7392 = ~n7390 & ~n7391 ;
  assign n7393 = \g1389_reg/NET0131  & ~n5445 ;
  assign n7394 = ~\g1319_reg/NET0131  & n5445 ;
  assign n7395 = ~n7393 & ~n7394 ;
  assign n7396 = \g1390_reg/NET0131  & ~n5383 ;
  assign n7397 = ~\g1339_reg/NET0131  & n5383 ;
  assign n7398 = ~n7396 & ~n7397 ;
  assign n7399 = \g1391_reg/NET0131  & ~n5453 ;
  assign n7400 = ~\g1339_reg/NET0131  & n5453 ;
  assign n7401 = ~n7399 & ~n7400 ;
  assign n7402 = \g1392_reg/NET0131  & ~n5445 ;
  assign n7403 = ~\g1339_reg/NET0131  & n5445 ;
  assign n7404 = ~n7402 & ~n7403 ;
  assign n7405 = \g1393_reg/NET0131  & ~n5383 ;
  assign n7406 = ~\g1332_reg/NET0131  & n5383 ;
  assign n7407 = ~n7405 & ~n7406 ;
  assign n7408 = \g1394_reg/NET0131  & ~n5453 ;
  assign n7409 = ~\g1332_reg/NET0131  & n5453 ;
  assign n7410 = ~n7408 & ~n7409 ;
  assign n7411 = \g1395_reg/NET0131  & ~n5445 ;
  assign n7412 = ~\g1332_reg/NET0131  & n5445 ;
  assign n7413 = ~n7411 & ~n7412 ;
  assign n7414 = \g1396_reg/NET0131  & ~n5383 ;
  assign n7415 = ~\g1346_reg/NET0131  & n5383 ;
  assign n7416 = ~n7414 & ~n7415 ;
  assign n7417 = \g1397_reg/NET0131  & ~n5453 ;
  assign n7418 = ~\g1346_reg/NET0131  & n5453 ;
  assign n7419 = ~n7417 & ~n7418 ;
  assign n7420 = \g1398_reg/NET0131  & ~n5445 ;
  assign n7421 = ~\g1346_reg/NET0131  & n5445 ;
  assign n7422 = ~n7420 & ~n7421 ;
  assign n7423 = \g1399_reg/NET0131  & ~n5383 ;
  assign n7424 = ~\g1358_reg/NET0131  & n5383 ;
  assign n7425 = ~n7423 & ~n7424 ;
  assign n7426 = \g1400_reg/NET0131  & ~n5453 ;
  assign n7427 = ~\g1358_reg/NET0131  & n5453 ;
  assign n7428 = ~n7426 & ~n7427 ;
  assign n7429 = \g1401_reg/NET0131  & ~n5445 ;
  assign n7430 = ~\g1358_reg/NET0131  & n5445 ;
  assign n7431 = ~n7429 & ~n7430 ;
  assign n7432 = \g1402_reg/NET0131  & ~n5383 ;
  assign n7433 = ~\g1352_reg/NET0131  & n5383 ;
  assign n7434 = ~n7432 & ~n7433 ;
  assign n7435 = \g1403_reg/NET0131  & ~n5453 ;
  assign n7436 = ~\g1352_reg/NET0131  & n5453 ;
  assign n7437 = ~n7435 & ~n7436 ;
  assign n7438 = \g1404_reg/NET0131  & ~n5445 ;
  assign n7439 = ~\g1352_reg/NET0131  & n5445 ;
  assign n7440 = ~n7438 & ~n7439 ;
  assign n7441 = \g1405_reg/NET0131  & ~n5383 ;
  assign n7442 = ~\g1365_reg/NET0131  & n5383 ;
  assign n7443 = ~n7441 & ~n7442 ;
  assign n7444 = \g1406_reg/NET0131  & ~n5453 ;
  assign n7445 = ~\g1365_reg/NET0131  & n5453 ;
  assign n7446 = ~n7444 & ~n7445 ;
  assign n7447 = \g1407_reg/NET0131  & ~n5445 ;
  assign n7448 = ~\g1365_reg/NET0131  & n5445 ;
  assign n7449 = ~n7447 & ~n7448 ;
  assign n7450 = \g1408_reg/NET0131  & ~n5383 ;
  assign n7451 = ~\g1372_reg/NET0131  & n5383 ;
  assign n7452 = ~n7450 & ~n7451 ;
  assign n7453 = \g1409_reg/NET0131  & ~n5453 ;
  assign n7454 = ~\g1372_reg/NET0131  & n5453 ;
  assign n7455 = ~n7453 & ~n7454 ;
  assign n7456 = \g1410_reg/NET0131  & ~n5445 ;
  assign n7457 = ~\g1372_reg/NET0131  & n5445 ;
  assign n7458 = ~n7456 & ~n7457 ;
  assign n7459 = \g1411_reg/NET0131  & ~n5383 ;
  assign n7460 = ~\g1378_reg/NET0131  & n5383 ;
  assign n7461 = ~n7459 & ~n7460 ;
  assign n7462 = \g1412_reg/NET0131  & ~n5453 ;
  assign n7463 = ~\g1378_reg/NET0131  & n5453 ;
  assign n7464 = ~n7462 & ~n7463 ;
  assign n7465 = \g1413_reg/NET0131  & ~n5445 ;
  assign n7466 = ~\g1378_reg/NET0131  & n5445 ;
  assign n7467 = ~n7465 & ~n7466 ;
  assign n7468 = \g2232_reg/NET0131  & ~n5952 ;
  assign n7469 = ~\g2200_reg/NET0131  & n5952 ;
  assign n7470 = ~n7468 & ~n7469 ;
  assign n7471 = \g1511_reg/NET0131  & ~n5952 ;
  assign n7472 = ~\g1471_reg/NET0131  & n5952 ;
  assign n7473 = ~n7471 & ~n7472 ;
  assign n7474 = \g1512_reg/NET0131  & ~n5958 ;
  assign n7475 = ~\g1471_reg/NET0131  & n5958 ;
  assign n7476 = ~n7474 & ~n7475 ;
  assign n7477 = \g1513_reg/NET0131  & ~n5960 ;
  assign n7478 = ~\g1471_reg/NET0131  & n5960 ;
  assign n7479 = ~n7477 & ~n7478 ;
  assign n7480 = \g1529_reg/NET0131  & ~n5952 ;
  assign n7481 = ~\g1491_reg/NET0131  & n5952 ;
  assign n7482 = ~n7480 & ~n7481 ;
  assign n7483 = \g1531_reg/NET0131  & ~n5960 ;
  assign n7484 = ~\g1491_reg/NET0131  & n5960 ;
  assign n7485 = ~n7483 & ~n7484 ;
  assign n7486 = \g1530_reg/NET0131  & ~n5958 ;
  assign n7487 = ~\g1491_reg/NET0131  & n5958 ;
  assign n7488 = ~n7486 & ~n7487 ;
  assign n7489 = \g1532_reg/NET0131  & ~n5952 ;
  assign n7490 = ~\g1496_reg/NET0131  & n5952 ;
  assign n7491 = ~n7489 & ~n7490 ;
  assign n7492 = \g1533_reg/NET0131  & ~n5958 ;
  assign n7493 = ~\g1496_reg/NET0131  & n5958 ;
  assign n7494 = ~n7492 & ~n7493 ;
  assign n7495 = \g1534_reg/NET0131  & ~n5960 ;
  assign n7496 = ~\g1496_reg/NET0131  & n5960 ;
  assign n7497 = ~n7495 & ~n7496 ;
  assign n7498 = \g1535_reg/NET0131  & ~n5952 ;
  assign n7499 = ~\g1501_reg/NET0131  & n5952 ;
  assign n7500 = ~n7498 & ~n7499 ;
  assign n7501 = \g1536_reg/NET0131  & ~n5958 ;
  assign n7502 = ~\g1501_reg/NET0131  & n5958 ;
  assign n7503 = ~n7501 & ~n7502 ;
  assign n7504 = \g1537_reg/NET0131  & ~n5960 ;
  assign n7505 = ~\g1501_reg/NET0131  & n5960 ;
  assign n7506 = ~n7504 & ~n7505 ;
  assign n7507 = \g1538_reg/NET0131  & ~n5952 ;
  assign n7508 = ~\g1506_reg/NET0131  & n5952 ;
  assign n7509 = ~n7507 & ~n7508 ;
  assign n7510 = \g1539_reg/NET0131  & ~n5958 ;
  assign n7511 = ~\g1506_reg/NET0131  & n5958 ;
  assign n7512 = ~n7510 & ~n7511 ;
  assign n7513 = \g698_reg/NET0131  & ~n5525 ;
  assign n7514 = ~\g1326_reg/NET0131  & n5525 ;
  assign n7515 = ~n7513 & ~n7514 ;
  assign n7516 = \g699_reg/NET0131  & ~n5587 ;
  assign n7517 = ~\g1326_reg/NET0131  & n5587 ;
  assign n7518 = ~n7516 & ~n7517 ;
  assign n7519 = \g700_reg/NET0131  & ~n5595 ;
  assign n7520 = ~\g1326_reg/NET0131  & n5595 ;
  assign n7521 = ~n7519 & ~n7520 ;
  assign n7522 = \g701_reg/NET0131  & ~n5525 ;
  assign n7523 = ~\g1319_reg/NET0131  & n5525 ;
  assign n7524 = ~n7522 & ~n7523 ;
  assign n7525 = \g702_reg/NET0131  & ~n5587 ;
  assign n7526 = ~\g1319_reg/NET0131  & n5587 ;
  assign n7527 = ~n7525 & ~n7526 ;
  assign n7528 = \g703_reg/NET0131  & ~n5595 ;
  assign n7529 = ~\g1319_reg/NET0131  & n5595 ;
  assign n7530 = ~n7528 & ~n7529 ;
  assign n7531 = \g704_reg/NET0131  & ~n5525 ;
  assign n7532 = ~\g1339_reg/NET0131  & n5525 ;
  assign n7533 = ~n7531 & ~n7532 ;
  assign n7534 = \g705_reg/NET0131  & ~n5587 ;
  assign n7535 = ~\g1339_reg/NET0131  & n5587 ;
  assign n7536 = ~n7534 & ~n7535 ;
  assign n7537 = \g706_reg/NET0131  & ~n5595 ;
  assign n7538 = ~\g1339_reg/NET0131  & n5595 ;
  assign n7539 = ~n7537 & ~n7538 ;
  assign n7540 = \g707_reg/NET0131  & ~n5525 ;
  assign n7541 = ~\g1332_reg/NET0131  & n5525 ;
  assign n7542 = ~n7540 & ~n7541 ;
  assign n7543 = \g708_reg/NET0131  & ~n5587 ;
  assign n7544 = ~\g1332_reg/NET0131  & n5587 ;
  assign n7545 = ~n7543 & ~n7544 ;
  assign n7546 = \g709_reg/NET0131  & ~n5595 ;
  assign n7547 = ~\g1332_reg/NET0131  & n5595 ;
  assign n7548 = ~n7546 & ~n7547 ;
  assign n7549 = \g710_reg/NET0131  & ~n5525 ;
  assign n7550 = ~\g1346_reg/NET0131  & n5525 ;
  assign n7551 = ~n7549 & ~n7550 ;
  assign n7552 = \g711_reg/NET0131  & ~n5587 ;
  assign n7553 = ~\g1346_reg/NET0131  & n5587 ;
  assign n7554 = ~n7552 & ~n7553 ;
  assign n7555 = \g712_reg/NET0131  & ~n5595 ;
  assign n7556 = ~\g1346_reg/NET0131  & n5595 ;
  assign n7557 = ~n7555 & ~n7556 ;
  assign n7558 = \g713_reg/NET0131  & ~n5525 ;
  assign n7559 = ~\g1358_reg/NET0131  & n5525 ;
  assign n7560 = ~n7558 & ~n7559 ;
  assign n7561 = \g714_reg/NET0131  & ~n5587 ;
  assign n7562 = ~\g1358_reg/NET0131  & n5587 ;
  assign n7563 = ~n7561 & ~n7562 ;
  assign n7564 = \g715_reg/NET0131  & ~n5595 ;
  assign n7565 = ~\g1358_reg/NET0131  & n5595 ;
  assign n7566 = ~n7564 & ~n7565 ;
  assign n7567 = \g716_reg/NET0131  & ~n5525 ;
  assign n7568 = ~\g1352_reg/NET0131  & n5525 ;
  assign n7569 = ~n7567 & ~n7568 ;
  assign n7570 = \g717_reg/NET0131  & ~n5587 ;
  assign n7571 = ~\g1352_reg/NET0131  & n5587 ;
  assign n7572 = ~n7570 & ~n7571 ;
  assign n7573 = \g718_reg/NET0131  & ~n5595 ;
  assign n7574 = ~\g1352_reg/NET0131  & n5595 ;
  assign n7575 = ~n7573 & ~n7574 ;
  assign n7576 = \g719_reg/NET0131  & ~n5525 ;
  assign n7577 = ~\g1365_reg/NET0131  & n5525 ;
  assign n7578 = ~n7576 & ~n7577 ;
  assign n7579 = \g720_reg/NET0131  & ~n5587 ;
  assign n7580 = ~\g1365_reg/NET0131  & n5587 ;
  assign n7581 = ~n7579 & ~n7580 ;
  assign n7582 = \g721_reg/NET0131  & ~n5595 ;
  assign n7583 = ~\g1365_reg/NET0131  & n5595 ;
  assign n7584 = ~n7582 & ~n7583 ;
  assign n7585 = \g722_reg/NET0131  & ~n5525 ;
  assign n7586 = ~\g1372_reg/NET0131  & n5525 ;
  assign n7587 = ~n7585 & ~n7586 ;
  assign n7588 = \g723_reg/NET0131  & ~n5587 ;
  assign n7589 = ~\g1372_reg/NET0131  & n5587 ;
  assign n7590 = ~n7588 & ~n7589 ;
  assign n7591 = \g724_reg/NET0131  & ~n5595 ;
  assign n7592 = ~\g1372_reg/NET0131  & n5595 ;
  assign n7593 = ~n7591 & ~n7592 ;
  assign n7594 = \g725_reg/NET0131  & ~n5525 ;
  assign n7595 = ~\g1378_reg/NET0131  & n5525 ;
  assign n7596 = ~n7594 & ~n7595 ;
  assign n7597 = \g726_reg/NET0131  & ~n5587 ;
  assign n7598 = ~\g1378_reg/NET0131  & n5587 ;
  assign n7599 = ~n7597 & ~n7598 ;
  assign n7600 = \g727_reg/NET0131  & ~n5595 ;
  assign n7601 = ~\g1378_reg/NET0131  & n5595 ;
  assign n7602 = ~n7600 & ~n7601 ;
  assign n7603 = ~\g2118_reg/NET0131  & ~n5611 ;
  assign n7604 = ~n7285 & ~n7603 ;
  assign n7605 = \g2229_reg/NET0131  & ~n5952 ;
  assign n7606 = ~\g2195_reg/NET0131  & n5952 ;
  assign n7607 = ~n7605 & ~n7606 ;
  assign n7608 = \g1540_reg/NET0131  & ~n5960 ;
  assign n7609 = ~\g1506_reg/NET0131  & n5960 ;
  assign n7610 = ~n7608 & ~n7609 ;
  assign n7611 = ~\g2117_reg/NET0131  & ~n5462 ;
  assign n7612 = ~n7282 & ~n7611 ;
  assign n7613 = \g1846_reg/NET0131  & ~\g7961_pad  ;
  assign n7614 = ~\g1846_reg/NET0131  & ~\g7961_pad  ;
  assign n7615 = ~n3016 & ~n7614 ;
  assign n7616 = n3019 & n7615 ;
  assign n7617 = n3036 & n7616 ;
  assign n7618 = n3048 & n7617 ;
  assign n7619 = ~n7613 & ~n7618 ;
  assign n7620 = ~\g1092_reg/NET0131  & \g1849_reg/NET0131  ;
  assign n7621 = ~\g1092_reg/NET0131  & ~\g1849_reg/NET0131  ;
  assign n7622 = ~n3016 & ~n7621 ;
  assign n7623 = n3019 & n7622 ;
  assign n7624 = n3036 & n7623 ;
  assign n7625 = n3048 & n7624 ;
  assign n7626 = ~n7620 & ~n7625 ;
  assign n7627 = ~\g1088_reg/NET0131  & \g1852_reg/NET0131  ;
  assign n7628 = ~\g1088_reg/NET0131  & ~\g1852_reg/NET0131  ;
  assign n7629 = ~n3016 & ~n7628 ;
  assign n7630 = n3019 & n7629 ;
  assign n7631 = n3036 & n7630 ;
  assign n7632 = n3048 & n7631 ;
  assign n7633 = ~n7627 & ~n7632 ;
  assign n7634 = \g465_reg/NET0131  & ~\g7961_pad  ;
  assign n7635 = ~\g465_reg/NET0131  & ~\g7961_pad  ;
  assign n7636 = ~n2147 & ~n7635 ;
  assign n7637 = n2150 & n7636 ;
  assign n7638 = n2269 & n7637 ;
  assign n7639 = n2146 & n7638 ;
  assign n7640 = ~n7634 & ~n7639 ;
  assign n7641 = ~\g1092_reg/NET0131  & \g468_reg/NET0131  ;
  assign n7642 = ~\g1092_reg/NET0131  & ~\g468_reg/NET0131  ;
  assign n7643 = ~n2147 & ~n7642 ;
  assign n7644 = n2150 & n7643 ;
  assign n7645 = n2269 & n7644 ;
  assign n7646 = n2146 & n7645 ;
  assign n7647 = ~n7641 & ~n7646 ;
  assign n7648 = ~\g1088_reg/NET0131  & \g471_reg/NET0131  ;
  assign n7649 = ~\g1088_reg/NET0131  & ~\g471_reg/NET0131  ;
  assign n7650 = ~n2147 & ~n7649 ;
  assign n7651 = n2150 & n7650 ;
  assign n7652 = n2269 & n7651 ;
  assign n7653 = n2146 & n7652 ;
  assign n7654 = ~n7648 & ~n7653 ;
  assign n7655 = \g2540_reg/NET0131  & ~\g7961_pad  ;
  assign n7656 = ~\g2540_reg/NET0131  & ~\g7961_pad  ;
  assign n7657 = ~n1182 & ~n7656 ;
  assign n7658 = n1185 & n7657 ;
  assign n7659 = n1437 & n7658 ;
  assign n7660 = n1444 & n7659 ;
  assign n7661 = ~n7655 & ~n7660 ;
  assign n7662 = ~\g1092_reg/NET0131  & \g2543_reg/NET0131  ;
  assign n7663 = ~\g1092_reg/NET0131  & ~\g2543_reg/NET0131  ;
  assign n7664 = ~n1182 & ~n7663 ;
  assign n7665 = n1185 & n7664 ;
  assign n7666 = n1437 & n7665 ;
  assign n7667 = n1444 & n7666 ;
  assign n7668 = ~n7662 & ~n7667 ;
  assign n7669 = ~\g1088_reg/NET0131  & \g2546_reg/NET0131  ;
  assign n7670 = ~\g1088_reg/NET0131  & ~\g2546_reg/NET0131  ;
  assign n7671 = ~n1182 & ~n7670 ;
  assign n7672 = n1185 & n7671 ;
  assign n7673 = n1437 & n7672 ;
  assign n7674 = n1444 & n7673 ;
  assign n7675 = ~n7669 & ~n7674 ;
  assign n7676 = \g847_reg/NET0131  & ~n5952 ;
  assign n7677 = ~n2557 & n5952 ;
  assign n7678 = n2560 & n7677 ;
  assign n7679 = ~n7676 & ~n7678 ;
  assign n7680 = \g848_reg/NET0131  & ~n5958 ;
  assign n7681 = ~n2557 & n5958 ;
  assign n7682 = n2560 & n7681 ;
  assign n7683 = ~n7680 & ~n7682 ;
  assign n7684 = \g849_reg/NET0131  & ~n5960 ;
  assign n7685 = ~n2557 & n5960 ;
  assign n7686 = n2560 & n7685 ;
  assign n7687 = ~n7684 & ~n7686 ;
  assign n7688 = \g850_reg/NET0131  & ~n5952 ;
  assign n7689 = ~n2511 & n5952 ;
  assign n7690 = n2514 & n7689 ;
  assign n7691 = ~n7688 & ~n7690 ;
  assign n7692 = \g851_reg/NET0131  & ~n5958 ;
  assign n7693 = ~n2511 & n5958 ;
  assign n7694 = n2514 & n7693 ;
  assign n7695 = ~n7692 & ~n7694 ;
  assign n7696 = \g852_reg/NET0131  & ~n5960 ;
  assign n7697 = ~n2511 & n5960 ;
  assign n7698 = n2514 & n7697 ;
  assign n7699 = ~n7696 & ~n7698 ;
  assign n7700 = \g159_reg/NET0131  & ~n5952 ;
  assign n7701 = ~n2251 & n5952 ;
  assign n7702 = n2254 & n7701 ;
  assign n7703 = ~n7700 & ~n7702 ;
  assign n7704 = \g160_reg/NET0131  & ~n5958 ;
  assign n7705 = ~n2251 & n5958 ;
  assign n7706 = n2254 & n7705 ;
  assign n7707 = ~n7704 & ~n7706 ;
  assign n7708 = \g161_reg/NET0131  & ~n5960 ;
  assign n7709 = ~n2251 & n5960 ;
  assign n7710 = n2254 & n7709 ;
  assign n7711 = ~n7708 & ~n7710 ;
  assign n7712 = \g162_reg/NET0131  & ~n5952 ;
  assign n7713 = ~n2231 & n5952 ;
  assign n7714 = n2234 & n7713 ;
  assign n7715 = ~n7712 & ~n7714 ;
  assign n7716 = \g163_reg/NET0131  & ~n5958 ;
  assign n7717 = ~n2231 & n5958 ;
  assign n7718 = n2234 & n7717 ;
  assign n7719 = ~n7716 & ~n7718 ;
  assign n7720 = \g164_reg/NET0131  & ~n5960 ;
  assign n7721 = ~n2231 & n5960 ;
  assign n7722 = n2234 & n7721 ;
  assign n7723 = ~n7720 & ~n7722 ;
  assign n7724 = \g838_reg/NET0131  & ~n5952 ;
  assign n7725 = ~\g805_reg/NET0131  & n5952 ;
  assign n7726 = ~n7724 & ~n7725 ;
  assign n7727 = \g150_reg/NET0131  & ~n5952 ;
  assign n7728 = ~\g117_reg/NET0131  & n5952 ;
  assign n7729 = ~n7727 & ~n7728 ;
  assign n7730 = \g151_reg/NET0131  & ~n5958 ;
  assign n7731 = ~\g117_reg/NET0131  & n5958 ;
  assign n7732 = ~n7730 & ~n7731 ;
  assign n7733 = \g152_reg/NET0131  & ~n5960 ;
  assign n7734 = ~\g117_reg/NET0131  & n5960 ;
  assign n7735 = ~n7733 & ~n7734 ;
  assign n7736 = \g839_reg/NET0131  & ~n5958 ;
  assign n7737 = ~\g805_reg/NET0131  & n5958 ;
  assign n7738 = ~n7736 & ~n7737 ;
  assign n7739 = \g840_reg/NET0131  & ~n5960 ;
  assign n7740 = ~\g805_reg/NET0131  & n5960 ;
  assign n7741 = ~n7739 & ~n7740 ;
  assign n7742 = \g844_reg/NET0131  & ~n5952 ;
  assign n7743 = ~\g813_reg/NET0131  & n5952 ;
  assign n7744 = ~n7742 & ~n7743 ;
  assign n7745 = \g845_reg/NET0131  & ~n5958 ;
  assign n7746 = ~\g813_reg/NET0131  & n5958 ;
  assign n7747 = ~n7745 & ~n7746 ;
  assign n7748 = \g846_reg/NET0131  & ~n5960 ;
  assign n7749 = ~\g813_reg/NET0131  & n5960 ;
  assign n7750 = ~n7748 & ~n7749 ;
  assign n7751 = \g156_reg/NET0131  & ~n5952 ;
  assign n7752 = ~\g125_reg/NET0131  & n5952 ;
  assign n7753 = ~n7751 & ~n7752 ;
  assign n7754 = \g157_reg/NET0131  & ~n5958 ;
  assign n7755 = ~\g125_reg/NET0131  & n5958 ;
  assign n7756 = ~n7754 & ~n7755 ;
  assign n7757 = \g158_reg/NET0131  & ~n5960 ;
  assign n7758 = ~\g125_reg/NET0131  & n5960 ;
  assign n7759 = ~n7757 & ~n7758 ;
  assign n7760 = \g1196_reg/NET0131  & ~n1901 ;
  assign n7761 = n1904 & n7760 ;
  assign n7762 = n6704 & n7761 ;
  assign n7763 = \g1196_reg/NET0131  & ~n4321 ;
  assign n7764 = n4324 & n7763 ;
  assign n7765 = n6810 & n7764 ;
  assign n7766 = n3176 & n6844 ;
  assign n7767 = \g1196_reg/NET0131  & ~n1585 ;
  assign n7768 = n1588 & n7767 ;
  assign n7769 = n6976 & n7768 ;
  assign n7770 = \g1339_reg/NET0131  & n5997 ;
  assign n7771 = ~\g1332_reg/NET0131  & ~n7770 ;
  assign n7772 = ~n6004 & ~n7317 ;
  assign n7773 = ~n7771 & n7772 ;
  assign n7774 = n7186 & n7187 ;
  assign n7775 = ~\g3010_reg/NET0131  & ~n7774 ;
  assign n7776 = ~n7192 & ~n7775 ;
  assign n7777 = n7183 & n7776 ;
  assign n7778 = ~n6762 & ~n6789 ;
  assign n7779 = ~n6763 & ~n7778 ;
  assign n7780 = \g3229_pad  & n5736 ;
  assign n7781 = ~\g3229_pad  & ~n5657 ;
  assign n7782 = n5660 & n7781 ;
  assign n7783 = ~n5652 & n7782 ;
  assign n7784 = ~n5679 & ~n7783 ;
  assign n7785 = ~n7780 & n7784 ;
  assign n7786 = \g3229_pad  & n5012 ;
  assign n7787 = ~\g3229_pad  & ~n4915 ;
  assign n7788 = n4918 & n7787 ;
  assign n7789 = ~n4938 & n7788 ;
  assign n7790 = ~n4996 & ~n7789 ;
  assign n7791 = ~n7786 & n7790 ;
  assign n7792 = ~n6906 & ~n6939 ;
  assign n7793 = ~n6907 & ~n7792 ;
  assign n7794 = ~\g3229_pad  & n5773 ;
  assign n7795 = ~n7242 & ~n7794 ;
  assign n7796 = ~\g3229_pad  & ~n5776 ;
  assign n7797 = ~n5801 & ~n7796 ;
  assign n7798 = n7795 & n7797 ;
  assign n7799 = ~n5842 & ~n7798 ;
  assign n7800 = ~n7014 & ~n7075 ;
  assign n7801 = ~n7015 & ~n7800 ;
  assign n7802 = \g1339_reg/NET0131  & ~n6004 ;
  assign n7803 = ~n5997 & n7802 ;
  assign n7804 = ~\g1339_reg/NET0131  & ~n6004 ;
  assign n7805 = n5997 & n7804 ;
  assign n7806 = ~n7803 & ~n7805 ;
  assign n7807 = ~n6674 & ~n6957 ;
  assign n7808 = ~n6958 & ~n7807 ;
  assign n7809 = ~\g2814_reg/NET0131  & ~n7264 ;
  assign n7810 = \g2883_reg/NET0131  & \g2950_reg/NET0131  ;
  assign n7811 = \g2888_reg/NET0131  & \g2896_reg/NET0131  ;
  assign n7812 = n7810 & n7811 ;
  assign n7813 = \g2900_reg/NET0131  & \g2908_reg/NET0131  ;
  assign n7814 = n7261 & n7813 ;
  assign n7815 = n7812 & n7814 ;
  assign n7816 = \g2900_reg/NET0131  & n7261 ;
  assign n7817 = n7812 & n7816 ;
  assign n7818 = ~\g2908_reg/NET0131  & ~n7817 ;
  assign n7819 = ~n7815 & ~n7818 ;
  assign n7820 = n7809 & n7819 ;
  assign n7821 = \g2080_reg/NET0131  & ~n5603 ;
  assign n7822 = ~\g1326_reg/NET0131  & n5603 ;
  assign n7823 = ~n7821 & ~n7822 ;
  assign n7824 = \g2103_reg/NET0131  & ~n5611 ;
  assign n7825 = ~\g1372_reg/NET0131  & n5611 ;
  assign n7826 = ~n7824 & ~n7825 ;
  assign n7827 = \g2092_reg/NET0131  & ~n5603 ;
  assign n7828 = ~\g1346_reg/NET0131  & n5603 ;
  assign n7829 = ~n7827 & ~n7828 ;
  assign n7830 = \g2078_reg/NET0131  & ~n5462 ;
  assign n7831 = ~\g1326_reg/NET0131  & n5462 ;
  assign n7832 = ~n7830 & ~n7831 ;
  assign n7833 = \g2079_reg/NET0131  & ~n5611 ;
  assign n7834 = ~\g1326_reg/NET0131  & n5611 ;
  assign n7835 = ~n7833 & ~n7834 ;
  assign n7836 = \g2081_reg/NET0131  & ~n5462 ;
  assign n7837 = ~\g1319_reg/NET0131  & n5462 ;
  assign n7838 = ~n7836 & ~n7837 ;
  assign n7839 = \g2082_reg/NET0131  & ~n5611 ;
  assign n7840 = ~\g1319_reg/NET0131  & n5611 ;
  assign n7841 = ~n7839 & ~n7840 ;
  assign n7842 = \g2083_reg/NET0131  & ~n5603 ;
  assign n7843 = ~\g1319_reg/NET0131  & n5603 ;
  assign n7844 = ~n7842 & ~n7843 ;
  assign n7845 = \g2084_reg/NET0131  & ~n5462 ;
  assign n7846 = ~\g1339_reg/NET0131  & n5462 ;
  assign n7847 = ~n7845 & ~n7846 ;
  assign n7848 = \g2085_reg/NET0131  & ~n5611 ;
  assign n7849 = ~\g1339_reg/NET0131  & n5611 ;
  assign n7850 = ~n7848 & ~n7849 ;
  assign n7851 = \g2087_reg/NET0131  & ~n5462 ;
  assign n7852 = ~\g1332_reg/NET0131  & n5462 ;
  assign n7853 = ~n7851 & ~n7852 ;
  assign n7854 = \g2089_reg/NET0131  & ~n5603 ;
  assign n7855 = ~\g1332_reg/NET0131  & n5603 ;
  assign n7856 = ~n7854 & ~n7855 ;
  assign n7857 = \g2093_reg/NET0131  & ~n5462 ;
  assign n7858 = ~\g1358_reg/NET0131  & n5462 ;
  assign n7859 = ~n7857 & ~n7858 ;
  assign n7860 = \g2095_reg/NET0131  & ~n5603 ;
  assign n7861 = ~\g1358_reg/NET0131  & n5603 ;
  assign n7862 = ~n7860 & ~n7861 ;
  assign n7863 = \g2097_reg/NET0131  & ~n5611 ;
  assign n7864 = ~\g1352_reg/NET0131  & n5611 ;
  assign n7865 = ~n7863 & ~n7864 ;
  assign n7866 = \g2099_reg/NET0131  & ~n5462 ;
  assign n7867 = ~\g1365_reg/NET0131  & n5462 ;
  assign n7868 = ~n7866 & ~n7867 ;
  assign n7869 = \g2100_reg/NET0131  & ~n5611 ;
  assign n7870 = ~\g1365_reg/NET0131  & n5611 ;
  assign n7871 = ~n7869 & ~n7870 ;
  assign n7872 = \g2101_reg/NET0131  & ~n5603 ;
  assign n7873 = ~\g1365_reg/NET0131  & n5603 ;
  assign n7874 = ~n7872 & ~n7873 ;
  assign n7875 = \g2102_reg/NET0131  & ~n5462 ;
  assign n7876 = ~\g1372_reg/NET0131  & n5462 ;
  assign n7877 = ~n7875 & ~n7876 ;
  assign n7878 = \g2104_reg/NET0131  & ~n5603 ;
  assign n7879 = ~\g1372_reg/NET0131  & n5603 ;
  assign n7880 = ~n7878 & ~n7879 ;
  assign n7881 = \g2106_reg/NET0131  & ~n5611 ;
  assign n7882 = ~\g1378_reg/NET0131  & n5611 ;
  assign n7883 = ~n7881 & ~n7882 ;
  assign n7884 = \g2107_reg/NET0131  & ~n5603 ;
  assign n7885 = ~\g1378_reg/NET0131  & n5603 ;
  assign n7886 = ~n7884 & ~n7885 ;
  assign n7887 = \g2091_reg/NET0131  & ~n5611 ;
  assign n7888 = ~\g1346_reg/NET0131  & n5611 ;
  assign n7889 = ~n7887 & ~n7888 ;
  assign n7890 = \g2090_reg/NET0131  & ~n5462 ;
  assign n7891 = ~\g1346_reg/NET0131  & n5462 ;
  assign n7892 = ~n7890 & ~n7891 ;
  assign n7893 = \g2086_reg/NET0131  & ~n5603 ;
  assign n7894 = ~\g1339_reg/NET0131  & n5603 ;
  assign n7895 = ~n7893 & ~n7894 ;
  assign n7896 = \g2788_reg/NET0131  & ~n5312 ;
  assign n7897 = ~\g1358_reg/NET0131  & n5312 ;
  assign n7898 = ~n7896 & ~n7897 ;
  assign n7899 = \g2105_reg/NET0131  & ~n5462 ;
  assign n7900 = ~\g1378_reg/NET0131  & n5462 ;
  assign n7901 = ~n7899 & ~n7900 ;
  assign n7902 = \g2088_reg/NET0131  & ~n5611 ;
  assign n7903 = ~\g1332_reg/NET0131  & n5611 ;
  assign n7904 = ~n7902 & ~n7903 ;
  assign n7905 = \g2098_reg/NET0131  & ~n5603 ;
  assign n7906 = ~\g1352_reg/NET0131  & n5603 ;
  assign n7907 = ~n7905 & ~n7906 ;
  assign n7908 = \g2094_reg/NET0131  & ~n5611 ;
  assign n7909 = ~\g1358_reg/NET0131  & n5611 ;
  assign n7910 = ~n7908 & ~n7909 ;
  assign n7911 = \g2772_reg/NET0131  & ~n5619 ;
  assign n7912 = ~\g1326_reg/NET0131  & n5619 ;
  assign n7913 = ~n7911 & ~n7912 ;
  assign n7914 = \g2773_reg/NET0131  & ~n5312 ;
  assign n7915 = ~\g1326_reg/NET0131  & n5312 ;
  assign n7916 = ~n7914 & ~n7915 ;
  assign n7917 = \g2774_reg/NET0131  & ~n5374 ;
  assign n7918 = ~\g1326_reg/NET0131  & n5374 ;
  assign n7919 = ~n7917 & ~n7918 ;
  assign n7920 = \g2775_reg/NET0131  & ~n5619 ;
  assign n7921 = ~\g1319_reg/NET0131  & n5619 ;
  assign n7922 = ~n7920 & ~n7921 ;
  assign n7923 = \g2776_reg/NET0131  & ~n5312 ;
  assign n7924 = ~\g1319_reg/NET0131  & n5312 ;
  assign n7925 = ~n7923 & ~n7924 ;
  assign n7926 = \g2777_reg/NET0131  & ~n5374 ;
  assign n7927 = ~\g1319_reg/NET0131  & n5374 ;
  assign n7928 = ~n7926 & ~n7927 ;
  assign n7929 = \g2778_reg/NET0131  & ~n5619 ;
  assign n7930 = ~\g1339_reg/NET0131  & n5619 ;
  assign n7931 = ~n7929 & ~n7930 ;
  assign n7932 = \g2779_reg/NET0131  & ~n5312 ;
  assign n7933 = ~\g1339_reg/NET0131  & n5312 ;
  assign n7934 = ~n7932 & ~n7933 ;
  assign n7935 = \g2780_reg/NET0131  & ~n5374 ;
  assign n7936 = ~\g1339_reg/NET0131  & n5374 ;
  assign n7937 = ~n7935 & ~n7936 ;
  assign n7938 = \g2781_reg/NET0131  & ~n5619 ;
  assign n7939 = ~\g1332_reg/NET0131  & n5619 ;
  assign n7940 = ~n7938 & ~n7939 ;
  assign n7941 = \g2782_reg/NET0131  & ~n5312 ;
  assign n7942 = ~\g1332_reg/NET0131  & n5312 ;
  assign n7943 = ~n7941 & ~n7942 ;
  assign n7944 = \g2783_reg/NET0131  & ~n5374 ;
  assign n7945 = ~\g1332_reg/NET0131  & n5374 ;
  assign n7946 = ~n7944 & ~n7945 ;
  assign n7947 = \g2784_reg/NET0131  & ~n5619 ;
  assign n7948 = ~\g1346_reg/NET0131  & n5619 ;
  assign n7949 = ~n7947 & ~n7948 ;
  assign n7950 = \g2785_reg/NET0131  & ~n5312 ;
  assign n7951 = ~\g1346_reg/NET0131  & n5312 ;
  assign n7952 = ~n7950 & ~n7951 ;
  assign n7953 = \g2786_reg/NET0131  & ~n5374 ;
  assign n7954 = ~\g1346_reg/NET0131  & n5374 ;
  assign n7955 = ~n7953 & ~n7954 ;
  assign n7956 = \g2787_reg/NET0131  & ~n5619 ;
  assign n7957 = ~\g1358_reg/NET0131  & n5619 ;
  assign n7958 = ~n7956 & ~n7957 ;
  assign n7959 = \g2789_reg/NET0131  & ~n5374 ;
  assign n7960 = ~\g1358_reg/NET0131  & n5374 ;
  assign n7961 = ~n7959 & ~n7960 ;
  assign n7962 = \g2790_reg/NET0131  & ~n5619 ;
  assign n7963 = ~\g1352_reg/NET0131  & n5619 ;
  assign n7964 = ~n7962 & ~n7963 ;
  assign n7965 = \g2791_reg/NET0131  & ~n5312 ;
  assign n7966 = ~\g1352_reg/NET0131  & n5312 ;
  assign n7967 = ~n7965 & ~n7966 ;
  assign n7968 = \g2792_reg/NET0131  & ~n5374 ;
  assign n7969 = ~\g1352_reg/NET0131  & n5374 ;
  assign n7970 = ~n7968 & ~n7969 ;
  assign n7971 = \g2793_reg/NET0131  & ~n5619 ;
  assign n7972 = ~\g1365_reg/NET0131  & n5619 ;
  assign n7973 = ~n7971 & ~n7972 ;
  assign n7974 = \g2096_reg/NET0131  & ~n5462 ;
  assign n7975 = ~\g1352_reg/NET0131  & n5462 ;
  assign n7976 = ~n7974 & ~n7975 ;
  assign n7977 = \g2794_reg/NET0131  & ~n5312 ;
  assign n7978 = ~\g1365_reg/NET0131  & n5312 ;
  assign n7979 = ~n7977 & ~n7978 ;
  assign n7980 = \g2795_reg/NET0131  & ~n5374 ;
  assign n7981 = ~\g1365_reg/NET0131  & n5374 ;
  assign n7982 = ~n7980 & ~n7981 ;
  assign n7983 = \g2796_reg/NET0131  & ~n5619 ;
  assign n7984 = ~\g1372_reg/NET0131  & n5619 ;
  assign n7985 = ~n7983 & ~n7984 ;
  assign n7986 = \g2797_reg/NET0131  & ~n5312 ;
  assign n7987 = ~\g1372_reg/NET0131  & n5312 ;
  assign n7988 = ~n7986 & ~n7987 ;
  assign n7989 = \g2798_reg/NET0131  & ~n5374 ;
  assign n7990 = ~\g1372_reg/NET0131  & n5374 ;
  assign n7991 = ~n7989 & ~n7990 ;
  assign n7992 = \g2799_reg/NET0131  & ~n5619 ;
  assign n7993 = ~\g1378_reg/NET0131  & n5619 ;
  assign n7994 = ~n7992 & ~n7993 ;
  assign n7995 = \g2800_reg/NET0131  & ~n5312 ;
  assign n7996 = ~\g1378_reg/NET0131  & n5312 ;
  assign n7997 = ~n7995 & ~n7996 ;
  assign n7998 = \g2801_reg/NET0131  & ~n5374 ;
  assign n7999 = ~\g1378_reg/NET0131  & n5374 ;
  assign n8000 = ~n7998 & ~n7999 ;
  assign n8001 = ~\g1164_reg/NET0131  & ~\g7961_pad  ;
  assign n8002 = ~n2470 & ~n8001 ;
  assign n8003 = n3456 & n8002 ;
  assign n8004 = \g1164_reg/NET0131  & ~\g7961_pad  ;
  assign n8005 = ~n8003 & ~n8004 ;
  assign n8006 = n7261 & n7812 ;
  assign n8007 = ~\g2900_reg/NET0131  & ~n8006 ;
  assign n8008 = ~n7817 & ~n8007 ;
  assign n8009 = n7809 & n8008 ;
  assign n8010 = \g2912_reg/NET0131  & \g2917_reg/NET0131  ;
  assign n8011 = n7264 & n8010 ;
  assign n8012 = ~\g2924_reg/NET0131  & ~n8011 ;
  assign n8013 = n7269 & ~n7274 ;
  assign n8014 = ~n8012 & n8013 ;
  assign n8015 = ~\g1319_reg/NET0131  & ~n7374 ;
  assign n8016 = ~n5997 & ~n6004 ;
  assign n8017 = ~n8015 & n8016 ;
  assign n8018 = ~\g2814_reg/NET0131  & ~\g2917_reg/NET0131  ;
  assign n8019 = \g2912_reg/NET0131  & n8018 ;
  assign n8020 = ~n7266 & n8019 ;
  assign n8021 = n7264 & n8020 ;
  assign n8022 = \g2912_reg/NET0131  & n7264 ;
  assign n8023 = ~\g2814_reg/NET0131  & \g2917_reg/NET0131  ;
  assign n8024 = ~n8022 & n8023 ;
  assign n8025 = ~n8021 & ~n8024 ;
  assign n8026 = ~\g2975_reg/NET0131  & ~\g2978_reg/NET0131  ;
  assign n8027 = \g2975_reg/NET0131  & \g2978_reg/NET0131  ;
  assign n8028 = ~n8026 & ~n8027 ;
  assign n8029 = \g2963_reg/NET0131  & ~\g2966_reg/NET0131  ;
  assign n8030 = ~n8028 & n8029 ;
  assign n8031 = \g2963_reg/NET0131  & \g2966_reg/NET0131  ;
  assign n8032 = n8028 & n8031 ;
  assign n8033 = ~n8030 & ~n8032 ;
  assign n8034 = ~\g2963_reg/NET0131  & \g2966_reg/NET0131  ;
  assign n8035 = ~n8028 & n8034 ;
  assign n8036 = ~\g2963_reg/NET0131  & ~\g2966_reg/NET0131  ;
  assign n8037 = n8028 & n8036 ;
  assign n8038 = ~n8035 & ~n8037 ;
  assign n8039 = n8033 & n8038 ;
  assign n8040 = \g2969_reg/NET0131  & ~\g2972_reg/NET0131  ;
  assign n8041 = ~\g2969_reg/NET0131  & \g2972_reg/NET0131  ;
  assign n8042 = ~n8040 & ~n8041 ;
  assign n8043 = \g3139_reg/NET0131  & ~\g3231_pad  ;
  assign n8044 = \g2874_reg/NET0131  & ~\g2981_reg/NET0131  ;
  assign n8045 = ~\g2874_reg/NET0131  & \g2981_reg/NET0131  ;
  assign n8046 = ~n8044 & ~n8045 ;
  assign n8047 = n8043 & n8046 ;
  assign n8048 = ~n8042 & n8047 ;
  assign n8049 = ~n8039 & n8048 ;
  assign n8050 = n8043 & ~n8046 ;
  assign n8051 = n8042 & n8050 ;
  assign n8052 = ~n8039 & n8051 ;
  assign n8053 = ~n8049 & ~n8052 ;
  assign n8054 = ~n8042 & n8050 ;
  assign n8055 = n8039 & n8054 ;
  assign n8056 = n8042 & n8047 ;
  assign n8057 = n8039 & n8056 ;
  assign n8058 = ~n8055 & ~n8057 ;
  assign n8059 = n8053 & n8058 ;
  assign n8060 = ~n8043 & ~n8046 ;
  assign n8061 = ~n8042 & n8060 ;
  assign n8062 = ~n8039 & n8061 ;
  assign n8063 = ~n8043 & n8046 ;
  assign n8064 = n8042 & n8063 ;
  assign n8065 = ~n8039 & n8064 ;
  assign n8066 = ~n8062 & ~n8065 ;
  assign n8067 = ~n8042 & n8063 ;
  assign n8068 = n8039 & n8067 ;
  assign n8069 = n8042 & n8060 ;
  assign n8070 = n8039 & n8069 ;
  assign n8071 = ~n8068 & ~n8070 ;
  assign n8072 = n8066 & n8071 ;
  assign n8073 = n8059 & n8072 ;
  assign n8074 = ~\g2935_reg/NET0131  & ~\g2938_reg/NET0131  ;
  assign n8075 = \g2935_reg/NET0131  & \g2938_reg/NET0131  ;
  assign n8076 = ~n8074 & ~n8075 ;
  assign n8077 = \g2959_reg/NET0131  & n8076 ;
  assign n8078 = ~\g2959_reg/NET0131  & ~n8076 ;
  assign n8079 = ~n8077 & ~n8078 ;
  assign n8080 = \g2941_reg/NET0131  & ~\g2944_reg/NET0131  ;
  assign n8081 = ~\g2941_reg/NET0131  & \g2944_reg/NET0131  ;
  assign n8082 = ~n8080 & ~n8081 ;
  assign n8083 = \g2956_reg/NET0131  & n8082 ;
  assign n8084 = ~\g2956_reg/NET0131  & ~n8082 ;
  assign n8085 = ~n8083 & ~n8084 ;
  assign n8086 = n8079 & n8085 ;
  assign n8087 = ~n8079 & ~n8085 ;
  assign n8088 = ~n8086 & ~n8087 ;
  assign n8089 = \g2947_reg/NET0131  & ~\g2953_reg/NET0131  ;
  assign n8090 = ~\g2947_reg/NET0131  & \g2953_reg/NET0131  ;
  assign n8091 = ~n8089 & ~n8090 ;
  assign n8092 = ~n8043 & ~n8091 ;
  assign n8093 = n8043 & n8091 ;
  assign n8094 = ~n8092 & ~n8093 ;
  assign n8095 = ~n8088 & n8094 ;
  assign n8096 = n8088 & ~n8094 ;
  assign n8097 = ~n8095 & ~n8096 ;
  assign n8098 = \g2934_reg/NET0131  & n8091 ;
  assign n8099 = n8088 & n8098 ;
  assign n8100 = \g2934_reg/NET0131  & ~n8091 ;
  assign n8101 = ~n8088 & n8100 ;
  assign n8102 = ~n8099 & ~n8101 ;
  assign n8103 = ~\g2934_reg/NET0131  & ~n8091 ;
  assign n8104 = n8088 & n8103 ;
  assign n8105 = ~\g2934_reg/NET0131  & n8091 ;
  assign n8106 = ~n8088 & n8105 ;
  assign n8107 = ~n8104 & ~n8106 ;
  assign n8108 = n8102 & n8107 ;
  assign n8109 = \g2962_reg/NET0131  & n8042 ;
  assign n8110 = ~n8046 & n8109 ;
  assign n8111 = ~n8039 & n8110 ;
  assign n8112 = n8046 & n8109 ;
  assign n8113 = n8039 & n8112 ;
  assign n8114 = ~n8111 & ~n8113 ;
  assign n8115 = \g2962_reg/NET0131  & n8046 ;
  assign n8116 = ~n8042 & n8115 ;
  assign n8117 = ~n8039 & n8116 ;
  assign n8118 = \g2962_reg/NET0131  & ~n8046 ;
  assign n8119 = ~n8042 & n8118 ;
  assign n8120 = n8039 & n8119 ;
  assign n8121 = ~n8117 & ~n8120 ;
  assign n8122 = n8114 & n8121 ;
  assign n8123 = ~\g2962_reg/NET0131  & ~n8046 ;
  assign n8124 = ~n8042 & n8123 ;
  assign n8125 = ~n8039 & n8124 ;
  assign n8126 = ~\g2962_reg/NET0131  & n8046 ;
  assign n8127 = ~n8042 & n8126 ;
  assign n8128 = n8039 & n8127 ;
  assign n8129 = ~n8125 & ~n8128 ;
  assign n8130 = ~\g2962_reg/NET0131  & n8042 ;
  assign n8131 = n8046 & n8130 ;
  assign n8132 = ~n8039 & n8131 ;
  assign n8133 = ~n8046 & n8130 ;
  assign n8134 = n8039 & n8133 ;
  assign n8135 = ~n8132 & ~n8134 ;
  assign n8136 = n8129 & n8135 ;
  assign n8137 = n8122 & n8136 ;
  assign n8138 = ~\g2814_reg/NET0131  & \g2912_reg/NET0131  ;
  assign n8139 = ~n7266 & n8138 ;
  assign n8140 = n7264 & n8139 ;
  assign n8141 = ~\g2814_reg/NET0131  & ~\g2912_reg/NET0131  ;
  assign n8142 = ~n7264 & n8141 ;
  assign n8143 = ~n8140 & ~n8142 ;
  assign n8144 = \g3002_reg/NET0131  & n7186 ;
  assign n8145 = ~\g3002_reg/NET0131  & ~n7186 ;
  assign n8146 = ~n8144 & ~n8145 ;
  assign n8147 = n7183 & n8146 ;
  assign n8148 = \g3080_reg/NET0131  & n7184 ;
  assign n8149 = \g2993_reg/NET0131  & \g3080_reg/NET0131  ;
  assign n8150 = ~\g2998_reg/NET0131  & ~n8149 ;
  assign n8151 = ~n8148 & ~n8150 ;
  assign n8152 = ~n7132 & n8151 ;
  assign n8153 = ~\g3234_pad  & ~n8152 ;
  assign n8154 = ~\g1869_reg/NET0131  & \g5657_pad  ;
  assign n8155 = \g1018_reg/NET0131  & ~\g1867_reg/NET0131  ;
  assign n8156 = \g1024_reg/NET0131  & ~\g1868_reg/NET0131  ;
  assign n8157 = ~n8155 & ~n8156 ;
  assign n8158 = ~n8154 & n8157 ;
  assign n8159 = ~\g488_reg/NET0131  & \g5657_pad  ;
  assign n8160 = \g1018_reg/NET0131  & ~\g486_reg/NET0131  ;
  assign n8161 = \g1024_reg/NET0131  & ~\g487_reg/NET0131  ;
  assign n8162 = ~n8160 & ~n8161 ;
  assign n8163 = ~n8159 & n8162 ;
  assign n8164 = ~\g1860_reg/NET0131  & \g5657_pad  ;
  assign n8165 = \g1018_reg/NET0131  & ~\g1858_reg/NET0131  ;
  assign n8166 = \g1024_reg/NET0131  & ~\g1859_reg/NET0131  ;
  assign n8167 = ~n8165 & ~n8166 ;
  assign n8168 = ~n8164 & n8167 ;
  assign n8169 = ~\g2920_reg/NET0131  & \g2924_reg/NET0131  ;
  assign n8170 = ~\g2912_reg/NET0131  & n8169 ;
  assign n8171 = \g2883_reg/NET0131  & ~\g2888_reg/NET0131  ;
  assign n8172 = \g1088_reg/NET0131  & ~\g2917_reg/NET0131  ;
  assign n8173 = n8171 & n8172 ;
  assign n8174 = n8170 & n8173 ;
  assign n8175 = n6243 & n8174 ;
  assign n8176 = \g856_reg/NET0131  & ~n8175 ;
  assign n8177 = ~\g805_reg/NET0131  & ~\g809_reg/NET0131  ;
  assign n8178 = n6034 & n8177 ;
  assign n8179 = n8175 & n8178 ;
  assign n8180 = ~n8176 & ~n8179 ;
  assign n8181 = ~\g2917_reg/NET0131  & \g7961_pad  ;
  assign n8182 = n8171 & n8181 ;
  assign n8183 = n8170 & n8182 ;
  assign n8184 = n6243 & n8183 ;
  assign n8185 = \g857_reg/NET0131  & ~n8184 ;
  assign n8186 = n8178 & n8184 ;
  assign n8187 = ~n8185 & ~n8186 ;
  assign n8188 = \g1092_reg/NET0131  & ~\g2917_reg/NET0131  ;
  assign n8189 = n8171 & n8188 ;
  assign n8190 = n8170 & n8189 ;
  assign n8191 = n6243 & n8190 ;
  assign n8192 = \g858_reg/NET0131  & ~n8191 ;
  assign n8193 = n8178 & n8191 ;
  assign n8194 = ~n8192 & ~n8193 ;
  assign n8195 = ~\g479_reg/NET0131  & \g5657_pad  ;
  assign n8196 = \g1018_reg/NET0131  & ~\g477_reg/NET0131  ;
  assign n8197 = \g1024_reg/NET0131  & ~\g478_reg/NET0131  ;
  assign n8198 = ~n8196 & ~n8197 ;
  assign n8199 = ~n8195 & n8198 ;
  assign n8200 = \g2244_reg/NET0131  & ~n8175 ;
  assign n8201 = ~\g2190_reg/NET0131  & ~\g2195_reg/NET0131  ;
  assign n8202 = n6096 & n8201 ;
  assign n8203 = n8175 & n8202 ;
  assign n8204 = ~n8200 & ~n8203 ;
  assign n8205 = \g2245_reg/NET0131  & ~n8184 ;
  assign n8206 = n8184 & n8202 ;
  assign n8207 = ~n8205 & ~n8206 ;
  assign n8208 = \g2246_reg/NET0131  & ~n8191 ;
  assign n8209 = n8191 & n8202 ;
  assign n8210 = ~n8208 & ~n8209 ;
  assign n8211 = ~\g1166_reg/NET0131  & \g5657_pad  ;
  assign n8212 = \g1024_reg/NET0131  & ~\g1165_reg/NET0131  ;
  assign n8213 = \g1018_reg/NET0131  & ~\g1164_reg/NET0131  ;
  assign n8214 = ~n8212 & ~n8213 ;
  assign n8215 = ~n8211 & n8214 ;
  assign n8216 = ~\g464_reg/NET0131  & \g5657_pad  ;
  assign n8217 = \g1018_reg/NET0131  & ~\g480_reg/NET0131  ;
  assign n8218 = \g1024_reg/NET0131  & ~\g484_reg/NET0131  ;
  assign n8219 = ~n8217 & ~n8218 ;
  assign n8220 = ~n8216 & n8219 ;
  assign n8221 = ~\g1151_reg/NET0131  & \g5657_pad  ;
  assign n8222 = \g1018_reg/NET0131  & ~\g1167_reg/NET0131  ;
  assign n8223 = \g1024_reg/NET0131  & ~\g1171_reg/NET0131  ;
  assign n8224 = ~n8222 & ~n8223 ;
  assign n8225 = ~n8221 & n8224 ;
  assign n8226 = ~\g1175_reg/NET0131  & \g5657_pad  ;
  assign n8227 = \g1018_reg/NET0131  & ~\g1173_reg/NET0131  ;
  assign n8228 = \g1024_reg/NET0131  & ~\g1174_reg/NET0131  ;
  assign n8229 = ~n8227 & ~n8228 ;
  assign n8230 = ~n8226 & n8229 ;
  assign n8231 = ~\g2993_reg/NET0131  & ~\g3080_reg/NET0131  ;
  assign n8232 = ~\g3234_pad  & ~n8149 ;
  assign n8233 = ~n8231 & n8232 ;
  assign n8234 = ~\g2554_reg/NET0131  & \g5657_pad  ;
  assign n8235 = \g1018_reg/NET0131  & ~\g2552_reg/NET0131  ;
  assign n8236 = \g1024_reg/NET0131  & ~\g2553_reg/NET0131  ;
  assign n8237 = ~n8235 & ~n8236 ;
  assign n8238 = ~n8234 & n8237 ;
  assign n8239 = ~\g2539_reg/NET0131  & \g5657_pad  ;
  assign n8240 = \g1018_reg/NET0131  & ~\g2555_reg/NET0131  ;
  assign n8241 = \g1024_reg/NET0131  & ~\g2559_reg/NET0131  ;
  assign n8242 = ~n8240 & ~n8241 ;
  assign n8243 = ~n8239 & n8242 ;
  assign n8244 = ~\g2563_reg/NET0131  & \g5657_pad  ;
  assign n8245 = \g1018_reg/NET0131  & ~\g2561_reg/NET0131  ;
  assign n8246 = \g1024_reg/NET0131  & ~\g2562_reg/NET0131  ;
  assign n8247 = ~n8245 & ~n8246 ;
  assign n8248 = ~n8244 & n8247 ;
  assign n8249 = ~\g1845_reg/NET0131  & \g5657_pad  ;
  assign n8250 = \g1018_reg/NET0131  & ~\g1861_reg/NET0131  ;
  assign n8251 = \g1024_reg/NET0131  & ~\g1865_reg/NET0131  ;
  assign n8252 = ~n8250 & ~n8251 ;
  assign n8253 = ~n8249 & n8252 ;
  assign n8254 = ~n6099 & n8175 ;
  assign n8255 = \g2253_reg/NET0131  & ~n8175 ;
  assign n8256 = ~n8254 & ~n8255 ;
  assign n8257 = ~n6099 & n8184 ;
  assign n8258 = \g2254_reg/NET0131  & ~n8184 ;
  assign n8259 = ~n8257 & ~n8258 ;
  assign n8260 = ~n6099 & n8191 ;
  assign n8261 = \g2255_reg/NET0131  & ~n8191 ;
  assign n8262 = ~n8260 & ~n8261 ;
  assign n8263 = ~\g3006_reg/NET0131  & ~n8148 ;
  assign n8264 = ~n7186 & ~n8263 ;
  assign n8265 = n7183 & n8264 ;
  assign n8266 = ~\g2883_reg/NET0131  & ~\g2950_reg/NET0131  ;
  assign n8267 = ~n7810 & ~n8266 ;
  assign n8268 = ~\g2814_reg/NET0131  & ~n8267 ;
  assign n8269 = ~n7264 & n8268 ;
  assign n8270 = \g2892_reg/NET0131  & n7812 ;
  assign n8271 = ~\g2892_reg/NET0131  & ~n7812 ;
  assign n8272 = ~n8270 & ~n8271 ;
  assign n8273 = n7809 & n8272 ;
  assign n8274 = ~\g2903_reg/NET0131  & ~n8270 ;
  assign n8275 = ~n8006 & ~n8274 ;
  assign n8276 = n7809 & n8275 ;
  assign n8277 = ~\g3013_reg/NET0131  & ~n8144 ;
  assign n8278 = ~n7774 & ~n8277 ;
  assign n8279 = n7183 & n8278 ;
  assign n8280 = ~\g1326_reg/NET0131  & ~n5382 ;
  assign n8281 = ~n6004 & ~n7374 ;
  assign n8282 = ~n8280 & n8281 ;
  assign n8283 = \g2888_reg/NET0131  & n7810 ;
  assign n8284 = ~\g2888_reg/NET0131  & ~n7810 ;
  assign n8285 = ~n8283 & ~n8284 ;
  assign n8286 = n7809 & n8285 ;
  assign n8287 = ~\g2896_reg/NET0131  & ~n8283 ;
  assign n8288 = ~n7812 & ~n8287 ;
  assign n8289 = n7809 & n8288 ;
  assign n8290 = ~\g2933_reg/NET0131  & ~\g51_pad  ;
  assign n8291 = ~\g2917_reg/NET0131  & n8171 ;
  assign n8292 = n8170 & n8291 ;
  assign n8293 = n6243 & n8292 ;
  assign n8294 = ~\g3079_reg/NET0131  & ~\g3234_pad  ;
  assign n8295 = ~\g1024_reg/NET0131  & \g1345_reg/NET0131  ;
  assign n8296 = ~\g1024_reg/NET0131  & ~\g1345_reg/NET0131  ;
  assign n8297 = n6706 & ~n8296 ;
  assign n8298 = n6708 & n8297 ;
  assign n8299 = ~n8295 & ~n8298 ;
  assign n8300 = \g1024_reg/NET0131  & ~\g1240_reg/NET0131  ;
  assign n8301 = ~\g1024_reg/NET0131  & \g1243_reg/NET0131  ;
  assign n8302 = ~n8300 & ~n8301 ;
  assign n8303 = ~\g291_reg/NET0131  & \g3229_pad  ;
  assign n8304 = \g305_reg/NET0131  & ~\g3229_pad  ;
  assign n8305 = ~n8303 & ~n8304 ;
  assign n8306 = \g3229_pad  & ~\g978_reg/NET0131  ;
  assign n8307 = ~\g3229_pad  & \g992_reg/NET0131  ;
  assign n8308 = ~n8306 & ~n8307 ;
  assign n8309 = \g2814_reg/NET0131  & ~\g2929_reg/NET0131  ;
  assign n8310 = \g2879_reg/NET0131  & ~n8309 ;
  assign n8311 = ~\g1672_reg/NET0131  & \g3229_pad  ;
  assign n8312 = \g1686_reg/NET0131  & ~\g3229_pad  ;
  assign n8313 = ~n8311 & ~n8312 ;
  assign n8314 = ~\g2366_reg/NET0131  & \g3229_pad  ;
  assign n8315 = \g2380_reg/NET0131  & ~\g3229_pad  ;
  assign n8316 = ~n8314 & ~n8315 ;
  assign n8317 = \g2817_reg/NET0131  & ~\g51_pad  ;
  assign n8318 = \g3054_reg/NET0131  & ~\g3234_pad  ;
  assign n8319 = ~\g117_reg/NET0131  & ~\g121_reg/NET0131  ;
  assign n8320 = n6065 & n8319 ;
  assign n8321 = ~\g1496_reg/NET0131  & ~\g1501_reg/NET0131  ;
  assign n8322 = n6127 & n8321 ;
  assign n8323 = \g2950_reg/NET0131  & ~\g51_pad  ;
  assign n8324 = \g3080_reg/NET0131  & ~\g3234_pad  ;
  assign n8325 = \g121_reg/NET0131  & ~n3411 ;
  assign n8326 = \g121_reg/NET0131  & n3406 ;
  assign n8327 = ~n3400 & n8326 ;
  assign n8328 = ~n8325 & ~n8327 ;
  assign n8329 = ~n4081 & ~n4085 ;
  assign n8330 = ~n4080 & n8329 ;
  assign n8331 = n3989 & n8330 ;
  assign n8332 = ~n2349 & ~n8331 ;
  assign n8333 = n2349 & ~n4085 ;
  assign n8334 = ~n4081 & n8333 ;
  assign n8335 = ~n4080 & n8334 ;
  assign n8336 = n3989 & n8335 ;
  assign n8337 = ~n8332 & ~n8336 ;
  assign n8338 = ~n3430 & ~n8337 ;
  assign n8339 = n3411 & n8338 ;
  assign n8340 = ~n3410 & n8339 ;
  assign n8341 = n8328 & ~n8340 ;
  assign n8342 = ~n1752 & ~n4425 ;
  assign n8343 = \g2190_reg/NET0131  & ~n3739 ;
  assign n8344 = n3807 & ~n3809 ;
  assign n8345 = n3867 & n8344 ;
  assign n8346 = n1212 & ~n8345 ;
  assign n8347 = n1234 & n1254 ;
  assign n8348 = ~n1212 & n8347 ;
  assign n8349 = ~n3705 & n8348 ;
  assign n8350 = ~n1234 & ~n1254 ;
  assign n8351 = ~n1212 & n8350 ;
  assign n8352 = n3705 & n8351 ;
  assign n8353 = ~n8349 & ~n8352 ;
  assign n8354 = n8344 & ~n8353 ;
  assign n8355 = ~n8346 & ~n8354 ;
  assign n8356 = n3859 & n8355 ;
  assign n8357 = ~n3694 & n8356 ;
  assign n8358 = ~n8343 & ~n8357 ;
  assign n8359 = ~\g1088_reg/NET0131  & ~\g246_reg/NET0131  ;
  assign n8360 = ~\g1088_reg/NET0131  & ~n8359 ;
  assign n8361 = ~n3410 & n3976 ;
  assign n8362 = ~n3974 & ~n8361 ;
  assign n8363 = ~n3995 & ~n8359 ;
  assign n8364 = ~n8362 & n8363 ;
  assign n8365 = ~n8360 & ~n8364 ;
  assign \_al_n0  = 1'b0 ;
  assign \_al_n1  = ~1'b0 ;
  assign \g101_reg/P0001  = ~\g101_reg/NET0131  ;
  assign \g105_reg/P0001  = ~\g105_reg/NET0131  ;
  assign \g109_reg/P0001  = ~\g109_reg/NET0131  ;
  assign \g1138_reg/P0001  = ~\g1138_reg/NET0131  ;
  assign \g113_reg/P0001  = ~\g113_reg/NET0131  ;
  assign \g1140_reg/P0001  = ~\g1140_reg/NET0131  ;
  assign \g117_reg/P0001  = ~\g117_reg/NET0131  ;
  assign \g121_reg/P0001  = ~\g121_reg/NET0131  ;
  assign \g125_reg/P0001  = ~\g125_reg/NET0131  ;
  assign \g1471_reg/P0001  = ~\g1471_reg/NET0131  ;
  assign \g1476_reg/P0001  = ~\g1476_reg/NET0131  ;
  assign \g1481_reg/P0001  = ~\g1481_reg/NET0131  ;
  assign \g1486_reg/P0001  = ~\g1486_reg/NET0131  ;
  assign \g1491_reg/P0001  = ~\g1491_reg/NET0131  ;
  assign \g1496_reg/P0001  = ~\g1496_reg/NET0131  ;
  assign \g1501_reg/P0001  = ~\g1501_reg/NET0131  ;
  assign \g1506_reg/P0001  = ~\g1506_reg/NET0131  ;
  assign \g16496_pad  = ~n1181 ;
  assign \g1660_reg/P0001  = ~\g1660_reg/NET0131  ;
  assign \g1662_reg/P0001  = ~\g1662_reg/NET0131  ;
  assign \g1664_reg/P0001  = ~\g1664_reg/NET0131  ;
  assign \g1666_reg/P0001  = ~\g1666_reg/NET0131  ;
  assign \g1668_reg/P0001  = ~\g1668_reg/NET0131  ;
  assign \g1670_reg/P0001  = ~\g1670_reg/NET0131  ;
  assign \g1672_reg/P0001  = ~\g1672_reg/NET0131  ;
  assign \g18/_0_  = n1476 ;
  assign \g1832_reg/P0001  = ~\g1832_reg/NET0131  ;
  assign \g1834_reg/P0001  = ~\g1834_reg/NET0131  ;
  assign \g2165_reg/P0001  = ~\g2165_reg/NET0131  ;
  assign \g2170_reg/P0001  = ~\g2170_reg/NET0131  ;
  assign \g2175_reg/P0001  = ~\g2175_reg/NET0131  ;
  assign \g2180_reg/P0001  = ~\g2180_reg/NET0131  ;
  assign \g2185_reg/P0001  = ~\g2185_reg/NET0131  ;
  assign \g2190_reg/P0001  = ~\g2190_reg/NET0131  ;
  assign \g2195_reg/P0001  = ~\g2195_reg/NET0131  ;
  assign \g2200_reg/P0001  = ~\g2200_reg/NET0131  ;
  assign \g2354_reg/P0001  = ~\g2354_reg/NET0131  ;
  assign \g2356_reg/P0001  = ~\g2356_reg/NET0131  ;
  assign \g2358_reg/P0001  = ~\g2358_reg/NET0131  ;
  assign \g2360_reg/P0001  = ~\g2360_reg/NET0131  ;
  assign \g2362_reg/P0001  = ~\g2362_reg/NET0131  ;
  assign \g2364_reg/P0001  = ~\g2364_reg/NET0131  ;
  assign \g2366_reg/P0001  = ~\g2366_reg/NET0131  ;
  assign \g2526_reg/P0001  = ~\g2526_reg/NET0131  ;
  assign \g2528_reg/P0001  = ~\g2528_reg/NET0131  ;
  assign \g25489_pad  = n1488 ;
  assign \g279_reg/P0001  = ~\g279_reg/NET0131  ;
  assign \g281_reg/P0001  = ~\g281_reg/NET0131  ;
  assign \g283_reg/P0001  = ~\g283_reg/NET0131  ;
  assign \g285_reg/P0001  = ~\g285_reg/NET0131  ;
  assign \g2879_reg/NET0131_syn_2  = ~\g2879_reg/NET0131  ;
  assign \g287_reg/P0001  = ~\g287_reg/NET0131  ;
  assign \g289_reg/P0001  = ~\g289_reg/NET0131  ;
  assign \g291_reg/P0001  = ~\g291_reg/NET0131  ;
  assign \g451_reg/P0001  = ~\g451_reg/NET0131  ;
  assign \g453_reg/P0001  = ~\g453_reg/NET0131  ;
  assign \g59421/_3_  = n1493 ;
  assign \g59425/_1_  = ~n1497 ;
  assign \g59435/_0_  = ~n1526 ;
  assign \g59436/_0_  = n1538 ;
  assign \g59441/_3_  = ~n1541 ;
  assign \g59442/_0_  = ~n1570 ;
  assign \g59445/_0_  = ~n1581 ;
  assign \g59453/_0_  = ~n1786 ;
  assign \g59462/_3_  = ~n1789 ;
  assign \g59466/_3_  = ~n1792 ;
  assign \g59467/_3_  = ~n1795 ;
  assign \g59468/_3_  = ~n1798 ;
  assign \g59469/_3_  = ~n1801 ;
  assign \g59470/_3_  = ~n1804 ;
  assign \g59471/_3_  = ~n1807 ;
  assign \g59472/_3_  = ~n1810 ;
  assign \g59473/_3_  = ~n1813 ;
  assign \g59489/_0_  = ~n2004 ;
  assign \g59498/_0_  = ~n2030 ;
  assign \g59499/_0_  = ~n2038 ;
  assign \g59500/_0_  = ~n2048 ;
  assign \g59502/_2_  = ~n2059 ;
  assign \g59503/_0_  = ~n2067 ;
  assign \g59505/_2_  = ~n2075 ;
  assign \g59507/_0_  = ~n2085 ;
  assign \g59508/_0_  = n2096 ;
  assign \g59533/_3_  = ~n2099 ;
  assign \g59534/_3_  = ~n2102 ;
  assign \g59535/_3_  = ~n2105 ;
  assign \g59536/_3_  = ~n2108 ;
  assign \g59537/_3_  = ~n2111 ;
  assign \g59538/_3_  = ~n2114 ;
  assign \g59539/_3_  = ~n2117 ;
  assign \g59540/_3_  = ~n2120 ;
  assign \g59548/_0_  = ~n2140 ;
  assign \g59550/_0_  = ~n2435 ;
  assign \g59551/_0_  = ~n2441 ;
  assign \g59552/_0_  = ~n2447 ;
  assign \g59554/_0_  = ~n2756 ;
  assign \g59555/_0_  = n2760 ;
  assign \g59556/_0_  = n2764 ;
  assign \g59557/_0_  = ~n2769 ;
  assign \g59558/_0_  = ~n2774 ;
  assign \g59559/_0_  = n3076 ;
  assign \g59560/_0_  = n3084 ;
  assign \g59561/_0_  = n3092 ;
  assign \g59639/_0_  = ~n3291 ;
  assign \g59694/_2_  = n3318 ;
  assign \g59695/_0_  = n3329 ;
  assign \g59697/_2_  = n3340 ;
  assign \g59698/_0_  = n3351 ;
  assign \g59699/_0_  = ~n3365 ;
  assign \g59700/_0_  = ~n3373 ;
  assign \g59705/_0_  = n3441 ;
  assign \g59706/_0_  = n3444 ;
  assign \g59707/_0_  = n3447 ;
  assign \g59708/_0_  = n3503 ;
  assign \g59709/_0_  = n3509 ;
  assign \g59710/_0_  = n3515 ;
  assign \g59711/_0_  = n3533 ;
  assign \g59712/_0_  = n3539 ;
  assign \g59713/_0_  = n3545 ;
  assign \g59714/_0_  = n3564 ;
  assign \g59715/_0_  = n3570 ;
  assign \g59716/_0_  = n3576 ;
  assign \g59717/_0_  = ~n3619 ;
  assign \g59718/_0_  = ~n3624 ;
  assign \g59719/_0_  = ~n3629 ;
  assign \g59720/_0_  = n3685 ;
  assign \g59721/_0_  = n3744 ;
  assign \g59722/_0_  = n3750 ;
  assign \g59723/_0_  = n3756 ;
  assign \g59724/_0_  = n3762 ;
  assign \g59725/_0_  = n3780 ;
  assign \g59726/_0_  = n3786 ;
  assign \g59727/_0_  = n3792 ;
  assign \g59728/_0_  = n3798 ;
  assign \g59729/_0_  = n3822 ;
  assign \g59730/_0_  = n3828 ;
  assign \g59731/_0_  = n3845 ;
  assign \g59732/_0_  = n3851 ;
  assign \g59733/_0_  = ~n3894 ;
  assign \g59734/_0_  = ~n3899 ;
  assign \g59735/_0_  = ~n3904 ;
  assign \g59736/_0_  = n3907 ;
  assign \g59737/_0_  = n3910 ;
  assign \g59738/_0_  = n3926 ;
  assign \g59739/_0_  = n3932 ;
  assign \g59740/_0_  = n3938 ;
  assign \g59741/_0_  = n3962 ;
  assign \g59742/_0_  = n3968 ;
  assign \g59743/_0_  = n3999 ;
  assign \g59744/_0_  = n4005 ;
  assign \g59745/_0_  = n4014 ;
  assign \g59747/_0_  = ~n4055 ;
  assign \g59748/_0_  = ~n4060 ;
  assign \g59749/_0_  = ~n4065 ;
  assign \g59750/_0_  = ~n4108 ;
  assign \g59751/_0_  = ~n4113 ;
  assign \g59752/_0_  = ~n4118 ;
  assign \g59753/_0_  = ~n4128 ;
  assign \g59754/_0_  = n4139 ;
  assign \g59755/_0_  = ~n4154 ;
  assign \g59756/_0_  = ~n4159 ;
  assign \g59757/_0_  = ~n4164 ;
  assign \g59758/_0_  = ~n4181 ;
  assign \g59759/_0_  = ~n4186 ;
  assign \g59760/_0_  = ~n4191 ;
  assign \g59761/_0_  = n4202 ;
  assign \g59762/_0_  = n4205 ;
  assign \g59763/_0_  = n4208 ;
  assign \g59764/_0_  = ~n4223 ;
  assign \g59765/_0_  = ~n4228 ;
  assign \g59766/_0_  = ~n4233 ;
  assign \g59915/_0_  = ~n4437 ;
  assign \g59952/_2_  = n4441 ;
  assign \g60046/_0_  = n4453 ;
  assign \g60048/_0_  = n4468 ;
  assign \g60049/_0_  = n4481 ;
  assign \g60051/_0_  = n4497 ;
  assign \g60063/_0_  = ~n4514 ;
  assign \g60103/_0_  = ~n4521 ;
  assign \g60104/_0_  = n4534 ;
  assign \g60105/_0_  = ~n4560 ;
  assign \g60107/_2_  = ~n4576 ;
  assign \g60108/_0_  = ~n4583 ;
  assign \g60109/_0_  = n4595 ;
  assign \g60110/_0_  = n4602 ;
  assign \g60112/_2_  = ~n4609 ;
  assign \g60119/_0_  = ~n4619 ;
  assign \g60120/_0_  = n4634 ;
  assign \g60121/_0_  = n4651 ;
  assign \g60122/_0_  = ~n4659 ;
  assign \g60123/_0_  = ~n4666 ;
  assign \g60124/_0_  = ~n4676 ;
  assign \g60126/_0_  = ~n4684 ;
  assign \g60127/_0_  = n4700 ;
  assign \g60128/_0_  = ~n4709 ;
  assign \g60129/_0_  = ~n4717 ;
  assign \g60130/_0_  = ~n4731 ;
  assign \g60135/_0_  = n4743 ;
  assign \g60136/_0_  = ~n4753 ;
  assign \g60137/_0_  = ~n4762 ;
  assign \g60138/_0_  = ~n4771 ;
  assign \g60139/_0_  = ~n4784 ;
  assign \g60143/_3_  = ~n4785 ;
  assign \g60144/_0_  = ~n4798 ;
  assign \g60145/_0_  = n4808 ;
  assign \g60339/_0_  = ~n4809 ;
  assign \g60404/_0_  = n4814 ;
  assign \g60427/_0_  = ~n4819 ;
  assign \g60428/_0_  = ~n4825 ;
  assign \g60429/_0_  = n4832 ;
  assign \g60434/_0_  = n4856 ;
  assign \g60435/_0_  = n4866 ;
  assign \g60437/_0_  = n4876 ;
  assign \g60438/_0_  = n4886 ;
  assign \g60439/_0_  = n4895 ;
  assign \g60440/_0_  = n4902 ;
  assign \g60441/_0_  = ~n4903 ;
  assign \g60448/_0_  = n5064 ;
  assign \g60451/_0_  = n5217 ;
  assign \g60452/_0_  = n5226 ;
  assign \g60453/_0_  = n5232 ;
  assign \g60459/_0_  = ~n5241 ;
  assign \g60460/_0_  = n5251 ;
  assign \g60523/_0_  = ~n5252 ;
  assign \g60534/_0_  = n5267 ;
  assign \g60535/_0_  = n5272 ;
  assign \g60536/_0_  = n5277 ;
  assign \g60585/_0_  = ~n5286 ;
  assign \g60586/_0_  = ~n5294 ;
  assign \g60587/_0_  = n5304 ;
  assign \g60588/_0_  = n5309 ;
  assign \g60591/_0_  = n5372 ;
  assign \g60592/_0_  = n5380 ;
  assign \g60599/_0_  = n5443 ;
  assign \g60601/_0_  = n5451 ;
  assign \g60602/_0_  = n5459 ;
  assign \g60603/_0_  = n5522 ;
  assign \g60604/_0_  = n5585 ;
  assign \g60605/_0_  = n5593 ;
  assign \g60606/_0_  = n5601 ;
  assign \g60607/_0_  = n5609 ;
  assign \g60608/_0_  = n5617 ;
  assign \g60609/_0_  = n5625 ;
  assign \g60613/_0_  = ~n5771 ;
  assign \g60614/_0_  = ~n5917 ;
  assign \g60615/_0_  = n5920 ;
  assign \g60694/_0_  = ~n5923 ;
  assign \g60708/_0_  = ~n5933 ;
  assign \g60709/_0_  = ~n5944 ;
  assign \g60710/_0_  = ~n5951 ;
  assign \g60785/_0_  = n5957 ;
  assign \g60787/_0_  = n5959 ;
  assign \g60788/_0_  = n5961 ;
  assign \g60799/_0_  = n5966 ;
  assign \g60801/_0_  = n5968 ;
  assign \g60802/_0_  = n5970 ;
  assign \g60803/_1__syn_2  = n5977 ;
  assign \g60805/_1__syn_2  = n5979 ;
  assign \g60806/_1__syn_2  = n5981 ;
  assign \g60808/_0_  = n5986 ;
  assign \g60810/_0_  = n5987 ;
  assign \g60811/_0_  = n5988 ;
  assign \g60825/_3_  = n5993 ;
  assign \g60896/_0_  = n6010 ;
  assign \g60980/_0_  = ~n6041 ;
  assign \g60981/_0_  = ~n6072 ;
  assign \g60985/_0_  = ~n6103 ;
  assign \g60986/_0_  = ~n6134 ;
  assign \g61012/_0_  = ~n6137 ;
  assign \g61013/_0_  = ~n6138 ;
  assign \g61015/_0_  = ~n6141 ;
  assign \g61017/_0_  = ~n6143 ;
  assign \g61122/_0_  = ~n6152 ;
  assign \g61123/_0_  = ~n6161 ;
  assign \g61124/_0_  = ~n6170 ;
  assign \g61125/_0_  = ~n6179 ;
  assign \g61222/_0_  = n6180 ;
  assign \g61223/_0_  = n6181 ;
  assign \g61224/_0_  = n6182 ;
  assign \g61225/_0_  = n6183 ;
  assign \g61228/_0_  = n6184 ;
  assign \g61229/_0_  = n6185 ;
  assign \g61230/_0_  = n6186 ;
  assign \g61231/_0_  = n6187 ;
  assign \g61281/_0_  = ~n6193 ;
  assign \g61293/_1_  = ~n6195 ;
  assign \g61307/_0__syn_2  = n6197 ;
  assign \g61309/_0__syn_2  = n6199 ;
  assign \g61310/_0__syn_2  = n6201 ;
  assign \g61311/_1_  = n6203 ;
  assign \g61312/_1_  = n6205 ;
  assign \g61313/_1_  = n6207 ;
  assign \g61324/_1_  = n6209 ;
  assign \g61325/_1_  = n6211 ;
  assign \g61326/_1_  = n6213 ;
  assign \g61328/_1_  = n6215 ;
  assign \g61329/_1_  = n6217 ;
  assign \g61330/_1_  = n6219 ;
  assign \g61332/_1_  = n6282 ;
  assign \g61333/_1_  = n6339 ;
  assign \g61334/_1_  = n6396 ;
  assign \g61335/_1_  = n6453 ;
  assign \g61336/_0_  = n6469 ;
  assign \g61338/_0_  = n6485 ;
  assign \g61339/_0_  = n6494 ;
  assign \g61340/_0_  = n6501 ;
  assign \g61377/_1_  = n6529 ;
  assign \g61378/_1_  = n6530 ;
  assign \g61379/_1_  = n6531 ;
  assign \g61388/_1_  = n6565 ;
  assign \g61391/_0_  = n6584 ;
  assign \g61394/_1_  = n6585 ;
  assign \g61395/_1_  = n6586 ;
  assign \g61396/_1_  = n6612 ;
  assign \g61398/_1_  = n6613 ;
  assign \g61399/_1_  = n6614 ;
  assign \g61421/_1_  = n6648 ;
  assign \g61422/_1_  = n6649 ;
  assign \g61423/_1_  = n6650 ;
  assign \g61524/_0_  = ~n6681 ;
  assign \g61525/_0_  = ~n6688 ;
  assign \g61526/_0_  = ~n6695 ;
  assign \g61527/_0_  = ~n6722 ;
  assign \g61528/_0_  = ~n6729 ;
  assign \g61529/_0_  = ~n6736 ;
  assign \g61530/_0_  = ~n6772 ;
  assign \g61531/_0_  = ~n6778 ;
  assign \g61532/_0_  = ~n6784 ;
  assign \g61533/_0_  = ~n6795 ;
  assign \g61534/_0_  = ~n6798 ;
  assign \g61535/_0_  = ~n6801 ;
  assign \g61536/_0_  = ~n6823 ;
  assign \g61537/_0_  = ~n6829 ;
  assign \g61538/_0_  = ~n6835 ;
  assign \g61539/_0_  = n6838 ;
  assign \g61540/_0_  = ~n6859 ;
  assign \g61541/_0_  = ~n6865 ;
  assign \g61542/_0_  = ~n6871 ;
  assign \g61543/_0_  = ~n6881 ;
  assign \g61544/_0_  = ~n6916 ;
  assign \g61545/_0_  = ~n6919 ;
  assign \g61546/_0_  = ~n6922 ;
  assign \g61547/_0_  = ~n6928 ;
  assign \g61548/_0_  = ~n6934 ;
  assign \g61549/_0_  = ~n6945 ;
  assign \g61550/_0_  = ~n6948 ;
  assign \g61551/_0_  = ~n6951 ;
  assign \g61552/_0_  = ~n6967 ;
  assign \g61553/_0_  = ~n6988 ;
  assign \g61554/_0_  = ~n7024 ;
  assign \g61555/_0_  = ~n7030 ;
  assign \g61556/_0_  = ~n7036 ;
  assign \g61557/_0_  = ~n7052 ;
  assign \g61558/_0_  = ~n7055 ;
  assign \g61559/_0_  = ~n7058 ;
  assign \g61560/_0_  = ~n7064 ;
  assign \g61561/_0_  = ~n7070 ;
  assign \g61562/_0_  = ~n7081 ;
  assign \g61563/_0_  = ~n7084 ;
  assign \g61564/_0_  = ~n7087 ;
  assign \g61565/_0_  = ~n7090 ;
  assign \g61566/_0_  = ~n7093 ;
  assign \g61620/_0_  = ~n7099 ;
  assign \g61621/_0_  = ~n7105 ;
  assign \g61622/_0_  = n7113 ;
  assign \g61623/_0_  = n7121 ;
  assign \g61753/_0_  = ~n7123 ;
  assign \g61764/_0_  = ~n7125 ;
  assign \g61786/_0_  = ~n7127 ;
  assign \g61795/_0_  = ~n7129 ;
  assign \g61801/_0_  = ~n7142 ;
  assign \g61803/_0_  = n7144 ;
  assign \g61808/_0_  = n7146 ;
  assign \g61848/_0_  = n7150 ;
  assign \g61850/_0_  = n7154 ;
  assign \g61851/_0_  = n7157 ;
  assign \g62097/_0_  = n7167 ;
  assign \g62102/_0_  = n7171 ;
  assign \g62115/_0_  = n7176 ;
  assign \g62119/_0_  = ~n6522 ;
  assign \g62130/_1_  = ~n6781 ;
  assign \g62131/_0_  = n7182 ;
  assign \g62132/_0_  = n7195 ;
  assign \g62139/_1_  = ~n6826 ;
  assign \g62140/_1_  = ~n6712 ;
  assign \g62141/_1_  = ~n6726 ;
  assign \g62144/_0_  = n7208 ;
  assign \g62145/_0_  = ~n7215 ;
  assign \g62146/_0_  = n7220 ;
  assign \g62147/_0_  = ~n7225 ;
  assign \g62150/_0_  = n7233 ;
  assign \g62151/_1_  = ~n6740 ;
  assign \g62152/_0_  = n7240 ;
  assign \g62153/_1_  = ~n6775 ;
  assign \g62156/_1_  = ~n6733 ;
  assign \g62157/_0_  = ~n6559 ;
  assign \g62159/_0_  = ~n6605 ;
  assign \g62161/_0_  = n7254 ;
  assign \g62187/_1_  = ~n6850 ;
  assign \g62190/_1_  = ~n6862 ;
  assign \g62191/_1_  = ~n6813 ;
  assign \g62192/_1_  = ~n6868 ;
  assign \g62194/_1_  = ~n6884 ;
  assign \g62195/_1_  = ~n6925 ;
  assign \g62196/_1_  = ~n6931 ;
  assign \g62203/_0_  = ~n6642 ;
  assign \g62204/_1_  = ~n6832 ;
  assign \g62207/_0__syn_2  = ~n6979 ;
  assign \g62208/_1_  = ~n6992 ;
  assign \g62209/_1_  = ~n7027 ;
  assign \g62210/_1_  = ~n7033 ;
  assign \g62211/_1_  = ~n7061 ;
  assign \g62212/_1_  = ~n7067 ;
  assign \g62217/_0_  = n7258 ;
  assign \g62286/_0_  = n7279 ;
  assign \g62287/_0_  = n7281 ;
  assign \g62288/_0_  = n7284 ;
  assign \g62289/_0_  = n7287 ;
  assign \g62290/_0_  = n7289 ;
  assign \g62291/_0_  = n7291 ;
  assign \g62292/_0_  = n7293 ;
  assign \g62435/_0_  = n7297 ;
  assign \g62436/_0_  = n7300 ;
  assign \g62439/_0_  = n7307 ;
  assign \g62456/_0_  = ~n7315 ;
  assign \g62486/_1_  = ~n6654 ;
  assign \g62492/_1_  = ~n6685 ;
  assign \g62494/_0_  = n7320 ;
  assign \g62495/_1_  = ~n6692 ;
  assign \g62497/_0_  = ~n7325 ;
  assign \g62537/_0_  = n7332 ;
  assign \g62544/_0_  = ~n7334 ;
  assign \g62546/_0_  = ~n7336 ;
  assign \g62547/_0_  = ~n7338 ;
  assign \g62549/_3_  = ~n7340 ;
  assign \g62552/_0_  = ~n7341 ;
  assign \g62554/_0_  = n7348 ;
  assign \g62555/_0_  = ~n7349 ;
  assign \g62556/_0_  = n7356 ;
  assign \g62558/_0_  = n7363 ;
  assign \g62559/_0_  = ~n7364 ;
  assign \g62561/_0_  = n7371 ;
  assign \g62562/_0_  = ~n7372 ;
  assign \g62566/_0_  = n7376 ;
  assign \g62567/_0_  = ~n7379 ;
  assign \g62568/_0_  = n7381 ;
  assign \g62569/_0_  = ~n7384 ;
  assign \g62570/_0_  = n7386 ;
  assign \g62571/_0_  = ~n7389 ;
  assign \g62572/_0_  = ~n7392 ;
  assign \g62573/_0_  = ~n7395 ;
  assign \g62574/_0_  = ~n7398 ;
  assign \g62575/_0_  = ~n7401 ;
  assign \g62576/_0_  = ~n7404 ;
  assign \g62577/_0_  = ~n7407 ;
  assign \g62578/_0_  = ~n7410 ;
  assign \g62579/_0_  = ~n7413 ;
  assign \g62580/_0_  = ~n7416 ;
  assign \g62581/_0_  = ~n7419 ;
  assign \g62582/_0_  = ~n7422 ;
  assign \g62583/_0_  = ~n7425 ;
  assign \g62584/_0_  = ~n7428 ;
  assign \g62585/_0_  = ~n7431 ;
  assign \g62586/_0_  = ~n7434 ;
  assign \g62587/_0_  = ~n7437 ;
  assign \g62588/_0_  = ~n7440 ;
  assign \g62589/_0_  = ~n7443 ;
  assign \g62590/_0_  = ~n7446 ;
  assign \g62591/_0_  = ~n7449 ;
  assign \g62592/_0_  = ~n7452 ;
  assign \g62593/_0_  = ~n7455 ;
  assign \g62594/_0_  = ~n7458 ;
  assign \g62595/_0_  = ~n7461 ;
  assign \g62596/_0_  = ~n7464 ;
  assign \g62597/_0_  = ~n7467 ;
  assign \g62602/_0_  = ~n7470 ;
  assign \g62607/_0_  = ~n7473 ;
  assign \g62608/_0_  = ~n7476 ;
  assign \g62609/_0_  = ~n7479 ;
  assign \g62619/_0_  = ~n7482 ;
  assign \g62620/_0_  = ~n7485 ;
  assign \g62621/_0_  = ~n7488 ;
  assign \g62622/_0_  = ~n7491 ;
  assign \g62623/_0_  = ~n7494 ;
  assign \g62624/_0_  = ~n7497 ;
  assign \g62626/_0_  = ~n7500 ;
  assign \g62627/_0_  = ~n7503 ;
  assign \g62628/_0_  = ~n7506 ;
  assign \g62629/_0_  = ~n7509 ;
  assign \g62630/_0_  = ~n7512 ;
  assign \g62631/_0_  = ~n7515 ;
  assign \g62632/_0_  = ~n7518 ;
  assign \g62633/_0_  = ~n7521 ;
  assign \g62634/_0_  = ~n7524 ;
  assign \g62635/_0_  = ~n7527 ;
  assign \g62636/_0_  = ~n7530 ;
  assign \g62637/_0_  = ~n7533 ;
  assign \g62638/_0_  = ~n7536 ;
  assign \g62639/_0_  = ~n7539 ;
  assign \g62640/_0_  = ~n7542 ;
  assign \g62641/_0_  = ~n7545 ;
  assign \g62642/_0_  = ~n7548 ;
  assign \g62643/_0_  = ~n7551 ;
  assign \g62644/_0_  = ~n7554 ;
  assign \g62645/_0_  = ~n7557 ;
  assign \g62646/_0_  = ~n7560 ;
  assign \g62647/_0_  = ~n7563 ;
  assign \g62648/_0_  = ~n7566 ;
  assign \g62649/_0_  = ~n7569 ;
  assign \g62650/_0_  = ~n7572 ;
  assign \g62651/_0_  = ~n7575 ;
  assign \g62652/_0_  = ~n7578 ;
  assign \g62653/_0_  = ~n7581 ;
  assign \g62654/_0_  = ~n7584 ;
  assign \g62655/_0_  = ~n7587 ;
  assign \g62656/_0_  = ~n7590 ;
  assign \g62657/_0_  = ~n7593 ;
  assign \g62658/_0_  = ~n7596 ;
  assign \g62659/_0_  = ~n7599 ;
  assign \g62660/_0_  = ~n7602 ;
  assign \g62661/_0_  = n7604 ;
  assign \g62674/_0_  = ~n7607 ;
  assign \g62682/_0_  = ~n7610 ;
  assign \g62683/_0_  = n7612 ;
  assign \g62689/_0_  = ~n7619 ;
  assign \g62690/_0_  = ~n7626 ;
  assign \g62691/_0_  = ~n7633 ;
  assign \g62694/_0_  = ~n7640 ;
  assign \g62695/_0_  = ~n7647 ;
  assign \g62696/_0_  = ~n7654 ;
  assign \g62698/_0_  = ~n7661 ;
  assign \g62699/_0_  = ~n7668 ;
  assign \g62700/_0_  = ~n7675 ;
  assign \g62723/_0_  = ~n7679 ;
  assign \g62724/_0_  = ~n7683 ;
  assign \g62725/_0_  = ~n7687 ;
  assign \g62726/_0_  = ~n7691 ;
  assign \g62727/_0_  = ~n7695 ;
  assign \g62728/_0_  = ~n7699 ;
  assign \g62735/_0_  = ~n7703 ;
  assign \g62736/_0_  = ~n7707 ;
  assign \g62737/_0_  = ~n7711 ;
  assign \g62738/_0_  = ~n7715 ;
  assign \g62739/_0_  = ~n7719 ;
  assign \g62740/_0_  = ~n7723 ;
  assign \g62754/_0_  = ~n7726 ;
  assign \g62762/_0_  = ~n7729 ;
  assign \g62763/_0_  = ~n7732 ;
  assign \g62764/_0_  = ~n7735 ;
  assign \g62780/_0_  = ~n7738 ;
  assign \g62781/_0_  = ~n7741 ;
  assign \g62785/_0_  = ~n7744 ;
  assign \g62786/_0_  = ~n7747 ;
  assign \g62787/_0_  = ~n7750 ;
  assign \g62791/_0_  = ~n7753 ;
  assign \g62792/_0_  = ~n7756 ;
  assign \g62794/_0_  = ~n7759 ;
  assign \g62804/_0_  = n7762 ;
  assign \g62806/_0_  = n7765 ;
  assign \g62807/_0_  = n7766 ;
  assign \g62811/_0_  = n7769 ;
  assign \g62968/_0_  = n7773 ;
  assign \g63005/_0_  = n7777 ;
  assign \g63041/_0_  = n7779 ;
  assign \g63116/_0_  = n7785 ;
  assign \g63157/_0_  = n7791 ;
  assign \g63164/_0_  = n7793 ;
  assign \g63170/_0_  = n7799 ;
  assign \g63189/_0_  = n7801 ;
  assign \g63202/_0_  = ~n7806 ;
  assign \g63206/_0_  = n7808 ;
  assign \g63207/_0_  = n7820 ;
  assign \g63265/_0_  = ~n7823 ;
  assign \g63266/_0_  = ~n7826 ;
  assign \g63269/_0_  = ~n7829 ;
  assign \g63271/_0_  = ~n7832 ;
  assign \g63272/_0_  = ~n7835 ;
  assign \g63273/_0_  = ~n7838 ;
  assign \g63274/_0_  = ~n7841 ;
  assign \g63275/_0_  = ~n7844 ;
  assign \g63276/_0_  = ~n7847 ;
  assign \g63277/_0_  = ~n7850 ;
  assign \g63278/_0_  = ~n7853 ;
  assign \g63280/_0_  = ~n7856 ;
  assign \g63281/_0_  = ~n7859 ;
  assign \g63282/_0_  = ~n7862 ;
  assign \g63283/_0_  = ~n7865 ;
  assign \g63284/_0_  = ~n7868 ;
  assign \g63285/_0_  = ~n7871 ;
  assign \g63286/_0_  = ~n7874 ;
  assign \g63287/_0_  = ~n7877 ;
  assign \g63288/_0_  = ~n7880 ;
  assign \g63289/_0_  = ~n7883 ;
  assign \g63290/_0_  = ~n7886 ;
  assign \g63292/_0_  = ~n7889 ;
  assign \g63293/_0_  = ~n7892 ;
  assign \g63294/_0_  = ~n7895 ;
  assign \g63295/_0_  = ~n7898 ;
  assign \g63296/_0_  = ~n7901 ;
  assign \g63297/_0_  = ~n7904 ;
  assign \g63298/_0_  = ~n7907 ;
  assign \g63299/_0_  = ~n7910 ;
  assign \g63302/_0_  = ~n7913 ;
  assign \g63303/_0_  = ~n7916 ;
  assign \g63304/_0_  = ~n7919 ;
  assign \g63305/_0_  = ~n7922 ;
  assign \g63306/_0_  = ~n7925 ;
  assign \g63307/_0_  = ~n7928 ;
  assign \g63308/_0_  = ~n7931 ;
  assign \g63309/_0_  = ~n7934 ;
  assign \g63310/_0_  = ~n7937 ;
  assign \g63311/_0_  = ~n7940 ;
  assign \g63312/_0_  = ~n7943 ;
  assign \g63313/_0_  = ~n7946 ;
  assign \g63314/_0_  = ~n7949 ;
  assign \g63315/_0_  = ~n7952 ;
  assign \g63316/_0_  = ~n7955 ;
  assign \g63317/_0_  = ~n7958 ;
  assign \g63318/_0_  = ~n7961 ;
  assign \g63319/_0_  = ~n7964 ;
  assign \g63320/_0_  = ~n7967 ;
  assign \g63321/_0_  = ~n7970 ;
  assign \g63322/_0_  = ~n7973 ;
  assign \g63323/_0_  = ~n7976 ;
  assign \g63324/_0_  = ~n7979 ;
  assign \g63325/_0_  = ~n7982 ;
  assign \g63326/_0_  = ~n7985 ;
  assign \g63327/_0_  = ~n7988 ;
  assign \g63328/_0_  = ~n7991 ;
  assign \g63329/_0_  = ~n7994 ;
  assign \g63330/_0_  = ~n7997 ;
  assign \g63331/_0_  = ~n8000 ;
  assign \g63339/_0_  = ~n8005 ;
  assign \g63505/_0_  = n8009 ;
  assign \g63525/_0_  = n6245 ;
  assign \g63543/_1_  = n5278 ;
  assign \g63602/_0_  = n8014 ;
  assign \g63653/_0_  = n5287 ;
  assign \g63663/_1_  = n5306 ;
  assign \g63677/_0_  = n6378 ;
  assign \g63694/_0_  = n6415 ;
  assign \g63729/_0_  = n8017 ;
  assign \g63766/_0_  = ~n8025 ;
  assign \g63771/_1_  = n5952 ;
  assign \g63773/_1_  = n5960 ;
  assign \g63784/_1_  = n5958 ;
  assign \g63964/_0_  = n8073 ;
  assign \g63965/_0_  = n8097 ;
  assign \g63966/_0_  = ~n8108 ;
  assign \g63967/_0_  = ~n8137 ;
  assign \g64257/_1_  = n2600 ;
  assign \g64266/_0_  = n8143 ;
  assign \g64275/_0_  = n8147 ;
  assign \g64400/_0_  = n5971 ;
  assign \g64416/_0_  = n6320 ;
  assign \g64470/_3_  = ~n8153 ;
  assign \g64473/_0_  = n8158 ;
  assign \g64474/_0_  = n8163 ;
  assign \g64475/_0_  = n8168 ;
  assign \g64479/_0_  = ~n8180 ;
  assign \g64480/_0_  = ~n8187 ;
  assign \g64481/_0_  = ~n8194 ;
  assign \g64483/_0_  = n8199 ;
  assign \g64484/_0_  = ~n8204 ;
  assign \g64485/_0_  = ~n8207 ;
  assign \g64486/_0_  = ~n8210 ;
  assign \g64493/_0_  = n8215 ;
  assign \g64494/_0_  = n8220 ;
  assign \g64495/_0_  = n8225 ;
  assign \g64496/_0_  = n8230 ;
  assign \g64505/_3_  = n8233 ;
  assign \g64507/_0_  = n8238 ;
  assign \g64508/_0_  = n8243 ;
  assign \g64510/_0_  = n8248 ;
  assign \g64511/_0_  = n8253 ;
  assign \g64544/_0_  = ~n8256 ;
  assign \g64545/_0_  = ~n8259 ;
  assign \g64546/_0_  = ~n8262 ;
  assign \g64639/_0_  = n8265 ;
  assign \g64641/_0_  = ~n8269 ;
  assign \g64642/_0_  = n8273 ;
  assign \g64645/_0_  = n8276 ;
  assign \g64650/_0_  = n8279 ;
  assign \g64737/_0_  = n8282 ;
  assign \g64738/_0_  = n8286 ;
  assign \g65066/_0_  = n5903 ;
  assign \g65070/_0_  = n4325 ;
  assign \g65090/_0_  = n1892 ;
  assign \g65102/_0_  = n6027 ;
  assign \g65102/_3_  = ~n6027 ;
  assign \g65126/_3_  = ~n6511 ;
  assign \g65147/_3_  = ~n6541 ;
  assign \g65163/_0_  = n5758 ;
  assign \g65176/_3_  = ~n6596 ;
  assign \g65178/_0_  = n5152 ;
  assign \g65182/_0_  = n5713 ;
  assign \g65190/_1_  = n1905 ;
  assign \g65191/_0_  = n5032 ;
  assign \g65196/_0_  = n4974 ;
  assign \g65268/_0_  = n1673 ;
  assign \g65275/_0_  = n3176 ;
  assign \g65290/_0_  = n6089 ;
  assign \g65290/_3_  = ~n6089 ;
  assign \g65291/_0_  = n3188 ;
  assign \g65292/_0_  = n4312 ;
  assign \g65298/_0_  = n6058 ;
  assign \g65298/_3_  = ~n6058 ;
  assign \g65314/_0_  = n6120 ;
  assign \g65314/_3_  = ~n6120 ;
  assign \g65319/_3_  = ~n6624 ;
  assign \g65335/_0_  = n5853 ;
  assign \g65342/_0_  = n1589 ;
  assign \g65348/_0_  = n5195 ;
  assign \g65422/_0_  = n8289 ;
  assign \g65465/_1_  = n8184 ;
  assign \g65469/_1_  = n8191 ;
  assign \g65478/_1_  = n8175 ;
  assign \g65507/_0_  = ~n5059 ;
  assign \g65548/_0_  = ~n6037 ;
  assign \g65699/_1_  = n1274 ;
  assign \g65713/_1_  = n2785 ;
  assign \g65835/_0_  = ~n8290 ;
  assign \g65860/_0_  = n8293 ;
  assign \g65863/_0_  = ~n8294 ;
  assign \g66094/_1_  = ~n6068 ;
  assign \g66102/_0_  = ~n8299 ;
  assign \g66107/_0_  = ~n8302 ;
  assign \g66130/_3_  = ~n8305 ;
  assign \g66131/_3_  = ~n8308 ;
  assign \g66228/_1_  = n7282 ;
  assign \g66348/_1_  = ~n1493 ;
  assign \g66543/_0_  = ~n8310 ;
  assign \g66549/_1_  = ~n6130 ;
  assign \g66640/_3_  = ~n8313 ;
  assign \g66641/_3_  = ~n8316 ;
  assign \g66950/_1_  = n6004 ;
  assign \g67111/_0_  = n8317 ;
  assign \g67219/_0_  = n8318 ;
  assign \g67263/_0_  = n8320 ;
  assign \g67909/_1_  = n7285 ;
  assign \g68049/_0_  = n8322 ;
  assign \g68220/_0_  = ~\g805_reg/NET0131  ;
  assign \g68413/_0_  = ~\g801_reg/NET0131  ;
  assign \g68511/_0_  = ~\g97_reg/NET0131  ;
  assign \g68536/_0_  = ~\g793_reg/NET0131  ;
  assign \g68543/_1_  = ~n1489 ;
  assign \g68554/_0_  = n8323 ;
  assign \g68559/_0_  = n8324 ;
  assign \g70915/_0_  = ~n8341 ;
  assign \g71108/_1_  = n3097 ;
  assign \g71115/_2_  = ~n8342 ;
  assign \g71244_dup/_0_  = n2928 ;
  assign \g71368/_0_  = ~n8358 ;
  assign \g71581/_0_  = ~n8365 ;
  assign \g71720/_0_  = n1219 ;
  assign \g785_reg/P0001  = ~\g785_reg/NET0131  ;
  assign \g789_reg/P0001  = ~\g789_reg/NET0131  ;
  assign \g797_reg/P0001  = ~\g797_reg/NET0131  ;
  assign \g809_reg/P0001  = ~\g809_reg/NET0131  ;
  assign \g813_reg/P0001  = ~\g813_reg/NET0131  ;
  assign \g966_reg/P0001  = ~\g966_reg/NET0131  ;
  assign \g968_reg/P0001  = ~\g968_reg/NET0131  ;
  assign \g970_reg/P0001  = ~\g970_reg/NET0131  ;
  assign \g972_reg/P0001  = ~\g972_reg/NET0131  ;
  assign \g974_reg/P0001  = ~\g974_reg/NET0131  ;
  assign \g976_reg/P0001  = ~\g976_reg/NET0131  ;
  assign \g978_reg/P0001  = ~\g978_reg/NET0131  ;
endmodule
