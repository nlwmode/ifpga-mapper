module top( a_pad , b_pad , c_pad , d_pad , e_pad , f_pad , g_pad , h_pad , i_pad , j_pad , k_pad , m_pad , n_pad , o_pad , p_pad , q_pad , \u247_syn_3  );
  input a_pad ;
  input b_pad ;
  input c_pad ;
  input d_pad ;
  input e_pad ;
  input f_pad ;
  input g_pad ;
  input h_pad ;
  input i_pad ;
  input j_pad ;
  output k_pad ;
  output m_pad ;
  output n_pad ;
  output o_pad ;
  output p_pad ;
  output q_pad ;
  output \u247_syn_3  ;
  wire n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 ;
  assign n11 = h_pad & i_pad ;
  assign n12 = ~j_pad & n11 ;
  assign n13 = ~i_pad & ~j_pad ;
  assign n14 = ~h_pad & n13 ;
  assign n16 = ~a_pad & ~b_pad ;
  assign n17 = ~c_pad & n16 ;
  assign n15 = ~h_pad & i_pad ;
  assign n18 = ~j_pad & n15 ;
  assign n19 = n17 & n18 ;
  assign n20 = i_pad & j_pad ;
  assign n21 = g_pad & h_pad ;
  assign n22 = ~n20 & n21 ;
  assign n23 = c_pad & n16 ;
  assign n29 = ~i_pad & n23 ;
  assign n30 = f_pad & n20 ;
  assign n31 = ~n29 & ~n30 ;
  assign n32 = ~h_pad & ~n31 ;
  assign n24 = n20 & n23 ;
  assign n25 = d_pad & ~e_pad ;
  assign n26 = ~j_pad & n25 ;
  assign n27 = ~n24 & ~n26 ;
  assign n28 = h_pad & ~n27 ;
  assign n33 = g_pad & ~n13 ;
  assign n34 = ~n28 & n33 ;
  assign n35 = ~n32 & n34 ;
  assign n36 = i_pad & ~n17 ;
  assign n37 = h_pad & ~n36 ;
  assign n38 = f_pad & n15 ;
  assign n39 = ~n37 & ~n38 ;
  assign n40 = j_pad & ~n39 ;
  assign n42 = d_pad & e_pad ;
  assign n43 = h_pad & ~n42 ;
  assign n41 = h_pad & ~i_pad ;
  assign n44 = ~j_pad & ~n15 ;
  assign n45 = ~n41 & n44 ;
  assign n46 = ~n43 & n45 ;
  assign n47 = g_pad & ~n46 ;
  assign n48 = ~n40 & n47 ;
  assign n49 = j_pad & n41 ;
  assign n50 = ~n14 & ~n49 ;
  assign k_pad = ~n12 ;
  assign m_pad = n14 ;
  assign n_pad = ~n19 ;
  assign o_pad = ~n22 ;
  assign p_pad = ~n35 ;
  assign q_pad = ~n48 ;
  assign \u247_syn_3  = n50 ;
endmodule
