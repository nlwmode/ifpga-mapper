module top (\G10_pad , \G11_pad , \G12_pad , \G13_pad , \G14_pad , \G15_pad , \G16_pad , \G18_pad , \G19_pad , \G20_pad , \G22_pad , \G23_pad , \G24_pad , \G25_pad , \G26_pad , \G28_pad , \G2_pad , \G30_pad , \G31_pad , \G32_pad , \G33_pad , \G34_pad , \G35_pad , \G3_pad , \G4_pad , \G5_pad , \G64_reg/NET0131 , \G65_reg/NET0131 , \G66_reg/NET0131 , \G69_reg/NET0131 , \G6_pad , \G70_reg/NET0131 , \G71_reg/NET0131 , \G72_reg/NET0131 , \G73_reg/NET0131 , \G74_reg/NET0131 , \G75_reg/NET0131 , \G76_reg/NET0131 , \G77_reg/NET0131 , \G79_reg/NET0131 , \G81_reg/NET0131 , \G8_pad , \G9_pad , \G100BF_pad , \G103BF_pad , \G104BF_pad , \G105BF_pad , \G107_pad , \G83_pad , \G84_pad , \G86BF_pad , \G87BF_pad , \G88BF_pad , \G89BF_pad , \G90_pad , \G95BF_pad , \G96BF_pad , \G97BF_pad , \G98BF_pad , \G99BF_pad , \_al_n0 , \_al_n1 , \g1049/_0_ , \g1081/_0_ , \g1115/_0_ , \g13/_1_ , \g809/_0_ , \g810/_0_ , \g814/_0_ , \g825/_2_ , \g834/_0_ , \g863/_0_ , \g870/_0_ , \g871/_0_ , \g916/_0_ , \g917/_0_ , \g940/_3_ );
	input \G10_pad  ;
	input \G11_pad  ;
	input \G12_pad  ;
	input \G13_pad  ;
	input \G14_pad  ;
	input \G15_pad  ;
	input \G16_pad  ;
	input \G18_pad  ;
	input \G19_pad  ;
	input \G20_pad  ;
	input \G22_pad  ;
	input \G23_pad  ;
	input \G24_pad  ;
	input \G25_pad  ;
	input \G26_pad  ;
	input \G28_pad  ;
	input \G2_pad  ;
	input \G30_pad  ;
	input \G31_pad  ;
	input \G32_pad  ;
	input \G33_pad  ;
	input \G34_pad  ;
	input \G35_pad  ;
	input \G3_pad  ;
	input \G4_pad  ;
	input \G5_pad  ;
	input \G64_reg/NET0131  ;
	input \G65_reg/NET0131  ;
	input \G66_reg/NET0131  ;
	input \G69_reg/NET0131  ;
	input \G6_pad  ;
	input \G70_reg/NET0131  ;
	input \G71_reg/NET0131  ;
	input \G72_reg/NET0131  ;
	input \G73_reg/NET0131  ;
	input \G74_reg/NET0131  ;
	input \G75_reg/NET0131  ;
	input \G76_reg/NET0131  ;
	input \G77_reg/NET0131  ;
	input \G79_reg/NET0131  ;
	input \G81_reg/NET0131  ;
	input \G8_pad  ;
	input \G9_pad  ;
	output \G100BF_pad  ;
	output \G103BF_pad  ;
	output \G104BF_pad  ;
	output \G105BF_pad  ;
	output \G107_pad  ;
	output \G83_pad  ;
	output \G84_pad  ;
	output \G86BF_pad  ;
	output \G87BF_pad  ;
	output \G88BF_pad  ;
	output \G89BF_pad  ;
	output \G90_pad  ;
	output \G95BF_pad  ;
	output \G96BF_pad  ;
	output \G97BF_pad  ;
	output \G98BF_pad  ;
	output \G99BF_pad  ;
	output \_al_n0  ;
	output \_al_n1  ;
	output \g1049/_0_  ;
	output \g1081/_0_  ;
	output \g1115/_0_  ;
	output \g13/_1_  ;
	output \g809/_0_  ;
	output \g810/_0_  ;
	output \g814/_0_  ;
	output \g825/_2_  ;
	output \g834/_0_  ;
	output \g863/_0_  ;
	output \g870/_0_  ;
	output \g871/_0_  ;
	output \g916/_0_  ;
	output \g917/_0_  ;
	output \g940/_3_  ;
	wire _w121_ ;
	wire _w120_ ;
	wire _w119_ ;
	wire _w118_ ;
	wire _w117_ ;
	wire _w116_ ;
	wire _w115_ ;
	wire _w114_ ;
	wire _w113_ ;
	wire _w112_ ;
	wire _w111_ ;
	wire _w110_ ;
	wire _w109_ ;
	wire _w108_ ;
	wire _w107_ ;
	wire _w106_ ;
	wire _w105_ ;
	wire _w104_ ;
	wire _w73_ ;
	wire _w72_ ;
	wire _w71_ ;
	wire _w70_ ;
	wire _w69_ ;
	wire _w68_ ;
	wire _w67_ ;
	wire _w66_ ;
	wire _w65_ ;
	wire _w64_ ;
	wire _w63_ ;
	wire _w62_ ;
	wire _w61_ ;
	wire _w60_ ;
	wire _w59_ ;
	wire _w58_ ;
	wire _w45_ ;
	wire _w46_ ;
	wire _w47_ ;
	wire _w48_ ;
	wire _w49_ ;
	wire _w50_ ;
	wire _w51_ ;
	wire _w52_ ;
	wire _w53_ ;
	wire _w54_ ;
	wire _w55_ ;
	wire _w56_ ;
	wire _w57_ ;
	wire _w74_ ;
	wire _w75_ ;
	wire _w76_ ;
	wire _w77_ ;
	wire _w78_ ;
	wire _w79_ ;
	wire _w80_ ;
	wire _w81_ ;
	wire _w82_ ;
	wire _w83_ ;
	wire _w84_ ;
	wire _w85_ ;
	wire _w86_ ;
	wire _w87_ ;
	wire _w88_ ;
	wire _w89_ ;
	wire _w90_ ;
	wire _w91_ ;
	wire _w92_ ;
	wire _w93_ ;
	wire _w94_ ;
	wire _w95_ ;
	wire _w96_ ;
	wire _w97_ ;
	wire _w98_ ;
	wire _w99_ ;
	wire _w100_ ;
	wire _w101_ ;
	wire _w102_ ;
	wire _w103_ ;
	LUT2 #(
		.INIT('h4)
	) name0 (
		\G4_pad ,
		\G69_reg/NET0131 ,
		_w45_
	);
	LUT3 #(
		.INIT('hdf)
	) name1 (
		\G35_pad ,
		\G4_pad ,
		\G69_reg/NET0131 ,
		_w46_
	);
	LUT2 #(
		.INIT('h1)
	) name2 (
		\G10_pad ,
		\G13_pad ,
		_w47_
	);
	LUT4 #(
		.INIT('h0100)
	) name3 (
		\G10_pad ,
		\G13_pad ,
		\G3_pad ,
		\G9_pad ,
		_w48_
	);
	LUT2 #(
		.INIT('h1)
	) name4 (
		\G11_pad ,
		\G3_pad ,
		_w49_
	);
	LUT3 #(
		.INIT('h8a)
	) name5 (
		\G24_pad ,
		\G2_pad ,
		\G66_reg/NET0131 ,
		_w50_
	);
	LUT3 #(
		.INIT('hef)
	) name6 (
		_w48_,
		_w49_,
		_w50_,
		_w51_
	);
	LUT4 #(
		.INIT('h3133)
	) name7 (
		\G11_pad ,
		\G3_pad ,
		_w48_,
		_w50_,
		_w52_
	);
	LUT2 #(
		.INIT('h2)
	) name8 (
		\G77_reg/NET0131 ,
		_w52_,
		_w53_
	);
	LUT4 #(
		.INIT('h0002)
	) name9 (
		\G10_pad ,
		\G13_pad ,
		\G3_pad ,
		\G9_pad ,
		_w54_
	);
	LUT4 #(
		.INIT('h00c8)
	) name10 (
		\G11_pad ,
		\G23_pad ,
		\G3_pad ,
		\G65_reg/NET0131 ,
		_w55_
	);
	LUT2 #(
		.INIT('hb)
	) name11 (
		_w54_,
		_w55_,
		_w56_
	);
	LUT4 #(
		.INIT('h8c88)
	) name12 (
		\G3_pad ,
		\G76_reg/NET0131 ,
		_w54_,
		_w55_,
		_w57_
	);
	LUT2 #(
		.INIT('h4)
	) name13 (
		\G2_pad ,
		\G64_reg/NET0131 ,
		_w58_
	);
	LUT4 #(
		.INIT('h0d00)
	) name14 (
		\G77_reg/NET0131 ,
		_w52_,
		_w57_,
		_w58_,
		_w59_
	);
	LUT3 #(
		.INIT('h01)
	) name15 (
		\G10_pad ,
		\G13_pad ,
		\G9_pad ,
		_w60_
	);
	LUT4 #(
		.INIT('hccc8)
	) name16 (
		\G10_pad ,
		\G11_pad ,
		\G13_pad ,
		\G9_pad ,
		_w61_
	);
	LUT3 #(
		.INIT('ha8)
	) name17 (
		\G22_pad ,
		\G3_pad ,
		_w61_,
		_w62_
	);
	LUT2 #(
		.INIT('hb)
	) name18 (
		_w59_,
		_w62_,
		_w63_
	);
	LUT4 #(
		.INIT('h8c88)
	) name19 (
		\G3_pad ,
		\G75_reg/NET0131 ,
		_w59_,
		_w62_,
		_w64_
	);
	LUT2 #(
		.INIT('h7)
	) name20 (
		\G14_pad ,
		_w64_,
		_w65_
	);
	LUT2 #(
		.INIT('h7)
	) name21 (
		\G15_pad ,
		_w57_,
		_w66_
	);
	LUT3 #(
		.INIT('hf7)
	) name22 (
		\G16_pad ,
		\G77_reg/NET0131 ,
		_w52_,
		_w67_
	);
	LUT3 #(
		.INIT('h20)
	) name23 (
		\G18_pad ,
		\G4_pad ,
		\G79_reg/NET0131 ,
		_w68_
	);
	LUT3 #(
		.INIT('h20)
	) name24 (
		\G19_pad ,
		\G4_pad ,
		\G65_reg/NET0131 ,
		_w69_
	);
	LUT3 #(
		.INIT('h20)
	) name25 (
		\G20_pad ,
		\G4_pad ,
		\G81_reg/NET0131 ,
		_w70_
	);
	LUT4 #(
		.INIT('h0200)
	) name26 (
		\G10_pad ,
		\G13_pad ,
		\G3_pad ,
		\G9_pad ,
		_w71_
	);
	LUT3 #(
		.INIT('hc8)
	) name27 (
		\G11_pad ,
		\G25_pad ,
		\G3_pad ,
		_w72_
	);
	LUT2 #(
		.INIT('hb)
	) name28 (
		_w71_,
		_w72_,
		_w73_
	);
	LUT2 #(
		.INIT('h4)
	) name29 (
		\G4_pad ,
		\G73_reg/NET0131 ,
		_w74_
	);
	LUT2 #(
		.INIT('h8)
	) name30 (
		_w60_,
		_w74_,
		_w75_
	);
	LUT4 #(
		.INIT('h2000)
	) name31 (
		\G74_reg/NET0131 ,
		_w59_,
		_w62_,
		_w75_,
		_w76_
	);
	LUT4 #(
		.INIT('h0200)
	) name32 (
		\G70_reg/NET0131 ,
		_w48_,
		_w49_,
		_w50_,
		_w77_
	);
	LUT3 #(
		.INIT('h40)
	) name33 (
		\G4_pad ,
		\G69_reg/NET0131 ,
		\G9_pad ,
		_w78_
	);
	LUT2 #(
		.INIT('h8)
	) name34 (
		_w47_,
		_w78_,
		_w79_
	);
	LUT2 #(
		.INIT('h8)
	) name35 (
		_w77_,
		_w79_,
		_w80_
	);
	LUT3 #(
		.INIT('h20)
	) name36 (
		\G72_reg/NET0131 ,
		_w54_,
		_w55_,
		_w81_
	);
	LUT2 #(
		.INIT('h4)
	) name37 (
		\G4_pad ,
		\G71_reg/NET0131 ,
		_w82_
	);
	LUT3 #(
		.INIT('h02)
	) name38 (
		\G10_pad ,
		\G13_pad ,
		\G9_pad ,
		_w83_
	);
	LUT2 #(
		.INIT('h8)
	) name39 (
		_w82_,
		_w83_,
		_w84_
	);
	LUT2 #(
		.INIT('h8)
	) name40 (
		\G12_pad ,
		\G26_pad ,
		_w85_
	);
	LUT3 #(
		.INIT('h70)
	) name41 (
		_w81_,
		_w84_,
		_w85_,
		_w86_
	);
	LUT2 #(
		.INIT('h4)
	) name42 (
		_w80_,
		_w86_,
		_w87_
	);
	LUT2 #(
		.INIT('h4)
	) name43 (
		_w76_,
		_w87_,
		_w88_
	);
	LUT4 #(
		.INIT('hf7ff)
	) name44 (
		\G30_pad ,
		\G74_reg/NET0131 ,
		_w59_,
		_w62_,
		_w89_
	);
	LUT3 #(
		.INIT('hdf)
	) name45 (
		\G31_pad ,
		\G4_pad ,
		\G73_reg/NET0131 ,
		_w90_
	);
	LUT4 #(
		.INIT('hf7ff)
	) name46 (
		\G32_pad ,
		\G72_reg/NET0131 ,
		_w54_,
		_w55_,
		_w91_
	);
	LUT3 #(
		.INIT('hdf)
	) name47 (
		\G33_pad ,
		\G4_pad ,
		\G71_reg/NET0131 ,
		_w92_
	);
	LUT2 #(
		.INIT('h7)
	) name48 (
		\G34_pad ,
		_w77_,
		_w93_
	);
	LUT4 #(
		.INIT('h5100)
	) name49 (
		\G2_pad ,
		\G77_reg/NET0131 ,
		_w52_,
		_w57_,
		_w94_
	);
	LUT4 #(
		.INIT('hef20)
	) name50 (
		\G74_reg/NET0131 ,
		_w59_,
		_w62_,
		_w74_,
		_w95_
	);
	LUT2 #(
		.INIT('h2)
	) name51 (
		\G2_pad ,
		\G5_pad ,
		_w96_
	);
	LUT2 #(
		.INIT('h2)
	) name52 (
		_w57_,
		_w96_,
		_w97_
	);
	LUT3 #(
		.INIT('h40)
	) name53 (
		\G4_pad ,
		\G5_pad ,
		\G71_reg/NET0131 ,
		_w98_
	);
	LUT4 #(
		.INIT('h2000)
	) name54 (
		\G72_reg/NET0131 ,
		_w54_,
		_w55_,
		_w98_,
		_w99_
	);
	LUT3 #(
		.INIT('hd0)
	) name55 (
		\G77_reg/NET0131 ,
		_w52_,
		_w99_,
		_w100_
	);
	LUT3 #(
		.INIT('hdc)
	) name56 (
		_w64_,
		_w97_,
		_w100_,
		_w101_
	);
	LUT2 #(
		.INIT('h2)
	) name57 (
		\G2_pad ,
		\G6_pad ,
		_w102_
	);
	LUT3 #(
		.INIT('h02)
	) name58 (
		\G77_reg/NET0131 ,
		_w52_,
		_w102_,
		_w103_
	);
	LUT3 #(
		.INIT('h40)
	) name59 (
		\G4_pad ,
		\G69_reg/NET0131 ,
		\G6_pad ,
		_w104_
	);
	LUT3 #(
		.INIT('h40)
	) name60 (
		_w57_,
		_w77_,
		_w104_,
		_w105_
	);
	LUT3 #(
		.INIT('hdc)
	) name61 (
		_w64_,
		_w103_,
		_w105_,
		_w106_
	);
	LUT2 #(
		.INIT('h2)
	) name62 (
		\G2_pad ,
		\G8_pad ,
		_w107_
	);
	LUT3 #(
		.INIT('h40)
	) name63 (
		\G4_pad ,
		\G73_reg/NET0131 ,
		\G8_pad ,
		_w108_
	);
	LUT4 #(
		.INIT('h0d00)
	) name64 (
		\G77_reg/NET0131 ,
		_w52_,
		_w57_,
		_w108_,
		_w109_
	);
	LUT4 #(
		.INIT('h2000)
	) name65 (
		\G74_reg/NET0131 ,
		_w59_,
		_w62_,
		_w109_,
		_w110_
	);
	LUT3 #(
		.INIT('hf2)
	) name66 (
		_w64_,
		_w107_,
		_w110_,
		_w111_
	);
	LUT4 #(
		.INIT('h0051)
	) name67 (
		\G2_pad ,
		\G77_reg/NET0131 ,
		_w52_,
		_w57_,
		_w112_
	);
	LUT2 #(
		.INIT('h8)
	) name68 (
		_w64_,
		_w112_,
		_w113_
	);
	LUT4 #(
		.INIT('h20ff)
	) name69 (
		\G74_reg/NET0131 ,
		_w59_,
		_w62_,
		_w74_,
		_w114_
	);
	LUT3 #(
		.INIT('h04)
	) name70 (
		\G2_pad ,
		\G77_reg/NET0131 ,
		_w52_,
		_w115_
	);
	LUT4 #(
		.INIT('ha8aa)
	) name71 (
		_w45_,
		_w48_,
		_w49_,
		_w50_,
		_w116_
	);
	LUT2 #(
		.INIT('he)
	) name72 (
		_w77_,
		_w116_,
		_w117_
	);
	LUT2 #(
		.INIT('hd)
	) name73 (
		_w45_,
		_w77_,
		_w118_
	);
	LUT4 #(
		.INIT('h20ff)
	) name74 (
		\G72_reg/NET0131 ,
		_w54_,
		_w55_,
		_w82_,
		_w119_
	);
	LUT4 #(
		.INIT('hef20)
	) name75 (
		\G72_reg/NET0131 ,
		_w54_,
		_w55_,
		_w82_,
		_w120_
	);
	LUT4 #(
		.INIT('h8000)
	) name76 (
		\G11_pad ,
		\G12_pad ,
		\G13_pad ,
		\G28_pad ,
		_w121_
	);
	assign \G100BF_pad  = _w46_ ;
	assign \G103BF_pad  = _w65_ ;
	assign \G104BF_pad  = _w66_ ;
	assign \G105BF_pad  = _w67_ ;
	assign \G107_pad  = _w68_ ;
	assign \G83_pad  = _w69_ ;
	assign \G84_pad  = _w70_ ;
	assign \G86BF_pad  = _w63_ ;
	assign \G87BF_pad  = _w56_ ;
	assign \G88BF_pad  = _w51_ ;
	assign \G89BF_pad  = _w73_ ;
	assign \G90_pad  = _w88_ ;
	assign \G95BF_pad  = _w89_ ;
	assign \G96BF_pad  = _w90_ ;
	assign \G97BF_pad  = _w91_ ;
	assign \G98BF_pad  = _w92_ ;
	assign \G99BF_pad  = _w93_ ;
	assign \_al_n0  = 1'b0;
	assign \_al_n1  = 1'b1;
	assign \g1049/_0_  = _w94_ ;
	assign \g1081/_0_  = _w64_ ;
	assign \g1115/_0_  = _w95_ ;
	assign \g13/_1_  = _w53_ ;
	assign \g809/_0_  = _w101_ ;
	assign \g810/_0_  = _w106_ ;
	assign \g814/_0_  = _w111_ ;
	assign \g825/_2_  = _w113_ ;
	assign \g834/_0_  = _w114_ ;
	assign \g863/_0_  = _w115_ ;
	assign \g870/_0_  = _w117_ ;
	assign \g871/_0_  = _w118_ ;
	assign \g916/_0_  = _w119_ ;
	assign \g917/_0_  = _w120_ ;
	assign \g940/_3_  = _w121_ ;
endmodule;